// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CtZF8PV4MMAmfaOBtXmyVSJt7kD0oANehf4VlUpMqsLkv9FePciGttZV7giD
z0F4CrNcDCx/3a/5a7/BIvcPRkBxr1Ij1WyKEchYtufZsUl63zSZQnUoNtLf
pL9P4N2rnPDCPy+w4fZ//5XpdXTzV2YunWkuqg4+4+j8SHlEzQcrCqd5ZHB8
bmZCzMFUfmd4fJN3mJ99clmcjKtU7I5zfekli0tnMjtK97BZUHaCW8vM1TAR
Drn4g/qX9b0MTJ0MpDQdbtxC5ubY8vhlCX0m3uOTDGRj1mK10servvnpAfIn
9smBs27lG1GdFgPj5G6GPPVo1aVy0wRSmGSHqDaG+Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Y7j/gf+hRTkZ1S2QQFTUloxiuXa/SVBPvhaiRPo8lPFTikyJypyE2mjzTAxB
DehxYYX27Pzoi0wXUWS2MlHWS2a165Zi3SRkIXlaytnbi0FWCG6GOoy6Mpds
QFsH4luHCNN7ARdfCcGBScZP7U24gaxSlRvbkyAhQV9wrOJbKj3soBLZEp+S
MY9qe0A3JZxOu7Mz1YsELQ828XNjfgZQ8tqgv0xror6OzSC80O/+nzun8KKT
KAl0NRni+lwqqdXy1XAln9/tX/ABvbqhdBmzTEl9nUvrHVeKfl887kT7lDpu
5hD4gKwniCH74igWN0Aad7+zMRGMK0I/zyo4rC6bLQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PoGtYh3oyIhGaIe8/LdpC5r8cC6XUm23KicCrDu15+Bon75YC2Cu1tQa+jE5
78oJ0LuoD2VF8WannCuxE+sJ8m1zNZKp5YCzrmbaBaIScp9z/N/OtK+PyzuX
1IJ0lrEN+MG/c/94/oV+htHZF1j2BFJugWH6ibWFlmtdPmfquGyt+WbpF/ux
/MdFl9E/KoqchXkA08uECT22HppJISEQXDnOlDuyh46Pe1/VPQ8bopGRUNW3
k8gkC1Mr4+JveE1Z1CnG7X4YSdsIzqjOzgZ7L8b8kcbtSygJCDChCYZZDo3B
03jrvqHVqVUYSLBWpshIp2REKCglMLXatfICia8CQQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BWN9EQSSk8cnBDhoT3WgCMRR1Vjbpqmn7/OmjpIuUIYc6iqHsgPhS7nfvk9b
eVl/+4wxnhvmMbRufodw+lDsYk+K4X0Ckp+G1om9GmuZGkPOjmDVJXdTY/34
xstzx34P8a9FfN03v2etv4D3pFPkgYbVov/5RAIMxOAPDDrtjyYzlc2VTICh
MRke6SJT4JWc2goJv/kx2qJBoP/4bkbRMxYUxsb/vT/gwy2asxAQ1ClFCJJ9
lB91EiNHBxndLvnZRDj124JI+uXzHTMck1qRgLcs0cFNXmI15Rpkquv9EPlR
dEGqICbSqDlB7LA6nGMyx4kqKGRTmW3pZ2Rs5u2WIA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Pz6W5VinuqCNyx99hq3fXlX7CIuOwHjuBpHpeXAkKfyGiKyN6X5HSmI8/9/p
uyv+jBc1jwH5fdzgWoDTMMexMmOAEzEP1rP37hjpWwbvbXeMzjIOz3U5Dcgf
uGlvsLexgC2XVO7k97eRhOgUgrIt3TWGvmPdkNXCuxmlll2tNTo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
FVcoTbx7m7KoMJcQfDhDuNSGBqFf8RtQ9vl671rO7ZBG0WasoAdvqlt/r6Gf
BxC6fmVASyOB1AyffPnGC6qotWC+pM0adW9Dw3L29T62OHPXz2jjKMPK173Y
SWDAdbhIO+mTmFmwANPrO8gVpvIADkE2RGEZv67nRkZcglAO9lDX5v2twwMM
FOhdsWF4XIBvlgiRHbQKcNxFqXDqMrBHJthnke6jOVXifI/+Wncj0NVs0K/f
a1s1Tb0D4A6TZmD98tVP6cNphrHxGHFrs009r7LnLSSEBTPAdGHd7mgtLDXY
1GxaDWqh3iawCMkO99EP14lxeLGqRg48IGS1VN1JyLdKrIxf3Yc9Bmz5bUbx
kmyRa3VRhiMtSI8T9JDkN2XasZpyO4S0teaM+lfS5jYP47Zb+4nbp74d6/Tw
s/R7lNbfjbUC2j6+4eAPIpV5DrxD08Sg4t4xNfpzKFItlDG1HfUTsb0r7q0w
udMkvlcaDxQ0kqfXWgkYdKxW6C81j97D


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sxWeFGen3ThEUQQLAgZuPklEoNMvA+inUZTxgPzRt+uckD5KP3q4q6KNrEew
05NSrrP882cVZWxZ8//uLAG54JxDgzN+NdI6vAccSacxMtLNctSiRr3nuShE
67b32PTZy+kqY8ydRzyk5BEdd1DQ6Ez8Xl64wRdqjnVrZ1pHYGY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QLiXBV/qxgCKuyd4cSXkCCIP15ZpLp6f6DvriZZQpfwFO5d/pWZIq67YIhK3
jlrWhii67qWbT5HenAz6FqYGB+tyIB9/TsNUh+H/C9X8/vadTpjzvoN2sS1R
kDQG2hA63u8G6KNJcY5RaTa2UqomaAcxGtshov1w0UgxYTMEnqs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1012928)
`pragma protect data_block
lGcvGSjyduVooRbNq3+HQ60idfKjN/YhB78H9ykgZNrkb4KDfelkPlPj59mm
5lVmH+kuhqznWbzA89aFKOZaEZv3jMWbXDG4XvKLTAFo+pJh0tLVrFar3USa
rw7AcHQIDGl+njcpGdCVnFovBlVx/1/fdi/OlR7WczuPK/bMPJjttrKOk2av
OkAiUp3nAsEK+hDtRsugjAwICt6YNGTCCzsLHJtnknbT9h9TVFw7MRGnNGDO
R+t06aPokZ0UzVyzPdPyHGEUtHnvMk+9NtnWGyrvH0AAmdty1kcRRxHvw9GJ
jn4l+phEMXcXQ28ejdzWTPhFnbL5JSjYO04PVdGj6iNGmcRGeMOBAbCGq9jB
q5K0qVWDfWTKmV5pO/ShS4AZquoM9v+XMcof13zf2fRtZbqDnaTd2dkCMhb2
wNgqxfO1nxYzxffx00sWmRXcmqICDsdJ7OpcvVRb1iQ7fXRpED8J2C2YLZ1q
kHxlW9VoJ/s3u3YrRYX3puLfZ5jReaFrrWGOz9qxGUESjLY7oHuYsrTpSRju
nKVas26QCCG/esOOf7H/TbvAkgu/sPQziuZT8x7JTk8dhSH+BLKaSoDMMaxE
SQR6BvlgjQqgwokw2k0qKloLdi9mCVjfg/cVUyEanpy4Fj6D4gqr6FeV7VUG
m1pP8OWwmBvINpe7AFGhPtsNA3MLRmKPmyWnb/5Ryx5U5aNFw+6uVeVUyUAv
Al8+CrHooGpkRhzjkbh7jH6mZHHfMQVCFQTds/SZqNs8sHIPvDTHG8EPB3pr
PtZ/9gjKeItemH7XEI9mxSnVUvu6hmIeqmokS3YubrKD3ycyOMMxhrdXx9dg
gYnZgNeGscwHlf8tepu/0BYML77MS5zXbqNhdL5BcvC0AUTXllnWQQS6ahrW
NdZB1PX83GLfjfs9LrSkuXiy+4rxJmuoBuajBiR+RtFXWHIeDlFQD0Fb0S9D
9GydVtCBO7PicVkAHV6zZV9Kf6DigwYE5L19OsGKF48mf8xoV1mWY55RbvJX
IJ0RAiui/FY5shPsd2ZRmR+YRiwvLS3/GZEAouf/hKRTzv2wxOZtZd7c+BzI
k7N3Ts2Q7tAsr1FfiNmQ3/mOpJ0c0OexXAyya5+oIhFuqArSOGSZS5lxLDrK
l+kkQ4yoKW7dxCS2+pkE4FsR5dyy2AwpELJM15ja8Bns6pS2Br39T8Euzo6C
FE5VsbCXHPHaefdvSV874TtF6Zy8wqTh30kmGk12UgXvtZmT0VjBSfU8ycNb
Ax1h0iV9Hj0eDGvUkOP0SS22je44a6FTBzdpsV9QEuF4geYcNiPzOZDFtnlH
tljZV1SN0+mrpUY5JxBfsH2YW6A/TZZ8r/mor6hNE3lXld+YlLObJ39C2Kdr
NUvPMcJ6QhStn0qE43/QF0peeqRdup0YSj9Ykciu/chwk1Zt4fTw8WPiTSM/
lPqPJPcuQ7AnP2WjWMFL/1Jt9NP9ss3Ksm38GxdW/3eW5SDLlYHJyktvUnJC
qGcF02nuKNfphPJh4s1yZdZ+tQgKMRem1Ja2cYETUyxZYWZRmhAsoyDFEFCd
FKo1rrYugOEn4pK0N2pioCdft5G60RoZXISR3XtMk8gBu4Af4fIjiMSO8LA3
vMpX2TOWBKMU9w8rJXT+8512KGQwhPYA4Yk6qeQlAmOoOiCGpoaC3bQzhQJV
62cBhV39oxFiVK7+fuxYv3wQ41gA17pfF0ZqcMOJW9VJ4wlHEBV2QR/aZ2Fu
gxzPzldBWnPz3ipV4xuF7ntEG/7j6dpk1P6O8U2KNR/T4CpqONNT7gxyK8bs
IR0Pw7JOqShpOIaV3S6zyhqb4PKrLZNdGV5KWxMPi50CvrXmeC58QYC9C+ra
uafxaZI08frzFaGhKX+JNMQRqMNINn/VFzi0mtsDOHVVgmAyccwom51ckgJn
DPrJOc7QhgEIcOSAYzn+nHgVdNVbQ0RlSS8sOXJAvGDAUeiRIh2jIEkF03SU
ov8LzcoTcNpegLM5tC3aeYM6vvFG0pU1YQ5THAr3NwnH+zsl/EHXwrO/xA9C
GrNDajv+3ZucEWCEAKlkDffs0tx+k1pKT+4zwIVUk5ixD1ToRsSSFL8x66KE
BnJ1vrrbHdZXQkPhvqS845JmXIFKBM/lkYjmYbvJED1i6TE4l9Mct82lQE/O
iXRHdGzyk+I1/q18vI6suaWs/zeilNPOUZao+gMPYpR5prnJuD6BgSy467OW
9Vcy0ndNBlLFWPnO9Lwdbz3TeptTibKCbDIs4IRVGFR578wp2Cgs0K97svRW
0OhITyI+LS+dPta97yRgVVxqiYhqRDFpmZD+UrOO2oA5UDWBMaKbdUKLiX91
GzFcF5oii0widlBacYOWOOCutE+tjbS0rMj26CADrsK0KzeNHZR5fhTG+3hj
3Cbpt3VnwEXcyAFsOeZgUDmMuljit9SlGEW97DXuGb6udkaTrNkMuyRhYHzz
PYd46ClFCdANrD0pvML6g7DMjk/C1cFJFPk+O/yMn2HgCmhwDeUl1DrMhgdh
2pamS9J+p//SuYsoVRwk6hKsQcUZh1rQqZI2eSkmxgXoqT1kXc4OsDflQPqq
KqY7RdFHmCx6VHXC90AKqnFbZc1H3dM94ANGCvdWBQ7KclqgEWVdQEKcc9HY
5PMVTb5/k19olWT4aHVeeAvHn4Vmeatn2Okymuma+qBOaM41vEGVawjZEPCl
quwsuO6NNdmARBGC/RueTCk4JUh0UGXOp24Ir9MQziPE3SWeIJc1ac7v3ldc
qP6jv/CMrCVIWM/Q92BTuhWbA4+uU8Zq8G1mfHVrUe0Z+puubJYU+oemnh+R
c6iy4skNsXWTmI0Cjte1d5EvFN305edaS0Ix+ctJW7AMKyTU/VC0CRnEMM/K
fHPaEJEJsFfUW456GkpWRKEQC8QDch/eaN3QiBTCRGgJnT5mAf+hOBmR0rCZ
wUNzLcMOwIEhawHVNLKaWmxqF8U/brkzKbGYwD1xO9etEvGYq61fSwD3usSx
ZmzzrlKT2gspZUdKVm5ObgtdqXBNNPCco/jZGza7ITkxX7dN6K+DRV7Qvnfk
tlFOiaywXXqtuNODP3qKD0FyrFHeTOjxVpVTPMzz58hyLbhIM/EV7vw1+deX
OJTU/pFD9KxLXmMk8WQ1PM8cYGQeNX3H5hnMtu6E4SvG37A69QzUpdcGFhjP
o4ChAJyAQfYRt0ng7UR0MkqSRDThgfRKCA+k/pBLiHWKk6bGvoGdtNiK/aof
QO88+qbaEISfOdwgOpjwCqE/VK3W6nd1jfzjQkGU2jyLO8iW23McruIXQHTB
bY/hSUO4NHzKy5sNvzFJGbRTc+suurCPATHbJWus+2nH+k8nzzV5WklU0Fto
rPcBOzmdLPBIgce+skGQUGKj1QlqmJ+w2o8liFBeV8r1hDG2ShcjQdB1XBUm
fBFrQp4sL5Y0pL2dttXfkGMD2j9oxVfIS7nNWjgwX+AeuVTRljNN4kXpHkEu
ygE+Y91c+c1hz32d7mmqT3JUpiRDThJmMBdKLiqNkS9QYzuHbVssJq7DXvPN
UlTYnT1pP6mm8nxKS1mvOv31SL6jpyg02tKrAR+aMmhTXPRPbpzFx7BoVOrE
x3BzYe51tb9f/w8sak56RJFMou98ZFhSsYmCAhSsaBHPggMzLI+tW5hdrfqF
clNF4yb0YmsIIkVcmYZtYUYssP+rGpXDNmBm4ZoxAVK/ucT0g7pFA0qcd8DS
e/r3mEWehp84jRxQ9+4gFfHcMKIsEhr/29467QvlAu0gol7/xeVrWWMeEJOa
EZmTWs9g4NiPhOYhncEqsZO5G+LrdP2T8msw+W338SVQM4eiCmtSm58+Ewq/
8xiBzfCSRq3QHT+PYU+2bCxd+AQzZiUAlvbGBpQiZYQhQ+QKwNq0ZtIBcLEF
/5Hk/V6g3mFsLXBSRZVP5iD+YdK7gfWjCS6tUxjR+neAlgh3LWabgfkN8/28
q+1o6Up0/1PHxEa6/t2Y7xNkogaaEP/V0yjchFxLDQzpRgb/oVqIr3QyPC8O
rtL1zRKOVvJ6KtVLr30hJ/yD0XDg9ZUeD63RCRYD9CrsvPbCf3P63jAQNMhp
uziCbxXsDqPhUL/y1OqyUGERkrYbX3PJezJ7uF1p/FJCoZzauTrYljXZRTMd
wmHOVvEMTL9tWWwZSDV6TfRnlxyc9PGcXJRpn+MvNieO6sbve9o4tQ5imYpQ
sWVSvNOZo97SXzJhExRXEkz6Vfl9eE9isgoGbFk1gS8Ue+K4dBr0QBv9b2eI
uuPGfNc9ssNCVH8ixGegU9KeomVxCR+YCw0eiN7Z3ETEV/O9hzF56eGVYJIO
fx1EXELiY8ifgL83+Ip4Fkul2ffpajQXm0ti/e1OHxHa+rP20GqLKr1loIyc
TIJTL2Psb5snhSNT58Izb8zjotwPJmq1o0xwq1JeJ1HBdNg3Q33pCYGJxTvJ
sxTYjUUwzHQodPK0W0/mouIVyIjk1em05qC2lEqqx9yGQgeayfG+2Z6EcDPg
IsVuGJ3I99mhnnSTJIBy1/9yi82O+2ep4LhTCnMAEEMnbrL51d187fXuk6mR
EVac4KxYtVWIMphMf8z+6+Y3i6xzBVVpDidBjnnNFcpn0u/NmpGnbVvZ/GlB
yLinooA/CkDbqdHILz+cozo0k02OomTmTovQCoD8T3hZVem+mxzY/iNNglUz
QIdUEp2mJP8OhFj1lNSEIwS8Aj5nWzFVp2Y4eBXKMfLEol0t7ZcKZWDzjGfP
ljJ4tvawsVTB1f0Dwn8hsqRduzowZGDo/DeMLKLdSNUkjfQL6zEJwbtw8VQj
VKv0GyS+fvPyuN0QEGGzA+/T9gMaYz3oNm3emsYEuZVdFQG8qD0YuU25QLTk
EV5GFgTwGQ4lUZA8vXmoxXFgFGsW1tbnjMlW6usfH0ri68TUXDJSe/B4fTou
djKtZNp/9pe1GEXExF3Fb1WkDi/xJwQavCyez6ShO11p1wq2+xy+Y2ZqFkHZ
YZqcNzHX+t9OEvXNdgmEOiyDavEsLykdX7HpjQdHV219GmO2TrTLLefjXjil
TvGolHU7p4SD9hIs2zeS9tG/bY8eAq+IoY8VtP7TZThG4Sg8+feyHAd4CBFj
ATXvWl/DhNcuOtai1YymEAB/QfPXVmh9FI/doC2znR0LKKwmldgvsTpRZJQT
Ak8YlZGDy6+9oiVD/GMsjqtnuLP2ZkPkWwzrpTMdvYWlG3aflPWKKte68IH7
W8TJrTOn1j2bpXcpVroTfOdtYi99Txp/mD1g4vluO/kzGlxKL/9OHDgeOiW4
G8r0cRYgjKqxDIjYD8igLodAWJpGhjQNjS0FpAJNf67n+0At7AO03vsfSFIF
mzo1/uKGLzXWPFKm8FTCi6ZrlyQq9bfHjZYmw5KE0m6vF98PgbSVY62afIo0
x6tPJ0hOpL+ESH5zSaf0mx4I4JuxYC0qOdmBHhMD2rfHIcqDbTKy1Xg1NjO0
/2AlEpU0qX5jTWdBK2wBwnx0T0GXeI6CFLfSK6GVQeeowR6vCxcxJ7LCXTrr
/3RLQuDxh6ej5+PZA4E1FZZ0zLhoqaBwLT38suOcchTmmA7Lc5kAxabhzq4I
Bwx8diHfkfQV/hYvc5jaoahihmBnLCk3rPY+HSwc3/SB28nNm3iPZJL7Hq20
hEOQS783y3Goz7fSc6XatXwb176S16wW+zs1dH3mHWdSLhrlD/20OJHzkYw0
otgcMCOpIH2q4kacXTAq5jJHdqiucYTQvh5BZHQlCW+snTdmOlxysCNKef2N
TSAoIDqiccRcv2ItsHBqhllfz4zaYLlC1htHnBMXtvJjT0wSlzFR+3mQNIAD
A2/tadD8T9Ovtf3T+NJCnrMXsQyx0l/tXYtkfPsgi79Lm/WHDQp55RVpEaCL
NP0nUg0gEjvjRDluKu0l6To+eM0S+leFHBNe//8KFQQRunz7UqlvXf2zzzEd
AgBjxjtNt+3gLZfroDUEBdyVq7u0QSPXBfiLefpVH2PcEUKH2PFPpMquMfJJ
jNtfg1heOMdvV+tOM7ZHELuxPlm6wlJ4zvxwaVSIWOVev0/5MvO2jfdDUmfS
OhHhvRF3ie5CFNSIxwaLqt1zzav3diPnxZimxrWCEMiHGXYuyA44nrTmkrV5
OLEaOiQzBgp0wnJrp8nZUQJfRiPA4FzDZFNPM8K10cWF+rFtou5QdZETZmHx
dSo3uMHMbZYb3YdfsPW3fWkzxYLDa/RQBHomYzOJAwBiRT29SV7hyURVnsSr
U7cyDHJzdcrrD+8sy7gbmdEW3J6tKSuWUGuMm6IYNPsYrKg+u4Aqv3TYOhWv
CvuGag4z53VrC9L2LVKYm9okg0hAIhCfV6SJnUKB3WnrsCKREXwCCv8vqRQJ
cx6YSL2QNuGTg8JCMugaFTpT9OstbKdyIWeMlImzO4YyA2OteWWz/YMi12yT
rC0vqNsWp+2J5KvScaMlvv7jhWgKwernKngQkW4/iO3aQLmBIGHVkBL8o8WX
dY6uPh/VXzj797lyZaNprr80XD8T1cmKIzKHvGX4lGAUxPVt6IffW2kAMSL3
zriIxqUO9JMnBWjBghVSI/rZDDj282zlyCz+ykgk4GIIqz2ePtZU8vE4Xn0h
Njx3eeximpmgMZyK4M3GzBF7W+zP2IwZ2tmr47KFzvI4uEdHuZP/43j6oiEV
s1Sbpg3BpF+ummivpcuygn2jPemO5N8cD5vrcwAvI1wqNXonv4YppVSscPIG
oRP+37tRhXUYNWL1aIV7+L5H1ysewZO7WJoaBRI5HyS90H1/OKMs301WsSuZ
FcseBYknTSal2hgPmj4jMBqxExaBUEfOfyMss6suOVv40VYFZvigb2MytBuq
rvp3eu8HjnXF9HN+Gk9zVpwCP0Xa7YUZM/qRTvj1/U5a4lg1dJHDReNMGQrg
kwEiA+z+W7J0+ds5STR07sFOJppT/Yq2P3bbXpKI/5ObxAbSVZTmJy2/Xk0j
cA7Xy3uEJIskAHH5r90vMFUk8r8YvhZ7qgkgfdL4r8gvhTttn7muqF/GMdgc
BChZF/oYz303gDqjuMY10BVT3vLUH0QNErrjCSix+rECVub9rc01Bke0JT9a
zYNLi2n9OvZqmj2ojQUTm/5D3C5pYTO87aqXqCWA+oEyxkW40x3EURs4uvVi
maXp659JO6IKuJ1mPxkrQXLXpwNTaMwS254/sReGFNu6PkGnGupQhzL65THJ
A006rNJUKlpNfgsUGAQwjO5K7XVQJyekrB8c1wwA3NuGxkfm5oDjFQj4E+/H
eEruk2s+waN6QwXIP/jY287k21KXZBtiGTbnisOqJ/p3uuP9IHSbTyXFyGDm
nW0hxViU5BO4jOOUnI8uZwb5z5m8ldd4JN2bMepOK6SxhBwChYsy3tDtPs+z
tf4sq5C4HlBASbRgS+biZEmzojyVSoFAjwL9BTr6m2ogv89l6xocwuzSSrFJ
A9x76JT37pTWmqnnhct3ga5Egh2wKXAE+84cGX+0rpye7fwQu3rSfEjlQN9i
RtHQLSMtIl/j+8VvFEho5W+v+hWMxRaubw7S+oZVVvqyjMGhJcQjy/Lb+UI/
xKTSdbdqeM3ciwAsyuCJri6AARgxUFDMWz1mY3KDvsq+5q8rhppmZinBuLcB
7M4NCXbp7DCTuNJwq1tUbc3nxe1WELJgZZRt8DrciuERXqXnxOESRqeAntCW
ZNN96GVyE14Lfcse2uo1Y6QC9XD0r+PPGreMzYA2ahYr3qmnYbRQUOyEISzX
P1cSheMtTOr+GXTL56FJkDux0tT52D/z8PQcXF9nWWfZkhHrpPEWxmif6WuL
pQoyIis1YM8atADO8mAEdN4u8+xfbd6OpRMZxJ441yTlJi8L6xAAHHdvR9gB
4rLCncOBFbI5gaGObISSLujl2wXQbBvLpgeZ9qJHnaOO2FaaoFyWYKGStDGI
8YZ0LWnmElYIMGqmJsZEcU2OGjY0Zjx4312RETfC8O4TSVQS0uFdZkh9TYKp
ONk3ca8kQMQDtCptMLe0TZocWyJ73NibOmvluUt9TOYOGg7OxfeD2tHzb60+
JLq1xDyMJqyT1/0nBhgUWD8grHpnqYxd9vM2/DI4zoUeaw8C9tR2/iMvGjf5
4A7eNRZ99I9IKAI94Onn08wlwZO+3wHL9zOF3T1Fsng/5TRvzcfQEduxVZFC
KLpn7l6yjChDnmJo2Sr3yzbViYZVRqvj4Bv9xeucMZLV7hDUh2DYUyDeJh+c
X5wXHXKcw/r+J+j6gycGCT3G5vOGhAhdEm0LlkPVlDqTlheVkvQJ8eICeT6E
cLXt72Q8ECmVLo3Nqyge7BrqlIwTNIVi7pwIkqRgGL9qqvte99zxRhUDRwW8
tm8L3IkjtNo6zkwId490JOsCanoregK1Vz4wR9m/asZwohxFExCk366AgZPF
4YU2PtXRzLG59j9EhGW0P2aKE7V5a1GrYMpGR11OaD1TJHcplYKgKYJ31/VJ
R8R2dfww8ZHyBFohMdHrCaQCq7zU/5oVsvRso5Kiex4CHhlziY1QPCvjBPUs
GorUbnk+9y8+xAaiges4Ee1nAts8X9iIlD41eBXEi4aja8FbFEOC3Ev7/MZX
06YplNR+zsT0OZ5wDHAIcPj8HfFhXYk+c7KvOJ5gq7EuDJHyLu5MqttCC1mu
saoFuW95XlXvTqSfLczlq3OOUy1YycSLuQ/9xGRp4wV6/yMumznJJupi4aCD
YMLLCZCo3D8hj1M/5ta6Y1s6qu5MAx+boxgVDEqamMoz4HrEMMTAwbtjtUd6
/tSDGyOLmF1spqgKgSjjPzQV/Pw/Xi8oJtGpdfiKSSjU3PVgNWqcwizwE2Fd
stYIO2TKB8N5nYV9Xa7RSTA4A0yD+klHQmj4egqSMCeBteS/MlAjKLBtIhZd
MXzWYp4YiJdcQBsgDolzlgQU0/bcTsF328+NVSsvitl/1F0MiMYjNoQBRZvD
B+bzPCs/DwP2ixwLMJ7J/ljevcUOl4wBzCM29MeE1m5JfRGARgeQmOnuHWS5
rbCdxjUbA3rOSqQZSSufcL2bhgg1awSOvaHUH6tLIEe1R3WBVYK/Y+ALLfs6
g7ejRVUNY9gAQuE0AyC5eBCi9x9eFppkJcXElc5twhit2gSd/DOUEsRDBgAE
ywnhVBTL0veE6/Pg+uR7sBdx15kUv8GDiP1IBjKtcrOZsu6lilkU634AYMtr
3aUv43ZPHM3WHQm15UK3nOR32mcgGLZnL5St4YNZ/KuILJrnKjdlj80ozIK7
nNbOkRbXBOu093Pjyx8bfan3LNoJUF8/KmWxA8B6VxVwmnKLMJjGwsHKEVzT
QxAOsoUajHxbf+njMYT02L96Y/Q68M7Mhuu0BWgU/gA2KKYHztxaxC3a5sqi
Z96k4ixH7723JbidM9Ux8zGjYgC0uLo6ddozTZXKMeIxbs5RGujGvjidFOtp
vGbMrO+JsKuI95gj1fcoZ7NGbE/DIbKx0DpbePSog2Jy4QKSZpLxYglbRmYu
PUNua64DuygO4JNgMNi8TE6fz81oohcR0p4z81jvxK4JfRF2ACoCf8r7pB2x
bYXbYVaYG8Pc9vcq1h194oVOtyVHl28J5xKEwD/DKGfMzSgs03306WlvPGLb
7i34ByBtKePfK/Cn9NSvA0HhzYRm20MuOkTtYs/b8XmDQIHZaFWUahqLlqRG
s0cs7036rlKB6uENrBirhowqJOwF/McrcFWEF6/99SAXaEswPBNwZhVSjMfL
h8vXik7S31JDIWRLTQYelqvEbNUdU5ltpIn0ygVgdH92LI2mdgsnN0u0eBbV
D2ygn0HZptTMerzXIpHybcrHbUT5BqHH+gzdmYfafhu3h8AsfnmwDMpiyZR7
bS7/jbJO4lekGlwSEuUoZNnrl+D8SGCiN9gx3TIi1TYf6+osBj/DDbBQLrRy
8lW3vdUbP0evD7USaj8gvhZfB46DCslhkmrY6W2jrL3i8KYINT8/tF6rTiDk
KTE3tVC5WZ+AEUCDbfJ0RyqqrHSwIwc1m+Kg0OH/5CO5QUclyxf4rZhgTK2g
Ss8Nt7KbEVH74yf6hysroxOVmWMQ64lxcd+5BTtCTJPFFbrMXCO7Exzc7GWC
T7aheUVHzfjhktFlqhXHZgpP3ldTOeD2LLctaV0vZhEcQ5c/ZhuEP2OoB2ML
9cmzTOwy6bTqj4tUQTVLs546Q69S+8lHjZrGDOSOLs+7CFyQlLPYTfDZOLO2
SyikaUdno6D6OWrX6nYnoAtS3fjVQab4KGd665DGZwzve9fKYuEz6X2FfCY+
mpI/QBlqT5ord/Tw6q39N6Szk/xiB+QwvvsxKuQ6vSPJOv6hwDNGklVHygmi
+8Gb/UZY0NOny41HTMN0IWMVzpE6H2VzNCcWqP9AlgXu5Kcoi10e0HgtXB0L
8Ti4w9lWEdAutt1y3l2rQDK8s/q+wlZGMyzo/UHlTAaXjyRqeqVL/UwrKrNB
YHAfIseO5TZcOcjUhyDddLgenMOouidS9UbmFhbmQHS/OFNeLvkDMYxrMjzs
4RWC/rZGHVFrcDVt8+RcNGHZ4wiX1HEdNFw/rzPGYL1ueWhC74AzV8M3XlRT
ihp0LsqENXq4t3s3jqkpSv0IAiL6B9yGC0ElvigjpeNGaJg46LVbSz/ZVNcO
1W2uhNhyJwwv4GySI+lnjAEtR+tqokjXh/AODEOdV5aFlvQI2dcqthgsn09A
Jp+erLF7gMlpyUM3p7JQdrv8cuc6iO4f3cFRzUNZz29iCCx28b74nlrtfFbJ
ImZ+mw2AJIzNo4O0aKPEOCqEUy0Zk67zat3WqQANCM75SdprVj+8yfEFFlJH
fgLfF1xuL4hrDpxxfiUAd9ec9S4/OEdijhqLHsiy1sg80hvUkoA7vFxK/TlK
5v0o3ag6SfMULy6vpRtu4NhKe2pFAslKhkVgw7m3hFe+K69C75KnqzRhxoh7
GXdOKpAb6L49G5WKPK/jU/R6asD1iaN1bFh4D/Cj8+cRFWznXuholvBppt/j
NPbUtLYkkIFaiz+Cy+LIzZYPNJ9r+Q1nXx4WZUy4NWwP9QqKwgrmjZwBFPfL
7NOO1rF2aHXshkZbfhJiL9wGkNVSpnl6NhvVnKvDyUFLxt75EfhieKab2qXH
kvSYzL1W/0ajmDyQFBgMIUxHf2OIJc0QP5XO3oGfoIdCxq1DtSk6vgONMooH
kltrTQwJLqbxS0BmdmsN9A7pbNTkTzj6viE3D3KScoYajVTu5iilMVSJWtgW
VdOq4xma4z90C0ZsThLctYcmqvgJCd5MSfXQI6LmBTKAdfpJI36ygRiLtXWy
PIc4Ub0jnok4JwchGUa+VIAzFM8hLeEPoYTk9PzZdjtky7J51oxhn5tUCdEL
kF99i4nl2i+zk969U6uZCLMjAyvJNhQx9+V6keIMa7kfEk3vNoGZibui65y4
Bw8IrB9hunTExNHqYN6jsCNAd9JicxHkU66PaBBSga759j20AqaAlmkfD7dF
M/TDjYKBeAB+E7OFhneCCIw9cimWAxqip6PJMXkLN96YTqzhy8Hq56uhZakN
A6NFLjUIG76UeWYnEgYWp2SC+EDxAXVCoLU8cZCMxJuwjCtiBLETBNPqVqx+
LArasQqbJhnRGgBnRz815+mO152qh05UNkETVaVMxU7vepDkeK+BbqPVAEdR
C2786BSSjxPpP4W+P52Ck2/Pbls/WwLnkzPCoIgTN5uLVGKv3oiNpYYmwewP
XQHrN9xyT6J+JvHva4ET50vXir4KGQXcPBrRwZhW4zWKtA+h8eaj1Bm7dvCh
q/D+xscXwSvXUSzEXClSa419fEnw5Q559MNxQO2NJNcHz0CjXpavd2autPOZ
tpLKxuvo0Ys9ej0Z8+1rF0TYLZBHg3TtspFoqF8f6Mr17+CfafTWQNk8B4en
enEieFIGRAp8a2SFu9uMWgyetcPWGQzeCjP4NvMSwHP25++1vDrDukIfeKrj
vyPJBbS79h+FNFrcelo0htYyjkhUA2xCIrFsfkg1bCk6CcaaOjxbWxbxhKcV
/XvnMkyBfcQhgt+RA2MqCCr1XqjZfRo5reLP0tPttFFDmbh0D3CgMxPxnF0l
a7DAd7L4UZcq6IRAtpJ2j9KLJLyclhFkn0xdCUzIp8P9P6IdVJmRaQ9bTRdD
aJH5M/wlLU7V5nhDGVIuOHVLo3hYNWS1dwf3TO9lDzA7HR2e21/QP0z8yljj
in4pkzMksupTQnKdhe/mSbjMF/r1El8jd0eurz6SBSVXcZ2WGkj50JANlkJ+
B78gv64QmdZMFH1BbQADy7EBUO5WUguWuSroqE95vLh4vMK3kPpqQzgcGdJn
UG/nqMvPOhvUBOZd5dCbynRd0zGoycRCOZ4GFCop8h4s8Aio5kKJQuepgj/Q
3HV09DKl8ok76nYICAoadCSugNkjf0RnB5E+WjFECVwqWYtWMb0DhdJCfIaV
83C2u1CK6A/d7o2e0hSKXVZZM4qowDIuaQ3u7CkTyw2YByAY+xFKFHozSvL+
MrkwhT/oD6rxE1vP78QxLakWhRoevaf3daMKvBvQIuChkM56O/fmksGTndPb
g+9Em4DTfo1cFD09BawptaNiv0nD+YAuI0NSQQ5S3xYoAjD71/4cRYY9SonL
TIwL1cAwjbitf612jSaRD/qHU+8+no9qXsp3ERKG3xB79sXV0ylASWoOJjOa
dbuLuak3iXJBvslrY32i72+whqABopn1EeX5xqip0xVC0r8UPNlNQg2Djy2w
oIDOGBRnPHi92I/g5cQLBZAPG4cs0fPx9w/9n04h4bH6G8plweiX2Dd/EsZW
E9Xj8qABwgSN2ZoetTDtFAWf4RccU1/Ixl0XQ3AT06NCe6QD8g29jsx4utEc
H2qy3R7icbhmYMDMTNomnvKdS2C74E+/srwI7CKzC+ATYJ5bUiBJFGeqaCgm
w0W5girYD4Ae/cziDA0fqSXBb1rKQovzuOs+r5+M5tC8/jtDJIexAJ3Of3Tq
Arqnh24nISmddOEgtlLi3wR11FLRD6TtN//MnjANORO0VX2ZcoyfWCU0mmgC
K0OcJ5ehgtz/50Y8HPo+tfDmQBtaZt//Mx9QSlp0kHoJOk+ApEGlE/IpBc/D
3wEQ/ncLpLOPIXHer6xbiwVNkS15es1zxKasZ7R0kaFl4l8icoH46ZdhUKCt
EtGLA2paO3f7AH03S4OxdG8bGObz+0vIQbafujbLoq4hPP5KMllHVd+6zCEQ
NDB0zrqvG4Q1NtXTYOa1J7J2M9Xme+LWxxuN7tcJ+Qqpl+v5bgipa5n4VhhI
3dvpWHBgi5q1nI70oNVaPdERqLQiHC0S5s9UppSXhfjpezkuM+Kb9eU67grf
qljdDZuF2fu7qxIy+BWsC8UNxlGnrul4Q6Cij/E1U40uOjth8xZqNI6mhx+4
jws0u6Z91cyQEPWEpLfNQ3nT9m8qaMydUnrUf4SWl6JP0WCtZnQB7YVr7zSw
Jjmz9VaV/SbvipNpkxPYbEDQv7OghZ7OXqPvpNGnABrW/sVHY5/8yIbtEdnQ
BNjBiiKLn3ZOkguRc6l30nG2RcwnK8HT1VDt2MZ2Ze5BmQ9JvvPnDq8zfhPv
EkN4qSI3UsAqLVJjjtI+p06+2c/2x9BO5ydVyvIihofdSthVkoZgYekIjCUJ
wDN7x6LfmPVjH8k/u7CicHKCdOoHg3XVvZv9Vb5fSQgivZFPZtD7vab6peZq
VaxbVd5QG7C45sNeGnv1A+AZzra8HgR5c7mddnAsJd28b6+0IhhoSDCHFyxU
F47+ewOOCDSgm5sLb+hieMEnnd/llnfXUem1P+n1l14bH99yUQvyDEBtq/BA
qJCvp56GPi0Y7mGu7Yk9Xu4LFNZ1M8SuH+IAZ2dUR3LTn4aZ9/Jpwk9uBam2
mFpJHQMCdSOSk+Y2qqOGm0HUB3Lu9rSdUGQVNT2hTR4eO++6w9TDCWNdRcHc
xJjXK/RtuM0Z6ra/nVqx2V4EF2H19rmaKKd5rhTscSi+NxvRRNyWo0Y0C5Qx
3Q4bE+JPRfpilhY+IGfZLpR5Zqw7g3ucUhJ/A7TfWEWXVfblG6GH3DUNpCZe
7v6MO8ObaOy7QssK96LdbRFui+3h56Qprcg5zB2Tac2Se8P2Q4dA7efDMGp8
b3Vkgq74Tr8aUrqWF9hihLij5eW9HCxER5DjwrY70uL9ahCiNjmK0G3E9sX5
udhsVaZbsET7hrKa2rQtWJq1rbtyQexIxfXPvB3XGkem47HGQxZtpEUf9xSs
TCdZDXK7T+B5HMrnysnODUlRXxqeI+DaJlgauRRPzyAFpv0lZ3CX7MUgd2AW
ZwbdovJBwDem3mlGjJeP4PaS/HRflXzHJkf7yCW8bhh4UuoouTexG+0jWDiM
dIb/HEhJNg71S2uh83Ve2PRLb+a6a0snAkqZj/n3uszit2p1Xhm5AtntAzm2
T4FmwMGjT29W1yF2KXE2JovOvD7899Gyl6FIkISbuMTlNcVnolnH+FBTTUTT
AAE8Vg/q72T5ySVxjY3EI0aU21SfoQKTtPejabKdrdyYY8aYSJRVVySMYfIK
xL773uWvewiYjVY8gQbdyFpruqaIAXZpvPxhwywAxMrJUFHDlBPcIYPC0gMj
1QqqQFDH0mpvyvdjg5dgWdYYu529ICQ6Jz2OvYrdfgEye3ypyBySdoqttt/i
GTMNuOK2Zl4YjImn9Bc8gL7Ef1eHJTeblfFvLDfsbhw2C4/gKg/RVa/bDPGp
E3bXeF2UFTQy/iH30iYXR4ufItzFnTC29Bssys2bNKFUeMWMCJ/XquL8FNgx
HuiBrPBf3CYjtHAPx8kxVsFdyyQPHbMdjMs2tc0NRn9xmH8uXsJU6sR4uR00
9TEq7LI+dWEzL3hfhCP0sNtS9Xc5j2Dy0tC1abVFMqO7HyAeowktMqwQBqFS
2CNMQs6uLvDfMCIbIp02HkyHG8082h4uj2BCWnEktTmmoQxOWku3Fi+4XAi5
MQd0tXRaAIHuPvev/wb+hidfTZ2cemh9WrrM9KTsCsk3Dbxx36Vaopb8iTjL
Eqm7r3txngcTlCEpMWRh8zkPbah9lF5LSk4lEiM7hILX8N7iLPBhXOr7Co+C
6LfF6pE/lGT5r93XUSCi7AaOnxC7RFWsnZV6eyI8QxIAB0cg/g28CLRPg4G/
0ABBCO735vySGbbA/Zx2WsW+wzTNtDbc30ybpOQ5NYtpgY1qNBZEZonNPiZl
FDz1KuS5cQTyyDAi9P6RE2XcFEN969f/J21b7bN57MvUvEMFMWG/DVGXkFLC
LWAMV0wXGE03WOR7iCGaToTvs8nydcfEYTGlZRtJBkfYDDjV+B0gQYwVSw6S
+oYFE0HOgmJQl7+Sel8b+sxvVwRGyOiNVP1MNE6AiTKRTJiRW4UlhQAKxCvV
z4jDh3VlHwQaczYb/cJzL3ST14sOUGXT6K8eVQDrNUTs0ge2WXEGLwX9p0Da
icQeH6mbWZ5K+XmRwXt9g/LILHoV2YskSsZWHbsXP1WFbZseXOTNEATLb+BD
9dIe6Q+0gSlMq82hcqfqmyDugH7H7vDfwsDrRjSC0VGr0dHQ4cBBiQkfEeA0
6Wi502Lvy38ThBLgWuvsdLCGV0f0HSmQFh6UpsMxEO8JhFuR6IHPPEQUiQRO
VyFbU8JZibReREQDueCuKY2zl/ZJuVrnVR14DX2EJilx9pa2Cit8k/WfvGBR
0Dm7QC2sTcxN3aFtHrnBGIRPL6Wse4Wl1olCc9fpY6ozrni439mFcGNGToVv
6M+LR2LajysiHIwFxcdfmOs3lBNjFzrswOzvIgn+L0Bb0GhSnk2KiW5y8Hwx
xVjCB+4d1o0p7yoXoc+uvM3BrApfeeADE66dwov89HW8fPW2WarH2nAomM6E
Ff6LXNH4dDEuwtuwzSxzs5Jihdy7l51h+MVjtchhHJWKHMW7IgazvAsfj3Si
r7h5WLiayKA8x6hTmQ9mbsfb1B2rta/q+l5GLymcxhMs1qBUPzFDufnIiYpk
MGO/zO9HrcaWIOSek2N2HpeGH+XZ9LI7c1Z/qqG3skTayVjUSMXglYvRrfn3
0ikg5udNLc/WS8In31Z/VHcEtLp4AoDAk83fyh3YEMeBRYEAWDrQ/43qT9pW
wFYpVRQSg/gCu56RIEHNLlpODWFOQ0Y1PHEbPisMF9riS49lotAvNe0wtHT1
cp7T6USH6HNH54ceLNFznq2XfoSZ6c9f9uiGLeeDuwzqPUkU6gExU13fTlX2
T4CAcRV0wSHzImifs8AhMRJnc8bklRtXVTiWWVcekFxi6GeUTVbRGvczVX1u
g8eVrsC8AMsZPZ7+c9aD3VTCw9DXMLlBC+5nEAvKAJBSju1me3J/aV86FBUv
Rme9YiIpFv8E6NRKdMx8xLnJjk0QRKoV3yQ94bM2fz0b4Y9YMBVvCbKCu010
6ZkgWontdzrTy+EROnyCHaUkceDcfEET2Oq9yEIBluAmNzVkS3x8nq68eu3Z
BG8o87bh4LhAUULX9raHOQz8YVn84Xcuk4mzt8nAGxhAuXj0Zh3vZL2WDpKd
ivkirw8UWuBwBqyBqlQXiztJ/JbKiTazIrp45VOTR7rF03oqxfSLgk99LeSj
psqteyCt1x4PxBhaYgQsrOCtDqyJa5KL4yiH62KMajAMdYMPa/m0ZqXJnVZH
JqNQj0naJS62U2MTGstpA+C4XMmcRa9bm4jtzt9uQk+MGREG+bzSJEOhzei7
giHBP+cKkjNeEjns1IRVFJn3FTdTJKkI6Eq+inPnWyg/PPWlhxdgdSdUPF99
mp4aiIVzk0X9L9fJSOGYtmhxBBd2fMhUpB5T6grvMC/HwNM7Sd48vG7Yw+iK
ZSF+4hFHVPnWQm/WyvaxwBbj70q9zblT8XGJSM/cxlkPWaDSm97ul/bzxDCZ
x8b4GI2g7K/7aBngH3s4EfJP08XY5iH5ZsmOjoKD7+Q6D0dk7kqwrTWU9pVi
vMXFN3+20olWOYKjiMDFgjsaaqYsGeSIgzpTpCczsCOMmpIy3RpF73qbOIEo
0EpKoF03iYsd9nQQQzK6U74drWuK51c8mk0Wj2ZzRVR31Uw2Nv888ViRK/bj
ZU1Qse1BfOVyqBe/rlj6HZFf9grh3L25YxIX/qDyjgU53zWeSEUz4EMAHuqL
Bq7b1jpeCI8IIsuSwNZ8sr1CqZQf0aU3qLjXcFufIF5PlZnq2JsmiOMaiyUM
2x4fCUDkukKvpl8phw8eHbSV+UFNp1BQ2NwFjCaoXCaZcDG9ryo0RH3Q24E8
7Bh0gAlAvMWqGmtwYqbim6y0u8shApR126y4YIqD6En4nAqiXuuVf/SUimmS
VcyO6pbb6q19q0ex4Qv/ppCzpKKOjmT07qXmZg/XAazjzUiTPFI+CaKleoEm
5qJGVAuyHocY/g9BqfFEjv0JTQ4YxQzwDj8wUzGXCqNRCMIebDRHGSn6npCE
OM2DqSSJJ/6mFtu3YkWb5GW98YYrqwF/iV/w5aYRd+UqCT/54XLyMUrFj00i
SE+mzdgkJsK45VCxbFBiIoQDCpJrxm5dINuIEyIBVEcB+R8/ATzsM2tbJ3em
gZ2hBq0f5jmsL919mtLjsPtTCZCY1CXtY9WYQknN6N10yO4vZvET0/Lw+055
9x47N/jRgJRuYc/7+DA8WBfp3QtlI9VIj4tMkPAqHJrAWO/geWvUBwXnA+lD
noiktIzFJGxgDUgPbmVQAcmFzCHaKMy0iLR1T970jtCegmRc1A2ttYPDcWb+
wr/tZS7MMKeouV9OxdDolXEmVIboTfFRGPVHwnw81/4IdKOiirrEeAyOS1nZ
8WL/rRgTliuoC6k5XE6Be/o2BV3IifKYxQDH7//KlEh0I7eufOfaKO0rxzaN
Tx67eNcViVH5s6X+1sO5Lu0fLYtNoxqEJsr1hdwNFjIQc9i+J9L9Me1EhRUz
5iVM9n3Oe/fbc3+h9NtXiBvWTfZRUN/GIIfWUAHoGLAdBO5XkQYA1iR3zGb9
MJGf+wvwR7icJC/eJpugKAnyrE+lvA3FaPWfCVZlKoYWjxVXuQhFDx/FZ/04
4XMR3ZyoFIJpKJY6kZxhxBQb09yw8s9yhtWKMM6OSR/negOqLrrO/FzHXBFL
e5RkxEeUyhv9Tncq2QfWwzget0EBWDaClntiX/Q4OgP7pQCBntbhhk7qV2vz
D9kP/sNRsB5sFi6Dfh0CinRo3Sd/H/4rVRdyo1jIqWco9UYuNrpSYPXZZHmU
ekWBK3QAC4Jhx7Y+1UbO2+tdm5AWRLujzbqHGph75N30BawcCwM2Qswvwda8
PwLPvzojBhcawehv8BpiIq6uQVcImb+lvLUwfkNZiYWfqSFEJImJWDJacm/0
xMCW3qm2CUYg5DUlrcND+yfUPjLtac9o/u9UJRyyYVNHK5gnDU9Fue0PZJUl
UkM/f81V0R1BenEa5mfmg5XSbkRFri6L8N7mfjUGULjoSB6edtGMpDDi1Vw4
pMX64Ev+OcAxauaT1A5mBeBDHQpkHWO9WyRllB5+My6Uc+Dq3FwGoCeFpOV1
MRdIzTDW5/GwDoKnDYenmBegCLkzi0SpWh/9lwpF1yi7qIMCcoORcOsxR5eq
E6Ag0vBzn4x/6tIxwBjCk/3cpwtH/0lNqXG25LKDkygWP1oY1LHnkmRIsngc
fXBqDbqe4w5/eyIQXaFRYycuEsRz1yf+diLFQvgtd5AP1oeqUCnGxpQLhwI4
TQdD9qZg2nXygC+9bYtdQjqiS4olLmj6wooKpdOgVZ11dbCwBVH3vjuVlKz1
Lz3DmWdPqkEnxwVW6B88QuvHHaM77Ojsqcv2l/UkWNdC9qwglQkHm1qcfFKO
UudzaiB/EULQ4WO7YDn4uizzuaZ1nDWh6l/T/viLxEVeapD2/G7GJxu1wB9o
6BdR4/upy5CBltYOPgX57rsGnuGURFF27/yiul21IZJ832w8Gn2AunwY/Hod
r50BROPTU078PIgLPBLRwwD5R9wefiuZqQpwKQ/DOWUZ+fLwqI2CAekJDCX0
BBcKCq3kb1OwtskOktqW5xIkiVaDVmkEbB8V7OmHvdVVdIw/s9/01AOqxouD
yWAnLsF1rebh9+fSEl1AFfr7IT6meyTxjs3fhcVbSsUmyiMQwnPHH3ah4q1z
TEEwLFOiUUmUcEphANPm9dtv9YEE+ZKCpd7bVoDsav/R7NEiegcb6FamgIcf
mQZktfzTAgCzv3kupcIVnaA6Q+l6QtQ34mFCGCB2S+duV5AdRebfTZyY8iL8
hPsnqa8E2yhjMvYqHd8qFunBWlDzvawks++CH7Q0eMpF/ZNMAuYHFmXHOYEb
DMzV6I9b0/DpaRkB2tB5rcVcRLSW/gQ9iu9LTUfAMPGWnEQIpupl6GQbPkts
Xo8fsqIzotyvshV02GpNNzzI7djZ7VJTWuK41XDt9UoCn+4TKxWrq/voMRKN
iyuBVHM8vGMLngExozCJ/Q/j6clpqn8SVFETIBxet+7O4N+EtOZ63a1SZhGn
r46TPiQ7tEBepfGUuUk8NGmHyPI+TGKuJlYhP8eh3e+RBNQ/XUvhpCZf5e8T
B8vhGs+WA6TRWR5sb7JAYFsQ5R72F2juz1W15At9uDHcuJlwg89Wtw4YKbnx
qyHDhTY+rXq2cK6a2XpO6j/mIWLnpaqw7hwGg+GUhcNlnEKNSbQDkxXSPOkT
MqaXHRhaaYjuE840QThD9WQrW4dsaL55hbywDIIC6YLX0fZEBaWRQwMrBwzA
8dzFGTO08l0kjsZHnbDjpEOURMZDCGLNMQnkBE9UDuQp2zHlEvhchJ6fDT+L
j7oGS/EtGr5YOG7Fronp5cYZNAzV/O/BJVQ8IRymAzs4vNOPClhvBooWK0zb
3vxPgdKbCl+fwJLQDBo3cVVnXmD3V1WCnRDznXGf1AFRU1u9aNlvB23NCFy9
w/Iacu54faQZEe4Bb3M/JBiD+3k0iPTCSNC3UK3KJOElMuLczXpEDgpCaSgw
hjQyVj4VkAoEAN7EvDJ+qK9V4PiHpiRNSiDhJxW1JM7qnZs6ICwI+fd/mVF9
H3XACA1To5WALaHySbzdP4hZ56xthPpKhowOkPnbNpfWW9GFPFkC9yklcM8h
S/i3mgjqUDdhrfpcqVMfZlTtWEyCWRQeTQAAc53cXNI8d5DfodU+1QJo8W9P
uBvvfgrhRCJ9aRz4+9qWcVrPMrLkqa3MKJsVWGGdVr/NEmw5eCdnAU7DI2aa
rDPuNsGmFm+49TF8nTIkf0TX5T0lku3uetvY9O5ccUf/tTAjdIMrNLDlLwMv
GehSrHNyFoMyZtNG/2OvpuDG/pJzEOobJvCSjxeIyv7iYa7KuIjLE2fr+3Lc
P+Gxs9A3vpxilRFy1YvVPi/zSs8jP6fTor29PKMjU/sMVbvGOoP3OS5yDSR2
jK4TCy59qVNL3HiNPuHCrP7lFWeP+PAGGTmgJYOk9MSXymQZKI+Ua/1OEuoC
l6swG/RtNk0FSMI34fyHZFj2QVv398PfzsYFnLAjulC4dGpWuye6a+Bo0Vd0
aqoyOAWyptPFI2Feid9fvk8qfwGKQXr7V0gEDIa1tUt/sygsCxttnczC0+cg
TF5EvA5Ryr9YuRP+m6jB/Io/l51+f42gRGWRajszxs/dmf8FJd8NGiJbE3Dm
l4e72JDnHeeMvU+nA/RhG6joJVKSyiOi/3VJMrgvIhbJxNp5SYn8+s+GoVoR
sFLuB87oXTKZ9AnZ+zbtSm5oG1trdejUeaDhFTE1B8R1BuplaS4DvCMqzDJF
NhDDMWwJQb1Ay9o25R5UKQ3a7usbWodLp9ZAZJwqkq6j4kFjdnKImP1w1Jz1
FvBqncRdVkKWxEUZzT7/0YSuw5xGB4t9E1WP00WpNAXh2M2vD+7ScYgkwDrM
W276igeEyRmt3EgSCD2dfkgjVo3GqhBjG8lmIVZ7cKSVQ/4L72JnRzkch91s
mC8zLJ4+opUmQ6Py4kQfGhTYYgJGnwKmpEUZg7oqWTh/CaPvXpUJhx9e4Dld
63TwxzL3i2gTSOxV0XEAMC9KjcR8sNdax6MrImZMcMcx6moMoeD7Wj42Lc7Q
v5XclFLV767RMnUIvsP3QGjhkba2X9dwoOsop2CA/f1q+PZS0usWqMgr5V+c
WIf00aPSsZV8W8y24PH1+4QI1wITgQfymd1WCKuZSqQ9wJq3CPVxlk/gVYKa
obOxSKLoVCVO9RxQ2pNYFexl7Rhh4Z2OKGOUwAZt4c8RrptjqrWLhhBnFmh7
h+qhmKMLjOU3f77b02K/UKfL/2/71DpMCsnk3vEmYh0QuRyATNzX7/zU9Q/V
Pm4gnr4jEF5rMAWS0wh9AwGH4Tcp3Qm4Qwt7o2ktvdntRtMiW1ejKv/CCszf
NUQJE+0WXeLIlEFyrrU15sWpP4e2Nm6+wgprykqQ2in1feQ3gb0Xg9pQuqOD
9YoFKMr1afSYiJtn3S91mr2391q1SfxCpoEwzEiIPKuN0pR7UxnR1Cm5KCwK
NDDkXvxJSiMY993GSMwgtKritBTM/bI/RZaxZoLJccFReHc6iaDs6A5erPLt
Hwv8iaoylKr38dpYZ/T7kbpoLAI4mM72TALST8Q/wErjQ28nhRttOhAUOME2
BXvdkZFXTALMbYKzfigJzf80g4j6QL+ZDB3LflcvIZNS9O0BrX2rPNjFezIK
20T9fYhDYNzdQML9Uh52BmTan27ARdSs2QcTmIDAOSSt1gbaTJnwjKmvOb0g
LQyYvGXTnvx0UR4GUtYfX8gaEHryEd+vmyemR2gLDeMgsD8h2T6KQSkbtLN1
UuhrdkSbxBqwkLKeqaca7eDG30bN95CI5Q02Uw08UGLXisrqroQhiOLNHc4g
iZqbuhA2DHjj7+h9BcWukdm7RcEHRKlxnJA2oqxaTgmROhtfNcOcXrQ9uXeK
iPF9JIEcrZ5ABZr9L0cJFOqFSWli9n9mBN6zVxr+A9stNM3xaCSfH9oOFj0y
zOsMtn1dSWvBZOcgavf53RZNTBcLk0kyUjWsKw4LZCTyix/P30/BvsYMUFil
v0QOMLtjNItjHmU1NPA+LxH0ZQ+BSnP2U7XIuXILiO/D2k3mEqNBZ/r/5Ih5
S1g6Tyk9APsQnYg7LLk9wmkc+zl1wYhmU59hd+l/Rc3Otm0mhqSHYyL0Mjx4
rPiJoUnkvVzYpDpXQza33056MQhNJOseDEqmbWQpcMKqMue9IA+JxMIE3qKN
xG+5bIKI0LxbYNZNRWBlbDvJt6prutfuQUCgWKRbtggJUvCgounL5WKrcS3c
iZtmeis+OORbIrYPYEQfW9yCVMXUIHJcRV1ov7+RgIENAqhsuOH6IS7oVAwo
NgKeG+m8LgkYxpFJTTYT+8ZN/mFKA9xh2akRgXLPIGEOdQjxdCi8v5I9t9h8
zXwzOJaPhhT0UH0aPDnnGI62z0XEA+FQXEyG/iKGmzIQWJSjWZe+glfDoUcr
zB5xnWvqbMQ7ew8cTaw5gMf0X8ib8wRHozOh9I3fHLlX6yvvl4NuLxNMF3aI
MBV9AbF2BA9yV38tvoezmX62EJU1KiJJVrYA2OSd22EhQKJDTxmPKb2LG+rB
JX4//O73B6+LqwUHvf0OAwR4mmscm5A7XeI+UwRhmh6hQYB4/gp7dl/thz7e
5X9K0luqAe4i9KSHmE1SZZylKdetoIKC3lTQ4bt2xFDuMGY9U/UGDhK4HfzR
KA+FxNRA7Sq+v3iyCZKmyb+r42TRsPlRnFimU7Z6w9QNtQ8Q7R94GjqPlUzI
yT6TcVkKCOGJwT9EEl25LHKFpFOUMdxOFebdfwtSARFiUdEcBFz3zkJluvDD
RTZMspwM11InW9KOmsN3kKtkw1VFHgBPybpQPcQrDLQpZ7iUDvfRWfl8SHTw
QGgeUjlx4/2ahNvZngA46SJO/lV+Ae2LXKzFmJv4Afb6Jk100rErga9yc8L8
lYp3NSLiZkudw7Gm2rdUTrqaxUi4m2vgbL5BO/EvT11GfhCMGyHqFZhTdexS
IYO+Epu3Oz/PS7SniN+4DVks9L9Fx6tw2VDUIwxaCU9nt3AkLobBj0qGI4/M
qm1lTEdAAcz0gpuA1A6RMWUnJlPwPPvzQt5fj6OIzvcy6h2AnqQtlZs49IS6
p3Y1TF8SpKmWtNvgcSDJcyriVyuoUND+tU9NK8/JxS6X5eiLq0tJHw2nHvVS
K/ht4y25CaASDIreG9vI6Ynxy2m9hOGn6f7P/5XwsGA/mb4IiIAYoRN/BmE7
rXJnBhYCVX/TYhLCzXCLUbWKzyKNVOGiCvFJ7XACOyFQQ5oKTGMQ04Lf3gYv
YQb/O5gqsjNM3p77IbKiNF/nJUTcBKHG2hfaB1BI81giI7oFemE1iWqPCreI
KGjIspHIBRm2FSGs3Ux/sK6r7poMcDpzrceG/iCIKAiQT8qgbqVmLPg3tLWS
YJAz/bhbm3URz0uIvADljQHbEfyU+Sb1EOfIoztnIRi00u9GCCTuJ8zIor3B
MLrr4rzrmTESzGMSpdJjLpVMwV6LqqRWrqBfbjFIUZLPkX16/h5O0iZ31CP/
1jNNzHhrPK34MNChfW2cj2xq8imasyUrMmx5S7KtliXHGIlzFk4twt1yUU1z
7HnURWEhjFklAxA3DfV6p9ubyGfybMfe9qawo41aY1PSfPsPfrUZ3yGYCxK8
6MgzHVPPxUg9s6OfLO/F3nEWyXiUd0WhWU1bos+eQ4173cV456T/Seep/20o
EHMYWFQGCw9KQjnnFF9ZgjQ2/L0WljFtJv4Taov2AT6uRUp8lloCQJLeyqZp
TfWRx/1X6hLarcane88dRccHfDhFEafcI2oz5CVi6dOS5NIm80b/5cdceDp8
237zieHNfGsfpvz4pszp+ppyB5DIiBXD2OHL/3OGMltF7GmAWhfbiAolYrmH
8M4fLy9ZV3MsQBqfIieRS6Huy+OTQi2BYYfVu4AZ6ubAJ1Ngj/2OoZxxrVJT
32LuSVPVRnu0oKa072pTwszFfdH3vQ2VTOT3t5JaEW/5+/H2QhlLaIy45jtP
4EJWdntEflKRL3+fOvQWtjyJ/rksWPp77weA8pXcoUb2TsUWBmjGdNGw/bjH
2dvL9nr7kdX+lKfrDPupKRPzJpQ/JOE8MEMJE/zlHNK18554x7eJReALssYC
jecXf48deNwOV/SbY75F8S9nYciG5ByRPo71IzK10LCN10w8YMXWzH+Eqqis
XZeuUNbUHF4OrkCCZ6DGS7zu5WEt0o6zbCra4RXTHVIrmizA/iTcNrTssVCr
yoqnbGgUqimlmh65uxm9u06uc3aObCqSSt1HvpwGwxUcwwbuuzYePmkZ/nMN
5dqJWj237Cq29IulT/SQ2JJyugMRuOha8auqrQzCy4MNS5Hvnz/G34f4AwcN
zjHV2kAggHgXGZdSwMj1ASTBG56xCxPyaeQlerHFfgBAVRbQwydYRgrUUmdg
FArSWUFhEZkL3N6UCt7n0OvJoD5gDBNFha9UMsCO/88jgRvSiFfDavIU3Sbr
ZW7NTrRKTndyyjXnHCLYRnAG+uxQ4obVeVXjPHoTTau9E7jTFcMdexqq95Y4
ZnuRqX+jyDuohEMTwpnlnlUEYHf9t0kQfpm+c2gT1F5YmZmg7uiKZZVxeuax
nrwC1YB99TSxwom8s1ev0n/J4I3KeTz83UfURb7XyRe2vp6jlsZcLgx8+gUQ
UX7fkgE1nuBB3ERc58aaXJdpA19hDDqaRszWOeI6h8Qb8MseJBT68P36ACC6
pYNGpI0mUOfGAKidtW+fNL4F0sXKorKPYY/C1BThd1690kYmei4iwY5jItWU
3VZY+UQlKhsfLhMjSf4+NeUdrUHZW2lrBT9FREMNjh5QFOL/MY1kwoH+b/v0
Vqz0zLr3fO+DRVgzNN2wjx5qbRPKjEstn5qXFxXkOoqJvnYLYUqfd6kuDY+F
Vq5/2elp0uSWVT1tMGZW4rTRJEatAhw+kdfvwN1Xpitm5OXrCw5vGLrFBBgy
tDcVr9OI0QMzffKp7NeIgVcFH4HCEmiCWok7iYg+8284JkjVL8EXqLacT5HV
p3gvTFvJnSd7Ub6Ikxp0sxZD13S8l5hxGz6DntOpPQAMIEPXL8vTPnGp/LL9
Q8ASIgZheKhk7montBw4Werq/BW/vzAHsf3HcyMwgMD+89dzR0lcX63P6Etv
GAAeRF30M7+9cBd5fBgZgcPAPY9AZ7MQId8P49Z4iN5ZBHP71JjGZdLPQJD/
t825cy0r1pcwZSpPULXK46WRUjSS+OWd3KDi+bsVumOqFxXk07Fln/YHy0EB
eDTJuCAjY5nzwsAjnAR2zYwYVWQtyYF/HT/w5omHvU515D2sRLpX7PjIge93
XY1HaaNf6L/EJ5iuyWzZIC2uXtgUZTAIMFvceCFIB99PjUGMDh8iYi47qmA6
6gJi9yZ+tlkXxdWicSBmkV9sHj5/XreWWzyTaeXy4vndgRbFnBIA5rgMhFiS
RneshUdAKd9YSPQafilX4dkskYbk4yhHoHfgeN8QMVgf1ZxVBw5gvrxAWRjl
fcjpTdRTZo9lu7sJC/oBZr1VWZg2WL1joxR3rMy9pfwUVcn3+Zn8e4ngMWLO
zeL+ul7KBltxJw72NnCyrzGTMAini49Rh+YAdsCLi5t9taFlju8s0crZ9mpr
hc3fSbC5oN9EdIPuK+7428vKf5hdE0nZu76rkgegqox6o/OujpW3eEOe+1MR
78fIHUwc+nd1BL7N+M34fuDmoAxXmLlVKgu0CRJV1+lzbtz5watbepEY6L/h
0lRieBQ2ObNKkDFC/4LyEbht4nfVb+3XHNnPnEQBxHc3ruR83pIgl+5rx7Pz
6UQz8OCazPWVTqHOVbVXAX1FYVLIkXnXpp2MlIowcC2Z/tVAyGUQD2T8Zi3s
R/4sjA3tC3rjQOo8Hkj4HCql2kXanoZuNfNHPQ1WZxf568+J5kuB7VKbOJCJ
bM3P1XbrWnr4M2H2VB5fFWM5HCXSioGrbhqD5S/BYq+FjJlgorXa2gLEJ5lX
Liyn0GvqaR7vkjUfibY4kYTkL82i0kmRCOME0CprubBKAPRTvLGfrmgxfW8o
AxyLASQTCo5Q/IvRI/xnGoxPqnksUbhFxhcllZL/GTEI19ZXwOECkCqX6mP1
+ZTwCGlLIOtxm+sYX0PLC5sH5nzTstlqbdkhw5IDjsE7F8qd3m8X+mgMGjdZ
y5R8YWEb0w8wlFxj6olBvYi5RUyCTboHq2s4zMACb28bF547BAC3UfJPLQY0
SP4LyohG10pWr/iRIL7ZAkvaD50AeN1UMiZCQqMfC0NmuM9aPTP1cRCZiP2V
dQqD/t05eAduWgBuDC67mAsaxPgt5VQYaehb8cFufy6cWP53N05cGJJgh/t8
m10S0oiXuBnKWwZf3DyHTRKHU+W2keX6LlK8jsl99jjBaJ6EzJ1m7sBRleEQ
mVMM3Uq45mutHL614P8mBYaeq1RfecY4HE1y9iPRnbt/wouY/+bgpC5UXlDi
yNTRMwIZRQPhAE8sbBzwUE9exnJEMMUD5g+a/inBgtYlnu10cgIDOq0LY/vl
6E3orCG4/NM65eXYQJjvfOnoKgEg65BakQDtiWtWKsjcHxwvYI+tWBLEChQF
9huQYLRnL1NCxgDc1WGQcarq6T0YPzue5FAgzX6Xmvgod63/hHGN00t4U9TX
Rksoj9j6MX6KwuTdu62qJvlqKfCQ6OSLmw/BnwZ1RhuEtVE6sPA1Ybjq8lmy
7Nu/PcQPlnutecXcivskb5F2TuQtke7QlgK1C2CZTPCpTG9zwDck+74l1tFZ
jAFulZcbm1eLVoXa8Wbu4yekjHK2g7Ps07lZeXGAkQBG28u9/SKVaQGOZdV1
cYWAHxzncdGYObnOCX81oVtwRTZNeMTdRyYSIyNmxqKrbF9Cf6ZW09bsmxeH
3kDKv/Jm2erQ4lC0Las/fLXy+2f7NUHpHxnU4vmMFNIvFlLNGVZ2pn+P8T/V
iHcwjcz8GwieHlkSv4CUiEnKGo02EFEHuz3FCjLPCjaBrrvEkKafZXllhzCc
4tIg/qgzALOR55cpzSRWG5PiSMTjz0PAfb9hesUYQkcHKTGp1xZCf5rjV0kb
drSfy4eBu4Gw0GS7vGJrbCvSYh8lroT9fUuz+lES4448g2mrwVCL2NqNuvwN
x6tHOqlNQH8ykxL08wrzRpu9qLKsKjjBE64nmOXo3KLkSdil/e0sTyHGkYni
nDCk3ISS1rbwOAlm5SfyH/sDhEcdcom83ImJEYeCLT4KjBg/f1Wp0FRFYDTp
Au9T8Za/0TIPuVbyNY5e54V+mAT04mGcQI7bvtOJM3KPw3y25QbAL5HuGD6s
CKYr7raBkW/Z+e3RhOrRQix4Dj7CKBuz1s0Z33Oiw35opvjzLkevS5r9IywX
5bmebIKZTSPOHP1q2H0hE6d66dUNknF3dLzmecqQ+SDa/Tc3iC6EsElKqzm4
U1hy5tV/Xx3Id8ikkueEQmTJL4NLGPPM8B32webASrWnrbogJMf06qW0SBH7
RicCXvg4ziYZSzYpZFkXB5chdbFidgoP2ml39X+/43+Ay7lGsBRdAj+jL8Qd
W2J7vD4F3sQ7B3mxmochjzFiata7MZx7r+aNlwq04bY/NOj7XQ6uAZkHPUki
AkdxeAAoS8RE45pF+6Jil10TVOnfjtNCW2hbGh8xXfdeHB56FOII2WrnBxPO
LWO+ybLUhmQd0pRllrfm3McgESPMCJKbhbaCfJao0ke4pkKy1zTfYYhJFEdq
hr72HgIpfDYt+toefrN5/ToLw+veYKPrDQYOkjyY6vEQOdmedB3Dy+pwNoM3
HdFmMCYzYIGUqlfN7EQCDafiNmhZJatmtD0p47g4uZejoG8u/gAnoSLWVAqP
z+N3m6bAJnRqWW8PyuTKtWfxkn7bGAMI2eWQ75IHExJKGs1Iu8o/2l5kDLn9
e7o1gvKpW3p3K4TAbPrMw9bZ9S5D2SaxUNF6FOGKLsiKOhn8epGZgg6Fx6oG
w4NwKZhRWFN7CJNLkBG6S6DWrBIYM43aLNyW9yv7Wo9jgW96WJhZXwKVSAeg
UGf6knnjuVfm3FbNoL5Hq2c4vwlDGfORiSs/lAM/wZ8sPPVvWUfR/k/E0x+/
ZdyjMQnGwWSnK+gwKoUwdEpZafTUUJcJvHAbB65IopFseH4BigCDLtkI0O7K
93Wv4I7dvNWA7QGBie7JCbK3Gj9C82gL7nz/sKj6nKQu8ytafyQnb9HV46qk
ExSIkp5QZeow2gFyXdbrjR1mKacvUlo1aZMHQ8lobRiwAzve0jAg36WnoEri
MbTyslr43YwgyAZ967/oJ5R35LfWTteAt7EQEWWrDvPpt2pB9yYWSIDMZPbV
6xw4YbUt7hfuna+LpX+InR4lNWP1YMbQrTh2cMc4U3evAs/6VTXIT8RE0lyG
WYNJNCHUFKY5Tvh4ZPCakWlBqk/e8AsRyB+4FVcNIaL4fmSreW7iipUsz9BM
GS9CQJtue+sa0+0Oy6PRcEywDEdXcuV3l1NpnsLqF8F0z7mhaI7sWgnHrDA6
gpyGXANqf/O/laIv4V+R30CCSHGwbeUlBJfoIUQMUH+mhDEMk3HsJ1CwCP/y
q5SEkeJonnuGGcO/lB2BYii78l+IktXzwX6lhx9mPzGUibfDt8J28iKsBWgn
Wawivt9sbB7MhLxi1Sh4hv2XX7uNV463jJz94nJ66f+14zhAoVuqZlORD5nz
RU6eTD38oQu53HAHYyTQ22px77hrboIuTu4R3PtKQX/nVH+0TgTIoL1BwcO6
peLQsZzYD/4usurjx1eJ3Vb7kvw6IQ6VUu4+t8lyilI2XuhBrJ9sVpHItw/7
jscs5IyjfBUIJv4SyIsLsijLvNiYJTX3h/JjhJR5smFt/VXiOjmldXL49pgL
a09rfZv/NJY3PZbQrY/Ze6xAmOFL9u7ntznwsg+Cyl3+nj3nVpDs912n0HJC
3b4oexbkB4c5LdPty/1W5py+GvXaH6vJTGGgWvnQYDItf1zHrUIFvCsSOIP2
nxhzp+tugXFM5pvlWlPZk/LpUG3tibdLoqW0vrIc1qR7pKZXZZ0Q7WTCAxzH
/CaODpWFotRCSsPb5Qn0I32vYvmLxdFeRYGhFBYmDRruSx4mnGVNmVVhkBg3
uew6AugtW+gW6aNRV/hkTMZBbeS40zmGpg/oRmz+nL2QpyDQR2GEoChE0L2n
hxGFpDEA+m+Y44/eVoWDw0rsqMpYrGfty0tw6G3R13pEmyDLWlyj/LsGJEdN
yCYDuaxNuIrvLzjjOiRL6xfcGAsUao5OYM07eEslTVJIqhvb9+kd3cfF2QOH
qlBEIid7o+DbiD4uErLdvih4GK43JTscGYXtKWGjhmgTR1iJ4gFev1h5ghLD
z5l6HsbibhVBws6zGqoYtK8C+lZ2LuISwOe2vcn7QR8XrWbaP1A6S3zO5Xdo
h8Q3ggs/MDuyalyKmEMLwGxGivrvbKU2oBEUVXZIcFSiMbnWY8+Rc4g5Yc5K
XLt4KQLvvzi372pTtfmnC1xQmiIQ2gPXPUBdyd8FyL1rE2TLOFjdTCT5Nhwy
ZbmQEGBX9DEQbIiwogtsmd2UTEBVOadH81N0bYBy+Z/S//jQSct5E12eva7K
xGTR13B1wbVqTtHJZQMJrp9XvWlvBCCRT/lmR77atDaWNxuMLWPG1fk4liia
hvLHaYUn2L4tVu4ZcTghgtM5tVI02QPcmJCfyycERPtJABvtgLboC1v9jfL3
g8bxT+tiVugNVoBrLnKd6RLgZ6LQOq3xEgIgElzjEpKFx4n0Pjfk4Vq1xl6Q
RcuHI2ImXf7yuNqdh+RFO+sGpPBGIxevLsEAeHVwv3/HfjSJySMSjBfBFvBk
WxtjUCrOn1xBlgoP0MiOmRgdOQozmGbjcDl4nVUIDAQ0IYhIhyTA9AsViSP+
ygwSrrPoXxsygLP6zKpr6z52cYQlZPMsNQd7Ju7AXSQXwmBdbOXZThaNxR0z
EtOC8DL8hD7g8tTKL37YSXfp5U0jFKIrK9SOQ3fp0b4ZigxhDUVgXe3RO884
bkyHOrNjbuycE2ivSta3ZSooZ8/JGuain9B/ydCoRMlWVyTe9BPtbo6rb9HN
aOGSUORAXnVHFVdB6Ipnm5PwNrk8P61h1oiHWSYkzIJldc8/ifecec0cgZUW
LOR1bi6M97ecrmOf/1TDEnFcOkfYxfiAf2RW/2l6Uwb32jeS1Cay3DEz5njo
6CF0V8bVvnDkHVwOvWn4ClbeI2WUEorU/cD8gOCkoOG8C1wVlBW6IlybQt1/
7ejtbNT68IoaMKLfZGblmNFrozbEJVX7UFqN4d45xJCpNTg1k2+1sMnpe87k
/j5dj+VTz4fg9EYmGZXb8DBUy9dQcuwB9CM7z9aJOOBILLSntrIHlxo29osI
L461HAnFKT7rDHYGNIGf4Lc915j04tyM0WsDFt2Q4olrZXHvceqMMm5cuDHZ
ap+sDuxLhKqX395NPofnktCyIcw5N9ePc85F/YpHny3mt7Yf2CgPVJfspV/1
xPb6mIypXdb6iL1kMr4wkx67rZeLOHDE/rsAu1VJgqdkS9Cc70z94kUomKZK
2xcERSTcjHq5Ol3JPTkBD4MF+uigAAtYuaK5yHMxtytGcK0YQLjMGTKh97Cm
sixxz1bY1rO5stBIHzO+QsLFAPF2BRtrGfpHwsUqe45X6+prEhQ+ShPYY2S0
hWkMuhnZsdPJvssoKCUvwAAouV63dtjt1hyf/eGHUOxh+NCCqaUkSq4A7Hqo
C0S/VeOqxofa/z9gvEpZW8OEJsxH5FgeD7QI6YjGrodnsTpZ/OO02iyBzESz
2Ngb4Qg3VX/5HgpGpgkzH267V1faD+OkMx2XmKc3Tg0gNIDERtVv+AIAtgCU
NNBuFjqdFkVIjftGxpFXo+P8R5vd6Zr0pVDXU+ti3JwHQ0iOirbrFH8DlhRi
RyggpMVqQWNAGk1fHYZph7IXS1MAvvZV96dGUqhKQSXdzYJ7dmj2EbEZ0fJv
JbN8q/R4fU0fm0J5AHd7YHvqM69Yx2im371g/q1hOzLotTZbEEdrSBtLsrqa
y9QaiB/lY2OIDXFw5SP6jE56FLNnGyF2l0jlwoWzROj0JLYmkr+R7pmLi+Lm
i1gQqMWawZSqz+OzwQ37cZQnZo9jX8957KeLstebdyuMVNXB23jcZVNMWBre
/XgluNO8HMFrMqDhUnhtzHTGaf3CTrR0qFFrt6iwKOuFuU8sXhVCd0eIYYNP
2EjcIgWi1OT1z4n5WSsHbjNUd2R9nl5ZP1+vnW2WPLVlzJ36qziEBFEb+yKI
xl+0kmoj3BH3uIYS97no+m4MXKbPTQoa4IV9W4/YQtOWIRS988Cf622R2Y0V
z6INLWkjeZg811fJY21wsKj0Pob8NNTgvW441Ck92P6vgpXya7N5zIcypFt2
8Sfr/+5nPUQdrZ192ABE7asPwg6YK5GX67WfZ+ovZvAE0/1jdmNKJ+8Bg8sT
zQE8Zsym2Zmh0bUPWB/Bwde7TzSP4ghaxV3gdhCO4svTNSALjwg9CHEH0UFx
11sSqE6WcUPp4MZm6b7jKUCeDJe36j/mUoIoBqLcGTzMmOWW/aNe7fW1OA04
qBofTc9SvwH8ufHzjpYkK4yrEzmetGp0XmiUAevf1dVQb3J9s3JtJL9SYzbT
DkV3dEQFj65CQbG+gQMwUt+fpEcvdDlU9ipMMXACssBfhvqxqfYv4rye6TR9
D9Tvwte0ZiwrqRCTgdW3YF5kiRwsrUeAIjpZhDteQrcvYa/oZ2gBAKhGjchs
b5E2MG7Wq0FXyGg2CWQtBHiM5S7dk1FJDK1QpahK5MEl9cc/uhAP4cPxy49f
z28O2kYtyqUD/kvgs+KD+1Ta43lAhQZMhoU/Ix5vKxYOOIyLLji1eCK50OEC
YQlQaBNXGmFt1+EAIhXB/nrSMsoGol/g60uDSRJCbCNdY+wiBkknDLV8mDwo
ony2u3/x/jQSrrExHb4nwHyHS5YtiYvwqBpTbc2m1uniWoJr/gR+Pr9793/4
Lg9tKgWEZ0to3lAPBbzDMeZ0gkMGCmPFFB85UaKDGSDHbpBd7XT4VPisKsET
/BD1hMzRuCRyGyzTa/k+3OFTP2+wdLXB82/xHM1Qm28iIkUyLk/8yd9UAtmQ
xqhzIGWay7HN8z5EU+V0wDwGCYXKyHOj47sj3bIHOLvXTre+/6CFjZEy96+p
hDGKNSM0Vb/R3S788C/hdbaC3iLbu9WMEsuAEXh+a5k24khtIiffIdEiLdyR
EWQHvtax9xMiemsX62Zysi/yeaQtYioShfOVbQ5NZYlCpgdfz/Tmn7pzIwjR
N/8/SqLJs/hssLzE/VY1mxTRdccDgNR7IQicJv9VU2Q8iV1I/tVh4ibfWzzA
GsgbioqNZ359bEbJS4Hou5Hq5mrVdV+VIzHiLE1uqDM/8wXqvv12KQNg0SHZ
bpAH2UJw84OL/QDOkytflndjB8BjxUQISJ+UsyBLxuRH3O/SY0KwWcn2yqpY
v8sADFUxz+ChMMGlHDsP3zprCVGGJxaQQs20HrmCZ5d3rPiEKV0zZNiCr7HE
R+a3MULINqTtG8DAfwX7T+d4cw3naL6jwKj3zNRH+SewjDRVdH7mDECa1uAX
1ysOl+MJ+Ebz5swCENmYckafRbE0hriAF71uJUeLvdQ12onCKNy5ZDQ1CdCF
iW2IUG0CMTbKHQ16jgLuWX+f1vTn6UXInuN/1m62G465OuFwUZLQ9wanQWSj
IfZ/EYdbC3hZQK20V/4zto3d6jLi1N6wbNDWM83GT0+OmKkulz74MX618UZf
KVyD49YogfmrBV+74vcs56YuAizwwdz+2oF/IvcLrt+riu4aVLvFLeegRmIB
+pSncnEkPrpu8tfqxd/OE3jlJd2rQssZ83Syy0HkhCZBXU4aYK045qRDPgfS
o9FV1xT+PJ0XJzL8Rr1mT1QxBigtr5pPzz86qn2ZZ/BtSe6n2ZoU7M7izG9+
+rQanx2O/R2HXzc3EBYul1U7pEPZd3D8Xj8EsDz5vYRGi2jyKx0O2XuU0blY
Wv2VtzstloH9K0PkEs65rv01XYrI7utK9NvdpH5fY1Cdl2ZQsXhomq2l3gqh
mYFfaf8jEYYUBYj2CwD0E0iT523Yv546kSgvBV7/iP7EFhgA6a9txE4EbF3M
eAmkKJ6y5hOfUt6MgqVfhBfyjQMzdnh9TkzTkmaejVRfAxpW4oTF+Mdr12+L
V2le0FiYUt7lWsSOd+gHurCNYabsjez7lqAybIhqdEQPNlIC/cSeqlW/4q5j
iYayhHoj3tCx1rIKZeuhgaXDEJeAt+C+7ZWkdo8cDvSqFxRFcPP5Rdy36NPN
eywPUh3LhDRWeb4vNwqtUMqDESdtrdIe7FgFxVrVQ1wP70/MsS+qWPY90UzL
AOHV9gPwRPxtvjb7aZLEW0+ZYxQ4UfmVJt/HTqHRlnOIkHGOftGJy9Gvx805
YHZiQrSf+LQBnD3OkBtJYwhUqzQZgP3r15MPPJN3w7G+U7NKNUdpz9YiFFyg
19s7KZ5yzqN2Fwl6UgprEWKah4+TvYbugU/zIS3s7BpyJ7hzqHkl/iek0lD5
rXJne8YKbuTazHhgFeuUquTAomjZt3HyQBZ7h1EjVnG8eHgf05pJ5/SVsP19
QCXDsqOzgmbxobMZYMukgkimtfOCaFbKmUXEhu/7SoNmKd2ajW9hDc2wtY26
kVrZrDX3jxc2T+0R0TbJUql1B33JMdqOYNrCryKyT8VioTVBb3gQ2kV5C19r
Gl83EKpmVCfuThREnUhurmKfClLxK4qLIsX5i+6EaDJ94VF4+qyqcNAkHIUY
rjNZhyP7/2v90tcwcYvRIL+srDt+Y72bay7fJZAHLSZn52da0hNR0TieAfLQ
1tlihs8Ql5UuNlUgmiY7ZrmNQh7qhGZUoNBQlzFrhswIF0hVaiA2gZ7GvaWb
eOuUf+wcX3mmrnJpPpjdoPO0ZGnmgyyHCCTUx5C5NbTAQFIm6guY4rizcWRp
sButR43PRBJhukn3uHjwM/7Di4AT5gGLSEePQ+WAKQi3YTYILgaAF4V5QLBt
sH8rSPYUyk6Udc/9S0DlLKE0OPvXdz53mrG/yxm0/fd/qr6vb7hKqIMEEwpe
vqFQpAmAY0Z1vJfPszzAuFyWT2oih2DjZS7qKu24giHLiDm1hB9zvbxSkFjv
Nz4AGhaeBV5foAubDRVtMZpHYs3svOxZU9IfiTpR1pMGnsdWLfDdnmteX13v
zAiU95CCZMA5FGCiUD9cwZi83OOgPOc6fS2W6JBhpgcs30/mgrRaaEeEkI1O
9j1nKHYJ32QlKnRQPUuQhXfh2EXIcJIiAockWTYTQXK1hoxAeXxfF0+nl9Fd
0EhzKfqu7PvnigOK2wnvCKSZKT8LT9G6/Wy4pN8lcqKwDeybYuAYxG04CL+I
+p4MhnSnlILXmNitJXe4i8aKiQ0p7w5Y8cUNwuS9Eq2HdoBMkPfAnNiN9OpT
+sJQ/BMjPKVZvXvpCOFzyg31Y5JO760UdYjqsVY+t5wzksfYLfYFEkoVr0xI
mHu+zLGNakficMufvOFHtYW7NO+fCwmvxq4YcqoCjSYbYyKNquTW2so5uGrX
j3LixB0DaPS0RyVb/fs4MgayKmZNqueqnbdxC02hosX9WKKfbxS+tIslKhEZ
QZzV+wSZUCLgMPtOySlvhFMOw5Vgj6mFLVD67qPSt3zHP6MXTqv/uLqoZsn1
rt9iMPs4RFVWHRbb6zK5e8qgf/VeNtdPsn87q6gxlzPGKK+qa76FODGbJGMj
teS9TDJk7LQ8tyLWVgCRsojhL6+TfZHy68biln2xItOxYSMMCJQoaeb4CVpG
vBIscmVYDuy6SDmtQKOK6TV2h5Vc+phpayrxOgLZ5/EXuSkmRt58/bTdAfU/
KciZRSBB/qiIqwguFoDnUhdykLcij546G5iWLrMktVpVJUIs9YxlhK7e8ySF
tBCIRRSu3ygCEOOtD+8FzNdkgUZlOQmYNB1qLMzoBqdJ0i8gzBMrufpLhu6k
5V96gQ2TRR3O7sXRhyYE1orYDkMMZep/SEowJnInQiGmnrlUGdbIDRz4N/UO
TBBbZsbsLusUtERXcIMZhE7Ibt41dRLJr+e1Z2BwlS12Q8RnB5FHsgwhk8yx
NCVGAf7mpKjIKRN6FJxY+ChuF1/dOAG2f0z40u1SW13E6VsJAwf4xglFu/4l
2dsv1wVs3Tb5QcZ6TKsxwMf1Sm+WOh+tHVKcZMO0tW+bf5AE4CAVVcOGkVxR
v7DOnsGQe5fz1T2F6UJtC5u9MPJc/i4kEFgy95CWR4zDdmjGa+NtB4JnGAMe
anB+eNPwApY1lR46nG8pG2rLPQJ2teyEixhQRTspt7ficEbdN9Rn58VK7ctY
8BCDaDe8yWF0rLzM5CUmfz7huWpjnqxBkCBjAsayxVdKQsRlsf2nApUZ8+44
D8Ef+zr2IaJyimnh1NEsKPuL4jksYEMUMkJMmYOqOg7KkFg8K+q6BgLh71ZU
nzKJdt29lKrVZFuZtoR1+0Ji19R+3lrBAoPlMx+QAgyWcsbF3Zhln3LlSJvS
uvfVZO6zpZEOL+M2h+NJculPFcGZMWhENqTHV6l8zkAdDO8dRvgJNLiN1xxg
yXSacvX2XUE1aEvmj6ufd2mdRdWlKcBo0wN3RuSfcul/wkStXTFf8j/PZ5nf
Ze0nxJmromhftNXs1rOEaNXfMc64ZkkvWbmGQegp5V/XdWeGY+obq2oTBRv0
nBsDCu1UGg7w9cTXYoj+kPe9yFLXUm7w0HMXtAQJFtxOA7t2YvcTETh2FUAA
MT2pyM7bfsBciH1PgVGphCYJOr5lgpsr0JMo9LzsnPyiOwz+D38750vRZSQb
2p3BDs0EfmjgEOIE1/jd1iNk2zfe6CeJ9usNwvaCFFLwbPcllPIHhG7pry6c
hoURzDZsW9ofky/ytsNonqHw3kenaoUhCOOXxPA9lwhUEw5edr4wnw/diMej
xG6AfoCqlJVBLZZrBbm6RHUq4TKK8SBiUkUT6x5NR/f03xdZtm7VP0UYZbj9
RtFVjmqMyXXgsfaOB/FXLc9UhrGS7/Hj0UN9d8GGzOSYxuzctm0jPPK7j+rP
CoAS0cSOE7qPX7Hns0KHjYAMXB7JjOqECbL9l+F7RFdRmp1MD76aasuFLLZ7
IR7T4BHn/KcElyCEQEvmxtDa3r26CXHhcBDEihHOx+fxrR3cZ8S/8cNbQaY8
dX9VNsWYX1hdMarFD4AEjUIKe9rX0naPARmVSobGnQkliOpAWNwuI2hTUCFi
6/M5g+xnu5bI7g4LHQ2rq0dfvgNJRh8pL27BdM5UGY72H3VO682jS0m/92/T
20bcta0iT2dMLm+osAk5Fmk/jSdM0fNuefe60RrsUU81a/xZLWg3EMzQVURx
kE8u0bWOs1FT+sE0ncxz0GchqENdyBNhw8b3iWGUYZhuvk3tIT7/1x/ut5sU
UIuksCO1HKotWcxLzEkYu0FMwsHfjSko4aOmE+ych406b3koWS6asVJmlyoG
kRN0IsMfkhrQrhvFomXJWvVOAQwZ1Hhz9d5OXarmpRbJOCV2EZIAtxqjjWiC
K4lTpaV7aHUir+FIY8t3ntzb3U518ct5IJVhIiq1cldH7scW8bZC4zVBUGuK
sAdb33zQhi2ax3Zcgoi7VFQutcsvso5sgp5NgBSVM9sofex9SRn09gsA4LF+
09gS8j7bAxED/gLI9A2DhVTFpPEHLK6EB3uU73iOKO4WMW58Tu5ba7c4LeLz
AAis87MdCt7gxpi/gDdLulzABcpi4IzkFvwd0l6VcmR6wRL9QH2gy2M0XUXY
MclQtrKRzgfG1dAbSGVOICncZvbngPqAF3YSfklUcR4LDog80CHFZMoOR5Jp
rcxot2teK4wa/J1KY3ydP4RW59OrPSL+tTTCzHC7edduWHak76hFPmhed6le
1BYbXP76wp5sbBpjtHWstYwPExzXy5zRrYZ1vWeo6ZEhjbxYCotjc053ZDUz
+HsscTuoRyJROPlLX1mkbuynP9LEBP5UvGAB6rj70/5wwJOlK4pbCxhPMxBV
RHTdo5Wjm4NjDV8rEGC/kiOSMO98Oz3zh5qLJyZ92g0Fv9HhWeNHiVatKFBy
dN0lpVknsiFDbL35Sfkgx+tgj7mFbHVCers7inkDxcSaFgi0qzkYJI01zzwh
mMZSI393nUkj0QqHQYTz3rHNxegXPaDdZ4jOxMrfs9PEo/Ekj+Sk42cJtzOJ
htCRHNHc4bv5JOkfxnSzFrNpKAIuLb3ILUaSrG3Sn0A7blNiexRoe1eQvZ+M
qZyp/3tN/7GUezF5lvjDmhu5aSZD8qGXq7HzsRr6bw8dhaH/lQZnOWCIpwaC
L5+MK7HmWMv7ogOUuJpL57q/SBIZttQniFKk/bvfLJ5GKVtqKcMj4uaCQKTo
lgexuMJ47m/RkMhGAmhfs15XS0KkKKjBtOtjvS53P5HuQxHIq218H6VeAqp3
VEJlSlQGRL9jsh9qYpOWUzENekaQrEQyII3kWjqnbHmpp0AuCJY0T9mh3XyH
i3b1pcvpqebR0tBTK/Ab8yJnmxyAF29idWRJTYDA+FWHGZRgm1TKxoG6tZrX
FdrenGWe0MrhD/sZOD/3LxeoTbslCqvK5/zD4cS4X6IgVJUXP7E2YE/d5BnF
FVYNHxj8nUZMo9Pf5jKUuwJbezk/Z6wK0M2snD2y/bA+Ro7ex+kTXKA/Lt7p
Jck2Jhvq3YNxNYR0Wj8fNXy2gnMnI2Wztr6nRQWU88EvtMkwMqh2YZpINjBF
MQ9cootJ5WOiT24tljxG3GiUfniVI7pxlNxPYWsyjc7iFgCO+ZFr+DURSJEN
m17UpGf/upPM6VOv0NlQgI8HQoPjm+cGCl6iIqOWT7lPYzeR8HgP+elRVOQj
mjhBQndZf6XF5Tz6S+xyI9jyhkHQCjhfxtqM6+C7XsOwMttF6DgFLifSe1NK
glZ0KgAEV91uFpZEouXTvPlBlbMOHEDXQcAn1r5/7wQB403IjNv3Ty9R4AkA
oSG14DkhgnNH0dKhewIXgnOSp3WnmRgJKz6JPU/AqVQXwnvkx3tIL0u9bUAo
aEmot2XESGo3vczCks+0nGpparrIIBljq339LN+xViPls6+6iXm5VxvC6UEW
ZcSTuf1rwAp6f0lFcBk2zLzxkZgY/hs3tq5W4i4ufzWIqYFp2lIvO6HYc4ya
GT8h2Po+Hk41QTsRKX3UVWRbakfEvxCnXVs/ZaPHicSdgH6k09Io+vUDRvIC
5s32lqmpEztn1pTec4M2xW2d/tHu5+2m1HkaHhUJtbEDqfSCOcx8anUHLtAt
teCn/KXZKqUmt4XcCzD65LL/aQnba3Xz+tWauZFIZUFsQNnwnYUWo7pYCnJv
VJdTMotao1moewGMRrtUT9dY26yO8EPKekvTrEv2EtOWpJjUnDgosDXEq/sD
IHXS+JNaUefdkn36Aa7Y8tzbL2T3XM/cbQEtHGYg1wVLSIZ6MB35xhDcmNhc
PF3f1Ro2hhtRl8KAanwNIle0DiqYXAlw3ul2GU3SlCM8Lxxf9TeXxcCFIC1m
dlUTX3o4t9eDoVC/Zvdv4v65ifIIAPEMuPp043QmKRGS9KTdRHeQyKj4xRXv
Lq+J7a5I3k9L3EwlL2SeKTUkuJXo5/cS+Ycm1uQum+RDlvNE6zvkjWmhD5lK
krOvKKn7K6FSH0EORFEVWfA1PkcTBa3rV81S7oYhlFFdSoMUYZUCs1AxqcDZ
F48v5Mc9QniQQEhpX9V0aV8ObAmyAPzZG7yR7GgEFuKczScW6gZjEVnRpj3u
B5x3LngwjUykC27cNOxnJgfRVau8t6Q38W4zuYs7gnbM82YbsnDPLux5HTsc
Qy6a26SPpex5aICjQ17J6Aem0a2Adp7LqXcsh+wEP4S0lC+yTqq671C4p3Sv
Sl27S2K/wqGJ7CtHB4f5U/+qFtvFZmyHZsCOaBiybFvbc3RML+01XBWBGUp7
UMRkyfIi8QQOWd/BizkCK4FP90eFnDs8bxNccuuZ06cZuMOk49kMLKSYMfx7
5jOsL83sbYLrXFIiwl+LkAlvgwjWhUA26sEd9A79hjn6VOPvzo0nI6NEslKN
Ryx2GNh3j8zMiJ1lMvIzLLtKT+OAHfrBFAS8ziOB6j/dEJzEk5JWscoOqT4x
6/ePwc4j0JX43Z+G7NoNjCCOe0AlGkpJ3/imFq+5joKIZq3n/mhO0BOHJubQ
JOKiDwu1j6XMTWCC/XtAkPsmDp7GaTlwVzdnKvHF2XEXNhXbKJva4tB57Wdn
7Zp0YMaE/f2Bw+2+fYTTMQFz9DsbY8RNf7xjeiLmiQAyCOt05UnqdVeEwQkh
NJE8cmIUAdsiuM2OYE620BxF0ZOQDZo8lt+ypvjTLzclvKt4kUGtANep0Bry
fIiStOLGouuNaiwDJFx2q7dHRHQS6zN/dRAh6S1eOeZIHlFqDAR7/NVoG+lp
mpb3AFr2Q3HEM0aqge4d25pJP+izDPtWXfCFATmMRtH3bbXvdO9ggxMKASuG
eKbuTYT77Cvi1bBDDFw/o9opqYsCdwi4DGBGmc3gTGW4Wh0/bDKjiiM8OreL
FRN+Y488jGaggk9rYEE0tkx93m8APSODprkBkUm2sTgv4SGbffGbPNvOFCHD
LmAmkKBEV5MvvxjoEWvBVysOFexq1MZEsGStE0x6z2T0WRondVW7TcT5DMUz
vAgsVTVkRwE+45Y/kxBaYlQsjEw+ioxcTCMnAhrUwAV28ubV9AmobC3F4q56
nXczZP6yMGCrS75tX69+YHCBMMPIewB2R2OKbdBeFDSD9/0vqf61eb2gqgBo
B2AGXSZOkPHlSIhM8Nf7m6D4VdOFCYctBkZjirE/+U/6r1pzAA3GNlAWTHuc
+jGNUZ/WBpv8Skzx71oiZ0Iw1aSNsBxJfpS/l9cTFhkeTBE4WrVp+k36MhD/
1rJFtCwU/cpurtNR2FLxOlIOEb/gFWp9DvsSpAfaIMPhL+Ck81YmzmIAqtq5
GvxF5OFQyxMEPETJ5ii6nTIJkxQ+UsBwIWEO2jbB4EgQlSr1rAToR/K/GB5M
meF4mC/Fx/5yjCQKip2DLD94FgQDq54u/wbfXseqMlmrw8UfhtYzzL6rqP9d
Alzd1n8U/StgzMCAEC1af9dNkWXyv/CrK5OzcjLFcVG0EGh5XV2RgpYRLF96
4s8M4Peyt4oFubpkSXqxh3Vi7Dxw/XYl0CYIWlLb8sGz4hXxHi8GpO3fYalH
AGIGRfIZr8VzD1i7JojLan0PmMeTslgMyoFD7MlNjhIMgEl/e35hUT4fB/gu
K2Zr0JRmCNRiHxUgWpVCYJIJMbHDXiyjsiOCzfe6+UKMrmHcrt2ftAHqenzV
drusc8AhPBJrK7QRl7Zfn+kgw29lf2QNFQEfEzyZrUm+rSNVD+Etyppl8jxt
6kops6uvNyBs+jDOGtrEduqsp+Ghe3bj4Kf/SVXef90OJS+F6tOmcQSYy6Mp
b/PQg3EQfJI5VPL/uNXFt68QwBe0prPJWJe0HdIhOI9cpu68k5BAFwFCz2Ca
JfYMKuUbDJksYzaw0e4uGdFPPHlAJsbFPw1qqctwYF57ejl0kzOm9+1lYmOk
Nw34dt0RBjlkHaabAQwgWHhj69k6gPUyjp/TLYvurT7HtrGqBRFPvWLTBxRf
WM1fkMoyrCH0l1g9LqH0Dz/j3aM+R23qfX1VTqpHLn3BAF4hz8jn91AQgZgV
YJQY3FDGGwP2W/5nlkFUGbba0k+BG+EnwOUHpSnKgQaC+BfBXLLzns2sL0aR
CmPK4AGgEKOaSrHvEKNlq1rv75jOG0TPyldFX5ctkStAy2R79f3y0197zcsu
rei59kfEIOxyh3qq1qYKIRfuA+ylEVFxZTU+5xGmunuBZTQSSZ2O6L9I2K31
QLblUDx5ysfU+1RFAJvZ4l0bynaxigWq0EbKNVRw2IrjEhbPb1h34TxEoAWw
VuOsPoBfhgD4Pv1myxnYnLgqV/pY/rlbDj/tdEikPfyh+/+pPeHpiYLAxKcW
DiH7vhVZzx5/ww6T13HiJIC9ClqZgQS3dusoLgIS5ZGLYryhBIJX9WDUG3+c
2pTrxfnxM7qIbibL9Hi4LcwSo8K8lbl3oDf7ol11QF7aUyFKGDiScv4hk4OM
GeAhSJQLY1cuSMmrIrt+qvl7qv6POjgkMKS9iv6se/z70HZiFvXk8o6Rlv+U
QiSGUflmxDvufhz9mwo6yvL/cXFxfpaKBm+MtXohSedMwwppDPd3o0+DwwUG
Pok2dutEM07Yg+4KJn4NP/6cP5mRire04Du86GlEVbwOtW74d4MYGcWynoi9
GH4axZOPQUAB9Oy7DOz0bYQk3WC4KcEk2SxoE0g0mKsDt3N/1jgUAzSCuHws
Ujz0dPUSyBW330tfQ7dndYazZ1ho+hxODPiDyBOoeTZ4ISGiPLcmanZtaZ8h
LyP81NAMSy28Lq8W5VTe4F0tfULrM9aIgUkRP5l4MBlHd2raC2At4+zVCuA7
Lz162QVIZ3Si9rsJpNR+uQlqj+VTkviHamEIsCSD79f0gMsheffyFTh6oicT
BEO03eFxBp7Dk7yXLHguTJjMVhkyR5Yo3mtNl+lDeiO5iQ6DxoeGiQMXb/vT
+TH6+GWzsvyU5RZtcMvhOaziHpYyyQV1ZUkY1CD2DmJZ1DF19Pu081VWLllB
T8OOGx93buPO4wdw+heRif7zFN5vp95LNRtrJVwb944c+vvXYkVgdf47IAnG
fMmqmHxnJhd5um7qv/5vZRu7JvpGzuUIQF/vkCu+U0UQKjVSExoZ02zQGQ3/
9v9P5tJz5gZz5TWMwMjXz3ybzOyckjS5PDf6tqOsd+kWhJi0dAQHsW7WR+62
bRqw+iXK8MphX9PO6WR/90qtUmPp6A5GEYQQCyWZnvRczp/S0ADbVb/WBT4h
g8ALKlU0fqKPmvcMHdjpaFTurAfiiyPWV3lSpUZithatlBOFBkXWaefprW0K
lq8ipDw7pdo/Ohv/B1pZIebXoIRCoc8S4q5qnGxvA4bZeyW9QbKpMY4ZIejp
ZF/eCpLMmfejXiweEtZMGW+oTkwnDCXvwwPB0MWvOdluU0qhvhmPbaTxv0hs
53tDyK0Gg1P59mJJ/nggl/oDsQOTRPpKjr86rqijduTv4wB+ITwqUQCQ/fpZ
6VJRhz4ShPFZ5gNYlqjVyMO3GJBx0A0Gr5MOXhm4WmMjQ24Pa8x9wQvAI6o0
I6APW9dk96GGnM2biGsFiPssXg00AtTsaraPAuTpLe2Xvb8HQkFjgV8LafCm
FQsA6gDbuE/T7DACa8o3COckfJy0YldxLbr/RZVopV+Hxksvhjq5ZBv87q7B
xNNZaxGjLb3zyAZqiTbKFyk+NIRVcZwn0GI/BXEgpFkJ4m27+ritJzpxi8l6
ECqTySvTm1TSCI+u+ngymq9lp2YS+Hd8IIxjNSAM2QNw6yqTQ1miU+dnpCFv
Eoq4jPP5jOFaBC4klO0LcKC9AVvpiqI7L/EumX3PPqR5q1O941lY8bxl4sT+
dVibUOgUXrnckEwEnapE5Vi4BoLJtlaHNMCdPhLvRzAIOdbSYlUA0xLaow4A
Ns4Zd7zhHJFoATr7YpPRujcpo8VXsfUa5gFJC9S+srUM419xstc2yJtQtWZU
/Vw7V9KSPdDL7vW3F+qNWXQoPNS8/KbWeuayKWttABOGvdcFAiFi66Y3m+QF
l1mbH/gpIJlQy91VyCki+4jWx6RdcdFfWLVOatnwPih/t5lo3qpDNpzX/d6A
+T9sJRpINMh/BKO+kfOCyzqiqAWXWD/c1wA3+4ERdVOTmsk3aPAIRMjm355V
MzFR8Bn9ogFJuhttTyw23D9aYS+ZFz+m5l7+5Hhl09ir+B5s3TedFyvvDwA+
b7uskEXExBlnqOo+qvQ0EhjugnkN8fQyT4dFGW8NKs8sAda6f3bqmdbojYNJ
w4H1D84r0xJMYLEiBooDQidnz3gU1RDWULbBqwkzasZpos5DglMuhOrR9Fqd
23ZUOSrI/LNonyGPz7ySQvYBkLWQ2Ygtf8KdBKx+2Zp3cUvn+fhBkTtA/Iwo
C7xVqifZ6YUSFFIqNKvw7TmzKB30zLfwRAhN2m1Ef1lunBBsSUPPDAy1vmqh
xTL8L7plDa1+NaQyIgNDH3VWqpOm7kAl8UzVSJCs0A/9KVtUC7Rz2dXxvGEm
gbXYAETszpmNwIyGfv4EzKeIrfjgCkPCVkLYYyeqFw1YjdV3BqTZ6SoMe4CE
9COuNzOd44OeL8geoU0Yg7Lr94kS6lCnwKPlQ9gOz48IFECehoNFORwjUO4b
Jh2d1tqbmzNk8hMoIzEdjjAQgDH2JE3TnD2JzN+LKQqa+5uqci/M0x0kkObk
o+Me+lwxW9F0jjqLuU9karPU5WQ4P0F4iQlsPPyjAMLic/prL1MWI+riMKxr
YWG/qmiCxnMH+42wp4goa3bAxVEeMrWXuPUQVpelD2Lqq4IoOIKVevx+AoDp
86bjEh31sIE6FBwYdMdK34CI3OsWVbgQVbbhdNaelX3iZ7RTeWOZK71Ldidc
BFvbSu9YD51gHuBDAEiF+9Z0pzk1znnszT/AKGycyBIKsxZwrH/26C6wDx4V
2iVXLvib3PbNL5axBYp6FKNk2uVvuDcXJCHinaf0hSZpZlsUpn/XXFeBmxCN
xRqO4yCd5fx+gRZdj3QIVkFK4lIyu+3hmKVqLriMM1Gqa+9KL+UqL8dwVdwl
x+ks7rOCoz55aOQ/HqjkzUjLPLCw38Fe+C9iZa5ghsaUydDkUnRMwvdKIsnQ
yDRrxAGPrzdNJC8XGAB39356cAo2cXqHDWJkWc/P8Z1xTqIxU7eWGN1+YYl6
OUSq3ct5ZDGelUYeUq+oKQiN/e0uVGvIeB4aiaG4JdsCORQb/pYF+0eO1nky
eHlnEsu9x/vB+DDCwOTG+y01k8FpiACmyOcOqBIbyzEXoB2C+yPEWzeKLyyY
ZbXbYl1kI2n45Ry5XLgrTZRYQXo6DCqQnytGJGMBOez6yckrUxWDe5RCZzZV
G11mlo330hfGxV8LSPpALvYBQcLXQxLAbMys7wgYmb1HQCc252ZtPwMX/nNf
rb9V+mvvzcYelKWv28B7HRZVv7yRA6XSuFy+2lzscVi2oynZHZiSKYDygVIb
KG23bE9ivlhXA1P3+g0oVhiZaPYzTQ5HtQ6fZAX3KO4an/ZfQSeqTcysY5vy
SwqFASbRqRZUqnkNsaTvKyRiFW6vmMwg2vLwpTYiBAVgqPtoQtOtqAc5526F
ynYpJIAtfvTM3UM2FD3hEFHLddddAsm1gMD2Sx58jdqQ7kycLyApPW/Ai79T
vD8oihITpmCaw5KBBZ8jCXQ1Tww2pf5082aTMwOkyBpVZ7+rvEiHtT107Rbf
dA5inttWkSW8kOUsoLHSURH9J9iZj+iZ11AzTxYCUEmVAZO/eHC31K4rZRpz
GYdfvej95ZbUhe07TYTluk2iiimY+Jz5OVk8KmZL/FjTS3Kjsu8v89gDzL1d
9Rh7Kn15tSJ2VBS8U1TaW9xd7ze/o5uPOgyePuTSgGsKyvTRMUsVA1Hjq1cP
b0HLwOGSo3tW5vkQk8f/dDhiEdze1OnzJIH+YSdkYBTLfAmEDCFAqaSzhCXs
OqhbfgXvxuVrwXrjigOGbdsWENKEP7TZNLLoG93cef7IrKhSL/RBJQ7uibp8
4advDicAyOGtyaD4trQqzxH0B1YTV4gnZF8qiz3UOq42Pwp7qRABePuWdkd8
gQhRPhoYaflElpbbq7c0TffcMDCEbs9QjFmGN8cGJ/N3cB71DQdbSECGbVe/
cuw0s3WsZyqjhlQSwyfmzuJbq5B9KojGyI446wC2WLwGHMx2WMiJI0SZ48HX
WkaaSLupm4dHcdoqqX1IHdwaLB+EjIS21kRc6fcVC9ig25DYUWjY9wL/bz9T
kjIg3ekn7oAuH4jhE6DayUofYFxQagafmUQxKldjaRzPeBqTWu0J6bsc3rq4
bwGdnQLh/p3WZIOm6sif0hfbwZLgc5jgv+zoim3a015C0UIhpQeRhbAQdMjX
xJLCPWVNZVtsFRXB86KnQCqj0lobnQXzGrUT3zV7zwIrE1FyOsnTZg9T9+NV
0z49hBgp17kcPnTSfgEpa1xsG+PxEC8o9mdI0Zcw0QwhxzT32sQwXgkaCRdD
P5MUeq/HZ0tOaatAvZCf/gTRJe0LrkySUAbQYG8dprduRqHnqOraxCaiV8JM
jGN8+KDN/OQauR737c2NYKdWpK9HaqyzXAva5nmxYsqUGxab59PX7Wa70KSN
gfxuOTcG54Fr9d1oPFBjt6F2wkUzNWmpNfZC4NYyqc/wQ207yWF60LL4ExQn
3PFiisQv8g7OCK/XP52T4dsPFBiTvUb3ar3RkAaxnq8kIMOArUQJBM1FAg+4
Hxve2XeXZGEEqDDlH8V6JXlcBPnBDS0IC8j1IxWLlCSzUQ5zWZBJgNWfuLq8
sNHRAGdvXKlGWebftTaIa/NKkEjgUiqQUZ8J4zaslU+K9fiUUQc3OJFKBbj2
EQ8skcZPqTJHPxtFR+0c+z3UiImC69a3CVlR95pS08otjF1HLtgGej1T5VmW
fQQrYhbibKjgA8liTzUMJewyRlLG87raxEFNQ7ct9p734kjqvfqfdRG7I5ct
wKOJ2PQ9wL4vZ9Yui7R4b313ESdmsdfQgeaY3PtubADf/A2i3feEQeZazYF4
ggaWGjFg0HXka5TMMBNA0tURb66zD/tGYN0428jiY3t3YwVWqXEL8rA5oQ66
Ndh0hvBLwySnlKta4paKfzCHRZz04sdlF7KgDqQuAIaYM9x3MV+V8LuEama2
LpVTkZ/QuZutKqVBw2axIPpFGBpQeJsUbQfnWUKOOG2WfbJJMLmFSySgsUJt
2GhZ9LB+yTp54j2cUvFL6nrkXCssXe2SytHR+/SbWVOtEl/P1Oe/YYCKssIm
vQjrjA78P+z2b2IRWZlZEycnYNd/yeZLYrKR764oW0gHqncMv5uf/pWcI5yC
ElNF9ArXkPs0uE6USpsBkyaDg5CPiguDNqoXHFljfPxSNLjfUmL5cNb65hvm
SFCbPZLrV73jhyNqxmnRqaUu0ef3L0J2uLV/if3qIKMJFYw5AbxzX3fkQLht
Pg34H3k3hiuQtHKfFRqMUYcAbxRcUVW7kDTcx1g+9RGZ1aNPVSEQGU4+T95m
sidP2rU1oLWZLhTPX3FMxlQ3t1wkVLM56XQNd4gKlhb2E04r9KJStJqSJBZo
hB/BbdFHbj1mS+wwMSuM/b5FImkJLbLkXIOA9X7ib01wRcRwfCywZZOn6Qif
S7Wy2Ff2OzCj4urVpSjFgpEHrAISPJnNbHe2IKkRmfrDFGsernl5ZSQYg7PO
x9I4Sh8EWX/Rc1UOaatyfrKKTAC7mmhsJgqb66yobnN3oNHAszwIkh8GsY+u
eGjCkf/vHSDbwIMGbOFn+AQMvT4DbssHwcvKNoT2W6G2tdzsOUc+BtNTjL9s
Q9dK3xxSWItHjeWVaIF8iIGwiZ8oJkd8fQnEaBB1zFwULHRvfF4gMTIlzspr
W7iFEba12Q57eE7T6EIKudr8IKjhue7wFZZqPnJJTglwNlAb188jRwgejRQu
kffqbhfjKtj3iyhAGq5rqrvyy9OZM29J0AVPGFUFlVrDSRuRbwjflaRI7Ixd
yuTtTV4MEVeGi9ZWxZ1hZnvNBWbcE3Ueo8e4ndDoYzNN77on45eNqnTrUvTa
RgCsWckUFdPcnWZ1r3/PV6cwhAUDV0EhcrMT8aXlbReJ4w06W0OzUtU6NbEL
9j9OtpxLgG4c91NN3I5pKY3dsaY9Vrj/eXF0A5IF5nRac+iyCkqmpz2zRldr
RNuEmm2ju0/syo4giY2z8a8KChO7S2hT00y2sc4vcxIFpZthJgYH6kTb6Rk7
Z/IIvCn1cxN4mQ+50oOTOl0/o0mD83CgACMVBVekfbKF4T8Tb/Y4TByR5upW
UPBF8896yxOOaB4cHx62E5bmCXHBoqw7kwvANh474Gyq77I6+GlwRULUAL5w
wL312hzy0X3wCd8lAUQLzITsmJlkaggxDcQKm8xsD37iGqivL6o5i91Ik31l
PJzgRdWxbSv/BKSLQjQ1sk78R6R02NpliQmAsQJbnZQVFF6H+Fo1HmiAyOoW
N5FIrmDBy9k3xO35LdYBSaQsxZTdhdfmxw+RtKWkKXrJksEyaO5mnxnv3oR1
Sll3UKswohP4AXR/c78qQEwrcqY72FiLQKLEyRMfGA3yE83Kn2RY63Mj9DIN
wVXsHo6Ezl3/Y3pKE5IJdRULxhFDUwIl5WqUB7mgBk5ooBpqbgQ59/o69PX+
HSuTWtk/8QUpyqTKXpgmgsbxFCNLoHkFBRlnrg4q7ncHNvAyTB6MauRUG/TX
WCdoxtIF8H51hiJnx4SRjI9fNPULyeoWDyF9GcAtaG0LPtyIS84+jn2VvyS7
hpPwUlZ3X6KT7PE+rAfnScDxfGAm/t399xRLnrk5IOMr5uN2TsZmYkgebsog
Ycxk8Z0C6h5M+4LtIqoll6X+3Hc1S9s5WbdMTmxfkYSScVUZ8xoMOZMrTGVl
er6J+LPDt6xQ+SXmxu7wK/pRoGzrvKkKTrYX1+o5cF1nVr0baVH0h8+zIT3x
qpkHzt6FYBeIRTFTv9nyvAt//U9/1Hwv3LeK4SNlIVqSF4hJoJDzKPRXLBTh
7gyZw5uei3M3NQV53Kkh5fWuz5GPQMGFuE9O0DPOAmIK1GHlYh1LDV0b0Fql
RNkL9Qa5bfaNJ0SGFY8ycVo95yG1lE/nW+Y/Q2R97FQ2x0xWzfqpcY0vwzTZ
LeyPhfjPHHjEZLAxPbebFABnMpHHnipp2NhsWBZKwBzbyDonY2Aa8ucemiMX
aYGbGY+P13NE3TuiJgVlpRSIiloPbgoeP2sZq0FmYYaGccmf2Rb0JeCgnWyU
nuJD2Xm1A4p4M+G41zQbugJ0FCbi1LvaB2WOvYahIvXzsviMesF5knWQrspV
KNb5KxMKUpxZT0aVw8B4Wjp7i5+EdoiOY4BKPphePowsSRi2+6l3mqBo7gJ6
wsPxWdbBR4FLDBBBR3uRfV1MV+cj2sZGeucIdDd5WNKzuImGdjldyGASQIjG
4P2Qh0IO3uzmu20TV+YjJofT5sS4c2+Wf6P4AXsIxIB6UilwbFM/RCjuzb0K
BHGErq6iGGDhhIM1fcmDQjt/rsM38eNnBxVTcxn+kC6/2Oe9t+voX+7RodtJ
zcMxNXh5s3AaRnIUO8d2cBA00Sf90A3xXNJ3YAdsubKKu7EnIfFHhYKRC9ps
WpfB8zmSVxcX3KeO21WFtciV/v3cvYcDPYSzjtqPEfpTP1N8wC9VsF3bA3kk
uIGacQnTxeZ7OOsgrHU2M+HU2T5o0rztHaahiUx6VPoOnxN4SY/0Vb0C9MYR
V3Pq8xBgfUbgra8qaWE+vyf+GdDsdrcnqtSrNOb4itG3d1I5U8epdhvC+grU
csInLRzN2E7NEa680MfWJ5dq5n95Ttxc+s1enh+wYmuVHVev/SWSIaCeKNjL
HUMJvnwQlF0+4iG1YpZDlbbsmdPi/V8xgSPWu7Ap5m2eG6ayLmpprphBEr+7
QEgUDuB3MEsJnU3OlyrWRxM6ITw2F0nXng3ZcrpfoqfFpB8RUl6fKlB62wgb
VO1DpIkdUeBVc6AZnW46Xs42bdnnGYH5SNnI6ebVj6jMVb0VWH3Flq17rHoK
EqrDiouXXKjTvl1Lo6xZuSyUNVHT0Fzjtec363I3qE5YsOnxAySNIFIt7ZSg
mc+ViLZJdTgBgWDe39+WRUvvMjVjehQ/dWKxz7DA3pZPRTK0CwQ7+etV6LIZ
mbaT1p+5kul+mWeCycc/O9BV5CDKz+IpcAp8n/LwIGe1YMqGqEQSmXwxG8go
3cWadoMQJtw0sIyRofelMtd7l/7smz+o88NxwNWxSOBruoL6Kf9UGMKPZXDv
f/VbTMB97hnTTU2w6w1zlKAr/64geenquSUBhuleaPhmRFlymMG+q0yizbYB
JRz3oK/gEKyrHSvm/h9EZGZqOjMVXHxdYeFbfAf8g9TO3VpgBqqBqh2bmW2f
o/RidWmi7fWfUb6E2XM2TnHg686IM0TA0nhC4GcminfEp9toINEGQnR9mYqU
1xXv5wyfJP1lQ7/yknvUf4dEsKhx8Ctb5oJ1Z5sLSV5rKabP7jk9jr5ItDCM
kr+aAkHq8D7rE7cZbiTQeeLLqX3g5rxzR3SzqGyqCFetctXHX5deEGGhb7RU
UQQXXuXz7MYqVE+KHinJEVsRuqoqYF6N1UAKqnrX7xzR/e0mud6c6PlFhyrZ
of/NK+Yu/rqtEUgHwVojJWPKgXmuyy5bQc63L3WCM3olJgwNQbz06reGXFWO
wdlB9g8tFz74py5S8HFNxdz0m83M/qu8kd5C4qJWZGC/ESukutiotim+wyGl
SdupVtMjsXe8hfQLz80FURlF9+ye3cUz/b7J3vaoUq2lU4qTHvKLFy34q1Sf
+Jv156o4GOvJN8cA07aSp/wtQbcPZ7YidE7IPoxvlj7LKct4dJLY2eEjQk+t
DCBI00k5zwORT+RbS16CgX/duu5C9FJhYQ3eJFU3Rza7+RilwNduoKc3XxYK
gLVLHH6Fc97JJH4HotgRYs77sqO22r5OAnuL4OXvqQe5+Vy80QQXTZDdu2Cs
BKHyd6tThtJdKjEcwG6wbKKTRGFRAdAP283R940AXPfVdMiBk8eBxh9K11qo
GLuhABOBybR7ROtppd7gRmEZK9yQf4yvc9MAtnzq6Upk8rDxvNF2ZY2yp8gf
JgEDZtpdhm2fabPQJKZX/Ej6ourb9dX7U/vvrwv/RvMmT+kqt3gJ6thBERzL
trZ5uQPjwuKVvYkwT6eG+Ud+4l2ouzWrIOHeaKCQNpcVrYYaqRoCZdkrL18e
hzQnEO6rgGPw8wq6Bf+k6+yebjxt+gGEkYSqBheqP6bOXd+lK0L5TVLPulKJ
dYroFkQ9NQaaZUXRBkb/pu01+pQw/ryv/XWXG9aZrQ8le1kKWJbKWtN6PWe7
CeNB5VlDCSDPpO+wkOuk3miVD1/jdUmMMuGQgj5QZOZO9CMxM5RgNzBfeiiv
jWC/+tyhz2NHgw7QzV/ySnxvIOA2sJrVF4/vDOR7abZ1+pjAH8vaH+vPdjyp
LX8kBV7oK/UW3NNCDztFOugfMFppCBw+aouFQdKEY4hEU0KO7U4j6fYHbUwt
KOSLCWp45yDlpeH0HM48u8Z6g4VLgjwfX4C+kWxaBNpUla7iFzE+cDTC7UAG
q9h1kOJezKyMgsl0RaonNdnlSLPYIhcSI8gxy492llI2hpC23WR0153DWmNJ
OPqVx2MMCugUXoxs9zOoR94QlOL+7eH8tfewp/TsgU/RxSIRXKGJMxPFoyWn
wrIGic+d0l0PXtD4svejXrprRMsVFGa5bg33IDFIfUj2x1NidhUgUUFBLUCI
QOUnGULwBnRTKFZfYvqVckp46zcbF2zNrU3KO7NCr1a4/OmLHfjv0kjuBkpd
s4JqwSSdLOjAn84yZItbbAK3WGtDLGKyrbH6/PccZh++7Hu62LVYVOV/0ehW
TjSkQpXPtdKWa+IeevMj5I/GE0o1/9GlTNwSAFYJah1HEUbkGO9McyLu7bNL
E7AjqTnKZrtn0DD9z3urKrqwuwQPaxMuu9BTDxRW+hEM/vacMQjfbvbk1MLj
OcG+HxTq7R/VUSFedJh7wk4xaBPN2ir0oWOdyQ8XVpccFBG2HIr0jDUHmFC9
MjD72TtUrrl/ClU9xbJnDk/rczIAiO/T13OjxnIIyx4uMDWG4d0Sp0/jF4Ci
KlttKfr0bigtO344cFOa9aEL7FdpHo0eGC8vekRc5u61wP6dVA+WbcCZBnP9
g2Ctl3dSBLk7TSc2kpZlQMXZAc9EbAmJPssUoPB6aUTp0CHhRpQJhMHixPTX
bkuVdjgxdyJseYqIhGQdC74gCJM8In8gWYMKKVAptCIbgiDxUwES/7hinjl3
Z3ALQUb9ExGksHPEPWnTtqSeIHMKQ+8kZCiy5blPPHQ22U89exsQWvpnDpkg
aa5YH/vYeYR6oxIjYocIQZ2vIzPTUjbot3cgSX03aneLWNaKIluURaL6muYH
hWuPqsleAJE5Ou32upQlFMwxNrJSWq6wZDKhwCOCXlU8YGydJwGS5c7cAyLG
MlqCkThNBDyeh33Ao7qiYmq6mBU/0in96QQNcijwkBXPJaaMRaojdS+UeLYq
wYpb5c2lVRQKO9PEPNERYNzJxs8VSnB1PUVF44E7l/xvx+Jf3BmETuKd1bKf
rXkrYDKkkGMYrgISUdElaHLZeS8numvWNiOGcnsBZrFVRtxI5xYx+n7mYXwD
HNlLYi2pnCifDuR+O9ho/43Iroq2mrhqQSIaiFyAh4bnOjnT9d0D1IOM6kCv
BNPIRHCE5d/aWef1LJq1CzS6zOPNF7dWWtbkHFibm+OtGeyHK6okYqKvucsS
oFWa8fC1KjahxgO6MQ1q7bVksOfllms2VZpXDab+Tni0UxJ7L+NHR9AdSsvg
lR9lYB0QIFmr2WxKzCz7J1fJUn5qxaEfhCnz4BNW2V032qgpd9b7xpQJPv5M
U/HyenEHs5vk37oKBd40/c6oHXu+WoQGqBpF1T6XLpmLkMlDb0Z3im9cjX52
92a6oEq3R7YuToG1soAMNObfYZQjan8y23CQpRfmK4RluNQKU0Mrsjof4eMD
ISzEwX/SSegNHb7ZmKQ0Jif/yE0mrQM7NLyBk9nvmEIowDyo0O4ZjfWjguaZ
6M12v/5EUuvdoEqVj+ISqNGsgBFxNKi5GERE+WTOTJTfyZ3kbZTKHNWNVVXN
kW0E3X201LyRzcddY0xgHQ4UzdB7pclEDcxNQV93o2VeGyP2t4j5Y7fFEavj
2SZNcHI5GqyYRb+3hqkISApg8i4chedGbTnTDluLmkh+L1yfOBfbTxm6A/xX
7IiQsSSXSNDErZ3N6iSLmTSSNj1bepUsaG4+thDSJ/ODlmQFVbJE0YIbVIFh
41/RWNQrWq/1gRRWqrAsqIEiFbGvJ3nvsTxcQMlpfqSAdAc6hwD+YyishXgq
wexHmQqxTNHEj46ksu1dtpM56h0w3ZXVvbnR+3ikEpwPyRumX4afsR15P8g+
y9gkoBnMMb7HBGYr0y2b9u+D5jXwzuJ1oUws0GnTmD9LaV8Y0DU/p20sb8fV
gtrl/CPZLqQaYsplyKSK9LI1vay4fNuew12hJRmmz1bQIqvBD3S/pkjZBjUV
PX7cZzi6zZftCB9q6zU2wwQZx3HzojToys3AK7HtTZ68Yj8afJvzGTO/UKz4
u8/bWhdhUvfqnEMvj0AR87dMPd5eS+WJlq+kE5q4eAKR40vGHP8VRcSm9iy/
s8ZQOl2lyZohwAjIUK9aTYHfcIrTroVwVnC74kFv5+Q/EmFsBPXNAPsTylpK
monmbsSmUwUg419gGsduRs6LkzBHRLL9Q43HrUsQRUXwH5HtegyIz/wHTH8V
Kou/krirHHekUokRlRXZV4+oLSy5h4ZfuwImOZ1DPdA4/IDm8gJ2JBIy75nx
XQu8FqIFa9b/Sa9IArrHlBxMogpCAyv5+asgf8gCDJNkcBfRhCtgtESBJa06
ozPuAYJYC2jRjUhSw7XIuhTVrgLDb83dKOllny4VMLEIvpkC09Zs+qzLiolQ
FQTKrkQDeJxguSNnBDJKUtdux9f01Nn5aYX4hqVpn2N1+1W5/5spBICwz6uY
R2aZ17yOSjTrJGBic1GPFCglNP4gdh5t1tk+QTe2JZYps/3qe/LIuCyqqBTf
batd7jBr7YRXZYPpEHgC0NXDP8SHTgRnP1LCWEZ5BSsYHnrjF+DnCiEX2yPs
8NEckVkJQPBDjnBr8bo6n/epp1JdNa7UDf4HqVmOtYEM7xLGB2dujeyDUY0K
iSk/XtyTaNtMHruyjmWYJRV0DUAwk/b1+3yew+BRSS3f6z+NxGn824MlA1cA
fJWefXoyujaMdjG5hQe0jpHEeTY+ecrWW6cDvoTAngKUeSCrdfQQXrBOEsw8
eqYBNw551KMl2WC12337+UQyzy5UEDvETcN9dDGTnJwubZBvvoB8E3676+dx
tOsUYL7jWGLv84vyumHtsu81WBGYTzP+WQdUZfnGA0wx909BQ0rusfXl+gD2
ORbvUzIMDly2+84479tOmDNudz4lyJfhVPAQVK8p7fQ9pXULKkxADsB0xwPb
srfiu/V4JwLtaHI49WLYl+PCkTk06bWPOjEMRH4nnUxvEKj8GYMB6W9fWLpx
8ZmI7+1tKokUrvD0ux46ONBZxmKgyJTQaaSgw4JwTS5Lf5fNf2+T9O3CQqMB
8D+YxltgpWyDmXtrn3+xzTKBR1geNxSeT0NT1JIuQc4dyd0CZQYK8bYLCWEz
Hvii54aWgjuf51WLk+CvufmT3XZBp0xVdYMPBA6DBQlPbhRQjS3RO9l8v5Kb
GPlnhM57CtZWN9iYVwwnYeUu861hegeV3aoevKT4VfEaUuOlVFDzCPJIHt3x
GvBa8t36BaxpNZxdX7T6hbBesJFEogcgK+ucjFvn+qwjdSAB7D5ldl7x1yhz
z1q8PkiMD9bRFCHPho0MfW6qJq/Gc+20QXFFtQ1X3iWcDfrl/L+H0E0iixhS
lKgHbfwFhf+9cpWXieZLCmXinBO+gYwT+wlHYNNiwyOnclkVNsXjP+eNvgMD
Rfk7wYvqPsSWf6H2+7OBgio5SIOXDQh2z8qLjnLM9OGJVNom5PQiVjXhBbvG
UO6EoVyDCVFHQch9F2WeSfDolqiibFXYtp5nyswr9QOIFZKyzEE5shLFvypj
mBXDOxRlBI6FePapk304NEOlWD8KEYBsM6ztX/pArZdTnSHi2rZKmsFuoH4g
ocQX0dI7iZj/4bWJyjuRSdOe0kX1Hhk/grx4ztvh+oVZjPPU9y0Wv6jcFVIT
z7FFhAaPm7RNvtL76Y3KOVHmf7g+Q1xp7mS7X5pDjqkA41WI+cQ0D0S+mGRR
lfr3HA2BrUUnCEMjIMCTfq8+gtruuKQFNoeebn+kALnGav4tbsjyYcbaa0w/
hq+NqlkSwETEj/Umf/lVo7vMQ5YQqRZ0jYIPA/IslTUHWW0Lf/46HSmfR+CI
UX4dMxhWk3yyu98PmfvQJqMLHZ+N2/dw0LrA6HAgtJCZhStp9y+iMcGcsiQc
O0fKmm5Z4jLxlYW20q7jo3RLrQB2SPN0eePFEItRgriD01hY4S/wmv22MplF
LNDcCTmgvRywG9OmjMe1fuhJ38GBwtk9DdQRUKbyJqWBbF/5XAhxMKCV63nZ
GoFQ7NPqWAoYiF7VTW0Z+iPMaQCPk6Hq8gvwJtng8TJSfk8kRW3EClEykEgi
ElvfVahI1Ccez+7FkTKfUOPDYyny55RhulTMA5dxkmtaQX/Eiqx6WBWgnE4m
2NUtERlXvvwCO2B8VuzYaqpQWtlH5WdN5WyVpP956EikY4iuA0CL5N3OO2nj
tC1idBEhQUHbgV5/50LfBMkE/taJSZvvf3y20tJ8GEt2czKkWJLrSKF9JxN+
MRfQttAnJjzdwlhnzPwtxAlOFDCjp5kj+rVPefGv7nxUghieHPXU//0SSX5W
iMRfz4gXZflY2aXpBioXwX1jDx0/miRHonuAGxUGCyWOPwvK0eMlrZpzP7NN
O7GPFkkrUe4dzVbe2myNUlVoyG3W1xKLv7GqdieKw+VueSyNtYwdlIHclrbR
42VQzrWUqCZFHBUVbWFiP01ZKIpEpZgkv2jn4fqM8NI/FaNhfn0mExTAlsiP
Yd9cfNipk8uiTxfLjp0jzZqKU9x0E97rQ18HSb9O6oHpIR75uG61DRh4Yxll
gJonCvJ3cEUwKoGLLRy1uGQgCpUoNfx7phaHkwNIm1W41n9Ul/mDGpnmZgse
m1HaI2F64mOM5/Msa0H60nlF1E5m/KPxYIzZlCx3rb76k9Xx20j4+DCXVyf6
1VDNCUZfxw7JJlMYUxqqzM2bVbZW85ykHRcw3qppR18yuOu066HJ0DKQyKKM
wNKiH8Fo204TCbZB3YIyHEK3/V9T+cZ60ExflcUCM4/LrQM2gFplpzbK1uwz
DwywIzHfJrFOD+ntFqqZwQb11KvnVIUG17EXwuocySLY4vp0InHiUZUxHJ5L
wKZzwLwxufHbHUVDHcQCVlQLj4154mwi609leFIQ6RA+bXRtSsBBMUpwVXmx
KwdPP6RsNWteYYYHtbBXr6iBlbbcA6R9fxQjlU45TqIz0MMdcJvW3/GITmE7
YNhBziGA+TaIfssUfdj4pC2J6uB1oBN7dKZ8hYZROl1eq+ne8XAiB18XqGjt
rVRSo1s1x3LaS4SYfwnVjGftoK8jQfujqjsWKBxrLBkupzfjjbRYILbfaEQG
mixBdL6Fok8G6yUzIRMnu4lRsvasoU2t6PUSdDpCBFGwQwT4sJ2sJ8Wn8XSJ
GtlZ+YedenCwGY+wGsDZFJ6tRIrKFsjeFGhrGULkJim6akcri71GFugQ9+gE
PJ6itSLqJUHa/PJKgc+I2nbfSQl+UWEPJHKbNSoRCoWTdzKMsOaC2wER9H/f
M1oRWhM/IM/DJwoOzyW7rgapGFdZbe03HBokFzy9WnJq4HOUF6FoYe58Dmd9
mSoCDoZXVzJnf/IDUZphBxJxjc40ZYJ90GLbn/3nKtzp67c2Nb/6YXV5nXmf
XObDXrLJoh0kQS7YHNwJk4P3elf6DPdOAXHgHGOIWxECX7yBgjp600JG7+xs
wMR35xG328lRwduENiqdP4oY3hd64w1vjuhrTOJFFWfpb6zgFHywUbkjCezk
NSFS4KeTzVIglNVQJkS9gK06mUQ3YVgwtT3zeoR5yGf+qRpA853r9pPaaYFg
hpLlfZNpXJnLHbuOzO2/YgyVjJk3jmakT9t3P1WFaF2fOK5rZEpH7s/oAk2t
tLmLYGXmb38VdFVaVe5pvlY9DjqqWBkBcOB5CqaFsjy/4uYNpKS3AgYudF5r
IStZMYkeLBDn7FO+8AnX4HqG6rwz6nbnySUhhPzzwFsKuM2gItgQT/UCOeM0
jOA9EPQCjD26/05PYmuBrSI4253lu1qRUUSG2tmz67/jK3/Tk83TMXsu8m/5
VZchks8Wfekk2GGH5EH+4WmDSpZBF7m1DEae1K/kCRhMuCCq8lNlnzlNzi6m
IHe8m9Valf47Wk3GnkjKnblXBUhnX79XCHBH9oqWpkDb2yPvra39BE9T0spH
/FRyptvlE0RW7oTTEWYd8Zp8CT9XBLJvjB7A5PkzyL8krgHO+Fz/8RVBNJRG
puUcM5TegGDSN9DQ+yHyVWHBva5m/38xM8vyLPtB70stqSg+MGKamt6wnMu5
yB70LMjnaiySaJyZhecEDM0rPDnvGNPuV6zKhT4Fo0lfwQJz0uKz88g2gR9S
QzZUOUaTUBfjJiQ6axCPDUIZxwaVAEIPyWAu321MQ8tDesiSf2Kuycl/M5a4
WKXvBFx7Y4z7rboGsFHHz7Iqjf8sYKQbpCnWFWafu7/Qzk5lW4dAxj6fdBB2
8YHzveEkhq/xq7HNmVX39qKYvu2XyqpPRnzcjHqyrYF+61Jyg0sC1gCGt5Eo
7yQ422P8saFFa9RNx4MOH+lFbb9+wT20E0VptMTyN2xKpWJ+SliQa5E+C17o
PVjaSh1Fbdtew7aQXQYER5qvFVaGieyIk1VjAUkJxFlFnu8IrrWmFZ2KwNiP
X+rcxixNesZCSImvKLmRLh9gpzgk568Ta6BVS8qDhcGPJSh37TSARWjdjaOE
CqLJN0nY+90BNQZs47IgoVPiKgf6TTrY5jlWPeeYuet/C26ueJCbcSLeRORa
EsbjzSm7iwDVACoCixmasMz4gSJVaCo68ZCsKgTH7AoHrFZKBKi7Zey1q4bP
Gf0wUrDxz6rXstNy9eUjhnqEkNC1BRnIzE/RUpie3I2B9UHWI0hnKPGO60Sf
UbiK1+/me3+zCHUntyDyEqAsD9zKzIf9uxl67287gP018WQ6/Puo7y5tu9d2
C5zJsD8iluym1DjCETF52y3GHs80zPMlDcueYIKQTwmYcUT1RebDLCL55r3k
tl+TObj2UpRm8QhvSBb+qB2Vt82+uPJcv+cvn6ec8C+YKg5tCQZEd4B02jyt
UwmjHnF08aWXs9LUqC0jW3Yc4ncflluWMijCbLdJJC/57EeJj9IPuzPoNrOq
FqIl86dPMJ179wymCHXf4ihxMiZZR1jXxS+6lMZfzswl0nbgRVSH8LQPU1eN
1DDHn2pI74SyjIWlF7PZsQmO1zY8cYdfRo2W7mVDt3LWG4QEWnSc2vLXdst6
KfVkicBMBGJxvUzaDJQ3V8Eu0hlZFhdgYdsjekuCOPMST8f5DiwjYk34KLfr
HsppLQ+ksmWvyO8QHgJyDYmI3DEbOoWf/maCqTGcNS8QXy4guXBUlBjIJxFp
pLWag7XQdiLKShLJYyRyjtWcrYuTTpulluLl4VtMz7hpaTX+ZCY/6KrU7Gog
WWwHUYj2N24pZl891Q5BaCoPqoQd+s8isVc/l6ZKOdc5XyeXM8HTOxJ4OEU9
kp0RiKTPKqEkDaZr/fF7hOQNPgBVT1yFR85Ad45ZUAIwiefTHttnZRe4qwO/
NGMtEz9oy36vJ8F41G3F0G7l4/sPLyEnKKB0rwqu9P5MSxR+N7WJG16vKG6b
N3c6kdQakHiUZ2vRxEbSPlyZJPxl7YSWlukqGeQ2jBCkPEJ/YwyxzlIr2wa3
jrAuLYkg3j5X/0Kzk4OUIYbygBpgJfJ18Ua3MtAkYWGghEGKm8yAp9BmRI73
G6fLQEBotDyy7+e+tx07u2o+CCdtDxyCahMoKstoVVvAWpSQFjLvWYl3CtTS
bEUl0vavvEhUxA1M96tYGvgNsCEVpnF/fi+S/4vem8BoqEpvm94ulNPsyrrI
RNIKJp9c7iJdXj5mrel0Pc3JtW/59qLVma3jLMret4Y477NSyMbLJLBFnql2
9QWRLc2a3Chq1luwjwrvrQuC9nb8n1JLZetSSfWOzwfL6cb292jygJznTJub
ZvA5WyRe5S4i5K4tJUUVMppWxRpFO5EE9UZDvX2+C6bfK6jyfHSIPIELl/iH
gYrB9qLkVU4nFXB2/H9O/ZLlQ2yyUgRQA5o74qJGatQ2hB01gntN2GhDw9Oq
F/hdnIK0XuDNMxvrAW12txvMTwHABKHM/x70bAknYIHIbYZa6cO/aITLmHDy
wcW+4CUqJKhKlDayQf/vsqSmQsoz/kMxL1Ol3cMgKI1GeTfrrIbItk/OcG1z
awwLnxkLY3ruyftn2yj46eIS92X/jmi7BPX4/9DhY+/pes8+pVacBh34GiaJ
XiuRndO/CBeMFjRHXtLVyDA2HITwN6crmoJW87kkxAJ/Jfzw9AZPTE0GAZuR
kw3z4pxZHHFD50bCYvtBdhJbAHvJng8i68r+vKIsWNC4YILCEhx5sGRMRDCj
3BMde4l6ZhyisCx64g5Xk1zf9Ger8BO7KAOhZyln4VQuTQ1AsF6pp/KY4+gX
cr1o8dNpY8rVgYsa2SHNoEUzrLTJPEGVyA/mzPuY13IED+8dG03LCmzlfIe1
1DsJt/xkM+nUXx3suzR/6NXQwXmjYI2r9M/ZrAQBMaiB3jYpvur6pQjwYbHd
q99M6bEV4lnRPCkXA7/DW0AarWm5tg6r53U4IBwMtdpR9AoxH0nu4CtkXy+7
mjLi8Zuf9I97byDAxV+OZZsKZOZNb3UGEyuXj6VBZNBLHz3AL3Im/04/VE1x
jJE1gFybWTERdcVPSnPc/mg1tNxe2W4+Kqn0fyDe1GLQOQ7inFQV0UtQqwz8
6Xu7Ffer+JFEz3ymTJa1gNrXM+OaMOAbS/ex9KB/y3+ipJmjglHZ/szpe9yO
4DCZcQCAPcawVIjmP+TV8NP9gw8uHlyUWbOJ8GZODWrZU1/BjdiB07khEQqP
LEiehOlEfhBhY20CLCdknK5a02K9FEPf5Wlfaxx8mvMVv+h/pYWMTFY0+sr5
evacEUepJcVWaQ43PuSTwtzzUKhwegoRop9uJn96JJo/UrcKc/iA8ioPxwyo
5ByT/MosL1cIHk0L9V8AfgCjhbxe7Tme+N/qzPjnbB9f4a3rpe9aOZgOr3Fy
/CAzykPJmKuG5AUcdpYBGS8m7hVxv2pD5vvruIIKCUt4o/YArG3nQ1spGME+
+oGNrQOBKVpF2M9Ir93jGie7Lo6nf/ieqhm9Q+LlZ9BOp34Un10jlaV3LACS
8xO+kPeByw2bnyoFRPvRKscmTPNNv6698nEFWbcsEBEgVtH01xeQvjZzd8sb
mfyj6k+at18y6JvkYWHVd+Xzrh4qnH/E4OLnLvAHRoLN+ii8fnoULcf0aQLl
sMUYrj2DNFnL8BQVczEBzljpCVkXls5ACl4cZ6WhvV1sMZLmDYDuyuPaRhid
25+pv4NSJvU4cSEw9vez/YLazPZELniartcJI0OX8el6q8ExXOi7wnzu8/dv
XedR4028gyq0aNZ0pAD9cbZ7pAT2e1XY+3qyy2+/D8PZez/U+UByvlcHKe5F
prGuUiW+N+ysBahcbL7iJAHZNcvbFdNVVizdD0aJRbOgRap9kE0ZpJMjmIp1
rkhE+u2Q98N03iQYskhWW0Qm3FK+w/VQx/noKscefmoPaueQtd4oI6NKbh3L
omTBzUekER8ksvlFNd1SlHN4Frwz4r/I4jpqm0XV/CxX1YdQxPO90/m8nMUI
vZFGl2pjYFlbu1hhm8bWLUgg5estG4ZqM2z84o1DvyE53Nprdf3V4L10GeQC
sPumM80e7iHitku368mkDIY2cIisHmcpDSkIXq047y+mmtPF1JkBoAl3fLgo
ek7wbMpaAYDo2ectxrnRr6wM45j/Kc0WLZMetLc7cTbsgKl4xfvCMWj4xHqS
P5gPYzhe2UDTjSqnBtrzPWcmJKl3Eq/CjhxESQT5nZHn4BldGnBqfd+u4GwE
ylt2yyFRgxPLlHqi3aDgDQKbMDf4GwbFNbzM4ut3sp1Loeg77d/nGVBjsDNP
sId8tqAUKU4+IaqqBwrmSVUgUzyI7pqtTxMSpRjTVOuDQEu9qDwDfCL6kFT1
HE1gtVhmSRaTh9kvlEk82uRNqbD8fexeRn5S+d85AeC1qW6mykW9melOMRH+
pBmRIKm8zIgGNtt/qdsMPNTicF799QYuHGl1536RCojfSuJdVGv5Eji3Sn64
y9IY3whSXmpDuz2zHz5JlsBNb9RtfP/4+jaNV/oyiaKm4lPuV6vNhYGZfrBz
Hiqrx8HXbhMaFnHIXNBjcvuIZr3+qtxx5lcHvV8iNJhg5/FrY4WbtX4zRMai
M6Jpo46vDZTCt4UUVG9rXF5X92+k21w0zq844vjmsPSig3Klej/d5uVW6hjV
c8WvTO4VTeJu14BZ6jqUOV6dsK3IeJsgfJk+R75+I1SuyU6uNRtCoIWsHPwL
LaCKAXObcRsIda+1m0YycNH76Fc9aiACCqDwL3SdOLEwavvm+/VE4yNF9sVo
QoNRHMZYpdqGvfCFjDGXF+yyRXHXtBqM8BYAmqeMr46bg1Vhm7g5Wimz2las
sKGpRsiwVtLLFTEc+/vArzsyFLgKLWIc5qJwOsTdjasTlBbhd7xmORFe6p/l
3X+ymDtqWm2jHLSIvQhtrhUfafA7nONPqR3DFlKbKurkhW0i6BO4okXoCEn5
sdssU89ldM92yfBspNnYnl335jIP/61ieW5O9JMOejeYgnBhnI0g08BQ6eeK
f66vBLkFAypvEAULXBfrkjprg3FGbKuI8XoQmu2ow9ul/c7maYHF47S1Wvsz
irwvj6h7FDVm8WKhrdMNbqFACQ9crlCB+lfIjt/VV7t/4+SWj8nJOxnXdMzk
XFs6Cux9nDOEYblfy0acSR2rZBgLsId3SvavYWHq1rcKWx7Quly7DABmsZHB
8pYotcoYmwADfqt/dSve7JpSVCyFSK6ii3vC6y/z6t0imXtNHYl90CQWDUpa
mM5KbOLUhCF5Yw/DlbILzpyAO4QIrdMSvbbL5VZqM5/RMsONeFCDGJ3Xf4eX
Fyrsaeze/SJf3kSRhsgsh05GMXmTRSSFPxUabm/tQt9o7C4Ox94PWFEU0ynr
rd2Eh5cm9NxbnFM5i+qwdInryQCLIIJJAtwpi8bOBYncoopN19P9K+j/KHMH
H0nlzKF4eAIuD3AfiY/T7eJ/wDuPwT13h2wjAR4ElpnA5izr5nS8CuCfj7c0
fm9aWUPFi11Kl5+fvKvJP0o7hal4zcmGjf/QtClcFWeW+ih6480c0KsgpaO5
DMYmw7taGY9egr7rfln9LL2qrx1hz0j8nTukGgAkqK9v35VW2mXv9Tzp1OTQ
A9ovHi35Wt/M2+xC6TdDIbZpPNvTZ18h1T42EEONh4NLsnNB7PEyi5YBNq9Y
Dpu03vYIF64gifKbimPdhcbvw4Vj/t8raj7wUu3bAHq0z2GBDhJ7HE4WBpoz
1utgauaOwiC0WX+5YnGqy55Gokf2jb3PnEuaTc62dq8q5IBi8utS9ZNgcTjA
OySqnL63IdoQYwLY5nO9wtkmgzNHY8l/SV6kplvsRs4uncI8/d5cvtWlZCwv
lGOdyPvLifJJ7jdq3oE8hQtSz+JhAV6EBW2Sx1/wYOV1It1/sA33AMbOX4Rd
bpCvFHzQAi4JMPD34G3GtM1hFboqG6PUt7lBs/Dnk5yjSDL127WSHdffvSCY
8hlwpbHxYdA7pmTMpjWiwdl84RAT7z5n1DYX5mNg7OGgBK3/ktQh5LllHSzI
n8mJ6wRAIS4R4ntTX6K/o6KznJzlwbacItNGiE8S7DqpKqRn59Oa1e80Wy4f
dcw+ITtrPud1ft1TYe/VHjMtsAoLXv5n/PrwFS+6HCbedSF7SXos+qM19Tn0
KaKRsHUcjMldEu/+Kxd6NHxnEcFUB3Rh0Dfn+MbAyZAaFQVIYBRaRDymFaNL
K2eibeaVpz2ML9Z7oxCaaj4wHa5s0DA0kYR7wFJN+cFRgSOn+yVqQp3vt+Vc
YxAsvSIZKJHzJNeB8mn5xqj6xoJP2URXLYkZnf8cje8ydLKk20FRo23TFjAa
JXf/woze2rgdCfjAPiX45K9MGIop0sXrRCT5uzwZ1p379sWj7aB0PlmJ+MSK
PYyoKpFFQlLC8B8XpSRgwDLh0NoVeyIztrzdyrB+UXAu4SOUQCBEdxQUqkze
wDcBXuvPUT0mHt0jtfEd1HxsnW+uBvFT/ExnMxjSZ73qOH0u8KJ8lFeI4O/N
Oj1az2wAjBnZ5gfrgatS2kEwxegUDsrdeedAN0GwMM/rcDsRbrBN8b39PJ1v
Ex3+r4DmEUkqlzknEHSBUdodR74NjHbDWTEGEq03q8yyXi3G6yaF3puP7L/1
946Adwv3ry04dRTpQF34k6f656xGj6u0Sdf1O8wTh7KN5Jlepu2zwxAJlS1e
pHkEeSmISGVcp23NiQtsbPT7BRt2gBZiVqCsC2HwpqWrCF2uWwTahjtbLwED
dLZNAzXOydkWfHCYmZ064BmkwrYh9GgFf8XgbWW0i5RfJP42ehCLSLbwTuhC
EUV+3Wm60+13D5ZK4sxIzibRX9ehj1WlWn62XbM0jBgWRcLIfZDZ+sZdTwyH
cMeCnW6Y5VULhMQTAgsenMVX40KG8KevDI28CqWArEfG0dcM3Ns7ImXU8h5v
JYJB+ImxRIh888L3xwAzwb1gjBWBU0ZWCeMtqk5gyKTd4Fxlrko1+VZ6dAFk
T3qNqMNuzJ28Aakqlg3wEK+jg52A3taaOycK+tNsfX5az9c1DNkVkZt+n+oF
PFrDvKPu3BK/R3yOXSjpkDeyxlp78kyueyASipQsWlI7XJIB0aCJGbD3G+Ts
z7clOZWPopj1HlIe5vgcsJWWqt1qTMjMgAPjc9jbxUs81IMRnaebvLe7Vswi
e78quOMTQMRjlZPUXUaSpvzNX2j5ng6wA4v2JSXe6saGqiXesUV9GjJ2xBuL
bp2n60lbsIg9m9H8RFq0g47kynyuM1qvQ1S/T62cikrGqy0EnITyyBct5xEs
NAJ2j7xF58J7h94q5pFzUq7gpCYIyYI5wCrwiWrvsh45ZiR8gCYSODsOBrC1
vHmUWwEh4pSI8ry11HEsDKNhq4ithGoRRcj8lcYISYqqtANUC74Fdr18xF8P
ZZhf+fgT8x9k4owZnHdkAcYiTN5yd1ogNzdQiUsL02G0/VWOzOA5PdIX1SLH
pBTw6QkTSpB8uvfDvQtv86QOGjVK0Hzx1P/fAGNqN+0P4f63e/fytQxwVdLM
Oay5chURJhOU8ekBxdPKvivljOb0jCHm4/fY0/ui80/dB6yN+q6spwr89G5h
rm8uw7F7/0mH/yV9qM2RceiS09HLVWnl5faJUUXuQCgddTBBn1AhJJFVnv0S
vNnBgAwVfV5sdMFx1c8zDwmt1I7wmx4JTPc8lMa+zqADE7kHosD5oxhRYls0
WfA3vwffLoW1NuvtPIwc7jhwOEr08qlHlcghMM0F8CJZtOcAp6cW18hThBWJ
+cCbmLoyFVM5T2BFdjWY0b+VpoQSTzDttYJ0kTLaKXXAnstkASBE+8C/mvZi
V+/Tsk8QJEM4XVGpqo6dnrlRYtQsN9wR5hBysHsqI6PUDzP/b8dvJ1JebRV9
Mhv8DDlC4f+m0q6DjTMKltI8oTqGa73kn7RloOWDzz9BkG8MQOccMh90lkj+
U8nHi5jMke/EwWvQ6B8l57XJyKsR1VnZKjIovyUMa3WRoCncPs01dPY5Xi3t
6bI/cSSkLtVh84gspUthkYQlRmrQbv4JfhrmrGqNDO2XQR0PZip+IPWSMsuo
nKACaqsJIkFGTh6VwBDMekdStC9GKXhHtIqdrA5NA9ixJpCB9FV2phR36TZ9
WYcMkG0ulJSsyR/0wPS+eSTgIDR0tWzNtkHXFkSKPGLA9b/4ew7qQamk5wmg
k6BlaX6mCC04+5ODnlk9OMQrBENwZZEiima9jzWMdbzUHxD9WHL24glhjcEn
aecw32G0G41VP09LuVbPtXkgPV39X3e/R9mHYvGPfwT1zxOzu1rjSwHeKzaW
fv/LCcuaRpMWXo1Kn5WfcOdPRQAzdoXIbO6WIiaFrr6+GqmFKVBxTBsa96/X
zwHfnkSgd0tQoHn0VDgxArvYWdRvosypqx0wEvdKwyZRPwmBLZx803QpPWDu
jCzgXLlREXt5tqT17smEjsr0WmKtASiXMe9b5kdJoMKxcT7QMmywldsYhSMZ
VfFwc2nT/FlH5zA8ZI8RcELXTedjuwYTNdutFjOmMgCCLAqva+6QPi2VsOag
+bCfgs2h+cvSg6czE2yqQ+CQQroiB8Yd7tCU77ifvlfV1gncdcjPmWo3Nrsh
KPnOba2D6fH/xCVBOhN4XUflL6qg5L3HvbY+JDI/epqGvlmPe4MM5x2Hcs0c
IHI8BbVB/+0O7EwK3cjrMSv5BIo3PuOSlaT/5yL3dMLIuWPQdyOdorXXqSNW
OvAuwJfB7tEu4UKtQnUNfnlcuQuQXD2cTV9yOiTDHrY29PPm5rQcI9NFdhmd
49odRQi1ucw6CxJI63ywg3v1B5zbxw6sZQmgRlw2CrEsqa2VxUxG8nfJZJe2
TX7nR9XQenfCp5tJWQ25nwb2yVgZ/8kxs4LkA76L5+IO1/OXgv5dWgnNW6nP
jjAOe6rILLaKBdxvygs0dp6fgNEEBjo9FO06ZGTmI/JW6hsskAX+SUKooyIs
GFvR3ZQE1G9jAadan3aZtpa5hNhbjhyBw7a0DWoJ2OkDohbjcQ1kGiiK/U5p
aT5L/j3WUz94nnBTqxNJ39Be6aUPBZN63rnV+vXd5LdqgsqumtK/yV75nlxL
XIe/rnOLpBlrjzp1NdO4viDRpTwd3m6UVszwvlKualDuucZUdteja1HuH/7l
Bo8RBwbCft4kPqOs4+SLVWmNK7T52wDqRL6pQstX9ff5FUVdao+4PMsWFLor
7K1p96+J8RLklrHIRE/+Z6eAiXI733IN1503hwh1q5iGYQj6bQV/qmm1xB96
l8shhi7pIpfrQqHbu8/AjNExc2cuN+r7MZexWNTQPfCBK5aePCXgLhQxa/ZB
+AhKANau9pvuUO56RoXwNwUwXlZSThMOg79wWoy1YsS2N5FOB4y9XDslN+PI
GKY7W9bhBBZ5EWcIQ9p0TRNyfBtM4Bkorenfrux3wjyQ3fz5NvYxHO7QTqWJ
tP+iOCCzNTVio2XWwgNKFaEajdfZCiBMvwQmxInR/leuSpsDtM7AJyQqNRJO
X8NzlD+nIRXME6KXmi7RRRDObbU7fHV8Rcqjv2MSN36SQNbfutVOkHcu+e6Y
1s4RgHiDZmO4biHn4A0EEaDN8tNH5R6hmETGXR3VpB2RAa3N7g4luguMOmdH
jmd/kPU0dqi11cikStnLhGKQxDruxTsIRtLkIbJErIG9z+Dk+eUGrTAWyIj/
OJudLTmBDxiqrdWtwVnT+vyiEkaq/FE0jcYaVbEJe6kUXlvD/4Wxz1pf+3TV
O3gi5m7yXg/n23SRXsKiGX6SpQ7gQTUoYcozM7fOhnx8SAMW3z+3Qj26DXK6
51O3BQgBh67tnXjf3MmvUfj7HnRdT1n5dj6rY5cK6BDPEU3DYbdJRvM1Ho39
cFIsRpFZYYwUbDmcxmgUFQNnPasCZfW2fbJGsPP4Fca+j75svx92RaNyMSQ9
CsnaHoFLlXJA4Bs6B6koPzBAJPsI2iSQCsQ6OntF41eGDJPhRJIO0TvLWDBZ
N+YEeQw+B7aUciGZvxfq6sK0Jhp96y5mb+R5FS9NaC1WE9tm8/VkGKldfMJ4
qqKdOw5QmicO9VYAg0GW5T7jBouODuAwAgc7aiVYFYKAsHKADXbo+Zgjpkcr
YH71sMgWXGBxit4my8WTuquR4q1m0FZfCKinTziPZd5Y7egV0a32U17dPX2W
VNm0AyNT4d9FigBmhVAmzzk1X5dLgkcfOXnP+nYUdIF/b/3pik2On6Ej4wUx
KyPmbicCk/F+iPW+4Iuk/GGeCwb3sSnTLobNjMO5/07VkLPNXWjV8X0auMWH
qCCrsjUokbTHwGLizG1TDqwwYgdT20cvHHiWQPiDO3K+gkAXVQTzkuirz6oo
+X5lnHytZOE8h+ax39vn3CIWzbB/IYgTyGfXu/qdTLtwmcd8vSmuFJbIIOIP
1G3RFOEUsRCTlYOP4X838SNOgclOi9MiZ0R8jrzdxa7qsi2V33wLtdu8ahEw
WTvIClr5i45CSSiIDq5tCnFHhN0M4syu/7pb+trBWMurYeqUl/0ACAGyrLqa
N6fEeIRae7Xv6rxWFidhi4XJ65P9G12eGi5J+3EgS29/2h0AIRQOafj6Awd/
jz9yqZufagMYlcR8/k0sOzd7a7nh2YTB38TvXxsvH62XptS2uGtZlMTFQyTu
CbvZ+k2fB4CnWNZUCGcA1yITqyXMlpdpr1+MPZt6e7JtebkCldA8tab9WkKS
l3Tl0puGg1KBbhYAiRYeMtOPwrZmcfjvXDVgkP91ovswfMr477emw9TTKoM3
y8Ez5SWm6J+B/6aN47lRRfVCbmppXeIBLJiy4S+Jax2MYWCGo8b7+qVna5d4
wHF96CpFIjUob2cdX0Lwj9Ki9TXMLY1UDUbH62pkcUypQPHsJYNmdXiiVVV8
FSlqHZoKR3foYXl1/+ZCiDpQbGg879UfiNibCRkS/BuAXmR4sp55WXue9UL4
fyxQr8eaEdQijAq9dzBeQV8J966U+FI01I5pvmuc8onNjr1sr1hDg8G6TP4S
sYfUu7O25fKG7Mt+BeHExM2U+NTkdthZSKC4I+SEAO//3xENDnztz1twT8hs
pCaXhyXX78tHRYWVoJoGt8NXCNBf/Hs21GKtwNyD3CEaMzKHVn0oRKFDOeFH
LoKhc7phKyDjMtUVxBNd+E/3jlDmdOGtCFCeDEJ88oD6MmMeMIXU6DIUadu6
ZaqHwXD+nQ0HbjDDcbfV1SIy3Z8rZeq5Ai7eHsERK8GYgR9POPs1km/w+q9T
exx1s43bcByNMCl8n1IK/CaGEnyxCkRABNrchW2fg2gzwSONF2WwmYIed4LH
3dc3HsJVFfJMRcWP7zECLm/zm9FJkPM3N7ghOFMVOmhdQVVOIrF8TpX8AmR3
q0QT2UUVdD9rZAIAmiy9Y6xMHn9o9ezIDmoKAJQBESRr0Tj3Ogbaz9xXLqvP
QFyLyZwzHjP0fr1n8QdGEVtDUeCa01hnYFSmPTkIbEyEyw52iqJxfZeb1cIt
AFT18lDd6w40X5Iscohb4+DXzyXekMz96hmx9M8YNsNE3e8uG0Oi0nUKf0UD
8Ocx7nPx35sXdVmvSsmhpun+Aqi3nFnuSlbN4+OtQRgpSxfn7vNcW5Dy1sd8
LfU8oNIJbUGzavSwYWg7XwIg7/lGVqX1U1puGZoc4RplH3mL9ls8D8wdgyJv
0EH5PpaFKItm/r1z8CZ3ynRrfsGKtjzBoCXRSU6MbMQk8MH9epDAWtR4gpT/
uy1ISwFGfcaz9o8vqZQOdMM9FKqBcoHV6Hxj0AvPd+OMQpX70YciOeYRsee6
yP8MXItljcHU3I+ArCoLmpt4B3EH9sDCJbeT6Uk2IPp0Tk4ja70cy8PA2fmq
xeHf3mYay2EOwDAeZGCEz/L40hHDwcR8FkGwMIqAGQ7ajWzptDbehbDVFvcq
ebq5zFy6A4CRCw5u7LNEZ/h4SFUqbcROOcsm93B7ee049GV/f09jrkEDieE8
XtfVWaMG2oUYTYiCtcBMDzyUliyRALkWHUSoXx/FjtRihtTOiQ58uNz+FDSy
jTpdVvhVWYVCN0j8eBqkqoqp7uLgfiZdeqxPpuWbQfyIy+ygKNO/npvJF9IW
9GlQK3NcnyjCGdXzE94iecQfHn74u79GHu91rR0+trYYrcwKvIKhEOAnbjWB
Dc1hhS9xnvstaV+HMxA+e6dYRDMpmVO5mbZL0yGR3sXRQO+yCtXK1+IY7Fbb
iCyiN/XSOaQfrx907x50ixxQ9BTcK2iGgXw9NJyaW5mvnGTfmTO7CuweWyB8
Lj7kuslwrSefAkxAx1pb8dLANb/akwtc1C2lhhn2R55GE1IB4oBYM2HJaQNx
WQ6ZrhKMbAJL775JlJlAs5HycG7O8RToeYyYWRoElODFb2bxrLbtQLIp8R4o
xKAKugVT/8YUtG2jyoQI8pEqQGx426vx47utfcnz5neHwNqiRLO3jpTaBn3l
Xk3F7Q/d17OONgxbvE1RCWqnbAvg8GAeXoRQ1n88R/tZh5cqJhRW1dgsL6MD
QfijCIHZrntw65KzobHNIwQXMz7YSlSEUgev/1VsdVQK9AdOUrMcseSSFSE+
XVTR7MI2eRepIp+MSE6BtWVaehdLR65LN+xVjrr9CErpfTnuQr8RYd9KNYCz
mF2y2c76qXvLquuB6ADxQYxTX0cIjYd+g5UI8ESdCTNXEz7JlcTvlVK8dPQ+
W+dsFbvpwsj4zhmVhpJZAomloUQvcFTgkV9Sv/RDDeyEm5yrfgMKUZwBoE6U
kLjClGJOjBgkvhA5bHwUuEFGu2rxItD28l4IOsCsvTHc2u0iXJpEHNeU14yJ
aIgZ0EBUmmzJC1oPcsFeetISEObL5d7CxwWHJaup3ahW9oTt+9iJlf+SvaKD
nMQKmCkv+TAhAur5e33sgaOSd5x7sItXvg7lkKC5UI9uwjvFYBo40UIq6Gok
aDFOHLnpbXVofcqQ+hjNJZ1Bj4Lu0V/FhvNXpmxg3+o7DvqQP/naqKsJdrxh
VbgS+SHg0ZG+ru0dpfqFkhrXgYZIeMGhGwtzwlBa3hNnHqu6WWalxPvY5vR1
KS1MTsdF7+P36bAjKta2lh3ICCQJN8UqHUC59vfmQFd8SJVFVC7yF2uw4Tr+
7Y3FqAfUjDWCoISxjXzxgi5BMAkzrnm7hBi6opGpKeKA9CFAeV4yMrqzBL4k
H8P2LnusJe6x5zRBanedbMfsktPf9pJ5heNaCIgTYUNlC5KMtHCUGOYcnYve
J0b95PNtuJCGKORLsSmoPD9yu+pu9F1wRFIwyHvutsM29ddKHXlJddjqcp36
jyQbosFC3tIwF4+yeHnV37EiBiyAiUnjSlhA2JjglojUxm39SCGasBhVxIi8
FP1FGWz+wlZg7CgyxM/zehOBxMlxf2exej18bqLqXNbXwO7GuX6wMnxVlzr9
doGNUzsTC7M171obucm7EmDiG22JE73FRpoJ8YwXH8karoO2Ggb+sfYkmkva
CJBcWSwkSjsiIyar35V3at8j4Rt191I9MIOBen8/JqjH2oDXXXSDIaoy38Dz
HptvYMVvbNW6mMgSFt3I3/t8OaFEdzOxOpBPKtzqul04iR2ec3M3DKp3vIn8
zOpELhSD8ToonKRG1dmBgfrUXHRNSrl+AmXjYlCP/6XtwDkAhXFmAL8PbeaO
tQfJZfuHbckmdrqRIng4Lzy5e+mU5AqCy9rD6wH8OjFgc/A+q61LHVSd7LSI
gG/fP5NsNg9Gyz7fHebCBClLH4x1gZcCUXqmf8EX0sOUo1aWK8a4wcO/EQC4
lmCenPS+7OkDy/BTTP/JR+vpX0Lo2LiGyP+GL2HPbmBw/kSo9jXNotr0ggIo
tvWwo8wByoU26gjuOlNIYWs9AURmX5/JV4ncKa0IKpv6+pJkZu3wHqVVetcD
fA8WDMWZWPtZB2dkYGa2WX3DPj5AHC/gy2CpkrPxrmDsB9OPCpk6MPEWFz/Y
MgSdcVcRwKGDQZ9psUc2clITo/BBcRqnAWWJQKZjZLKcOHXGFJESH3eH++bI
9bLniluflSFsWlqNBuxT0bxTyrCNzCm9fQ0LdlcHqj4wb6EyUuKDGQ+7nw39
/sV0wwXTNujkW5LHDCA4Zuq/ZVWomXY4W/UNQxZOJesmofH0k7q4nPevjtRa
MKaiz2I7P/02ND2zFgqUymsNW2DmXRthcMjrk18HE0cBU378lAuQyDx/jeLl
h10bypKNTN/1pfF/hcxCJcU78xeWYvVvCa+R6hCwrfn8SI6CoRzBE8IBHlF8
k2Dqe+hAtFarm2YriVwJhnlsSGAdqKQyZ+8tCiJ+SNdb2kVewR3v6hsJpphM
i2PRmKSLkrdBEZEDoKu2A153opX33hqYEt7gbhWMoE3xE4qV8qveHq2zmpfm
5hAAlVLMEmVJIgIVuWT0SJFQ1RZ8gtd32DI2qkfGkKpLtieVY3Et06KEmPsM
7hjK7RzX/ewrn3i3hbdk3g+saPgbxlj8ul1Vzn4fM6MgcTzhtYGyFW+i0HKQ
axyqZVnRl7SN6CjveKVDos0vnqMhjimr+JS8EJZ54GYqDkzZQ7UWL66xUx4P
Wpv4U3gE6cR+tZwpBvfg+XDUbnYu/sKUgSQ1Epvtv0q5dVhkXekq5WShCKzd
yw7M+f86hGGhdjvewFYi5ozQ07vTLETxqrUKUT/POBrom8tpACl+yleXr1CW
qimR882Hm87ZbAlhlx65zPencjKLbcEmOS0LDzZBEalIDUJUaqnqukl3ekxA
1BG6Jnt76HUlmQWwS4jItse+evwDBIcBzwYvBE3wUfrAJsAVMveCyn+a5ZSE
wXU+GQ+wWY/MAf1dPVTA/EcXpDEtWHLSFarATG36TgWH9b+khMaFTqFUGP5j
9oqaMdHnT/ocU/ITjvIEfzlK6+/qnENA+jnyJYmhfHL7Jhxa3jwUCFNPrIdJ
6GN+hUXFmmyV1SCr3ieJFr53uU3i+7kKKAoZ/2LK7VovYq2io4Yj0z8K6WiJ
+aZqj/3/LYedrnyPZMUwBHB6QeCCIcgViq4ID99fWAW/rBmnAQvJlPeck6vw
/fDL08XZ1oSLFqcxAfMrvUna8OL0pcJAkrU4N+DYGKnfMRQ5wMLksUhhgpR1
ztMfVWZBWupzG9hK65v8eHQlK8DPFcvnzt1sj2wQjpS09QtwOQQ5NJNunsJ/
m/G5KE3jTpS1OO1IYmFvdn4uNbSw1aQdFdXpk8/C0BhmSPPS9eaUD8sXy3qq
taMcd1LKX5f0jxKA0EmFrNXgVlrKAa/2u41DDYyENagxWRwp+a2PMung1NJq
6RJBJK/3PiGml56ozGlyHaZXknp+SlNYDGx4sVrXAoNUvtwgHpBv1+cFv1lE
JC4SepYdTL+HjmQJyYg0Ss0ju+8JWnxzmCDPfiofGp2tRmeQL+QQJ83Ig04h
33o+VLICSIR2Hnzzs8fCVFXMpS42VWS183csTGPrVImY7rZUZ4gnfidZ5Q19
J4YNJ3/jd0qBn2SJtXnmv+26f9EuXg3c4JnCvGAJLT4cQdOB+U0xwx/fvTG1
7hDIf4kVq4Q8DqhPbRXokEyZkVsNppP+o579HadPgS3yqQjwoBkFM9SZDmfV
//q3GrB8nAxRRO8Bkb8h2qco3K1fzc4lL+mo8w/b+Urn2EFOzKkjmfxSqg6t
IcBh8IRPAgMR7jfows3KpxLPeTsBrpt32VYDFopotdPPLLj/JoOd1JBMdW9C
4a6SiyvGx5EUDHxy5AvX62vawPMDcHiFzMITs/xiWZv1NvZo8F6iMOZ64sST
FFJ+G4xPoC30HT1cyvMn+kJ+87skjmC/Q/4NewgbTY2JnKkSz2Dvp6AWCGYu
p4yfClZ2xfnIl7/bsYpmyvo1dsyhFHkGNNuIx6uVs7gIczxnomVxNBwS/RBa
bvBeF28lj6GpujXRE4m3LxPHVOiIvNjlr1FvI5rSitpbVePjPqohHdAV5t7e
ViE5iualKUrNdK/Zmjm2qBlcAVc6L6E0Ty7kfw45riBLiYvnUDTLciWWhFdg
jdK87IqHcJnTU++LZk6lc8QfP+mG8fdCMpXYnFgueWi9Emm9l8v557Xq/gxN
BCqJpVDmXwJNpcbDdr4Cinskm6UZYbo04VhJ7weli9zBYbrJvYZXUcKCvho+
VfhipcaeaLoi24G6m5vMtyVwfPkAIAXUdX6XBI05OyYXf1bjpwoPAEX5uhJV
Q2c1cFZ9uMLjZSMYEl+0NRScI3rw4qcP8Q5wvYcpUsIfx2aRqbTWurR0QfBE
p9usid2/G7/cf27sWW/TCcdHUvC3SM8O53bwJknkXGOJ8XCTkc2qWTPy4jll
ihbD6Ey9KZw3+auPnQfO0znfI13YaLG6oTR135/kHoIwTAtpxSaEcDPNIHGQ
CvL44fTEE7N/7YGFDlnv8WSvz69ow/ZHA/mLTlfalMMAshR6eHwRqZPBP7j5
II8LPerhGLbGU167eVx6G82aIAvRnhEnVWGlejNKi1Qcor/Yjotgk9yMaYol
JLVDi9wjM6smL5O3y5F7Ig60iWsbXkh6o1d/R+WEEp3NC7l9k1L30+yXFbl1
NFtSrTWuln+SOJVXL/m6BaAs3OJnpjgDWq3xoAQ2F0k5pBj9Vvf2/bZAgdC3
C++WrZacOb8fDr7leVf+7XlX8OSTtO1qaD4NYvB7k/w1G5cmdjJQpC814Bru
Xg2AJAoRsZ3blCfn60zye+v4XY9w6L59k0+emmCXzEsJTd87J5FSQHgY1lbt
WZ0JwUSeztXpC4WeyN9Ws16lhSu1mGzjv5y7QhvoZAlH4o/gwScnC6E7QCgq
qSH7jj/wjnJLZ7TFlPkJWUw/sUe8XZnlalaguk1TGQKl/AMC1djKldv1Eil1
1FGyuDUaR4mDmmnNph/gfie2NxLFxBmpOHo4QpZKb0FcwWdozLlbujZ3y3Cy
5btatDsYT7VfIgaN/2uIh3DNKwB2W/UPakHX8L5fSIsuTXy21ZfpmT1UX9VN
tzRHIepDVmZ9xlbN4bSqfefGHPMiRVIDRHs4IpdKLjPc1uYeJTDY2mrSeoNw
NDmotNQPsb86/zpt5Q2SQc0VWDw6OhMwJwozEfhi/R1SbuVZpQomPJEgMnRX
bAd34/O8ylGcjPC1kKLpOgk6S1qfi/p0wV8SmakYBKBR7SlhN8HHUde82UmW
YNNDARmOZoWYOfrthxHHuZz5FwTarTFdBewRdPDu9gG9HtPEBtSMCw819jL0
xNM8u5vIRscZS5oL2/UqAVCwxo/2hNrxP2DHh/K8eXFbLzhIfOJKa5s6I5QV
P1nnlDdvh2MQhoCVKEnYru6iPRKD2mR//T18pvDgd31yKXzxw/42JyQb0kHf
Uan4hndDBQwj/hpzbJ9TtTR7SN5p/+E5rpNc5CqkCbpvI2C0OaUMoanMcPjd
2F/K9K1FvBdjb12KFxtNhKcmujBVTIRs8QxNowx605f5ewpE50EGqVxlY3hR
6zX6laHCg6pgYEOHJwMR71Wd2aQnSfn2HNVWDi0+Wxjd3yurQzvcU4h/xpNt
UTy4ja9QnjWyocjeohm31gmfGS64D7FVyrxYzMXY8hp8M/w50FKWXLC43lgO
H6jrjO8X+lsbbedgmHUrZxX1/JpJaLEVCdguHnDu5X4ShUF4w+o6URRx/L90
YI9A1ZFvAocJ/l956dP8BvtTnRTYNCxdY5n1gB1LAUR/Px4QJFjVLzSVgoI2
OxpSl0FCBXhL5olRzK4tiPuC5e7IYBFgpMkHLz1NdL+VgI54VhWcJ/De7DcJ
ea1QCPr96/G0hBvm8f8/M//uew53o0VHtXSJDupE4sXpz6mz2FoUjZNorUz6
AajWvKu+18yM+pbXAHU9UQoqGD1pF5GHs/wPfUIeu2U6h5YLrpKbd8os768j
BvSNirOq0qZ6OLwiVFz/lRb2RuDHummHO5ktaQajaktNXSBeaf8oOjuu1RN0
Ps5Sqn56/lHefHikmvLeADwCY7d8QoC5+6A33QcWWrzTzxDUKBy1sJsKERNS
A5uEzBzWY+uppb+dY0OHk+156GLEJdNNLnOKz9AZRH595aSqsguWw8iUi02F
Tg5Ji4RQrU4uot2mWcisOS2r3J1UMv3Zdr5krMZaZ5u4s/4yWnCl+4yP0t5H
9TdiMgKsuIdnrrRBLbF807DUYuT3a5uGAS/7BkTTMcfWlr4g+c/Kq4SzWCOe
pYxxp2/y8eF0zwV5oL8cbfB2qMTVsKRux0D3q1CXG3ICXlCgtnJd4BNSMMZN
I6Pj7poraFOyNaPj63J/4afAp/cvB+b+GBQGsj2Z2ZffgwcbRVl5fMtmBsxj
S4K4ObF7IWiopBX0+KqfYYO89RRpgz1peBb0iTtpyl2HcnBnJ0IHysdhkN4S
95DfAtm6evBKNeXfg3TwsMQQPfLCnbhZI9z26xMI0NdqsgsQgq/GYF+7bu2C
XldmV5zS9qgwC9U17acknG+IWRVx5M/xdLmj8hrYM+vDLgGd40IGouuDIJel
Gpmrv/OcBJYpbM20/LHrESYxRO+RMzqT40hhpsTWrAPVD/ctl/LWCOzIFk3Q
CESDNRzT32gzogqa9jPulyCSZ91TdjW4RsyG404U9zKIUJ7UTIsjK7NAC1cM
LolJCSAHThazwGuYh0g1zL2W+O8bLxw+U893CoWmKqWwcXQiP6STJc7oUbEN
VLeASrjGl/TSA+8924rmCZgk9zz42GBSpE3CxOdB46mTmVatpU7myr88wV4H
JxmS95rjjnQkd1maDHR0RggzBl3+nVK925h7akudlS0tEApz68FlCX3+3HiN
Qm/AxZAxoi4mDY9Mv7Pg8eauEaK89OGjM57G7+PIGLS3BDEY2wOJK8GLhrVC
6Ig0490a+Ksl9F5RtM5I+AUQAWM3H4B5enaUbcuarpBQCsw0A+D6maTC/vbg
hjj33uPxJDtNxbGdShgOFLx72+u5siMdS8Ms3TzLmnP+yuJ+6NLqviQzrsYV
r/TOJSIsYGpF8Lp3djyz0+toT1WXRoXhaN7Ou//Bg5WXGYgPqmzyfI0WfVg6
W11/MF4lyrziCbzrdZdJy1MZ33FiJ37n4+Si9Elqsh5vYb4NlEenXNqtQH3O
pSvEnlfE4oQtpNq7fq8G06CKrA7utmvuc/CdwX0m1u36lI/koPZe/6S4sobv
YY+KMQJgk/U/q392YmWmXwErmiGC9U0pZFlL2D02akZoZhdbYUPjRWJU2vCI
21qqNq1Voe9Wrhoh4cXkDC/ZkK1Vl8fxbccti45YVwNqbbjXfWjThNj4DCkJ
Mw8vjzzauH2taDl8spuy2oEw0d+yF+48YYoJNsKQ0pkmR9B0Mhws90sOWlnk
aBV/3EzDFWbi0J9xixbN4qkmz1w/cXlTnnYCrMz2HDqSdq7k9HJ7r0CBPz2T
xUcMd1zsLLAC/k4nDNj5nW2MbB5Ojd9tYSdMyPJ5OXagvjAEF4xf7QBmeE2M
faTw+vZoLP2ftWlmZGYJJFFHU2PUC6ClQkZarTjqMy76IKDhsCPylhkHLmAp
B59Gwau9Hg8ogYrcYNiWAeTZ8mGwNsW2ILhzlJ0l0RiXNH3D/rrfFDdvo2Ko
8sFiGZv09R8I4uGEIzwtVgdVftQGwJTUuVZWB5e69nk+ElTq9szAfaqVi3MT
/QrmIna0jGkBva0ZWZONGK/Ebt6Ukg4YE0RRYqW5S+C2BcfddbjItqt3ptWM
7v4Cvb3y+K3Zi5YFVkWJF+lVP1jzEOddTgLH8ZOgyz7vpOTJ7gQtNVMXDIjF
HkYfT8HArawSo8Qisnf1IeIv7WQa9ht57ADM3AViPpb9xbrCEYEgZkBiEuIp
zFCJt4e92rW5NCBkEB23pU3Dij+IasDVIJocI4xRe+mMpSWeKIacAUBMRhTF
CXZmQTNnKxGYsGQtGKqiSniJWNXylYXO+C4tuDXbx+6wSmIqUdldwvHon0I7
+4HSXMCBsCmdMfBwl8cEfbJA+zqklhOKx9ROaOLuCvKLHXQ9Fw8LdYUY9550
9qUpGPQh6V2+Kb6vBDSp5VX247K29baNA52CqDcL05sZ2LRTzCd1Gq5D1Y4K
uuZdl5kb9B2VYoSA5jNGN/nNEEg0VHneiZC0lhY5RmtnNP0KWT32Ik532aSz
7wDKwp4HO4uMtuwgkSjwdJusKrLPiGmD8U4Obi1GgUaf78KKyGxjyNaYMelN
AlMVkgcYtqbB5ttnVf/64dnQnrnYE/oOr+C70cyQxOHq/+lHTrcUm4Ztp3wC
yK8TOmvlNaPdP9Dr/O0k7fpaJovrJnRrEmJIseA3WiLsTUwBHjmydvqvM3bV
Gpd9HN+IvAKbZuvPMUF8faloCvKzNvazmj4JOIM5b+q3jF9mGxbxM5gXb4hO
VyyZL1PtGoZeCHtCSU5lXxbx6ui3l23I1bgQ87SWi8A2byQChJyRphz4R1mA
BpHebQR6NzKXifu1XP0MlwkI7Iu3WgB1n2p86qpYA1gSvn0kPmNElrPUE986
D64zVA2PgPP3+LCZ6+GzoGP/JkXOYScgHiPR+Pvura/z7X8OKBm8nChPm8uZ
o6Widypl6gJGt40Qmh80TlJSuduYgAy6dVu2Ogyv0pRfW6OL8qUTQppzzleM
dIKSKQPiUGiYxWO4AF1NjzWgkFLqawW84qnww9Upl1UyDq/bXefj3Dix7GF9
fMe+BavITMPD1iwFkZfIoFXHAdXY89EnpZxveGMmazC9ki1X47NKTuyknuk3
YFrnjytjHRTni+LxX8VUTQM8Fc23LASMmnHFU96qQg1Ohw2fynfHuD9PYhWp
Jq298erQD7wj8Wzg8JDbwHFtVR1Q341p1vebFKUYjGgxzRVANKpsDuKKay8B
m8GNFhKnXyRCYrTSwxuVnH/YEozM3U/PpAOjFMnZ/fPaLt/NvQ6oEBzzwtw1
xwKiaXpOzYENaEvF9C+nT5pX3zwj0vPFDaECLR5RLPULh9HS4afUdGZvCPf4
g7AtZ7NL3yYIebP7zaODGE+VSMQ/KJLRW93en6pzW0zO55tAGGGuqmeHzdWS
2PNOjxHSbZfgtS+PuVKdU3UB7ofotfOpP0etlu3QcilTqubUZyq2QpFLIWDP
jMdX3dlu/9zcz7W9/ZkKt7TDyMz7JN+/m3t4tQxbwnLgzrqvHOzfkC3G0XfZ
fiMgWkM7dPaxxlNrAXM9NLV2GwcxCP7yx/lKZN7Gof9MdPQ+t6Q77aYaJibR
9FCDCQRpExSFHLola9ujQGcUtRNOlppO4f7N3D1hIrvsexCEemHxsaouipVX
3uu8WnWJVq0rCENZDDQmN/RdAwabZWKuD0nfy9Beh+fUTEv6dRZTPLEc+BIn
8yDI+yGVXEmaTB4qJHrcj5vai1MfcXkk3b7novgf5FOXo1axpKuEOMFhMyXg
NGwzPDjeNZO1+NpB/MES9/Na7uOcHTeSftmyKaeXwe9G3yAyHJGrFHyROumR
SxoD5ETdZC6aWEzsz3j0+zRyGYcHhgjMnAkc4QADQmhfUzt3kQrr5E4sh7nM
QzQN/jQ+f2MWwO1Sw6zaWPj1nHINVc8/5sNUkeJJlNjP20D8sfMN1V+jLfIh
ap6Hr6Bv8mKdEWQsjuif1KnJ4WyTMBLU/aPLkiQHR7nVLbIc1vsgN5fB5vj5
lBjTkLz3Bbn0g8bM1VoiEpIZVXRsZhgdUsbtLDzTYq/a9gfX/K3EzE8zLLE/
eeH14VtjjI6fak5UFf6yHF6As9znqzFlXqTI69i+rp/+ivRkUZuarkbCeWwp
mDV7V8Owb4JnfZMncVnZFgqy7Z0+Mghgh+hkSXb5ElMgbWcdylIG+PkvQJm3
pl19p6lZL5FQndzS7E37fH42O54YxOzRYuaZXAsABK/20WcfxZmpWDA0sTTp
nFumZyw//mMnEC070BiJjXo76pdl6zFd75K4izl4Zk8Pn2Q+bnkgfavKeDCu
yux3oFrAaiOQSGgYPPuGkVEnw1PhZEbfOFM98ITsFYhl8c0LyFLKhNBF4fes
bs7BMWl+yHAQ72ImZ8OWM4V2daAjXUat+CMnkRjpWIhgChsXCkF/DtkDTuu4
rothnO9RwGmFKmD614/fJuer3A3JgSaXbB5hIEn/QASclqDQ7FmAROBxXOTq
gth1EIRpxIyLiLTQR/1FrhncEGkt7seog7TgEa6IhgolFxgAI/7y/+arGUyh
Ri735zH/9HHGPesRkyv5otYwXV89TdnCLI58HLlg/W+Zf0J9xNLSc5EHOctp
72GTU6nxNiCVkA15fXmERU8ti5z/EvsAj3fWXXwqVyJCR+jxXY+FC8UcsyA9
Zg48tRDM59JXEXyO0xWWxJd+pDGoMOIm4abjNGiiFKc0nzpaqOh/Ndc5kRA+
8xZ3zB7kt+ZJax8VDZGZtrl/fqo2Q8fnWu0ZNT9e5oi+HOe/hCy7+Ko8xzlT
j1rH4c1fyX8Qggpf2XiVmEqRWQAXNkDYZVRmpLNJ+EDKo7Iah4Q1aqMDIfjq
bDYBcfnNWLMjjMureyl6HTVnek0MHMt+zvBlW7585tltOmZB1R8Hyvq7jsAC
174pEifIGv8RK5zduIFkyUNLhdMCNptHLJgA7OeBkr+o/jEIOMJEsf0OurbL
nBwtzW4ZgM6tEK1dxjNgB+B1FegGaxops1VGCIhTchB/R1y0osGQox6KS6/e
PO/UmYZgNpw0iTGZfYsx71Jyw6RGUV+NdPR2Ry7pgEgXp0eNTAjS0V/6YDvX
DWfxWOyB6WP3Y/vdrEEWXjb9klAhTt9XCIWSS7SlZFkWLw1aGLjPEPBhAcx3
+rgvRMvCioT1pSKr2M4NUtUcWJsmGQ3eThrxI4F+V0jA+jgTPBPvPUpDb1ai
ucCDkMq7iMIueHh8PCcitzb2s1ydl4gL31KvJyAg59KWNUib57YedHB6f58e
1Wfo9bxNStBpNKgz2X7PoSogq/CLTyo9u2r7Ktx9KqBwl6nxzUepYMLi7qus
/hFB4UY5NvDgOxU50VfLwqH2VIB3xSLN4my1qXE1Ug5v736+0aXpe0BAd78F
zEB5mTZ24RzJGAoRraWB7Ky6Lb9GGDhwQ4zBbLU33YO2/+/g+dLkMTaHAcV4
J7e3HHVxFUxN01NrFQcqpAVn19+8oCK08PUOJAqRvuQQ5kkIJ4442mYR9U4x
xF6GJXt3YCdBV+sTnAIV8spWZbdh1xM85nTff0nP7vfIUIBuC3o78B01it2M
Cx1tagt8kn5w3hh2CMqv9R1GhrtK6K3Xq7CX1t07d55PuqKWv6yU6mNhZYH0
TqVa5+HepTznLaeOxqSPpqN9XgvkVg4s16PMLDt3WjD+uqA859WAVDkSs9Gh
efAtZ5OHrJu+ydsHKAj0eON0tMg+a7xJVCZQrFuVov8zIJJ0oahdWU2IS2ou
J1lZA36jESVAbMnRIYz8rbiI5KOPDJxL8mC6DQo2A+GMnOtljLRSne7ukKn9
Unl6zPBNDUjNQj+E96LPpCN1AoOUpm0+4E9vYTAWrDdfU2x83hoCfj7av4ku
TVNB8uMYb9TuJgJbdSr4wnYAv9fEESjO6gSN9dAou4gdLzmQO4+HEn1GPNuR
lTCy8n66whG668J0aq/bpn0LZ/YTOQR+EvKh/dojPcjtt2dF2zjPmNbdfyMV
F7AgMc0vh5j6qk5hmLuDcD0+zpyaTBc0wi9dbTqyTuY9D0HExQx46NES7/Bk
ZUv+8o+ziSdsRjpfD5LcrZz1tsKExQZ1SAog/s6osq3X+FR15Wuisq6EDnCU
YNniuw52z1ip7M9zNExDWpRPw1Ey9RBvLhQxRg5GWvEljo0wNsORjv1N44Wa
xznqFaUznu9McZ0MAQPNcJMby5h/iznBEIzDAkRnyQObLuy2RIND9cfocIqr
FnXVrvW6gTX3xeIGkcdXXdH8wWABODXDEgBpoT8JaBet/4nMu3Ui2CrSfb3S
hQecUPRXElzJV4Xgfxys53hYpa/F+FN+uKmOcNuOM15O4hZ7NqL+BAxcIsSi
KTD3pGD+a2BeUWa/oBH4u+WB4z/umDYwMtL44a9tGQU5ven6ynJFypLyzvcF
dOXMFH/aI7eMVh7dVCq+sdaPQ0Lp74L7VnnKk4qgdXRbdmYoCXYlkOlUqQBZ
0Tqmirr6WOTY+pZ3ys1GZpAvmehp+a50L8GYusrvi/uRMZS0EveTdrnTzF7F
XsIRjNdck3tuj3KlbPRA8zrqJOouer5bQuueodUDhIlgJERu8wlOBwcyIR5o
k9N9hOwmKMLuMARou3k7MHx4rJkb1ydY5s+xTkmE2SnVYB2jxm0JdYWSvxgd
biaadQvNriEluyO832NmwQYSS8rkQHyh1SPPH54rlJsEi80V7E1miKDz+eve
TjBgczFFAZ7i87tGL4Q0yuednqb4ebzXPMNST0zvnhww4CoKyv4Dutk4P8zu
xe9lSdLyo1NQVk31sKne3ER4Zk6lZUX49SETqPWO8OhMA0RW/alD02VNgGcR
DOji1iy6s3SHPcgVhymk7gN/GsFlR7xB6RsBX0gcy0hxU4BqO1kxls3L7D3Y
pNbXyGTXQte4maV5/vfn3j4h5ieZ9A64L89fcCLgcTMsYDc9g3oOV7jRjOaV
dNI5agkygEy0u9Qpjqt/kq6uLkJp/BCkAXcxdO2u6eGpjNeDj1N1N+jnTIO8
ci2hwMVqbNYI4R+OGAbMSSPNeCOttsrsyT1cmF+PmYQXhMtyyO4hKWfsXxG4
05TQxop8ouY6ussEdFaFWwYVghx+rsUmT+TaP6e5OQBHvEerSzM26Lpe75Zd
7UXrt2F59tkOfSONIa49DHep4a2TC7v3W4namkaWpit9V+jk61xmKoI7A6Rv
8Z+THFgS/wfZcsYIvzmWc535lx0FOUQTQOCp/qA5+pIkxMX3H4Ca8sxILRPR
eR7u+wr/IdyE7jU0dd3tkUKrwunCjWT9DKfpeD96UVdgWi6nyr3cB26HW4Ya
CyUiJKbR8aMGH/t5PYnMuXwSRXSPDQdovUvLQ/dJdfFis4Wwr38Q/57smseb
8dGNBLvHCydl7ECnadeWoFr52JK8hbBzIrhS9dC4/v0U3hn75B/q931Cuyrb
0J7kJZXhTfjY4lxoZSgNByJCDontIyrFeS96VhrIkXpIqAww6xowM3QA+aVw
8FcfIjDYGFnTlBTqW0+LOIAYAnW+VrZ5CWaok1i69Hs9Nsu9qMC1hRU/5bNs
q//CSbwBuZCV595eZSjH3e0jClnAGX4pjbpHhmDMVUtqOWgSl4EL0qGkoJ0X
YjM+Xw5uvlb9Hat1V85Q+kG+9EndCux7H78VXNnfZgrUXcNoQElqu7FAwl7v
MnwxpAO52kcZavU9YPNo0hwUS0dEBuaY0mwGdGWt69dlw9iN/pUyoSNupFsK
s64l0sgSuBWk9qA/QiBx3yVOO+lp7dO5IQEPxO+Sy5J2wVDU9sIQFrydsqet
ZAnjcXpVtfieBY9SqqPzihoJlkHX04rVQl0rNIlJYFEXFZUFJ0wYjqpd0sx3
0TyQB1/KIqOoeylletbXjphm0G2j+gDw6w8IN5UXMojq7DfSaAdPsCD8fCg3
Hyv7tNi1cefeDkMe9m5BybOw3F/1oOS3Qxn1QlX0lkN6sqByi3NPt/aVHQpB
em2ceq6eQaOsG2FQKQ+PRJFIJa5xnvRum5sbDENE7hvW/Y9fSKbch+JOtKHX
YoxPpw8fgLlBGja65HkuhsIP1kxGrT9zU+yn7jmKYgsWaGGu2U4dLt52k7nv
KhHJUE6dOEnIRIjMzltQb+IL8ZgSwSFkbyyuzC8SyQxFggD8Vhu8lxaneYIA
6W/Yx65vjYKEv/PqVirA37B8sxs7ADVIpQuJecDAiLXlpGQxIP+Bh9PFadbn
AoR5YSxj1/C4Cn1YlYsfqrAUzjmYAUbTuUyLr+PUEaekgZAtnIcZevO3K6od
S47Yn4mKfpDU48lyczXhzQS7GuWppXTXAXtKkv5hBqAh3O+QMaD0sywwfFOs
l/Y8mlAdTRJMqfaHUFsTdXp9Pn1X/Ov4cB+gcBvDqHRS5kss8jOSFR2iwYXF
zjRe0zMqkkNEsDWAXu7Qej3Y2H081g2XA5RvOiN8KLK1bfF+ITCEVWkb8G3R
cvgOLaBipiGHHUx4x+/4zplRIwPRQ0Zjwu8+0QlUv8pkXBAIDW2fssfpY/C6
x9rpPZern+JqWd2Kxzvxgto9El7I38ldmEzsOhSCCojqJHLDzY78b9UZEmB5
q8Zf36ZiHkhYCe02FTklsJdinzrVCR5xny4iKQuEniEYoju60gglZkkMkkSP
wF3PKghI5cYf7FiLh93rVbuVK9BqIqui3/9kcbLJ+bxi1uQAxh9YUbm4gfed
P70Qe2SAjZAj5I+FL+gRPD+NRiez83BWt+MaRAyBk0gRCbiuW3Z1XlG5huWw
cGNJRGTP/Hh53ypMaDb6iuOVqgXqBBFTgi5Uh8vY5/yWqtvXBhrm8jmY2BhY
eue/1nbohveGhd7yx77Ebj1cQiPjaxyLadatXqf9tfj78b8LzoWvSjZcJMKR
N5nCZAS82C9tFlF4kchoxf6xrPbw3lPXoZ2qUfpkKCl9htLcduT4QYJKYeiC
B3p3iMTjKc27DHgerEwrujyf/UyWGZuV6EmQu2WYa5uulLCQzh+qxqquzOVk
mfDm+cVyazKTofSft8H2U40ijIcqdqPGxOroLTUJ+4JEFfIFq2jKtRYb8D3Z
NcR4fkJlwcpRJRAW0SQNuUOGUuID1wdPeNmogpq6TOJd1kmaXKsLyloxha+8
Dm0gy/DEdWI5brKNqHD6aCa5vlJdkr707lgiQ/8JMfJNlc1sk/8pWrSUFAx7
2m017fmchMJuKLZ3JPJsF4ZrdFWehdHnGuHa0saOWNYgTrWMF9H26a2oa8kW
V2vnrjwvekG2aZXHlaGO5oJgMkPcSmsLdKhmtNQZYYZYdTTITuvgwJTIqttn
XUUDxcfiHefhu7hISNoSWzWipkdYzb7DH6dh0JRy5+G616x3dnHJe0+7a+bp
pCQfrZLXUOBURJlGS3IwP24gsEgCzopajHC1ODEnDi80us2Gd0ySNhZt51vp
oanvB8FNqI4bNoRi1MMzi/amzgadEc8qxmU/FHYRyVBrVWv1MZ1rtOEyYefM
UHhc3GH0/dCo3ANQ57hi4X+KODCUrGeQl4ep/CIwNPESLgz3sgq4kjgCdMfZ
HelVZDnscxezKN3a5QS8W8Pjjzt8XuH85/A3HuY4eImI0maJCXgUQ+WLXRdo
oFbumAvq2m8EGvEyycVji18e8GHgtN3Wlpp4GEr59uacL7uox57VeBNT/5Bx
bvA+Zy14Jmt8x418872lfAO+PiXPpAHmQ5CQQdlpqokm/ZtO1CLsjiBShvkj
Qo/RiZtaa3SIdmCo8rNUbah0m4H1b6a+VHSGxt+bhURZLcQJgUN0w3Uoq5We
YZRf4+r0Tc3R3DV4RPgHwdTSbdHJeISP8UjwD4bvwqWCNQR9tlxM3vxY6WXT
uQdewfsWdI8Rh22FTP4oOewo0KPjTID94p0RCaOwhMEqwG3FMiSSrk+IV0EY
ax5vRn3WGD4ek5Uo1p4OyKVBpecgTh29dYj9XG06Xw6DY/M4p6ytvbmc9T+7
iprva47Ye8STdN0zWYp/L6DKmv9P4i1q1dHkydk47/TBxBbDGK5vcomc2ChG
cRRyvPl5783Bc5wIL7hvJmLmkmQfye8zCyDi6ALWtjTlfIJ1oEn/OfgwrVkL
j857OEkyzt9B1OfkxQ7GsZBFuPBhG6fb0UNM96G9VjNnwi0qFAlnrjTb2eMy
ZSoKZ+oCeVuHNBzoFF8KsZoLxqXgg7wiODdc0+pxajuqYQ0GllyAowlb/nTk
mIPPxDakhJ/s5OdUqOpyIXzyxxzpxmNKxKRYmPNUicwQ2CL7Z8+p96JJOQFo
G4xca/DNf24O7D/PtuFAMKLhOpAio9EMZRjJQdXv6yuma5N3OZsPkiHfYI+m
HiN/xQ1cFbb/fwpUGYhB6rSHzAC2oRfmS44eu//S8CIHx97xtpbMInX8CzoQ
JA/xzrtvFIIy1rzzsUSvO/kWQti/hH2BgBGSmatjoTPQpBab5SR8Zbu2ffs1
/TQSh4EmXRTdzEvYVV3A5erwWC5B74EFLns4RqFu+BuAi71zAE6+OCBZszdZ
bU/ldI9venFL0RMUJodLLMnTXWo8/ljgrXgT11oeoz8shSWLnmbpkm62MAaK
0BLPMVPmNnaZtLg9HPKeimhpKV6Hprt4F11zlmz+ybyXuTOJDO+2Gjmn+BZv
p8x4Q24i9ITEQnTsIcKLw/8OAGmSMo0n0coDWlwIJjWNpIM2w8WQ6e3R9Fx5
PT2FO55XKGkPOs86WxT98BkIxRcf8Al9AFvND6vpcCECCYBQrBHUIetcmsGf
2Su1Hxj0TCTeog+il7mPxk7m5KRmddhh6UgC3xiM9R9dbgU0luFE0xxNeC3A
IDsV18RgNsLfUyVX93OGlxoDgEd+0pBx2hHY8/ocIz1ZfLVx18qGcS15toii
RXO5UlQ3vbH5DmeIyZqeX0WdXrrQiE0n2MQrHVN8FsaYwxMYjqf5kcsgexeB
b0qWBHhYiCcpvmM4C2hO8bbjZo1L3KSBZsKQFSArTsjO3wHjMLCGJa0RfsKK
kAaamqb2e5a4yUyPbedjAxHNueyT4G/672rypZC3akwzDteiXwnT/uDrpCvE
mSnpWHhI/8xaRQpNMon0/ggnsgMnvuRODfBZNlb0a5nif2wXl/37uY5LH3r7
3CJ2O9xU8KeQGHEt8gwgjRqAAAk4wrJAgwiDdilleMw+8omItnrSI6GAaod3
fUaERW2uabnX1o+eidw/DWhv1H/iW8L7lIn9p3UIn35VoeFKboZDyM+ojzi9
a3A4PZx9xiTtDG3iEklxwoiTMzj4lt6BZaL28MWl7uoRpJDtXPPV10BG3ihj
X6KIxIb2AHgMI0+m2lSzYg6byai9J0MnXT5Q/5nWMKVWF7E6P7Jfl4/RU3//
3wcK1GrI4PAzqSrE1p3+nylMlvifdnGfbZRkD/bbqIA4Bl8deXFqx8U+ZJQS
IxbMjtKx6QPX4TqWmqqd26dMuoOrw28QWsjyCU34Scv8r8Btv3h59wi9ahn7
BYPisPX2ab+2dyOf1qmFabGrMNDYoXluPlRyzbXBwquxfajVZveKzZFqZ+GI
GiEuUt2Cfuv+AJKrBQcMr5t2/UqLshQVCH3tbRS5MPTdmqJ5m9sdtGKO2N6S
Hv27VDAnmOQc8nlyrU0ijoBU9ne9eHbTmIIJVgUo2HfPXy1i6Mnrc4isW37k
QHsjMnzxFG9NJrWc9cLpkmZ9PeB1VqZfbKEU0YySE6wHZJLUtkwdu2OE+9p7
NMMb2t78cn0yI25fL+tqYzR4C3VYLb0Q8kLbHCs+zSkrzLVfRmnnyph7PnJi
otkOsp0MrFBJOsp+YdxAL+WafEbwa1+rGlK0P0Fb6PC+ZOX7XggJclWv1UJy
E06+vbM8tHm7+apr/x9tWbq0IqTGlD5Tvyk4Uq11YRiHsAaW/nahPNLu43WA
16n3BzYHPgrrLGd3CREr/kJ0zNyTpTJnetxK9DuQImOG9P1ye9uMY7NbV3aG
deQXP8Pv7KtqnEGaY8t6NIoR5+W4DATVbDgFYn3YUXQvv12FEshWhJ5KVsRK
D6FGqMxzwfpAS0G5BcavupeA81lk+HUdg+3kAV91EUR9uhJGY78xrC6YGgn6
2ZQStZhhbRuK3Laly6V3uPSlooXlxyFrpDAv6WogkP/oAaabyC4mp9GUFYDJ
i9Qd5nO9yjy2j+Kffz4NGz6KOsMl2YwwuanQ9FfFLxG1HuivlfCleIt3kzHe
LxCe8c5MjzEM0svpXQABMF6G2OlysnG/ND3sYfJ3/xUw4EQ2X6DSE8O4v01N
HYwshd/MRzXwxGUd4ml6+qqnN6OZXroqrBFJqEuuFJyidmeVIf1HKQmc4zm7
q4ZQxnVDSzFsuoI9XIX7K05dz0QnfVHnqpzAwNEZFuO69xffz/YewHutCLl5
N18LIKAafH32Jz2TGDmrwRl3QuMixtuBjeXrjmjbZcDwnApAPMYHwQ+Xah4x
5KlHOlQk0grvXOzNLfAr/GpI1bc7BjlwK61Mhhy+sc7kWof/zD0zy4iGXpaH
MpCyqWF56/8+GlTvhBMM2hr3IGxqMJTSXQPNQ2PZ5uoqEh5FeKa76rwDD31n
yrktrpemy2sq7X7tL1NN5S77JhmlVkcDa3LrC8oi4wRME3fNicR0HLAx+nmh
T3/p2WdjwqJKhoiYUgVfFIuIANS4FFNL88u0hBWzMut9Yfwy4p5BtaDkoyHW
FID+FodMFmHaFl/8f6kNExp9nGhtTPIgB6d0AFhMPSDpj3AvMHiMr3GWpj/f
XYOARIkOPw+R3EgGqrObPxxuITVQJC0zVX2ldTXUGGMTeSNp4Rtl3BU7hyDM
gclbeky5RNUXTyBGcd0U+ge52rVSEgIHKl8wQ1DJvVenVSL9lSXU/aG2/t+9
Fy7ZKFk/8F4Fxp9xS9//wBgalpuC/HRXQs+syR0nVVHrLNTLaxMzj0C1xaxS
N510dHVbjvHjikTRQMQK95kk4Jwv1u+LZSzZU+jhlqHejdtrh7y1o1aItPg4
aFFyyQeIv7wMB/85cVy7mbYS/1SUlRYM+KYs5eo/+ImRYJoVJFcCxKmj+Nap
so+u01kwT8LCdbym+em7gAL9J6WizHhskQfXE18xCsz5ImgiFISiKct7EfWk
0AWhb2dXkRkhqMwDqlSnGWwE7ve0Irv6h7NQeLmtbmWvf/f9K9F7GD79cOYF
eRZzUC3ZNON8LguvmQJ//Kqz+Z4ty2E56sdPk5GJ+fkIcDQHUjVnBkdyfuck
zbL3htNplT59MpKpBtDm+h3/fgE2RYBIDq1jHZ+TaEICl7OBNPsPCjv9s3fS
p0WpYQizrTaZICw5jxMM/+j0pq8QOyWjeR4G71JitySxvBTRI3mW4jtHKf0a
e4c5XGrlaHj9iDnlyMej4MkKzPZ6taOUiF81eM4fHhh8KOjbxOKP/dEhbiiV
o7UvEkgosw4h89Xn7Uei0ZKjwU4MdgpDxkPTeYo6jNPMtGMKZMqZq7mzvpOu
6cPAg+NVE5UbSiAy+yyETb96hQqsZW2qnsyppx9m38dLj4Lmz/UN8pfPuOwG
6yuSEclkKZMyY7dlzam0ZecB+clbgf88MTq0wbuHjixBO8IIk8JSdrYPGUVv
C2qumU2/yMDigM3OQ+0Tiu7Ql1Iget+iBBYekPDvzgHS7A98pvysmVSYe0Ts
2jlhRDhK3ZiRap1hsPr/z/Sxqh9LinkX1nJcXGY8kZsokSsAW+rNEKlLEGNV
HnGUmAWDHk4nKNCwaNXXsCZcPy2iIkg2sUsYiAFG3Hbt2D9G6f3owFA0HYse
SrM5YFKbniU73wVwIr5Pr7b0CxzPjSjC5q1gLBZTZgywDQBGW8ZYV53uXtdF
bu8tjo8VWiUXLt4DCYYTPF5gWPUvGYERM+ZIJBjGSoClleirSNCdHnDRCh8l
lrzQ96H4u/2mRROJKnhtNKlxnkyDdeO8vZE896F2BZ5z7O+WFuCi7hBSSp+X
h+6v3zcqbxOJ1Ta/ZO3QZv7G0gR8QURzWeAB1I2dU6Ck7yB5q5eVYBhzVmOr
JSfWKbuN1zsWLXPfJV4JoVo3vRJlsrp0lSeBnsEb7TSbjcrSTxKfQlH2XxtF
3st/meoGxe6IB2xH2fAgiJzJf/OuNZ6m2XxfgGz2Ecg0LoZ+YM5oFw1TVvuM
szQzEHHUGfPyZH7Gjpr3PhUGjgyadqVnGFfHGeZxIED8U0pbyQq1G7ZsPz9u
41mD2pcA3ekjUIlOql8/qlWVjAnxGwZfAy/QYsIQwpBN6WAP2w30WmcZ/6Rb
OfRqu0Q02r2pXODmIV9P6+9FsOcpoLDUIimnRtNyUtRKHB15AOj0DDklVZKm
AXM9DUdyzy4zWRnuleKawKayA/I5gjtubFnUI9Rc3+0AjE620Yb7J2A3WZcn
CwEHJgoCjoOQST2UthjE4aQIzxEq1ZOX38vCUm48Fd87wBCJ2YGdpYyrywAV
YHr4s+sLeym0C9rANiKHaqJcpZOrQJBdr0EupAR1vW+c9XTLnqnpMLutoU7r
2sgoN2a8J6mtjTgrDIygp4cUERy4DyZX7AoQ6FX7jw8JNrB4QUtASSuK+LJg
554D4YuHhDuagsl3dcQopXM7uxYYG6IQBeYF/2iPAmqTj3vgDdHefpUtc5/g
Ts8voJV68VDeF/ePBXpw6vKA3RpA+wbrZ2thaPbX+MzihFWnKKJdS2C77utn
A4kgKRgf9LDYGzsGLaPfF05Nkeg50UPS7T6NxHb8dKCkzkwj7AoB/zHGMgKq
AdG9f9hea8ZvO0ELMxFUY7sSBPSu2uI/yPJKw6BeOTNKafy9FzVsQ97fcDb8
EES2mygPrB+9JkWYC0GwRfbW+HUEAPyLQvUBMS7XhLEX2WmVF4PNRcjOWe84
71seeEdIrFk9LrYPa+H/omaXvdn0sdPOW0R03boTY7kveHGCKYve3N7SrvUD
iVyRCRnBTIYxbW3kN7DkgQUnT96LE63nN3XbTz6ooM4KAdGLH5e3OnphE8N2
kD0veNZE1Y6PCnBwMnuLMt/2ec26ghBXrkdU5E9T62XtbEdtXoTXCDJIS1sk
LhwXl6YStNExU4c+Llf7/473qtlCU8it6Fmbw35VqO9E+FNdOw+XwXaHrjiF
/bMBlK04QjwpfpdpERgNZcB//XPFqiZXOvG7adRaQ7QOyT/+MW53DxgStWAO
qtv0rGnN+3Z0zZhjbZibHeaAGoN1LnHPw4PvT05GMaUvAtUFQU2WNU1WqO7d
m95QkBKMWpPt+MRJE44rn91/aReRDPx0K0ArekdbN0SZ3tlwsw/2TFrfN2VD
1Ze5HRFWrHrcO74Y36xpucmfws4rUHBW/mvWeLC9Mzhk9Y4OGGaKjBD52GS6
+VyOsd8dApntOs76aJRmkl8hDwMTs57enxHZXlUArvLCGjWOzgh0CmahGQ4d
/d6PaAPfOA+KcfKGvclJ388hLlR6DrGESls4C5q6M2gve9qRxUA35rDPKg9Q
QGmhFO2Ki9fmmiW45sx6XQcSm+5cTY+2NCFWY3MlDp1NJBaleguAMD/gwvbm
2pDhGGRZ6pP7Z4xX9wfWRD9TYj4hQ0neDDrKRv1Oi86us3bBuIuBz3QFrIYt
1Dxe+TIRk3kxuGauFDmem3uJKgCXYITqQX1QmuIcsiGI8Ep4lU7VX4wnkqet
Oebe+pFiIVZJtRq+lKSqmK6IT80gRHE6JTkv6phMlkhaDY2YqXNkFk9ZVwve
5obyilhOq0viFUHcBORdDviwDvcmrL8MWD203iZlsR6plzOPtQTGpR3oxdKq
zW+1XGBRVrUTk8L4T8BHV//T3g0QxU32XX0GjcM8XGZ27PYlcsTb4u4XbYHb
Szteewc4ok0AV/hv2Ng3fru1eS+1Qqzw5WJq3djTqqe2UBdy/JkWOUXQp3qx
ylkER8ldOahbJxsNiLgja5hIQNM8v3QXLL5To7KK0dm3Qx8FVwRFXF79W2BU
MFbBTqyENZ3PeSGUodEJO1THtsO6vHkeVDBN4cnId5j5FyqroN2t3DuvxTQQ
zBOdkDbyen4Yarq2yHYKM6gGXWrx0DKj3yeJUn/IIRjEeagosSPPQQtQ9xlk
4jBMSYs/c980cRA3476+SM3lm1+GYGfwsvp+Y0GaCmfKlaL5JVrnKC/nNTie
HpN+B9BYHHpWW5tOsBbKOHstYHr69T4J2hlcBA1btCcGLxCxhmyh2aNjunBU
ZYir6Mnvd7gNrS9RAHOCk/XiAAHsaB2wrfn/NmDU5RyL0JNi0xD1UJ3CuBmS
p5wCzrBFcfrdjJsEXVe2fxGFfzgQ9pNocB0hMwmto8ZNrbrqShExBCjbGfcm
M14yU1kZRhctnP8Cq0tRJK2ftmxgL5U6/wiBEfb/VDbU85y1VFUu7iW2kFQl
8ap4Zg74muBKWKyfh+2ngw6x73zc25xjpuS/lMTFdeOutfHWE6lXJ1Zk5ISh
b9nanoo0+u1eYNE1VRpUNFD3jQeumIG5o6kMrWv/XkAcDloz/HaUrUNXLI+R
4rNYZgHO0eJ7fB6gBLsMZ5lIwxE/vHRyYSc+UM+fXXUkmVtzqs65fl6c++9X
h75rDNiz6T6BaDzoo9Udul7Yq6s3wi/R9VRH6rM3/EsGoSTwz1rB/yomi0CB
HvSTZVHuNx3BaXtk1q8MXVG9rBqQQRt94CWXt+KqHnj74X0PG8cy+4JUSmTz
w6XwufSXO6WqBbg35I8aALm1h03FQccjh4BddtxO84qQs25wH1kASHW/LOSi
BjTUxBQwZorIAsrA+Y81uxud5x+UO7m8MstzbYuYh3tb84FxSZIJ3YFIDep2
Whq4yA9DsnRUBJmdvP8ImcwgCE7ZSti9s3wspX5tze7r1qWiEPytco9Cez98
YPA82ilDcfk8q0cWgizMPeeXZ8N0cg1gRkwj5LXQpbEGgY0GypTPgiQG4dLe
0NCyOwsgN6QKCpyLzEqsJr7j+EW3eczZmPAAp9syAACBzUojQ3QCWJjJnswm
I+qo+MZ3OppLe6d63iR0JddS6wYjuOqxYLUJEXKCoinyLrcCquI9j61Gxnjb
tgqqhditZhNYh1iIkFGElzcv44PmN0csHdB8mSR5pG/euqRgkAbMr+j9n2EF
nF81tds/BEsxeMX4X7q9bUo0vQl0nERBRLJbVFD5uG86rKRdIdpM6UKU04m3
fYzNzY9ieBoT7MfOYIHL0LPFJyM4J9Dj0UzYsxzJtbT8K2uTfJ/EkGIsRLvt
IzbnkmOXzWvi3/TJnGEBKHyG+Bj7XkDznkLODLPzXxwKpOfm0+EcjLOl+ZWY
nYNZsZPMfWamXql6Abghzh7bP1TmO9DprWL9JkcrzfNgGLaq8n5SjWMTISn0
q2EdXqb3SovRjDdW9666YXWFc0G+X49Ji74zXJmdwZ78HlE1eLCMVXurSHmG
VmLbSbC8KfyEEnIm61jvAb4JvO6cUdQSlu7c2RtFhanYoTwOyeq81preIDvz
cpciFndVqI90o0YD5bh6dNq0Bt0yXKy1VQ11zvPwcad/z8iadoRiqzJsY9fc
K2yZAtqRcqJWDPGjqsbi9SxzxR/aiHv+rdIXQSVRYAxvBR9MeZy91EgY7bjg
u6+gyC4PJlGYGPftYQ178qMmySYphmNhDrBY6C+dwuMJ6VxhgOEHjhcOGTmV
POC093Q9y/2bJsijlnJYNAEKvxF2/f8xDE7H5tu9SaWFIKixFbKCSJIoJBfx
83SGG7EBkkOO28m01SfShy5xDpPJ/iAJqiaMCyhVKkgI1bz8P02jD5C3pMXV
RspmkcJhbsIRGkbFmoTQdNfWoGDbdv5ljxvz7pmf7JSppJhOKBaukTawb0rU
7fs9OjZyoaUtFx7a7vTJsYxCf/3arOwE6KkV1ghaskrrd7Qj/YikREryKmxm
ksZFbLE4TPrbx3cz9mQT54bqqHcUDzefBDeWCgwHg4wkhFWbSAjJZ8sHqTBb
VBq6oF0YevPykZCuTIHCDTWr7ZC99JSSyLHGwCHxXrmGXiwPJQ1YcgpxtL4N
YdXCdOD6ntsqx6tbUvUNl6geYEEL1Zt0m1jbZqsN8sSfmuc/SQPxRNns5F3V
FXGlymxAxs0asC/jausG5suoRtqFjrDzG07Ow7BalG4n8VwZhdbUiKdqC+bH
lec1Yzf30h8w2j+4YGkFRrppifR40ckhFdVVTlJVEQe5EjU9XGHZFotkzTt/
Jpiwyb0piyqsroJmkY/cpqHdX0hQabk+Gf8Qn7HpH1XTa5Hjkgk0cc5/9T24
qNwmCz84O/q8kNgXQseEGyJqqK7G4jzTYrPT/OGcStHUsG1/MZv+a6tWAutm
y4CKkI5+0wfqk/Pp74WqYGToh6M6HWEUIQnjY7G1ZgdA83H5C6Z2FqbDCRh7
rE21oxH9yj3TZwaWagFb9mnSmJ2nOdTiN/ggRNQmFFDZ+Qesk7opvJ2dYJHd
f7LjD1q5QyBuz4vnchWxF9bkCF9n+OuDrZUoajp0r50SlIEFI70HSKU9qnN9
/zdKHUjJUDMStAQ2egHvpvZf398VUnzBBBgO4GuBYqn1wzcIFiJIBi8uadHs
OIJPhLkwyvoY+VlDCnqwK7EUpX5rL51JpMwPLI5Rr+DKRtCFp7wuM3cyggqZ
RRW3juczh5iqIU9muGLDzKFUsg8xHlGwgvoLbPil7ve37RZlfy3kntn681zK
X2INBoc/XVTGMW1VrvN8UikPfJqJc4Ip8ZI8xSBR4/DTRC4qjaECYGKjZlUh
AYDfEEeVFDGo0CYK2pMiPjinz61oCvtkrgyDmiE8kxwH29TYXmI7LpJUB16V
+2QpM/e/fWhIAXUO51StuCF9IGqcjkeThOc+umOlPdt5KZMQwLyRk2UY5GzX
Ign/GzBYXW621lgZDgYqT4dlUYI4fqnS22Uu90dFbqFiswfjnnWnKNMI6n5g
jv4dUG/MLF1CTMZLIHnxKEWMZ9SKi3d5WqSoBJluv+3qbcWEXdjrlUpwTgvb
lW4OryddigHqLZRxWYri1ivu7TNq2DkyDx1zurC1273nlsI7L2UqsclwY5/G
kYeVop2zbDEnOFiaF2mbufdBekL/ie06l86WiatQuB1NuSH/VPZXgYSLfd/T
dTbFGbLd6vfESBDWsz6ItNHEFQCdDRbCeygo3pulGIjzW7wzT1y3ZHUnWEjt
riSHHTaEjAU9yN79SWKeCG6+jnq9o7JU0ajfUq/mo2Sh7p3FOK30tygA2QBh
XWqbDc+NRnf24Qo4JqOUxSlvMt2mYx7CAJ6xff5/wtFeDqpenPDZsR86AME1
g9bqVHGkUig6FfvtjNGg+Zjzbvw3p3zrNhlOE9cA/RkJkZwXPwbxofHRYS7j
LEx8OhiL1ax1an2qO6yh32syosmgG9txh816/xemhOYFUpvB/j+6jzAWHk9B
/nvfYkK5pVgHV46utbgd7gMbamRYcGvBwr1vfuYnYEkcGpFG2eIHZJQFRNeQ
1Vd53XeEX5WEpZfHwOiPq3b3sUbMNCNSz9y6t/izHT10vJNPogjMcehMLq1d
sxAKA1CRc0gkTOdUattRcHTjJiXUl1Sc+WPzuiLzIqNNrhXvSLQVrLU6Z7vR
dfaCmf8oPKCiNH3XS07SgRZCiXFnMHrxiaRzkQJWSZXDVMDla8Kr+ZoNswFG
IuotcUTWmcwTrDRcs0CEUIuxvFr9We6jfZYplBPSwuWzW2BNvwCPND+ehnaf
4B+4ZoEIbOsB8+uekdnCnBWQD4zbJqkOgihC1ehprcPxQMojyEuqeHf+DfI6
7TL29nxqruHUmpV6KFXGFa5XUP04c+texiKxxT6YrS6m/BfKqKt2KZ3jqXd9
HOplJRu7n79B5KX5VMmJYWC1E/l66lQ6JSbeHq4Dkm8lF352lVqWWKIuSdBL
sL99Pf8qHj1cqN7PZo8I/REQZvbe2KwfPib2R/9Zr9hYavlZzpq2pG5qbUxo
dg/S8181pwvbe6/WUM8JR8aH+GAC6qLOVtEsT9+XQEm30tZUBnuG/1ChqGnd
iYZ7DnWJvtUkgr56AD486l7alwngT2Tb4WD1jJf9ZiPJekwDw4KHcnedaEVG
bpaJDPUOhBIGeNmT88IdXfJv0u6o2fKXAkNmdJEW8d9aosZkW3u55+p4Bswa
fTRc1uWrxwtSOMAAtc74NbnN93Hv9LF3xwfd+/R1AifhU5nhV8aN8sUZqFt9
tdl/YQavVafLDQ/q/inF0zXszShNDLF4XuzpaJL8pLjUDgGAtLiB7B6jxrlU
6qtLnKKJeKj22JI4yvnQaIQKa3yDLapQZyhGN9clEONZXHkd766/RR9xOcaZ
WbwgrVnXJvw5Q5KemSChzXtrQiYxiBCBMuabTF+R2rlnuQtRhPN28CGp/ns3
0gOhA41OvBB0R/9PFUy1nG5h9lWAKUQg8ablSoxB6IbbN5ZncBlFBqXwgeLH
oTmwI8VH4AJat+Tsu1UnYJNp/gN1uzjVJfay282YnIi/MqX0/l+q5iuTFohQ
qlgrXZ5UqkrBWKlrRum8lIHTplBDLLocAtU2a7HddWDQd3gdplOQk0HhOMuM
NMqHDtRfErwqLedKRwqLHaXWDwKTpYFvI1uFK+LFCtXG5DLzy+nX7ZD18N2E
Lpn3XZa2h4TwtUerDnGKi85RuW0QmUJTtbjpcF4R/jyo/Ih5AiivEGP6IQK+
q4RbIYCdKZtFTCbcWPnm9rGNZKO3SB3FvcHgDvrK8YCN/Spu5nEojuFcHQ5k
j/uabjIA9cW/b4CZ9ku6oHX+wgrd0xLryZCT0F/5rpRoisAJAaG9jnW7DdLj
+nlhEdEPK8ARr7/8QgM598MWCGqzlLNOCXI9ZQWRZ8y/YNx4G8godCnAI9q/
Me32K+vmgKFidC4Ny8lpdbz77UqM/YR41sHSFzRrvoTyMeWHs4/00tCG2xpw
ON/tjHjpy4CyJh3Dg1YskTJd7gev8H08onP3Faeay5CP6BUs6GPkpWooVirp
xFR9tfcAvnvxKi3GjYMjiJX2JHye3VwtPF6miMfBmofsf1CtKeiy+gRcTmKa
RnTjbD8TaRaafMbvGQfcXMQCO6no1yDkZVYj3cq2lPNNmHFGSrQ+j9iEQdvE
bB6Z+sVwFPzVmpWt7FF5zXd1xPHiqQLeDi2uItEupPa3NqIEd3FK//W7koat
lfsD3bHL44ydVlCZYW4sS2MPTu3CWG4Cgk1zPOSou832dwJyM3x42s+Xp7Ts
MzzQPYK17WBYyc3hH6Xwo09wGTzC15sAUUfa8s9tJd8lk4xVoIF1e4ymmrGf
WcrGQ0aTJ9vWbn9Cb8Se7TTROb9sAh67FRCW81WmxFEUs4LyDuaurDYWVMuF
lmwqhoCcJz1KM18g4JUd7Au5k1w1NJ0Xhz2Cx2vPknWOQgRxJRCMau7Vso82
7xLqs70u/W3uBO3G1FNeyDkJEU3ysMxSBX0VFxCXFSnPGPI/wJNdDBJKueLg
N3yYvO1/qyjowaphSg/mdzqR0e4h1SPPYHqRpPHD1GzsmPAB6uG0IADxjAie
grj5dLU/vJHV0SVnN6Wn43fatHLsMfq0TtTR90h+UjXjIKGGJUxlnO0G4WXc
cJ04HJyZSBcs3mh+Cn8REej4lg9CYNtEQpX+DZHjYzGXAov4576rtah6tkjU
v3zoKs9dZckTHQydH979LsNb4lhrMES8aw3maUMkJH3EMWof8XH5DRpDN3Ox
H2IRBOYtRQZbP43xkKCv57MamNqsc/TVGzxLNVB30MRzAhBC9T1tJfm13dWc
5TRRZTt4BzxwK0Kghbu7/VSPnu/tmfHtm/h58qzXuGjBtjZHEMv8ZdS8ktnE
xreSnj+SaI9WefLouG24VsBYBtddx1Jfm3r/B3KHj+BshZbg12oID0PvY2xc
b5BnOdDBg6nIJLL3ra0ISOawEfsCWrf6FlkvJJAL/n0NSe7/T/DKen67lbBQ
8X8MyJth7oVl2YD6ffKAXjOjWJglRUv+hXCpTC6UC8XK999G8vzfpAfgHLDJ
JZzLw8ye1j/cUvZ4qerfg24bE0wUBBrxtOm/OXtFjAmll2m10YkZs3lUumg+
rN8gMOv0YCU5lu/DaLC2Xb0X1aHb1y3idazmUPPgqvnboAAuRDCm4i736jCR
/PNaQUJqhTJ8GAa+AwrxirsxJVrYhOm07kCyd3pAFOMcgiPIRwOn0WtsV1Tq
/k32GHipLgFNj7QaRFHa9fnKn7mysbyIWGb8kxrUFPpBU7mfSDrZQ3enPYHL
ifqHhVZVjam2EYOw9zZi+n9y1mUHNyY4jW85azUemqRBLLYwoon8lvLGS1h4
OkV9vGUA4NyQqlz2d8FwVQf085temDw/49HLef5YVAHXYrkNi0XOBmmvjJKI
9uCNu2faOxyvq7pcqTRDduppJm6QjV3Cqiuvbt8J/C2x9ZZ8wgEkFObWHX0u
MFBIoTGiGiSNBdTZIfnqnCxd5z/Z8WFKaYN8nLB8UFKY2ozX92hkDXhBROxx
YhMdErER5725C4klBm31QzmIzjnTfB1vCLl/5aRRdwV5Kiph4ysg+ZTXLL+L
J9L81r0RMIEEcFva0H6UgTAYMtAcY3jMKDd+urElJMQK2WIDXbH455XIXk4k
9v0vdL3vmLb/F2XJcDH96v+EhzSA3qJvwzoODSOEL0d6+BF2iXom3Zdx1PBA
gBVY67Kcf70oJjn2g1UnKgYD9zHG3oeyJNy22j5ml+7WJwpzprBn+Ts+u0KR
zCAgQMK0wDQTnyWzdRnZYk5ObHCFRdHB5KpZRDpa0Mz650a+TTAxnOwyx9Ch
IvgA82sNx8U4DCeq8Kl4hehYoMBAVgD/vql8zkEyE4nuIg4DLFyNvi9Hf74o
b9dFcIQQA7n/cxEqhfRBYPOV9R9sx/oQ60ydsxhGBD+ZlR3HD59lekbXSkDI
iHUesMj7t+aoBhhmD782eTb5DZImnFidsM/TA8ERS+XD3NarkfMuZ542Ri/4
T33Ev5eSUCd9n6SwpHDDEwhOClpIQjdib66MPZZwlvbNHi8BJKlopf9BNWCK
U/PY3ONYMInyzsj1OyM9PvKzWPZWGx1Be4AosnRJyCjHiGpcGLV5u3yNKpfJ
A7/ZkbeYbvza+jTNMgkmJMcJq8D6n8PORSmvQGtbYCVybhqRctcoRb6+WWSf
hQKNo8ZLPl5S5TQwm/YfWRNrTRE+FsED6LKVBq5a/BbIwl+qzqnsBk+rpDml
76SRGQd5POqIZWYKqo8pEQmYw/OxeRyO6J4dQMskh2L88Kme93HfIwgf6AhT
Kw60keEiUT2M3WoK0KfME3rqIg6I5z0XNM8aE9mnecGs7bsXE8VyatD+7uwo
FeyL7OwUlMY0vWMX2ZF9GS8MVBi/r+sIWC8Z3PIymLt98WK2ojimjhu9NWQZ
619bsmY8//M3AirVrjyNvqsmygHXxcfRSqOMBggctwpaDYAgSt5TLJaniLcv
PyNmClBEYtR7i/Jp3/SG28RUzYsoK3DHEoacssYVq12rPzXb2bL47LKE/s75
POucShRjnBD9Ml493VLaY0I8ogS2RrF4qQ51hfp5bkExwubaSGsxU5ywR+sq
LKAaYl26y54DCP6mRPhakczdoZ/lIe0LYZ1R36npBg3R2jb3nOZgqUFwJXk4
uZCt6LNKBv61iTBu4lqbxNJv4217cBwus0PBjQqmy9uIHhcNpoR496Zc1smV
jANZs7q151Bfe9TvsTieCsHB8rSynLgdojooZw8Rgm7DspBm8JkHaONbSa3G
6sagpC4QR0qqzbaU55sqRXFbc3WHIl1e7w09D0O7XgXdFKMcJuROBV2qwRWN
KvTHhXyH2T9NAojl25JdTO34N3rf7lAtvztErcbMod2qLPPGFWVBxAelKGNp
7h/vMGSRJV3WJy0R0qUF0iXTl78gFQhgEAToau68DLd6syjPVMqnixv9Un0E
CDtRX8JElmwW2unw/7d+lqQCfqk4E/ugqZcoEUcWTF9TaLyXrMbVkuWcazR7
OMJjaf6KyhcoBK9w5EMQJPZV8mxXmMuaS6dZRZPr1FhFtab7BSXJCe8cLCQ+
wDTCmshT8eQKn3qsH6/soOIwV6V6g80GG1SKJyK+1liF1c7E2Xm2hTR9W5Is
OXstlAd+bzBhA1q6hlmgKp/3c+hQ0EiGEf8bgx5VY/v/sjKidapVb87MDxY0
Lnm9hvFjQ6PQOcxtC+VKFBq/81Zos/uwQEJWIsvWAqYebicrnG4dnwl6Ejtu
djmCFCcKT3zBADXotw4xIFXliwS//YWsZSF0UicnjMWJyhkM3PRqFO7ZEyDo
oUwvfcthC7lzs0YB+IKQP069NHYgGQhgvd9/+v7D8DxVWlfd5fzPTvqm20d9
JnYOLrHBUHBqIIT/nbxNDFKoMvqx0Z2aEKDt9w+EnDQizW660aLbqB4hkaKy
gRpyk0GrPRgK2taZ0hp5f3fIglCPduaGUxwpz0CNq3RpM72lF1/wy582V6rl
Niv1Gw+bbouB8JD5Oh3K5QvVyH5BoIFAqZ6udItBUCif+x9XYkVP8aB1I3x5
wk0J88eWJS2HZ4fpkxAsuSWrml0y/evoQ4Dbbyot1Mq01HC/HkjAi9wpHL4s
e/RUepZSPmy1K+numS2JJNjWAAG2t8wDMXrVTBja3YZL2Mvz+K2NV4MdKA4p
3c8er0OlHkZsq7JE9bPnEmi8PzbcHTqlgRFwMPjFP3Cyrht16vLBtpyEsY5v
geeJ4AeLUJH6RE9oRC/7jI+5xC+AmtgyLvmIYKqfWFkby9Yd/5U7K18SD5Gy
lAShe0V9TtVy+nTe8k4xxHxtrlzpRtH/brvPqm4OJ5zoHrzoyAeBYnLnnpVv
z/90eFMzlX8g3QpTg1wS8RINC20vOYA5CDkBUamF4wAVdfxULHF51u+0oAOF
QSmqQdU+4ge1zO1CSab1xnO4xHHM2Gm8Tob3XbhQi6Qs79W0Sd463Emzfdtf
fwfi8/ZNgvCjurvsDGa62OI6ynNgahQEzCmoWsENmUSTZXbOBGYRDGPGHZte
W5vnppkYDSC9CQsFvpjVeLoh8EUbRc7rwJnsZXldW0W7p/H3IT5uidAboyXG
hAnOUst2tnAOJDzyfD+ulGLeDfmmdHd0orNSnlpfjzD1rpMrNgz+R0mt2mjD
cFU8I/dmNLV/JZOekzLHiol5XdxvwxmteMv/TlkWx7RPLSftvM5+Ro43QA42
hvCbKhaa/QEOaRb7Zeo36X/IveSkvPolQg/DtlhESOEPz5z8WXv98UUVcCU+
vMm1g44A1deFg+kAPZR8BY4WFNKLjxE6wKOnc0vbBRm+IyHSwEjjddXRSe1Z
4nGb/spSN7dVS4hof4bToeQW7seQl2/2MNohcagrCa2ADJSs4PO8mia4m4CC
JdSJnWipz0p12JRn/Dkl00tVAAi5SrBBMxjCsRIW4NnoarOTZ2V3kCzrLZ95
POXQO37s1q0KdlRwOGVNOUOF5Z574FqKogTe0MuhtQrYKU5qfHEXl2eD4qTd
KWlOUpWHELotQsNFMwam2shgur2PYH4FfrWYZkXjtqBVPokcdw25k7Sj60JU
ozNi8p2NSdAAH1IGxs+xDFtRvwUogZNqkjLlaYecHNWY+NVjNuMpumatORwk
3QcHljmt0TjxmlqqpV15YTTEUHT+1CWqMRixnZRESxmNzzCsGb+T4Gay8AlJ
Ba7Y4nmB6uF83Pkl/C+k7EcvNantFMZ0v8v2ZN/zEqXURc6k/QIaqbRX/Dxv
GNDj8ednsoyd6gLdx9+3ecMHvEuHtmEKCsNxkCepOg3BQ8ILsAOCxjPSe0AN
PCEDOf47rzWPMfE1S8by7PaymBQVmW5DEtw0OUYdEsreLgFU83l2jddfiAZd
UMHT8bzvzDrxrLfbpsivzivoAbdBoo/0gw/AGMzFbXcefKPx4qY1B7/mBjak
OMx6gt1Eq/wgQzZqILd3ljDPtXKclXfB9zA6F66YTBMGPeSlnjsaoYGRQSHJ
fZ50rHd33ig2D5B02UayBWFUOMoc8hgxBnvccoctqgZVfPi9Fc+FqylfJ9/P
LQqkDDvotot8cf0OpQmKte38T8DP9HAw3IPSeR/pwAYzdQvLlTO88ouY5CJA
x4u22llIrtEs5WASqpXba0s3NzXe+b0Xt7aU6HIB+Vv47L0ihy50Op0ZONcE
82qWZJywKXIt3E8OeVyKCwWF/xyoycXmv2gYYf2YKsN4zJ79KcSPloNbvjpj
PE63D0hEPtkW89DGw3xgf5p3pCC5ACENQkf7nSxHyM0rf1l1Op55dnpenoGL
K60lOR6x8ny4g1SGU/nacf5AL9yBY/GEKeCkY9JeIr1TVpNQRuojn/DIlDPA
3dXdA4XvHRgyZVFNZljPiXHZqrSw1g0gpp+RB35HJyky5INrsDwhVwkcQbN9
0tdmY8Zb+LbKxMXUy7uNwxraFKbtmVHGoYhbBjLRfn56WGTfqLG4tq8fXj+p
n9IrIFjZDiv7qyDWd9f93a+viMBTunEYnCbUimdwMYc7O3+8OYezTqCIPQfC
3qho0me6SpBC1BClGW9zCdOAezkbs14OfUt65wkS+95rxA4NlELg01XHjVmr
qUtwLr0LPoAMB7FN03rgjovJ54K2V6XTXbfW5bFmuZHbiCt7qs/Jou1U1KQR
Gb2yXfmLgYjixfY7F2wRod2wJ70yOnouuj+imUYatKmN+P/dyl1yR8+6h65+
maTBd1x1QempWPb/PFYMVx/AsQ916mJhyH/qCFeuBb4QH7v1h4jUxe4HMlEG
7m+a69NFym8VFiohk7+DkXDs0rPHiXPWd59vCGu+3YVFNcmRl0hjrBdjiyg6
mAYN73OpDo4+SXeWns/bKs5hhGZgax9cUEuZvYC7jdcfu9+0+9MrAaP8cxS2
HT0fNCGS9ujXDkFSC8KVXlQFLXgPCNstadvM9guQdq659BPvNZqLWZS+mCe+
wqVAiwfw52356OWkXZyFhwb7i3088sI+NuuvfzdIuSS6l/PhY1FoerUPp0By
un0tTdpr5VaPISdf5or4VJtgKZ4jqkweL4i8bRlEm3/m9Tu6zHSYKrxs0q2u
99HSfMVY5EMukOwTkT6swLDiXdGBQK1OfWcYbrhsRkGEKk3kf2a766N4si80
FOstQTaipYFZnjezooCjJukiteDv6VUpkLOryy+X+DKLwKyZCSii5QCjv+42
wVgd5E7Z7ZXm6e4Q9mFYPlzaZdXg3dwRtURkL9zEBVDJjtVjGB7ZVmaS9sJK
UTm/FlmJ2RB7+C9xR3hEd3uuMzvGj5mnajvZOwBfaREJ22+1ddZnxRfa1aut
BP9tkP6kXo8vD1D5OXM7eg3lkTz0f9Jrcqq14RE7bXfeIyCd2IraknqK9io8
2ukewisKOlcadUO+ktxcnypeTD/qGfMUwgfP9PwsKSMB+8fSiKeHyWdc3WQs
k7JwtOECvFgB/F0nZ3FvomIy3C811BGiQHQZn8+nwq82BfxqTzKhfa7Io/2b
TgG9aKGBdpuq1WGq38inZ3dNRNODS3vw16MifQaRQ9IukbyuJM0QlJNltnOg
oQtLzmnLq7bIrAcSOjFb8j8HC6n6iMcad/9nL0WCujtlHl8PhrmothKQwr2G
bwHFr8Ek34uX9XCXkKRhMmlKMXLd9ha/RWazFzitlZa6TiM1Ug4+fckSL3e5
XWA7tczvsoiidzAy8y719sSdH0xzaJiuz0JdilrqkKHFHMcx7qw3lkP/pL7R
MNBmx10VQMEEB5zjOYsRMqmbbhjK8w7uZEOGc+n90TK3HbJVrbC1uLYteHR/
7yybdUbLxt41gsE89gGCq3CwBzfsUK4yYPUz5yWF5/tkTfYGBNkkWRBTBbop
1QKe+04nWWM0Ndsyy1KNoLbyDp8gcJZGhJHdKjO2pKQZqZEl1pdEE9Nf1hiO
mBWdbjOTjXih4l+ZsIfyzkutxbLcZs3Tqm7tS9D8yDXP8hEsWvG1Roo7P7hC
mtsgKvrZIXkkm+ujjkYwBQeTjyrOOhUO/tWHsFor48TPMzfuNq7FUV+wgnMj
xk0tVNuRdYdxadVnmxtKVpvvzHi3rqGCHpLlM9iDfz8jwr4KUqrehcnadxq2
zy/gf2D2mMcZwob8qEs+eEsr156gMIREhitvNUNRyEcDu8sV0IHCp7Kwdb3F
ox229wcgHbC5AADkUEVMkQ10HLMkxNqcG3cSVwvjgwduHiqUq2cEk1PBGCLE
QuBhbCQqIhN8ZNH0nNvZdAwEpYMej4BcN4wkChjp2Isq/ekmij7rRgNBCGDg
GqgjoEb2x0zBlHfn8HU9qCxL2qfU9KR8z5RLmvNy0Nl41a6LxF0VQnSscNE7
0ZRS/BOgIX5pD+z4VRVSFXzf6JOKKuWPyOfc1WXsxBj4jW4dOmKAucMsqTUY
XvgKs9qvjNvMpR87bq0ZeoyI2ou5FJKppCBSZGNdL/F252TmWfiiPV+t62Lm
4kIGWX0OcHKc2d5EZcgVvl8Ju+lT/mHqLFIJkg5UGXuAws0vk5SeqC9u0hhF
8/uwGPxEqYgJ7LmoN34Q/b5RSTAI2XAeZV4OB86RQhe4gPIW1PRxc7K3G5iE
gKkjBvdGX5vLNDF16JdTRQmrLHWOSiUCJOFrWuX2h1wsKgn0CjvP7pLmbaxE
Xe3TmRLSgs3xEZ9+OnfUhrBjjfRaJvseAKF2F82m3uwJJWBBrYCEVBk7Ho+b
ws3YkBK7/7C3myDAULmgDnu30PAwTpf2owXdRZKr2v8u/5ZvEqexBhmjYpKl
IJo0Udf5PEF0MJHdgD5xi5oOWJACOSddT1Noph4X6ey9y9s091sqx44YjSFE
Lgadnr16TpuLjUHLngS9HXFXdlqhgZLF2Flt62LJMNZ3NmfM/4RcXsM3kxO+
acDUuWhA0RGoGqUh6V1ulgk3ZtUX5aDOByk7SXT+mUTCxyNZX5NscoxWGoyb
7SEKEBHv8woT2YWWeErUe7/bqDoISDZb5kmgZMQckji98mN2l+7oQv2/R/tg
jYJYNUH9CXdM+dlnEvJQ+Cu89mhuD8dYfGdz6jbEL6/VRYW8O5BSO233f2Am
ym3CIL44TH3dsps9dFLAwRtq6pPOp2BjfV54Sbk/pi23XIFnHlfgps8G2Yz1
cyqPbYQ73jM00nCAIogda3oTUUFxDUHRpoz6TyHMrJfGh/TC3+EwQnq9NAcp
c2trQokl46Vp+mWYYYkZKuF6s4F8CUU1OvYtYRkl09H+2LaOjIlivkUW7Srn
sj7HmD+fSN3DoQ2W89z0up0BYA9XM6sYO2VkuNUgiuFoUTEAj6BL6vtyI0bo
ar1wL71qAeATDQBBAnwmc8z5+dMDwYEgF4dcCSDs+WRC8CiaN91enHS/kmRz
LFzwWRW5fGjsBGNp8oFuMpjc4BCYw8t3qmi9CM6suTV9ipojCgScc+S2mcnv
7+vmL9Y7prvd88fb6jDPGBqqiDTjOKzzu8TbIqi0nvZI4UojPoVRMO57562y
qdJCG2q/+z7332BrVpaHYwfXugvNvJlnNIStKUjT9J4t0j3472G3yvzq9Xhe
nDAVfQHouRhrQNgGZzRazzPTbXdCToBXO3qPmNE5wziPXhBO/nYIiX9vXgUf
NC5GSaOMZlHZf3UXWsIV0rPP9wyu/Nc0ZiTJsl9zDGw9D2i5fU1PSySLdDxo
M8RjXaSEgR4/KaNtlrqqaQ26kLcgbjSzQM1Vbz7l5NtbXeJOJEMg7Q5EOubf
b28iDedLj8OY0kzK5G3x8r2f+vI0qlAhCZ4eOoS7h1d9s+8NAgSPsJh6p1ss
4YEUSvZWQze4TfSF8gmPQM6Aiy2fKJmS6qXL8OY/bsqeVbBMmGxf6jWoyPYO
B4sjr3knNu6QGClx8xYJXbgZXUINdVclLwOZlFfo0Sekofbgtqz3YbRPdkjV
lP5ZF2myYagQ2l+TIsVu1iFiaDoo3FF6bt/XdzpRzjmlkCdON+D5VkclX/ln
pStEVlnjibvRkjBVk5S8fTSkJqr94e8il8vDfMv69ZXOdmLdGgprbZcBI483
EPjjdYzWg7x8uHbP17tRD/ssnlPyDIwNO31MmzTsw/88erM9xqmnBCus2s5z
gF1nkytaE53fpzQ/+8x6F4xTYdhYMvRjyOS2qMnwtcBTuDKO3331wCpmqaNB
1eJ94Odi+97L2wWW7VW46HIMmHCgVXY9vPUPyghr/ZObIm8ZbEAOxZp8iJZH
ELapI1DFcMEOqUHuIMK5oAQ9nDRXiUggVGKbKDBK8ZWcme2IyG8WHK1wugrv
0volLUqV9EA8YAq22WQhlKOVbcup+eUuOyOl8a0Tl5fCi1AyL4wVkC8+C9lK
U3fm6/Y5qwWUV42WFmCn06gCd7D3a7IVhGq5lfV13sgeAUlhgMXY0TQOTXIC
2r8RUbMjRQnNA/v5ObzPkHQiXKqvCVnCveSjEiP7eQKocrsyrRB4trphJ9as
qtTlJ7HdL0I57Grxh0Fm0Q6v7nJ7TMs8CjRbhLh+J7j1NjRVDvZ15vjO3/h4
Y7QkYLykk5fFYPzkgfMAAtL3fDKO0ZN5KrJ/hAMDPL0jc1enbLO4yKchkQTs
DTcRwaecM8s7xEH0mfK/Lm0F+heTScZjDnlaar9TJ90HAUtLduC9vSm3FiMy
0G+2HCYIlg8lYRgMuL95k5B360LFs+n/LBt1jCltna/qqeLgEPmX05eOIzV9
HAjI5+GihulOzDw+xaubDASvMuNc4MRRg1/dVYTErXfsOP4pyPrKISehFbVK
H3b7B1da0PCDre5hYmAIIIBdoaX4+4ylThxTavnQcglKuAU5npaVEH3ZpxuV
mDZlWndZsvvI+q9nR2dlmcsB/SshuvckHc+seZyFMmdP55/Qnu890RgwsJaY
TYYfpbiXeTv/LB9blFPyIolLMHULc2KIzx4yav83u0hWlhVJV+fPX/yOgBoG
5q1x8nugCXKUHI7iH1/MSSInzls7rugFMKkFeQtrEKDjh/hMokOi3RyC22+M
ZsezFoQSOr+r801eLqBRB81Tbov/S/6Ns79Y7+FxWQ5bGudBGGrJtFo+Vqtz
lQu2o5fY1f0OAzNP0ImkdtddVwE5/zP+uFAb42JLkbNsz19aNVoNl1SFJvWU
bKpSIrVVHsVi1cb90TTS/vTIwDnUb42XTkGIPDj4gc9p89YoS/wEpejsc2Qt
thrgVNVmT1AoBPBgFeJsQxl3VYL8z77PnIsFoB+BFu5g668nyBUyDSrYKbFt
c1dy16SfSwve4URQPrOnrFQsjPIsLR7O9YaVqWVGJAbrpewz7/XiXurtMWkX
ofwIWIbSu19f2C63hNi/Z/ZzzYzJ8847ibk3GFt1QxxTdywY2a2h/dgLGHME
QLoiwZ51vbcGlQWWRlp+96hNjYSwHInoCFPpuyjtBEoHfR3tdBjQweOLnsEt
W6hMG+mDb+MFVK1nhXNcmFtaBfrPQ493IAA+GV6ap64CKlCeTnqZ9ZGszoMs
IHEjVQmtuJwtv4wsuGWgemxY64fb+H21zv0kdwOc/coUg7KRs4f0i/yDUIBM
pDV3gSDbScAQFLup62Z3GjTmfk9FVcsVmN2JoSRszZJsVo1t2KyNAm0JHlgW
CqPutiLtvrGGraqqrljVKDqm7DLA8mw1v/T5GWUYPwBYA9xewgA2R4fhqyte
NKBdw+khJC9lshmCCn8JKPIapNSLlf5PneGit3H7z5wROqaodoCp0mzuAX12
HJGvaWm7uL9p+wNYSaFzbRPQ56sSUNuY4Z/nH2Zk1jqS3Z1CpZM+Nf45wqfG
0fq2U/wQ2Xa4kkN3Cn++vHELpuD1KVRSpB/cTPI5cNgBrU9Nd7yfQbMBRxtp
V2BXPtmD62l4GBhe9OXOjJoXS+dGBxh0r9oWw1ByIxcOj+bip4iH/0WN4ilx
FGu/JgvXKRQJIZ0UahqYhRr36+YhcW/0qks7TCS2A0Egdi4XrSffS5Z/UMP3
6mLrwcHJhbv2T+2GPFKN1RM6a7fU1m4sneDiJaUgoFmogWU3y8Vls/6WLuCE
baW6/sxJDGFM+fQSPJT5ANib6aJoAAMNzsFpVsQcsVg+dWByVUCmMjz/AeD3
B33+o88MAqpEyZ1WLQDuKiWrDfbCa8noT+uP/ki5glwsGLRokvwwitGfSJq0
w8CQVxfLWFiXRxubI4rjO8zlBcFbZ3G9bV/kdFIkwrdjzIwHGyNB6mzLEWkS
ogky8zggjvTe4Hz5zYVjZH+VOg/tCdo7/EFnBdftuvLhIJqGyYJjhPISIIrY
9BTLTBrCcK8UE9D2wk8MuQGBeJ1zLcIh3fvju0NOMYXpLaHof7dqFk3eVLx3
3bGyR4v7aESSGz1iqYNzsjYNLOwJSWyQIB2EIz+IZQQ+WD3hW76YKQNqm3Ns
O8kqoY4yGNW0N+YiTz8ZFCpK8VZ51r1sSXRq1EKmaitRZeTnuD1kH0YtuzS8
nt/lNwH8I8iismuyhLL9YlACWyF1e4ccF8tgRxt1PpvsMxv2rWEPSsQZDy3m
fbwIvE1qGAuQvqdK+aBTKM50fY6aTCI8CR16VIL4UTz2sv6sHZNEv0w1ah2T
iClo55dV991u2a2B525zT6jTi3zH+OrKEurIG4ktN8QS7WpG2A9vwBF5sPOq
zezBhuRb+8sF1vW4drNCD1+Cl3Lem7inYlvuPjzqGrKywrM9hA1LJiwUperi
OVjHCLwe7+ZeKD5IpgY53oIaasx8COlOG7Y5Mk3WAWmB4TFngOzk7RMfCEhG
vJFe3uBKZUbBxgRrBKLbP4SAtC4pfLhN5FbjORmQEAqWKguq0frjg2gECB/a
DdDhHNZhbIJrD1XrkM8hGvtNe+yU3owFD/XgfDAKe4wxCRwpGpBOos6CVFGV
Z+/BWhQrJtyYeHyn0M6DW+gOUc9RmArTZ10bn79wcAwK3Bvpe/DUKm9WbQdG
sZi+KrJ1o4K00TOlxNXZn9bT5cOcKcj+8Wc6ikxFIE5vg2mbbZ3xIbb1frEV
WVhC5DOqka+TgX3pQHGSZO2GpRD4nkYLnjOZuEQ0245AoQmmhsD7mrYR6j/P
3mMw3VP1yDAz/8zsPWECWejdhOs10LioirSmJMgvQ/BboO0o9USDbv8E1bvZ
BIRIo6UUvD5du6RqWne4K+PNR0vFoilKkcr7cPCwlxPa/2r0CJ5axHXwOHwJ
inHWFFkbZystAH8ndgaBOHMkfKHa8MoHb0IOjhrz8ruJOQ8b3jRqA1ybFSBM
/uFvuEeRcDAYP9B0dPCsHVwarMnsN7cNNM7wSO0VtgNLSuBDPt6eI3042cm1
jD8WPsdH3dQIQ9mz5QA8eHK2CR0spWKgSbEI0mh35Zgn4DCOLFZsBiH7mAex
VOVQYzb9cLZ1h9yu8yAr6SGqHQXxIjHcYcw55JlaFuffNR30YXC2tyDHgU8k
klaE1X/M47YP1ATX800K94ZaE7kXv+F38pqtOuz7f/w5xc2iWCZOz9DyMU/r
wBdbYZF/e7Dn9Id8cIGeQsWlQ+7fu/I0hKt+Mg6vmEFMkF3Gi29+xDAQUCtT
R+E/14UXkzdFC7QFL/JfNXx+MVuuSZmZeC8NQfV6O/a1ri+2MyE4IOUX8ZeE
/el5mDBP9uLTJjfOiv764IRwggUTTRcT7ohf6u9yhKoq7luC7kI32sNGVEZA
DNH/XWbuIwCmPeGHKPZykV7561lISSomFB8Fla8C5eyvyc1QUKAU9qVuVSLp
XaFQLZIhle2NBTOLAVvbOBbusqo7qxktp5LzNuBNjvKsCXrWl4fYJ+f0KEoA
yLhkBpPUmL3R51kM2RnyebpZU/6WWFiQw2qVxr7QCh1MSdPyWeMD9BGI6DiV
0xzghA0AJi1bASlnqgNDISNOSQ1eD+R4GRsPmL6naRVM8rS1T+6JpSuyb7wf
QjmYkfqqjUIj/nibR5AIqT36CfiOyaXG5PeJcy4fZwEfJ23HC9C5/ZftRMIj
ayfFOW0fqu3ffJAXaNTpz+5kVk6GOu6xERBJ3/bk/fpCrOtoXzhzPgg0FCi/
Zhm93rIydUojGaLbo9Q7pG4lTy68/ozhLmv0ddPmJ1fJVMivITCjVkE+9gnF
TUmDTFs8m1YKULIm8lHhJeQ7+CaV7zpXQUvQKTxqH1wnY0JLS9M8TZOSFg8l
IB7qU4+cFs8924kI+qK7UhcQUfFQL1/RMUhnGxWZ2gKWlv75MpXduoJsrg0y
f3SP253kgMERlMeGqsONdYosPt0t9nSd31UfzjVvQjV/+pfGtL5gWmfL0Gyo
dZs64DrPHwmnsuqUzZe2l+MKQQ73vdSrhW6OIw3KleF65LMzJYgiaVhDowDV
iqlFO1a6cmmMpPg3Gb+eYDJXB1f7i+iZoM4VX5h/mjg3iLYkSBvddRIWVTRg
CYPf799akRy0aQTupvGPNst573kBCuABOHikHUmrztFyBgDsoSd47fvb4CT6
LoODQ0hTVgTxihhuyLLIdvXsVaJgLwSMQVkNM4eW98unnc/4ZwdNXDTGCxyE
0+j2ufykJNWh5U3Z/IjBOETwkJeKf0aXYNDOWpUiQTwmAyRRvzgZda/ipBhW
Gp+uYJlh98D/EyMF4fZq05t3IF5eMsgtDk7MxTdSBRId/Rz4anIzJkesh6Z+
7yotrKlHzcbJBFYzuRdfefyHci334V/bofb574vIluUi0FJzykNg9gqtN4pq
/T17u7QFX7d9MtGeUPCywgkaV3pr4Tqz0cJgXj9b4iffV5iJb0sksn1pP3A4
QxzHKqIhclVHTZlXjXpo+yHUMyK39rrDC5QbvWyA33RVWQUdB5FGlXddyapt
iGXHASNFwNiZSR2F+r9lC3enxC0KIEhgd5rhZw5telEYcifKjqF495RdNcb3
G42uTYvYN6R88d6BkrmC+IvJZHqQvsq7e67M9EdyDNkS8bHG7oNQkb/s5Ip9
VnkprniaH9nb3v6ecwTr990ZFkKt/dtwo3yA68oigTTrGDeGcB4au44EGvYm
ZVq02KfQ/bRNaPpxatKOJ9fjy2IHEw2sDq7Hs3s+rWYZRnF7pChXJANcKko9
QdRzLWGnlhxsmJRWaBK0zY3Dekuaxe/a9WlOwSLEGwmPquOku+Q6RbouLTg5
n/4KBW0H530cziBIHOvFJLeTN57n6zdDvdK33tgV8qNRR1XBo+MfyLyVxS6I
OA3UyLT+yZwYuYagVOzVuq/zr788WpBhZ+Ex6RoTfVE4Dl8fV4EY3zOn0kwk
e+vbI7GNHBb0u0zvuE39g08aWevvz2a5GBLlsL03Wu0kp5qrS7FWVeyo9GKx
Avb0QBeQmGhc0xz74PpQueQrvV+WkXMx6jepHa838Wy5q0UpcGVXNQIwLlCT
jZE4APkfRhtzhz9rLSEq7uM6BmPoiewM/zNpV4oKoT/nKbXqH+pomo8kwbi/
7LsC99bhNZWNWL26MkCaZ+TdOE+n+3EktzAq/h6Nq38SjJJpcb1XPiCugxVd
orqZJWpxsXYf7u9uHsZDneR9rdagBP4MIbjj/bycF1UtUCZNp3IkWivp8R0V
+7pQ0q5jAm3pShD8VJ6tTe2DkK6vGVUGa7CqtCHVfdWnuPHCeXgJ9UgmkFK2
BGqnZ9qJLQh5H/xl4oIUH6lerQIxbZJGMmm6+RgLyDS/Ao3RElwANUidHoLu
odfKRAuqaD/eq6Z9dasNMoqzo+O0Y7ClqL561lRmjCZMmELrghcwP/cxTs6i
psPBUKBLe5bw9xIcqWzLzQBd3Rpg3onDKECAHV+3nmTUQQ1yJ/xY2FQA5HLH
ydjo62tLmcbKTlTPl/mmxg8DCm+pmasQL2cTqPgctoJ0zoeLd4vw7l0i+pO0
MNYyf40hmjpgakjUWsX/bssq6JKliRKw/VeIs/giQLr1tK2a8xstQ9Cz5Cy4
/phaqeKYIVnqhJEhnjttc3eCBvL5Pnu+0tK7OIPcCmPJfW35hXs5bGvzlUlD
cEg0R/mw/jVkhMdtdCDV1B7omHfU+gz/EQ8kLANypn+vhsi+rVoG3SUnnVeZ
DMvNoG1D+VNDD+rEGnq4irRhZLce8CIKLpTlnbkR8c7q4wlMHJwvck5x+A9E
DHqGnGK/PQqnRdxltErHMvBAkZ/SABmHZdtQys8xmfmr0RPb6tqC8k2PhB65
kX18w2BsgWgZvGnZ081V3bqufyIoNVJlvjGu1KdCNSwBLPZYXyGBJiw2BtG2
6fIyE4HdBzrubyUwC+b0Z/sRxjE++KAzSdsLkXBusC9SProB0jX9fEBGqsvE
W5Pp8kQqJcdIaQDbB+Yw4WsXjDvDMCf1tG6aTm8Kh6PwZFzBRmC8m3KO1QtG
h7FKVwd6e9zVIP1w/lNwwRUPhYuoaOPALd9Pvqvd4kn44sByVTjNwLIBaTWY
BUmJTvfof+JZ02BEigw2OJ8XYtpc1uaRpyu7TESmjmrMCGzvRXcHI2nZV2Uh
h9dVKHw6Rvc1/ZNTmNOsjb8025+qGLAwgaLTxQ1O77buqxW4tG6umehJ5GOL
Nh4l+8ekWsoa8aWQdO0c6klEViSXgSSFbFpfQGC2vNJ4/VP+oO0VJjHR/sXe
7bmatEEzpQMXGooqVna8AUs5m0eFIo3A7Y2Z05FB/F0vr4SRrXX2N6C2+qp5
RAiPymc2I1pLFi64Rs1dH+F/TJu1qwg+j3E6CopBlyfQVRy1xY9Uw2f5DL4X
Ohh5xNKv7OeLsgOxpVLU84CMI4BdgwXOXL9dj0lbHlPP/BVYrJIUEHLyJ+B/
8lbJHxnAHSqD6kYG+ulsWz8JAKYVOfwYNECIur/+jH3fEPvFoVHKLwm1hMgX
rrdPyqVmYs2fRXJSwZA6ldOR2fCrRDKP7wUTcQbMU2rPU5obvZWLGGjKXvxY
X3M56VBqcywU0xoSeGFitD5pY8nxKI6UaYa1eG9wkyE0hlKginLMlKF3EXoX
ajNKFg/RCHr52SBPotUcw1vgFU2lGtQeo43V4AaV7nd9WB6XDrPYe++u5eOm
fsm5Ds0aHHFjRsnJTgrt76hTvlPLjkHO0oso307IbagBbSYtGjo2BdKd4dev
aKc1rEui1gaaw+fVu3Kywod8HhOGsgUBoOJPq95CgozlwZLJBnxxdrgCwT3m
yNiwSe/QWU4BQxwt5R2GOIfy5o3FmQji7PcATKsGHRNaFS1mwZd83mLnk6X1
kEhdBeN0/imIn8Gen9t6BcUUcxQs0AvS3AQBMjGSaeo/XFPl7DnEymIGR6ok
BN/b+pw/27AncwQKGOMoih7urmE1kC5iM3b0HdQCniOJ/04Y9sFcjrFl/4GE
6ORm0/mJwzUmQLFy8c9l/YiSfyTZaw4CrzQxdCso483r6Hfp4QgZn8YpFKa5
xq3/3KFwUmckJnxyOjjHEjOJTRw8k3EfEhHDrHJD5+hES/5mbYY2/1s7WSJp
0mmj99OzwzC43NJJkIRvKU38TDxBPOZEpL+1wRwUq8NcBymPLtPZikT2MSFY
ikSfrwEd+sVs58sKLLiF8GR1eLajGvmrwj3QGfDl7s9kYFYrvuf5xvtZj3Pr
zfNE0bZxKF/pHdgszwHoFOgVIWxBAKLddzq497UwfhhDvTZ37Pre5x5BSGAK
Lm2vbd8qDBNpRPyrs+RcFDWWK0g0odXePFyuV0jFUsfD1mnNLY7amNr3rsoR
qlCRYqs+zE7uM9luj5kwkMylBg13hvwGxmjCCWv4PnQ5vtqc5Z1PnRJh3ryj
VnjdyTWI7BwDTm5SegMy/Zk9TWqZmIlmjLfcUxVuAJ+Xe1HFTmPQKZDwts86
a8ivs6VX6qfHnkXEekbVxGrlqjSdPnMiJRGAXdOoawHbtDAiihcPXuzcIwIk
LKsHaK0RwNypaS17VOfv6ZupIWn3rvhEtl7uYFUncO5cLMs0IkjjBZWuf2ax
+RPgrDx2/V7LaM5Dl2wVGTDxNbkq6hc3zPi0lRpfY7PGlbeAUgqWmC8JptPU
JjHXVTUfRj4ylLuCPUtgx0EUMQS2n02xN0O0uae0PUXHw7sdSALrUMnVGfRa
OS12nBqopDbr4v24r93TLw2lqVoPEAyvJTHwg1RwZRosFDGl1Mfo9uswu19A
ux0i2RazzIoRRIieq4Iio17/3LGuHkdGCo6ymnhSn2TmmViblfLqgcQb/DYr
3O7j3+Cpo7t5zCWLrQfCe0hecvGe9s1XwYje06Iqi7i1H28GXYp1CawKsAiD
raM+WzeKB2erllrXmnEt+87RX3AVx5JsBmdJr6kYz4gQPZ8/0aNbt9hHsg+x
YW6uC2zlFtLiMsmjyfMqNaP/O1M7Ompg7ddg/lXSeQKvRd2hZpzZiDWmNRYK
5osZh65dcI2rADwHEVqul7JRJvYyzoYvZM/+AJxLWpjSSiv/RQB8UATo7EDu
s5eOMpRiNDfMZQs3w/ZaDIna2kECwbq3Z1hmKup08Tbea+Etko601jB0E8qs
OJzO7jormp4Jtl7j8SdOnKqM7Wp9wBJbSFNPFQdltvTgS6OlBynrkEpKAfiB
JyJlETB6rQD0NeWU2TpOO8+Omwg7PL2GmFjsNLDwvUm3uRCP8R2L4n2nKYoF
ltAF9RXEyjjUpv2PjElIToV0FypLiAEdDBLEAtrGlDNEPstaxNKsb9CKwHRy
7gIFI7grkfZ1Y+C9P2T3J0hPV9/J9rtaGRfnx9BF47G6NG9F5nUlFT/UJlO5
y3yz467ms58IWWSPcdsr3sxbGt5xTUsXpKE/y8VNSS0+EZmd6PJx+KxicKvG
aclj+cfIzSY9YFFlXHXnRpFxs5HTVOeRWs6m1MxI2NEnYncmHJoErKcrwbLq
qTdXxncgVZc/mLa+hSmSH6KyVDhTXkWu1VE1ROPiTqZVb0+2cWCdV05NmUgC
dfRwCvdQff627R9qjWDnpcaXQ75pPRQ01MNtGezuNTVNJom1TEpY5owk2Fh7
1jIpMWWZLfnyaRF+Hjbveo1PVGVVviwb5DUN4/lvoIBwDYJw53dXrtVph7nT
C5Tivp1uCtIub8Y66otBcjIQ49k9xYWo9Ll8TkwVJdTE/jK4H5N70tZFIiQP
bC895veyK8uraCGvoS6AGxGBWLha9ZjDl1lLQsmXjZC2jn3H+gt2cZDICWWJ
39RRqso7rwmr3HO+Ey/NnfH5ZiZsGEG06LBYQUKg9PRwRnyZgMOeBe+cRD6E
qEkVoZihE+RjvC5g2dfmDrISwKWCnOIW0It46/mwV9EgqMqh8+RBP2DDRFv8
rZk2IW53v1mv1TMhuZiSXCf64vs7OMTT1efYlyxmTLd9MSNGl7oH3rqQ8xrf
So2JRnFkLz5VUKK99IPlaTX3Cx2r0u7T4wVXnsZugzghp5wClpX+Mk2CxmYr
jXwnoyIbq3+WnMDTzTw7ZvUiPLLqKddc60KgBMhIgXFCy/jFNDMVgrao10lM
Ged51dyyVEHOrMDza7RQ7/y0+2UkWF0WMUDLLeyi2iweub/GySgaSoRgmLWl
445JA+DqFm3FIUWmfkKSLt1Umz4ROHLA1svj6r5xlZycUsPiQMK+9ULzhHPz
Od7hxHQ2SwEtSMFOZTuA3S6sGrXyU3w3x6zFMhS0/wBPgJNMQ4m1Fgl1w6Vi
nCrCZfyrTmN52J7sQHt1EvaeLgOsFbJYLgTtkaCUOUTXetImNNOKRQPgicsp
Vpkso0v3fIqwh3qy+66S/hyh/U9UJ05AbFp6fkWtL5H+pggppGgb+HOxTKaL
raHfLqj0FTw8WtSLsE7+7uPQpK0ZKZyph0tGYZ1oCVoayIfUr3AKWHTTey+1
bN2kVtSdpWMlV1t2wf19GuHL6ccSuIJJNpEnJA40OmvRYFCp0v5T+gLy5qv4
EwUHMtMZiB3GxUXMKzba42/m6cBe03gAL7x3jS0Ya9bBUVl4sRtnXs7LDbK6
eDuz4ovbywAMnkWnHG3M2hJ5Mpr2WWvgnys4XXA0e6uVER+JHOBHOel2VPCn
ffkST0sLCXR5SwKe7rr/EwBcpd5vCaZsH674Ppwy9YFGxdSuEmXInTJZLEEC
TKGYgUVV62WT7E++vWIfni8uswSp1jSiA0/ktnHCXFQQKb1RrJezt7iMNcl9
bzc58TVmJxFqZdkjTsQvUZC1u02XsMNq8OFpzDNxmOHPUTcnwHHKHto7oPKY
TcRJ5GHcD6z9qNOfUPJdlZOJFodWQmO4ZPAIIAfHzlZ6bhDMVuutUJs1bAIS
n3eR6GIRLozxsbpH+IdugiDVhgDopaKTgidULyKrJ0qM4eH0d3TvYFCd2N7y
2Uo8c4awt/MicLzQHbkUVibPCl357t0RMi+Sv57omsQDvXL1hBBqqR+X/vLQ
+7MYRp6WbUsHN5BJncH4lNY0HSBbUGjFxAQ8Kiyk2Ly+fdJWPuFroShnv0UX
jxQaxHsrINgdxB7MyzpzdlTNMiqrG7dSiJvXu3fcok2wGwZCIjZ6NOBmJwY9
EP1kX/JnL4IWVuPcINPn+cxtAErOgCzBcEqQ1283Y+Lu+PbRYKOlVZKoeOj/
S/+6slDyUR4+rbln8SHMW+wwvW/n1Lkz9QHA4PbNVWkizDg+OtwAUaZrMyRu
C5KxEFaEWWwcwLHIzVWUMdscJSWZEVmjAu/knKSY6zel/vygUmvpQDEVbmM2
c8rCATtt84BuhV+sF+r0B7AS1lhyvi6z0T1f+fx5yeuTyyNylrm906ZqBSwm
rFHisMOKhmPR2gS1xM1XCD7n1lQ+Czvn/5VHmB3l7hAyfg5NyCllKILM/GEW
EaCszpM8KZ2FmJZhWf1DEa7POy0x3lvsOHnqydZeYvsSQpkCnQIr/s3rwlfr
FPw/NRatfboaFWeIZPKEtE5uakPRiF9wBzBY0YyQZ1X/hAn2lQTZcxoYzY2+
4L3dY41yUnVFMBOKjbm4wKf6Z1j95pLIjVZDup4NT32K24P4JM/6KaU/BLgM
XPfz3DHRHIbMu1JrKa79nPFHSZHuEH48W8/7BwhfOPmxKrX8QVKZPAsJBNA9
advHj2i1FduYcMzm8Pl5ZLvg7A8bZ5dYTmGLduT9MoN0HrO4xKwbHGcrDNc5
Y7Bo54JHdrlQSUuQRLGza2CpzlKMbm1l0uzRyERnILRexy17eW90Xa+QfsXz
EBc4R/NRJHSqcDxfV5CEtcIodxyvW6XKzkkJI+cP2Pf59Dlu/r17573h2d17
ZCi4wI6A3CG6/lUu87VNcXDcJswHmNK+PW5FYrHbawa2liR5dqQDimcZFImy
MiiKJOwGvDbpyeUjR6nP6bx7oOx7otU3D2rk6GzA5yFmJ/IwGkxOuD3UoczG
5h5Xn9ni3dudmqeYPoV6vI0SoVs9aAmrxvyU7gb8iG3RQXp8ziG3xmcnlPag
xA2G7Duv/QTOuq3JWFTqY+wRPAaowxFAxmEtTX+TZNzUO6HztDd5m7y2rOy/
sMjLwjQBCubllBip3NGOCp5CR4rT+Bb5iv9tKWbe9Sj4x1IipAbWCu3OJ2zL
n6TFZHHl237CLyF8YK4cVHASo49OBUghCxTVSOQwSLs+TYKxX6dBy3Qpk5zb
opyX4WGAmUxUGZeh71W+aW2wV3YX6kIcsuCG9JY0wXU5JyyDtbpRTsrdpk9J
0JXulCBS4m6JoQl2B9MtnfqRAy2r+XXTbwTqcogkcBoP+/MG0JfaPmWF9Ler
/WVz7w73THzlHSAJFBsDhkUVoJmlapfN6Z1wa66OgrNP13LuXtKvxGhcBkkf
iev3BZsLXN8spwl637XO3cP4CcJfVn0BEJBI2Di6ppXY/LRu+k0WYrIrL4Go
X3XBLj0NoEmlxfI94EDcs7FTL1Bs/gAlsz6olKQvjwHhY8NPsy1sNb7yGWtI
3EjGK2uSsze5YGOx6c89vH5Qdl/wAOVyLvOePrn4ANAtFhh54GmnIos9lgvL
yWvOfPrBu/kH4RBosKlkcYu/42lGaRA69JvBioDKV2th7sa7OYRNwj67BV8O
bGwTJghhcAHFFibjdWKmPYsxHm0QWNj/paGxgJCl2CWQPP1blG+fH4CbGEQU
a/rSX+RTwTHKWGUEcvf8tLsYsABjr47rLIDRVpBUt7+BSzIQtuGhlS+eY+OT
yI1CZOWHrBbhuNCljTTDD2aQKs1ia8MJWrtMRkGxwSzc1sb2yjZGuQ39Ibha
jYPR0X2IhIs2hTrxH0DbJGEVyerGTMX+3Eyalp11UburRq3Gm9KJY1vWneDN
tXmuIrWdhYTxaA9DApVreHB5Cq2MO+eXGDREolu2OwmnUg5Xlq44Xa2NX2fk
XJ3/ych8Ga/uUuZk9ZCfIkDbX9fRXjvl9RAibg2KUCI8BBJmW1dArEOY1Q7x
pujqLoDkLs2srbwhPjseUnAt4XbyLQdIfQU2z8E+6xBt6o4NxRc7XoJsWyAX
CYnL9oTlCq0OE/acB85/f8PEXmFl025Bca3x5ZGmod7tY6GQaUlUUVkWJuvY
sqiqnbEd6fnZxSf4xErbuwlFNYpYWalbDb+m2iNBVmvlZjHuVcMVGzFHPRuT
eUsRbTpXfw16dF2WSjQGmylmZ6XaYhUnUbvDrgezDHGB7xi/ClyUdZFZWtn0
+AnA/r0l17/aVl7O7jcIypbElTJFqrfKTPZfUX0R8g2KkyWUF0Scfb4N7uvx
0shLYw8NAjpKPU2K0HzcvmO1kWtHnHgFQ3RKLMO0HVJDp6MVi9mgehnuaO79
cXeBdEU4HkO+RBUGwLjCNPL7iVDaG4YD/MwBzlWZZ8zZhs+y01umX12H20em
DamA5az1HKlxRbAst92BwHWHU+guooXvowRjDtwSTQPD5NwPYJrzc7FqaNCG
zjJKawFe7MQXSmCMZbQQjW/9ZGf+pZN88vpoplo8kQd+Dv/JVDdaBoUIiatU
3WFFsrqbtZCu9J6EProOiLaj/t5AIjEwSu0f7fKAc+k2c69+z9ib4/K/PzuI
ilHQPK6etUzcdWmPSI6mlNj/MysBgbbMeUg8DKNKw2GSfLtY7Nx5nnVVamgU
Uzds6G6iJpPnlf32Mh1LYillrQ17OlzDBIMfxicVxKkFP4L5Vq2eaWZM1JBk
ZRxa2T8J/4Aa0c+uIHWKyOj/8bZwFoywc+VKWK6rMCVg+Ps9haFQdZ4VGIrA
2/LoCG/Gok5tR26x2rUdhXCY6SWPaZHKQyk0VbUrBZ94mRaEk2sYNhum9kVa
YheaeeK2hGeksTseNpoc8mGQ6+pLy4QXg/mJr0fac7YXwRcWkbNhTkQoY/h/
KIkQufW8sPya3zmgkYAVnE7cH4rkwbQl4HirKCqtuREoBFir97uDKl/XmLeH
g/X8AnBrNct9rv/ghBHiJf/ZEd1vIkCsNCkyMMoX15yA9TUCY3Q0qpCkv8IF
BDoFIQf+wZByrIjY9OmMNmIne6w6kUqnn7+oXM2sIpmdgsFaRQ/Op+X9YVdE
TqD9PKimtqfYOvR7GovucTKiKYJ1DcGx2Kyku+UX3ldgXpf4AaVuWxSKxPUJ
Vv/k5Z+ucjqh3vZL6vnV8/N07HhlmBzlm7ZlPw6YslDLfQFC7Od0wTRsDYHj
u9CwrIfpKEHXCy0rF4KzN/Lceipr9tmeP+YxtHeAY6PRrdmaheRMEXP10/xJ
3RSU32gWl12IjWTH7JNEGIuJY44LQirRP5+WsAQ46xQBeroc0tZkdlEuztuE
xm99wX7hq4uGThtWXyvTvV4xGXKXfC5gpL3Fxam/tCjOb5rPueIfhfr/PuMD
HoF9gG+qNZkdCu4mweAcFTmEURmMEThh+KyARWXXieeNIiABxXW7QOeQ+kz3
pRaFEqhghE227t3PbOwKt0NS2PojL+9rJly7AbSSvZ4a0qzzOPYhPA/65nTK
CdPn5S+TtaTTgOhCq5CU1O5nOGVbdb23Lptg1AIbYX/X1a+E3xXZtDQYETWc
XBn4dYweGsKPmw3+jPC9ocbamK3lssGWMUqrOvH1achyuBPCJ75xvw4/J4jK
KBoomqHrU+WeCgYCQrM5BbVVflFJaP3AMlxg9Cas+Bfgp2rqAGPlqMvdm8PD
d2SboLzvraZOX5V5ujTuOZB52LQxf804crZMZpxxf7tVdRM3huYUDy2qDBap
hGH9E73dvskJ/tSXkEOIqUze8FuOWjBN8KeeFBkoOyelehK0PwChV4BcB5wj
5eX+vbduESkTfnNOHxKjFnqIAN9TzLHIBsP5GeKnipIu3tgDa3aI2g5Cz05M
UjAn6ftlFEL+0eqVnew4IOBZLBvdaxg4Zs8Cw8tVd3zslzLne3YgfYpdybUM
geKwItu3i5ktwRxQ8pVxY3OXwK7qbBOGhUr6Q2HNlvEeDttrlLkO+mYkbc1G
3ZjoZ6ePWXYbM5cO28JvHBwvN6pSI4l5FxU+SX31ARV5xk3sIClBBpFRTqDt
wr+wR47p+sjtk3+qFdTKZghakBJIYg7lyB1SwbDk6lLJJjJHmB6CnsUh9StK
jhz3QqNIg5a0Joh4xVGcaGHgHnWya1A58BBLY8ts9UrlE19uGMEC3b6Fffx+
R76nyVY1GPd7s1TKKNH448i1DjgvYMqP3VZoqZXXRxxmFM9xLKNf0Ok863tm
8M07zrQLaGrdF49t3UCEPFmM926uBg8COvgYQKB9ECJCl2Rvp1Q5+bN+lxOj
PUplEuu8pKEBRZUNJwxJ6laoYNxS+3vGzBBi9wiKNWs5xOmHOM3ef7rAlGlH
t+Cyv5PoVoKWIHPudMtF7AnQUfX+5u+oih1EL/VP/kF+1lrctHzJnUoTb56C
NtLrl5dD3FjQ4VJ4INlG4BXLSCqFR3JtuXRPTDa1+4dzCPVlo2dzaoDQNNxb
cQtL2UFPKo8cCFBlNu6xdENzaJ8mqGqYX/1CJ4EOpn3e6pH7IkTsLawUhhrO
NzuiK0wb4SLtnoZbVccW+6hJKKNqXcaE2Em0ud0zsD3mW2zisFsP+f6y45Fj
okoBKPuyKuoWloWQ1wjaZBCF6/RtVgfxyfdSgveB8owC+Of8QB+8Ij+lwNSH
cGOniRCWaogEjWkLknU2aANKMHuER8nJEGNP+Q5ha5N1huF0Tcu1UWykkzmD
NYlOwU8h/XFbYR2efDinzBxDsyzglLFJiW63nJk5KFsn5HwCSSvM1wnHW0Vl
wxoK5RzjVCip3i07crG4gXDNQF6wcvkwgl4mCUjVZBhS826ja363SYTzsZ3D
Tdx/yn2juyYbeoFuagUUa7IVh1nr63klPoI44dQ/2alP7DwIZuunG4M8KWmI
4gIYivFmjviLHIZS7pVgCP+qKdvk2tnZdtRsIJKipT/sAVKQ4mKfT7Kl5TDQ
u3Ueu9Iu4vWHmlTEuiw2kMuXMF8ZGYF3QJ5v4LNgXjg9QZebRM4WD0rCPqEg
/B/39eMvgI1Dn3gFngvduFaYluk6m/fZCssw3FrO5fcrdiUpjJUHoKC9woD4
94mP6Qe1vfrNKvCafEA4brUwosvKf1WtHjakKnL1rR3pKRIC0EXFAEqQwaL0
h929LGvhEOkCMunOtXlo0BZeqvHamsEwVhcGJ+zLb4FdBrhgmSb31aFZ6kUc
yLe3VWDQ1V6Ufw28Kybq5G9xqLYaz8OyUuzKiH4InJfV09WM8iQmKlQ4gd8w
UFhRLlT+VVL/0EuFD6Y7PdKfduUoHR1ZSsJ0ArEhkPa75muoNKsmDAqBu8v1
dmPNUiHogwbA/yugFonvaugBwifMP0iW5nwF7F9NGjJwcjLGgsF1CJfMGX+s
XZPMQpeA3XwiiBinbRHAX/vx2r3FMLoxOQ0Ear1HgRIsAgf/o5SCWEoonlmz
J8bM954ihO0ORa3Er1ElGhH41t9GKjpdGttDsqmy64a1cWtF4ofzvK1S2hhj
qCn541baDClbct5E6WobAf7yqRjsxhvTzWPqZ3B91TwFoLOfhBScuzGUlEh/
9cecg9gp00BF+RQcjCxxrHN6XK/+MCjOA8hZJ1NYxcuCju+hV+vtyyaBH3rK
FpLeqBDkrU0zqIxffDPPUVPZgyHsWMDgQc/LNPaJajcZqk6nNlB0wMnjSM2I
d7MGAcPR/9a3fj3o+gXtjXUD45eYM3KtqkO40KYr99lErdZFIoO1haF5ukOO
wkcWzF2nVk5JXVfSvSjJxiicFIcoAQvlZxjyCOHCjEXFhR1IfJA3vTSJw7UL
ZRzEmtcr78bkENnoighDLrmQ9RQgBp1eEKCc/rybPfZAgNfZknOfiiR7A33B
bH6Zc73cNykyL+0w3E1r3u90Xq0lUd7jN541tD9iDImWOMcqrOP4h7Yih9bq
EBfw4dooCTggReVP28yrp/+sQsuy6kEoTT1zMbCzaSbjT8MROs2+dokCOQF4
t3Whj1UGoDsTBtYdZoBbhcLh4O9Wg1JOw7MK7AeHCu8ToVOr8ko34o/SJjRW
5juh69Miv+KzBMFzAA971th91rPVm3cIpPDLzopA4eg/gibqdiXbTQI3hJgc
9nvNbxQZ1c6WP/l7rwaKKg10dCHpc5NrvvOpUO4yTao8kWkQhR9NPEqlRYse
IbmnRMrAfJpGgds8yIDur7ZLKs8ysRDBLRY/InmUXb+3S7ID533VfmcaedCA
z+3RBrmU6t5YOEZ2GC955hYVJC0//0IeRhIKUrSmo3f/EbcKaQ0pMx9XKI8S
SRiC8HG8YMQexZSHPbZfPqwavlP3XygW3vWsocMMegwsm80Y9wph/nFKE41V
hjF6bCFeMtwELp6bTSMJEdN60YlyMIFtoqZ6zIQuKNoz//sFwHLx/+6OkIyd
DFXMbkZVP6A7hhwDaVSfmAzOFFjckpdP6y4nwO5mo4oLWCh/IEJoCjUL/88s
BsgcTw7czGPztlB6wZ47dPKTMNoYvNJ9hp0IWBbx43atlpPw15nUIAV2oJ5N
LZGY5n05QvKp7aEqmv8AhTXeTWP1fSzV6lx6WjCiBjQYZDy+9Lj7n/+OZmyI
e3lD+RDqroEzMFQ8uQRVFafHBMbNfVj+6VLLAQJyosOOIF0R7U7pUI9u8kCQ
CBI6ZOqwKCnLGcGrLCZuwX49t4/7tHDeinvJxt1QryK4FAYshvlpZfvjH1gY
vJFuaUL9qzR3sZBBi6gbgOZd8ICIXW2au/Dbs5KgO6K2cT8pLQDQVYz2hf/B
WLx7+axPqAWw9AWwvWGqdlFGN0zyjF3WrLULvqqhzq8+q5ofoDayyPdt01jm
PaFY6ZZ6jbNtk50+3wmHyEQpdtNIouqrV85d9rpLchjo22R2H07eUdBglFg9
jAZoJSYqz4IHE0vbxGfnrufmNlEg2o4a90RTdzTbM+161TMGsJe+KkAMjKzX
IY2U4ywS4a7kTdKxBL8Yn4AJZ5H/+vbZb9z+lAJyIfvtRYTws+8Ql/JYtoyT
Rtvc4uHNTRzVSeaY1BUDPbbTLwaCbM3eW+G5EVOYt+LRY4TtM7I6uxiwBYP7
zfXNe8uWj7JOZ2BIMCWSg15APZHhnDbRiHhWF7HsXlBWbizeGCf/vGvA4op4
c5hgjtb+f5po9zDX5YJMczAYTj6uS1AXHqd6Dq35Po/RbUpNZQC2TpYUhN45
331LI/kdtaM4ncdarhSxZLyFupWerkqSNazREK584dwtjAyM9FbU6uy7b/Xe
2qo6sdcV3znBisbXyZuI+QbXLH8UrK2+43UwFjFup9uoZLszv6sw08P+0JoY
OrydTwT1jY+ezvJxyTqP4aw7XTOBggIkSxcfUs0x4H53LwkKeSOxjVmJZHnM
xIN5T58tzzN9O8rvU/0/b9mfFVRvTy/K0Is2xm4BD18Q1aGDwevDYkSxyLj5
h45gpFhmSfUzoQV+C28F11V+lcjk+OPcAu5ug5A5RdQYQs+dRrQC/3+mHRic
oMlWIm7YoWgLnZTtt9TT5j7Oirpy8YGLFpHXqknb1ugpU16o5KyHRycOx4ep
EAxZg+b+v8bkWcBPMsTVF75sYgS8xAAE7uHsCJJAZkS5LVfUaOjairtuUgsm
oc0DWE0i+OrotG7iEHtHr5PEaCKXD0F0Ial/7OAQ7lrRC1/fTVUhbLg1NS1L
RuuIKM2dVMnInL+7DuHVFLNUY5BtQxyEuk12Baq5x0Ug4Jn0RMoTXFcgzNEc
CcG9bfF2m4mGn45eLl4yWSA4kyFCP+a05j4OrbvK1zAeAVwuE64uHO8ZCIl3
97EQ2fPBEviwvy8RPqs7Y7mTJzo2/ec5KVor0k5lRh6Ent1hlglDAw5emKmy
wzxiVfNJaOWEtrgqye+CObOlpSb/kO65/75ZwdP4mwpiINY2BUjkkvS9znjD
BxDQ+JH272ZR/XdC9ozQdLs0/hXB+kBrThOqng6TKTnCyp6zIZtJJUGv6me1
82RvmX88oHmiE4l/dWFlHK7IapGgfGM3DAl81h5l1Sfzw68x6o70ZAQDwQHK
9fE/U4AMEDECXMYeQfpk9T8WoNy57TtV38Fju697yyYohyhCGL4XZlCwGIi+
qO2S6rqaSvZNe0NE7Rr3HS6JHz0JIyCMzgcotFWQEKRt6kmtXrgs4nOaoh/D
OG0MUAaQ9m2qguLPILItv/ceWkrKfFSda2y/X2UZrirHPqjsGeqvtDK6K7Eq
i37POt9dxd8MFl/+cYJ+M0Rfjm2U1It1LHKVu7dhqpLe2u8jnixX2ZEZiNuv
VtPUToc4yT5VbqZ+bnF8We+Zcz+MOegITrpXcK1d2mjmfR76tzEANLy8oeEO
XHUNuSrv9cSLZavOAjYlxFeCbsO+F67WJ3kNFukRjTa4CRawP7bmglMys5mF
H+aialW1+j7HHDf5HaNvJ07XXKhUE1rxQXWuBTBHFMcDTIlwL/STKBbCay1B
bV/AyLP5PeuQwszeZQCSMRHDZokf/T5egdT/WVoVicmwEDA4AX58GRlCpXew
/D7xWTJ4mylGsJA2M7flKP7I3SyBY8HlHrrvQXC4wM8FU67VdtjDviEK8/tH
mOf1LgsEMTmnNsuIGFYkgwk07aw0GWJELoXh5jgftUooX48GQ0Szs78Q9ibq
nWhiSrI153lkxCPqDnk2z7zMexoKxV/Hen80XajPu4cauiCUd4AJEvfesdou
EieitEP7D6bEVznP7TVaVIuv5AxYaLS5c8AJ/SZgM1Rg1qElw96XYHqltsMq
ggCQbEZVzf0rFDHm5MugfvY1LJUQg2x7QgIt13GBjuDuY+jlkLuyi6ZFspgJ
YfCK+vWV1gL0PTB4jaRzvZIduHghX1mnm+VZyrS8DE05p9WOen6BoVgbdmcJ
QovnBoQO4mq+OFUdkFlMPEWsL7Qmof0aR8eyJxNFhBL/hWQi7zOItYBpdLUD
7iEC9zkKiLA36me/4YiQB4efT+PQX1hKg3ekdI34snNzxZ3/TPMcviUzq+70
wzuHAmAP1K6D4DB/EyPL5rTJGcKoLgb1cNroNZ6JRB7i2XVyXv1XQXzuseFL
ZZDsS/fr/tRrQcrWQfnnVq/djHmGgkkEUEukgLuZp7OgfWAB3ytCSPiQMU5O
4pYAgCaHxdgUrxR4XzSukIK0v/24IgfyrD11u9Gb6UHBWH7BeZM9oekgqPd9
J+YC31fy9I4WHL/+SRhh5kX5fxHUlSr08+NbXZ7wYdl4f3Utcq6huQ5jff0a
uoXpVrWW/owP0ZOqQfLnQEft8WK4cNq8nDvXcppq+VYYP5ekMAr5jdcjUMgm
j+C07y2zjUuoJFoN70t2Vmn+HainmqHz1V94dlfEJTeAa+TruD8SoU2Jq2fs
EV1R8OL6oNvhP4noySKdLecfdl+z951LbOrqtZ1UFuS1t/CytttIHZ13/nfk
uhQMiGth4aVsQ0oeL50LDrFsNF+FACzpCu21XDhORHmVdalPEODdajFZRs8n
dlFC+9VzFbC4gavOWm+2IWcLP8CMqZcjJueIGJVBz8TGjjBD9rbCdrbhQ3L+
xmjEmU8ZSfvQuct/0KVRVSrhhuYmPfLG8j96FN1WIHEL1Y/m1oOMcv0mfUZW
jo2QEcbAitdaVr3cRsyCoNjA+2Fn9OlzfN898I5Pt493AoVFR/HoxiGzyQvP
1U8Rjw9mFu3oJ6S6lieefG8HPxc8kzcko0eI5C2dDDI1Vn194EfLpyRxF8cw
bSnsy9wQfvrIMGOVN6U8t06aUMzuu49R9EEZrrivc/Xq7M7XOOoHFichhLwq
DE1aasBqfzQhuKY64XRKnscXkh4xescA4Hua7nx4N9yJjQV2+isthkKi8+VT
v1NplO3d3cA1upwS4k3jaNVxbzQm4OQE3na3D3OyJP4LTrPdUM++g239HGan
mfXuJcjOndVqjPeTMboSvRlzDYuIt/SDC6wCbpOQFbd5mfKtzo27Tmp4aQY0
BdqGlGnu73gmUJjsZUSgXllqVHJ5ljrHhr36+AJUzO0IJwOgHyo76GOYshvF
RBA3+76HPm8MRTyppYTBy36dhFYg3j8pYe+sOePSwyQOYWJka7NeCTljSySk
o2dwCaeWSma+OxxWA3w4r3UUGzD+GJj/W/QI+ik5ZfTgWHStMFX73/NEZAfu
eyawrLZyPI61hUTtpUoS8/1HobI5z1nPONK2eF/JqhynsCrIvpDDGOUx5Ytz
yKfoU9MGix4XaaA3ghLvhb/UJ7uJ5z9ckowc+DISeFdwicv0GsQGGpPibRrs
S60y0RrEf2EaMh639jSc9dDQwKdgy5g6GStPqXuRVvDfna5JFr+ua+5OtAcP
F7s8qQExrMMMAnFs2oikTRSOq57MmuytAPhWd+o1oY6oPmlHjoLi6mB/GGwl
m1x5t6ti0nDdf/evVn+Hvd27w14L9a26xws7xRqRoayuQ3+NTRV2IgUrEb8s
pxFTbEBmsNH2PMlPjTRlAsYO4pNJVSc5s4FAPCJrZiGN2CUEGpR1wPEHHacJ
DUl+kgl6/feto8wB5gU96qCtR4YvbZ3a+0kUtdiludRCWDC9GPhMWGNYzg75
iVzOOA4HgViXUbjoV0j4jtHG1zRwQrrP6Oq+QeLLnui69pkVni9UVM16W2DK
Xcmq19z/EGdkrlHjPhhiGE1WywMIEcwB7A/3PTvRvlu7ZKv7tUMLEIf2nEhU
jggCp3OWn6e4FOmC1s2A6GTO0Br1jnqCE6NbchJoI++DvUXhxlpiR4yrfrkT
icA5soi8guZG+4rYWoVoI5wOQOLyqLwFyeQtNa1oSKXfaufoHhkmPRDTzZ9E
kaevwYwhh1kNtZ+G+4cqEMzGmtWmrUe/dnsEyteFhDJOLg7TEccAjiBbJpe2
Dk6BJEV1v8weemzxN+P1j5H5uVlLufb3xUlumV4E7seIV713CVi9DD7S0/s3
TTtCkr/9wYny5jYAMt/b/0ja5km5u3LU5OgYg3UKlUaDWVqte17f39xJgnQi
DGmSXW4sPkIH0Jtodz3yj1LHcm5W7eFq+v11wAUlm08Q214w9Fs+ESjhjrd1
95HKUQCHHYNkdFFJuif81YDVVPCxUiOMSxFVLUxAUjDZcoOhx+8ZN0emzQzC
BV/BhcrG7UJQnEWiZ1jMtkb8z7GSx0wV0jkpok/ZABhdQLT7Zsbea2+dPIow
wgwjh/AFAExR+sm2QXj8ab6WumnIrieqdcG4H5ksaW9x1QTbRahCwesvn8VI
iVbzSmeOcMtC94tpoL2Ismsyx579eIcF8qFoqmFOZHQ3tz+nxJSNIl8bcKED
KTwkomVpKrSRqUXSbI0737noJ4T7SaOdBPv7ziJdvYLSBd3f18cbPBg5P9ZJ
Z7fWpVxQKI5TMU7vni/ymz3rZ4Yv/eYgF94hkbEGvJeEv/MIljjCFjQSZwVT
4bjjZvbvWlO1R0xJiRiHYU6Wnekyzn5Nq2XhPE3ggCSG9aABN8toig8epJ7O
RN72ryIUaD3htKC6xJQZWG0I96iIWsoff0VtxeWHNm9TUttn4vfT69AXE2HO
Ag7MvylXjBurmr0n+YKxGnpFRtitK18x3bIhkMHRNHI9KBvrRhXVMHorfBK8
UrRQiHv4LbBEIf9xzZVhzylBOMIMbAZ50RhnOkq2baNszcspjrYb4aWsTyEO
arUDM5J5YOhV7Cr5EDEx420006hIIbDcI78ptJC56rNfeyB/q6g/9wGZDPr5
Ntib2aGfLNi4U+wwKbMNGT4jJh4BYVkuUnwxt8hiAWmnAyx7EI21DXb3+zWC
uc8Z0j/XOm1FAYI4yXAhvFvAQVQ7f/JCuEzwUnbC3eyxbmWNpZ85rpck1mQJ
NOuQJUmu1gf4EMTa4/FqNZEEJ0xKTzmbhwLanB8SXoLyb+9OLNDDD6t3gWCV
hKKFy2UG1SBlSe7CrBOrjNnhojRI8s0KLLJSMgRk1SldLWvN0YY+ez3xqR17
iSbSbU1aeuIKvesWNycmkOp8d/lMVS9TjzYm07mxFjQ8W76TKxDQjLswNA2+
qZRbjRMS7OvfmBROfyDO0RMooPkR3O2fWMl44KNZoNPRcZWXpRXTl4M7sNmt
+lOdAklehVMxwYfhUBpZqu2nPAF3VboDvOWJQfriYzPTxwgS5oOpOnU6GSjV
lSkVMQhRjqq4ETRhMuBZdaggLK7PY8EIJHQqPZri66Xf2nVxYK/LWfQOo9p6
iTo965/CQ0vQsBcbvXFO41pM7iudUMFcykoSkFVGtmCW832Vo0U6rOmt9xnx
VowYLQbm0E40hmHOy6Ee7f239/Th/6NPD3+P8i+yP2KaYR8ngpA4sJ+ljOlH
KoZf+lbRIXeLPkkwjBm0sAl0YkNKxN5vMMoKA3HefFYo5MATYw9n7ol0ow7X
WBSV0mEfAlIIZRTKWIpZ6podUtdj78o7dogndcWad9kW1TioZbkwAFkvJZLH
y+KOPWc+eHknpDx5aIxqJYSDGF1HcS7ub+gAkNoRqmDOHt+3lWpgZnOFSxYQ
imikki1vRqfBW0Y53LSn1unvRtBvdvMmeF8BIzg/y5OCSBMP7X0hSxvVqEFI
uYTn1ingcCPGdippG21v9eAITl9rvsDxopdyKKK15a62tnPw8uV1kaZ0LZUW
yBw62/yKJCyycsyPR90PjtuB6pweVZUR+typsGDxzqYid5mdaNTsDNObOVdW
BPXVeaUskZHEZdWo5XyJUptmhX8v1oCUBGvpWkK+drCCsYWlJfH9BbWa+C50
jewMe3TH4ApcbSJSUpzVy4uhaC4yaZBzdD82LUZNz4Fv9Nf5Z0cEOm9bHJFy
LI9doJzBa/lGUajuEXeBQCetWV+HANxwcvs2pY5yGjm+B3y/fiZ6f7mzIcbz
UQlpT3Xxb02rgTN7FnWgWvIpu7IyidQhYRhvUB46qFUK4HRTKP48UEP1E3fc
N/R5waBmXb2DhQYJRdTw5yawSm2ffCcNPmqc1YT5QHhfqnI/RW4w/rW2Al9p
mZReKGP6Qzgj01wpMEex6VLXZIGbgb1NEbcPkITD3N8AMLHSv1MU9v6K66qH
MnGya0TWzXcJSCmsCKYK9+9B+/z52iK+rNgnWyaTDZ02yIR7tDyzVnYrjZVn
2WjZZ5WzfCqLo3BVuv2ay5Kco5jM8itGTf5G4rme+bhmaLW+Qd3CsMKKMnX1
w3l9h6QOd97YtKA3oiolyrRrlVkgvKy1I2PYgAr6f+x/e7s7h7dcMB7/PfOz
mGyahR/RcoxtrcQf2OKluK1cz0cZGmuanVSLxlkGLIQG1cL+BIE0Y5/FGEr7
49QuGSGVna0BDeNwT0QaM+vRqlqhkvdTVzLrMLGJGnMH3mjqtoVJfISeCKZU
BBvKZdw3pF6GDxK+Itay2AlS6U/txPy4b2mIQiMFdsyH4KAh8FOn8gzZrUaR
vdKjo2H7sOQg/F9OPyuri2Cf22Z6XRwtpbm/HDqdw9keWGE0mNgZZfdLhdoa
lfllGy9IPA/ukBdVWLvxYHmhBcIXoZAImkmX5KBgfCzH9TZ8iG6Pr6yyTXYW
85w+cwMgO+l2FVqqKhANZCsw+J8OU/83SfRmJ9lTRLeMHfBZL5RU9bwhjz1x
Mf5UVYUi+N1y86bTuwccDHeQiiwDa5juIiELtbCQIXm8Bu4T7rG3uV8tRFqC
6LNF1P/+VqzzK9l6DCPWEc6BXdrk8TCmjwwrk9gslE10RPv5Yffq9dV3ocRz
aFCFLHJHTnYJBRjdpOY0g8sPNmk22ic9OnFXZryccFz/N3GTd/1s+ioHwAEP
/a4K+buJRDM/7aPKCiwMxGgD6Co9UXMzOqLTppoRxuvYy/NHQmzh/4o9FMDS
LWJoTmzVC9eC/Tl5/kyjU4IaZ1tKBNKGQ9f9h+pg765TyAr2NXMU5RFmCb4u
f+uTC9hWjQaAXP1XpBcw2dyKGZj1VvsTYQWnMqovNPV8mLWM4e19IQoI36XC
qF4JfVxA99fE37SLVwiE3zLokAkxQKkqg88ZqIsXNpVtYzPPfb3X4C0ZaQYZ
i4q654bUfkUXc8ZAOzOCh/WGoCEu8cv7RKKaHgV4H1PWbJ61z+syesXvKC/q
zLgThQ8PMQHtjwVy85qvhAiwQO2vSgaMgT6I8kntzcRUt9Y0S4ooQMBBGXjw
R/6TKbJEc0shyMBqDLG2mhTxKTHi5r0ykoglZjtF6dwgJUnFjB147oiqBhjh
ALLukkzSb8+g0+RLTZHx7BBrwdNflApadfOdfLE/HyNK2i9tnie+HjjhCGNq
vtsiZU97Dc+L5KFzQT/S2nGAfTsKAvL7bdvoUvWvQG96b6HeoudUq3OSCNQi
EENd0xo9HD81PZY8TWrzjCm2Oy2vXJE+1/sudwgL45BKz1net3B0N4cMzEaE
iLoG27ObSXdz+gU4OsNKdcfRznXcFtUbnH3JhE47ewg6NAev/hQRmbnwt+gD
l4Wvn8bb80eVTDYzk9lsW8uqI6jVyKNDE2vqi/LHWSDlo+8MLvXMy1K3c+tC
Bwh+h+epCXg+BWOhQRrvY+fXsqumoZbR79DBpwXqnjFzi7TVK28xuJzrnM01
wDls5BzSoX5FxQXWYjJ300wmwnhkFTXxjjeWL4jbH6fZEz6Qn7F6G4BOds/L
SPx96rJpfo3TsfzRlI3zWu0w6OlaLDz67ZAICoTB+ASCUkNV6K+yVwKvyVm+
WB3W20M3QxRlhnpQlKqV/SIrKfcgTedpiydvFFfFvUoHyeGneXnbSTbFt5Cy
m6KsipvndBKCd6YdExODOYF3zkz3A6Wm25L4lg5mz5gkdA9zgB9xaeHuCfWV
AirEZ+oO/EDRZYpmUnVLdUvQ32rS/qEX2kmiDKoF9/R/+MUDOn48R7+SsuGl
yuhr2mOCy/6PddE+8cr1ELOO4tKIw06DE+KyhFnRpsXtLXz3SGbQwx/jowL0
FnZKN5KrHbCTEF8tnQS00xVxOFS6v0ywh7NriOlzLmDR/t4v696rTAG2bqXN
khBv4jBnNeiBPe57negywpV3OqTpNJS4Z0AsglorVH/xE7G0XnaqiESkOaV0
isOW4vZiyhYCFAYcQIGD7nWuGbFceN0r/8ad0pOq1QgUSp9BQVpWGPxBIVy8
ktowcx9ryNMvBIXKjgkKP68O6UvrEgTepji/BNG/+as2lbsgtUB49163jRKF
YmMwcbyBb6dE70COMXmRy8RiGET7Ynpjs3B2Gq1PltJNWvhtWMc7UasCk5qF
d5xf6ZszKpwcfflBp74W/BQMIisiJnz0pGjqWG689K6ioGul0i7VoZ6rrQmN
/d91NQDrkp72ItlXHeYJt0m4gmXrNaDxSAVQup1mK8cubW0qVjiMpRFTHBfM
Yz4WLOAE5xZWYJ7N6pjqJf61dp8E8Ko+3vA/sEr2dB8Y314IzXOrb/exXTDN
qXfJUqmbhpt0Rs2v3Zn4FARPsPPD+KRaDJm7UpAYZqx1078BekgNwGsqwiT2
zFe3FR8f36JMwXAIF9oB6iNhcvqGqmW2GJJkZNa7ZLarxJVqGMTD47Lh00Lw
3s8gMsymF98C8+/b2MnYEaEAPAcgrlHtiDKdyUUkhFOJJ7MS+EpASlMoCakq
1Y0GGFAAPKXsnhbBainSDpI/TWHkUrlVi10itfN679u4HXje8kr4QBsQblns
FEbOVjXTAToJVYIMk+7pUMetEPtTDED99Help8XNrCsP1r7EI6F+3CWN0weP
fcKycB/GmdWoHKnX4+885rqdr9CXJte9Q0RmTd8jyJJrYe1iQmZcUgrAk2S1
pS5dWqrrVSUssGiNJgeFpimBnFaRkkqqDR8YLiJL0vm+33LeaSbAoeoljr7Z
0wIu64koEZ56mlgnoeag2TOUha6M/cJ4b/QZsDnKyEAVeqgmaDe0IVrNXgaw
S04XcnbWFCGFeOjAosTqYdmsFicvT4NAbvsF9j56jK8bH9Li5ccMnHkOVx/Z
omqiDQ8chyh6x79wSAzaUZEwPhrvb6jvJfnVA/7Dduo7ZeAwPQZ0u3Qsx7wC
n1VK/mT8IDewcU1rp7Jbk3OLjARJ4MSNlUZBHz1Gk8J2UHpRaZEYJ/xFkg0e
puURqoR02mzfdUghYPaOMnh2/MWEFOBGivmoZS71E0MdNUWiEgjO4R/X4e2p
j0g4I9RHC3zm4RSKr5JBRcMJdwk+fE63Sa4DB5V8AWdJVxuTn1lNaJG2j5ZJ
u6z1w14n7fxGmUyso9G5B+dtfOpf8hcczOV5NthS4urdf7FT32bNSPDRCSgD
jHgHCgIaEfGKaYOZrVALjDLGAP8Q+q8VX0HkJCV2F6IAjH1T5sFqCESCudQT
zU8qlqxNE1LPIwi+PJ5gS0srX05UGEpegwSAC6Hnxix5eF0RS4aA4X1+Z/Qn
otsMfw0a7+JRwmYHdZ7bnDzzDsMpsojfttssvKZRxBSMBxVGqx7iNTa+9Ck/
5vh2gG0OTppiOU6X1C0UFvW6p2f1T9o4OD3aFzpSKMDltacOIrGLSzG11N87
BDISfCRSSRNNPmtrjaZJtBEru/aDx8OzYpYUN2Q4GQlzDdDGjsp6vY29nAtx
IQrsCER0oQWmJusLvifg4GtuHiPd0kC6rPw1L9LDevflxIZysGvYJn1tmIPo
9g0y8bIGdetAUcdeWM2Xql4VsP2swl0t3wMsRn0Rx54rkOlvdtaQ9AoM4vad
7G4rN/Yyd+4THdnSGNCU45mba1VUGTmgqcdPZn7E0bOBzuzxXfbUWoqQfNdr
ZfevotVJYXdC6dKzf+k5tdUtdr7thGaek5g+SgZGzcnqSKk6dQ75xxLpYJ0D
OnoykHjv9msEXtw6AuClqrOYKSkGYPxhOrT2NW6BO5uMwBa22BSqjt1BW0HZ
/MnQjsDWamtXBBBMI3bmOUlFtyJPYD4isDZ3vkgiWlifSA31+KAzgvYQR9UX
3FcOvopi+Gb3exZImhNse7qgUEoLDWdsXOQpdmZaSGrjc/9/C4ORS82B4BoR
o3V30auMVAfuOK/oYA2WT5IlE2VucqZlK+LaNOg5fkIgxNbdyji0PBwfJsL1
tYSfsJec44zP/eWEhlgkovuhyWILuEphHOA1jaCP6x8OBfsWkkhW/BSu3ltw
Gr8MGGgYQGt0eSz/CnWPszC3L5iEjXe0bZtqjYoagxjcjm+s667EKyoI3zCn
6RRkpqzNZ/NBmAdJYYsFhuMpOdYqeTCcH6A6bBLQxzAumDhTrAmfOa8ze4tO
sAtPyAn/qscrJEu9Xxj2fvceNqFeEKY94F57v1g/OdDr1izSYF4fpzK3UYQv
pDSO6xnEcMUean8Z9xjrAMdp6PbupQCbimQoeJrSAqH8PgnoQmBfuGUT0bLP
ovyG1e1cJRGFMZ1Q7TADD9FE5RPr0XZZHBrZBCi8wIcpfCZIvXS5R+LwHlHH
l+mnfJf7rY924aJGTWOv1GajTW234gz79JokWJXg+htif8ePhIb1ycAS8nPd
H0udzFST16Ihxwe5v9m60Dlj0wWYM0pb2yXZIH7pI43Mkw+w6HmMqWnOcfkd
VsLzEeFMJcMWzwGnLVr2mvs2jMwBzuPrg3oRR8Lz4skqr2xZ+7BkIp2Xdygm
cGC1/01BPKxArZvJxIkstQqgQsWpYyp55mWqDJEZuxT1f5hM0X8WfM8TWjhv
PuEZPOHq5z/QZwgK9e8I6klKF7jDE+ImLVgDcWqXCl36w4xObZJRe0sZKHzI
Ww0/Jho6EMq+98Vk0eE7ccStPLn5wO9DT6XEbrZP1Wtel03gC3crfw3UTfRQ
xBu6Zf+uPVnGGRu4tDeEzsMrnPxCvWr+Ticczct0AWM4DTj6K66mHubOPMx9
f2SJMSzKFGH4ZHvCiDD4SBXj5zB1AAytmfonjOLym69owMEajm7NX3iLhhVS
1Nnm5fmOqA0KtPOvXUrveCpK2TpPPaM3K5Y97fEbQzpGGxVi1zITucTKL+a9
c+EBXdKiR7mLCkzCZSRuZ+S8SoDh3GAIadC7RbdIP//cKVefxlr1edY77az4
5hTwsQ5MN8erieGgfqlVBmuhOAU4uWGqf+Gd0SzZAj83HvII90k/pjE0M4ne
uIoRYjzolRiFbfHwrfyCl2QkTeCIi7DHFL6LuyeCtaTQJIsxPLIIpfnUdSN7
8mUQAuTf4G5GLnHGIxMSexN/gB9OAP2ZoTcfaAMMWQbABeF1TmRIUJq7E6XE
+pMlinHwfqEvEpC4/Ab+QcRAFCVt76jvwV79j+gkh2g1eVDEK3/1n2H+vvO+
qgSUwoUj/Ibgb7I+fUdzB2oPuq3yMMNSLKdortL2D1meEn32ck+RBHQj6Q9g
1KIJz6sbo6Zm6PNe6HH8aI3LLDfbvM4mJQBrEZHprRORiSdgR2bDMriwqZqz
bo4kIqtKTI3Ka2ynmijxsKJvKnfisl/POoLrCYWRQf+Xs095iP4Gp4G6lj4u
7oj6PIh7na6IyuTYEGtZA5hUzH3GO1HdSn5iHqogsr4IeErFsFgikEk2J0g/
ghUFOqrIFeG1xQKrk7p4xkxcXp0MQL3kEV2rhE/aDHBdMm9VxkBBaNnHhJ5Z
uohgGCxBwOht42Tp9d/ImXxm4OC12yrrITweluFzhHfqniK6ZWbsaMQ2SjNj
BLvVeKtDMeD0624mf+LzzxM/0Sjo920Z+0CaQSQju7kinZVI4qjIPc6AQgGb
lNrxS4spyVjht88h8PrKekbl/+JLwufVFesYK//pvKrAyiqMzB7eqVTH9ovz
HLIJ8RxSLU6zqUxtLQtrQS+0g7bO/wUgRsXjSSIVcvHOGmiA+DjXvCe3cWJ9
ms5q+/qwZsZHooObQAh9rO/NyI4G/7clNL+99gGBMejf0uZGB7Tyt898Mn+a
JVVAQ/6sGa0HZYFRLqTT0JovkZpKCXcdJfPOOEQ8pqHeajmoCXIUFklE3Q9b
WAPVxCQcvYGVUDhavzATs2S44WUSHSZLLut6LFq7Iji4lm9yQgbQpBUnHAFs
hNrF82rzjVYLKrDb9Q6I1uE1QZjFwtXgYoTMdcY/yd/SFFNi/gy+AJFenh86
g156bnv6NLdPHU8KIdhGMXSRiMVh3zWsikjVBdhrtBBx7tpwcqQEq3gJx11y
HTpe6s0OEJOXacfiji+OsmgIYoxlsyeIBFI3v3Ew8yaxJO8LBwoMsSfQQERL
CeaiJL8bHlQXfOgR3AvFyyCuZGmoM6C4k554ItaXhxBalQbRZNTQV2RsI90M
U0K/hREfJ8z1eewP2bV42pkmE3MEay5pw72WkA52jg9NGhRMPIyDmEQcpDjc
t3/okvnR0HKj07bHxDGcCuJsW7F7iAz41//0UwQWDjmrUzFDrl2KsH9qbmNX
lKqeQ00azGiReVpklahFHjQdB3wOxTulZDAGJGEiohbL5gEWc1zOg+edFqTH
1HLuPvez0jBdjImCEQqnSuktcBKsx8INsv5rZAmYaoPXtXMhFF6OBXY+Uzhv
hniIo5ORtkVHn0T7XoLq0cQwuyEBt5uPsIKKtWphvZes3QWBHup4IdYimF4g
tLesxDLUmngSX7Dqq9+C2a8dxQcD9UuKTtL2p/aXAKMc9887DedeUMHXeSlS
NCMn33fwGfrzmgZUTup4kHF8a2RJQ5IQTtrdGjmaaA74rQ6TckboE/p6W42A
qb3fQPf6My1DHHp9I3Pi1WmOmxJ0PDnlWT0NMUZ6GRDncKVFPzcUN1lG/oYM
c30Z5kRCSn4v3A4OAXvR352hdbDurbX778r2BOHgzBoaY1qb3sXBy8sYZOA/
N5bX5Aj/TVutvUq0jhscx/hR2d1HeUW8VO1cbIO9b0Fin6BzFZN6E7e2BVGN
838BcDXWLFw9bcXDYJu4Vq42YYHiA+cBBVHhaHAoyrwVSZDe4yyy1hjPe6uY
g1j3WNtmYprvIKPqe6rib9d2yd9BrjgHXy89dlArdLRUPpg3VHUUMARb+SoR
JIq3Das+XV8FhCGdiDaB4sEJOMp57mUxzzsHNLCBbXvRc4pdTWrVBxx/fInA
1B3YwmWK4k7OPCvLyK9+8xEiIHJup0wn7gadgZEWZ5YK7rSk0gcvxH8Dm7Lg
99G/qGWMKyg7e4ZmGxReICUlNwIj95O0UfbxEqedSVl3cwCcn8Rot+Cfa3kg
Lz/N1pdJnOUkoj3Rkz1++OzCJ5HGZZBFy4qA+iuSZ6cn/hA5WnCyf1wlMXR6
t2IX2y48MvJnk9uv4eDK+vCxFbDOYnpulHgmQ98/51Tkq/GsS61OK971Fn+N
sZzl93Xm7QkjNcxVjxRQq4+h4nPGds73SNOJ1EvS5q6KbjTtgwKD/nz+Cugh
kBVLDh5lnaAq3DdQnTgqnD+bZU7uIng22amq4qXJ/ObCn5oHPtXlSLtjVfFD
TfNpoR7dpCc/97TAFOe3Tw+nGDqsiq7Lb1/LFOcyT47C6CokkHQ+6WUnTy0E
6c8WFRAwVKCTNDLedYPv/Z6mV52BZJTjMrsjwCQ1yWAJY3vbNrM+JtsnBzGD
szVtrylEHiJkpScgavIAOgUG18idJtTRj5EdnE0lP/0OmsnOjbQw22arZg1p
NmTwODGvYs6JbyzcgEQP97ucR+/Q8HHCSt9r/BOX/K7Hx8E5UCPGUOLTMpgq
uiVyKElRNPLBh+CIuz2oHbMIp9ac3ARexnUtl8Dc5fzSbQlF8P4Ex//62hfd
49Bv+hTTypn3dLqrAKR5UyZg7ffcwgkCY0jBop4lK33jdD6cfIpbC5nlfpew
h/cRzQ199p2Sg1ULMP+NSjNx+I7d9yHsgFD4v8lIMDnZWtxOT2Iy/RMV1O28
t/mBaui4/82v4XIxCL9VtUKmGQkx7gKG/lkXsvRKEC2WkAJVp5lPw+FXvKqI
Hcv4HEiUtoM+WvkQjjzPXT34Kr2JxY7Pe/1ZZrTZK3Y4z9RA1TcjExu+GzUW
QTfFcb4hm3ToLi+Uqrd6DkEYOEDv5++OY9UOziwXA3fb5JPQXKwHw2djI/J4
EG0XOlVktgaa31DK8SXcLZv/DnIEnsBNIjLfS2VzOLJ2YGApOSfzYbXuJ+CV
1vBumXfc2Mj/E9mrDSPIdPIUrWMDbMHrNVLpDFUSSQObjlg/fHuoDApCYROi
2/oU8jJZ2SVDv6BxpIGPARZtXsjz+/EzedJtpKPaX0B9lvsjlyILpxvneva3
0FkfLuXIcm4HKPeq4sIL2j0UHDFeD4BPTj88BzcqcG715GVGcQgPl8scpfNM
95k7JroqFWsy8pM47jfNneW0DvgSEBIOm3vYkHUgcje90aoFvPw4nSLRNzV/
bniUjnuUg/qQp/z8+mApFCFTyjfENFJLjxXij1RjrAoYIQ0i4xzCEdYY6y31
MgIQ2KdLxEKwNXWGDplJjUN3uZh02yYc5eSBwKgQ3DDa2BN/idaMiZRLCrUD
n1SGNoVylFKCP59G3gu08jf9DS3LkcFchlYlRt+3xWKkJKBowO3Mthb6lYsm
qwUbqR5/duZYbkKJwmtMz+Mkez6DkKKTqA/B4qwBPp9X7T1BjATkYbkozriF
YmqazCJ401ti772qcXRRahfzAQQAaGgg2a8Zz5vxDg2JcJwNVle+bcNIS0Ly
uxoaFq2MUKeds8EJLxfon73xalSy8fhoSxhYO5ZidfvA1p4A+pvgG6V8x6z1
yPTDZBuGuvl4Q1r0UKjRYBDwrhoiftbAM+S/BZDWSxz9Q7SgKU4tHfx2XvkD
CjreSVTeKI7sh+xDoCoNGR4TOdz6MIaUDsgk9kmnR1BacmEw8Xy8e4XNeNzp
8gO2l2c1qGzouKEO4zq8STdRgj1XJAevBGegTxEYXyDfiPcj+9PttOF545Zw
8s/SB24lsKA7rD2pwaROrJPRgw0ExanbzPAOE/WJ100IGsdWg4n3yjln48a8
tJU6eKGNLsm/Zemh54Il00csUw8H1zc99pmugEHDbpkzK7vAMFvmRiHn0uHX
BfMebCm/BrPUSbdIAy/ef5X628v7DrIuvwU/vqSgdqNk9/wgKeGjLZ0j2e0K
VhRV738pQ5cvymdSulO0lJ6NwIlmTfhN0+9uQvzJtiOXIgi4MTOphAFu+vMb
ijCTEtZ/WLhTLOIxm6ukdFls1+0mtBBLptcSsX2dnDaZDk8UOClntjfTSD+s
yqjo00At4lm8rXS4dbkRIfNJri6YAsgPvBtVDQoCmVig220B3NNzNTAa5ISJ
10vEne2cUvFBd3D6+1vqApZJc/DDtJMbZsjuY25wiWOElXmzgJPY4CSCjhan
YJktI5czSHPh1A/ESD64LIXHHI0P0OeZlCl1lPL2oCdrFuJUxWKYf1hWWbQp
478e64XOfQNzUbP8H5JvJWjoAoRt0SrOUMK66zGen3bRHjw+J+vu9ebB9PT0
eiB1psxNC4B+2fWSOKBVvTYofqXyEy7XWJEPGHlnFAMV6vWXZzrDgTQoBBNd
sKx9wHawtVVWuGfFf5rzOSe5q4vzkko2YdYYac1o2ww7BvkmX+nx3nG9Ac0u
CsxKL6zLZiYUjLAJ9FsBs1taLQIaTA8NDN+ztbgEZFEbg9X8H3IbKpBmomEK
HAAgXd4xERXRVekQbPbqW0+Wzuh7PWQ0r1ZMSYf9io0W39tIp5Atd3qwtJ2a
3fMJurOx0XFM5aTzqY9zGcobxHOB5lM+p0VSbNCX5XOdHyomrMBwb3FbJDd8
HuTCoJH04ODeOmRZIphoAPKF/vNJdUkvz4NCI6D36reY9PULhPLBG2cdHerL
Um2KOmOv7UIqrZqFfR4iic4hZ8RoVEXoZ4k7tb/YkdewZ6s+t3LTG/svPirg
fn+3LLEQkMRd+YQVhbWfvLqQ72v2SgJe0J7SxHTH/XUu4dasy10+vTNe0yZc
F6tJjAzFWtzAOaI+/dkben0oI2gHQc0pCHjW6ll0tjoXQkInjfSo+z563rHm
gqcwqwBI7cOCuYJCKw57Pnvfk/P0fckWwl6h8jvAhxQYAEiiHFkx8TFdT+bC
OOcvxGh9TQTVRexCdPtsVmY7DO80awpy4uCenXkK6cQ8PFfmKA6RoxzceAN5
e90DdwzfPg0za7stopm8UzM5PwIcTtiioQfTr8LEZEsbxSfiL3RIbAiEZJOj
KZ1e0ZaHaAkUR81XrbN72ovJwjBVbWEDbVD07Mq8mJRDNO5beRyzvDqTImyq
DsMxmxefLDWZHdmhBnmmjFsciUbnDI9R/Y7qvCUNuXFpTITo4WVZZghdsS62
mNSFnJqMSj1QPPEmBeQ9iscwPNmChH83ZbSCjgmd/QjA+gaDlXziCncZN2+N
RcHkBOwmMAdHiCxFePF6zuIcJIQpdmDJBTkouqs4PhhybZd2zAR4HzQFz+dQ
0shptkIoed9/3r00HdCrAQ2eUMdzYjHtIxC5cP6xGtu7GEvJU1BYhYuD32Ui
p5Ssfgt9F8QWwxP9dOfq7DM3Xwuh4YkI5zBNgQ1oJxDzENforw/a/qdDBNam
fvClmKhuqCYqtks5lrb/GHLdNsP5k4qrlK5f0bByH7V7aBcz1Ll/LrOVEbbl
X2k2ayJ8W62MgWBe4FIz9ygeUHDFp7HD9q8cDfoS8XI6KhrDwpfFUbZlA3sA
wbFDkqK7JOeYp9Gw6FTE5+IHg4M7MdKdSDto3f9UQWzcR1gMpYo01VrkjPJk
FBmgmSNjdvWjWO5P+mYwBmdnnASlXtGHujSXXPkNLpu9UUOpbqDAjYfu0GFj
hC6NxY//9lG6WJuZYGHFAo16RTl4U4MI/1Nv2YZKMJTtLpMsPc1GTZ9K7tgD
m8VPUTJ21IHerKMgd87YumJ6d6jU3LThj0yxLjS+oTSNoGy4ejdVjo/eqUAq
HY1H8NHem9b+Py/SZ+FohRNHDi8UnHYKA9ODdC0FfdVFxW9bpEZQKst6y2TB
ycXO0GAs4wybaZXHx+NtnAyRuqXsM0sIB9dzYuitKPbDLANMzSQYkoqpmznu
7H566AbAkbKgWM8+8mgoge6f1IILE11vDtKYM4AAajIXO5MWVCyXJ0680P6L
EUzusDVLWRuctSYufP6GqNOLXqEIyHgMTyW2WoLFGB3Qky0tvFiHQjpkfMLp
uz4lNWTl9RQbJZUHGBsKyO2W20RPxpp3zFvCeGJ3GKNXsqywXTI5R/EcHKhQ
FHhSVFvXvQlq8zEAdxpbg+5qRLIavYmYc8jSujW4Y/fU6D0D8P7fO/FlDJ1y
q9E2QHAHHmlgRyZu1VhVo1DuR0R8cjYPizN7VkT0XOp/zGEww7cZEJ3N5fE0
bqMBuG4y5lLzAIYlfsUEo1rZIlb2gMXwbZCwFMUNI3yJu6eA2gzROc0Mi2YC
c8j2YJAHxKtcn3JMu3Wg6AG/Mv9wUoVA3M6U2+WAnJ2hHF19Y4l5JDcuoLKu
FAlLZ4U9DOzjarcHVtSZVqN/38AasYeEsUOJ7R61nUY2vtRFhaPGmVPUIzIX
sIB/l4aw/cmPTRTosgjxLgSigy5QnSeGSpMAeI8HfRvO7gtCv+0DF7bQmZpo
P8g/tBOdT8BShykOZH6IuLnZXhfF5BBtIWk8IzDVgZ90CRmYetPj/exAICE5
7ALNWa+aMVdxYqBC8Uvli2Ugvq8apWPGA0BRoWF3cVZEaOpB9yhlbDi6mZlP
ZUZFswxv9H2XeeawDTUKsfdHahC83hZX4czUb+EqnKyCXEZAuv/yxk8XQegE
gmXuzuNs50aTmnPtwSf3c9ykatQF+nasTaoHgAVveJfZzwCMJSx6dGoV87Fo
o++56cPfI7TF+FdfH+6sIvG0pi5D8LsvK+NOxHKlI73fxDPwFVQNyUGoH/1X
nzkeeTY+ohbQ2z8NQElapfGHu0yprFsjaHb7hm3nH6w/5YI2SxJNprCV8Kbs
OaDTkXaF9qViGBvSRH/wNyOkztlIjRTITS4rR5e0gKRdC+/JpKBXcmBSMsB/
3nq6cvIGvR7G/BXfZveXO8Sjgg4AYM+7EFV/RG7/IqiEhRwJkV469Qukn2yM
/nY1rWYz/oAQPS8u3GqUCfjgoVcIhl14GoDk1l9/LTufRD8M9M7qzh+gxV0a
TCRicsKWc4tuhHSURwrbBhZcw3VgKvyf9AncuVa8N0ngnrzgXVsxp08hTTxo
jyCAMiDS+XV+0iH4WAtvQyAY7/3fDd2ik0M+xDl4Byuh/SveqtMfnG84WxaD
y4eRaTzog4+Oszpjn+d5VW0kXGgC+shrQO7zJK29oAqSVb7a9qvbYIcvO9CA
i4hvsZbcV474amsopa901SnyyEps1X2hxZzqbckCBUU5Yy+iHITY9n1RjqOd
QCICdNKl6dkoNUR6x8cyOGDcmeOqAamjoAzJ5lkAiGnEN7P5gfE8G5asV9LY
soBrlYkivDq1HYmp0YHi/uF7e3gsu3PDYZzUiEC8Nakt4yViB599DH28ZGAL
oU7Hhbu6exLvFDJuFONx3c88e2ogbTzAn3cifsgo49KZQkz45zbiExq7HnAd
jJniVdGrO5/f0o6EGxR9z031gFC5a9d++f5rKTARNer1dmnNtg2TAf3ccwgq
5JrWOwznZG0kPKIvsOvRVucInbieNff9vxmul5puYXhSL+BNy8MQQ3z4Xy2j
tOsMN9lI6YGYQZlpKoijfOznhJhFrWU5qB/V3taWtgKvHZyv4WZUPAwrGYKq
ESFYvMoEjTdBAtH1UyItBZN3EuHp24pSgG0eQ/gO5rQ3u7UeOFe1iTRfV4Oz
A7MR+VtcADdtOSKDlH2Y395UJxo1pvjkB+ytjgzT/cIEN6dC8PyotyVlhTDX
FOxBhNka201C93Hcm1nV787apCHzMKCBx5qFq/pTsr5KB3ijHON/b2LhW/91
jQfVcO/C7yk0ujP2pVTfM6kGWVB9l7SUA/8ixagvH7GQLq8pqU+jeN+P0Gju
Pm4y8iqOyzMf4H8X5t5gCNxmQw6pToi0m3N4W5aKWvs6iaLIscgZQO1NEgOF
v3KNudVEa9tlidFcE9EGPWNUK49Qqg2zcuWpAwZ77yzEiTzc1DxYQHGTKQUZ
bPQGyrfT88/PdaKd2TfOYRgBVJv/faopfFzI4dFXeWgN19ZldcXdk1/gkr+n
pUFqYftLgGX+hWrHBkSxHaz+zpTLE6QVajRMfRLeLwQ8Q7q6HOvfmtmYKN3F
++fEqQk8dpvQneNyH8QVX9TbxtJROypCAK69fJXmZYXBOzdI+fC3wOMZ714w
OJmfzb7yUZ8q7zwAYZFqMdZrLYVDz6acUMcS78ljMuaYE6IrygWDYtJaw3O7
Plxoe/OmPUkjJfSphrQFse/SpdVaB1PyGCMPWkQr6TPh18V7no+DzcaspzNO
O2Nwm7vPWfYpLFs90oNEWiNvnU/oZfpH3kU+1xCaXKFITlt/0xwedV8x2/bt
2PJr+OhOGH4X8UfFgKCRf80NZvLbFBVgCy8xneb1E+qvfrSO4OAW8VY65tf/
LPdYX7WIm08Xti1qVpX2pNk/hIXzNaTVyN7zr8Lur4p7VVRXHrByJphjIpbZ
UyT9FD0nqLZE04PWfRR2/ZIzptd2Rs7ZqZYwNL0QR3AnMWabwG8dKshOd6di
+m0nak3uQEh9i7AehwtL42W/4ex+nf0ydJ5c+T0trioHF0hbU62so6xhsGgr
iqp3IBWAsLBI9GObUhTKtq/gS47I1Zwq8l8f/cIE1Blg40f52wYWqbIV8vId
kMtIBJwrrY9Bhhl/A7hX3AvuPf2uxddWBY9J6S8/AATqSlZh56aVGmLMb6x+
/4cYCtjpLY1X/upxsrZob4fU1ZDPzrsfGpXmZ33hduQBhjcntDNTQqXJ6EvW
kNr40a5Z+e17GEJYYB7lVLUa/x+7XDZfRXD++x6eMLlLnWIbDs3F3LmOBlSn
i245wqYA3l6JOGjC/LtKyDI78r8ifNUQjWR5Ng1c17z3vsYraY8LiQG8OwbY
QIiV+lxbKw7S5Mtf+X5HiBtmW6Q5QfezbGUkdQYUORq092RDKspEvXXEWEe0
A/8wEXvrTzg+YlUTm5sG6sDvsuDr90lHvnS/v1s7L9ULY4g5dTFOcHeqkRhc
nPNFva5sMSHhJCcUOx/STtE6HVmyvhBZ1I+ZPRXJYWnTgEtf/Z4cEVwUtmqX
R7nrlZ0313EVCDUL+JIMaFEwBpp53dhS9F96RHLGkB/DIrRn9U7vMJ0R3Ua8
gt++kha7LFHoFgeox8KGyYZ5yF0NUTzqBYDex07MmO/mBBDkNJBY4YWgcxNr
DzHW+UxWUm/MMbUVt6VWZa383P969lvXkgBkypkmo8uZbYMpaD+dR+aQLa7j
Ing5VthoxeXQ0zUOYE05/B2AHymH26Kptb7349G9pIHuxIVhdR3F+4zB7dM0
k/CvoFhlySt0uepkAo1oXWnGy03afMvzZnO0PDascLtSuQSbwjuH9O5HJPVP
yVhMeMNGLHi7DGvdGV/Ukx+eDcLRj/6+fXGUFrGYoZ1uCvlgMMXxBRXMaumR
9kq2iHOI8AZvwVdQpg2ZtJ1GE3S4RZRlAYfEkLEKcc1fNMHhjBlKp1CsNAG0
CXkAmbbFbuRoyl++riOTyZ/nrWosbItlpCnkKR+FSI5wykXBY/tPTQUKemHf
EMfvuelG9m3Z5MF96lXy5gPpQgq2YeYK0eubtnQpWaC70XsSzY4fT+F9QT0i
YMHgu7r01w2ym6XaV/fSI8OcETwJ4I9EnoYbk17mhkzEnhazlOfLSG4dN380
ldiMNeGzyTAcvylxcbJw8vTN9x2S8Uz2KlOGaaVUIXocrq2+00bvuI9f2Y8B
M5pAQXUHhmPOTGAHQrYFF/OFBjimT/9XJLJOqyhXfcFmHcCbVz/KStaKsbiM
SMifllfuFMREFEa7q4c+WSuernof/zdfFZ0j58XqhlDA90i/y1EvwLQyrDbw
pGfTWnWCNODG4bLMx7iwHkme2E1G9u+OaLQKPDDFyh2bEGVVXVPwOEzWe9E3
cZf2K6u0acQhWyfn8WRqG9fkOWiWIn3Jr5fEit6AWmUSvd3eG3XVyAWBU2Jt
NIlohwsNbBpl/TNHwAq+4iKR6Pif3pr6tcYQ4KCo9/Srqc0vIOgcKHwUnwSe
GD49BDkM0SHm64el/EgWUode1TOnpFZ2vC2BjuMVEtXQCNA9L7UeXzXMLVvZ
8YVCBVnaTXOcP6rJmXgGxWlypL9Vz2+QHTxYuNyiGN6VzuFZUX+61pJp1gM/
dm2FlD88oMa4PyCe4tkUMQJAknInoaBArsZw2LpCO150eDOI8gyC71xpYLX1
Kac1VaX7xAAX3iRsqQsKMmjGz4QNLoGbwqAPf6Ai1hlR5VrwxM8YoYmR2Fb/
GgZ9LNpQw2k/T8/+PvlY9UUX3uysp+OpRcT2++vJYFvJTyDFHE4VngfJlnRd
ZTn3TimVoq9OulSF2JAQejAsFlHctquxzuKWfrLabPskBT6NZUFjjfHH3D+H
HhYUYL1mfT6IRSnFCBO9R3M+EdZT14Oghx0QW5cvV0xextPkQsP5S4Y/7lcv
Y6G4jbDq49pYZjuzy0YX5WNNwIVHKHRhMDEYfqYLrackjjHlsXTVkd1Dy7xU
tg2JANJrLyZr9b7UX8ssVPY+3J4cyBRD4IOXj8wsWye/81+C+79pwnUl0VWz
h+Z2w+3y+obo+n69NHXytg5xYElZ57cVLnDHccQCGh5uEVJ7ep6AWogwFTJy
QDCeBxs1le5P33JcDtZxB0OrQLIVhbWBUT8cBBObDf7mPW5ma2P3DbWRSNPo
Slhr7Fm74k4WQvGswt5zz1XsCSnEl4N8MF1snMsFPp+DvJc0jK8hrDD6WWVU
bzsyVxOHvmWQ7dQl/9SjpGdnTEKtuXhiWTsM+RIvqStBCCut1oPEi+yncdCc
hZDr5zr0kpq/vJtSEPR3fHcHwiQ26fcELebUgvBOLYN2vx9eBm2KzS9M9EuK
NTSY9ufyfVn1kZNW1trFs9WwJJVvdegpTpAM4fcuO9tMht1HOjH3InfbcsYt
D0i1yOhOF7aN9H907zeMq8bTI3qSOE8vOb7UT4Lp+ePIOK6+Jy4Xuvw2DXla
9XytbPiniLuI0l+l+JDP8GE3w5XdKto/MV4v2bax0oW9Mp92iZgG7aT59vHs
aYy11V0AJdFUwML43E3R24+Qq0AnlmJKtc+Nn6Rd1ucFMxOajkLC6LY83xnL
77ZDxEfm1uwysWIgRyEf4UX++dDorsb0h/nEvU1sCXTXNgJO82rdEYQUp2Kr
Nb38mvTiXV/HyKhlN1LDOuqOpem2Ig0swqPlmIOJ6HXk/jdNV0XedVs3vPW1
Z5snVEUE+bfDGd9Q8ySCYCosbPenP0sqHDCD7xntTFmKcy73AcsTL0zJ8O9c
RqCG01tjvTT3JlMobBDfa7wMELctO8quwXOgZoAtLtjg33fJNBe37vX8n/b7
e1kztFc80l/IOllBwNgIJ1roluQThzV1dywPAxV/AO7Rk+LTd9hHdu8NstxK
6LEcSduML1LT03YFQ6BE3b3qwieuDQznHpzBVwT5FlP9wI0QbZxa/fIUGfJv
PyLyY+uqZsg5JsKFtGPSBXtp/2RZxR/eF01U/tqhxVZAgOhUqmBv12W7EGf7
3EEqG9p62VOkbPKXK1MXYEIpw/G4inJRdJuvPu4yQhcVaCtesnlr3G0WooCJ
MbpVddrd0HxaYhGNUdVBuIyZx3H0QRP/PLGDLLz7KAWLwJ4O1xnq0yCpkf/l
g4R1DPQl3oKC8kU339bY5tVf9jGWLz0ciGjwzEV41YP2lZDiIwrJmIuZenvE
iVaq5Qw055Ql5J47v2b6Qq0NPe4Su4Edc7J/7+JZzZMixo5+QoaG7J3y5LBY
eDZu4oKKVB0rZzQgHfiUT6D36Wkyf19BtMoU8gmaiw0Qch+bSgS56jbOvKbK
v6ks8RyQvXAIQEKe0dwxGac6nnHjPdbQeg8UrkBe0GHi6Qn2RPbI9G6X2AxZ
F0IR+CFiUDixYQCu5Qo8uxyE/XsUO5CCsPWR68qUZndisXqhYJHfFvKmn6gq
6OuM+is8d4UjIMBGMa/AWdj2Sh45aa+C08JONzEMWB8ons+8odZ+iC17K7dm
jasdwSRljZbWwjlbtvRkRxRRRtaS+bSx2X67cjQ03Dd2eVXgcZaOY7aVLWV/
jAK46lHmJ4xV+FU0HkPHgy8E6YGlgD/6gOK0eUyltBrhxJF3767Wg4M1pM+p
iDGKZDp736JUNG6QzRAtE8GxRR7Zd7PM8hcYHXQCEJwF/VaSctkXsTDmsHsT
f58P3XlbbsD2Mpasgadr+zGP0ZBk1UiBhk3ZdfHITumzbxDUyIqOV3VAr65r
EOots/tE0jmt8NQHeydRlsUfHVGCrdzoe7yR3uFde83esvkwTnxJKxKHMlGI
/abhhGKbWsL9lwP7Jn7DjT653/dTS/4uD+ucny2hbcOcPcnQcQr46HHB8GWB
d0/pyj32TSw9Du23iz8P2DpC4TUXEWjQ+pTmRMs67rGWpquWzhR6i1Q6hrYQ
YpeQWvZo9Nz41oia+WXslp8aRnyD9X9C5tiZSknWe5EHNeg+xR6jjaoOR7MG
WFO34hxEkNo71FxJDVUkazki0n8Mtk3xttsqy2cwOn1rpG7kpHfjBUUJPf7t
AR1q/pxxi6h88im3GYfBisLkj68r58Osq2aTGltchrd7yX9g27pQPhLVl+Nv
UlAhQU87PaqtSyY0tVzSLEmwJ69iGn2qvfnzrdWjH35Av3qdhGP/RvCzSrBw
tgKzDT9ChKPGq6gW/rDAKhyeKuMTxombHVEKNQDE+wdyqhODca6Y9Q4dQz/f
v9eUVQ94usNoocer+5za5UNDPdcvf+pS8uwBpEumGOif7013ooEayYUxTeJU
CZ3kNYYXWXV8M6jL0IQSFQyCB8XaMAj6cpuVeJk0US/pLEFBI6fy0Aykgbtm
cRfHG1uIgmlJfkD/S6X/uIVwb2SftONJM9a7b6uT3KxbzOzodV93J5N9oO8T
jtx7Hei4GgA9PDav8qkM5Rjja3h3m2fX/mhfGckJ+JOSu6MwYsK1opf5aKzt
Z3QBT394R0wINgEdNVtIVI36ls3OGCtMHUuEJ37BXZvkRTMLmJlsGP0B+tIk
X5tRA8Uun3N/mITj/dZaxTij+Wd3giXqht16PxiAZyspSLNfeRhzxe3by4/V
CvT59wn2iuHb1ceLIfxThq2T2pQK21tJPYeUqWczy03K3A3/BuxQbCStuDWn
/LpImRxNvqEIvBOEhxNeaGgBcVkEMZ35iWaNGfnofgSFpaRN8upHcx0ybYx1
x/jg5T114Id2cQ5aqyClKnYMSa/1W+nKYnkUFmPiS9Llgs26pBxbx6Q+WS9n
dMJVZRfrqb0FS+SgA69gJwzyUqaE9mYAZ86ALrETXwoGsYHnbvhgr2/HVDwg
B2ZjV7SW8B+gqLAsTtCUK5zfW6FignHAFOSDnoejC5dvQScB+n2ZebQmlkeN
N7zUPlkj0z3Vp7PuUJl+q2MfFgf9UAddAnA0thSiaVvhXDdoB6+Gd9aYWfh6
by1AYYe9qErQgkavgcXIMEtuqRrIlke6gazxM4mEvj2a8dEJg55M7GKVRIX3
GLkYBdREdmrsXlkinFsqKv0IIgkq7TUvnlUO2zr5rVDatoMwgAs6EXIQrhse
/uTty6sHuUAtDBvUTXuA9LV0Ig0TKrQMq8A5KA8jstmcpCDJ79caHcAyEqe7
DZYZfs63Ix4xSbTGMdHb24TDY0SabkMmE1ONJlwNpSTLJ0Lg0pvSaWcpIziP
3Y6beQRrnZsYdyLZaFcONk1qodMzmMlIu9CdMtVSpVQXM/jjJn/65BY6h2l1
aFb3r4HWGOxARg9pmwilrSVSjziopiKcf6UJR34wEx0ex4dmw75Wr5HCTBER
kYbwpKqUm1j3+sVh5fubYBItG7XUxnTFOp5tviyNFJ/GEq4/8REaGyc0+b2L
yRfsrbu9VzOOT8Cwy1OkWTKXjlH7lKIcfCkz2JmyypVCE2TmrKgKrVKMwuh1
3lEpWzdODMv2DA6EqEze3ysfqMUqRNAeusTAWHnMLpKa6cTkNFGpZiCScSix
7XNj8xUxG591Wsr0nB0VuA/CmusRuFiWnF8h72U6LjuyiIToylHhJCla/wv0
KSjV+nP1WKI/Qr/e9iJYgr+CWG4rwymFdTX7uRLjWtx962alddKfaYAeZRRm
tTG1pI4a4Ucj/3rUtMMNlTnEt6CvXjTuqykcan5Yr9Y8JdwyTyJQEWoRIPLN
pNdJ3bVFiq6BH86LQZFiIcBCGoNFif50tu15ea9j8sJZ7/90eY8b1suxS591
UZ62u7hFh2CW6/hkQE7NGQcOE9Azx7CUTY6trjgA+HM6KUdyhaFI5lY1a56b
5f0sygslFRgtd8q8sjq6aslHNuO3KqdmLGx0TPGn9YiTf0Vp1wiZjbF32wA4
Ya4bKSD9ZiU1hZ2yEbwlCqisccTBBEFx+52KZVbsCULLZ5v4jj9rtLAZsOBh
UxRR2Q2EEnNNcvplFFHNj199I8UNeFY/srLQSMjCrqsnNU97i6o2zBIytDaw
nkMOxcBUQH6LS74cBqnSqIVFSkwRKmsHe78W1DZGNSnwuePGjoCZfp5UobYX
cXHe+079jiBxERDrDZPt5AT7Xf35o8fQ6XH1pY6Cd5KSxt84r7LuMqDItUyZ
4tnedMAI9hGYmRqN5Qs9OAm0g9ZxYyRs6oTxtjzt/juctBN2xtC/04YcdWlO
6GZK5QDniVsuqhaFpGfY3TCykUsULd01RRnnHdQPQn0shejecwLD2nN1oHy0
jvM9tH6O6ETebnmMAPcaLoKv+8YvYmPHlNKWPntjHGk6aMqJzjd4iOkRA9XK
q/AQupXrR3F7vyTE5smp8Xf/gnBzC7tZGcGo8uF+bcK/4vbNBE4TTAgD8tGN
4ajtNQ11opiP6uE76YFLbYocXJ2NIzX7Ced3HEdxnPvTBkY2oD2QLJTGMPsy
slhQlygHjHQIiTTQfYKysNaoA0O2DDWIgDs1vYQfrcP0U1iGQYJbfzSjRigm
jNgReeyCnRCI8Xjk+Jj+TCY9BtxyTc+j5mx2kUZW4aIdsVW9MZX3CiMPgFZM
Dv3IWC8G75LX4Q5O5VJDhTSvYN2Ebea9fCfCziyoc1lpg6miOaTMFakKiaFq
HBXyASDlUMPQ50Hs6/Jqa6mg4LNt5oYcUBZQhNJQu3OW8IHQAZn68S0Fh1hC
Mi+xy8LyTzJar+NvT9wDdrcIMw0gjMhEjVwnJiQ8+ldx3FuNheXD+1S4AtiN
e04ekuYc6oPjO+KUOQaBxCB8Roe6djiIEHrsIHe1o0B2Ptfvg0P3vpYGJtZT
89rWvoaXi3cgIxSBrxqXUSspoXUTT10bXrWQCBLc7aMceYyOfX9gZ7i5AKt+
bI8UiHAopegPTz66+5lVKe2sCe+a7c34iB4cFNgtxXQGlIqcg17T43EgChoE
NG5pRxh1UWvjdO7edg01R/ewBCpHxUmyIG98Jc3XEM5DVwGANH5zHvCQU0qR
y6cW06XwkfFlvsq2ZUaY4NkFtdFRnk1BBtcUNrMOfvEw1z7cN5sUb4qcdVrc
2lKlH6qrwB0UKUiRUMoFtn48CQ7CQfgDDmyLYaRRsEGmUGjpKQ7d5vElF9Wc
ng81FaKnSeXSRzwpCo13FQmOkAfqrkQK7qTMmoNrNap4cGUJpiNS9psf+5vJ
Qz0K0jBFCN5SxTBD02nSt+q6We//l16Izquze6042tMPfOsRIdHuELsclrNz
24XQ9dQNcNFs6yK3nSqqfLwQtqaw6A/XL3lXssMOxfv44Km5JgOrpDLHY+pv
4YaNCQsXdYQHTchrQ3xZqD6XTXmn3dGspplOlc1fTst3KKoxQTewoF4AmUCA
CQhCIxBYm5z61NitfkHN+sPByvX2g+pWVp/KMuxyn6MqdidoWsbUpQrVfX3r
DiH25Q/flEwy4cWpgU7wr92n1NVuRoY6FxKhxJ6wqn9MyNzP5CyKryxTZEJ9
XaMKpo2GT9RC3W+Yx9I34/bH9oky2W70bnEV7zdvshET3s/B1cZwy3FzzJJA
XsPjDsQsnQ89xVALd6+HXdzVO5AD6Y6Uu7MosyinyjwvVHWdeNleFkkWCC2x
nPNLP5ge2ck42Azvg0KTphfOpvWKvSL9lPh/piyfOEWXVE/vclZELDnlUmka
TloYoIgK7+0PIKKs2bPyhRp+XMlZABqgyovg42PQCslWdxkM1+pHe9IHHOFo
mjbokkL4mcLTjJlO5OZ1rKs3eX/yUrgs2I9vR6Ps88JdJu9CLqZKF03/OxOv
IKVnlwhlS+oPkmHk3PfOyf3lLca1dskYazhF78B3OwOaSZJcdHcJfQEnTAqd
q1c1JcErXOC+CBgncK5ehRARbq8UxR9hQ9Oam6vgHI//xQoE2PYmBl5WuEHI
ocNaa2jT0hJCHcKpF/QMbobqsrs+pNUsHaJCGW0CokcSk3g5dJ5/tgVmf5mk
9Zuk+2mBqQYJ6XOyx0n56JFzQ+L8RMFucBXIjeb1qvzrYoiu1HxBLAvHBnvb
k2qkFbX2Fb7mwi0Up7rBi/IaW3R++Cx9EqE7nioaiUzNi8ge65QKtq8VaLOI
Jog9rShOIr16aRSqleslf7ahFn8qAohIXgStilwvKmRLtpQZHHIujDKqAzRK
1HrqJjV5wbnBnDSrXfA/0RvYjMpWsthVWg0dj/P86O8pAFQwV/sR5JGoHbml
yaCE9UbXQXa4bYDbnURiyZga0UtlmmH06tYtqurW5TYvi47YSe3PMGbcgtra
uBcXETmNep+nceHjq9zniLzIU9WXPjRKhUbz4YJGSReCO1ynNECvTnmlRYT9
MMnjf++i64OPRnyIpEMdPbA4RiXV7FysXGw/mfx6OH62XfgahvGOHqNgWUJE
92ngHe8ohhN0GP9a6wKGNo5oRTyVlf16SCJQz2aii6TaW18Bkk6f/2dnrFyh
ZxPgf/kyTnTxhdfsmhYv+bSYhNz+GGCp8zmNhYU75R4WK8aaBUfhMNA7bPU9
QvY7JHqy0tortchENIGZQmwK28Zk7bW78dJ5iGf0fNZwJDUCJZdWrH/6cnii
1wAB/vAzd4tYBcakF9RxJcWUQnIowKdY0B+vNcWp49FoXL1f8898WEGjT0G9
VChWztB+sL4KrA5Z3sHYcQbjPfgLpE67oFtVlC9ZaV/GwIxuSRg9+XvT8zIK
T+iTLhMqtcR412eHsOfve4tXiY84bo77QyOh7Re851dqDh3x0Nb85GAywHmF
24JHAaMartAjVYhrFAR4uj40vtfhe3zoq060I2E8ihUHl+c0fNU8k/nNokvR
pT7PrNTYuz9qHP4D4pBASzXBBMxxj8FpiIapSxgCJaOEWN8MwbK1N6N/qXbU
MPyyJKnkjN9WvUtQSlhFBLGV58MedF1fePdiu+6w8RTm5X6ng2Cjv3FkCAmE
PzRXxIhNxQRlCKxqg1SHkm/G2Y7hN+fE0CqjySvWMaA9lcpKm7EiT4NYEdWe
GkzYj38NSeL9EVubTbA3uL0yUrsTmef5OSh8K6G0Z5mHcwdUQTuLuaIBaArd
T9ssWeH5+DDBm9rd5TfE6x0BFVDdZTq9+ZXKkplZL/8t5SnPdFhN1+I0hTsG
O0adRD9nkZCuJwgZm5VKmL/X6AuiyYYeVY6zrnSWgMiMfH+GQ9DoAa6Om9iS
DZPCnH6tmg407J0x0exDx+FL++H1SAzGC2tMYpPvaAw75MEjHeJ59xzeBNmd
3pQALhDKvemGc5IOTzttXGBF1CmUl/XvYq+RLLjN7u6ztdfIDc64/tSrA1JP
wiixLdzV91vgvUtm3dlenJVN8bvASqQn5Gh/oz9FyaX8jH3aLw/xukF2F9Kl
0Z5PKc6oF14C/UNnr1+az3xa6FgzNOxBKRtw19aPZQdx5iuVCqN6uwdAKSm9
PRI9gd1gavZHVdLiclsSKQZni6OeXSrLaNCPKO1rYX04eyiz2t5Sa/AOy3VC
2Kn7vjVs4PuimblIHSivDZqTod+DzbfYcRL9OurTGTjH3E9Qk+jU0kR0vJY9
e/eBHmp3Uq4FB8a7farZQ9Vl55tQ7tgmwE8WsB9+kHx1Z8HPQgiLKIVsIn34
vK8lzFspsNlp+bwyjNajNm7xs8BrZv+BU6VOTnnkPpkzN473ePHC5mcoPaOs
JaJEbfCJr58nroryU1KLX6+VUdNpEQs1ONbsxqNTPkgu8/zdlK7a0EkLLVNr
3avZtaUfQkk9R7L8K3ESHeH/QAddyGtcpCkZ0gbO8evT6UD2DHjc8K05lf3S
V7c+Gw0yvVlOu0TkA86u2nmJswuWTJOGjqQu0gHCzmYwBDN39DDm4yP+1ScU
Y512+PiOEFPTsj6p8osVugpWEvAmnLuoWgl8unIMSH2mhUeN5IVNNr8tpZXE
9C/ei08uJv2pj9vsmCGsOB96KYJqh++N2XCcW+GnDYYe4tqS/uzBjISk2AGR
YLv6VvW7raXEA+p5Nx17ZAp/s+16AG+DMme0i+7A6GxRx/u2AgkEHdN8lFs2
jkIJMK/nZQ64r330G1xrPQs8K6xXTm9KpnSdzj5doz9Ad6stGHnMb9qQ6fem
n6rY+OLBwTlF6Q3+WDm90FQbZCyt0bam7GXp3XGwa5qgYh2Hd4H59S+X6fCo
nwyXozDPo0LEYBdF5byguiv9j83xNyvVMaagsNyfMCA2VtgricSaG+YtXrtQ
m1u41Mx9mzDoZ8e3TvCPmb2AXBPyfc+JO/u0qcx6on1aOkjC/wwQ1bvjSI4J
3+ev24E2w6G9q9J6yd/EE/2r8ko6KQh7y0m2xcx+1wVN2GMGsX+HzO+UDdgy
GJhG5Fy96Es3Bw79+XIbldMOeGVm695WEfW2LDweAzFvhMEDbcyCtbup34UW
vcOS0z5zGiG1UD05mZCeUeZbpeMCpTUF/Tx2bGMSqF6pXm9y5R4yzB9IoPmC
ax1THeikv7Z0ogaZu38qg84+YO5xAVeNsDhr7xhuh9NWak7l6mCZ/aCWpL25
E3XaEF57Vw9CwCs9Jab7Uc4LazqvM8Cgz7fQpTsGR60HqYSB2y2APJ2af4MQ
6p5XFDsFaDY+wQopmLGOS7OlBfYTFlwMph/h320S/hvpIhzyoRdTmvd/Uuoh
pLGJeN4gjqg0jppU3JLn5JEKQX0z07dxiEGwSagnzdW0BUZ7wnn50PWwkdW3
9kQS0/FEjd+fl6EIcGswPbi5evDOoR79KG6e+jwNfX4acQAYVsDazlHtrOf0
H8cSKYfbdBlrrZfgq86WGOZUtzqCenNYv0PafavjaWkLrtMGOwhDFYHWrF6z
sawTAGtHAVmMrYLIMdJ4eNzPsSQEW6oOx+ebCsT5GSA5sT9LIpSp9Gog3Z4x
wJnuIB9RWqLm1FrUVbgDqq0MWbXwBp5zLxsGhrCnyoiyxrgG/F4MVuUL3Zv7
RKDWODJXlLojaQ149K4KQcbHZy4ElhazZDI9EYpMqFMsDX4ICbv7LumER+zU
nWG26dI/oM32j1sB9+eIlHUDBHX79XZAGj5BFcHzF8elFj1ujf6KWp5wtFK4
JE47OorewjyzifP4ZER4IcvezOTzhy8COjzgDK/yYzelmJOGt6NBgO1qfJab
tp9MRgE18zkLWgNw8V3pvRoe6sCbnX7V+x1BAccSfXEw4CcJNT+8TPTl4tET
9ces+wL63040NMYvxaqhgHLrxdsWONNkIvH/bhKJipLq+MpJZyFtJ6lV+sxG
DqRGbhmgYCJWYhLC4Sx03DdyVaILmLS/KbQ7PuZOAa5jAGRAYCbaHPE9krMK
zSTdII83vOJDZr0Si8e4zgLXi1o3BuhKpX1d5CG7z3opHcd15HsSOtLgYX7j
chjaGkkJUI/4wNc1iJGtFbqyGbjwo6dp0hOCKWxqoR2hxvsEOgNs6F82KnaZ
80RI7pECwb4WC3iYk8qYrVltI/kmb4e7WD6SS+QYH4JuEqv91vdkudM6rC2g
M4Uz7zVNmO0cvjHLNYMmwOHeZIo8cMGo2LiDXRuneQyWuKvCWPeywA00t9HH
br9sE/N18IWpoRJaKV373YqgGXingWpwnyuY7+X8/TVPMB6TQEiKtUoa9PtG
K73rnAzMYqEvirkvtlT9WTUxo6GzBqBLdTEmjIrhp2SAlFYo74BfoEdUrgfE
2LteDcwVC8gEABsJo+kjx13Y0C6nHWI/0y2VIKmR+sGn+MPNC7EzdiuD75yZ
QQfzgAIXdIjAR9boS1kWLRrpQSYKI3iq7XDbdhJrF8KDOn7JefFUQ9NYD6bI
38yMfDu6S0jkA2H6P6wKXa3pSWiDbXaGnKMGyN2xcMk2S4FiSM9ilsLVl2qY
nkbrHtwbH9f/9Id+vFqtCxZCxlcKYYzdZRf++c8CgqUEoGSeI4fSjqe55WeD
o8op6NSAar4r5U9f0R5kTT0mP6jVtGLIhcwpLwNYscQDMHtMsHIzbURPFSW3
HYVM9PyV9QoJGdYmohcUZBQJqcog5lU7g0P2hlKWW+jcCVcaLmdtUKQ04zUJ
+CklAAqlad9ZKqHZsgS6eNUnBISPctwncZ4vShfi7HxkJZ+7DDHK+eMfYxZ8
tX248O0eDLGdfgxrtkAxcFm2A6yGtLw/06alaxmqXsHa+a1QFwwhJBgq1kMP
6poIpEXtktBNWKFp/PyL+6HvE0EQmZr0MFHD3jfxzI8sfG80o1jWEzLxxIkB
IoyFa6QCspv+3K+EslwPzWd8QoctB2m9tcUO0w5WHpg+JxHk39aDIzs8KQy0
QCwiBTfriwzl/r4WbqaHD+/1+lfC9wvIkPmnlrUKJps+3BqgtnhLgMt8JyjM
ACSEIh6vpuhafXtBvuq+J+BqsOM/9ODnRwCfA9KK0x8mKUUWFDfxp/kYmSi5
NUfyH6BGVzRTVPLIHX8pGIWsIXz4fA38aJBYpbroKUAq8yiRWFji6sKPV+bs
A4mqSsWwACLuriMYSTRb9N2fc6iMmYU+fYmSgUSo18y+VtshS0tgAt4X7suz
aAWita8QIAqNkaye44DbMxOslaBO0to/8lexiqUakz48YZDdOS7Hs1TSMGHy
Ps4EZzkls5vvygKalLDdkM6RtPfvul8hsSlssQ8unZHC6imedzCNRf0nUQDJ
bpdoawujas2hvebPCtvhWCIwMXBJSUMnRRMcjzKh0KhN0eRqnYgd0SQGHGhe
JhApS0/ESzp/wkv1MVjtKEqiInMrESKPqdyIglRK/9f1zO06b9ymZ5m9ivfy
fHZLLgjyoXuIxaj2maxYrFJAAk0hnvowVt/LjDJTBGqlyY3Kl8+NzKfDkDNM
xcmc3+4p+EZiFBz0mlL6mTlMcHSQUWHhirTSOBINApLWxcmi4FADxJPOkIl/
54awWQtu6xhzWMMf9MKL0vrBaF9HbRny6oI9YAxOot77KX4oDgFa0oqvPHJD
87jrsGgr9jIA+ycqCi8wMJwnxz+OGJWX5X9jD3dqnVP/MJ7VEZJXnn8rh/9Y
nuxdLADMzhxIHpYok/xmuQJI4IgOyLbeo+oWmi5BxwPKkpL/vKU1woBA4/Gb
ZWoJ7RX/UgtX4dmNuoyHSX0amxz2mREN39HAQVgAQHaowV3pVvuJJDqT1Rm/
4x2gn3qHIsIGrdTGyRtmSuZH0JCrDOvmXurqnAVZpdYxo1ClycOCLyoEfLfI
RCtnLNOBQEEtkhLY3MQ9N1Yhs7IVF7/7Zsqq0mVKDPcD1UT8OBR3eu11soLA
pfLaaNGsAilIxhlRNxtzFJlJbh+mpfk+UmXhwCcWKVP0R63LRX1B1nlVsK6j
fUZUA72tW8OhGrTiaiHLJw18WfW2QJi2mFB42yoovRk3tZ4gGVcTz+eoQCC5
G85/pFGXjBh6ZlhFSd3vtz4W+/r+nMekFdyB8sPmdCrOjrcNqXWFKN5DOiE9
7XyxF2t6SdWsYzHrCt0hgY5Bql89r/iNfOa8wij7nuC/UBASzJq368MQK3kn
rIxcaPKHl2JB15crvE1z3VnwTEDNTHKsVPdZ9yY027ueyYHT8eevIcxY2EEa
8RcljdUVT3d78LC6FOz7ZbrR/wyZuDyzGmMprJoX+zuf/sC2Yidkteicf6oj
gapZkz8ZFI+Q7B9WgtlY87dT4P2gdGsQUSwkK4yrnP4qgeT368ByzJxrTwJ1
5bULnCLUvpVmXYe9LAze6EE+TvAPUS7jsboNrgo2h/HJAU3gS4wZ/meBB1sN
LD3yUMLiz7Doiud/7Ar+LkZg+/cl6kbRybRTI4PzsBzh7ap4QrHOCnh5+rqm
PmEmUPZeoYU11JBS0tNdr8idpES8WAOrvdDg/zqCKBk++oeNDG+MVmXfY8sN
BvmnuQpOhIrVlnb6QrhRelKi++h1P6cxqsenW6Nw/BC/Q+80urBC4zBRmsoa
+TLd4yE1eV5fsKaj7d/tSnbJ939oz6NOJirkSb/DCZCInPNcd6TafkVIYEZB
pSdyjZZvMsk9XrxicMtjsnr1FSUe525VkzPhtJnTZAXCpO3RHhLBBmVZz07h
Iy3nOyDvqdvQ/C/z14ysw79OYBG9xVa4EgJpTVgr9+8D6RW47Raety+UNxfZ
3Q+Jd4fennLOS7m9Liq/73gYI3yzRd4Eqia3pGYbZrV6Hy/gYNGdCPwb52me
v96dZqxxeSCBeGoKfi6WzBLsrEnezWWGH4sXlT4yFhrwy+ZmfyCheYO3k/+r
cAxF5TRYFhAHsvfGTFx/NZ1tRkJ7O2P47tk9jXi0o4aPOlUVpVMLFRuRkfGI
M5/M040QIE0qVPxrBJhBawZfd8Gdb/eecWUL43ETCvqPDLFirmG37WAT3zJ2
tWZ0UU+2uXEbv/GBOK6xQCqj7Eb91mjs8eh5Q3ed7bgoFJLwrrO1MQoLV0wQ
osXr3D+2g95ZSWMTXmj8zFD2kI7px8U8ziXkb/RJM3vvmkKHTOwrs5t/uMVL
grJEGQWHpcHBeqilToN+6vTeHLAhRP94G9NP1u2eylyA9P9Zs8ff+UTpko9Q
3XPPZLHLqvtv99t3fm9U1mfl+7P6PsEHSUFWxvYEIphk+aPUOki8VUKz5NgP
cdXyyWpCzDteaxwf/zMZC/cNfotxFWTTNmqMWtrREML4/pLGIBX0u4GLbcbn
mPVG5/Ne6bEYsuxPWR/ejcJKCRbqh0DyoPgcjUmdEhPUGgQ+oa2yTqlNR2iN
jWFM7nJslu+7uSy2dPhIsrbiTr969F/8aBAskLLvauMENHqsHbGgoA+3Opzc
WGAeg7x+/njS+DFTedFEd5jVZIaDDPMbNFRC0aqKyiPcfanIQLWKJbcJUGLl
BUZddRUioI3QiYh+Je5vkeBWDM6KUS353twKGrNWMNvbAU6QCK8lL11Wcan6
Q+t6sKVkmQcPGfl8MR+oi/OnJBW2Sz7+RMmsLt2spuoW8hT9pP9iYlvOpgBl
PW7LRcmzq/dkzgFsnkJm84xNmbfUgE6lzSwox4JibDGF13n840LhgEYAUjzv
kLkgxb+/Fi/tS1x7eRJThzsImZrAlICzPnbAABteE0EmXfcGamv37MmcxoIV
vN0ql4lViKshx1jbZx8uUG7COQCEYlm92rBH3ajApVPnql0uNvhdciM36Yhs
RtbCKwVuOWSlpHu0uhZGv7xHwxlI7/4rUI89AFSzPT+Bmj475XUsKXecfWg3
vhIhKQPMH2q0hYBcJgg5JUM9+mY0+RDOOYesbXqT8aalw3xxpv6NCstGsmVQ
26PWhgrGnb5d3HmA91XGHDKEfzWgUn/3Yk8Ec80u0uW07nOP3RMSkfia9Iv5
5UgD/PU2gstNoeWN9IDxGZ/bYzpiQiLi/zYa0sCjybt94RSizDAiPbgjpuO/
2mBkn5FM0yxQydS/LHSGA17OgjtkdmFXcae4jmwp9nRpVbARb+OYXSf96jtI
Q767zA7L49uK7oYjHpu/OuoNDM+8DDSA+84qBVjqIOCqy69sr6ylwYiov2Jo
Uil7/qHzpdPqTK7K1MJxXf/OTn+QTUkaY5RIl5jo4MSI5HR5KxA80qs6XJmV
KV/4K5FtFS68Fbn85h1FSruYAJhhaZmaB3V2EH74woWKuuPa0rYJY11MfiGF
JmC24Vh+o4t/GGssKfVlSkyTxKI3oChcicMTs9Uv8iRfNW/dI+e1uCmhf21K
s4ba6BUVg6OlmzMGlaUBbqFJcNgkBLgidV6rMBRkmyx/CW3UfmniXa+SbR2K
e487350Fx+vryT1UisrD1ENMsK0QL3mWB/NpJDNm0xRJq1U+TaLaHnEkfK0r
bVHr0FGsqg6UWxrdxLujUvgsT/2/W7P2tGLcifDxm1zGuMGOqXbVq5D3cYqB
DMoFeSzWhSknwo642xIrevfcqB2ptDlncfk8etWyRrGJXY2HkNl1iEyDX9Lt
zIg7EVRcgB2LgAlQSMGN6cPc3xVBDpW+qSkpFQ/XQJ75YgNS7oXaVCnedMmr
doNE5kw6M56F6FlTbN2kFLUz+goH30jm0GIGyo5TMybyUJ80QdfAS9PkAfdV
/ALmpMYcoDatLcxnRmEK8wjDARZP8i9VecaijFCaagHqSBqzGPRdltD2mA6M
uMzxD5bNkAXRpSreaYtP1mvWt3USN7VRbSW9hdfUD2LaYYvMrA41B6YHivkF
9ctCwZDUdPVMvnBCZRg1cFSaenSm8PBZ58yfvoCuUDYOSyoYzL1tYFh2kOIZ
QNGocHYdBa+AnbMaWuUdD/FDMdji5hAG3KXz8cK9fZmcSroR0UbryNvDX04+
YNdrQe4g0MHhJ7TuDUQtFTHV2/yhFikpJDYsH2lMtxirCd/yWvjww6rwqjxw
3KSpjmpNv47C+n80S3Mal1jhkxUZc/mSvK+j9VEdETcFoWA2B96egUBeSfFa
D2WieTasJGwXXXynTyaIDvZBMWtUjGaolnTf/97UR5VOTZdcHJqr+uhnPLuq
/VqhC/4c+88gIDpPwWl3VBIxk1zC5RafPX1a7liYkPVnVfiOwj+J7HXgJyU1
lOTV6h2oicTShKhrACRwdgaQwldRRhXHjE8zc0wnIJXlx2m1efSN7wo5GMXU
IFmbKv4V23+DhXjIfrN4x+V0pMbA8pWT6L4vjdqOY18A4CPr8LnhVIoYhpcp
jQVSyE1AwiC2BVwoql+1INqApasayr8je1S2V33suMuPFRA51HXLUbzFDVsG
FHi9GGfbAraaZbb5hqa1WAvUc/TOGEa8Heyo6zJxJjcUV1ZQgkaxRi8o12SP
xIT/9fIYynr3LylkwX9ZPc+98xjkt9YeyMVXyQyBBrermP9RNmR+fe17dJgx
uhFBrVNJdUcy5r2qYPDL3e0TR+qq0i3swR15R/dR+Rmf8ft3N/gJwx87ocNv
hWiFBlPoU/vOdOeDQjRaMlT/Y5X5/HuMonLYSeZRiZKb8aHq7DOA4+rzMB1I
mMnMCOOR5JcSgiMV6HfFUJs7G80J8zUy+jq+n6p9uNfrT375ks0NSPdyf/w7
QziNeUm2F3j3PbyffbeIAxXs25nJxNxLJiqgUbs6qnXmrq0K94YzmXsN15lC
Y1YKBsN++xWmC29LyBsOPcszgFGPWIHM2W2VcNa7GLIR/HUaTDsL1vp/GeYo
WJ1k8OhbUHmmbrz0gemBn1SBSS4RtuyjJIIj8AYYkhUOqy/+gvhibPVO2mmI
zu48J0IiZjGUgAePqa6qwOIJb15dUHX0837YhiPUpH8Yl4WTNzDT1BN3AswD
4X8q1BXMmzn1L4XZKT7liUEtreqbdqYV6UF8o0NFxWXiSQEL+UgEKnw+vFk0
EemIDc181+AygALQaArmd+ZiUlXwgjzOmJYUZbMSICXd/4c27/0WsdKF7PDd
OzWvoEx4bXvc7LVynLfKm75S7Mm+dToAdMsoymOw8HJs3g2VASdHBKQaQGBI
JAcrv/5Pt+z2XcSTpsNpg63YWisSkuAyRO0WHmevhTr01Ms0W0WhO+Cs4o/B
W5M4Le43GDTd6ihGwazSeNO4RydI+dzmoJByvIAzAyZY3FI5HKmFJcD9z9nL
FGYMtqYn8P7pF7I+chWmB0Ne6/9exAA5YRpipAXgdbmaMKE8CGttgy0RGuJy
SCJoad+ysk4KIaznDljDNorPeyleptJZWfZ5TYfTa85D8QO2ELbQU3wagyE5
i9vqXf+EC1WwGJln/daAiv3TKyAtXHtITjPkuC25GNCDgY5yzfHqan7NqdR4
6IfdFOLVKvYVFsW79WIrYCCCcS6aMmGlIcKnMomwmk4KQJZfHWdh4KVMFYWQ
9J6eoxjsDPYuxOiK8BrWjWxbMJvSmEJUTGQCd68uiOvo3i6BhZmwto1I27FB
ti6o1Rc9FDhIQDKa74uwh3ntSm+s8nfsP37HT56CkiaVk36YT7du+c4XYktD
n+rPvrt6QchXn6e9Q7MlFXa+4R/bpa8t6smBBoprSpXBuLWldd7zyKo5OGHs
SjnrtkESo5XWpuPp2ryiTnHhOeBrj3ulx/jf980cZnqwnxqthe+TkAAqvGxe
vLfqtUQy1lpnGnnuhAZEUMqcg5kuzogJtoZiE5Y9bFGE821UMaXvU3RtMN+A
thb0lMoAAZbq1CasApKQialWMUFcebDNTCyeGxc2f9s3naw/p0ivUe0sUG8T
FaBZix6UGKhCEW92xT48hS6HBDB3qY0cdAiDnri5E/bF0dpKgjISQcaQblj5
Ec4lD921btQwZIhNUTrhRT4QgTFRVY6+hE5256/5xXMuVb1M+/AbFhm21Yzs
Zl6bl8NIbOGVtvCHrG94NFcUl0ix8qbokilpkAvmrjjbXX5h99j5HEO8JyCf
ckoi+ELQRX8axAx6CwbT0wayLiQnR2UOL+cGL80YMF+Qkrx2Eq+vT2UbQ/V5
EIqPo6dciBek7/cChjXUe5xCyD0m+eGx1KTdVQWKOryRhjiQvM1mLyYdxbZp
O69Jp8e4ljqsOsfpfcNd/draGZl/ar3MKjFA3DDI6iDOiICjEQ0dDds7tVkR
hGN1g2TTmvRoPY6k3Ogp6EyuEImxRXVoEN2f96PQ9I2cwt5Tw+lUJM7UtTGd
FRHkB4pAzsQWU0Y6MXqxawSrwLX45d50Srqk8pGtc5JJYRjW+vCSalhnJCvI
KHRTi0cS8J/a4YbuNPJy0UFQA4IXxY7vMTovKTXc63UfIbA1FrvVek7PccK2
1htMiu6hWUknWFlNMe8t1JF1CGocjYASkWiRN6YF1mXSF92MFCjLZLfnPEdT
p+7KHfFgDKyKgyZNMhoT0T6MtvfeCDDU5Cr8JAbvUrjErFhnkA3nVY/KDMX7
pLOfUwRYc4vPGCgs0mTVT3/LawMPALJiqB7VQmTN/6VglNF0347LbPfYD5Le
1ajJQhMy1WX+j/yo2MFUfVtW9EyPG1ipNgfyCY7ANwFPKxdGkCq+dDeroIIG
NbLB5PPlyVhay3btRa5LI5/81QwpvkaH9RgRKJthwEgADa5N2/Nw27B0lXgl
COqeDmBpwzBeSwxvi4bUyrVoekX40q+8Konc2HHHuQ/HCiprG8/wW0JP2MrS
rgWLxg9IeKUwmFTFpQaxAt16ss8AxJcvevmAokcaBeri1u7is5TbHQ2FjmHC
m648lY4VNwj9K5bvZpMfztRUknJy+0eT2ZOUZ8E+px6IW+EOxsCj9y+ZSr4W
y6Yb1lEsQ3sY0qmwZ3YHoS1A2Roi1Quf5q88L0jLngxTm11Iije+cEzTxlhk
OXD0yPeWm9MVQDJjvnBdF6GyW/YSsxEos4Qgaj9HMncVsA45HL8NEEZaUbLL
QAjT2IBtPmh+negwFC/96dm2bzG5rxxxrKKPwCtaYiTxhK4Dv+J9pW2r+7Wn
ISXsCUodNG60MEqgmDKQmi9HQNJXbgQ3oJov5uOCbjcyaKlOZuaXv7aSCYRo
Stq6dYj6ZU2doSniQkGP0YI28ovfQBlEP5T+ZG3wyZSWPwXC/Q2Er1f66AZF
zVUNoYXd8+dOMoDgs8O5egszHh51SLgpCSVzMKyvl1JGt/qseiSlcLjgDS1X
jnlc2FZ3TnH0UqUsXDnxwUTWycBVR3Wv4F8gwyEsB8JTlra4naqDETgWGqxu
YKHTP+WoiBSYMNyKJmiKzCzTqvggDkofhLMnMxcNAoqclHm5oTA4EFfYiFRK
KApCDd6ad/dZS081BiNKgSrmYc65wgKsxMsfbbNZ1DQbQ6cWkIkguZWm1LEe
Ye+7118Yi0tHt+ZmMsfOK2rpCapE9b/HpuBidZN29erbF4vDNAeLgyj16fMZ
nHZPpJjWv1Cj8daNNSzF3bLEIDBn5DfVRAkvoWBi6pZl5aPZ+Rwgx8tgSA3U
fP23GJI5KE6M24fquGL8ltFEhRTyW8+5xUlw9uA1JN59/j9OM4qjA5V5EOke
xgxGduwHFXfE3NbXGxG3QeyZSi4YcqowBqC8R0EFURoe6hRuZOsNru3VEJVD
2nH65rcQWq+rxdDKOSas+SpBKzyhubCfyyhP0bN7C8MPErSf/5tEydb2aCjp
6RpkgQ/+dzCDlEElBLJw/ufcgA4nkAvyxolvELG+diJJqJIyMHlCQfLyA2VM
9HUXEZyUfdRMRiTj4Y+OR2R+0mvwkpsKl+zIU0nD2CLiVwwzBzUliinsETrg
uNGN49rz3mLsgSU3pxBRRju1AMJGTnQufVkdjXiNhIc9lDXInpKwnrXO8pnb
t0obHYdsQC0wrKQsAZN/UuJeFpHcAg1vMMgxkQ8W1RDr2WP1gnV1rKpSwMjt
cCKHKGKsXL3Hh3TVKUF0aW7YNJqrw5eS4OVcaXolu39EZgQqTEkoIJXIAdQc
a+zDuD/sE2DQhn4oiIz7lqr/wRyEsxTNvNxVLpQwK6bqkHlI8pT5U/sMBWCH
hyXhqKlUzHXzzUA1kJvG9V8Nyfe5yGpWnPOhXXk2JW8dsOBUG0ZKfFyGHHj/
kvAFzMKB0RTmisV2urlcYfDbJSgIqJVxtFcp9K4l4ZDKPyedGr3jAKRd3Wor
2iyKOYdHI10qehD1ZPcm3lekKZQ8LVqin7dprFhhBNv8WV8i9tiUJnSL+6Jz
4dHyECHKjDVUB5oKw8/04lr6myih00veDpQf0lKq/oJG+PodPrc9Mo558WcC
hZwo6L2BASYmO09xM97Z4shbO3ahxAWg9Dy/bNM1QTIURFg9PNAUe0N57BQT
zeNdbXP3/zwyLnHZ8poR6O7LShuWT+fTjzn32hOV70TH2/A8NjsLMMUmPF0n
35bhBAVpXsHSixNaIveRxU8OJTkhFmBZCqqAY9mED/NWco8+NIRjl55gXCGh
e6Lmbut20K5+PMI3nYsr/7j8eLP/FUnBW7XxW5FDN3oYeEiuSLR90/TPeWfA
AHIW5JHRHf5AcmeKpOv8G8wTsNAiAREFaBLi8cP2fLotA62hWiXgeIaU3kzv
9JPMBNkNpCGK2tFD1D7ib3q0NzuCv0v//QB0eFEgvwaNN8FZnmtlIhZgXqyC
yjChbnP5knMbILoU941pQfO5842D2GEOYyYBZTniodvFW14t/JCEdEznaZGt
Na1xBbEE1GUnpdWzFsG7JzaKOYAHT/gPUcFzh+qwpWhgadhnwyF8hkLbmgTh
g7QuLZHUTEOgmWSZACC6NkUSmB+ORJiI3OoQZt269LOsHnMUr34DeqCcO+8S
f124ZqVA43/MddUTkrGUgFLC3sDO/LlZSKU0NqoiFr/CqdPFD5xheSFciWez
+2luh/oCC3GQfYfyfjs4ENoBmFq4tFwNsuoDPl7H/7xJewZQusx1o/6L0Zkd
XdUed1bFUtrQe2r6lx5kdnUqmx8vnaVlBYu5WtGn7Nj1O2iKBbI5bx582FMt
P86N1AqU/zSk+UJu3mxG7CS7hhc374nrZNVOC0svp1cI9qNOkSCwwiLP4/pX
3DSf0ChWwEoGH535L8c0I56UnMzGxdhrNV6639T//V/XA34e+G4V0Raa50eO
Vov/pWSMAG4Fr4FWtbKQU3/0QCEvvRgpikwMAyXzzyJaj1M2rn+gN9YyH6N8
vVtWSvtQOe6QLboU8GIqyxe6y13jYJ1sw8ei7FYQaHqSpoZ6/Ki0d4WL+sFt
94BIM/kWU9rPaf1sXXVhfgYIrnMs7wUrP+8jB0EriqIVXgX76qfzMwM/uz6/
e5DKqJ58X67uyjZpIEsScX3L44OZwCRE/Bh1ic9TcfNBR2spFwaiD7AjshZH
nWmFPYHe0qg7P347iFnqU1gtL6Xp3ihkUIllHPy1GnLICUAPX+zXYCPS4j0T
wH/DHkT+gKJhX4t79Mom9dhhlfr6f1QOqwimBCs4AfaQXtkfQBAO1z6kk9d2
yD25Mv9J0BVdMXRzPT2UWKLtjAadgJpWQ9WMvP4eT8OPp4sDRJXwNKOSA+pT
zzdMwNcqISq9YEUEoroV5hXfe2P7TxyFDsbTvXfUj5vnILrSwTAy8L0sXA+l
jh/h6Jk9jhV/6JhI5IKA25fb/zS+At+zF2SdF+eWNgybZDQXdds5EQwq1TfN
bPIPdtlFV+ceTsb9IZFXsxCyteu8Vxc5y/MRSmAkjCjh8PdSroUWt+erfkkU
/cBTtjfwwYjKKviUAUpT3a/1yU8r/nAgzxJoUL3tF/Lo+iywR2+LDplAaw2+
+FlFr5hdo7jRHYFPd3M65JmAJe6Vd97il5YXiSN0epLcjhb+qQMr9ICW1TQS
f2WAaRIQ3mEaa60oysteu1EV8nJ/suSR6S+ltadN4guoi0meKEaTChLRjWuf
QzUhgy8URfxxTIY/bNcbAgZsP1ADP2TXv6Z6s5zJWgjiFWy/6zfQVlYoFne4
CXy7rLxf/ZLJrG3s3wRpjDKve0bTmNkRco1Br7AHyxDvB1n5Z5zSLkp+hBo/
qNkcqRV5loHr0IIqLnEwuSgFFKD+J3ybHiiu6ZqoD3zq+UNQeYK9yvsQX2ay
UY+frER88EG7fLpdlAVcjkS9/FU9OLmxdUiX295eSeHRNq8fM5Za9KfqyzjT
PrC+xjP9yO+NGxFWWPicmeHeru4Huh2Qg/S4iBtCUwB8JdNZku1b/ivB2B/X
/9ELzmZt7m7M//HZlXaAb/uxRpEBmmkudv6adWPOqP/XA5LtfDf9KJctu0ss
j5UqEpqhqISDhzhBXzEwqMlzDC0ORbLqxr4CjnVaYiMyrYosf41zvToJkReN
YdI7gEppGBUbCvl0k/0YqEpeOaXcie3EB2iZPOJA7morMiF9lTLl6kvBuPLK
HgXXp/+tUlj2dBqDASiw2V5FCB44pGsVXPmcm/ZCxoNLxPqjhtOs4tIWpNTg
5sSG4z25MrcTd1BssUcnuZFQk6lC6TpZm+lJbj1y+/w8e+gv9vleqY7LAEo7
Q9xjaxq8ymaRcEuNZ1C3Bpm7X+yvbSKmOOssUMpbU/kmY5nOKL/ItqtDER8D
eKVVvXz+EiBqHlUdZpvxOnaiA2g7N7wqDu7Hl2hgkEEiFz7twyyJLUE8Q8/N
ci1YBHZ41QEsOJQBJmGBA0h150jsro8fasJdpcI3ggedtf6K01p+6V09K07C
fjq58/ZxGy+DpcXtGwxjv1QRLYdlDFNpFxpvQID8pGkBBER/EpZ/yd2MiGfe
2OoNdI1etKR9XbFvChd/IbcrzrI4RR00tfGJTjUh5rqQkQMl+BvpHplt59oR
hlGehiyPQRXz1VfrNzy/nViVmGAVavfLp0sh5hjzYPAoGdpN0jb+ajUh9X8x
2eXa2/8wQMQUnEj5zY/8NdSw2fdqr3yoaTj9lWy+xuWJ72xBhWnj+X6CUMKM
wcEcOq3njcNUijVbVCSsbudBgjYl1nj6pQooJUi9Yzl+Yi+HqOappePNBlvU
JOVOGCRUmPL5uxlunpr/B+XDdRR2CX+Ii6/ccTYguQDfjKA0lgVkIsGxdft/
+OmOJa/hWpB70fWN+XJcuOY3hdm5fvu546WkU0yrELYQqMFUXmLw+dguMZOU
5UKGWbuKGggE+Of66Gas06Batmf7HPcW5mLgFzD1pqFM9o8l1YBXv6guuObg
vfu9TN9U4hxPM3RuytVLL2aiCE3Mkz5yuASBK7pRnyL4pdSrOQAhoVCOHnsZ
bJ5OTcYpnGCPYlZji0CKDqSqo7tLQCsIiOonqcfNciBZPO8gyimLECK55gbN
ao12S4Gh84ngrA0HYbtdXRjrMhz0QVk6WraaoWzbgayQ4jv583I0nQhOb9pM
8+45Ukqr/7BnhIRqxgYh64FtywXZEU3vIrrABwD8jIgUuBtywqNeT8+6ZqZM
QcNfPIgeae7S7BrP9VvmEyW+93qz0qWrV9Qmy6RqQfpSQc5XBsJ7nugmjmRl
2oUWpVFjlm/hFnMUXz/uVFEpRrW42GGHqBhupcL3KYNNHXVoBeVr0ECCXFKp
IPNRHZZj9eabPqSl9dA7dBNUwbfcmjcgG5vxpV4Hm2bBxDEDDkefNAvb3nr6
RlhLYhl6+SayT423ZHyCMULwf7KAJwxv6CSdgnyZETyQtr5wIrL64hySThLd
6xPy2+tgGyyI+7NKVdOodW7RY9WtxwRbNHmDwsv2s4+Ary4JQqBTG0kxLb4Q
oMXMI+O4c6iirRqQ2YAFDQix0AHQ9m73MuD050s45HgQmMm0RevJAWYOFRno
xTIjnpr35ESxqokv1+Z/PV8QhkV8AI9Q/UYVLKSRNF7LPglaxUMkYz4puQor
4iuYg2SZPXSLqgTPmsFbhapZyGjuB7IHCbQsxl+vQRTVZqWfczfXvVlVoSib
G3qP01Edanvu/gr4GuLVW4gIOqXU+80F0EitIN6Z0brSpCYsOeMbr1YUnjUM
SCeTPBUQh1+B3hvOufUO+VTNA/YH3BMkPiEfmDrc8nAql5GHOhrpy7YjuPS8
FuGeKdIHwMyP9VG/EUyCtsAooQNmQggqX7uFcFe3p8XoZlMn1iTzLDtUHLuu
d2JyxeVqscdLkWqimGqNtTx1H/LnDntv5nEx7DQ7e1Q3cvNlaUVI0/Lbbi+m
Gc+H1y50A5taAq4X5W2l3INNEWxDAv6u/X6XpYqHzuTwbOfvjZcikd9ao1Bf
7rfL4kQKxx15my2Lmwzh1jSIhIvj5n2ZJJFqPYJIf489N32hFsUx9mXBbRak
cCIK2/T5fEeNgzXxRGXvKZz0SkbAmX6n2o6SSpHxkONoOPkj6GsGnB2UwnPS
dyOx+OsR9Mxbpx0wDFocAEDLMXqOXAPMM2R2P9lci/AZrluNDTgSybQ6ENMy
zHiI23UhxZ7DTjm/P0UmnLLZzWfiD7/74PxLUDoh8bV0tiiZ7zI9j/+mCPBL
KIh4BbIXSiYn8pq6tsA9optJDUD6ELG15b6k2knSKxqP13XNrpe3f7ceDYC0
KPG3y05K7UHhv2nDjAEdo3qAfwJCo6MSrfXbfQptl7JMM2yMZ7FNpKHJn7PL
184d1HJsYK646Sm2dDjbrxGU7bFOm2uD3NZgl2uUPvbjJ4WCGeoTxPm8JQvg
KtLr91z3ElIlUcLJeIG/x5+j1ZMYKZ1KbQNNOzx/Mhfh3o+OCM/8oE1MGHc7
wooTLICAZpKe/3hXWBuqhCtmBPII7o0hlXRxpOgTNdiR59Ni6W9xUQV+/sd5
TwmEjTLd91Hmg1gGnN+sMnnddmEpnWr+agfzOAvMHh1dbXpWnQY6j4HAPpw0
L1ftCmXy/CKO5Z1OCy0JgNv4ThkiRV/1XBZ7CCynaFJE5cLGirZvTqvBwB3E
1MoLuP+6q0KNcJRpqqjMxXgk2ICFrlPLDza8eHOA3hVpGVAj17g3ICKnmFeA
vEexT4dYGfsLHHuQ/JtWa5jPrNi1e1DnxKsMOzZPl6j4mcYc6RZYYfi8DyVn
raTXtMm6dIHsMCgXIMBapAYBUdN/VaJQ4B7OQgLleP7aPSIFxicUFHi+g7KI
pcorVLA09o/AeQ7l8M4CfjzTO8y1oKJouj+HkQXIWGs5WTJsbFCmRtOtGZI6
5PaQfR6c9eyi767y9IPYetL3SN5Jqdtyd9gheTuuQNkLiw2oxR22utKtC7D5
t85UgY1+ZyIMt4C5Pr0BOAtrgwxtDKRLYhJ5tSUnUYSm2PDD+AILRaFhizv3
B5OKe9OKWq8/Ip+a3VLBSlBKdBpCVg1nmWfR2BU3ypU3kCCnt3KZj0prCAA9
qvm553h/DxUHyDIFb3jS/TqlV0nBtdfd7h7txbdBY9nuQAiS+GL9eFQZ8JNY
Rri3MuJPJqW1dU6SBg3XC+90/zaoiKAlIpthoMlXK+JqFEa+LbXAc7vIrla8
LkeFLj3Q0EdYs8OKiC19zoLqEFaV3RZ9lH58FpUEctGyaIu40ogJRB47LUPR
cSRM/EbIuI1BiC92OQ9RkJlvRsW6HWWpx35OM+LQitRZQ4q2DnNMpYypQFnO
T+hzks1kRcTDhganAN35gm0suGOZOlSCaqxVpiw+4aOKjk/XHx6evgjfuu+X
V8JQJWjVw0WDR5dL+uoMkfoUgkoY60I2hqmqGuBOoM+/JyB2rCfXRfhdXhCS
9C3mZSdpFG/Hbi1K5rBSEU6zce4+Ea8vvvIeW9Vz1RHXGV52aNFNtefhrpyw
FR6l5P4KLl7QQKmlZrwdaZgexr9XmF7c/NlnFINVP2f0kFA65R6Yo/p9PqNf
3ZFKiyrDwjlBpmjvNkM29cfmhxcJ8ndKlmWK84EVf1hv9VEXXMplXAOqGJOe
BbThOYfi/1aT9EACL3fdnemTe4d80JBHv7vCBJGbT8jciPni0RBYKvskaeUI
ptfeRopjfdd7AEiCGSAU7oZduww660hOHE9R4e0eWwy96SCOWuA5xl/rr/eG
qWqq4r9WtaMjxi9kTrhiNktROLue19apeogStenBHdXgNyviDv0Kj0sKS4/A
toX8SEtN2b5zNriGvF0eUw40zb4qbe90Wr7Aq9sia/ssw3q/Z1JuHI3u9MXO
hgs54FNzTYWe+3PhMTs+mC8SouC26clUWje4O/xevyNz21eATev4MA1f+AeK
ZRYvFmu1uCMRdo4R4Wq2R9GqDVBK0O3Wjbs3zB/a9aNx7JGbirIKcIiu2jSx
JDyvJYzZvHU6Ki0HggZkJ58nrSlfmD6sdeOGgIVXP9wf3N0rKKYHxIl23s4Y
20/Cv31V/4vXN/4dGuqOCxAof+h56o7GOirImMKBaxCJ3sgxgeFTAV2TRSKq
bmH9RWmaRXA7tUgAKvzdZt3C+RHe+bgsc+qGiLMumZBf+h0E0OE/bsdiurtR
jOWSajAWrWtPvFXvgePIuotQekvKmLnzEjcdAG4exEeWb0EF5JaRREcUcmof
0Z4/1y2jr5wF9bAW6c+qK68SmiHOltD6M9sjxnSSq8l4xu+bfcra98fJVfde
Wal2k+c1Gn6MUsOyWtWgMdyAhnqui1PlkjX6FHyesyDTTbcm7Gpg9SkKQVVf
80S/gAt7IpDcE1U7DJnhw+WjK3yqXbAa87fHV9MpHq6EhRzieTnKh/oKC1m0
InajeQt1+kl6fQ1s9H+5W5POZ+iUHrzBBkmBkd9DVppj+n0R6orTLmti9i7p
g/W6Ui0UcYTqvB+9SxN0D45cxocNzcDe+yKmWcwOjSUUN2jOGdXBfimFEPE9
gRjyRNeQXYi1Ti8BYJpkpIc2WVj33DFdw5iyUdkV/cIS/3Psx7v5jYshwrG2
3PIO1E1yAw7GMSa13MsfNYsfxmQN4aGv5m2R68COs6liM+FAieCAcCrYySRM
tRuqHck3PMEOOErlV72XDsiJKCGAvwaO0xUeLhJMWrYF/QvUcgw5ZffecRis
9SFI5YcnhAZnVyXO3taMUWbWsxixU4AFktPUEZgg8SHWrWOkUzeRtNClRFv8
2BQmI5EC7DaBW3kubSQoHQMZ06up279/UQ4qoeFeMeEaexo2wPnlCPVnRLGh
Wy8uSYN7tFLZ+RYqGWC9fPoT2q5HcWRVFeEJ2w911NvnNBvUOAEfoQRm0mEA
Mp4IeukzX2W64hUuQlgVu9g8di3Ob8SP8+2Fs/nrY140Gr7mvuvDGeojAHcV
6kns/apAOntM9MzumKWr5VKDv9yl/shPMMcM/eEMBy8sieIkovQMjdRjv6l+
kG427c3oTEoRy1rwIiDBAiBgNs4+5kaYRQmIyoGiVdmYMIdlLL/1FkAjd4U1
2VCaO0qEKYwvKZ5mx79kEWu8rAD+rs2AGzGk3WQmtOCG+ljauzu5VRycTnry
Q2che7kkA+no6A4O9ts4mbdVPqr2xxp+LrJ+pg7j1KmJSsNlj6J7cUayTMr9
8MAH6q8HfkAO4q7efJCqd9I6TR7xouD8c2F3BH5Ereb42hGMzKOubnjlfJyM
eR72ac2xvcMQg+GtTfK6mX5FcZdu1zK7TnbIJ898TxgpDgv42KmZyb1s+Q29
7mEpDeW+LQ1PhaDGUOq2np+TL6zNIpTlsHlEUh2hPthurKl4eCquTTxn18Lo
pHQ+XcqK1eL880sJ8a/JqVEZHjTC1oLnvmtOAl1JcFpXS6zhLoi/ft/6lWPY
5JFPhbc/pV5+BBfH0Ooktn7yDfcgn2oBReeOblDY9CmRthFXf22jTMZWBYhJ
tq+PDcMG+xQARju2VwerSamisYP9AdlliQF22ELVSfB30XKekvyuZNmCyW54
ixDCgJtLOgb3wobsuCpVgj9YseeaoFcsk1EuxdTb4pGVK1oRT0wwHcgTCH8m
7BZy4jmmNrphCLoLUrSEXOBHKOjKS7wiFO/YQ0eaaJig3FfyKw2aCrcoWfvS
Sy4rzKGyfJYOn3l+B9UyteLHXEEN5bDaq2mThxBembC0PvSdu7zAEA7NWVtY
JRwXawPbJxO4oftdw5YQZrPHtYwsNZD0OuAT6iUXrglrPbeDqZSHp+MXS4qr
HR/UFXV+vNZ/ANOKujilugygXSUvRcMY6TEG6FExRgKXET6bQSVm1bn4ozAu
fMwmtGes2frFt1X2hfympfPZSI9CXPY0DJIh29zZzNZ3cH7c/w93R/0QS2xU
wM6s0Ro4kaCTFAu1DW7A+MABhr3ZhaYWZ96yVbMI9bzXdeeCycFnV1yGfwHs
EwDnpNnfORs9D8KzlKdTVucb1Ru4G6BPOK0UC0ToBiSuoWrc6bDPzpUaR5P4
cMnS8VT8JA3qrh1ShipyscIoapFaXTUIdlvCHGnQzJoZMQPFUiKmu4xaha2m
97iLE+9A+qRBjE1oD8xrzCe64XfA+T/ZFvIFHcOGGE65TaFgq5X9KP0RHs5j
h1AyRD/gtEToE75RsLotSh/j3fksbh3O+/4zBVxu+TniPYaOhNrA5iX2NtAn
9RA6wtrylXxDLZTAIpGvOkkn8zi5vaRIAlQXyhKfElhbb/BQkut/7jqTnfo9
0LQSndBNBqzFrYRzgdl3XnKRj6VUPi4ojTRUK+3o6BJa3wjT3jCfZfgtwRLI
LsgZ6WBPuI5mt58re1AsBds9Olgj23OOQfOVLAsayAXYV90pkfVOxrfFNMQc
4d83jZIsrntRee0Pej/qBTpRBgP7lxgamzfBoCiVn5NkHupJlTY5+VAWWOPj
x0nsMLhc05lBhJ7GIBWvLftIt4E6zjGoDD3NIEA16ZW56Uu21dH+LgaP3DkZ
wJxMDQ6bVI7vLAJeFkmMfpBPWBXTQLylR+2SoQTMpdY5cmX1uHpIxQt8XfDo
m8JVzVeGiW2+nC7TVJTeAhZ4mqzX+8rtpUbQ+dxOyixienmxIX3z/6knBaVp
Ol9jYys9q+BLw6Qolsk8FdLJFcOxPfOA36V4LQLuYU/jKNCpsyRyIoF+mkdP
Ndt2zhyu8lmZNZVNqc+pVDx3J2vHkwZV+OUoI+qFZhpi/r3MyGOJzCZZG/4I
21pt7LuBAJEAhY6/GaefFDbZ8k+xcAFicLpY82ApjQwtXTurMSHuK+NxSi5L
gS+KF1tvezRjaP6OhFpTiuwMV0jqvHCgzT29JKEDtxHTmT7ld8Jpqu8iRADE
ttqQYPqTzC9TrgmcAQW6TtesIfUEMadlvu3E35uU9NAwEEvsqTCbLlX50hII
w/d1p+Tlz4X+T8uqL0kiBD7wl+kKzzUXhKXZ13H8VnQBBSFjy+7DEFMtKGBE
Ir6RKxN2aBjDqaNquOubKFqziFgXvFeFsCd6hg/sCADoFHDVtIJ0fAXQdh9M
6Uuu9OVsxLlscVGikqI3fFTviIXgcZf4b3DkvHaH5hyEGkkchTjl1/K7WKjT
FwefRql/uD5Z/pvZ733WzrVEfUvWJMxUziwJvAAbC1hMl1e0tqm8K73XtVWn
SBkl6eTzDlOqm1drhkFgeaVgPIBISd4izPC32XBjTL8nfBXJ+Q8YfyGo2LI8
7x9I5gNPBshqY2yQeMFXxXSablVz5crTg5eEmCxmbh+eV3t9M+ix2i/NmecH
iAM9AkNRaIOgikps0xCkB8wh9Wvqg2eETmZHYc1CTPUlSlcFkEj4qX7zyJeG
1K+zO6D+ucb2TtkGDgixGWHmSZmj3tfI8HzvdnDsCeWT2SVET7JakuP3lQLr
iaQIOlB8Dr0s3sT7tIzvvS+Scj2OB4fOYBf1SmJ3U12k+5+/aqTZDS4cNQ3X
4rVHm+B72gGCqELSQDf/t7LctVmtDGw6bjItUfQE4Dr0xtAN7aP0Lv9mcyKK
IHmYROlWO7RyDb2vd+QXuT1hCdSQrld6Yw0qgwaNoviUt9vuMOtlFw3T6PKj
ccXV7PzdHg0p2bz95NtfzWqHQMcJbd8WdMdw6ClfabvFhuO+tTKnpG9ZsyZ1
k+L7n2myfuieQp6j0AeWTi2xB80qgTe5S1WKfRHuuN5PNSQsc0YCXQ6kFAr5
Wh+178Ze9QdpoTxGuCIRvJGZmOm8Mim5u7HKs5j+wX3LR07vLsJXJmA82Xq7
g2cPkh+bjrwXAlFBwljQ54eyQu2vZXKefXShU419xsW/CJmu7LPcvQQxTH8e
Awxv6tX8NKoSI1LiNat869peQFjsVmTiB5yPhvAhjnFsGo9CIjO5sFX8X6Xc
p5o10baZzarqDufhHbhzAgKemM80Fg7aa3rBzJbdWo/KkiVULx/Yl+m288nH
vLgG38MhZ/w0/HcKOCNrTpSs5H4LxOyoPJJqGnFmi3rOAG314nEgm6EwDRU0
2nNxuwms2K7B3RvD2BOsfkPVIhtgoOLYjWePb5mj3QFFjcN+2TKhy2GUyPBr
ZpehyGrgeW8Xqz1k8HL6Od/N21D1yX0wNAZGbOENKWMK1kTxSFYWrxxP5Sgh
t8GU2s/cpDer1hBroFFrAhIie2XmBeyeoZoB9oWHo/PAh4+2BOHEUnCp3guH
1AfZgKrmGVgL32wx+lWyb4ZmMISOPHaPgGSkCAtO7L5FqwgahwW2n8XQZ2po
5W4F6fGddeZggJNndxO2rVG8znkUQDHQzgjWczvKpZWXJvSPzjBHdySVekjw
rYwtbkQksRs39Yr7LTPblOKfzjp21cYwgChylP2P85Cugu2C4+oY6FBvtBcB
Bq3nNITOlBSKQ4OqD0wu3OM7ZswB3YiV4RSs0H8TmcRmsY6XU2s+nTM+kryN
QXWKpfhsyVkAJU3BBfH1GTIRMNlQIGtkOrPppRDxsdpWDDtN2TzbaJwo13ec
m8AaTKrFMCGbJoQc9zbzcqTdZ3fcT2y/NB7LCUHdpUv8w1T5JenKPoj9zeMc
B/NDUDC2Dy2IXd6Ock7NwSt25hz4biR4cIoj4yrPGHLzTf0o4H5ZeAqiEWIO
7pnF+SIenUYaKsn9GoVpOEDv4rlXyYZa9Ou31vJf4dxu8JOWZtE2KPp866zn
YCAop8l3d8hTVtEwnT1ih55NFkUB70aJeZ8NsG7envN6g8toyW3EzXdJSmgn
46Sixbch7AIn7S06RP8SC/L/ZRWOBhhXld1JEkSHZS8tJZip4+zNxaOSEXXf
Am9f8OkL4s6PKsq/w2dtLhG25+4AtocBtyoJ66iq0bDt8WBf2A4DnMrH5xgV
HqwC+VwUcsd6xO5IOp1lPykxh+HNPspAzC3E4SZphcZtRp7W1BIbtSiYUsKX
Uk7m/ZHQEPmDIx7F+9nfrvMUEG5n4ZSquDOwtUXnM926VVExQQjzO5vTmOs8
eOT2jOSg762YXpiiBUez9Wwq3r25iTeacOEk5Pw2KbVIYQBfspD3vi8xd7NO
VEIArz2txu9tNUqII3JwNyVVIKGlRhV//uCCjji9aYwFr0fq7PVBqqaXDVLh
Q6q0/GmV+FL8+bN7nGwSxD1ExRtvv+2gt92XZKRusVXAJDDgcFgBOqMJMSGN
jRAmctkjZ9x3sZM4VjyqlmspOKqZjVD2nwrOCm+1FnApg64m548ssnBKbGZ6
FlpApCqiwf34u1s2JQGY9M7EQg+UajWNOzkabvEpgMHHZwNo7p0+Yu7G9BOD
8rCP19Jrvil1xE/BM0+qCYo0MCYSET5Msce7BiU0u09pXmgwRgOKZYKZaRCV
YP87RoIMxJzsshphV6lw7Q2bJ8CJrMu0UVAfP7EZU4bjbaain9hU49orCG5J
LeQgvOXWZ+lbzet0zU++bhxf4qJjTvXJF/5EVtv3YIx8Qc2Ts+EvdxFu2kNO
6O29JNxbip2bWosm8A3diyZzfHlvbgZD1/DZhnZ4n+x3W6nbWWnqPLU0iitf
kPgLEDoUKlyjwIcGkRZ7PIhOouZMowKDm9ff4jQVR4ssdGJOEqZIk/pMVj/3
SJM4aulUlhKmm46wkFETyyTBZ9Q2m6VUuFnFwTO0ufqDBZygnDPiwI6NQLDB
poaqWU10FFuytutFFgkC4Fcu0YuiaDty92EnPs409KX0N0ZTM8dgySZqWzpK
LwsS6q3YmSGMp4OiAumgzFFEADzIktAfwgdANMoShbxw6Nqjt2JGvmA2Y81+
luTinDFceVvbE960IzorYcZ8Os6xxJiypegDNIDeO1zBEcVqlD5AWN+16a04
4i5mr6XVhjJ1iG4s7Zlcjw6mRIQ9SFfwMcc3kytVytZnuRXwpJTof8YCkeTV
92HI374U6Cg842OLSHmthDfT4VXM51ZS5MIUS8ibNYi98N368JS2hBe4Rwps
3sP028iHWO8tiCZ/orD06QKxlp1gi/CiJ30kM17gUwuMq7UUqcJXiSypmpNz
xvVr7qZnwUMEaxWEP6GNpBOkxJ9ld6cJs8cV3KJK2fugBoioFyCbQTlndFxq
cxchjl1znG3HZBpNFnv1CbyVVUzDA03srlJcSt4HXyA9ZukSH8Bs23NogVMh
5ckmXgDVV0TKiVS1cG3kWux93HQA6FhwT6tuoshOfZSM6+MylcRmbOYY3W2l
G/8iGclI18kXkg8xXYuRE+XllqHIxkl4Mt/N6E7VKljWCrY9J4qjIuAj7Uhy
WaRKHP7mauBXSptg494Vps++KRwmjjVk59BkE/MLi6HrXDA9hY1VjgnyyV4V
xODzTJL4xge7Y6HpB/4KQT3ck1PtOWtnPWKVQFpMuuieli2z4zUJVwHDEWH0
MGh9/bS2TILBPRWLRJ/iqWrBXiQfyy1CvKIKW2mZKhXUYlqeOrE08Ih2xlKm
pRXT6QucYJ3o9biwvXR5ezpqlaTT54ucP7hDCQr1w6rSwEPKhWsaDPrzbkPI
kalC+mJux0EXDZFe+AWNZ97/cl2meP3UCmZuT9iWBdGWkOkzPZ8CitR/hoSw
xWHqS+A4eyngAx9SfRhPTHeexNSRTl1wjiRNVzjirB4nf8M4yKaiO+W+soFS
VFzsgPquhGWwJi5IwrlFZr9rEHklZZKDUMebSZ0wodr3/0r/ALT2XqBTyUkX
Ws+392Kpgjg+sWNQawdfisc1odosNW38N8ZZaTZIFx8eOOvPWYOYPWe9ue+9
dlWxJKdDHRfJmMR2AX/p6EWvMYCWMmqw4voXynx1KHcCKs0m/M81JFYl/Jtf
A6TVzeyCqnt4cwm0isxFh7/sS8DDRW4N4rsu2NbCPAgFPMmO+amGrDfox1xa
k65b9eMSpw+Jg/YK3SHAs3Z29sunccWJd07vzpw0/4gs3GUCbuxZacQX2GDf
ALNJI8545UUPW++uuk/77AP02XztJwNFz1+u5caIDG/4jzinqmCZLOVS4QjF
R4YxhqAjbqv0XmTW9Fli2Iqpi0psHjSGpHlMw/qvlxZPMYpK03fPYIL+TvDY
6bWuSMB9xoG81tgXZgouwU1OUIlJvpVLCyAcDUnsnCgQ68p3LFU0mjAXI717
Z6FTs/HVOYdVBMuAO9N8cskOgzrmJ2EgnE12qSDFFL2j7mDuaS1qw+eKAop5
bPC1N3BbSeefFtjnyqQfe9tajJWCP4lwJdzS7F/BE1D0xw1hy4iBGecm3u5A
KdkCyPfvya3K/D5uWvyJRo614JfcQ299tMiGMAK4ujz/0XDMKo1F536kBgWn
UeXEsUiZylk1v0kdtkAjnFbmpiXz+SkcmHb2vpdEoz/VspFm4B2H+i8CVMuG
yK8UsUcnyWlviaTD+/51OBx7JBCWwZVr/nrG/Jc3TxYLJR3Kkp5FbGUiBKAl
4Vu1di2lrc/QYdcg2FZ8WXHYiYhgT7etPYSNMNtYuueNQ8t9xZqF8TI0pAeH
j3SrT43Nb3yNiPTriQrT5tdC7SVHynocX6uLRSSSUzuxa8P0lm4mdiOe3ivw
mkeyxjAULyWSNOoqh70neIUm95iAzAnB68CGJbPsSbNgDh1fcepFCEL1m6yf
mW+2RHgVQ328cRVfSD3hDsJyRxBMQXwBtBfmS91wunCZmX689POQ45qthJUk
+ClZXH4X4zA4BK89wPdtDEDkthkKIZ9IdIdhzTWRpWvR9+P6w4mNsfQ4hCTn
dIRCVcqdDrBfO1Xth7SDbcMSbKE0rL+XpHR0fs8zf8k8cr3bQdrenZeXxCYD
gMwcP2te0TwpIbG1zr7wECYecLhj7NUiJkg8Hq6m3XUVSYKn7f+n3OW6kpSw
Sleiy3HKjnhox01Hj4Fgid3xcBA44vY3O93hY/b6T9cHZlp9KEL3lzT7yQUO
vsUAozvHU7hxcOuwm7rA65d+//hlzlw0AULnkTI1HUgbrBEYIX7RV1Cyr2Vh
V5p4VkdZeHa+j497BUGIxSLKD1/vwkmKHJflwKIpffeGUBMT7gLSN3dawqQh
mJ5H+s6MJzrudtWpmsdjRo/I2XE2OyJ0KgyaH6R5KdOhgExWmxgr+Wp8BKgT
G01OLCtTTcf2hNAv/81b4C3PWy1/LYGO4JyoQ7NMQjzYtn1BSX+4jh+JWH+N
hP+8VMEbiRZrJUcp/+dVinyGtCv/XpAPUEseFhAnFu4U8EBNaxAZiXthI/Fw
QK44hQ8UPHo0115kiLYnveiZLPxp2CFdnBKzOB52ajFOhgmiYTEtGBmsL+AC
qcllQSMYVUWI6AruA3I7uIzjOpn19BFGK91TYyLlMWj5YDylxZu1+EUVNAWI
1qUv8BKF+9qhKlyonACv+saOQV5CaBfHbB4ZKbqN3yjZo0N50byaq9bd4ir9
/Te7bSIempl7skD8LR/qpFJI+7YTU71D2VYtSbgsEJHoYycciyxHQ3er+jz5
SX5XbwGXTEakR1j5+9arsWqM4leZDPE8xO8VzKjOULp8rxZyA0yIvy+uTjhv
mqCB9gldTYAUsM76cJrUdNwwbi/4RSonWMt0W7DXmG9+zsBUpwSHilNM9OHb
/UTXhQeVau263KDZwzbezz8Mzf+z1TMsW65O+OUBFOmTWcoClo+CnPSDYhBP
XCDpE4zYsB1A4naYotWWYORZZBAaCIeehA2BGtv3P9RgwtYN743FEmXs4bIM
QkN3IJDOesLNgGGEdpfiCU1yExZ141dRiOMoTqgHYUtRyg2KXgOQ2nRnkp++
5oqVkUc5W7AiWPOXnxtapk15xMUxol800ePewXX0yJonyk92Avk++d11kaXT
yI4U56Ck/7eltSxHcDwl6pMlQPTRkaPzM4GO8KiAWJPu7a98+5YRTSJ+H8pw
04vCN8Jx6YoF/kQ0o4u2XtRqEC7gkHjvApCoqZ46DkA/j3aJL2K1BupLN3BY
sTXnJaEPomKfyP2X/aKwC12+Q3UbvIA+5WkagCU9BkQVR5LZRSsB47dpHYCY
KEv2vA/BXW7AHdaQIkN80dWAmg2wtXTk7ctuIWqdvDbqaB690Bp1mBIHjfdR
6sroi2QAL3lV1TKlW5cCMYhh6ghMY6vcLrPMQvThq2UK1Av8ACxlQ3b1HxI4
40eViSlaYereeh1cOMtZfaO0LgVZQ1xMZORJnUG2FsW0b/rriwqsuHWh7RvB
sK7lMYDGNeITAFiS392DcklenZv7v5mVsPFQDUCudscvRFhsZP1mGgf4sZYZ
Olfy4c0xYBdIs4WaqtqDO/b1RpkItWoPjty05bgr2SuWt5vl4llECNSZlvFT
4iacdwP4IQJWaBZrKNYITN62QPdbrooN9uglwksoBC/bSqC1AFq6A5IOYmPR
er2nqF0BV0cQf8JTrwNX+FHcS8Hsz3+74OZsSMuBikA44rF4EuKqXI8GuZKO
vl5ZfG8t0HWHKnqFKcydna9MUoCpZM1YdVxR9SrH/LgzK9cp/316mXtKQ57h
4bX37WrWA7f8xFDkw4jqddbr/R3xR+aXyUr8pU2PP+oxXBA81/U72hgy8+ag
E8+K+1PdwHymiqrVXk2Rl/vLzYvvd9ZU1N09AGyo7SnDn1vi+67CFuEEAwup
QYzXsjHlnITZy5kOI0XerharGOZ+6d1IK+9119o0t/xhyYCmxEMmo2KAxVeY
NjCkbmjAEuwaSIr9t6G42dRKKXB4feKZ4iRXfJxwz3k0wCSbJ6GwFANHZOBU
9kc9oja+bkcW5Etdm/J1PmftK8aUFPsEMmGO+Zw2X2n4xLvX+nH5UzOAtsP9
vDeMZlpIc+e0KpHxUGMQpZAs7uzSqyufjyCgxlg6Vsqbu30yjIIu0CjCZYBv
u3kWkVmIyLx+uZinKKXMIg9bACP5WRhk+ygWOeYRkT55YO9pg1v4hP9SOifH
3UqT9R4q5a/AuOPRBmxNPJv8HIOidIRNbrc2dxUdVpGhasnILuSvf3CvZUI0
L5Lx0SlJy7a5Ad4Jd2E0mYTqOchK+s2uHo2TEVwczghwgbZi/Ee+1LMoAsiz
7ByygQxlvZyZ7+lTvdHlvUzEwuhh2muqQ6LJi/K3Duyz+gTFZs21jjNoK8Ux
IHoPJPORMnq4gkpLdBkE84v/vGNMGKz1x9hOns85d/rcZgy4BIEXBqpQj3Ud
R1gp91yjWvCrsiLCdxadjfjO2vOUh9MMX12EKEfiIpePjmOUSUu8KgPhyyRH
fnozv8eo8K2bvacJQ1U8ZSzQTaBqM2mfQEFYz+sx7p6ncePKkrfU589c9/VW
Q+5083qlV+wJVhb+v7DFea1nCr5RcpEMuE+SrdahoOymRAn93CDlPhlQuOHi
hETuGxomqMZoTt1yW8Iba6TDczAl/mJBqF8WJJwtbPqQ0f2qCRlrjn+MxtW2
EWJ8z2VFkWyiyTSnFWPcCREikQo3ce7+5gT+ZyzOKKcpgH8b3g1vdK2P8K4R
GwuIGvnta30SPPBAIR4mCu1/spXx3QVhf8nkkLWlbfECITqh+Mjhe0gO6kWQ
AEk7JJt4smViFCMzRK5I6DGbELrQV+74Y/1OOMx5mQAxb4CEJSxto8IVA/Mh
6LL5IdV/o4kgFzy63JMbqqmIv+9J2e1Mcl+VdCBoB8bac8lgAx5Sfv1WFwSL
dlnKaj0mxw/RkiC2qm48RJADwQuE31SzI8tFLPE1JHNPgNDpOTsCDwSnxBiC
AtUzUgTcNsdz0oGFYSQG6N/YM2OUGlJ2RwTNRPxQubOpL05xaRmUrVeHDfqE
4uwmtwHOXsnFS0baMywDkDfcA4v0HGxSrwNkmNLnW0qkyocCSZrNRK5lXhBh
ezmIV9BGihSS0rre8hbmTFpJlc/tv8JhZlAOR819Tv4Zv2TCSqsLfrH00YFT
2p8mZRjs2xzvZG5YO18CD2AI7bSLhf8jt9+wM5EZXb3cqILuuI3dYLELLhTg
x92d+WhdaISWRcaIR93ObtJgWRQffNMh3yPfPFfm+KFDom1Uf4fxrt5SU/Z+
Czi9xquljPuqD7JC8Vq9QjMvdll8wLV4Y8bLH49IK4Ml4ztRpXZ4SqusWs/j
6s641SFaboKWOE1nSrA1nC2cD0NCsuqYrjuatz2hcTMEa2V1DpQaepyhDH5v
IWJ9+7bs2pnEYJprLQV5r1G6JWyTThhc5E70GR2Vn8c0NbzGo3G2UiDc4YMf
Aai4g46EiYcdlEzNI0byX6emnstf4nfvRGxFLLD8qZtwKHXb320z2SjQWHUh
FBg0CcHoBq40d0vl3XudC7fHpZxBpXGR1QjY+4RyBsoWerY8Q05QZP0hDJoe
NWGpyG/tDKlS2yFNX/5U6b4GLwL+LftABCXQnCOmpO3ZmYLE6741jsF0U0Jh
aRh1UJ14kOVd7rpA7vae4xwudLkyXK52u/pa38/4fqnNQ+Oi+45nb8Ci11dr
nz5HQR2MG7PpxJvCn/eW1joEEDuLdNQGVd507dUhA1iCUJtU6MP8b/k2XDOy
hhOih42FhHxW6TVvlAZY8DeoL2hiY/+pD+5uRKbR5LufvSRfFYzAkeQzHMDb
y6nwtP9MaVDLQJakQiHjg6DS0wNX8eI/5VlAqsQYsSst7v2GW4GHAzoXfK2y
8LxD8gB8HwMevDRFcgLZHhFl2Kk1ZqvKSICLNiNrTtk1Cqo9Bl3Zlnz/WJRx
RNjFhI+ERDiSxGvG3YXaRbMUKZUVLlQX0pZylbJ50s1LkOBafLLD5cc7IImw
3lWmfS9g41YRmyXMJFv3hmVPZdtLxXSYlg+NGVNmHG4m92pi5F/U175IK5hN
s1W9MLvl5qPAq7bp0X60G7QjDVCcLhBsHFhwYHgUUS82xKAk9XtgMnNfNV2F
b4gHZfomgLQVgHFhtvVm+8ZVHgye095af6pkl+kf36tkss55crX/Y9wcqhrR
dlvCq+aHzkUC0jk8IICDPSL/AGrTIaZkWuF3Mpix+3cw4tPvfoBoiI8nnHC/
wsOXs6GaqOMwQ+818O6HYkqee1ycEWwrBvGfW13ZxJ6QK3mBDkDn5KFDbP0z
TtPIDMXrF2MlRcQr8RrgpYg+40MaJzCH0oSs/x+CnLZfCoC4uG6dfGT3cvFa
3KLYAmqeuq9C8TZEedtw1R/MzSkXOfkzX1NdSKTvKwRuRny1tT7i+75NOnDE
I3eac6RtovCZixTo6ZK6rvPgrI97+VQj1/qviuzNLlAzeFNLpNm2ol4Yg5E8
n8dxz20Ry2SXK/koQ74fEbQlGgxHn7Yy+7O8v5t8LCapM+d2ptbDFCKWxgKM
2oG0KGl3qafK9WopooXiesj92PbWTkduxDFkziwMfNEGfBaXFenf5zswnGx9
AXba1SLXcAoVUIPjCkffO0ZTTFM/ixnG9xlpof6yODW/7E/jhBC5jCcPNWt6
Noe5N/SkxjcMsDGz4YnIW7v1c9LcdofsuiZrSTl2v9vOtYKo07SS65Bm/qbz
NJWLXkbi7A/Z2W+2k8IeqSf+k1piHBhmfmV3YqR3lIf5A06sOJCelBRYnYMY
GTi4j6GjVQJqBs0dUnJqhpAVzzgMiu6DcgLnypEDFBoqeqBMsGoIvWujfARv
C8AkSR5GD6u80PoML+Q9ttIS/ZmWofiYCbCS2o7Yo08ONqhwiQePuxDgq1z4
DcVSx4tXGwjMCj65NyKCopUcAQSnyHz6smqDAiuYc6veLMD9ZuuN6XKVB9q1
1Sh+GFsBDvf9sh16QVTXSvF924IE2ljI/m7DMc5g6gGV6oidWhq153Uxai5w
XoKy4pmO3eB8a2BXUnseI/MRoTY40XNGtbq/JkCHYeZ2RMq2x8IWWXT8UHmS
r54iVkxbcMjYzRASbGwyNuuEe/VKpC4wspjnQwPsXMIuAQNLy5EZ/Y9ASt3r
li07d658k/z5xcnqg9Rw3kOIWQcoEG3nZwoZ5lL0P/5d+fb7OztaY8qWHlvy
xGKTvURH+WcHA3emp3nwm7LiW/M3TOnNdEPIyfujuY2g0Uj2zRvrmXrTIWks
HVwrYPJ4EvTdGmhv/6uayaEuOHgAjQnkXY5VFlOsQdkvW1VjjFwf4bt57Rd5
9gNXUl8VAsvmOWdCahX5Yy3iYN2+oJqMlv7fb2UM/XkpKQp30LnqBySLBhxA
S6rHgqC+nt29hD7TZ1Em2Sofpj/ZMrYsfM1453ITVTI+HgIz+3twFVXyB3Nf
lOCRdA8uCv9VrWS3C4Zyq5oIRSFKaIVkhVzGgVEO2jyHqx8KelU/xkHgozHk
B+GbiyWs4uPzOhOyI/HVOHbQDLjKbF/394XyQfga2cT8AAkmdn6TpGMbR4St
ZCg6h49LvqqBdDvP9FFAosaiP7wB83VUbjhvbdSqGZ+8UQ4cqmQlYeXzLpX0
vI48w1jnYcIQWnHPis7ULL2585hgoIN01oQrqy+RU7FQwyUJZUyHjVvwVGH0
euoFPrAxyaMUYR4xbxXNXbJ6DpdoSc/Icun97OKH+O3Z0w/ugGV1+hubRk38
aAuEGGIK26IG6N2uLZBokc9eEGXdo8FGDc7epfFMyd1zk1UjpG5YlLufEroI
/UG4NlBrE5wRplx8MTefuO+zEmiGVYNavLZ4fAKO1pLN97sPrQn7QuaPOAmJ
XDQyhVIR0g1gzSdKOAC9LnIy9bwCw6Ni3RwQJUdaJdK9j0sBCxttPhIGGqHp
8ocJ5CrCfDmCNlzqtFJtUFeiLm6qG0lVLXcPe3S6nDNTlEbo+5+UhAnmpBD1
bDLasksuAIMdgPeMPBFqsSpUzPXy+CUQPUxgAd1Q8hm6m7d1+S+vCDdTkCgI
ml1SpFMRyZtjDctWkCf0RUqKMWcY3tBYia2E+bIUdzvBGbmenRG5oF+AxTp7
Rnupd25alPKRHEesEUhgVf6I7z5l9LLHex4Ez1N0f9axqociiLZjv6oKFOOf
HEsd6ii0AgCaRcFPCqE+bQpcbHV2uVkzU9566j9hoq0oaqgnJJIU1YuHm2PA
uPZcWv6H2TqwRcY/GwZL43AaIUQZZMunNxQwF55SKHy/fU6Pg7Br0fsbdyam
NErm9Ldk4eye/k2jlr5fjITMDuwszKtH0+eWP+wQIcgYekSVaY3kGOJ5We2l
U03dv9lz0EoNBpGEnR5+OWZhsgwuJd3lMnaAYww987Sgw+WuheEENzIbvpvU
jfrmeKno3lLPzMQsbZNd7YaTVlFaks2SOfvnECxSLbO/NAiKtrBRhLadK4kH
Xb7oZj3GdKBbzVF9mfCKIIuxXvK0FOBRMqem8ziSJIrWvIUqf5gS+RUqk4dB
2BVZnVlkJTGWFgv5vis5L9pZjdWjhESEGo6ptMv0x1V4TNf9hGVchOHur5hy
ZXnUYi5YAPDasUlKr5oStglnXCKVkezYA3BsMBvT4cOnM8PStaVXbCcZ6p5Q
kReKJYD7MAzgGsWYPIM8vlD25jNvfvDxA2M5qTTvBcL8VaaaiYKxtUwkU/tx
baL8nG6j0XcoA03iC2K3PhZNopmx8VHAmKv9HmWZhJzxXQwd/4Wyu0eEmL0z
EOkcwTSmEvwhgkNzIdxYA33uggyx6bsh1Eai6a5hUQ5u7BeYz0CYgjW1fIOm
BEkE2ZPA+gqAv1cWnSbXsE7SvdNZEtHk7GpiUMm0eZgApfgTSKZhnPWvT2PS
3HyUUVHHdkmYfkVcZzLD+qgtG/X0KgNyh5aK3BOjMafzdLvKltxzfZ3Ezg+Z
ZNnhtLQNWNu0zEktkI95FN3y21KVLXw4bIqkv4XiQahsauxjPwfWDOzjAUmE
j8HuaweLkklmwBeB9ZnVYOpNrkRJ1K0CsgahamjLar1gVEbdgVNpotYcG/Kk
PAJ9v7IioIEZf0Qvc24wo5ekwoOExTqc6QN/zj3gKuF/TJ6LSkgT0SsvU/2r
WGk8LVEf0JBuAoqdgouelSYymItBzMOSxu9eGP7Ujwc9vg2DXZdMqz5WBX6X
zjmmMd3+jZTTt0d1vVoRcUOnuzzYKKpUp1vvN+DUeaQ0xAopXy+rgunUyPwh
1tV680VqNNXtDvadMnQJmXnJlmCXmPZEuUPRVJQANnAwDnUTjwzB31pZnoZp
WA1HYfRwbmNbg/WeH7snJiA65nHtds0lqJ6IQ7fsLijVVwT5VhSl2/4lGXOH
/RrmsCektTe8oLv+ti4rhpXQ9RO1G1hpf0YL00AlQ3PjNz9Jqu88iBy2O159
jMJ98MclKROupbCA4TyLoRXtD3vqGa/pLWFPxUeZiUlbBfMblMWKa/VpF49f
ajlT9tIoaXY60tUYKgJrVZ9cZFQbet1vAsWKXqtaRXqdN9+CPgYdh4PDCcU8
NWzoYjTc2YFu2iuO1ieETKyi3rgdB0zp1ITVcTjn1vptz+opxx8/P9NSLT2n
LB+0GYTWf0Qe+inQjfZRFOgnI1j84+XzW5mPVfueknpDcCLtoRhQlWNPK2mc
NZkYMRynGJrH7+3jRVTaberIqf0xWZtcYjQYZDKyso+tYEl/62S/atk899QP
CZgQ3HCovyYjOrWykLO/pvrYLRHEmX6RIvskFBLQQUyE7Ul3fOPMb5b6/4qz
dF82mHYS15YD2yPCH4ecJqYniGVNPkfVGJvw6vStHb5kxzcXSu8/crV5PfWW
FLsdysvEvO/6091V8UBJa4zOplPM4PDuTuOSdbChLbDpif5/YqHrlubgSyz5
8T3nFAtLem7yVH1IEqM2H7DSa+ir582Kf+eyZfBs6F4SUICJShdLHrdu7TLJ
WGMNfXg3z2boxjHMAcuEDWLqLxa+x7BrhhZGnBq73yHyWM8nsB1ujht4AwGN
SQuF6Erl5Cz23XKtn3+aXyv6h3bo4BnfAqCx3QXn+iauUPJXLYUZ/v1klBEt
F6AXTeYc1NIW5sRIT5Xh5TYA07/NdA6YPfxZ/MRg2ZvBkE7G5hkxsidVUQag
Qj0Ljh7YkCzxfZBNzX4KvIFDfLJ+Bu4W+u58dTlplKLbsa8g3pmae8n5gSPw
1IHjr4Le675lT/ee5FsdezCgkVn4weqoP32w8BOWOnyaO7fq0lkht3iCWcWW
f41uM0/vE9cnhifbQ4S3aVEL4CiggCOzR9rcRg20rF8BSOPu/T25FxH4j2W0
uGMvQGfSJug2I3d+fnyGrbrsBlwnUwUdd6RgbLIxGIDvVwQr14dtzfBTFVl+
la19LBTASiDSdFdbRF5ehbBtQzdT4RkxdLP2w6cZekh8TrTvgCyNuRgnpth2
tOc7iuUh00d8sGTcJc1kQZF6E1Zlku/XhhlizhRKK0mxTzyZjpOAckgAgXFR
CUxwNcpIn9INrUvchqTPFKQ3516NSyRv3dlX9A6A58tHk00rIWuR9lhpHPKY
uwLZ4PyZgMqXoD6s4bc4aebrJ/NAqv/vTvzPbf7gv4tp+UUQRk+hRHwfQSc9
bgNsf7Xwd+vbK9rr7y6oma6pccVQoiPSYvQmR+6g9+A5YuBw9Lms5vIFDjjD
1qplEo+oRH2WI+PoO6NWTa3D7OnW69sD+xvGFaa92m/uArWwoVgsaRLHrirw
ubwgxxi15hhfmMFvazLvv2ZeUnjvXYsRXtbOL+Whdh1z3x6uacFyB/Nbwt6I
HG+mZDRt22kCqYvP4iDx/VYXU98R5HH/0X2l3cbEeQdb0Vv8Py1DE0IS1P+0
+wdjQHPewKJk+E9dIfxEQ4rk1pW4T/R/1cdi+fnHD8FEe5h/FzTPx5VKxTJS
M9QGQRk/0IQbswcntmOq7u/E+7pWTGma8lJEa5g3QvSMbWTwAoy6/x4EiXk3
0va4JqGDfPqi0Sjwn8tGzT6CrCNQHrxHv9eXaj6rs42xZYwPKn8YwcXqYfEZ
MROlbrJJFLz4qG/EP8mESIIbMGeSZBKQIwdieqhROWx9LJrf9u2N74ufZgiy
jm/gM6ntGLH8pSgKccO+iyknqvQTAIpfNisXhAsqNl7H22pjtz4sDH4X9BNR
X1xTmKV014TRPU9WD/KWMOw3WlqQGYogrj8U4ooepIQnEdbil1gm5ovokaNQ
XpmUWACsHO3ZGeAO3kA8aIYeg5L53Cd/YRt/z5k6hWKIC5RdHxd5a2IFsEYC
y0TdfymYDbsSEUEKkvZaVspIrB7YYUP+O49Gtsp6l8qjsQErbH87UCpqws04
Hu+HyXu+NJ2VYVph1wAG69cUgGz/94z6XIHxl5pJyOBcR4BLdb8EmlB+fEap
pcjwhd4+yfy3FATN+TtaoagP+GJ8+0fRHHJ/i7lQ+BjkBAf4mNkLrxkRZfMC
K1sPDWz1y8ClOvOKVoWhlI3X1WMnVJ2OSPyNalb7qQNQTpsYK3p99zG5dmC8
jfUXFnTPfER9IvSNJwh0dBr7NYu6iRem1DPNbyrBCDIbTqN4zhq8Yo3t6rpv
i1YnpwPvBW/85/Qd4oQDae5VdXNxqtqP7IAQ0O3oMSFzTDZa6+DoZ4vov5tT
jsSQSimGA716hF8j/9lQlABLYQ7VjIN6tl0JqV1+CXuUewz521Bfi8OkfT4/
/RtZ9WGd1ue/jxFFiYkO4km4m4l/z+do7R0TrOLBA0j2jlWgIunxNsi7Emaa
JI7gZfs4huMZndyHXrMQ986Ir4fxIWLmAE8HDLocK+LCSqwPwsqPDpq6bb6F
by9kchkE1BPdymL9EONGF2LRKAm5UakKrdXbyHmVco0zFmtIPMJgkH8lRq24
exDPtHR6oJnHVzsRVkxQmoe33+pe7lBzNVrzhyytaXxQXEsSKCAIts9cHDZb
7GKI0yPAOa0vnMnqPHpMaRpQmDUL4g1+V6QOaD9qgUBm3K6EUWC/eMo6c7/Z
ESakln5rOgBBPJFJlfyB0H7a+63qyNy9mOpM4+GtYfTq2g/wcP+2cNeD7pps
gaS83J/p/9EfUuNiar4/IrSj1+s6UfhB0DLeM82RWssifssSH+mRuahOVX/d
+b6JFWie75sHXXV87+6AuRbY8PYi/lae95JId8XdNaV6eqGwEKsYEWh69ivO
YMbV6A+JF3QBiFRuCBgIbDPXZdY5EpPuMASUiqMoY05mT48nOr7MTp5F68x/
MOQFvdgYegVNoE0Knodzn0NphqIqlyCp61XDadOZKMcTmmSsmxmHSjrI51vV
yyZY+vgqs1U0AtSOKuygUD+5lCvuJcHAG6jlORlLVNlBDXrgeEY5yXaZ0Z+l
xZZQxtrvUMG6ARB8vRL6vEVFDGWPpleY4sGRnD+CmLAvX5B6lrceIaWG/ET7
ukNs7tlQbk/IKo7rh2xMRB6XvR+EeXJ8AsIuH7fdDznuSEwQXIYPGPlSciz/
o7OWVYu+YcaHCcqAzjNdEFkvPVdUvGScyxa4VicEPGP4mZcgoZLKAN+xxMP4
yUvRiUd/c3yUucmu+FHRq77OS3TlCCm5CrhekDZSq7RldAsF27a5mJM7Bp3C
FQAGEiDNNBH4bvtpyA1t5kEX2xo977VQyhpc0OsVQ788bDjFvF9uNkTlNO8s
jjn9T2AFjOGizZ9yMoKPSk2CPVft8zwWH32BMwnWWrCJ5u+whjTj6sCKfqWy
MwW4wJM1dq6lX7gLQf9eM4RhBVqMbWfdfBS4fvuMZRE4xQ9v2/HKTo5Hjx2N
6NSM9OMCfGeE1OtUYU4Eh4FWa+N9hNeG1lpfmRpBMrPU1frEyjoI8ZwpoGCb
dyQ7jY/cf7uA0mBRAfFn3T+yEDMXgP+oyIFHz35ehCQqV7RgvBvGEBfQ7gXo
431dTJKkLg4UH3Wz20v7t0okmIx1McMe+GFo8X3qXeASoRMvX5jZm/tgv6nd
rHu9EhiNBY/L9qFhDvldQpVbEFDlXDzVO608RrIxrA7B63u4WGMgCCR1VFvy
2VMfftraQG0Rn8vt9gfi47BOZgBnV94V6V5niDuvPbGsb9Z8Nn/tYNEbXyiM
JNjXwtzmiiDHwvv1VcBOiq/RqMtkZGSHscP+UOwrkNHqc3Wwm/ZxxzEJdjVH
IZtxV/5AeNjujnOOPaI06n0uMCYpvZwh8Zez74S9nvxzokQ7fuFiHqW7qh42
qORQckGNofQdl6hE+layNDdby8esCDF4X0Qh+lhcpr/+Ym2Gk+Yp0dreH0ZS
H07kbXFFOBJbG0aO2YsMOdMuWzjQXdOhCYwQKkEpwKd72ovvMDkhHFa5gfsO
JWf85E8hliuHRldXWAzmzI3aUi73AIz0RAXZxvcTNEu4SprzaIa9lAI3ODbj
SpCNMFJScjPURsshhiVnVyuDef393nyIljkzRagqek3p0ZGwpCHnZeQzZzqR
R+QO5N83ebKNmrY9cpQXMCZnZn8IBYTDs6zeFEKp2h3+APymx/wgv2uN51r/
2yV/6JG/c/zDB/WtY0blNpI+axFlxXjWwoQW9hJanf/N9xR789Suqr13/YYL
YT2dZc2w+ijSVKG+zsyAEbm3zQUjLajHKKEB5XhUA9qyWixVsnXRUL2Uf+Jm
9tdiOi0H5KvA0bFiVtUAyKECXDI8324TBKu6/TuWT3bBG/mgIWtDsK8+rykT
5oLXjSURitidNT8L1uXY5rNxce8c2izH5RhOL67XUTwXRtsGOvMiII7QefRX
F0dr4Ab4uMASrcc0Ca+u6k/RGuWZs8LB2+uhd5RgDP8GrktlbgVDngKKEMw0
3LflXM67Qv18+TSbczTFnTfXuF1GbAI9H0a4boYupaG/ac6t3pY1RbfS1SPC
l9MsAqaRZlaD/P7LVgt3TkQXmXF7VYaihav3rmCL0W3rxHfW+VarRPvb5aVN
3W29PE3Tsi8fbgPABwbZGTCPmJoIxvOqCq65Yz7JMUijzVhH9cWNlvwAaxD3
S64G1iGZgO15za856jgEwnKgnn5ekOLtUgRCn0OI4XbyEd7Ih/RWlQ8yQZhe
flUrvxWh/l7BXNpH6HULapfq9voBDBGy3i1jHWEma+9LcjJmsqsswImkIvh4
1lc8wgE5AmrKjnJ1fSgYofwL7c3UUEBpK+71mKWNhLIZ04WnHNybcTxov/6Z
hHPkyq+BGhr5y7/mn+9U5pro3wYyRffKz6FVK58ru0bJBUrGwOlNImZ2rOpa
+Fbjh7AZ8J/i1rplVAlmej2BgSw/qiilqN1ZFKY0kbY9+xP2BRaeVqWBCLxz
zRRu6wu6HNsOWNszC9c7fIsPbIy6jF0h0BHUSGkxChzG0HN5TII4G7Erd3bP
01SxETvP9ENPcs90si6oinWmUb+4Qf3i4s+jDMBGlVlMxsfjpzqduEt6dzOn
hb2/PnL+vZfIywROWFb48ImVAZpVQclPDB88yDoOQEGeFd4z7wSAILsADbIJ
08vJFbo3QLIAJ0VJD461TdZcZid6hQl6WSEJUiHIgbD9a/xVE/XPdsdEmquH
ESEDdrrNfdDKMZWADFOtLsLrdiYs9fWicyPtTKqwwQP0Gysfx0qWQcIYRWwO
+bdFS5wmn9/KHVx6tUdGQQFe5rYpA1SYIaV3yayrg4VewmVpa/A65QmJ4m4j
5OPueduPcXReG73ttn0UtRZcOdJX1kBbZV7tosuGw0heSKphYaYqhFikEd3S
TAWq8LsRyNEDG4Y153w9QTN/BU3vfK/TTYokXPyEiELqA+F6PXXawb1d3EaC
KWbxc7aCUg/hQmuYrM0q0PgGd2IGMNEjKIoHVCtv5cswN5v3PmDjOyQ6y1N3
icAIoyAbmnSiUsWuLmXkKsv6kePdnSQl2rvaa8t51e9IP2uncAHEHAOlpAx+
CTstKSp5UlWNTKv6KMhCtMpIlZfBTaqtnv+j9h0jVgLuYlXfSjoFp7L4HgkN
jErG5wHQMcH3yEpC3YD+Y18jKwjURKHttzD2Klnz6LWOj/sGrKVCTzg36mzf
xx6+o0sKYsFstXJpDYBRY+AxKdG8uYS2PQ7gmnLu1c+Z1OPewGPmyasslkut
MB15c5Be0zIY/kCWbTDRghJfm74Mv4dOao77ZLgHDx8BWxupAo6qUYKNhogG
eqsBc5Zq8Ua7w1+fsVZ/B4AiWoAaL++S22f3rOZ6deEsv65cC1GSbxjCmyH9
xoRMRmEszPJfBJ5HCIOgZDmH66wMHEdt4uudR/BUM+IF2tAxS3cZGWL10ic/
VMX73iDGH04wWOILIN6wsnYL8c+PmUloR/lQqcPo3Y50MvgcSeMpsqNHN4Z9
i3v979a6kfT4b3V2YFVrl/djuecChVJECxrWVXtTUMOxiT+r9vXwZ/eARrta
HvIYVg6y8fr6e4R1Xqt8V8GOyVdj/O8A28rmUOnVwxhFht2E0AnEgrGC5mxK
/K9BmSVp+L3bWQK9nzQJTb187rPhycGux+Vv+SFb75+FeoX+zdRAwNqQILOW
Qfpf+J5JbsHIf4rUPsF1XXfwZiCNQlrRl0lfunHjNWwgEE5fGeeqggttNUly
ei/5RCJR0h0Y2C4E8VzheXalyPL+x3DW/csiksSZYqHQaYd+MeuyGayD11kA
qnKNoIh1Nn2iuywLL28MUMXJvB0S9qi4ZVUw/JIA4lpBPLy8yogpMxZS9D6K
KpJvCc0d0wTQrbN3OdExdS7cPtC/DXv1Z6B8DAGQFCaJlUEKA4/RvRfrmlYk
b4+GggnPjKKkKi6fIjKvg05KoNTqWnKAmP0mtUKGN4H7RArUEtAB06gBx/Yf
bP8vqjN+c9QO6Q/lOqX9OYP7ZF7GSVvNev204pMYGHeuxOOujwjTPndOaDOH
Z6k3soWAmVlc4WD0Z93Q4Ka2S8KgNdUHz9sshRp1bYMo6NVvGvwzMisGyLu4
dLDiruqjyk8i3ZdEWzB3aKaBi8rSzvAJlPfev07s3PlBdKPl2UuvCb9P8+Vv
5xdWB4aIFYiqN5UX6SCBrN5Xu8YU3fmDypIhgpgFQjCEQCb8eYH+6itUyYuG
Y10HCXaD2UhPSkTTYXWrut1COYB3R864LDxV8QbuojIZaeKZ4R3vFbxk+WAr
yhraFt6w7WsHcLVPGVSP/fvAlkpQs72QWyz3mlymp/ZGeDShap6qjbo2DUTO
bNzsEJkbKZGHPVGv2OmarVUDTFUDg5YubPLfOQUCEwhT0KJxtYCFjegEMo+v
cy+MMc5j7jR5sLar2e7xFZGNOncpdRZDcXxOgNFLvB8wdErEk1EoummavumA
RWJyTBVDuTIN3wzQ0hb7eSBLqclLsDQcs/Ua2e8aTmZxM5oRmJ4g65HzCR+u
KpCrfW2ugYnYpgyt38XGkHePZm49IVupDpK55XOwL9abFD6BNvqzlt6vKqd4
UGSsuL4FC8fCwH0ekAQ+8zQGzvN53BPvU012kq3dbYOIYkKetLoeQGAR82Hq
QZmweSv50h4q3xKs3myrXSGJAAa8ElSpL6RbcnwwprM3W9Nckz1iIsOHAv/m
9klrw92XN7om1SYO4tEmafIXv6l8n5NdDArTeSatn8VIF9vcf3xswdEVEct/
8oBsbfuKbf0Ry2BKon0NEEej8S3hHMcEZi/8B3pi9nVD25GDHeu9WBPQtxXN
k2+temXwwWBCFcpMeQK/uFAfAhJVReg7WjduD7JQrWMVKjSLJuOlpEdmPlYv
I1vPJZNlmYVCtxna5KAKma/0ADbre9dhHJiSpbJdHX+ZSPaYmQhRxw8tz67/
cJR3bNyn8qkiwzyZj8BMgCjcZogWpF6PU32ZsOCsAZLqZ7fbkJPclFgba9m6
l0HOtuNNu9ME5q7Cz2qPqCvApdCr4tQt2xZEE71gTnyn29hrV0/adK/bP1PP
nl1DGojbel+ruXezBJza9FmJYszf0S5tcgdpT1BG5gr+Ot/V09dTHgbb+Ktx
dqxheCSll+pOsChlGb1fomdmIdSE35zA8biPohrhN/0sOBky0MAVhDfUD+lm
qN9qnYgvoo4XT7GIoR/uBmFU4oXns0lF/UGvW/iyCsOZun7P8TDg2MI4usNw
5X9vOjBy90+6Ww1Qws59Gpd2poEOuAmfLoHuZRYhOq8FOZ1oUe3hapz19ofI
Y4+WL1HJ6lGn2q3cWQrMhSRtcUvM2NxcPyaiB8mRjK8bnCYSaiN2TVVLIx/9
hMjW7a5V2R2mbHGfVpf1u6lySgwwL8WeOAQit8VffLAFdLVGkKrExnqF7Yof
7ajD4OdtYtHqrFEcEOu6afRQI7AeCNb162P3A2+pCaCUXR61XTTCSKsiH3Tg
RhlYNZ4ODZujEFQw48LlYTXKfeyk5ci/OF74tXn1PpuKPiV1kAEykXjTSJrH
xR/Lgq204gfKCoppxKKLypA676y7odDKkDC2vH3HXOWjj+S/sfnAZjqAt8fx
DTsBlNc1WKyzfiC97NHI+956aUQAK/rEGuhoCe/y2R8S9EUH25JADBpESI4r
pvcu0vO3qTY3w872Bpf5BmEM1RgBWvVImHdO9Oz89E8N9WQYw+7WnmMLgcK9
rBCOU8erdCdLv5M4R1Pu8TOV6DowUJyIjozQEmaqoLfSQTnXSinxbZrsRUMY
+70Ij1pxh87oZb0Y48+GpRjmFnpiPnv+sLZdFd9P3DNb/KBa1dPskFkJhwf+
y7b6t5eKnE67MOE9XHEhgzbRhp2mLo5o69EE12AkKwT2qhiV0tGbYzjGgdZs
JDruR8GmK3n1uY8ACzvuO1GqkMi+BZkyfPhMnpZaZ/rYcDoIG2+WNZKuRZW+
R0yVrqpAd9OzXoY4gHC5RjY98shDY3jU2h3WiJWh7t+8de+n9WvuE21ot0O2
IPpf6H/sDSjPBhStpsBVQd5mLAVLhpqG+dgKiy+/Co+gvVifrSYQO1TZOA1K
x6VOZEkTI/BfA5hYsqsMMD9Hq3z5buwD29nIQwU/f/ClfgzvIz/+54v+hHJP
F3kyjtFlEh0z1kUpyYB7yPoLeTYYj8KJARKaimMQI4cA7QBq1w+oyNKPd0Mm
g+BhGK86KVsedobNCqYyjHcTA8MATXfy/xKia93WZ1Oz1++Lhzc1vZ/5w8qe
Ehn3Fbe+4hsHxu5m+BFIS7p5BDvlaBpJGnqrpQIfrzjw3K+D3RTnVi6dXa1F
m2+OkezusoTmjb9WOOPc8qzfYKJRoAsw5ZjHqjnhig4dvUtHaUvyJtYbBnyR
tycf+0HdjzpwQca5xzv317rhLN5UPPgN6uJhg9DrHxwEwXrgTxiYvyuhyD0/
3thjsn7Uyv4+otATQd7f75rBNwOq3LUa8seIjgXyDu39tB2PApuaMHz6EEMx
mouogT1Cx2l/0CSOkewCnb50LJ7+hNHevTcJc2KzUKIXrkoRXbVJv6bKtyl2
Z3vCoAxNRCBjcSqyiDT4aob7Hr48BAKudathzqwozv7I16I6ZNOdRZZ7gZIW
lq02dq6XTBkt+b2Qj4iSjgRTgh1d61lRnvmXq2owXVfyPGDgU/SPyiQJ0DT7
mx8nRIZIm7w9vONYoNlcnxsU3ZkFwVDaiTFQj0goOpcbfyE4ITy6jnSXweNk
776f2ohdOZdE2Mf7dHfXhnDggko9wHq9puMmChGtQhfsTG1ncbL+dMgeL9ss
0R5Flr0Sn1Sxj/J9ykHPFzpFdjgZGAuTftkhNEXfWsc3bLfaNHK8nHmHPhQe
ObP73u+1rtrBHmedGW9PR71fyYy0hjeht1ptG/68hMo+LqIpGLCOGtaBql6t
wGd3OVCWlPz/r9b8F0K5vxMnBEsVzmRsnU2lX79QWPgnSVQQO9yvx97RrEso
JOiGKcK9tjFxkBTWHdO3hXtZxMiGcxmTrgwR7WTXaDBi9dVhRvW6Ry9aCABm
Qd9ZF4c0FwBonv7nLPRcu+UDRZeRB6y2Tq/txljGHRRtty9kUHo3LdAHC75b
QnXGAXVDd1x0KwVyG/YX0S4ZL3Oa4E+j4WCgdrHDd3JrZfsdRbt9eSdKQDAI
EKHL4ZkMe86NcB8FXxLC6ZkLrQspk+v8kvFYjZ01Ss6E6wWFsj58Yb5BddoV
/wT3eLrnGBsJbxQM//JKYpS2X+3HZJMifpktf29UK1S4e7Dv8E5u3IsZyRYY
/hqZhdq3IkSbizg/RHN2f5l6BWM78sSrScHtyuqdrei5LWM/HaS9fQHUOa9w
2zukIx8odILCBREC/dkXFUZPMEnVOhEW6FlE2EbarOd+yHLwp9oISggnAHzp
zLqEBj0fX1L4T+gRzHRjWkTAPmDQfceUlNsKAFb5cyvDr06F6ezvGtnVe/jV
HAi81VC8mXJ5evf201o9986UDFsJ5inI4ANoHSKtaar9vhU08LHXEB4mx8WP
A0VY58wEOgKqAM6U5zhjBmisKqB7SA7/sQ9geFeMCL49k7+19K9LWxHnCM8f
vkaTCgPbNxKvIKrQ0YPT656YTGhWaqoBml5v+3AQQmJV84hMzEdj58HTs9vj
OxuoF6fO/JpmI6qSUzJx6IIcra7AIMkkxg7LJGteucPb7WWlZEyCYhoc9HOx
e3sdfszef9xcOLIBIaDi8os6JLn42jsM1m/1AMgaVmrxIyW3irQJu1pQ70AS
Wp+wncuuDNx3rO1pu5zZxAGx6Y9tMELumJkxvO8PESBEUw7pRkqd1EiEjEAo
Hv5CuPQOM7rLgiWCWMColMlxE4RdDhU+QgtEPaZB9u6YEfdiTiPfNWgjatab
NUxYfAx8hx8nhk+EHeCu6qnQhSquTun29AU6OrPZHncUeomrjzwSZuR4rDnV
NY4HWbWm7E1ZUDsoY6yGjQHRfxL/HtZSvUsuekPpu5B1Bp6IzJCvxKHKPWJH
jKOogDsL/nZnANskVwvtG8OkjxeNcXQ7WycHNMT8KKLPrbgohm7eaTvXumRd
e1d7bq4tIpBCsjwIk6deKYWanuV9WZUJvd1ir/y/PT2scpMkhLWwuTzFRTet
Sso8DFwXlVra7bW/GhExKRMfLRcPUZVgnFj+0+Za1DnN47H4Qj8yweQB264/
Sb1oIpItAk9GbABEepoeomO3CynBBfDLcxokZ/fD1hOr+bM28rcj4iUKtGIl
qd0cSXdLWdpaFRLY5iWKC474AW6xxk2w+YrO6vQypCcId8oPTfZPZ0FyQ1oa
Yk3F9NSGfV4wjsE22OOvXvsMt8OGuMPlz5yDfGgwYO8nB5VJ/IjKE7NNrrRs
ux8TAd1hrF/xpuMSZxvqLiAQXpgLcw1gkIsO+dAFUhlT/AcZCcf9rdnYI404
qavmvpGk2Thi/+EcXm6hE3go1L4fl5+IC0UNOiLX9DwC9CGa6vwSPOQC1o4m
sX1qYLNRIHDAlMnMbpy9S/b1DNgorLXaXXbH+j7ii0Y3Of+B+gtkpUAND7yz
C7y+6N7T4NJxMHO2IVtucNYs1PipIglGxApF6JS4sJZVDz5qrr2dCWW/L20D
kcrDG1nDurdevxphUeRCKGr0f+qzHNOcCmV+FlRX4hjRqADCv7fK6xz5rZ2C
LL2VLoCcGn01Rq82NOPAmzxulZLZBfNOZUyLxc1xOu12ELbPGyAt1t+DO/sg
41pnFdIY0JIIkCA7IgL1MM5aPqjVJDJMA+zRjtwoGQpi21XIGMGMa7Jo+TCT
rTG+Y/Z0/7bbP69WStbHxX22vL5+oU0of7yGMyHUhnUQNcoEKbYgQrZqapdy
gFqlnmHIno2s8hbtGdvaJsBHfuvjztUJ0QpznA8QRYOBPSLk/5D+GvsUNa/u
QhV8l/OkMMXXkRP2lxBwFNXlcgKSgJmo5kSUWpVK1be5XoPW180u8z+qXGGW
QhDpEn1LFoGbzf/WWZ6yul+qPIiXuLyh3qZ+0Kl9zVM9GjgiR+E8wZdWH8DV
Bykbqu90PLAj72jb1vF+BphA6l0hcR0K6Ax7HWMlx4zBp3SiQPrNxUI4NQ0G
f+zm2sCwvLoyLD9PBnLCOrZ6rwcUXFyBUqMH0rrSOP8cG8rpy/NfhqPJx1jS
8arAm/Ec7p2zTOocEsnhEYQbVWNU+z2W5R1x3kvcIYBo5+L8XtQyXye/MFG4
xfRSf+4huwtGFTVziuOngVrqkvcIDBz8kWBrAN/233ug01JdWiyRo/moGmEK
RVGxc1KQYTfn9EGbjC/WdeAVWIiq9vkVfkHFJLnkI4rpRnz9/dQIStoYvgKN
2KFoml+q/KI6If+7tZkHKiSAIfl7hkNMIAoAWNIR5muqmXg/j7r6OxDOtKyh
oKXiQkWcm6NGOz+8OzFIX601UuoGBdJ0lrbpY9SZaV2iwsg2Zg9RyIWBCQ/p
dg7N3x6oH/xMasEEJ5ka/hd1yYVoGTxQKgqZyWJVnlCWJ2c8qnn8Al7U/JGH
2uqNBf7aZnW9aXEzFw4H1PANCwE2bT43UZg7RmC8GkzE4ZvoU9qgde4HMl8Z
6GHrackm41rYnhPbvsqb637T6sT8ah0fwLTVFr4VxqWgq70DILe8EC+8hPQS
rllKkhTl9vly24C2a8ZSSgLFYg+erRpplkOT/pC+fTdMcge/dg8CrR49gqmF
xM6OnGq/I0B+mIo2uITSD+aH0KV1sWQBa8TQct+KaC2XA9FdYVB1V1+zhwRc
axnjmXmqLGbpOBEa8PX+2TfG5sPNld2unnnK1vxD7DXz2jqS5IpyrArBhkdh
rz2WDWApFVf+I79whrobWIl6leX+yO81gToiRxZU1MTF6LB9MaQSIk9PgaQ4
PR3ex53KoKz5y5AA/X0viyQFOuVrzvEc3lrok/9SEg8MG4hDwgTKNJzUXzTS
EVV30SIxoToa24v9lP7TnsDS08ekGmlYJyXVYW9eT4nTeXl57EabgTdd35V6
oFrexlw1I0Ti1UnxofV5scN55wYT/Yj5Go0cmygfZgBUQEwrELKxH2Np8RyW
jZJeXTfEIFG4qfHgVZY8mobIKrkH4WohSHxIBdlBq2HuirFZFcIU3kBX5AVJ
1N36CSuetljKEs9LWV8eT4LGa2HHJSkHKhvEc/hvIGjLN2yy+VKvDnAD9G9g
sYJYfn6xHRlJ9Eta6RZvnqyML7ZENvenQjKCjIR4DjjyMNE1H1BOeEA5up0g
M/P+lfvBfp3VZOdwQkiYh3+enWO1wIJcHzb8IiX6NG3iUTNR6ELybNb85UKR
75QZZtJ6uAiODB8giiB4EtGzpCnDNgFlSFHQ7tEZ0toCWcESZp3XD7mgTZhU
XmfA9gTOHQJr+MRZGcKmuD687idHkQLsYPV5tZLDW2bf04zv1MusrocYbCet
jOOS/8JA4j0etUT6IyZnAgtpgppBgPf7qGGjw87LZck3UD7bC6FXNJKl9BJa
PG1ordWw4DUt0yJrtR2pirhBO6KztmA0D/1//SqVLwrrdD5vC28LnPoGGNzG
wOqm64oCF08Bp/F6fGle0+1YxN/DNDfhl4hIcpD5FLBn1h+MP8tdOuwIN+9H
M1/VSflhfRc5Suqmd7oMiv81gHArxKnHa9vAeksYOEe3cFVxegUSTcHchojv
2UQXls9gTTTmTovFK8vV8rEHMjkRvT2t8jfRBS4Dimv33b761vrzLXoj1KPQ
l5E+ZSQa2lMqydlxtRe8fDzxlH4/7/ypU0SSKBCJ6OP4SfwGKrGg/t2vm+GL
/wPr498Scf097kEQWwdbjf/QMIGYg5OhGcv37NOk2nPf1pGzpfgCUcROIXmr
sQmmy9j3GJKxcq3kN7eYQF6KDy1YePJl7/MUsZ3exYi0x3nmXIYksXKOCGkQ
ESs9u+AsA+FyltK4sawooNFfK7aaX2+CNDnsj9e492tM2l2zyyhIhOoxarI6
huV0FyWfUxZjSSjzZ86MaQRzMpFx1zdPZIjNvmkUGDN8sNTZTXk+JMh2jXwN
LhUtaCgb+efGEOgbeUiHTP5voL0u84Z9kZJTx19x6ykGgzGYsdW6O0ywNEfs
2Jgmk6o1pdBeRxKpiRw4vWkpVjaYggDRv2MCYJ9xQ5/dPtBmGKvPqLMn5Fij
V+Ce30IZ6WjkI6Shw08H7qtSjihs2g7M3gclBtdDTD9jkGTdd06XepKRLWC8
DJJ6kG3Q6J1oHz7h4FnFQ1O5+/AKdkLjAIqrmkKvcPg51RgrrjBKN7juciDy
LZdNhaaE8zAO4Z7eVfsBPFwh2l9u8WkPYqVfP4RzQIBy7RJIn0q6xoFInHmg
101CxI1UFYQeE8s7YHYd3KJ8TwPXzA6eXDYtbBHdWvO4FXuahJAqa0X8xApr
pz0V90wSkjaDbojCjV7HGszifah6jDGS4rNy96JkafvQqDivacHKQZelQJ0/
2QKWmTRZvAvUxgk/0Ocqh8hfBXWMjhf1MyVEQRgDzinnPvw4CPZZd/ZwUWu+
J2E0tBXKfutas53HYKTA9ywPIVBR/4BB6BJjBV+T9C3kK8Uui+b4H32hM3qm
T8CBr+FT0lZmFzk04L7oDx8L7FPqiFdRPvLjF9SdBnAKTgE2GorAa9WDePco
O+dL394bPdmqwjs/9hqmoecgv9B0BxyQgoD3LhXwabjv/pTMW6xogt3RGC2f
Vl7grI2vNlM1FtsZA5JvHsFc6I1pzdKGsCH0kYjPx/k708RqQsmUoYsMpZYK
Wgl3wp4vFxec+bDUEYpjPjJQkL2/XRuGkmfDgwamJQdU4+ebGnG0gJUGAwf/
K8LjswEFKXRBk/6SyY3Fo/ok6b5PVfd6sWNkfWOSifnYXcHg3SP4Ra3TQvk3
8GX/S9FhVrzwSXofuQ6J+gwcK+PqQEUv/Uwe0L8Drc8XwtQvL7xsf7VuhGkR
KZ8o4MovABM75+rslBFvuVF9E30vmcsBKDnZV+mqcrqMMOqzuf2khCwFnEuf
32s1NY8ETJYHPFLEQTuN1e/o1M/+2DFhLbwNc3HKoOrFYQH2ksYf7ckT/9NC
vbaxjhm/veWdNl1kfnRrUJWzGcKjknuQr7hbMv4znbWkuhtyiLuh5404e/et
ijJjOHxZY9sDYYxHgBy++MvXzXz6OAx+I2B4H1E8D6APojdvyNgDyt5tXee/
YH/eV8qgsWiShXsJNMIhq85h2oiOkJnDsRWwFU5mSmAYCSOyKHDIiCR37OGa
gekLzLyHHBPajqpn+tQRcFudDONDSivXd6RiW+ku3Nih6c3UhBliKDraizX0
acV4tmuQ0mnUN4ik9b7TwRWszpiwxybMtfbapJ0gGJDzgjcj2kzNpuBGctSt
iT2FEPBJYEta5KKHO/bHXN7AmqS3FHsTJHxYIHMAJMi2G0wKu5djPn/s+zPy
B8E7l7xeGb4ApspXvPFGIlLBb6uRQ5VrDGZjB49Bi1FVSJriXpYbtK9cEd+A
1yCHKVhaWF/t+8WbgaXTZsvRtwRNXkfUg1ilwXam7m0KzuW6jk5/XFGozVHv
U7HNoagXBb3DpjTR/xRGdYavRGFdkJTUE6S4sOBXiw/+dYS0sbWUd1gTn/Mb
As9HpeAjaWkxEGQmb1To/WtEjGEnzyvlFJC5QL2uWHddtOOqiUesBU83ZYKV
866LtbaB395qVuVmicRaRwpP+8ecrhgHc/V2iVU1Ec9Z80gzhpuvDcMsj3rx
9ZJwTUC6DrNXaBoJgR4yE/Xx+XfxYndhH7K+2NLiFaF6CmntdJCbISul5Rn+
xxv3kxPhp2UA5jSD9Ih5U203pdKZGkxF4MIbCeeO2yGfhJptEBqEKj34h7RL
sFaxR+3OF7pUaw85ixL4jGcfTOi9a5NpbLcct6yaqyaQzUn6AncAF+5JI1Qu
hjUmKI0Rbbsr3U7pek4cEoHKAAMjW+a72n4NQPN3RxmGunY+X1JFhsD/KgVh
4L240+86bqMnvrvLPcsJFLfxoOMjpMjh22mK9wW52pXYCzwjfn0YAmuoBvJj
zy7eaciXH/CPkJg4RRDjXLut2RkQsISIK8kfpdXce+1y4jzwpPneZjbpr6fg
BJHmx5VlFvkY6jSoIoKz4LqUpHEQDXGY+sDgcucg0Z03GMBbn4GZKmsHQf0w
A5Jssi+8Iq6v7tywVy2AKk0uD5CpBXpbKSzApEK9VkN+ZhbOPc6jVpXrB2xz
2eHq298ZMMnm1SWc7BqI/OWhCxKvTI3uehzkoHoZ6e8+dr5QrkFQ51c1b7My
hwAsBCntTcZHuhJdWsHUU/Wxx4m3bER0494aZejAx7b0fmjSOyt9XyZnCXPO
YJwxEcoE4rSW036dnDmZP6TJW2PNc3i+N/cWBz/xYspdlDfCZs71AWC6kMTz
XyAv8/Uj62FiZiXQJAbMG/ue2GGOBz11px3xUAk3Zk2g3PQJPw2SsZZqgh0w
GN0V7EhkqyLR4ppZe5H2w7JjGpa+G/strzh3Q60jbc0t3/avjnloGR2cwC94
5qI+0Zdx7ycrK3ccL/rPgN74Ei/QMqBM7QyQbXzD0BWPkU4tRVG7wf6C/Zw5
dlX0g+D3zhJW15pSIc2L8dtY+o40Mj3bh/yvYNuJkeONrmwDCWk0Maquar/w
GnNTenczt7nvE6bVnwxUUUwi56GhWLaZb9yNqEIT+85+K2wjDQ44ASX9PwYG
Yz6GxcZHmtP2njk5lSUxvMF43PJOj9q9VJSDR5HAnRUuMlJBPKhMyRP3Yjxj
9GTYsx8hOUw53yT04QhV6VACNk6vb77V5F+q2uGVAFxp0M5KX7itX9Sm6BLg
PkSP1/f2T2NjQjR0URgh5C9V8fOjStCZf/bViKPpBHJSlbg2+OqV5SKkDGGs
iNNhbLsiC5lNx+d5GWSZ1VtBQGVdWPX1t1a949mQHG173hml+QuA30bwyVxL
gICVX+kwIj0sw0XbmgF1w91gyk158NqsA5Ie4NAeIEzLM8uaAbJcz6KBnEzs
Y/2VIi3NfMvie1bWg72HFy2UCLUewy7f+N50FaJjqHU8rd816iU3gBSnD7LH
7xhnpcE+zJQ+iWgDl/v2ihJnPBDW2Ecr15UJUBssGp2JJI0Gz+rjLa/2Gyal
Ty3spgt8QpjnKxdaJATuSX6a8pKYtmdHiSm1TNsw+sAvLm6uDGRzHfgNxiDj
ZFY/1dEBHVrQ7SD8GjwnQoZKMuIPQKFPPXgU5hNsTgBdqmZjCDVZaVn3Z8sJ
XMt9olXqaeeFOi91vSuR4Nri0RpJ6CMRtlaQFt+J+6jHFV32a6hHQhroWilJ
agCqjgj0GFZrYbal6Cj7smPURya5gtGzvRO3z5Jw3YUbYMRXAkpQc+rdxlMH
h72GBgAJz4iYrBzt8LV+PtYJwA5zxomc7B3ja1SOPisMQPRaBSagkAPiMt2g
o3r0NBjEF55j0Hrkm5CUuSsJpKzbLVgIpJhKrPeHHLJKCltJ2DCgTHuRpbU7
3sszxe1H/T7z51jaBSvUI/If0zMbui9vJbqLWn8RylYy6nUcFziaFM+BFwcM
XoohTMeTS9RoK6xuOc1bx5c7TYyCx8grkz3VdtrZWMMFwY77lks0uEMHON87
1axP/b2T4OyWRj8C0j8UpBFAw911+myriDvTi4wM2LFASC4dSQPjivV105U9
fvFoCahBzCUCr2f3aCf/k2cxTgX6F60qbj8usQKeqlYfIXfhf9auPeSdNiNV
fJfc4Je8U/oq1tj77yNKbGefnwogIag3ZjeLE8NyRh10LcPLmOCUhm59hKtx
LHqSMBWN+cZJY3jd9KqVUewhADpsn0oyMSy5v4KnlJdIAM8ICbhdzN0VON9U
Xo3onT48qCvzIy2kfkGLIKLmBHBqBbxf9wIXaZwFhgoObqIWq5g2aLjy4L/2
E7AVUpJ3w97hL5EnDMncye02MqM8JO0RI1ne5uMm0qNEmzhT5SMcv0bm9M1W
ZbTjDMLYdCRkpv+ePZOWHxHVZgauABQ5qp7zTrP4aRWcKK4HKoJ++hOUWYSa
7KxEvRG9WeLic4D/TLM73f8eW6D6fdk8E8tmUfSLOpuFkP4ux5Xb0xGvz3i/
pnm51lgPSbaVIzoToB2lEvbnHDlq+LPSrEIBHDexSvPSwawR6ufd+bi/YOaN
NXbHf/QgMn75MyVN8bIYJ/5+DfI3uL0Fi2L0KfYDTluYVoFNeY1PK4onlf35
iT6zdwKnlSkDS8Kob9FCmD4I3NNNNU+BFynp8Mg2QpdZn+jsWuGOIUZ2SNaJ
To8qugn84rl7k83O6jaQhXPmeSLQgTH5cVzLaa1Xy8LObj8m5trRWqIS8N3O
TQNYAY6aqYQ5hJ9dtidTczMBgG+sFAbczGxTNA8I75BZjYzkZny7mav7ZZNW
K6pYrKJDOxORKC9v0sEVFnN7sxLJZM8V1c7OT20gIZGSEhTbQ84fHuXOZM52
i+6DbWHCVJdeHfOE7kgAc1jWmFd8WPqlywYck/xMl/ugwQNKNxFko1D7xcs4
BTYASxiTDi+kSLKWZ35LHVCZ/6JR4ooV+N5ybRmgnoDt7JvyliQjSnKNTsbo
LnFNN8xJ1ol6+gnx3786kcbtFFew8s3VcpcKDAMgF/8GR/iKhUvXMEdtfJ9Q
3s+WmyQgzhP7PByNF1Hk+23SpeyTtHQuR+eqG+wIoid4wSck6ApXzZCHcDhI
lmpdOFP1UUUlRK5qPbHshYK+E3F2Zm/m+Ja3FEhod0tQ/RdD/Vha8Hr+gVkN
NP3Zdf1TWamEGdv2LOKAYBG30BLga3sv2ZIBAlM7r+EWm4IbkDf6Rs4KHbkh
MQRgAuGDPu7X8OrJifhuOtsF1lfZqh1zFUUsH1qMK+XY0aqN2heHi1O264u1
ijhcoZclR2BeYOm78Eq2eJtlK4EHQWwvEjTeG9XN2ViCP/d921BSgzdVSZHd
1TLL1t9PUqEnJqB4qqi3OiYuVKddTwua8OXJzII52DUo1PApy0yzPBWs4zJc
5bRIm6WNZXfVNkSluNgvEHTG7yd6YGMcHnzi4jzc8Bz4JY8Pz13gx+Qbh7bY
MNUJKgaSIntDuTLexjJL8GDGlQ7Xkw7ALmXPJFgBes9sHySHtcavhX/6O2dO
Rh0GW89pKOWxIiAZHE94zGBdwFH+SPpfIGU4oPomCfkmMctFaV2nMTRLqLIQ
1gG+iO4xrWHxCTrPiB7HSM43+NI2QJp90A+/y3DshScLJqw+uCxPNwt8F9cR
CjIA0h2TW78R51IvA87346Ci+z4vjgnFw3yGqfaLp0y39hItLlmuPJ6YNb98
Mn40Y39V/D9w4FSfrZeti0oswzAY7izPTbHsVXQ3Yz+Tnx9382d5PdcbLXTO
uxxKyXT8vcXNnFEqp18F09Lk82zlZ1MNVKh8C/SofpCBMShruRCMezuGZ/1u
3HLPlq7V39R9tJvX157muYRy0CSK8iEOU+RC0eJYqOjYb6Pd3IM4lrIakRQW
mkBTNLkZyqDZskKLSLl9KyEhqVxraVAf+o6eeqLGGkD2FpEaamIAguHCY1wg
14EcDI8LQL0Ni6wP272ZfC9s2FHfISPynQS9uwDgQjHyhUEAuEBG0ByejGtr
3lghRbQzvhQ47HixH1zfaER0EyBfQbDtrvUd0ApN8FYWitkQhytB6Gmd5pTk
RfkoLDsgs76raTqWZEgV9xuYWwsL8OFt5xkAON5rLHAhedUcBhBHm2zEuaKH
Nv/ANvzRL+6VqXGjioJ4a8WLR0RNcwQmG+pEjuwonEuZ8EeyBAbm65WSZ/VG
StAIghRwwRwdtInXXv9wVgxaJ+ZRhE/wpv8zrFfAb0xhPdSWaSoTkLNm8ke8
a6UQSxWHLEeMEVhuPsEMAyH2p5S6fbbTLiMo1QGvuCaLjRk/o9Jlf+CNvaYM
0aA6ZwFTUWcpES1p0j94cvuJuyTWjY4L55oKpnK+mgbJmnXi0Ti4uaUg4Fni
mBX2RskhTv/Z0wauKKBNRqZcNfYmdJQa8ajDPienes7Jw3SSpix2c5A/qmAJ
Ubjy637V7oZVp060qpR7OIPVfTNs6ehi/E5WB7CYh7Cv2c9bNlBtb5YKvCmw
vx6JaWMTC25rb81+i3s4/a0Cgkwe9d9eDN4ZMZi9JKUEacbSQ0XnW8WHz/6A
6HuYZ0loGvdECj+WOsoDeY0tmZtIX76Qb7WR6ImNihpsFxi8rEEnommZGsim
jNlKfd5Q6CMXanSHdxHjJMMY1xTqxt+b9RPPXWoN7lGWSriauYQW3FEusumO
rHQr6xSeT0E2SYTEmW+2NvOJY42SJEW4GyPgHUTCj82/SpiDjj6BOExnPy1p
FkVjeft9VFoFxqkJoLYoPn27/VH3eSkQgI3nGhh/130IdRvU4SXh4LN1O1O0
pFGDBrk5fPNYkTkEmg5bEeoqt8dg7iuUUTe3Qn1X1DERf5csui7AozfCoIZ7
JEQNPO39UdiVXzXejCvxAgZN6Oy9UHktWlkU5EPVUYifeLSMdLvWjVpUmJMC
PE7x0kxZXPcjWHJdUebDNSujwfiZ4Y0AHKVmE6k+9kQ2eymn0uKRlsVhah5+
g/iwHv5RJRcksizQ+8jMuuR3S7jxPB25TggLt/IqvPBWlkLTYZz6aSz6qAjA
EL8A+T5aMCeR7iBE4zPZZxDWCeDuTBmroZCRQXST4e67dq8YX5/CJdop2KIL
CgnNekVMqkzohmB9UYPhChEqkC3ph6j9w/4eHodjSbr+7o64DvmJgiVLwkBp
54ejtzbusVosbBepmcJU7qVh+bRsPm1zAypIR6zusBz4KHPTDmOO6rl3ZiNQ
ycNMsG52KQVlq6azRolFq50l7YYmm5uk4ziKGsGVNCbJXqJkCviOMwI4dIKG
FN5YjfmHnizEiv7pGREuU2SGplHlNdZgG1X5WDiXRgc/M6+z+aoQ3Jz5CtUr
yYcGoe2ONFQuLYeZPSUiggrTG1mBLLxV6auRVsbR/3ii3bGijjKmQeaQHHH+
qLBJ5OclwFREtK4Ax67QgkGtA4vdql2SjSxKWWDnOoekKpzvZZ1jkEAdCmmQ
KJEwd1KoGsOqQFF2iB536hWNIjiBNhH+FdDc9BHUaLhYZCKj4x88l7P+XkHQ
PcVb8hd7BG3r1zcCTmYnKyjJa5H144Zvj+EYUyNyX4h0XEwajM8yI/rFseAv
WrHXFYhhkdyxD0qwZlOOb6F7UCKQlGsieN4OiFnft5j360761ilgz7Nw1ip8
YL30QUoIQFthqh57pOE3d8yM6Fwu3uA0xwroPr/rV010yoxfyixRhIpf8AoY
qn6S1TSVFN/EZsoKrxrpPpB0nngWtm5DHWpJKAjGcqMHQxbu4qRZPv6VL+u6
lI83IydK60qRb3cuSSt2XJHi8tYld0tmWSSJoZ3b9ngp6i1eYKu/P3ZnkvPt
7EAJM/feubm3b4kR79kR42yzgNGkpq1mMz0buxmPNchHvleW3GJgeIWKd1Fq
YvaX5d5TqXCfCPZ1KmWJQUbEc2TDGRpVx/maXxRFUhKUTYYhikkILsEEVNEu
cbDyOk1sJ31UYB+H9AQvuiYd+d/y9ZXUi9IMuhp20mR3xx7+4zeEw5jdpxDr
MYYAQWKUWpQZVsCfCyz48b2amDeaWfj01qCt5ybVcHeyRDEYH+89WiBoCwKT
YdJa6OxWokTYWf9/54A3KgSA1fBt+3lWQgIMolRLS7i4WPJD5zFORCnh0BcL
CLt1LXnqLind03BbVpJJV24c56StPqB9Ok8+fcUMPcrsGzM2GWW6KyLXIoHs
+A2rSLVgLFtWHN54o+FM485bxztKaeoPRNyO87rVez9Nm2W46/rQRvNhzJM/
ktVZqzYc+FIHispE11VyVAv/LVm953mxi8e1PjP+/WHNoiQBTJg6O2oiEQqe
zAY8yX6o0qf3b5pieVUdBn9BkVL5KFTOE3sP7Hc1DDjVrbmdPZyzFB9+Tyr4
uOFBzYBXkuIjX024RN8s7m+ktB1oBUw6J0LZlLrjxu4GscoKFn7Bc9EvnGE9
LzlAjx6vxG2W/bGYlmm8B5pCDEDIVHWVzBlusIwldwAvDUXI2I+8uW25JcYw
mQM9Rg6P4iyOjLX2hyFnpyrJ4XHT0mvNwFY4vWB81R7SmRJ88DF5Daiqjtbc
dP/+VYRbv+5QlSu8CWUuG7opkcGCd4Mc08W+DPXg1xjC3sz3CVPp/voSO/AH
XR/x+lqcoIktnW8YclEp48YJRT8PuzohFAVOyHdlaP+NiX4DkXgG2RyQNL+0
Ev8VEACSRSK+fnK9+JArbszZCRp+Xj8qH/4gu8/l1BjM7fMoG5Z8BG08ilLI
y3SAAhvz+tn/2Tp07iQM7w1kF0mwNY67do9qPcNnHqaToQM/bHhoKFfery/S
bmNfQYnkPqmQhN50UoZ5nMuJxrvR22iFa+uY1zDvnHJVJpcDb4eLzbQOgoY0
dPQKhBZkjXApvh3+hxfsDNeDsn6HEUkJjJeJkG19guq012T0eDQi0en7Kaxo
dKfcU08PQjWnwlJZZIlvKAKwatQv2y0AjvPK+fspPX7+en+fJWi2I3qFt9YL
OOW3ArVNmNOXVGQLm9HIvtfE3eD6oK/IIqPKZxnXSflr6TlptLjb4ZAshEqU
TIO/Dxvm4GyC90kQIVvDHyRUES1/4nnqqV7cEYYkb8YobhPgID9carqFi3Ny
kFQiwfU2vHoC/naQh7VWcFCsyj3ncubFQ8AVLry38ljQ6p6yMvOAtEnxNscv
UkcsCMXtO9WV1pS2Prrz9qT77ajrKaAYnk9NsM/YThgZHGxQyPWePYa55OOl
T49t4sr/FHsl8qSiSXqOz10aebh605fewElwfEzYsoWOeL0ElD9atEdp/sUs
sqRGMSx6t0fCTmCGBfbvo5n2xtcqyewLTfjTJj3iFqvZ3GyqJqMXlfFY/Ncb
u2a4mcQejPs/Ki4eqOMGdfJjbvXakOJtj9jgYi8PoOKoqVu/ZgwNEh4WYGZ1
X/7T5e1QlR1fuMZTmgdaoWgFui71QgHA3LsHPZJhGPlWhRvPjm5dwDDSFYBw
mjAPc2AdCXbXhPsYpwLUW+4KxzuvxT5hQJDnO2EjwopaB2vmlquEr2owTc1O
jxtOurfCwrzy1M+Za04vzoRQAG2Y4X3SidPInU5hNQWk45CLvqIWvM5kbXfK
NZop/LKOWWsHTpHHJakKvh0AyYRA8vxoh/kqnZ2SoNHMvvE6vJ2WWxjDPPnd
cB5yN57nAB8r0G4njjgeeG0vjnfFWp4C/7JHl6pjSJJL6Nbr0GtmHtQfDlTm
yQ9wME5Osyih1ZvKIA4eVdi3qoEuWkIft8rB9bXewafLS4ViglzGu2kd1DTE
Qm9FdWyt9P5qM7n6ugRM4VzgsfVFIoscf/NZBrmTdhGxioeXEY84WEBDaV00
pMFjkbDgk5a4374SZCOtAumomBnW+E/Vxhc7ge3NpSeilsK/QJNrHx3EC7pF
Bn0UnWFoMkNq67x86lLBlhlfbd9Th1NZum1rmcica44ivBxixldPOBHshVjB
BD8BGFfTWkZueAzmMF6Yyl3qrwsZLUDWcrrvjYNloI+funUvcGJwTr9drZJw
L+edDflv2MK7fiFwPeMMjzFj213jsqzfhMXGXajcqztfBRAtkUXbtLszXGnm
0/PpDCnW9HSEpDxLgYcFeCkOqOxsfybSY4I0p5clZjpHbHFpT1/HghTOvewZ
jEcfSsaM1W6e47wrPH2WFpI670qmxpKI1HI2KNdfZuUCF3jpup8zLULViOWT
Cw+pNLyytPVco8zKjKD59ktLCyzVggAJfk+9fg+lmOuaIYkGn0tsFvmYXUaG
HER0FfdB7ItIuCsC44wLyoNQzx6+i4wUpH0OtdfQSIftVfcnQmHXFzPKWfRT
xzKdwLOiU06VCmGYqqzkARkmk4xsd/NomEadmb7/fHBgn/s+LG9tQBaATWd2
LOiBerKbfeG9EjM8f8AZcOkvX4BoRd7meFP2Z0XuveboMphbUnYXuwlK5mRZ
zZizgMIRex6LvdEPdd0R1rmK/2ENjHgVmmfxXBfr/GbDgqRP1FTSCNqiplOq
/tPlmubduja5xuqGXl4841d3EDbk6F3CZqFa706QW59n+B50uRlmvzdANsOP
233/YTe8kjq66/miUuNLUcQDYPsgNPuVMjE1aIh0zxpZBnrTA3olPxkLUzhN
IP93gDh3TLD7axrjuyFxlGotTPF0pdYZ0qeBeSmEiOfjI+h3veQj0jN3Jq7D
fYpfYOIuCFF1B2oQBaFaxeNHfcH1yRsMC154WskEqoE3t2EYvR51DuqZQEyy
yLHKH/StP9er1bftWnoCuV162Di5XYUkRl7yHsLpvFyTEynRCJ6Jy0y0d7vZ
no/lmY+noXRWAnf07Qg2XZFUvEsotZxGgs97AMhRvph3HF7RQ4eDa6LomDAP
mXVy/RezJQki+nQEL4rkrzZnEyCITk/8fjeF5cZTnz4fOyZ2Se8lll5xYqJ6
KFf6m3DW8NpbPcDiWfmFCRkS0/+HqwrxFbDdXwG7vfMZivPZ7vgOsi1QClkI
C2auN/YotDeoVXBlPsA4BhO0TS23dq9+rpjs4kh1b0my8ZGj+4oHmVLtz7Gs
5WGPPwTBwLY/xIfvlBp4td2WhaK5rppJewyVnKrGGdDTObDTk5duACIUlZNW
b2Iuq8hU8QXzKhy6bNMGRLpral7Xo7U3dbhj3szxNIekI5LxPQgGd3UFthRE
zmPZf0LuUoP0/AlfXnyNkvugEucMo/O35poCT2eidrtG9DZg4p2Zg2FILSBb
hpiILgFHzOt8l4dvGh7orZpGPxG8PPPPcBhEkkp58J9nZiVz6gj7scrsWtCv
HDrg/M0XtmIqdjXmbIUHt/F2OuUq5LggQMOuMM2Rkyw+hd6xDqcHoB/ehQzl
xX3GANKxBZltnaWyDJ7D0NkWQk4MArtM/h4f24dhy+9VpJlSmODCHz2/4UCP
7Y7TlF5qsoNEN2FgFFfoCEl634AK+sSZZTzruYnprQVf5rzgeSMJ/s1CUcwu
EH7vZhsJ/vgOI7KrdXedO0ASow+f93jUmttjztpfbUMzecZcNsDNou5xE9hp
jzgSEOVUBe5toLG6bUq3KxUBwnj/vRnjs0JfxWae0BBP5bDSpoi2QVyxdha8
ABl3VmMnh6ecgBSADmGP8PuTsZ9ZyFpAVXs49ssD0RJMvRXClkR1YX1dcoa9
1AKI0XZTZqEDSJ2eY5mKe8/vEI8u4Eff21d2s+pl4A2za+oOlDMD/YoDl/Z+
ROxb2AYr8Mp8U/x5TaE1rsPs1pdoBjU8isbpUpiqx7uHzKX3uG1Yg66JfqOc
Uz9aWZW+lQd6ybumc/91B+2+EE8XLe42JYmnDZLcGoaFBj1iMo3eaPgBzU9L
yG37B99b0caSGr4xsRH4B2lz3PjUlx0lqIGaozRPb7zROeUO8jVkhNxXR0VF
3w5t1WoHMJGski+Ly0zZ/Hleeq1igKopqugZHnyE0pz8x+ByD97KXfYo33Xs
+dBjMSKlm1MLQp3+YkVN/q1w3r8CjGCm8ak8h7vMiSe4NQRlFFSPN7v+Ylxi
rULYJ5S38DoroqXeEe9uosbbRCsEF775IErHUo7EM6e1pv/nfG8/qnnGXefa
Z9HzT2xS5ixUwS81ah3SHzglgQhndmNRi8zu5htBBLAdUdwNBlFZhO8/wXE3
sK0CB78YBWywVMkgzblo2rJlfYdcnar1oifaGO9lb/UgaUTgRSI6/be6CAQy
WotPBX4jj9+h3+hrE+VWM7rca4Qcc4wCuxeqvjGHsEORW9e5BmZL8QykwLWi
NrHvhDIZ3Lbu5RqsHbYBMbzHrAHh/3VljQuhBMs6aFIZiusGFcg98p/e6UCb
RDz+WmNqVllm7osUsakG+wHLf4dioj2W91W2Bm06cniwHRGAgKNRr/X18pk/
E/zxDo0/LGPdQIfxFwxyN63omM1eyBSIL/Ye/YnmxCmc6sx9glPTIyT1uIhE
K8sCa3OigH8uESzM6xVxsFlcA+f2hxEEs3S+2BagQx+VACSKe9Lu7qRY2TyI
w+Vo3Hr55vjtWBtyFT3M8cCETnQimaKtqLpsn6dHdEcrmWbwd+WLgfNO0I9x
RUUoG+/l8DpySy7JVQ0Rwep2JOIbU6OfXiyyGtCx5Kotum25msG2xj7BCLTu
wZcxDayqXNM7wJMRXC5dqUuFsRfBYDxgVP525YcQ13l0GEORAacSb72Dp29V
tACyEYjMoujXJWMi9BUv17dI9QO2/Fldbp/qaiNzbJKhVeyyZfJtXhMhNNcn
ntDNpTHmlCje0pklp3HL1FjogQQjdpBgcD4mEWjoIYIQAZLtZOQsmKPixasi
RvCWZH4pMd7sJMj+GdcVwFoXA14B2hPZctAVPIdJx498kwyBf6uBd1xexwCX
z6srdFOcXvyyihPZGJK+vOqJ3l0Kv/8ZNiBTp5t9+MIv2Yfc37y2o5CdpDT6
50pKLMWCahsFIcT2HJ6rxzC+kF5A5n4yPMzGCqR+ndiA0AH0knkWeGrYtEXi
ovqrHh4/bBR+OVy/ug5a9hZlTWxp7avdRSd/41GK+5HKOvyHzcsHRD2Qq+l+
7vKz0+zCoSCD0EqMVMZlPoUiFz4C3r7rO6UnJB3EBj1SHaL3z1ZSuxypqBkX
3a9OPBUhzPJSLPsqyG/Qy0oBMxXbGZV+lw6XbyP3tF+izPzmqzYK28DApHWb
X01vjlaUk6GAvvvI2zoOEvcoGK0rpZ1Q8vOlyn2+hygcOeetV2OZCKN9t+sK
YY29QPgeMVJ7XPkFHySmunyLlQuN72MiWQIYUvANkfBowIhX+5D5rEBf0Ako
ZAwkhFUotf97JjNlAdWzAYXfimEmT0pDOFGoFvXaSm5PYdjQY38wlIQdqZ4i
0ScK0Y8zelp9QBh8KmulFWENhx5xRA6Rrkb0L3lu0f3xaHGVyc3D0ag6RvPk
MaVmjf3oTBm/NOg1j0FZ36K3Iz1PUoMqnWcjcRbBWQkDIXYdM625aB7o23pR
b6Icjxg6A8xijeGIiivHQ+a2Kcq5r0ZvhHQi0Bb8MUJD9udFg/eaOyuowAzj
3QCjXR+EXGC5hQ4ykti1JHzVnIzboqACIEL8+tVvrp33f4LCN7+a438NNBhj
UR3b7hR4AESZIt4M3WaTzoAsZlEl6DH1Ahtww0Daz1ewmrAiLFFCVpKttZRd
z7pXY2TBGCFQ6uNVnyjz6fb4+JDjjeLwBm4VBtklgynzibPGfDuNFBOsujKL
tYGVSyh4lrlB/cSamn20o/hEqZA/7vyZU4QaTaq7Rb0LW8sG4vEfkASqi5ud
wDvyu2c+Fmbswz8XCXZWOFeqAXzWRemi4sxKDCTEgid0vmmTKOHrxMbC1Jvd
1fOEb/APvewfAGBmPttHSbHP0IeP8b41DItEKknJEu5ht/VOK00VteMPwPWd
ZPjQQRtNVKQF2sN9KKcaF8+P+VYIvz2tplgpFfQKXfdDBj4u09bVUxtvPHf7
VMygDxRRnsAptRi4/ZBfrpp4MSJV4u4tb2Krt8QmZ+z/8z+d6yPnUL4w67Jc
OE9/l7oln9UpkWuwGhDoS5Yzr9grre/TB6tKLZBEWmNK3meA3qwLF5rG2mq3
ftxYoUhGqYIk04+C3LruAU4mMa+4BnAGsszhMCENcwumcD04ZFtjEIorxAZf
6DNMXihdQXv3FO0jmYgnoF3pkHHW59iawimjgH2aOpvnRNoFyfqKX10q6Pkz
y23G6fqUmyfB4fATP9dSbRbaHBKmWDc2p68RS27Kyrkad1UFj/wbHZQjrOec
iNVRyhX5P4WFesJQpNLGcfEd1eUd4aghHlqRaAkI33YKxwD75/Pql35ZzpaD
RO1Pwi1k6U0D0Flepoqan+sLXVs3L2msatUE7n5wzrzS1tD0C6HvUgSYFSrW
dR3wBcFsFL/TmzYwC2t8JU2ZuUtdbAW/9M7FHyxAxOH3T/n/Cc8EwyDmuq7x
yfQpj+CQuquQnoGyGD+czGT+trphzAt3u0XZfIW3ygFMSYaVk1VnnT3U5XE+
sPqbw6LJk8FJgmjLcU2tVB3lCzaRNCqDy7Y+nEMUBTeQe7LorTCJsJt4kWR6
c0I0sKs9lcEIef8jmx7qbjn+rJe0c8Ar0hVR3xCufByyk4eUFH09tJMCAKCD
RwepjfrTAW/m2d9tGw7LLwbHg20VpiGNR4xedEPg0NXwxOK62abvOb/80Pox
KbHzJT9e3E00bDTSKuZB3bME8Ue1gL27HinUFql02LfSIj0lMfB15t78V+fa
TJFcJKAOYtDrGDTNh9mJRb/FDqINcYtBQkVa5XVxn9BJcpwnSRrrQnZCdXUF
zpR0yDzCWy5aobaayYdTXdyqy7QG5ZXPRrFMBdlIvKXz/tBQHFeoLXZbj9oO
ck8tkBTcatQhAji3Vaz8hBrPWfllDEr88agfDuUUdHmhG59RQBS58QLCG6GT
/kLLMuIuSLpDQZIe7CshgN0RmnT70ICcwK4GgfI6ndE8sZ5J0ihRd2ftAPDO
P0N/i4fclTQQ+WCrDIWHjsjLDm2XDv2aP6tgEmHbEDJcV9xU3jHiD17kpkBB
aPl3d1WZDCLMFgeFaOq+eusCgVM3YjwA7JrPVqWo8ofZOljJ1NfpvqHt5hPm
N2jzTRK+2cd94aGu5YcLf6wBmoXK6OfruHCQdQnYzO5nwGsSe+smZj9PiWEV
nDtm7iCWtcHiljEDycrnaC3ByQrWlQj/jvAZrX4kdiJ0p+fcepoRJ8pN9R2i
4Ww+GBFKu4yn4sCv9LS6daPfxYI+3w5JEzPNoU/waiuh2HfDED0ZZj70AwLA
XHtjPci39cKlPk6Gya4K3fe9sF0aWBDW5m9kwhr5MmWlo39Z6CcA94KHxfVQ
D9i9Yx8ZJ4MK5PEaHQa9tUxAQ07wbDievOREBIFm9jTTiCSXFOWDe45IlVVZ
1vxoZmU3t1C9PJ5QT6gHVRtCL+vLAUt3j8Cfftw+F2Hrmu/2YDumPsHunyLh
XQEZxGVU1Sf0wnV4UaGZe/Z+UxdHIN64ouPn+JOGYg4uhcvgbFLLsgmoQEfF
4F1t9a/RXHr5QUdablsD7OJcje8yPyknVYCEZqUrUAndCexgBi1QGm8+P8nL
wvkO4R11l3Y0Tvt8Lqf6/XvC4ySGBZ/fs8a/+K9ryBhtj+s6QvpPigTmCHNt
KPhbhmUQto+r/1i8MeyYskBZ5u7M4Aqiz+14AjOMEnIZeT/3NBWC/94XNelF
FZ3oVlGBBzVOHE6KX6WG6K48r8s7FIlE10jn7FA+M2ZV6g6trOCegoUZMtxA
w1+zv5RqpOkEfviDAJpbZAvAqf+6gX3ieqjum5LHPyfPA2H3Ko1qRVjpiGbg
Cbo/U+e0I6PFuo7JvWYUgekoBR4eKqKJFJmMUpb0zRh3NNd1l1WZ2NszglA0
lqFJWPaE2w3mb8TPx2C8NypZyStqL4QeZnt5b/ltaMeayuM6vwjrAxjpZdoc
SjjLihzWeGTyv0+aRMYuQmACQQBp9+PIv2T6NDvW9Hii+jbLGyTIMAxxjTIs
ohBM/n77f5kpn1kD7yE+zhDf2bDX/lbkKAqUjWIxynKAbaYX3zQwQwpfRrIN
eLcuXEtBgBtiF1QBFwUhB5REOHdMdcrk6WzfPZ9Zl4HW4jFr5oOEAbvEF9xC
4zQ1OFWfnHhRWW2OBU6aZdg41C5NlwJMOWwZCcLX9+R4ShA6cCx2GwGYQV9v
0l/EAqBLnizFqWZtyY0jKN+LlIGYeOm4PP8ITarKXel+hGuzOuSCO6RsRtuy
v54lWsBZy9Axql2klixBrsjIaqjMHp//6nTCnlROq8hq7qx5Od1CLs5H3GMP
WmUTIWnXAp0Fl/P8krx5PZy02mYZXCIVdQA+ustRkB26oonkNKJViDUWMytM
VCZkBoHt+r7PXDiHs5zLdjsFC/rqgXux4Kx6Nl22lu/J4IC6R7Tl4k3qY4yt
kR9ObkS5vRfeQ330cmP4JKkDxYRffnK0GxXgRx1RTkbMDAScj1gps3xrn6ek
xKgSbfNrax2AazPxHyO+V2tZdufqY86GL0/OAlpMjKOIUoqckFZdRtHB1X/0
urJVkM0qgPDI+eSZZkqqz2LnwKUTeWK0Nw4dhFxBf3Gv9Ih1h7LXhEadhv+k
14pJ/srwqZargVa0l9QPqux2tJlFl6LY2tRFeDAj6JtnQduOKgfkWqLqZImD
H9wC/+YyOADmnm+gIwH7viG9Cq+kpJ2fwRWSrEfg6707R+KtJGaGCNP3XXPg
6zTZKSUkzCh9OoZysOOUjyDW/TSIzkYW1dUMiPR3Z9ZPJmcPGyawcGWTVwe3
ZcTN/2W01sFAS1yqcqO8649lSpeR6Sx43aQRO+KybB5XANrVqszMWf9F9HB1
0zc3wv+lNPpc2BAjjtuumSPyckf77TRTf5uYLS7TdpEdAIrMDLXvB7/0MoSD
eXR2aOSFVwA9Imzt3yH5UTIHY4i6vX4T6eaEDWma2QjZJsMp5Oq4irzHg7ck
ng6crlnUjRwhlR3KbLz6RjH1J0Pr53pdT7JFozeoBHowlwW5sLNb+T80gkz8
yRWXbdDzl2J5EZ6BEsUArhoWppJQVH4FlLibsh3KHPK9AdUBerklER0xfK8F
4Zyl/Kqqr+e/aYkMgovtzUmFmhvgM8sC2FX4ykqWuW0ACsWH2fO790VUgs/z
0S4VGkTLefNQ2XIuxK7nCJiUG4wIALqlR8/sw96DWcK88fO6PzTCEnDJlw/v
qWOh35YRPKUqUFG9olTS4aO3mR4crnUx6JbRe9MhkmzZAOxHAy0ZWpFmBOsz
6gy16GXsW1rGS68WwW2axojx4AW93uUrnHpMnkvFF7LH099IyC35eB1ZHKIY
1FDULjHcnGC8cL7Kuszy464g+6/htumcK3WmjmB7SaWS6AXfRqp3GdA+2Abu
q5PyhxPJonMY9/v2ZsKfRMmZ7t+uUaLoGGfVeFiExezAQd9bTX7Y+8ViSzSs
4sOwZMaFPOI5Iafy1Zsajszd4C7lk/wLwKycaI/Eykzi0Z9Zs5iq0lhKL8iy
WV8phBFgooww3UBUP16FQz/54oOUXJBeV2yLqoLNkxFiEV1bvETJnm9//aWx
9jDYQ7OInF3tIJSLth3br1LbmNqoqAROibVm20DUin9UL41glzPH8fVgChu6
kytIQ/T21947wMG8jVoE1xYkLTx/4JsTfEtE/caRLhSC30jegd33r++/UHkm
PvXh+qrjpvLhW5daupedkRTwuKS4wasE8ZGfgcHlFTWxjSBQfdLU1HIH4/sc
CAOat2t5TLP9j7YABclQvMjY4IDHLVKMTg5rvAwWebR4BfihMvei86m7RfsU
SqVZYa3VPujlA4ws7RTAdCjgrqu7znUUMdlA9LXK7izfPT+5oG3kta/wpiX8
LPSNMhu68Q+n17/tE8irTwavBKCqoWN3CRLXPjA5ctknHW7WAhOHIjTA1gAL
cJjjq/cP4mDoQerv6DNiFbnVM9JPUEmNhHBY4noGHgtYVEYUyjewjWZFp9ER
dsR0ROgMUau4yGfhFvYm3mhrlat8/NvwvKXUYFsEhRzSdSQA5sQg6rUX+AzU
7ufMjECahL/9DbACEIl2LnT8LYYMo0ImLiBn4GCKimf82bIiggJ5eh7IPCML
l+ZQEjdCvy6yLzToa+jvn1EmYtGB+c58qEAhRlFTuXiCSatHB4DcdPYLkUFV
tDnNfwGKGpkGeVewenAw4sLz5rbDiCrgML8ULbYhU/z8PhbZlP4gqUpA1X6w
fGrkXq9TAp8LomyzeLNf/QTed6NVGW38QXlioPVGtecH4yW1TvS100/Camou
dXkx0zMxrPnXKqBkh4/jpan2+Qwfpg4x8erumH0g0AA2mh+bmjVfYcLNOJc3
pJtn+Rd4Xc5qM4ARaXHvbe7WU8w5FJI3hTfhYxZzmk5VZMAT/UZCg6OgNd/x
BhOETBgmDhOLsjIBa8vajFyFlyY5D8U/imIXQIvD07Xyiet/BQIfAO/Jz1Tn
Nl96FlxUrPjVfs4EbAPDxmMKds4yp0cdSbqdX8VSbIV14gk3AsC7keog7abc
Fl15P/PlkM3Ajar+tF+a0Jy6d8VXCvLtl+1GxoJepYtWEV/UniDCU0xPutkQ
+/Xg9krJdEvVCMBii5UBsJ3GDH25Iv2S9ceC2BW7hFzhXXh7/uMchu3brgeF
Bs29gicibI4iqGCKIW4YythaoWEWJ1rzGPhkrxq+NE+GSYQKeNrCtT11LaUD
GNza3WKLmYmgMNe8vbJLcMPtLNL6fNUNIpYfYKGwCeWJu/c2rPTRB/tVX1Zv
ZJ7U3Q/7qyP9b6yLGHmhcG8XRlrLpTeI4p1kPiIqwCaN2wqIefzldNyFFa6p
DKzEXDDj853SY7Q+fK2Vsl314bymhquNdDOltmHXli4aFU7FkZbi+8IpFDRU
5nQrxfwy9xpDs2LQwCcRzh0WYrNy/WDnTlBGx3euea5tx5zdvVRFLebmhjD7
Zf80tYxK4KW3mc9fC1fCGod3brltpRt6szYXzMjLjR7MlL8huCVtGRFpsHyu
Cl8iEhnrQRsqpM+LlfSTby3SayX3ATFvSDjiFp0uBhwGSF6rjm6o5bztwPfh
5nTBS76YWTNgpOFraC4b/dU5Jzn9IET7RIsqNdfuk4WAWWDUG2AISctBLuiL
ZYeiIdytWhyw06PR4H68yqXCQg7mAK6R9EC24v8xEglH1H1PDEkdJboMCboy
Kbo5gz07N98iPvEnrZV2E6hqYT9mzqMHeYrXybr/NhlYWJ4heStvgSJYnw4e
aEwtUaR8kRvaPIFx2LlisV2B29+PYg4BYOm0yXoaUQlBYV2HAo/F296+kPxL
i89mIOGpOiBYQt1hp5tsdaUszazyiZLyrETdknWGUaek0kJIKerq286cKLBH
fu5u1w3l/Q6PiZTRBSBhpKhmH/k/nBys2D3GaUpuEB4QB//xipfG6YU6M5jq
d39SfVSuxzqmxxLYe2omOBTxYfyfjGm8n6Ve0SaDJ4txEgavSfUCtDOhEGX5
dboDJ+GtQoZC+diyQrlTEZb5BBIe5lIniBjs6i4Gb/TQbiGg0lV6CVhZMU5j
LQOCMt3Juw32ZSe+lH2JtoMX7pKLAGycKjcQTQBIxS0+57Ozktmx+O1VoJcc
FZQVIp5asbiiDxar8zqoqEidFLLMzLTXIlAnSUclTcMkPO+4KoaT1ttl9yYH
kMgDxpFQVBXJk35xOawH6yF9s8t14UCdGaT7PCJG1VcEbpfXXydmvyPhs8PL
XQSwdSEJecip3KcP1tu/dGFrQgrCuValpW2v0wVdsl3tKWjFaV2oB2FHP25k
REtfl8Bo0SrVDhr+WAGvqCVEZlfMYMbkYnha/yxfw9/nKEbrUG3PUtTWmFeN
wXY/ZTDQCd60SIyOp+AC4jpKCqjaydXxCBM5DE7KNsumb+x1t/IkDZoM2JSg
HoNx/DHoVxBVSo9Jf3PwKgywKFZ1bnqH0Pz8J++7r3D52WivdYls9pq4zA+X
iQCIa4i/UK8TwDGZVKJDVhKdWa/w4VfW1bR6BP1BfkKobokQLOy2mNuJlgRG
HCtrcTgzr2x6gykV7Gse2VvjpI1s2i6mctOglzdlIkp3GfI/Ygn92NNgvix3
F9QMHiTjxUYAfNwliDk47D7Mf6A6hlQXe2g5oIqBkquoCVdDM6GQPPoZOEDI
ztoW/kIp35xUfINdwokqRMcfq6LWUBygihBhr5nLVSexopfq5E7J4BmozNlt
XNNwwL9wWT6GuSPWuaIiKqFGcaiV8xHEFo1vVMwa7SeNpgetJs597crg+hl0
Qe/lzgzbobaUtkOmV7LbA6Z31p+xOtz/y0eVhxXSfoIZ+mV8dqi3i2AZIQ5U
MSpbHbwhTb32BWcfvPLNitGIc4aqu0fgxEek1rYXspO090LsQN005IEmwVKf
qJIx+IKXp4Lvz00K0Zaw38kHFYB2ntKRnsKGzx9Fsj9r7LCW5XBCraQlKMuJ
lvpqMR9rmtxwiKA3yEYyJ94ACVUFHLLNeeOml3NQCJ0htmeEpojnn8lvioF8
zhK5QV31dVj0MJF5NFoS5COltU9qLaIzbMaeiBMsl5YvvKnLD2NfG9OOV4h6
o6WT6onb+831/t83nSTNeirFocXQ4r54peyc8ti9t1Tw6JvZ0mNWh3H2KzZn
ffEXRIcJk5+FCpxNfbhoWqzRIXGjaVNwqyyfQZEwum7MsrEemQsShnrmQU94
Z/gexmchlpkAY5byGGTfLD/Dfyk2JKI3e7Wxwhld8LC5s75MRHVgqLg5bHER
zvniM0YKnplUcoWStFXaW5OJyagPAz1X2Hk8UC8friRCCWjEJNBGGqTQLuUI
4mPW0dGPfZ3wwFTE+BZuqLphOFqyJC54QsXDfMxvXk9ViAm3eneeKXoZHvNX
/nZwxxfQ5q587KQnuKF3jORS1ZIFRQjPodYUyjwXs+OFYix4GS/oi8j+y1rE
mXJYtfIBB1nFtJ04R05mMm7yiosJCbU1zYKo6ZJl9qgoyR+bRVvi8I7Z4D2g
NtvdzAZzx27n7rJVSj3zx17J7kCfeCl0hW2yk0EvaBxSpIFETgBrO7mQeLk4
W4draw19ve/jjTUhi5I93aFjOoKKw6D9hfhw4sH9Ev4ohVvuo9T/mSx9aEtm
iLkWxP58dlTxN+boCAFL13Bv/iTkfQoVdgAEukpVQFnHNKN/ChVluyW99q4+
9eNT7G7KH5nHSEsGPqzuij9TQG6ZK3AszWcchfmWbz/9HxpB0WlT45VjQ0Oh
MjwSo/6Wl0YJQ0j/CbDUXVIECVTgoxwqNFJD9D42fTyifKoVNL5CcvFiOq70
IgMficNR4f9GnOgpwcns5afEuZj31EkR1p3T2xkuEfpMC+a6GChSKFNC5j/d
KrgYAALlya04AvSvbt+uM4nMno06wVuifP0uJdupbuajR2TTCBT5HMRTfNgi
Pi5+QUYQDTZMo+TLGn8DWQ3p1KxlH5vbY1A/lR8njiVtY6Rbrzp/aaPxcbJ/
aZvNUs204t8ApJv/VZSqZpAt+cd7WtkF8tBhJDpB7iSUR0VvkrolIgOFI8/T
+0xoqpYRnNrQQCtW64zcluhSBDhK8thjVyQTx9sRpR9bIHqF0a6oRqgxEIlE
PFTYkwpeLJ+PDLPBUQsQmiLpRtEpJN1S/GgjpNf4jvZQJOvmO/1ezAeOvSe1
N3mO4/EPGAD2GlvfBVr5BWeH7GYqjjJ9mzHtaQlNz4+HVZs5fYwplz6jx2VC
zkiejVLooGCZs19FIY3ZF7MDIAQ5pG+dTcTYNnM2HvP3FpWxr657R4NJaGPD
WoHFLqSIRQOUioul62rSEmAn9iOoEMR+T4XnkkR2fTJuOG7LHRSJ06gYNCdH
zqxUOl/XLDmRH80qsRe44G10WLVVTM7rkMIzqY8GUWCiajOS+N3dSEi7qB4f
i5qmuWTpXSGnjdHxBu5iXLcoxtMXUUt58WG9PdfWp/DOsZ/YOU39F/cdFGPh
zyvWl4Atc0Opp0ji15+rPDawvsbnOyAYmTBuWTkRa36Lb1nBAQLonDNFy37V
cm0e+CFsabnUzvM6c+nTDmMsKbc+RdFN3kX0CPR/TcsB62K8PqVg8iO8HLYW
I4ivFVj9sDZU0HthvoaM5ds7yMV4SDrIToEO8yJy66zS68wmFdD9UBXO5YZ9
8xzw3UdccenL+KFYhbFLEe73oqSLj9mTwblDYY30l/SxsnxAkxFISD5bRj/p
Zt+vDxRL27oyJgeJ9FbJ7uW81QfAG0j0pqTlg/w7a1CkDDNhi0wsdZXtTvQ9
o8WuQuFPM2v8OZN0ivg88vi79CwXIlzO22yoC60A3bG7SkcXHAzO3b6AMTUP
ykXZc38PQByraS16x7iYf4f5P/nxm/Nv2mdOhHy8l44HF6SwVQmJJozE/IDj
lCeL86zZbSNJpXTDBogMf5UqkaL0DvzMzoIkekmfyYrVO65SLNCwct1I8M+v
v5rK/oozAHtfnjuH7oDmQj2Tbque8zQbvULSDcVGc/n+dsXXQO/rqwsjLFTt
OqDecxRTbRfaRlwXm7flQe8msdNxtmAl5e+8TjSXH/yBcmMrT5YxI+LHdtVz
VtBRIzQ94rQkXNzdrXa5ktDc/1QReMq6xSRL0zLMTDeqdCEnaGEuYf7LlT9e
ze3+TD9a7rTnAowdUuvqUKrjtNRUiC4d2sJ++kn5Q2LiIKEJdYBleAnkyKFc
BsYqZyaubLxFyos6B7JNZh6YcY/YCXDD5evfbOAPolvbLcSPbdqlvPACfoWb
KBCyYdejkFrOOz0PiUSwELnoKyCIV3SGx0QRS8jZIBhwDOmIA29rN3Std1vW
YEfl117gENAHNRg9SOYGTNQhVPJqgvQ+YzckCfrZviExc7NASQ+gSYtFj2RX
OYb7tHtEn+DaHmuIMDXQ7f1pLWvqEXWO0brvqTiaEdB+NheEOz4QhLwLCVC8
e4hB5SVGATxNxf3f9uT2dPuynjJhzbnYXN3wMeKJpB/0IuWGMAhD9yzkQWZa
zpLsYyb946ZfulZg6XnNuBRQQCFcQKYfaBorrRqBg3HwtSCpKvfbxHQJIvyC
B02t1hJT1PoWUxaNXFRhubRhTUFzOpxz9eAEZOVwGr9kfVZpqPmKRj+3Rnvf
9D1nQAw59Gqm7QKRsQasSYeGPWaIFlKoKwjjzMdBGf8IiRjCiM1Mi+NArwev
kLNAZ/1ml/QivL6gPip2tyQ3MNW/JwMYoZ4WgtndNaWPHB6ETUHLCNKfduhx
TQ/j4ZkNdwMVkiA+C6q+XCYobbDF3UOwxiEHKlaLusd78gCZTv1J3JH0g6yc
u0LeEhTOeEjD9yRIHnC5tcuopvgaCPaXOUHPPzGlIKV+nly2iG++Q6FpO44R
d9bV8J/mE65YWhqMvAt1XykK0p6RTDMgDmUWztwMqGUy6W46Iq+i7+YbR6BW
/bXeXfv+U66Eh5JyraIlvt4FXNBsnWNeGND+8TV/3ln2AGNFQ+Ma6dTjFAM2
g3W9Ci5PcCmx7zCp0AZYL2Bgm/GaDrIAYaXIaIsOjcmxiC4fuhugP6251Fev
DtVllK8F0bcxMmcaczSWaThgW/NGnPOq9++sxkN6XL5BwEQ9hcmP3by/fEsA
Mg8q3Nsc5EsRwtUVEsUYiWZz8Pfin2cTWJE3BkQvwTiVTpKblIwDQY8tqncK
JfahtSeJaz32xkBzXoFRE1hO3N7JHD1Izc5MJqy6rbEWcyWctnVK7LSEobYX
Oq4NFYwg4AtUYPnzhNVLL0QskahUyIyrRatsQh5RLNkENk6WuUTPuA1J69/3
0LMrZlQdDQRZV3yqlz4bi2R87u0qvxolMIO61FU678fNCLVeBDkMdW0dP0Ru
+zh4+J5ZDq/M9ionQR84dmhM2L484xTHtMS+bG8jyPZAda+PClvDou5uxovd
YUWURwqHa7om6xPCQCDtHsK//KQCVnOxAeyR2n0MBm+8ehMr36xGT1XVMaY8
Z+kO6iS3hS3XqcTikrtVgS4T0vrVlLWV6ZkkJMCWMTwAzDTx9OYVCS13gCS/
9xeGeIpq6whkEa5Ms5EeShGTQeA8wZjPUNHYpThtgqrm1JgD02R/H60bSDRd
ngL83ZamJTz37kPU5utIrj+eHN+4qk9mzkQyfogzzwIah77zsa+FJGieFe/F
k16/pyr/Ve3bss7kMbs3HQRdBI1cwTQIetHkisGYzRLrQqTEe16ihJ69ALom
+J5JwLG2HsLeZcsSe2Lo2S8xcjzvSfj67juLM4Xbhfus9uqvdz1lXp8TDdb0
OmrB9AmEyjEbOnnAyTWcsNLU5MB4W7xZtTSMDbRFsCaaCaOAB0bsistukIYg
imyWkifVQsfTBwFIoCoA/LbjcjXEfxuaB5e/K4FQSUXLTI9XsoNkepchwtxP
F/f+xzEGMq+LM3GMUg9t6VTBNhyK0soDNuN6gFaaTGe3I1ZA7Jjg+5XDub2C
WXbXxH3bZ5FwPUgIo7z/ItUcD7EIjhJYsv5fHMIprqwVYtuy2cqjJgqcGHio
DcvUwkOxLQ/NqG3q2/CKBn3w3o2TWhP7PjdiO9c8qu//1N5NbDXNScsyh3z4
iF5Jjw3noB63fSy7QRdz1UrdBHKPFOOo1Z030qwIYqAdJ1Hc/bpZnPKtGUJC
YQR2SYae8fKwkXFpta1iIGE2JjgkocZKjtMpwL6SjJel13s+Z6ZQZpV7UK/N
GDylUmkX0cKy+lAlVaQSsBHgv2Sk/h2RNsG/LWoj4I3mqvbL+Cjbzoqpa5wl
uobkrGZgpQBCyrRKDz/Uy9B9tn+lPxBDbj96NbtoJQgndVjGzfobuQVmzrmo
Q3vlRvCvHMGjU0nZO09rv1dO/wmc9pMVP7n7oRmLTkX2Lpya/n7mxjBlnryM
xKHBfWTHauWh8kmJaZXRgRHdT8Ntvd6k0Mzl64ckraNqYF2PAABPUbTMZ4QW
xf2SdJ/G1/vQp/MpXj1hYWgwLY623WFh/P0p60nGhInhc/2OMoG9sMTW7fbA
JpyS3JN4l8XQlWrHjBe8IJfM+P1qr1shGBBamnNsTOsmyyBRopXcZLh4ssv9
TF+ZNiGq0C/LnYJVEp61K4uvuGzPA6qYG4E+goPmelouOaX3JqpVovgtN9M8
wYM9C5EA5kFkE7gmxdtdEeCXiiNz1hgnetF4Aev0UiSjfjOJa2IGWBFSyrFn
+OxENXQIhf9M+iM1dN4qEFTCPkrk4nLxE9RS4Ade44TXcRreYm1V/Gg0+dp4
ti6a8RdgwxQhF/Fm00g3WcMdtavYqh8MouxzETwcCUMWKzu+1T/rd9+kDYxF
gg+DvX3Ax1PfgkZ0dYxUxazQ9xVw15RjpJWTX1PyAhv0LB1tyRlGOTisXTsJ
2L9iOdbBsTCt8iSCf8JQAlvwV6uOQ3IiaCaGs+eop3zuVKC4rv1UGRiZu7G5
+zTY/WeNi31LYALJoDYXCgqnV8m1wM8Tel8mTWc1cpdHX/ytRkE+5qY455Yf
Zai1hb7L4zzY5F8570bQKgp/PYIttSo4oqBUUAoRIpmMjgCSGHbQsH3m8zNV
zv0HFI4ntA5tSIAeyEEaBWMewjjXusJIct+viTYZ8npt04BGTxL0lWy2wyyw
kllPOJA5ofOwTyY2MApQlRf3MAuh0iYXLsGEMXGKV1/lyZ/QXyV6tc6MTxUb
NWdsSUe/jKuJw+Memnih+hNR2FywXULuLzwueh6aht0b+QCXrn/z0+nLI9pK
RD3vqpVvQx0ibZDT3BeLwTD2vEUQZagbZD9VSVaTTxKZaERxdVwzNLQh92+f
9iURjQhHCXSDUH628HWiaZBvxrNNreR5PYOX+tmI50PegWSgHDrxUz/qQikI
TSpOkf7HugdDnarqj1/fX4VW0NCUuEPvRbqOMM12sKG+jaZJasv2zH07IsP0
y7G5Oj5lfcYVui7s1XONIlpX1vFIa/EPnIABt4lB/cljWGvO+aJZBWYVx8Ic
LRO1tQF8F8+13kqOCvfIpv9x5LGUXhS0cbvFoa+AoreVnzhdRB9CPs5TbIZe
8pBnQZfdBtp1U3yp3+QOSIwrQ85Se2kcFt2LKgUXxRf9PQbH/KiL+n2KnXuf
I/4lyGQYplEPgdr8ltGJMHg1evx+VVhz84S10vp79CE7/EyytQdJCrng3rV0
JZgFhZRfJbJR+2ceFH1BTCc1F0w21QmLs9XPJVz71K8NB9/AVF5ccL/MSYMW
aXr3Z5uTmVVUFrHg3/GTFntdZ/TuDPpaGG2Z4+ZLWwMuQRWXI5K/1gROxy68
R639N3QtYoZz/FTztyzhiig1/+ed1CRt8/BoOCekPtwSrk/M7uzmv2ozDBn7
eBf7H0bMUg9iqt1DIF0uP5MyaTltoEGU047P4NzZLiSZFRNHPBlPWZ85TDaO
SmW2M9A5KSDRjX0rvziktrbPcsb+B+CGMSer/1M/DYWtpL1hwKKinP6tq7P/
wRekIFKodQ0kXsObk7WyONknXZNrIIDQJ5K9bx4QBJIE53zBhWglS4qUNbRX
byV0zdijcN3n1eHWRh833hBvMl91nPZb5B4z4iHB7BpmaYaClipj0DzYxNH8
Yv4k2VVtxR45OnpLFHRsfAX3nMWKcx0CkGGavZbNExJdIwXSqjpiF+YpPGUu
ymUq3T1mhVKYvKa0ods4DgTrCqzl4ulEI9tCOI+CMoz5qmTjASFnERkxS4I8
IGxl2f1+licrkwm/UeQSQIyJYTYZrMCC8Qcmu8GeSjzvB+3rmYJFaq20/V4o
HkH1ZtaIlQUGZmQlskEY+k79B7u66r4m38v3faVhBbgaAdsBUTVLofgW3yRd
QK7PeIIBdETjp90mJOZ1MXSXH/Vdwd8TgVQaPBNWy2jmh0buJjDFGKsovFfW
eAtmZwHvCPaopBh3smXlID+Fg6P3WbNzVSeCLKqryZS5oKuW43WufWujNmjq
gSYei7lKcsvA/+gR0MvuPUEPW2/qf6D5yIYl7lXw1rqbOBih6vpf+8JDOdjn
Zvd7V10NSJ5gpEwYpo/yyloxSTMzfQmCKwkVvRwprI4WTczShti+8LM6Hvu2
hJXOvOJVn1OwOEGaaN08WgpA5Qlvm1krH7qEXhH2L9DUKcmGQsgeXMAH0BdZ
sSb6DGGuf6ydpececjVKFnwoqZeJDQ/iNOFFCw/D5TqIeY3uN35jBNRk+ZR/
5ERaf+ZwuHTwsMEwDUYTjYyxRexVxBJN3By6T/0vmZ3DGlanlMP1SCJ8xf2J
U0BEkJWL02C0urn43b/mBWmql7IJSA/01EJNUBrGbbi0O/0+g7xeHFCEitbI
k0Nxj10k3R4KxGHmGkrCawU+dbZa5yPw2g1GwFO7BLVJpFHZ/JJIt2z/XMyf
7TVJPoVMORUBIegSfu8g2oNVV/q4dPs5g6xsj09e35gWwVzU6ENnnTk2pmUY
mQBDBHWj6il6PpsF/R2MOYESOGM3n2BwzfqRXGundBscwhgM6ifqmgGkI6/y
P85hlMZ1gljb7P0+xPOa7mmb6ug5E/zCTROCo3XXM+hksnCNfakqOEzztWE+
aWbCA2gtS5sUYngveuI3CqjSLOneeKnZcXXxL8l/ZQ7afNNXe7h+O6iPx16P
kvun6UUH8nom5UoFpEk9qa85F47PUbzLwZI3wu5bsMtiI918PlEtGP1FM4KD
yg/myLJ7m25RX+77jGGFIesPLu7SN9S/bOhFjUFNS10W93yYmgA1GC5BtGZj
uWUYxYraiychLJt0Is7CYsO3Oer/KizSdK62yF3pqPpiLZIm/swiKPdnzgwC
ZZq38nYWXHAH8sAur/m7ELh/N+ztFejM2br7V+uO0aGZMoFkqgjmWObIm6YN
EIYWOTSpOjXTLeTNJ7/mjTVLueTV4vlLcvsV0jylxlOl/Y2OQFRzQe/04d1c
+PxrxYzVWTcdn6ewE71hso2Y6hIENF4KJmM1rHxEgvpdLkr+kSRq6b72i69a
XJQTcvLdR2t4lqiMpEn2Dp06bn/QqJsvnE3JnQfaCzkOrcAaVPdpM3DwFkWX
ZhOaaHy/UjS++/1bn5hNtrOkfCTLDHRo+1lhMBy8LqeEqKsGuQ2+V60O1QCR
wDnH5LftihJRL3bQWG2DPrb5+W0OqJckBsAvqgMxBUuaM9NSrWCm/8LMZEVJ
RFfM5amrNdrAH7wSBRcxESwwjX4lnC7iQo4a47e0bhQLbIk638Gq+oRbMxLN
Mb3DWgEi0XEb2pYd0c/gZPkCVY0aSi81Z/gP/El5ezNJUnQ7RBiyNwl3um5A
CSdnRhLfLgjFAnXD1p+9Snrnwks67Lr3oJqgTH4kbq/rUl4NYHeqFyX1aBhF
zUdLmj0KXjwdu6fKZh8wyM9dOH8XP+XGbdGgJFLv1wtdtIneLiMDl1pYm6kW
klmo34SORSQWXRTlqdT0ATwbwU3rgtjiRvOPSKHqWn5Ji4ROrYGVtDsahiqR
ew2XuNP5shVPH3jFIbxez1fo0RX1pD2ULuZgejzUVM3YF6BFQWyMWR0mNpBD
08DKZyj0y/cUWNQE5LzeXQx2tuY2POxWDdMMAkKLBm5zbt+hAiwuJqt/iUbp
7e+rMjhn1pbx3HX3XWIUXhYyLgH43H5h+FORcNwoV/BnzRxMaJCThwIWfMoj
vNGR26hvgb6cwx4idGZ0OUVPIu0A0Ucrm7QrtCQjmA/Ux4mYd2kv9MGTzGsO
Bm0BaSYe4mJAZRG2KkO0wVQ3YLhzc1lOOoSNRZK9Ll8YBItO6OPlWIMNoLAo
3RFORYSc9AHHRc1YuPrNxjGwPPHMKfV+4ZaLCCoiWzD/xpekvKjHzEJy+1Zw
ZJ+7K6EVFK56mkd+vxeWYqmojR+BvrpJiLZODYKUPz+NlXNd/bk0H7HlX9pb
uPxwIeyKBVLdJcoXfAvB5jascG9xq00Mpfwq9mWptMpQDCwNIqH3BcdY/QFS
+Q++l/baMn8tIYLWQ6XCN8/JI9IJAp/+fK7PsQCXW9ZfKq59e8XC1O9ALi8t
geo0CD+jTFxK+bBTvvG/TiUlBFDSQMqZhxbE9FS2nnw3yDTzfjAk2aMUDPK2
PHKQjtVlpc452yFe5V5APDEzY25y496IuX+ZnawkQYj7sios7bCgB3jiA9PF
s354maZ4wdGIUeksPG+kpMQm2dfvhNeYprmvKuzt05T+ilIb4wOql/wg1vL0
Oy6TD76qyk1u9XgFhkH89k36H3JHtZsrtt/ff9NpHNzo1i2ajVPODZ4mH7W8
iMD074DD7JdX+aRQ0jUiMHdRaV5WMJcx9ZRur53qrle7DjxHRxQ8MPcUL32O
QNd25sh/izjH06cZPdhs6LTC4szde/pEIGfZWmt42soCmJOYA0VwQcUnsNz6
qQhwi5zqZlN/upFvu8+o0/b9FxWttjzhKDtO2mHQMOYRYzWHlk+/Arlilxzd
6wsuMwMkfZhFp8u7rNznRv/u03NJhJOxCG7CTPpgpxv0Gy7m0CX16eLqphmU
TZHLpCApNjifQbPgOhj8ezd1t/fIoDOjSBV3q2ueY4wqPW86Tp0z3g73wkIS
0o9zZTlL9d8DaSDLcKBbKirosW9x6hZCHDve4Iw6+NAqDvxou6Hh9H7RShBS
NcLoEYkqa5SskYqbgTQ+8KMR2f77Dxn/kzY3DpVICC8wHeQH1kK3DhBPUKm4
wnipZpbOcvkayu8dKi4haLXFZEHxf74H9+YaDT0WE9qSQH07R/dEFKDUC8aN
EWwasDJBtN/KM8+lmN+Fmu2yh0LCbTvMJx5i3XYll9vCHBIUcR1270r6S5cv
D4p+F5nXtxqvXky8fqpbEHbDxwvf64K4ilqzMf7xnbw+7vJsCTa/+MG50pH+
cs56nQ0OXR5tI3YDqw+FdEp/moseZaPyx6UUrwb996RrD3NEDZXDDc6BkF4B
0eGluQPE6nXl6U0ysBpy/i1tene1olkg3EulHBMCLBd+941wOROkBgD6HeRi
+CztyQh4QjU3uUBR7ua3o6FNAZTZI+rgLsXXRIQz6OLqq8I7AleP4fmn5BuF
TZMKm8zSbpwyu7wCEay7/xSDOaBktEDQk7mx1BjdUL9GpxBisldB7FA2KaE5
VeIyr7aiJUbyJEUq18VBHpP3cUL7jIfGiWXu8YdsRc69FQrIL1V/2CStcOQD
JbRmZCP3U3WM/WfQzsSd8sv8cY9OHQI8z9LACnVVcsvThitk8j+WWP2u3437
wILMfV5gDN+jhQHXCyAv2i554U7ww/1UCMrDXZ36zUz/1ewYm9RABgNKJvLU
YVW6gfwcAKBeUyTaWLSQcqkfoeudnagq3qHcQ2AMFHqWlZP4fHH93zIkE9wC
vnrpAIrptodHTJNDXpvNXOjtZaom+CgSpWCA+vPmFQScj74pvhKPO6GDcUMT
3mESzXWZZ92b3zIRJCQamVkfeNdu7JbpXUWst3br422ZQxJtwf5NBvNmELlW
ZstJnYOFhoQOmwFiZX659AJNKg9WWKVLwIbVJZtwtgQZ895nNccVkWmVdZZI
4rTeEdy3v0Q9qAaIfXrPmWAsCRgKuiPq+ttQmoR5OIfENx8B0O3xJX/KPB2c
n1uEiCNlHqQjR5/Vl8fE2w5wZEPNFANfoRFnFfyn0z0sH8ng7p4Ngt4JYRLn
moSSvjmqVRSzsqQAYlfUIPI4nu/5TlYmHb0RHuFajbEnM/L4Dv7ALKm6ZEOT
XG2CirN0uuXy9gsVEpEkygVZJB5g0jqADy4H7T7YqgZ8Woe+f27HUJVmqQvO
ulatqb8VJ5Zwg9Vk/OHrxSSbsgO/YHRPMovJqDH85b960grQ8MOPi7I9KkSf
Zq4sfti6SIR7F6OJH+nkFwAvowsz2itGqQ3bQVMfEzQpRiuGpOtEfwyJLU6+
ote8DXsBKpww6ozRN5SPn+Exd4AsiUZlxgNqinLRaaDgh6u6wvYJFQgzsfUQ
8UsRXwwmvTwl/wySKmsNPjnaMZYSN5ZnVJuSS3S+UnC41g6tMBd5QLViiweT
YZkN43evg030aeNbm1uS+sBbiR9Ch95FhwiEI0Vk1bfB0SQk07ySFgam1bWs
gk/VH6lIK4xFVuGxYSV395nRq5rVzHhyfb0YHNG4uAcRBZqcHpLjw+zXqFTW
a1X+PDM9I8FLfGfJWKd4+i7Dwu4EJTDNKHD+0K+dG2hITHkJb0y8xUyVOyZW
wYNI1CJgH58uoC9fg8GmLTKq+eJ6G0Q+khI4fM52ogxrl8TAifhArDRQziwp
fbLVLmd6js6NsCqNNuwGn5wrID4C4RrlGbp95HsgFM0E48WEsAiA01JwJdDu
LlgYPaYPaVYK4pSIhRT4HYa4+gIM4UghU3TP/WAni9okcyeDeTpkr1w9usll
ylJx+h9AxCiH1x3m3tIiXE4CVh4IcU3TB2ADJ+NuEd2ZHWEDngzQkKxhE8gp
wLqGrov0JBG9j9LVDzRmgUpppIIVcN2QuNiVDA7lxxKiWQ+lRQlfoS1bo5OF
4C84PfVOjDaTGxdPj051DPd9E0rZUljI+oLw9JNMale1Ysoc0IWS5r6o7KPK
V/CjNoM7lIiwPEfkIWWKxMZnMiXeTskz45LSO3//jXIlH555L5QF3+cGgn+s
dz4eqZKVLVn4mnV8cvFljPCEiSCUWPsRnObedi/urgbqvMCnu/pXsDY6wFz5
MU4oOshaNEKopjWYgbLsuhpUsaKNLyGinIvitGfxBnj/mKhFD6EO4wdYN1fO
af7UK0h1ZSTN3GYuFAq3Aph/ny2kc3JWXzI5zaVlXA304oKcRatQse91EoO1
GapQ8LVunB7GseTTspDn6qcwe85ZxqUqvfTDPP/AVls/vh7fr5HxJ1ej8Euq
V9t3E3cn50Xg0yyqJcmBnWxK8Xr7FYiCEU4LLBdmwE4dYZa6KQRK3xSUnjFm
4RwotmI+E2domMRjBm0wU3WQuVmKAbbd4r8wguT1Ay46O9vPlFuEsYBG0EGq
0/g0ewSrLRWEcQUmI4TOXRmRkCJI6Wn1hdCyfXEYgoQw3a3mEk0xaqUlwlgK
nCvI3tNciBJtJIc6mxi19KKC/c3FOY/PZ9LZLwKIut/cZWBSpRCGuNXRXZkc
p0Ub7pX+127PIGmBqbS5vz5YomITk8GcleaIHlO+wHrVAfUnWWsRx+ItYqmo
3c5HoE0cXvVGZrXfq7ERhQYHrpXEYid7z5tnHGl1/i/wgGrf568FmfTrDzg4
oLQxIYRXYepzLpHUh5/yPoZxQOIOG+Vfo+XxVXm8EAUbr2xe6281Tc1BkR4I
evtpVHqahRMmfjIdqlssOM0rILs+AjRZyEqc3uzQIYN7CsH4ceDgzVoRQa9/
IkKrDYmXR6spTyzJULaj5WHRD8ar2OP6V0bwQM9KC6kPP3FlvJ4hcah+IYFF
fGDba7mnv+gsjLaHPuOV5FakRl+lYKvfg1RZVQ91KnpAvQpZP2tDyJ6rgrV3
oyx5JnoSc84Ul/UgQRqDmHBsQpIxHCh6PbbG59IJ+onmMvQKJdsqQhIDYXnr
nuGrUTzhR+O1NZ/GK7GLFW85jyWS8Om/e16K+srIaJYPkpVEby0223R9/W25
5qyf1kCUow4mNGvf0sj0h4OFvURHWZ+mb7H+TVxI2PPb/Ia0zF+9fRRg3c4Q
RQKnZvWxQl2tcytzFAQPWxj7kXGErvdUi6ZhAeWTaOIyLc/5ZXN1XTMyeMK0
JA7TltOnxPWiQrd6ElWvMZ9/4XE9rjTWylvWIPtU/ST5Qkm18sQemOifUFgF
4sNY+RZ9+kyj4hod1xKlh3aI/1A4Y7eYmSNHtQZt/4RWg1s4Wq2FAaJMYfzL
Ozv0QD2UGZC+mULFTX3CzWWsga8g0CbIHirlZDmMYMSbJI9Q2Foc1mjODcOS
XkOH/jStZ789tLl6A7D6yM/XvoFZuaAgFON4Hijy35JdcQaFgHCrpWm8VTzP
u1KfFujIUQkJj4eBGmiEtA+8QLY3hWp8KYD/Swca8c2RTZ5jSASAofegfFT3
XIPsV2ZRnkM8jOjPQrLLbOWpBInlzDr37n9m9CNBTZHgLk2pmjIJq5DjIC+O
OqK8ThPclo+wZgyfTwR8UMBsXWiQdzkfBxd4Lo67GKKb7fETSw0tUZZN4OF/
CXsD8QhiKrIVyK3TyBBhL9qpyyU/gJRpXLZAD0s6uw6A5KdxhigmbEj8Q/cj
/5dDMc4t0F1+xV1xJl+ENkQDoNPz6tmZtZaIJGifqR8dGPZFx2EbL91/ErhP
tccYMfF0HLEr9ZNO2dIxKusG9lId0Vcf+Riq9vo8LZ5Gt1MdDRsgBGl57UKH
QqJkdU6FM96aKfFvlq1FPXzyBi2m+HXKbZIlyxDSsij6rKxG8Q7d2S5tkNNX
qxhAukFs2oFl8kVqW4bycK5Cjr8a6ZJ9wbLtMmmkEqJos98+JEWwsit1Egvy
LchPw0gIUlRzyA9DVeyPB7CKde1ris9AGQLoeTWsl9s7aEJUl313nkrrg+u0
4W4w1JzefW7Kl5x3CwaytCVFnIFiP0gBLU4Rc7DTK6EeWObPDmh1x2gjpFz5
AKmgF5Epz3hIYse+k6DtzczRYdipc7JGoD1mwZg94eVbAS+nA1WMeQ9eNa2K
xfjYs/+KWM2ydsTLLpRai+VhOlXHopdaU4VUiXJS7v390sGSfx9Uc6pl4bcu
UwL+a1zv24FM51QEE1QdTmP8seh9SvKptoJEcLEQszfIQQcM/bTnAtrUoGX9
M4Cyy+PkRGpiydfyhsKlv2SlRPoihWKHjgWEwqJ1wreNEdKMgsHl6N5mysDv
LIcn9c71i8ow9i9JJGDhaK/JpDGv9g/8KWwHccMsCPmC3JUVcNSgdsQ/3Vmx
8CvhhvgjG21KKLWogYKuBcZ5/KC3EfHyVMPDjV+djn1xzUPPLRiU4dNojb+d
Hj+Rry0RZepdSfAn8ZSBCPv4QigEZjUQkOiW6hvdw7Wje9AiUIRb4nxPJB/J
B+LX+cUz5JrXuDcr94Pd4/HnYa3LW9qWYLdzMW+MaGYC64Ty0dy7sdW0ri19
u10WWuYefMrUcIfFXF2KSclZz28+XQKWg1QW2lii+kSGOOVkDG3yvpo11yXx
Qn11T0Q3U7zVw3ONKcyzRvHSA1vvubzDV0MtgrXudvbEp4fpuwf7zZpWoKRs
Z8aM9CWXwwboXbtwKNY6wbRiz7tiLKyJPFER+H89GuGE0UyJQ9JLu3NNXdJp
j7mKYSlVdN6WWjJcT0O4/WjfnWAZX26M9fcdYZW2u0MO0A1O5csmfOuWW6aa
nSoYkuSiyysnnl+A7VKzYJljTXnxejzSIED47/4u1Al2GQzM4zre6ssUxsD1
WEnzChV+mXhEROfxzHX1fpxCuIgx52mgmBGolV4bfim8qm7Idi0V5DQ6Rsk+
FVlc1DjFJ9S/J/zJOW3UxDZxGUGwp0QG4WXpLLd/WO7I4FvZqZ/iYFZNRx2F
TnL69lfT8+djs2Z8F9ho66OGslcftI0lOiwYxPTJdaJ82GihUfj6PrbgMRKR
OLaES4kX5mP5Yus0FIaKETNSd1bgIHLL2mOjhharDMJlpplDj0vPSK+k4hlB
Jy/PhFqHKbM+ixW/13BK41N7saMJtLKmYfYli4XM6ShlqD4llXKI4fI30pyg
+gnHgdv7F42zXEXvD8+bM4x/omaAfX2TAL5yi0vsSmYpKIzTkDfslrkDuIzv
sCAQxmlZfZ+i+UKjVTb+KZSHLvgJSDdPp0XNTI8LHNYd60NshdKrQSWAveGv
2XdlOkaxQ8IMWNEEXcHqW2PneiW1EhAlp1HjwUu0yVjSfjSvgEVS5Bj9O6+9
T7vkxWzmg1pz0bAzzI1w0QNGI/4kilgkWK82YYb4BQquTWrP37dGtyEcS4UR
FF/puW9eEcPh5to+eAWrtgpRpWb7M2isIPXt1GF2hkS4IC8fU+TQ9WWbG/U1
n9y0mFHs3GAQqgp20Aha2BKgiXeg5nzquBiABeNtpZrbOtMcUmFMeIhDouw7
tFPFvaot48Pr73J5N1txeY6uK1Z4dmmehw+NuIsdaFk/TSh4iBTcCLHpTSpL
tTA8HsjZ82/VdIEyQTGHaUWIxiGGYNvFufHk2H3xmW71Hq069LaJ/NBQAnk8
e0P7nbOHoI0ZcsPRo3Dn+sgs9rfALlNU+ClJW7r2Bx7DvKxxKFXyWConE7EH
aCfo6HxC8Ko//8ExdQvSVCshSqXlzSluL1KMcRvD4jSOG1AuL7rXv56oz1wI
GV2kDbSVc46y2zE1Q9aDv/Bg8fpz9c2SM7YbhnglKtJlEMkIsjbw0BND9OTt
2GaRcMfp3VD9JRvo2DeLLML4/pGl3nNJlx2aj6f3GdMe+hf4ZkItmpkIQsJ3
SXYsFq+HNv4tl7k133Mr9vhuL2F8QIn9/IDDshcYH1FJdPG//NlLYQN3J3Op
JuC9dhV7HIkou23VzGy3J8kvAvgZTEgz/HyAjnSkdy4PYQTx/mpueX7NvzfC
+9ct97HKqST39+cbiGPdS37CK3upO1Mw+nsx4C7Z1Nl0zxDMKWw67fhJHia/
ye0m0jjk/DKB5xCwXRPmcvpBJFIAEPYAyCDlK996W7fOjAwTdlSqAhhb+3dC
L59jbC8newbx+ZinhyJxauhiOnIq9i2+zkOGkTHh+H+hazFsQ+AJxSMc5ehx
NFulR39T4NXQ2skdvYr7P06xzyNIgm0J8TsSgKqiWpyDOeIs+5GQpnt0v5Ok
jb9BFIQaXoLsJAydMCNtosFkmokhCr2Hzl+8K6SvF6vRPGWRPZ3v/3lFFLQq
0/P2DvGMAOPXZSIxVXBl7ypnfzoDnWspBJLbZjAYNZbUPeZ5zP3h2Z++RG/I
5UWNYVnEHXMkFzb+u/rGJZJcwINdSS+R1ADbFWZ6uxqTO3dDuNwI5eR+ThT4
kYJZS6NeP2klL4rN3fCEo3v/7D6euAw5KNnlT7uZslRS6Nni4Gsrt28koN7m
uUUo71RNQL38PHOVzXjXUqeJI+DtQVgLMJiVn+uxScgF/o4SqQdWrJB+WJwi
P9la4ADORv+RSfe5FD+4XlvQSmu1kQL99AN69i/Qr9Pd0EWDPhoxprhWyiV9
DWZu7Ja7fr5+B1LdOauDaPSneTMj3kRAlspGsIDqFEHjF2VubxEeXIExCPNt
pdGGveHpaRPAGGqEOduTq4y92rjGyxqA+zmZGvSLTJHjmfZCtupgG1NlwvZo
NT0xTcDhg88l3//HN/EQndRPBhCWJ0CB3l9bkOPzyYMQ7p9aKULXA6SQqKm2
+xHCrParX7kxgpK2I7DFebYDr01oO4TbGNzcMBZXJLD8+mSdT6et5VYOt4wj
QDA0yI/mzLgLdo+cDCtA0n9kyArhFRdel+UKm1Cffm14fddV2hsVTkF2vCxg
gP2Oeh+lfN56cIb4uE3j+r0R9QuYNPTuvzQ9pAD1QT1gjbVwj/tlwYVNntPU
JkJVaI7sYiibdgCniLiv1z/JgUQFeiQFinjeymadyc/cnOfIHb9ZCVMTk8DC
/z0q1FFqUQJjZa0x+qpQ4QhZ/qpOkQuYuEKEK4/mNVh25O/AfPK76aCLB/uX
MXf0EJNDtbl4AXgR+80pgsoQVLrEUHrruw++JXpTFTk9Z+KX9WBXj3wqh6ev
gxeblKZPAJPKMo6ZGwS3jWK0gwDWjEUnr6PS2WuWak1O/a+Dy9qCFBCpt7+O
0ylqgI+Gn0zT1Gze+AX9xDyLoIx9tqn6JOjyOxWQ1kKPsurR997oS8Tp8rvu
gozinwB6adHogI6dDS8ggit3OXcXjeCRpSPNYPhu7+iWHnSSwfWh1loMX7LL
TJUpbEUYSPsUR1xUexhsbPpU3mVgUvj20E2H3qkEPwXGt2TEEUbr3KuoO1eC
GTgXU+4+Ffl6RV44KbFPkCefP85n44Nl3vni5QpkcraPIjMWJHYDL7sEautx
y7bQFpW4hbUjjEr+F+n0gGCA3nCEFQGTq52k+CAhZ11KS+xlUxQCh+jVAXUo
RrscH2j4A6iK1lZpUTaIH67n0NBRwSB1ezUxoUTOAn1fTtCbZHHOWpo8gAja
nPrGwDjSqbjJcQg8LXQbI5t38Xy0Sxae/bHu3j30jioMNK1sjVaxiDclz//e
Q38pu4JaB/ulYHQW6J86BJbGl+8N7sUeGOli9ippl/D4PNLm+ID6Vb8sR5FK
lK4GZhOHVAbDgt1CzHiY6q2Q10g5uxzxrETLPHBTTQjbLVQfCO9PAZGRGlmK
qbIQ5+U/VLrmV9EWFFmOWHVkg3Khsz+fV0n3iMRX3l64zfT0eSS8xnqDudwu
oGIiknl4GhSxwFzCU58EDEht3agiRO+QtI4jH4ciTjD50nKGQZ1uvsM8fKwP
0vxZRolFCJMzjKhR3CP14CywN0VytWoIE4qtoV/Bf59yTq1lun/pIuqHaq5m
/qgY/2xxyS1bgZfJ1fMM/+gvStXyJ4gKRpj2soyzTKHfRLzmNi5jMtyP4Xvu
//erjXJdNOffmsfX1KPAZhMUjtIZpJi3NjSClLXMqXup9QqEWWE/eef0Y91A
Z/f8g/ujNytvBVyvyIqq7P3Fk0UcrsPUyfX5FTcRxFzIg8WRt7359+GtOdQa
MlkFbPGCMrpKuzZuyxLiBkj9q4ssBeYsP4mksmI4cbjlm+BuktNYGew3dZv5
wVsRyxZL9iau/mavY5bRlcIE7gXW1FOc/VcZ6A/aadjCI8BRi3cuAMKExVxI
cO6XO9qWW/k1IeBWVNsyCIG70Rp+RoeMZizRkDFPeQ3SL6ukmkO2fLdo/13G
5862BlxOjLZaiiE0ErwcSIni10PeXBOcU51EdRDGgcPDiA0alpZtBLn0iFli
s3Oma0AAhX1Jkq49iGy77nKAGf4ro+HZO0yTKzqY+5zxcnbjlImId/bV99FG
61Imw2VTStbkeQVhJnBXrQDPUpiesAQ9lGLY5XGmqz/+eEkoFntiyNUCxJxP
n5ZzQM+CJsgpalfrjhUBfavYKU44rUrVnZSNe/eMqj3zYk9ZYt07wuXZn8aL
JzWLfwVOKf/SSQOUb9avUvWmcLT7KTeTuV1GS+4VUOA14c22hA4t3i/Cui1P
J2DXQ5y3Ha7FX0oiH3x/OV2J2k95ug4xKd/i2SbDJ5yOenImKnyV6KTvBW+j
b+QTG9kOIqf+2AB4VGxP1z6f6EMFciKtgECDaPJDwFEMPRibmEEAmydzlxyj
/s+p9Bu2M+Hg8i1Qv846ns1IMKaV8TTHI0Dc9IxEsLqAqR1FyO1kCb7Prnwg
0c/B5cfO4HkIEroiTCxZMi9jWcp9kRIY+R7YOO7w+w1jBWbD7lxZ0hheUz9N
9q1ZB149LKl92OdTo3pPbQAZ30p7jJO2Fh2abKhXdiY8w8rt2SR66FR8oFwI
v+RHCrJUxEi4kisgOEQUr83ANbnvseo4zqIJshx6OFhpWzJjVtP6n2XsosS6
zNFAtK3jgCcfrHqNnU514uv5qitutH0KFPqgHgAp7ilDMxumJBksSdvmqUUG
HwFA9fJIv97kHmJkfvYAy38RZiqwOPUmEh4Zx1ElV8509ZqyJ81S5UPplW/v
h8neV2bMv9ASZ5UNleyILnFTVXVR59W8Tp6W3KSvuxN74k2j2McexQc++I+Y
zuQA4HXO5tdrKtzExO5qcrVcz3jYGVKHIqMkmVeacrE9QkNJp2/bOF+9du+Y
Ul51ZLJlCelRiq0EIjQSB4JRpqNUQMOQUjfpHtuedPFUmBwqi8Awv57YkMBR
iaamRbNq22S0UNjmWrUS0BZgs4kJA54ZkUVEKsGU1VieQsk70uhaUw9aBsKJ
RVMXJ5TE8SukzuiOk5gu0IZoATajqDmE813XhlWn4GFiYFTNt6fqMPn9RTZz
afB0bH06IlV7S1DO4PvT4y5uYU3cRkFngd832TNDmF/R/VNnjQ7SaLA4mXxw
X9Z31+fhpfqshcgsLKaNnj67i7qIHf/A6YcKqboR3O751lT8c0WytIye0HYl
p2ZkhZKDzjEZtupSm2n29ioVx64ulmZRd1Zk7uXZFtKTwou4BOYPvcmrQ8lk
AGT+WL5srEGd4TUT8bSKQP7RARKl+hIfHa0SAcssXAQB7JMxig6a/Hcx8L+E
7PTvGf8UETXe1W8YMStf0QpBz36qJxSuUK9CEXm8XzJx/uiVV2i/8CfRqGcQ
0r0aW8qHYaYy9WArXfBZcTQPfGcLMVB/fotG3feutvtC/sD30F5Bw8pY+3FU
JKkVkEUFpFyuxjlDoq+iygi2YAdmxZsggznzFdMtqcweb+Dx6cPr//SLtseU
VjCS9l9TJWAskWhsuOcubfiWQoN/srnjizolsXpaRUcIId3pld/MxWjkN5uJ
7SO3oCTUJXh8Z2EC5R8WCVy+ZXOe+0uf+eMyJG7lOJb16H4tQ8q19fn+oZw3
SNHp2yL6t+X6s5A9OaPJF61lk3ynouVSQavufx61GwJ2DZdjDZTMnB89EvxP
yXhqpgPyNFMrKypZejYGibzM9YIx82v96orImPwzw9tSS2MIzS/IR7UfeJIR
AA73Cm0U7Yo4gUZDZ9OYc3rSc1qLaF5sDNMdEohkkPE8TKngWwSVsqLpyaoa
ZuxE2NgEgE3MO18G/kJKObDRoQaj2FbviJ7sDHf4oDnPbjh6BB2rqmgOb+g7
NrJXV0YmoisA7wsUfBGtnzDfVee2kzYNaMdN64VNXG7Ctaq4J9zdN6tV6GHr
QeTk4yBTAdjgxvSsKh9ds6z/RUMRNmHG8GARC4yrJwdaz9kMjvEpzV5tkcyu
lD+gssoNTOaajAJNGgzGyMtOU/bOyZFJ+nlLH8qsGCYIqvCUdbs5RPmIclnF
mFqZWUi30TBC6eFjpFP7HuQs282MpBVmwUY18Fr4jywe2M5tYbota0qioC70
gK2BQadfWQCIw389lbml7o9127S2mfZMmarMqItmO6EkbgmfsOLhZre0bF4G
7hBQVZxcYpBibprRNB2ThIRL7hrhXLX0L66/WtfJuk5855V3eMHdKyYqTCQy
8TktZD1QMVAyx+OeqVH9bw76pkUL0jxdhSgaLF0zAk1f9+T8N6DJnET1GRje
lw8pMJejbj30C8Dp6FRi9A8I+ZkQGaAyVnN0eiflGJ1Sng3cg/K4mRCjhaHO
t9+l1DRWuTiQ/sQo+l70fVaVGKAJCaYt5QSnIdpd1RU8geZd3N3nk71+9Lil
Afqi2dm1+9jp5De8I7Lesj/REoPRTQtasj0nQjc9YgmuyEHIRPzv7RGQ4rXp
SGqGlGNIf+p0pRtIm2kN66YU3HNustbW3iTztKbAXtpO9PWnMmiC8dMbHTpy
8hzt1T3nQa0O18/UW0qUIWalnfLTDdXZclMs7yAUeJsLxaOOUCfuXZBQDcti
xxtTp2KoYfR9IRMHIks/4gcPBeztVFU66PsgEfCnw7liXOBqcTqqrBaKSH1V
3zHJ/ytAuKXLXHkqG+hhli5N/HF6eZZygB708jZbMRldRJ11/onO+rRH6hnC
m7Iaq3rpsMYK34s5QXKR0HI+vfR3nEQkZGx9SfTDpdDgf2GXcZKbt0dawfWV
hVrVxdCYIKkK2yt+S2lyVlMNb/HQDO6W35T6MYs74r1o7uGHOlLzmiiDJ8/E
NfAyuaERm0QZsHb6DFN3pANFIYRPwjY8ljwpTZAnOPesYfO50oJd4/JK8iqy
OdNbYOJXFDv0hLr9Ze054o5gVFE6bxdDid6WPDrlBf2yUc+oIlZlFAstThNe
VsQeiK2GfxjfrVNZJDUPHOx2/lrAL65Y68ufhGpr7qsDB4zthpGWyP7x7W6Y
/4gOE0TEZNvWkmOF4eAXLzwRjDZDio9fMMEE9uOnEyFTxrLiDZwKhdFFsPLE
Y+4i/hckTFP+v6IgwlDGi+mu8Fqc8XCZd8R4SVVruHA3VIDOU07qBEPSW40/
WRGPbTq/pxd9OO+0QveNVi6+Y0fRn9XdYC5sBfif1FybRbpBTEDiygGFKlAs
r4VlaztJlVcf0c+xKVI8i7WnoPHVHPoPwha0QG324ZnzFrmb9uLSgUnpUwN7
WOw4YedMdF8rUVaKJWSNU6T9AAycWnjGmG7Zu6SSuqOVqdCqlqED2LPj5NZQ
PnSNNj9jKyKXgcMUFHHqp0DdR2Li7azrVQx1qmYNwtqUhCAKeRiMJxEepx8b
hhyQUiuGuVo5Vnqsk+lc38dKy5kV/CpiDIextlVTmxUBEmqVD60BfX5En/u3
i7RytV8PpqO31IO+ItZQY3Bdn1a8FAvBuJG3X65wvITxq95vMhjvhvEhhDLn
ZI2NgWQUDI7RhQbqImAHhrzcaLuWu3E7HjN+DkTLUQvLfjUNEuv7UCAMK6ze
kDZJ0M9GiuCv4Xk6A/wpiKcsHGcAI87xSiCFp6L/TG9HZeBndRciv+JrNYhM
G4OMSEliIJaqtK3MaeyKHqDKiGUM++OZKqlgVG6zsQWWFeb6XRG2CtqVxvt8
1oQAa/bBA8/R0ufh37Nt+9V1BsGqzC9hcGYV+iEoYZxdPdZBbm1p51Z6z1wZ
G7+aZMat0emOx7+ajPgNkGKUMz2M3pKz4CD164OnJcnbxWIva5tnLTUATbjs
MAC3ZkcA9WoQ6d95Epj0isG0GaC5YsE8QSmrGtHx4I5BcpnVTayP9r9NPpDW
Z9Ch2HAlluBT1mYNh2NvCG6sS4GmJ/4MAuv2a7vYo0DWReojEOhyoXHH3Kpa
/bTMbx91+lZdaB0UOkEQvqJbFv1UU+4YvcW7DizpDOFZKzxPaEOdV8/bFuCv
nXr99DDCK1iomSs0WedlNdyhcxrE7rCnUI4KX1CpJHjws43/3x4Ud6k2fLQJ
74FdAOzaItrnWWbFF2w/oxbQYEjHyYNb+lrB5LGHaWGtZcUCnGOobye5bu2o
JofZc1fhg601fSvlI6FB7F4BwOHvYJswQkaw5ovUaI9pwVbzt7sTm+1DwfPU
XsdT2iGdAZy2vuVWFPtSV+DOfaOPXwhPWD16VpSs55geLuzdFitYdRHSyqpO
xhQXgUrwoJQOGuR/5FE1HlMd8v9k4i16cx6l/gL54CVZLcjP5k4MyqV86sXw
Q3wsem1Q28Xpbm9swQu9qc2Pzs5YUq0+5ING+rDRPW+hvwv/jIDv2kZJW5hC
49LBytUslF6ecYe+w9QfhWskMOhwE+20kR5cXZb3j4LAGWBPjvjcf2bEPtu4
Wqe35MHc8WPMU8LxrWSnXi3umrpraynnRuC9dDud7RyLzVk276Cp+K02eeDc
G44/PxAvdqpUUMYios5g1SxNa2klJ+iZEp8g47UV/OhBhVjwmHG9gj4mlM7s
4H10A3I6z/6/YLKFNA4lbJpKkTvuWkRgSTlKe3b8XBrXJMsum9PnAWTGCdUg
6sygajJ9SekVYZpLV5h2E1ZOxb73VmpCJmSu1s/tJvJQuu3wreet+laCrqQt
UPAJxsK2WQ+2C/Bg+vTzIsAXD6FKVlamDftm/uD4qqhlQrYPeYLVT4iojuyB
hN7U4l79ct4VbTL8LS/rh67tX9QOYFB2XDDtrLa+wz5K402xTh8lDGZ0spMy
2O2zxBjaWlF0eO4tfvtczjEnxjwSY+l4VTNxB3UoANzJUbjmIhVSiQQQXnLY
EGAHPVnY96wVi23L2EoKh3xH+Dv3XION+HFKVJ7Rh+WbD8/sqQL3EyqEaR25
eRCu3x28QTX9epiq694zP1+RJ0pSzX8fY37N3JA7yObNUlK98Xy4fmY3rAs/
ucIbG2k6Gw1C0ooKVD6wX4vWLeGNKVkJZcVA0Y4oe1FtfdkTZH9allUaNyEh
sQSYWZgjQA5bl78Hq2s0iZta6EbbNFQXC2VAvYeSOnqWY9d6+fW/B/Qg7fqp
lJlaU/riMyoPeYWyd967oFXRTpiP15kYYrZurDM9B4uQUBxhoDQ/wgnW92pq
x/eiD33tKfvrr5kMIbrBTvRyPpCK7Rsqjz0B1j6gWP4MX0IFuNq8qvfKfdL4
ZREBdrioLfTR3Lgnc7rePbrx7U4hYUOwi+n/0AE8m2P0xyA3mkQ4f0+jRTIn
8dZCswU+IDzG/A15ArhOqQyC3wQaygk8PA/4pszlld4kTHrdX8477WJ8r4pD
yYxVxrJdQLlZwuJzkLIrCvrqwTPPrM0SGfXWpZAkKR/sUyf6SVqAQ0g1EmgS
2kQsG304hdsL55RrDPK7namZjRm/DotSJNepKCFpMJ4qzqjx6YDVdDfiBFw6
DNC1udfDsZqjBwnU7qO72MuDpjkdrQ2mrgy7krjmtqugsOBzC6/Km5lQwpZ2
fytrKlKQL6/LEL2hH86Ct/kxFsY5Y4J42iwE4kD4G8idf6hY+cYPM7Uw7z6g
V/+kBgBrekHMFuIYKKRJ17Flu4yqCK+Hn0dG1q8DVm8sHc0GYpE58OPJY7+d
xP19xMmnD+ClNm4NljP/gsHwzbv/9aTkJYCS2nGjNJuLvoH8KHwk5SooLNTx
iKvuirtGxhSaSr0kfFRgGvl3ncedfoqqnN6UCuu0sinacnZD/l9+dPapZfs2
UbwOQOjrpXI1AxpUPaWZyCZjngUlc9UY50rEbnVYcJYaGfNf5fige3cOi79b
086sMIv2Gb7T5WVeo4UrYrksBGkZnwDx7rDpNBBOvEEfzHDMV6em57pqxshZ
2YSti229oWW5Fne+oOstyUZ2+SQSaWGXyD5Hbt6wYvBpjH2iDSkO5Z7zE+oN
xgVRNqusk8z+JNtJyZtaov0ujcvsh8MjRh7WxjquA9R9+GSSY0lOYBemC5qP
TJ/py3wdrCrzCd/HGrgWrPGR5nOZVWkfjKrD5oqhnfPLNODVTbEpFnF2r0ta
fyVG6cP4a3S2aD6Pncb6DtuLfSYfEMyjrEtwUBtgcnMPO+IxTBRYVOt3OH7g
xJJG72kmzF33yjP0EhU1jUteAmxQk3EEOYF1lz8RU0NoofjDNTwP6oAKsiYV
azKd/HoEoJxfS9z28KSjFU3oYCezT9Dv3PN7flMamyXBuHQ8FGzkXxLXMKsH
Sk5RXLHtqSTt1uWASajmDTBCV/eGmhlb87ml9fnKaRDXggnFSbcEBSt+cK/+
eO6ElxgteZOgcbydNaXJ2up9dfrmDDO0Ii+HdPc3q4g125D5CEPDEGwo9yMb
6QhRmkRtuz5ohnsDuiTNE9MVvnJTml2OOOnocUd4BA82DaLLBJWxK2pvx9fG
O4AHvbpf1g1J/fS90xNpf7XG5XsxA3xqLsLMpnagfJjvpNZRpizAm94fXxCk
DxvfFDqyEzKZZvxN/4seqTQ55ANzuLls3ipykTS4Sq20tZsBuLv/0ZXQyiI9
i2jwCKWBqk+6mKH5gRArtwzGI/5IcNI/VF+PMTWu2oD0PNIn/FlsomHQFsTz
n7JCJea5dWfe/VyeZGp9Z6FGg+FZK1Qzt9aOcaJZ51Rw6tVqg8kH5Y2Fbux3
HGnizSAqPuAnm4s9Y37Uj2ld0nlGX6ciJcnoucg6NyVeM9+FziY9/0r1RcL7
tRnI3vkNli+UXLm6JJvSzmHEH31L78Dnq9o0dyEPXYxFJqTgpEBrSyjcfXiT
taj8SiPcHHzVVLAJI2R76bQNvo+yBuRibHE5SI1w5DdLA2NytRGa9JQ8qi9e
5cuhreAjx7b4N/x6kPbM/LHVboW7aR9zuQNTdJGKXKMTVE0dKCpixwkCZZP/
x5ZTVS866WuYE3xKIPhBv5k851WpWg5ITApRYDk/ub7PhPTP7zo80YuZ9r0s
oGjDPHicvHD0tMinRMiVySBdUirNMcE3pNTu0g+CCR1YtHNSAYlbenj9LAtk
xk/8Acqn98tKmKosT5zZJzdxiDgNnZxWYdtt80N17paIDRuBj+rn7jDb5LTn
R+e179tcorgk5J5Stn5yjbNRxQn2gT/oadbuOjS9A9gEYsXFSmnZrr2Gusej
L5izxgT4y7x+DL4FAPWhGuZH7uy+9l4hkUjL4cW8Qx9gBj13vqb8xbMFtA6Y
mwKJVDRul2Zasb6lIlgK+RAHp7o6TrbssBSW8dvLvGTBJnAZLN1esNuAjf0R
+DGxI+I3nk8ei5BBrffzgGSn2DlXhIE07EObBLHlmuR+wXy9TnsHA2PynnIb
pwneZ3y6Id2mFYUPH2HtaB2BWwYk5X4cIZlwU7RBP2j5K6FdxZVP3WSK87/V
Xa/6pwIl1nU7qPhFhRGkKBDBmIM+Ysd4pWVi7BGy9LzNtJ5ST7XEAbSLeqX9
kXi1+CvP/jsfKd9uOyblPpb39ZGwkvfhfMiCBO6B3Qxxef1BQvtI7NG0D9Sm
9U5RwPaxamRutPTS5AfEt1GJ+OINQek7xdndxY6h8ilU1PfmRF5VjwqyxsJT
x6Ceph7YAsljBOa+x1cLok9QySAp0w8VOEwIFB9MxsLaa7U7YwWN4iQDqNzE
THgU3tDSnHatWO62HXXAyAuVYgGjsXvfinE+epCZWqEhGYZq00buvKKIaM/5
8XMmj9djBqTljMjMCP4ki+aMtmHEJfNPNiQ681EiVd7ravXrhXvTdgGyS318
7L2sQC7GW41z/XjLroRVfXceb5VyAYGvqHqKbDiak7sHjKk8OfCafhqtBUbb
CV5U4pPmb2+gbEqQhM1IT1sIKSavqetX6C1Frf8XiBN8nfSTKKbqYAX9CvsE
LLQOkr9DzsR/UgIVjZaCe8Ktv8hPjBl5Q+AY1wbWP54QiXN0ifBGstHolDgN
O6v0CMQAkobvcwHTR9YCnShjDntMFYInaSEaEKeZSNOz7/KHlmC1s4lETZnT
eZ+W4hb19Cv6MRBIjnRIu/8Ey5tbFupR0zhjNhUIHUaCaG83Sz91hzZqKdkJ
ArKdq3IU1pmeVE35dW1pcm7dOPxQTlgHGLlgKeS3iV23XQlM1enF16WaEknf
N9XwBIFtg8BqI440Z6xyVqAE3mjeEOyBjMB5Q0KRRTim0g3NRCxJga9Pbtr0
t1MNF1DfBTTqy7sdecijkVbpogZlO3TqQdXM2LDm8LbYrDIbjBGXSH2WzKjS
z5IEIEYNp0qcrGYWDgQJ19jHKOtWRXx3X9viLexncRcIubtlOrr7Zs9p1NpO
65Xt8k5YtBJdFGPOVPPxdcIR8UUjP2keGepCtdQn3INewodIIoV2MfJNN3pU
O1Q6vytukoYAJnh8XhiZMe8B2DyMAhWXfjuT42ZnZSow8drX4T2uOaBSP9MD
CPAT8M3471uHm/bTRVNDsvcOgsa/iW6ghZk9WjhRJYfKZtkNk3svnVI3LWiH
fLvZlX+LjRud1QhX3C+lE2FbD32Hca7h0kEo0bb+nlqAmO4HfQEYRh2V2Mqd
lOoc2eNEcm6Ri0aveGTsIQoNjsGH37M0mmNJ8VaCqua7lmhDzSz1IEcZ1/k7
/jzrQnm+/shrBqSWoK8YX72EwEhLOirWnaiiE4oSpQJwq0R2lhN3sOW/QdHr
mibpiJqBrquD3I/7UXDP2pgJSrSHG+UQPBcQ+JxEExdR9b6irA27q0RodNMY
fDaYuNB83cTz54agEryEev0yOctpm7NRfHxVzQwMSiHNBg4C2GsPFulioL/5
B+8dIHNjA9KBinjy0fHKxGjIEqdj4qajdSc8ao1SfvJOo7iVlSmQcix7gu41
K7zKYwb79DL9Bu9ezFBmv+luQFbKQlAIFqf9pk+vVJk5Om+tz2cR7Z6g7NTs
E/ZThqihRnZl/iPabOPs+pinLUiqOVawRhyn9Wz4BCqE+DQ6eU2IE34t5WSL
kEGZP0ueGDaHmHFTJQp+GBRJSUjcEb5PPVOXyLJSOOYOs2wX6TvxxYfKXEzL
FkvWXeNi28Ou51nqWq2/+r/SWfeM1d1gWQ7meVwx4u2M0eH5KjeGX66CRVtE
bQ9D6FblDpkAIXwTxirwRu5ynyTzYUwJ+K2Gnt9xmL/2Omsgpd8gV+1PKnnJ
GbBhl8e3ab7exKzUYG/MJ0075OGvSU8+zEv1bEy0BlS1rTwL+g/aOXSS/xZT
B9Tzunm53PHE4n0E9f3egOO5kGORXlCXKCo4jrIZ2G0sAhEJT5zrXfw8y9TB
2cSRMMAuWJmnOyxL+F2YXuWuwh2qYW7T/K4RhMeiv5QmUommSKVeY6v6G2bJ
BCnWPCbs22WFHflUe1WwP0FeC4SL/oYzIELB7FKl9GdYiXsOs3lScowbkDvM
jrPLigMIkZYI7Es9NeWrIM7N+5yHVVBgMTjYPxQtzc5AhgebkMCDN265GJEx
xbqMaIpXu9YplSuGg0cwoQvfZftqnzYKuu7eeHaaZBsH2mwHsZFNhwz07Zp4
fYvFg3W5B/g4BCt+6CNCLARtdSkC0PeFiTADmcob1QmLiW40b+NJKVxmoQCa
kiOCHKPzh9Z6IJu+8VESyqaTLIDFUtpGWuXxhMBYDbZLaiw0AS1KVE9pYadi
5P0DJTjBGnvHLTD5i0XWiYQ2mWT8hSPdCYFzcMQAD4lJ8DTaYD5KVrwOx2G5
qhXVSGKnBrYjp/rAWWcPVabx4nOS37BeeReZ9p5//UnXi+Hd3DVkSOEVwcg2
XAB3bnywprRicVn/AAftk8leuRMcf4EODMnRBP5mDFpEURvhrXWk0pRitfAR
Kd8kIbbX631IG6E8ytkMQT+O4eCCLBFrjruRgzZsQvSJ7avP4Vt1oJU7rxqF
0hJtz/PcjwoK/UVupbFg2Cptf9GAUFxwk5Na5X5cdc7ubpA+k2Xcj+ceVZxA
N8Dyq1JQn1HMjyto3dF66APCWtnfbT5lwSNvBV2wL9f2AZ0hs0wZhN5oRX6D
frsOarEXhvQPUfE2CFv7160QblliukX44FlpS46qnI2FJAWfePNQ4H/NC1KK
xTEWCf/LRghdvcILS+HPQp/eq9Jpw6nW2lnNZa56kUFtyzQ49dh7Hi420pEB
8P8ng2aovmZM7xdFwtam2CKHI03IKzU0V3q5OGfTKzCiYQPrE3stDEve98mm
jE93RU45DX0V7K4dTBjTggdL4GTERSS2Lp8dIT6K4xWTfuhK8nQCRqYmWqlz
cOpJ3A3wZezLTZDBoynzRVVC3VmdKtiHIy4LIdSqCWpfGITEdtTsE9+M51rB
Sj6q/bZy6hcwpNm6V9CumeVWSrzUbmjiT4AjG6zMcJURzi2WhkC3mY57q88s
VFEVRPmSI/XPAOIChdS517bFEu/2KMOh5uJOnlbX/j3fuxoSCdGb+ZHjeInG
0LhOUZAqgMJFaZjqKFB0aErlVEipN3t7qn6VgNFkcBJa5OH7WPY9VcGynghi
bku8tlqMrfoCAJ9KadgdCjrXQvvzU17EvILkmwuH2IhySruZEOue+z+ent2X
vB/DhD3m7fY+7pMoN3jZ0Vf+4Txr92pj0kdHCYTYYAN5HC3VR4toFY/OGhMn
OK1R974KxntANzbOYk+NiLps1CIAy+B7dDhBLKMBTEnU92GCx7H2Yg1qRNbo
nlBOhnO90FxrA94UkWo+Fp+ZcRNTtsEa0sh7tYhlQ6UKpJOzxh2v0LPTI37h
NZwyflMRs88uoYrvX2J5AeBqm2bW+Jl2MbRa3FdA3Hk8IKxtERg8lYf7P6/H
gCTWcNPD4qCTgSd+ysJ1zd60tVBH5t2ZjmxJV8UIpUr4xiryEtpUxqOrivoI
/r6+KiglOlYhEevgU11uWLj374LgItV31OeKn4tEDjNO08h1RLojtLEJBQp2
9EwrDE3q26a8aWxPHaumxVEOWoD7tuAJJlBovmKUF2YWxmuO3XriprF2HEe7
ax+PdKbLb1cdflaDXUhSZJoQ0DPTHv+27vik33vvA967lSWLodYv5LP6I9RL
1MDdohMxyOWZ3Z6bz9f6fgKwBrrqxmuok9ZpjtDWTbgqAoDprrbLtOcCr2mR
LgymyhfM8Os3qk7xuAYm2HEXfPsMvk0Q+LFamzuk7BRz3wj9RMxYkRVxlzNq
Op4MN7bDPTqZjvA2VE6vTRKImCn2eerYBAZpLTv7uCmBPWuLUoLnS83qWyhC
owzKO/uR3lVIRh1wHifYN0VJaoPKQtG3t384pxyI1HpqCrZ6vwXL42Z916bb
2wbycE1oaesc2GTlIKM5ZsnVW9vwI67p7kotddWsGu+QLqBXHIdfvmH2/EVh
2LwoDJfdm0R7Ti+70eck6g3MqxWKLRdJgR8HMFClF9A5bzOo+rUmlzPImTv5
xdM1iPAQF2KZk1ZOO5bv3/nEe0VrjRvUiPqG01ckurcTjcvNhqnddXgKILda
wG3tFKar0Sp3w7kQzIOxtBm7tBbM7KUNN1NcCE1OCoJk63ubN5vwxBagqYmg
bbngqP3pv7DWHxwWnDeiisYBvukB73cHuxHXSTJ5iDAXV6cINuyI9OP51rZW
qIwzVIaNrE37h+sn4WaZvCj9kd1F8HA8HFCU3I1C/Mw6l3z76eoG61q56p0O
hGLA5C6PB01iEC2ITSkkSX7vfkJnQti6x5vlIhfbeg9Iak2RqCzTXoIT508Y
mZgoHRHEr8XrozjAfBojp7NJSOYthAuJRlLQcs3i6DAaTuXgu9j2e5sBBske
jFL0r8hiQjUL8VphXyM1vhWNiMeH/Dqlg4rFNdW5V8lOKIaNrVoInDAR0PbO
SJkLrr18RuBD1tpeedoSQBE5XYaPki8c+mDZehGlGo0sX+QPaiJaqKbbfmox
RpSmw/8dt4UYs2+SmjOa3immoYQdUKtCHJDrQc8P/9t4YmPF5KrS767L9Mfl
+zcu7y2d4X9gIlhluZrNv+XmAEKEMuJsagIKmKFbdzQ/E8FjJ17LPK1HWm6j
+wP1qCeE6YNQsN60OnI/W7U3Asyp8Wr8nATSVJ54sF1G9LlQotjH3JBb8iQQ
y5YS+Wlt8TlYF76J21rYuAb/8r6/f1U5wPLtcER7tltgHSiBWGtIMBbn8Xsw
q1rdEAmSw+ZNdQZPf7PwpiVcMk8Z8fE7AC/SPyAJ4XZd43nY4M4w6hNRIv8n
XDqSXM8XqJo51U+zvnLIQr+EKpZd9Rf8Q0OpRtiVeaFvjH4EqnxciiniZlY2
UWQ8JhCtpkdoHWjvESqHj1aiR6yz6vwVLRqHPPf1C2v6Ci9bKjnOlQ2Ofi2b
wneZTeaXionuqQINlocqt3wNI9RKY8ArhGzJN3Bo1FdTBYm0JK6HJPknmxVO
5QrElZ2U7s8c7RuJR4JkPvIry7w+U4JkW386PeRJviE5My6QdDqZdzmbbbIP
jj3sNJ8ja8mGiSAWeTS5wRvUMUnNJuGpWHY9e795jAG3enCaCe7boh1/jit4
dF7Nhoc7t3GDCi5d1qUhSlHr38l3/T7ZbTu4HDzjyNig4vpl0cefctHtnn/o
0HlxW5vry+mXp5fsEUnP8irvK61Ajb5dsGjHXvesp2rqKBqu5W2+ZDojjJ+E
5uJW7jIBbjATvJrdUM6GwurAcqWsrcVC34+Ur/FRfZXccLXbj3BfdbdAlFXO
jcgN9GsqQrrAHm/P4V3m00z0CUQlTYwAFjixIuTFVOxGE76t0kMSvfvGoDfw
S0IHlIUb+K6/C+hlVuGQeVSTTImYGiTuU2yrX4Yv6/H++/Pdo38fcp23dPUh
ripT2HGXIfB+UIBchafkendXZzY3CfShUcSggS34XUVvATgiVy4fy06Aco+A
aVYH2uVmV/n2mlEveDAMVn8j4Swg9hOSj6BVZ4PrilQMldOU7nhNnvnbmnq9
LsLWWTS+xT1TX45MZUNSYyYnUk8IQOvI+CPI6odLiYIdGxo9+DkX6HAJLzo0
Q5xc5/e9SAcO91ArQDLqLOg0EaQfcW+OsbJeAk+kXAK0c+Xy23cw+9J0eAY+
a/FICiIjzWx+XRtcqanzEXIhp2D/sRP7HxFqlBfsAAa9WFnIWsnETHb2t2WK
ybqtPUHj5hop3Jmbdc1Tzbvg9NoW/0yb//XRCPqmHCHtob5VojbfAID8FMIh
tFz7mrPxvYKr8pAHV7tjUcNhcEPSGz+Wr7V29MPWCsAXc7yLguS/LAi7XYFF
6//XYDjQs3+P/N2LKJkVjgk/BWFJrNBScJag7qMr3NpaEqO3etLE7jBk/egw
7gT4GPQmRJMOnRAjE0Pf+a1sVJ27HUOv6BEahsUc/MjShSF7Uc7te4Qr31g8
MFu/qSyw5qm6s08PXnoYegC/WEJOSeOTbI2ruIjuQ55RD4x3Jpg+vC/yyosX
nUI8MeOctPp7F3C2Y1JP6bKZZ/+rK72SF60fZptPUTN6dnPvUvn3iS/o+GmI
spLxphV043S01pYPM0DnHCgP4TEq6ynhHt4MDLz/51krXUITgL5oFwkkAk/j
JGhbhw7UlCKRmEfjm5lIpp2IGNurYD2cZxvwKgygeWZl6g7YXcCywUhWT0zP
DoHg1+ZLSHm+iNrg5bjH/l2GVe0Ogddbx2MZDF+hlKDPkL8VuxT8sLbT9Yg4
Wo7a3RNtNgdlxt6oKgml18o0Py9Y4/xFasSVGlr3P6cvinyMDC3Oj456uAuh
H6aDDlpBbUKtLzCzdOL4ZgoSGw+/jDEX5a5qEGfwKk0tQjBGG+TQmUXDD0Z3
YF6Gn9PpHanuFbikKndXyF7dh8HwQhkyJupExLZNSzRv3K/zSaRjljrHNqab
PrQnYb1IaG+nByDEnGez2qvWuzLvV1bMiDijQphZOrEdhKgwTemGlV8XnjoD
BugB4LtRv3T0KL/RnXei5cWueEfxmFKR3hOIgUhR4DWJg+sFUOeqpZnAsCKO
nZq1PivJAcSfvCZOYENzOXWSyHo39fOwUsqcAuZ6jcG2I7NOBb5WMKpOmqbY
c56CQURrFgcGTZcq/X2tFHwrRY7/whUUwXagZ7FnXEQhwNtj0SRjnh9ZYCWG
ZsROgUzph/e5/G1x84sGkRJGlVVrApfu63emj83LO/EtftdsVVjO7NrrqHod
R4l6ZSzP7x6p16LCWq2fpErH98jlGZV0ezcmtXsEC6KyJt/b/HbqKS9ofGpY
YOazFNncKSJMqyW9jSk7nwy8lJusRpZLqMvrsMTDJg0OAzkIydaHixjyGdjo
NyeNoN2BsUTCAoR3f02EhmbUckuCOT3Gv6QZJsyaP0cCUPeWIXrqseaQv5ZJ
nJPa/n6zMWBsNQKeQWt9kB8aiHzL4r7m5tDopV189H3f0JVZNARThj5UuDsx
F8ExqnkkMIpS9yZ/ZaYRzODyrixBU5Uw6tfqmxXrbEQa9rDDr7AQc8mI4Cea
akla5jD27IlpyVS/r1jbQqLLRZxXVVBLszSDyV8KXhRtNkDeuTCM6WLDc58M
vUa8vGr/6J8igLrFFFYpgE/F/BSwP/5+/jmWMQCuN4FdHyZa3DEkPbiK6tNW
p3bJTaKr0ptPTPxk2qiz8Y7tl7f1to4LJu+w9JB51N/nixU5/DbdRAkYZ/Eo
DhDKzokYgCNYrgkbYmu9+8ePBE+JuuErsbzUBYf3cBMQtij/vfVk4Lews4oH
kUJlIttrlyEXoWsb8mcEFHZCfqPUYH2lNW4yBhpf5A2CNJagcal2EcDjyA0n
/43IAMg7206MpDnsCRJSKBN47tB/y8cPxYTBaiiLN+DWle8AeusD082sBJbm
1Vzj8Nb/VKnhbgM4/XViXXsKezJv5ArjwpLnKTcLuV2lVCfgog5CHNu3+Z/P
6jbyVc2oELj+ryovmoVzrJ9pK/hmyCIPY42iVbZXBhjyghuGUMFo9Tljyoy0
vdCqUSapNNJ4vC0YNHY3MWoNn59v8jQIc/M6uTIITq67VilQ8tUaq+43/UJI
x2fDzk50NCkRarcJA8mZ4LiZ1CIX68IjhHvAZDINaQK7EoKRnN15JwYn4eBY
Kg4pvwaW/mlSF+lnrl/BwhT3UjlcKXXwZ5TdFPMuOs+5JwpDYl9mFtF4dXlh
+tfSZCaa1nPcDNEw5XvtlLdAOa0jP4LaaTRZOOjE250s2CE6RfHs//zJaN68
HOIN384no99I1eNINS6vBr7l3td2fR+i1qrBNad3QNam+7AfD1Py7UliQzWq
w1fuIAQ0HD8NHI3dHdWsApR33G70n7vLEJts+W97apK7buU9Qx9Lh1QSWDjE
2nQz0UATKT8vsH59jGjaMes52sWunf5RADWySYqInojw02TIZiTr1tv9L/9d
2HsSC5C3ykiqf0igl4RcXyJhhsIBtz0V48D4KNWAg8zpGKyHDLulf9t1m8TX
uRVknTGtObiaoe/pJz06rYP3DVFzHvpxsaaRndBsb9oZOlSLke6iec57O3Tp
iZHsLGRdVFrbCTFBV2IyAhmCa2ltJppiOaN9uKWSU13e2xUvLkNZmEceAYGB
+zRAxo+Jz3320SVqBv3RDN3ELCCB3URYppeYQPq8mdZufPiz0oWIuzUjOBkg
46lasYaXdwkfyZntRMEG+M96qc74FkyQBib7srDH7Y5+XKwOtBu4IUbXqlkA
4qEd4p/JfR5p81/m/2KKvv8tB1UMV1fRIKmDUHc6/a8grO7xP/cJ9BDEdBaE
4Mj/VYD6DVCYYAUt1I0C4tlbC1LejiQBJguEtFJOxfOLfWBLsmqOwOgdaDkf
RWAqHG/efURymkG5spWrFKGIcgY7xCcsTD6OwAAtyZVWEt1fMgVT6qVMZq2r
Vw6WCanm9RrLKDLPFg80CdL+HFXWZHONqzpxUZHnXFmkOMdCznBEkKS4Cd6B
wB6rnTM6xWcxU6GlIx+WkRIewgMrN7a6UJVZlppch6narqaoooi6Z3LEtG6T
tust5P345Iwy6zo3+5LBvS0lAw38c60cUpmxPE7nz79nztBaUuAvKvJKHynr
e6XZ/QDAt87qCcU7LNOLYUN1u/Fomr1wZfgXCLVBdBPlmzXuTXEC2EydW5qa
RcpP1XM1+4LbF/ouUkd4e2wH3sCyR/1vGBtUXmK1NXg7Pz+UBMcnet9YoiU+
ac9V1oMDMd4SysO3/x+iDC+STjf2sbcsSYzwhqdWVAHI8MteSCNA6fehGvUz
DsTlOPr2h0Q690E5SNoy9QAvT7/4DMjnE00pd8SSjlLb6+aq6TmcpaEvFnq/
GylPC88/Z7dlGoSAeldxp6SnZ5ItvDSXN2i7Qsgs8lRwlHlAfHG4Up5pwwrL
rHIDqdtkg62KNaCj9BlGIt61tCI0B5zcsgHJh8N+M7LzURH6agAtZvWVbUlB
rPbs1EGv+qcC8j50Rc4okbgprIBUb9OBkjGbgacQJC+yLu4muEpYeUdYozBI
0EBMoU2TTHl3wNXc/I69yyiDTZAlS7fBUnOa0fPCRc9yuwTRahDfudhkTSr0
MGR/wJLLljJzWRDl7TgZZNuDSoP6lHM3CDr/JPj781UxtdjeeJKgIPTPpOyF
s1jKOr6s3zlKD0b6PmaPnGh4CfHkzNX63WhIxY6E16FjqUVYNobK/tYcylKy
wjQezcApVQ7c5+qVLs3qijnRR80YBOTdh/cOEtnEKIWWyfKrzZUW1dTuklyl
X4UH/YJL4tNRbp/YOdxT9LcasyxeBLLwgTcF6YMqWbJnz3MPIgrT1vBJYvZT
yIKHydizYQE4pS07B3hMqFB2FkpmIkYPtD+gxXb7SGmMwtmAIHXHYpPlTHfP
VOzWFCbVexTcRAlz8FW8COfCxzyZIU2GKkJhGBjaRhtVV/LrS7/MpjB1fTq4
6ttOt0xu19udHAavaYSSLHW4VnqQje1EnhFQ/oHToM1zEH9TcXJ5+5lYMdNa
u0M4PEdxpWEZeZ6MoNLPh3Dtfh+RgIbIzwtU/sNd6ToJtVDSLA52OnDcu3wQ
ygAzR6nhmZKPY42twZabXgtWmroOhWO00WkpdqSgvSablNNIMQawtRnqLLrW
Lgq0CC//9l8OjpBb3URfRwuIv6i3bHlVtKi7wxG9O6xz0JlP6GpBshc/zYNW
PDd9/Uj10vacp2rGACHjWPQhdHQjcjByJlrlOh7auV5c8hsvEGJYzXH30BRM
+6Zpx3/hS8mhzQz9y+K7H3TkjDPdmyXInP7c6CcpvxZXlTorw/lZ4tnEwt4S
3H+w9PvxoIPt8EyyJEfbSejLDfPVgnCyqByQyEDApE9RLxMk4EbP/Rqrq8hu
J4FR0Vy56AlDmPkO3ZvtrMIyyYnkbN2tSeOH0befE+rQHfe2jYeLADeainG0
e+CcZWDER+XLtIZbNuKXNrWq5odBzhTqtxnfZ4WbT5YMQzhoN9PLubFY9yFj
iFTEfjTTzT+HfghF6tGZiROGTJ3i0Chs9OT7phBgiyMd0i4KthKXiq5n4Ezf
+2OnlWy8NQm1IKL1YzMI2B0WhG/Hxo/3Odm9FVhklmJO3k7YhxRWI9dgRLku
54mUD41K56wJUYV0qt2LoAsfVrzERxioZ7ZoDYDoolDhZt+nI8MtL+CF6lFu
xkrlVCtKFovsNFqnAa0k0kIBpuszsfRlkhQoJcTmZ2CnbfxLNUgWOMVO6SHl
j/ypiAUK6ftzpLjomjc5cwd6Qm16xM5Dli6XNkLnnF01ZBTgTXfkvzHRahj2
6UE/cV62bDsc8UR6ULVPCCHeXuc0K2meg8d/mI7YNPKk37s5pby/D0umz3eT
upRBWaAYWk79R/q0lVT/+2u6us2SsDscxHcbCIKVLJcxbuKK85xEmZoe7/lW
Bk2kmE3PZitZcvb9XmKNY2UT/tV132Wucja0K0JY+xUBgaM06JB79mk+cf9W
kNXShi4YotLTo/CAm5ArGWpb/oisIviqy7WwqIb27DHwQdIk65K4x5m6XP6V
k0Tqfk/q1tbwN0SkkCEt8renofVT8vmZ8CM++Nbhy7usvxwER/p4HtRl4PvA
KzIowC7tH4IgjIQIqv062vsjCmxIYLBo905R7dRJ6uqwuVlJKSa53P1lIRH1
FWzuoAyTVBw4whqaOMkZl8wkD+JjAbDTx2VipPSF10wlNWlC7ZvF5cx5IWnO
yC8qiDo0VZhNuXjETJNKzx1aYz9mtBdW9Ot4t75Yi1yr+PfpMbFfEq5hcYtA
wi1tSFgP8/asqNQefqgi40IM1/gANQ48Q3Whf2tQmLYKSRATegGBjVns4+Ze
wU0AOG1/Mk2nNx27F2+gIBQDa1G5uqwN0WVMwH4Di0Nzl57TsBc7VVrXsKFZ
vdFxE7y8cGgniCtgymgc4pwXMd6c54osupmPBx4AvVnSUHaalx+wEaY8jSMG
WwST/Sz2rg/mpPI8XCoiftb6lZ2o+pr+auM/77BTJClNqobmRIRRIoP6QQdS
PsvqOUCz/txuB+msN1xFfVo4HYjPNnGOuV9x0rfjEdXmxNP4ZWWt97Gj4Ofj
7n7cGj/6ER0TGN60wMCATzWc4Rmyk6Pfg6dCMYCx3oV6C/EdBMHlLkLU6eUg
LJMYPnXyuVde5XlYQGTtPZJd3+yDIIIphm4lRFvi+teJgFfaAzrccFDIYmr5
S8fGRYQcYwl3AX7KdWoFi5rCTXsWFLyBUsufed7sOrFWAQI8rFmIpJzioGvV
Y7DPUtfc290jjJz5Hx5zsUGzYp3YfWiGQn/J1QBd9OvdS/qcuXB54n29JYFl
ua+YONrFnWP5DyARpOIhpiN/b4mn+Lq/a/P1aMboCxHITUD1M8jpuke9erGj
NznTLx4lFzFbEzJXOoR2mJBflbIc42H2F6RHmP+NdgALLaMrmsCsr6y5QLXf
cHnF6hdAUuxYe4PsV37tMgJcvTCrWrINg0s1hhZTWYQCIQpeYAfE38Sg8wzC
4c/n0bjrAJcdQ6bf3BfaMpGkPLhj5rVJ7MfmAHv8/11uMR2oGrK8Rd7UL0Ow
CDbj+ZLpoo5ojrTcq38z2zB7Unr0/hBIrNqhoRHL3zV+3UVTZ0WUXx7bWYP2
F+SWJAiETW0Rvsna5UdQn/WHhX8lBp/jOLlekEnY/eFgCYfWRsJT7NzgNnaH
ZxJMbk3fpY6JzAv2yQsjwwSsDUIdDivYmbkKmT8CCxVhBovQRzN02/TEOJnx
JWsAwv0yj9iW+kP7hiyhILUAOWDsw5Hu9JmDNfkMW1EjNUcA17Z6iQWYkCYt
LMy9bckmJ1bCdvc7C9Y9ZahW0jLxFFXrgxjsfrfjW40UYC/kGKBdxZY6AoP/
z+AUoIPbAKca84iE1M3Xi8PowmE0H6PB1K2Cc0C2nvwyWTOpkf5zQ9WyH1Dz
Y/tWPiYurODWmpcf1cfThsL7mQIDYxQWeCGjQh5HZ6eMXiVQwmsbeABu7wlA
Zra9spLD/tltvtQVJtziD3yvv9ymvXdOJ8G7H8apFWyaV2KDKLHRcKIP58C+
tgcUctREXATCeX+xGdYwIZqWhqhuQ/kiIQXksEBYofVvreOZ4jjwE2pMEkwX
0oC0OksDlEm2dNgen4784+LJTUkhuNjYZFXrUxdTETmRXFsmj6vqm1UvitN9
aOoguN/k5gIykk+dK8rjLTG4tPtTmOpm/ELxaK/iwFuE01UPMGIk+yZ2NTey
+8o6O+/rcE61HeKDDBCQ9wRhMpExjsPvvMQrL2EEhPWHhWXwSI5DBBq5zcll
R7+8UTex+j/z8iDaaIF2odTSdysAfwroFVoI/1lS4l1WOEH4szAN10NMHZ3r
AITbkAWsFZXoVXC8oPb1EJyUOkZ/Qj4nTA6MBk4yRzbcuMby54hkC9NLsUmO
sPFiwobbDKWGXQsv4jKEGJP7hRgPUQwVXZ+qMzmZhg9UBferkJEmw9CrGS8L
WS3FjAl56Al5u20dcBnSuusQHAHuO7u3BEMeW/2ALf0L+pINelBD9a5YWW1p
Nq/HJKejULnVEM9TLs4UYIrcswWiEK3bKwo0+W6ZTaBVJBGQbwc86YxBQ0fl
ScEuL8SO5Wwmbt6X7BEN+ObISxOKDMc7rkaVXtch0w4Bmy4klO86pM1XdDDK
DBKVPTk8+MKhlKp1MptZ9N6AF+q9DTvOGVgvKNrRSzDvqKmnQZzknu1L8hq4
ndmrFd9z14vgGnkOVuxCtSa1EDczfXeoUBYYn2mGIgtrBLx02tIbl80aTgFM
m09Jh5GLhwHtfK7YE8iaynCOmzHm1Zgb0vXQsJgTbrECLEg9JcRtjcxRHbRU
ORC/1ZGLmvKdN995zT0pdbfccd0g38oMDv8gFWWBs0aTSnJDG2336thwkb8/
Nsd0UMTqKjexe3rfmJDadnb80Edqvp9hRz+mjLvGVPjvPNvk66/X0IkOt4JT
jNWE02fh9ZQhttet6PVQmOSdSsETneuIXUSZxwKMYxFPfNMYbHLsUTPLnnLy
ioNJzkVBxFv5VlulS95qFEsZwPF/pJFwxtTHz0saE5pShULNpND9Su3mCsJt
9u1cXiH+wORyaXM2rAbFkAssHAJSABqWHcTJe352qHN324loIOOTzs3djThz
Hmf24JxlviKHjs3h1y0ZYMM10HnM8Easa8u32ZhPZARsflTvgddclqnoXa5g
M4tkNOewpP+75vwsuGla3bbYwQWZcoib07B+O/2W6/baUXYIukFihYwnlfvs
IPFyWekxB75C8cp+UtVKBWM7cB7whSmZR3xBorWYZn9dJrl/GHNKx6xHwsZg
jvDysx4X1HiECc/k9zQbN179KKe5aV3RHxq0NU+PwiJKOq6Z3fOT8BUsEgCA
eJSYSPzdZ3HDT+4jBB5pmT9IL9HCZqJm4tpjaiyRbx0Q6+OHA1lVt4bUU6Q+
ttFfG7jpL3/zdB1U1SBRqMcEjHqWpbV2xwxz1449fxtyRZgmapvincQpzA0d
g9xtZIX4lsqb+hcTlcdIcFQqz81lzAs/ErPmcd1uGhqDesE9Til3xey2ZJN8
CRTbNvi6ZpcqnKU1agyGkLaBeTeNY9cmrxJ2CSYb1HfgyUqO3FK/UuwoBexX
v06NkR3SDQNiM8F9yXgiCKL9g/lFg46SGYsLxnNVoPOuCI3SaL6VcsKzrTAW
HYchZESnZ17reOSpj9/7CroZEl80232tN6ILwSd4Fk04fOL+J6kyPrLnf1YA
MIYLle+O0zqoN3dwCRl5+vaO2Bdghvj/OFidcHFXLilDrHfkgOgfDa5Jyc9Z
G6bYLmCJvzS6XFcj7RINY1/CKriVRurJN1iC4yRad0neim8IU6epCClL9k9x
y3aEbiijrT2e9//KplWm3nLE31L1miEdnRzVNGqLhbRhFDq44ZkOE3HCFaqF
5F8fCZWfrtgrdRs6iOsXrR4LVq6fyW27NkVuRl2Qjc6VbF0dUUSuNZ5cnr8x
YVGWXMz54e85FY24mm5PQMEegTjUsEAFMo/FgVs+cjolhiSWsOiFZ2BW3T+J
yX7WFoeukf74L8ta2wJKnL/QcTEHb53P7tY7FlouF9zhUZMRMH570P0p9xk2
6wLIVZHjTn+rgtT5GbEZShCmfmETOwDvCOmc9bmT1Oh5sR9yw414tEgN1urv
wP072XgWLHiCJG4CRjSB/1rGjTsnPdWp3nKi2yulBRG1rdc4dhtsJeNGrOUG
PoRFnxMhFe+3jErRrCjnsQS/xiFda0v2HPnQCbF+b7EhhFG7b33N6y1aVWT8
V4pIAQZTVkW5GaMdUGnZX/eYrHLbAiucukVaCR4A6AL/b6rs6P2jC/zuso2T
DjyAYs4EqT4SWlSdyXq89eFe1yuagOn3rb9KRfyYMb/CwffggNlblhSCd/Mq
Jz2qimczEt7qEC65EH0WvwvYuvd+N2GzWd3OBIsVZ0n9oZdl62sEaO1U+1XE
rWHHZAi7OjSADuLZ/aVEbh6wUyG2STZ3ETtRYvbaF18B769UsGBPfiJ0Mn6H
bPrcdPooEMK83Hoh2qY9VOh83QF+yLxyqcJC6wx1e/o1xr7Vd8sARbnhKirc
MkFePbUBHqudyNfY0mo9j9GWFvRsHG9s4JlVDH/dXkJaR1jYwh6EvNIjBomN
HqjuHLUs6pzQua0U+tl3PH88ef31oIm7Tla7KKnKQWMHJG1NtUqrz+87G+6i
lpyGVC+sYtj0b+ILuR6PR8NHQFlPbugYO/hHnIDsnIweCbqco5BxQeC5i34c
UgXWc6VGgAyh/fuxtFeI9XE3lMyvdWJxvYI5ozW4nnUZsyUTD03uRrAKSOHj
761R0Thn+qUCKvu/bGK1UuUocmQUiUh4jrHAaUECR/3qY0ONAbJeuu+enbcB
zMrcMf2k74KD3ZcCdds7Kb/NUVZcZqtZhbsV66zOmUuFpVZ7nvHa97DoJX2v
Q7teUghyiMWyiapudLZkZeRlPSL8dGkMmSS38kOqBIb80ldF/giaoesaUMdR
c0KZjmJIccxyh2tF5ZpFs5apYymNYXdfJRJhynV9iLUvFId05O2cwdWrN1nP
S7L46KxrglPlkqL58MyiNrKkRlQkODwolBo+OyAmXRmXFinBNvJdUJeAhyig
1749jf5jiivEGgbZZw/QOvxWyDy/Se2wZWlu5LpMz6wPcrvVBc+zveTzPHJD
YmtQUm9i+Kj9A3ZhMj2Tf3QCqvdMeQ9H6jIzMA9w3FVZKGJyQ6szNtfLy62i
wYerIPSG58jag0OofmY+QQcBw9ZA1yd/88Ox8+3YTAT9naBu/FuhtKhybPYa
PnGAIt5lvN1uKxzMziT7A3EkrT9JctNx6er8J3dszwVe8OryOdP0nTKYXEah
Om+U2vr9hwkuWLd5arbSmll6yE4OuGNDcHBJIHtBsAiF0eXESfF61v+iRmcP
n0IYyK/WJ271fejAMHc0TzdYF+SaGp2NGezh9Dh7VitSMfKa1tYRzymBCNZd
diN4FsMD8BF9qxPBWKBWTwjsaWjlpgy+bHJRvhDSW2Oxje7ckBmsbi9P0hv/
reljbaO2qLjihvM5PiWXdh/ghPlircyC3WaqxKpBDtbK2yF9ZbT2lIzJqfst
KeP3q8dwv1k6SZdQ+1JwdGAnJ9gQ6RMZDbWJgV8J/bPOdulgK47kAxnsC5I7
GpguEsqm6LvZASAtGPqYS+fhoMEbwYCZiHIuKX1c5Dps+Mb0JZr6ATaVVLcQ
/wN02Jxu21bnu3Lk8wQKKJdbNz93EEMuLW8WS6qdjG50nBUJhCgBIFC70ikO
F2cizF6CHOa1xYJ0jGAIMhh3bscbh1iZS90Yg5SfmaiKUZlUDRXNsyT7D6lj
RTcLN5bkzI55RBbD0OfXlxHat+eC66X04L2iCvC5PxRPSCTjCR1QiM8AboJD
nvKH3vz9oGItmOmX/KeclaJx1myrgJp+NFU8q0JPmzkbbgP8pUnbucFYYQQ4
nDJM7DONvPkQ5Q9mVpcvei1RZcAeK3DAwNsxWagj+njN3QaEwrBV0caFOc4m
wQsph/GhI2UXdCaxzkhZwE7lceTt6TboRtzzbaJ6VYuXZ0gqASm2b0MWTY+u
RBFxvIA7e83q06Aymg1PIH24JOh2Na79qebnXtP8p2xOoCOXZDg4qv/YJ7Hr
GWjKZSUb79PkLfSBEe+vReOZmcgKqVCO+JmcJmVOYfVZbkO/HKIkvLSY0ZTR
3qVhQwRvHpylxBJhlkNejoVIm3WUEx3H0QX8o9gXL9FNnUlQs+Tw04HVBGzP
LVKW8ChAOrpAcPNIHOrE/0KCGYo2mszX2Ym7axlaIhctJcqMbcXXPHzyjy2r
VhdOlPLyYIjaSCVweY2GOpCXQ5ixfl42vRewTXEUfNJmc/cR0BOdKvOW//Bp
UCWWlRl3CcLWhHcmUC+/LMRM0oZWojGR1WZ8ER/m4/WUu9y5SSdaDVZMVzrc
88VHIJfuA0HJEGLP8tOywPUAChIQ2Dm0MkAUHsp9GmGSfeCD3vbqbzyxSreK
0R8YF4YAtxfHP9IdOPFx+014i2adLsTTnZR0ORldsth97sD8DviirgNVkCai
LutwEIigX7UnS+4g6525PesCZJO2i6wMwk/HSDrwclBfLXBY279T0M6BXUTW
EYbfKSEgiRuow0ncJzArT5PjTkJnlNrrO6U8TePqsvvjmrTRraeG4CekLR9r
rPhR5oYdopubv4zgvAqrzMN5/PxvGPK9KmwGvwjFdYHhgO20jfsYYgqyqtRJ
7DwvA3MAiuKF7DviamJcY8QGp9pX/Gf3IhQ8TD+luBkYDQmzoO19t8LAEsz+
A3PtV7MO7yc8ItI9ZnUuYN5xjs/Ix566d0Wuq8Ze/l5EVfj3FDXn733354Nc
IQrMk66JhonIqnblBWQNjsvlPhsVi19j0pn3BH4b66rYXxdIw8W/U8GdRYBo
iW83D60F1bXovbb//e70pXFyXxWOwJ6DiAFh/efHeb2sWIjSKEPuNDYJfgnA
fZcH1eQg1f7BPkpHSlmpLPmA1Rbj5JAmo1Xmgy6Zyde3HYkRBnSejfySOSsB
9i5n7TuJD4BsbqjyqKV9sAm0MLUjgLwla+rRCx4bV4gd8T9CaJP/xjcychQJ
4DZTJWJeGKpjJQtbGZlcjVMWbo9fHoyFer2a0zhmfd+J2qxzHQjR9DTR1A+B
FrJzatumrsj9ifYS1VySTtw1W76VMGJp/pEy2PIi66k+37/CaCk4a/njxvWN
4RaDm5LIdD1Ryonud/Yrfzfuh/Qwe+YwfIOTATZQLupGzOND+ILGSqBxdqnh
oJPRpYFZNDjXMl7KTkXiPg2OZqNIs2N3Tz8p6cHs1sTZlcNSh8hwuDEZW7gM
L0zizLN9k3h+SqTJ/U0ZQTFeMQU5PpvM9UehjFQcIyu7+qz3BbUduXE+DO5h
TbqcXerVhhCfEfKkHVB4a+45iLaQbnzJsxireNF2BN+Ik/00HQN80SevwO57
GW35GmMB+AV5buCchURpM/QzbEmiTqBVnh8GJ+BWSSqFpZWLU1Yw9oNNm8GQ
PHNLWHLZNtcSqeK4/0bZ40AFhbDU1/kIpdhk18pDcl8WYXds2wTdGSvdJNNn
v9A7jnxUaXGMhTr/p8rNEstUMuzOfxasgRXGfqw16tjbkS6nlN6GV/M3W5Ia
ycF8RHiDEipG6rnbiblblmIImhntz7ZhBDnQPgx7ol9GxbvxXdMju/DPJOII
P7HPy3wXMKucT84bV5T6lEdG4vDmnjHIQGLNMsFOPVBkbNvsPDB1VAkzgMXC
gRxXuRMfmn4ykeUsC9m2Eh4wVZlC7NbdgmJa93ug8tiBntxDImi17gkEu6lM
JweJ1taNfq/RUTz/TuMTw8hgZEo2IsjrjbikZr2SJWDRFs1REPxDZkvpTEDz
GaRxO9zNHwYWWinEOs9wKpbI9KEpCEoKuOvhUhxE88P8yf+Gogb/70g3gOzJ
mkHuNGd1tvwiwvAmIlmiraBjCDxE5duZMdIXvlbjx5eJ5Or20Nx4uM9p/b/t
2VMghs60NXXaCYaFLu2t1PpDLLrM9+lPy3Bqu5bmKKZmjSwMKnnqaGECOkDj
OwW8q7gKgrQj9HnPcPIoKzbl0B15ZNuT1IY3Mynt6JqHKIM1vt1p6VHVhkpC
7sslicqwjm5vswY9hc3pHIZ2xMCXLDChqMhlNrShKN5tOifPp751air+R0d/
KKyTwKHHvpZNIINsMpdT76/J0yhxvD64YNUy59PZhmAV9Gs2OibeS4wad1Mx
shKVqMobhS5aoh57cfQZczqnfgn+co7DMeVQwPg8LZSvDIxLE0aIllp1nTPn
L2b0KOITkVSdzHCdw4FwKaVmutj065A3AiaoB1IJQ9E+9YWlBkDa0h8/sowB
x6rGvGOtwmvCb959cHtaVq4KtKaavAI163gjTh0I4nyPUosMyXTZLWxqc5gA
uQWAQaUSosB812M01d1wIKkMSAP0KxwArpQBX46nk4xqvDdYHrs6mE8djLwA
QZzdueptPbqdUnMlcp/3Gy0b6/wfAN5O3ucA6sQz4Zxq2Y/VI4WMaqirajhm
3gEQ7ULxj5Ek9no1mhapln5lyJOKNA7O6oGauRbdi3b/hSUkQYcgyHgaezDw
YSAHZeZUXwHSGvVtDQ1LToahSTJpdn1CaBDYagFg0DcHqxmpWbH8qvX4wfsU
pFBfoARG/AiuZDRJ7WMwYhuANn7vWIOclGJCurOkrtQV1dqScZG58GrQy73d
ekk66sUyf96uoihMTURBOZxIRqxoIRmimT9AOdq+3a8Tg6Bym+aAzUg4m1xJ
1/sNxD38iG1mJhKZR/8S6Qnw9d725vfv00Bgj5lZbJvDFpMYX235Of42nyay
XtVwahFsnb/qbSj1+z296XyZr0OwGyUCn2EbfvLqy7OustDuXyF8PBUfI9Ke
qh+XjW072HgbXY3tEKUoxRm2rmvNZ0Ky4yykKzUMWCGkqrP5jG9H8TCUGD2y
HxzzkdikKbgZPqyg3roCQB1gYKs8BEf6JoXuym9UuwopHHfgISq/34CsPRer
Nu6WFs0CrsBbsRSrPN+5ohgPT7Jjbb5/7QChePL+mX8gbIGqxerAFA1r9sXF
eObhQW9IlQVB0Pm1yWrmPDCLcOCgVjnf62cLV2FmO74VdRBFt4BywUTC1J9R
j16ldgvcIupuxnCUWHy9lv3qRD/TK6Rt7VwN9bBmsumJIhRPQetc8MDBJZht
sVV76zHIiM00+b5F76OpZHCGuGgp7sbPr0OeDP7UAqr/wCV+0AK4uAveq7Vw
JfZej32r98I3WRuQqUxBqLA9K8dc+nK9eBQDs2kSWD85H3WTryF9LnbHtMov
pAg/YIyif+s8F581U4kp7hMdvd/U71H8Sy2ezleghaaFzBcqk5P73cTwliKc
xN4GR5rmf3pNfcp07qzuX8HGQl/jlBBrpr5z2TX+pQUHELp3za5laVcbAgCv
IDkeLo+h7sBZXMIsgAsDY/z6t4B/N/FNpexXwxVePZ2MoYtC6WlNCWiTp70y
V1K+p98krxHEfhMeVdEl+Iss3+67eCZBZvmtOt7JTrM2ZU+HtjHGCCeqvfBS
ojDh8Ju1cTBhluTLVCEf1P/f2tn6cqrwEpsw00EynkJyWhxdQQLE2zFa0EIj
cemGLr5VfsZo+f/vEO5Os5s8tzrlj135ngo7ku7O919LIEhVE44YXVvAFFqc
0KW98v6lNVlA/QvBTk37ouCJLgHcUFUvgKml9zPv13t6C4A7TM4JbKUD6M8l
lsOU2JMUUON1QBJAcXi7XbWcpZ7kD4IDQS63rc88qs6pXmZMrZi4/eT9B408
6J1qG4ToN+TUhcFX0j0qHyRiDqpsNbs8Ggx9Jjj8izmq4EtvW6nfFPIofDDN
mZb09kLTbm9ealOIj4PO2x5xvzvWWf4A8AuwqQrCym55uOt2bJYKMuQ9Uvts
PE3Dwjg1sXEzy3VMQQATNB3cKampVWJ69Bv8Te6mLceRThh1RgVkAshb8lO1
2AW5nMGtqSYcWxA0ucc9i1lqbWdGuBZIuEQ68YrkhlcfpYJo0Fubf0RXujpX
fXKtNjmJvjDAUPAIBEyYt/Vd4nnk13X2ZC69eHGz2r5s7D+Q83/qrxOo0uIc
PDv1adXNrWyiOyGh0xH/RYbjtCpq1CGYtB3W4YTotTFGa3H90dQmwYc7rHs9
v359cnOaWbRLCpfk1OBDvHFP9WWs/nL70hIYDXetZ220GAyZFf9YsRlTxrwP
WNb7RMtBWmMXowYTxJMJG6U8LQ/+85o/UWnXXHuqAVpHt8lJjUmOw62UWAch
cszyGbUgLpSEIxQqH8UpKn4urOWL3sp0c8ItHKF8KDUd+Ag23J3O1P7x3/9x
NcVrsR9Qv4gF4ZaWMbmw+Qb7roS0yAB81zNsCieCPnq5nNc7AnomXQkDrDAO
j7zAa4tSYdWq7l9Oplrl+QWXGcEI9E15nc3L+CO9LXues/3k9GrmSccHS4C/
kHuUYpszDx3ouAEJ7Yuu1cNh7ya5VlObByoV3bWN6NHe03nndRGI9XNzCRod
UtCjfeIOUS+T5gsHFpG6cU3FTSEQYme1PosjkKiUBvuAYcbBr2QL2CKgWeM4
w9ZUoxwdWtKaNdkwbZzEWzl2EVweTUwRBlaFOUUUiv2hv/xA6sOnlSiC1esd
VSzvQ+QJdgBKvKIU1fCaIrtrgApRxj/5bwnAGDfW97misdKCWHEqCcJppKVl
4fvP49zlQt83w4YvBCOv6S6MXweUyHXFw1HofisVKJf6zLAsHS7Zi9ImHRhU
3VorJsCfcAWokVLnwZ7ug9HK+fiOzYZMBHjdIgMBCF99pU40MySto8HCreY8
AjwLQyGRoVa7ij4J95nhpRV6436pbooxrnWM5/NouXWyq8PNtftdmChw+bmY
B9whSmXTRE7Z2kgQZSGpjGO7zleR/monV5gykofcdYG/pJy36XLyP2Ngx4Mo
Dm/HVD5x9gfWk/jh/LtTv8NRWUNF5bWUckNJ/Y0xT6mgvWglNEwbsd43Q11T
IjG2Yuj4FvtokfaJjFUpjOxcAagIaeRTXGhlcCkYzMRitsPhpS+jP6dl+8mq
6n1cMEZJqmTaUhugMdQjp+oSAUknJFob634Y148ag5m9f1oyuAjtO5aTWq9O
Z1mAfg9mPQQAiENJDNGCI4eAj05HcLNmk2mVgw9vm/Mj4Nu0lpnkElHitriv
3eKJTQnDo+Ihjd0kWUxjO+MHfkP4loYlIQdWB2yqseB8g3MqZKE9HHC4MxFp
cOoDiFakXfHoxlTV4RCw7s7znveFfXBNHet7TI4kiWhOsSSLQoG45ALQg7cP
t+0f37bH7PjARJW+uMcJseD3wvXG8rfrp0fDQBj6uOLT7A632IrmIToK4nVR
Lij3MWw+OpVsrhmNys7qH6p4yjH/PYkBQ3CswBItTgMbxpOOra2wOkBQ8aFG
p0OammeR0K2PgHQGMCmzQGgj90XWuNQMnJQbmCIr1yFiNouELFC/ha1DREIu
BwbQsIyoasiGgPFU2yEFmIJ086EzjRxFcTl0BfzKipo9zTFMI+vPBXQoPtrS
ZGAaNjpjuS7cPjERv+EepQvx/2K3T4B+GkhRZzqg82RQ5Rb+p8RRtH4v6fEQ
SZ2iU/UGAiIbfUZwenWlXMWceQ0iZOurZW8V9Zx5n3MYmp+vb1XUM87kfvpq
ZtGy7REW07PBBSkUlob5gewPfI/SLQnCDRAva24MUt5Br4hsjPRZR3de4cPa
bw4szFxHlLRR9PlUp3UBmngFhnKq9fKjGd/iWavV4rJECW35yEP4Ypj9SSaO
kLIG6VfJhEDMcBtXQLISs6ymOK1sbS/bOxlJV9dmBu5l3T84BDqiJcrG0y6x
BbhNgtp2r11KaOXNBf9G5Ga40+QiySTZ/MsQ9apKLH0rnVmQG2u58ioCtV+B
mOXEza2RRAbk5jGLQAZMFL3E/n0BksGWTFteK7Z5mkllhs3Dipw56ATE/uLT
CY/aRq2vLYQN16qs1h+F4Nbmj7fkEMqQTfVx54JQF/a6vwibXsrEbGWs3J8J
oz9nGgH0gIC4BbvVkhcS1BLgvIA/2HE4TMlW6Au/SHmSaL1ElPKtXuobMxND
VvcriQfRXJrEuQ/RdfEdxlkX8vIYw+7ao2pvrIaVofAMbBI0ZjYer7w3QTRz
DrZUYcHrhbqg21Nh+PyXyqbwPNIiX0PudRBc7wHD6NR8XIiDVwDdyNBbcOuq
uBxiqjB2RCrBumZSzfT08Ia3f7v//kpAnjzZFneLKXT5OAc+QlkBOidXSg0i
DiLXdnofvrT7nTUFFaeLHyXrdB6AvHP2eJ7oMS8nzNhuBk2Pb1a1GwZtD/CC
f8a7RN+msDfNXfiULWYmhi/NPRyqO609JhTRz9cYoVttyrn6pIkNfXNdI5gw
6vMT+EIFVjw57WYQOCNOaedcTs9u00T9CbgsdR6guY7uERY1MiB3wM5fdv5f
GwDJWuawUJkbPmsbjks0F43lEdvM1HUP+MHvaPr4/AoZeN0dWPvz8KL4N+SU
Fu2RuZQo56rcmbrQX2JGnoU7LcdZKoPqod7ReXIseZsfF1nNe1gLVTAeX59I
sqDBewOw1CdleAYybG7+GU3qGBd5xlEjDL9rD4jwiBd6uyDGnAkvIb3QVFuV
3tmD3+ayM21akSVA2o3i8gHCCtGz2/yMIrD/YbwyASvRbZGMQ8LPz670ZZu2
zrAc1YslH+syBg62wXlgHuaw/dm+KvYtag1tWVt69LY4YkQ5RLt+lz/Z97te
7dUzF5eIyaRm4EZaKurUJMfCV+Fz/l1RmjGjmXxYrX0dr4xGT4xNQvV6BFBY
hZuiLi/TbEf0Dqf6VQwDeofcC3exV8+EJW3Sl3GrF1ot7lfzztYfGPi7dVb0
8Y21a1PcRfazpYV3WuAaRTd4kVkDvsr45B+8L3jsa8NUFWUCYBA6Z5ykLa/Z
WnWxaakw8DBmLNx5K/MjxHe7OO0CLFBmlkCHgQFn7cOU7f445MpFN/9HSMUH
BniaDkUTkj8W38RRouPSegs2yq2PsN9qkAct3lO+ktKJuSn+ylU4kTPim7mU
RadIbD9zQHqth2oNlbHoqqi7SiKP0dh37HW37SYCpJdqVuirUwOOOSCZv03m
zQmkbn+wlqcywY6MTKc1H6+VoagXlgVdp3578QeijGnSFIgSp0GkB28CN0Xu
Gyg3bdL5lJ1Jn0Vv7x0X3N1HEslWotQy1vBMDglPmiq0Fcw2tU37pA/m+bOo
yCNT3kaGCL9iIxLRqcodGT00TAsjeUKfAmBBM34kGYveP5S5sMyBeSHQ859Q
BeJCjD6gBZY6y1gEYQaJGycCNUXXUORmiMVFswSDHwilutdqD5zby8EQaJD+
bZKqhtW/FhzFKFoAzxnw/b4lK7NDcfr8aRQlBZlHL5OAy14xaXDk1IjfV9ob
OgE3mVOlZIVKXFRGe8BgqHxycsmYUttZ9os3ctcDjL7wpbF/QcpEuRpLo67v
7mnpnBEXJSVM/0CW/tZzdY/NjRDQAqyn1E/8RSj4gD2tMzl9C2L8OogHrFwT
MrapPySs0diaSHrPI6CszSDzAROldZayCpRuNYUf9cxWNSTL7GYc8Zch659g
/+KY6mkAhyF6OesBosx0c7U1wOuSrnxaXrHRjDRDtwXi4BwQhbbE0A1YYKiP
grIZOK9+dhUrQork1p5PiqLN105ujYlBc0EV/nvCKo/snHGquAP3gIxjNPe7
XXveW+TJzVnb5WcKNHWPCFs8J4IK3Fp9raOcWE7VQKjBIjiSy61c7yv7ARsk
abWmTxOX0p9O7AOV5Z6TZEpunK27zgq3lsWbile1U6F20Vf7tpSLmOuwW60+
K9A3rrQQVZk44hvXjjV73ASfd4umBymvodwCJ89IyuIKj1C2OQTI0xrP6WBJ
Jahvb2/+oForS7YNCsx4k9W6TLpWbOgTtMlQJ7opQ+e3p9PglqbBVUC/urgM
CEvW7tG5+dTGhxm6mJcRnTxWhDwAsTjNNz3Yy9C2zg0RWfigtwElqyzV+iY+
oNZbCW4LuMTUegKCWNEL7XqiTnwXpMRm/MLa8UoZ0fOewzTOH8lnP0SaZGVL
i6bKWKhG9GGJTT1I+Ue9FVBVWomi/LQKF+2yRgOM4+wVvduWR3zkhdwGqHcU
5xBU+V2abFOtWv7TBh+X7YPY+Zo3YPFJ8+69oaicOgqvczJ5IC6nVNt1nDob
iSJwzqopH1KU6xQr9LKHrhdt7YN6y7KsyTNEZbvfTSkibZcE1jFoTq1xQmis
mYhv1IF/dfqUeakiVKX2UDmpEWKyrdBf+j9P1TBc7QxKUge16U093UeBuFfT
/zchhxKaDs2GLBSV43aByS8073G61/kcbSrGRytLkVnyV3+ynWVDGnqzljzB
gkbbnr7Z+Y1k5Fm6QgIRdWc7wKZLLXE+Ybu/aeMEnD+uCW4IdPqkRRll2q8N
PccloyMSu1ZZz87SfPLH6Zx7D10EudBxjEHjjKBs/VHz0wc8p1aIuQZyIeW3
hrea/J+8xQn8NLKX1j7f4YNbBFy8yn10iRQa8tkh+rrww2TcTePIz3WxtOXB
mERPAJ1IMSQLEMO9Lgm+tlnV4mkk7yYpmIt7VV1bbyQ67zEPj2KWsDvZ8sO+
fP8PngpCazTMIyM4vDqH1+y3dIrtP765aefFWGXz0Qec1TZ9wOFpY2XMBnwf
OyFdW7TQA++X1kXdFosKv3QDQ/6ZMzBraUSL6jciWo7EnsdJyn7guEMlGfFw
tazawsglYNtwt9Ox5r/5fIDmiw8z9H9SLKOPlBev9fn1Bl1p25GGBeYp+bXI
iycWoXmA0vCe7njPD2sarNbq5nbPpzoEX5JhzAA2d/CaClqDMf6GRRNluHuL
9zUVlOo2xdLeA4dOXWAhLF1qD0qBy6fEC2Jw7xLogiaEDUtu1q9731Hx02nY
q/N3s5SPF52sJ+OXO1pzOpNZE8zGHpoud7qLqqL2cssJhRSRn2eZ5VCOJlCU
oPb1yYP2+kGsv5BJvLh16FwEA9HRTkHbu4kdKbyStapnoCxPVoL3VTA/ReBi
gqAmtPOX+so1mtBC5aBzvngSDxH2JO1OmhEfzql0ukXIECb7vofKHOgeHb3U
oGrJ/4LwgwqsVH+dv6WC+ASYBFsbjhW/lMXp7J8ni30qeVvkADOHgiHXKwDj
aFHR7JbIwX+oHuPYKlvtz2DSXesAa+lNPKvyfgEmSYhZ5sAB2FmgRX+plmOz
78fR4W35TghI4MqbmZU6MPfyG2uB6X4qbafyPuCItMsq3+yQSGntBKb7o5FD
8fKYzA761ayOGFT7Hqt59S9GSmVQjUx/fiaO2zyigUZaN61QJDqzqj6qi2Mh
DA4OtiWSOZFaCk5SHFRBf7FcU5UgJ7S3IuWGi6kPCeS4/4WAtamX1SKKD1ii
VouMgy91bWtK1oP3nlu47El/XcU6Grx7n+pm5KH+qB999tY3kvL64WyiO3+z
LtpH66dw7HFCmRZkh25gwgYWBEbqixVwRXfHGH/QugCOFSKjYCj8gXCHwamR
1QQni4dlth6JGWIG3nPUFwyqmOkQps91j7+580sZS99PCJt/l6cBHFigUNAO
tNG/aRoG2xD95UioWhefoQV+le1cfGXeohHLqNMheg3hm4/bnhSHnTmPpt7g
lLoyx93NigbBT9HDVjS7aQ8kDdeA5T2lvYeUGgrw6jttfnt6qoFF+DAbBnWY
avXo54kYxJ3Kt2NB6Ghn3fqDwpXz2RYN5nZLT0j5fNrLCPvZVZ2KJUpXNZDT
8kK1eBcVS6hUERnr1KeaS/D4GGMEc5fZS2uaUUX7zewfhyz0+NWcuwWduJMo
qomQrnyUx0KNWZw8vu+mA+wxtF3tuy3xQxzSXwuI+8+rhbnf23YkXjcKYM1h
uJt3wcTjs7hr3LxUW99GyR4jzlJozYfAS9fShqH3Gp0gjBMKgRzeDElN3fE8
9zK/GF4qyCl/JXRnmUDchuWw6B81dxPLD7B9kCK9bmh+awwXiWsL8apk/cxy
+s/uYarguUS9aiKAHNzzHULoInR6E4qkZu52K/ZWGysNAW3C8H8CuiSR2vqe
beNZ5NpdmxYWRUGQn/CruUNlqK9meSgV0i0b+1b4rJjcZ4ScEEA8CZh6w5sx
8XmMSdSGCs/krJxgP/MdU/c5zEqxhnAYcwwNmGo+TDO2gg1NenRRy9OxQdNw
lEy3hFkmbTA2BYyH+Yr3sqb4M4Fa+g2XTLPLm5wbB7GqK0oh419VUZtx2Ho1
p1PrOdRkS15iC7EGu+LDjo9oneZEbI1PNM+I2Y16pOxip8MbPryWSy9CFFVY
BDL5bX4bJWdLyv1MtHSbI+V/1AX1OadiL0zrK9rWyxAARj3aqIQc05miONiA
f1XdnqBYTtEtReCSBn+ifx6/+ivpxA8sIWHYLjObo7bRyQdAzxgFty29oPr3
/pXZtU3CMm0U4bpr9Xh8th/chLFA3f/8WYQs5txtKG6trnolSXsjCOqb+1X/
DpjUvjn7LZxyaUTyPRBWVJGmkhtbfG9wS49RbEQ9nckbD5ffWr/f4iq/NwmH
LcMRTqpKn48CeGC7HsVP5PnfUBlIvpU5N9nJmEkYkzXZx6dRfMU7XIE630hT
zM96fFRFyi6/A60NrGy/H9DZ0IDts6pq7tyWIS35esU2/LE18RaKnytq2bEp
Vp0FUY+m+tVfBBdLw2vX0s3+502/aneoeKYAOVpZ+1A5ukaNCrZEeFzEIKN9
MbXZsYFWB6Hk5BfPigcKmlVRUsJZopFjkACTEk1PUqN3jEj0iII9Y06LNArY
2sCWkW+Dkb01gEP9ZXDy30xtMQqF0lyE1jlL5GqnGiNZZlIwHoLqG+keLy3I
pqxyYpFi+NBe16S+2BCeM51o+6UPRZJdvgtCR94y/sLInJNRGYWbSJ6Zqcxr
jdNhv/6YqVWEJnDqhaVCAzXjCdr0UOnSUkj7BQyPqOsRluEu7lHi/HvOmCjo
areP20Hhh/jWz9UemWpSI8Da2pu9oAosrx1BJZr0YPdr7MQggnZ8c3QM8iBJ
vlsPuDSWLTPCWK+WWdB9NzlvCxgZRAbZsNi76PeVbwFoMGqR9pYVF+pAb/J9
scWzsHOkFj9VyMv1NjMJ/V+JqZVu4hgJgiTYNdWCJntIXbiAOcGmg4h63Hoo
FVtjTKYzLCeutgWl8Xd1R8gxwemcKYSeUNlxcgxm9OgTcy8lKh7TuSpXKcuE
KndN+EHDqMvlDE0w8XNs0tX2ng0fpfVrwKNHdAmUxzwINVjsOKFZiJudz/+e
n2l8eMRd/hrzO+hefR/yVo3ijF2osSKaODCWKVs2hObF/1i5T4siaMTyS1LF
UX+rVPNL7AzMY6yHC6Tw18lhXGz2Fi2wXWUadAwrSxdez/Mw1HZm18/T1aV6
/qRUpuwjU+vk9HunKZk/9fkOfEPHfgfvAwgh7FRGLzox+s0fAqwIyIkoKWJf
3Kbsxu30LqjPbRJEg4zIDw0aPebo29opAjNBqF2PzIfySExa4POClNOhMxtc
XxX1tqdYP/SmokaQa1EzcS7N9iAnvO11136MHc+rYFFtUekKviGZ809aKOmv
5Dft/2+ZMdfv+7XpTijlBBUZOKFR9MzzsYIzL9k6MxUkKWsw/85MDr6VkSeq
9eQ5A/TcOB8CGYAVx17Ii7RmhxjNLV7bx7g7G2KdFDOm1/uZjBzbcBVGCLdu
GRJ6PpNCrH8X2MQ3aPJN4MGHrabUYUG3vBtXfJPe2iIXg3FJSw8N8rgrceIn
Z17MVxU/fpUgHBICo+BMft2WIepAShdkCN4TuANEsK+oVT/fN4Y3yp/QsMT8
mBMBuD4J6BVVETlfpZzPDGg70ph65Hj4mbrxSVFFjeSH6vClbQMEMAYfRZxS
21SZsuUHz6WheOzErunQSUugZLrEbEVoRbvPNYz5EAXzUpX/BpRz0E7Mj8rI
gWMgZ1qUxpTRLK0MqHINPc18T+AaBAnaByoD1VjJbh/Uacm/tiHFz7fAh8p2
KeMt/Q9S+HGSXda9+lYYlXR7IVUbsWxhCD5jxf9ged0AnKlACS4ddnNaE7bW
XRs8tUVJurCGr+sfFoxtmcm+DW4LpDIReaJbqShSelCK7ynGnNbbkzSwH/sd
Kb6CKWAiP6kW1eVAR2xR0vHhM00AhQiN7TytGt8AiL/RPlEJWhe5gELcCZIL
Ul+ZzadCciYitoA7VwcBw9ats0H4dp7si8Tt+ZduGPqU6HvSsAEbRAuwNdLY
eaFPuNx+EL4aiEbCBSmhBAr0r0Jg5pWFdMAqLkjknQYjom9Uc8Tg/C6Z2H0P
3ZogOZQt04X1S4QTqrzgf1W5vA22LerRIFueAA0GeO6yohNMx/uads99P4BL
YmuaOpv7npIQYQz8pgDPjk8hVNxe4/04Do9cR4+MrUZcdvbgMptd3YBpv3fT
gxtMMStXdxfRlYEt4Qgif2RnTZU7nlKT/Nq2JHWSDSMAQjXp2hnDySnotX2u
MBoM2perrIte5J53y7A+vrlJgGs7MV90waJn3e988DPNPZ/qQZyvWoyxKlN+
BYHWSxpE3P8qyGLsZRIQA3frV79Bwyc+YEVPtNGUKvNDoP2JLoYwhgpKplKj
lANvGclEsIHHmaA7S7HG6GVR3Cb9ZHH8xtN0uPzzqvdD4mXxNw7I8DBekYKR
R7orgx25jVlHO/n+5uJk/HjYeAzk7MKfKJZiNYZRQigvAN5SeYzc5akvNW5/
kOuj+UGR+0HksvDD9GcCBR5kPgGULkQgny9YGkNRIpkfYretZKOlZWc1m0vF
Es5CSefv+5rFs4ju9AZ06Brd8Mr4hWgnAE6g3u7R+arloFQVhVhp7HEl6CJl
wS2xaCPanxeO2wFF4e/O4JsEIwUPnvuEl5Iam6VXJQDoYxGRbabQwm3KMQsa
WJzhwyG7Zx9MQ/Wqi4qaq9wk6Z+5P7/DgkufDlnSlwXko8gkh6buIR4n0Ony
ldhBFP8VzFlTPJKN/wS+KmfCTfNs+lG2Eb7Zohh0Z0a1PENsIvSz8QyQqM3Q
khhzexE0ehZ4fCBHCfCz1qJOmd4dMEhDL7qQ5MW77hmHWPSrDPLxb3dL/cUo
GWYaoyJyxXLYLivlUWre1N5u7UnnR+n3LMQU7axDAVuj/EPkPw8znICwb7NJ
1C0Kvu7Q3t7gERvrU3rZLGQNYSWs3zPT1pY5dSm/H1C9i38txXaHbkBKMgSc
7irSl0rptoiNFToqs+kp5a9SzY/bRXVqeMoz5MY+vTVFQPboluF7H95aUJDw
SWcpNItQ3AuvRCL0Q1gESP4WveON9DfPGFXoH7s9VReGtj8X494utYLN/1hA
c3MnIP8TepNbOwejLKL1VaSKfWSZGbh0n6TFgJoXeH8MKwWAbxb7hAjb8AhX
iQBlTokRhu5tHKV+Zlw5AUkZuAe3LLT9VzhoYt898JVK2qEZuyJXbDL4MbuV
FjT/In6M85F9NLusc90gi2TLM80qLaZUt9ZXijY46w7XwV+gV9LRkawYUjTN
tiwrZ+VYDDqjr1NWpvXJ97qnNpUSF3p9BqE++Uhfe58IWT4oCPzt9dxgcaq2
3iCf9SKFhaNRvRyC6oTNbFubVtq6G1WgBCMicIeRygpdhTaRGqT4vK0WZRzc
NTZDCMPImitmpPKE4oy/7XrVfDiBvYoVovHPGAJzHFlwBBDa/MvJHbv3DRRi
XxqWeeuwddED5CHLDnuTEnxpw7/3CFjuwxgYDWjoT+2EpjI4X/Db2+jCGWAM
6hfHKbOJdKZqN3TarLwoKbvf3DMSh7fA8aZ4uk5s17HI4Do60qzRP6CBEEUZ
sIFZlr7YF+2bWa1qxEZpmuxHRf7NVQx4OgxeuY6cRb0UNTOm2ojHNvGw6KfM
6GOf34E++5gJjRp7PkQJ9kAB+TN0qn30kUOsb3U7FZCsqA4N80MKHAbqsd+Y
buczrdULs2u4l+vc3LJ40eepj3y4SJihtTK/zKf+gf7OrAAiu/md4qLk+8Sh
LeT+VRCpgUNKj/rx0uA9ZuMHjldFbrnr41qcDeqy1CYC1ldIJHpvau8/nIiz
jw/wkdDv0K5XLL4e2PNZZi/NCxNcDlhCoAnKGW+kRKVIK+pfZ+zjquXVpIjI
UTi9qG06ikN+shaNdxDjeLNNJDNFbYpkqb1amWFlhTS15RZ5lzFcuKiJ1n7s
CYgtb8+Q9f7uUMCjDEZIx9cEguv+hcy2T8wvlNSmRcmiGH0ZBP1xlQNz2K9Z
HAoswe45vwpYZNoXHMObPJkkmUoTVirSZQvVD638bk8Euu/MTOq+CraPlSon
zALDO8MQKrCp1M7r291gQ5tmaMDvLPIe7htHz9jn51NMFJkf4d0Uz/BV0JXz
68RWGF9NzKytzOIOOrvhRDFe081oPnS25YC6vvLw4zYDlFRN2KGrDJynFOOC
diy7ilB1EdtdBXmwsuE2g6LYyQhRzJUxNGxkf++w6l9SVbvj11Ni8Cxxvem+
HSWjgFgSAJ9SnZLOOX/ikcZQ+aPO3pi8JYpOfr+6/Kr56jM8adfCI6n+cd5G
yE1KgFdhyUXyTZLEC1edrNbOP1PeZQ67Sau/nqeBbdG9FHLvnvk8LNvuNYsp
OoUXtGarHNYbEqfhbamuyfuclCud1DczIEKNkQoUc4avB9E7uPKwqy6kxsaP
mj1reGD4cej6TqzYsz8z2aqE8Kqttn0rVrxVo728oGmJTV5wGOF4kfrjZA87
ZIw4mEZya1WZpp0gEb6KC7QVDGxXpSpv0q0+ivl4EYJ2zBkkyv73Ll4U+RNu
W2kEHXO/Ca0IVJvFK/cgISGWlYaWH+Kr6dDtN6St6ZmF+Fm881V8hww4xCcP
QsE698PfbQjZ2CYLSeqH4f4qDjK+6Qjt/9DTJzaM9nGGITyPnzAu4YTh6CBi
mT+yGEZ+bcAPW5yoUcx3ZqSVe6lVFJ1/AWwzP9y0sAwcm8KiebrThb/qzmKa
2jwkQX+xGrtPGaviddbab3TtdvaEctpPR2yv01EqYaDkEroXjV3NhgWr+W1Y
CMCrOjh4luTao0fULarsviY3gAzJgEQuyaodLd+kVAQb13rIPM8jMLG9I4ne
3smBtmWjlRDhhXXq2sGBcU5V211JM4DZ4Zco02Xf28nBdN1cpFN3mSdqmmRR
0mYfvHpXIZkvH02OsKVV1/F+F+DoxSeEeNgG8Z4JeMU3aiSA1kmk42qh3+oC
J8sAYY2M7FPPXyOAnZVvpbQaHrP5ikqmE8Pn27wFY79DXs/ti1HCtyi861X/
bzIFRdx4dnS/3K6T0A1JiC+ij5ChxKb2bEMHBS27EQ0n8C0DCsctvYxNdwbJ
EvwlxJS9DPpGZlz1NHq/1bdWO70zEzvHzD21w/74mFM7CPOo8V8nDukX1j38
YwmNVQCGglce5W8I//pGByA8Et1qTZmsfNF4KtyWPQYtfsy8Ms8Z9xB87/Sk
U47+4hhCaNdom+hPP42bVn14qnd4IvrvM3vwd0bE4VywIqCpISRYb/HDhL3a
FaThDUrK5MfKl+ec90m3Jqmo5owOZVhLriRAycFqh6rpkYlpmdZgAyuujNQD
Kaf5hdy41TwG9+M8yDCjxxFnmYfpnu7vrlWq7X4lcmMpBqqizweKFXaXdAqq
s4yO84DgSf5xhTD3kaoeuR3yKr2qf/AQgpxI8ISKt73Hu/nTJcAlSdWnjLf/
+ZDap8grFjOB4RlOD6ByKawIASeDBBAAiAQaO97uSnJUTh8eCZ7rWNWJEcfy
G7sEFcEVdLpcW2LNYBRq7tjuLlRHkzU/tgA87kxzWTm4g5q/+RMyfB/1M5wg
Fp8joDhA7QmTbcpckdVytJ7TOm2MTQ4y1D8TuT/f8HYaUejvMzZv/cgkRjXE
7T1JgzpVPH8nyv5DaK7Pv4ory4Q3e3oy19Lyzi1Fg48CBHo5Au653+3ByFjf
q8n2FGTnWhCAZoV4YZ/+YqvlIMawtqNWOClRDdLGuRhcl5Y21INdwiTknbaI
m6fCbfUYcEpA0FRZHjWWPzecP9f9/fCxwnBs5uKwWEJfveQV4l89oOzAl9eY
hH020UaPYPDcVYf9VJEvekL4oZD+RX17jWRkjOSz4mtPbKVZ9EOrk/wA5KdU
UpQNWIbZW6VdhLd2qkw84n1H2BxP4z+87UloXy8xSdxiiX2YU737y6GH4ayg
8Ccwp2VeT97cP2OcWYfVi5eMLErTTs+KKI4OarPyDFHA/OSXnDXcvM30A7Lc
L4dtw9pKPXPQLj5DmvvC89gSwk4JDfhsa5noraC/1YSmWezRGGrkG3CsnO23
lCbCjuuGcneGJFBELQNQM5DrEIWnj5qPTECUL5Tu2BxYKTQB7YpB0YEzr7Se
XXRePuN5ikyk+iUstbKvwjoAv4mGiirE/uAWoMG3z8kDhsgAHnGJMVbDlZH6
evqY1kNO7edoVTT4KxszRvzwu/bso1RJguD8G/u8unz9oGcw1pRr4XLNp9W/
T7zGHMCV4wyyCLcNJr8Ttc1F+eokYCJFMdcFQh5KHxS052wHjr1pWLpgTj/y
p+PbjQ2TZKX8NRfGvOFu5JY9BCva9IQDv4Snoz9QlgZZLxKEG5wCRsE44E0q
No0b257Bbl4jZhgcJqlRnFtP3fdWldpc/UX9fMrkZEcuEKjxeQYl1xjAh2p/
8MoAcrjtEHh1m9MO3jqtRchFm7bK8gVrZJQz2iPOuwd8vtrl428kpPiFfYZ5
7gpZ6XcOP/k60pVIt61c4rO79GFCWxkrpAPDTkJquQ5rAY6GlB17SdAA6dmF
SAr5FRCOE4YJ/PGYZ1xv6KMVeDrWeW/5UWteUcrUd6gs2/oxhDAsGFCN0HI0
MoCn8iFWP8EMktwLRRtxJqs56QMDZUcQGLohZ1/zkbcigGZC27DVDiAuCfGT
iyKFLHECkcf+ujR5jJ5e4wISIQj8v4a9bwBLbXeQrUxFQ9UYSsKzblSFHwZx
AA6nyt6kTla7j82Md+5ruBXmBO7LptxYUWU3l9LmWFNCmMdFTuyFacNyuLk1
lXAg73Y+a3c0M1tSVFSxYJhh3fCRrvwxKy7/DbF+Md9pINTZoQ7VzW4wIUoP
v1948BEHJI4zLS11WKb9YlMD+VP0M478H0botd88Lhm86BCmZnuzgLSmr7jt
YO6o06KwNVpfRciRM3zQEqb2VvqWfMPWjTCriy7weTLThDTFZ6Rwnx1rC13z
snmcOl3CJRkR2q1b1iKTg6qNzeKxKDNUFnTy/mnP9CGHZ5Fj4JKZ0RGAVk0R
RC9FCf1XhNIsbi1jLctl/JdmXngkhjVydAfdwYjtG3qJWp1uLebNSZCR/2eH
6qxz0IEz0SAgmKJF+C1RUYO52GeydUzitrI+Arr6dPIqrnz+muBnE3+IJVu4
HfbiaYX6egKiss8InWRhvN1sHq5wxislh0YQEgrKGBV3fz7+Gj+cP4wjN/Bw
E3h7L3W+w4V6SzVM0AJSc6FPbTUgMBaIZL2lcb6JYASwhXK7edeCxi9AcX+o
NldiT9qjPuD5M4l7gbGaSpqvfUiHSqRozt90CrxVYhsnJIFZ+8AeDrrn18Wi
LVRn/S1dkk86QF5w0a+arIGHwEOZ5l3qAF9Aa2nTbB/5Yt8HF4Jtir5YAXko
QP7uABSqyAndt9rP5WFVbmnAWX+7S9875YleMKFFsZxfUzNTTtkV4TnWRtJJ
ireHJoqfPWjDFn2f5r5lpGCDVVWk4tEpethOAtirlMTpO2gwDIltqoBKC3Rq
oj88ElLfGakLGmC15Cxx3/np8om1waCAvxEOaCNI7RM7pQOV/kpk5scp+6ST
dOsCw2DqgT6f8sZYV3kaVh9eOvwZ5CzTlUT0Dep4kez/XqV41UcDzEqmLONQ
nWqR0vtZ/w+c6DGJHUwsm0mnuGiR5hMH0FDPwcZblpNfN9+ZbofkGzRT2rM2
6lqBm8csVJHPcwqQmElcFBQXDvh8xSNXOOsKH4ybEvf2JRyXnh2duQmWtWWh
i37DdK12VLAjAeSeuAJqHZhkrTBTYi/Yb7UvB4T33xrc6nIouoVYrk+t2u5z
hrmZ17Cdm7lAbYKARmWkbi3odDYBF+uG1JPV/Q33TO8SuFQ1C3z7aFpKFmf/
gthm23lHgJxVwyfi4pAGNEMm+rouNDNwbm5P9WrqHcB/cvecKbmWfxZ0uZyp
3jxaRW3gnxBrYC0s4kgNjoDLET+PFh3rW8FVHVNnTYSg5dY0RLPA8uyT5GSb
VZn265gSE0amVdGrZ3TGEHgnM645V1w77GOrS5ta25/256VY+cIl8mVXpqAS
uzCm+K0MTx7AIXUrp5V00jNiDvaGh5C/CKyRiALawcfnzfwqEsrcnMnGlMnK
GBBVoBz/wl5DgxVJIRDBzPIQJFawTt8HdygsZFnCyJzNWrDvBWtvqthEH7ID
JZAE5fEP7rEQUfcfbbPZLGCCDVDk4nbeEMHgsJfqig5VQXnvqqhYtvnFMMKw
9Pvb+Rb4uOM1TmySdUgc/GRmsLFAFk7qTlc8R12TJr0EpoKqAD7C7CCnM4vn
rUs33EBxUrXdTrizWh6b0N1+rZ9xxh9xwtvo6IJ5FYFtHaNGTnoGQ6mqz4bm
yjSkru3dMAbuAAz+sA5Q1y54jEWJ9pRjjNkQ0t9VPw5YXEMmU5vVATdGGaaz
w56OYArAreJxEIwU3bnPnMC7QQ0HZDKbU36bJd3mR/4B4csMFjOTQXwity1n
tkHu5WrA7s/z742EQZQZsfknWMvjF4eOn2sjoG6SNK/tZGzf7BWQKPI/sy/0
vJ4JA1SHAfRmd5e/IsWka7KmaOJUjQeSoWNQH7iMhQxCd41kGRb+AgtjY59H
1BpLFQlrBxukpafrsWmLGkSaRUtiu2Qy659WK7YlqGWXurJCf6EuE2jRdGVs
6+F1AhUOOzLdOhzo0vJMOyPDjLv9wjEdELBylomPRs0RBV26XQrEmA7wRz60
wLPr1iOudVmo7xRthy8eVGvw2ZA+7XAT53662sciX+BvZZzqCNNgcUHsLiOK
EFlpxzJe6TBCWEqhS9Jjh7iYTUrfBA34MYy0wK1C84v5f18Hc6icabtM6UcC
9rszMzYLFZm/T9Vpf0DM6wAy/FuVQ57nJe0Dkl90toIhD5MFzJyxP1JN+U3n
7DfQGnjtMtP0yHKvHmSHQLoiYfaEg+HxmKAsQcZaep+9nQegUbnMevIUBpha
Pmn29HziQxCFtdgMYZKnVgAYrq688YD+xKtLVqkKivuwkrhkyU6Xbn/dpJdl
8xpSUt/XfLfUE8unGP2sXoRcvCyNIfsT0okXrCOVPWJ7ff51k6vU2J0LkWoT
RXdcgAB/Cw6X54sDYTQTtmTVkMCKhjpcMBB/Agv1N8Y+zxvucHFLl6ws/MEM
rq4xLE3kI7L8G/GPBeG2z8rruMRa6RNKzCt8NbuQmpLjoEix2Ya9NOQFkW7A
X7nIeucFPJYqRAS526cfQGcguVuNUbNDnURLE47UzSUTq2GOHdmk//BZJfU/
HveetXR3oBJomWTOWepoBVOqWhoawhqz+vkQxgSfaNq78hktNDPbxXEb0EuP
e0MzJNAAZ1vss3DmUi6WClpRogX+1oji8vBAhZPosLZWgZABvLPCclI4t1hb
C2u/kU0b7te18aE/58Wkxp/SMJRmPPyVdpk8lrreyYQs9obpWdlRxDHbXOB8
l+mvRAF6ESBlHQpv3SvMQRXELrVrwlNVpAyLZ3DsIcbQBrjgWPiV5Nkr3UXr
kT88YddHDfI5KZFlqF9iNS32XDIffKFxQrEr/Z+H2ujtEtV43F4Tuc4aTU8G
yxcX4ahgJx5iEFCLmjOMAV5IVYabLyQQEXvmvRU+KbDTi2qMNt0MZaO6QI4T
RnYadELS7Ta2oXCuBjAQ/12O6B6g2YUZ1wmqlHPuWzMorofLfnpnT9ukq0qX
3TcaHxZCj/l/grEfWo6zXL7TWyrOxXcvKKOyCUEDmRxNE3hsgM8LVdWhblfm
4723SLz3SQ1nyyM9Rmqc+RzimZy5WtIQyKW6dLYTopXCQYIw2Ssl0FJpVuyI
SlxaH3CZiIdGKFoMkXHyrZuMsPD4ksKcdJFBGFsrIsgmRw5pgZtOfR9Mq8ih
JabSfp8IsdNuA5ZcO/SrDJZWNPBpzA7RHILHHzV6hFnjr4P6fhdd9Azg9Kdz
+DNws7CbmhOiCrVU8B70iztfQnxN4MeB3FllIYzKZ5p0Jogx2qNfnDfqBG6i
SGRtZVv5hvSjTjKPWyzgCdxiIVBOyIhzoCqRJ5vl10ZSCB7G7/zO1hGfUp3K
DL7eKtXaqgwaBaz5V3MvCDjwsBzdwIFdQN1SbiMrn2jEjI/cWG73U1ZsTVAG
l/YNZOwAEYyp0nyeFqO6aNU9sNPuLkN+Z4iolJD0UJo0YefOog4dWEf9Wav0
cjSaMGt5z0u2XyyYYUjofPHEDLPIe77d/CLifLvRYYgACOdqH2aCShfzC2ks
GxaN0RHiav3GLwV0CO3HkZQpEb8WJqnpaPs6e5p9vwtL2lvz/w+mM/y+fQ6U
KKh+5vytShk46Lc93on+tQ/V9o4/ZbDmEyZ3COejqQK9ISQtogFzkqNSJPD2
+NccnWiFcWg7HYqOzd5b7F94jm3LyUSR2zroPTs15QnuUU0Cb0ijOy0HB/1I
IcEeVEHuOUnF7QtpDJl2sDeeO7JvaLZs9BMVutf9+EAtEx5LpVGLSxShBDaS
xcja47FhI0HXB4DxUbPQ/3ocL+/ewpm/9UFNDMAXwyEKXkXHS9s6InIYq4hY
Es80uRXVHNpf7obfenQcrBgZ+nr00CFLw5Mvzqcamjcs2vlUVTqz/n+wY4hL
26Uug/3X3K8Rz8OcarLUqTmWsShVRLofL2OYq77cRRZNl+YG3JUg5B3dph3r
oi22+hANfmrCEWUoOg0Xyzqj3wDMCnubIXnp5N13RyWiB3fPMCmydgwXsSPi
u8jHavYIoRbfDc+CSNuf62er8U1IPWawyam4b+3NIt7gaDGJtx8Ed1v57X02
qeeWFDY5yA7ovNSIc2MXXSCBHR9hNnoffMUingw4a2A6P+YHW9cTGVU+jY+b
oqeDkRScGaF97TM+T4gBE/DndQibnotInaudOnm0pTaNnZDf0/gsukZd59MW
jHkCY7y9J5u3X6537HTeZs1c3aG6GUlOgRKk4tLSxR+Pzi6PDEZ6Js9Cei5c
zOH732cXa4Et3m9epd9ZrtTXE75emoqCkwL8VagHWY+rma1n2nwoVG8f5jSE
rKA60DUoytx11ncylrL9B5OJ5pn890BOkJqHLs2A+8SoXhHwM3JQOyd4lY3j
FubFxmIxe5dE63OopH0tvR7gCn2qllnGzGSGSHaAiJJc62mIFVbAlj36J3AS
Ic5JKiXdU4IE00QUb0irEhL3M4B5O0dm+oZnPuaPM+zaTTdixm7439bR7s0A
bWHsx1Nvd5dCA2dB7Tj0XF1KfksKQsz/27UTjgJvw+gJqCyJfP1tarPpZFs0
qS36UWXrEdylTfUyywqYAx35JtpawcMUdIxHTroKDtK/rJF1ia1H44krbEST
PvjFKAlMgteKeuhEOnYunBjVwqfFJvRgBE4d8roBsx47p0oMtSC/mswE6z19
HZQ9HOprs+z0c955uy/6/7lh+tEJ3UycpPsdlQ31uiVdwRV9OA0461sppdg4
exGEW2kP34EA51BMFl4fMIWjAWz5NO67DERxp5jyd96r6M5465q0dJG1u8vj
XmtI12nogdj5LwRLrgUGcFAYGQKeMrZVVwigsQu6JRCnY1+hzSBlVaekRLKN
Gk0WJMIIVAWHJ5v6VffbyotRcd2JIqVNLXbWpmc1m7fgfB7OQ7bmh7EWWsqo
EXXI/udx5l548JaBiVOv+k60jaWpID0Km6fNIRfirZheRZCcxla5q6EMEjW2
Lky83gtJEkl+3RxN9ZPXU0Vi3Ob2w/TVTgLlJg9IarPgofIyWt5PIMeCXBpJ
SyPVJszIteRQdDp/reXvKLInoDzOIMXB3sJzwRigQW+/64TGwG9VWS7hcmpw
Bt6ISRQvLEPdthMmfIQMfvADIImy9DXH3MQ/RDy+kj7amNQGb7kZsYSJtxqO
/fXj/VTvYjt9KHUUVpb1r5tqYDWEOR8l59zbujo3BAwnwyecX+aFxLouwFEm
xtX3LLX1XQxGiEmIk4hrSVOWZ5Qqt9BqeR1snw+VWIRMpRgyKzHvX5HF1jwZ
UaWcKbBRsj+dPId311+8WtI8mZA8F29qspUIZBECA+Q9o1S5ZEVuyjB34aTZ
LYlf0u+/ZmcEZu5AmItIUBMi2oJ9rp5hNIlpFWW5IhpoCZ3DsjWyJoeHB8fO
09XkMk3K2yIEsYrAomJjkn7Lv7b6iOZbkJ6Y3JmG59puo4q5CffYZZeP6XES
WeEp4jXM733udx7KNlP76yzBpXp1FQHCa6iY8BxBp/gdwvUmm3sdP5B1Yf5N
+cC3ansIKYYNGch+MBBUlNADqh7+MMxg3zKmvAT5QFU+6xnqlFfO2XizSYqI
9VSAiXbk8xM85Fblyin+gxD2hajjJTX1/MkFBFlYEASS0WNzZ/dPD9lXFp7T
YLCXaFBrkYO/I/YyN/M/QHM7UqjR+IE1H9anTtc0bGCTsMWTxbnwWeM5vss/
LPqVUEdrTioF8mUsQR2hfuVqWFGddXDmJhzSduZj3xIzZCSPQrRg2XM91VDi
2/nCYJedgqJdtr19mhKRrqlMc1ZvA+iFe4ZntIgSOyxFw7cuTcfctyereKyZ
20V4jKCGl3gjgCkUEswqp3gpbjtHFcq8exWcvrouCvcx9fAK59yPDpVFpAtk
9wUCBor+AW9d+HWsNKTuVZAcXUdF94bZ0fu4pWz1IIXFKxxqcx3r6wz2yLAK
7O6DGhIkTFbrwINHE6ihEqlMw+elHHBBj0N4ar3YfElJH/c9pWBqZqIhmmas
ys/e37cZXMjBzzhkOPfriweEPy2P3R4hBVUmLxIj+pAh0B4OYwVKeUdWvZgO
C7tbjtlwaQmPWbspnSUAslHTZ3MEuD+OSt2nBsM/fzdsZZ70liY5k85zf0ND
72OUZ6UV/AIqjruHuEpu9q8MoW3S9yXQo3oFiP5QXeguo7WVDXwfs/Tz088m
V597j/NytE6fDsXjEQTu2VAKEE6m53s4nN/HhvB1uiiJx39Uq8NYVPqYON0D
pyZ5CFK0gj+r7Mdy9qQQW3QUqpAz6ABdnOsLJvKa5EzTYI3Z5D3fFaycJWvu
vlGl8aUQ8jW9HC5pgT6p450DVG6ECWJWqfmnyJGfufOZFM60IV8rDZm5KnCE
Na1ae9X8XQTpC2YnV4E3GnbLZ5bmzm5KlM3EvLAaojFjTPe82s4d+NKvXSTO
wts7kaVF790mU7FWRk3EeGCnINln7XazTJDPGIMlxhNmThvmVAXiu5H1J6ZE
Wz3rkPPx3Rn29Z3wfaPwHoyj2ZXGFjSRur3atG9sMxGTW0y/ZYGrk8HktKyl
VKL/BLSDC0zcAhtipsWBoO6evpdfItkFjHJKiX/CDpOXC6q/S6tDRKBLUE1D
+pGH5VVY2yi5W/oW5SnESLGGGwuISvmVHu6US4pJwlhFhg2M9pq1je7TTnur
lZJ1fMCHnRbtPqY0+lYVetf+Gq1EPZJQ5kXGpfWNmoqfY7O03ilNGtPpX4we
UscGQsk7mrQtV/QImjEIeO4MLVyDtMCwk2nS+Z96MVz5M+sWJQtQVEV7lROn
vB891syy+saDffU6ug1STfoMSAEh3ajwdsAzKZVSHu0wfX2HSOO0/DudxihD
cX2vlVjspkeIprboQ6ovREeZSbdXKkmJLj7mSy5nJuWJpA8/E5aw6Hev6JAf
zJ0xvLRONFhuF0wM/92tzsP5zsv9eJ4irHxBunksWiocMxIkYFgGWqF9Djjz
KkB1qKa5GssjU5O5tvgNu47NlR8KoVTq3GP9AlNjzaJWqovlBRVD83xDEDeO
+jN/kY4HCUQo0udUvbxsddbGmuQJSpGnHJ+jW24qSNQNlTPGHrxErcCDCzsC
izp63P7ksFVj0ENLFG/BtsSmLGTh43HIc5R1kBpE20OI2DLRNcNwqBXimyWp
vk+0xeBUJVrFvL/tupIGhB/o/qFc3ZTXW3WSnshZwTsglLu1mLhWsy8LHEio
jPJRxiYQ0vKGvjsaV4331dGkZvCaD/APeHEkdC5pmvfGxRtby1sj4OGTfjZA
e0zTLUAaxnJL9ghnDRBlYeEeI7juDUurEjpGhlkVnof+lz4mfYpM3KUr8eF5
XXgeFGNJd0tGGH5pUYlMPTrYvcFU2djlYYjGhop/CFsqLajgTxsgeo6hMm/B
Ip/0HMeOKtX0WOxmwiLzz1DXUkXDGddcdVJ2P9RMaeJp2loLqn43bMNoCUXS
ziL9wfOcyVeLTNKIqoZrzOdZljS2EAkXH2+MyxrLEnG2oQ96DGPljgOhCMij
Ac2Sk38KUo44xTR1VnwMChbDymIxPbQUWcx7MaRttoe7MmdB0VZDcN1MQSlF
dZwrFj2MnJ0IYylyecDWEz8r91QQq40EBMEfDYCvdc68RPqdCV4dJBp9JK+r
s5gOTSvOr/sBB0PcjrYw7VgYs8PNkrrLETwSYpe28PgwSE82epKVoB60DdkW
BOO7uFoNB2CtkevqXndH5XHgJzNSl82Jiwpp5ReYR+BkdNDUJiIuZgQn2AW3
mIJZOKTWI2S5ikn1vFEmdiKW9W3rCXIGrYsJMzcui/bVxMt3agtkB3Plndq7
efXY4aSdbBDGrDpZYzfMsyQhKCqGGd/adDTGzTJaToio0rp/UBj7os3MaMsP
1STlNvu4irCRZnfhGfPvb8PD9CzBGjbX746/tONrpJTOUYYD+7H8/H7maiuv
OCDtERWZbU1rYKvQq/pRddfBigRV3GUFEaHiaGm90jtJ5RPde2FqIznmjykW
+T/y9DLwQbj258Lv2b/5PEZXjET1vOZmrnjZfPuM/xPcjPdV6gI6BFeH7xo5
F4e4Vxlwh2pRlN1gS7qKtVfCuVPD8o8uzT7owOK1YZKwQWV/Zvej0vCHXW7a
u9TP+h0TQuRBa3qNr5+zHI2ret/gvloufpeyLw1gGwJtVP2qZSllOopaegEl
sTyBg0rJ3ehOG+j952lN4/Rj490DnsJGkcxjV2JIRL6JVksXLimlME3/2G4O
TpXto7NZc3lcT0rYFNMEvZ+pjj6gjQjbgc2h6F22fhGgXVp7tl9/ArQQqD+Q
kpT5DmHnMaZn58Ld8c8f2cYjBpLNtzSbZ50N17YmYC1DDJP/SDW9E3e9Nis0
hF3gVoMrXsuaidpHAzgAyRopqdooZiT0y2So364rvNlnU4MRbQx0tzvTvnaY
bTaq3N6sDeqpTZHtsoHyqN2UfUWHWkl2fdN2MCCcOibBd2abb2DKWbXz32uI
1oB9JGpEAFHkseU182FSvci7RTctCKU5vJvpw2wHuWc+FZRzd8Vt4ZdvPg7L
3WZCWossoW/e66pGg7aNPFe6v30T2GACUVh617pHBI2vrZ1+WhE3c/CbGgJ6
yZEdGafKNAVMp6t79twvKIDa0sTaJD6pql5KuuJpkYYvx9u845x8g7SlYrQy
Tp27G2qqFTiodVE8csJafvYIqlfEDxD11XCDvrLbADElDoLQHL2L8kE57Nkd
Ri60LFTUIsS+Vrv2I6EAYJoakwGvkZ3uFjr7r//G4O5tU6cKThT4EXwf7zvS
LMO7g9ZKEr7ZCAuHmj0nqiiVrfdRRX8RnmmGYoJ+KE+8AFkCLyuJe8pQ0v3M
m/ssMRGu+WOBebxKw3K1SUqy2dsrBVu/1NH/2xepDgoGs+Ncec0evcMMJozo
RZrnVy/WDwOyLkNwkFTXgXq1DrClYY/oRoddmyB22f6EkavPSTvzjC9ezmO/
4oQiKsW2t0fOUuqvndd3u+f9pG6Z8f8yza+lDiRbEp9n4+roS2ZFdTreNQDv
IQRBOKmvKkSv+xKFt1loiKgxAOL2lwwe7yyQt4j9NNLwd3QIRXkvAuP2wvA+
YhQrWwLh/KdDXJ/4oQ++3vO/jhGEUHg1w4YnB4fgv5Y105fgqOakxySwExYu
lXECeWfEDz5orTjHfoUaGcbpk85UkS7O9iHB21IjxUT7bR/Q4MGyWzGB4PHK
OE1UeZbWuHMMzZFB+Z+At94Dl0HSqZxlA0zsf1n5lECus54D6sbX7L6af2Tv
fKEHSxdECW9QGR5jZTamnJrtmu1yERrvPGfF5DV3abhdrw31lRTb5tCHW3nY
VhWwkaXMTWBbPDxj5VUqQ4xs2468+/Wsxe2yW4P/6tTryS4NFSocA/YuAQy1
S2zWkmvhTgClZJgS+XmvTJHv+Hflz0yPeTgCbOLWn8pxo9RH2K60uaIASBOh
rTLOiA9ENCSeNLjROvtYXbdfKaVKsVILiCgNevQZkXRhrda66W5cDhctJUlJ
n/uUIpDfV3zpv6nGCR9v9KUmGZxKkePS6AuX6gSK81QsNUORNu3K6kA6MdP6
Z6qLpD5XfvEBpeGQApECl1TrnWf8in1t03XGPa2+AXb7nw0BZYRGv0AvfqaZ
gKfw7i61PBdG2ZtoiSmAMJQow+krTfcFWsRcohNX0URT01YspuZJpX0VyePp
rJoceheVLtNPl5idN9oaW1bJkeM5ELYXQ2hGcRqfyMADOW+S05Kd3FzLu1Oi
cM1CRU8fi3xCsTE65j2zhHVYgcIs2LT33Xq40wq7sMl49yp4xfC5pj4+OhLF
S5dMushfJSfRfM8Wrzpt/qoIY3Gs8k5JlLggEEbizdMfvkCjz6u4b4+15hGZ
KFO9XA9cby/p5mBfyP+5ubB49TIiNtbPps5fH5SD7sHeQ5OUILq7bV+z1tKD
a65WbWJ+IbHUYKJUwOlKkG17Q3NUgmmggeRvxUYWxqSlh9YOSwefSMAvIQHs
I+iW7Usk1hbx6fIktHJAgysBI8SUUYSnP2okXEL/m+Beg9n5wD/aoBj8t+ny
QdaXIEUtu5o4yahyXB6czw194338IOMl/quR590bDyOUD7LxJziqn6tFt904
shKcVOdoZHSt/f9tNvQHDaGPdRFadX3Oml2uY3H/vxxKmsk62bFleiQZw1f2
26HmjtWCE1W+B0i+fRo8IzU6e7hW8rBKn6iuYUKOpiWqQDncXPdMTayzb7uA
5kE/yqFXV63AoLOFB75sjis6321Ahlaj8fgKWcthIHVpapgLYo5bQZ5dr2JV
2n6qOx7BNmqV7uJlD9kHp/sv2WE0+079KIFvMiCLqw01CLwEXD4pSC3VS7RC
oqa65r5SFgXijIW2onF9KJ2jEKeEOyi/KxMRu5xklD2PsEWzXwjII0cqpkIH
64+dts/4LHBmFvjHlPL5ep4mu5gPE5v1fc5fUB/9IWSWQN+CGB10MYuy3CO7
yNI2eVA2gOB3KXOLmbciqOQXBMmE0ri9VW4pu+OVqzaUu54HgDbH3T6TF2aH
4Z1d/gwM0Bc8ITDI/NnEVP90Z/CCeaaEco9zoH0VZ/NNlisJpeXw+HcS1ATk
Ec82GVbyj+hgjhfnseHRzORS5btmEDDIlw0mz5PyM7vPl2l4J0E54Hdcm4t9
nl5hkXZl4P3GKj4UaAERaoZBzXucmcbb97hG8FscLqQFgZbqNSdY3gQlsTfw
+Lj4xnxiYYlBsFSZYexbYdYPBhhpQdodBhz6yEo9SKq84oNSqioBHUqZK2N2
YVxGbIRz+NhNBOLDTt4F+CxvY88nkINGPgw698oZ3QJyN67zKP6QUju/OSMz
hzgpaVH9enP6NWG+az9C/PX/Z+IuvJrWjzfedYlZojSoAhfSJ0W2NacaLZQz
ZC5Gv6B/0tyNNA9adQEkGu4JzGHl24ZZ6tfKb+4/6eoWVIqMpZH/eJ489Zyd
FEtPOOu4RfM7z53IU+zfebn5BRyvLG/0lrTYtuLFaV5cP2sCSNLC5lv12hdQ
jYjkWzXYYZFK7jGGPWf8G3u5agZlYtZvyoFmA5V00oVefXhAksBrtdls/oBV
L/8nzQZ9enSC4S24mlxTt32iBy3Aa+znmY56Pb+ys72xNpyM+j6fpTU/rBBm
83vbETTftRl8Ug3aCXe3I61KGN2W30kkqn7CDKGLLzFNyFdsxETpKnvsf1af
jSVi2eft3krhutOUbVs3VF/3VXvxc4JAtfP4a/N4WtPmB8/UR4Evoci1aAL4
XJoU5AhjajOXQSw/jVv5iMqzrgFec/hHUS0pGCrurYBvjZRraNy1DrGS0kaF
ZKvHOhQmYX2BwJZjuiJzpmC0Hsp24XMC/6gtIh09U0OIajM8jtDA0ZxtuArN
CAvVAkY3/0E8JEMhzqn8njY9OWA8rIdPnHxk3H/B35ZsfS+SImpwve8Xlq7z
eY5bQuphCnMwpj4uW2D0e4hOldUIvTMPhpaI/RXXXgm+hqWa0ggJPxpBA37D
BQqeQGOSvxGyN9cYCu7WD7qD8a2VR87lKoRgVPHDfKxCI2mwfPMOTSzd9srv
1v8P7R7kMbh6AzLmxQF2XM4FSR8OTELSGyIwH9JXslPFfII6aAHC9GWVrg68
W6EEmFgsxnqUe7DztpIyVeQUa6FM5PrqQz0a+tIm+qvua/yGytrW8mjJrPgf
3t0H8qY8eB+80joWV0dWgMcTYxp9ZV+uOewljtDnt6z8PXgjreAdQ3Yqdc84
foo7CKy3m7dQfsT5/bW+sbp8KAsbjoJo0ot2xKJLQadAFi0XdVOaBGOcZ7JE
iSadMNC2oNUpnkO95MI/9mkVOmTPlv3s95hGK4XNxstrY7Fwcm8Nv7gGsUP7
od9gmhiDhIR5yThKhSZckffyIrntZawzLMgXHwdIL1FICAZAS45KI1f54x4G
t0PYwBRe4++DYc+CFzdFRsomiQHx11uJZUSjKYGA3NwsAXRMV7Uu6PcO845r
I26IFE/LbEFYH25bCbCEgeqdxWIlKKeiN1EU/v+beUQecW7Xl2K1ipsINLQC
OCAg5nd6HXHZbJym6yy5+rkiB2eaVAXCgi/yw1xrQAakHNix27p6x4Bz9a0S
7JGU/JOWCK1Z9cwAMCSqQOHBQkdC8rl59Z1g/CGn6Axe11FYhUHBUOFpLlLS
Ep/lu8CGio/XzkztMaRFc+J0FJ4pj81efsSpfilh/5s/pz17KmNqvi4ylT2U
dZBMTdbvjGaQJK7WNufsOzzInmMuobYLSQ300O59ZwgGPLx5jjuu1iKmbana
0k+5QyCHmmIFNvSSUDtOFx6mGAbNMl974UxG9SHB5qAgZ95xYI4esibgKCPz
77w6qN7cg1o/6DzCjC0vJX+6u6WATwYkcKvsmP0Jz48M1mZW/WX2xL/ehfHe
umStIHUJgethRdpfJ98dcyfSxn5FB1Cm46SkBoCk7dDuckARZvuWWjhkIkdS
pGRf/p9lnv4TuESZKTAAguleuy91StqzubyQlerQbBGcSFsdLu/6mJKsaTuZ
N8JVUzR534CAyDyCSAyAb+5ZNuP4hMRt73mBwgVKNa8EBehijGtmNXQ/8t5l
jschOuZt8i9TtHrvQ1B5Mf3zcbHMwAsXkXbZnKoaw7k/UEIPGzu44pwcLX4n
ZHV41ikll9dYGsGfROoWg9+aZp695Ub86l08Dv4Bp1WG1XrtteyZwNZzQ2V4
HRviF+ql0cmdjtMQeVYsO5yz5iAYQhwjHkzvJE3r+hBdHXSmzLJSzufoXtzx
L/EznxTAUebqVOoN1rsrXpD7l/on6S2jbrD8tkUPgQhaUhK+J1ybM2zJZyj/
iIT9g6nCfwWolOk6jjKkD04XwXbbgspkgzUvzW3n8LGKtDoQxz9uk+q/wk/P
o/xVXMr4F8CIvGsVcawBdGC5/Y8WGyIXNhq6KVJPJkI63TshQRl+JzspMAG1
NTNn8ope9VIXhemeCaoexyJTQ5WO2Tj26bQ/CGNlxBQijbMd6g/lRPxZzva/
d3bBSkRntYnE0EKQvQ9pOuvXPs9/Oas1VHVbNwejxStTqdiXTyzedqsUv1PV
AgyTlb1w5QEvWJ2W7sjwy4tzFeIfRsXNonrRW8i7DzmjVXCh9xow2jMBfuPG
yibFvoMb8D/IH7Hlxv/bIL1yFPePsGF/5FIXEUYlwRvX9N6IpwmwDvvvm08D
f7Ejb0ZlWpCL/6rBsPU/5s9IuM53ZcyJsXX7nx0Dq6NjWWDC4q3NT/0yhkH8
UXIQb+FA3Cv8T34WLewhqETIM1yj1bj6J3oFbNF8ISZtvqh3mIvDEpNyRou2
FTsJRtMbRpT81ezzi06HFKWn2HoplT8en/O2mxfFO4d5dnEr7xtnH7MNyJZk
uAuoVuxs2DSU04BennuWBRjqcTRc7idtgR92aY5NJcvmohdhwaBvdtY9bDMa
G4MIDNAw6N/DpyzdyDMOY17Ymgd0eBx2RlZ47yvPb2Mg9pLLqLTpm8c580F7
eXDOooyMWdS0DAjrMN5QTbQ2hMAxk0DBL9K3NZK1Uei4yVrDNMUMH7pJIE4j
QvrCdFbSTzSK9Kp1CYAsPorbJAVsiyPiA7opAqAl/COX8fj8bsalIK85pFcW
3KGKocmb+A4wRGZM3EVxiGeyCLDMWkZpW7RtAp4ROfokb0sOEyPmBXGmwtfN
w/5M1HDxiWJ67ZybsFmEBgtIvG9oszqfeUv4Qh+PrBLyx73k0K8OYHXK7rzJ
WDxktB9cFxJjvyQhgh+kDR5KELPWEGPIi5tgnfDc4Hbpv38ZxFIpBNg6jARo
s9GBZFnxWC45+grRZLE30EzF3DM8SgE0P5PpHac6ZXyLejyGOiCLax0QXh/9
02zrcp4HOrHZlKuNq8ICWLDY1Pfn9IVLpZLCrQ1gup6GlVzmiKamofQ5SlA7
I/OMuYjPe+bD2SDjJn5wQarNuyDHVJ9CtWT4UH4QjmE2O0rWKP48Ubq7MWuR
IEtkuHC+J6So2QoEbtAAejgf57x56ZVX68I8Mvcch48sVs/VgOdkKXzkPOyS
k70BRqbDxmvxXnPluKgIEbII2NybciOB17AiYVxnDh4BVxH/bM1+6mzHSBuk
fppnGzp16Re9eaYjFC10lMrk4rryKpr38SXIOsZO7jdqKrRn68MYraUQh6/7
gSjc/tmy6Az81ITcJcNigR3wSmmVJcCbLnbI+iTDyKhSfX7hZkcfhhlIZrUX
2ijqUuW0pZLhd/y8rzN+Xcob1Ptt75kjY7nejklO0lvRfda61OggLTga8MBG
ePZHVGKvluurtPNRQ7tuz7ORj4PeHaeepJXIUPXRCnptjYiC9qQXHkovbyVY
7bl2kTGLoo5MD6dgF1Ng2BYqkUEKfiSIApZzeey/R5+5AjvFnrALYg/xHFxY
FFOJdc/9JTpKfPN6B5O5mgCKA9DdOGUlDtTnhZC1iYky60aK+ZvS3CMQQY4t
IVSNiT5RmWl4qLLuqpWqxvhZj5x5mQyC7/rDsNvZORQQTZ18yXdRmkTLcQ3Z
yv3vAoQCxvtSmaZ/htr4obxpZdOPOCYvp2B6Bhnyd24igJLL0RkiQcCGHdoJ
57tvrajv9kAR0I+wHc/7OIPDeH+pz3MVQMgrErtXuqCLFq+HWMbpcXZmgfFu
ft2LDAyxgNBFwzsurmOSKNbKVzYvzKob7ZaduzZo0/vPfkh19zJ3jZS/VQ1l
J4H4EeffoPjoS9WnRGkykwX8oducIg3vNzhlXeCfhKrchw3id/sqSxNnNLgX
OoI2J+38OW93tHPIRNQLil7DHtQsa1e0a67D7l4jNGociwTXN8X7aydYp9fb
K0wzGtLDYuBponG37CnGq62A4CUgLy5599R6oj+Ieai5ft+l+uKnifrHFPfs
NZ6mLrbNTaszHmgX1OU/Hx/zLbJ0CDvJZRoR9ppEFQSsqjR9yGx05aOJHYlz
ERD0qNWy4C+UJmIuUWrzAuekcafiNLR3AJkpT1+MnM1Gw5nRTwDwMmRcylh5
Oze7UU6LM40YYlttPIhj1NbCSGWOgtroz58mRV7QdmxJrF4ZPj7APkSPCM18
XXuZmk9mru2GF7x94b/kBpz/FeIPUbHk2bYE1Cj6l0dzvpyFL3n+2G7cj3fM
MskVbc/QV9aBvTesTiyZkaFKgAaXOLxETJBCb7fZg6lLMJMN0qphzraKgRSZ
4aBGtKlxfWy4xKer9rR39nq/0j8/0OV5spYITYDxfR2eg6/K6bL8FgEaCWzA
I3Ch1HDTp2ITeM8QUyt9tBWo9t2eiW71z3c7UE+qNN4+NV2J30fb6VeGNauP
c4HPHrP40HUQyS0axS1lBmbYPU9Zg/6rD+dwgVX+UfgfQFx5g3+bk2dOwGZh
CfeO5c5iYU/J46BqwJk7CZRXgm86TO3QI6ZcWJxNZMxdmj6lrFlN1yV0jlRS
PiA689BwaZcD/Ze4yC3YV02D1zCdQf/lp9/My42vOpfKmGDDpmH617duzz+0
bsJkErpqGzZ93fmzFzUyCnTXWTMmkywwtd4/lB9bYUwBjeV3JVLfvoOduBC+
5pnJj44zfI1wfPRUR1rrGE3fi7JLfow0r/JkeFOmiKUU/WCq5pAKUB+F0xrl
NHZX37tMYsYeGbnR93I43JLwUs/wdqSzMMQ1Y9kxvO04hyoNHADpL1LGlbVr
ibA7HxVqvJ3CbeD6gcPjjnr0UX1FCI0+HlJRHOv+BLmY0u1rt/64zeby9N5D
BL0D3GtBDzwHxS+fMGzBvXp3yj3LMJOFdrOdwv6Zfa6VHrO2RbVTKWdYBIFE
fMOaxgFdEiJVDYdgYfLYZVL8IActK/8Au/ma/19XlxI9SLnXNvdX4o9/70EE
7ZrLJQw26itwP8COavt+DXIbE+jFt+cZ/kXJRUmDVD629ZOQWh9OhA3NKJer
mZf8Yn7VWabpTdJG/a5rmAk3scgJsTN7iehJ0FzlgfE4nGDrTjMq8Kt4KiRk
PV7z7gBnMgFpkccOuQPy+FudUnRZ8XVgLlde2qst8f2DBi2IrljFie/SK737
AaLhxKdPaYhy/wazAcCjWXAhGkWQ6hSzGYsZ3uyFKASxCWwuWD2fZj1kDPYZ
pZ5M01KCWAmVxYBr8+s2MZ0t6Vw5DfZ6uSmtgwHNQAzADjivrvQPoyM3vTuT
eOd6oQXsS33eVONM/JwvRdSOEJb1+bNwc8YP7soEVldHbK9YAXejNBc+D1Nh
sSsB/X/7f7Sk25H5yNcUBaCFMgeApCRI+AVVzaN+2eSKLVlwPzV21Pj0QdSD
07oVWhKiB2TIcI4W1zIpCrR3m0ZVg5SYt7cqoiiBouDrBiFdPRJPjBH92CfC
jOn/DQVimPLhUmlKW/idTbrWCtG7AgO/W21ei7m2jx5inoI7bOXe4v8UKOHb
Vx6aAZ3VopWMvzegK5yyAxGiHA3gn9SN1FSWxAq2IJePZlq15B21+ldqNcwT
aTCVq15xpe/LyonSO3XQeokzhnBY2hrRnLqNpBO71zWK6Xo+3YdFynDY6wts
avNorwgWZavKU0xbBtX2ZYtSHuVsoNrd1TkKbBh9Roozs65MSkU60Wx1wWeS
310TqjD1VRcc9eupjSIzF0ndQdpX9cR2BiXTqRNvCVfEc8X3NMSOIHosniaw
b/g4iVNo+6QauaDa6EWdyWRhs1HZ7NeNx4cyT8zQ3zG4bAvFNuNtv11NSuOd
TZGRMtk6LhMepB/qgyW7XBoTRy+k4stjel8ZvmLZmNatNO89w8r9lQtF30FG
yWOwfT/TDUgEx/zBX6E/W2VV2PjOrDlQwbh7Kvyk5RiNg83160fYRUU5L4XG
KLBvdaRb4amjgsaZccNNcmOfFxLY1sbhPsidhE+ERj8aff3QdZk+i9+/azEP
W8ZFQhxlg5RS9hityiMPna+z0MptCgvsWg7AEQ35KnjcZcAopw/wamU51arO
hrzZBueHCyGeN9CdZlmAIi2AxOvRz5nItcc3DBuIawsLIp35MZtccZOQm5s/
eoAAFHb9coSwy0MVfOaTHyd+S0zFrMKYjzkLmCFxJBlyYqNvZWuyeo4bGjHa
Ue/rSRAy+BDE1g1aCcU7aZa5a3U68gtICHh9YqImCuG174Qi0JOR0rF1R2Lq
zuIjFCRbyYNXCnd4jajrNpEgD4sRbL3qensNSUiuSereGPMWG9eEQh1JReX2
8XH9L/yDCKhypU/KYrxh8vsacrN6gJUW3Tf332enH/skb3IFSQs3Kw5CDhOu
udrSLtA2sk/yeKs2nmtP+/YkLOSx0eNngrQTyTD+jZYHHNbgcuD+mEc5vJY8
EbFvHYpfLXEPphAeZLTrsFggIGJfKbkjT4HSTsB7fzLUkSh8o95OAme7Uz95
dKZ2tBNPC/f4UTEKmip3bEsfR2TBnqCbGxiTbLpqOsPM9zx3h9ta/lL5PCAj
Br+fzqwKBeelkxd6idOUKNscFmBSaCLwEbWqiLps2Bf+knyIooaTqW2CZbKg
+vBPnj++PkLqCo8FwrS1t68USChn/q0v8HxfU7mLTKH52gQd9iWIdqL7rgb4
LuvAbxFk8jMthor9RkUBm1GEs8yO3S0jvxhf8xXhOWivfcgxo7kTBFPHHE4J
W2iPKj8/NA8ItYCWKcFaNIcuDNAAboEODGWbbuLBd/venM6zW5L6Qhx7+KGP
PblEaujrlrfMSiZ27EkboRcu38Jw/MmzXesDfKaRtj7lXVqqrqZ7Zx4PuRvk
wYGhZUfyweBBRt0secHKz2kpGCWGqoL/p+s0h/IysLsEwrTZLJKHZILeb1Ig
iEmlXoSc+6FVJAE5CuSiD128pFjyhR5TbzAvLg28RePsP/yJs77Hkt/LTS34
J83nWBN4qVK4aiDNHzX8Y/n7EEWe0mMyM1tcDceSI0iacGEWIghS9PtdijLK
ZrBPRXj/ycxCCK25VyOeQSMANO+v+XPJlsYVrb/sjG09N/HxQw2cDREqkTwA
AscCLy3mc5kUdNoUDQcxRuZjMUAKXIPBjNTZzCNv6OiNI+k6UsrwIRMi4ZeB
TvdaveKBINIxImurVOO+4xw6BEgIV69rHsHiXt1nj62alQcvjjp8+KQwmC4i
0PehaRD3deoVBipe5m5IKMLoot1uYUAcNtqydMn6tyXd/1CT8234bt5/g5GQ
IkA4ZzHFIcsIbh9UG3pIB4HEaKLx0HrrEqS7D2/nxC0E6udcvOa4k5/DJMIG
5MGBnDQ9Mwwy+3s5EnUe6Cnz/Zv9odvZDRPDUSaNRwajL8NFlz302luw1Tfe
PoHR/xsReIGdeG5OwjooTDkcbHdWKfWKRP/PgcEAiyiX+sAmzAkvD9G4OJDr
x576U2O/THdoSRzvX3uqMBl59+8z9hgwDAb62Z9iBZzFxqJPBZd6HLjHz9+L
CN7LMsyzF3gn0H+3SQREIYRSLq2nqv7lio5YHCn+OUCOhebGkjjUa7U7ACva
/d9a/ftTsdgBZGIykjdxL6v9IoaLUC9CXj3wHMrr1VzogjlXxArhuqfKLD/m
kjOubq0JJf+xWkivNP/zrWIpin8hJHEUNBEl9Fb0Xoi/syCvzi7sLwcRfvD6
sCf4yIuppPHVgNj2lszElSGIudDh+IhD7pOW0G7B/RYPFhZujuvojo1pjp7V
/yworvgImJadU/B8ByVKHFsxXm8Pzyw3gG92zuvJnobYm5wjQ73Bxi7/QW5O
qpxCnR37jV9kh4Hfx3Q0TVQQoPf7w3ptQuXNbvg1nBZ2W1lqOmNrboCswNdI
H5S5V0fBrI4Q4cXWk2g/xo8bkepUm+SxaUjlROVEZIbdxUR2s+4SVBRh8nrf
emnC4n+LAc67HB6sxdcxQ1e5hWFeW5huBUXHDuyaVMxPsdkmGAqSQJcLrVbm
P0l3lZoGTQ5i2cujSt+HOD3KekbRBXJeu+zFU6eTO38JwZgRhlhRro0n9N7o
FpZkHagNg8VYs4Mcu6V6pFv+lRRrU6F87Uo9HafhFmGAFQRbgTld8RANUxT3
NxoUt5rA16ndnu+CjBmSEFQV5E2lkd+4hLJDe0W+Y6jSU8HhxPoGuCt77RkQ
6QytgFWk3tigRPpIyLq/LDbA9LIfL9c/99mLn1UMkMlaOkgX+xb35EOBzpz9
pLANEZ9HjhFrilEaicZ/pWEW6wu2gQw72cdbc3WrtBJbRx/EgKjgEUQh//RW
RyNmBeHLx/lg31hyKNURvcuWAmFcNiQOR6pdNg4UBkSaEEWV/KZlc3yHmg3J
UfFQiU6k7rEMhF8xdO3gsW7Gd7Y0+9BL0h0QEqfvPcz98Ohg9oGz7BcjVDbl
AZvUfgFAIf+lyxh1pRUOOKJNYPIOmK27pX1rXnWno0oR0ApFBJeu6ioQgYjj
mDGjKuHqlh0F0jTMPpKGNAcQfGbr993VCF0MNan34xsYFtYdd87X3qORdZsE
Q7gdWxhPcGZfSXlYI4fdin+8a4c1vGxg3Yy2wHSmR498zVSR6Z3isAE/Q4bI
Qh8a/xPTFyU2r2QdrZtBulSfCXtC7p3YRv5rFcIH2b6vfPo1DtgN4q55G7nc
kRSil9GBdbNoNaHyJ6kWHEARH8tIeJv0su0UanxDqD1GO/5kCjZCAgd9LhNM
2HGx5BEw5vwT5TOmhxnXg1+iSkIAIl27JMBr7HNt7M1JSRTE5IsSwyz6wgLp
oZhz4TK3MF8S5/UuVgLGCogXx5OAm7ujIGpbBO9nWQrzauqjKVJPri9kgTRT
SdJKjHfu8Vkx58wj3LRN4zWDvQDbS91ehPyPGT4btguIshcagfhOkhY8a4mN
sMDB8T///Zoy97zgYMlw0DWpEFZtEE79J4GtJx1GJZ43+BK5jr2lhLJC6Ulo
k8WD1KDgQP6/9eA6mx1Y9O4pKVM2ON93DsJSww3gWwg1mbJm18ij1xAyGaYw
SyJ2TJoxSTZTeqj9fWVYuGtMmfPMLM4xRsnIfmz5ptJinSsEfsaZ9q/d8tVq
GiTz5Lx+zVPEZq83xjAf/MMbmf4c79l9zOi8tmsldZbomD/JwswonXztrr8L
vJFuf3TbuFV5VBWhTLdxBpvFO2+ZeVY41XwfErYKCuFpgZbIhZukZm3UBu+j
BFcp8S1S5BuR636Ur9mbxphTJ6MhIhsaeb3FNd2P9LFHuWve4rzmt8yiBO1D
d6LXDEPkpB3fYG0xBqd/1OnfreJ+ahUVqXpe9voFanXxVTR/XHaPH5M1kZhM
r/EIAwubMw2SK3jvmMPZbCshejF0OHFuIZSF9g2XlWn6Pi/ObiTiMUnQLeQr
s4PSrWE125U5vaKRewLFrVa//UZIu76C7324mk0yEliWniY+4nWZ2Q2Q40E1
bMw8/fvNlQZqTWGuU8RnFmRbpGzbbDlIgPQTSXc0MkVSKiC7Zice1vmRRoxx
mSaf51nem3U4mnVXU1763jGFlts35JmMTQCLUJzYWqyNUf9vUvgLhPrGJnNy
y/A87PwePsQXOc0pvkECdUgXziEwODVd74WS6ejFVFUV+MWEgtCQRe2QZVYF
rM1Wznd4IphJQTFMULOfRlbZNCp75JvSFyE+5Fy/p7vkg1O0x1kzvmOjf8le
y5JzTC5eSUphBpH3hg9V6nxrDY39d6szdxqWy0yHPW6Io0Fbehxhz6OOohgM
eSIGrzY9V7qgOcSwJ7Pga5jH3uZPqm99RM4jfV+MvXqgKSy0l2qpiDtOp9+e
xy1UOji+4ueRtRZ96DjjFoMKURSRkMu/M4vyIuycQBPJ9KKIVqQgNCneNyd/
BiFiDpxeeEjQvTwgJBTmS/BVPxW5UGKlw7r7QSubQg8Re+r28WT552z6GXk9
x9QreDid3PZzFnC2pvpqcDQtYD8n+keAJI8Qxl662jXeJHw7Uq1ZSk8+GdKy
A7s8OgrYsPjRkpyH4Gfeg0ZWdJfC+/KUhCLufTqis+4sP2WLFZc2R9wV6cy5
YYcNsn+6pfn/r5nFWSFRmLPb6/CG/Q1mdJHIe+iECndS85XorQAki704WbuS
tvKbNOPugorMARk3yetBem8KjNQ6ccTIdzk5KD+BgE3Oc3ytbjlnBkxqEyiK
cZfgkCCVY/5hrji3Mj6UeLFZQKuvwQQAqoCiz/+lVcWV2l+H8/7oaCRua3Ps
9Cg+vTHXi+5rzYR/PiyZ28b4kxcCFt3G+xrKDENU/lIlE/U0DAlITAzVymUK
fNMuVUQ/zBQCT9X6zVyoDX2iWUCt/YJsfZHsCVIhuAOLSqy54UgfKSkoJLv5
qgkNAYD9l/UJiODfppObK8fPD1T2DmE5lS5Id0HdXsD+3g8uCgshiZsvSKTP
+uzbcjg57OpPxc76qqP7/QQS1wCOlGo2GS87YGn+i31s0y4jkeOrSHri+5V/
LJeVXf9xFzOIAgQaxNHOFtqZeexywM4o8hEf82ISOPclLUdea9Deh7eaWhKO
JZhxhkGb6JHwMheKrDywflTHw8rIFIipmQkmouu7fTloHBjkzhFaD0h/tg/M
TEVpTPADXFM/8ZxOfIJI3gfL/SKBYTY1Z5aWSUAbHrsCypYAzHzjAM71zTxI
PYAcpd9wXkmcP3dByVX0L6PYkIPci69RAP5DXeoHySHrxfF07kJmOrBAMyg3
3e2Dvk1QwYhiwyrYKu7Q7GE809yaikui/blYPNPZ+iX1Ul01CGoCRxFfz+dt
dEhYR0ySs/zTDQ3Sspf4Qyqio7L4+YzKA5yONUqKl5QcCbPRtwjGLaWc49SB
V46iwsBIyrdyj2qXSuTNpsZwYzvi7JD24gfYzxyL00I6ih8DnYhePByIHYtj
cElCCILzSz9kyuKtl1evChBpJh0B4IXJsrIHiXBzLotGJ/w+kzi8TxsUczKQ
YV7NAOrH9s8u7YINz6QHb2ZqwvcW58KxjvY5qDFFBu7H/O5XiQad0PGvwjU0
SXCOK17SER02M7TQxlWUW6KYNqkFzgdGeHeJAax/3a2qOHmqkPyWI0w4H1Dw
GKZ6oA1bh0YFwiwAYPt9CTgL1xnYcjuXpLeNuA5dJ9KhD99bdoC6UWL0V7T6
hmF1XASDbhA5qc1LMC5zYy1jNJBZ5lMguls2csSBbMYTzop7BoaI+c8FtJpV
9kA0Msxib8aju9lBaQDdnoTBBthJT65csnNePmRFk0FS0eaqv6mr77DnmPZT
znN5NUMeqtD6P7KQRVx6gUwSCcLcy3owhNlz7WiK7lYnFup80lu36tysMiIH
ReDGxKP5sNGFlgJtTJvnltGAaMKVqkcnz0BcpwifbnwVIrDSDHxoiMV/IXlS
B/dCPoE5DkIjjwjHp+nKK7VJpueOjMWaIWhqJ4Z8ugl25XvQZnEYCXWXc1dL
ag93bTscVKY0drMYaPkKTgXtNeQvMLcWe7T74Bbq57+JXrZvQTJMx7ZexrWh
zNHPtzfr1X7FoLZXva1Qj/rRU6fy2yVBxPQeJG/2l//KystQ2xLK25p9DlCQ
Fzacp4jZQt1HqlTEzn3Im8C+rhCfVmFEF415gU3bwvWb1g4O9498itRUfsAv
E0i7tnd7MkZjCi4XLCafyVlqwnWIQRMArWBBkMHjzWqtEGwkD7bRtQKuIZXg
jI0+d5JM4vwnQ+oZS4k7rJWMPHdC5q0jeIkAvxifp/uBnQwisYgrewpFsIJ4
OxXIT9pjtXWVP1fCKgH6CmkP4wv4Oztg/hY2RWOp0XohL7vVwXS2q1m6SBoO
rNMxVPqEPk2PSa34okvzm2aeDHg/Dr/ILtv2lKuNR2zssfDpIIFWRoPQXkAe
NBftKqInkpr+pkQzhdsd+P9YN0S78ezt8bmR9vqOaxkR6/Nqqvj2nU4bitF0
GV2M0YB4L8CvnWt4skyGnQYs/Kmf0hjaCkDjyBN1MFfJybRIllRwyeZeomPl
s00Li+lRzfk6D7ccsVD/dAazIYalWY0WpnA64ZiUtlF9UZv+wiZVhMtlArlU
upCNjLyihP4cLCXh0DfS+lPUp9+FE0koH14wqFNn+pXvNwHeXS+kbd1JKeP+
4MJMx25+5TJc9jskQ/uSezC+WCo+F6C2fT9mZA7b+Epxc0H6tUPx7rASeQR6
lxvfwP49ZiScXQbhGXUfgPt0Qhc5SQN2ouG1GnPZCUXvTxQ5FB3LFr7wW+7E
Uqv8VdYBYYtKnUuPPBlpwiXiSPBYiQt/2oqXJp+23JkP/Xlxh5f1xBx1hAUW
M4BXqOzM2yGhbK3k3BfMmjv5Nzz5wFqjZgIiJ1S/tE4moTr2M6rT/wd9HnPy
/XVTn+Nrw4crywoZRHy2+cUzXPfscvolJEP87NsyflKhkLH/cB0IfvQvONZ/
HEQtmiMyU+jfO7OyeFChVIm6QGH8esFMnhNtPq46t6tq5JyqT7BPLqtI54H1
403ddC4IJjBH3Vr7JF/LUe1hN1fk5ahGZpH0rDQfmO6qAWdCaL4W3Fdr8kq/
hxw4mKuvl2Pc5BrNFwLOVAA91GY4GFwhT+5W5rcAWjIN1hqQpT3d6dNPKUtN
vP6XymK7pMx7PMVCJw2dPN10rwY7UXr4KpPUhRp+fJds9dLiS6jwN0AJEVbk
t2MjEDCiW4rEXy138OHhkllwapByMcEPmYZWv1aHGpk113QtsFFwn6jQVpIh
qwp3zX13rdyE5cfKE+FWFC49Yub4P5JnmCiReZHNn0nVSfBg/i8iPKD9RoAE
Bh/JRPbhRlDqae9SHHT0nj+lkQVkYPL0vxIY4colnBIWMBQlWx2Wa+0aWfCy
Fnl3fE6GDJAY8W/8HMTyrcTRQGlUZigQ4fmD0FRv5Fv4aUehgpFsHPoQKvZj
NImrEd9TMtJhYjd3nZ9Ax3B4p1GE7WN5FGVLZtRsStXlX1KlggYqydvCko2p
G+kXMLD0TAyk+qfThRTgfZe6Ueqe4X16aKcko2vZawCa88J/ZvE512TQ21eJ
xV4DA+rx/OEOEt0pBpLih9tvaHOrUH//8y0dIsZRmW0PHtTdXhcaS/hcFYmb
/ySCfQtxZe/s3Oul+W4u1j1wmnZEn571EwNs6nTLI1oGDCEp7/bdfKc9vUtH
UsgHey+M55LChITZ74rrAfLf8OzrvT5YMIqB1baSQ+77vdAz+zZ8/wKS6tIt
27zE/9HwjrG9p5OJ0lYU0/+wgDIGBNEM+CjlZW+kLrD1n+RELoWIiXWLjX2Q
XgMXDQ8wOJHInyyzOwsY9PxekgwM9TKehujOKB/B+oM5yBht/jqxSCL/dFk2
5XSPxz359hkR1l4ynnsc9/ePBjd6gLkomU8VVhtW+B0zu5BjGuF6KK1EvxgZ
+N1vSffh4rqO4gILdGDqCQY46n6M2OxD+MlP019n1AUWb0qskKdkjIcV0o0a
pJH9uYZuXvJDID9JBBh0rf3ubk5KeVWVpUNsrGB6Kw7meYKspMSOHv1ZAad9
AdDcHaudwcihPxz3m6aldj3aA4AeeYJLMl6LIKsw6VqdB5qNAJvyrVKTlIbG
cjXdeMfWBNlXGLP5vKHINV6br+zi4uLnMh09e8LqRnjHfjyH9WF7C2nfTKNW
12tJB6igigBHS4qdmX8854+c5cIDQ2ovPq1YWowdObIXLlFYkraMDqGvVnK4
U2OgUTl+jQzQh+3BxsH7Mrld6lT40bG3IEbzvm3KBDb16siuiqEc2jhxNPZ7
d1fbwsGWqeA+/pPyiRWbROfgG25+kpZDJXvZ3Y5imfKNgHpo9V9BwWHdyGFt
WFGocRoPpqP/g89IKmF7ZhbNG19odZrWaFctAFhmGDv/8nU5uY/HPP6RZABX
Nfdpi2soW23nvfgMrosC7EbJMNNBtXI4s5sG+bqwhvztbS48ip26F/dj+W6I
SS/S0vlINeOM04e/G1PgxqyYZM5V78K3nqmgzz62jaOa9xYTUqTridWNFX4w
onsm3aIVQa2tvTiK+RCwdahhZ7BzIp6p261shiZDy/YfH9My1fISsP+T44ov
2n4iuFVA2g+GsXrH1ODFvMhkWu6HeZ0EHP4oEjwjeU0GCVyKsJXBNNgqAHg4
avtVzBJSkmHbnuxUXg5g9XPz6Bb76qDi74Iiq5B9k1bSCtnU2NFabrTPGMMz
wFmz7Nz2nwXFmy0p51ZHbiFAvRiy4Bn9IIHDs1pmCe1gB2SGhlGDOZNZvd4y
onaaaNtwx7gsLVcxDw/302Ftd4APeUQ9TI75irlA/qTxhB+TtnbJ9cCNPdqn
xmINCvWe20h/0wgX7PxVpa+t0Y307NqxQjseOM/GB3Ncmx/+R0RZ4qA065oF
RQjVaN/l8MNTw2ooT+ytNm/Kggd2fEZJ/tyq9y9sXOOpsNDcQBaKXEAOYw0x
2S82dxRP+XXQF4Ta3DZFjHKSBDi3GXlJr4rZKJnhlVAUBza4d9hTwuY5p5vM
Ufuk7mYTLryMQvzrFXdxJ7HOmWsz6Y79i2PgUZiiMYIgudcLNg5+/89iFINL
wa/aKH9CkxbCg+IGQAOFly8HUzRds2HGD4q5clx2gYiqCs54wh+VK2uylEe8
0Kl6hIAhY501qLP+i3vXt0qNkNAW5KNuqiZzW6hoo9f2P5HonphoX3ESLzMM
i6FWJsZww0iRS8b6POpu+N+fricdWSTbWbFDrUeUP/xUDy45blFd0/2JsD8n
9TDzDCiHyGjmIfqmKd4cvrZWKUmfMV4ZhCayzhatAbahNk+2AelanTCEylup
ZlghriZD2q2e1jrAkMlJZ2krLqzxORH1Uwag37HRNj2JmApta9NHBmpeSmYI
N4QLBV/uuu8Z/SVxW+CW+gRam6hGZDQWgAifRg/nYnOmzlumf+PGnxNiNhkc
xUeUm87OtTMwZD56ItJCye8P9jqu0XocRDGYNB4tIIX/FgZ0Vz1+i2NOzKV7
S2CftqM35z31seJYoMhUlRwP52rlcopFYV4B7m3NtM0G835rQ9UZHsQWwzss
HjHV9wsysmGLdvSIJw0I8YRc/DO8UMLZEmVdIkgy/RVWRlXJjK55TZUb6LPR
1YlYbfVIsdTmz89vCR3Fb0YhVeSkSwKm1bEwAC7Vx+i1tMvhQgqUMgWAD+4b
8D/fOXyXrKcb7R8ks1o0c9MErxfSs1Du3AuaBJokOMB5Sw6/dc6y5BxneCHn
jl3JvnG3xzpgV+hLClqJfnVknL66bKCPKeWFIMxQ1551GElYKhbYvvwwqNBG
iv7E8qaauzROjBB31TigIi2L4jKWR21qZL+RE5ssSnC7yl4Rbe6zZ53zXLLH
c5I5hovbNSqmalsBdBLoc2EkdR+1cqGqCJTwG+YPltR/QxFZjEucSYOMwsSK
TpNgb/D1nfcpY52ZJLV3lw9bBHUpoRRf+wRoYYIIj4QhI49b1WQaHXY2oaYo
0brdteXHYuCcC86QE0rvKUTiHSKviJO860JqacMZ6uGaY5gWCsiwEZTcQE4n
TCmeaO38nEqrIekDOuxfMWHK/5rwH3gu8YYpyje3hy6YSxq9t/E+oHw4DfbL
mEQFBthHNO28P/ZVzqhlWCoFDt/8xq4VVXs5FNjYaVRUj/qjBmXSaUlbw69I
kpBRrE6zOjdIRmMnW2FPsViY/P8uuf7OG1Rmd4mrkKa0GayEmLC7V1Sv53CV
VNOJUUOWkRKfuJeU27EYvqWmWv702FWM/C3zI5u5YSye/aKn8JoNUdHJOrRG
KFFxBwYabM91D0lMEA1NqXcG0GxyoRfmoc4/a9HkjTpyyC4Yf2g8KOKH0EbN
x0VpULXs1xwABhgEra00GfYhRl0lVs/5b/Nw5jjQEvpV+lSj0UqyejkAYFYz
c6rAnDPgHnyK5fRXfbhlEmbDKI43fd4H7b6ezHXVKQFriEsyf68pP0bIzJ8M
ctq2U+f0a1s19plcxgv8TyD8rTRsdJ9ROQdpHcV+35USv42hSmm4jTTCN/ad
fKgNtrxEJWGqo/P3b2CkF0klb1zuWgwtByuBl1e59+N8rc+AUyGuGZy+1gI6
GWgAyr5PUt3w+aOkj6QuD8kJl6e7Q7jXvQStg3dnV2e2V1abG6Bkfx2dta3G
oWgZJGxCcWO2S3e3NzkjZ90gXsu1cydRlm7Tmlq5b5KGS8mdcxPOeeHdCc6T
5aNVXW/j7WcWJGmBPmcWtJnaDlR043dLcLz2wAn5SNrm1xUuAuCHRq/EaLIs
saaaR8/RqtwPYFYw2QDMltPiqwaseWIiTabhWxturIiWN4fcbsXs2dSzjtrU
tQY8AJp/y/92B8WefFT+PjF612LOSx3zAqtdTwi+f7lG6hEZ/bp/aSxLQdT5
rLfUx6EjEACYwb02054ChPCCoNDYuUOWuI1ujIoKh1MkhlTha24Ald3MQEt8
sCjO97NzofUYKRO7oAhpz4I0j1ntfnMQ1LSfLNh0WxG3Ham67cNBRzpy4yBJ
4kJkpfYHLO+3z422BNiI9tQ3uLAisAZcdmNcyZPMDmy3z3h/GhFodWZQaMNJ
VyVTEE8igh0ZJkJqhYlufytiO7HZLjtzZQQ1HM7bwycXrMEhE20V+D+WJ2W/
p8o6hDwnvoLIJ3Y+h4m13ju1wkRWKQOiOP8uh1QLfelGoFm6BKUDTanxhxS6
LmnLnaXQMVEvpys9FpDnyvEiqOjXfbBTsc/NR0GSF4gaJhktYCQhetZua54E
EEtVmPzmq+6IRB308fifcfZqzxGLPRcpvH6ewOu9MiIL4SdIef65jM228E2z
r0hjqPKfDpiPo/5mh5vKXasmrrauonxZkTGQDaSCy9+6cXcK1HsRZ4hafz9z
+y7r4+yeZWhEhljfw09tsY0kH/OpS48Dh2buUNu7JFoZtaF404tFMwBpFHB3
g8J0fYaz8SfBmiFdPlUo9gJyKV21e24sPrD7i11G1VEk6Jr5ZKntug2TysCF
bHafx/61e+bYM5b/84q9g31HcljgEnig/AP4PtoIo4qZzuDhBS9pqa9oOIoD
eow4r5AcEiDiLDdg3Sr/R4G/X1FGRgpomTfMq2nK7iFuDbId0KhCcDD20au+
ZgzDvsMTO+6D2sDO9Mm9RCd6LgAc1+GfCTuuMR6p+yIFCt1vjB7I05n00kUy
P9+eVostliLp6r6AFSaFAT233xV0Fprv6+S9hdfP0Xyhqrc4Lh0tuRXS7SYn
/PbgCJcvFVWF5I8nl+3fgf5DAiLUXoQ446QCFfV912/OswrgCMyKh+j9MCQH
7uQBWoFxb5ji5zOwPe5CPMhdCGJhQFoV+gO8mUnDKQwhfBET4eUcU7gLvwhT
NAc4b9iyQGvo8sXT+EBG4e6h7f/Qz/2++erTK/BZykEV4YcWOhp5yXYvqdSR
2r39wihfgNFR66UUXffptoTO+lVqIxUifDtq8vy19DpG7OBDxWkF9ptRJKyN
JLwSQAbFfOeuw22nZg+IYrjFqZypflYCsD0fQlAbyACTXcyRstci5f/Sonum
BYl9fW1Vt9vNARLz3fhNV9E44JWHZvmTKlk5J6CYmRH2kBfLMmEbanSmbEWO
3vu40MFWUP+Z2oD3ngQuF/aQc87JZq6ZbIrKGlCaqxRYTLHQMghnd8ySd0Na
sM6uOzEZb/Mc1f/VpjbB14QZVBOtA7LEmb81/x//qCbFR5YbyAUifLHaPyMq
AByJarCuSRzF5GNlk+cQvx8ZCLdI6yz94Ew0p46FnGHPSYnB1L7hqtHCP3L5
IMYx//n+55RatC23HMSb6pNVAEqommVqOIO4K3mcHZAbdOO67QZ8SjT7cYGO
AIPnmwRRYG85g1o6A2+a2mVYFsw8Kw+g1Mxy0GHfpzLyAPVRzCU6T8jgVOhX
Vr2rCtadfRD4NOLrNcykK4FtykSL10PQzSUqG+EwC1MbMmcBwJzWlXJvGCO5
if442UQVaZ5w5uVxvW3f7m7RqhG4L+LLi2hXplWP6pHfZDcQ7murMCmBB/8R
y4kke+MdXGzXag7aHwb8+nO735W/WWISOP9MkUOrrmbIwtHwwrwhSRzFdegy
MLjKTyk/KhK0LeH9e842OKF0p3iNidyAbctkFHv1VG5G9SP1fjBKZc/ZZTqY
kBHO8LEKTgH5xvl/TfoHrAVeIMuPCarvlnzT9pF5Px56Bj64gL/ByDK+wWOk
JgVJK/bI5HDPfDzUpI7hd31GdDlFmerhEujnvSNt9ci/2nUYyDWhQYb6afsU
J95RweEw//Flt6z5x3a5/F6O2Cj4iXZv3fmdTVbt+eu9Hq7LPCPEOlXfScBY
9k20B9oyAA5uK5sRvA2chySe/WpD2GyQ096tLLxKNMt65GryU490o+5kOVjx
3RnWkks3JjSGD0eC6x8HoHki8DamaaKVUIEIYlMuAden5I6E2xPIymiIPjb1
NfD+9R/oThF1X/XI4Io0ZeXMPs0GINaJzl2Nus1Kj0y1TlIZiWBUKdbZ+0SB
vsfFFNXmJNXp7k/zra7sBnHh9I/Mc2of4t2R35vjDD+FJirH1EeRonH1xSgo
PIknZcYIJyNonmTsymfzdljwj4i+EX5EerYi0diGw1GwLA0P1wkh27k1Mqxo
pKojLBuffX/e5dSaw3FgizZJwC1DQvecfEVGFCHvRDseCnAo2EvSZyj7/owG
0R7L0UtT6sFXJa/6iy6/Ml6gvKgLYte5ROUKAkmpeRJbB29FfmgaXTb13AfB
majaYnKGKbVcv8WYEAD2qpgqzOZloWhJkqjqWfgr9r6WpjJxHuQJsNJ7ACgF
Gq+OrYx/N35NL+GESM2kBCk3S5gOymhbyhubN6Y2NhQ3EFl83FnVcY/nqGN3
2QmRfQqyUXoztgkLTF1YrwQtOz1Uu0Q71l7cXAmXGy2BWuOyD5cxumuOrwQ1
tFvAn1d3ZMIfTPGKGMv26S6UpQc1fk+0l+6z8Y2zpxc3CRPJB746ziBIACWr
AK60V9myw1NcBjYCwfq7nZqOJefL0KhX4WvBG8yhN8gBBzLZfsxD0tWSd9/R
Qnw38qDaziHc4TlJo0ccdGVKibI16Fq+TjEv0lOn/UIGZIDM/zmG7pDt9aqw
bjGp8xz6J+8j/L21egFzK1+9bRbeBmntzPS5A2drp9KUfbzUZFi58ESNk2BR
Casjx4sXJxaa7CKKLvbjhjY+VMrYojX1g9Jf/wUdhcwlcvqI5cK/E28lWscx
RysRBHAU0IdpNQvZVR+AjkGAmhzun4137KG0NiSySNBfrk9aalT/J8kHOfHA
o1XI2UyOuD9vU2txeTF9pAh2To6mR1gZxrRAtrZ5oOpk3S5i87mvcByoR+gD
VLksTUAS8tEEfaE19RdG849t+UBEAT+7fcqZu1qnWYT70zVlL1HQ0wk/wrIK
ljSxKL+jAvG8RP/bvK9A86R0dgQ/KjHbtZBe4J9+waIYKr+JchrR0w3dPFlJ
kofeGDLvfQXhAmYUj8sdr6FMOnlqeaFb/vx93ytjPu7hI8Ngeh9jdLt1Xkcs
bHclqyqQZnwWlKQyA5aX0NO/DhcZA4O9ZAsaJkb4ZOLv12XiyyscgU8ZRVmv
ofpm45xMILdF2skP1q0NnRMob7KILM5pYu0quRpp78xLtu1+bA+TaQzLzePL
xBbWWwgavWUeEarv2ZjvZ9/yNW/Kfnngtivj3L26ZAbQ38F55K7kXpYOZPLG
MmRmedKQHHbMLJ2JYZcTXWfGnSAgEmq6aRKgC6YMcJVmOPoZebIvsHA/Op7R
HVlo7ei43eFbh3m2A4a08UdLQCJK6fVYt03jTpgwpeJIn2r0cVkRn6LCI/vO
PXq9QRQ7XI2IBQCBufOD6eydy/hxaGJeVgWPnO7gvrJaf3bo768yASErAL9d
Mi9cuOE2hoPPt2adJP8+5q+e6nGWdDJ2QwukBX8ZJHKZD05dNZOsYnFIA21Q
kx4U3x99/qMrOhukNVMvRQF4pYN6cDqJ6EJdnO5bk1JDn664a8aka3cYuPCP
04hcm67AaVMr/GKTaKxpVjqKUegP2CmoWKKbB92fdh6JpQTcywUm6bcQqXZA
PjMeiUnUbw0bZAVJE8OnNFie89XACrJa15kTpfG4rVmQu6yE8umPwxYqXFoo
2JLZj9ZYyaHSn9B6819h/c9dms2oc3o97LQu/NDbAGEJlLsBlYU0Ey8bNdBd
Z0kkBRcShDmDcE3D5abv1zfPZv5MO2t+erxF9gWLhx4JfrEjZiCGhK5/NL5e
MvGQFpBCVVNnlaNiN81081NKVERKUDs1SbYsOepdv/2tzT03LBavmZvBs/aM
KkvAXB0UBUe6dklumhYgIuz2+lkjB1aYDEfLbGTcQDn13thOoEBURzhP8Be4
Wl4tQ2zU40UcWotaaE6/v1GQH1lErzCYaZ5iL5KZotpOnLK5yzsWtFpFU11O
mE+dFJMoojBXwPVZXSvvTHdJW447uTawAAFewm1Z+fSysr9RVINtFgGy1Os0
XUyY0aQ+R/x7rALCij8Pel699q4y48Sbk8Y0VW9Z9LLTjEY+HRBy4xZhgQdO
V2q2mCouXoTFz0kUFuKEbbMBEJf8hYur8B930OYJ7TZEreyYiuSx8k2LXDT3
EDI80vHUz6qJvQ5OUrpDAykvR5Fr7u14IX0ur/9WvU6OY+DMYh8XPnPyo+/k
w16mx4El7BX62PJpJfpAA62E8gz1DOq6QKDV4rruZda8CYPOP9HTRTxP94Yf
M8iSokSz3QFonXDF7HNxtOt8uQ4B1o21HqJgDeM/HYKRa4kAahErok6iQAY1
kCbgO/Wp9ylCf2G4240gMJt6/QqmZqTFK1r81qD1/0V/PWUic9W7qLie3za/
vabm2NU/Nb/XxzObijYTWPLqmiyHhssHwip0+lvhC8c4PKUC2zzRf9CA0ozH
kzV3O8ca54QmXYNNnNeH82i4XzS5RV57QErG4Lj7PduFrUBcsuJfPwLuNwMj
S//YxygoxrrAY5hAMBOEGbHV7+cGQ9PpQv7NubAXALRg+/yffwDFPr1dY4IK
JGhYFyiBZwLAoZ0cX3Aq/gywNx2P8C6O+LFXHG9jwU3XT9VVMXsZuz+QCVdu
9U9qC8GP1ixbbggkqdmbePtBYeC93K9Hv0Q7bc2sUvBVZ1hh8l9Yk6oI13Pa
CiLFFCgZN4ZyyJvzTTjZUG07DQuoD9C9xjmVqdoClABGCw1ykDIXJCyyZ0fi
zt5kPpvIR2HbUmxNgYZ9lv69pSxug53q4+eE18cGyk9ejdvoESxoNkhtCLz5
N3pq7exK1auW5BP/YUuMxPU3qvJufZVQW+YQEd0qwkAuEogEYLjt5Zq2Lh87
xF5itHj7rQseYyoSam8YdOy24sYUy23XCEs8KE+3cGuKjSbI6JrQKqF1sETX
VYfZKd/MOKRsqOUutttQATkMQA2wpySMYLuG8kwfzFo98rCZgiUf0XwACXcm
gPBCStgE2FcaVBBFeIJ4JSVqeOiI87Ht1oDZeYuSEqYUB6B1cLPY7QrF8wEb
R0DyCiCtWQTn2/fV44F6vJxK0yMXAAEgpOISXRleqmjxq0w9s0gmN/fjb7jz
dhnuywWBQ4ih3+2IGea9MKIFQ8019th656tNz/JuN9p2HoV/Wh8LNEYTU7fB
2I/Ag2lFd4fWvdfUBMlYjlS2sS7UFJspW3tpi0qr6lvKrrjwEnF1I++8lZ+F
b83Re2Bhodbq2oa3/OcFXzJ9A7uTBGAFc8LAORn+Fm9ktvZqeREJylUzpoUx
RIIfmULSqVHAhPSONbuj0INp548KfrPcSbEM0iJ6lS1osVm3pwjRLKAR3Auw
qv1XOgkTrKahTIiELOBSi1SaiTW8b5AROW4CbjUP/Cn9iCBeuztxN1C9xbs1
LgUDgpDD1LqRYFK/FF+JJPYJlpR0f8FtLhTNpi+FM0yWBWv2pQqfd5cr3S7t
P9HZjDP0d4kaScaqQxjtykz64ovzo5VshpK13HCggu0FXYtmaA8iEe2svR1w
KEPi5L+zoOhxeNiZjGR+WHb5aHtaLYHK23NCE0juBio4m5A7DUYEhx9I/tNu
4A7Ia9Pz7sON7DPrrn+rv/lrdrukJ1636pqUtk5uyXjQni8+nW1Xxy909clJ
8WKMKZ/P5bzOSen01PadhMfdGgSK1GWaUVjPKuA8WfjQ0bbg6xJvjOqfoR4D
s/LakyysXB/onrKFwNldv842GdbE4KM4bhhJ1PjpVkOnpcHix9QqSPZuNe1N
DvZ/M1pAXHmzF/YU0oDnl+ZnEgbMIFUXyhz9GxM+lzUnhcwVhVByH06BdrFE
xtZ7WbiQP5iGCSo8BnNDnjvE/Pn4Fi3+fzk+MAD2oK6QR+ZkODK9Lf6eJiaw
8LIb1wtYpGCIWRyvAIooXBRNV2/Cs+MAH20ZWH86hhNK/R8kpsgzQjE4z9d5
XgWtRZOBfRA1GfXfOr5rY2+GwGHjdiscSx6dnXTHBp9Oz74YGvi0IxpD7jfJ
+gWYoFMX8CTWBbqUyA83W1NOgFnr1omQlb/exnkG7zrYz3kr4vnKcuIV2Xzs
f+MaUsMqVNn9LNsYsK1xU61mnJEBzlAdtgC1MV6T7XbeUhFjV499fAacKiqi
lgLl9rT0k4LwqFsdEAiAR7DpbwovhscCZ7LQ+RqHP7J+HmQu7gTV2pEIEnw0
RYei0Qw8K/vO9O1anu29HOVt28bW/NBYBJCwrJI3Pn38P8+YfZrEIUEnoCnq
sJnS8wwHQ9MtWFWvjeQca4W0Isz17Q8AfEVlLipLu0jBaG4IlE4DvuxlUmZD
lr4Fe2NQWDkKpoJ6ANRmE0yT56r4aQ1jo1Okv7R6t8Vv7DYlMA11wVpr8OKP
9OL54k8Q20n5s9oHuNg0XTn0/+EX8Hrho1g7O3CvrkPHDdk6++tEzabhiGe9
79j5duxLQZmpTUABlVn651R+k2qcNDCa7OVY+AXOqTHNf3kS6gPt3bzLCSOz
3KYKkZGMCrNk0x8nV72rXA3TR8evi+S7KeRZR8H+240INCnL5157mWhvMgkR
4EUO5j12n3a5TE1W5BL5C+wq/j1fYK3OGmZY1Uz+xS9tWEWjSGSzQs3nsp+5
u2ioXR/3nQ0mKA1ZfjaNsNCGk1xm+wqGPIQZYwHhzTir9tnEUpaOEhCl+2uy
d97JH0iuD15kl0/t63v5zhG9BhcCWHEAFQRgEu++oT8cT8Ba2HgBXocQzFnR
dcHGz/nTGzs0yKnZzdndOVMVw8rA8YO6xae+18Xn0xkGWATfYVLXFPxXHuEa
hFD5yVioGt146QVEtM64R7/AQN0BdZ62jhYhf8WH2WKj4dHdpYNNDCIrlTgi
HhqXeXznDlEsCA8VQ8+GLbT1wGJascVkfg1c8Pd51oOl6QqgFXVTqsRfTAz5
yeFDDIi+jaza1P6SI7XE3o8EdCpHlNRG3OZ9EC0qhUm1LTB9xlKlwXC84NNF
GWiL01KQZkjC6fQ/acsgkCxZrsUuiwseghDubnh3fCH5A7/xF0f/6VYNEmpa
o22k/z45xPSEzSXgW4n4lVggze1d4bYuiJMFHWAGYeiXXlxw3adwAPsxtSBP
0GUMEh9eormlivMC44L2oD6GRJa0ju2440WoEUU/PHjLxMjjopA9cnQEgaV6
N9H7xaJ70va9KzEX5GksoXnVFIVLUwbulObV6cuJMyIBVJjtboT/OwNkzSf7
oX6XD7ujHyK4og7OA1dsTiypZqBnFPv3QD78E7rJxMkvbqk2To7CdlpY77XN
juCGTV85lk7mNqURkVIsGBDba/N3CT4JJ6KM4znZCy0Yd7gIkeJLpT5GUfmU
dmQstFYDpgX/kMvzhxsx+TqBl2Kd9ELH8vyYCFxtZaPUKULwkgcIfs2HtLCV
O6WkC+kUFODcNcPtw7FC1TjhtIFcQ/gx3YqJM7WbeREfvx0sK6Mur7ZUR9d1
qu3Z1KNWhVgp1fXkaNjemifcZb7bAH4oMLqo6wNMP7ue41CJViVbyb+D/ZLc
VlHgxKWNHybbUG4jFhKGWr1p1Tvxznw3jDF/mQRzRhxBRyhS3NJ2zyqGZpkf
4Ixv31MPPl4y6FR7jJZeNyCFmYXbHZeTV7N0HloJ8vrwC76yn9O52wd3Ja/D
5JL1aztzOhJg5ywCdhl23xBv0q3qya79pQuYw/hDGMhoSSlzIddBvlAHIBB0
+yLA61MXTuwYe6IeETXHkjRBq53PPf/Kkcn560l98kghZouxidR0Wt+bCOVy
NK+RPUYbr9XljlH1TXTXIjguJvrep32F8omYPdVDSkQA9WeZhHNCIIZkfAJp
q2+ChkkKlbnm1ejiEgL0Y4RCgB9PH6EUu5/pVCrMq5Vf1KIEF7KuOKbnq1Wr
1mDi6jFRwK0Owzo81dWYUM250K0G3gfdL/wiEeI5hh8o2+kZjhEjEHwkT6DN
y+j2PtcYIiOVJ7W3Qae8hwOi8AgWl/T2uRAigyi1HR2XjAaapPi/wjkFpnBF
1nAStduA9aHbjT1xyNp6WLZgC33k1ZqrSNu3Td0Ti9q90qVMj5hA/uPQkKsi
Uvhd56okMSIQxU2Xfv8nQOhXhMXk8WrSBRLBt074fbcAyKxSOYo0bdNWWvCP
Aev28+ri4MDqMHgOcYnZAaEZ4w4tiFrxkfmGhb8aKu4N2ZEfxVlh9C5a38KN
d/YMuzM7j17ganMChravXTApLt7K/WLpfdeFTuR0x4y/wtl/qv3XnYxAJDlb
JHjEZ0pdpzt2ilUU806yTvnCTkbczXuZHhBsv6sc6ND5E8grm84JVYe+Oi1K
2Tjz34elfIebsiKapRFiR3nC09trgcfGhiyHhc1QHyee3xkIorlQbcn3KylL
vnSoZWOJcmv3SGpxoBkptbh5qtAIAl36jzSOd0OljSpsy0nnzwmzdlXI3cnd
CZVc4HD57YlanFz1Aa+IrwCl4Fqoyx1vtWmhD00csNmc8/lkRkS4YVF6e/SH
HWBLyU/x6jDMfAHj7J7OuPph+3NQ2RNYrjU0vhPQxep5U4xWvNeWR/brno5E
TokT+e+FzW5QKKg8Woosdx403pngQcOZcWACnXWihHb5Y2CyAqRftfTV1yok
dgRLZvSGxPjMHorkn4SelcFR5UI3aSpViUoQLCEENksXyBMGVlSmVT1F4b2j
aqBydinOzxMkboUiZ37P69tJqsxJAmQiSwCyg3xDMBnhw3BoLyjo1MTVK1BE
cBYENY/e1sBaaoD1z7MfblEohdLDZk9T+teNutCzN1lMDEDYgasTU/CLeajV
mUqAJVw+lcP59orZjByO8nc+URh70b8wjXFQCcMeGbMy8t/qD1dBR5KEtxUf
iesAj9Wzed6R+k/p3pJg/Jo1ZOKiylbWcpw4xnSzMMq9ImuaErDcBLGpBMin
gNpw2NautdpXEN+I+qZ/H+lU7odvv5JOx4sQJ4RhhgiIQUhf3N4PXH2JkTxq
Vt7FV2Jssms8u20MByAZAGle4Azchrj/j6M0kHK06P9dq0G6/ZpHblWpZN7X
jngXPqvmHDML5FfIKj1EeDMuBfJjm+pXVa7Eblm4Rnn3UNN7da3n3z+lRojA
hJffnmWAnvsgtCpc5bcqIbHv/LFGoo5bdNMoIX9IyAUlQ8nSJaSrLGlGB6oN
3Bu8/O+EQoCNFEMr0ngrVOlrE54qtS9oxR/oCSL0P4ufH4BD9hl89a7DG0rx
CV3DSk738xltGMn+qVpLSE8tG5OrcpcZCsSeLgEjN9d3dLHwzGRkMNQ0NSD+
iU8CtXCrtd2fbUqH3siR0RG6D8Nn4D03C14E91X0BkmLyIy1Oqp3cHaoTmdx
ioCRuEpcwLEKksSveygdKfPKBtHQVBkebANJ7HtZPLweOjuNeiuU+jCxz5wt
g1rAEeOe/dpbLRC7jVtdeCxEXlRNFTJBHeKgVbkxv7WJ8zy3FJlpo3SJnF2T
fj7GXZC8MO4adQ10dE5gmzzDZVJm24YwVsrxfsBinmZSw8mNFWE0Joo1Z4og
lb4+64tROVTjSe1tcyFqmoTjlYZP1qdWv9utw3TgMWkCG7+ksebyUSigE2Jv
fvwiNOY0DI61Pkt54K+3BdberSxuav0OwM8rf3jX684qnrxbdEHq6rKurcGt
ObBlh2XtqpYqsa4AOzspGXH6ZfoVm5BWEo7aeTh9F/n9TLag8wot9FbegYST
ItSaPzZ0NiuwbIQu9zqNRFMY5+CWCeOCt/z7xtEXkh7F97eGble7f8neI6VN
ORGzHbWtH4/y/hPxZ65sKtyI4abcSCicWe1d8y2GO7PNMaovnmstsKKhON7B
vHYUFqHo1nRPjDSVGE4lFkP53+YfrqmmdO8c0BhqeyZubJGwakxMB7n0G1VT
hw9iqVQ11XNVt03epdtdbch94pDRjDmae0WdipvOl0qzNBTz5w9aVYBDPLis
W+go/AlAJSnx/TJjgDf6If2vLyAkaaeKmoJkgs7mWIJoo/onRb+SrvStfm6E
k7rw4nLBbCdvefx7LPlq0LVw0EN3M3h5KhTWrsi5Jdy5SZwvJVQUPlGnXFpj
uCLT4H5hKaONu4HO0UsCscQLcS1jYReODHkF+lBrfxqUvFMY2drEbqe+XS4X
35inndFuKfyGwvxqXliKvOh5Nme+B2JUhIiwtRvyfqKcqMHUEAq++q3k7FsO
Obunhv0a+W3MQPHFjVBYNqXlw9zqrD3by1hdAF3Z1sMzy1DEY5zZLKwSX2Pj
uu13pHBXX+5DC0QQiraMp9MVh6nvcvzHT7KNxBImm1WJ/s2w5wYyVQ5FJGrl
5I6OHQY1GB2iH5U+YtAIraHWLd77swNC6ozY9UAawBg/xK8GXOuYh7cftxh6
8h1REfQC2mq7Z/JvxuRGRnMSAaPBtC/T+gUxTq6SKoQ8WwnZ5/30ZjEghr5O
whz+MpXEmvatFer94A45YRYxzriynqDCHFWg6BNV/1y3Tax724BG1nag1TQ4
jmSbejkCg5rhrMr/AUySJ4RWJtmITnYt3WLOIF7kvQm5x3Q1yIxWy9cYsY6f
g/3Cq8zk0EfDJVKtipCAdovXNlhz2xRAx8Y4Bhiufzwn+gJuIxjW7wVJT5Nh
rNVxCesa2OoQVlygerdiUojMOI/YUrwnotA8MBdArrYhBJh2cdwTov3ZdqHY
1DIz5hB3xujbRj9oFwdMSM1fTM/LxEbcSMdHkvv62tA6JhnjKhkT32dVWQ6E
k1RdBf4CavgLwaO3M6O1ZTNxZfK8kDQ7++GYMTwnl/aCmPh6KncjgyvAQ94P
D04j9cf0jAJGzPmq2teBZtOA6aGBb5eSTGzOkwtJgjXU27RzAg41YTqBgq8y
R/xykfUrWm2FjYFuTT2M21Nmi7wJ0e6RVeb+8QnGf6X6+Lpcbzps1wuetki7
Z6B+7/2y3LTjQJO1eo0vUmdEdayvxgY/n8XmrdfZeFdnD4lyfaezNS27dBaK
VI4FyKQCx7QH7iI010Mp7/6owxswLTxsu4TPBTIA2PneucBe1RSlc/a7ij8M
x9T+0jzQ5+ghyn493lLaHQ2Ybg4IsoedEOaUZsz9klxIOIG8CBf6yAx+vOxA
nkVPJRn96ToWZlCu2kHPcFkAg90SeRWAi13Ch15xULBUrlIZ74ywKA5Cu9uW
0lsBO2Ap2wJH1ob6oyQEifjrhiuHeZS3Hqz+tl23rq/aORC+86zz2oyX7ep3
UL1tvQM850McXyATQFtGTHhXJmoR8r9OHJ+Ll08QeFjrf3aeFePMG+Nu/lQO
h8Wiq9KIXzD4MVdVo0iLsDTdbD4jJC5xCDauysqLusSDft+Piv1mnLm3fd0c
LOvLHFqUyYSWX28nB2AnAoZC/ZP0DB3VCAvn2eCUcNe6j+yNUu5xQNU/7Ern
C4cYqsKL5u7q94c8yhzmXTrzF8i5u9tbyLBPseSaCPFuo/Sjte7T24l0y7Wc
zDJcEIIu/byXaj0nWHwiaqPAdpHKMFtcQWyGwePyVEdq7GWL4fZgfwBLQtOx
4D5qAeOl1JjJmEJ5Vt2NQPn0IbxuT2xEvS7cV6XpgRom2sPfMWbiiH37LF16
4dznJ0T/15L0AVYVrn2ACsMpzBvVxcDee/KUvrWkk7g3MrT7rYfDAJZgFffq
Gh+V6JfZT1eDaOYh8m9zoe28EllSlenm0yLVF8pP9M6KA1ho8j3vnqs6hYsj
khbOo6aJMrYlU2rEK6rFwmYdT5/Cwb2OVDOTEmGUJvOKlFusRGFvnOLc/EuV
UJS1MBnwJMsPMTakNIqh24/21qTcYn5n1QmFTFdBBR07s0v1f7bidKzXt/kE
HcWV1/0+5+HedZPKLVdh4EsfHRgabzncprKR0pY02fp8SBc+1ZwBYavBhFpc
sNjgxPVu6JtCrv8rgJz4bVzfDE2jo7Le4nHflaY4NzVw02U/IY8VGxAerKVH
VszvW/jRK4H2vzHHI2q+HbDs7A89LLVj6TogUj+89dvoL1+2lceifhG5FcEV
s97q8XxQtnRvas1RDdUpYgbH+YC/IS09GiYZqDZP8Fp8wdlHaptMM7PeBLao
7nfLIajNL5UUyyfo6cyXT9MOaOmHwya7+Vd0WK5efH3y4xynYUe0j0SMOMvv
S1aAG5v+fJirZY763mc33/6fbhRIQUVsE2eBk1vpDILIwpsZTQvgey1dD/MO
H0tqzLPvLChMagnyOK37QfpVn5ZXxk2/dGhDkH8VKGnWxGxTzs8yFrivdzNX
TI1Mhepm4CQdt6HLURcbbMmzWMEnBpLPR1VCJCO6dWWiWuy9WOuco3EUSYWT
fmx1SYX9oGhu1Bq7yGUd6YY8dQJvZDXP3RIaf4bopPkGcbYrzIPdFH9crS89
3q70ryNWazi/u5lHws6KCi7Pw6o8RBoGHHQ0ISvAfhYs5xCBdNqyzYBXRyvh
XxN/W+8KkA+I0WPn+nl9Joh3K9ffkSocQeeUfdAp1SmA0T5K94A7oEgGrxSH
7t/2UKC3mC/gjSF7F30ZH8Sk6MQSAWHNvzFFaAwG9SbHuGI5nHhMJppuS6f5
Tll6hXWMWPkUIkIX/WMIsaG7glwbom+IHob2DtF3jPthkXnbxOLuxjPXuQdy
rwPp2/oiOczmcGKX7QjSKmhfjXOC4dAW2X9LDhMd95ZgIAL/UjtkwJ671ta3
Gu27cwC+Ky6w3iTpWuOk20SLRcA+JACxmwr8YkMlHyfjhQSVJiEvDsM1K32z
jCFoB4QKiYUBvWt9mvEYrJ/okcZxQF2vaxwzrhxI2KgK4Sn/uj8KjTt1wIRM
gKjD/GZLOCwWlmMF3ew+Gur5CHfUEi6jLUq+baWRm7pyVZnmQfwRKMC2SFtz
QzBycLBLqvNGFuG9UHnWdIGapf+wtHrGNP0bi6Doghb2fs3fAm0pDxG4OFoa
EkYdTnKJDW7/jsj4GPLwKEclu812dPbG6uQ8lfWr3L+q8SiyrYiuLFD4nBM6
nA5vRAZPqszkVnneWirSJZh4Lx1zFIKexT5vT42CGuJL9U8dj0jDDtNqiLvt
XzCJK6KnkKobZevnRrLP9ZwBpIIyKWw/4BxK1TP7+Ju/JYs6hqi2mwvd6zQX
kVvSNqbVDoVkLLys4+6jDSPWrRTb/qRhmmr/jz3bNCSq5r06EFsSFxutPKPS
4KnE3+S8Zb8MG+Fc47HocBvXCBfSzYyYZbYzQ+VUO2YDhOKX74UoFtXOfH/R
TlVmbl4nJ9OMxJxw41WRrlWjJx5vvH3e2BHu8nIldeKC20TurxqzLGgR6n/O
TzdwaWwah8vAnr4YfCUR3bs1I+Uk6TGBy4qk6OM1A0uQI+a0bBt2stMdcoBY
BXi+SxnPKLLd99skLOLFqgypReDuobn8HOruCJsNAhiJ577D08fSUger6rb3
Pi/ap2eKn38jl1sSZ8VhHy+jun37EhuU/FAbCj3OixZe2KkO5WCyBLUpt8lP
75nWpxgKLek0AGwfjV2QhtX2nYT0jov4GQzCGJXx3LojkjChm57N1CfNC+ee
zELs/3U9IuHdPNEllT4LarX+i42CyaTyCaU6VGvf2u9btsbMZBCex54e4dLu
pErP5qE6wOMxK6hHMDVx6c2UaUBMFOY9V4vOw7esZnI+OiOpPkiKnRm5UWic
OdkVEw/2wQ4c7VXYLeI5ELSLweArIPzFDmx3RnNk1TJdPp2JqTRXu+POmlxO
s8o5K9l6EsO7mwsJBoFqDKuuhtJNzOQnwcOzRGXVS2pRwEZ7EXRTXfRgV70m
pL/d7NexDEcJawGKiCMkH2opx+k9RAdzPP04Cp8vQUP06skpm0P4N9vzFBv5
ug53r1wPRYuPWU0egCzJZ3swsNAvXqojqcxxgPZCkDV9pqTmmOoDLI1uxKEh
ZPAyoT+eCC41VamohecNQL3E3yjogd1lLXAd65zYtDXWlvGqezI+uug3BSkw
756Y2dwSPE81j3CczO6uivGXgzBQOgB4KuORhMb6KRDbfT1eS2LjECWN4Lw1
kQFDlfHe6Rmwv7ObCSWxlhEPtVaZUDGviDltoBea0QZ2e74y6watzStlR1zG
iopJ3R7+iUoNfdfk97rLv6Y7pgguBFRokQRpNYnSEdJ5Fb/XA5JUlPvt3NQQ
n8BXy+mAAvNLCwxADJ+qAXMkjkL1DMghefaceMUb9rPd09KsPGDsGoblvyoP
G5y1mcyYVB47C0O8IdfyljLTeRjlwAqGVwoBj784e39ucy4Krl0JU62K3SP9
tnQndlimwCOL0SWk9E5XaHFq6c0KXxPciwC2J6FmIXaVZCLARLwr/GBjg7u5
IWfsCBci9gsgiffx4QFguL2KF0XA6/NpngNHzl2PJFAXOQ2sEiyCcSVDto6X
Ux10fRBl5iLejqP9smcQhW/milpZWoDTXwu1H00uUC2XRxuHVg8CikJZ2mXI
P3J0c0GduqQI4qs0xnuzAJiv3hQSSUByRF4uVDUOa/g1sIS/qYU5XEswDhQG
kCMuv2G/HH3o+/+2Vwa2bQRr66oPQkLE8FruackcxeAtUAfYM3KPby4xjgs0
Ag/e/R2/tuCDyq7d+KDoZgo8157Wx7tXb0DxHSBMwT0xLOtDi7iXxV1wMZ7N
ZjEGLX5MEXHnfy3g32+1zhsF9Wvp1IU1Zb2Jzu1lDvGnN+lbz6DnAVGcZyZI
2SCxbpDLPnbK/OMZNe1yNl81788m96edqjLYc13aIYHA82SmZ5/OJSIyJXLW
Fse/7MxEuph5+AyOas0oR2bYDk3oSOyMHC82jeQ0XzSgA6IbtuOG1cfYxKKl
pjvGDdk/vrOXaxMRGdeIy5cwk4cnfQvvj1EOPUM2Z2gdR9RH/TY2zq2rlcJE
F6LwM/WI76a+UvW6bcf7wr4Vk0KHbxz/3YDqV3Rne4eqKRNZ5eeizBQL+rO4
uUE1LyTLhBYV2gABjMS+BEIp/yO1hG6XydU0qZt7KxQ41VCVqFPg8D9qqRlN
KtfjT1mbWk0jF54Y888Y4S+2C3Nx98R9yAsOC5wgVZpTTlIcycJdYFomGi59
Khey/m4rcGbu8xYjRhLzWHDCW8P8+/JCZ8ZPaVuEWyS5gaKcSbOqG/KPtEh4
ePtiieEXqy30kT6MSjfTaCOoyrJ5/fdlF1xnnEkjfxdwt6PlNwlbZ9vMAT4E
s8R6R7Ep5oo/qZEJ9ZEnr5fNNpO/aSGOa7/B3Bv28xt+MOgf8wSQt9YVIeIQ
3aND6wcAKrUBK+jXeqEbs2fHFNo2tg2RRkOvCUkq0BIWWPsJks60xHojCbN5
rY4hC3cklpB0FhdrsqV1p+jieqSF8GOnAzORLjC4gh9zmAD/ef+epqASRIEK
H3oYlcbQaKmYfSiHw6JwIhMGRGMv7MQUKSZ+PhJxGyuXCdkOYFnDtKfiGR9P
sfbbGOEdf0YorxlWD/q15wVrkq8EtB/fuk61T4K1w9rL39GykCu7hBnHqnK0
+sbbQyZbvqwa7RbISo55Gvcb6msVzyooWRXjoLyTxFDgIP9Flh0A/Ib6rHmq
lp6IWAxBhFy55fRdceOssrBXgEjfnStaAzVaAphpuIHG+jV8P8HDTYRk2Z1w
mJFlqh2JA6Vfr0Tjx0F5wggQ23LoUBLcLZvreSaGbIr24KVkTs4gCP/+37yq
hO5JkeQdZjxn/tBAIOwttTWeN4x8Em5H18ZxZfRSs/6xRf9ezAQ4WOjHhplp
V4wj7E/L2NwPc5jAzXjtirrWrXfaUKofjim0CIH7qWKBj07pjdDW75NLOtqs
QdB7ONMPf6r1PH1C8XVC6OP92k1c0r2dTbiQOR9Pz1rTb3GdVeTBpRnctnyX
zclGc6sN5LCUm23xgYN1H8js2hg3os7dgcP2oWYogkQKYZkB+Zb9cGX0R7f3
vT91eNKPcyOg18obVhoihlTYql5lBclwgIBcpoZW2ALgEQzuxpeK+TJxTTP+
DN6lRAL64sytEe5d8YUNPjhmEHNWj+BiUumZb3h3LZ/SkLU2k0EYv3pL6EZ/
B6eH4lwR2wli136g18bQMWMxFRMVogalA3Rx2iyE/S0iL5IT4k1B5e24Ag0k
AZhjx7sGfTD6MeI2184a29Lse7NHA+P2Z1H5H48ldJv17xpFqQbdyNSwQUCl
Og8NZXvGw1FZWI49DIqLeMU/7JPRWsH7dBUn2N3TcZo9I5BcM7b54AFWbiOF
siaVv5E3XWEkHk8MHeVdK36wxPSxIU4TMQAWwK04Y5L5n40eeTVVJvOovX/v
EZnvcb4z7gCL/c3LZzoGpml5VSYK7PURA0reI15tgblS1dWl2P0rQx08Zs8M
iX2KoX3Ei9SqXWE5M5O8jW9yx/MjC++a+mg4rNZhRxdAR8BlarGZFFtsFNVl
VbmJWRbR9YkxAaU3v9vZ87xoVryRk/66oexYjdBRR3uXsF0o7QUJ34btVKhZ
lHgUG75j1CNMxhnNCaT6CFh8/lMqpzV81VqV+aggF8HC/ZTGfASvlLFKc+t2
+8cvAp45p+d6cvdbkFvqSzYpu2Ohr4WZ0Qhl1ZQajc//IUwO9eet7kRsu5Lr
z5Pk3szn2ymREMI6zwnEgFEYZYEFymlF2z3a6VkbbLqlbTABntWcApn8fVtA
xJ3W9rV2a9T+FvHLUf8xY5henKjXY2FaLGqbVtCQvyjb3mmXMiA9xlBo0wV1
jPZaSSurTTewLfcHxu7e+1PB3h6oz2XtzbBwS3eisnxU7mubvxGcODpU/seD
PyTbt57PKjH6Rhhfdkb7UE+D+KoS32n5v/Ddhe273Kt0J2zM7TXeE6HKCHDS
3nBs3T+U1MSDpMzGHtccGWYB5ktC+WJwNnzwUaTrCZFFtFEKfWp25tKMLkTs
6jefhI6vVCkIvNrUADwzcLyckK4ZWXTcK3uSAi61IxtTEAqxgFUnLu2s1s2U
Y8ri2F/HluXL0j42o1iho4rsq498xGipF/kE1+7QFsW0MhXPbJITT+PGOKe5
WKUQAg1QSlthASXPThanueCjUPeoqDwnAYLbg5UyY6GhJhOcfw/uu3PJbquP
wXJkHVEjN6AhkaCBpQay3PDUNlXwEwdDfyQluBsk5RKTDKmeUnldlLKh/rOo
vTP+VF5rAj3xJ5ad3JQzEEj4FuTAHnDkTjHXz1/JUe1Q9kXg+DFjOGb2ZNdm
53fFl2CK72GtHzmUzRyuoCqD3YGR/QU/GjUZ3L14DzXEQOE5gt7qJ/IOWhph
dzs6KWdQqCV6E11C6/IUuNAHJHxq8RGjbjgLMHSkpQLeS2Pg8KR5HY69wudB
tV+oIQewz9p2xNw/+3noJ+txjJPVC3nwsY+9KOvW6S9e030binOz+HB28V6r
SiQok/k1y1U0H1SkvZrw8J7GzScCyLdE/myOK561Of7afhLa+nDm7qjzI2I2
uRdsLUFXN+EUovwkVOtz37P74Magodkd2NWNe/ZGbh0CzfMZBtylnv8f2fbw
kjt8uu/tfTKV7BmM5fyCPPTq/sdSx0Gz0H1Yf+FceU0C2Jl9+Nw3tg/O+sVA
IW0GiT4Dg4IeQ5RtBudqqhYvTS99WP0o/35qNsuApDOzL2jPEgqGPjgs7GFi
wapIhDBVHXljuFA75t1bzkJRTZm070n3/BZzIwAzi6WjOvl7Ni5CXah9Cahy
2/8KIDU3rNe52oCOcSzOFd45ptNFkpj6Ke9qKfwU+GyS9MPK7C0IzV0LidZ1
ZPHl+l2z+83JfEAXBftZh4mopa+Hnj/uSO2EAoqyoe4PGl5U7ytdZl+HP0+V
bs7CGsrUdD7y8KSNBxQttpl1z5I5V6vZypLA4KGYn6Y4RBc41H4Nu+Gx3hZM
EpyqNn9LTpnbbn4hCkAoCJWyKuUebtdGh4+5qReIDUcgXB88Nwe5wSA1LC1O
V8hwGNCFjXclAmlTrX0lC85m+zUtEVZi6TzA7/PNNdRy7GyjjwzqToMU2Ygy
SGa8ANm6US/tHtQ/kz0Ljc4Zqj6mg5eHptpyAxf95QSrK1623v4Djgz047Jo
6HfEGBGcvRODq47m9MwFJXwwq96UdUZ581kCywdJkSCCbAU//w9rYSa+QMs7
TtdJpt0jQF/yko48fqotybHi0e/YrQR8K/TTtwItRdRP9vIWl9/CC1u8d3D0
Wo3ua/11b1r/e5I2l0qxYcIC4N4ETYXmaplYwxP/nRrAoyxcCyowTodIvFFe
HO9tFuF8CgZzUwkwk7QymYXDFXVqLFwn79UosMqfvPrmAalymLXd/eTXpgTK
tNxDD0mdn9ON5zy6ILuow/B1mmtrgVqN9rQPHEXeLuAEmaUtzMFX59qcPBE0
XLiCd58VNLtW1pUbXeoAf00NM0yRwrKl874y8aTIvlI54WHM3JqiJ5WwHFRZ
wTNHqpwOyWQsN1ZdDxEgPCnmuJOvbAR5+W9aTrY2zkbWBU7FOd9F1BmUOtAR
tVHq3nWz6CQxFe+KMnDxotQ1Oc/i1WXUQ309s/erGGGG4B+3AgwRqnzPaBYJ
Hg8/nzquWrSwI/o50X0yoah/hYwA5CSqJPJ6ErZRo2t5hgBF+DC0JTbyDdhC
YqOHPnw0tLQb0z2VjfhgItFnYcVvrb/GQvM7jKTArwaFki7o8sTYNRpSbIzQ
O5+nJ0fL1N1xYLWJCc3VJ+UEwwSrZZVICTIG+7gYgfjSfmp+99HKJXBDqMZM
v7ZvpCRywfNbEahRAx9HU1xGEf+r72gJ+72zani5it7s/MCjaXK/Rx/qBUrV
w89j4RbWtm9zu8lWQWX1zD+c9+KzEqehcWlMJYOExyP+R50ikXT7BGBZatFq
v7w93nbkZiBVruY34vldh9nRutsi27Cio9/wMMikOdS0HjtEsLq15+Ako+Yc
KX9n4+DlmVlCxvIVDawMBV5VM3hb4cqLp26SbYNRXCKbg4eVtQYQl2gYtUen
WVMsdCCI7FgKv3XmyA47fcxKMsEx/MTgmSetaVxoFRS4yPomzjQP4YSGpVnZ
AB+k6aBnnE7YqZcLoLs9w2VEZfmfRu/Z8ve8mdUNOkZIgM1YOYs2x9k1WIgH
M2dfXNqX7pH7y0BwUx7aB3n5yrkjLBsmg6cj7GNMXwRcKX+sUcg+bZPq/VCn
VkmSk+oyyRpWSw/0inu1MKaIrwytqrI8bKAyOV3IupdG0Y/GjOILaNpebxuQ
pq5LpSfM7F8UO16b+c+rIkD//72DmI+vE2uMGvjDfEAMu5rns7YZg0W9MqNs
hDW4zPcCd+xuTwo4uS/q47zXamh5ensZMjABJ0S0efvc+SWjhpXchPgdxQmb
SD146+4T4ZwEpS5q9tOcCCFz/WvgBt3ni9QmhVGvrk1LQWdbOu9NMK2cEaRj
gei2ASx9DhcxOYOSy2K+L66vLCfaKKY3aENy5+tsljMy2YyGfH5Lh+vweWBd
bvh1b3h025xfKtn4uIUYeplVSivs86mZ1TtGC4NI1aRCJXBhdbWRlnIXVQkA
v3AGks3WHgw8LR/MtjxROIXl9Semb/NE5t44A0dATvyESDL1tAqXMZ5YcggB
KjsbmucaY1IKuRAKjdTTyxMtNH263w2HRgCwP6UOh8Me0QglVf1l01G+uy26
zt5bBIUFWfwTJgDgZpV6A/XFgh3tGfcUbeCAPCqutgeKW0wrJTfd9725qjgJ
N+G36EpE6wvD0N1owxeMH21exbdEfaZ5ok8fOA3l0kcRPCpjsI5T474PY8Xx
kXZ8iWp4a+KDE9zVvkL/UXXS4+GPipsgCdlwJlkVAhxNxHnZqOiV0O/CrLWY
zXJ6MUVlXEtT0RInVI1hzOhPoOgn0jgXAcGZ+LaZNJIZATlU0LuBYWffzE7B
BnCV1sy/zvwRtssqUN004BP7kY+9Ap0mgVVKoXgAl0P+ky3TROy59woNkqK+
YOfEkM8Zk5WzVkLmhx7MbKR6JEjbROTiXyTVbB2JFWcrtOQEi5T53ZH9h/qk
SrLhq7alNhvP3a3yK6+OWY0wNwB90WHjtvOGXUNnV0l11fX8VFAxD4Wt1Ucu
MeQ38Wew5NlDNCdewNO3qXKcWXneiscI3XSRsemUU8Kcu64YGXSZAGu/kIKI
T6cYwqpmA886aeFunBFBzh1q0s1mu98eHR2Fmlxdfuy4lUEklKyb5JjOtM60
D2KpU/B3BXbCiPgW7CzY+J0dAEyXjagXgUQmae43Yps/WNupJtSanFc3w5HN
JHPDaoJGsvt2A4t3Fiwgp/G6ccLjVlZo0OvT/QJwakKqrLtmwkHIoPsQM+AW
Awk4nVLMcQwlS34VQSr2MKC5yWylFvgejku1OHAtLT+ZUy4l2xusCjpuVEkG
yVwccQZkfGbH0R8EzwENA2hA+/FcP2bHw2sMd5GI+T1Mdf6BtUkjUDbn9jxj
qnNm9ducCXNQU3gx+yl8ZKSVPIb9s7tAUBKIITvUABRRY/a4UVsWwmasBt0x
/4oNx3eYVh6czy+b6rEkWAThzO+Ib2U/RiKc9r3lb5/u+5IDzc5gnzN51pMU
ciBS26SjxAH0clnUa4pyeCkRpyTJq21GZRh4prRpuA2zoh+8/ocUNVhug/03
bq7+6H+ZAQIUCV6XZMjK6mEDBoaMtb223cQ5bA8ocy1JxUheqJmBjDfFHzmM
LvyZeoQJJF3zHcFm1UqRFH+oVTGG2mumVPV7CFTBt2pij9CtqFHrucSas4yj
7nsR98egQn6w2uP+N4R6VKUCsGEv6db9GzYx0LPCwX5+QNQEB+X6K+u6L5Pa
RXziHdUk8K4yxhnSAU+U1NEKurosFzmeYp3O+hNV/e6og8fNkT+et+bvx6kv
JHd/xLag1BwipDYU30Y8Y7IuEuNcGTs6HRL9xS3cn7Gc8H+vAGCpneQl6Bv+
JHXyLlK9Bdh9zjp3H5RYlWvd884TU2akzu50A8Tkz3cfc9bT8njVC2nsXB4/
Ln91LSIFjjSL02lDs+Mz3RTnPzFL5mLWwZEs8Nx2G5wff2enHyvuk9iiTGKq
n/+HhPkdZs/kdhoHRwNKJoj6tO/G8/12R1kyaUtsqyaI710v+y5VnyiUtbUh
Vla0VL2uK9r5gr4lNI2picTy76U9TiqRljXH+HUq/HGrbKMItlfE2x58gLfB
UKSkD2ryCQZ5cj0T/XkHi8mcVpDzvsxJiyW+epEODYEzLLAFTevsM3IeFty1
x9yr9gguryESgdwfs1qXkk8IFi06Pht8ITQqvF7rR75VORaDltq+iL1Up7Oc
/vqGmyM0pkLhkZ1yYHxBjyPBYRCfyXcFbeG7a/3V0wusIf2dWbn+5kTdGYTC
os0oYwIEoOrN2ZCm2XUcj3zX+6mvt4+v3OPEq+1pMN4/201VWHiUmkUZX7bB
LHTIqxvSsYzDZu0J3LEFNMU0K0GCIo68DFgzUgC75IP129iGFF4KxcgNCKeM
xrFBww9PPbZ8QJSYbx258WNRCUhrINWRDLHcESBLlSNYrEbFT6F2idcOfukr
Af11jOtvRiMzJYw5MahvHSmlD1Zq27LXc0H5jUnE7SRSN15NuOjkuPOqohNz
w96flryXmjys+oCffjCyje/ksY8EHSYcfHtlmlVsOtpJIPitMM91hJzy0FNa
3Hae0XRpoCAN5qvmPuWqU+DNSD993ZnGnYVzWIfRkaWJ6egSoHfDNWxhcLKK
cjxAPBvZjIaj+OCyQiEnnF+q7D3Q5+sN1l/8cd0Zlyrzb07ZBxl0IK9RMgB9
aTYe+ueC0w5WsXR3KapjsH/oloIGTYGXStE2NBlEGibOn3zg3QRFxKuZdjhX
XDmAaLjNRfMU1OTBXvSO5+PENVGFyNM2jWLXQijDzuAqJgHOD2EJctE4HkkQ
qcIv8B58Zvk6TNpyPFTkNEFaL4q2rrs4BVdSvaELtg/sz/sQIRMec5TzC5xz
7p0FOi6OTsbpBuDv7irVaJFD8x7zlXjquWVaIqIMOe2Dr0YWErIoeaE3z85c
AlMXuWZLAc0a08qaDg3N015wqx4KNYVSWCQqBZBIuyiNuz7cJFLa5yW4W93Y
pdZbR2BTbuMDtwvBXBL3mvmODWhHABuMSGew8GI4cne0MgiRLyUibitM4dwU
1boJDJ6idkCMZJwyGULTZ0m75YqXlJZ8YkYBTUPem2H8JEobrhYgHMH4KWvM
BRwzbt9q9SgGwQ8Js7ArfFD4zRtMgZyKOXm5nMiLdByWZrL9O+6MAK+geSGV
Z96TuSJp9JMN70qeJE2L4XR8EbN2PuDcG7AklYRC6pgNLXciMvz0sGqR1UgD
78oi36VJIwYiX3j+AmfvpE6pXgAsz2GhhbmciQ0tvvfEbWvKRb6DYSr3fTbl
mnEvs7Kjl3Egf+1OGQKuEwS7qAK5n37PKP9uRzOWJld/ny8LgFzAkAVl546A
3yyIOKSZW/r+9hE6eT/azm95Tr3rPXhXAMB3U9xSjXfAVMG2ObsaRQgWWB5L
4De7rfzWQM84dMdAA2/9uvW0VZ1ra4fxmPI8ApZQpsDzBNwdKEl0oF3Vn/HV
b8ovTE8CHV7c528cSaCcK2dBwr7qqZjU9+nF3aWy1GGsdNf3Q0PVe8rPF5Zl
didcWkHUnFYtJbbPn75W9ey2+IipwN7m/JUNYx4+8gK+htEpBgj0TRlVaelt
FJ86vGOZxXrhw13PLH99q/BYI+NnKxgATThE2Br3Ej1no3JHmqssrFczw5cN
5AtZpsgv582AVfqP2gDeoj1KmFBnjlEwDI67x+Sj4hUYUDyfW4WaXcR0uKRG
QqnnnUMyyVbmlydJY0NY9fjrQ4703IezHXoTUBMwQoAo5bxOGNWdOTrzObVL
F63Hh0DamEAyuY0DutUDjMNvIB5hkTto+aBpl8B6+Wbxnj1pjpnTpooWgNG4
w3zNaWobz/3tfBbj6WqQ+/U/YQLitt14rWqlXJF/vEM5qrPeg4WdJo8+yrv8
b8yNKG+wttMeXyVbtkdDm61yHsXFjcAEZQPSdjMV83CA0eh1J/xv1RLDeL/y
qwrBGD1RxxPhXaUjNWrIxPDAxwYk+ExDf7JEekse93qBuWSrUQcthdfPVCFj
LHJANn1CmbXj3ntPO+u6ri4VaWrXojGHMKRh48O1zSfM9Vez2jREhXTzYgUN
wG2+P50qTCFaBCF1eca611eV48R57zfqWToR4SakLIR1Sjdm4ZVoiNWl72wx
M+F7nu5lod0NgKs8q5NdubXPrmwJbRD8iLozDYOUkxUyfB4iJgaSf1f+zbX0
kr6y/BKHTBvjPbjd79yFrg6CInjcf4F+ecqDnldDifCQ1FriOWohWxmOQkOY
nVUXtEyd5mvXfYOUct3xhkVpUEaVZu9LR58QQQ4zMjqHssPsItcCk+myS1Zs
pVJVvXjCD3WAO3uJyJeLUp+wMr4rgKCLY1qF+Ja4HT5fpR+m7vcvuOim/R8P
Puv8+9HcErbYuIg1NzTOowHU23R96oXhW78EqxlL0BBWB4XJUD5z0gm7g4xD
hcvNS+rHmHvL99gavaRSKpmTaPHXCGwjBqjVPDnwx7gnjTMuFVRUKFKAqgs2
3VQ7ILJt4ZNQBaL5B5IQlQQV27ACsYROCCbMxX3PnMc862UNLZ11JaGUjK3B
RKL3L+oYPD9M7985haWU/sE3ov9Ko2Er6/yKwT8/wQqKevGEMJbhB4l99mWr
cCL7g68C7nM0J7lGwCfrPtHIKtEmOsWnkQmlz4B6iRw9sQml0nJ7J2sDubNi
eK6S+XzB129kLU7AowcyjCjdTNZJ/Op5WkECrSg+83dynlgHJhdQmOr8kcas
jGdLS/ggdL9VXQvZ220tzwh0TsDqnOk/eJpUctD66VLlnGhugvCbh1tk3E58
C6qAkQW+EMeQxcuGYnl1S5hu5OUvT8ybfKsWS1UZmJ8EvzYnigwUQB5avY9L
e9AXUQFVSOKmrCKU82porcaa8pou9aW+YIbTxRXrY3K0cp7h1x+RhiCb8myY
pfMQy2wJAtYL312Ju064slYPKQFqvX6ENjGgssc+xrtQOoljYZvnBIlea2Wv
pxJj9FW8O3D0vSlJUjO5x38/a2asxETFIVsYokfI5jXFkaIxfvMf9Y658gHy
eYc4/Z9LIvFWE6p4P9kHM4nnw5KAETUsNYUgOhQoNnOho/GLhWKrZYMhRsFh
0W1rNea27aXMXcp32zB2PWaS+oK4qIKqtOqOnfP8j8xTXhr7fBiWnq7E0yKL
OGE1X30uNubsSmFsYw5RC5IsIHyeq/zQo8rUM3e7CHGPE4q9552kjMYJlsp5
4U2KuXxElli0Ypngogp245T1LEXaymCPSHpzNyP50+zmUCtLQwCgizEJQ45g
3Nn/3ybATjIbWs8hcxIT+86uqBmjHs+vkDPtwCWLz5o7kW10oF4PxZVJEkuE
QvgUdHwAukmeiTQbXS9B/ws30EuwuhMi1DjYbHVM2JQoNz/e4SMxFRjlZcjs
M625DEbvhMGRa/7VvK+hSO/Ta6ldrOwlBweIpIqptryP+ZjIwruIaXqsocKp
zklRiNaF80mfbU+mvxHrHQPhYRIQ1bm0y103e/1j3nzNWpeBkmObKwgLFG+A
6O76NZeWHwTXbBcRkceGB9bE9FSyjpV11mIUVCr1mrVTAmInmiZjvLDsDBwV
EAc/1mRcaf2JIy6Yuy7G3zxE59ZlzOsJIqd8eQTo8kYQ9cyAXkOi2Rd5l1L1
Fn200hS5W9YwT1tqeakU9cAV2ZFwqYVP2N3J9HN0tYwFZ4ZOxGZ0q560kUAJ
0hmTdbCH5jgftcy/joenJCLXEhLsM2vj/UdTjKG6IFmNpZK7RCZ45JdlZx7J
ZSajI0vWSh6jeJcs7I0/MIGfJQJtu5syVOZm6MPfuhyc/6k0OKGi/7v4uV3V
+fOLboYmid6Fb6GewTUf6sqokm8+KG+K+rAxAk/GtvYJoxH2CPogo4qVZ/1g
gs0NTr6+Nm6qNjSCsBOEqh4Xn5eyVznQn9bh7RNTl172GCBkkWrpiNA5Saq8
wlX3g8759PF5Zdl8Yip36t98uF237k/XIycMoVJD8WI6TxOhTcGdLxMHgAar
EEUG1hPvbUj0KE4GlRvdYXeK+f8DxhDSPwr26Q3PbAVk33b4nvaafkjompcs
4Y3AiR4bXyoZYjDDnAbFN5jzg6UgaEKuHKi8FU1KeUmCP92kuhdvfXj6jutJ
U79w4PTjs+hcxIs8QRimHnSGPX96s06/zCpCbNh/GT491DoWNmpucIhXDysp
2oetN+h8+IuiY8yDUJiNpfbu1De9PGlkWA1L587AFrNOQfu2w1Kuez24fI0x
Rhn2kUISFSE3RBMlNgY2ongKKpZh3ZTCTJthvFOqLFD4hajiJ8BHQXQQwkoI
NR8n/R6DYSWLY/DmU/TOu3qbK6ZtzXQqX0Klk1j3xnbajg+f4g6LmYy5Opb4
BhERXkhHVXlria6VpXA5ysPsmSAWGzgHHCFj1adTEkrsuD+4jLjmaJhM6Z4C
Ty9+FwVe9wb3NBUWoggqr9Oz92zK9fEEBdy1o6I0a9EgRthey3Y2/9NQw1KH
lYuHwubquUjVwvbVE+gjl3CkzcZP2fxO7VQP76QzPn7VKSyZiS09LO8TBBdK
CQyEHf3vBjmc/l5IfYReKK0lpoklULcui+qQJILXLU5MvG5BmX2/O/QO4BPZ
YlYXz1+zRey7W6ngvLp73asUS41qJ6DqP4QElP8ANeDRiVe4/v7+ROxtbkXh
kOUI1q/sBksDH292OBS5JoQWdQfY09w7s/ml6FkfSEIKvt7nv6apra2aEPhf
pmi7Xrrrvg6psBFesalfDclZCELyFBffwNOokVgc1ZkMnE0WIAlsgEmEMv6P
MzQTh61gM+fv5su4brgEy5nu1Rm6nMP3JbeYf2Ho/C4xD1s8r08WbSVtaqPU
m5HDJwYwSmUzJj1zfI+R/drK8XuXo1oAzXv+HMF/ABbYuMO/CCedTSaqXK98
e8iQmiwihb5XK/yniPbyQexzZp0huDvpPvH01KpZE1GksMsJ7b5nuSAUh/eD
yRbNPIRxta2IkOKvK9HBAmjfo98TrOmwVLo6Ap3A3hN7Z0dBzZeIBYYPghY/
Ko02ihYf6hsxfXC2wYFS0jBT6vnbKq5+T0XvVSvIpP08gmjnzVPpd6tb59fp
fFq4D2ga6EqUUqNUBebvz7FA/bD6GsYALfv1iPoFrNBihNsiSSnAWce65NQ3
REpI1T5AWLtU3hGwsj7b6ubqKvRagOtYJqYwb5KJk+Y/X+4MQPlVKPxRr/jH
cHrauIY/6sWLVNtDd0gAAsmN3W2UqvUMDeRqcKaL89A/ordt4mHsQJzsuJYS
oGdXicTrxJAv0alPy4Cq4ui+UlH4L2zmE8q5Nza93hX6VRHzOrZiKeHGfrJW
kjT5BsXUR9yx5W/NOVoXeG5QTKTGKzqPqzgk+qv87ZY82I+s8s2AJNRxuR2T
UItwE5HA0WkHgcN1BHCk70nkiuIBrsHkkdlyguParAIH5ekOq6nLXehVg9N6
j/MhBw1xUPaqTba27wuUD7obxI8j04s3IMfUwJawGMNwA9qHa8I2W+k63/Gv
SN05+g3t6z+MfT1gNMDJVHDnnD5VB2+qr/u7xDklmzxDDJ1IFybulMiD21Om
Lk7DENdWMEunhKXtkdMSxZI6yJAz692IPR1HT1rYWJZb54l8mX3QW5JKYA7Q
3HKe72QWkN4o9lc0+DHOhUH6NN/U6tS/wblD9I29kEwNU5cA8OTViZ04PgjU
XaFjli6t9FW26HxR7/T9PJX4bakJUK25a5SeA/JmbSw7Rwdwy1EmNSCTuV8P
BrzRcsfIm0rGUk413V/I+bkEMxVQ6b1ExhxyHMQxC6eOYpbpjnxIvM96yxgM
nYQDcOwpBlPm9t8ewb/4F9x96c+b72hQF7uO55Epn23Dfy6MIZ05SmEo3cHL
QGTVg63ffz9H1gk5rPSNHvE+jHRCfq7PWMwYl5l3Y2UWwFeD7/Dlf+ezoh4o
GzjgF+mBQBs5zWnptABrY1kNd6aSPNNbhA1upP2ufnf5qUZsDLD87x8Ca/38
dLsHCs1kdiN4zhOOoBKXuGrn6S3nULaS5F7o50EVDfBPkkmlh/XK9RiDIKAB
apl47S6lqqKnYf4TvvT6c7K5IKBZw9kc5QI6VYTDvs3ZAkQpVwgm0cT2qXsT
ZToPCDuDdN4AgrpESOGDsxf6ay6g2EFWwzlb+T3+qAOVrY/AXiWrwcwJsAeb
ktiuyA/y17cjnHow2kSqrVItJAHza+lUsndYU85KjJVicPakArXYouW8RBnz
KejberAhCrgB+ALQXGQXDf+tlGfTkU9NGHUlua6OpB/I5GsSd2kGeSYpEXcD
0faSqcpeShD5v845WHw5xFJiPT0J+t7OK4hdUD+EZ3IX1TUy/Uh27LY8tfeI
yifdge+Tq0s20eEvBuWwXqic7lER/x/GcUNuYxAsoyv2U4XwH1oj0PPvyDW5
NrQyZJE3R9roTwNWSNziaOGwRtTveljuCZJWhWUrvivSsyV+QdpV1iuPGcdC
oODJdDvyWXqFN2ZKmc7H8Q++H1KgR5fyRmSR6138WVMaEwACSK3eK6ku/U6L
JHPJV+NazGU/d8y/gjSl/0wo00pgFwA5wFJg+K/73onZ+qOhwSllG9IRjwSY
I4TE1p/qdkcXyJOUmxkcBSORSS0R1V0r7sDIuBEv1NeMb5TFFbA+IQGGGKqO
zky09/GSKYxEFgSIIjEraLOYvqss9GB2V1DpUsLnD+Ya1rihDuPxr6zCVTaS
tycjqUkTgE9ebr7NMKVj6R2CE70QTT1054mPDTm+nYGcWNJzkJG+kldu6WPb
yEKSaKL4zcEBlyNw2ZT2MDPg/+UF2dtq+OF+1r8VwN5g/WysfSx3AT7fgBWY
Ikvftt00sH4RsWnLN3D3bMC4fdMe6k0G+71Ti6hR8A8GgkDTr/0ILQ2pHRxV
ifK52ibGRiT3jOJ+G4848gi9B8Dv22y2bIwdP2eWgqGB0ds3rBw8K2DpHtdV
73CJZVoh6L/7P8QqyfmH/mwvSXz/zTUrxafWaS1BYz5TZPqP7/Nh+7oA09HE
B+3tsa74f6KmT35/BF+vst+pPxK4BWIG3rgy4FubHGg/SThVWd7DReBV8uZ8
/2SmYInvZCibfNgq92HWLzDPl3E6IYNsA5FrAtoWkS1pnh/0RXN9hbtBjF0U
q9HzCdb7Pr/AXut0Gj3Wq5xzZcJYnaWHmEpMHQV5vVZ18e154BoaWDSCnTW5
YiSxEAg+X0hd9JB/dICd0o0HsxFrjAd+t3Bk4YQPd4t7LU96dWYFxaAqvxXI
t17sKE2MdI8dUsp+2AtgLbpg+205CWBAW1b4zfGEcM4dTlQ5V1Zl3mpjwoWC
iQLoqsUmZy+Ya0EaDb2DnhaeTtg0OIqCyvctwjgEyrJ850I/KzigeT6kq95V
1kdzELaUO+8pMbYC43pX3XAw36oNTWukAdTIUBe80bO2oonwubFvxPUEIFKQ
rVVFcDV/e6WYHepM/0mWtIim4Q7qYcSTD0LRvIS3SSNqhTqK/1tSszyEKIZ7
uDzQ8t3TTAmJ9ISsZ+GOD42kery8LW71sCsMQAQYlIkn3ir2x3HyH5Cl3rYE
d6rdv45zsry4ZlEvvaxkHEvCRPSemGppwukW0PgwBtqNceS3VWoHFWqEz3yF
FcU2h4PgMEP94uUmABqr1gKSGsAToSWxCAzj45qyQPS6LfxBLSRTTHD/562d
VEOnJ7Ao4v0NkvZtiFKmivBZwEDhacLxfqP+6OADPeQF6EKcpa/+0Qv8sqK+
UpVjXDnIWiyEgh5qRTwfbY1liK8CBrpB7lhitV9ZiNOUGVDVxywYhjUHZraA
5NyFd+Tz3WjJDvbBzpczyt2PzzpdML6op/OxVY+zGJKDvHqgXBQsM5jl8b/j
CUL3GtAJQ4e5Lz13T/YFLmkzY/J22DmqSGG9pEcuC3bUyF1xztOuC1xkdvxz
cc82fxa6huXaa3lkvNurBUgXfFvaYoU/9RVCEmHBgGsbe7m3kFW5lk38DFLk
dzCCWDyRqpklESMD7QvUSIHPlT61hzfdr1gzUe6mpQEJVqgBbEWpmB2HyMmb
ocyNZzPDsK1j7axpAeKRrPK7xVn3qbcwaBB/ayScnLneoRQupRUOE+X6mQ7P
UzzZtiLAID7QDGaLb7G+KO5eHrHHkgmCCzEN6sY6HOajfrkvyO6oMJUOfLem
kHN1j7bJjQ40gm+AqkUCnSmVvz+qlMyclDqApgVGEmAuN0zemwohbLsQ7lfH
GYeYlL7mpvMtbjYy5h92Hwd3NhjxD3evfdJ3Yq+Oi3zgCNqGD2vxDVWYBv1r
B1UqycxBW0eQ+esu4o/P4bOg/uwB63EhgrkmihpPJAdeuyFU9sAIjn4jXypZ
ReC82FBB7tqsjW6PJsak9HT/hWszuPyAmCB1irjQCdXvczLmYJc5zO2dUmlb
foXnkW+/lQKt0qqs6paOC6Mg4992xtvse8cNW1PFXRHN8hll7Unsuv8oJ6Nx
BkxCDBpnJNdjJoSfj0bVUcE0+Swmyic/Lm2oRZHEpabq82bdCS3KQneZUMm9
QzhMJyGb9KpXuqpWk7J1P9RRGw9tKSa8+7rvFipo8eLdRfc6zoCDN58RARiN
hcZFcO6mSDBhV7dcDNCt1mI7qgzG1+QV6yX03aBEzbhgoTbGzhR/9ownuMpc
CO2Ax8Dpo9Qthmcf3lXxTIhI00HO/TIQ70erPmEjfN3nExsJbAXhDNoH0wfi
V2XL6Qu4Voq4juxx4veGCT3tcvdhEsUqRxudmU/cdSkYdl4bD7VIHgy55AeN
a+IyTe4gAMjalyCC5W2EZM3ZJRttbdH+6NcPXD4I6rSuP0MilATguq6dXrPZ
t+eRbaCVLnhUbmNW0IpwQTgz9VWIVh/lyyT9Dwu4log9k3Ip9QXXHMlr94Ne
dZs8b7ySuaPf6M1dQ9Up3X9V+/t7xp5jFdovcteQ86D7uWl0XH0w0t2KuKt0
Lt36uDJ4ML2LFTY5IIkDo7ATywBGWEBlBU1xf5PPjO1dcpZ/BbuYFgQ4TaII
OrmY+TPjYJzopj8DWsV4d03LTTgOpC0jDN1KImIRQDDUjCTkKvfQnO5IsVsl
R6a8nrDXS/ZnH5s1j8Xlqqn0Mt/EK7KvtYvMFSXwrg3ay/BUZpU+gXil5dO4
Srh6yMNNycHgMpwUTGTyinbkreXkI2dPTMHKDWsdvUWRPA0LpLZHG3DMFBgA
YUVI2mUNgesg0kqYv1Oi4lmq9hsLlJP1LvJXZllxEz6RPQVVRA0q6Tak6f7c
nlYvVIkCXqkXnTydqrnn1JHvjBp7+S+62wYYcxubMQRDR+IPMJ948d/l/Hiw
dFOwQqngCP8xplhQ/1Ew9UL5qJKM6wyaU82JkCkm/5ehH/ej13lvtKTnB6SF
fKY7QawgOwhqLJfGKeebm4un20y71E8Vg1fzuNI7C5kB40AvbjfXUDx3opVU
J9H6ySa/XZ5OQaAfqTRADPbloaz2DRtRvAHISpZvPI0frsv6v8S+DG3h1InD
+Th8YYnMIlLTE1CXAdAYpAGkaBeZ3J2OIYmSOiaXzoFmk1g0P2TJspN5chZq
JMHbQJ+WBCyfHMrLPqAATYjN06y9dC8aoY39AG8/SRAOK4/MjpH79eOc47gM
YMd4L+IlnN1czChQuT+csNTHaBByJgCKmhjkZgY5gH16FbcYLJ9LVQBtytDp
XVil/L67STGhGvofI8+SqPnlC0pYt7TXKtvOVlZuD9VD+AVVTgMpFgMtPiyp
HHt42ImFaJu/ww31V5MHC8G5jZRSNZts37YNR9euBE2bChvOhfPeh8m8b4sl
yv3TQWdT9nOd5+jaJYC3TMYhk1Zetuo3ESV2oRDIJx2uplT0XUgkkpA2uVNz
8jXAV/T3M3LqGWb5WZF4mEx/UE49XrxL5oxWyG/Ic9D49gaP3mRYVib9Mq+5
GJU4ROMhD2THTYwQbWaH29uuwXI+CkMquJnhdlr8XOm6uLzXK0iWQ7WVvugP
2eXw8wjdKto9nCA7P/af89MfnLKGDlwbUeT4JhK5c1qjOo+YV5pmmnej4sMZ
rC+rlgTRTrRSSVhLOF1wkghp+mhmtISU2xYhw6R9bgevnyTAcywlvGylLuf1
ZUFCGzukA2M1ctDnEnv/jfOa2u0Hrugd0MmW15Pcglk9TwXxvJ0AtJJyQk4R
SIL93mGr2zKN9g9NoRiJy6Rv+3vjqhLGx7bjunnfJmPwIWHtwqGYV8vbAVjL
B1NuKBo3Y4+n/PHllmOZKjhvNZUd+vbA5VRatHZf56uqRrA7WEJ/sGMfxjD9
qugHgh9Khnog0+ryJKgK9iXkToK5lTEOKx/bDTsO8CCR5ZV2BCGC4DVtLO7n
sHwQ54AvKn9iQUH14MiAMdgWfninHkC1CM4yluOoGdMyuxfs6GKmfZMw45rL
fWHAlJ6ltGuz8j0GK99ksmiPvzthE/1QU3cJ4T28MrlEC8U4jK05iZT217BS
cxIgJYB5fnyK18KOzSfhCGWT0+HoKgUrKQOndwT3jh3jLuulKwELgoDdOl2h
vg16B6VvHcKlLcCvwu3jUmmSRNvf2SV/6u9pqkg6o2Inf7fUZvwUK5Mx7746
Tydb/3k/CyNlgFr43hL/UOvQTWO3XGD7ZewCuwKFl/0Om9zrPkkucrdrVU/O
7iFOQbE8HoLvN4KIZhc9AYSag9LGRvjF/e2Tf0LsBRc/QZ6s1d6JyphJmOw0
JJ+LXW2WZux2nO8Fz/Q/VsqUSrcP0kRHV2wTXocKwoWJWFbKA27LHjx34nWJ
9WkSpGiCDggaY4IhyuBmI/lvJm3uqtw7BSSIb8x6ojLxuDNWw8AcNriA37JK
1af1Vci7XPLjsN9ttmxC+ajqL4sKasFypduOsVLR6PcCg0zmlMxRNqlYW1/A
hnRljrgAdkg9zeijRMzh8U34926zPYRVhoLRTwkYY8GBuiLyqbXYbUn5x3lr
qLWGlTxE48Ay/lvYPY7kX2uaX3fIdf3H/3lqYXIblHWMf1r6yTh2m4miFxu/
I5bKevaWbdpOjU/j+f1CnY3Wn00mZDQg9Z9AAXOx/lXSKpodbEXSiJO4tRP0
tJTQdWMFmUd6gez0WAA2J9quigN7C6oOKAEAZ1aC/sCxggbdatjC2bEGSJ06
y5zIt3mbiOYjeXvujJ6aEn0gVJdaJ0LdyRCiPMkA7n2rhS/z1wTa+M+kk/fP
rICe9Nlho4SOt73HfoV5Yx+woiXMB/PRQPRpBlU0QmF+3e6EOqr1qP0YtJsu
dArPl8jGuwwah/l7VMH73CYJSZVveFRfXCthXMTu5EMFZwn+X7wRhjZuHQ30
Y3kjIazp0RzGXdfP6sdiPF7kNwO/ehc7vu04KLZreDELfE5EEuLvVAZy/Hxq
JFXKMW0xAan8ZmHodTMrs/z+G9Giy6PEwRqu+sJw5+qqpOK8JhSTJcZ8/JMA
Id0BJmDB/YjqxU9tL/P2hysaCroGyv3I6ysFmLDeL6O++6DyUaigGRg6mReq
rwBNOOTv0/0pAFdyCaEzsV1fq+eQ1jTNolUrbjRtDrvnlV/Vjkp32NT5jiUL
gV2bFoawWMsplg3SZOC0jUlGK97bt4NeYuNKJ9XB49upYu07qBPlapc8c7sE
bHbuUVDpAiIhM/g8P2WPbOpFUZIeKhQ3UtyoG5F0865MXE7pvXIcxj8Osbx7
B0NYQER1Bn384Qc3G7Gii3Ks833P7OYt1fPBNyaLTCYmaopVnUFK2YcXvGQT
eU2zhOnnBvwETmVETK8q4VwTR6KE5GgHwA4JGpnVr4duzbbbD1xljUp/ji3H
ifQHsJxcXBwpAYSt8YA9CLqYfhtEXS40ngsU6kTH7l8NYPEYo9NhVJEVhbGG
vRzo8nVRSwDW8D/zA6q3ddAAzy/yxvriGIxHlKixDMAV1E0xwoK8ID20mTeY
QUgoLYNT1E2Nwf/wSyLbEJrdWO2F57ziZmXARVIg8AlKQR/e14O5ncaIaBmS
JXhtnJ2kH/CZab0Eb+XsMvBJzwDDQOknDE97zHmAwmW9huk5ZGxiWN/Ied88
uwGaiIy8HW/t7Fery0qbeCIKepEXPeWoXLB9Zb0XZx40FtetlPqlKQlcqZwW
rF5ipqUv1OglOF7O+PADlgFWphU1z874gAyx7vGhInfIbgimjy2+HFzJOmz9
DICa3wTWg/RS1fw03UMb8lQjFE1Dgb+jSVJqe1YUeSfrmsw9xIjce4oyZbvu
hrN3UJOibQDoPCi6V+8++rHWPGKIkDY/JeHS13FLb3WpGTqzAaT6ijCkPHTG
AA4LtHFGnIcA7fzwjh4Q+jl85tmMUbxLHCc0VPZpgEpZ75pzjOfCS9go0ZnQ
tb5cfAbHt9PHo9nIsMS+HI2bS8BYQxQX1W1CgUQ4O19n9DoSY3Y6IhypR2e5
4bML/QA2a8bdqiG6cSZCMltLmL5WOj0UWI45B9Znu0YxVrDMvnqQYpxW0sD8
SLoGBiKbuADcc5VHf8Nm/wAM3rJTJQck41EFVL8uIRhcFGptNayCDw4jqYnz
FD6n/y3+sUBgO9HVHVo9kLJwFd/2vWWNCpcxb3F7O4J6IqzUktn/HvQbDCl6
LYdUulx0kht9aXneFV92MC8gHMRB5p5bzyE+J0ll0+et3N8buGD9mlm00TYf
Hgc9+Ub+En/Vh/r7z1sT6/P8gwv2uDEZ1aGII5Rg2VWhnVNWU/KVI2rGuU9j
2lYht1qU71MUiOBhVbMgyY52u2o3IYGuovdi6I9bKkRsIAdq31S3ioFvLCj/
cGxUS+2+1aa2CW3j4FI4R+Ny3tv2E/Dcd5ThPN+Svp77bfTQ4hSwL7ndmZr0
95HQPbF82OyhZ4KmUZapNuF6ZTZkKD63EYbn9T2EZxTBH2q/DVGBsJdR/Ywt
OodJwz/hi2u2uK4jCUfM5fX+eXjDix6AIqakpzPSft+F2B1aTiUcYnCQQYX5
j7h9M1SRnxba4VqEKSw8Piy+M6iRO77rqJk6G8cZGrCymbbKG46M/NniNF1q
WJlzEc02r3RLjwk49LTmykgTEWi91BXbCDVDmhRe9VLi1PSVDwqRFmvQ2rTB
DgkwMitJi4F4whUXuC65eJmJAuWtqPsL/deg9ASiN16J7iE8gqONr3f0DQne
CY5XPHYcf32S7e5EVPRowRRMgPftHStlm5jApxvs5q9qQv3cRzMh3iUePaY/
Q3y5arag5o2ZgQ0ZpFB8zttPUZYbkk8x4NmPaOcjMH8TsLMIn9zATCP+hlRH
j2rKoWgZpztx1T/7D4rQnJu3aZ1PfTfvqQ9uI/FDfLFFzwopfRynj/4s/k+t
Hye3/okgW3gFUb2RT/MpYK80JqORSLASzFh8zh/y+MYq0yyNrwDrdsw/mNGv
T+9iHvaaz4eXqHGdZScXATS1YcyYPDhCfBHTMGmFKKJNShES7YgNawceQEhB
wxjQCmZnGKDlfYS2yUEV+0nHAMW8ukC3CRgpNehWvMXz580LTDafw3gWYkVh
zQMM8XWkWWWutP2sz7efy5wvHirmCevj4hB+qLtqfCdmmbtjYFUuOCjHnYmT
WeMeCCMDaUXtbviab/uUSvED+ap/ZnIMc/u77Jaw+p9IPNIZLvg/MH5ZEhpr
5tnDSmpE9r+HlxFQ9MqQPmdGxy2JwNS87sWeMjGru6mS/4YuyNuJ+TUjJqRW
FPBHK+TOOo0LMklTugMOVh9mC5MagX96nPBtdnoOcgDKE8YOmyKF8PvOchyM
yqrpB5YyCT28DDLo35DHFxrGBRYGmDN9HZGjlyfqQWw/qw/nlX4G9Kocl2ft
HfvjtuU0LhlOzwt0l6I/tgECdSBhMM5/9yNzr09KstOd564mlKv9Mb3OGqEG
Ju7QQtbEZ2wZad8j8AJ7z904RcxmOUkHB7R4ldr2Pqp+v/YkwHZJu6udjGj6
dnTHt+ipY/RR8AUUZ8I3vyVqJaDfzEvli9GqdDNFzbrLEsmlLPLUHZGUwur/
jYWEVhV8jHYVwDPCiVVAYTBjB8ea4ZGk2kgAMzOXTyAdXO/Ws1bfVbgwa0h0
z+g7ULJzjDvNFFO1S3+WW/yDcClBKiwlSHd05UCsofUTGMM3sCrL8VqV2F89
knsq8mCQU+1Cypxxg6QATKHF0zhca+xq+/BattVb84J1XS5R6KGWokanLbqB
hDZFo15HBdMk1o3TsAt9ab4xE/3U6crPYeQw3LWybFTkrJo1i5GzNL54HzNn
yXm6pZBdzoX6tr3A51VeLxE0usCYLr9v0EA51dMRb549vfNBps5qZ9ztpNDr
WNYeqq93sKXFoh+4rUxDRVTLVxSIfEZhrDaWgxO36RHTk4PP5W3CzxUYIe8y
C7nw0Z3yt52h1V6+htI846LnvxpI7QEV1F6XZdo+yvppbrOyph2axaZKXQ2z
GRBi+HrrFqXJfPe8OO7dy9LBZ9DpQ7C3n2mS1DsppE8O+IUNhCq8HoUklBb3
lK8Va9x4eN0VgmUTkBlxcQqRwD4TdJ+R7qMf7bahI9QyntRQZZnEcArgQ5QO
sFbmmOpuwZz6ChURzfbxZLsB+nCzT7RBD4agOzuHCBjGK0fAhDp6/N3vwfaj
3rQx4o9/8uZDjFXl/g6hMVGuyduXRPKL03fL6JFSCjnSDiCt28/mOI+KOtvi
vvUVn/4UYSNAYAqXGFAck00VvtEDNiVuFVq+THN6a8zYN9YfMU9o1b0wwhf2
omzl5/Js+zqEN2mExRdveTU7MP/nVwAH8+kjn2RWWuBpdRO0oPpyVtBFnNkq
Q7WNCG51lW38RNFp7fnzqXi9YD83i5RQ0O9/a/vx7h29lSzG8W62K/8GE+uE
FwUakA44go1LRv3bzpPWnzC7201Lx8PiyJRVXPR1pgyLa3amlhN5UEoCG8+Q
Huig7CC6wfjYr8aQmF/wIYkIZ1lVyaE4vz5NhjDY27anjX1cc8vrzZe+z3v8
96b0b3yfAqU3mNjk2hwzS+TdqSEAsJV3c8WyBZHG/4Dob5mo+XetXfL50dBt
G01077SiEYYEHCFX0PLlbBayJmHiJA/P2t1SHJ2LNaSkchUHJ/30dTsmEdH0
m4qdqGyxyCJcexplXZEApd8fYmFFY5yV/2HjvtLZtgUsxiFQvTEOwo8Pta2p
HwcUUA0iytp8j12vNEgsvfOLozaxnOf9hziowoJXQ1XhnHp1EUKm24YGk+k6
iv/Ny01eTCiwIYqaXbMl5xLybSjbosTGEBkf1cFJBE5OFPiRWV3o2Mews44Y
BWAhdtY5tNOiY3ZdkiTvri/irCdKJLumv+19WBh+b9baPbLNtETqgK6dVgkK
m7BF1oFzIMr4J0frog+Cexg3llCeE9pLY/orQuAcHD6JbbwonAwCMgRnfbSq
cKUTGUJi1jbTavCvvFMUMn2rbh1qjKJI2Vb5mYCqFxEdmBqUz2O8LnPqWyLU
6D6CpWr1wi8ea3uE0N9bTpdcDOgLEVrlpH9j3w76Bg+ESPol/ebRRmqP6Tmv
Sk8Hx67R7S/ceOyaBadFP2gp4yyxKQTEkMkHubDxJ/5LggCX3RFRianPrGSZ
DFrPBE5MkpYy+k8l0oXBECzCibpKdqPtBrUwk09eqm0GNHPEYgP2FPL24Osz
J46MZ03otxdxOAKMRebVGQ23lg8loMyNshCg1EKIDB1ViF8cBXvVjNqwYrfB
IVSzs4m4TANlWADkf9WxRYntgu9ZdDvyPNPdvWVt3ecsekp2HCW1pZSHk9Wk
uF1eIIBXvD93yggIjN/jEFinpiHW2uOQRH1l/0x13qGmxCNP6bVidSj8QNXi
6KQERxr2ScoUxJOYGkRjS7dPHJd5R3q4OYZGH2F7z1JjtENnRLc2epIV0eUJ
i6hy7kwCEdpcw0/YtG5kmlIPg/mbmvJilORRH7HMGi6BMP5Ch0/aFPKV1Q1N
+tAQxAdevMC9iTapbWwvH2KpBLhJswnVEpttb+EL9C0ed7YwSJquVneqHGjK
t83Tygy0G5Ify9GCMSYto3ud0rShS8MEy56iPSr+SiDC/oJKULq5RWPVWjsL
EZ+hIsaATPy30e9ygK1HpXz5YaRYS0AXJKDcOS5YFAuFPCEWFcS6rx3S/9ya
Q1OvnyQwCJQlpy+QolJE6vqqoCT4anCfLCIeEumMJF/oTc6mw8tI10AAikeY
kr6S2IAFpZmA6occDglgnWRq221AvFw6ebrcidaelXRE836mKSobe79mac25
jev7vdKzDzRwPnWXGsJZ/Q/AqqQfbE2puV3/fXri3+/RgpLJTWRjIP9IuElJ
eHtZ2zA/QVtTOJKszw+vfM8H53nBT+6Lj09HERgMbdpbv1YpTmrcfPUB/fQ5
TTqXY4j/0H5IcQpcyCIj0UNyZxRjEnWJyFEwpSXUaxKwzMeECWSG2FzJeos2
hwWsFm275F/4s2mx2Qi5W6DZjyB2x0VwBdz3m3EAYg7IC4Ltk2LN6YRxMu79
/f/8FHbgUEWPMvldhXD/E0rrlz2vzinqoi4kwC8thEqRo4UAjjxBBsyilKmi
kbr9JZFScIwQwZKbs9qyyZT2czxED7e4UD/pp45S/7Yap0y6B5ym6Td0ymA5
8yPAqbXkgVbPkcSlFraU92/ARHtDmSBJ7q8FCF3JhM+Z+zINHficcGEHEDEK
Pd0BU52CCGp3MFRZQ0WnrKiujF6OvGzsW0/5L7KnBGngyFzFlg0w7CWItHMY
zoAb0uoQHNRlIPjudOKyAEXhv/gomOOB/YGPK6bc55ZeqE7JcKywDOlNWDPR
9VVvJ0axpoAQ8K97yv9W5BL7IiILyeSBqN1ppxHLRfJaie0E5E+OFAlGa+ua
VUKk6lbNjfCEad9FIqdU9zLJD1nqy6jA2ue3cl8yTGPcDDTTUydYQlCZ2q1g
KikSLKHDyB9iXObOgTFmdEiURd9i3wdKaNTM5YSUx9ak/9tMET3i89YccSb4
DTA9TE3CJ+1sgDIiLx3T0Bvw+UnQl+h/8GbfSdbmfe38NsJVwvDt8ZU9jVv9
QezK/taxQG9Ax/0tpxGpVIinefj3nvHaLZ7+19SitKoMDBIKUkqMAW7eZ9QN
Cj/ta6mH8cYSKRBBr6G2jcd2oox8EbrNusG9ZPKyDIlhMHt260eNR+PGlpzf
IB3/NNVfStnqG4bKUoTBFb7HZ9YtJI+PFDg9h6o5xNWQgYb37bbT0FUvxGVH
eZ9JLV7xM6ONq5Mn9fCZsW0032JUGpFxZqgYcrsY2YtvcPrt6ecRMsRw7h3R
6nAGSRf+vIf2fFzF89JBj9fzm0axbl1F/w3DcZdQqJ8UbWx9LI/KSOA9RAVK
iGHVV46MP3n/InzTRpB8ipv1v+e7KUB5H0CHsBmi9Nggh0fb0LrreKdQBMxl
irVkAtjMgnyZn/1c1aMqDHQN1wsm4ZtmbIR4bNujABeIkEfkfsQhs6dwVs1U
f5ha9YzVBoxkThokCFiSG+p6ICZ7SIlaRD4jN3t/99yEcqslGn7M/L64sc4H
c7p8gwePgaTTejIdc/wDXqaR1PKyEgGG7bDpZbw6O8IgynDVDNe8VQV1zIE9
6lCYeZjF5VdK9+XLscgBTX/9LpvR47zPeIrKIn36IQlR31W88JqJa97+lWUT
nkBusumf/BOn316fFc6daW9VfQ+GaG3dfuLBIRPTTdnCFGpE4RbR7PtKUeyF
2ml0oD47DHPuOypx0Gsh8MuJCo46M5IVycj48thHbpBh37m7oPq933D25+sX
UiTVrUpbn0/8mVIdhhKLOoHRK4F2mUcB/nP4uXccH88Fe4k28wW3EnFolPKw
PZbPpFwh4pswss+qwkSiM70kFIOkLLSUmsB37ejfnLjlP5cNMLDI81T8Y9YS
LT+jSrNjqdD6+7S/mvjXiFpLY5zEBg71haWnRgzCDuW6EgOHPsl+YpHvUWQ0
Jkt8JR6FCdV/WsPOXnKoaSyxJDHAy008iehXA2lXDLg8t7GJetFpP6e0jEwY
owjDCU/9pBvoI30XcuNCkB9tVW4Lnq3Zsgl66uYib63WUmDGFoPW3+Gav43U
D9SInQ1RM0RdsOttevtPiNKUqUN6oarz1o5kxQaSjA1cqKkn53CZWtm6994I
8w8wjxmaGAbg4z/AFP4yB3Aa1a9VuiuROuFZFcLO00XCgXmowuJNUkTwsfHN
7PXe9uLVlXzQoAlVQSzLkumyKiwzlVDhL/syKC9pqgKO08aVeAwltCYw7oMh
qZQ2w0RJ8TGDF0wkkxNfyJs4SHxcP/mmiNdeM4jwG1ZaZgxhQE2zGSe4Z1Qu
CZ9HOUdq0eywmxeRJN4dMjp604IesepMAQqddrimzk1pgzZCVjwz3WetyncR
yYe3vuhzNv+V3Rz2LbxSAM8OYvEeQEqAJ3ppqwzpEY1xJYkuJKYk2qhFLZUb
Y6bWJv2CzUPO3Vd4D65xDovOJ1rMlOCq5rySUv+jbvw8GnY23IiqAuTnYShY
AYl9u16/VToQmd9Zp4wQ3ghli9/XCI3ClWum+AtnFedFX8NXX5ag9b6Se2US
Cf1Ig+E43WsU/AV5FjGTBbzgLjD51II69+NqUhVswvA49u1P5jW3BbdwUJul
72AiD9/tLkRUgG1cM3JSp9CaHKEceILTV5W9e2fnzk9WVxGXXoxc4nDVY14P
Wi0bU+HTHXMrE3xMQocNG3GSmJ5a7RNlU49x5wYOZtXpDh7pFMQFqQwoJC3s
GfZ5ZgphxKysx229+r7qhnUeV8U1kdtKuiIkQfl51fqytxhozxrhd1LJCcc7
yC2iAyFJdT8g2Ux+T0+wNfh/6ACgA2qzHk8/zuRLsVzlWmdqO5evydXxaCuj
3CvXuBGXhonHhjIMPplOS86ObSTl9Pt8zarmWEr/UK7VWm+/ZRwQG1n3mV8d
bvPFsmNhzPjZ9VdH9C0Y4hy/Pm+8Jy66Wc2ixshYBScJrphqIUtWTo2Cwwzf
m60DbonNBpvsMapEjAEaehKKz8qoSeQsHbTFD66R11Ws0dBjZgmsvgB0fJe0
E+jrpkVrnHppd8VOeq4Z4Y3wdsa/E39SNuib4O5xCA6/6IHQO4phzlkcQQj7
yu+mAV7mHVGuuiv+MN94OuzACanBgWllz8pqmXinB9588WDlziz1fhIkcyOY
I9VLdDZ01AVDLGq7sCT0OQkmV9PIskDuwOb/rusb1RAePv3IbeBkELvy85Kx
EM0Dl3mkiUAvOCMi3mdVT1ruWc6/bswaJA0cOgnsdH2mdzZFKD/pJwPOb0nT
Ej9O/lSBFQzaqdzQnhIyGrsGoEq0qbBgiudirVL3tht9+eDTEY/OFgSPPZvu
MOzIau1EvQDOYLBhG8BtpAZhtXbcv3WEeGpHaBFNsEtcL8XbERSWZL4rGdTX
SUY3tBdEpv6WHNcor2nrzXqyeENQfGjSUb/soBX1T6dnEfCeHIwkgXV9y4cf
7dBqmAbX6enAw8RqzrTF3vtZBj/wKinSMrDKEI2drxxSBCndNTbTcMZg4OTz
NMrfGlj3GxST3mi/s+myzypv04lhSs/B0WgyUbnTxfkZN6xfrd5L5qPCvz6m
IVpcCALRTaDwSxBcCbTkjY4Q3jDh4PPwqipspiPKy971aGDB2NOrebjB54H7
C1oTgZI0WSP8iwqfl1stzzL/fCD4LlR9ahre+1weiMCKgep/9+SoAi/dgWm4
/Rw7PQ8/VMn4hFVVK2NDBqUHeERKk7aLrH1fLlySvmPh+2jNwqAQ84BcKVvL
fNOq/xn4LldAGbGpDz5kyZvKeyO1xAKeemAaNSIH9RYMLYfhlKJ+Li66A0Cs
b29DDWCiDl153SMZ8pIh+xtOjUH+57UTGNWq4pIm+wfkodR+Iy+ME4cPEGUa
4yRdwTOETraM3F4c4FLWCyJD5gqzVaZk7gQBTQIA+nITED1EPxGX5Tj5VH2U
SHTtwu7TCbGAi3ypgmlfmsvPTscYofuXOYcUisQB/+ejJYxVcFWsle4yXFk4
aHlwBX6dxwjnQ8Y8Xeq7f2Dfqtj7nDJohcQenVgAeW7KQ9jaVdyAmLJdRIAc
dcK+15TPPcOFu9w8lFjMsHzUebBl6liIoMJ/AqVwfb0zMVY+699ktt7A0GtS
k8htz2WBDZp7PNKXHdySKMzM0euAnT5OxmkCt0yr1tf6qcWqh7c153RVg4My
3i9haLF7YNILtxeeNtzsYsGASq4OcD7HF0+Tf7aS7xGWJhDH3cpQRAwzpaPT
rmJGAmGYm/H9w7MdVavg0AyIDkSqeDppc/48Cly3PK1kWV5YtNKKxXnEezJ0
sub685jrxYD6Y6XraFW2wB71Req1+UnYVlkl4xA3+M/HVLYH6hPML4fPTPVa
69S4d5DF7xpIx5mlhsbOkF9uecixtoCBlGGGsAVJnxA5LH+srthRuvSg4c21
lBPLLCUPCwOH3wPkrD61XCu7ZYbVaRohztW2iUZo290WuAShLejCdGMsk6/8
hVCnMROd9oxgTgVSm9lyfa7FQHerevjp6GtD3IMvM9lIjAzZovmD2t4EF8P0
Byf/ExCC51vtfd0l2tVHy3g2vbmeSqMCs4Wes1a/xy+VpbfiPpxNtxo3kpgQ
DjKekfZaQhMRIxxDb3uCwMeXFMAmmOdsE7B2o89rsNbKOZzi3w24KGiD8jWd
OGemdkkns8Jbqu5M7PVgCgWahBW5xBGVL5FAzWQnaETIngJl6U115w0Ab1cq
/hsjbvk3b3TsVILe/4OGq/rrW1hEYhg1OhJUjqmrrphrO+VJiMfrm/4nOid/
Nj0Sj6e4rH14luQmNmHF13+962AV+c/upyWTAsSaPfQ8hA+jonqy1X2KxsPv
DDOPn5bTqYdJZvBLm7o3q3iV27+9r38Fz5Uo1a8VWcwT52r4eXxwFPStMlVB
DCIMv05P3LCSWkBYwG7UWRjiEZMzglj+6UwUtFZOGZjZpZadI/1ghJvbxVJa
/MfvjnV3r5iuxjwfKeTyk4BBYCoROW6fUF7vg9ciRZb0ood6o4Qy1jD5YHF7
CJunye6GPqMBwTx2LAW/0D32XRCkQQ6n3UK7qtyVhxVxk87wJHpPbgYW3Ux9
z9ULfuVZ5UB/D7u2xHQnBxtnn73EgBX2SgfiL6BHKfzdNQV84QkVqqPA3A30
oDN9CUCuV1P6unSSFX4HTtbRzHo6oXO8HTq39SW1e7qc5Yauc/suTrS8obXo
JdIpslZHSygBbfM3v/8bETpEH6X519YzvtgRniZS6VSg7HlAirt8wvhs0fDU
jJomcrnTMNT1oTT+dBjSA/tnFGmA7ow/D/vMYJazm8NBWlDBUDwxBQttiZsi
uRzTIJaXJihrLlJBJicmL83Bn+ttcPtTkhx3h50fpN3gmiBRlK68rLP5ME1o
kV1RbwrtDtDEaP5kpqNLEfvG1BkUqHbsm5MIVjcL9iuhEqxsYegjx9fWl2XC
DLNx9hiDTcdDXRYVi4VaFK3Q1/jda5hkg/CXAg8rncw0KbpTq4dpm0bMTLKY
taO6NfPcxDPQjB/SESmNlJkNFS23BC9k9/1spuf9EHJ7qHcfzJ3UCx5Ug8Sy
WG7XWoHa0A1dbsiv36OniPa7WetEzJkauMjlfSUY+nZLqmroi9N6PjtpT1Xd
e4YWYqS+vazes+BPX9L7aOkj4wgxSQJrZFhKLL8NgcnabEEWsfA6fJ1UuOLZ
ptJmEoGxLJ5TdYoQvnfOaLxgFxrmQbb4bqatlz0VmBKeyXE7YkcNmKaQwxKD
MFisf4pwpHlWnTJrlhjP3/eDWzwd5bhOPN0d1vn910I8Laja56QlvEwqEnoG
ATCu6ylRQKozki9lCnf/LJyya5mhWi7xXSXJyQFuO2BuiSwqt0FYnJPuMGFr
mWZ+BiIRYx2zM3JuWWC+R52UjyQcDiJd08WVMBGD7QhuzzGfkLta5N/bMBqi
rG+ACn4DiAZj9/gIKM1gf6cIoLHUM2ZUvhynKsGtPDx/FK3OcH8unA+FCYsw
eVU2h4CEyA7O5HBH8AQPFEc3ov63MPfPkfC1aKwXiLcAJKBNFjNrde+cG9ij
VH/lkbLYBaUrcFjkLb7sJ2kWkBkjkupWzRq6oWa2nA/bEXhN/uTFVwovjina
IqHgVyCgk+48w92DNpk9QEWG8UJD/CLITo9vJHVmCXUN6vE0gxTh1MYe3k1w
50LB2IhWVuFDrBUrX8NSuFecZf9b1uDrcLfAV0vLJ/GAG/6eGWBfQGlTUFaU
6e9nBT7/51Nfh/BztnwYtzna6Qw1WfpSZESVYQMf/ZjarVrAcY0IE8G5YZRX
1319VjUpyqsLGVj5LM8NGQjjLU7NPKagTzX3a8EERosCl5OyzjgWYckV7qoC
Vv9DIN52vaC3fxCjz7//o9DqV4HCd1YxIs3L5HEdShZJmIYOdp5104b+L0ir
I6TYMWE2ZtpfzEXS4R/A+Bw0OSn/4S5i67h2HRt61BvEXhqQF6Nt7x0n4iez
zCX1Cc3LabSP1sazbUsnJ9nN4qr+VxJ9wCX4m1J41+eyG4mKW6G+PK/iJce+
Co0aGvsmDBmYsRFIUDYRglM/rv87qTOMl87u7XjpHWTGsfUBEpOXv26sgPUX
wMo3bDvRLxqT0r6RO7F0zhouZ28cDmS0bfaFsttd5M0GTQ0T41P3JzBjbZ/C
reAlU0si/6CrXLCrgbwcU2swWdqWlVNpJIzIEa5FKNHCvMknWHzMHOR9NCiM
eSfkvb2eDz42AgEWKa051paopwORLtFyaOO3XE5FmrS5RhzVSGj0hGRHLA5K
20io8vj3TPefgs5l46bE8IClZLy9LtIS/xYPj6974eh7Y1eVy8insrMoDUi8
MR3sp2H4+iBPtMupL3fMpZ9Cr0FJn67PqB4ArWMFkQ4B/tI30Fl4e8aRrvyq
5BNIrez+wenuZUXPnLFHpFZ4Pq/xXbJ/+frIRwbt4JVEbwuAlaVTD8uvK+Vc
oYOrjC2/MdEJKPgHwvTqdfHuVZtcJGllYaF8xcP3A7bcnTE6ecQ/y7I5A1eA
WZHhKgSpToy2RUGBIztN2kM8AnS7ba42whtcfATqa60t2ELNbysROpwhhPx6
f801ItMEwVrcXlgEGIru/avoY774vjdT6L6KUZnxHxEheInfGMHooBIwPucW
6gELcUunsQpjw0Rs9gkjD1KxSaAc0pGh292smwKEyDCNKmkLpmr9bSalsIcY
YhF/MmYTaNJnT9/LVXCRELBpriipMbuhLNWdzJhx9lLj4QfI0vD3FdzOnFgG
8IF73oy7MajziTDNljELKmITtXGk169WvsXn/33kxsx67eQNBH1Y9BCN+DkK
wm3bvQgI1eGTi/3x9XL+8wEZlIi7TiJO99XVEcWPuc9F9FH7iGi9TFRm/LY0
MVcqNpO8bXO2x2gX4deFI+kRg/vpVK8rFETxf1wgnF/OMQnW6h+y+uJ5vRdx
47kAP5+GFMpzoEkSTevPF5aZ3OlvFlJUCAxfjD4AOV9rp+gggeM1abmw1KHu
mBPNnZMtFOa3907Pmm7GCoswOIxVBie5cgWJMSAPka8xonO3KWqNIPIguGzC
yX2ISAmCQu8Iek4TmyAWdhPELI1cUVZC7bo01eylLJ97zf6+mZokwqKReMiO
FyhrGL7RcXl4OPZiCh0mH5OuTr/Tj9pzR1R8RbFQDXEal8h22XEivbuNKsOe
jP5x/d+FCdyXlzbTI+YTIUvIWi465P/XlgY+M/AGJTQJMvrMpNGr73DxICSP
X6/E6MI932ee5zW0Nv9LHVT8QeRob2nasSyFkHVZrqdzr8pAAkUyy0gVxXpy
5VfolCYJLzBleF91cIo8YEUsPZJrG7ZGOxkEwfAa/MDyWnljDkehnEHcMMZ5
0r3rswACdbczObjxJ9mAjTcKIjQ9Y14oEciRHTGz9YaOn0l0GTT66TQ3TpzQ
gOhDLPO8n/ImzrsOZKFU+9l2nnSDrJkxQJiGjHP4sR+etkMZTTYK4S02pEk5
917iFbHvHASGxIbCfA2UG5fvNvDG5qX8wKzqRP2/ddn6ZrNBtuC6E/qgpJyD
dk/M5gT3v925qyadcDnJFS+36AuuE0DVkCWxoMRkufmP9R1mDavIYcHl3OJs
Ue9JVWzH3Ird/Wk/B22rn3j36RckT5T1ICcPI9taM4Jy4zwWQNdQhSfxu7q8
gnzK3ICb9BL3d++D4rr6Lk7hRds2P6j/ARcmqAB7YQ5yk+OYogU6Ttnm2PYf
v4JFC717YHzC9a7cEhPe+o14QAfSNvSLEQDfeuG9O3n9mBi+A0YL0SG1kaYj
QripmGWEEqGNDqBqfIYR+uu0lBPVuby3OXAlayP6l9iNOw7HxLn/inSFVpAQ
d/aYQvDgo3+vc2Fy6uzf2Atr8cIkzbXvH5XR2vospMP/afKF7hiiSRtf9oyY
c9B99rdHp3ZSJbqgGzla9JBobsxePZ5KIBGJgMF4a10qr/NiX+aRKlu8CIno
ofHW6UlfEynlTVpE/LEzYH+p0Lvm8htQkyHRXDSUiWmF0QLmIllN/zLpqyZ0
+8FXx5QeS+zSXlpTHBsp7P63GOfqeq+eAD2p+oidCmEz+fcCdN5JKyvUOf6p
RMzlKp17WOR+eXkBfEVd19ehPLBBsapss/rJHy2TyYyj82IXrphKO+WqDo5/
d8p1T4ZIL/02Tfd6zK8ignnCKYocEZVlc7RKuSsnXQFmSR8vUI8v2Km8zZzn
G/46MsEajfOSCxoBiKAspL5kQREXAh+/lo9j8K3J27/vAxkKtXNU1NRnWODV
W9E5s68kHcBXw47NISbYGr92ICh0R9FR9GUyy3PwPl2pzj9Gxj1PS6ExXpZM
hsOyVwrQjB2qvcpS4/kcaQ/D4zDsldMJ8tjeg79KyT/ivO783r3ukjHa7e/B
0+junseUzUq7zJyEX1szMIV4FVYzWJW/87iWL1A8i9Pzyq2vsqtRAaxO2Jj7
Ua7CkNoOWAlbf0HDsA7TYBcbqYx3/L2eBO7fx0U2ELbsf8llAtdDEqtzAbHe
QPojX8dOcuHgjX+VDrvgEj0Hb1Mu/ePXscJibIfGIMyr3A01AcJNlhP4dF1r
rpktLZOzL/tWIL76NKBmT67NQDeubYWXo/5nxhvxdU6D1Gt+Ktxu0FyOalyu
hgEyxL8yxr6AoqhWK3c2gsPZ9ugazmKx6PJ+B+jC22MF3+0RM2GO/5xol94/
3zBVOBlwlE+7sZDvGtHSwbtOZBuxm3kQTTvB63krlygwRjLsBh61lcbXDdnS
/iCoQ/wBJofF5E7qBFXbTFJVvNgARGPsJO8I/6nPHgZgn9h7laz9Kv1Xqx8o
Td37TdzWUbOOh8DDG7ROEGxYcvereq49ElKFse3ZfuYnPaiwcTG9EGlPhMxG
K1PB6sb/dfTzRQBv5tGVYFelVSgMCaJVryl7Kl/cV8VjEJkioReI40lsW/Z6
fPJvkIj3GPt6x+gtxQ2jdob5qZeZvkv8iiZvlvUDx7rSETC3MPQDBkkOopTS
JaTKX3dNGUdqqCGqcrUK1gJj3s44j6suEJrI7H0nXvAS6ydbXKFHHJQSzBfB
nPmR8vGPbUAM7CtJ/8cGEv/yLN7g0OhLhzdAhriZaoJsA3iLe6s5ZEaldWKy
lVs9XFyXZmnb+TX+I3MOo7qOvMnYWYMML0STx9evZIKG8UmzsegFNUjS9l2B
+fj055vziI7TboKmbQ9CUtsW/I4iU2ZSLRqWlM5XZcTRaiT+RurtnDHtD371
7COzsb2keKzxnR/B3oP/wTK/OuYxtxD4x6oC3fo8e66/Qm5h3ZjBo3ABZ4jj
mzusXzPnBHUVaPMOvPCk+vW9ixeSLgJEVUfQevVEzTmCKZjt48Iva+iaQJmT
4d2KHcwRidhelKDxQFOsAgO25m7fQZOqS1SMMWPRNjAEV4NxyaqN+8qbAoZV
sFc/ScjhJUnXoI0a/BItBTjeiJJZdeggRPGAIC5jxI0ELluXQxa1H5u4DIJ7
hqJD7iDNMPFP8aNWDGmq02j/udoneshhR+RuMGBCj5Sr6++TKEnGrmjfqHnb
S2v33yY05p0qtpiOvM2Rj4YtS1GHUkB9qbxwawoGe6L2BgzsSlPPYP31Mdvk
C34RilNLoJXRZsVNtkCbfaBCwH/KXQ0LY7hVb7GbPqoPc5cHuNSGXk7IVq2r
QN/X7vLwY8ZPDkX8GFPL38WFC+8VfXBktAxTlmV8TscSSGQqipLpmoNfSegM
nBa5P3hAWpHDAxVJmhMaXvovtvGT8yhxIQjOqY+NPWw55qSTOmOkBnj3nwR8
i6q/PV5UdU510PgdISly4j0pp3uTejGmgnSeQXB4jh5V39imJxt1iuGf9Ao6
4C8ZuYOOSZztRqtTomYs9uJjdVX5DQIwbNHfuZaVANUUTWRsLP/AEMhr3c/5
lpnJxBOOo4/wOI80JkDnqQK1gsYVkMLzDU7i+TaZ55d99HhnTB6sB0xeDcrQ
Dnip+/kHgOduvZQrhydldk2v40lAcj2yBUd1qXFZUF07SjTC8UlZyTrNgXUz
fOuh464qqwKFpuMrzcXwYjEicJ6DJ4+xkp8ZR0MlJvaPIRuK46ii2hseZLHq
8Ri7v+YY4bDXKN93U85aaRq6smoGJY7P5/hw4pVDLHCOtXdKPzCI265ArBL/
QsMA/++D0WuZi5onA9By1rDKMHxc/6YKxurlOJCf/vmZ7Zv2+eTHrsNHP1jr
cj1Bx60f4Yv4sbmwYmfJkRqRbWT9j6qDH0DZhCfqBS4/g8DFcMwW2QELcKPY
NEov8r3H1P6vZJ2SE94n3uh6Pf0DjKgWcFfNJyRlkwUJ1ifAsdGe3IeHbwLq
w6uLO9gccDDyTqlNyEnY476z5FSU2Mjf9T+n3YjQPaGB01w4ql+Mip/HulHR
g+CBEAWR4c+btu+KI+u+GYFFmZ+gUZ9iosUJ0I9XragaWPkLil+sNQizH8/K
XI1cfqYxE7whGnpqdec8vsH64WfvOA/m7zPXefJI42KWYxz5jq46HtI9MWnh
t2kbUVwbuxpLsHyVhTl1dEN4N3Shb2YRYgnxM1ZygVqZ9Dh60OnBpUWMZxc/
My0FZpIbYvdNSh3Wc3W1WHvbtE2DoGRzCQG5JDG6aECen65uMMqpHp/qQyAD
GNocr9HsPPoxRTJ9G1ai+jpPIPTOpfffG9EekeEjp3rduOJNwqayXdZoyelI
5crsM6zQfF6OpQG+BVZhQ4yCFqXK2xDA3+XYeSGByz0IAlde3OWGam1Ss+mJ
qw+JClD1L8cq8le28/drynU28kNoD8UHecEYZKJ7ctp2BUDx001ToG/zlbdb
SjSGHby67ulsG5zIJkCGXEepExYWrz0oCs8L+HAMJBQy1MTnt05kLI7ta6QH
45el2dPAxWU4n5JsbnXEhCYWkTvDZF5oYwZMCvvSCBn/45SzMXbCsSUIcNXp
44wq7IJOYF+tvZm1vuKqXXgnYkLEmcDIVCs6ZOws8bB5UhUF31mFsjqlBAgs
HDLSp97r9YsVu4TgL4OE6Id5Rimgni2f/3x6/DONOXU7f3UToXpfnlF7KJqE
7kyBoiz+/51ZVUGm4bFQP0K8XFW9jH+NHT8arnt2mEp09hzuQjEIfMNlOzUc
umb7VvFnOQ56ogWIryO95dbwNqp2jQkKdODe1OnN/dMNebjobONIhDxWYLpv
EsGu6NMrwxWWAsJTt7SPDYjr7H2WmDpwZQbu/00xEFzQHkoT40mG8BHB/gdk
Sm1Eozjp2bnnDA05jK55m0OZuYeha8H4bwLXe7ziHvOY24Gy7tukd+0OzUa5
zs2MhfFJBPxyi7Nc/IRg9iR6aWdMvPmSz7nLnsZDHEuGePKTC3sGuuVGZ5hg
U0KJ8vP6zpyU+UIDGI2F1oUG7Vm+8QPTEcRjs7WfPyyVsGqNbpagsIOSYbp6
QfkYYpzmFxaPr+sGSQNigl3/ZkgkKbr/JHdCAbfK6BIxOS8UpZGCvrUzGFFk
a/CRlTuu6/oVk0Rj73FDR+n/NBpFhY2L1FmPYqnPZ365dDuMtXzDj1fpM4IN
qISf0RJPtpCtfA6esDfIO7gvziyfqpwyn9IuPAaUQgLGLZYMeiCMWk1PVkxb
8OxaDqx5TI6BYRYbdRjMh8506AS4CkiFeNYrXL8MhJnF2MyOS8/mY3v8Kt9E
DWW5PfdFcu9u4yIOrXwFsRUzNm0JxhrKMXakgRelvcb4MHNa/7xnnIvvmARq
hhJRHLdWLo3/SAnXOetScKSo1sD7hWihSAh3DtHTb8frsy4kx1a96cR4LuLr
YCPytfYSq76x8JWIKFK4bZOyhLbGx0QhOYlqwE5gQ8t+odlCJIScAZPLlck4
WbKG0iIYIvHitCmDV0sSIvkBPgcQ6SVUNcfol1QBxwE94r0VU9pC3gxxrGdC
14feKT14PMM23uvMF3LuFkSC+QzYhXSuPtNiEU1ir4q0jJAGc+maPcx1rw3c
wZvPSTC5tcbvpcG3PYuFFKlER0aV6PYMRx33fUaBbKPLz7oKPJ5nKVQsNR8D
myv4mjoJw+1J4R+6smfqFF+TMV/9w+gOxKDCjz3+OMeRsfwTKiKEiqRbq2+1
/OcdVFuM4ssOTcDtFjOJ3BBfoAShWrEDsCUflkD8qBPtWscoP8OVMqLPjxQ+
WQm9EQAYA81jS16xc31RxPfwbhK2r5DmONnI/89moHSklxyTPtzPXQhoibJT
c6ZP9p1dKPAXn5qW9PARYWR6t3euIneaSeLJiedREzTRVZbzW4daDbT9KZzQ
o/8FwL44dIEo1K15RsUBYZE5X2+0s0PtD70tOeLRVI+V+Mz/ITFQA2No4sju
WUQGTU31iQffNkB2HeE3jv6RBugHILCHDok+ltDYXUzQsy2+3xeSwV6H+z7L
YKv9PZfOAO/T8PrDcwAG1v/GslZYAzARqJqbyHyWekG+1rZN5P4pO80WiFKL
aIXcG8JY4w2dihhF3OobBZRTzUKZwNjeP+unXSXgVovXiUIogRm/kuKHBdrN
dXSSEmdry9ElA2OjMNmi6NiXSc9dYwERF5/XLWq8qpS/VaXTAGmpqpi9EYk1
AWeuKuqcfxxQBSYgqpd0g/soZD70g6wOr5HOjfU6Bpi7CHJ8kwKLOaCa59h1
UEC4RKJNQRXtO+ebE5WBnd3BoUQFm5QLNxLYG9WUI8nF/LfqLWhJvhBHeDER
Skmy+69YDE/VsduL5DmdfpTkYQkbfK9vcJvKRN0gl79OJAknEuvK+zaOQ0wf
MXP15NkVhUzcatE3lekfHFuwTeHpCBWUhOSrPHVW3nLSmUxjlLgjCWmEYA6p
DH2i82ya2qSsTg1uQnOSJzyFDeFpoco2ciTWU+hfnd/JPV4CL7GyRcXlEHQo
1ckFesDWk4qZyEf0vrUXLhyK09TINX6x2R1WqWeBt2Y7986TKQaY04JG07E3
pET/WJt94RNE1YzsJpZXq8UkS0dR3TTc41wHaf73hxnRJ4kq8BGI/Ex2rk6e
IeE3DK7JYVk2j+uUgLbnIiSeZVRdZa8B8BtT2TigVenuTmrPpWmvwOSPOWh5
OPMv0zZ+zAaSYIPeAdPz444uIH3A5apshaoFPAKLxAkbj8ZWmltYCDC1GrUA
c0HDo4mT0l9Vg2O4L0v+kxfI3NrIfoL6tiyV66eeAt4VZv6wVgVt458GNAho
P13wFqmCfjgE294tAabl2JADrV/VEaE5rpS2mKqtOvAG2+M4ce3TNbCPulca
wfi5Jn/trmzrQWsWGq/y/cxOkWObl/acvDQwMb8OVTF9+TF56VdYOOHTRtXu
JzyKgFA9wMycKwRVd2sB2sjKGlCIc6X2Hp+17D5UV1f/ygyqHIzQMrz/WqHi
TWRMVkxT5Pq03ai9B1zrTOPt737B49xue6gs5a6IBeYjLYbjnO5D6/T8/4/u
A/D7tM4F2eJXpwI19sO+abm6lQRC92HjTLC5prNyabjHlRTwS8h4pYmXKkWE
VT2ARH86lyDMMzaazq5fHq5dUeXw0uGZa5kaeso0cci74LBoQecm8OC50bIN
aDlYZf44GTUBJZfmH7NhaGwH3M5wEp4b5XclHSTHGYdGLKKrTD6gvpaqFhe3
oAezgbuih80PScui2kRx+RMZ6eMItMH5uU2wEDE0r48zXdL6RXC3VuzAj8K2
7p6ZitjUKDXkxCjCUb+Akg++OCoCgTk4n+6iDECJ6R0vSRufqVC+4oEl9xo2
4AwXNPicEMpfhIU5OyrsztE1OG8E42XWTUrpByflvHS1nOv0Dv97V7QqYR1q
ZocOfwqnam8kU1twRQSVqj2JvWR05NT5Fjz/0dMNuwe5aBAV3H1fyZ6Ylt29
Tk7TowOK+Dw/lkyhCv2ihu3Le55Y+w66L+MnmAubJlsYfK94JObzzJvK343+
J11Cuoe3RRLjxO6rjj6UhwSUhhSPq4nWHX6Y7uRqjRZUdVQShRxf2T5POPBF
S4c+SZOwigNtG3k0eGw9kR9v/MFgBbJnqDY0kyDL2+WGK2U1ceFBa9CzFwfO
9POpnc6PfVGTT57NI9+dexNCSYjEgctRMW2nTGOBGoyniEOXoQe4t6fNAFGM
28b+zEI+zdQUuMPmwuxX2uqn+fBhcOS2FT9FW9no/wPo0fHYZOA+Q10izvvY
hHiABgV+JrSHf60XGyrZkYIS0HaSJ6Pk7butFubx+8r5ZPlPbV/X0TCUYVzm
BxkjnLrqkKI2W8koPlT3rtCvozipAAetXoWvqzjxHrRjKqXJxqaXBfCna8lK
9LVHhzOUssIEJX67GFjJh8ikTGN/ukqmTswQ6ToNLrQZ4uRnpLo6cMO9jS+d
dFOMgPT/u/zLH+6lqfgzH2NHRGKVkQINcElnPxeGnh9ouqPJ8FNpSl0VvK3X
tLG+xtLi9p2BgxLHZ2lSDgtR5FlANqUjXGzTu5AuTmifV+ThepFHL3Z/voLI
S5B4MNOj/vM/c2sjQWdbQGAs8wZ3YxwBmyou3LyNO3pPOudZFd7IgIyhihXb
Z7N448xaDDYItmRDdLRX5NZqfmauP3hpYRUK0/itVCRGND39JyVxZPsln7rz
GIONKq3FZEIaZV28brolTPRTcWrgdEiqYC4UPYnfsqb4if2nGCmtun22q9KL
jWq+nJCM57Ys/00+d4Yie7p/10E6JHPrnMdkCl48+MJ5E1HOfQXnie6g/FSM
YCwSutm2d6nPtavb713r1gZde/q9IqrZbUYThdEUYefBO9ZCdagvhHVcvwMk
XCa2BQ/QDI+LxWc/ElDGpa+Vu2Tj+Kr1+h8y2DVxS2/mdk7oOgMzD8sWoaxQ
VH4YgRNdMtG5iubcyerA625WJAUFxxJ/Ru9jnOj7RLHmiypybVXdM2G30Qq5
8ce+9tQ1u+XlLOTH5V/cKbMuxlSoGu59I852+CsvDTINd/f6PpHcNXMYGTCI
qURRtVQ1bRuZzCKTaIfeNfK3OYqYqg/qrqUg9+W1jw/Sr2C7FhR0isTucLV+
xfw9GjCgXmmkSGVVhqCD9+VvB8rzcOHposWrpO5swOQ67AzohL/o+oDH2ZNt
yr0pnV/06djgX8WtIkZbDlyUkpbGqY1A/+U2BDhEm5U3iK5Q64/oQ9ajRlCt
8J99O6KfTJMWD5zncAXdxH3U8RfLAMIHijom+G9op/i8Jn57jbCM4sNxC3Rw
AKkaNtB+tkeI5xpEhbCXH36vafFsHRHZHD+tW/ujwi/SW9OlQUam4CeCE5zv
LZAm97bfWRhRYqxOdQbY65rWxJ+N18Xs2dBZ9+b+ZPcFjKH77i9hLkosOgLr
encdI3lrV3rRn9J58GpPDZAUJtbGjJArfsrA05rol3Q0EhKTXX/0+0RcBD63
JvggtCQw20QugPkFJro9NDQbm+VbRFE/Qw2zNQ/G+mc6eQNeKH5lNJeM9hMG
0OjipE9tjcGXMAYRMTwfxVxJmlbd+jPrAbXzJmA7HEnnTFyBx/BbCvxisXRt
iE7vVeIYCCjiXza/uG+cOacpW5nGkjpewMCb56o2BYnclOT+kXfbAOkLhHfB
kvZKFDPU9JIR8ehpH5JcUiz0hENQ/kqH0LRS6mrmbWcbPX8RqRj0WE7PhloV
ZbD6GuHcOoNKT9sPNr/28aN+bY/XOFK+rlD6MszgEKo/21RqS7N4Z6ye3mdM
AI5vra5M+CmuwOX78pVBXsKM2EJdhsNYf8b3W+J4QfRuF7s0GiVchqqJdX5y
Wj8Xxuhlnmj8nut39aPy0DFBYjVddE8iA0+byV49IXqGFCNM1g7I/au/tR+H
9IGgQu7DhmjoOoiNnH9bOlWe09zKDfGf975WAc9A2Pqm51VSO4f0hay1MXgb
wRMAFSOUguu3gNRvOyeTsUZ12ZBaxEe1C4TIULfjtZ/+lKai4kBajAZbwVy3
pziMStRQJaZY6T6hgHEPq30gtCCfReszikFH6zAkQ0637vTy2ppsIXzJyhaG
cceL319nEP/djMsnG3B+qZOUxIc7X37gO+G5yBsYK/s5uoWbOH5SFxsK1J9y
h7cOEZwbZkc7L9XhLU+qAg6VQNTf9GPNVvE4ZEB96+WIVxVaIXLbUeq1QM8b
z7te4ffCjIu0FaWmFidp9MbbJXfcuYIiTtiVbSo01Z7y8I4nEfIakM2Zb4At
ITxzJYwByqZqEWY6pRiBbLVci005mGht+ab+GO1dL9ICXD3JJZszshyiJ7Bs
yMeoT/4raz7/T+OltKvljXQY0e8o0aXr7LRftJEl6mLh+yiZKIlGHOzKqjai
vw2xQC/SeJ0zpM7dM0vEUGTFDD5ZVFsV0J6DKKmyIaEMIIUk43gfDoa6lL2h
8FLQwVbfbEwQPK4z4MielYP4Lo1/IBgfgBn/pWyO+c+xUGkjfjjClCwdpqLX
3+yJxg2ZK6s5W1pDhwsWPs7AXa6C3LbxYEzKNpgBLwaqMvJu0VJDU8UZDikQ
kfLlEfIIj+XmfM96KSYAVm62/tQb5mzOiF1vnwApWbJrG34KvPK3AIFR3ncH
nn/cfeQXKUfh9A6T3PGJCHVhO2puyUdg9yidzBy3rNHAzd6JUvtVgHPTO+W/
Bp8leEFrrtB+HgrNxAnQMRbZMJ/BiY6CgY44I8QiaP8qhEg4duiH7npYXmYT
iFBc1riZXFttLFrf+CupvlCBcTMkZhfyb3znpWz5a1Q+Wz6dYrtYfAKn0qtH
lVLfFsSymi2IRzAtbkNy9fx4XI8e+6qPjLUinwA41XbudNJ+lh4naGpaXpJG
oY79Bp/Sfp7xe7UodZO1uV8dC6p2GZ23ZzwTHqygeNNT97SpKbWNmB4ZVOg6
zGoYvLHeUtx3JXgKCEZUZ645W7DkHPmDUzcW10R3lIyrtckb9q8PSl14bVRG
eCsmS9mVqYnmoz+zD6/s2A4WM41LYptp6/d4tofIVAHH54o0kgiNSwitb9VC
iY/oGdGOeIi3tr4InN1Mlki4Wn01GZJ6B9F4jCPxXX/WIIqFnxCJ0grzuHWZ
5gkJ/3Pywltxc42WSFivytQBAvBGTu70w4GqFK3fbqYrtkpZ67E8qoZOs7kc
vjWYY7uKJ1KtPtPf38Cox9vAa6D/fg5pGu1wjlZ6F2tJMA7Qc/C3mBHvpFRs
7FktWRw4IxoZfegMWtL9NRCH7q9aTFyIgTN2314dLBmi/PsprvQieFw40E4q
ad/taao8B7EBQDazfP40uh2IfKaz9pUA8/tlp+WmyE4JdRvPV7rMNYVsIlhD
+1gph9gLxg6/78KwqRZgLl6DxVvACA21B7VUXdIcrJWTWX14BJRxfWZpX4CN
FHp8xW8LdwMiE0nXkeYcrvqK6dtmRtFw/gfQYf1p3firhJyjeq8hm8vKvktE
wqwihkD2rMaS+M4BV5Utz/je5ywJP9KcbzKyDmlPLMnYbMnCWS5RTALHfB+3
342XJJqQgwQuYYghdu5VfqaJnHhnXJKQ7GXtotu3vvO2f9U2BAwSxPsIfXiK
VXlDw4w0J8Mc7WKzukIwjR9IFmA9FgVGEZjaT+tyVoQ3RuynG+HqhgZ3ftro
5H6jRDy/6IJ0lHRKoucimh/ZSIDVvCHiwl9pOnVc0LlqQInUuF/pacjX/gXY
u0AGIu+mrjmoUMWdj2vXpIVJLcAtI74aY3wTSBvxzBES38f4ByoinANHVSnz
aBthIUJCYWqLpsd4QVE/ZCw5TgtO/Q743hU2AJy0xAlc/RhLshyj/8ZRzoL4
98UicxU+hxBAIzHRiJT+2blxU/wWUqPjhgOAKe/m0IoDKLF5h7ayxYVaL4fT
Cvqo+7Ynu0L1bPNkQdQVS08C+PvSxu8ekBPLv//S4oa+CIjVfZr25OMKM65B
kA+wcaa5x2RAgsXB2AyhnNNDx+pPsa56xF0Ofx/CqWHyzZUi3tArm3S6unfG
JWH47eal3Unv0wMOGLMNt0LIn3gWF8BXFAUx+6eVtt0b+9gCOG1wJKDs//bL
W2mM9/DGPEwUUH6tOmdO5OrETK3U+FZ2MxBhqadNl/rZoCzuL9U/1UtXFDsh
zDLYUjH0B9tPDd2+1VqIJak6PFN4E0GspCmx9vLyExJ7EGYfMp5ih/3dwElg
BT/UQE7pYCKFpw84tH27ann4Uwy2hHdGfEiezss1+//nE5vsbQfb8A+I0FUU
2agYa0KQHbSV30ZulfmeEIobjpKMH5UZu6YqGrkSL34GClbm/DWhT2eqCp+E
7cmUoIGivYMYEDYvHG5m5DQ88Q+C/oWdFljNHlWfhfTUPXYZ1gVJiyr1GifI
2CU6UpK/Xuyt/G58hXaLs6P4Wg/QHazRisQHKmJjy1titoc9qiKS6jZRKvZq
hq2Jwdy0ZNentbnkJ4fRY5y4hO/JFXnHHzTiNNnp176Xq1oesQjbQABuDvoY
fLyjnDrqFSxU63GXq2MTjSHcST3pSlOrxCDORP8hvybHpRLPiXyvTdo7mhHz
aTmy2kPQTqvPKxvkp1Btul/rMz1SmQPYQdynjKSL4vJ7JfJQ6GNisXKRfPIC
bf9ltCg+V7qW7IfN0kPMQhDFoD6m39ukRDe7Rbou159987lWJ78VqkcV+5jz
fhuX7b+O9TnAkPHAjeOhi/PWypB3dXRQAHvwTuLrFM1a2jOxDKNpx90txCyL
TrjqE9vIbY5CNOvPVZKlFDT+R4byUYOugpP9AsHxgjCyImtK71PJIoVD5McC
EQElLPyIxY1u1SqlX352XtLiOwh9Eop9BeKwN8cLdM6vdGHa+BQzDHjtem+r
rs/FXvKE/XIkO9pvd+LDQ/PtKSpFMFK5r8CBLMpdsHGyghChBGR38ra1fy8j
c8V/mWLR5+JYKT4HBU8KjxNquj1bxcX7pWaOB5XwPzvQheX8Cw7IFoJ4sEAd
WhdK0PJhPEqAGeTbgrVeyVMtuZyJaniEhkEaM6FIJB6xlEMwCGXQT80KbdeD
Lj8viK/VMHeM9k3jFJMXNApyGb58BMp0wdcqP2yBCsQkAPLkfpFr6M20uDD5
3d4NsKU33xUth51Bw04qqp43FhsXFbc9PBQ8D5AvwBTk+V8nq2Ahd8L53zpE
9HkE+t6SF1scXSrrRyOD+HbWPm9VkpFFgB+BuLHAkJIYSRA+7wk2U3kxhS4s
5lHMse2TBsQUE8ayN8afMKK3qKMICDsrEcrKVaquWqP6yIizkCN1o3LBRI0r
zljLcwhzMOFtfiWlLnTQrsx7g+0p0PuY3cr4HVlAqj00S5MXXzExcVzN6US1
f1AyWDmv0RHLURc+8cJm6ofMTAs1obKcHm1Zh4JZJOSbWME0uAubmnN5ES80
sRhV6M5/ZiymSGSYPbmX5kTPlitYWx0d2khuPnDFcePROT/o2ZZ6HzygCTW3
HHSdXocx81ewB1A/sFZ141f04Gv4I3svp2KwpbUSk3zs8MVogbKswZfk2Wsu
H75J8LvCKCWP6t83sSWfGTM8fnB3Gkda8cFx/J6a/pv9PNm3/qGC76c/2Guy
lePuw0IZWQuszwsqA5k4uijH+vx4DVibK/CUhQ3Qkky+1dW9tXd1CvDxtymH
tbJQk/poGRXckTWa8dyi1AorBxC547VOC/ViO+qUHgTY7oGf0cqA7LjtO7uf
XNbuEwAToOsMTv5dhHwRBNu0ZRjjMvEVPOvgIYDdeiTxMMCVhjQ0bV67ejR4
6y/ipZGOArlMd3JfM+R1ClN4dr5KgK6twWyRPTnKYNPYCFBCmrcZjcWOkZPq
fLeSQnIlJXU2AdpU/sMP9SIg2/s4AwNc5qNA9o3bkwO3KfHDJw+dFLdx7hxi
YOqQHcN0XDvdrhpXjjaJODWDhproabCY34Cho4AEmFb+ufFlNlLZd28DqiKJ
CejpOt1BQ12RAWn3iG32SLJsFRuXRGUK+MAmd5TaM1xb3F18yVPOq64xExNJ
h3z7wUMR31kthP96ZHNXP4zfbsayTDudYF/A1S8ZRMExdD8aHYTCvmGS5eNR
Zp7RY8OXoI48OkMtthi3ZGo32o8AOhp3xzpNffNctqBOCMhGYPm/HmGr57lM
mjA6DsYlz06gRKQnm2fcC2eills1Yjyf2YxXj+ssoAec/gBVCydtsOTDRxhH
AqBEEdWS1Yuyo6zG3iGOmz2/q4ZJvjkzuKgh5UuPG9grYLXKwAhKl0z5x/xu
QNaZFizfOYSKDFG378z3RxQZTK6uhzRdfutb6VAdFzfXZ48GvIl99RQU1Lmj
PMtoxZCgEF8Zp2XQXeQbV/3tmvoJWW7Fw8FTl2C4JDup0kaPlOOrbCZvAe7q
OD++4BcN5LdK1J+M6WNaapUj7T7W7kw7kCk6B1uaBvu65mKkr2CuupxjcmQe
C7/N8C2IWHlfz068H/gYRNUWaYDdTY4cD4sdzT7Th012IHFmeAJ1KGh0GU/t
eDzV1u/RBIjflCaeDZ+cvNcE7aZtF+kaQyvbfJD/bD+sJYnAhUZRCGuHm0mj
maL47EwCHhXIbjmRFvcKdU69sHx3nhBtnxewENzrBmJqc7odYja8mIeOfb7p
sK5g2qcuk6efPTU+UDbWtK/Fm9JzclJUOptgxYFY4ztLm8QqV9TpJ1RcbIQJ
XPWZqC5vRTQY1BTwU/fxqQ3N5U4hVeukJXTMf0dNuumKlNHEGfDigHYlZcBl
7z/8l0oAfaiKqHNaudcKpI1Wq3UPkO5UtdMas+3tEEgisItKYgP8iXWSRuAd
OqxWTMw3NjNbUJPrLVjpwzEZx5qLnKHAOQ6UaDadhlRvFSOu54AAHhhhKo1I
UEeD6ypzgwdYzzC9WXH1ZsXGaU7X6Vglm1g1EcZjZ9jh7gISc5p9NZa0kvkf
lrFyw7dW6PrKkKiELmCPkiyT8j10Yy64SZBMiwSYfnOIBGbErohCQuKTQ4f2
5x2y0K8qE5cpr35RoJvvfy/93jF+uCF6LPv2ZaP4cdlCVngLXkox+HP4J1Gm
X4Bs9AMnCyKVgD+7sJnfGbjPBm1CIjzorNao0+w68LE91h+z0SgnAGnnV6nF
uxfpWs7WUGsM14CK/dL7m/mKBPDBeOjzsr+6LNMnn95gbBqyuh8aS0gT+dUj
W/EklWP4M45GV6HSgX4y/OxcIbs7rgFQeIzwq6CiTQuPs2vDrAOLr3HTXrgs
twHn8o96O+9/ZLALNXjP9WfFpygYLEhCFT0Jl3CMWlXAJkfzCaOkpVVFmjoO
Wh4H14I/zNfM0N1vJ04OnkgYsOADHoYH33z43BvXZt/dII87Z/vnLqzEt+JU
TkCBiyiufkY8aooVwPkYvzgTYIgqnR4QrNqID6Hk2dwfdZ3dlMPvs0Uv4L+7
ML+EX43zePY+U6wmR7J57VBrmuyDY6dYV9NkK/5BktUbm6KD6k/VUSloI0Wd
X9rt4uS7ih7UafXFm6sYjWqSIbmqdkedyPEpo8rJ4E2M37aDAzzTGkmZK5BZ
0+D/N2vD93q2Y7a/ZWLGxe7RIT5Ngbb+tktvQ92weuO3a9aKllDiTwF7Xv7w
Qfl8HHDXEUv0bErwDX7DcP2za9xpKM4UDR3kW596/65igsACo+VtFjUdovnc
mBowKcqFzxhTU38OxCSBHde9rdFCDaCQ7AhE1rIsYsgTlOgvvNnKGTZ66gAp
JJ58ODjp87oAo52tigtAtxBiIzXlIvDHesdYwW6lPA7FYRVez0tG63oPheF2
pkr8cG6gzaYvpw/uflrtyM8G2eH6R4lsBjRaQuOm2SZxalwbtlUXy3zmAdVy
W46dcWMM5XmQHTAhYsq6su410VvLHvu6IF+qFhACnIBdslBU/hQYvZW0KJxu
KJSDZX1n3rwB2Nbr1/fSyirjYPRZd4v5kmLLFnAIR7RpjW9fgWykN2waoBmQ
eSMwa/KhQbnDaJid4ACebfl5vUpGZ7MwbaZ7dwjp+MJn9I3lEm0aNXyeu0Cy
sUSGvjgVwM8PKKfdtu9tNhnYHxpNPSn2ERC56Tk9crSsWTG0mxG4InD4Dc1Y
EMyFKXrfg+Bx+a7qHwouK+wFsZHy/gwBgnN6Y5OTL4GTz+3+rfEGwPAapgNK
JOMnfuKnKLhmZtT/p9Un5U83IubGMiJn6WTAmFTN+kpDfwtddtscu7oP1aow
IsvILoZ7xTH2CS7xjCI14vkLWfhZ/ZGLawVg0ILYbNcEVUoZyeYuObW0kCZj
UgQr84/EK27+fGfVii3lSl6GbnYKZnkUB+Xl4Op4FvrskU62K7BsIEP19EsR
QATSwoVDQ0kBx3szA4u8d/AjCV8I1e2E+MNxNG6nr3rzaX6UfDLtA/MVEPYj
gvNRO3j0NLcvOb22pVvKUzcmsAEpl294V+aLVXnV0+Ih8xOFtRaGOfNgZxNw
n4lLS4gYOv/M0941eL3OwNtkS+XL2WTFZ1h7+4eWAz4yKjdre+eejQiq2aX2
vzrbx4hjlL5/eWZmtbfA2f1L8bNpRQWf60/5ObfYzzq0SAz8OlE/kRWKkbTb
FWKW8enyIFkQVO6Lo+D+82OnMyXQHUn/xTbge0QWQtCLpxQ88nTxdsHkLbha
dokZnlcty9znEoUL7+bDkIwOpdx20aIIq+lnh4vD7O+U0IMMqoWcU+Z27r4y
WPfWinRT6BM9uHtNcBYJhs+VqNtFTSRzII4JYV1cmzfKKDjQIJX7i7SzNeCp
Fw5r0Unr2LUEl8haAny5Q81sIp4Y7Uj19Gm3/bW+uKmu8+Vt5AbI32UWG5X2
YwmXfrHDvU2p3NzYFopKGer6fb8RoEDs3Q8WS9n5SDSSY6jjEki7T8eWX2Z9
FS4TOC6MY3A2ii/1SDr6aE6hCpQDVNokdaMzRx0FGCqQ2pK0HfqO8S2Fh1Lo
yMEqua80xebm0THUVwWJIta7ZA+UhCJgYTl1pOVLSOv+GeDXBkvpnw9kLIsS
TpOxeoypqzFh5QysDMrzvaJ8JKjynMtF9uEug+yumoJ7WlTfNQs6YtQdpNYX
hJXHluMgnfIhIphiWReVXZsg5WpfCmv5kUT5K+LpE4UHQPfrxRnHxh6Gy29L
w2EGemWcJ291H5Q1xbO4uXWnV9QhmMb60ErUPPuTUIP2MqpvcVtBBvph9c87
boz7YDn4v0ZZc8y5XIGFBrNLy7Ovu4MgjAqy+shDGHx8ISyTXVTR8b7cuay9
R+OBTeg5Xfw2VZbfVNtulQb5IWBMsrZvnIbENsIvR1hg7o0/mP8ulqwfLHhg
ADxam3igimotg5jxzsay25fHTcJqFcIuHHlgQqpb04kR3C/xnscGA3Kq9ZZ+
Mix2YB1cWYYFfR4Krsd5m+O+zS75jVzmkxr6Jo5UCX0hH+IB3//kvyDoC1/e
sQRRioi/d9LSwCDvjAJyVQ6LUeLIF+lDo4eMkSwLJv+3/5lm2mBHUTUlZ7Y5
MMzROttmn+fEeOQMo0VGiywRr81jgjtCPYMN7kwq6QPA0/S2BvyFqf7Xd8NN
sWUd3IRXHB7VoNMx75eVUFPaGs4KvlbgDN2Ox9rGFTTr2jzxyQv9Mrx/ukMZ
qDx7kgn4rbm/FWAohf7ux8bkE2SDWUu4jQ9X25orXWJCFCJha7neVTja8/fz
DqMomvNTW1YwvYvpjEub/r5oFIkHycAdIPl2ElVnekCrNMYJftW8bqTIAh4+
72+sN/6g7pbvjHyFHaqOTglR3LPjUn1wXF4Q0r+00o7kx2iC2A/mpFHjsRT7
1fdxti2e/I7DQqR1ZDUgZT6CnFE7bc6qlDLigbFV6eY6qnkvvgqA+L9Dk6yw
f4Eqjd++NlezoDUjjkYjzZOd6kUjuCgTgOptjtysUjJvVfDt0h3leIm2C9lb
CraMkphul0vAMn5xqjK0Xj76Cr7a4scuL8dFOssLB+NfhdOlxaWHRikLdaVZ
6AyAoG7xIatFy+gnu0AURySguIkPUZzuPjlb364nMCKnroR+gEUEO9ZGB+pL
CmQWW9c3bZ031IlrSWo6R8zmY9K1+kp1M3IFcFwPbyF6tV5W5bXo4Hey9XFK
wIaXvtoT4VCl5Fx8YoKvTniDDyn3GPlCvZsGHGEGmHJ8lyJfJ2DK6du7FUwE
fVp89LptxjjqTagUkyTNpzXp7hi8b1eNbydkL9yDaUVTNRfPo9N3IgCnrbOX
D7WoZQqviR9XMPOzTLtimhY6wcIomJLrTT9SmA/0yItLO9PUqSBPbIhH3umZ
S57P8Sr55/zQlUh3BldkU7679aXPs1hV6Q9KNkmKMO3Z0+N7wYDTVfnsIXgu
29lgeSyBoXuoYjD9S+qtjAevhqmmygLUwkLngv8ANQDQK9IFjsAAdC7/aQHM
duyvsoh5O85SWBxt3lpZS1RVaoyatmDJARF/EVtwtaKL/WPl1HX7AOhcJN3k
Q6TNVqzoXd2pd5ikXCRs0dxmW1uhM6bhdWTtLbhr1uRrbQqJwuozby7Rsr0s
U4cY3wsrpxU0wb6RtG/LwPrB7rptJNloI7FiRK9of+hKJJ2O1tgWXQqQ5+w3
/CA81w5fQteW5of5gqaz5FV+yXbfC4KiVTWItA4iutscb/kHutLI8mPLASaA
9no0PAnnNVb+x9wLvbXIBYMJcgJHjYPJm+Q9MeZeruApKFCIRkmnwGmGn44P
kDwqGIoEQUUIUjRSrYCXDOOB05q4Vu4DopgI4L8fy6jsJ9kZqArOWqP4lEUt
OmGtLga1VQPWFa0ZeqC1QjiSF4BNQuHg//YZzpZwS4N/LjnSso7dzvnhx5/s
+aMK/c9/FR4jXz96JzZ8ox3djpZX5X4xCqeakFM7p8b9zb9lYCrzsBMewgeO
4UzVeyf1r0DjRyB4ttHnvbnEZnhGCZjPDsJhBdBllY0W19rsO5VlNtSQ3p37
pH7Exw+y6vRFHt17SbAaIEeaTS+mpuqHsszQKCvUAZotANr4bYb4PwJpU0h0
x0jHSWfrOY3D5DXasvcm4M3gHRSzhurNzpEhbsJ2IQ7d7P/oCCN79Y1+ulvS
PI6pZfwJlk+sLBZ+vyYfyOxY3sUMsXr3X2WvbQpRccZ/jAyu+cHVKbiSYhyd
DIVXMPQK3ckdYF9xLSoJXuVc5867vLa1ZH/JDCTqGKskUXbWaTXKi17LT4gK
rked4NRar1WnFuNS/HkfCP7P/cPr2+FIqViC4I1Nwey+q4UBV54Fz6H3jR8P
28tfXykalrYjOw+BFMgJSLMBbEV1ylHnKSBzvuuXnhTL8Mj3Wi4Bq5BITWSV
yEUZvx8TYEeNptlHpq1nR2nycMJSmhE91Ip2nYAcS0cE3sZmULzMUruBr6xO
sIn6387VQEFFauIDXEi6RBShgW2mGJzTv1OLmryuH3EuGuYFtnV+0FBtPa8r
z5x0u0f+mDCONJ/hhKJ8hm4wJcTSDSLkFUQMo6O7vh+2CxmZRCh6hpBk1Isg
3v8I6xYGsYlhClcC+6fxvQOnlWNBZfSlCtHAT9w2XDXJdsDOQsGtZeQfOKB5
KdwcGSHDil+nYHapksdMMV79W51sZxSfCzb4nTcB5cIMomtv0+b4GN3M8S1y
vSH7x7vOcYfEgoJQ56DL6b/Fk3YaQPZXk/soYRE44VF1g16dwBY4iCJW5y+w
4wW+pAK0pgsKUK/wwzdtFrrxzGeKleZNVQulOpSzN2pL5DMEj/9e4z+w3Usu
u3/SsFHdm0LMt2ZZ1Pr85EbX3SxxX/njnJgX66UOKFctlgrroXn+/z8568vJ
K25yN9hZDP9q6X3lL4imwOJhkpMUahDb7fyZebZ4UV0tGc/1Bfxd8zEr20tT
GL6K3hJffdC07MGTIRYh5gnmijRWUgFQaxqSgH/s+iPbkDcCNTvTHQNyk02/
XbKhjM7FZM3+w5pI1avNpUKj3bL2S/iQ65fU2xtToBopc4wc9E2WPMGJwiNC
eRrkOUJahbouTJayFF5XmDj2M75qTrh1exyKlS+BG2vEjN0sp0gpc02QiCV7
lwDOvb+PciyBkSxvp3FH5cr/cla4Suay+Zh2HM2pvXjrgfmef9WmPQh2Ve1/
eaVDnjnetyt1J+6SCWF93G/GpFvu0JKE/vFMNIxQS5FWR/gmoBADhVlXlg15
VB2v/UmuXupvDaULw3TG7+USZI0m6PJI7uS07wtwR4L+fTZvzqwpKRzsF4xB
kLFK4QyIl731qcPNrYFPuBzU+qJeyUWHAHK80hUqMQkVjQmLm5yGWtffmfni
cUATR/4uFPdik2lbJliXC1mBzQbW3hwjQHaLYiwXObiDapeWZ5o9nxNNPoW1
dY7cuUX1dIev3qIiEpazd50QaSXaDQUAbduQcliJW1fEHMT8gOQr5Qlo3Fv1
hQacleNdWRMo2K62+GuBQWkchbJ5eMjY13qYmBQREe601IT+ai7rgAank+jh
1wSL/kXTm+hv5vbP8GiZWYox+FubfN25YaRtIsiGhqKvz2MRfDeG8SciSJ8Q
eU5wNGVo9rTO0OCj1xOQenqYQN5nDt3+ytw8P9QxS+lXJ9cbUjIEKaqafSvG
wYG+s8iZl+VRNXjCDcq2MIruENyj8OcHz24S0HW744cI9dmWF6h7v4/X1Yuk
P25ro7iAM47QpiBrBXsFmG5W90WSs5o1T2IL91y5bH7YK+67Bs0vBlRhUH0n
H//AWPqc3QiL8O5st3RFMnQvsrx9Z0IVdIP6/LiDaPKRsybApZnGjaoYoAtb
D963SwrOOogI/2KJxkC/XdHdNS+zP8oKTkFildttg8sDXRgUNxBuGCyhXqEe
40YgeOr3bYXLkBVoxg7jMNZf6OGSSROoSJ6kUhdAFztmxaaz7xlZ7jqSJg4M
TQwZBQmzvpPknJ64qWk2yIk87qHgwK+wgNLWCKmJTlJkFYvopcKCqhfRy5yr
FbJ1lY+rMW5TaUAyTb8Uv53n/xSGFKOwd6eTXzlU9OeuhhDBe2SUhZSJMlH8
tKDeKLOdf7lZx0Ab8U9xEIXSpwg6SzWu6FtwkS3qICZL9rAelokp3p7r0lpY
C3OdGSCqoqtGfbublM0yLKnD3/Uy6ACZInYEJGeU36DBzXPz5ox1vQpsFdW8
iTB13AxpqoLXngKir9gmgiknYcJMu/fGMEh4kT1NaMba6htm/Kfi8RSPwbD6
6g3gRG7im684jlkRRlcuQulVvNfIoh6i6ex2a4PksuvxYrxvGK1Qd9VoD1RZ
cjiQ0Mri4BlHih+u89093X+L+pT9bie/7rKoH0ZvAUwD5uU6YawyJk6mTNvy
ym0K6ji4Ayh/GCyoGudWVM4uq+8xBvxJps9A9xw4ByMUQ3TmwO+8XotvjgqC
ggEKTQhAiItPWnfx1LFzqqhFPAzoSzLsf7GVPjCiEJNuAeozWaeXaPZRA/1p
p4Rk66FDrxWL+prE4+QiP6wlHEZUk7qbHROv/+DNmDookdideeOEtZmoVK6D
xlXKyPXCQwOXxvA6KdEiefPTW+29idQyu68uOHO5bGMWdtM2q0R8pPAgtHt1
mbok+fTjHNBdhyMcxS4KRuNhdQPgblq8PskCgAL/OhxMvu9R4Y75PBJrrdOv
N9zVxDfAwpTAHLui4fD9YYU862jh6hvetPL4pXuf6vMvOzmnBkze38kZGvDr
zUUXTnSGIF/K9JurxXepWijz6oNYyTLMOBFuMsBJpc5R++KZrbqoM4hZxqma
z1s9Eynmxkc5zcEZLf0gCD1xGgsQfLuJq6XsijBw4iZZGNFJw/tVrdp9CLD7
widcpHVvDCmO8W7kXqVQgiGGAEZpMMHAT0H94ZTJQyXb+gdVGQXjIfmlSSrT
tH4Q6kCVP744NgVenUKn8r6viqT7pgbHmXB4X6gB5CUnTHbQS5E8vvnIMhnz
xf4OLAtUMzEtScEhN5C+hG9GhnZAevJ75Hw7zWKZT1ALCuQ+qWwTGacg+9Bq
3p4YexlmrP7k1Gbv64Ab3l8BCuF/rEGXIqWNDVUhd0FT2FTF1N7L1MCte3sQ
zjs5IRyrjqp+ozC3/lKP57bPYc3ub792Fdp6YITm8aTuhyNk4u3gX7utU0BA
gHyyhnOV3EA81c5N7rJjJc381JRmmfGf6tb42IXkj2GnIfZHH/QgmNfXxUJq
5hDJSQblaH8hVV6A5Yvm0jLdYS06g0GZUtX+0GMKuDsrX7KNMlSPJ+IHH2yp
Aii/DPvehmmGtl4C+e2G9IgLjxPwaHYVMLNfz57NL1Wj+oii37Quu8Opqo88
oQ1G2LjU1W2otBAe4Wol6t9niGGJpvXwwYutra8xkOw1t/61jR9tB9eaFel6
mkSBjjjCA25wCOwTrCo6eSZAUgIK9xqgmq74PXthZnycZc9+JfPdhGHOD8Jl
DmLIZgG7qpzCWziJUMuq+ONrFtYpXekp+5rdo1iH3bSzwclh/xOnSmYImu+E
gEMWYl/WzhumQz0xVkIUPRvLBiktP0FyL6BgQAXrt0EKidiqcmGKqRlkZYP0
d/1w6/PlAnmmRdLynm+oXuy9lMZlbL445OJ4XKQzKVjnYHvqMKGdZze2zscW
ivt9mGuky8kFeeP0fVDYSBW7t7k/EN3cmJ2hnxGFaIhF/yoGONO0lbk78miu
nkwtbJ2kdAoqJd+NfyoFN5+7GgVYh4q9GneltPycNacOL2zJSqTGKruWh4Cn
lxh+Lhhwv+GMjOckM22UiiNSeDjkXF2ywxmLKDxTASxVTSSFrUVdeIRW5qC+
YIS2WeKeKbsDxbY54uQDfJ39UkinShBqFGhsnRE/dKVGCCWSHuvxKJfwLEkD
j4BHE7XciKjc2jyn/5TUJMOSg19ZHkfFssiqThAyq7Gw2B5+5zQPeZXX+qjI
GQe6heajuGHL7ExhSNzCSPn93gc98amPRWwAriJuV4/aTm9rp83rA8NdA8dT
kb8TWbjJWGmt0Zv3tOQVMbNkg8ZOY4p+b4k8zXOMgHjER0Rg/L/B2zARmYDh
BoiJT+FX+bwgK707Jm53ela6QHfgjDiY5/G+fdBTfr/YAOrM99SDkfGzvXYF
aPgtVJS8vGvZprDGek+jfmqwwX++8tt/rIM/kvfqP7awzaNKpAUs9v5ipV1I
4/SkEd0W77hWyLBWtl6PtAqH7d5Gp9vM5ORt0bsjGlnIrBy+H7s0IZY66v+S
DbSU/Pnp+EeOgNIS6FMXJfVLxn7vyZO9LXWw1f+K/6J2dyQp1F9ER7L0EzTt
w/Z+tX6ylYhsspTJkCX+70xsfzL4oIHHWjpz9nABeFVr7KTVAxyNhFO9rZh2
UQd+8ZQR7AwLoGJTvnh4TBxNblcxXUsBs04xxIULLFXhZ27Z/V2Emtz8V0jR
IrQOqVS1UqPKKsG4TGPj7Y6WRGeBc4XibRNww+fMId3F3ZwZEKyB/y/BKEwH
f+Qp0yKeU6I8eZlRM9Fz3hCsBWblUE2o6Sx/ONUpf0fvGVqLjiMt/LZ7xTLa
hcTj44s3aLWN+RqdhaC30xf4soQYQ3u/OnxImahojaZ4aFm9Q5JAanJz1gOt
rxKS8zyQos4XydKEHpKI1NTkSNLWyRz4k8XK9YJpNAJendbXyWvcdsYk2DIl
4/t5xUo+oVacTlULPgSHrSdXj33VSHekvjkKX0Yo67eHGe6+h0fu7citQfnH
dfh8Lzg/lsFfAOBqxNyGUaEJertiSVRl3nO+62RQMaIUvNj+NWxja1csA+5W
7OjeN30JwUdzmU6ZfRmxWHPtbW5LjB3Lp54a0oVgO5xhrqYHJRejycoPqgYT
/mYCvt5vIAqdtTL1hNfwOOGrShXWf2naCwj2DikheC35yag2OA+aLTjQytQE
Z1oOHnvSe+kf5hIKuH5KCNH4XAMyFk4dWRjXQMxSLJsmSfKh7Xid8keN9b14
kw8SVUcLn5zzQ2xNmTTEXkiU9C5kqTPY0XRhcwK/hWWyo6QBi2RRXc8hWVzv
at6fMdoPMTDol2F/rUqOa9WMxVs49PRrG7beu5PGzNW+vcLQze0q/F9fKkt4
/w8TlQ8cD6IFDQyyFfsWT6kc/FQOC/syQHsDwpwmRkJ8hTxX1j3tsl1fujHy
DO1sRs0gkRupzZL3MH5WKiFI6LyGNe7mfbO/xnp8Jb1AZvwo+cpJt3oyhc4R
akZnQ6X3uXs1rjSIEn2m2NfI5GOp2X+8JjsiGhrchUGhXHKbsGzcU+YmpETr
jh5STJeu7FnEB4iwWGIIzpSTZobTdMUFwhDQ3XJMJDZgAimuXFwqgUNLAdp7
Lzpon2itIgW8ZMzU9q4mO3zkS7BAE5CpisJV23BslcBxsYMCMTTCsvCMxfFi
oqxOF2uZUY3p90xozXcdcsAQ6SDhFAS13LTulP3JkjtBVaV8INN3y0CxHdHi
mrFeJ9gbh8cWcgKsxXOUzdYtPk8AXm+aXiPcpxGMaoBghLbUGgjtKoBvHEc7
rKJ5ud+s0YCAEaEKbidydyhkIrg3SriVtvo5IMbQ+gLYldOU3rFFAjdFsegD
+aV+OxwRHXIdr++yr4rJ71mKs2cnfAgMASuw+Zx4PGaRi/cBNxyNdPJdSLYF
rZazy8ZekJnw/YCI5k9IfhCh89tPHyVqzJ1ZzrQtoTZARSiOVh7Z+314bXl9
cCdhrJfrczG8sCBi1DXzwynbtKSpRzCaObbVRnEniagQO4UErzx3kuOIB2ch
PD0fh71jV5pSTPCqMiE6nUSw0f1sttWbMIPQUJz85mrNKlbXoeO81TpbWZjo
ciX9gmGYZlgceeI4IFDXuUKmMu+mQwEDI1NOrFyKixzhGlRxcQ9VKItyBNdm
2mrAc2eXNfZlqYG2Zi8Ji+g8AmOjf9u4qiwkysUwAG1GrzribXtNXJaP0r6/
IqHvOZ6P0CIfUXp5tGF5C4W+T7kwan+OZ5FFX22fnDRicSR1gCPRFFGv/Gru
IdOmbJ/u+VVmCKgJuKpDs+AS1z+UBCjE7qNjAamDU5j/2o9e9sFBk5fCQZ9N
3cNe8MINvEkzfecqkxsZes4kuTmGTT+lsbrjbn9fYn5Xnky/Gwp0tTWPC2ep
K44J8023cKMbiVtryRTXLjo1hzwHSrdVeTEmI8lE6+pbsCFSmBIEiy/Cmkls
enQi0t3o+hB1ToI9iCbrIXnirIxXeQFt5z4frOD4CWs6bVQyyykmyIraWPbM
U7y6XRAfhcfpguiLICcyGEaaEC4W5iPc38l8h/DhLqtf74dGcFXR8I0ITqQV
mMEO48/ojOcbaN2fGsnK3ZvGQxWfmTZKIYxWIGtx41UEdyzAJqfSjGmqW1ne
1HzPSwkHlwA4dm7px90EfUxh39uGf5XDiHk6KNZmg/RkwsbZADkW902AbqVJ
h4Xr1gN3FG4tm5pTEssdIQs7utZ/bgzkgvlj1fDI34M1MDo2N54uxR/BmKAI
ZMJAWWGsoV1Bp/wCdg89c1W/zyjzMrx2K/zkAAmxob3v517ouipQRSVkbGMs
OTDnQ0wkcYasiIKH4sewNFzkOYdGdtLSW/6kBnmgBOQ7lJjfAXnKXfr4mdHg
9NG5+aYon3ULMjQf9a6yAhrIqAfk0LBMXmmo+wZNBKeJxxP0LHodT6pU7TZr
gNpkWOjNdCbNuwV5J1pusFORObln6DtyjSUP1rDbmUwZwfwquQbdrhTyZFKE
digE+8W4DHsdWVra4hdd7tlEe6AkV0ZQqAu7Coho5eigy4B9xlogK6adoGfF
ZDKC/RqcKqB2Hj8UZIsrhmR1DpVcrPd1P48HbIXy0Zzp6mk9XuyT32/ZG+aH
r+qNZ7YZlZgl8HEb9X88PDASJhGJARHa9xJ5mvvFltm5f47H7tC65CAxXfXh
KjRpany/z2CSTYkVreo+Spp+17FyHUEFSPQGgSJtRdUdRdimm2KrmOmKa6tM
5YgUSIs+M6gK5TvSTtDOFxm8eRPW4AhOyys6bJARCpk5IL6nFVV1Wq/en5D3
J6P1JP3ZRTvoXdo7X5O1wMzj+pDAAZjG0J/bx42BgNonQZxURdXT9rb6eg/3
alP3SkPzywF9T46R8ncPKxr3ul6LxrNsDtTFBpTxKsQ5KOJwlmniN8XoV+tL
ksMsw8XBYBZNcXXEqE2n21615gythlr36fvhqVkqRnrm9kneGmTOnWIkOuo7
EBpY7VRwKpHVHJf3Dv7m/1ZwpPGJCB4A9bdAjm+QLjye8v3o/12RfvQF6zS1
AJvJfA6QLisACM/H/mrSMGXGfgjP330JAVsP4pyDJk96NQ3nicHmKpf2whwR
OFfjcgPP2vNGluZCUuRqb9gyGCv+361bcwWuh5R+CDR/VZerkn4hNMzlnn9e
xhVQrXovyHHFdeqCyYrC2BiuFxJy1xTUzjP7bYg+LpuPQG1NZGv3KGKNVJ5F
cuT8WSkQaHlkr4AHC/Di6hNZn1bXE6zEkUDKECGPIFdNKHXaR6vDKwyRQRSv
wEKTJiCvxeeSD5+WDsw/JpXiUInDToiZAI3WggVRd+y9bMOp61iHK3nkd190
M0xLqWhvEaIsgrp9cEZS1qMVJCN1AWpo02ZaM4Q7TE4xd83Fruz7i4rvlFlb
Jo2pvI7ryT/Y8ObUS1LL0mUPUylQH3EPykHUKBN5XED2o+G6YWZ4n9b+8FpA
Xmh0aMBvlI1fIkJfzyRW5mcO4DVjX3C/iH5P/dq33Gj4BLLvABPfipqyOYWw
8fx70Ouj8KUYGIi1/3n6RS6fjB1No9GoqarsnEzkh6NBYCzwkb36IcRWxpNF
rhgn+kQID6o9cENsYrkeqs9uZ0axcPOO2bi+NYiz5fejs1FgvwoqN7Nk3vD9
k4NavUUA//Hr9arOc3kOwTo/03PMQlr5OIhaUNxibsCNZlvnuEnbQlJmO5Tv
KOr7zsjJIE7E6+PnhiRKperpu9g2p3aQD4lUWR584AnvqdrBJnUV9GazJv03
QN4o7gQmxam984EfbvpY2bUJPD0nq+5ZM0clV9aL6RB/tXaeujNFxQptiZHI
Z+tuno0vdWFNJQvaEpSgSZJ0ZvKsQmGoOJFC0fQgWEWtpPCiJB4p5A/6xnsQ
6Nq9GFeNo3JK2TM5Sdm1VnFRe/msoI4hMMTGiZt2pinQYWn2dBnuVvqQhF7z
PDt5Afnz1qEnN2iKQ1Bqdqk2O7weLkXHJC9YMIt+sLZicRdeh/MGIsfvksrY
4QslhkN6QkFYijxR7f0UE0NAD9HbOroM2EDxAOqoTgw9DI93tHVGWVYSXt08
pOwPQ5lMTQEc2gB2XaPQHhhoYPhgzoMHoJtuWrPw/y9CDUhUcdq2VJ+rXWsX
SEBlfNv5O9lcD4IZQdA6hGsU8x9uO075LaiOoc8zyvu4aOBOBzw5aalSyhG9
6zKXBjpu0lUktv50g2sLIhzcbvWtfc7wdnonR061UkgFFGxMiKzzmC5QXq8c
78rkf1uUnPiApgsZlWt+v89AqH1Pl20hzmWO8ZPoLcGWZEnkAEHyIP9tZVH7
i/kxkx/2+rJ75MXk6uzSL15igmWuA/MYwFruGE6o/jpPd8tIJAWEiOa97GmA
Aj695O7miEdyoK29ukGrIwdHTS2UXDLnn2BQPsRLRn5VM0TTdyfKqZ2/WAn1
Pmbn79CQ3OFgfFuV3sU/eLRp8ky8M2cfglg+52zId3/xMlJzeuGhwi6zvK4C
a9sqkApt7iDVGfbZjflDajm7rlmhtjlGM/XmlSOToqmVbWWL+LBCyacg9Z7I
hU742HU8k1kY+qcEdKIm/tzTA07f4QoEZH24YuJUgvmu93i9S/wkZe/0kMV8
bOpUEcK7LYG+Ikzt0E7ZVqwfiUnWsPj7erlCTaOus5xpzu2Gzf33c+S60sxw
CSeYHIy24D4IhXgZHf4Iom7euJQMX6molFjKn66WFmmvWco8KpeIUC3yFBrD
ivOAJYijxfjLCRlzRMtE+ACLOFL02u4I/iGk1J+ELDG0BZ1GdOu3m1cYBV2P
oFkQGmuLJ9vf9vxYk+2ka2V8UQ2vlup6uMrJ45+NCXselESognAlh/72ewmc
aQHK6RRo/qGkgLdeJcZVCuU9ckcZPeu/yINvO/2ydby1EBo5flnsnld98L8D
J8zQBewEMBdjLfN73XZNKNqDONoTR+Ovl/jRxnCbVP2N2Mgu+0NUbJfrhegm
NMN+GlhYetSqND3vl6Cgi+RTGtm73SjomWNDM4CLz6ZcPIWm7bypNNDl4xmF
Zle+HyhERvHf+p1M1zwa3iew1CAX9+QmyTtleRKWnVDaR1hC2DNzO3bLwhGU
Eu5azuoHb4DX64NsLsC8ypOfsUzTB2Pf0YFWnRJji2I0aQdeB8T/pP8bYe1/
deVRThaNfgO0fWzrL/HKIADZdLdtTGc7P/9393zDbeLheyPv3KhT5chGQ7L7
aAf0e7B44U/5h0VVD8Vmk9K8NUvLOeeTqfcKAjenwBuCICx67yAACt9Z1JLb
0kbB+0JaVu5RhnOAhKpp1RyNDRaeIZY/CCMRsPkO9pBs8gLY0+Rax30Ov8k7
mtatQFNJHCPhtuYpv9olIlRaU71VprP9u5ammktaQfOl1XSW+cYWtcuL94iF
S/tmGTc6uDMdi1/FnaOJg+YZWcZJxPyavF7beUvtNwGRR/OAOm5LqbHt7l8A
qwwp5H9Fsaji0rvw6AwlVwwps0BFMMfUkbTW5+vazd/1rwXfHnf4dmv8kg4v
keVtEEPbaJpDECp4UI7/YByPW46AwNyqVJo7T+k6jrkKUaWnrVKqXwGn5Dci
SoVKzLzXXRoLC6dMP199+OD8peb+TF60U/UZtAqndoog0/u7z9CnCmYvGsSo
oCHjCWWqoRhYjoslcSMsRWCbhpC22XQ1zU5kDw7nWZSSJu0TICm6oKUdg3GI
2XY6JucH1C0ZoPUxNU6lx4HsCRnE5YE5it1SvCOKlU+gcv7QzukjeRbSCMCP
G6/Lrud+lAcWYTjeVx02v8UhQtayKF02AOA64EKtfMBrQJxA5M1+G8CQftfW
Q88JeyLnb6Xt3XjX+190VhnnD6SNTarp3dBgU2pS+5CDvVuOZcg1HVHHVSyD
5qeerhbyAOHZW8gWxcjrSTtcKfmUI8s4wYc8CqpeFBpCyjKGEfEYchF0taK0
QbMVudOJAgNUb/DOHF8GOldJMqniI36gYiuqvzh8Nm4mzph4miVWA2G0NX/C
ujU7lEctkT1rFjDK4iJVmmHIrwGvcN7wzjlJV51sueiUlDo0Sav08ggZR02D
mrPP6GFLxUz60ZYkYo13WFjqjkb7yJ4SgQv6IxMoWkxbbwvN8qG/1j3EiwoQ
DDBZ6DTqBzIMejtE+bWru0xFUQ2EQLr6+vG29LAt93BZmBSp3nIVbng4FR9u
uhlwrDUKfK2/dzD+kX8M4A1hX7pQ9ijvnWX1wNBSrV7JenXrlPPB55eVtiml
aYQ48aMQxWy1anZW5G0L0PIBo4sVblWRRzXwQdrK7Z4qv0haLXMyUxPg8XQY
3FSHefxLBXV0JnTCGBiZhe/3TDoyPIW5Hzruv87YEJuAG/J4HAkUXPIitD9a
DTgtck6+x4e/5L0fGA39SpOJloPQNUDEi7jzvmtNEyzmBwpmk6scUDNjSd+X
5nOm0mtkKwkkTMyh+36XVkhN1Zbs5qu8lXiBaO/aHsh2HN9IJ1cg7qjFmCB9
LVeK0S9ywHeD3xpTdOJTynrdc9LyjW1WisTbYQhU5MvWbPqlzJJxvJHwKnDN
AIdNgvY2LMHi9niHRYB9y4aBW+hjlceSc5z6aN665bW8gtYLcNR0iku/pZD5
fUcU6TlIjHSoMecDdupqVCxfYcpbdUd7Wdmp9BocuVNZGJdEAihueJ+V8O3W
oCWEE8Acb+rfs2h3Knlms0kTC5CLAfxUebLs9WuR3Yktt3znQ7OR3++vz7RN
SUGPtV622o6VHXd6WwZZLeJ8ujut6EFgQNSJBKGOJHzRGFZDsxQfpqsVbQE9
o+nlZeacIDq8z4GqlSSbatJ/xRKDub08R47eQfr3eTKRX8U8EhhthLPqnw7F
jxi1MsslIU75WcAelTugeUkHw10ttH8eB0CXsPCf1GRHEhKUtfqQkE6cFJvm
wnvmLKBeyPjqnLV+Enow9bx3qe2DQxLlG6yoKCst+McuG96mJ827R46X9+gB
Yu1PzvLk2u341u+IO4VCT49n1Daz3OK0OuQKFWGsi0q94iMB3vP006GJ4U9j
/wV6hc6hWLb06oLO0Nc7lVx/Zf54eLgMjY6vq0UG36/RNSVPCflFkmh/7lu4
YX/0O6pMV1sr4vdYDd579GQS7fzR1xJJrR99gA+ydZOdYzrrl7JM2VkeWTBl
5VAaGKWciH6N48/mv6bmnSHwTwc2h9SNx1h5DWwNyW0RlkSYqxbrbfLZ0/vX
WXEt4he/kh3MunjOhGpYpjrqCPT+0vuBHHJ/FvkrgsiPVrmwY2tVQHbbYPb4
PbAz3nJptepqOjToImT2/h+pzclyVh17bXIDUO3KNlYHHQ+fYaMkADaJHH6P
ejFdD0KEQ1w3WR68+8z7afXW8k4W4Dcm5rKd4ZxR8RJH2fri8gFoBnU++KmL
Q8vPloq4t7kvxbM3/2MklG/w+V2E5mWrFE10sSzGh/ZYhtfbSYMDO7W3czxC
jFRv8C8qM81Ft7QjYtfsLOrix5MJlZIzafrlcTwPx19UC4l8NvaIeRARTqV/
EKdTaHl50GifVAE3FDXkwTTD58Sr62UPWF/uAPhekGZWNEM+MTSWTVTrdRAF
+3CzUDB8jXVy4SXhl7UrJ01jolAXcxIax/pqkYQZZVME3nm77jbQNieNdPz7
iVXGHhYXZrPcjt1cwPocCredD/cw9LlS9EQJEiqVzr7gMt0cPO7Wb8wRBITV
iQlokgtUje0Ehqq/fvYIGUSjJMW76IjK+feI1jPg2MPKytRbMlNpo6q9fdBu
+fNIzowgD7WzcGsYmHKr4/S6kqaWdRciSOTvWnKwyTxgu6+oMxR0rFQGEJCx
ADXv6LO/erurSVACCUGzrgQbjvB9E+C3GQw5wFnbqXLzyHVCSP+bowlAD2ff
YQXant5A9AOntKt7+6eeWk6mMKC8kKR4g1/CjGafITfAaKqyr1OqImNVokUz
mgh2QJ9vVkq8wYJyOwVoQCr3puC6iI64SlZ8QFke2huiPCs4jyDJm0tnD3JP
kwCd4HZtr6lIqIias5HkMj8UVL6rr+V58Qd5tsDEZH8BkKFECzviG0EtuRvN
NciI4wlZpCe3CZ5GzP8HmxUKffj9VVQy31oK3EohqFz+AnUPdXz0/bemM465
+9qgZGEO97Z1pu8ScBTBK+2XYgrV+UC7771k0bR/h4/ZcTj7TU3PqLBXHpH1
DsPw8hg5kVQ7dQPnKkXnn1Fr5pNUqMUSgxjvf4zVqPwNEcGldF71Gu4sj9w8
2pGH+y4Dx5qy6K34J5DQJJypv0h8Q2vFdpu+vQ6SkWcxM501ixVg0/5cSn/v
SvnzmGXvwFjDffTLaGRqPjcCYEAQ0hDgedvD+faEDRau8ThQyBxCGo0THcZM
DDvOn8YLdOOTLGuOB0khanmzf0OCf5nTyM4FsqH6VCNv8eppxgq+OyMCAQY5
fvEOC+rgQn5AeGeRTB2EY6dxRg98UUBpK6ObVCqgnnpFRM1WhTpuKp9zU1UY
wyO3BK5uWGoUUnxT/pBBwvDrJhpWAyGd6ZEw+aei/OZeYQGgCPGFqGogHeO4
b+s3il5ntKODPI7QQ5Rhdsp7K1dD5jasVoimHgiM2XOVzfe4NPPlwjrEi7Df
cYbIokuXJYc5Yq2Sz2e9woxPWN1XHQxfxn4fI2nLRho4mRHy6qPYOdEee9um
/rGDxvM8ftkj505d+oZMyz95XhgqHPNXFBD8QAIp0RcBuvDOI12A176HHy3e
EzJQGrizPEilGkdpEfE8/dlKyx7J31GWoyqrzHW1UAAFPhrWYod3z3ZO2XXe
WPpj8S3ESyakkpljmV77hMrXu/+AkrT056eAlOvsLbpSog8ql9U76NoWLR+v
v3EtC6xWibZd5ams2znaVdOt4trgLqm6EPZbDTyi4F+fDDRJ8XNAqTqaPCCJ
OtWnuVgRZgsE41kVJOFmnK4DMlgRbX0NrFrHYpNse91y5J0oR8+CZawzh4P6
kQk7X9FHtk6n9SZjS9QYy9l/h3rEjeQ5iWh9SMCrKsM826zgYL3LWOzfDzvU
8xyhJ2x6f7ZZGaPC4uAjw1qDgAK15rTSWKuTTyw5jVS5+GcwLiV407GOYAh/
pzK6T8DxkY4Jdf0moyybGVLhrqa6O9fJ4PmVDrdlGEa5Zpb30rBYZ5e0R/cm
WSZx5dSscLNjzJyk1iiMOi68Dhj8OSmxa3wi/MEtoSVzNgDvkN2rjIpKot5C
dwjAR6VaH6Nu1EcRXl1dxW3ZG7SVQi50mruuMf3NHiE35+z1ZejODlTGpS/+
9PCbyfbh+X31FVwGd89ae35iMQDpC7LfL4n27CZAPrbR05/Vemb6WzGW/0pV
6I5DT7ATy7rUTLu7C6B5TZqQI/JCWY4LZKZTSEfcH6JEPbG/nJASPlAgMMXe
vYZTQLi8May2AC/usXARSNkl1ikxcv4NrLHFZkp41Qt10Nrxh7lYYHEK7E9H
9ooJ5OlJ4XZ0h8zPOQhWy3SU3Eamec4piSDEz9vsBsMQc9H3Hl4ZDJWYS0/N
F+G7OztUlQrfJoZfi0YuFUiMsEuJKtTKucWs7uFzNzPww10TW3pEfRIPHMaM
PjOUeP1dgwOa0dJlP1kZLj2enTLOa5dLw7MZ+ok3I31l+zReVDbbdUm7SFDj
KqVNalLWdHMwvZsM9EDGBie0qB46hH1OXpAaAb778fL1eKOibAsbPaEmcrKR
Tx236McReDSd+bdwQMQ9G/A3VR+xvSx2H5py6mrBG/iLBBnTRO5bkh3Q3CP6
PnURuV1f3qQ7temRFsZldulDozC9b4r1WeeLzUs4PAbr2RO9m78ON/uaGip3
TQBOkOtKgvqkw1V3ICDRR9BntX7c3iiNIhvBdhY2F5uPRq8u4/GTvXYVKkq2
s+grY/0FTMUz7AMSoJc3fK4DUeDoUPGEiC53M3RLr3aFepLnDMcZuIVGpULP
kR6EMgcaA4iHVzd8BcyEhITiFbUL0OZ8W2LBCo42RswWkeaGqxYFEnmRqLS+
YmrHGCXg4nu8KlqbGIgP4eYnhCSd90GI8O7BWUtCcIKfXAku38I94EsIbhn1
mpSe6JboLw5/5p+l6H9J+WFyV/zUqE/IB4PuzBP+8GAZ9zPVXoMO3I6hoQTt
7ZTIFZCC4vKp3rBMCOtr8bJguHYYg21qUxklCratbQEtQ9RWz5mOj9OnuSho
jUNs60aP+7hwKPP1ICnTY2LwdUgO0S8w/7RqmdWoFTMjTcMzAx/lcnYB7JwP
wKeeEWGWNUcb4rcugwZz2Zkbmgyok1wf+7GFbXhltP08ARAZa4AH5nsnFBxd
b3I9X0ofze1ZwWDfd/KqPvoSUBi4r3FDMSFnBuvjKYWLPvbKfaBZPPzd78+Y
Aij9CPIXQiY6lxy+xNNR0TQumvOytrDol4aF29pID5FhJJOfq25pw7keV1RA
fb/yXd6fMHTKPy2/OqrPhB8Nrq/A4EO0jCiz/FQASAnFY2/xc/fy0IH5xW1K
0zBIC+K48+bvsPt7B/yafJPzIsqvajObMKvr+0qFYG8ShCXnFjrka7l0veL1
AzfiGJZ3VPxXnFenJWZJZAjALKpQuuG/XNTfe5K+B0oMrsI8Iu7UM11e4WFG
G00nFYwm6d6qRCc8EmtOAUbllWI05ll0M/UAKV2nscuKUY4JznIivC92f0UG
ViT+0rO+hV81rcK0hBesDKD6l/Hn37ipcrF8P2DhnTq7reIhptBIQ7h2osLd
KmL1rGLMxlTM26ddbMnrwWwi68RVESNDUUBGbf4qAVL778FJORzvNGrAHQsB
k/aHv1TqvJ8zq/+BYAB6pmnvfxmVaAPrmxZG7Jupi6wbff9jKB03IcOuwaDz
azDfGDIJ4H4RZkc5f7w96KOw6Au/4TnIzQjk/6Y3A0WPLYc7ki97u+TCw6Md
PIsLKIoYBeMXLgRyg5ILrXcV2HlBzL8k+OuITuIvej3k92fhIbT2A9H0eyaM
u5Fg6B3j4RB/D1EIT4o8N2VS8+E9gc0932DBSGgh6M306LaWfXSuizLtZtsr
iQY3kpL4mtCbzibV7nJn90SfQ+t2NLjE3MzrLqyYy8FRQfjtreW5dQr5ZKwJ
aw/pOHmdm0NIwd4QSK9YwCG9OPJovauZcCEzcxyhenh7Y7qf6bFoEx0OZvgY
bVFbd0JeEEkWpycINjzPVvhg7jKSICFL8ruPsUAZVacuw2SE3Gl7K7mjisqw
6/cEFAWACGk7zM5lQ/WPIAB2NcIuNTc+y2QlCoxDZqNZYTgTyxb0axCobdr5
MhNZbL3GbwEepbsAEFZwfYImPnmLx6n66inhaC52ehDXOCYTd5qX6OCkjjI1
D20DQIXRgNoXgQqojKEVCZb7pO0fMJwfqXqYEF2F4ENiW9lRMfKlF1YZnike
YjICycU0DLNzKla92zHK5ide4tJcWYDAB4DG0gzHX4QRRN1gl0YuXlT0aWIw
ZQ/u0spAaDE0IXtwPeHHyLVF5v1Wsukgtrm8fLmP1aoYD237c4prc5+8cx+i
2MYuNy2hYiLBbr9YrYT8B9ZnEacaKjE60dcauvRRgTZxwZ8GAnND8PiZJb1J
LSIeLcolSKwJnILASKSEGolpWEvHp+HiQTq4ampF+TR+s7kcjHatp0MWVZoO
l+cDTv/TIlcZ6aEqSw76ME8gBlZts35sG0m/KKSAm0AgsI4fp9o1PZ+eRl4n
KB9rgYAUJHaV9LMoJz1+uJzGaxHzh+LH+WmlwL8WkanH1mrAojbXLAmYLRSo
UsTQqScPLh+2BFQknKze3lnmHynMz9Vvmn1iMVcq3n9gaIKkIs0H1LQ75PdA
IL0FegplTe89pyomnCh9KeOZjRFR3WcxxF+s4AmAGp/CM2FvRzWzn/9QWSI3
2e6Tr5QalCE5RnFtDKd6zp2xH7iu/ViqfRUYytS5/wj2OHwQ30vOQtbwA8TR
xOiUjljKvfU9CYaXF4itYoznn7S+Zdvrqbqjv2HXDgzC+M1pTmOoA/LAJdl7
S0PtKtRWDYJkFGSAtbn1U1pvqUNorCAndKDdBB/mFkXO0R39h/5STkEBII1m
z+euQW+9FSyg/9mIfwNwMpAnb+eM5FQE35HEH19CWZo7of2xmw609B3BqPh/
FXAeoSjEwfCtG/c/zSuIaDtLR//r5D0VJ5h28ecXlw82rL1uUImKS1b6KoaL
8/vMNbCJx2d8vDa7+I/dYojVwnb1/oJV4sos0Wu3/q5F4UEDfZJ3t+oPip9q
dQxT+Ad+O1YxYqwOluPY1KyxhRoFn4a62XA2EDwC67nVHy73hYaAMzVDTSNe
pcNsPmQUVR3WldqxWmkdP/V9+IJOcTv8p3uuFDn910fSuE2MomcMp5xAT0Vo
CMeLK1GLLLm2z5fGlRNpHZVGAZ7pgkHa+y7yucBSTraCweWJ3XDunvDn1V0j
QPpqV3I0WQxbXyn14dzZbf7Wq5xya+k1A0AosaEintDprXg6WCwafYCUlM2/
y/3kGEaIE1MU9p0cY2IbA3wnqJK1wnlmAOklQVvsgmzCKp4D43wLnPjUcdHb
3YQXwndEwW8F3VpauAGhsonoFjsQzUiVlDVB2HyeiQjufKPoJCmuRzse/qwC
Bo9nADIschNxiJtasCuZJtbrmi5ElII5MMcB4Tg2GJWIfhUWN5312vf3YqOo
3QdojVJYYU6UEuyJfH945GAD8WEZutQX3SwgMEyQ+jTk7yg3mEgI1p7BjRc3
ipvgdV4UqPXUkLLHUbP0cpRZyaWLAG6/M2pFIuvi/RsoP6VWYO+gaMK48ouW
9XEzDe+PBp1cUIR4YFlhVJ4nouIqtoH8Yx5ypS6weTEHtvMvxzw+KQQZyeag
1ciHNs3jBUQ8kDrPskfb6W4InD4d4A6kY2VmQIoKbT5Yx9dNmOi0hOvisN+K
OMWmYfJPAHki6dzaq/ia/Ovdwz2eXuGndsxV+PB8fSH+n3G72T6yGlWZdPh0
58eYhHMhpRHGaMz394DZkwn18JVaUoBqU/C5bXLUYOOx4qto0BS2IoX/qGYf
ZHTJ63b/KLoioxykTuPjX3RKFF4um8Q+M+/DKd+FlHOdnPVzt5M0a5XtcNUR
fk7icUfL4Os5rOJVpBiv484DSy66297xW+ttd93ra/q8LYkzp1lQDdurQeGM
QvBLdfDNGUEhz9hTAxaCBgOXh/tdXqeCpyq7+T5IBbO3nDU3dTU77uvM74AH
X66oEgoqcbP/fkTp4/onSAuHL0FE64VnIGQ1ACU5G8uuQIVD30BZ4ZCT0ZHv
9+JCAYAHfr7TTBqkMVZr99cpTNsmdlZ6ZhgfkJYnhQS0X65UMLgba3ErhaZm
LedwJ8QiSK+8nwiYgDgkLCQmrElxPxAc1l5TsdJShhGm09ladRvyN/vQyTXQ
d+Jw+7fbMG0imS3X3QF/eUsylpWazeVxJ3qBmC26IT96yJYYScNtnjmvrJzX
HYrQVnPkgDG5IYf9i4ju6knXrbC1sxrdTlK2Y7kzfx0rPPWTs/GQ9E7xqEcK
TyllJQp1i6QIkf9ZUdMt1DlBhYY6peZMvCLkYr+4PE3CE2jtLXj2lGLR2KrK
reozwcE9YkX1CQcroAavTBjK/fblw8eisXTDg5tUIWbORzixwlKZvv++FjrS
2WNL5VtNPaAtC2gTYVYC2qmPYemrANSaHDygYHZOYONDL5r4oDOxZzQGyApn
TvD5pBpFv+/5pWf/Lx7O2Q6JhvwGGo47hw+FCYNUU4D1YMr0IBcZ7L1/k5ZB
+wnmAQLw8H4OEdP6dbedHPvJH7GukWTsl9qgh3vB7olGlvlgTRy8NMpDIVPY
/omFnJZFAyBfHh5h2fehMVE8U83ISmB8YcOBUNzFzVKPbhQkI9i/DPi1YPte
0a5KN2daVt0tRQIr3/vP5TPkxkgHrKwVZ/H4evxC0fOoEzBd2S65jaii98g2
MCJ/Wk+V8Wxdx8C6N/E5CEgZfVhwlir5maMWsEKoQWQP9ZLFs/gubeyyWxky
eF7uMZl+lape3mtes7gEtKHIJFURMCOTP9u7jJ89pgaqm5UtkXEY1IA4Kcb1
DCRvUHbVQWfAT1g2D64P9uaBCpX7DW2nshOoKIAOA64ybzTId358C3414NPj
oL70pUNqpwLVHNLORtR5HI/x/+1L3MDD/VqCC9Ea3fwSJMO3KfWWy6gK0h7D
flDu4GE+ZFKfdxltdlOXWDaFgyF2XKEKR7nbWSJDQdAWHV9J6MIuawGgfeYs
bbVZMmuauTW6sjpmAMbpqzw1nQVSme7fKnE2Fusf/YY1C7w1E5F0mZR/6N0T
y1RUVnzjXIQygeBZ+CszlWG4mmJnoC301zaHyUpDddCLRwbxqbRI1GlcZeeF
HdjnAC5/4J+ibyZxKFSHXjmIgFuF1zwuKhlBOqHXc44aKHByW4oh9xUdHOHv
v4T5GtYliH0zZzprkkkclUotHJnyPl3575e5RLcIv83F37w/aF1aF85PiUx0
M+fCHMCGZE53q2K7Ix1tPRbT67W7R2K6Tnt2g3QAMmhoI3Zu1WgL5AA/5EZ3
nhhresANkN6My9ENjnCWzRMJWyVfB2Oa+I8QJrIyuK2uTWjZMG2Js65RjDaP
CdBb/4vR/wtOB36PoO4VESMvxojm4zCNWTqQP8uWgfLZ1hW6CHWkEHJkf1aC
H40FZmNR5c0DBAP8fAYA411ePYpb2rA8YtoLokkTPeatntG13O2tVulmXpv/
QtzzZTap22I6aP4XunnoDaNogbJDmHHy+fct6Se2mThLI6UYlk07I3K9vEES
qgQUVA8zGFVIyztyExrzqkyPN2xS9Sge86GllLxD2dkUxIBygrD7Kp0vzY7K
UAoAULvc854PB4e7DrA295SnGMlksgkXvmDkqgDSuqun3doJfvg3Kzqdpteq
IWToEHmavfOP481dazEQ4YyA/OZXcSQ6ag8uABD/RP31b9zUtbeEqtcTWTHS
mOdf4jrp2OHiRmjvID0Bhr2ZlSNuzMkZB3GxcVNpv3QC6pC0+tc7Ea9DloNp
1PZLwF0o66UDrvmhSfeSZNtgAx3egDzppBaCEJsLjiY/jYUwvp7X3h3p5dBl
xbmWbznhwKhUdsI2nex8oSdKZjrEItCxk6wMlgH6OU3IJFvVV5O7A0psZSJx
JZKEviNulCh/9JTV/65K1M82JvMMzvJshjCvqEa8wh34tbiVcMQIjtJvZSro
MxoKPhpTVyC2FKOxmOFN/7mtqnthdZAMpBTIpbyhCq4a8YeQha+NE+s0n0hf
wjE2kY162VO3Tm25IewB5DAYihNKMlPLg43dCX69CfYhCIw+odkfpI6QT9Q/
fzZGLbnR1NqfqpcB7AQGdsgDJ31NN1rf7ptAimMHJnwUBgyDh2hmvj3XmAt0
may9gciuEQGxSrmIPr2hlCZ3OnGDgEyfPJqaiA4IW6lIjs4zLxOy1JjhW+Iv
acibPvr5cFLmBS8MGWaNuB/YQ19vgXAZp8x5TSM3vGZ5EjzBNHPAdbXpq3+d
SLu4rkgN6Rjl0acQWJ3Bsqa7jPUnTcB2XZ4GNKBwWLrwRNIfu0333l+ssCRr
AwJHHoOrdPfjLE4OOwYumhAYHNjcOpeLWUPMqEsV6BdMTX+26LILIeIwnUZo
+7FmvVAskPq0IbQp2vrxW50YVe7lT+3NW9JHaWdb6tPDCCjfJgcbEQ++Zr9y
m/zaunfKR/nlpR0BuluWk1ZNEbNT7+6cPRO53l9simmMDosZLOC1K2wGUu7f
IyGaRAQcWzGDPQuF8ApS/IiGo2bcl66xh+aU4fURb/tI6fYo3f78lUKVNMn5
Fx/Q4Ko1i6p1wZPRxziRWH/cAFI3dRnIFkJK+1NI3Mh/R25zhC1fX6bD0Kpc
LrYe17JJDnxMHfpGtMW+KjMG1vIRieDZVmGdKEfWzqDiVzGXB8pdaJJIjm5U
gwC1WXNC+sl37vSsuMBY2xd+mlIYVJZ8MsAx6s1ZF61jw/9uNg2MLirDbt3f
vqZh7yqzmpLkj6yi1nzcklmIRHyHEbbugM0T0oLVuFe3givtijii5fGwKkIq
OsTxMTvfO0bCQ/CAZQ+fzsJus07sakKVWy63rN0/SU/FeAYAkMj0kmy2OMwN
PZ/0D4Ssj90snxWC1LoLLawqkaYfWGaHELJSjjNPpQcqgDFJFgxCexJy/+gK
Ig1bvqhaO1pSTExlM1BaIdD6OvAiQy88/I7If7Ja5GLcn9OAun8gDCRVCBCa
9yyrzP+L1ImqX0S7+NqXYm2DG0vtV7HtenZon0XHgOPaIJ5qrArm9CyUIip0
t8pPA00/7mJiUp6EBPtBJE/BX3Hp/0/cLW0iVFaUMd41c7KwuzlJksKVtLcQ
JTPpHp3H7jqyClLITQyNuXiKPi6xlxpnis5iqok/9O8iz7JAkLfVeFEnsRiK
sgHFBemBPVy8pV2vomKu4lv/PHR0NTacnj1n+7+WxmItqmsDadL1B+zJP6Em
GCHmXBOmROcEciYSKrvYY/HFRmICgC9LWjtdxTl5T9nnTAY6cEoaoT136Pci
VAm0eRKAwopmVAkGhgr6i0zzs3zcTrIvjPO6+CcZ+l+f9ZsE+VSEmBHwdyo8
NdcQfxiqKj57nhO7/U+sfmREuEeZR1tCywfqnAIkxlpYE7v11rsTIg3u+YRU
aQl4WLxy/fkyhx3HSQ3TJVIyPM3GDIJ0I1ZfTsgq6GV8XdkG3eunqQa5bqmX
ptGzHmn0Tfhg2PEmfK9FinlnCnck27h9T9nr6klOIBrCH0/x9MXBF1afvI2K
Xo3eyIxkvNNh1g6eZ8x/JPxu09PygYu3nPr0HRWyfEwsCthiSKfIxuJwLi93
GHGes1b5/OABM25z65017amCvPRYJA5qc55t2jYCrCHxE99KY1urC8bN4gly
hTWydtmRWualkvGI9q6hbagrK2FjZKBU7IklBCU0dqJUP99BINWKcFJKIM0/
DeM0TfyuxFzrGjZS/EH48Jn8V9zBLuN1kGQvRUldNZRrzuu5TeoCwONz8ZNS
b18kwIpc7tsTgBLQSg4/+lWaq3CF/V8f5+gpQ1/btchO88bJtZW/aofnb6td
RS8fexX/FAq45nYQ25ZlBPRKLZ1RWngfykAWJK6tuwba+fOE2bzvz6mImz2Q
6t7SaXgKPZ8Ji2vHz5gGAPHeTJA4UVN8qSRzOvkpXvPML5XaMWV+DUDJ9JUJ
b6v1h+IrwKDnWQQVpOjkEy/VWL3FJNZWVmI6YLtIJDk0dLJUG+F2APJtzd/0
hTUXvP5qN1vc0hLRwxNlC71DCLgee9pGRTxfnlSo7w95Jj9hiJbJNGHaJ1DT
wBM8DrvoVdyfbWyjPsTNBNiX1pHdNe+0PcEmEPGjYbBrp8VV1Vc1AZFg1Zen
kXVg/i+TnQ6gLGxIO16yRJ3x8spOrBRg+cflVlocQH1swMoOI74yd1T+9C04
MaABKPycKQjV4MWLLFxuisGvWg1QQjbPsVBbd4d3nVyyixrzthCihyz2rfwA
cPQ1Rk7rWDpkZmhSTdRRDUVI9Yh7lcHA8vXJyTEejmv1zk/feE6vRBbeth98
PdooK5YagIc90sb4/ELDyGZOR1+CU3rRUHisXh4yxgI+IB3Hiw0o+VxwtUDJ
5Pihf5iDQeOW5Ej8TnToaZN9jyQwexb8Jb3S4wgWWx3fEyCBBtz+h6dIMpq+
XyVkMyMnYS1+VGtCp75fmrI2qqzxxisFHhxaeXsWOp9YPdqsERAHvdxtoLKT
Vo32pN8TwWZP5l5MfJWVQgpelAIJHii0xQRla+LUNVly6efj12vDHeP51L8A
RKln9kuAVssBf38IDHkoq0wbUpysVe8En6pMvaiWoaSUVds0d3VE11/tPKze
xhv8Z74uWSui6bcd10PZRjsldPeBmUKD+s6Toj31vBsgPZnXyTANLcL1LaAf
hTUzSZpEt332H6KvMhCiRGjwLu3ubtWt91WcwVyZ8nY3/bRFKYchTzAlkAwB
iSjMHz/Q45MuyLMH2Ef14waXCPSchsPX/KfiiIaEpLJmw27V5w1+1ovpxqqP
DWH90r+XU+C+kg578K9vquhv7HCvjZIEK+WRQ1ZCRfeN4ySs4SrObA+4CYJk
UVZi4Irxu8UctFIN33wMDEjmRX8gXC7XVgLApg3wn1Y0ivFhsaB8qQxCTEiR
2mz+eDk+CN9lRUYpablet2PH9xrsVDjgluXqG6iuI/UKx33GAIJ4aoo3Mb3X
By7JOj63vJ39Kw6uknCUiGsC/k2c+1WNMJCMLXQ6AHBxPio5Xtc48FihQOhh
pzJdqpKfVgpq+/xY8u3uxSxwYg5kDbt/ON1M6UTjSJ1L35dwAzlV+UE9BHeD
wYjs1CJmZkqDbUqZaY18RlyCrdN3beUEkiWUTXTXbVovtc7TUb8rLZbdoDmK
SaKkEpWOcajqzMFMtgo4fCUYioWx0PPvYN+WPeePjkXI32pPrit6L3B665/7
S/Myv18Ecs/5IPANhbAxZWECf1r9Qtb9Svh4I7jr49Y6lPJG4oRCJlJcCRyq
bPxmQmbfVZGQ+YdMNXEBhbwYHJT8qlZaJXlYAthrdpzivo7BZk5Fv2jfz8Dx
pOLml0hoE9pmDQmNAXb2Umhc2Bg33u2kR53O5zW7EMOrBXcrQIR1tom4qKMY
zh1h16gnrLwQGNAIGUZ4fj2sf6Km4FxYr/2amVwiTEuQnxvluQxnyANzTOR2
9g1ant3kPPYbGuF2L19kGMGByGXfq+fBmIsvj6fh2aTKmfsz7xjKIi+lgDsj
hnMkObi+UZEvWPk9fgXX9VmCVFfUaSZgy3B8k5fRDEhQZmYc4rvaEMLL7hK6
MpZiKYrpo2/AgKmgynw19IHtd0l+d+MChqjn2ZWN7fK0qz5p0HRMuNdVQlS4
nt7SeBRi27HSR4bvPxSYzExlFTeqm4QyI/8bQT1gcAPoRgocssgniHo6+XI4
vq9IpjL8Cry9He8BLs5yu9m71Ob5y+CvkKaSeNCsq3naB7hG7vk9cz3IN1Jd
Um1qeE9vBfn0BgyX9hdl+uR3XaaO/2gshSmJpCrzQ7Lj2H8EEwK9pzNJzcyl
MQwH2H+j4+ES891L6oPNtjuxXtoZKL0zWyaYXKcp9OppF5qzLgjJjUpp5sTd
JJnbnYvefH1mjR5oyywEym68e8HGQBeZOpmqhmgEkpNEt3DrkwSgIXjbkCjQ
9W5d9bmA02/FvPHNjRap6rHRH4hd8qHsE5xJUKUsXhECLuy3EMZuWII5ZtzC
WNfjkLc+pA9S5jNO3b/gdjuX97m/MdO5XqD7i4t2hGQsNuqPiy2d2m+e8czD
TOLiVDU1Rwjr2Eomi5uCS3yea6/Sa1ULcMGZPVJmYbCW7ka0LJ7sjaME5wLv
RYOf1ZLtXNZ4Go1Dm3sNjeeiCV/5kKrb2tjKJVoZkyR++lW05IuVkNkzeIHZ
TRBmvg/ud3wopE1psfgkyAjhim9m+ERgDfGiqRUqGWPJIayxC3nztBEPLLxg
V2a496ZGmjrsdX3gitrkMZLh8ENeroV1O1hqYuYXSeTqFjoj7jlXSCunrEKe
gOW/ybJaoKTMx62HYqaT8qk9OqOcXUIDVkD2oeqqSdYAeKFa2cnjIL3p68TC
COzrich1pPCQ+iQvdQmhwyc4NUmXoX9UwCzUyY+HtmjNVZmPstKLpIWxaLwT
qRqW9pltlcl3fVuZtZIVQz4cNkiMfz+j7R1HRUSkG71hVWCJVcEloi/vfpTH
fOOzPYk0koHaQ8pwlCTqonqWFqsiZyYUbczuiX9rOI9hi9JZC1bzw6jBjSLY
hnMv+ZBBCSvKNuen194auJNKWl31RKd5yOPiIzCC9kb3d0wjVRe/mBuS+rlR
pvfX1kK3/YOM/4msSm9C+BDU1ulN4K7DFPbw1V8AVuIHSu786582LmMpB2xy
ijWtXqv1gEVWY85qx/GMLlGgeLiNl55kUxqexXHf7qTgAaTBdHWesczcO4sN
RzvKv190YxFUVaRno4DYL0HPhsywqlUaJNhIhVe7BFS7gL12tHYnqoOJn9D3
MnoTHMzO/AHP+HoJ95pxUI8rzkEhlg3JLD3vTIRa8Nqd2JjkAkA9uIg/JywW
gUHWIzUuDn/RhZwj4Kid91BcsVKBWV/e76CZjW4avL9nx8RuwVHc3xzvPrPD
17uF6WEvkx02XmnAVNtFMZg/RiPkg9K4TxDHpUW4g62EQK19hAnjPlaeCmkE
LdWcV5hiIDG+J6hG+BKswRZNEisvxswXGnpyBTQr+A6ucqvFqq0ZZEY2s8np
4Q6W/MBX16HT5Mfm1cqJsSfA+TSujY+SsBg0Z4Klu3LzRIMDJfI10i581jDV
ECr2NOLW5jBYpW/yRGZx+Kdn772WZH4zNXg4i6HcMqxFvdjMlKZ//+LMwzP3
/wG5qviDA7C2O2XK7cH67OPH6Mue62aYQgZXRoaisJOpX6ZP0/NECTU4m4IW
fS2NNXkZd7L1zHy4Us3d6bxUeer8then+9wyGXAZbyLvL99IrlvBaLeXGK3P
0cA6BqkQIVPlZIe4iYmfYyi3HJlb1e61s4Xq6iwWVizeF3f7ARRW969D6fTU
VNm344MdQtM4k9MmMnG7NquKd+SxS6fwnBxhmuCyZUMZcsDMiHehnyHrR8BL
X34m2+IZbBJSh8xXi/W2NNWT2DH/OqQxaQqwF5qTxck45H+OxO65Kq5tHKmA
mTNj1sNWOvvqfeUmKOH9lBjJ+la8faq3N3Hl1+nt1HjZ+m1n7RDBkeRWqxJm
JVA+sr/0Cn+F1WhiLjWA1ym2lRYmcV9AtB8eTuGTSaNeyu5CXF9xZdl7fgP+
vohSbgtvcv0fqx5A2iuZMiWis6egYFn6PErdIoAaAbZXiTA6bk3mGG6d6e1Q
h7D1R33b3wbFYy1Vt8nhjtw6CTmvV6mTJk4d4UXJqwwUjw1xkB5Wh42Gaohy
0bGx8NvwJph9vyYxqk71nlCX2OWqr5bquh+Jg3CNSETz1lnyOAu3GLDM1Z9D
reWx6ym75DAfR6MM1tw+9Z7uGON88Jj50lOofrqGx56HIT3XqUqeHNjY2MdW
Z3Xl9JbsAz9i0dcc8K+aRL9ulnGRuCMtwBNHN0UvE9ly+CRQf/bEB9miYFrM
FObyD3KZPezMWBqAJGTqpYAU6KYtd+psOheMMjgJzzilFikom5KZGpT3w/Hr
SMxZINgk4v31AyNLE3WqC6GtkPumvCH/HjT01Ui3LVhVwoCOmVgUirxEyWCN
YA+W0s11IELA/O6le+g059cVzqEqzSPjLADqPy8cKBkv5lu2TG4BRk+SyxBY
yOWlfjeg1W013OvByD874JD/j0YCVCgmrZN02u45osl8ZjFoPDR7UeC0ywHX
RmN7BeIofEdc/1n/yZ061IoryvzgN1S2qiV8UsGOMwg/UIuw+OpaD8DsjW3J
CpyHI2HbBnxmRCqAnQ8cbe95ZT8/X2RcmZvvHSx4xv2EDsrBDpPu1Qex2p+w
Wuj/p9+8YUj/yFMfPIrNEADqxGXpmNmxL/L7neWatPqxqpVjPr0yB8/3/ea7
YhqdVaqkpWpUFYFQPzH4f585EUBb3ryH9Pk97VQTSiCNM9uhp4bdggiHOpG4
eif9F+capfiD9Q8+Qnr7gBf7jFfZ5XS4blOW0kGtPPawS/UuA55B0MBPZNw8
10QQoYeLGh/Zcri/hgD3ZzLzH2N44JQYxj3ygfuGNRabDhWeJEc4MKhLhIwj
lOpC45biX8kMrxH8V3hHm2GWYx1Ig1zDZ+G2M4QvUaoAvx6vuJ0wTxlNtK9T
tIFQ8NgywVJQOdSKS8PM7spiRBrwfyUefPamQ3A0ah85JAkLk8m+kLZ7dtRT
NVfun8TLdisz+W3fjq5j86PgLRRzvPMUMaP1G0kGkNqFKHX5DdZEuixmAA/h
7Dx/MQtbl58KJs7xWGW01Oo5pLEJsbaQdr2dhcLAi6j3/UWF4S9WgHvkM9w3
FmGurNFiVX1F/bSKn/hDwa+MrdMc8tsltOj+36CR7F2aR9j40jqk0z2TIpJf
GXXrKa/0QeM8E7Ayu7s9UgICj29jcXEiV+JN3qhlBbMYf9+n7wmJWCU1AGfp
e9i3tArirc3og6ztKCoLgJZ9Oh5Tm4NHRjD+3cfKp2S2PVcD6eqji+KQwcJt
UUet2WhPLMzVOG78M6RNC4jBGrnbBdtDDUOFq+stHUI37udE0OpfNjirwrEa
X2/aQbPsNIrHi+3NSJaUzNMRK2OLGQH7TRs6ALF+MzTvSN69SnSzU0Hai+jS
S5D9FMCQGU9AlCGcLGIKkiIsvE6uszMFaLZM9gf8U1k+SLK6raB/Har8KUAo
SwLN4LJ2Nh2ZVfHvAuynJdyvNttdBloSXLvE6q7gCMkakTIImAfxvTnXcotm
OhKbxn03nPW7742+zqPZJ4t2F7/gHbebVF5rRDRJZCAOJB6LIXFosyIPsr/1
KsroamehxmrS9XjpdbbysNjyhsQT0JpFXkqTmoZWHakcUDwocaTey8mqUJgx
MAdza9tUZMwCobrIDT6RVlelLq1p18AHZAz9RTZoQIb0sUReijJgq/XthePs
/W4AIf/AAp5t7t6gT8+W1iRe08Zkz6QBMMkqgSAxrrH2679mG5BV7sjCIRhX
vjBXYUpLVTKp037ApH8sZ9xeziPGLiBExiy/lUSWtpNN41U7oizkW9MfYbik
OnLFDk5ot8V3UhYfN65B03Y47WOlntyAFZXTZr7Nv7/spUK0mc8vFM5AWSRg
9Saiy3g5jv7d0M2I50dJDRSByMf7+jGn/JLvC0eyIol0kudgVZsRQNx9B+19
ajyrJsiL2by+MNPl7gLrWQkn9TYUzrTmfFIMJqUry7lS7ZrFVHBPfNTBolVJ
vv72sAVIEL3A/CsjVktf+qP3h3mv5Ye02usK4oYYD6j7jI6W2ybJIrQSp0FV
SAtjdsdAlspWklcXIFCas0jxsy2dD7qMcgPk6h0RQssjeJ8QUVAqlN4UpPYl
z/nXxoZ9WGBT/3luHfOAytdvnsW+0inmTSZADNdswgu0ivjVD01yYEmW02YW
45knDyzI+f+A4EHzTX0xTfeRVT2762zJ7YoWOybfIimE6pmqys13v5+L4CC5
zn9Wp64sOmxUW4Okln8ElZQ5FBzjveuklq+2tEMJBmq4nryUVNmJklQ2FkMp
A6/5ZC6srg8DOwjKuQKoO26SD9REdXkyXnRYde8QYsvcG3igg4ObNhA2wjFo
P2wjwzZ3MVNEp1QRyA11Dbv7RXhfqJrJ/NGHH3r6h6vVdFL3Zen5DXzxM9uK
zmOHh43F2x8w8o4URl2BvbGpM9wophNkypaXzVUdT18l7JZTjuohf2LleE9c
D8aMBzcq8RMxm0XuppXOZBDWONhxT9kj3JMlzjMC41lIBIYxBgRj7d5S+pqz
kZbVkuR/2MTCb/hnsXC28QQyUAgX3FfmrxEUTQGNvuPMW9YBKDG27NIJIACu
a429urVg4YYG9LJhejgEnUnWMVAbpOwkLwzJ6Z8Bf0BEms/lyygjrNhCLIQp
nrBm7c6AcwhHmNvsuhZm7xtFDWeQhG0vqCxueX6d5mIfNyH25nQP7K71dnxP
9FQNlXWV0Yu5GgBBPosy91ftfGUgmHxF5vZFfjqCPDdL2/OqIrEsoN1e2+3i
IM5hP64fEmJk8FxZ5TH5CcDHsd1mTeu/klX2fW+lEMIzrdlySVWtG2UGqUbt
0K+DaY/Rt3tQH2f3t1ge6HINzXriRpBcA7F3GiA/5RbD5PQ6LfQOM/oiW4Bw
uJnds3Gi5QGECuiF5+wDDE8FvASUIcrdFN6R4/+7TyGVbjdCE6BhyXxHVg7z
/mBh+6DushNSTrmRNi70xZaRfg9Q9bBnnOj49BCXNtc5NXJ88zzYFJWzCTjy
pB3LJnra4NF5Y9U/V52arePeA+zCKblxc5fqtY5QqdFCv/cF3xUFMnCnPH06
Q9yb7Ryeq/q314FVVEERQScibFISMz2EQbX74dxrdZ9Kke5IXj8RsdQFvEXZ
jCQuZtd5S2E6NqGiTZIyJACo35g44yAP2LqfB3cTlEJP5j7C1Fluip0e4tZf
gaSxSwsvhlTpJK+t75Qu3xxcMBKE6k8jDXs6zPZwYXHGiPYLCNq8l3UvQqyu
qM3i34Xc9UeSzTKhJ8SYKN00CMSCQCQc/c2GP44vcyWl2DI1zrS2ZDDfGvfr
0jN8GAJiCWUY0tW/u3Pz3PMzUGBrBClQZgLeSs2IRfDDowyV1jgiGWnSJAOY
doJCAa2x3kI1ukgtABJydyEengdMdNut494AT4i/qNom1JYkrhD6wXntdK/f
O+gtZFU21sJa9D/iWA0BypCtE7JXmwOsfWN6Grzt0gs7fEWCbEwx1FnB1bti
a3h1Cxg5fD0KuDdNlbv+BuBIcOsG41i5yp6Xm2QsI2jsYeXAqI1GfpzxD4vs
gxLkaeOQ9/QbtI7oL5/DZAPiYBzCqeyWSDNee8JYEqsWDMaqHjUp9klErPLB
6vhvhPZOcwaQboWlSuKMjgieNZCxcLwUxw8XcGcUMsJrQu0C5uNEJZtB05aZ
beNTQpY0e8vtDPJJmcjR8/sChE2MoydjMrzGdR53jR6nQ4b7kT41uBkxEGyT
HdGi1PvBgyS3qJscqeJAdYUMYiQajuID8oM7btNN76HFiNxAgKxhbOprqzE0
b5u31x+4RYJm7ELF0MuHYUMDm5SMBMIzTLDH6+YLTNHIiQZ4d+hUvDXnbr+a
Xfolvyufo3RbgVV8vREXbTddBF6xtDOY3DsBoTcWLirSUrrDI4LRB/ck2kbt
1whk9Rw79JczST6Rf+DLRPrWNTXPfPrh+2Wv6RPE5H9KNUvfpkduY1KRi8SS
YkQmDm4sv9AATdyBRKqWvmpgf+hXcHOkiSYfDE23eWWBZKHN9yDsIvSbizGi
ExwDli9kAhRYcDm8zyx6mMXKGWKRE2xVexvHSY4YRgD4goZ01z8bCuXUPFBZ
PD7SkBlZXtb1vreG7KLmSdwgi34fT3mL42WqlQMoWT23lUo47IC3HVgIrVpu
w0/K1NGc7Fvj7W/LYmxV4/Ag+2CF3osZ7VG+/5urM+E2k7EaViNFUa2VoPSR
YDdKCFXK+tfKApnmVMSHjH0xryP1zuDhiWpbdchVoTJgRy95kyJSaHa1SXE4
yUszKRmTZmWa3wrSlWm9KN7tZomwoDLfKD+Xs6BCceGyWMrf204CBEI5x73c
AMpXmkp05Ih71M3Z/HEh/vLhH9UVSCaaR8XfkemIgvL+OxRUfem0HrsNNSDf
IwlCmZaVZ1QuJhEbwIS/sNduvj6vhvV1YrqZjWRZXMc2T0Q1xHbvIOSLmEdu
l8bJ2gczxRpXgvm6DEXj4XUnSiwAcomM3et5ErYWXQhJvpi3/lKe0RliD8ri
2lKLUz/U7rCRH6MZ7ab0OhDSZD+cLsz3ZvZEx1Mflegluuf6RBQ3CO80k8uw
ICfEvOvoo/abQB2iyO+ViuEWhiQylQeKuSraeyKNCQl7kFAsg0AWO162lNNq
YLQ8mKE4NeCvg1i4d6G/LKhsL70hFH3O/sfZfAA44aF53eiffeJBXHoR7b4s
waEJTfEinFPR/X6gx1OBJ5JSknMjHzNFQrVEq4sFd+3MVaXLgiXsav1hZKmJ
+GEHKgk44qOEUPRzJA4ESEzmJ3m/pGRQSHg42FL6EgnadahbffMXnEO9VXT3
lCyASEB7As+DDJl0JRIkQS/3lbpdGeEQD7qfar22WOyYw5v0DVOoJQKeFklF
SP0xuaHDlTwuZm+JEQXKPJPN94ZwhTKxto5sGJOP5fLryeg0oPMFlpZEyI8K
StUy3SdULYO59OELqdCTWzzZOWt8GuzjOsM+2omTMz4DWjZSLwfVjeH0IrVn
1WU2dhLKMla24VEb4LJLu0t18XXbYp0nol10wFvJ7S/9OuBmAd0iq/QMftSP
h7flMjaZrV78JMMLnfGl1U0L/ZpUKPwXpcAupbHzmZP41YHIb6wEFOlE6khY
waKNO3/4fH2XKNZLkE+2tZdUUBLyx5WmyJBMuGWr2cY1j6pfL7/Clj7APlF8
ILu4rDRgzkuheSyDZCyUPNOBbe9omby/bDsdB0EGjOog2V/7Yn+egLXKv0Hq
6YfRWs12G9ZQwso86YCAWLAllYWkgaO8+hBcCQcIWNilE7a3fym7k27G+LUs
gPf62ciaoBqlPUCj7W7B94ILUVfQrqdN/vz7MA5GljUyXrsDajliN7/kJKyC
WxKnzUlr3HoyTzF3tmsG8GJSmh5Ta0cp1oT3liZnri4/8v5Ud2l42wfJRJ2e
rZ3fdLCEYi06krkoR2Wo4N92+B3f2Qx4yujftomB5EQLaxFpRhiHlhgF//vb
UZs6sObeZd/TXNJ/dwe+yQF9D0EaWCbnNRYrP8vFvcTx17TXdIIFpS0YJ9oD
VEDVrxl9RQ2yilJUK8qIS+jQFIcULmJybL4IaqTPQ0HN3sPB6wjQH7FN3lQ7
oJQplMFu9xlADPfWZFEC/Dj7U43gfsODjPhmX9JFQ2H9rYpMnlUhNxbVlH50
/U9gl5SkgAPwGmXATE5HveWkBmoet+W6HsuWpA5NEItUWlIg3rN8IwWrrx1b
v5K4SlwPsJuUggGomunZzs+LldjbX72R9mAIGk4nAYMGYMpwUw1gaLSkFshu
MB0lVCyz5n+l855m/9HBqhWxctuZDluPyZEtZUYmtT85Wdrqyc4BicqFHUhK
3/T104sxAqleVLo1BcHkNf4gXc+ZDrUV65jO4a2vKD/UHZkiFVmJFe9GGWbq
6MNi4wtumtG27ilh25Noc8QpClWGBIDmo2Px4LB3fmquRuNAhUum0CmgmX2c
wEdJ8K/0/kitWd2FxQdB9oDDJbmBouNKkzkoLjzeVaYYCWza5M0/7VpCZGWz
GzzSKgqOGGzyVZk1JDxEi5ujylNFrW9DQ6e06OzbX8GAHe0s2EpoRTd91gZK
pSL4IfV6V9S2p27VPJY2SM0Uar8RXsVycWuBlmQXvlW/4Rm7vzDubviSkco4
rYPkku2tenVTYnlbSO1x6T4Nq0oA45pkHpq3HuyYQNz150ZXz0cVtfHuKeBo
KE4AnF99ZR8Dw8a1UjNFFObT6X7o2WosA+nfw/2eC+2GDuHwfInG24maJjEk
XR/m9jgsAN3ffLm3I6oeqacmTNQ/OEs49+Xb8ynPGgd1nbhjpH/jo43yi5Xs
t/jEJvTeuBbOkmbhG1Z6ppjfTjA1d6RWzpghO+25OP7rXQeh+POgqjF7YEvE
myP7TUMoLWBazfunau41kxybLhDaFNE9vJC/9C1PWcCW7wrrv50gFGOc4Mgt
uwXHZL7H0UW0w5ctefbtT+ArCmobb3a/cZh+Gev8k1cHU/1Jqhf1O336gQxK
nfPMxTx1RE3/ua4o9MZfrQF49TP0GkC2+ZO26sDwiv0ueaKn4kqg7L46TJGB
41TUfiPHqbq69FNRhy1ppr2gO6yCO0WFKebGFJ7yV8pDzglmrLbS8EQ8ix52
QaauxEf0I6FcIhV536ej9mSfhae5fYfPG24C8WQOoHG3w57YjDtAFO2qmlQ4
MB2W/a+iyGGX2w2aLre7FM20c1MRDBdy5ZIyzKd5Xz6Q9cypNKR/khMrFQCt
R04p7UJVx84epyhNL9zKk5AlQV8QNTmGOA4bS55CsMZ2X6W8aZYO47tnxHjD
GBQ4REvlkBhHpkL+QTvE4vd+5QeNmneCoGQTERHMNGNPHrjvu5XiudqEHKh+
WbE+UlGH+abl5BWOH+lcr9hKh3xw8JmmRy6+aS5ZluPGMviqyinPlFDd4knQ
LexDfn2fNbBcr8Jdn0ln3kEbo/LzE+ZQp3phLipAHOzGetIo2sdH3tmmNkZj
Q35SD9hxAxR/PjOsERfu7PSYGefLvQuxvGRMcOeUm/aeEqr2bQHR0vajMqnL
uMz8LlCKfQqw4ok2MTaPFgAFMi1fiZtWXZI/fSnuiyVnJbOSPw6feTsaCV4A
QoYepbENksKA7X9nbaJJvCIm7wIFfAnY2IpQ8mVd5cnrLBcMn3NOM3+XB9MC
+7WlvzbAl18O7Z2PPFpUrOJ/2v2XkccpYJq0Fa+M+cXDkk4ews47ep7eD4hB
1qLmDnBuFjeGfAu3Nbtn8krIyy8YMXLBYcP93tI18vc3gI6xKw/ESbHI1ret
wJlOchzAzvq7SemMQlhJ+XwefkzpfB/4gVc50hIkajfJdfEWaa+prNKKH7Qg
S7FBzGOL7qs296KeQSCfEOSkFqc7ixFMKMbRoAwfk0nc8FHY10o5hRBOT9Hn
VA8F2cIPIjII+5jcViy0itqKDIcNXImHPj1O2nfXAa+uZ1+8YQAjY+fEBDn9
PYm/T6aIXevdUqT4vd3MM87BtXZH+lKuRHFQJvYpV+5fCrtRa5TjO9DKq/oz
wsWjOxjZfVBIpqSmMkhx8qLvvJ+kwkJftJiXV2CQeiDER2dn4T0Hx3wQUHKq
XzPbEw1xQ226IKrfmTyklQi8A4tMcQsieiLW23Qbn1MI/I62m6PQPExej/jC
igipgIwKeSI66fQuHfd4yL2Qkyxe2csbZ1QWA9Fb/3vtkArFBlSlYY0zbzxb
/cCd+uKMyVmch1Pi3OV2h91NNZpfz6GSUuqhF6yygGPfRAnmnoueAEPArsVE
1dl9rH38N/rQmmpXqBHiPub/R37pDurArNQHStZTXEjE+mi16VMbOilfZWBI
evzVX35/ZdXr9NQkQxtKTI1piTH6Tw7zzn1uH3auZHKN9Fhs+mLN2MjMYOqH
6HVQB1YIyod5PNoOZTdu97r81oAOOuTXsmyJnKX1CbbNjTMjb3ydnLdeQyyd
1Olj1bqCM9/r/0AO6FGDy13xDcxzLN3zrsojcaCguMcRvBowB/O9Wzmi74Sp
G323Td2KOQFTzXtkrOijcQPbVbQje2m57L9B8gGwbnpDaOaQA4n/sot6YfKa
yDUtLMFk3+nWVNM7tY5ZuAIcIp7VFcQcjTys5AfwDSXzeS6HmgU+cgG/25/H
j/oXuMwKuqu0zZtufJ77Bul+wf87KgPJFsgiOEOPhayThqz3VdFXra9WcPWZ
N0Kq2sSpKcCyZklh9rD0oC6VlwHWoZXzV3hG7Ysy+s2xATAWQGl3qcn44VmT
P9PfeJRA+F18x7XkPiIO3TevmCbKZfK5+vOAUrLrb3nb98yrWh7AGUgtuJe1
lUEM1oRsoc99RGel9atbCOyO2LCIkMw0fZ7GecUPnKwt0xRAFphI5pui10PB
qUxev7qQ/zg1alkqGUfipMWcFg6RD5QCecqCrF0cg80GQQSNtyG+OUYtmNZJ
egAV8Y8XoFYj3N5cJXLmiYjCnZwgoAqshTSBwMu5NBc6P3lEHVNXjyBKqldK
9Psjunw1v6OvZfNaUEZv0C5GARFv8kaeXkBYBUgqsW1ZidI6kcvmGPHy1FFa
ZJmp/TD5+leYbFLlc8KmczYreI1QAhMP6aHm9IfHgT7oOevQqZUq013wtq+Z
sRKVeEUquBiyOYmrU1XxRICckEGk2PNpuiYPMAUevbFsCCHm0zssISG27CKx
6bV9UDkkinwjxYFy/YwiJH1HbaQhUDTw+1VIwwYplGfeKOBrzPFuH7jKCJ1s
4tDOEatqecfgu9Bib6+EcuQgvmMNDhPahETxkfcoBjuG8VcHhsW1nkcv2Fmj
arW+2vaC1IgZKnPuImBYRfL3RXXbFXjjB2gB1Q9A9o9weTyCoD9wX6LivRPB
QQolDwAe3vUEkL7IcR8IuFjKGv6FAoRdLKyZ/zwly2ykC/t1Z9nJOwrMzeN4
hIH+uVp56Z5X5ODaaxzPkuqcTHVgKoWuNIN8+mNchpSQQfy7SdvWq8AuRvMO
pM7eVk+w6nETCMICusNhE5hWbAbnQWQd43/+bG8fXx55zS87RdBeNhia0pKQ
6I+x7MJ7IHj+Ipsq845b4Czc4baisGnLH9bYT7fSQH9veH05h5roPEwP+H35
ahA9rxCEf0ukocRGMKRzt1jB6WI+Y3B48zTSU6QL7hl6QM0SXtIWWUZ6OqRq
pmrZPWSSShrFig8wF2of8111tDJA5wwnQHfh4XKoCcsUyWG1HtBIyuGMNp+9
GK4yRjLJ+LUGxJ6dboKcg7PqDZPvNh7UfTcA+ptRrsSiNtT0vaU8RQuH7vj6
L7AmNv+sQpVRz3I2qzCuOMxAwPfCA1RISKVI+9KLfLa6F8PVzW0PpbB38gqj
WT+l6/u2Uqrk2xTDFc4peAvcKqWkqwcVkdjwOAmMeOoqNvZC06yS9CbdTVNz
yWXq7YglKkXkqfgYuQJyei2g9IDRRzezQ4V2kjQ5UE0ncq9eK9uF5DGimjKg
KBdvsw3BJC411Njhh1Q91BCHkxK9QytmG8aBQObeiWEBLNENOkMay4unE+iJ
0VsOPK3Li6tSHJIvS249kPOdgK1gRvyUkA3DOPD2GEqyaNeV3yOA/rISPxAA
pnZ6NdSK/11E2ySE76x4eUgRIwvfqpzzXh8agYkk59yR9ue6HITZasz+dI2z
Rlom57CebeU8zsYOjlJ8cXCXYPpJE8VpPjwNvqtSsml8WVej+7sZGt/UUQ5u
OyuPWBz7Gu5KoZ83pVT9igIxc1FnMJLiZGAgUVPogzDtHnL76/IvpeS7PR+J
1SBvCmu/dEoKVZeFsQPtU/U8d1wTzXIY7vjxlSrl9kMFSjaGK+pkq4NsodhF
5Wh57LwQqzhoTwJTEMq3VPKY9spuEMz1KvbY2zvbqhZvOZZmr9qnzhduHtVE
l2rlRZ3hR/RDrwK8+NMlILw4RNwK36s9qb+YVcWZGT/olA+JPtmQHEnFem2i
LS80gi16DiCCvbIlumPFDv/F8pSqXTw8pNiHgUnaaecA0kQvM8NkGpihdE3I
i7uCNgfsPnB/nfe5r6iao/wR8EebjAVqkZZBxBnzdzOiIN50Wv+Uz53Hkd24
CSeibDUVy0zhU4LtDvIVumlfPw06IYlTgESw4QpjSyvkIoyVhhIaeMs+OvRU
0ACKQoVL/9qLp/P++A3sqpj/SCh5sb2BA/vNLCLLqa+Q/j6xVwEn0h0hKcCB
m8tY/zkp9V6bQ7Rbgt+oDTAb+uwr83v8Ou8DED9X0gDjqFgiaxhpGxZ5opWn
GO8N3uWrr2TVGmbuUfdwE3uvlA354OCvo57/Yw11sXi2+6AqQfHsI3O7G5Kw
ZBhrNMClgeK+yI+r9WvEMOpDZGJ4RXqcQSMsKDkudtTjoKnbjT4IttlX/FHL
0iUO0xGUrwDOpjySWGw5asI4lkKnnqMsfO/ZdpMqPCPXpdBev35jVaecbMum
IpYRmgcv68AeInMvK/bUuN940edibKZbi0HdumAGzkkZ9N0A/PDxbsYQ+90s
3ioGuaBXz7KpmCVpjcLF2MqfhC/sXuc/+/Yl6Ei1oMXmB/gVnBQ1nKB/Bgdq
+Bv6N8U95N1g4AmOJN9yiMiM3RzYL8zUxaeHpptNdICyw5rcPTWWR0OFjQ5T
pCJ6mqOlRsGgr2qqY7PX2YUTe33fOvAEB3X7MdkaqSPb94jQ25jSH2fcPNtK
RrfgIu9xnh2gxDfoFm26jjBmVpNwkQ1vzThrv9X8YsIvydXx6ilv0Tdbp92C
KxgE9ZsPwS9chD4bMuocHTZ7K6yIR3PVr/WHlaEX+/jS+Vu75AUmdxvnzKwu
dTh6HqfLsfQWqyuhGLQEG0dVff7ij2YQeJO0lFUfD5Uq+1rKZP1uzi33FY8j
SxZo7C8C3bDtl6j5bIQu0CVfPstO8yq4NSKkuk96i0Myl5OoKK6o7Yjm6p70
0ZY5p//eGHInAfKo91YBtr719sio4H2uxTwjtdKt9mHzEIP2DbiYixTy5e9V
UtAZQ1TAIKoblrPqyf/m8rrriYig+1ikKm/+H3vrRzG4NOShmGquYdDX/wG2
Hu7ZB2ve6HD/azT/xbkBBgrdNwLYOoCQdpDGmbLhrrQBEkWys0QwKuElQTGY
mIgqosNa2vpsBt0U7JDg5r0BhDXNkw56TrV1pMuYOMIr1xF3VffF/rwy2M+w
sAxAxb1R0eevpMFHuvgoCxbfzPtz2pn84SIpBj2cR3WzdUsjc7An2lWOVPrK
ovZGVeDKCgrL+qsJzU2j8FB3rLhCRtHC90S/GDFxeDRR6NX8XRShmnXh09eM
N7u/4/sjoEY+/UolJiieKBHyYLraLngEGTe3OiWiySKYy0h4p6ERm1LYm3zt
8+vgd3eduGIDXXr+b5nDRmjqFXScLQZ4ngXBzXApntFIY2IT/MnVLdQq/toG
6gIE2IeI+byV2CmEnGzdIVZzSwSc1E35h+bGwJpApdgDQjX19e512OS1lMNm
u1G9OELLcNPo0+8sgRaSHv/rBdcgucT+DqIxrbcZCuFUBAT04ja3M2fhD+NQ
GCjGP2+gTh9Ng8BsJn6cBcUtf04gQhfONeJ2ZhLoND/VOTmFWOSukamUvS0I
0fQidkyLEN+h9BaZFBuZJjxjQdvl/u0j0aPaXOyO0hOsDq+ZnNha6EHlYUoa
s6SzVxt5R9uHJ+dlHog2jBTZrnO/JunVXymqTIIS2NPkURCDAsJMZJ+z+vPa
K1JZTzdFYn2M8sAFM9sbOUMhvPc1AEr/9Z5JPRxoDFdYK2oWCmdznPK7UMuY
BH7XhF81bBtdl2RYnnCvGimop8PP2zfEFP9rz340RHpPNfGox+OTHSgtFwid
gOqKip0OMPMhM9JIVpiWIh5ze0JWjY4zND+oSd/qRXQWeR8RsMjdIdCkX0KB
AKBwbsM34rRxtYOaVikCLT/kFsV3BQvFPCqnKz5RprzcLnn7MQkG3+5cAR8q
lP0A/qNyy8n6Vh4C8zMeTC/v1DqOiNy4O099hfaRUNyRiy5dOO6dlp9F3Kv/
a0BjDq3o9wmORcFzIH5XletoqSISMqJ1d8jgIJRK0IhIeyhTBP/mo5Mg/4bm
5RxFWQ79DSQdgul7lnrFemzRMjVaz+5ZlFx9LfhfIyb0aL88lUI/H6ngZXAX
87R6kMk3W8+6bd/IcEe7yPZX0pnfkwxZgZm0OBPTY9w32Jr0UfXbsN2n4+QZ
HlwU/x96iiIZXA1z0azjQwnk1nqtUcat4aw3+se5T5eEJDT/s43yYg+mhtkZ
T3T2iGUeUJFPgap0IHN6qRGuiZUttjkl1hLkhALzCbihad4try4O6Ul/q8Q/
lFUyDymKR0o+PdFl1EzugeJHaDDTpUjhUio3H76Ukrvkb8VCYraIlgbC9J+G
tiq5LuYnoPW4csu7IylOaim6ZamcsLVih9CdfE7VLfSSf6mDOfr2zyvr8g2n
JmjICLUryN4/0K+c/L+VUrmdwuzJGGHZoYnfMC+sE78eH1oGSalsrJChweAE
dzeYZNBUTEM+Hx2s7rw7vdyX07KoCfNOFpniip4t8mLckiTJSk4lI/zHpMmV
km0fpztQTniqSdGlyu5cUaGHF6yrh//U/h5udar2NCa3hxnBcV63Vu1j3bLj
ymhmDOHO31+ComqlTVgalXpau8NvG7RbwjKOrRQIs+pZAERh7dvZa+uHOi0o
lYRJwXUv46/uCI0yTaKPHgjwZkwG2YaESJuFyOO3vZEkLVU6KSNYW/0XDXp3
Bno7jjbOrYOTOaLxXIlhUGJ0hHm+DAVLo08F39HFk9xLYpq3OAMhpkKCN/CD
dF66jnw7IGYs8VsXi6wB32D416yBm2mb2Enzn62tmRWpb90bnb0bEeiKbhYv
TIv8o03s5zr807JrmkAaZCm2Y4L4swxLV9NO4cOHX7hCXnuFLMkNPhdKIItw
mVYbpwy5X2nV4oYJGaXrK9YnP1l3NFJSM5dV0iFkp5twX3Afy3Afjbj8ETYI
+sSGaZAfqF0cw7iWqsNyom8BHS5agJYJ1kZF8Zus8Ee9zi+rpcjMHwaVlMyP
lrMzBRLCT/L+2LF272z0VCebPU961zaruS8MlkaCMfALqL6qgJ1Af0m32ZtA
2Y38wlEKnmPpC0dD0cCCYEyd9h7wAnijTMBYTVvMukWf7Io2fv5INyQEIRSZ
lLt09kNQWxMaKMKT7Sx1iBKwxrOCLugBnnSqdStsbcOFxt0HJEnMlQ/3So9p
tZaOm9nUu+BdW+yUOhYTEzjGU1sndEtdTbsdwoS6wm5CYAUwZHzReLS+bEjl
SsUkLwi95kXwWv/hgUjuQ66TLNJvlfxafAS/SjkPdGlXWcGKUV4kFcLy90nM
x3c2/mgGIiX9XxTEDMx/S7pF55S4FYHt9BQiBJa4Y0zkRdCpmcaToY3HZLaj
zUzvRcCVhcH4kqSfvSluw16MjcuytIzlLd/Xv/PxALwXXqdvnP3XY54NrM8v
2zSmdtjLmN+Z/H/UWNTgvV+VxkYqLmpZeI4GMnGDo+AdDYa3oemn0ueLuKCC
iYmF2OxQZp8L2yBttN9LXa4PlCMaG7fd8llBLxnpc2SMlf1bP9l/ma2sdaab
zORTky1rj4dtY69EfZkz8pfXLaLgXnXM9Yq0r7w18wRCd+SK6ua734lTzAlv
VXErOJGVmseNXqQjLC+qZC3lHn1q5OKH9AOMW6TZ9iHFKBwe2QcnNozCL/x+
5UOjPjLYwjS9tv/jZPn2cyibvdBEGFxgoid8X0dL2DaL05uUpfNR/PTjrTnJ
MAyD3n0SAZAgqogTk1DJ6O9qpR8XJwJZHVeXAgjVknP/+72GMTNUFn4zgaRG
MBwdpTcb+eiHdr2duMEK9vrkjrDdabmsn6B89ttvKOwhTZoCMEyIrm5DHet8
oIbM0FnKdRqnkLrmwc+ZT/Q5vaArz7Z1Qh/CCX3C9PJ5+T/xE2nmkniD7apt
SxaiXTvL9+fHNXwGSG1ONanu8adNgMvK0cKno0U8PfU3FcSkj2rfAEIm9naQ
BF7EzVppvR6Txmf3R59hAIvBg1Emqw6zsCWGxnwbAJEfqvmA7xzVN7gwgCoB
3zr9d3teiOh6oQZAAEJJuN0f9u0ya43JaA8jFCWX4zjeYvT6XF3QI6EQuvI6
zii0yhJqGnCNAadcz642UtkLaWF64V9049r8SKi8fdGtwfR4UCtHxEhjA1sd
Y5klvHuEp7zUOvqIWUEmVVM3h25XH2tJKyQVmysfPpqC9erxHh+ADAAo0hda
mlW6iHhUxHI653GVDpP7mgJcUxe1WMFWfylVjfalnQVVHff2yAdKLtnQMjkP
GxxmpXFD/HnSphhc2dleHzF+5UF/2r2inIlZrmIUts9eZWHoZfpUq8ziL54R
TeFJMQMs5vd01XSOnkn4gFzIpXaGkP/6BIYPLegopRFFi7frWtjF57vl+Fmp
+V+mxwn/WQ1i9/k0Ok0pfaOWpPVyDPDp8x71d9XK6ga88qlMawwV8l20vkmm
Tlcma9sHAQiU8+/j0TCQ0lggGbrR78Vo47TpqKRu63w4UAja5T9L2u4B57HB
VZcLylmKPtfzwlBvODAzoKRqbUoeAdcHyWWUXxArTCO2El8zld2yGsjth68L
HrLi+yg/zRJuloxkvoAiPFdbjA5U/x0gUr7HW+jlPAygSalqWAXVrew+rMp8
XOa5q6DvCVZ5vEctkvlXyXpCtWAD6v0VBNM5ef8xC3AOPUHnS4/+uoP4IGLK
g4fTqQrULYKIcXNKX++lraSnNo17U+l5L4oS2R4De2wTnx64pTFkWxhr3CNp
EcaFcUePudTNaZbob9K4y2e1cY50wZCcts+CG8Y6Tp2cxAlaPw6tberRP8pO
kOf9MRubUsnQSe0UrcVz200zQWo00b1JGMabnsAkTQPZXetB6wyYRy9bSsmA
hUC75fzEbYHqBHeHlDPDStG4J28k6urqkMFWv6/sxhsEI3uE8nmAvgDvbaJQ
jWwIS/WDkWayCqHrGn7Xx8MOP29uGPYGhnPt2xmiqX81PLPXSjWf4TiNwPZf
X1TypkpPp4kq5HjeNUa5QlicfpZMp06/Vi1VvYcyLqRV1pKw2RvC+VtRnqch
o+s5NZsCYlWi58PmZsFVB/SEnyWFvYWXs/tamsjWxOIefB1TWOgGbfiwiccc
tGPy2JTE5UyIn/wlpvV7yL/sYZqW6SThV7Jy2G8y3Tm1lZg/Cx7PfVJlBuzf
DiA1w6HZx0byckIZfQ+usg7AJPQ+vzEZ2dq7JyLtJOmn6LiHqbDg93IvdxfN
QNFrnyVpdkEKh2nDtc1bWHvp49ldRjY/joKojceglkWpLfJsBZYYuQV9tUtV
6Ij3HRvctMBaw88hNXxxa4Vpyw/T4zOK+wWtZOteyoDIwy7ZcKgbadM5qRQm
pVjZAnQH1hHx883TosQ0wcAaxTWhI9nQxbz8+PPvXPJVt7zQVizsMJm2dMC9
JTgOvg39nLeSAnWSEfISXYX/5Bv4cvt2qAALvhfL0mOZ5x6xmvElHbc2zqbw
B9Gu0bYgrDJDmxJLzXiiW4SqEqYYByxMFD5qw895ylHr4d6bZuN9fhrzFOl8
RzT+kE7JyM5cyYKEv2O4avorS/Esx7Y4IGs1sjxpwr6U/zdw7bvpcS6BQmMj
5swg6jnzr/Jr/cd6CMX/4t0mlbc/8ZAhCLaD7DmZBjZT8Gra16Wq99JXlSBv
dV4n5A6l3sMRf6VBtc7KjL0c89ZY7XfEAvDxw8gZyt7nOU+CS0UjkgxAOEue
vV8rGe8FYxSZOaRJq4Ve5XWePRQ6xOH5e/QEKWnQBhD2wV9WxqeUJZNzOJK4
eMnJLlu4FI6vwNC/NhF9aq4KgBzzgcuK1dIMtb5xFxPvJmO6pmj2hKEhGoOC
dvr0z/NWNcWGR6dGIHDP1dodg5nFI2udvs2XqazsEtIqyfPU0PGxof5IzpDH
Em7BblVXHQuHCBaHCadIESRi4HKN95V4vLhzyL1mhE5lRTu2Xj2HyccVEQuF
TZMUcmYsTdrTpaj6K+1SUzA0vsHLkFl0Fy0lY34GH/kYMVENUE+CLKk9G44F
fsh6xTIXtR88TmRcwWvI965j3uFHjdI503k3hVBE0lEcPFyIqcw2o/+7y6+j
m4Zpjun5LX4Z3a5E3yeSxraVkNocUWvCPGBBVjo2a+0gLbQqVNHFgSXvlgJc
6bZkZ2U7+nFj7h3WsYzNt8PG7P2oI5pKgp2KDMss0yxb1Lr2AIAIjFeVvsc9
qyIsBtZgXKVLEmqa/T1FNP/pPsgsyix4IARtTU0TUDtAwbTTxhXXefLXkvsP
OmFEslBqn30nDWU3X9woeqryZkXF3sc9DVyHfU46UBnRIuLGxpRc/LtbgRfV
6Sn4wATnG9doK2dRk5ecgjWDiz7Grl7ifh07JxglT/FlgO/Q6zicUbP9+euO
rZHEoPj+3I7EwK3EgQpAJIjPp2iyOk0z31JOvPZjsfsay25N5JSf1rPJ2Y2z
ppvxn2VI/iO6hmcTzYrYgLfom4HLi2RYDKff53+cZ5ZKtZYcJ02HydHDUvfl
Bcn6Hh/1ushd13GVagDYXqN+HytmBhDS/59jamEUT9CWR9DO0Eiv3O/8AhVw
MCA1pJyk1F5EFVKs1DZBE1SxbO23RCjpLdL9yqWV8hC62TdntNiECNXgtcKX
4YFKgucPIsG3cFJxkrmeFbLklTusnvX80GuG855XcawNmYMe/q3+K1BbXEwJ
lyMS16CCtNQ+bYjrPRKghcvM97kK//loTV0UuEYz4iiAhNe30qe2CBatT6t9
P2gRyD189bT7MhwuA8zYT3ovDGOkXiKze4SqFqPZFFqocTtWro4nKsB7qNXM
kkIgRYxlNn4RjTmKYjdQ4MtJpiGALBozMISBwYhcNi0FMt50AiUvGahNDuMm
+QkSe0sBENYaGT7kk7uy9aNBNla67Thq66h4cAnyljrBuH/hhajW9MJGVUQs
lDiZNjy8YmsvB030XB2gn/BdMceg94Af/CXtaj8WThQq+O11nA8FHl/U6ByS
Pz3ZM6dt2IFsFypXLyl9mTiTGSGMVUMRkqtuiolB0fHGtrjQ7JrhxcLknYkY
xFJ4Ii97rO5w4FnfuvgGrIGpdQcpFJ+F9OjynLNQarvZ/UvtkY0/kbN+G3lM
K8QMQvtR8/3W8FsthLUZAaLRaCnKTdo3IC8rNbyxkFmmD3YSoq68UHvbOgmJ
jwMfPgQF5ErCMyRXuFTVU5Di5SnCGbf1ZKys1BTsUzMzyf1zqZ2qRsC9k17o
vrQE5QlXTuBcwk43aFWAKn1BciZYYEoAJOwGtcAGUcruDuVYfuSBvQJWyMII
zSGktrzzCvrBXqhsGUY4m7a4S1xoi/BBU40Hw8pBEmt2x9gmD6y7ea0B83Na
i90n5ojCh3i3rFBLJHTRlcpD8+lGAOIrx+Cs+WSYiu5jjIGf0qDISgDIrNWX
0QR34+7NybSbuqpqaT5jU3ZevIEH19aaSit+sBBs+7P/idgsU7xn4WWiXjiD
oEnGkt1/SsEuZSu/Opl5hC+3yDo896aXD1+wsY8drfx1nQvyZd2qa3YYdbAC
Tl++KYPo1hyNWVvbuInAPnvs2hl1eX3J0/21j97VF9Bzh8TQTE8sNASGRoZl
mLxqxdGHXgu5kLtWnFemyCcHSQH14NgIBy9AYsBFCw2w8JZTq3zeBv/08MBS
NUoBEHx5GTxYc4sgpPPySMeBhVci3hMDKVdlpIx9K2VEZLBeXyz+2tDyylfc
WVShjmlGPzkpL4B8vFwWihDOA0P/rO4SQL5EZemLV+2LaPtEhmJr2ncBYEWc
rqfdk8h9I3G4MzieCbUecuE+Iw8JaDAfHiC8t3Gt29R696xascyYE5ARBCKa
S9qfkqVIDnplXh+RJjElcS16eU2DdeWc43QO0P9SMCD6NFK3BuaVS3v1nAKF
VCP7dmvP4Ty6Mw09M6WAY4X33AjSZAxbTDGjIXY4LxI2JjGqrsZHl39faaBE
wdDgEXxDJttJ4dYYQoQEAOveLns+QSeZd2gbESvoJKUsC1OgcWtY3DrxzTxm
20aHUGR9X7TLdv5Mm6shCOzP0S+47cQD4BGnEQnfe+3X9Oq37rNzHzdALk19
uanFqvq3sjptPzd2EjzRxxZgngiOxunkyJm65B/82L9++6WhJlnEtKLKq9W/
Ta0YhJaXM+ZMqQKmmKFC7ZxooirTYTgerK8D/Z5ivNk/4yd3F99E5AOqw67W
sEIH816gcA+G9DA40nNsleXsXH98eS1AIq2TfvVyb7lz86bAyZrdNAtvQ3rg
mvYYT/9+06nExHzq8KpUnHYNKnn7PVeGAAbBG+CpmFyD4JUraSvBRJmzhAYT
mkhu05Jht49PCOrZumirTdMofUxw06MiuhRYHKKqHCn6SEJez0/AyDfRzjRm
Av0hbfV5Iq9HjHyofaOxi9J5Rw/8Fp+YKw8HTTtOGjheLYClOOLQvTV5WkWG
3ZKVQQMA2/d78iWQgkN2/N3gC1mYVjoZAdLlp9P9oUI0jLv88+cv2+QTNNBx
FyAv6swuhC/DfZ3OP524hOofrp4nGuTy/INpooRHzv7iybCKFf2FRsPWAU8T
5j/T5N1vTgDsHzFqMgAeT/CLdIZ+T/XIvOE+Thp5ePJbA6YpJp+SwIocpgaM
9dlFRFholncv4Mb44NJEyO5DFOMXgd4pSYnkz2H+113PmILh8+VqS+UmP8hh
/CMlrG+/q7+XSSFrxwqnckQg39hQ6UUSB+oy+dCgB/a0McoD8J5pf01JgsV6
o4dw8o/QzaiVLBZycCoM1GCUdzvsIwQK1ROIcc/LCYct/NjhrE1mP2S1ew4d
1LsYXK7oJ02pCE+4Xs7TJ49OH9f8nMgSWGeE5b/8PRguZKzoSonsB0LVlAzq
KwE8cbZZy5soW6Io/YJ4676ZAS+qbFxDv6JwSHp9c/WvgN/fjvfWIXFSXGRZ
W3TmgObfr8OPiVQQIxSXBw85SXKcZx4fbVqf53rv7b19BJYyZmvjEOxyGKED
Jng+wealUIAcmfPJz/qGHzHZDDbE3GfU5+cyn49F7a6H/eWoDg9n4eJSw6Am
AjG2kr2F/wOsWJHUc5CBa9EVjVRZOitRq7rleWT7Y87QUeo4VVrRlaPT/HQi
q/P1dzMosIv0zLr2gpesoADgP4IYRF6O8+svDiY2qTdxNIRVuDK3NTLJ8Dy4
iVZtD7f0iIzT4k3qrEvP787pAPRosDV5IYHt1pNLY3H0y8mscqUYBmLDWT/U
ASdSUO5osCutxPiwOP+qN6YjsIKXaFpaJmEp87liW1n7/LG6gYyd1ZqxV8Ct
cYg1ZtaFsZ9P+8E83Ac5qGbDFAB0LGXIBvDYa24LVSQSuRaycNp7EZaTKo6j
qoBnb6Ey7xNNM8ETqPIlZBZJ/xJF21IfD8EWKckyEU3B4S4fGtrwjCJ+VOzr
6Qdi+EnaG8RHVDT4ijdBmkyQjRokx8gpZT+M/blW3MgHeu1jASG2S9ti11Cp
GsE+OcGizv2/tXZP6gJag2K/WqP/7UL1FobCUL7DYvvD6ZmLcBouj2myj0oT
F7BlCw+88tvnjuFUSIJc5HGgtvORkL1D4c8kfiFZyuqqf9JXXHqRj5wJH+KZ
rwlkE5+slY2Uu1g3QI0j5SCN1/PLV37jZGo8AfzMN0e05xpDVYG9eLu3KRoV
+8mmoQstFnpIAhvWYdeAyuMv51voSr4TmaYIvRd1fy+zOO4HNcdkAh5efiOS
4aBPwIr9MvtCXGSeLTKObexe9EEa6omILTw//V0980lVo3mxr4Yzcwu8Vv9U
d8AB3MtaUldisM8uvo9GHJoAocziBRYPlNTIgAbyYntV1N5pGQuCI1N7XQlc
zRFECi5cC/0e1sGYbbnMy673k1b1BJI36prv/kHVfcu+KEQatYIxZ1qqJmdF
LprFg96cEC/lhghgyPMPRUhjqudoj6is8XOqsv4hfsoS8slQERU/ohyvrn47
c8lB3QcGVW9h34Sy3QagclVQydNFBCfIVf9zV0jkxSC5YzNiwz6Tp0t05Ep7
FYiN7XsI+7dC2EH7DsUcpp3x/NP6UEyE+qoS8XZSrYa1+/bVLmKrUX+agory
d5Gm+qhqO2kNGM1itEDkn47fWOi9H1VAoaiAk7h3X5/o/yCsuzHYTcP7U2wr
bzQGUBW4LlliSeXx59jfaTM/+a9I5eNMJIV7cJakv2I6ZMjM9OkY3Cdyn8zE
t9nUXFu9EQ2FWv9DGkgsv4ulb36G+Mw+Nc+WNw3lmTdTkviZcAVK92AMy3O+
cGXDh0Vlby6g4XZXkL5EqN6MtCzF/QclSNMG00cJE1zgD/OGJuupYloUAqFG
WXp+NyD/lfGaEiF/DwatUhL68LPBVJuOxDASFuRap0IOsaRATXnLxn4mdO5J
NW4/g5cKxX2+edyq1B6NgzhG6iCLxRDdoM+wAvTV5RNocwPI7EemVfopq/0U
Bu9PkuWEaXVW1v0d8KVDgK2fvib3CbM50UmlvH/ofZh7tgyHpx31SgmLHg/W
Y4jJHkHdiCWYIho6MwPAzo/rw7U6imOAJHtwhm6B/61wZMbaSAAY/C4yPpe7
Q/zdb37Yhabh8AjLmfV443K3rjvJGyZRQhpqNBCwEwln094Xq10Iax+0K4Wt
Nc1+kiQdRHIWcZDNcDqj6gcp0xYbWZgjOHdpGEbXNQslYNNefS1vWYWoZAMo
8m2a+Qhlh85QbnkYaBhpqqUs37L/Ab9wgabDZHHNObYwfFeeDqm7qzGNuu48
DsiIA+j1of2lazdQLsfReeVyH80EPIdbzny2kU2JM4ZTQz/jhDpvleIsiy2u
cKhtkGUlTShpcdZjYK81CPxCKq49ENeiNWuqHhlK1LiIr685JeFVJ+FJ8v1E
VSY/c7v5G2m9wbBRqgKYE3zV0kLu0Kig4ISeKcKwo1D9+QJV2k1W062WJIsA
zmoI9eG0221GJwPvq+STRMukMYrkv/Of0Z8hm4UEpBg5tNoJJ+ybUWWLrElQ
/aNZA4nM/65xnyP56OhwiKXpXVR+lmMvHgm5Ta/7PkHKDTryfZsjlGvLlGtN
C7rbhMRQskJzqnwbCj3IOgHKdgRliHDJu4Hq3H0PHKizy3kg1f9ynXc9Big1
Z3a87mBH314LomSG2nD9I2kt1uefGTsh8k8dPe7qw2ud86SMIuv70lfol6K0
IMFyIj3Orj9cII/5OQQAFNQOcuc3MU9gSIiuc8h2yq4ggXDuom6OGzvYT5W0
A9EiKVs/uUJIJoF9HPJ16Zg14UYzdiV6qMIBZpHJpu2q4hxWkesmV4B0tGSn
JzUSclzFyYbIVo2XgWVlCqjfhhp4EgVi/Ud1kcBz7dS7b+qfiE74FqD2Qh8/
qoC9+HKqD7igfFg2/jaDUsmZ2+9bBjUC70gB4OO1T5nSS8fadTFFwfYjx1IZ
M+wXJ9Q5PGy6Y/ZPvCM9ldNAjDenj1lfb85e2fhypfbpEE3r5KMj+sGCYrY7
dZF5vy6GnVXLciliuQkCRGgTP94MUuS+FnVpx7OzuRnpzV43q56Xa1DACx0X
HRYsCJvgtnAD5bd4PAo9XNwfTRIzEzlmo0c6V9pKrh6l5oNT/01Cz11TJl5G
0UkppFy3a2OMHQJ4dkCJLJ0JwyyUqJ/NofD1NxNwmMtghCjgMYRwSII2qGhZ
zjXqwzJ0VKvRo4p0ltiUHrWRMsILJfkeo9mTCQ0aGeiirgFhJmDCd7KaF6xD
n9Rm6dRLpdifrjia7+jJzyEExbVhDBBwS3GLfQpO+d1d9SwvcFSUYt0Eq+Oo
1fzcSdzzwgWSRECS1Tg/0hdCXjw+4VbKZW4DXEp8ngymuTqfDXAROcyrqRj2
e4AbPrm0CpPeDX7BUH23QPmT4Yp/YSjO5Ki5Q7BCdDhc5evzP/1e5XIlvu0a
mNv9PSRZLAPBygfXOPpsjodpftgoT15sWhMZ24qP7S29k/4c7eDu79mrL+UO
W0Qo0sS8lAxj4S6lXQURfbffA2Fp7hOXEUFxjKIJebyZZKTHYs+5sN+0gR5f
H0fhpo5VlEgH4/lSuP6Fwl3uooVOo+fHGMkVwLEh1ttjQVPNXkEP44U4uZG0
FO4oW3uV5sS2yekFXazVQpmisuVwWKtnhdcB1EYtVSX/AF8eof4QUJo6v3ci
NEC+H0WEk00FjSmfdAMQfnbpmDJoXX7Ca9wnckESAx48yttJnjrSLGoU0rXz
MGQDn7MFObJzNPQkpU5nAMg8JGLdlxA1WBLgUA6ZWDafaSnI3UJFpdZQWq67
ZL28DZBi9y/H96/RKhkzn4c+MLYsLG7Q+Lk7PgKfsLFxf/LnZNNc11J+C1r4
H0iM+8KupeuNtcmL0hpmmclBSdGRFUqBzwEKBUr+8Qc2aUSvs+NUE7fS9fq0
+TGCAZX4vskbJPPHVL7C4Eo/TWgsC8+e+EZwduzFEhdz7glbx/o2ZENQ+zPP
Ey0CofqdHxOX+Ar7A42ckrkedh/WhJU2yMUcXCRKxZU4pbOVmqnv00fKyZTP
gMGbzCt315KlhL8eIxjrd5tF4gFFaH2ADrnHWlq5UWBG/TktqRm7AOebda73
kJVX00A691NgzY+yWQVBksmLWso2OOy//ExUxHQcTG9r1QhBk7hDREQNIyWL
a3TIiNEVMyQH2Sp+NZ37LjAoH6y9l6HqxhHtNM0ny8EST3Lic6ju4z1L/aVq
20u+1lkPDUrzFpI9ub1RtMJ7JttOPybrzv/1V1KYA5SndNF0cOBn17U/FGEA
CJvH0o4Ngw2deE02ncwY5IhrsxJzP8MBYWhCU0rHqClYTqGLgCEmTjo3iYFI
Rl0bQ4OKn9er23Y6WMVLQaU7182UmDoj45HoSm0psuzrbGmV7y/69RmET0HT
WXqeoSZuw8b+ja6HggSf5VBfnpRrnW3tcIuLxlof5k8curuy2+nF0hRKodIS
PbMweUHsx4a+Udfdp7bhuf/Z/EsGsDwEthez37xFnE0pv78C+Q+8SP3Cq7//
M/ucgd++uOqvWsziy83knosM22eIoI1qwLC/fRktVWmuci/zxqPhXQ20vML3
amkTh4o/1EgcXqZK8UL07M1IzM2AVfvp4dVsx5YXSJWbDlSRj8yeG4XnkbGH
3IaUohUrmXRxNi/dQR6KdN1SJjUZr+Nfnkk7sKRqHrNx7BfKaBrC6huNj/oE
No5kNZiXq83QfobVlz6bpTWuom3ax/rGgLz07k3TDrux9vOklSkbPORMxx0K
3G0R9ir2yEmz3uP84DkAIgjwL04VvBk4cwoAvuJ2yDXfI83W/vcy4NzIoKCE
t4DMV2PzSHn49f7ftfqc1zHstRgqAEQVwQTlEKn0B6YlT/5rKfcAlRWyEQjw
FeOlV4dml8wzKBIezPtOqHPw4ru3n9wuP+xa+EWooP3cMs2m2FTu4rtGOJGc
IPqNVntPAog7SmTZdfT5e3NlGHCggLG19pE3YSsWKD+0/1sPPFaP9lZmEmCf
R1KYZMYxocaCZ/dq2PQDclQPE3GYSu3XBR1PHoM1YQxzbPc2TxPJ+Ai31TlC
ATKnBB69Ycy3GRCLSIqIrzb/RU0cEmDuwMJcEnzhsrWcnZ/gyjqUTrkEupc6
KVWQstl5gu5r4mJY+B5oFZV/uXWgJzgmqegToErL70Ybhy+a3iGJmmN5lsl3
RmMMIE9j5/EN//jHPrfENJBedBbjmdIr0u9Y9Wow/46gqyo0Ki+9h7skoInc
EGSq/hADwKbLNeeNQZJXRf10ghHcspsbNtpcBIJLhoqXKQxqHMIn3mBKYbiL
Hh7+KU4fs0EHuRWTneUtjQNwf2k5ar3pz1B7K/dp82IgjKWjXGmTYZeMwoa+
ZWuA3A+MLQA6xlmqVz30hS2EN1qy9FlaUeC8RFsOBem0+dJJoNQlJf0JaTBl
iZsbZrvDshu0ysSJ6pM8bs7Ti8r7mLqW/N81ovo0Uz157jTIOEHVNeXvLqUl
1Ih2NNlHgEQxbo6rKmM2aBKBU47GOACaAHhkkSBxV+XkYBJh+6sJzac+XyRT
E2xb/2ftF/ZQSE9viAy4fElxU4taWcxNpVnfXzHk2LaLuywyFQIeH+HhVCZm
gId1+HS8mJ202e34T95qpVh6HTaLFFK3Psec96FMPU6J6UYm3pLawn3qHHGb
wVest3YcUBJNIVWd8YzZoFgaFfTcBtJ1IRolbP+EONNW9DUspPhMaVP1XyeO
Ku0PgEvOWLetSrTfEOZfZx5r5yP5AR1WcV+8clBdx6YHA0Teup1nnoNHMmdP
XLYwxfO6RI8dJ7OkfhWkZHIgOciXb993I7MAUJ3i4+k17ijqtCwrrQHh26ih
iZosH/IdVUWZ84fpbI5ZiT7+3o6PiSEG2HfbkJQT7TDb5o3OxaiSp2QZu7Ib
axpluM3mZB4k/x2x4Oh61bXhi4g5lHVcEEtq7o+ERwjvMO5wG6n+PIXLYlzi
s8KCQFmtj4KfGPjLQnTrIsShmR+I+rjkXcB02Cj5+xDJcfWmVK6tPjOUgueo
ZRsLTpvM2svF4D+ssTZbzMI5+Hzq/EcWJitlf6mQD7dYMvC2yaFvt9oTeYIt
tETPXF03Zmrtshw2olEEAzqXPm64hwOaFnWHFusA0gJhlUFj1fF7CQ3pLhEv
CytSWc1VnFqlAHc/QW0cS6HS8av8o0/6J98iStq2A9zZwXbtyKpYPLQSUkE4
akWRVwfDGwkJGCPIDydkLISc9eLSU5lmvUUt+yxhSRWld2YDAlglkmLS//X9
LHGQg2cWG24L57aeViUhRiU9p+1DmcDwdEJauYgCZSQ3eLsK6p1jtHaRiPVv
429ZVmyJyx/dg64Kp05yHmVp1Z7xff/H5LaaaPrJGhV5eAyprq7/KSMMIBnI
Ztvjn3AxGDhWMT6jz7RQvCkL52IxnS9DUfKqUADztw4UOTcRFIU/NpIn/txF
BWYZx0SNyJQLAxxEpyRXNKdJot/nn7Mz9wdwt4GjaoUVmC1MN8++EAkhAG1Z
f1wJpdR3g8KmuO8Zk0dZFU4SZiZCSN8rjxt/X9mJryZM8jsyzRemSK2kdjWq
U8PGpfQKTk2ojqIKEsP2wH3u3J5ZOceMKpuxk9yBQh+kORggtydBbWnywQaX
QAs5VhwDZl8zxLDPRQjuw4aFQwztzS4/d6QrpXEVmOUq3UtuHJWp6pMRbAC9
+3zGqwK+Dv6lxA2eNCJJhS3pP81WGohkbcLUv6pqcHw/XGxsC4H2LhTw828q
0lWoewosQcyT9EH8uUtInHJMikzgo8tzQTPrhdXJeM5tXVckVLuEMSrFGTU2
4bi/ErazQzjfvfnD9T4szElSbQXrLdIevy7slPqmKu8x2hY6KRKScLqy83tu
7i4jZkI4Zqp8/gJzY592QspwT8DMa0vW6qosVtzx5aGTWhgs+vqM9mRcWp7F
/eIvr7/QQEJ0bGn5hiXUZbMFgwDf1NXGSdEGZTMBscynUxfPk9fcwOP08Ojg
1fVewetnne1aJ3JmRuGFXBZUg4KWDcRATSM8gGRrGRXgwzqiZWv0sFFm0roV
e7MkyBUp0JF/4bWR16vtQnxLunrWTah50Kh/GOZlFYwVrkE+z0qyh+KFgKCE
+wUhKsq8k5+EAb+2KlLmY8seFivISlrInJ8opP2ONS0IkMxvjf1wOG+2qFb8
Mn3rpGLmnIxtjiQECNlCYCFXrxoCZSgua3Vm0D70rxTPYuL1wyQji6+OsIC8
fUWZcCoukWPAu02J/WCltHrTt5VSvxMGcMrTc0IfhkTp7mdQjP+WlaxXxfdB
+zkZam0kjRwzajJqQROlDHYXeUYDhIPgDjARM3vhUb6aiQcXWkbilL5+akie
01GPIKzCrrrP0GYDeeKmMa5coYxO6je2+M1HCGeaeEceeMhx7MFVyxJz1wrC
yIts7uIgv/RRzhE9jDFGnQBG+7YZcCuG/WOUqix0/8m9M7cAR01w3+0U9lHU
N3qb9a1oXp5/FQF4e9BMEUGpdcMY/7HCRH3FIdQrGwNiWIZ5sl58VqgJGbO6
6+pfNnPKDeGJqoms/WC/CeD9AV12gDS5oo/x3y2g8TUYXFLJnfwzsp9pbGjK
wvTkMMuySfLN5u+fFz+cXvL8bQbe55N5BayblP1OxpjLDpmPXZaJH/JSgNmk
//Afknc4q9LLPClCEnMjc0Jvb38lMwJJgGPcGG7mooBeg78C3TiylvqaNxeO
ZXlFz9hp0kenB15x53kCgXtt/dgJc7VlscQLgrMZU7pzduFNcmn6udjKmty/
FTpSdWIA3fBsr5v7Ac49S+ZW/crDCaIkuI5MKuOsRUOWRP27WcsXRIG3qXFP
AwjCdcccrabe9otMi5sQrbP5kxULKkFgPSz/2nWVSGAMp21dBP+17ZY1jcp1
p2GiQSfamXMW+9GqHZxho920GLRpeLQSuht2AxHlDOVWIsF/b21FQCvn6xfq
0cnGg03LMYsNn2kgoEhZ2SKxXtgeqfMytz0ThYmV5AZbvNJTn4+qNaHoHiR5
eHp+IzbMwR6rUsV+KiJb6X4GbPqPewclvMHy6iLcTKDQVcj2P+u1OZbNpKNP
MIRfU8Yvd893GWgbYD0CoOnum52gjTaOeeTKzWUV5IQDrayVCvAIGyESNram
QpXA8boixYXmP4Akt2Oo/3hI2LZzCa65KRAQ9KbCxQeje6BJvzWPTqO57kNR
1tUmliJgXXwXIXVwHq+ew6wjaKMwknQGpFFHL1v7L8nIaivz5qfQaDh6AFvY
rmdjvS6VCCKPCMMZfQ6xj+IYAdj6wMjdeRep1ZFAJswq61AZgwjf0WLLowHm
t9cEDK0c7vuOrfbNv5/Ez8YLg3KsreRtjWqJCq/gyZV+5Og1pqGgyQNr8Von
k/iOQJJ/j8BrnnSgbCwPnjsqzhRLmt2UXCCipxNGR6AukTZtLxlK8bb+cKqh
JRcSqE0y/IrHlOg8hUn3jGHJEKLaVzSn7zqj17YUOMcZdyjVj0fGVIJ3LVL9
WapE0obqL4w6Qh7ARYhmbXMh1EaneGt91wpLRPwFoBMNyZwwIZvaQSkGxbIi
gICKMUt1UqXdnWo+uXfg1LmKkmmS0HOod3845y+AuW8YUFYf1eQZTuCEkrli
ukj6gUh4qyCQMSkbfXBH92oTXbBdCHfkEjIdT8AOTfkRhy8I3Ml6H0+7jAdL
f6K5hwoJ/nzwJTWVgOt1uY/UIkDM4ktn6XFxkrB4P7yebNHWda8ei4wjLA1d
PEBaFxNLhi8ZvyyL08ORzGrQn2up/vryaPkwdJ8HYo8Wn0bv/jJMFRevCTmN
vpSwzCwzkl3z0Dlg05X9fsmr2A+SThTvPrp/gf+QZe6yBqiIWulhVdFDMQuP
G5tyJysUE7dw+aVl7JXy54eSB2UyRgwNRDs4IZ/PjLzlrNHBIEZ4lea8D/CV
0hFkuynJx6AtUDhCZJg0kIImdsgQ05/PLzWmk5J7M9CiB0UO2QQOPRjuAYNu
GlJNvqg2TXCfdviFLKbSIA5faiKCqOzQU50nSpLxOA6vobpTNLT7jPSoPmsV
jnb4PDOlkxST9flpj9NKYJjgPw3S7IOfKEMZYPdYTeyYo0YDGImeA/iCghnK
LgonD8ADpMeUgcJtunIzMpMDf35pie81zhzAQpbJuTMJ/seoAb4pTDZKgpRD
q0gb+SHV52/2oDEt83mckTyRJoqkA2gHnTgaiItlGvvHFfPkUe87AeJlB76y
CYtzjoJRy8RXVYa/dhvQzh8OtorjSISFJfdc5LGzMkgn3ehi7zx9VP35zL8D
Ap56h1uIqr+xSOrfgkw2I7jJW3cFj1RFTqXa4S5G3irhtyduyF26tEoKHyTt
GDbGfvD8ynVsk8hr0/oWGc16DEiY4Yy6XWxO0+b8ZnI3JLaRxFtaps0RIYut
GZh1d6xXZkCrqVzaYfv5n4ePaEgH3YSbT7ancoMkKC2NYKlFSfykH6TMz5EX
ZIDh8FhqZrVVIlV4h5JkRWkfUpBy83U/NyFEOnOHdjKvt4WskLQvGiIxJnNT
3/hzlVIUqaon2lrdHep4VK93EzKMoJIZn6plZ6I6pzsUL/l4grwEfaf8y+Ls
9+qzNvPFOjYzkQZYgxMIkPafWGzLD1qhje4hNDtwApTqQSBbRmkeUEOmqyMV
VwLbvpUNN8GeCNT/oMRaQWsH70wpRw343bfw8YSGjCkmcc5hMhfPqu/uFQTW
PyysGmAbbYyK8IUQJH8Bwt3hR0G/ojYdw1nbrFZFEXayh6aBrXHzMg6Vx1it
z7oJOb8Ui2HuPw4IzFqNI8M0TtqS8pdJDKKX8T8DaziksIlrILjwzLemzudI
29UevImRerke7BwZAQ1gKfv0z2/N/c0gDSznea0TNx4TvakdGo09/wfbsW3o
vnJ76HHDVUqFs2MGTEhSaz29q/4OPWlOWfLd/DqL+5nkpfGqIg3+JO6rRvSj
hVAwvWv/mCDQ86cXsEPRoRUoBzJPUehTDP2QPJGub1240API60d0Do7ft1JF
wWtYbo2mTwILeZ/23B2VXEhpVmlWT5xboqfxRpR53tS0fMeUcByYuZsIsuWM
JfHPlW1mTHuGP9dYyFSFekb7LSPkiK6wl4yACgFdr/hI4Ax7nzeGGfDZFbki
W/nJ3IQg+zGdJVFEl+Zb8J/zEgkqwg3CNs3lizO4nMC2BWU+FvNP/TNM2P1e
YQ3pLyU9CRcnICvvmSUlCwXKDDckj55zlDLvx3kuEvkfPXjRUghRoMwoofC8
TJBfgMJnYPRcVyc9Q/zYrF6CP4BYHtvBP6SxeACDJsW0XnLEj8PldsvdjFIV
R1hDxl8jWefOZ/vg2MX7Q8g2EEsOAz2WOIeen6/UkrcXOySV3XKE7jpclvNw
avuCEMAM+LjDfHWtXt2bdXEk1XffTYaUs6fGz3Zx6/n/ajEWUoStLDOEouMi
xTNx6ybBkN7ERTesP58c2c2phlc2etT/thj4VCrD27UCTEFuR3AeSokoIC4o
9Rjy2TzRcjILOkeyAT6RkULwv7CsCdaiaK8XTIv0PSSaeH4OrxawO3072wZ8
XAfxsUnOEimE4Wrri29LaXVpX7X+cQ72bat+A/54hgDFcoyA9I/LB4odqrPh
uAM3RfM7blhkRluQneeB8ZRGPFOrID1le5a+BSJ6ZOfPWIYsA6BjYqscfu15
5kNBhCC0+K58e1G43JdqPmhL4PPS8WkM8IM+zpMfS+hdGO70LZgpG/pgYZlo
kGnLmXI0iIXoRT3pw2uClOUsME0Cp2sjHMkyxalb4HBgn22x3QS3TPHsWt59
4PgbjNhfkIrgz3DQ56nD6fZyA/YQc810aaNCJ3lE5tjv/cdsPfz3sYz1D8Yn
NwPZGQAbHqv+pLYcL9U2guAbMJmeutmQ9EW/J57zptMw2pY1SH6FtekMdvpk
be/VgFfdG3oCLVXmMhFJMNuq1q0w8DVZWPeSYFrYvzfi+WbF/iHonfJ17mOi
/BFjtCCxl52YTg+IkZzURA7aQCi09ciDFCdMT0XeF50sZkjDIbpKG+WSwqLJ
bdsvygMPlO76ZtnCuUFuff7caKRHDz5VERXpiGb+GkmuWcPcYT1Yfy0LjAlK
POHyH3RaFoaNDIyMV8m5s9n/zvwVurfJbTQIK5MvkOts5rU/wV4Nd+vBypJ3
CpX86xrRvHgsPkNRIuSX4Eo1J5UK6sm2gG9oee5KathaC57fzWrDgVOFXuwK
pIR9iSHejkoL49OqE1Obig54VJRvUI5jie9YphoHAVXJecWHOoBKAQOo5wZg
8jBf8/z+BGBRMgsrbi+VSlh/iABBCWhjiyYLSTr5/HIVOtzR0Pv3hpzOv3oH
Jg7Yd0NrooADNfncVKYWCIq7SG6sHyhkZZe0lLEyJEtg74J047tlTmaGkSEU
0c/ztHYdTbq1lxso10KqK6H36gzjAV2j+KpFdWXDyU0oq/UGaQuY4iPsTDVH
H3SHlvdQCnD8DwzICi64ET5SYUZvpCeeL6dQJebmfJFn71xH68bQBwW2Jnun
bKjqDPMZHeXvTWbfcvIOGcrG1P+cFCOsjkS+uo4RmRf+SdpG1UdlWnH4yItJ
2q3WKOEJWUHRZ4caBS1NfLTMxPGa/MZ5IHUMvGo6dok1LcC29UyBtVYquGi6
evb/r7blPquMpq6ZLBBKTVVprYKCPY3UGfJd9sFh9UC3K8lSBj3MGDTxBP/u
xs/m6Yfp6CEicvHUd3Ob8tf5gTRiko8hj9QX2z7OkhmTGldxs148hWFSQgFt
O3m3ASLgWqeiLTOgkLe3S5fOVTDKA9t/sUTA5HxMc6y8ZWv76+VAQgoOMgVe
N0YN8cDTCd77JJg6LT2u3sqgGRgKm1q5abbeuq27DdLDYOxCbrdgmuI3mnZO
oevea8meyw6DFsBQnZMUq1K1ITcRh3aOAB16t8G0J43AoCdwLtCo6frVZdNW
yAgD+MSQtZRrBtUiFTO6NtzRVdD5GJo8qa4qeX3BtFm7FVj9Gc/Hp7Psnm4p
ssKulU5YQRtdCodzjivwUkmqeOfJv1ydocElS40xwVAZ8gpVOawRFA4Gmonu
0JV/V9ZzCH7/FOVRCNGqV7z4sF5gCM9J1JKSQghScsF89tcBNnWpgigr0Ooq
pXYitIfpvLwQTnX2XWwMPcxgcs0X66kWI78Yddg1IBzVfgI7r9PrFTZw2rjl
v7tqPvRTdd8MDLO++hjDv0RwkRWCb47mj+1YNcm+LqigsynXujCXkFF4xnsp
odaP/DZbMUdAPgHtt7PtX8SRaziP6l747Eo4f7DswLGUQjaVpLGtrcadYMRq
httK2GqrRPP5sJ7dv5rXe+48GpwkdK3G7tMPMM172Z6tqFNmNu4WY9Nwny8Z
OiALifJBYGrnZBIr8quZbaYQi5Y4MmcGwooHZEbueZRG1a/FrmdORLFVTHmz
knNudUnKU4cvpIWV31+63AnpbC0dXQj3XAMKPJqO3MeNcPlhP1dHdBaN7Wqi
ZoBfNvWrKfK9t6njIsQ/xhRllraOkc92DM5+QuXCzxoh1wFydb/wPrTGcswy
D8dXzCU/rgSsOEcJbjfptEaOqZhFN/T/LBENabcL5zqs8gec9V17KcUlaNLf
lHcb5sajdH3/MW9NQm0yVpMn9y9ZvyhItxx9yCWzT1jdqDS2R6mMPpUsNAs4
b6L/bb8onTqMP+81dqAuc1ugDGdQXhF0JyJKMG6JrxSwOB0+PqtSvtz7+lWw
D+6PvjykoYGVQhm6E94fCOlOuj2XL8XHXorJpxFYS7NTi13YVuxenkQtdT9U
XFyhTggZLGV7sOGnSjNO7/B/5mftJ37NZrHYxJBEOTESVN6THpcen8Bzy0PO
wv5cr7ufzQb/9CuaAO0/l1VVSx1SFqQmkTWk+K28bXF2UuV5Ke8iaHM9fAcV
G9dqQbkfs3aEXqMsvx65HS+32u2qjr8Q1TIuvZ2oLSop4c8kqv51LqcDZBWS
emSu3qF+DRAp7wF46ZeEr3Km3+1Gcewkz/DLmfP2Ftdw7AHqSYqa+BADuGUy
H8XJL7NNnuyrc87oOR5tY+NrEUqN9lUR0DP6rkDCbHH+WEdXH852dwjG1H3Z
WH98vgT/9AXowKE2bZ3cB0IpV0wqVcPJBg0az9kF+rsm/qEKoZdFw+5GmkNc
RrxHc5LkD2i2sY1J8SzIUEm01qRN6Y0Ke7DM5yJ3NhgmWIF++W+WX6ucq0Ka
QMhN1AIVMhDRw2ChhOHwwK8AtVTMTNN6QspyeGn3q9xbtNiKnliWVdXDzpzG
Hc4FjE5d91RkUDG0xIlh2KOoVjG1YYxT1VNXKCldlFWoDH7naiEGB8wiLs94
5ODsFyGqSkw30wvtWhw/X7UsMOVvzzO5Kb7TZ2dCJtLHvJrNA8nBZGvMTvZh
ukqK4LnRqj3LAxtOU4cGC+HT7fJ5MQNWJT55fMewhKiSTzJuTnBvVagrN10b
r/IOwRvVP5so4rXdffk2oNrbs/4X1i5k7F6SerKbCNaJBi6Mz2qCSot3Po22
GSHsT9MHlIjTa2asmouOgQy9nsTpyYlN49S+HuZ5/B91YaNkwQWz2wMFidKI
rghwNIOQ1epSCQv6TQLnv+UtgsqVgkSGWlWHB+LgTDWcDl3E5O9l8E4bVLkI
cGWaHw53f5fc6tiju3OKhI0DuAWOjdU1nRl8O9+NSoJfW5CH6kA6Frnv2EAk
p0cn8dDs5oZDmk5VT4NTfy/1sbz2aQdhg13UTvXXuf1r7Us7xQjNlcCLUcsv
h1BluSzGJtHjgOswLD0DpCCVniMTHUI8KS/mdHjMggn6mqXfGMV/XpT6RF0E
+J6z32/hP06vnu1YdwzktSnhvBmHcWJEVngTUfwvcc4PJRytYlZm1UbMozAw
ASvAy7GC2+UB1SgtrqNpaensbNS8gBubP2hoEgcrdjKntXPufjWoAuHGrTVH
z+McqJTvBR968kZmXS9ALq+BwXACv2gJAtDtb0q7D3DFnbsS3Yo9GKbLLAdT
pdrt9XQ131Za7QzzvbqMg1GUsoUCM72aHKLyD87azmeb3vpy+Z2A8u+ceI2u
EftChDwan8111ZeUfDlir8qU+BZOIjsWHFXSCZjxfXG2Zk7l81KBB9vTfArY
t7Qw11uvhZC+moyUWM99zXG93Ka6YLnqmzaMeZm3hvNrBjefaC22DL0vSUzA
wFk5dsyS7ITQ4kye3/En7KSrDmK5Vp3RWlpwIMKOBtUl/awYvxCTHGrJefm+
WW74osDtjmCoOwE7QU4l0hJg/GZv++8tPtRhF5Ov+QR1GyGawYi8fZe1uwJ+
YbhvirI6hlACXXkVwLmNgwLhLVm/nez56efkYl4izCCe2yQJ6nZ1SzaukDxc
Rr/61ey2boj5YZKdBdH05WrD7b6xiPRraLe/cIlBwq3c6Ro2qR9/nw422X4Z
E918HHYNE9sP87f2JaBW3fC4bY8fj4bFn0J+md/Xh5TfqumD4dwTKWwcEcRR
0I4MuEhwyXTlGCml9ZIDQmHb8CGVb2ae42mzlOjxLSLyk/UqkK3/+ZDT9ys3
BLnY+4snkiEZ1oQ4j9XL85ZSRnvi7mqWIhUS7XiCwi+he7K9mCz5InQEMwPA
UC97Bt2aJC/M9ESBhUP9QxO2jSrQa37jiuFoYlTsKERo1GodgPkRL2lE7Rpi
aGhBuLZ2QzVeYr/+09BxU5rAFqwildN0vTyNyh/cJ0WiQroZRenyWu5rTJue
7l+InikQmVVBWbChg4UnmQlGfDlDvHmGPc47F/1Xpw//OC7hNIheGsYzber5
C3SKuFMmg+rKDgClzNmxJioJQskVhNApQHJqPHDAqGEK+WRxOFxUD7SaAlRx
jbhK3vyzU8shiV9u/0ffRb8r8YOa6VH2AHm44HYZQQeCSL1r/whKmgRbaBuu
LdX4GZFhYJ+g9t3qwSbiJtwp/uC0aYXVY7v6nHvPsa6UKzr/+neZ8VJCizKV
3nHr9uUswovH/8aXq6HnorsfEnyvjbHUaDRfpW2S/z+FfMn1NHsv1Fip2oBi
k3yFBfgYiLFmyUXP7QZHIfycd5MUGt0eWGj90pxWVmXIqihRyVinrB+D81hd
IvXwFs0zt0Qu7M3UR8a4DihazdU63qHzitCpgPlRkt/WXl9YzAbGlEX8POTh
i1ogLPvBL3AQf4LqjwpxnJ7emZVfDu98boIgHF/p8Y5RtfzYG2Lu7MyFgUf4
mlj2EA8yOCa+PeUpVkWlD+EffgeiVBcVMUFrhSUCz3n3mydtDBCzI0r0TVz6
15anHnYqbbP2uboTTi34W0qXmFm0YTcMgFmkWOPaKIzXskDyIbvt4T/Vu8EK
dybkwYRrIYilPKG93a20bWvcLjKhpetBJhhjmLXPJLs/XlnPYoWf9zhmBKMS
+Qa1UyyDBr4a7zo9b/6RvzRMSNGKAU/lghSRUP5SZoYRPmNDGdE3W95Bizc7
0RfFeeMMX9M2Pa9mITax+KjfdK3pf+EeZbdWjQa8sidHUKUCom8bOsMhxxBV
YAl55JOsOyGTtnwfVeTFAOqS7ny99W9t1NSVaFxxjGb+HWF+AVRMZ2hDQR8H
AL+vRLyL2MUWpxspcbXJzWKxn8K3XSegcXCHgY6dzFhq/KJC4c0WQPY27x3x
n7g58RzdeAq2yuFRR8MyQe3+v9qvPhKh8zGTAe7CtrT6Zprdh8bjD1SwKSOV
xvoX5Is8EifRKtBwkUo/weY9pDh13aHrvAHaLrMIkQ8aOIQSy6rlckzx6Kpj
arAIBiKyOeOHmg09xAELuzD9ZsMqGmO3+YygS/Zf96iZUOV/cn9QuPXxsn0e
vmWcGmJN/UKTm3ll4cq4qnLq/JlOypp097M2XOgifqJXguZwY0GBl0adFNCs
9HgKvIrQJ+/m+8uHdBvYkKKWDOemQVm4wk6/3xrfC+TJ4wzawkdr5WJsQD+z
T/Usb4iD+hMIAVbSeaoZULlenfDgaiTQr2Ey7t17+ZJMTyIsx4vi91FSEZJr
KkcYj9j3RDyGkEFQA3RzD8/QraO0r/KUNxkbCm6S1rsdyBj+qIfy3ZZsgZW+
4NnhAULUISrs3xwikrTR18RvzaPw1UoCu9f00bRR8cuJoDloEn9b2LJlPyLF
BsBSEDFA2JKLUksYWreoJWVxoKQlRU3dw0E8XJ//cq4ZBOXWq3RibHr7OgDL
umseXoUCDCufyGv+A7qMCZpy5RwxuXEfT3M6AnTvMcx542RrCIsmz525X8B4
AAFBXI2TcBiPU+MR+oTCzNTnWFkkUp4Pg4l+PPvb7S1nLYcxyR2yFItuZp7d
XTb6IbvCXPr7OZlZJWgFZ/WguwHKNTAd9YXTe+r3w9ZgoZeyLio28JV81/uZ
36Zi3RTdIU9VDqOyBSS+p+3d0dpGEl+SSc4dhZAEx17pxeu/Pnsn0LbonkFe
qCZQ6whCLyvTzLpMMDn6CUfg52pY11lWzjmfqS0z61lNIEIOOhB4XozpUHod
xWNB8Gw63bVCYKIOFmASV61x+kJ9Vx3aJAgSHDOHPMBqDru5u/q9yZI4KeZ+
jly12K23HaFiJyH6PF1ZMpMmHVD4Cn+C3lqkjp+XFCEIS3+5jqtp7dc1L4yR
/VDlhI506lsuw1O/PW48Vqa9xgyxCvUVdHiFHtapB8JeRSC2CpAOQjPwUJeV
Ipw49yuheiykoXC9T9cpAT80JBeZ5tEwzmHRm6Gp/NDPauKpec9jDoCHDy6D
E0vTuiN9gdMvVbi7Zkne0svAJWGPqz2WAIvqvBAO7KaIMRZ/oTK4NUbcACe8
oVdfCddsGswHBO7Vc6eqD4p9ipKwz9Bnzo3tUxBTpPYhvOtGRNx1z2Ft5PQ+
akKAL2fStYOBVScfdMoDMiIVtjhgMRGDWXFPLezHAI8aDiupsgy92sMrYjt7
iaSnn9DAK9WB+czsxI62OzpK+2gHyLcZPDVHFslFZXZTKBfelxa5zBjYJorQ
rfJiBvOl/ZAQC48q5Z22h9q/ndimOmoiiuAVWO3R3nvOke4q1Gd75/w9cjmD
O4bojkOKQFl6rBYXj+W29h6c2ukyzKV8RPROkICvjY7xmdLfa6Iymk1AVwfo
HYcZFst0We5a72kwpeDZvO64jRwJDBWCJMDd0kPHmQ0GmvD8vLC/lpxAxpkr
9CXAlYHL2QowMUSIOfzYovmvti9ZoGTehi1BOjbg+9RFpD86NymVH0TsuFas
OEbxIqvuza0xeAfxbWQAanmRwCFbn+iU8WKARLlAXEM9iAoTIxeZ7b7kypiq
AZheUMF17qhhM20DAmsECEnjGxsi0VGTkyLMrh+oGMI0h4TlHlGHJjxeWJON
oYDKhkWHj4GrwPBM4I7iSWfbAYtPvg9Xi20Ygs2YWD3Q9PxybJWIAX4Dg+eE
pmtaGudzyPzKKTlus5zNUxBhK1pCFSNoQH5kHon6uAuSRp21IrY2gDIsbqh2
5GYY4Llo/eZzz1PnRXp/v3UaAjWArg8XTVr6pbV0oAu00NLYGB6plEaAG8Lb
S4aVfnvdreWDtudTwhBIigQq8yYyDuhgjkmj/Y1Foo4Dv5TjZu3aYTrnLj+G
I81nFeUIcXlOSN311ycGGc7GlqteaYS4XUjx59PIdbpDKzZoD4Lh7lVdI8Gy
jdfLBkZ1pX/5jHBph44EqaCHygQ7It+VL2uLEffdsbEENozKHnuqFFZbTgTW
ufTDCUs62YzJX2++TIDCpWEkXCGBct1ZyzaheyC9m4N0BRyTpKG+pxUkLvEx
rVijR9rwhCJwSio1BeBRijaFmtIKP/tOdHG2che8EMpDDXBKENg0JlAoEyOE
FCK0l+9QtvARX2wMqGvzs12yAduxcivDL0opbO9Xs6fGHqXzdxx7bpz7hn7l
uNWsWuqUeUqgS1848XhoB9hZcw2wKiSXQ5JWX2jaGJiYIgHdo8sKByKYudV/
0Fiq9bhe0K150px2TP7PRZlzOL5hzFLktniBIhyunymqhg472IGwelLJe1fy
V6Boy+0QE7v1davN/fxTt78G5Z4luwNu3bBOmGSHEiIEe2wJUSmnjYs4LQll
mRcmRtTlXURj+etpTFC4lKOpG8YdaiRMnE9rjzp1AuhGQsvXLvz/igUCOX9W
+Ah7jt3h9qb6mJftfIu3LJgZuFFeFTfCeDL2PMFfICRmt6HWaxheZT+Rbwql
1HaGpL3Tr96WJCmvDQl7i8xwetoaVAf1aiOLO0TreaoWzS9YuUQis0uPceMT
oRuvNVfSIs97F1Vlb3lyYS+aH1AW0tTMLtPEkbbuNaaeC/lOs9sK++7LiP+b
39u+u9hVAlLbuFc/WhlKWFzGRGCqU8FgFCNAAoRQCMLLz+iEINjJbZQXWpIm
0MXpzyxAby2s/yf0CbR21e6qeinzOV2t0jhrxEp1GjaUmf2lqgyyKW1cq4ML
poP4vbwc/qhQXlWGa6nPzdBg6c1oJGlC4Ew2tGv5h3hm/BeBrxoqT1HzcdQB
fsQKmi9qD+o4ImLM7jcUfSygBnwmz1AfQk5hQefwZaMaudB7LRpWfKEZS4J+
0EwTTKNRE9VDXe5zkyLMSvE2vHJ1Za/dqNdYMP8VO/bgmbgxUsENyipgZZbu
8hHLO+fGtVJXValXD65ZMhkvpIhFlOq48QOHwXLXzAsHl457ImZDQPlksqWF
I9p7FA2Fynw32lN77wxLCXqwtGNtvyRisvPqMqmHgL6BSBRXQOfsWFMH9SI3
PLa1I4aGXRVK3suurdvg5fpJtJ7gy+giwe7mq3Q2rAyCYSdTskJN+O8zTmox
x3RhznAMy+2F/7B/rHDaITCVZ60E9qPSnckI2aXMTiJ3TjB9VKBs68aPbZQ+
7IAGn9+Jz8aTRKJSKG3Zg3DilMZqtcHd/yopfIe+pnN+GC4dObkvBd5KQ7nz
JIPY8o7odYHFa5yhewgfmwZMxDxVz/Zmr5VQVws0JyjWgpA0A1yE9vLrULL+
7E2AfIa3lGTvP8RSkWWrRayraMU2txOEnoYVcnonZHFzituWVkkrOS+I1Esd
M8SqGYIjNGTXvvjN3i/JVSuW7Nn+Nessd6lkqXTvJUe5Slt4LdyWVSdEKMnc
zSpgx4Jt8wTGiWKKFPh44La1bNMUYL4nh1hJmwbK/BwJeQfPRL6DfmlpkavL
vV8aDjL8Vq+o++FZpoVDzMcjjd5qLjdO3+2cWtE7IXmqwpxbMrI9uVWVOUch
w/wsMobeDeBFXJDnkavKjMLyPVjMKRU1lF64zZQfgRgGj2qD5f3QGovSXAXI
qCgc6lbjd1JJEqNQhIy394Hw6E/CP5RQob3/kA2kiIst/hOwNqQlFcvICi49
XcrmrSreIHAhW4LpC+rN1CXx1c9QDx+nmIgNSJFVy2P3WhSkxWp7DYhV3cHZ
VGXcf7HlOg7EwnrU/Ck/F1Ttnp836VGprw0crAw5y19Vi/HNX/2pdkQ5MzGD
GkJnIwpGmbg/EyegFUdZnRi+SgLMahBp2MsiltDGx+hGbLQlvJq2GLa73vzL
w2XhS+ctmSJ4I8TkDUuSjSK7+PkRLOGmKnVuOkVe54q9aNaUHu7YFr2QUdWp
S5LmStjvAnvNiUuD0MlRybE5+OQweUv9aysSDET5Sw4LhcecgnCIn1ZylVxy
jcTQ675IofslbBVYebLcwrgK5Ye5ptLFICmzSYsZ3I4E0F1gF3KF0Ar2MCcN
iyJSYDYQc78uND4RL1KJk+8Y4ekwC4cQmNwS9aDCah4VaEtII5d3pLppJfd7
heLitKmWq41ID3QKjyGXmrVAGbuTy7hfZHRMgDycIbkWjIk81ulbi2DGlr9r
IzyBSyn+yP22Io8XnSRGIHvsd2JJfnoA6PXEbgMpyAcGoNUh5PEj+GBxlwxQ
Cj3u7eQ1A8xQeI5u6cA9KfxB0oHLuwy1HCwaPhd3gHB7KHclj+CKoLU4Jwe3
COYzgav3MVZzQ06V2+UdYAt4XTgGyn6uOm+oYQpOFiscwOqFFGnUft6KJYNH
pH2jJQi0Cw+QwvgKIW/jLpNA+P4HTOYQHaaceTiK36onqAkyds20ZBunu6DG
k2fe0by8jbb2jD2sIzw6OkvGyx2Z3qGMhwXU1y3nZd3OQFPEO5K+8tHJ+4uK
nNjZQjWg2WPJ9g7D6cJoWCeosHBcFzak4h53MHJVgOxJKgiK+LPoQjZOnJSp
lJcl96II37R/Bnuq4uM0xGJE0IyCwj4IvYC28nXaxI0du9YBy/7XCZ1WHZlP
Bslw0PWt+vMf2lYZba6ratUHm9AI3YP1oIyMMIRHpEza1V6LaJr4Pgtxe2zX
Ac1ywiUWHTsIot9DCw4Ttg/4ENrYY+tZky1a/xRvfA+WkLVIktxbzIcbHDWe
bfoYB2iYcvuG67w9VTBEOhy1WdGp18/WwVl5ULmkMq6ps2kwdWOE50bpsEyd
5hz1dztBDLmasYXbCnrxcrnFMMI5GmJswTJ1ZmrIK4CSgqhktC45iGDw9WgP
pp0sKydBjNTUIZBxWvCNk50pPxGacmBUTeEjQ7JD/u4EqKpr2Bz9+6sS+1N2
w+GzwhOaBToICLfOQ6RcPZXRz4ZSZ0K6ZJD1zmRZoPDLnT6LyNEJ3BWpCnaY
u1XI5hzPPZtRSl0e9S2ARArBuyQFHlY8zxZgc0rm4F2ONyYcjtJvMs48vE77
pNY94mzJduagppMrPqdLQW/NeVvFMPql7I2ibyvmC4nA1DYfCxrWHfObSfrQ
GQHAuL6bF/ZcYMij7VyyymtZL2wqm31eZYHUBrtye0Z7yRrhZTlYBNH4xw30
petMphx6ATRGs+q3en2Lg67NrHxNmmK/3xLbx3i1+o6LJCpkgFUXnF1DjfQM
dFx2Spr4aFxvyePRQjdIoaZ3UAJrECQcWZ9nHWy8jLj1VJ1Im5Sl1O/4CISi
LTmX5CpPhhWZ2R9pEvhvErW7AlZzsAeYBkUtqKj8PoubZcznYsorSu7SAYKK
PSxomt+CLJp0wyOdM2K0EkbejXnHlE86g8SLe5X833YerYho7SnMB9zdgOyU
AiRRjCaOOYb1e88jQLcpbPIQueRoqhsuyORpfSzQ0PtVZM4fOomuWA7WVFK2
mi9MgCGgCFTSfDgsvdn926XFT4VQrzXiIhBxaPGkxZaLDq7HZinOjME7dIIc
titL0o9/gbeV4lKLHK7cD0fVl/S7RJ2VzZ90zEri/+sQR4IY22gYBTY7w1cD
mTNV0mGPJ239G05q3KRlm24YWrQIH86MElXOfutxrA/e94kU0UaZfFnvmqUT
cyOmgSUYjyhMkuywMrCBDRyeBKMLcD4sh4iaRL2KVkDxhL3gmLX666gnRKMa
DOWm+YZlavzb00UJ479lYJopvV3emd3S+HHmUBoWocgZ5UVftLe9KfO+Qt+3
Y1/FCQ68L1nx8PtUCTgYz5ATM7BOAl/Ee0Qo1N6ayBXO2EyN4jbRs7zXz9pQ
RwzunRWldJ96F5oiYpofEL50Y1Sxaf4aZ5CLzLnpiCRPMnXZmlcPdTZLD2g+
O12/8JUBEbXIQD1/v3aAB0D/42wsj8EqM2P4M0a0sKnOH9hxcRJvRIrBvKpe
UTt9CI6eNd2XQj58LLfNagT+CEwWatPCdnPmzuXEUedyDQy3Sf5SgwgBi8PR
kbCjC4ivMlLEZUSd5RSOrP95sAKVcT8hYAyNMP1FgBpWH9KllSepoiCnjY+g
+qeKI7UtIUPBcslg60yIeKYa4bo2dhDxh5MPqeEEtf+C6sBmDjlWxoQvwv+O
jm0MmIS7kOBmHgDr4aWNBgxxxI9zTREoV5HTKpC6DXjPnFZzWBiOvR9llGcv
3Bhp8BNcvX6++EbVvW22k1XYOUfK8SNrk5UuYe3EO9M1Bg5UpDS7OO7AQK8b
edM4sErZiihZkyHl/y1Y0EZedemXM9ZUO+tEGaegMMpeIgaSkIPz8L4CQKL8
2L5LxDFqdrn5YZ+490xcdHuL6kHpA5wrshPaQwUj7gdJxqgna15OPZHNVt6r
Yca8lP2G9TBTPVTwP3qwnkzBqRODzXSEMoQFYGAuFphB+bWjSUheXhmf6B5I
tbQT1U0s3k2KnPxyjfgBFiRFAS7shSzBG2l5CTo1TcFUepaxIDg5a2bh4HnA
IbslDfAKcD6YgbFNcLvhkMYmG2VxqJ6LgRIJ65lvxtMMbcJbH+o8khoTxZS2
90lvHnLYIWceDI9+7x35o0bY+34D8QQpBGIANCfftCZ5ofIdfFNVRMJM99IQ
OX7x4lE8l9dz/iwan9TT/sKGnwxgdka+ma6IXwJtdF8td2bHpmK4hylDPEXF
s9+dJ5J+QYY+316zogJJ/S0D5Z2za8/sN+Ju1pwM3fpAPB60AqlLvA+B92z/
zpfLiZRsURj6ihx5Wlu2P7q59H5SD0oD/BPsYJEjas8Pj33oEb4IdE7UcPN4
Lh5LYCn9k8IhRKpJU40x10sJbRSdhN7PWEBze/sr4DwXjHWxRZV8ry7WB1bZ
39aIDqVlc5q1bbjcPjCkTb2h859W4cyzq7XoKEyegWSGEx9esNVNi13y77BF
CPxrLy6S2brmzeXs9fa89lYlsyBNWm0NsIZ8BzgvwGJJbZkImskX+1Mzofwe
t6f2+SPl6vDLUDR9SZ4yAdqE/ODaP0g0cpTsQdtdkyvYmNTk2i1y7pG2BOaX
M2+g6wgxUvw0lGloYKDiwVwOAYiBLVxie3izxxBUhmdfrzxvzPhAFPi0JWMx
ZpzeuVRlXcmt8Afh1xToRxDLWuSjhAfiPOWbzVB4jwTnJzTbKWL/g+r+xLzS
94n1xwWxZ4EY02TB1xLiabcUnOwSz8puyncHgNDK45DtjXkkFhNRBACDn+D3
m60LsFCiM2rbZNRbH9lArqiDhnfJQZlc0kpwwqiFGtK7VqmOhG0H+BsfB/xw
s0kdEBvBAc3+ZEJieO+foyr2wiSIJB91iMXNw1axU0X+v2KB/0xcXa8dh5IV
QmuNWWnYLOpoIBE/+z8joLQ/pU+oysmaLhFnqZ63kZs4Rn1S1Hwb8GxAQyZ3
cR8hSThR8Hu1W/tlwGn4o457T0LPmM+ajzCvEXoAutKlkVeNs3EfxpwNKrBo
jEoLK794VGkqN0bJnyBwz5m5XZMA1TRKztuJelzmHcVuPGmyJ/ivSVp9vVx9
hFKLx9Obm3RQtVgHuI46LaAA36bGI5jy8pacTiCmfBTEIbHDq3jn+p/oUnrQ
FH/5mW8/xt4+wlx0GgVjv+als1BmAmuLscd1Kl7S05wnwXjJct6p8AslIa9K
JYQ7/s7Gb8bxsARJDtJhwtLqAalqmC4mmI8qs7JPW9wNwTg4/Hx5BM0YWYy5
X5EDERdFZsOCJZZwCWOpT4jFBxWrVcTNzMJbXjCJfRV4rFMsIuwgQb7v3Msk
vVv81Lq36yqVRvTEShrLXBvPOAV1yISN2UNuRj8RdKXdMA5ufu9QEMjhKQLU
doCqsIgn0fpAmTOVOwaA8MGyEjmozAXR7KKt5m1megmEj7iDsneVfMDyuPMB
JaYimKlRrMnqCGV1h6EYFCKlhvacL0ik6JAQ1B60NtD7aMg28le9kfVYjwgv
TIhTTzFzjIBZPVmEiQ/zu69h5fr4tRCQdR92SIgDnIDnky5gS8eYkq6Suawm
x/Mg1B3PqwkUA5fufvlmAVylz171rwZvna1+nFxkc1R+wVShd6RrS6l8Y0+q
pCtUjL8rmBR8+q50GCBRqUsbZUAQPDLiOl4Zw7NAfCfeh9wYhtJSMtPJcytn
ktw41/X84m/gR62Sl9u5LtSkYMpUlwiQlgEvRlzGkqQ2EhUBVRxtEJXrbr2W
DxxTh7HaTBpczIpAY+P2OudDQEksD7+UkdByd7seSj2vKHjcqYGKtrOWLDRv
6QahLvSA9cqNSd74jMNPXwrka7c6wb6JlmK3lPfRwOViE78oiPGaAJN6ax3J
AFhJ3CcqL5S1+3rYW1xUT+eq9w5oEhjsd2xERhyhAuU7HyZwSAP1E5aTeRRH
bgpfDbq2q6rw96MeK0g8titT8Do2RRO/GK9aayUqUsiQNCOE7TLRDJrDW/gs
lLFCTaYDoXRTNpVYW32AlQpqZbnz4FlnCZeqDzQyoET32+n4ZRwavMcwCN2v
ohjM3Xw8uQiu90fYTTDzTdsi7poC0DnXNLLIpA6ai/n5VIDliEBzWiCdmwPG
OWe6MWSOpNn27+tdSB/5nLE67hW1NDNOqTsI8FUAosW+wAtggIWZmdZ3GaUm
bdMLLzyLQMYKZb7HU0xjEExKCWA9hnhBdYvsdzRgQEUWwNobMW+PiPR2Jz0w
7vi1SmD0KDHwbsbwPmeJixDJxq2PLYXWAf3cCn68aD4xyOkuySeo8zNzBbi9
beFSu6vnvc3iz8kkWPXn8GiTU4sFWW36RXqPZ7vdX247KBf59i0nUMfX9vdP
c860Cwn3LhrBFQu/6gTBy2d1Dc33wQTxy6wawe9XKQbv8Cuw7rPJbZmAXeVS
xYXSN0/Wkxc+BIjkxTHRF7YHg8ocZkBRzWL4YyUzjSglCJgS/pYDVDJULdww
6IOQDnQ5oVUt5rdy8DjbriyLMJxN/l2SV/KELgBnRki0N2tehwu25mCcbGMY
Jsms5s3X9Y50ZYmOG+UOVxt7jhkAvS1JfqGtL6TOUpjBeTYB3jcJWISC9I2U
f/RX38RRTJ9TdY1BwbkYVQgNzTRJW5yK74LrD7pd+FwrqWTIeQTHCcocaE/D
BRNNiBhzfBgn16lOD6QpIkxFgcgyDhvNZAlivKCrq4OLBX73t+lC+Pd2OXy4
AdsvHfYquQgFrlDL9CQqs/qDHU8j35h1lLjQrqyqSkdFWhOYJ8KDdSBbsd0q
XTionmH4uSeyQxoTmZZPkHXStQ+PXujnx+waVXvZjuYcNUOD32Dw83XpBF/1
jLM62RGaPLp+BWXVmH9Vxakpx0lxlLIMp4mmkjjRctpF+OfMePZcHn4QoZua
fui+Kb7VQ0x1avZGdsxmLtzwQAf5bM4nzIrLKCp+KSRjxZKHiCA5X+9e/Czd
Fn0VQwGouNXU8sls8N+kd8kHQax8+lyXnB3G9lQoRvaNHpQYroKCi75HF39N
bSvsrB1c+hDOWOuYg9S7wRpaxh3b2gdlZkgCPFDSlsmXnCZne52KlaXH5Qdt
CjETj2rnUChxfsnr+w5tVHtxlR4q3cdm4JmbT+ZufIbCMi0tZ0DmZj3blYtX
tSSXEmAHLZI2im2F7RYeMG5kKxaw890rZF5p40+QUUDWKD297aUyy1mxftRd
hCn+XbmDFuaw7WwfO+g3EOeHiIwnLupbdO55b7goKtlid+GrJRS7vWKo0Fyj
oz4Mj66q03W771l48mDAFKmiB4HLyEkN/t7ykcDgR5ESG/xe+nYYjpso4Qi+
+btkULBaD+BPICh3wUft8yHmPZ3y85N3AOfHu1ZXR2zxwhcHMD3h+oHf8zKr
VBXw+dIIBN94xnQ0ln/xnfuAwgjO72i7AGFQnH5bAVoWp+wmB2fOHN35EtZh
oyoClBmrOpamtch6hQRxLL9fHVz1U1kUWaYjXv8o8s7cq59q+6Cqe7T2dM3n
U9hm4nuSQOa+ju+Yhwsc3eRt/7Hvz+C68fLiQE49g3bWaWEC2BifcYCc0JER
ef/e1Kcc05BQ+RVu1lKpswSTneitsHBw075lvjZ3u16dVGEjI3Dk2zV1Uxml
NEXhWEhEstztPcsBe4ObjJi3RUgZjuFJg9qUrdO6D9jzDL7fzCnl4KKycPZv
BFx0n/E7/Oa2NSAOgwVryG0/3S+2kI3IjerryDEH8mM7kmHvL1SjbX7MiP8h
O9L5HfnDscGjmMtr0sxMg88DqRPutO1v88OH3r4NHAYPQpOjJmNyOM8raCag
6mYKsy0DYtJKqESrz47lJdhtdfewY4AAlu8yH/Z5NxwtHSZexyOmh4McV4a7
mr/y0ihcLO3WteMGa4T7gjZs6noz9v6/sgCJ+/ekL1+DqrCUWyIi8rF5LVte
IpnhEWvijo5TehgoJsXyZQWHBaAiJEG5dH3BKeLidfXL0i7h1rcrjKZBLMu4
9lpdfFOcSeCDcFkXBBThIwn7zK7IPo/idwXxnLH93vgX0s/h3mdJ81lHDbSC
3NcXmpMxEW58+2qrvrWv0gBtOHKenidfZL5mo+NhaFUWIpVXHqq5J38qK04r
DZugEnroww1k9LigkcjZRFd/if05MuY2G29iUsXQycMsUOSj+ZtjZEivhYK4
Abu3KQDnrRAw5iC+b039x4YFra0dBhyxdlOUeRhgDJU1lBRCERspD97OKLOK
jR1If8gMjhinkkYwip/UW39YgWgNjeZPQ64+ttawYE7SQyBg+UxfHJEiIGPJ
rWTtgUzVKtW/U0RblvI+RckYKSxHv5yKQlXvyLAyK4z3eVPfo5x9usx7omJx
Bj3boggajmHYWHvWWNXvGgDOs2ARjvJpWuR747Ts00mtUOla+XWX1Wwsc5vM
04tT8updq1PN3zlYLhKuGM8emnvyewX+t5MnyJEcJAmJkg4Kss0e8Z2ekSxo
kzLRBgxDmgN3BzqlDLkoNG+QCQkt9aEzfZjcCeg9zX0CC55kPtXiwyY2qTsV
OOAaUVoNshe8UzNy/RMZ6PJdhXA4dndB1SuOk3IB+pGv85lRPIhvRiPxlBiG
W11Va0admdUgtLClY3lmPAr3pQfqAegPDinZPnPtEGboSJXpnbcObfdUg+G4
fVzQBeVrenbCj9RhNIzLwVtMayz/RvAtmtkwG3VqZDcMy2L4mOaOz1HGC2OC
c9HDqZO6aCYNhPpNbwvEdYLTFpHw28H3/HtaZ3p0xYh4hVTJpNPPQQsFRQFr
FR2Q4vuCMYPL/UTrY8o4x4MtZ9sme/C9mUShitMxf75ON7/mYqN8lzR9Kudj
NkdRakNpNEcPukc+Bd/AdJ8Rvu1hp2GNjYMUiivlTBevUj/oOv45OuQwzqrC
a5QcYl6G5N73aVG+Ws7nt00Euf4ieiqLc19jhqw/q+O+LOwvDojCc85Mad6c
UwkujIYFjtv5hCYaZJZYJJtgfKXbyzCcYKckke7u70s4tjf7LfhGC+H6+ms5
rOD4DMb8tun3bvwnfXyYcAWk/9ozmU2SYRxq7YVdLDvg2B1VOtk3/OfJjYAB
3j2GBVrjhHptPXu1I/RN+JvZIugMhkcV9zAMSPwO1IBg86Jgtiaa2XjemIEx
dlOwTztUFuABqBW89wbcXimCvsJLFqU9BKmORVhHiGHZmZeFxFzTZs4g+vyZ
Knr1VB0wYyVa4mznhGff6m5rhCTFueiz9OMdLcNkFvFEybhnEiSGZGg3U4zP
99nF+WnRq9i1W/kcQflvSyTwrvLR6T8stD8Sy151qm57KYBFRj9yyh7+H35U
xTCKdM/nBPflhr2rnEE8R/HFROjJ4kI5WCS3kGNkbKPjZujMFXnq8FeOcY96
/SpA2u3wRVl0LUoXFXxcs6ZfJydNEinpiKNx1S/MI0o0q5G4DnnMOPmWaSuh
lDMffm0sG24Gd4+UKBihAzJz0N0SkyysjT8l4e32CVxo3wHbID5Z9ljExD5s
FZ4iPnZstw0m5yeA4f2FX/h5rvTd1ERzwv8YntPkjkqedlmUJi9gg6sZSsan
tvDQV8KBA1UKBIA6Y8Zy6CgkkuELmwuB96i0mgfXOWE1GrytuJTgZOtEaPtV
wt6dI+AQ0QoC9UiEg24RidWR3i6PNktGrwpR6ceJIOvv1TipNjZ7acNNYCoB
9G6FWSQnVYLFIZtgAtct4VvDao41bZoC/MGqcjdlpiqwYijS8cdY/4CFTqhm
EUJQoiuw9RFvPm7Ti8OIXOC8oNGFWVmiCsRetUUdo49X+nh909mEcaZrFjpI
mipRapGHmrWKIWRm3I9uKuRS76HRfp/XqrNd4sy79jayhM4++/tiFo9MWYuL
8yM3JBPR9EIccedRnN4mESp1yn8uLZQuracOKB+U/gnmAtZeJ8FWoY53s2oD
CuHPVOjtKEH3HL7ggn9MO8ayMS0qbMTxskWzYerc3U2fBrPU97jfJ17sKjX1
b3MNax6nB7ieSqExrU/uLkY4gRqFK5tFaDy3lgpUyv0MX0opGQg5hJLQvexp
Ohy1PY3m7AAVOH/pmzmSxqvRVbYrJfvyKNPyfpnxKDUJs8+60Xt/RZImnuRL
886vLPevlZ+imG3y5SYe8flov7itUVFUqmqUk/e0Gi7/Q3DXhvyrmmCSn+WJ
b8Xb4l6TZzGlm2Hq65tp6zeKllBsSl6rzh/XVJOfOW2afK/ZMFOZsGxZXnDB
OXyx7fdze8M+KpILv6ne41f9mSb5gzoT/LEQzXfLFsfBRkUaeiniKPF864Yz
7W3mDkL79ZkSP8cJe7iPWVZXByNRnQfazDiiGPyXVpva4tBBQofbJmJw65bi
MHldv1qkCUJEbsZBZOz9czPYfy+PmoyNsGgPAtVtcIfJ9fGOpCsfQs/WtyKN
UIaSMVh0cajwYK2MeSr2Qe32MXB2WvSSgteJFckHytNmXPLvoiHPKklEZucN
ijxza+wu7PO/nX2/E/M5IkcJoDIoOTDHZAQ5GAKQ6B2avdwpvdUuVCnTxWTV
ceMrl0BjD6rPk+4XbEzkTHvYeJU9V/pPDBXrCaXtyf5/9uxbmwuEIfLVx7MZ
1B0yT4wFNeJO9Ybo2LQK7uC7/+uGLq6Eu/1nX2HFKQoFkNHMzfNFRcJHHvWy
/XTNzacNeAdu9SAqZFl+f0ToNe18SfdUCSbp+JWR7g0PAtvQx4Dk5lDHGFiE
iKcn7dgOFaDB+3I8p2TchNN+/I/Xg07kTAPgqD45Njja/7JNdimv8tLwOPgE
dyBoaEqUniPSJE7EnhINhUuZvvXVh+g2azK2RdFBM7GmigAcU/DhkP0M7Dd+
QqbByw/fLLSggQE8TgmBS8vzeHbVdtpobIuxCPpWto1gz7cVCIgowgowGjk3
6Rx1zXGEY8NiU4W1iNkjtywCNI3Ghn1RvTH3SgpgJhYDznrOn7S711LOB+4u
Sb08wDnbEMJEDWREE+OZojHNzk37onSYyz7GuG+rrHdaGIGW9JIw+VODFANy
R1/0EQ7ToDIfsx0suqAcMehzlyZy7dLjm3pGs3/OpA4AwgKZb2jRCqNx59kv
+QP7uerMnIHwa29iO6dXrH+vc69gYlXYagXKMiNftGtnH1lgG3RlACjlawbS
orzmIDemImosB3BjGZGjuz0OtZ1Kp9nhyiU9tmEBQWf0CvIujekGfAm52lUW
vFqrPgKeGi595GOeCWT61jRQmvV1Ij/JqHGCQo9SiiVsI8UaCm7N1osv5qyy
dYpD4C7OBH109BnnE2wQPLu52+E7itiSLz98/rQupcpJ2Te44KErEOBXrP37
xpuleve6zwGIYlo2aZob6XE3zfsqI2DSZ1poWZxgOLtYhO6oefQDCGOxzw2q
cS7hc5h6egef8WDvtOH2ZjQMCa/ywRePY0hxeMhjlFuFe+BPwBLJWLiHzT9z
oBJR07puDeMlWDHvNOB8KtNYITVdM7w9S+7mpuP4N4+eBque/JQOWGC71qOM
o2i0wpJb9Ck5cPnXTf5OUoEO/u0bJT+shOk5oP0DPDNx4MKeVWsZMOriLoD5
GKHDiwVseobix8j7tQTi3WrV8DjIVmR+aEAUqSmWNNQd49uWIX+FbgInbjyJ
NR5SyG9ASjsVzTh7MKFIt97gT90D69CIUIQBCGPnr3QE5xzNXGMF64pYywwe
N9JARdaWiDNPD4pzyKnUmZR5m+oT/j3Vpc5CdI5C/KtLoddVq2Zd3usIV/Au
T3icZeArMctpKMnWoSBGeQvSEAaThMl412l4j1rVWhKcxjKgyBFR84uPKSKG
lY9XjI3EZsiH+MOJdRARRsWDLe4JjrpxPtwG8YgGpdQm92dwlUxM4wPvzov0
eslFORJ30qKzMN0tsrRBq07ep7D7emgfDuMRP8I3FYu40vmRsAe8Z6k2QYaA
8EmNXT8VBe4iYYBGJ4nisVvmaTq5HOWadATNAo0mWD77Nc8uymFOQAzQ1Klp
dXYUyCUak9tpHo+Jch+22hsl1AtavLsxjXOZAOoTuNyEM3u2thCrLiJ+inMa
TIB9izRib5C2BnyfMy5+HM9+NwUWrs8slj283Ibb2I1qmKQIg5T3zWaLbK0x
piYCIj7UACYPa5A/ss0Sd5WHaOMdMj3QFE+lksR5+NqHjLbioV7u02Td3SBM
4GKMXtKnD/UM8c5JGRzJMUPJPbIeWq10+K85JKtrOqMvt7bxiKxGf+zLjb4i
CZmAeKoihTLdjAVVCYv7s0c70ntnXmbWcGPaeEy/Fhdo64gt6BwTemoAdjZj
tEp98cZGXJleG398KyIlO3dqO+L6HxN+SlJit2Xgbj1cmZo0c4ngY8iyVZgm
/Ca1KxhJSdpYaTmM0YSG33QFjqZ/Jdl4+uN9MCbPpSiJwhc1LAY7duFuCwPx
BiDJpXlBSApJO9n/c2Dq5v2OOOOF/Gldha7qJBthux6kIBIWbKmZGLrl/XBT
32o7W+7Oud7NiKstQm5je1BT66ZFA00xWJoFcCZg+UKSUgMbhzeRwKGy6amO
5Ed4Cf/t68xv/dA2+azINLPqdC4PvKjr3Tb/Wbsmd1tFecdGg8QWZZLy8Le9
bw0yG1bOzwp1VTf1Awk2ALGpYcjjoTATYeQAxQqidQQFF9h+6rbBt63kDdDt
RT3BGbGW27KKbxbTxuEHoPfaoTt9nH8h8te5gqPcw/A4cm4L7UgjqoaxzcUp
48K691fvzpxpy41daMxDGz3PEZ/KRXZWFM2IkhfFVXg4+JcKuuhpmi60fgEm
nYPb3ZimghklzYBt+ozL4jeF7mokU725w5WZHv7QZ1bvGU+p0zocLFY31F/o
0mV2CdD/ZSE69BWMyovPZEWAKjR1ekyYwiSL0FRd4GxWJeVOm6sF1KhvIMBH
WAhIaelMvQfgNa+8LuUG94Q5kg5rhiB62nqr7afFGtEDODvrRJTzicUXVajS
ZKUgAImbSbZHDvhRaTaoumz0P9BagMLpGvEX0nUftjqhCgNp/fz0Ipd6baPz
+JlWlH6wl81uw0nBdaCE1gXmZkc8OwmCEuYok2DgXVZmv0hFGr2xCoOWaQln
2AwHuH0ZK7fq9ZOdy1fISIR7tk4OReRMuD9Q1yrzXz80BKLDeTVsNwY18gxo
bLkxMT1+xchoYfUWSPAPgkUNytHNAVCF1zEOShV/iWdBkQ1Fm6TdO+8zFTuD
l49F+Wz78lKpiPQoRBaKBv2r+OHNXMDm1GUFanf8wz0WFmogWEL7f2ht9UZC
kPniEM5BklznzvDQ114BOdCatrykcVZDz92RAFlWmKe4QpqEUOmzH6ZraX3F
bsAlbpZhnYA9hbH/WDM4eM7hkyEcpUOQ7QgXCyQzCsO54SkRsXhWMrVmOwiF
ba9wbJsX5N9NE22NEmFcHhcLmH1FbWbh0Hof8RWR/XOz5j1OU7ClGkOSx7rZ
B1BqIikHYvaZ1z439O8TAlJ1zYPgaaAOXeFZEslPaAwCR1Rd0UBCwLmd67A1
ZqGrChoS/Wt9js9NkdzXQjxz/PYjTgEdyheoyrrnFlXE+04cDxA9SUjsHD8F
iSNtMGZ4C2wXF/ESQkxmkfaMJdteLKalT6WB8cd4Bj+oOEvnPsVTLmtxgJtz
6LarAiCcG05rVD052mn5Fn/Mt+k3H0zRLtE29hAwYRzEpPRHmaYVl3H943AI
Cg2tvNRWomhLY6dja9u9wZ4ZaQaOVXyYEICmb4bm8LODx2h8pMbBX7p/N/YP
MRcL3HPGJfa5DPIF4g6bbCNk5ZYtK+QpZXAwwHs39bnFGR/l3y58NpYQHIC/
wL0f3iVaAakFYCs7aThlHAhC+rYH6UX0J/ne1OfGdM4f+/8Lr3nFCl85Eh1O
dhzZmg9ldMeBPA58CsoUYeKF7NJ5/SAV56LxlDyRGdR82dVJIyOyfgCVA+Kb
tSvWRjd9ogaDCA7e7ygSxPEGSqiNiXd/jd4NAWQfR8LIVNpmCvdnjX5GppBG
4afUxSDy2i47PmAjrwl9/TnIwtXDVfvc9RXiLCcp9E+IaPWqTOemx8QxQIwR
RY2V16sT4kBMR6llJ4MMpX+1IuMWVy9le8PleENz9rX5NVUeSWpGmYEEG52J
OVauKCuEFEDH7+DYsafj/ayMcSwhYzgt2gcq4douqQWreKqKK9DpWXFJ4gxA
a14JBzfsNz5awtFbRmc6uDI5/0f9w015DncAccCTUpsPNNo7C7UI/QLuyu5P
akO1PC5n+Ad+NvKXp4TzsLPV0o+wKz79uPefPyeoORhEqE8rYe7IE7G5623y
KoPZaHAR8NTrNhjlzqSDDfFmZKyGCWmdi3Ko2RnM5EhxVS2DVRkVSTZ7YGYV
jZUc06iRZEdM6TDsGXEIK1b3RNW/G8YrILjSJmcYQu9WirhWkoAnUw+X+Mmt
NW9kRME/Klpeps0ok+b1UTu4DkI5Eahh9KLLGb9DTrF1XFHOaA5Oy/8q2f6z
EqlEGSCJnVEUjsFcwvEc+JsYP1WUQNYRkYgglDzwr0CTGiXntwe1usz4RMXD
C9mGsFx1hhQ50dg5cQfmt5mw2I953xuyEB4wI4csvHQnlonp2kwyMNw6T1Q8
nTXnuHYFF3CAoEOBHnUyGGn3pYqlHz3V4s6w8K0qSQTDR8ePBluziEyucurK
U8O7RpDDnNN58kovWyDFzAaL8lKM5P0MHZpB0JKvScBxnu9jfGzJt2J0R6sE
t5P4zOxt+jyihEVEUnxr8AidTZJCwLWhsPCGHKwj69U1L8JMKfNxm5QLZhbj
PpVxHU8SkuXI+LQWOGA+GeFrmJgsQx3iDnXSBSl46sIoJHwUAF0prsSbjK12
pUZ9GDwmabrRnfoaL2F9fWCE8moZZA7AwxxGAF1gxHTv+zU/BqP2asnaun6T
pNHHZ4BvTUOayhdPjfKrHYeMOkkmdbMGAlaWECsHdcbekTlqnym2twRU1jK6
TsHIkNdnxIBoCFJTOmOwRQ4+cFvfXt7NHt0bo7OeBwuo8Yesamm1q1VcBera
0CsSrPzLbABnTQQ96QuqNI7KkR5QvQx3qWLfKHylyTN/oZuiXOKlOv66Up6f
m8Bwka/Vcrf+MaxGNXVMt+VWlt6xkW2jqawB+Al/hEex0khwmB0S4qkaBRJs
ghdWpkV2i6yGNIeEHOBhxljqe7OW+2GNgFwdNfGc878f7IVbhgKHvUeu9cBu
geQXyEzqYXyFIF1cPMTzeUKXvJxsHVIZv2P6RyDqhzhPabFDPZ3OCfICYuTd
MaYVrtT0QcPItH3hIcE83qC9R6A2yMrqyBsgnMuUACtlmRTyQuhHbgGc3TBa
wFRoawJGcbay/U06dBlwkmobko+7mc4yD4AimTz0VBU3CrchrqmjjMrsSJ3z
iqVTIBBTodE/Iv9gBFR9fzEqYstpR5HEr2+C2PoQbGQ6TO1JuBHYt2+/zt5/
amCaeQqr7jZZ2CFY7rDWovwnmy6tMh2ZBvkOmlQMsb8rCCD9CJl5fRUYSFHz
ffoN+yFJev+FlMtW8iPw9DKXYlr2yWCp/XCodVB3tqgMsoQwLKBT0YZ+d13M
FxfUaGU/i2VwNficopmsGcy7t0JZ5cHmVD7vHzq3CFuv5trO2QF8C4SW1/C6
kbDE3mv2abfDQ3bZSk2AJrddKyWeqG7IFcrDMTc3D0/KQ4s6Ngh9Ys8g4KIH
TgJDRnPQRn9C+cuSECxn6LDXkNr9PU+a92C0/T7YQ6Kf8jvt6gDs92zx2HER
gxfKuQ89cPNVdGUG9sHpGLn507At9iYePseP4Z4b8RTgHnD7jlnw7GqzzxF7
bTmL76fF7mSeVWOrjU5jhg/mkgsmgD27zMn3sFMcDwwuAkgGC4uXFcpY9jrW
QK0ReF9HnuvRzZ/3o4Rkvve/78VJbYIWE+BmitynrXj+YauLWPmYoYuXk5s5
qCf1/IExFGirN3g9+NQA8nx027E3k52JBXAQa5dO5FBGDVqYZqU47ccjBV8G
rQ7TNI6njjnL9//5MqYhR6gDP2mx1gtKdf0DP8jqoI21qn/xbYxJpK2CPhC1
hnX967chmyKE31RF/DK+o1IEZKG6RmII8RrDDknjOcCqjJbJ9lox4Can6r5j
LNti05hNVFn23UsiZau0RU5lkE/PmZi77qbqoWekITtRqUuPKVfUAqulMVJ7
902Mm+1rBKKilw6dZaYVECttvMEWXCXZ78kT/R+uoT68NPgj4o2iAx0Dp8/p
JkQ+FGhr+Ovj+iyMtrSDyLy3CILosGPMytGmkOetbhZdFOozY9JN5YnKiAiI
xZXXQyt9rfOo/fWxy3ieUt6y/Su/Ww1v0yyCV8D/YdxuHrnRYI2PGLmNRAFq
iuEhGfYDWf2nkRvEKy/ItSNXlbYPdaDCL0pSmdnOFplTb9aQ2KDWDksEJBxV
SnkGqYbjXTb/6sE2T/fvzPVEkbMuErA5FawmRniQiuxCgy1/4XWapnjW9RMw
mi+UBvoAJsNne6FmjM6l4kY2SK8JGUgv5OLckAV7m1QHZx0CfB/3lCiGeTKB
YFwO5O+HAeE1Q9YOQ4yFTDsncPjuhUttuKAoNfWrd4oT80twZtoW+h7K4QuV
hP8VyhkzGewwHAJ8npuKBNF630GyB4Hhq/ylaKQV2o7hEBdz0ocf6lZmX67u
CqNUo/VLhuKnqctalvJ8+wQSYdyxLNRsqU/+Oy1/4AR9jvLTwvH5W//RpPwY
1vwKzNlpgBaHs6Z45R+pZyO7g86jeVipevBqEEuQP/YkwdZ17fY8CLsMuwPW
xllq5L+3fTZgGyBI8Txv2Gx5XKwc+Qtj6vFvMEUwhs+1KrMTwj8L3I8YsiZS
5n26mbwgWSA0B7GJX5NPUWm19Yr48W5ApyJ6zQ3UueMfA3Hgdjm6DkwHW4Xw
7IdaVTy6orzhAFyEK5Gmj6XTzjSCEnaItusuu7ABGfTNKE7bFbEqHQhGBA/g
ni6yIc+L1CvnLSPIiQ4QjA2DJEBuOHzhcsILnJmaFODRkCtT8XqszzTGLqB+
fkM97iNVZHHkMcdQhCbvp4MSMRG0OZq0xBO8YJxxum1auHwzzX3iHKXG6Tyc
g1yEwmUbSnSSHsWc/jk31XK1e+HC4Wbwp8quYBw7WhRphb2HQaLD+zNbQdnq
PRefG7MJQ2yUwqNL5p4WnO9ylfXVEb49bX4QtUuF7XD7W28gxEn/QE5UuXHZ
yXpOGnAb0G5SQIviZvJGCOtUXKlL/ey5ZvhhODyYtnm8WcshNdw/XLIRlxVc
XWaFSq7/cZah6qlIFmT2RxQmst/03qvkGL1JKsMRWU/1mzM5rDoXzvyvmzpR
cdvlT/sFhmD7WgoY6FAsNbZH4WbKvNTpqB4vev89h7dvyZFuXch3akEWiavB
nwS8fxIb7HHAk5O+V1hn6EzeopQKXEN5f3vUAvzsBXpspg2NECSP9+h3Zk5X
be5peY1Bh51ltcTFyMUXRZ9BoLNTyqgEfbtmDSefzdgI1LEFS73FCixpSAvn
KKgORz11gC5GPh84gqONTkbEtdxk3RYRAI8nFkiTkmQ569VfJ1RA/u2mxrFn
M5zJ2MzmpwVfm2A6sElQKaVx/siDLhoKQhhKxeg6QwF0Zk7Qo+xmsjL10zpT
+3FTIRH7TniMQLQpSS4qDaz8XMHECA5LZvLI5NII/zTyXm0/UjbZxdUaJPLX
NVlQC1tIvXZp5YwGSo0oRx2T2KqTSHhxamjabnC/FF21/kMU+F6sN4jp5/vc
TqW/sFbo3Bl8FcoTEyW5FUCG/RNpBWtkKz6JqHA/VOjHpsMHJPPi2VpuSS0A
atEnXj+EWG3WBWs3VGZtUPD/NPRcRbhf5ROAnyJXMEFoCK2RoRbNDdIc7Gxn
FPn3LH5pxsbhZ58erjoHG5Kp1t0TpAWtj4CbJMI355D/1jGR5ED9VkTt3y5c
CRKUEvdU/7T+9maAoBKZ6fz4DJECIrf54bsc6tfdvUbID0HMtXH1+4YpBoI5
9EDULAKzTSvH7Ui18eu9t4WWDEFdhN4t+ecPgfWyvhGX/KdSJKzejDOKUPjX
21t5sCGx0c6iHw28Y1u90ZEhtaq+X1gJcTJ4ECximthRvwdgw+pCA6MHppYF
TCKLcYU6nQzobGNQxvbHu1A6msrYrWpga4JR70SS6zEsn1bFAeyW50hk3zpY
5MWsAAip6z7eA43oTrT0CGaHuTLMXceJa8lL4eOEVGY77eQLhmVauOcpLxOv
2DDgyhWR9b7CvKSqYorCpLClKjXmwUgkx3wba2AOrkCOvMa56+HsLm9W95pA
fEIVpmlpivAwfciw3VBJchw5t5ZYp8a+k8wZLImqV08jIvvyHS2ibx60rfSE
AMWMKop8C7I7jlUkhx8iWcikPvFgVzrAHzK6qIrJb1/XUZbVpLb46Z5ouxsl
qcQ6Nx31nMtUQ6s5WmU8QzXr6dyACG/H/gpUoGxoP9/u1Bo8kQK4w/ufm15x
TSaLdPjGvrDCMkPw1dtgCq4sJ/8dcPQTniTmYMFzwjkwd2iJk+egseeBCud4
eFkZMQWjErnxHTtFgCfYzpH+OyK03DM6tc7JUuez9tQQq9EbUzJ5oEDdip+o
IAspZDrtBnjedwXqwlyVnbVlOkL7mCaGtC08U7BoLosUQE8I7nAAN4amgy7X
ALzSuTKc4Ho/TNUE6Y7sNqEbrSVSLdRo+uYAFuRJepuZrrtQNId8ZbDaD31G
OJ80j7rWaxs56CO5IM/mT3piL3nPRMkOMLCGngArQbANKPuKjxz9rSFefY8g
TlBwffLyEl/iPMs14jnL1VyFFBPomJqTb760aneKw2DOcTwXC9kciOHyMtGX
PWoyyFaTH10i/GYpHIpJKOXL3aW/qUxGH5S4RfVWYNMXAqOCAuETR6ZPnUqd
TfpP6oPCKL5W7tH90lm2pL2jmxtqCgEckq3wOEYQuvugO8J4j/dkgLXNMKJH
bfiNx/sjrApolLx/PYPRoixJG5SctyOfM4RG/jVgNbWBYOUi4jaNbqmbp5Zs
X5Pv2qFKJi6vzqnNcjuoyQ3kxvRCphW/0pA9q5DEqx1paR3D8yfOnm29Cclp
JPaifRHSMYvedYMutsNUuisN3cch9cgSeiuG6Yhvwis+zMnT49fJHXcgs8Aq
ONjV/Tnv/oioKg22aUbTn8JFhjhe1EjegO+7fw9eOkJfMgkwFQUqNBYaPvw7
GHhGJGseBndBWDuXvEeiFeeXn3FFAX9HiyD5eftuqF9CbEx9FtimUqilRNIU
U65IRn+RWVMdhyC/friEsj0cZd5sqvU+pSM62L6SpiHeOfM8+DaLu/iM2q3e
5O33RZ3BQBfpipJZ9g8meEvBJSZfjpuZmpKNnYtuZng/jUSvab7nKwfKVkYg
vewqtndgYYjLm42TEnPUpwuuqzvqej8ZcP2VhIYFww7dpIdei/py72rJL7Nw
iu68t1Y7U9WijTPTpamHWp/6V8TM3mpc+bIPJTAgSYWjsLIoo5b1RWjw8c8e
FvDMEtIDBp7l1qnmID03eYnYwbgG1VRuPA2OiCZGE4n2b7LAUkspfbYKQ7n4
p0NKT01psyr0K6cc1DWnHTjftnMi2RAzTwUJn9BgfK/MLvq+YN+nIBKDOy3N
LWv5zLKc9VK7TGyyOEcdj9PxDspH60AgGmCsR/hbcozBTphl7JCcULB0uc2l
W2WwemPTd96g/qg3QMa1fBsKbrjp9xn4psy4YVTkrpFWWEllWVGO3dFlYFF8
2LGfFKV+UGM7xk8JxwI+bgGcPHpIYtFMOAQRAAPnmUBhi0OTbQcFBAqbkpeG
x5yULKr83EzLfon3ok1X9eM2wNGy8B8RtNhhkkETZJKp8l/hoK0r99Ngc5+k
mAQWjre8x4OyoxV5PBUpwtpq8sdAU+A1baSSdwWKBhBhhZVjxsqMh+gj6lf1
K08OC1ZOlJ+Nw00dQUZmB+yn8NeGAbaCGG+cl0HTICyhEgBLfUqUhNDeK5aJ
FMrNzLgrVI3TDBVb73NuCgX5kilVTsvY1JvrevwtecnrDsMBPyxLjtRR9NPs
yYi6mrybZ1RTQ75rAfQFSE11fM+T9JlVJhUJ25+C6T0goM5EuezQI611JeNA
Ty+i/X9MvHoq0ierRe1cfZQAhhNR6vHYOlmQXISo3bg8DaNKv0i+E1/G2KV3
8fJu62nbvX/alsPhBvOcazsawdM+c/qKEnPwJ96wUuuTwRWpeEGW71m67Hw1
a/qLKHZWTL1rVLknEljANy0gcz21i5n+kmC7z5wWf/e6ak+RNzgR6vlOhbiI
0nISVHlA4ZKMowwtVBM4FX4qkN8M/UL4EVOFPJ0v8V1tO2rrejWb6niBI1un
kbiaNdJcT7IS8MzlgHCmwAYUoHkWXl9oDrixrRfRYILE/IgGIAqLQEZM5Yfl
tD9SHuI6AIKz0u0K6daj7d+JAeBPtiaGjzTed38DFMcSIbUCeLpnT+mgR6Mt
tH4r5shZ1rFvRC/oTg+oMQ+PFKtgQf3xCaSUbZJi6W4bBjw/mFlBvYlTwxLe
Hri8/bnQ8XPYypzjfauBZ5dDHcaH+Up7Cez4U45XTrEzbZ28WMZDdhPJMtQd
1ucAsDQIztls967AbqsCtAdk7vHI8+IaRRkIhxNbPh8vCxNtkk8Q4raHimOX
RN5l+0ALMTSSSEeyDxpdsH/Iefn35hqw3eh63RMixaPr4RQ3FzxWdj0cJ6Ms
E5CmLkw96ewFcxy/fXFyXE9Qoiael8saUTcLs8E0R6u6zM1KC9pr72RC8tCG
3ZgPoMVCkVobbznLyiK1gOP2M53zrU2XhBoyNafYSfOVyohW+l+mEUgk9sUZ
KugJicBSFgLCWzXp0Ac5kEBwQUOcAsTwB1oC8ieBBvD3O5BK+ZfzfzTcDpxC
HyqVQ1Vg9pEVfD+rbvqfJ52fkalMUy6AYcc+KI3eEvahs5q8cs26OCAoZw99
GzrO9knnCCnzGJDIE25h3Do8VePFjF99F2U5vp/CxKjAScXDeLgf4nnwQzev
cViGOZ3JMyUWUDo95QJVz+FxbLnoxo8KeKIAINWfTUEEot1yxu5ICS04GXqQ
QBF++X0eMjT7iJkiOXqrnBnvmIfzTjFVNJwTsWoMaAilqj7nPOakLHcULC4b
v5xpf8FqFs1gCFCTum/Q0lUkySAk9XQH46J1zGsq4Qz2nbLbdgRYzvitTt1r
WLGF0PO//35PBgkYwNb+K0GNsMhwKB0P9k3xMTYkRMgTYg1198eQXK3Pfz8L
mHk/RD+M1Vp1i6+4uDc0FKoC8ESCAXUE/McK6rAVaPsAfhvusrkIjuOvdxAn
bpgobu0Z7xR/S9C6qXDmmJbSyChvkNaxCq3PsTp29e1feFoxyffwN0+0F3At
YIOk5PmT5GKdgeDpQekabbBJ6Q7eqZUszwZkmubO2zLXpCyD9KjYvL7Uvs+/
nEFiVFvO3dbnG1mz6XEq+FjResCzobBVDiMHZl2a05Xkfqv0lZ6JyvG545Zw
wLP82qyKI97EC7dhUCAl4qdRUO3A3II5Pt1DmrXSiALSqtT77E1OlMCkWiEd
tKEaRK7VCihVFl+VrbAlCiSPBX5trj/82EBrw+Swi78IVmWIE7qs/8IZG2jJ
Pmqq7k3QLFL+JhB2izzGsUv1sxm/UPwTFfV2Kj8G4WmKHOv+CmAo5gxJLCpT
Gfa/WKuep5CX9cZ89m2hc5KBDtJCDJpurupinLMNNh4MRFgvJ8Pi+qJkzMbu
2q5dgVV4UHhIA1kvzn7RaE1YS2dihyeBJ7+RorCsM+C0H1PsvQrfIQveb9dM
8y9t5JHwuDgFhhEm/7I/VYqZISG5Bo0QPeQOavjumO3waI5zzdZhj+z1v2Y0
Fdl1A3g197nv2f8aoLcvpUxAeDxarrUNLHmjGZIHxUdfDWOnHcQD/NnDNmmw
0pyu/X6ZkQDvkGXtN5j4AIiZq16hIIc3G1lqjIR4l2feyEP6nGWdnULLslca
jK6kllqmErbH77L0SX/w2oaQIaDmHTPidGvQps3KgA5dkTwjmpWJK0LaUjIS
C1Gr88AW3J5HUasSlnE7RHSrTpel/pSOa9M5LtBIcRV5+RJSA443NZUcQxXp
Y7Kc3pYcCFytgRzxMcz1C17ad8ddOHJYkKKFquZfaruaUlDf1lSRpt1bAXRZ
CJvNJZix9o07QnLkqHnaRtsOjiKeQHtwiihsmRUfNykaJverOdA5WiV3oyBK
/ZQ8FOgMn1e6gxtrLIwg8dbb5Aih1sBQmD+44M3Mjr8YsFH3lJcdOe3icbTc
4mgShag9TpcY6CjzSj0q5SLFOm9WIJXrX8PzR3qhoGlSFwp+v+HtGBlX/XV9
YlkDRo0ObDI9XaXR9fP90wsjIQOhS50uqMHW9qcA3mSyJc6re4WJNvhsyI9j
i0R+ZDfuc329BvYcz//cN1O3Ns4bwhPiWqbs5dv6Dz0cShM2FdCL8bRt4FRj
WHpjSf+sAqrQqtWYKHfrMwt4+SamCmttkZgQI/ifTM+eGrJ2PRguY0nKLbFc
pwXOURe+UptgrFe+xoGLUTT/4XtI3h/t2VjHEGR0LpT3XEKYnmIZf/K3W337
slaXu/Imq7LGHzWjCHNTa5bnNK+BHpXU0LybxVL3Gd8pTYcoRkTKI3RvJ+V2
JQOke//e2XWxEM2OJE8N0RABBavhcZMqY6CArS/LPyaTFHmXrPCMIG5nIUwK
CbUthJwtEtg9KQJiplVNJv8ZzaMhzeYQq6qAsK3Dpar9HPbq9yku2+/l9UFK
dH8ywhQuo3z7ArZWOAQm3F+dWRhOIGBK979+u/tFoX9HAYOcK8oBXjH5NrBP
5JmopdD6ZW+Ln+epfe7fg/CikaFPG5kzBWj6ajff3rCIUp6ZAMZ0bgzqVJ6A
pfSOBQeGcGVxXSp5vAkcNfDWSQ3nuFZEoCh8SVggGs4No+U26AvZLokmSCkT
bzTRICVMOVCkNFN0DjWaHCJ78zmWg4myG63HQPTxhvIrVyTC4lmyNiRsNz/J
y2vod64IbZeHwaLRm5FusVi4f36xuR0Oj06VLCT/GBMNMHWhf0HKkZODtzuc
0NItoU0VCiFyM/UlzGz+r00ez4LQvqYFG3HQCpkaQeyBEFP47M9M9nxgO7MO
8v/ECiSAtLdg1KqHHCx24lelum8Eq2ej/hhJQvdt4YTViXaN2+tyDmbDBcgh
3gSTAIlAPOP+pQaXt3fqLjx1WpurixUY3Jz/4htHfTRLIA4KGi8NbSRtbARs
IkuZqdmmkCtpZxWQTsr53ZzuztaxpD0GUHQTPXJwbepHzA3Lgedib5iiC2Bp
FtfKsMu71yD6NA2XjNvbpQA9O5iPIeYqzFzq0H2Tf4HDUzcc4AnVjVs67Vix
PCE/H0Rxp+f3lTApyhQ8CUh/OWCqapLQAHprs880xAXLjB9i8KUEoYcDKOep
Cu3/vFkbtELfX24XjrE9MNgb3JNgTgrxU86VQSEvIL31pemLRtJPxpFhgr4Z
Oir99d7LdsTAz88hP8ATSfHjLD2iePlR+RmqFktouDBY6hDH9m69tCbAevZN
1kJFNxJGTj+7oBRhFZhFuEMB5cPPIPVjd86vaXVm2z26dPISQgazqKQ1XsKu
5MhLpFNT07NormupZLWDSJwrD8VlyDupozxdds2SnInIOUHtXRg5JnYmGOOT
rWyoVJMkbw16bC4mr00hrIsBSEHDd918NYkkIZdoyEj1gC17O9HH2T1HqvoU
01TFkE9laGGeFvNl8+5OBJgp9HJ6dVSctGUK2Z7f1uOctop8WQf2OdQH+P4E
Z3DualZag7/u5b/BkuZO/q4j3XFgxW6FGuQmEgWcc1gCVzFx1/0WcBQZa9ZX
H2vtvaWA6YAwGETt4oNxn/AORB8Nv5q5N4LF834UkLReZMh3C2HV/VR7UMCl
y2K7L6d2Rffr9LJPqBROjpwyPbdtNx8y2+vPxtn+CKrC0iFmn11dIRO856oV
OXexdpOGBOaWIfn2so1QpOC5LM0NlS/kcwNU2KwB8tRC+K/xWbCGaWZQku2M
8hilgFsKw2hFyjZI8gm0FaoBNRwNsiZGIL3B6x3AsspIvPo7glkaarNMGEWT
1V4NeH6k0KhrC4sZY3alXl7oLGrq7Esns2xjmBMllgKV5rXsTcNvM/R0cWWC
3xhTq8K1UNpqzNs0rbFto+Bqg+fvj7peFi5Rlbc76h1rj2BboUUwjoN6WYkh
dpZoCkSVf3qZdetCfmMlnGZ5o+YE+uo6BOb+yewNPxbas6mrJcEmCpB+D5dH
z5IZ0aXDpQKpVlmuXBOqK69g8X73BY6WEk6/usliwxsHCGxKPU4jB7pE32w+
VJFU1Y30rWpnjv0F6wmJOiTYA392yUvT01H9ucLkxtacroPh9bPxYXRxdXQ+
AVtbvsVyHpJuui3UXhjjh9wujNl6acccd7FbNFzvgHrb5NloKa3BQUYmgphG
rha/4zJQuuwFUQvF3g03ZeDz5hBzlPZyHqfzDpuoqGkPX5LYEDcVDXcANgEO
ska/WuPM32KLFshArFuCjk1R8XMUzXhyw9m3m/ymqsU/3OitA5tkIdKZZXJK
rtajvGHP6xs/Uwu9ZdXGqxK0j4BxBHwlCSA7ip9mDe3zSmkoxUxRow0NpugF
PuPHxm2VeHxhADNT4pbML4lvJSpIz4XeqddZtcJneC5vaJ5KOXRgV23mzn+n
KB80+Mlsl+4+bTjBmByAYEnFzXexcPkIIS1SFuHM1nXKgB2RmF2svpxaiWje
qtxTcKZCsEvzcUqCJNlFNpE0Fe5f39XK2F0cm5Dos86AUlhC+HSnNdzg5jVC
I/Ayj6mpgQfjKdCrY/eVqfnA4BSvyOmVrDkPeVlhkdTdat9nJP8dvvWJbXPk
w+w0lnNkpAkLiLhIZdsYCJTg0KMb59eOL8O/EJA830vbmAUfbVOp6IVmVJT4
rnBZwSE65WfryIML84KVlPw1/JY0EaTEOH9EzZ+MM79XJZYr1CmuwR+bs9vh
30PED+y4brKwTpOhbBOGgu8P0XX/WAiCETGpx8ZibmRMJmpSKWlTd42AOUGC
4u/tfFun7iwLkHcPAHYSddTTJSwasA/qwT6KDN7qVVSG89Gfy/MpiG6+Ii3Y
d3biINJi5tthIprMVlfZrAy4eLEqa6aSoH3hJEp4MJh4Z6JpKcbu2aGr+ynL
p/C2awXwnGOSoQpEN6Dstg0A362O0qpkklm/2Py0dTZYVlAVmOHwKOPoaKlg
NLK/X/a+/JwZCTHpTVAWQMm/VDtye5177hEWDpS7aFT4RLH47u0Dl/jCrYiq
CZrolvyenZQl/smitBYvZlCKVF4oSUFKF+M6Lqsvead8tfGWDCy7iWeqB+7p
98nZIywuaNXrh7D5zf7XARIcs/CJslImSJUbPt3VJ4y7tjyfya+1GbPPXA1I
fzf1dsc01YM8J7t+B9saJy70JFQvUUetriMTc11r37VFxPKgGW7PQ/X7AQip
wt8ClpaQ7wEMVXwmR+xPgG75lkdfZyXr7YShgm5c5q0AmKnc9Ai4HLsy43jg
IAdQS1W4dt0R3hE42fsDuU1eFzKwZlYMtptu8ImwnB/waXPMglo/abEqi4rx
us+nZze7t0+nsxySIT94PcDUqJ1PBsinV3Kwq22vFdOmDOaJ6rn7ftvdNYOH
nwbo1LVKr9Dk2sKMu+vGv7BVcrQhR8VTcdbDZrQfBB9gYyLNWzYewVpOeZbr
8WvYJEDABTTOq1LoF8a3LwEm99ulo0+fs1U9/v6DMFkmq3ANH0op349qvgFv
INhNB0dhSQ8CW7K++etqHV9qvY5vHyrDyh/djotXtp8ds0/16rCi4Aahq8UO
i3AdggpN8+yBdV4dePbqVWf1LDoU7U7vgUJtBngijxsp/KOE8JdZvH8viwx3
FDdfSM932N8Mly8bGEaMmJXvl45Kpj7TbbPL+zjovLhbkr71YdaSsPE4/pgK
SQJaTmg7zgHPwU1NZ6E6cYHNJOPKyw7XnchjyNpiGmve1zv7BHPQgxtvaAWz
pSm2HmwWz6Aa636GAzFdYGb8+Lxrey2gB59uhZRMMKt6wp+Oti63v47AZh7b
pWcdF1XHsUJKe9ZpsaCrhqJEhSvM3nHJU7JtSdCa/DRTDrHonBS0AY+AfPZf
HUuPDcDkVNQFAhpRM4nAyfG2Er0Lsv5WmaBYBorxnQhkfoy+1N1aBn20wO84
AxKtIhQqWLBPZsz5PtVWii2tp5j5K03yYQNcO5rvT9T1DyAOnLpZEYQGLRLl
P1C0rzj06sOYHHmP6SQQA4KngFKZlMHHdq5PKzsEjUinbI6Ilfjfp5q+oVZd
tAqs0O/Vr1N5u6go+OUg2q8akesf9hsGj1Hl2wLOjdcuwBmiKwFKm0IQQmXC
NRqzguu9vhxCFOCxRcX//qCteTvgvKhzIn90DVN37OXNeCLZnNz02deU0tnv
q3cNDLzDuU9gVo2IF2oDw6M3CvdxaylEh4eHxJWLrtfzTuIsoFWXihWSKSoG
7+VrifA8gTj/WexgAkHtjmkbZ+H965F3wTTd3fqcalnJEtd5cpI5HMD1CZGx
wPOapCIG0cI73X3FHQCHzn5xOnXldJtI6oO8DZD9pDqGJtrQhelyMe90WWQk
PqjD8lH0yM8vuipsdnwn9N8ycvubVh09hUv6ig9v0mkjf85YUL7B61Hzbg1k
TJPj/N/eaH4pAzrNHyiaShMYWhTjOO5AO/2GQqLoWkaf+sosGbw7AeTqWRp4
lxrdnc1l4Jb1pfvMe9XBC01Z5gf8jgS7ctlBs1aR3Impi4HN9IF0Fk0m/vAo
biunXZ5/1r83Jj2KbYClnD7t9t2epWWRNMROnylXubebxU3ruGIOannkloM7
aQDAI8OiqEkws1Xpmx/j031K1J45aCLPpha///EFRLKWVIfLrrU8fja3Sjih
31B5G/wJz8y6oLJI+gcnqfzxTqPHVH+am4iuSx0G1x/OeYV5Tnb3ESXEdh0e
y5MktNTammRSRoU1FoQocqjVWP+nRL+5pbi4NGLFUasaNNwu+G2StL4T7P+E
uEWXFqeuY8CcpB9BZcmkhbEu/gl4FJCP1zNZw7iQEmLCeTpS8BJsc+BNGXSq
XfcBIua9MgQOhcvJnoGMmLRTaRkLuY2mw8lbh/eFHaEWQAQBvCM1JFwxAzYM
ZUGk2hkrJeXiXOtFDU+z/R3DSTvHpurcF6KMWOypVT6SNGq9+zveOG2Shyuh
Oe/lZMOAs5odOGUbbdEGnCLnlPEm1YoVu/hadMikTmlX5i98+d6lxQK22zF5
WmsRMDQmXWOjc0T5V/XtJq5fK61zmmYTmD2WUdBqrMg2p2uGrBC99VWPZbUt
adBq0/89QC9OtooqKmpsEfoxBxaL0UN2o1+oSJiR2PlSDVXOhajsMDzMM4rp
S42Etz6bqno/mA/FbUFCCFwmR50FeS/pgTXYLELS8VBWLJq1v0xaMhCVTvdG
6ppjzMNujeMDd7kdYfqpQIQGktnbW0fHtzvQpw5Xfjg7bFHkYQjzF+/1pyrr
gpirLwg0FYftJc9zz0qR38F267hnQw45qR43VSomwyY1Pgta6HO4/LD7iT3J
3IT36CehiKlXP3ov6sDjqyPvqqfmmeObyd2325hiMnKc4TAjhWMrvxJC5bK4
S648AepKxihqi4+/RBHbJ5tc+qNl3/nbMG0Qz/Ygsl0LgmF1dt8YQwy0+NRt
eGYDj1H2nOurP8+GA/m1PwyfF40whoy2W4SstgphBkDyd1vRNhVD/XhM8mR+
0Y2Og/lJuWU3FuQC7P4BlwMnjuk9Mms8h0hBckGSG12V/T+h+DENib2WPCTg
pGkk391IhCpwCF0BlvBuQfsHAHBIwOgIGcbQf4HmZSkUCmC80eUZ4x+BEoaI
X18rNkllcybBoNPmSPG9HUbjXVWaqY4dPdCrwzIHc6IgwW8NxoOp2fAWzILH
9/vazfRiaXMg9EMENCIxjeSVsSc/sUZBeFO6Gqy+kGuQuWTrqsN63mXXg0LD
lzq7XcLvoONJfZPdsOg2DXn0ewIjy3a9UQiNjEvYtcWVHTdbGn0YddStEzN0
P4lnH1iObHHPqCu/0tHSPvC4DwEReUow0eDWOmaw6hraL/7mGVEB9y0n1INp
yGjIjH7v4TCRerFDDUpDYhW32qe7RQ8o0g8zJoabE3Rxop5a+en5JC7hi9XD
9XUrzIklpAB8w5M4g90mUAwPIERv+LOWYEzXJVi8clsbEzcdZXxQhTfkbhu5
lq2me9WNzcxEfGBoAi0p0wvQnPo/ebJZjhwQXw4h8pC0oT78bGwioJZxRNlo
ho0JI5/4OIZBI0mhBz3oTYuCD2DmMAzX2to81SZEyfEPQF53pd9y+J6F2KDw
Ki2te0oUAgBgdo/Q74hcwocPp5YluBOtwVEibOzVXREQwW16VqqlND/lqHp6
RjbMU2VsxTHwzv+HbppKV1EtUI6syiUQ3ipRuH7jyvv9bejTxYSDb5MaA40z
PwyDqg0xPfKuBBztsu45r5eyM+uTorijbRusKVvEr4vpcV336S+r20JS6LUp
nE27y7nFOknQ3gZHYvXfwRDT8tBUZ0ZdFpkVl3ODlBklWXpJxvzaNUOmybp9
uSO1g3RWKCLEc4mGoHNotTi6PZXA8J41QivqHHMyyOSZ+z+CDaDSZ5G1catx
7vqxcKFsmeceAWYuUWedcr5fo+E0kcjWGOxesXkhu8AswMMLPPzrzIna2DLo
6F7p738yZKPfRNkAFQJp+U3ert+xDYiwFaar1gLPeU8ecWi2wzrqqGCSbyqE
s0Zb5ipLNBl5F7bCR3DpoRlshiu15fVEisVetpv0ZaRN3ZkeJg716hsVgI1w
sjDANAfXATMewao0mZDcjJzyGDy+duEDvBkVglaIrsrRlRai4k3AQEVoKjUC
QdiAwAqmnBOmkaZ/yMJJO057SN2zMJW9QK3bVJcq5NyaMFKRU3LwW9J7AeC4
EufVRcnnPSAav7EpqWSDsG5BUGnGBmFGv6ZZQWtGoJKJsicNyaACv+oOj2zW
br9DjtKaCwceKwrQFvXGaR9mT6BN2I1vnAGbDhj8l1W0UsgYKOdsrxwc6Uf3
UEEt/OOkQrPIDoeP5TDa+NpTUdSzYaJn+LBdWL4G/Mfha3rqRzsjnjQhjx3y
DXY1M8Tr9/SwjyrZs+ygI96M3cjDAOnFIBii0j7LOG1zPazlnaKeifEoIuJm
nB7+ULcp2eH3KQQzZSWV0h77smBNe28TG+RAvlXjdlDycGzW7V6tYi+OAdLd
p3CO3zqe6BtOB71U8bZgurkxxJgGGV3Zh1xGIyyziyknEwJYK80z7QVXGMq2
c93YXZnkIRJpA3hXJ//ECt+OjIy6evXwyDY1QS8NePaxo1Jv/s/JIS3MO8FG
ZgahWFeLSBaRLD+YfwDScCP6qASfcus7rm1W/SJh0hcrHRocPve5p8eDOcqc
VspARGIvOkDNSKXngA/xfzH3+JDRehhxEYBY5r85jpcj5dKTkuj5tx4aVMg1
oDDG7znNEF40KssIaoaonKfZPRbXD+IbBrUuDQausXpMkwVV/aCBwgSkF0K6
0arhFWRiA6DjjFAu7+yhhNBAUS7agvu9pvbDI6WB4PcJ3E3wIPR3Q1OUlEwx
HEBXHOnQjPVCe8L569dH4RjmUJyRvFeI/D0ic+ymRiaFTlvBo/d2zB+y9VFb
R61SlPDzrf02tHplqDTJF3yvLbOXbx6+mL4j1ztnTL0EEmzv0h8BRPPsoM8O
KWKO39elri2KTtf7mBakuZZcqtN6IeN1RKniMwuZ6vqy4pjvK4SDzA2T+Uww
FlDj5JS3sEhtbDHXpLnSnzSZUTIijr8SwfU6aVDRusspvIlVmYjnMjgpv+I+
rHtzSQ591/GrwLRd/SnVAQdx46YlZM52QEGZZQfhzJ/UVLdLnx2uQJ3YV5a0
R+kfqpBTgh1Lcb9u9dwWweUX39+DUZn1oRK1/5EVf6ArXjlJUDdD4sfuZOS8
XvYLijY8WIecW7o8atFjYF6Zg9YOrVf+LzOjpAddH6crNAWsRreKaRHHQBCS
k/zaYR9AGe6H7pvwuRSE4Y92aPh0ug2GvKhlOHkLfqg4ilcl0ThuZ7plmTlW
R6S9F0o6rgdeoXtsx6EO+2XLwn9ZPqLnslkXat4RAZtC1eXAfZ6uRTeRyqDf
cX4ZPZKVSAVBUTn5lRtC89SulccxinCLoYf8TvAWrqNZ9HKpgkXgAuj4QHsV
ItLaxQeyh3zlP5bttmtXcHl3KlB1m1Dp+zEZKkdw4vQU5IJVRoa762px+fxM
SwwA9LdUYOAqS2UFsoq7l7nzAxtahdM9p0OH666xAwy5RjUlrHb0HQGeB+Rz
2Tku0J+SQxLI5YX8yp79db6z7gWmULI2wWMxAtYer3gI9TnSTbdg0U1h3r6J
mX5h77pb79vbfrIzG6PCJ7hZI46uoNfo3FL+3xtmbxxv4O0uJUkWxny3PfAM
6TNgCsiuYTIP23bajxg5FjcSiNc1d3uZfQLhJQ7KI5yrkb9W7tk23oUYtqwD
FxUGV0bdCBFL7tJfCRrAssEBxs5pnGzgTpF77uQD8S1XXydH4QqVffF3fnWP
kFbkGoxk22CeG4AQKVnh+KKL8WpXGFpkfTkLnSCznaSmVrJEoCBm3vMUTZtW
Thels6+PgUWhSh/kAYpOCAYwLaG3WerlbOJGkJJde1GiXRuaWLBjdL3Tss3/
3yX8y28G39if/52hlA6Wwk3PZm5erScvxni7S+QKSSp271iAaZpRH40At9/b
MRKw5B/Fd4Rq3fbEgF2S/iIhaXlJrAO2I97xHr42XXytyfEfR6i+hko8JN1j
efO0l3GvGDWLoGPOVLXT6WR8NBEy2Jcf4q/H5zVrP8BoG+TbSXqpYGGrAr7A
NYdbHlH1QvHlR5Iz/TRcMXJ0qR7GLELTxqTqGLlaubnQ6fk5G2EdvRCtddir
+XEVLMGNRb7YDomsCvaGsIpatXW8MMu7OU1868D3gpGtFxlPv/v/j+VpV0St
VIorCLOblcuAMw/E0tiTxAb4zHkNvbcrH0UkGz++DjW0yt3tpe7gIAzl0cjS
8O4ASRf30YVXAFj0nfQ037dghma0osNXDYzI0MmGfoVx+Q8NmhwoPZdjvmNq
LGeJAYNxA8YSrn1Xs/2GLb2zNRk7nUa3FgOADVuzqoJBqyKzOszlO0RjDn0J
6fYw4+O4+NfLejEzSuneeBQ5/9gMfzCO+575qHgjNZ7k9pOjnEVmNhZ3DSzZ
i4jFctuH2+em+FXXrPz4CN9EKnISbI1B8KR7P5Jp53LLrKPkr/cWB5/rBxbs
3JCfqp8lNxReWNVu7xvF2cJP7KaDEh7qOLIrYb3XrfPInVwj8RADjRnuc98r
Iu3oVIReOhADdxkH95wN9Z/d2nanannNXYLfah93Ccf7WiwdbMsUzN5OMSTD
oNOEwhIzrDj4OofdxZs0Fkb6fIt95bYwtrk0hz+cOj8jbmNVCoKGYXzKv7p9
eiXxR8vi/DXQKRH2NP8qsrDRwvh6oCEr/LF/y2Meoxite1PUWuUt0GMTlpjM
5C/JFIWL0aU9TL38C0qNp6uAnUeA0ERmApc3h8952w43BQ0/nHQ2GFMUq12r
3jCSdzGc9WTQmSEI8PRx3nwMvMuvEyPSiiLXR+5WgnNTO1i5IGb6beBb9RVc
FL3gWOvjow1QG3kfS8NUn90dxM0J3LrM5g2q/j8P9BtLuvIyF1JGl7Jh/+FG
9oKiIEutDkE2GmAYdlMsEP+UMdFBGQej4q1uv83bfgssq3Z9UIQJTjzf7yrY
AmASHG1qh/9IdQD/14izp7BNGCZqJ+9JXKD1m6+xizvvUKuIN6oRl+9AGlZS
kefRJhKnNmITV7/RnWAfvyFvKPA5OCvQUATpO9Bx1y3DCK24Z72UzwI8nWmq
omAKG6XFtpL/8WQ1Cc1ivPVv3JA3KACDr5NCQE5gxabj41gvYNbWhvhnHOIR
r/6199BNJ0pfJcUZCW6ZZz7smcDCI9Kx2Q1udEUT7az8pjRLnZAdbcGGI8dk
5zd6IYsOuXohJGOSMaFnL4wOdEZqQekF8ifUDxSJBkAh48Btts1YLhsAMYnw
p61X/oAUS6sFgp6qE9XnoUbUPqPVle4GVaNY6iVCv2bM89MB/WQK/Ar5TdZG
gCe1BRNPi0ZM+hk4XVdc8HkRi5dMZu7b0tD7aDf3AaLuSzB85VMmeTnVbqU3
WQuZVKML9UhF+O1dSserUqBEg4G66Pz7LEC9bzwboG/gk4yTJt/w152iMJHF
5eU1vj1aEhIL2uD6K0+tY/4uUEt5aJsm78iwMF0H/Jgc6LmS9qB4OJ2nwVXL
Jp4W6EKxssrBAvOKQfoPww2MLR1uD9AYo3yGyDksgejEga4K1HJ81mrKqy/3
Hkr8mTOsmB7JBcBvYmN9XIJeUNal8Rf1FnHUg4IukJHXQ0R4EpOYNCAqRTeb
dvM2I7s4yNX/HpIoomjamVk234bY7NBflglaAOCyaP2BeSLrcA9Ytyw+33wb
Wgwl+xqI700qeh+LItajiLLKZX5BFoVsYOx/D0WE2LlTVM9Qy/GPkA2+0dOk
AfehebA/HViU7o1pPcTZcK/wgaItzkF4I7hqyORib7KPrIo8jZqs3l5s4QRo
W7wWiYxnJJQVGxFTqF1658/hhO6mP3B+2T4cFmz9U3rLSUSK6UGlu3R+j27V
PAwDUnkEskr2h1M8MdTRmU3UDYd6Y+Elfm34CApdvMXf8xQktMkl2cAExsP2
ak2n/bBhfT3DNk11YRNQ9U5Q2l6rkPEoztYvrzjo6USRPIhlBmbulS5vVJnP
IdZykjHuyqLB1abOIdhCKvXoKGylyHY4KLQNpOWItejfZIjf/Zki6pXqM9H1
Oru8xCsYTD4Dm/RhztGTOa7KjbmmPWaDIvvFDWZiSRagxCSabFDcBAM2bVJh
YiBP43GdAnzO6bbFtJ1TEFrXLtN9+XE7y9W6cEqrUvSE1jwwHRF3cD62YMeT
8c1+Dch5y4hP+bG+NLqFHTCo0Mx7zMZjF/HWBsqWkT3t+CmFh3gEOscRCs1/
QtqqBcD76SJTTh+sBFdYxxkngD47fe7EHDnEHqWD8bXC4exAh5preyHrn3F3
HWGzMxJFFQVpLO5bv4rP36wsD65rVvwHJ05+XmV3ZZvlGDELMtVvCP4RF4Oj
Rn0+tYdxM7XDDohE3XhVWSBLHnL7oJCtayHr5CtedAYs+cbAjyqBYI4XrNlg
YLprT7KI/xn7yqrPWlsyF6KufnU7/E6Jj4/DrvgWXXCC8+f830JpoQKi2uzt
GolDsOCAVLNZWjS0aPA3IeZOlsFdfnBrOfGSItDEzeUmzVri7+TcIqOU6T2D
FSJMFwcbsGWs9H2qyo9BGdc6eY5j2rSRuJmRlcVhceCuwyNGTZmwYaa4m8Jd
aQUUUP0mPW+/TnB+Nay8ge3XcMsN2TPxF60xukmVyXwZOrmkaaXCMknPfktu
dS89rk+yF3hXzzwfb43/5qh8vYjF2xGg2pdm9cASo4dQ/f5WDChWJMxOgQT2
zynQ12x+UnJ4F1PyHcWfClv6MCmx+VjY4YAQUjOviTvMg1M7IERKU2q3KT0v
WWWuwK3y0LG1Li15XR0FbwShTn/YZkAZwdEqrxeDM5BmsYnoatI0Fz6gXXGl
YgUImA9TvP2WrKKnZ/gAzrXSqlNIL3ECVerCdIxDZZPaekxRjUH8js4+/mkR
FVgMGNRUWK4jsYFFU2PorRFtD+HO6Zk1u12dNddo1hHHDTjHf/fCdhe+5Csd
5KRqYDv20N/M4z5EREIZdgAEwSAXvQMhfhhwIfXejep0omfcO7MyL7QgFlaV
2xNO9cHQCCF1waHzSAPzGYpqothEZfODjIlYevSVFdtisjkh3QRxXlsGPsTY
3m3sZysFAuv+mJZWwX9vjQFPCfDdBCqqSBaduMdy+qV2NtRDunUIOvjKgVSP
oQv9S7qsAdx9sz/AOGY1RzEgUzslfWaY1y0b8F9n4Kf/dCcLXIf7kb9+ET2+
b0mTBAlp0czYvnclImL9evilnxUnGODFbzL+I6hm+jzb80rq2KYJP1ssd5zd
pW+v/x/NBOGmtpg7hdfgyI7yet8u4YOOeDN61+BgP/JMdrqeg3MIO1l4eLj/
xbiD5m02yRe3szJAYTJ3nRQJSaNjYKMbgsjeHbXDJIYwB1Xso9zs7O96x/Bb
rKlYe7eLSJb1tqko3S/88Q9r1NFywhQLvz1RC5D6fNlKG+RopZ+tmY14U+XA
jvlPjppAwooa1ngGOIySJNzXe47KPDJ7lRPx1gmlTuFfl8bUtPhPe7y4m3x2
4DPb18QqgFC8slCzlo1KDQm5TCftQC65tsC0RIQRAYDtOr6nNboCBDZVM/G5
DydYXn+cM0GntutxDZnz+4V8k2iMMOri68xMA5QYFSXnASiLkKqea9F05rlq
+xoqeu++/vB5uPYsXD/RvZ7mKCB7TjWi5u2wLt0vYtnOAg9yRpsSIYkYd2gu
6eQ0fvEZbqxLip1G60J8mo4RNrL9M+mLGAx3MkerPCQGK0v81V1Kwexvx9Mc
nq995MkHcwtZeNeMRmheMpETaffIuo7TWEEb7Ggh7S5/MPICXGSpho8VG9u0
hSRIkeGFwiQt5/j9OiHTOPyZG84khD6RTGAPv5qqjIQT7ztMYImx54/zZN/q
lOXZHMc5ZCmXiiL0Ou6FW5n/2MhLtS60GPkejJrWq3Ikk+Oyjga4alXU7Rgt
kRe58nIW0/YAwLoChl3PaivaDt56kgXdTZaYtsq9zgidKDKkicOFp4+eUbsR
Et0lrtoHjzU10+19DoT92LXgS7V0TvZLbprOecxPLuxPvIF4HG5G9v0ti1tz
bCV/Gh2ZAmZpvb41lQBkb/7qY+1FVFQsm8eu+bXvChs5uI1SqbB7EUqdQPuu
lJWRNA6Pqqjk69NFnqxshJHqheAbATpwvuxGH/L59cv4VjFWbjGi64kRarmP
dWa37IjOAYHCpol2adGJvbilEKGRSt///ZImdNClT9qX3WYVgZm9I50ZodFg
lC+eO5yowo7Ad8vshumPSa8/ZiumLrK53CuElXYeLFQcaDDvBUOldOTxbfY8
riWyR0weZ1eia+MmNx2xsktHwooG4wmOuZGrKUA1chHpmZZNCiu4FioUwC/E
5EHz7qlm3sQz2f8Rgf2tTa9DO/xLK+y71dRCZQiqxSfT8rNa3Q80A9T35/E2
rgfDbbCq6hUgTSM3xq31gxb8YKsQXYk4h4g+9bmR1eEuNoVdbA1EWFrNCYwK
VlZUNpygXLlAHi15iG1pQZ4/06FqKSlEdis+TOlgVMD9iasRlxZCBKspM4/k
+zRrv5bv4hXT9OdWSzWduly6K5uJ3wiH1wSFP1w4nTgHcpPeSwegHCZfSVQK
KKn5I5aXosQK++9rg4LUDZ9/ZMhBMXegng5O0zGe8nXZnrYt/DxNIzgVKB9Q
LYnscwKXWhNsZzw7OYx5Ogm2mkzh3Kp1fNO6TfH9GwVuRmG4UKV7Qy80QCXA
Vpe9Bug105ZgBAzSPuTOmDdhND+1uFAyCagMDotjXQpdAF9bfjktm2o1cbQD
3v3t4MEZ3M1AL99+cPcdbEJDaS4x+oDlffYTHq5vpJ6oJ/P9ES2hf4j2pWT/
qI5Q6qbUM0nKyk6s/0ApP6++0xaLqD98VLuNsVy8zP32HtMuvYHh9PNRNdEn
Nb/QDX5JFPnh5YADD7nf036iTiJ8k0YJ9Y6gCnor2NLSb26jnZ+GVoxriHiK
OQoGsBsWubePEO+hOpoYYOFRuZNAsJ5WQG0dNgWyP8NoLFVcxsCBwNrm2RJ+
8ecd+qGq0WQakm39JPrqpFw5MaZITXguRgz3DQC9p2tNEMIM7PjLl1oivXLC
KBoP1Yd1gyOS71ofl92+9NvFi8074gaZNEX0qn4vmAEoHBXooFGraEuOCoyB
jOFCRFs+9IGUKWkPMuofOHV1HZIbiX77VaQJT1bHw520+gUglj+xUg9PP7OL
mschQaYlcXDVOE1aFo90GS3wygMyHXhlaIhUyEKhnMnxK3uPc1K9/LhG3nzq
fCzd+g3AXcWnfw6YbclbAEsy0kI9LBAB/QFLnV42UmHCzM0E1/0X9C0dy0r+
Qp2W0l5LCZvovYD0dDeBPGD2HOYQbOyQOfg4q0vyd5k54ZQuMAwZmDVwZZxX
TtsNfBznNlAQVkyOS/MV+hFSeYZPcJQOKvc/8Gd0RiFnVS+5dRPtOKOLuQGN
kiUA+rInSTpmYKCj6TJUkL9Lp50NownKxPEPayT7AQcpsV2SQGZg3Vs3dJP3
XGV8Hrz60ME1FRqNy7mrCK0MRMBIjF1SaQwxVUFJ5svBPRsEI46ZF67m93eO
wZF01V9Qs//j7MK8kdql2VhONCCFFUOvdnmIIdeNLqkhybdUcMuszRR7yPrj
UjCdGaNo0PAr5N/emEYdcxPD4HrGYDXmSTK+UkWI1+XiiKZ5TAakiCurRPx6
slX4mENrBIoGjm4sh9uZlhH7ddicVKfbBIHPC3NoNsyymjwwcvBgXSFglX4l
2XtmYAytPLJZsZ0WfqW2l2m+TTcQIvqU958v87qLSK57lVR9+uBXU/1PZWE0
DccqYqoHo1E9bHVPU2z1BjGx/GqSmS5MQ226TjcUl+LW/G+nmdQjU9uZFSlu
0/Mmy5Ms5LUkRgMMWRvMB1c9HUzvsCe9UvjGDUmX3OdE0LFj5JstuRGLTO3V
8istHPO9kvJ1hUvXNyidp1JRR0K50G5By/uIKAxOBSawwViL2YadSUaE9hs5
x7oyUYot+VxvYW06TcpUeGChmRRUD63JtIQUXkZO1h5IQSs3ojZwcantao4I
HuLRrVWWPNAfrmNmIRiApNf4X2OdmHrzkf0Sh2wGdlAbZfy+Za5mjXrlbWYU
w1fVhG77SlW/EDXDq2fzF130kWAi34vTLSHQsHtUIQgoGvzufagFH8Edg5u5
eA6fG8HFHG6kLsw1M73w6ZOxYPrSs6UqIvyh3DfhRM+o7/HvaWgQu2FngxxQ
xqleIRzJcuJPZmZYX/ekO+WZO2WLHRZFR6etVddIy92n6p/pC44qkyzF0tYq
KNrkV964GHBISkRhm0hAFagSHwBA4xMo3+yXxm14ZnIPOPiBJWUQbMOYRuUs
+ZlH6FQwx13hWfz+ejo+2mwMR0STWyvnh/mrUSj+zZ+k51c6Dh1CGtIGtlaE
4e+hwME2evhtTDX8veVcsyhBwK/YX124BQ9xN9NsOpX4LEMX+c1DcTOUoJK+
FrT/RiyTCIBP3sqfbRCkyBS0DHDGb+6tVceDTp1laDT9h9Xpzj51slaBwldJ
Qj+7K/ENDKvv87LGpK9zEMr5aZUmH+FR3SwVJkflesVyXWsxxLcp4qxY1WSO
2JslwXhbRfcWJqOa2ODRw1e1fKI8mfr2QoZaO4RRi2g+gyjxqIe4FeYiJpWb
+r83RVfn0FJExnf+mT6AB2QrkzNzXq3kCMurHv+rUu9MN7T6iXbW0UB8V0oC
W1c4fhhcdtk8canEdpaxsvprKhSKv1joWR4kdsFOBn0qp5KMFm1P6g9eRUtn
omB5FjrBbm2ujnosutaVt22DM+vs1vVm0CgX4cA0eClOVw6UDbVO/dVybi2U
jua7fXZxuCddeWuAjHgmJF2FjxMrhTWPQEqxf+RBBAoI4jA2cHq5M+eJ5Q5e
YZQiLQJrREmqYEMZkCgNez2bRQlVeMH+hMQP1sxIRDDKN6fF7c5NequI2ulT
PKf/9xmt96Rxg+CPR/KPLFO1oYeqlwYdNXabNFWk0G0nWWvXXAhCqj7h3gdW
TbJ37W2Edj8CO/v0S+Wzc6gaTSyfhZOYuI1aWAkNTJKF/8zEgOW3ni+FpzzK
rLyZPqGwPIQHAcUxJqdEkZrhohKhlzAP4vYXlZTdK14Jp+7WgX4WGsNG06ub
wHm7mQyZNPJ2ZXjzs4yACBhMHGzShofq6ikELGp15Xvg28OWKSvDISZWoQV/
ISgZSoCAMg5+f7eZ6RGaCS6voQ1ay91JAt4dpEwzibnFkdDzvCjLmDEGkOo0
AYvnlF0ofXMB3Sh/RFomZK+sPCu+VMSuNbREQOpPgPjLFdBYwIN9Ccof+Mn8
qvvbIzqIBL/MUmJ3lu4IAjJx8Nz9bDKwUr8JwQlOhZzdctrGggJ9BuaFAMHw
WOGXGtxwsRz3sCrPCYFeRBa2oVJ2f2E3xhstEc6UmPQCiPmdg2gFd67xpVM7
KUILI5vaWJ6qnALl0HKXQkeymy/BcZqspsg+DaL8D+sGEeWCFXnT7HPRbHEl
Zx1bB5G+mIQ9XeJqZEsdHnKvTW6Y2ay2OurXteDB9P+ZFAbp9lKN8j+de2Y+
W8kUFTS/Sp4PR7452X7521xZJzBO1xoOcsFDVGkCh00f3rKQi+9d5Bgo+3qd
swfKqCfpln1N3kdXnVEFbvFuaxHOGRaxjwNhjqhWtKXcNfX0PIAE1F9lMTG5
93nyHbX4cpLal9QtpJtrXlkhNdtykhV4jErnl7GqcAP16sGSbIedBrqP7ON6
szJW58nw6Rz/i8W18PCttSTue5aqcTpAkALiPc1CucFpAIynqDGCoLxLPmVl
xDh3pYUl8qJ6vRtgkQOcej67pjwp390wE0EsQlBgcrSr4nonvvoJetHK27W3
9gzEnJSylKnVsdFocSwKPHFPcpGnwetcZ2wftKeOCgyD+ByECzf4u7OIN3q8
wZ8OAg1MV0Nrq4AyBVDqz4utUSzH8m6AdB+CY47Zg+3AYSjSNrOtEQvBMs5v
qS8zMehWDFq0se+2ziSpgC6d5VBP2F4TcW7fedtigfnjmLGGV346USpe0568
YoIlbQQGxApoDBmi05gKrNHNGZsPrdWXf/au9GRYpTt8eTR5Ap+DnhhO3O6K
+28iyM3Sv5Dtln/7C1FON8hkP/Zq7h/jlkIA5tLcgKtXpLxpWUGJowCQoY2s
3MY8Q92qrLHPVXA4k4cSGXmcJ0I4tAiUGkw6agMIZtlUHIscivQCwx1AdB1V
MahOYtwpYfYFlc/AbVt58yhO8HU0CccmHQwoFr23V9ElMVj/UIo/Q9K9AtKy
mu0LzSn1kjCpmA65JZEKxz4vxoBXAeL7FOsyh7Ss72h0c7UTx4SpO7hN4SuK
ONzDYykB1OIoA2QVeWFCLMZcZvAVidgk3s+gcY1QrDvwpz1x0/8UNKOaWvbn
JBdU3zNCbO9lQoFm5t6Y5AcvMFNeYrC1fymS5gOiKvmgqP3aZDrzYHZCo/Zl
+KPKZ9BgDyRACB7HGoLX5lH0DuZmib0UBQ/5Z2x0vIkLjZ9oceC8wzfK9fPH
WrQxX99f+QL8vn+tH5W4iwXWOIlqtl+GZk0kW2Yb756spX4FlTKKvKzbhK7S
6tVYkZx63yjFA6MSVdGM0uMnM1v7fGhD8ycfTBEx9iL4Y1CLGoRWSvLKPABa
iGsXtyzMj0/nWYGVLcXdO3wT20wl+hec/Lm1ZvxoB1Zv5902iSfxX3GEZglG
qu+FLQWWmDDzrOR1wgGfI/tCh7aIkwUi/a3TdyPCOZl4YdxZZb2d2/jksjqb
6opv1pi60wbEcZvNqHSOvk0ot/qWPypNAG1gFBYY7C34m1Lh4KBrooNwfurl
ZC6fh27qnO+uGFWD9DLpp8dglaZdfxOvtHNE89d7pSFetY1S2JWTnvtTHpov
TGgH1BFqV3BLcPoH1ZryXJDAz/TXtCiJZL8HMTMSms4VY1M3PbV8PsprAzS8
Hh5jdkQ35F9Tec1Q1XBC+evI5V3kQLGf9rIPF2RhoIyqgFQ+TEdGR4guLapl
dP9Nv+y/5oOLI8Jjb98KJ9TgvdwKL0vqb9nCVHN2+xM5RUApwjybkk87YUM/
NAZpcgKZ9qiJoDkMi1HlokRfP7xkJSoFSqiTzVEt4LM9oyNZ9tMffoBoljoQ
2ctUSY60XV00jHSDd5K3NiEIJjWAQeXJFq0DqpVtCaS0qDv3FhPNxFzOFgXw
fl6SJ+JKG3seoS30nl3nCdWc41mKy1lPL9em+uqnmCduJmrM6h1M99YltAbI
8a6sIjAxm7x1pbiJZcLe7KkxG2AQOCvqRe0II2o0wtaPApqI66K2nwiAXnK3
ArnyGjAbCXs451R2B2L1yz3f46tkh85wfGIycBWiIz5OXhnmSVxL0D9izkRy
aP88WnqRKPgaE5wEAddevZK9vRUpQd9Ja/onB7B/F8bIXGlVJaC09faK245y
uU06CXAcOo7KIgqJ0beoPROqpwPobCmK04ScvS7wduCvZ2JBMynQAetXuhay
ZahBOXhdlviBP2yaZLhfVUo5QaBGTDYadgoAj/5mYlpHUhYdr0xbGLy5DBQn
xpPjOxXPDve6De7PbM16CjMxaf0qIcNXAkRrLF0wDpZeaHxh729VM2j8s3PW
oiNdvz4+D7As2/HDkW8bAacUz00j6K4erf1P62CpTvIZwf7h58yrYmtn1Ldd
14uVneln+V51D/G4WJVQHa4nodCeGI1VOcGw3qGS84Xvb5MT83+Z7tXUpnlH
H9/ATsfBEn+/uTIatNMBaYXcluwQzoBV+uWvYEGz3BBWD1ZaVleXqHPEXLwu
0fi0ihQGbYYifE8UxLrFRVIsUXzOVmV7h9ordmWqz2w4NCBGElNkJGxek4yE
1sMbGY4kDcC0feNlJl4x1f3KqrKc+Ma7YN9GP94ucIE+wmllJymHpAcEe/+W
0M5y5aB5mu8UAb0fpP1yIeUrYVMYplqZzGk3Lx+OE0d7xwEcyp5gRA36YVV9
rQk9xRY6ZcoyyPOTb9UBZ719Bl1O14yL0gV76OpRZ5SQERUAsLcg1cVRdICt
CAiW/dLi0SzvVvrSAAjKxryLVrnEB7rA/DaRIcz/5owZNeN/Cqj22l+dZ++l
FCPcrWsplLcIMOetn1WZhxnkxae3QDfhIpaOrq9g6ZiMZmKoyYcw1xmiAm+i
Z3LTLNd9JP0p/lBpWVqef4Gh1WwQUqfLZnS58NyydM1ZsdnrrqPdxZPayHMd
5fcw0T/OXff5u2eUyjWLOO7nJev8GQ2gOwZ2NLtmXbZjRlhu7x7an35bkjNQ
il7hbHi84DnYcFsjs2NP0DPgR5c1erKKrsuliWiVxq/fD1eujJwbhCLoyj/u
ur29B2v4h6fSWczdtBfrxl2mE4tw3gxTDEIskcuLFXFv3DxTU+2AP4+dkGmr
I3sT2ZhN2zqJOL18TcWJSLpK/O33cUp96x/y2H906Jt96Tyy9NM6pUHU5k0t
dfwVEmYL9sgMGwCQYGmLjuZn/UssVFqTxMYsooiPq+tqng8iEqk/wP8Qmp1T
7PJGxRVT+DMETuTkJ0UmI5M20WUo22/dCfr+vk0QghL12550m4hiK/r+v0LG
zxEVMOsMYG5i4JQm9FO9+Fd2FupxpWk2pm257InMSd7WbR2KnZFk+dsWNJkj
KVvdIBu53W32+FpnjXadplTWVyOZCeR6/VPrdAEUh9OGHNoZMZCrH0YIAbXV
mVbsHm1EcWt7U8LKSXPlp4vJ7iMXv1nV3hR8EJnBwppVHFhMWzTkQ45Q922t
eyR8D9UweI2K7HwJ+4jFZWU/8FWdnj/kN6dFdeRznvGvzQZALkY2HGGsS/nJ
5ZILRyXBPNYFTzdSpZ9Bc6Y+6RB5pWIvnmxPkykLIaYA+GVl9zuobW5cceAS
9iO324Evl3P2cNscGv2mpcd9fqkDB720qGR7mK6FHnDZ0xHNMBSFn8eNUENm
xMSTKtZsy5kFmmi99eD1VtTpCrncUY5DWsczkjU+FKrLAsnz4ncFGc2SeSaG
mRJrAsSQwM9bc/vKkBLmU+bIWBhuHaoHGJuPFM+5UmR3f+7QA6ueLY7TwwIG
CYykhHGCFD3NmYMsxv9/X4OhWszonEjwegjV9YfmJMZG+p+qvw9DPnv4zoEq
qYahoPFSZuUVs8AZdv4FbPXZAZFcMQmuRMv3SzaHv0vOJa2ODPe+eg5TMdQK
k0z7D4G/2/P+aQIGPokLPgDiqE7nYUQ2bWfh3QiwBkcASGWeRJwh0OZ/j/N3
O8ny0Bou1JvfmpJExZfmv22Mhhx0rJueyzJUctyquhifXlu7ZfHCc5ld/glo
7zy5x49TILi66BdpwRi//nT5DZZvqsS0GZV9+kyGIaBzYWTmXDl+sD//olIy
hQZA+I7CyFYo5k2omYvc0axGqxrDxva4962b6oyYRtCjB6U3FxhFsaW4nRH0
eyiMK+mqfK284RLsijmUCxKKfUUg+XQ725f3EQmQQQwVzpWw71uWMurhcesw
9FdFVN0+7gbOVkiTL7eVo80TqbVywdwCxOqhg61ySan1MXxD6YWRP49OoVvL
9wYa3rQjJYLJR0CTJ12r0474f6bLxC6WLBisroa77t1eev+J5pKtic9/IDuc
Td9PPD0xMUEuilhPPAwuXQL3a22ELzxSUAhKUppOYHGoJ1aPTu5T1thA0dUU
F3BEwhDbPl1G0bZH78WAyqtluntLxKUpKDcm/MS8xKf+ITGq5Nhtc6AdhKwJ
S2n5fYKHhc0QUuYkJgtbn4HntSHCEQnRxdG64TpdT8QM4CFDvC6+TqwFUuOq
auWO1gtKfxWx5fb/NwuT/1MaWNqcvOj+JwveohSciq/0ISw7EW8xHfH8cgQi
JRFtGgMlKU6O2zxDeidLskNNngwkSObx2Qwy8lrgcI6ZS3lTTvSq3qlwrDT7
xiRx8KYFciSuK1JMXP9cgI+P2MBkmSxJI3V3CNQtcw4JR3s0bSuwiCyw4M1H
t/4Sy+f0XpAs8jv7TwENM+2q4/vxp9nbq4uUsqntB05Wu6ytmyJinLcRUMnb
kR5QUf+XXi1HXwOLX3f/Rt3I9H4FvRSQqG4PDM2akK8u0LjEyLgA6moYHfuo
6zBkXN37VEWG/1y3LIb29SlaHo36tc8Scgc79PKqTB/5qHchJC0aSxOWQUdN
S/0d4IA02gL/4wmqsTuqqSiEhVvOzxntawEqWCFDdjZ+g50h/BPgX1zGAxAK
pzzPkSrh9btbo8NjvKZVew2sAwsJdPjLMe5usJkTUbC8wyEhmqzLQcD+VmQ8
akzJwdmNJD8oRKS0Ffz2dU2qDxmh265Y4m5f/cOhxFQeD4EXQTjhyX3yqveo
0y3OODQzMsWpsEz+QlDuMwYd4oZ70Ky9CF7LkjRsS63EU2BxRJAzQPnbgs05
Lqls5DOHz8azbFUrDY4U1uyn//w4ufvW4xcabqNAJ9sCjv7DLzFr3qRvYapJ
GbFJJEWrldXZuBuX7qHMs4zUhpamOIB7knn3LVAC46LjMzDH4fl38B8HFNLQ
mfRDJ69UF3IjjGKHRd19BpiZJ75DKs+BY3hqdtBJSGjkX5+40khLkUiuPnp1
EimS1goKGvj7MfoSLtaF8MPiw7gTgJUI7tgUD/uOF9noCCiKocFjaMH927+u
wi1tNBlP5NPYFQIlRpGbVetoe0qgIq1NPQgH+spURVU9ZulBp7854IZ2+XQ3
ad0XyeXPx1icYKn6pNJ6lsKka2H6E7y83TkghR485/fvzwOYTbKtBuPo/BoQ
VMmLlTdrQafPn8X6E/Y74J6D+sO9IfSDG/BUG7zUw4wgyxdSu0pv2QWLsYTz
njj1TenD0kx5R1JdUiuChBVTvVaBaHv7G2rQfB6m3FM1A+sgXsqMulZoGvow
O8cgWtX68MAmL1VGYIctzuC6aKKbcbZvCcHG2Cn7Z+bqkwcqGcQ2tl5TXnBi
bxhl1FNjGILT5luMGezmbl7kwxic2d9p1cjsMRIn8Ay8gB5aSUSGEk9FLAlD
oa1KPwPYj5QMlgwkJ+2ezJLJvzdl+Py6FqGFDVcbXUMLKzpFrRzySRapi++x
EPj2uGTaGuaTxZY2dGVHQnfrCKAvnuK7DSxxNEg6rEq8qvp6hozbAGR4Zmhi
zSVOYoUvUpQZOr4RF3ITp4Kv5HNLTO2aaNIhGITQKpmu7cznnEyCVJhdY33Z
rpYt+KvU0o0mGNaAwllcAQO9si+/hQYxUik7xtrmaPheuj//YDtHMWmYUw77
A5gC5jNcUC3X9pI8OaMow/+NOSJ940vJGWMWmytWqyxLiBYUq4VA0GAoWsMM
NB3k6yBdwkMlgERwKDGNsqGIC+4sIeaKi8TVB7GlSOUqrK2LVwKFjotyhftC
Z2NUTv/b7FY41CrYdYNYbx2aOCAJkeUsrN1jy/17WXxYtb6e5AOxRcXr+qFO
ggyObAuGKqqtcAxKty76sVyNX3yxrxfCxoir+BYxBXjCw3R7Z2Ek3lJl9ApB
GIzFHlIhksZGF+nuOlKcXDf7CPJFcdyEWf4LoMtwt/dSbSxlm0NEghuLyzGr
TsY/UVEJ7QQ/wCSge5795UwlW074bKorJnhgwZaYpOUr6klDbfaVdruTpiC9
FVKwUGY5cBpfri+nGlY7pXzcop2SoLi8j92sG0SmrC+ARuYfwTudGkkwFQ8r
b6wjaIcC489c/v/OSyVhLblTOs+IFGlVQe+2qasMYyAH4ynpwOE1PKMRgENM
lRAJM+UZmy6yphRstVao9u7zqYZveYOiaO7+Ika+5LdMGJ77SxrVwrasz0Rc
MUVFqnyXo1YvGHJdtMuDhGmMynXh+684B3lEs0zrKvDe1ar55rG5Fdg9QrRN
If9IBqtTX4Wm5otn/czydXOE7ih/AO2vckwqIpH80cTqDAgHnHXpODYHo3qC
gajBBzH1uR95+B9QJIVC4EL+Sf5D+E/te8FE2Qs/1hiF2elkiTPrN3BM6w+I
c3GWLCCs+9jMzet6+7xVGlzgjdwuQy/y9Wjm2nGA/osRqwdijd64wBsqMmJF
kcc2WmOT7X9bByfYpIq5MOqpCE+ebaLg1HX71bhUaurTRoAiACC53C09ekcO
uzp5J9/VpNnL3UyBk7zCXTPZCeEJhdttGOE8LYwIQ10emppLC9SU5nOoYAUU
faXcU9/Njjt9sQcyGprYZpXFhKjXPnyvCHppPt24faB7qjZHyS0TiahlKovs
kww9oOkkmQlhi+gZId0hCMF6cZjYLzgpMsA9AsJM04zsyBcqZCRgFoLgpIKK
qU+mSPXBuC4UZxKCsSy2YrdeJrN/iQU6zf/GD2g7J9VDIRytzTf2c8wTsJCT
ABTDu/Q/mIlpewfckeQlnM1yTKCN/4vlG8EHCB6IdpwsoVNXpBfevUiWvXMj
qHwJd5TKXIHlJmE8m8MFmMIKRmcUkz76o6Fowfv6J8BVtWIxHqd/BFV2xS25
KDcMtnkCKpdR0n2/05oe1KlyGvveEpLJCwq7nDg/u5dQEfflWx4gWC5FETz/
RE7nnf9fI7U0Fu3Z7BSWN39Y5ZzCVTc8VM5yoqx38pDe6gL4eJecAljmV0Kq
Qwtp89eV+Z0Ms//0lSisxqMEk3l4x0Uml6sCdRNrs72dRzywKpsJmcbNWwNF
ej53nlFIID6AVamLa4qSqzi8hAV5Tk57iXHLK3mvoLq1uY6oAhtG/SnpsvaM
lDpy0mrwHqYv8jwfsMpez0yJVLPkBt2mo4YrIacpXAqkwp92cbYrmRc7C0bb
iyEPOAXcRpk5q+WVj/AkB64C9FONLY1pkscOKa90lQhTh3U1zxlsagCdMu9P
3cbWpzmTWQHnqRRNtp9WeQ/np88kz8TVeUJmDK8jeyCAskOGIdGpcd+1xJ/g
RhlmPT3Y9uWNXXQOAKf8NwvVZ8lG16WD5UenN938adFhgW6d2rwM1GEkTZlF
gceegsFgCQbNqol88QrjR7dBHMHbEJWgiXMxKJk4bM9RZp22aKbu64Bh/21y
Vbmcl2KhFObOwaU8ujbt2Ud3qrn1HnX/V8a05uDEk/SKCAFcvlWo5nS5uE7x
Xa/8T/q+5QoXsgZWbnxS3I+ZWUYfCTOLWJpu1vOLgPBzXrP/RCALa74pzqQt
bwNrUF2j8njEbyJjHIsteaN23TZfQm57g0o8gmbt5EjF/Kz/aZd+7mLc+iVq
bxj2m9vicP2Qw0uFRkqX6grZMmFt7tikM86aV4cKHlnyzvdYERTJSiLE9V3A
XlMOcnTm4aJx08Q68LHuT+UWCp2AmWMRpPnUaJVML+b3cLLOEFgR3vbGQhvU
CqkOdIw3hWf0Z/kJVDdXmw/CzFu4A+l+VRoHps45ufFaZ1vYH4/MHCZZ7yhQ
ADwg9F9KbzTPrEeUahgYs2ssaj2NwlTr/A43yVsxVwDnmnRS8lJX0/Ma1jQe
X3Xo1oOAwRlImzuJJczwnao7siHowzkPY4vH35YlT4bldS1wrsnX3vSXs7aA
maKT9qmXjW3xHdBApTSCytqRTenHh545ihrq/8jVcFEvB7PQsWixtCIECtfa
qtB1uTU0HaMz685fYmbxAbtFhUPJKArTueekfqoqTkGGBQ33lv8P5qUYevsF
YW4nG2dJYbwQ+UiO7dNvJp2tgFYewq180a9+qtULRLj6744iY+fZmSKHP70K
7ebQGMHbx+CnSMzsuiQkEOyl488O85m6Jm6x3fVi5YebX/H+BzdWEfy7Plgx
m9rQijTsSegNMHoD97N8dDdCqZBAYVO+pFrrKvSyiKhJffqWJZY84iKLOHBz
lQqcqYU6xiD+e21aWsP3aEays91CpCusgdaePhhlUbe6f3Qdk8GSgQ9bjQRA
NM+wjs88weUQWU0Kuc3bzbu8oBUBNGTeUN4nld9/sLhMOPaIJ7QtSscwkEYL
zNjJLs5/OXZjazuxk+vvi8TG/+BF7++OkS29DYUDpbUd8/rMKqz+HV3aIOs/
JVqqw8Ds37Vf8DqUL8zrPIIWYwTtks9uicOeoFFTeJECNP+qG0wvJZiLu390
SIhpFAQ08vOk8oOI4fi3F+021Lp5aX34yfhR3asuChcVVqUWKmOgRCGQmF8R
eXHY+kfQdzbSl1O4yyI9uxyp2sCxGeXJviiDjtrUFKyOGmjGNAC5zYAqzyWX
HGlQXqk32n55s3QmmFAzjv6IzCIC+YFaN0FtYkLQvnxjGz/9zH/nKhbb4rIC
TesRayqtWkM6y0Z+ApEUhoQMtezAU9EZXfwcxNYkBL8ObCzcQwnZNbF25wqC
z1S1r92rn63TZzUD/wQFfmO3ZUT6BtzsP+VOpD00IhQArV91G4B8n8swe6hh
Cn4OwrdHAUitvqmhxVoTXntGia/N8dQpE8QlkVLr+jeRwcIY8impDTR9v7DB
PjQMklWr1U17I8Yffj8RHSdQ+i5IomYkbM1Z1Od2VfCZbVEkBfzkmaefxeab
bY9v7dlsKvTIg7kNHvdyR33zREzFpYZWO8gvD+sS4BfoasQ4l65C8Zk17V6X
CDna5h89MS9g+lX0NbQFOMMCGcZ/CCu77G4Vmvf68fWJPHa4tICZJ0zlIlFy
TSRncAVCiR5XbWRYLGAZSRCpU7h1wbCZo+UNcl9eF0IJ1sPiqWyNTnxiBkma
fKJGehrM2xEfpEXjg0b36sVh4pT6Hg+c3922N42UJ3qe0eyywYvd+xz3/gZm
ZTpDgxEXdAiW+43Zowc+71LkAFXzlYXFyUllw+ox53G7OdB92SwYPqFv3tCs
BDt7TxN6r5d9dgwArQMDTgVQddCgu88945pqGOPJ9H49jcpsWjLOZc3MLj2v
Gj3rue2AVwuzfnjM11HYQrOu4t4BCt/JUe7VnkuJNw2cHiyll+m5YItyuuNA
cNUyCkk+G7XQS0yWMIfzi2R0ECwVfGlhkA/ZE7UZcB4CP+z7/EM5E2g+yxQn
ONfI2OmEOHCeP4Lkezp6+swCCfutt+s7LXIrGVq5NiRUlEJpD+7yx1thDcfL
z8kETHlAtNUJhuxKEyOkKJXkLqy+GTbnrcX910auJiktcRiDAewy8TCvziT2
AcN+d2tnYi8CKTRe5eYZlZRqhMLnN8/IknrEUzSmEHCcC8Vb+8EdbEPkWdJB
BpmtRixDsth9HnWycghO0dorlhHggcsUVSatJy+aiSMC2vE/leKEkOZHE4U5
eq5gPYxIqHD5IST5fqYfYUZOSgeWgkWLRZKb5+qAxZKH83mRB99PMdQeC6OB
NOdhAuIOs0mK22ShyqS5UFl5SNI9e6QG7IJVfbTOX6WQUOpfZUHMFZ8T5lVp
iDoqMwMBxEENwdfd11cFsvPe3Vlf6KjsFzYq4XBcjbPKJjFkPZPLRYhAc3aA
gGMLGQhXkDokxVrcGYMCjpXsYh0TluAWUqI8SGZNpLSGm2d8pVUiLEG7bk/8
gp5vc0UvTSSBNnIvwWgDe5UYjMS08JCFQfJFHYLbFDvSHA0qpvtH3vf737yr
YPNrumF6xDfZe1cll2xAojgjKIytAXAegHAkEyAm/5a3eIFavzaw7dbSVPL8
BP60279f8x/gaxufAPoCwhlE96wyAOOL9I0yqbUG6/NdPlevHF/jDFGsndJk
2X/sjMyXQjqmWKIvAMC632Nf29j21pkqu5ICj85g1Tf7NR9BerVi+BTnGtTp
EaiMO6zO0xaU9Ljws+hPCPKneV+fH19kSc/yCk+Ul8ltwQoMp/JgS4Rk87W1
hY9j31d1mETu6Dw46j4Har82SJoq+M8YLfhfB/1tq0KmnxVLOzCz/Rg2KJJ6
3nQivh7jTc3a+nVysNB3tvAby3IA6eDlGBgdkbOdU7Gawet7VpwiCfntesYi
OROH3rR/C43Xfpysaq8ZcTzcp7qczVkoeP14zQEW96ihUBjykhUR/JeRVKnD
lyq1Ia+EBtEGNrzDfJWK3kBfJU17vkLT0UCFiObqtr8YMldqIxYqLBN7k027
NEqiqLHEhGqmkTUV8beaiGpSGfH5CuvqKpCe5rm16Z294N886+eLOiR29ZEW
uPtRMR7D78Ai75+9aB9zINSQ6kyL7Gb03/wpIRehVxRq+SmDHwlC4+kSYnfa
kxHw0tB4ZEPowPLBIoFKySIWV7eOZi2D8quJT549e0O5scRBwbdesnShf7Gn
ags+VinHo4RZaVn5UAQKvvbuT/mZWsToYYmsysN1lPNo7cF5T7Z9F9f3E3/a
fzjRDx6BM4rARKMai9nwmviCuNEBRZ6f2Z6KSPFAKhU3wt9C0pwko9vUQ/X0
gOV/8DPSZBPNjDIYAlxGRyxEZFqECjAgYl4CTb7TBM7tqPe2kWiMtfLW055+
8ZCfCddnWV7VKWiPmcdktwnO5PiwREigyDzyMQ48UpQXyjLReqJ63n3vYyLH
tYbDvASZNHQq8+2NnDMKMXyNZ7HAWrG5rgM4ihXLIW+2+A6Y0If9Tt7nti/Y
RtBYLCiADHU4jzeew4+wJCXXyv0waqbXBpWgR3vUv/9ETUgD85ssd0a2kBec
KzGR+cjmgUwz8HZ2NFeq5QbCGMlKesX2zcpuFAM211QYBnMoiK4rBqEMTswq
dyBe6kyf1BYyF+JfexH7OHWkKV5j9k1qPFvianIIUFh+uC3iTjesSFvY/VCW
Jo4hv3DAz3xubhMLzFaWbJ/eIV7YwIPzaHLpfu9byS7BHTo1d47qy0pWbVNU
gSoGsXbY1pzYO5qznWxm0WlKm2tSfNKCNpFzNC4lwNlOgcD2jRu0PxoKFauE
ehO2N5/X+eeZF5CUExkxaeK/Sp6ey3Jpjw937Vk5cseXvj6YfmsqIisNua3R
ylWQMDB8I8jPvbRi3QNzYr3OCeEhJ06BjhSc4ujVNuOiqXPbaUCzpeeP2awV
N6WG1nroQx7ZsJMt8b9K5Lq028aM0vooDVwoceAMfXJOdTU3/y4fQgy1W8H5
ihMh/oBWOk5DK/abNy00THIBvuaKgBeIHsT9KDkalYoqcVimAVtJgaaxtkd+
zh7TDRNljTeLC5YI9o8ydXa07oae7qv7RMfnjTwwClq77GObP3Ch7KKcKKO3
dqZ3dwB3rhN7Cfo2zMP+Vkcbdo/XpywjSaZLq7n9Kf/bz78YT39Dqoyvpt4i
JVNLyun28EQA1iC2X55121nO7PI86WQJnyWrVNIrucsydCoLR5I8EfltUzMZ
Qq+s2xYQAOF4F3JrHVJ7uOLqIS9gzCR5cB1vbI7SYgOQpFbnGmcnjwEYti73
cj8mkx8EaDPmAY5BeS7GF7gX+W8QsnY90GpFd41qH9UIzT8lWdaw18YLmU7X
5EKEgOXm4trIe+SsnttnNbovAt0GDQ8HKbv4Rg9Q/kd/1NN2q2Yr3iGr7LBc
tq5UyAAEQJ/9t8OJPMPDaVv/fNK22ALSDG0g2LO3biIJFDoixxJCRDwG91T1
MdEnYNLpzpbrQqoYzkCqVqi8dDWas8evb57Wqt0exF25lSF8rCxWJ7hNhnwg
BfPXfxGNV+/VM6zb+3nJDkcKwXn0uBH593nCV9bZJmulsjAlLiv6IkWClyrS
CysRYmR54pfAG4Tw7c+56f3Gq/Y0EHmPFtcSR7FI6ja2reHR6m6VJs+TMhCW
u6PzNxhbThAdhW+qXBfDiUctFoHQnJAe4Aa7JcFElve21b9DYyfwf8VNZP10
fK362zPkCvy6SHbsEV9hpZvNFLNcN9M3IbHmUli7lYSZy+xFDjXxN3zbKe+H
lRq9LA0OgHdYiM4b306qSKAZhoPIpu/a8V61Z29veYYnH5QnsdrxFvykGPOK
jnecBaQFabYg0iehK0b3Wd5EuKSNljJnc9U3EJ60euPH87zr6/IaasOtruAz
RzsiWTFnr3wRNRYkYwtYuZM2VKutLRJAisdSJYSeH+Mlu/31hvO/0qMqLg9e
DuyFY+yOOLJEB77fXG8aLxZpEldIAV1tNDaaGQ/6q1fLBWBtjnI9mKCsmDyr
zNiBLrmcOF5Qx6bHFIws0D6rrpLl2KvQSqZ4OeOlbOYBwMQrQguSDC4FzNi2
K5jtErnLdYxbY2N7T3CbHW4AsFTc8ELIwCh6MhQKezBFCkXrLgzvrRASJIRn
Z9S3YhbMUoQ98odrd7/2VeYJeClARrVP+CEz/lcV1mUDO9e1fRaHPsVX4Yc7
qdZWe7NjkVzSHortTiTKklkNUf++v9X4NMLsJOuemL5kM0L35WPD4yQ7vUJ1
QWsixq2EzyzqjDnlGFDvK4d06s5rBQitRfETkO94iLOdUUkprOF+jh414w0Y
Wj+xxbCqZ1AlcbD7NM5pDQIMnLPeDmv4LwIXu8UIA8wpo5C8/tPOIX8ARl7U
UPLaAHZjqqzkgZblFU9+d33x7LQFyu/hMtWQ76FMw3FqLXKjyQRXqCcf7zhp
mD47H/kMwHL6cGSJm5qCKIlf+slkiInIZ1LXGyAPCVF0rXRj5FLJIXl0nhcU
N1gO3CPiPtbKzBevaA0BaFfYA8Avdh+rlS1co7ZyiFZWk7AVmMjU4V2bDhnz
99SJ1HO41eMjDWRZq6h6KkdPL6M8stghoFARYfLEgKlSJZB76/ts79iKQAIv
xqAIXR6aImbdXUGgMxe+kJVnnUjV2H1jkNpL2VzPhZNZdnx9SlKOOv3vlaYn
NnhtBTVpUBf5vuXR2IjiavemVKv0S+vGGagyi27JE2Ci6JFUSvHEKNRQoeJf
V225lm/+aCnKRdRKRk1Imi1bCGhEUS9hG9zXohQytPUHrEXnBHY822ERW54S
juoKC9FdPbLa3/FqU5u/KaJFlbMosX3R+nbO/U0a7ooCksshuaxkoLWOpa/n
v54JbCcdmLFWxWUQlrlVPQgO/JccQ8kHh9BHt7DD3xF3xdKGaGm8KfYhrf49
fUykjRCy3oTrbqHPNHM9/U/W6XjT6skie6At4aur6cwf62UiCSh4GQRdsBKw
/f3Ip+azcZAL+scP6TOToZ4jLi829quluSzmg8V0//FZsFwJvjO5+05r7ppn
IVwlZ6HA2VnMNtpI1iF+Ug3m6Pe8QpA/cRGCwaj6GPOhAhu3EMIMcjHxJsWv
zv0B6IrKJQEDg6Pc3QYrphSiJFf9rZ374ZWBSAyvIgJ5E2bRyFsCHqnVpXOS
pKRZfwjhNyy7FjSs1TEcPhqGk6gntOz6zIrsqv9LBnZ1aqkBRoMrwG5nsnvI
5jSLa+e75Aq0Lj+IK8zUpcegC0YIgOQi+el6+FM1dRXfSHMVnmVcwn9WSILM
I7fnsa/R0RVgiXmh3JmuifeT+NYuOn/up8DMei0iXajHA1jqjEBdYTHygdTX
XUMZVglriQPAGLsrH7g9mhVV/QsXLbyNgUeQtY5yU7GUwwFSS6savABrIS31
A57TGjhcHLZvfKdpbmcUhfsqxk/jW2L2LqiGFHARVD3EFfKeqy/dvpn0gdwE
l0zykUz7icMHWlpOuCYDr2DaAaOXWWBVG/QLYfFPPEMqcdkuncJOb3REtUZ5
wkqpySqOlAUkFm+6LQoJTBw2zGKPDjnB/92zcMFtVsGGKa+hCLNChoj3AL8x
9seM5kiY3tfiv3MrEcAICz36W4jwVZqfu+AczJDkdG8P7+cthQVv1qSCaMbl
2e7pxJjjBPf9rhpRrSTzmb/MJSiheqmmMYLdfLZpJ7aatR61zMIrGTr2DVfj
R1cmr/sji/cSx1/STD6qKX+cKplJSd6+ZA+phwClKS3ceZehWwCWjDudX8av
i50ZTe63tWzT8DGAelvmyCle8wovyjtxjOa/uWVF5CdCPtTEmr4chtQ2CjqZ
1u9qME+2TSw566toMzTXXBOyFIY/ueG+tGYpsJ+t5T4HbvzztG2X/VqCn9Tz
miHzm/SnkRHOAOFrPhNPerOdHnii0rPoNdl1f87OjlAu8HFJ75rJDtAdOXrK
mrY7w0+Un27AE7LVOkuK9nJarjnfpRpsO86PrulnYdfUwbhBrfTfcUiNECjh
ydRupvndeAXH0rWhPObFGZ2xzMXQzMgST9XBtpokWK/9IFSBTZV8Ks5ywmtR
fpi/eJegl9lsA5XglMjShFfzU9EM66mAWYgFuRC369WRn36Z7sCUrw54Lpb3
nBaNaklHo4jSNQkvprljTArgTo2/IdjS4NWthmyM/c6mLddM5rHD9kEYrfoE
XjChkuLgM6JAwByeBbT36+8aI8kLLj8rhMRkTjpWUh1U1VBDXwFILX8/qFJW
byscbjnoYKK57HjeZlRl3oeLL0fTsad04DOXZWnqFVIvpGDxo5Q4YkRfN+hb
mJMK91xUMRgB74aWI04ZRwoxrkE6AuIrxEU1eANXSdB9KrXt4Iql2l8cDqPM
dlsjLkUsdinRVHefJ5P3081LRzKzQtKqv+DSS7UKszCANVj7Cbi/Q+v1qaYS
iwdko5kEwgeXueqVqznaZAywiQShwiQn7GeS+kqbJ5KRHH8RQkyAuoYMiLwU
ANh628pr6SjFG12dxw7/DKLhUFBMikyVhI7efGNpNk4pKXpFxqRAEGcrrfsF
i/Ep5fGQjBZlaUbdLvoEu26AZ5yRcjYQ8okm8yJjPwWHL6Eg+Z1eQHj2r1km
9sPtcIY7hO8hV+aO0Rop9IyQQkTmuzq9mkXLTw9IBgJwwtUIJkqKQtdToFrq
I6RcRH3+wDIdJ82gC+sS/QzvWA4E8VtSLV/qx4woIRV/T36yqbu0l1amQvtq
WSW/LYEiTRc+yjeq/80HEYb8vu5LPoF76kAWV/jY1xh535Dk0jQHz0VBFw4C
HyHF3KZaTtEScfCj6WWF3ya8/aYe+eG6bx94n3J7QwUtFbS9SPyfzXWh+7MY
EsMXI3HWD672x0JEJFS0r8BCneazEmFExBlB7hiKugxjO+hyFRXpQrm8DQzv
6DZR9FO0bqpINOnscz0N4dm2F6AqJ16CkwWn/qeTrFSyqiOsQJlDuaLSoVvg
VDAHCCb8sLsjZ5NW5XCpcONh6NpDv36fYmT97Thy2UUItkxQ9civAPBZYW3Y
bS3ZhGfzBEyrNvilkQziHmR3HPu9rOHVI6MthBn5jHv1gZAxi6BnugwV7pz7
fEhH1PhGb+qjl6hlMaLzq7XBencRSrpJouLjCECfn+bjWH3QPoPmtEXmthke
trRQIZLnr6dvoF3QtlOedN2XNr5rBGa8LhaG2Qo4+zjpAkrY++gXNjYZ9CIo
MjliFj8FVInd3Ib9tx2BrExFKe/m2TrA6PbvKJO/EhP0tHqM54ADGAeU/snm
UEhFT0nAKU2cGQ/ks1v7Qr4sIC1tKDg+fDqKVMAXkrRBC8/pWOkIiPO7WKV4
M5vYKJxZYYawNrwLMmhxY7cqWjueRwg2Wjc/V2fWm8tIKtUmUbo4w0RZxViR
OiR2+3NBIBdOBWpPckUGIJt15K3x3ZiqIYh6B6Q3tLPtQRTZOoMVKT9rm2ok
uS/6efnhaByPnUzLQZgy7RakSnxpjqvunWRQizcvuC+5Vcme2/IcI+QiAhvE
GkhpGrDHg3Z96MZhtihmkd7MagHd9uZ96ndftdoAKiTrys7kkVARD7rPuopb
QOC1icZToOE8zNh6bIL+unl8l0b5yiKa66u3FK7ZSK3YVDUBisIjXE0zkEo8
SHJf7md9uny0FsxJDeuVN/+9OdlmXLZkpMrrQxJApqqO3r90dXtnJHSC9qfY
rhrZdrgyrtJmxE6uBVQkuDBmudN+IHuZWyaycpWWJb9VopLN3EOufCQCMUI4
v2jlOAf3za9yhcqfwno9bs1odbsCBzt++0YCZmgGkbF7v21A/3Dko527hBGv
eEx/QKFmV7ps8aVcL0vOtqONGLMPASI4YxSfpsih0FpAr3tZMcuaFQqDr+Xz
RpVbkY5dYC8jVCoVTuxcS6HvGg4HpkFeQcpUbzNnTWchpzlx7SpP6CwOEZeQ
4wrmxEZMuKcqPcs+vWFLVDrjoqZ5h/uculdNAACun1PZM7AncQBxgTUAwoCt
D+0S50t0NeT5due17UgBypPHcnzA1fA7CratEoT+d8mHSFWPM5Nwf0l3Yx2B
/NtwgSh4d/gAZWYJAe7UPnsutKPOozZ4+vXyB2sJ0ggp4V9OR/WYYRf2kwS4
KA7dZf8tZi9QJwKmL+c/fwpMJwgKYK4gyZBMdkygHU1+87v4IANNTC7pnBx/
imV7rcCdxJbvdLfd5Jp8c2HdfN+fvd9bJnXYB8yiqZZuYofvJtQowCO8cxvt
w55OG8F+f2A33ZlP70xLc8NlulyjmJBLQD8QNy5N852xOiVoGp2h28C2eOtX
bU9747cvGUv3mXXCTUxC2DsIOgzjCD9QsLBZWlDdgU6YKPo+Y8rDuPLtUXjz
6qW/vc0vq3VZm9BsL/6G+kPkQAYu5+SIJI3BHxH3bqR7m3J8KJjgTidiJjB1
6D/j4BQEzOAdvS9g/CeDl3ZBlzncNDLrjzzJSoat1sySm17dfoC74ZqOOMCt
ODblv+pyO5Rl7bYr5F0OyIskA5LcmJOp9tojMoo1DleT+JvwkUdlqNsW0Bj0
XnqE9+SOAryIgbj5EP/E4p7WGHE8RrhmhbaK1ZlxeCdaZS0gcGTBMvjNniNG
xYsb9M8/5PHtsvcOCyHwJx2DkdQ1ToiElT3qUVge3TNoXOPPCrW8i6sXO3H0
ju/DhBlSGIOzfACH8HJCjHKQ1osl/BCnYbX9rjzqP3WZ2NWZRAgc2Xz02TTh
7pKs0VnjGsGEZYkByFtU4D4aQrH0W5Wq3N4wDzKFHzZ7GOlFyI0hmIETO1os
NJmTuhTLCy8IRJiNzYq8E/MCQmcILfcN6Z11MH9uANgFvHLq/J5dAaEod8pM
JZZqb7HfPvuGABf+Cf7DGF34qDTCpJl6MOJvuKG/rl57Bu3Yyl5FmA0DGIGy
cjyvzeG6+NpVISwd54eJtFgZHsWhxGw7BrWzJ9nb6OwVOO6Dd1BlfG0kvXRD
bDb94n3hDvBKN3NoLJleoupuSF6TXKZztgG3UyTKTiPVzGfDVfTJ3iciANno
uwE6GlObQFzqx4HNPjmoCkpNVZPH31F6vza6DkEqFrVXKCmDSl4ooUqdGqXW
NSNmrTq6DwppyDj6P/0aIPpZcehQOKqQCFVuwlWT+U1txSYFTinZSLomYTdS
FuxkANAgl9sXIuNoewhVVasqDIIBIQ0+gtGvKgS8sd4AikFcw9/Kc6/t1qVB
rYtPG/iK7nreMRA7md/7FvHijlgP/E5iGmz141p9fjqiljGxbqr+vxhyOhO5
VDUWI7Oy+CVuyOE8uiv6jd4ZKyCGEzkk8UmPPFfDH/D1T+SVaAh3psbrwg4d
j9MeXt9igK6hQggx2KEs86PYs3pz3QsVMJUnOqxxOxJz2a3i5BtCxN30Eivq
MjsPbcw8TEND7imrmr6nUshVbXU1gvjseC+0HiMvUn1tRiVUSNAB2OfWronl
yYP8MnNKMvts16bPtqqztOtQUGYVSPEc9tOTo738KlJNeC9WcMEdizaR7z10
Sg3eyIDYj+gPqYpTuqi0eOqbARysMZPGMNM2nY6CJxEXP+rwpYdBdTcm/8xb
mJPBVwQx3/l7pvFwOI52GpsF995USjf0/0uQ0nU27AYTjaXnYQ4oQmrPMZy6
5GssPaYzsN77kwecxCgXnGuctaoaF5SXItDW0dcq7RuyJX8fJYfHjMObcPXd
GN047CD7cbjZ5JoAEjcEC8XPFEl9sBClyVkLfk6vWemvT+t/Su4AjeSDAur1
uaz+RYWZrPN2gbjxzIqdnNuFnbg1sfUPn1jhIkjmTFwlStW8xaRhlOcE1Efz
Ez41CAMW1YpHItCf9yd4MJmnmJe8jxPjPNduWflDnLUTcz1ME8Yo9R4t4awr
waaTIoz+YmEsgGejQQ0nd3DM9avo27OWIrRNyP51SVcivag1aug649ipEMHF
O2gCdlD3xTaUmORQGpaG6l7U3Akk7QAeiVrux2E74siFmG34IRzfp7cJ/wnr
bS3O1jBccDyeNsgiSykKDWnxB9GQRCeiZOkyNNbQw24iT/RI9aM6X1PuuEFN
8Ca6j2kYIaGquU1cWIomt8Fub6pFmxs7X1Dg+8tC59bAQ25602lHTOi0WUmY
t1eD7NSKLYP+qJKnDWFpkA/JuSGhg8JGlhWkpR45USiqVAChyO6ZKjgFFofm
lQkoN7VkSRLiqywNSECYgdyOhBqo/1N51u+GAkiDtPRWiQ3539nRfHIR+Y0K
1P7ZVYvTyUbudHUEU7+AmvMq+396i2NgVrEcnkYpamiUbuhvb3q+o1L2W30q
7TAq1k/+Ox5l9LNPjlyoK+XyRE9tw0BNAcDqMe92r/6lP3ltaHq5V7lzSYLj
5u19huY9+8Rxv2MyCMKAAZ9oWno+dMDu0PH1iOnQw07/x7BmfV6QiiRgGJM+
y1kkWFl4OoHtfXodpmceYvyvicd/68yr/0a9dPmwQVV+/ps0gwybdWxliwCm
ZBhZ7YZ8Un+VARKzeSEh5K/b2E1/KDgSFB8QtrIfAtVLzUNpxVYJk+S5UYzh
wyXb2j8JRY4wWFXFSGN0MNwhITAaJIyTnorbfUAOE2RS2N8vL3wNygRYeaqb
XwUVHmflRKWZllLhFBkRfXKP/4oUhf92mPXrtAua8SZxngtFzal93pNcxOq5
blUF18yujN7CrK/3nZLRfVkxPZNQxJy5RJyiNYTXKKXMWhGueybt2GF+C/6c
nrdPZxH8B5myPcTzwyxNJmD4LbX9O8XV07OiG6BFmJnEdPO1dHCLsGjBm0uz
yb3erRY4trlAZrmzSTMk6xBvieV54cNGup2yT2hdOqOx4M3zMXkSKSmqffKp
Vy0q0Lzzus8IMHBXvVJRBeVMiHb0LBK2WlockZrqyyFtr213w7FMFK9q1Uks
tFeweHUpTmCJLy2ur0MHloROOkaFmXFJoA8ryQpj9/sD7cN/nFhWn3o0wSn2
feylW7e+Zn1RxN/VCefrTImQi79PeWD8vIbN8X/MHprdbdlycu6C8xe37bn6
Gf31hLzmWeKikBw0EHYUiIaaoG1fnhDK0vpoL0574q4s686xB/onYE9GVA3n
kRDrR0ErGXZ4wIwXC4keN3aIMDpkQKtF47FA/NNSvoxZi5qSd/BzEn8tbHiN
iAlQDsDhWIRDqtioxahu39CbvNXJiChhV74mHnnX51HKE1jctVF35wR+YUGk
UC8+632PSndbM0sIpXLUWnSOVsKaQoalSTDm1yZ8AydP6UWOuIAWG5dJDuaT
LjBVkcRnHVspmrWdNHfLHPCAvQkw/2KjZE4ClFGre7MJugjr50zHfMRc+fiN
VjVqcq9V2gb/kn+6Zg9rpf8rHNJswe0o+bXdojh2OCMIy/1YY6w+RkaVzPB2
NrFoFaFPJPaZcJC/8l/9Zr+izwaFgfmrWMonolH4gLZTzvgI45T8gcPjX7A7
Zd/Rf9OKrDYRXhQk2qPHTFAdNunUeQFyLhLrdxHOaas9+j4Bo9/8lqWHckmM
3mA4BmpoD2RtUD4UJf2J7xdGGBupMm/3f3wVOsu3/uUqYZDnC/9Ncwy2JXxp
7cYlrDWG941zmdL4HoSzyB6x7DPVT3MmmqWGn6uOVs4n19N6YCLaZeQkd76R
m29I0utGMaTP/mquJ1pOzRbVvDGg1eWxgsZJOQXFU8BclkObGg0jTEQW2nSX
AYDbIJHyRLTpzbvaU21TF8bnEbRRE4g5MiMAT24aTRqaQPof1EiofZt68aQ3
EU+R2gWYmFoAWedBE6oaQlHdWwq2ENKLJnRWtFYLEOXxa0ARWBQcfwpWodKI
zBz2Vjhi20ELiTTgbVF/ns8oqga3CQpkxUGkmkVtfclDgYXiXlSG1mCbZ9dM
B78qfMaG/v3fZiiHr0JcoUeqEvG5Rol7iyGTSkA8VZtoX6UJ0vtHfY6wJBsw
/KFjSl3hJPOMyjSEEXncCnuaGr91VnMvAAJ2+MsIKGtJq5weD5/cOYBSaeiu
p1l6BiWtmIhqlosOAOlVSBD9IqB8gx2v6rgoVA8ilihGTeoEAZXZOOf5X81z
Ta4vw3yeozZSsJEJfr+sM6dVw7IKO5Qtxa2kLHp3bf4c4m9sajS+GJsGqA7n
MOeCyWi/P9Uwb6+6EgEWPzc9NAGSam9OMHPziXE9CFpbkiULNdd97gMNo0hc
RkmLUwTxxq8gw+gGMuEnMyBrVysFxGbA+i4yRfV1dyXBQGX1aOzSwFFdfBTB
F5AxRmv0yEYPS1EphphcpAvJCNV58YQ5XGXSua1OSWqQ0LeCx/UCcTXoMrAV
7r4tRg8n1ZVopcAlnIp08kqHYar/JurqS+zNKLZSZ3EkdVIXRG/tlnBGsaHU
GXOUfJbWHgIg6O4QlbzYLVe0yqkPXyBNeLR565KwKye396ZfeDX4Q3kL6cqn
U1iPGZYRoKS2bvgxxDvcQm/kUmPaXKsNVO+jamPzGGAvlDi5c4Lxi1yipUy5
7CoSIniFGw1KXVo/wrnwnwtto80zqjVkntC3OYR7PiFH5SJJybiGVG0Qn+xE
LKvLyciVvacLm4f6N3SEX50cwIbu54/ou5xeyHho3jXYsyKxBt986bTPMuHa
bHVdzgRnfCgUtP/NdcXy9pV2bCKwYlqEhF8DYVCmUs6MX0ijc4rTN4zrgtxI
rOZMnYVzeemILJGw9aDFjNUV67gbNPf86w/GMfGpT3SjtowigFYyik2LHdcP
nkIi1xQFijiAPvL6Nob7+qlZF9X583SsdvPuBP8p1fm718iQY3Fe5Boytzrd
BrBs6brc+XoduWRusaVxtYUJO5+rjv1El+fcxMjjU9jX6IQ1T1/xoZolt08q
1w+vRUdjXssbDBe7ofqNxrKAKhdOpCouiKhl5Go+qjgd8wjuTyrlPKE668kP
8TaEH0Wv+W2KFH/7ajWGN0uCn2BCNgcVpZJ14ORaAGghb4agcGxnX541cpXc
1/PndAUUshJFVUXxIdCpmmCL9Rq1UWJAGjItq+44PmTjBphfsU63n3PpnXdG
LAva6ONXlYyT8V4U+6u1C14IL0YIT11aG6413iuKjWF8gzndSIFuLo5WWOJJ
dGYBzKc4waeNSsoPGhxDAYom3viTDhdljdvlcW6BbxPbmJn2LyEKkLk9JEhv
xS14WzbnOTUyWmPZWbi3EohPpP8KPzMuWBJ+HnE5u2weh/oP/Pvk3ZQcGXTG
qTlD5p5BMZZ9DqB3cQOM/nb4buN22cYvGuaSch3VOryEwkKN15rsnM2nl4EH
o7KgM8gkWqgO0CMTJc+2zZWpOikuOOgXtRFzXlwfUR7CIPrXXZ3pk0uMzYk3
ZB1FX/5wH1Q8GYel7YBiuzeswcTM7R2e+b6yNj6rwnytFga5j7jKxJqhojBe
NZoxmDUatg6NLMpIjAVllgNtxcaEdM1+V3aIuxOkKtWt7Lp2JnNYTMQEXbN6
krzUdK5K7AARZbgfmIZXFpPAnfByvTJi6uAWQL3FJwW0+Vv+dMpGs6D4ZTP7
ojv6JXky4BvBvSLFvngLJ/krePy+S+wpQXQy10NvzZ7swOuCDfJLe+22rzGZ
pVl7E1rwiYjoMQWoVf/lDTVecn6zyqz3UEtkoOLSBdjSUf5M+GS5mbhUc3pI
cRuHs6bin5TQh5ZU0102LUmncx2ofzcH2VY1WTjbDB/RRsMCFowxKePGWIQr
eDzaEJHN1Sco0PdUOgQ3IKy5i+vimneM4kRIR/AJwk5LvjhZmbCUt2N5xEz8
fiO8+jPz+IU35ikXMrpZtihMdnuuyfFIIJPky57KS8Sl4IwLr5ccqSyQQ3n9
qmuV1ceEUC6cM6LGWsglpVpfksXyW37RNFahEo8GbL4lpJGo7SWykMck1qyX
3TFvzss26vuCB2SyDhEHC+NGEQ0y1/AXtbtC9bkYrWBgg9fJYo3OTR029yGc
IdOKFORYTqeBmMGfmymTpDfINd++LWTT36n8FedQWGyKiZh0f33OII7KZGSj
GT5uDu2bK8h4cTN579Ul0KFIgYNau6nzvC/nUPf4204bfQT9Fump0oyInz6w
PCdq8Jw4BUR0hfD4syVCp8iWBLQLJgw/XF5YmJ/4JCtuBnjOtDjzJvpZaMDK
aO9MoyuPqLx5x5ARNcr0OfvDtuz+s/fwtFYvNJ0cDwbuGVRrw46CcIhbBIsV
W9TSrwUtuhcANvRAcKoNlnTWalV0Halh6qAqCcU+JIJmDGiqg0TY+xOcM22f
5hx6+VWD1SIQaJGVny4AqDywB89uvAVx2t0KpNn1CzGdzSkw+p3ScH7BjaXA
6hj9/vFC9sE/fSn8EFvhpldB2OhDUpXw3im/JTPC+3RNzj6l5/TRIRNiY0wB
DV6YtpmJhPoS0e2yFrWK28V8e0KwoKXhWLk9tJIevrpJNXZM3Nwc3am+Kio0
gVCJkMJb+QcPWPmwZ6C5V/TArxrlzT3LmQc/5+LvUEw7409PV92DBH5bjpL7
wP35kOGxiuPt+D44j8Nfngr4yxVDzvuYncHkMqm1amcNybO6JMoTspw2WpW/
Rc6IXBCeLx35fFl95k9QN2NzzIcv2EzHdgFxJPycvoSeNePlZD+jLFawxzAm
f+eXlDYTnI+szc25VR+Oe+EVhwx5FZuZwEAokrK7Fhzo9WYGeqMThCDKbbnO
0PQFE5+QecU5uZkUn9C22buKRQxVq1V2Gq4Ooa1QlKmosTu8sFUpE+nv3lz0
7OmdVnYgimN8R8z3uqrjs88QEd5mYJjgacv42VLDtpRYX++I9k5pHOeGRezK
rSoGroUkxkeMZi7hV9odXKwi7TlzQAQWttlLWcsn5ZJfJb/oMcKna/ZuvtaR
9/T7ANQzApO+mN1tplJdM7vbuguXiuakCzJ/C9nJQcLdIpn62iTiswVery9i
VlSFN6W7I0x5ccy6LtvysPyEt3Wo3mhKOdJHLgm0wOXKB03SSH/dJ32M37jl
FrZc5NxY9mLX4PY5FZVWcPY0wICKVPp18KBywl7zkNaUkoYD4Fy05uISqAWx
vmJb2TKPwcU/LqpYo36k2aLn/JyIKupm3nU0kuIjof1sDxNF8MyeDWqEycbK
e91kKg7G4ifY7+vZ0WkVkLirsJv9G/RpNFdZxQOMG8oBo7X0uVbPmSF/WajJ
PxBf/Jc4y7reawtYf0FKaVplEN9dprQ36vogR7UUFaeoRL8FOq9hpOHHJh7k
mFfKOm13oOcdApXRC9mqKppURWL1VdTJzCsjKE5lAAP4wbM7YzxF14xFcz4J
7TK2yU5S5mQFH9w05bIAItPmWUjHQ/KDjQUkHzQgDtBIX7E9rNGQZvPxof5q
LhRXR8WIMLG0aD0gmerYAXvg8OqV26Kn84nzcZMJ0FPLzGwI7pnJZKVZwMFi
DweOjlieyk/pZdjuhccvtYk7WcJc5FPzK5GFIrJgPIFakLWvRkJ792Ri9/fz
eqSoJro1HebByMDeBKO/VljYFqD3oigFkPekyuAwCh4rWbeiuO3RYbFoYXRY
FT6BT/QtUoO3V5gsQ0bOUS3FPIHmO+W+sjFnozRIa+z1l/sWDFriS9ATxX7I
DazsvuMCbMm8jjphgfuxHAP8SXxhpu06Sri/OmW4eSx1Pcjz1ZpwulqD0vO2
6pQiOFavamkyetFppHanhuA/M6wSpO/JBNH+eUpQeIcpFYNeStyOh7FTD1vP
n/ZMhhoBgsM9vQEpnurS6x6qh3yP1cVHCAitw6Kk9FZXCaCQNfXTMH1P2Pp6
bLGum/xFU53qUU1nFdYmErX11n/hdNT5fEUTssoB/16nBNHADW9GWpLXjUda
7mjlnCBOJLrFeZwD9BUT3KFk7qqXVWRzl5z7YjM+CHK+ZtzYPHvUx20Npw4S
/cl383M2AeegvUS6JjNcQAL6dTbgfJWLtY/uEeczQRQfl4Z+chmftufLcEWU
iXtSiTCCeWWCKZNGPkg+VPPfWiszDQdo98lD9WNFwkL4SdD7xpBZVMw6W2cB
xJ71VYwP8MvsYgb9teHgh6nQZF4PAtosANEZSACyu5PnSz862j8SHBL5oEy+
+NU+gtJrud8lipc6OR5sHF9nR3GnVsiNjo3QDVq9Vj/eokHfD3p0jDDvl7n7
wY0D25Z2+OcYjudbOuHZdY1HA8byTEknwfUDeEr5G5sGi0uzMfp2uQcS+cMh
aaebwDCrHHeGN1K9rtl+6Vd6DsVJuwlC05ZWBy7VaoJwEed9bEWHr2sICg2B
6h3taxFPpsJI16rHvRvPa5dDIA2JclkrEQ05jXkiCI6L/wfQblZJi8hy43vE
gZfIaRteO8qHB3QnzV14D4X/7QKi9PsEGADJLhlK178LyBuizfgQjlziJQzd
HMHCiLKct1EGWKYTAFN3qhCfLPleowZJtQiTucaq7hu1H+3QeAJGmHJO5VYr
tSFxRsWpZ9hiKYtL/y0/lF5+8zO6okokqe03qXly05cDd6IZ602iDj1CWdjA
5yPoekmH+OPOkwtRt3rnEo+Geet7TTRb7RhIaKplwaUkb4sI9JIiS4zepnPQ
RVrYfN6x8eTPU8UEyuy5usErjVjCUQg1HtETz48cfQrJq8eLiokb6A76FD5c
XamOUpCnj0i+fsDt3H4CTQpBM1oNqc9fDbinPP3reeTE5GWy/Gmj7wZwg/qC
FBA0CaTFcpAHXP5phyH6Zov8F7YUY6T94PIURtQXDA1cgjIH4Pfk2+vb3yvF
/W/+rEWTiH38ioyZpDD5masgEDiJGvyfcbSXtatRZzOGCA4jw+FcVWyDrgM2
nfXK1hpaH8Sh93maa5gMwGh8VXsjxM8NdtkVUGZ94J/nOlxN7BFsXhOLxuX/
05Cv9OLUx3ErIvUu1LXgC1zxkxfKg6tciIPHVEdZKcIDAWgV5P3xNUmgFrGa
X4Of+5wcjWI/BRTci4EPYK9Ddy5SJpHgzXT70wALlUwmi483BCPJZO9Su4yw
hRNrqGIXV/vADW/PDUE7HnYIQ8bi9Nsnk7iObOZCNt41ExGzC7vy37YQ7rIW
/WgrW3qNExapexAdY+lAz8oLPMEcrrNeKp0HbLgCo1UamsUueLV2JDyVV2DN
VWxGnbeQIy+TxZYHKZ2EhIOEV200pnlXikiUnySojwyXyJKDH3Ej1aWbPoTE
T23zmvrngN70CXQRwkCeHiEOV4UVQiEA7rvpwBOjtqSJ82lTZL/hqjnaHkkD
pu/w0z5qDUksfVswRf6tbzTt1po5WFqN4QrlzAG1U6u6QxHltsbwFCaE7bCh
Od1psy/bZ6mFMa8WwaN9bx1nOTcJHbzmIzEXuHTfKZ9t2NZ8TzD6W83HW0Jp
BeO3Hk4oQZS0h0QBi89mFMdx6kiVG2DRSMuXuE2RS+j8XxVlJUoO9VQjqv/Z
ovFbtstvCq6gpdh1LH0Qlpk7u1Bu1+f66CvxMCUVma05VImveuc1fER/vd56
NG5bO7SBMhsA9bMQ1yIje9Pli8F6QgPspdWDmk+S97vZRC8Gz3ra9kk+SufA
NChykLRP896NhE1Wh7WaiGYYXQQrLrdSe9Tk0O4/090L/sITz2nD4ibZYVRT
h5W6tczuNStG6sDP8jrluAbjG6FTocJLkej6CEtCEJTIu+p1YaKSdImZWx+9
i3jas+pVfo7uGSVRmmBG7GsepsXusId2jIJo1O5kTgezjrptgPeli/ePmtpF
yggy6hMdA9Jnp2CsF8VYi5s1Xqr6VXk8/roS+R10Nqrcy8SQxILOhsZqmSDH
tkgzvoelcWt4QVG5zyhLTDzkAXAd06JEGzp5J76NnK9xrIR7Ds4nm3CMrTic
VsIIq/ETHpxd+5ysCwO+PPn0uGvsu0T+g24YePDoiqUc743FGA1kl5diVmDA
jvMX886kD2xu8TfuzfohST7g2Gqf8csNd0iFtXcxErBWKln869FYG9+kyClP
gDQwCpkeMJlNwpJJ1Hq4RqwiL49MGihvzPPRGmmg3QkuIsWkf0K/TWmtuW9s
goJgZkZXmY9GORZkems2D68YC77QzXYl4sBkfrjUCv1PJ7Yssv8WqS/Bq1nz
YZmbPklhYP8+q9YVCZdO1AzHqnRBCKm+SMw7bu9J5muHKfSiZF2dWGXxiUhf
rdGq0B1+Sv6u0zbdAhTSiXGz1orijnbEHTLD3ru3JXIwNrRedwcXkUoW+eqS
HpRf9Wvo8usff7I/VhsNl85JkD37L2KOBLqYmSiSGN5iAxwXcwzvXgfKI88V
mFt+Wo/Cdxngs7iN+cxT98QRyabCUveqcDq+GLHuw+MpIQRtsHJ8722AEj86
G2NKHkP1QVuaSUdWLFBkHQkcfU60G63J0rzfQEW+htnV9KKiUhraxAvj6mxD
eRXi0PnUZjYqEnwemObM70HL+69lKheLQhZsl6C8Jv+Sl2oBN/M/bFnEwr9B
FJzbkFMNkDwjigG0I+G2gmPmlCFkR566JViTwTtwmpD1g504yHadMOMPZj0q
YztMq+xtqLhE9E4H97eFuuUh3+/mFEm2KbLmoA915EMSaGkfVLNsp+u3nWQL
atFdaRXq0ajaNejFbv9cff2whhAaHLLNV77wCqT6Jk/NHgqT5r3dKujXB0TL
5kQBmQoyqVFVH3Z1tJiZeBgfkfdouYLy0tvi4B5TPCY6zUwdLHpNnLRD8THK
caCRT120aPWn4DjQFIMx/6NlYpX6q+SOMGTHq52DXCw7PX5VruD8+UMcnbGU
ntHvyq1YP5hFHvNKjbuga+u46WFKxjkX458I9CjCKB2+rE2MpyLySkM5631A
aeIEYL5acwobzCM1bF7sHUtOSFIFeT25Jc6N6NHltv4/tTJOX/YE4uZeUOTi
BvsEgrSKgmiMIV2joFu/EpKvTIIKojVBXKVEA83B/gNXM8Q/1b+/QhugvVtp
o26wVEoGpGkJIF6KrAnf4172+aCNQQUorYc0+Yh38ZjNVmgrseWQBEZcPub8
1fo3XzZee52+0WVxRAaPdcb2oFwV7bZvMJP2w6CrTfZ9QnOkFxtcA3V38II+
zucctjHB4fmspVqRezbYr2fI6fy+vtKk9s/6Uc6ue8wJvsfFIfYPw0RT2TVa
Qzya+F3rGl/nrBl1MYsjRq5Z3Noxu/fCeBHVuCBYJ17ks/s8z5a4J7iRgv2Q
SeQs+t+zDcRrFcGQHtUVpF65imwPJKt98TMROCWDFHAtFrlthLTrAiOOSURd
8EA5d3Mv8vrE6Fxrs7vV5SEjrEy9/vwL4lgcIyP/FD4b1AnuzeAu93R2b/YP
6kuKOgbXNTe74L+fgetSoaxJZPbg76LlXSU9Kfw9VtDDKWHKFpiNARhhs2Oq
TmK8WqWdSKNtjadgvdp69oTrB4TEO9TvXSxLeDv6D2wHlJkoPuac6LRxxCyt
7Pn7rw6HmZL+Ex04zsyPfH74GwlqzqEDSz0n/sXU0WNt+CtY0BT5oiR6UjIZ
vLo8+UnTeGH6f5AaPsn5PjXz7+12vffl77ddljnTWL+dDY2rQF/F5I3Moq1z
c6PvJVrQIYnBWq7HWW95rnHl/zhjANluQzG1ti09PZ+FL3yW02CvUdJcUwld
mxoKrKCKXV5M/CtrKT6/fQgqKyj93yCVM6gKjnJm8eitXbWtcFE+2Lo9abFq
y3b9mLLVpWtn4NZdI5yNNJmCRn3kobfoPWZwybhhaHtJVMxupz8yx8qc6QTa
YTyJWYaribt4czThyadfVtAt9HLLFnWNMzZRdze5LLSMIsJdKkDOzwB5LcBb
AqhYTYd/jLcUPS/ar+muEJc32HQubQJmqKpS/bGp9SrgeLnm/dlC+NyC/VCO
j7cc1aLYOv3ca1unufsaKTmypyRWt36w8RPhEgiMn6ybxhZ45RGKJvLvfio/
C3Abk70N7P1zYM0v1bVfI82MtvEtL6lc1iGvn8e1teNRHbvvVx60/HISVHtW
6y+iaf6BPqGrIFvJ1AlZjqrLnOANG41yLWYyAFni7m0vn9CZW7Lx8Ooy7u1k
qljJMWW693zZX70I2xGwGhf0x/wQwkXcz4TonEi9WDThxZtX4spiG/PkZfk2
iuofNCEsoUu6nLC+qXTNT0CAku63ch0MPU2R0NwYyjdxPkXQB+G5ceGkfh3M
8XaQxciTLus3ta8EGM7jxbM3015bMrDtFIVqNbd9XssSyBIU5kOLs6Fh2hOt
CFSFAwm6JC5KEq4OmlUvTgyTgtI09lzk2yzfP2FrBUyO4l6yAVyUygtrtx/v
Op2L8PQ+vZOLeV4tuxW64aur8hbn2XDVZpipKb4hBlQPuBCfeVNI9v2VVako
RSJCaOvyyy8lqpvEigV1fkV04JA10iDABzJw4bD+eZLt64aZAncaDHacpKsz
ieNx2JKw9fbDtQ6DcDHoJAdhn6t1ZBsqneBpTsuSii3LWGLb3c+p0AWbeGox
ohSNAbfs7ZS93VryCofjUHa32guh6b2faTvR6wbvNwi/J9jl8c+H6iqwl6KE
N6Z0Ndi+qyv1Lqdna+/35TQSRHTM+mhDvPE6BSYxEQEhXkAsd5VZ8XSrrTi4
NOXPwII1VhJvh5kZzRta2XEJ680IAFfhaM9LWoyV1ZFGQT67Bfq/CQ0c4s3r
wl6bP2cdk3Ik1ZAx5bMTuGIBH5LG+T63doV0cKnCezmUnLT67Ex3+foyyqHp
vSuZ4ggoFjGFbw6WyODc4V+8VFkgK/ZHTvhg8G0wraO4LxTmEeK6imXV3Pe/
mKXqXRfexE9jNh9u5QiXhbjMP67blYVvn7JTkMI2ENQI881gEfbvThvQkNZD
i0GfF+QNZx1PeKVJJnsr/r+d3WXnIe/SMqPiJM7DZ47n+UkbTl/emcP2Z4nd
QD6Yh3s007RPGwk4NisJzG8fAqFnt7Gg9AdQhIaSjXDYE4L/w/eqV2+eOOyG
JesLBhCKHRah1gG7ep1IL3nAo+U5Spgki/tEVEyrLH3QQ0jBvHRRTnytIpfo
tRWZXhMEKQdDYsE0/w6xj2BY73UH+Ia3e6DICmX7/NAeaEPSCIpWfviFtwta
WEYzz/EV7HSew/ruEm004mqmfhOxTlpBpyiSIDVRMPdTCYnHGz5QRSWOMeGG
sRBuGw+utpHZHuoFEB4hwD8yAfW8QojYzA6gObvmLRaYx0tzvDrO+pf5rAub
MBEWccaO+6daM1z1mBjCuzkXTCaJFI5NA3UBTKLTg2XitigA9rMQKsDmhrgC
6y2DGWfAGlZYq1J5WfQn1APnnAmyfh+K/SulPCLVsaJRNW9e71/5DH0D8++U
HJfrP1sJhIaQNSQZ7Oo5epMrZdrjMNtynnnNsp+AD+9JQJWGocvNCM/WvztE
Vwp0dzcMg8vzTE601G9jMtSKL+FqYh3KuHUqT8PTxCg1i7BUqWfhmc/eg1wo
3m41gBBsk9LtkdQQiaAncAKSFWUEzUgNQJpDlTGfl4WyvASBz+b92vF4DDMo
CNe9KeV5L1xeDVOr2jTUnc115T/oZj3vjIO/PlwQsa6Ccsq9pWS2Jk/pwenH
RAw4KmrXvpUqHHY0kfzckOTS8uqJBJhz/SUFET2lFJRUuSl+9rxNqxjGXAmw
yzH9xsEKyk/V0xfxRDrxTOOgHXAPEjxzGcE+oy4Px+2nbljEfGi+tzNNZR19
C+vxDraw6s9F7+F6O7EVK/AL8SkNdfK/h/6LGWsCeOkkao55si64az86HV1o
HUkK6wMGeXV2f0BrvApQ/GK1tg4dCoNVK3baU5qL3r2iFS1gP2oj7PzLqSnL
OsGrl0kRhWZ9etLqTeo3jGDcWDbPpHdiNSvMFQiy4xPjnIFTXHI+OOsuaJT5
wfOUNcccRiU98PcAALNkOCSvH+rnJivn6x157ToAxV8VhhW12GgtI8K7URpA
xc+pJItGLxonfjs3Vzs+9pX+8LtZfp1PFE3YMlW/moY/2FsjRe0kyWuztfu5
lK8Zjn4IBWBnQBzMdaph+jl3jTtKmiTAKAEREA7CWw7EgnN0hDvBEQsIiLXz
X+/tWldvrwVj9wCZ4abDVr7fExFffFSJjPfeO9pZGM0Em/dY79168H+AYPNV
VnTda1iclnxl4TKfZQ6t8iATxSgf1BhdN7AaOkM9DXG4h3OH8w/2tnDxwG8F
GKG8a1PQS/NAQbaOtMoPNkjv4PP/SxFG1YdblsJE7rD0lh0KJxRa2bRDj4VG
5TobiU8ZWf769BlsLnQsmOS/aLBoX52x+EptnnOFo5bpggFpUh9Be+iWvxT3
AkpINPE+oupY6uyDY8Mx0c0kNt3TKz4buCJpCN4sTZmW3BAREI0Z0BydWq9f
aGvqqNPU4wNGhsDrRGDVQy8LQNxsgEBBTEe0AmAhmhHKE6zl614EgWZkYbnT
htTuR6+98l2mabJcZEBlIw1pQKRFCJXxFKpUb5GShg54H5yz8QddfVwsWwuE
lmIVnMocA2//lSFckL9thFthBlJYP4XJAB986yqTbzUQldceVeo7fIGgaZv5
MN/2rlpBIFJBhXYE0bTI2HhyqsSsR2K9VEaiJ3lUIpZrnRdBRChBQeJsCJ81
6FUxkV0LOeI6Gf8pvWbUsAd5cv1Pbra23rjZ4KISbIIstidGGtfrqyc39t8/
CvBAXt+6F11/1fn2VUdceQsrM7mEDbKFbKSJAlNfauFUlQGioMREmaj8IhbF
dOGwsvhP5AJ15ksZNHt0Mdpjwkk1bzhOYzyqGFMgVZzLYGrFwQLd/QEeGQ7R
CDsfHNfL9xDPI0IVHt9A2g36hWD5xi2A8YcRnPLveEUOxTMCCnRHD6uDOhqb
zt/YiWHPNjAoOcJGpWBdnHN+iXO8MD7JPkb7xAJbsF7upnOV0flXaLa/hJqM
T7XB7FLKyiu5EzSMGptg/lFNJ5rbSwq/AzI2e5B+/DlC8HEw0BujkVZhoYVL
2B4+q88C0KUx+WhXgsjEDkINYwIff/L0ulsFd9qbxAeVbJ98w0kn89zY6TjC
Kdrh1RiDwNEwJ+2U940lKneEPtCYTFGBxiVNIug4N8RTWIkbhIgNpASLFNSG
rMMaTb0OgDYraWkl+SrrrsnNDCnwMvyhtjhR6fmqLVuqHJBEeG8LV36K4SLO
Ph/xEa7spV0NtCH0QE8ykjbruBx/Vq9doV9ZidMdzeE6ZB9Ja5d45mfhZD3i
np81PTPLP4cHVCzvXNYZFZJ+ZBVnFcj+ghgxpk99Gm0fOcK5NarPX53LwhFi
/lN5Kbz9GKq+E6xnuQqBRJUG+KoQN1y8CyEPeijuQURGkA5N3puLJqxkUJhY
idisJC1Su8isHsUrqjNcuR163/a945M1n5lXzRWWUQwstDSVk8+Ojr0cBQCJ
Y6pBrJARF2lTjHOdd2nRnEW7rUSVMM5WQL5j/yJ/4Bn23zWzEmGyUEygSwkM
sIMY5YkK0x/2C0Mtze0VTE0HT9z0R9FvIrxvsPDf0sADbU8zIz3EmkeU++RB
5mHEVZRglrTNVhLjBSO4wItlrboFpMqfPItcPS6jEj6T+If3+RNlRabXwpxS
hWZHyXg/+zJ/9oQO0vvyfFo4o8VcgfFC2z2V5fUyh58a2jw5973Pn+Jctl4a
uMLSAlXq6FmoIxMnMHdgPECOd5oE02b7AaJFOlWZ0JvE5J0xr7b4QMgNxZmA
emlWn3Cd+CgmfOIq9l0od4l8R8ggeCOJd3fGBNHudkFZvl6M7LXAbgpIsBxU
1/NVLHZcdGS+aP0NLbp6We0xYGhA9mZeIN+gqdmoEIBrCyPm6QQFPDN4fncC
7Yp9oHyotkdlC2y/kZztrhJGYH5mHxvoaHUB8WPXXxuoLdm/wE8cbL46gISg
x94c2stBwByIYCG+gaChDWYDJc3bq+mm8qMLJMcXJaRiaIwlYqM+73WX7fMJ
/dwPwETB75Rjnmfiuv8CUEQxNKQFTMtlBHqW7VbXEBbVrC/81oGvskhH6/sK
boWejUjQe8pRRP8aKqZ3Z+nVfzAFegDcnhF9qyKQTwvuiEB3rp1HiMzvlkKd
jFcnJi5U4TnDcQ9CX18pVmsqFV2DFpcVyATgcq2T5pjRDpgdoyjSC1dRne63
LpnyfBPYASM1pBnMn90teO/+2lCGDuHt+aUvg77GyMH2aRJM0S4mFPIz7XaO
HtSwhJ5JjxFv6qAgLgibUrBf7+zbUTSL2YR23CqkUAdNUWoJvsLSjJPn7ixm
7Uzohn+T+sfV7hdRh5z+/g2t/ct2QLSAAQPV6KUbmZlv7SdslOZw+vZLjvmQ
6BKNMyRjlkHS/msDnSIkrr9OucCvTtnDHIXC0jBulCYIYFOMosOhSWa48JwC
Vcr2HHn+O5815wjj1Es1X3uyvIVqIvgrfL/8uEaBkbFTD0wb++uU2NymFuJC
UtWLfHrjUv6ld1j2Y+cCxyuL30+XKBTOL6wc/bdRfKTXGVZUvb+x75KmBWis
06Uh43q6JvWyy88t8jonaHMSDMkHxBNk/YdI60JPZm/bnhb7l6paAXbhQQnT
u4TOFoUTtJGaqoGDizDb/CxO480/MygR4oSddq3U48nfwAsZa1Mq0xlpEX9z
phNBOFUFsrr7Gu6G5x3qkuTtiWEwW7EshTJta6ZEQIppQoCimsaHTEeg9cRV
0Aa43hXmKLHc8kur+oppeaLBbsCR7KdXPnpxSX2/JyphsBbCYwvMlFcVCpAn
ATqqjPw5K6FNWK+L48D+0rt4gkTYOREnQoHCmotn66Amq1sievu11i/qNpco
7yafWRm+PLPcm/hwUKu/irLZ2sIBXdJU8i05PcQYyosWj8IufpU91pNPE2bc
w57jlZBeLFWRM5vBmlRxy8FtB5RbFbZHRB1ItUsvzezg+22FzYI4Y8cRp5MS
VOJAl9uWH6NQhAUx2IHirm2JlVMDrIxBmajt6BoDx7sLmsXzow0iNrYIR1ak
/Li4ov85tEtN6kY3LsTd+8thA5VhL/3bCKfAhVNQgpt+mzz/Y0Xzm0pgGfrW
kje85uYk8wZgwffo9Ts2I8bBTzqUENIDdSLV5zh97TBz5y7ISl3drfeMDGS1
ArdI6He3FL99JTKhigCBcozwgwUYKcQhSzdOZGwO3M8bwpn9P8ubxDqQ0tp6
S3R0J/qSEb1NXfo31tRor9oJKYWvFl/kDD2UrC9gkFopycyQC28IatTzkRqv
L2yMgoveUYYxA+uyLvRmP9/6xyMvCWyy2r6ED4tqy5TewbwRsqzGmQKfkH62
zn+SGez0Qm1uIqhTvrx/+3/hypc8uz2r3UOuw3IMuDVH2V7pljHJFXMXvRF+
CeECmt+0TJsNasGiNhEz3Zz9tpKYX8/TlkkjMRUo9suu7X/TCjr/rycho2w6
JvOMrnMcBnOmwp/QvXQu7jKmubTfigqgyDc1oR7Hv97LkdL/CEj7NV/DWuLg
Po6E4o9lxPT8J23QyRn3k7+ldJauGuSGNRYleBYq9bdu2baikL4gwA6psnfa
WRZGKS5wZWuvLwF1kdRUq27HN6c2VkBciKsZRsNeZp6wiCLHUHRptzVpxj0k
HSrXTW1hJVuzogQPCbcni4Xy1P0Ni26cPBc3IV1TyOwFyDQPh/eEtCijRftD
UtMXkQ5eXhzZ9II4McpbNg0LdPNXD+W3pm+M/X+n+W4TrXbTyr8arRc1ezHo
fha5fv3le2u71N4OLi1g7Zbg/9WbuTtDj9G44GM+wsY+/zi7W9YIqSQl4g6V
1MEdMUdf1sOilG1HbeOUhu9jxAcXUsoD9RJuKh3AgefXeQJnGOvPrjsLDocU
TmrN5kgU2uTaETpC36MHJVvV1WXVfvEQFTFpWcu2C/qJczSC1HYKLozWmquR
mDzJUCPy1lK+aRHYy8XGlpBgJ0ksjYqvZmOg5C/ffyBhU3UcMZxmEQMBcaXR
s3mGmHavWRjVTAQe1UYTI39srC26Kq6R9X6RpOq++C9JNBFEOWuA6nQN27sO
ksKPeGnjgkNrzShuxQCaxZjH2JVJE45/FcMUYorwqz3pyDEi+AfdAk76VXhs
hOAJ8ZTr4fQ85nIf6f9TVEb46AM50CyGKVsosswOIyU+FFjxW8VP36LUGrrv
lVwlW6FPMzymtuhnEW+IWthVWOZPGVB80SA3bZL9vCY+Fr3FnuYh2lDmKgBN
Iqfl8gGk4+tqzV9yqKfM8sKcYW4hYC4ytGP//X0gZApk79u6/vfWY1upa1ja
GmzVHSRG1bJH8Cm4gawdddayifqiBiPIJ8rHXYv5Q45gOpzdord2MrDjb3BZ
VqyY9LSZKFybtD/zfbsKGll16fOoTTd9G0p/eMc3evUd/fbyxUxaJXCbUU6T
eFYcGNfQSUKQDrWwaisvsVswyjw27afv5Lx4UqVADmZeQkfXBUz2Tl11FwON
fVKphGMcwCuhs5e1UtuPF5cMTU2JMR5AvHFCJ4pvRyHYaE5fl7E+Ymli3lDc
XMmHyuknQwoq5J5l6PZl7NdqcgOw5MLvhUnUFrKbQuSXtyjDpt1KoB9kWXN3
pE0AF6BvXoVoT/dpX03Xok5x9SU+tSC/UkK8A3RYtchtpSlafRSeEiqUklvY
OgWuefakPrxGo4nfXB5iW0RjWQT7867HWCGANEnATnvzsarsJYsG+b6FuVfV
WJHG3dibOtA/ybdw/1OrzaLXQhTrNhLg1Vf5RlLj8cCgIOd6WTl8n5acn36N
q1F5GgXn3u2oJqif/5QcXGO/NHlVRAsMAgpFeQGe+ZqCuZDsSILWuefUchEq
pB6TGVFxO3eZcwVbf8dK7THq2tvOnIxdK4uf5eizYPKGhn0mO1zD2ha8+WNt
Fs7S+ZsGVO926JFhkQE3nJmwYM4V+1ZGh3qY0Oeh//MLmCjXF7JR7kROnjEu
tjhjdxdMcThWG4WJjBhodMYlXaJ4FLz8puwt8u+S4FbBiK4YMRWJb0cUEU7k
+rkcYpwYXBH8rE3NzrjHBwz6QV7g4UcyjXIHG53jpAMAy9tzgOUM89P1hVlN
1RaujGQBoCamxDiqUI/pC0oPGuFF2ZJJPWjuzGccpU9TbCoWRxLGXOLpPGcn
c3iI9c7fU4iurQVi1tSHXwYNbZ42Z6p93rFrWAJxzS8lQZlxkYs6wlYjvlVM
73KnVr0ZHr2x6JONwMSFe411u08o46XZ6+rIlXPibPZpqv+qZEpwR8ClxRHP
FnhZGEEpux5IQya6ZyZF9UY518edRRrNrL8a2RO2sEZLLFBZdImE1dCvqbbA
XfZAaQtIPWHxTz5MJyrkZwmxxUMcf4b4yBDQ4y5GI4sKf5eu0zMl5C0sjtvu
g9vT0mHBUwvEwpj2dOrOBXxDlVPtmYlyhkbBTwpfe7RBWV551c5ukZBrIUI+
O0+WfzAmpHDsita83DiV5CG4AC814tu5SeEE1qnc2CrLTiblEVAateEfCdj7
BA+jV42OPh/2tbe6qkIztkppHmA6tTHGV8a5qd4fjg4ooJet3CknbNE+r8h7
zZTDOJWo5zlgg7pNxR27/9fIrL7vIPNKwUY6Tzyty8m3WEZjiHIC/mfLpuPc
1FMtqpRJ2tqLJzZso6BuPuorALK+xwstbPAdHG7dSnj8kxhGg36XoCuhbPMK
iT5V6Ev+ui0qDS3N7ui0RgjLbnXGXKLy14nQCZLv4gZBDk8m4x7H4FMr6531
5VCjMvwmzB9NUe+OTKiHS5fzx0KktWYfaoqx1u9yMhnoiAC9qRJw3eAHf7t+
j0wIv5m7Fal2w+H0fabGDSuJTDXVIr8+pwiNC8y2IhSP7RYjX9wwV5tr0rAs
kz8lcGWvwYfBavoTJD1dYkVBha4suBCflmsYfpvW3GRU2Hyt+Eo4QuXGCc8P
ISFdtrrq6xtT07M4necMXUZ8nzxjQQfTXFPY9D1JRx/NsVeyvaNryKXqWuqZ
dDO8AkhjxVPRvy2/mGmg9MWZu48PXijrh2mRknVAhYhTnAJ/ZVg0ipFGcPRi
UlJKa9LizH3A07pL6DQr5g3qvvbbHbCnBU2TCEFsBWXBVsR77Te8wUPavDfL
KVlU2CgKNTqZqMEb4udGlI/fNSWuv7KIW+Rg7Bt3dp94Grxr2Jmd5GERzrKX
rO6zwGom9YJs7gvE/Ulqh7tOB3dm3AeWG8Q4Daq61u8TjgQjyV0GwrkGrIib
VjQtFyJinRpDYZQLiKiYMmLnj3c3wxWjAdmWSFGu9YvG1rPPse5mH4+0/XVS
6NTcLjGJqRtyJtHcpaTmQDHRM4vU93dVOTsjv4xQ9B8DUTOwltjo2rWbLZVf
Xe4K717tJw5feEJumLY1H0cixkJHcErz9j3EdQC0+4OXfQkzNdwGvXpVw77I
Q4ypLfKqWJIfntR9oLL+AUMyFPhgYSwe1cAiduceFu+wcZJJv3TdE2X1z5iu
GirTQ+Kp0EY9mvzhgqNb7AiqIK+u4H9WhjYe+4svZcAg5NAT5ajuS7R2yvVt
Q0B9BuKVFLQl+ocEBXCGzL0Jedp8ah9lMjNlnyNupVC0Kb0bPRzRTGI+GoGu
LlcvgJakbp8lrkUXcLNlC3fcm0tJGYzcjJmjcWwQCGke2fj6GNlH9tios+k6
nidqKFI2cYnFs1xcbiocv3cFA7z9ad8lTUHgds1Y80Y7GvFTYyn73l/RuJwE
uMLRbA8EQmI6TYsY3ipTL/cWAJhGK9AZ+ALBGgcUHAHjh3xoUlKVHhZv/wR/
HMwWmZ/7B5pESEkSSavmfiLCsSh7TD5wEq0buNVf8Yn8kqX4Ro0um3cH9DPl
G7hSzeghQM7hbPl5snlYWc5CMvRtJnSUoQIst//I3FBwhkh/RZYKp+me73SP
RJ/a4ErqA6nCQFvueOflu0QO57vRve/aY0asP7vNZdYxUmGs+BtsW/u6YK0X
tzs8a+PQZFBv/oXA6QtweW3h+gZEqLkTRfiICrriiIn+9EX5DfSRmvNAtQw7
3h89Gig52D6u1kQQekcz8rrAzlEDgSO4rLgsXEvGxBEwp15GSLP1Tj4di2K/
duaGCRYQwfSWpJeiEJLfUx4GbXPPk2etmtF6+7aJu33EiZ3BH2XusOr+R6na
0Wvc9fBSrbvridWImqbnYtwRCG3jk9pIUmIMLuTSytAF+ZCghrXTdLFwN9fm
7dNLp8sM5gGsJXuyav0rPLYL1GiWNIjI9R0a5kaEPlcxIukPEsTSQS6skR//
IP4i6YTjDx5HJPQIZDt+rUaYNA/Fvf2KudPolosN6rqLlm6dq+5qWhifRB19
bYJ6zSqDG2TYreHfH821QqRZqcRA9Gl4aDbrjvyGaCsquYX7DuhEhsS9XguF
dNHSkPrSFIHjdYzObp5DuNWUXoNGiESGgTws+DH7aPR6zRcPi+yHbhiweb+G
3Idd0MSW8SlrCAMZs9JwFyzNKHn8pxuu0EdGVNtfaFv9BDc6HKCQryjPBCHx
ZS+RPFaZwzWCnKrpyHMKYrkhOW+UF6mjtzHbQAI29pfZclUw9w0HoEufDm2V
yu55gVtujnZui2wTktTkBadJBhTP31Fx7HombXfAn4feAEhyecJcBqjoLUdj
bsk4NaETP5/QXeQdFbBoRLQRQRX86AZ2sVIzg7Z6BY+MKDiyuNJH9CzW1CVI
dxhL5ghm+XQoWReZtbS3is0rxsmyqoQ2gl95z46flP5vNK4qJaXZW6ujiHHY
7oMtesj02AFvuv8TeSwPINXHEYfcaH3ukm1jVBOkdCQcSlW3an8gGEO0iB1L
PddroKVTmfT89XSmLCeutzKNN2Y0S9/qlwmES7cP3yhqukUVol2KByPWGn06
zWnKF1MGNYZ6fskKqVUcz9aKnyQtF+roum78nB8p8ZYj4vYUfZZ4vkM6uwq0
REi9JgBtFz4OTdpQxjHAc/r5Ru6mEJKJ1EDFBnd6FOJYQNbzw4JlH+8v2PPF
39NvF5y+YCP9zNOYs2Gtd3TVcAMFTvxhLx6hD0jQSU7SkHXJPKu08yzCLyVC
mB8pQvY6JtZPfnRyidHycq/NB/Yh+znKOVR14CPmTyp5fdBBECs7J5e7SaCg
+kvKn8Gefj7TaSBltjPnDnaFXS3a27xFLU8xTTkhO0kG6gEcXTGAjEbBa4kT
j+KohPaxRKl1QOmLbepeD8DsF/Q239hLlh2B5acTV8lY7tVVeRHGzEDDsvsm
q7fa5ePdT8BpFAyhQDSW/EibNVjn7ukbawMm/0+8qyT38zkBYEQRJ9Hry4O2
dEmIkpkoNZ8QqY3GtxyG0sbAf9qjKcld6pGut4zp9tdXqtJner3QRBHjT44f
YHLohUoaroprw+HPbV9XsaVfapr69cNGl+aP0Shy+rueFd2/1+NOMHp77wfZ
zAXbtvPtiq8ahBwzrc8QLDl9uLQLm2ttxCz5PNZ3w8S6Yp5HwPa+1Wr1yFuL
xlkA+hzyxrrydvroEnt1nJj6YARxSX8l+lJAiMNF0jKf0CCsgibUfnW7B07h
29baPcwe7kw/85HmSGweXvN7ISHtjWdr29MQ9DXs2LtkG4ffflj25cqT0liF
SP5d6HRcyNrF2UzxeM0ciL17h3a4foKCA7Z8iuNFAjdPcAcxy/HKNlmx28Mu
kjwuz+cqupwRP8YpXDOzXJ9du3VJTvGw5QUIzRiln4FxJWiw7/B8HpAlZ+Zi
5c0MH4gtNNE7wJWYy6mymkbkS+lWu9GazC4jKxVpdCoa1Qc/BvkCsn/rAwNw
7Nz1N0lUJu7jMIlU8J4reXrsVo5l+GDjgTXnohQ/XSKh4767vaOxnR9WXQKC
GB6ItINm9XhIYoYyTds5BXvEWzU7O06VmPgOYoNZLbudHw+NkYFhrnRklg5K
GvPm8zUYsjX4CHPqDe3as+yND7ZUAPafBLLuaXc8jvNl7Drtq3fYJEVIzGUH
weHR+9h0K1L4OD8WRBCoWKVWNLcSWCy22d5ap4z3woVWxJW5QqgBTQQh0UDb
nThUp3roPV2K47G27NvTh+AGac0T4R4gtKqrAA5br9s/KD5kBiKMS3L4OWvw
zoSpVzsybpgU+g5unyWEoGbAMsmA8m3V2CnIus48XEPEXdDMfbptrZ63ocEQ
ffKmaFD6e+h7T67qppTB2PXPhZcZtKmx8mpYRl+lgEl001d+nqyvkr0QjAiF
qFK8UG7j5LL4jwZPg6DhFS/SQ0C3H483DqqudheFaBZF9wqh/pmRB7YiR7mJ
Go+F312/HyIJI2WUm/fSz9GGySakLpMA8kpQ/YrNzR3g124SqqCZeFc0Kbqo
pEO407yc19MvCinZ9oerpxjTcbL/Okm2SUrDdsMtWlQyi0DT2o2KhrmEhbRf
7tN2v/rGz/QjnSYXGu2QgT8hrdBH0652F4pW7GL2IPOsGVMCTDy03LhyLSMi
rw0dbgqluBuDVwu+I0DZgHcKqTRPummEJ/CR+vgNo/qm0GDT5Znwr/RbUm7v
h7Wam0fojVwODG6qV9WEr22uISpsZsrdBQBXpkDxE2IP4ldcoGmgVyOIrk85
tk+F2tTDDPkncuj7gVJYOoLQfbjZD+fiTdshMEaHE9pMk19JwWtyUi0AuhiU
NuUgXRwnGIdCJdArUI1+Ls9wJL2uP72rf1loQlQ3oJ13UECWtO3r8t5a6g00
VcpPNnD3pwbDI+04zZmuzsk6QwPgersvqL2soG92hemhn5LK9du0AdErW9cW
Rv6foEWuHV3ygMGZ4ypIUyLwU7C6a2AbFOj08wHbd549S/hE8vUlv9HrGL51
frUxqfcmc/bIwLMp7ZFBoPEHTf3TU9mGjIa8/m3au5m64zs1fDIIZ/uhVyL3
AbKezQP0yNTcyb3XuRr9kQtaNLHU2E0kJ4yZLlINsq9oRFCL83VukiPy07fJ
ZDOHuHNVdpM9EcfHaKaq7BvQuqu1RXJL1ZdUXGQ7ZNA4eVRZqJHg6Z5cd2jB
l/9wplAquVwVNvWL6QODgSaUxdf22OinkhGigD54bJ6NvFMJqC1ZSuBMGRhD
crcCBlEXtAgoHw0q5b77j6W5E4K926LBkXxRVaUzaTLXQz5tNgv2ExnQ/H+A
Rz5J2eJS7jkmszGJgcrZitrjiRIhQbuHiC1iO5H69S2hgzOKCFpCpdlfvLw6
DRzTssPV3bq4meHPon1mxxa5iB4qqWj212W0G5oeRBhomK/6OYWOxjA7aX1d
Kv0JNp1GaX3HWhKNrDYSiqEhbMAB3+XPVgZ4R+w3nIkkJhvVUR02W8jZ0VdH
8c/6P8YuAnsKYmuXNdomErlQ6uo54oovxtc2jN7dhZqRaXkV+5tbGiNxf/0i
jLZRsiwvpm6Jp1tHDosDFyUApkFXh/QLz9tQdBpoGkKi7cX6NkLE4l5HrRYw
qdLJWCdNlyJkKFDO6mxLBdLGPnf7h5GW+J0A6Z4Fpvo2QfyDKQhpRnvaLtk8
p7RkTEJH/uYHvf57vUAoMpfXZOzHuskmFFE8jTJT4HzU4qvn/Y8+pJeNdpeD
qCSNvjsRy+1aSLSY75JplzCNqTqkmoUpC1Z9NkJevJtIt/wcC8+ILapOmkNO
wVAc1YtrBsSLY7mB3hgdAYaBfbpbZpE1IBsCZ608XNQEkG2ZzV3dH/IkpavJ
OMQVOVzSR70WpmX9mSDpYQmXBU+PIqIZkX3Lk4UIqIxAO9VwEdBzaKAfDeao
pElBxg4Urc1kbHsRohc7HOu4INRloiQmuRjl2m/vSwxiRhYG9uaXCa5TOYKj
rgO03Sk8vY75KSMVFA00uRHimz2ut2daUfMXlOte6kKr3Jq+9whYcSwvR3PG
hFcDdeSUEjvTsSSXuAL1bSyjc4VB8ez9bXrFhiUF/nuPVapLp++8s6tslcCs
XHLZeK+VIhrTYgzE1KuczSdUoXbM3PsytvqJf2Wl3v64Bgmbwlz7mE63+RtR
Os9b6xlvMXLOIxh9+bK9AJ63CARQz2QqGvpGAYOVQPhkF4sUKDgVO0aig9Um
ubg0mHklfP+hL1aO40xPr//JjnOm7OkdGTvLQ5700TwjGxSt++uHGJ7j3LqN
DVlLIaRIleuQDX5XAGrRm8Ciq4EdilsFtdWTM0lvJe1HQA59oQNQ5Qk4iDWa
50MoxGSNArSi8Op9HV6BGkK48VX3J5c7UPH6darEBQVMVb8ZhcET0Q+NJA3r
9OlgL9QmCrenFh/KcbmcxkPD96S88Jk+AAtyNNcFZCmj0tRLYGgjumLhgZCx
NpQNrrHVDbCjefhg07F/3Xxaf62LEO+lvZzu+9KtYqbS6aJH9uffdoFY+vAx
hZiejdqe2k9y6xDgqI2AnJqyVt2as/QwX1C1T386e8zwN2e8NKJcUxYmNPKq
TRfOJ6/sZsLWP9jpJgi9Af1RoyNsnAayncA7s4JNU/CCqWnanCFu7gpTMEjK
iuAASApgReLca/dQNGfqvZkP205wZsJX5kXqetGET2nl1Ro7FQUQoAfb3SF+
PdAp4jk2rJXcImYOq4hAfWBHBe79qcBgWD7a3l9rGYcNhOVqTjWEIHXL08kr
07EtGIaTshktgve0ReH9qSr6fEuhit2rPKWpN9AbnPAZZLPql9qpOuUGa1xY
at+jMzDSfi5/mSaA1/+riNxOwFzT+1BC2xmM6S5b59zIUlsSL6lEuYp4lC/f
zGRwDZZHv8LWnb/sASit7uDWq+EPDdsnYvZg+cFK1MiR5sDZLV1wghzM2Z0S
q68TFvVMVz/jRuM70i9b0lwyeOOmL0Fi8WfbHOM9mgwR4dDzsaiqjufAEYN9
pwASHsg9sR/3BI0jLQYvmtXFK16B8xPU4Savb8bEu+X3n9rgzwVy4lvIT3+Q
Rf6BgGqqJf4sPaz/Xhs9bYiH4d28cnBhWddxp430aldgucijsYnKT9mQI7n+
jqAQ9y3liku4kYZwxKw4qw3zmqwP/55pkjWutgrks/iAlcmylshDjg7ft9gW
Z1s+NSDv2QYoHsOnPw3DDAMnS7W+0ROin8eu1W9Gc5/5TIZPoFK6Wfo6yDHj
k+xrCrtllNJVLqDAdgv7ttDKoNPgTw2ZnON69NfKI+XfkpEIq5ue87wFgv+8
78BBvkXkGp7UEWmb0ns4fuaycyzFLkc6UXlFJjEZA5m/yq3Kd7kQX5inK8/O
Xi+4e8gvD/iNtV2p1T4eWtvuxKs35YthyhLtAhTLAvL0X5jlszURw+priEyQ
VQkdvIsHW/N/3JwGSIBTZlv3D+L6sp+nc4mlzLUjMHU15VxEPqEZL27oYlab
Ogd1Iiq2yJ9yexpFzD+9uDO92TYZi32h8gFKrATh58/lSB4wOghmMSF9UqGe
g9WQbvC07/ASOrXfxTu/5SpOmSypoYutR984+AAlJcDuyoSDVechIwBJo3yX
lIOqwvzXHcYELAPqVRTQuQbRsnV1qLR9bd5/gZ7nVt94RkAxwZ1hQIgVKK/f
0lhYAmL45TUPra9FgHNCnE23JcYS4q6lJZGUlNHBV79NdMgcool/iUMaE2yL
gEOr1Yl5XNCEGTbd3+s1eRzG7F/X+U2SusfTL4GoHw/v8uYZk2/jCvm3Cyfh
be4g7K5A9DPNYrPS50BErulZMsRj140c/9tPy1gNJLJ1v5IlhMbXhpCOCtEx
9FGghSRB4KJUnRQinvezm/yUcbiBdYtImb1ZaBeMHbB0KayatiY+J24iZGvc
RK0SGJQ3QOxeka4SFhBu8s4vh+X1Ps6txdtc5Mk5mnE8nXs5kvG78lBe1xBC
4jqxPIODhF/l3pqLHcL3Ppnysh47MnVD9AZkU4mbd/+Jj82g2lyUz19tkmz7
rE+uJTjtPYLb1rfIfwsMNwfZnbWhApX8vF7xBVfEZHnocuZ5d/YdRmR26rbU
7kZ8l5aYlX5/JfcOCyvDtJER4+WxrNojrEjyF/HWuycPphRhwoE/4M7+B6ZV
yQsCyddbg6qKhZC6o9l0vCICIGLsLuPZlJW/Opnnz1S0dQNMK4E44T4a+7Sg
1Un9dFL7tMCGMeDEsqtgTs87ADjiyF7mTThDs3TIdykvV6JYjvtmWjc58Xiq
50g8aK93u9Got8ztgC7TF1AuMlFBJYTg+3HEM7LS+hymHUntGc08gg7FkgL3
u+HmJNVu5jKW36vfZj4B2Ea1YWZPJgjMv6tBbLtBOYVdck3P3m91bp+nza5J
fWOgal9FjuLP2epPfqcBh1PszmEntQCpu4I68eLamtUuR3YoIu7KcXtFMxwQ
sVbvpJogzZr6hsyQjo6a9DuD7odixOi+dVtTkBddu6Opv3znPnBWlmAofS0D
OnDS//2bqVKjnsngl6ZW84bTue+dELiccTUwOhmH5BNc1+7zvq6CSpGjS39X
4C4agCizrtUnPC1ZntQjetcwaJMJsllEyQUEfRGc2MMF34Thv/6fFMUz9GNa
BVzwTmj30v3fDeAxy5gWUg54MqCsU8mfvrUqtLE9Zzs2u0keeIoS5cUMYHpk
nEJG6Tskmt2jeqYpyCGLw5jovvD5blFZh1rYOBVtqTbG3pSCV0Zx1YzABjur
EorBCPp2rMx71i03RxiWOBxdpQj7y7HfriqNTSdM2bd/sbbQZ5v0493J0hjF
uMJ4MimzbpxrRasjqXUIS6zoLO/GIQFSXklZE5AGaOrcth/KmbhIYa2BURjL
fjsRw9CoUGIlbfPrGxETTIh8YV1TVa9+uFRosSzpJogkxWXGSTeUFhpK7KL/
dIofAXZhrG88g5tOr5j01pXuQQ39NDqme42fAHVQ2kOcuWMnTGGp8skTlMOh
F6BRU3Qv49r2WkYAYNHQLvPXb1stURuUgPA5jxF2Od9dZerTLyfKWIyX/XVp
BQrb/fnzlankvFs+smJdpFCjaSaNXfZIOzrp2Da2bhcgZiurIncR+el99S+f
f0oLK+wmlyuV/JeKVNUjKr6HmWvEwMi42OHpLVp4Vaetm/BLcS9Oci28vgll
tny+vGNQBUeW6ksrNIWp2IP2VaW1GoV4nDgTl7L0arGnkV4mBQ9uEVrey5B6
+cVrpIzAHvt8wakIRLzHutikJKLou0jSSm9KJrkmcqoMvJP1kWz4GYU85eUn
oKGWt3OYm2w5c/OENr0J085LkmWJ10OSYKUksfgYnTkHKeQqc4gz+8xpmKGl
J842HXGif9z1tgmzvKloaJYILpdnCprim6ReRmdJlXZ9xrMtrJVd94nf9+ER
kUsj2Bc0bSYQkusc4QvP8LWY2I0JG0lRUFKYC7/njx0sELUEc/7Aj9ZAlB7J
OnzezlTZHd+2ElfeUlI4TA/hQiJL90XlhC0tRZvzcG9VUbAfVr+Yy/gE9Fan
zghAOlLx/t5bsNxMNg+Gm91/A0RD5xt3CDQuhesBqZToYP/lfpoSe8nr3vHP
/0x/C6USDu7xQsCX12YUDjuMNxTd5G7ksJjvgqCxuvyMaqmTwCBuOr0UJep9
NaFfj0V4wWL7ZceILTR4Z9ODesRngNfOFbkpFXchr9cM8x0zEgXgv2VxAFVx
T5JQRcgXHHWYU/3AtieZNfLrj+Rvv5+W+zYEslqYAmwGXBxRUMeJRdaiDWbw
slDXHCZRpqkEMpHt100JOxP8ugT/3EOHZCW4Tc6eHiSZiwvMXGznEpvQJ8wk
bOb+18T2QWpskk9seWl48SdruvOxH4ZNTWDyAcobTFzIOn980MXNGJk7GWM7
2SKz1/FgMDc5EUISec9JgmIMN4vz9peYVLSaU0xokMn7ALRq5ji/pFzWOPpn
/ItShzlF7J/BnQmCGCeuVrlFGtKWXxkevGyBj2dMEo9dGm2KNwcCb+ZRHfb5
m6jUd7j8zyFqRZvJsRDldmzY9oP4WybJTbXSZ/1nJaNGsnM/G8O0HM0OyE++
rcQRWIi2IKeXqBb27/KGXoc3iGehwdbr5gQJh+xjelbFEQfrpS5rSaWM7mZf
k0jZa6V5qkGBMhBvuDv1vj+FcMCQOxQkqk/fCFRl8PLbq1esOiV2ItRFKYOr
kbDACicWdQbZgUfzUWetbt7PHW/0TmPOHYMKc4UamNL1UbPqxlQ+qK+Gzk8w
tmUaf5w3olnzw5l8BGZvl2Uq/QcXddozcmQLKG9jjiIdnQPoKO+HYSDoDwRE
1zn6QPnfwAaOcFpv86Je/ruJUasxNwTXgGVlZ/Rx/QStLmC/EI2zrIOZPA0/
Pm3DbGhyr9uvMhpfx31nLD62LjHDLWy5IhMncQhwrfbTru2rPnda8BVZAfJU
H7q/FbSnx3rjqc1ks2OGaNkPXipq2nf1ySxx+G6Pv+dGru1yT9vo9sGWlnEJ
BCOJ4TZSvP/LK6CfC1z5VX/cth7F85ucdztEF50LbElrhipcpGJyKLHCxuN7
Z5Ky1cjDtXHfdHZaG9wElqsPUd3LGM+d1zFf2ScBh1Spp9SYqlEoRbfIH+HR
v1XREe6OPWgtv78LNoTkZq1K6QiuFUIdXcxvw5cjDNQ+/iThLOS14YxrwSEG
lceQmnSudRm5G/0DYRXQQAOLVQkX1pqdcAiv4/b0YtVGemwQ41flYwEJYTUk
WuSpN1CmWWgIZnEiTcdNblsHIMok/5qsy1zXa+fvc52R7/ARVyuud8Mnort0
wpBORa/yuQB4MCucy+bLWD8fczTNWKU2BEf4UYOkArpO9B9amfDF75l/y/Rr
SzJzGgb+fK1B1axhEy6CxrR4l2MuY4svWxT3vSxrkww7ZW0C+onUwE9/5OIA
dP8/Ykgb3twGLVs1mNKdSDrxy4BcJKZxEYADpZ05+xhUATKFhTPorCHf/P2e
D2AIH07F7+5Rm5goStSutduINcOxdlu1hRP5HVIDhKDut2wpJZb6cmoxSlry
DpFmnTACG/pMRGvtqD1grh5bkDCNpAN120b+MuZ4yW2d9pWz9oBctPSmSqDs
ei7zlFcRVilYDFPyhv2rehJmFRW9g7Sb4AHshJZDWeGZMJrsmx/J8dXPceo4
y55F5JT5MF4jZCDlYHy0dDG4C6BUL7tBXwt8+MXlqRpDK/h9fO2lvDazqgL+
pIsI+6FglU4KvBGdS0bSpx2S2p7qcPqIMiWk2nOprWw2xVELu6EToxA9pmVE
fK7+x/FW+hlY44nQGgPyMFRqHbOngLosrSiWECUg3pZBJIdZ8AISv3MtktQ9
gvgQLmUiCIeuwD8elZI08dc4ZjvuMG4W105uhaQPufgQnUhSPNW8Qs5SXFe8
3OZtM/ZbkWLYVE/OR31gNDvmXxDkbF5i5QbFrgExvlIxcVevfZzfyCCP9HlQ
AO9KI2d4RfVLv9JkbSu/Z5NvIMvmRqrX8wqW95wDWgoLg2o751Gh4pVvwcmh
hevIIKtgdndvVIeTGS2d+d3HOJ94hqvhLw7BEbAGkUe/f0dPx0XXn+nXG4Vo
MrCgaVzo+hmhZcieCWGwQCAsHbsvXEBe2iSLBXsX/u07vhkfuhvInt/rZ71h
Q8VGrPo/5TL5imE7A7GzyilzFI0cfTNKP+fn6aXy4+FoWzKqZcwbD9a4txN0
1qYYw7+zWwXTK62PdSR7qo7QDgp2ybdpHzSbTdWuoSMDdxbNoJsUBkDJMZt4
d9FQfLs4TadxJ2LYjAvKcWiL+AkZ424hk72YlQ6culp62mh5fO2nUXcLnfcH
KbiztGI9GrSFdddQ+ulu+2GT6wb8XrSuMcBjPBtmCJD5YWN1VbRf97ewchIH
QigwY2yOtMk7xlQ5kvtAUoehnhHjggdOaQQqRvBrGIFpPwTIMj2OfIvWlGPj
6RL2iJP6DaF1jrCKtyhpnxwk5zyjS3bHXEgtWlSJyAtVxbXvpLriHS4sKWks
OksKcLM7mUaL1IMX8GmdVQm9QMxLKm8zn19xZ84eo2AxzTezT29RjHIu2iXU
MEcjzBiGEdTEW6eUTKha5YD/Et8/N/HMTYzwz7O5SNBEFt6F9lx4DJoR861D
GaBe19FYlwWJBAGbpaTBV4+U4jnX2SU3KXlY13kON7sBjjch8iMyNNFmKas4
Lv4sFzzb++2IKLdJnmXk9EuO64f3zGmeSGjIAxL/LchXfih+iUwXgDUzTop0
UMI+ZAPBhqmeLyTYLB2KaeR836Py58CHLP6+C+w7L9FQzuArarDp5ojIz3B3
D5qZ1noyVUZWaz/yrsbIjagYRGFzlV1imsICH2WBX/9Q0pS22lstW75S6KGp
N6ZgH7oW1UaMaasnkuv93rdf70MuWm9U3g6NsH4dc9tBLE+Rot5HbEYDivym
la1QH5C86DjggqP075/hu3/kWRFjfUNNHSGHU50sC9O1YKsFcHZBQ5cHNJSL
p7MA05vn5Kru2UqGrf6CxiDsDPW8LBSdfhe2eCJA4Ow8SIxevqed7nJw4wLA
LgE4j954dKKGpsuOoduW0mk/uxFG/GWWDqknQKGYA3Do3HR/6Btu3WlUjkl8
jSpD5fu6k0GSRrVZTifmDHPdv6SGHEkRgdg+3jzTMzjq1r04nIQop4tf2Cbu
J2rYbJqvMaF03yOfXgVPM0k4M1ktcs4OwxOtLBj7h/yu+HqHL8SjHW1/mNaj
3RgtIg3Qrrd+8lT8c0ocdN5jKuFCvntKpHtNdVqWoLTgH162d6rJPugSdGBe
YAmwE9F/8n6tWsG6qMnnT4amF7FJRCn6AFdcKb44QSYB18x1qeICgxfgVfcO
yqAFBPVu9wvVXnIf3dVl1VGbrhEuoMnM+SJFrD3FYmm6rKWgDwhxw9kx2XEz
ojHjuW2KCaXKWGN/KiJ4clxvn01Bz0qXhYabpM/keeqfp3j49OOYqip2xWxW
XL+xwrJq1VLzlI9zT+qFVKvAA0vZ0hDPwNLvCh7ygV83BzzeKhD4Qkdk6XDU
wIQt/1YODIlQrSDpuk0ZB6l0ri0EPtE8O1pDD6/MMzTN5Ae2wgItltdL7Zwu
KqF9rLi6IRRYO63toPj+UQm9omOoc7QhY+WPDHKeCBF5h56XOXha9D0iZx8y
UwL7W/d7K15wZd/rE+IIAjSpzwB9MsBg2GFt6it5y5iEqCm1txEQkdG8qwFY
EVIOt+uyH7iGE1Dcp/eeknJb2B3wKBL+PA/ymItHai0bLXzkIDGYItpiDsXK
TUDLdEnYATLojzLIl1YyCR9w49nf91x5jtFAQ2qJfyueKxUp/J8UoE/BRrka
6hbfJRe2MILEIRPCe+o6J6CTDewsKUl1bRODw/9erg2fNzA1hC9o9zjoyowV
MMzTbYFsB50+oAKo8IqBPSDJsT4bs1KXqWuQ9ioK8zTcd+hl+ilZw2rSmuB4
BrTkgfJJhIsa3Ui4J2yMPDcLkX6I7BNriTjDMGOeEz02KYCExc611QaGWFVo
pcZN46JebE6kGxnBetURh+hwFDGs6DmtdB0TISLNJkLK3rBqTrVPRtm5swDe
cOdmOqF0UzBbXz53Txe9F6GAi9bGioj+0nIutX14LUXXSQQjBru4LHg4ugaG
e8wYXzc32hgABWHRPaIFi3009jPUCfs03aac7Cc1WNt+Z+8cg5IKl7X7Jq6a
kAvuw8r2EUFj1U/Cv0wYBYPCR/dOFdaGjKeV3ka2fTExzMdRJJRun5X5o+LU
dN+BVI7yfiadCjOeoypNi1AmEQbuNPt5eEg6zgJsI0Uir217bWgl1JWTeoLe
sLlMQZOQ5WV60DSS1RyX7aI+QrVtKkL7qdgaVUDI8aV1Ks1GsbZJ0yJ1InCm
TgRHI1aFkpFhQKulaU5zcN6pn2dPdvyXNOao19CAt44AJOb3T1AvvLfFHFQ7
l9aNMPDmdAjoLHxli5Cekp61WkCQ+hPZGReN8D7W57NgQF32sLBWmG18KYBD
SYj6aSenLKDT9rRny+O7pwnQRapLaA8pZ6JNnVRFl3ogM7+Bv9ij/svfi9pv
2A11Y21mu3UmO+ieYveaF1e98qaUBoKQzFTuCp8fm4Bx1nNZBktGyfKiq5lg
G4tIXdAQ0IxWR/fQ5lrwS6VuQoj5fB9yRu+L4eKnZA8v8lqpAMB5Dd/WEqPz
w0c0KP69lVbrmuzSpMtQvyT6C3PlYZKPG/fxL/nwVgs0PAA8JLzSNpD3mktP
UdhirCDjs4eW1rLKftJRTQby7rZls52Isd6XMsSWtnDuWfldN8/eo+/TE2qa
qbMW5ykjgnRHOpYjnf3DTLDx0rjzk5Yn7NJRXQwwSJkboI9Y+Y86h2bvaJQT
IaSare3VbBZxE+4QrRwTQPYys/CtTMzKjaAnuY7pF70xEMtaNL550vFc997m
ZkgsK+TNShoSMQLD5IstFgX7mnN+jDSCrQquFno3d6GPUm9ZEPIeC5l1bqcj
K6XbrNEHZxlqDbeqhxY3dF1TWn9qDojX9DPTTgbQb9fSjTDDYhDx3/b6a50W
hTmeZh/Smapvs6de00VifxOGaA8+MofrdblR3LOZ0yLqbF7//yGf1E8z95Wj
+UuzOkRc72swJMy03ea5AzvWjMEFj+oUrdLnaG6k+bxBnjBCDg3jGGEmD1Rj
tw3Idd+1oK1/2fj2AkZskFKWfutHXzDmznFkGmEMo0ZwfCjdNiFAqMt12WtM
3IUlmDscmKNQGXTgt4ptCyDiVAghNjRSWYLkr6xSDknP3NM344LWFge/NKFg
vnYRr8Zo0GobkrwDxnYrdLQJKk4os59iQvV2VQehD9ewST13i3jWqvQIEwsP
nMEO8mQx8JDa9DCxG5YS2jGWBsJBDgwRpqxio9cKQBWJlatkoISGOgma5Xq5
ULTP+R5LnWPhiQ0xeVdL8hXILRAuTZrcV88yxWqAybDImXjWgU6T5Ai5iVF6
/dNkRe2ybS1QcY8zAdhw3qnqN8d0Qpsq81PP2YePcvcpxPS/4TY2n4eMyO3W
3Zy2GjZgkAAHNdxegiEY6IDBcvhWuuAduMXq3CFTaUsPDuyu7PqYySgZwxwB
eqJzyW1aWmk/SQm4KIYW213nb9qJDmgn64N7DB6QZL2CnEcIQDDVwczGgQyi
XsOIjVJdlv6YKEGoR2sU71BM+NbPDg5ZZwZHD8uDYWZB35vQcDeyIjlq0Pqa
mkWEAnFlr5jOgLLSYVH/Q+lpBpVS1oa5WVl/UU8HWrbHawgLhZVFrmKhMJ3N
WWlGuVqN56SAClD4qOz+2IgvkK7/aveeWipdkninDevoBzjAWYXUvSqDZ4P3
JX1jaWmflPZ96OSXG06pPfgOCTkTSUAfKqQ6ENgs6bsPFoI47s4Qxv90HFvJ
uClbB2m8efFWWdDmuRtuAYe8quIvOHDhN0dL0L3/0A9siJppVanUZw6xLehg
moPwvlZvxuAwknXUCoTFij8mP17+wa4l4DRMZnhKywQwZlZHa/P8bAQmqKYZ
1pzjVdIBrspFg8I6y2jjG/u4HN9gyiTQ4KmsoG8OjzPhn+BvSTJXsh7qWjex
d8N7jrhIZUMewRr4jrI+ioUawiWBsCFrvXK3YX/TT+GRa626MQbZr+KYLQuf
Dk0FcuoBFSt75CEytWdS/aaqoMHlwlHbX0iiUwyyXzoM0McNbvq/HQC9+Met
UOZ6fPeQ1ZUS4Effe2RhbAOB2lTRD+bMYAiYbz1Ty771ncj0K8wWkNwa4Es9
L5UMdnElV/DOhuEi30+JjTfs+oVDyXcGNSSqrQt8XAHAORxAtC8O+/TRV6tO
gqOs+7aN/9/xaNMioKJrSKoANOLsSwLQ0z8rrNS+hukQ3AlEhHPyJy4eyNjy
92FSTcYrt2o+9zTb1oRrdeLa1fBjxvHOPI/hnsA16O52QwChNIKb6Wxu3FTC
1JUL9Ruj/QQcT5x2hreSG+7CghhlRoLE6W0slniesfZ4JnY64bU8y40umnBt
dEzK16R4D1egFHuKkJZZ4pulBHj8BYAJryz1tF9P7sc9XNtc8UtzfqPHFnX6
1gzbuXTHDJduDw9AWM+kVYAdb0UJNM8hIsB2KPTxrWPtuyXFIH3ZXHsiPn9V
zpgC+FWHru6fgirdz9Pey8tDr1d32I4/bDO9d+zbqjNnWDIiAzPRTmgP/d0w
6Nkfyps5xaXc4GP2/REku6/BLN7lHaj8sdSaOxiDuLGZrQOpEndB4ZPenodt
J6BqduDxtXyZxHWS/EHmN9TImpiuPPhJG7d2mznu0EECB8fJJdl45MZuXEQl
mk5lo8v06H1Cm/5WB5npBnlcf5h1bna5Uf/wt8FFLrFm2ZfqVB0Un52wGLSz
yw+rU/j3UpXSG95tskPR6DeU0cGkIcs1BVZuPEtCdK8Vbi+LhStsOUa6owJe
EQNc90lTcxiEd43DSunKbwaTZUBH4OJQl6LeOVRgE2GykZ32FFhUe4FpiF/o
v2aPdFHqxKkUqq9y8WQ1vMn3DGA3jCY9GMFkbK6uTWPa+Jz8eO6jo/WucNIu
V97VQ8edaQQLZCt+5uQ8f/GtDSHXX7N+ceYVpxeYZmaMyvJCBko2SM3Y3X8g
LWORsGsA03qCJuSA5qBhSLFW6lvxDM13nlLIHuUsp+ypCN4xU/p+ug+WPbhK
ZzrN4/1zF+GdRQ3Hdt1o7aqXVxLTk4FHkM4AtyCM+CwgZApyJfF03KG1lQj7
XuSfi9pErvMYJBQUG+GMuWW8ZvRNmom6miUKvw4UzS5HE7Mz1nE8T2E40794
QUTz0jZQNcRdR+hTYWixkeAVQDcsT7hf/tu7+f/gb3JrSNYjiMKbOWr8s93b
ZpKBx9edbaaFoGymdAdE0z3pAU2RkgSc+8oQ78EDc2qrCTn8C2CJe7A5WRKJ
utsa/egyQofFNLxY66TqiueBsh0Q/3DP03y2eFCMjFQ17dPVFnyD8GWvhk2Y
6ou3aCHRhsBgbFGid6cjbDuiUhlWR5+L7PQ+16tzKHvog9G8OGNegf2gLSIb
LiakQkhkDXXWKjtd0UadjRM/U9YaK/qZi0HxrnG2DiCkuzrx93W2HPhqb191
PleuIzKjh/y7eInaDu6nRnoSj0AjEqXJeBFZMZLJEQ5TbJcWjrcQGxtvrf3C
yaS5Vjbe+oGvlIsfsb/Iq2DLR1MCMhMBoQLmByDA5wwQ18HxjGJxuXx1Mt1R
nDJpv5KgSBdkiYYOyreOHN7FScOH4Rgk/rzvt87sPwyIwUw8hDpJZqbNzCS+
8SPw8o48KFG+yrtt75jAvfUND63TDxw928JEt4Ox03Pzg7SYUp4F1YiDjyBN
sw00yl+XS91fIdte+o75JX3dzZ4m9xZOv37zuiyFaNf1yo1T/OsIbcD1BcE4
Q2vtetwUM6oxQ55SGPlT+jGsanO2bOkoCODhEfmMdzVYeWPwvH4+iVlknCwx
yOlf0MyJU77I4J3aQugECiy5DfLcYIKoF9L3s7+ojLccV/RVe8/ICVGeV+ak
fkKkIhYF7GhIq03ByiHe2mHIO5DyCPhK83wTY1UAxy3qkMZGGvdODb+XQoUF
je7UgYP2IjIG/+vWDhjyU+aTBjZsFvycKYldlBp0BsROguZSfRvBTQMqvdnj
z2ne4xMaxTkht3BxJjf9UanDbgdMpKsstEe5KMTac3F4flGoLn0BnL5I/uLu
TS5TCVIq0AE/8eibIwVOaiZzWB8lLuphiqCfIWRFkHRzLB+Kw6c5QaGgWGWe
vxb6xmBavefCSil4lrQbZs5AI+ASj+43QBr/b9nUPTYzIa9RLy0ezTdIhSkG
cYVgldw3QAxOTsDuBPG1yusiemgQju4gMOQSOIJtk9AxrdGMqV1K1zZk4yDb
cJBf49sZbZfIhzwfJv97K+vm7IFaxTxWvpulGIdjaopvhz0Q0InTFRhl8ck7
3plfjzsOOmheBkEk1TdhDWUxw1y6fGLt6f0iZsNmAU56THnZPki7NrS3PhPi
2E3C+sar0ZpT+SgJ8qSEH1UzmffSmVT/Hbf0AqywcuyJf98e22ye4bHyeILB
SAn5MHxWeF7dboHa0rXns08R7pSQXjx9peV9CX7HH1627QqtdxqptuksQ8hV
rSJrZ42KJu9vZUfbOOGlluGQEui+uLnQsWX3P9psQAgOqpCBu/XRnvVeQ/fy
w18/GrzqhQkmT322D1F/ApcrQQt3HWPHYlSxI039cp20WXs3pjXwCBrTtYuZ
x5eaebs6oNfY1wVTAc/lcl0jXVa6KP8KM6rrvt8Jmecto+gA5gqKF/jCBiq4
DaXQNgZufBwZOCQUeS3pJykMcYREl5Hf2zWlHMiCWdso42Hwy9Nu+dLrloA3
0kULG19ZQuw7PQaaP3lv+hEQxRRM/82/8Dblin0u2yNPvzh/CikVCU5nr4x+
lXJyUghXnzSijCxwqE29I+XlD+3z50Z7CCUTaOey4lkoYVmV+v8wVFzpos7B
tkGgmN+uEaCbWpfB5H+xN/RDGxKUBWgJGHfM1YXYRpjceRObw4qKIF2wgQKh
UsCYRi8hMzW7OSvQ2sYt8V0D91MfcMgd4TSK8RUYe5h8GkydTi4vQP0Y6o3b
GQlvaNFbMIK/qgHdLzaT6KyxcFBBSReW04OGAzVRhNcd6nkB5ZZXl7YfGr+6
GCJl8nVVV0pakRu89DgyCiU6o7S5+6SZlFbeLgUUXKyevc0QphzhLQsTsIXi
ChtFuhRblrONYurGeVxxI6T9pUi7TBmdwFV4w+h98dq88hsymF3BfdEOtwTP
CkVq/i10kZhn7lRhSMrpZ79OjysHHNjPa7uZNLm8NTDTK55vTX0Wry+Abu3M
qU7wlAjqsOG3Hkw2Fqquks+VAhJypNStGrxYaoqahdsKq5JKSmQZyv8QlwuY
slRPYXTbJFJZsIQqdhnWGoR84U8UYpf2mm7YZndQfRrGIlvlHBq1PD3eIPOI
kM1Hm6fbPNvLcQWsTGdtF/E0OTw+4rezExmdRe6VAQlPzFCZVkiSBwU4Bbm6
0T/HWvLnpRTVQOqrvt7xmGrcTqk8C60VPqeU7l5hjklLkgv7rrj8yiNJS8uZ
sL8qGkQTgWfqBa20MFuSW035bb0aiCMsGx4jyCzc+ILgDgEw4IS0ZDPj5+Ks
SwCH2xW8Lkhsom87t5KiDl4NCJtxfdY5k7QmwbPE9GkR41B2LaKyfSnvv4fK
BItbWo0Ow8kHcYh+vpWbOE6LO3XqngPwbYXoNmxM8R5vVU+RT8q2P2AMpk91
7zfigp9GtkUGCAk3zkp/yNNPqvhRgXzOma2TGgNHdw56nfOo2Q0BAnsrwC0+
p/pFK22MjK+GjXT7VjWvMgsQleN8JFnnS5ogR+bpn3TzNS1HHQlALbS5lfZo
ath5u24+r6ODq63FmiWhbFavKhyAcVhZXP8MFRe5whO63QAIAYH53m5qplUw
cly9tqkkNQnQ7ld68Qe5Qrj+czTz2F2yPzLjipOgY1sHAC/4t9RK43HjV2Ji
L048pcbmpNpY9Ms9BunMI3nKfaJCCf50uhm3MSCQQhhRcYVGnMFXq2oWJxnN
qyeGxVM8L8rAV/eFZT7y2Pw7TGig5sUGkYjbcStDaVb/9J6ImNLyFKxiNe3i
u7SeNPhRLIufhxa7QDFJfKa8utVpTVifVT0ASMOpJmPQhfMGVwB/GWJeiaf4
HBPzgbZwnOLAEhKh4+Kw4+CWSTa7qtPysHlG3ty90BO8z+bhc8NMnn+2PQlJ
yXuSdurub6ZBzB0hqyGLkswPreyzR3McVn9Sf3fxtRbcGySoNzp+/11MzDK2
swD74duGZQI5gyfFgosfhS84p5VjKamDkpMgPdC3TlKlfi4nxRuQ5W7omtmE
xnMeO5IdTiCVlhNKZe/wNB6I1lJveX/IA4wJp5wynn2oumr1b13rBdvGbtVN
5skLMsP/cmcf6cAO5rFlHFxZQTY1SuP2Xzq7p9/8GtRI9GLtZakqG6g33jRA
p5es6La2pGJECOeQR++TE6esrky5guHFY0u0kvRNjLetpEsiRt/lBr5+OM4N
YHUWBRNWUYUV13Kx0OHFjhHiPUcahJ6K9L9sbqzlGXcL1kC7P/uf9rO0M67w
KNW8NCyEpRyuOpWkVT5VVepufXL3puX43rS/nzcm8xePiMIDDi6jDhCLUEoo
rdpCsnXV52u4BpGCKUY4tzTpoF9vszXYjkNC668pVBsrvy/QpggPYBTNb1e3
yd8UD6qdubjsowQ7nCL3dHaLlcqmkBkws9kLImdjO4bjaWsgvpd2QDOXEs79
WMs6lAavvh+Jc4kKLGVSnlrPze7rDnRu9+nU/3ss7BI2LiaGYeIj3Jm4Yasj
gx0Cx+o0LO+gKZhGuKxiLc4kk947jD86AzMSlfg9G8itH+OLx3mBLmbTtnWO
gCuesg6YpmajYZOIQ5sUW9CyxZ1g7JPmKGjPFhWSEfsYHoW40Lxv70SBkqPn
hfM176+L84yl1V78YRF7InyLqR3KVBfrMHvms/8zfrOik7qnwfQfI/51Nb2c
ev3M8Z6lg+wj005w943rZW8XWVROFMiVeG2uHZG/sBFHiBVUpBVIq36Yedtx
cuMJXY7+GZaxZEGaLIsXlqWEKFojh/o6AfVq0lgK8GIILTj6fHGlsn9kvcg9
M/jrTZgyG0VN/PYGKBdNcZjSsoUAFg68K9qARNSSE5d9mYgS92YFGwezCHus
VSQKD5g4WHygv8tj2zPiQYOFR6uxskRUzrPm3w7cjMYiay5sYdNw4CnNehiB
3HZPiMhgFeH/bAYX86lUU5Z3U/pt+9Phv7yj50VL1FberLv9ue8gijqUOfzn
QBYeTqVirXIoGGCOjCmyGLcO358bIgJtZ7UgHi9h9BHBMQhWIRjAx9TfVvrk
BnrFrce89doTN9iuC3EZUqu2DkzaMjwvpY87kvUbNoRmjobVbAyFXyqi8oNc
UmEdTxGfbCkBGHM9AJYdtP2ycOfaEzmOkACzGbfoTyyKshyCmH82ok197H2C
aEUjniY/3bZvrU8KY0c9kKErKYCFzbkciqnOQ+ycGLaLmDzTI8W+HRstU7be
8IBBIaMdTFQnGxT6ROsWVC73jSXjqmf9pYBG1EcIps9xEEjkpSK15xYrZng8
sb4w4y7g45Av4fDcOvxFOOMgPap7H9DVxlMPpLlLzU0LbIn+lPYDZHjsdMTM
fGbbHuOomJix7Hc8D3Oadh+SFctGXQ7AFpoIofpWu2TzDFFFIu2UX56/H4s4
HvEeAr9B0bYfs29Yj1z2N2DuC/QgzfAZNJNZEGC1KXVtw/j1q0msGFACcyj0
V56Ik8ZhadNTuacTqJz237LMqI9bAsBZFuz81A98qFvu66Pbx+L/XdwNvrrL
6s+JftQI/j1zQyunxK9MxPwMFxszoFFVuQ980rKIxyZPM3K5l7NXjTFOgukS
nKyn/oDmyUXXIWFBs4AE5x8eAcv6OR1B3kB+IQ8SH7swvLfAL3SKy5emq2s7
zC+kaqjkEobT//x6ytCFTHkQOSC6CXbrcP0vIKwxdv+V+FChYi0YJG7jt+vP
RHiw5iMLba2k4gBsgEMrs+fFR8CDwtUM8fmf3SOmMO0QGEmla1I/gk606B3D
IDC/SYW4dHZLrZeF4VFrwrlG8tAj6rGDJBVSFIaj17R0Wc/bo6yhqMREQNGP
xHHpEwBVpWZPQ+jvj15SpWBtw4Te8CnL9QEFesuRG/+CZD66mg4P8YMJnPRc
mm+M+DPzTPvjqUfZTLFrTTNiZWj9CCb5Lkod7GABTlYMOK+m6L83nlpDVVsI
m68cTEupfDa5ILsHWesgz3VDVt57XKl/Oj/LCVoRf9yzJ25qrEFmWIFtXatQ
k6MmW6Jq3rn4BLMtZXvo2YhSp7ebAE8D+dqOTdamrxr5ZTPLv1gGudjibvz4
j0oqM+NYMSdQb7bCgDDl6EIGmKGbQuZvMetiiTbHsZThVx8zFCpT7pN/GcDj
CMPzMY5O1kPdBr9DZhqdZ6i6lndW+/nfz66S9frkWx4Jt4HcM7oBLhBSn+X8
qAO+fUvhOtIJrRY62HWS4i0Ox83ivvid704Qxc52i6FBUWXkTacyHhYsfVWO
/HIC1tBm3u7aTs6IEBNPQrSmfvRx6np+frN+hGiNip3zkdvFkPHVzClFkhGh
nikwv5+TdlgVSCxpvSXjfHo1aibqIqjHlu4cB4W00HC3jAfsa+1LoJZwtLV7
MRcLg0h03RrFx0nmwwtn3IctnsR5SPlDUhS7UdcYFkYrnv+fq5bOBPjAJAoE
ZcHACAGe6yRFhugqMc9yfzbNz9ivOQAfZd7S+hfAZ6NmMfZUfv3yj1Fx5kBZ
6KWyDTgkzpFczekPLYTJ3CUD5ZXPVY0axh4pYO9b+STbRo/mQVDEO+TeF3Eb
O1ju71Wuzhf18bmJx2CRroNEh1p6FhJtIBPNu+ttA8BXk9w99sl8ZVXBTIFe
Xuaa6t6z+7cotV4LKtdoWRDD9Qeds17BH/5tjdvM3AyDw0EC1mv0+AoBMdly
PSMgIgWaFMG7piE8z63oExBB8hSu4ry9b3cx6QferGdg/0zNwVVR5FXQnsWk
oUVr5ZTBJR6O9DQtdjMNdgYwVcDDmxfas34XK7834bS8yMgsvqAU2uSzG3yS
PVNNjEUmy0/Sd0NMdHW3XitdNBZLstUoyxTlcuf7WDtpMYpkuFIF2eCho8G5
36mJ5NpxsBKaSxtAwhPdmK3eCQWugnc1+5LdLaJPiip7HUhjolSfcKpY7POq
lNxMt5t835K0IWh4aPAnqsVsiD7cL/CpjJ76A5IOW6yAzRrrLjyN/brHGMbE
huiSusnyqj9P5AxrXfK5iYmVOYZrLxL4qFQaWyX42q7Yxok4RKEF1cl+QLnZ
jz2PTGBU0RDgl2iwIcPstW1hFMN+MOKFpzMZFa2Atj12yaSsZRr3K7teX790
al/blH4CerDCzBBaEH73GhC9ca+8UYzf7fhb8/jQ+oYcuOGG5y6uv6mEOVAy
MahdEaE+e8bDRLrTNuwZgwx0VTQYtdcQffBDRq5/371SYWnwdCbcHeXB17od
iE7OHxGpmgF+nt1ZeHK78iRgCAxyITfSBp8A66Gy+RA0E+IxSBNzKsvZw0cj
Vfyhh/te1RUwikYtnEI9NLhsq4NA0c26vverLBUag7Q286XzsfKvlkxRvRd+
8MqULjLu7o/rJQQ0C4sXP8iQkVJ5Gc0wnSXV5AWOC0mKwRsaQzorh7fvQUv/
OqgF1lgPVkpt4+YHi2pL4W8nnttG8wfGnRGQC5snbmPxWzWZaxiw51FgrEYs
uS8Z1TQlAZGHIfhfnh4GRGDE5GzOOujRwdHZuSAv/ecwkFrHnhniIpEASlqe
eAUBFhu+30WHNm2VpnaBrhh2Yh3TUVvMk20Jn9jcPNyWJVtFNPpMcjBwvmWM
+K7rV3bx3mPEthNYh1meYr53GJKawPN5rJFv6YlbLlHauZWIJX4TkBbAvJYB
AsrVTu9eupQnILNXJA6BXCHqek1HNDCcEHKw0hQEtEtbuZIYKoDODcRWOuXo
8aoeyH9+pLhMsYUDgCPJFZuKuUTtOiLaK4xecmYxoBIklmsTd4aa405Ym+gM
QMtQHgv/C4VvgeWrsODUfIQ0HuYDmMaQSx1T6Tebs0EbEmxXmpGzTLhwS28j
/dKmGR8wqq62JbJR1okaBix0iPBYzIjVf5kUuet03G8zy9df8R3+GeyiGxlX
SDDKGgqhhMB42UEMiJtLTBHLFN5jOw4z1HjyC3vQ8H6J75L944pZ6T/3RR9f
1hDgZAINVVoNo+ZsRe/Az3fRgNrU7YGr9JYH9YuYwVvfYrybflfo2+gZ8mqx
Te6/XpkDjOHsJ54EDDyKLbF7BfXoQXFvekxTKb0FEno8OG179Pey4Gs04WxW
/WysLiC2Ttnt0fhtsLyjcFWmfjb67OQKSImomef/kqZYgGTvhA33mxWGzVCj
d22NLbIavMhjKuli381fD7QsmuNoldrlfOTppYKrkHboQRgelJ4pcMNMKUTK
8vXfONS9uHX3P+JfWFewxnoYOqcFAOkD5jQcrUhNHaNfLXFR3Y+vYdcJ+Phk
7EZp6n5w0OtyaPg7jq6IqL1FTz/OBN8TIH8tyGxIY5dg+tkbGQx52Vb5TqLW
CvR6OibnJmu6bIbYSpdm0v+v6++b/M4k1knAMN0V4CJe0ilp96mTbXltm/TB
AOsaBe/RB1pOK0qi00mMtr32O+8VUkmtSYvRrwQPdXHLDh3weC/alofRHfEn
7ZDXulnsMrQMt5ZKifJDU7zsnPCz81YPCoB4Y55iOkzKZUqPLQ8yByGFOkVn
+65Itupvzg/8qESZR0VZ18nnjUexZJskxGveR6J4yzoyC434nQUBPK9mVln+
8XcJ2H/olUTqyJz2qYM/4QHXI/k2n8D6GL8G/5BN4jgriOyYfZI4D/klY7fv
HA7yYh4HxGwOIGUilPmCz+gB9v70L4p7/Fzy4PfmJi3FGx0ueOy8Rhh/SAyL
UGtwLvMYpn4vKX+2BLZv29MYeQ/5vhovWDn3c+ebjXjG5ABzXBT8rK/BqPZ0
uzc4z5iDVP6NsjgkoyzisH3x4lCaZXhWTPrAoK4LJ9tAXAnOp9qlhzo22Dt7
oiQhMxFIXsC5CSw0B/Pp1FNg9Eb52Oy2133oMhoCtLFnq5gti8+80YLXm249
BIMdxAyuP0QbS8kuk2RkvnT2sj2aCwZNjVOt2m+zaN9tUv+KqE5sI3AglZ1s
rOcYQJb/Cpme1uJyo9/cdFbwPqG6InDPjKLL5MSeJuAXbIpQ7Uhns2W2OG8b
rtQKLGOA7kJHE6MY/hnJEvh3ntlKAuageSKUS4a4phczCedXXG0od3LdHFL9
tcfZl3fmT9WwUjihgIgMIWW5eP3x2Uw53l0k5dY51GwTCuQcvEPyHH3uEWxs
ljXsFejmnJ9zd8oSokS4Da5vGs37YaK30a7h/ZUc4JlJHd8cY1mnGqx81Ld5
aDAwlb6UZX6eeiuzO5UksXPljGFDfQ5JGa1fUs9nXLqM2FH1e+v62/wvRsh3
PMbL4bQdS8JzY85Vyx2ik/e+uYzPDdhTlsZ7h211Ov0JoIcJf4nFJr6IiOaH
Tu6FfRVOOaUJkvwbnG03Q016S0w1ZmW4YymEwbdq2xKwZ2Efxmzef3L/gaCJ
/ZbfnF1pdEv7gp/092/Wmamvco2Yr+IXHakKJIByy2ZKI3UX0eTcWdh4BIgf
tkJSGcMkIaQbFgIs5UlR7OryKRn7hA4wF3eypDBU+kx/JEKbCNf1iHB0t7oK
nOTfa0l78Pg7PjhX21dLaz+6Mr+ZxrhNhBwp/TmKQSom95OEQw69nLqIBJ3O
4hCKrI/73n7QbflP4sxmaSGGiLVDXD+C6WtRlWmv28VWc/EcTpDSgFh8b9b9
DKp/gzHEnMvCE17A7zSrcBF34JpVwV4h1p5Ddz9SI6SglDBOqsmksn0LSSJb
Txg6bbl3BRE2kGOTA9EQ8LjBuNkjPGlF7PsYrin/He0endGWDikxxc2m6lY7
AlgBQ9dneOuhd+XWNGsdl/QeDRXAFfsvHTjUxno1LEBzGGxKZPHCA+qqcebl
lgp9s1bw5bema6jUVyCimQ2fXur86NAGg+OwjRvK7G3BchQL+gzKrOs0wZG+
yGOUj4aBUHxafETE/2O1MkGbJUJLhYS9E3njGfJ8CP6Pbg7zq+6G/RAJQSOS
al7R7p8wUr+Rl16U8Mwnroe6wAfVMLXxGhatxHvcLjBSygsfGxxhsTU+650E
WItSk9abS/FJ+bFLRDJQAc5ZkDO2+nQSUxXP+4IgLldcIhVP1MPO9ENMS2da
+Qy7bnj9/hMFBbRNs44t1uSmJ6z/2HBbUmYzqlC6WE1QF4eMhOC/iIafLsgD
hM1mFHxXVrB25tOyDJPxGAgJNgpK3oo4fiz0HFkBqzzCRB3YOWg8JrqdjS2h
Gv2OSAp+uGTL4yHFe0hmI58vEyeKVXMOZ4zgtJ3PMIK0odq9onHx8KOKvfm2
exez3WRzbe3ZvkaeHvCBCzj63PX2TvGkHy9U8nL58oEtLQsMKXDJQxWEYERH
HBrtgdCUHKvN/uu/e/xPNIQsf2FVKnkaRQsOsnkyTEv86eaphdkVIJXSDPd+
5FY53aZvICBkQhycG7LS1/16F4je28LI8XG9gWX8D104lWFV0VsU44ipviiR
K9UPFlTYj8DUucHPwCP695DjiTIpLxUqsiV0z6ZGHlCWJFNO6zoBxQi3EShm
oc0KfnfDF+VW86AkDivIc6WK8hCjAqovTtT2vbywx8Cm3xpDHFwFYZKmsPHU
6etpRFnvKacymQNxNlLU2YwjzsaeTe/ylPLp6rtTS33APuyYqB6nH39tOPJF
aQukP+bxRDMauhVh38dhql3osgV9qnioaV64yMmnPIcnTEArKkAK4Flx9ku4
U3BUPi59TEIm0a5qxr2QgXxe/Dr08PFgudFvW3WsCV91EDbj01E560AWjrX9
PrfOz26/WXfg+5AdlyniKx00x2bEK4eiUhYh1oFS4b+/SDp+D5SFLkv4SC31
41ci2d6/HSzwd1IE0J/BBG8piHBdmUS1bBXj/fwzptSWQAnuGpZOaJYJ6CFa
gzJ4rxhvbzEAYcRmNSMQXxX44llqtWRZIGTMvzgMHEVmqPgpPwU200kEYa9Q
aaO96U+zfxBvUvAu1fzeeQZ/P6vxFH8suSjnz9P5iIvri6EjCYy/c3mjla2X
j1WBW+Qbsai7+J/xJLgMuo27pNMr3BryzeLpUPsk+KnAKeksonfJJTtmyWAB
7QvkUo4qsy+tPxZVVH+eFHgRBm632fdxzGEpttprrF6UT+R5l31p2tAtPlGo
N/BmbHSqRnuWbXW+He7cMyZXkUtCutYfRB/qUM0iepvcap8obg+AqKbE/R35
d8fYScoqgntZTXugOC/knqNURaQclalXW9ODCZA57vZjhfh3+VC9X63fDd/9
LyDCYcOsMt9HhLssnwDopuBmTkADFM7tQ8E27dQT0OHirzBQfiOYUV/GN5B8
kxE9BBoo+BYrhT1W6Rt/kKKGAtXI6xD8dn6FBfGFwb0AI5zc54/8oAXhZEUK
BIr/v0xgJOibnNRz5lsn0G+nrhG6QtT2fU2UPxJb0Wm8AhxCQCP1fsdYz4gd
ljW82IIcyA9QEfevMmI9seTrSOYYIuUHQao3fEMjxoTXZpNOr1zfTcXF3+CA
T9K8NGlWDJclrjLxnJQ1jOFAdEfXiyygxiBvyCHMdt0SOmJMGS8nqIPyVMb8
v6qsvqPJj4cGsdhNBedPpMo6D8LhRREq/d72D5b3sRzpBnAQTbgc+xeL0gnr
sv54+a9ZU9nrx11uHc/amhV/sMk8Ecg/nYjbrB7b0Kpxj75/Z4xAKSzIPHtH
DBsCpZIJx3FglNGXaxhldcd3awklL7jfBsgGT0NqQDGQSJH8ynfeWH9La/B7
vBJtAFukYRr19TXeIy3WpeMvK12IJWjr82BHUp2Fl07c/M24bly17PyCMnu7
Z5Nr76U1ft6Hua8T8eA3UUy6Ui3rdi076RHD2m6j1QNB6EwCsIxp79sUoA3a
ReiLZWeioNBrSPTC4E6l7OB9iz+RdeZypoIqUFF9nmBhMraGYXNfgZfEdBk1
lT4iAOcMHciEeJjFvXem2AAMDgHADvGq2voQFvBytNC0XfMYDVY7OwiGNqPH
CK58IX0ecOFXu7ubkko2QCQ1I/xLjFOosXTMpnpLR3+OJU0RFq9kNdVSkrfd
XGX9FuAhamPIkVh1sGw4MTJwFQa+DHfj5DPS6xVPBlS16lai701Gd/JouBU4
5L4Q3gVlEyM1W6h6yp9Kmnu8dPt51Khl+mbEwkS6R2sfcjF/zaDeVPG6urPa
3wJBdoY4LegSjIXHMebPip7otxkM2S3aQIo0RWP16D24I3Ad7q9M15KXvx/e
t1MYgMZEJzThrzx94iRCMitZvTGRW5WsFnFC+58UoQstAtpRKmS4UAUQbuxl
QDVIW1uSiSEy/w5ZSbBeN3MsTbJgow+Fq/OP9aZp2UjWJ+n8wMZwSVZISWEp
Cl5XE4THWkKTigKSeWMPR8eY+0oecWHHiuzg9niVWpQnM8QmN36sf07YWdx6
ciA+I680Pak7VL9YhZQLrKJ5XlI+Qh5TvsWzALNrg0cFHfta85KZMrWswLuE
/WAPI1DP+bHKKS0aT9iurUYZsZrTBaYZu/lZ3xHFB9xt8+p3D++kvKRzwPrT
XLxcKeU98C896X5QBRcCzZF8Ktn+qbyHG/ISBD1TKt5ho4/v4lUd3MgBDtDC
9uoaMu8/FGA1dDkfFUmOWi3I8w2wfXGnT6u1jynJ2w03Yqn4AxbsOU5+vZlL
s/liOgtqKGHoiJ6WwGxIayQZ5UwCW6+UXez/pn2bHU9mAzFODCVoJfG4rpWA
XTG/bPeFPlj6FIzn2IBwTH9ZI/cBdBrwPqk4+jFJ+bjqVjCeK3U4j7IeIPFF
m/GwzSJH3ztRsZdis/TLBpR8I3lAD7OsfMk0RN2w6IhflLjfNudugkFHYhqA
+qNYD4RV/D6Ke1uzHjB93Yut+71SUYPxJVOAO7R0fTKV+mbyyFo6U8L44RMo
HrUzJjJ3dwjfUpGafrXCOjxQ7hB1xBbkIDrvxaiKQrZEOOlZeRoE+FevO1eO
8w7Mv8VlIOTDKwBpsxcvFi3APM/yvu7xbPWyTwvkgQz1iFEx8ZzXJ26SDVbF
uBsTOogmqVwRsCjmd84w5UgUskX4Y92da4kbhmMAeku3O2TFZcozY3cN+4tm
kFc7emDkNI0nFZTXZtwKC+gKSAGRqxxgOY3Pme0aKDO4Fl+HlrfoAZXLiKiU
jDRdCQO2rD5qohB/YFGzueZWdv6re3m4BU0lb0JhrBPcNLwN+jQvNcN6p66A
5v+tJar0fnmcOto+afi4hCONJQHK4IiUvQK7z1YiYUlJjw+6EuNLQ5U76eCT
w1OFoysiK4mqcj0t9MKKvERgUCXCDgnJGtp+tbZqTk/16QN+54J7uxvDascM
BC8QtfJ0akV2j0v+xVI7sp9/uP3aKuuxIg0n+Si3D8289LBIFfCakc4E3hwr
78BoyfRx7Zm7H39c+oFsSaMJqNNM4NQ5XALPZGzBK2by9tue2z6sg77DNiXw
paY+YiV5PqrrrEjYP6o/Qc8nH7nOrIkG8eHH+SdZqI/+EoBXiNSmmh1NaKAJ
tz2SDJsbHf5us+f0TK3oCytyxFrVEdRlLOkiy0iZYxpihrLh3IHlXSr+xb/g
IpPlTpB4saCJYqfCmTFtgVHY+SxhFsPIG9EfJAic4gUEWEXwip0jBZYy9N4D
ZbU5y7ashXcrR7E3i5WN1e6UDkXldrFBFnwjOyQ31YJ1TKtxzIrBz9QgdHTH
jGcwMQBbpoiLYBztCSkrWdw04dON6DBU7d8jp8OzflyFiv8GEP0ANIhyXP03
mGpWIlkiEPk3p+N1DagPnfYeWvlD7dd2E1TGeZ0moRUOrtvcJ3/g4Ec9OfAg
BtoP0FAU9MzyqylVjBnDauCD2Z7xqkuZxUFzIFgVGLJVZEe5NKIQACYdjinx
GBytflWpqyUs7iyb8TCp6DkVfs/JR+DZdRgMQp6rcb8GRlOTwCPp5Y1+2Tbq
JZMhIskkGa6pPIr/SZ9prcGHQ3bheJ50EFyNNiNPEhwIN1ikxJdDk00jARtv
prz4Wl4gz8XSqubKh1sbu76luFYSXcrp0fIKUFhMk4sY6DCTKCq4xPI9xm0P
LF5XVZkwPk5CcgecRGt6gCvM5KLEaKVxzAjbza3NAeBNSt/34aE+Zp4yIRKR
8YSUIe396vwCY2mOfCSk8Fr2ce4tha9mAv6et7Wl4cP9ZMm0eYr3DglkF0z6
STLQyP2GqZtUUYk+zQQR9DKCH1p4u6RdQBvGUr50qsf2H3xI4O3fiwyzQtQE
YPGhpOXwDRNeASmHl1IkEZiLH3fH6n9yGalq9O9lS8/FJwoXYA9MBaz+b3aC
Cp5zd0aCMmByrBw9tHEvbrvKaW4AqLzVMJUIpyE8GLRgqVSdKg+AFDW6mtu+
/aplNhdx1axuzHjdknbye7M2K2itmiAIeEK6lUtEujxSB6zGkHaALPESF+tt
b8azViVjpp+GuN5ak0h7oP9C0T3o9DLxyuu8EACsmhMJNdEvHzzUqw30ihZ3
Zp5bm+EyOs+hiwmVyDevrJbrM6GwhoSFhKypjUXMgBaP2NpG7t1uqJ1pQ5zY
EKVRZxuXFVLj8Z95hnQzFwJPrsYjX8W9qN3JGaUm7Be+gDoSbEi1w1nZHYhj
jtpMW3GxGrPstp5wtHfk/9AKogT9hwya4KsJ/N7cjBlGd6LEgs4LtS0aK8pa
I0xcHtGO+YQ5vqmfTBAavd8pZiQXdJn4zjMdZRNCsuIpmzoWoEQFfPfQV4qF
mzcKtNhhMR436bRJcSD7B/uqodgXgQ4Zrzo+3lwmHf76m1NBvn/1CV0FlTed
8QdmIKm57jKmJklMUzQzUvB5Hb6SlMI4V0hTas42UtzDHmUm+eNED0JWCA05
IzzlQU3IA5G7AkCmUXHdrYYgxliXs3wF/WhqWiDZ8eqYqWKO0gQEOTPlH/m/
gzytyFBgyztfiuHN+65z3Xm7nyqPzwsxwtJyYgQVtNynnE3HFjt9HGGzbQvF
eYhUsugyNZwBXZpWW2HX5ju/ZIQSBwekOl12iynwtPtadqOHjHACmpFZOeYA
MeJcR4m2Das38DU+92tYbdVjaIndbHMsjTHf1YE+4E+iJbGi2VlBnvKbbxCJ
zxKSEh+prtjx3cTKLhEL6b6HyxLvhJGu8JT14lDX2s3TXz1zIgT7E0o5SFrb
czpXQzqWv2wOSvLyQsCW6T9qyVSxYd9TCGcIhGIY3ixknJoMwTE0fSFQX+R2
sdEzJkucBScCWppOkB+XyIgckCh7QGOxBFCeVx0A0YhE8DFgdatcZhbu9bk2
HhyPb3KWsGyApNiFkplewMPJXZlRE+uBbBntu8xUKxIPW241LQeW5EGujE0x
zqZ7sL+IYPqHoofKV7H8CGcEn6vro6u150QYFwbkeEjEYo8GgSKwtYygcPCK
nHr5OrU//3/UzdKiqmB3uQu7ayEJ6zPY0W6W6ewPTvp9hSqWCqAIE+ODODl4
wmOXN0raNrifehlLkXtyJ8SXt8M4F4qW8djbtGBguX05jyrNacq2OpXxoN2V
SVt0gt0FqqcBEReYmDDZU8xjK0av36hyB08yyrydcI/7+TIlR09mcVoZ1gB2
UO7TreZFczEHpO3KKgn3eJYO+ZJeSu3W18ENvSKN7z+/cUpB/jFIKKoY+EQp
3+h0Z/cZyuosIy7IrbfD+tFCGkBcCA5HYr48ZkVzZ4cqQ2l47pVM+9Fd6pHs
JxtDhgCvReEcl9bZCxQ6UaMOD3zJH9jImOjWnO3d6HxAfvKaUhwKnJP4Qcvr
pJBMGmi6Du1XyWerOAFGntao+kJigGMvCVqNrF8pSZqs0C50yRsSlCDI7FqD
41YdiS9ffrpk51XWMZ017eol/D+kttDNW74Jzjh2DfWyc5ujb9lvYopu37tX
BQ5+GpmSELIT9lL3xjAqK6E1GHJul4GpZw7fHnDTVPygbYlY6xV8JmZp3N6a
2FrVucNCEZxlflR/GUab5uMJxT7uESPb4BIU5Dx68AqzMpa1/na0HOWc4IeX
EiGNqGbTRgf7dbWc+UKxrEDV0ZorenaLZSUresbPY5S1/7qqyfcbr8m5vpgs
SMhmhP5ncfa3ODQXw7he9AOv00EAxUi9K/Y8T5CQxqIuoDMnY71dkjpCYZHE
FjRV90abcXKV+VyoFs9g3zQvEfCoz5vgqnEIG2oG06gVb44B2B9jKdUZVD5o
XYyt1crcvAiqGeTsde299a23UeylzKaqMBazawNFXMnDS7gZu+JFphaMAEAx
QEg8A8cntBL16hdlDeNQLM19V7rZTD1FKiESXC3tVc8dyGOoPqJusxyXKOe3
J0duC/rhRaW3my6W4o91sqDosaNyifI6EnFwo3oyKPSSl8RsQrA3lu1pwBiG
z3WBLIFklim+k6F2UMQUzz0u3AIXRKTrLYhfs/46NTi9Yvu3ApgcDksXIOFk
Q3TjVLwhk5sZvGk51q0y6Xw03S8bgmEcFrQzBJpuvyKqiXXuMtwUv2kUYFMJ
cofJ80RXdX9lrhjv3l5wyAs8iu9i7bgGO8rIS1WOm8ij1XPMuK28cBH4FFlH
Lm1mrJBCoY+YJrceVp6HHhZv1XCAoekeJe7ikBIfUooiMPDJyGeygdU+maVn
rdgZZ5wgDFgG5cwgyXKpqesEcXRYezsHfeAWXHGRSA3vGTlvC18jwhHnfdPm
gJjVSok+18d/9Uh9L5rtelEGR7GiyWC/2v9XTrG/glYRcFBibVdevMcoUtMn
ZzPofaxVAunhlHqz0a5TaDEpOshU0CXuJdiXuOe77shh76cJLsnFW1ivqALX
l4I29N2OIQp42VSiPS4LmC4AoyJPtksgfyRl4pfa/UyuihV7uf29xHeDSOsv
bEIa2ndmFi9z9TdIlLv9B+bnKLd1ZB3xnfD1EAGAzbYI8uLdtM6Oh9Aqo0Yb
cwQszYtSfsWL1iYVgh+tM61bO1C0+VpYvTtoDQBKwEQUJAF1Zhn08pzvd5bS
mTVJj22c/UPZh1NOnEWxWM0ebIDQrPp7nrJxWNvcZjT2nO5RqS+UMgn20ZTS
r/WzaHEBkizkdRSnc1UnGEIpf6OfBIkbWxuRWsR7l9HzlG1Q9XiDW0A5OKjd
wITMzCCo9AIQ4zXzIwwVH813fdNWS5tcfeOP6281mVAyMxmcWYg5PrBilQ5S
7WT+DOv5sgBKLkDUPYsaIge/SPJ3BUFkcfQBsAifGroVVoUyv2d9FMaHC+Ua
81iltoPXxzyYqqlCKkIAVrxQMUHtdOsL+rpDe+PNEcXJZaz5FaqCYMRFbEk8
Y25PP+9OrmA6izEXtxflHFKSwJzuv8NYX2rAuLUdZ7P4S3GH4NbRS39v/Sk5
MAzBn8qAzPYfAzeQKJI2N2KDIPtI8/vUVeCfH2Fwe3EJ1qryKxhj6xnxGXiz
djiMU0xyX8EUcM1ZJPBj37fOmG3qN0Gkosa037Cu4IHDRwlHTccpeUc4KrW/
HO2MfHyInUXrpulNTM7DGbuyLaPdFB6/PivnJCviOvUnuCJQW14kAkYSmxXq
9TA3mfKs8MoLumbTgoFy+VtgZojLpi3i+w8r31XisfeYI/yBr9ZkSIGCEWuc
rnXtS+hpaZ7d4L22lt8ICHIyptQ3mk9Lkg2sPvZI/k4+8s1Skf8qU5buoX+T
SzHno6bRZpOwOKMGgRP0NPv/hER9dlHi2z8x9iSaOGpamoJjgaTrSzlqmwC5
GM6ZVhVz+TNEBYWbjexSGc9tkU9rGXM8Nn/hnsKjUN5RNiO/QRiL2o8vq00N
7JvAYUycdczO+Mjdl0q4+xaJowFpS45qbcliQTAbmNRtKSObNyJyoVDGH/1M
GPdqGM3UitWMIhN24Qz/yUd10rPxU9T+9E9cQMMNdu/AasLyWCigOFnLVFH8
rozihGeF6FE0MdVHhgT7GBPNPiL9IiJjObXqiLhSG0nbH8XVg7r4H/cFymqT
kSVv3Cpg0bqTmoMgkIrmtS2VN/swrDzy7kHKwV1qkYAOjM1v7Vujz6nNwuq1
wsr64uzu6bg/8kzBRUTyU9xpMpkUDi6HUKIMCI23qKzyMELk+o2VQgxCnKQo
q8eysj4KhS5xeW4+k6OqortJEpK9XgCmlm2wTO6hFdvo0tg2fBwjIePuMYeU
Y5jlqIBjKB1Vkj82L2bvo0mW1eCip8YcwOoUgvKxZJRiL9w5p8gcXSkKF9d7
Qh2bH5GxG1TubK02VqLOlJWHNKPXdVrI3ifzWNaHwEcXxu4KT+uYl3mt5Q8m
LtHVKduAj8JhVWqUj5chaQLUOpN1pRtOtExSULfDmKv8FXgCYWHQu48TCoLB
jXb+rZX784xG3rgnyTr8rn7R+13id3CPXdVGnT5Gpbv6QuwVTzOfEbPKbT3J
d2rPTDPnEw79GNALLynKrrklS0AgP9JZa7Y3+v/BP4X73AoDjgr05qn+CjKd
7liOPnGZdsf2PPBwQEaoZBCm59DAqi9B5l57RDmZS2lPVsbIJiRjng4TyYFB
nqwCUtSP3tVf0CWm0PkI8y1Sgr13Uv7z46WIzLsjZnm+GIz/KsIRaONnQvIk
EPIsod3StGQN1yU/JDCp0SAZFYzOIR96VOVN9Xvx1bHXDTLMXLB86VdrqvYz
GKrZjGbhMUEZmwreqdfDMhJ7viHuQoepG8AP7bHPZXzHjlPrvsa8YIcKwNRo
SwbzmdMZtm6FPxqsNW7zRoXntPD3dPE5Rn7cNNw8vZldpxZCp3b9Y4tR8zI6
mik9ACMug+lm9PTorS0T7/7sIgax+TYQS/A6LJlAP+urEr4b/lwwfw6dwq7S
Pf0BOLPpde00tCJW/i98wNe+MsvydKLji3DF9iHKVhfPYEu8xerQ2FInqCy2
WhOi1UVF97Xr0ocNN6YhHkDo04Cz3mh+OvhiidnRrGSK//ajVhShaKz1vp5N
FKqCcC3MXr7xip11ZcKCWHCtFis8Kznv7sXJvQ/1t9pQB6z1svrHUk6giRTX
0hdzmspKvmxBw+JQHIRzpUxTUPEeCx8wq9q2sjvuIvjhwp/B3Yb0Jz/8sY54
OCAsUiZht8DvKukr7xc+0dLr8giD7bJZ3nAXfn6CtvV8tvH27hmwlpqRWu2h
Fc4RGUsdkx0KwA6emwG2AD7fVgdKBbwWF1xDbmdpICA/rQerWPVMNG8WXYRs
1dO6Rm/oKD+0pykTJZSEgFiaEGX82b0e9BJV6WEuM+ikb+O60H9FyRMpR37/
14WIfUJL589VtcoDxb/71fYfYeyLmVvBEacObQeJan+/AMyKM0WAZnMZMwrM
OCCWbctXUzeE/T63XgHJXugA/+Ps4Qq9rCnAUraObLy747LhXoIONAVZgus4
+enG6DztuLMJz90YPEjNAwUyIej86bGdOMZbohfrCyUJzK8s+kGZIPbj7ENF
PmU3RGLDTYKGSgbijmUSyuxHcIYaABIcJha+8c+t3xfEfAOXIDQMtVJbUetw
OZcB94hwiVmniuMKXd8Vmq7qc5Fplm9ZPlHm/NkMHcTTjj6IUqP56ALFPQJQ
aOKJMZlZ7wiTyy0V9zEPnorJeDUyb4zTKk7wOQPeF7tGz19NKqAP3dfOw6Y/
ZOauet0aJoR5bNlKqhs996ql81HjWpt2f9uDg71T/OSPnmDfeCaLMsSdJDtM
O//dFpm3ccMTdicbDqKXsbcXSqYuhlgEa1JYbiabGLk8yeFj/SHKHPxxgiPE
ebXD71M7jkq6S3g91PP+KIFx9Hyvx8jnie3tk+VIeX1bcOtAFbOP4eYyqj/v
VwyuqibLpw9CeRW/qtOtYUK6877Q6eC+p4cqihtbSKkIWF3GDZrvZd3srsoT
9lDOVzKtxbltHHItWaKaoQ4rceYcgiSciP3tfMnDR93GMn5OVDRm8nnf121e
QpbzKERd6lu+Xwppt50Lo9gJezJsrgAkrc0v4iYvcmsiRMruul/LY/P0fg0x
cc8DIERG4iGnT952i4X57KkuTXXmW0raSXdFj+0cWR+9q7NUp9OmVK1dubon
He4j7iJG/meMcA6qggvI+EJRVR0MB3/O6Wch+3WtpH/cOenhxzs4olEGWAhF
Oy/h5vyCKGnhaDzJ8OsCgXHfQXk0eSZ0QW+7xMHjcvwntndPWH3yd7lDsvGu
aQ7EUEFujHdmiIdV5p43UNgn/0S9bFMX3VznuLZeZFMTamsqJzT0rjNjtTYC
/q/iW4rHykTB35sZ9g6rTYi6xg32Pg0mhRLldk8u/w5yZdVEiR5LjFq+V7aV
WNDNr4umzHBACzA1WYLRulsTYX9vzQUMSUQ9xC93yEruHod1xhMFAunSKkHn
q8P+lhMh5MHiL2eZ87VTtSZRqIz1I6axf8UKnck33DwfUOy4uh90S3fwFONe
wDMy2CnZO+pGpJFelYRceHhA7VoX9wmemA8vHsSiPSLCZirBW5jGnSF9MIoB
YUL6TnApC/Ahlip3QHaelb5+8mKj9tpsESjo9CNQ2UgGvCpjXWcpC1BCMwcZ
GiQCXRl3CskCEUA0j7XYJSgxbWwVCTbbUyWKTheyjIKHrxmQJof5+jlZKvC6
Tk4VuIgesQSzMW/R6j2Cr8xWNWi8YydY46e2BD8/BdoPXLkpzhqGZmtZVi6i
vDT7jknIZd4gPVsDS+hN93QZXF7woMupgdxn7UorN5e2kgM+mENDrnZwlWox
PXavHTspKTzZIxupWEuxA5zhVTs8mxdR6TRpeLEH1uSiEtCsWv40EU3sxcUI
JlOgTqci0TmZNiREFEwSGpB2C3X0wMGG4ZddnKAcc3lBj7KmWhCXlN2B7+Ro
f9UPIcIAzG8JICTLbT7vbcC4hUYAeCbbO8jWWsffvViE8VB3LtPPNjP9qlyw
9yXa1x1dgAqb9ZjyWQryzICdEhg9Kpvxqrh9pRX7MYnAZYbyTU5xFBrtUqSH
K7xX9QvYahoRwEHpxAxZt7GLV8knaipXr91Y8vPaQKO5FRIFHmNiuT5QWQC/
QmOy4iXz1bO5c7mRvmFuosGZE8qF0aT6gy0o2DT4/yGicndDjH4Q80rb74Vq
t7TuUwCVd20YDFjD4/meKewQqVsHWDA+U5CKGYlPxxrW7M1sLIyuatKoDYyf
cOBU555/ua0UuJOWX8W5UfF2cFavz9H4sN6thCSyKpq+oBLjlhlSH3M8W5Zs
TU66A59omKlQKncR6OCvzHXTaTaCNd5Ou+GxUoL3XRlWjUufowfOwyqRArps
rHUyosY+18uKnSkDJhO0Pcw3XBJB5+tws8RHeGnyRbIBGHPwuUuiwj2n0QzI
uK8Z6W3oCzUJx+ats8qllTCcKC+bIwvqxeOF8m/rAJNYTvO9LXYFDce6ifKb
SjH4v0OdJNUf9o2WhGnHKfoRyG0zy3UF16krYNdBHhGthi6+stahEK5A4uE/
ZEssE+5hgtjztjspQqLIiZR8lVU19/5MHPGXU3619G+fdYDxEhY8Xo8qcnFs
IjyTyFJQGuSqVYNd7jiZ1JWgomC6GmKl/SIe6zCDF1xEWwiigFT4OmyIfWjM
VNlX29Wf2WrgI/QTO0lq/KzAxU+XPKSqwDhkXbVRojRNc/ZF9LWygpJTFcHx
1ENA0r6zcMCx8eY1NKYOTRk91/TEGDH/rWnqaEXz9kDtZ7C+97vMDTvnY3kk
EApjMDIydkcApg9324UMk6uyAuq5OV/pWLtL2/dkaBGKdksGpW8xQHeahJGO
2ksW+4GCBVC9vaVVNf8oc+gYm6tDLaTij8lwJlvwe2ih8tQdHEkYEzaiJTz+
URo3nMZlxzqOKxGiWYE7DJBjLCYOX8TzthvI8hZ42oJT2Q+GKENt5l5aQsIi
cjbEUHVBe9Q1Y57f/u8Lm0RZN/rp20lY2VQwNIn3AsXFFpWTd1DJqqQLAMvC
uGGGiVEXW+JTw86FFF9iKBN4ieq+ppp/M+wNz7/c7YqyBh3DQA+uWQFRXYe8
+zDqwB8yzdMwZMk3lUKiUP4zKfbk5VnIXQzYwR/FrgKd8P3vGAs9ah+Sp5ls
kfndH2UxiONGOWrCxVq7pp2SV0Mg6K52Xp8QkTqdMOQdn8O+f2e/sqSAQuxi
soZezWGBD+I2tvakkSedgv7aEuP0Gm677UsVA1Pd+fCDzpB6vT2Nr+VU8g18
25MnYVdAdDqcEhm635Lmy80numdH2+Xxd04J1jhWGZt8W9gHfBkHxck73xI+
c1Lw4GBH+hI9EOqG2iyck2HiRt7clPxz2K/bkaSte4H265W6roh2xvj56brx
xIFJ3nVveAUa66WJmMek4z96xCsXq11RjKIR8b1h3dFal2ce9kACUQHppDI0
pYRY6ay1KCUlpCRq5Wz6TzUKFYQgmwvnVUdF86j8d0tXnPnvejoI/1HzDtME
mL+UGRFpCXdFbum1bCB8tOLznUqgZwMZcVIJ05XK8bu7fXnPLWadlBDeRU1u
oXl1VSt3goSax1cM0Qq8n113LCKnLEsY8zVo8nbqHEC7z1AJ0vKdTBFJ+Q1a
UqXw8tB1I6OIUaEY7agYxIbJ/EjRI7nOR02xjUAdEHxb+rQ0tF86H2LtVyIz
m32d0z7xjW0A8Sh3KZTV+XBIYR9brJsEYizjxEPaoOUw4uvuaeSo5Fkhbxnf
LCcaHDFjgtX3SoxZ7Y7IhYtFRTwIHrwQDfYhX2O4kbxer33LM5WJKy1AYn2M
qhJ6rz4rHjo2+tR69Ll/IqfvtPHv1h/d+ZUtrWaM2aBOIFk+lID3jayx3oZB
XSeF9pVr8DmggSB/h3jLkr/aLzxHA+MInGqZ0W7kM+oUDwdUpOa+RaYR2aRR
55WkGRbcDf/DkRDf6dqA1SK5x1pNu5vzgiyZnMazIJ/tKehrEDOSTNLaw93J
4qoZ/XBs7RKbjEkDXrsP9pM7pX+wRzW/uvxD0AZ1B3p5M/qRpP7/dpwu/Nty
8em2BWPvezXP93wmEqgO0IKeeVYELg9NxOYR9S3IaEm3URLYdbRSsGP9NqjS
iIvhwh1h4BkxCCXO0YgXfItn743mn04KhfM0dk05vbGoF93QbvmiP2/vRg9W
A3DNbAtHdsIwX72CyOUvn8YaVuMNsxVIsdU8DIDCN+fzjpnMH3ZbZFBvDw4g
HyDA1Il4RPhBNnGWxkBoJAGdeh0lSUQOq6Lv+SRz3uMOACkMrf4qoybFOw5q
fMU6bjnTxJsQuShJRoj3OeIXyEVJV+emn5yf/xhnJi/aGqUSHL2Vdhk/JSiQ
umn4t62V9x6nGT+B5k8/TA19NnOgaWxxawMxf4QhqqoL0MquHgHHwaoROU73
Yb1hiLwlxLtHKX+fVE50c3bX3PTTFx4z/pyq5gs/Vr4aQj0hC1t2f5f4UADm
pgzfBoKaPMC8B1D7a/2pj3zPNBt7RvMePuFgpAvwNBuQjVyE0KfY2RubcYNa
ZRHIAN0xc0zFKi31OJV1S3Hi/RVwTzjq+8uJ1PTOC3jV0/mxw0l63FDKLCnT
jhqc7UJSYPwJPf5qJ49oL3w2U3uow9Ji9eQpZvfTCDc6BVwZsLs3H1d+7sQ6
IsmuOnxwfA4BFQkAHlfUjvCwjw0fcC0u1wrAlrk9XgfKM1Y6hRCk4wJV8rNA
H7jCmTuiwMDJ3AkTgpozHIVZ4moe8J7VSDjRndjKO3Ue/OnPAJJH69vAJgH9
pdHCxwGu7hLIrEpCpxLe3LBpq4C+927UNLvfeCYHwwFefjUahJs64wrMl2N8
B4No7SFxvR92OmugGfsgEhN6Rj/BhdPtH182ZSCY7rF6t7AhF3TKfGHoinrw
yZCHrBqSVl/x/s+3w3RYwOeXPlMbmSQbayBwnbtvfykzWkSFWLTjKqLRS/tp
b8ov2LdONdg5ltfq2LZzsZZtF6MJHyhyRemy7iHJnPfuarhuHPeGw3NurR3q
DjW+uSxwSA5ELGJU0ekn2EH4jBfQlV0dkBUIVlckRvOGY9jPsAz0gH4xtd1C
v5iVNYWKrO/NzM2WZ+687AWJ5aeZkMO44wc7yfF4noGD+NgvyHGeNX2dbyrg
zqb4DB7hx5CU+NzyIWTKglki+Vk9bJQ43qOWcpj3EekOqTrKhRZ0zxo5TLiz
KdjM/K87Cy7QRvOzRpQlhxt/YmbiOqvofubYcFLlgFcCVFuT0PHdCu8bXY1o
GYwnC0xx1QJgjAi2RcjlmTUDCjT9xTE9FNb8jZMhKECPDi9zL+IujwyX6YGe
0Xlu06IPxHscWY4Z2jesKwa+ePtILeGamU8A35FizvWn0bHiJcVybbqEbiPA
XutAfmn8B3nDkn0JYTRaNCHD3bGBgZCsRKrgWPiIOKE+zhd3eH9g97FmtvQ2
29hIEO2MoPDAcQ8kYTvM3LTwcRb4trkFqofbYbjgzp11KKUD1tpW3WSY58x6
3/N+ynsbga54Uuacw4cPP9SJ6U3jOjYVWRaJXnuPyFeMAPCPldSjxIhBvGpD
er70ezo9u249/Uyx4B0KnqgoxZGkabamy9CMgrB2S6xqigOTpUDhwTPH+sRJ
K6+eqOTJ1s+LyhQr1pI2djr9FeDMxth/vNN3oSV2Z+4d7utLt2U12dCU1aQz
cSTK31TUzApmM+B9XJyBAhDjsBW+r8pRi8JuQENv7Ixo4J7pZZ4aeBJW9src
FYwIsG+sGSTAbU61ynDdVO6fWUa6JF2O3MzGiXQ9dun7wPC/K5kC2AF3l15/
bCs99ZtNT7oh8WqcxKfean1/7hNA4Pxc+fbw8v0KK3B1Y/0oU0LrErmBh5AA
oxhYSjcp2mIvtmNN1XEI61upkfiF/sa3ZpheNwUJgiShhAIFhOt8hmF1xU5y
vvZhztyC7q81YStNVXDWku5JBEUdP7jb47xDhOwvcYN5cPGplpNSJvUc6JQ0
shVzzhltobfkZeGB2kkYOx2bpWa9BwYWRcpQDdzTSGe8xOLsOOrTAIZ5KtMP
025iXW70euIDDVNINERtzFRG0MjKLzFyyyYWmcTDsKoYwvSM89DTOuPT5aSE
3Z/oC44yh4JvpB7pH61LO+JnrMCawtCAho1o6PefKAN3lj402ipVTTiEJiSx
wjGnzDvMfCmCSUuCmjT/kDk9Qu7qelrO5jM9/Hw9RCaABdqzYqXkHB5fhahv
fmqJTM87wYSWoQtDsRr7yb696zY3ydfC8/E4LUHBssoljL4jfBXcJPM5g3/E
8xcfq7zi6/C2i+is/6YgExYCeL5VdMuZluMTdVojX8wKANo0ipdwaIjqSmw3
jPmXxogfjS0bSa4X8ibLSB0hdIAUb+gJOPJKbkepdviup8UHLRrtfGdHnKnv
VepuLosRGg4tGzVhKLmOnSSRY5xCsBM/NEsRF7CrvYknhiG0H+XNELFodPs5
hxFdS/MoYHj/vdp2L+MU3UmEmAvCendp9gxWvhZkMDQR7o0i2G3qhk6o91+R
aErzHef70ARBUYaXH3l/QnKqg41R0dbqA1bS+9Fs1HbtVafM7psK97mpNIv3
lOSTP/vLAF3VEkFkCSCXcLnXfMJonx5qP1rhheB187YYkVcpVeV9WfOvHkPr
jNhhhc18d6CGWto7JXfFq1aSmrfbSuSxlQFVwOQ68SRB/GQnx0ivazybnKeR
YJEy+/WmRHUUuzY8r9k7O9wALUHmtPwvQwj1O2pJjEy3GEVCPRic3esy8cDM
ecin4E04pqHKoT+h8s78qz8ycdgCBuXT7BvwoeMDm4eIGIu3hTdpHbiZz6HR
dhmTWvsKq6fuEAfixjv246LO+7mS63GxewI2aD2HYx3WRrtxClPCOWYJxTld
TKfCr1KDzPnRTLv+yQIMYgWHcY4MY/J0DeSDFHgy8UgV1y2XBf8hqYZb1psw
Uxe1lC64BD294noXPT9pE0hATd1o449JrmyOsxnu4TCvbJjCuMEftly7Vvvj
dvcweFcheJyAit75QlsL3eZrYSOmD3UStwqqaJQ/e+hg7EaF1XbAaz1NYueK
uFAU3t2ucU7avZ+EsY4R0BMi72LRiKkuLUO25lgSx5iFfiIgzx8lwFOI9GcA
Y2iMAhgqg4pShquy/ux1HtFGVFzanSyvuJkXQ6dbtVxee5OEgKi7XahjsimP
1bTucyY9B/6PijMcyXsO8dT3iWwpJgpnshuIFFsF4cKfiy9x+ZD/Z/10u4DQ
S/bcqPS/bN+41wrtTK9zmEzrHoDVLv3Xp2J5ahpMRJnh91F+bvgwDWqjNxSq
r3vJ/f2TSKLLd/vYJCSQc9dXJ7SZ7hpJilLJEtnelY1QWyjL2zLNuIks3RjG
4XMOXaDCP9zpNplC8cHQOwN8d5Wh127WV2C+mFjgmtHvCE6YMaYW782xr4Ne
GUdJAyYPG2cGs6ZDRaCiBijD8bKJ/fcXpUA2YdrsKQnTkX0X6KwT1WJbbM6z
VVWnDLaqUNBE1kyTbpW+471SFMNW0FDAIFgWzq8t1FGGkzua+pFPGuSjmQA5
95VSEf8qJh+hBtfHwxBAc5j1hKCrf5P/YbSvkKrj8v91j3o3RDRc6JXkkmaz
Lrvmx/cM+eixtveV9xzBkVwYKFieQv+HkB2s2ImprIMdG1E4bkwwQqs3w6jn
lTpy3epEjilFy6qkb19tK6v/N9pVy5+g8lHHezpokTBu8T53U2RIhAGHGR3l
eMCmJc1Pqu5tlwtA06aDPuuDecM4JySURVm5l/M8dL8+0wj4DJRY2YJ35BkX
IJxB8nzwgBtjtDE0bU/Jd4dlBA0ZOFzK+IC+ZDPUZTDWsBzYiXpnpoROlQ9K
GA881kZV46Ef28KZNFKrjwscauHhIxQeit8xo++SQ7+K4byvCVIu+58x562t
TU8Ku8CGlN7dtGqcet0wUZS1iqns4iOnaeWjusAuDRn8wKYtLRUWinY9aX9W
a72BnmV6FPDXxr9VMGag2cmW1SnPq/bWwM+jJZh2lbAffUrDGBFHkT452Zyx
X4qfqiQ4MOW7cBHJlAfboJ4xaYo5opbLx37Xg8FmnEwmJ3CZgLslAOtyCrdC
9oAlDLHpHmXQvbLSWEKJrlaUep4PHDUyhCKL5SINK4Rmp8KAYjhgsQlENXbB
UzHfLRIZxQc8KHhWCKczyEu2XsgMRqbVLw7P9eXlJOL+R7hck/MzfWF52mGU
q8FmmW1HeFXSA8aTZ+SE6oStlZKlTHxEl0+EUasdAzREuojdmGxN7tfwtN3i
lAX0JIRZL0+uMIjbwzGLmDow0sKWPE8tu/h1CnwxxEfBJ4rrl+2YiLFI+CB3
RtXWsgBSotvseEDOMT43S4WI8LIHvGdccLu2HOaKrj/jDID5Gmo6tyCz7k0K
7zRQY68+WDEqQg8vZiwBr5ylTNW2xESqiiETSQN3efYzOz5xFADFfdohAGJc
Bfc26mFc9toimmmQUP3RRAP2+i2262HJUXGXDtxBI3yPcTCS4t/YriBQY2p8
oHBhyWxEqoIzCOGv0W2KMhETR1MgZ95ZgdOS137rDo4ybgc8PSUbJ5BqdLcB
XTVBP5tfKkZQsmrYNMHOozNdoaBjd0rWBf/BY9WPFKzjwiJJQRMato1hmygC
VfvffjIk9ypykLkpnKPKvwEKyo+SIeNTGzySZgTHIWmRjedx0gw4mhECTLrF
93rtyAK6+qIBgV9XAFS7D58EpWI3pBUNTSaQ5m7d9qR8g7ONEoYSLBuM9bw0
wcmtYgxLcpDO2MVxSVud1pR+nEVofEkOPkG+hDCJvYpl/xEXZ9G6qcMK/yOz
7KltwKi2y0mn37dBRusCIgF27fXwSpCw8ERUPV2wzsmZ2yOfd5Ch+eFFo8sE
kyKdAU7DmMhOM7NniHFFyAtYC2lAghRuQnqM17doDX0nhXGyW4Lb0jVLnpBQ
OKGWUX+rNRd0A+pDjzzUNR4Nj1nlrrogI/gwg9gWS6vJrTHNWPvTL34XUYy9
a2io4wQYZjVT/FwoCL2PZAFWU/Ic0x0h1kMUa7SvPtaDFT6TrlUEZSPiM1kX
2hcEmxx1LNuLejil7oN3tnTPqjrZEPlVL/NduzAdYiTVDAGV9B07JrTajWJf
nlRcdEx5weJawR8pWQlz4ZeYYdxkT2yGVtkPRDQax5kIZe85mgpSD+OAyH2H
n7+LdJ8YovIARF6ak6JlVY3CcGQzbMBNDWJ+JcuU4yAnv64x8dUZ6Jz/37Sl
c0VTCxsCpFPHySSfD16fGXnbeSlNLmPkQm8K+FNNdSZYjCLSSrO0ii7ZlRCp
vtQ9iNa+rG3+OHNM1l3ATo/b1I0ka3wjQ0A8hMy3HXbr6Mwdk+VHoAEkw+AW
IzaQiZq9qADkAvMgV4SRTDNi6UkiQTId/HVSDxfpQH3s/v7QroiavDLmZhsy
CYihYhTiGf65wriAGjxGs7ADG7kI2/clQg2LuSFCfVtVknMtpL8/l9qd7oF2
X404QHPGBKMaFqCZVXM2HYyK6/N9eeAVETZCneEO14+ngA0rp7YQwgyTDi5N
j2pZ92FCi+awV7mSGuxe3GUPebD6zXXYLsTv8NYgKrJI+gdy94S2LqOTonit
nI+9gdgZXRJgEfCwhLLRmcJrPHBP5bo4aU+z/q8TbTjb1U2Hb+8VzaRejvDY
FdGN8BK5YxhsTMJMb54E99PXO4yp0y1nayHgMPcDZu8X5hlYpOHS6zeigxYY
8hI4FcZ0fLzznCII8Sng6OIhdBSbMncmXoRmidSStx/6Kx3iTAhPQ+PUj1yA
DeIXfSjsio3LXzrf2pCg4a/lfarMFxcYy3P/lvPYZa+Lcf14YswuG7BJhNPR
HG/b9tx528A+saJ9jkJ0c3XzhFVd4Eq6/Y78JQj2+vhncFU99YHjT4EQpfex
smyWeI3TeZsnxGdwVQMOAKQUO1BQRU/AP7jlSihAIHqlT1epGkLbwHFHfYNN
CBJJ/KU3VjjuXMxGNrIo7EZ7akX7SJhpII/tYZurDFMqrjBSeNpoMsNUQjsS
RsRI9v+qpXMb2VtL3L8JFTY5r6XbZwK0V8/vM4B4OL+RQq+UHs8krRRDUg+J
D/E3UzW+v51j7HZSrRI/do8qFz1RuYNV+cvcC9d1pYyXRophrgG52hpztapx
ofXaBFQUiN8u8+7soNENr24L+4g5TcWEm1gCpn3CRIhpx6YxHlkjHE6zoBMt
5MomovMf3tlfmi5Pnu09zZv0fooR5ansomevKQNo0be4Xxx0J3p0X3BBXFn+
iOiF//UKWPjuehghISCCo19x4ECnfq+kZrcitiatzpqM7jj35CRfL4GcGW4X
Q50VASt5rY3b4aARfUelkQ1qyUh+zfiTc0m5sp4B+lMvkZpp1HZsWbPldSnE
rUwvylZ3vmnTYTgrYisZZ1KbgpSzrgZqu8ifxkA7R2YmGPU30lyho0ItNfxX
8W67CarVKFSDeg9CvFwZHHiDTmo/3elnVdQueivtMapUgsygAO9hl1u8Fp3k
E+/dgRpQXZM5DNTA9XiKVj+5pC4c9ljGncle/+GqwoFOuZJ2w1f3W1Y5BYNL
NlW+Lmx5A3F/Tam3oKYqV6LuTgDrXbh+3d6+1koiRZGYkeCN30stF9+0csSy
TKW8d+GdfiJCvjskAOdpExL2hFmx9WTXU/e8obNX0cvJto71rpJtovGSkx0P
UgPHl1FMj/s6G3XsVgBux/y+GMosTWnr8F9rBrwtaaleGsS2mmsXAJfXUDdH
PgMIIyqoqA6rMVuk/E6JlnrmBBUkzQdVp5GhH2VmWcMCwlwBvsvk4UzpUiim
yZUNxNouq9/k8NF7jG7tf3OEdHzs4s8L93POAzXBKEx4lu4ZQVS8DheGrbH+
xpW6NfrDa3nzhUc1v/+7JueVQjw373tWD2YjKYGkraYjidZjcZ8NnV3R26Am
040XQbtJauCyQdPAY+dNQcY3ZEc4gTBNtKewAH59v0DyUEGTqHZMMyAxrAA2
9NPA1Bru2KB66ooJEeczI7xD/cEZjeYE4LAPc4QdNQ3bTmi6gpBnO4LvB8jV
ApYvy6tJv5rD3PGyDBlpo8/W9b2A44Vnc/R/duAGA8Jp2FD4ENX9kdJWR4W2
efMjJOrEmI5O0FdFIz+pPmWn3BR15r+P8KqFKXkp6XInnKBbYSEhSB/LwI/U
BFZZRLYsgqWNGADDHBrWCKyKctR7nz7Kg5FiVJ7L4HaRUy4dV8HZQ9EwRw9j
7AAsGtzJxLGAQ7b2QZg48ot2VNAtypbpwdcFK/drX8nFjwcgm47RPLNzrga1
fOjaav29+RZucNo0di+HL/4ac/IxhUkkZp5evx4rqI6um8URW/TuDHf/l9Y0
6WQznCryi8HdP8VcxllJZ4X391Frq0CeDAIh+HF9r9aC8mYPE9sG7iDeXbsG
RUIl0E3fOaZlWB9Kk0b6pH1Mlqa8dQB93NCaDyhImm2dw/NKdlXsBYbHM5YC
u4hBvR4A0TLXUlSxix49cO09/79cdEbPN3It2cywZWgOktmqNFfDLNtrCEQp
o2VFmlnttyAwS2BaKhikUbOGiNClT7xqiZ3eAXVJoPtc4zD/smEqJgNtqcJs
Bg4LN17mYBP92RPuFpVDQswJ5fNKQrCSaAMut0ZKii/kygBJdTfFJE5eK9FZ
nApPi89F0VogvDp6q2r864zRpM5nay2hS6sfAc6+oKmPAtaJ5D8oaj+q5Apg
fV1CwKObAvmyRRvZYSAMzB3brhug9TtXd260jeC7LPhOa9JliHSpK99ZJRIP
WuyGV7IBpjMIgrG9BjZaJLkK1Md9W/7Huu33ShWZB17sJzq5ZBqmvXuQCVHE
tC3ULHban3Y6mZ37YeoFTHkb56/l8bNyb/LCtnrB+l4LyVAi+Z3DddXO8OzR
JUax9PznLA6Ys4IQ3LfgvsrCGQ84x3QE+6mPvWrAu+oWyKlvLVSWtp1P4i0I
75XKyocFVPJ2md6nOw+LpODy0lei0x0+5FnXDBcqkPFn8xPIJFXBgMOzMlxA
FQ0+Y3ZBqYDnxdzEBDYPK5sD6eyCITeG5Ds2Xtp/+WMkrlXEVpDnTZ8ScplF
whX0FJGsjbPvLE69EkLx6AywNC8x+cxPZFx/Ubg3IKJJV1uCN6jRoD/iUFY1
vZs5TTS/RPNlHh6XcBrQNYZt8w98fOYjNxN2T0uX1TK5xq1a8Os26YZKpqM0
BOcLSPRQOMfPUPmPA813/4x015DkemN9omxzA2RhAvYNIOcskzysWowZ52tG
gZ7xICNVLM0wHxBuEwtulmmB97jZI4Zz9nqKg1ZLq4mbnuxbnDp6ZA0cAkgS
GY3Vt1xuTpTOfSSnBZc20HKUg5YFfqF+u9VQAqNLTiGJaJqhzIqfXIwIBmEH
8dMkEJMwPwpJtHqECg07OCyQC0g4+Ia2qcp8//vY8vJusehG3P+HKcPBm6mj
HAeIPQ0MuhV3N1MaBIJjOs0dtkhsMsD0jWnzbyFiMO2wjTP92ZJG5mbOhgXb
pSlrV95mu0+UlwXhvtoh3gZHeY9tgcxzGyr9SkV1Nt0v0jQtNMlJpvg3lSHe
X+unEUTHpqdNc4eXSZSu/hnY/sERtRD1Q8DFwC3Drr+Vcpk3Kad51v0m8fYW
OYB9HpPgXU1oT+FZS/6XnRAQPMGUfCslSk+qamUD28t2R5AfYGkJQBuIA4Oa
gDW71gq8f8zWzZF1dGUMmrn7fsLn+OoWVCS/mSqCJGvLFsJllXHH9lnOhlk6
JEoXxsip4U/hSLb9WVEmgGxiutDCnMMjvu6OPv6Kw4gxO/aJAQC2qpD717on
rFUsSVP9MJzSSi0mfJMeAvR8gTEYleJDFWrOyHkKfUDEmFfKZhpoDkt4iJ+h
IKBCwsX9Zm7DCBlHtWEDvoir2RMiRNgsetXIxz43Us5othBYFufjooThA/ZW
N8ohy6K0qZwF+AI4eyDOm7ZsqXNWkPsbYGFY4Gsk6rs4t1WllFwCxmZEBTXA
IavOfupA7YrHFiTtgUtWO/8eOUsalm7NAuauhilsnyd3dElgd3wSDCjzJTsb
bfg2IWiqNwLJOysjqK6QQ27g/MZsfLP2WieDgxM+yKtuwWiysQVxVIaSs2rc
1L8i48h3XtvmAn6oBLQbZ0tqXd06cYgcq/YAyzOkARwEqnAkSme0156XlF5l
cweXQ3VDgWLvnyyG8wUQ1kqX5EgFXSxiOFx8w3sR9J+604bKP7DVfvUmsja7
uwIZgpsOksdPjZRnLx3HHELwtn1syQFbrZwdD3bjQsS5NVfpKhOMeT797Lb2
DmGfNCHYkJEiUgjn3Gxxq9IMmlN+2UGAP88S1x59TmXXVFLAhHeH/rge/s2B
eeNss+MvB7lc9NXRw3g3wgb9i8sZKtQw98/N997LSSh6rb4FvGpf9OouOMil
7FLA+DAxPjAR5YRHbF80cDgdvFQNhpXroxlx6/QEPHY625FlMi6necrczi/B
JBfVf+xTFKxXZTuDaSYnh1WbDIN58rPKj77Xg6IMBKCSxhDLBiOr1ARApzTi
P3wCoLAsSgHnbQcCmO6JFHMATbGnx2g9E07zowSEV9l7mb7YldORg5zfFa/I
btYXtqGlXdvwqFbLrhqd1f5t0+k/9z4JnJboGV9H2to9wUSmoa3Ueh4DfULC
6sTh/ZZ6p3Hvbk0AQ+r2ecQWMvobD8ezK5f5YAf9FIKXrHWZBIG8DbvqQJfA
VwdLl2DZ/JHJ3Nyx3nehkzNiLJspPnPaEyAVFaa2+lBdoHrc4l+EusBis26J
SN7ykJ7EWjGYlD3sWwows/tKzWYGNEeP+B9Vik7ZlDFVPEsUfrOfM5EPu1jh
/lTEkOV3Vqj1aY3bHgyLHsjPNRaL/G1GmXTCDH54z/24dr+QZs2frn+uhL+N
+S6d7iOJ7tXN6kb88PhyJrZHXEi5yRenYdtaN76KMhgpYEvmzd+zxNVWqqqH
K5N1mkf9E9j1T5GojGZHpiV06QlZIyDQEL1tpT0m6NCoJFy9D8uGeO/xcgdv
ZjDWaKzOnw+NJzPaJkHFfbI0Ljd3y/qQ8MjU6ZyspJlKMEsKPBrIEtOq+hKO
ZVQLxqRUA1nWLf5Mp+NSgQVtK2tvQJN++whA5G2t2PMEw4DrGzfjbX6AFjAU
A5yP7rGLKRiiWdCdr1YcMCVe3CRWrGmHtNRhaQU0TxLJOcaWo7fwsY2tqDDa
hOKZc7uFcFxI0ow7E/h7vAxbODAOusbs06+XuwJpfmM1Na4++ZnDtOZcFv1b
NfKFhTIvRUALQQvWsjJIbLAjFMsOz45Cysub4n6UpgGX38Tq9Y6E0zuhulte
1vXXtwc/e8k8HuKhYP1NnwrkLUrvqGT9w7EIORhQbMnzHRrYKj20ZDHA/gq3
YeRsPjvv4BUkmNI//uCZ4B01iAMF14am3Up9t2WPSZEQJuEAK668Tz/L8e54
fphicDFxTEt3PLFCbdwTsMJ+e9ymej491U8JaFAT0B8vJHAVwAtw2aw3tk9j
x5FLGPMeIG8QWLuPUJC2swBwYnAVQCLrvq7LI1jbhi5Bp8mmtyOz0oKEF794
G6ID6zijSCLAx3Oc8zLyVcWIHFg5n07W2KKKIqLFnurU6JJR6Rv5oitE4xbo
Bl4pSwW3B+fYbmpette8L9/m8jWODiYEwMZmV5vDdCrLdIHkygGNwT0sqDoh
rXyrtWunGfKCUqT/popsq/7hgdjmuS778jEZePueUrSZ5r4scvD1OqHGXces
KJlLJuatNf+8OV7Al83LgFk4i5KHJzghgNnACY6tnxtaHS4lmoSM8W71b/zn
3VwLbQY1I/SMOTFcQj3n6h1WfjYDbgHZ9Yuw+zbxVtGlyNR6pI5QAx64CaRV
Sc/aMFBdS09sdRSOFcJMSFMCaKYwxqINEu03+2pnpi64f7k1IFkkDCxwWLPR
CRcDEQSQzeYaWkf6MstHmjElU4W5iVBa/KxnaFC0hrsxJ5SlamP8WH9TEpLh
qISGHEuBzpbdZmIDzPCKzntJZiAfjXLZV3SDaIxj6DCmt/yHZNijM8i4HFGc
QvKOChoZ7KhRUIccT+chiRdCVhamtpTV2q8h9E8BbpQuKGZ+XT7xVPYdIudI
hegSAS+8iDoFb882jImZIFYuKVcLRwoJNyg5YpFHcLOZRWOenPpm0M61hcXN
PXcdhBvMOIYo1d85169DAO1O9iRI5cPXq9GOIXGcaxu3HQBrmiLJ5sgFtwch
tIAzp2P73JF8K9z+LEkdNULEtuZFJRTGlt8kSkye/Js3U7bbqbxjcAIR3GQ6
Mol+c2DG/Y6Vw5CwVf79zYmxg6gRGtb0SjTDhjlfmGk++mjU4dXwKBc/HZR/
z3qP8ENCe5AsXgmSsAh3mpdWkolxX9DfcVkMUKu7H4RQuS3eQ8Zd2Iq2B4VW
Tsg+NvzsbiNqVAa+7KTIoWVTLY+ldxqbH+FMfFMl/wBAQlHPc2HWHukFftxQ
kmlzUYkbfW5FflbjVgxxYOux8eGjrNYJ5ktPcsmGKSNmZ003IDcKvdhYsYrU
XaqN6W43g+2EQWmBnZEy+CKB0aCBZaeOlt55ybtL2VV+nYhJFL0afveFT4G3
upB6FlBpeFH0bMsLpEvHawQFJmr6cZxykF+qLuYgTCFZHiUB+QFLYroQrK6J
CVCf9eZ9JimGmS6Uwe94WTBKpRL1KUsoBNLZi/qyjJdcm1aaJQpb6iT8Qg6d
G+fh44tDK1r+9OYNKIsMWboY8Xoc/kqKcJNDa2C6BWYoq+KbQBIWa/cfbfkW
QBHLxTHUAH4e6ExKNeLpbDbV64rNauOStdgYRJfXbyolcULOEjAXIZ4IPUuJ
uQqAdUFmF14wig5NYaQ+bUWIrDkiDjeNxL6J6P86GXQzKieZ7hqPrk4ykMcH
uynmo/j7/SPsiZp+HGB+InxUvQltVr5gEs5oF/AfNDv1WS807/o1vDy/NNVy
aG2+KoCI+T0lEYIIa1dgVaPmpFQ7pNUcVTXbclpZDG5C9QAPCWpCZtxCaMRU
kZL1AZUXHjfgSWzlCY/jSc2icgztArM67i0diziU7TNzMVlRWr1IQdxrGZr1
SsQMDTOIr/Xq/geWMBmoHQ5r63HhqK4eO15WidmAYOaYsHiTAPq86jZH7Q1n
eF33WCly8CfxpYqe9ywQbuMQfo4BCM643qVdBTPNf54eNTl0ynW7HQgvi5ER
eqjyCOgeyt2mKoP1Fv5YAjD/dklW4QFzXwTShqnPdzevq8j6Hs9VHYUxf/Zt
ry/rB9u80kf+aG1f8v5jasNc6gTGMiTqZ23BkfqMVMLo9+nUz7LtfJM3I1Wb
uqZ24UuTgo/Vf66f4RUS7IC862elcMY0bhyOj+RKdxulv3s36w38Cp/fVTfs
mQzcfI715umWXCQ+KTRveLRNbFBudEv8zlC2ZwGsdFS/76/DAjYABgXhGLI1
rEMGkNk3pCy6AUFlNlk7EabqClB2JcqVQivmh0OeK+qMCkCZUSnwgfoJWb38
ma1zvbFKv5kA9JpRoZLiVISSK4QJGp1c6bda54LqUQOKXQAXgHhCy+gqLeAQ
3y5I0whMWGbF9Y2wmC1EM+9V7b7ai26/VUOwkmJmSJIAy67p4yEIkO73vsXy
NwM0CmkO/bXGPTfmfOT+Ft/p011L+i4VPkjGJ+qq9kYOi4FIl7HiWERs8U0+
CUxNKvVGsB7ZTorMgT8w+IK14WONrGXaCuwhjVVTDu2RFAl7UGU4vgZhutOV
PsgqfarL6eMK+A4Vd/isWVU+N+CMuprPbsN2Vgqp+jFlLw1yGEJj/GPH2LHo
5ud81ksNPPlCquugW8A3iAJKv+aw4SrNZbpWw9haYzn0PLzfV2om2e4Po0r7
TOoTA4K0a5uMMBO+auBOe29Tqto8xUpYrGilrWX1QlVb50Jm1jb0z3uS2ApF
98wnfpXBdGX6aUm5Lsg0HXuSb4zJHj1dbkRgiin8xO8zLq7WdEHlLyvbLste
HY4pKIiLrX4SrigbK6qzc0U/L7MzYX28GoGAFXRg8cchL/iXpkZ6qlnKpg4z
KqdWtFVG6YstzlsZSLleP9y5v5j1uBtoJB4c7S1+PPjJ0rya2n2Om/vpnZpP
VyP+5gMtuR2gagGtePAqWJehXp4FdTAOq1J/BGaR8U2AUpBDQX7o5X017QZG
T5AGJFWpAUMxdPJEgwYd8gBX0lcBQx7xV56JWyQGkKAfthrCdl8vIsNNu1+6
vd5GFxzxogn+78Wjq8Cj2wrAKrQ3bBhW+9NhGwKaP2kJbWo5ZZWeloGp6zsW
DVUs3e7L2J+n1JShrdrg1y74RRRP8JTv+JqgQ7sQ4UvoFld4KYJ71kmeC/1p
8PBM8LihWVn9uE/eLRu66lUi6xLR7oj0wT9LSq1+dkBADIQmtgMqlq5xk29Y
kNgNfESROAmz+uaQ4fyav9920W7l9fBdUp3dlThivcgAGTzMdYT4Tz5N4s+O
aAbRIozV1JsV8bmjYljzkFJRehkufbgSXfNPrtmHUzXPK24ULokUmhKq6Sdo
E7/4dCViQoiS/H/iBOibceolSgMSMyLx5GkWT+EBGmub1Sp7V+ULCYF6A8QD
Nc8xhJcGBlZCuuwdngxVYBuz51gGneNYca0OZzLyWRmDtCVvDzpkhwUuqhyc
DYHzrF7jkuxiRfdfTmkiIywPwpOgXtpOsQzsrPIZiuwUX1srSoPHEFA9veEy
0sOo2O8Gq1LC8fKLtdpembRholnBSi+CpHUr0pB+LfLF1G8h9l4zJ0HKO/j0
Fw5ty9CN1Nvc/Ax28uZUYugN6nreNCrhL/x3GFzxVE97CNAO/HquDJYNxMRf
G11sNc0Kgh43zdPdaATR9oXka0OdB68NxluwBnUYVjCpRtqlxGi61PBUwrPj
bN3H+u2o7E6kmOQPedg9gl0bK0yPhtvKL0jxXBtL9NlPnPyG1oMxYC3ZZ98L
bHcE9tFxFJRh8KhC/4nY55u/muL6tfZeWyoIKM+htztDcEKH1db5QzV6Dkdt
F+pDjWC+JTgK+RjYS5l8ETu4SAhy7vIL9hShSW+eem3gbkvBc4G61lP4h9qw
OZWvguhffD9KqjvBNLjGqIhgoeQq9cym/zBNtB+0gGVJjqc/diRVT+aATIDk
kvnblgR3QTSzLSMl7dOT6QRfnbZ87j/nmgG8yLMriCKWm5BvIViP8HcDhfRN
NPS9JyACkgjtn7S1tXeLF+S1xImc86ufdWhSK//gweaZr+IPmlXMhRcK1LHv
s57jGqRAEEx1vKg0xqHP1ns/HVhYJAeFcE3yKFzNcqKaMcxdr59+1ZvZa2IJ
EO+TDNI26FtqL26mcmJ6efE/rFQmBWKW1x0mWaJU3+vCo3bb6pYMz8xw5taH
I0B3X3nLaIhr+xJmhgFLZ3wxyo2xaBWs4CrD3CtGcBr6t3rObPK/jGCIYIc2
Vf6huazNjZnAku1RNTcfB6tJVfRZGrA95O9n2U5gZpVZat0hDTYQL+JzlHYw
99m+ETAqK6StNTd2OZqyeiK9C7E9/0nJWPddbimxQeNJhQPwiDbS7PJQbxs3
1DePaipGknbxc8xOtBukbXLAVSu59y0yoGvUeCvHCyTc4KP6tOwH0uq5/Y8O
m7/3yHwcI/1mHmw5VNVwA8TEz2HpANrWvo69nG3myN0b99FMiFxQ1KMRb888
lyHV/AFIjuyNlSZPltQathQtdZYFoj9t23Kfkjha6ne5MtoCS6ysmxQLyxmc
CEh641TLqiP7aFzZh+GimwR3tTGNJrj7U+rIiLzouTlHVPvUHn6IPdMfiZuF
C/hbGFon+7kLrbIEA58MRzoAGVyP+GvsvFqh3xll0MrtFB9uDqbOk7irLec0
zT8jP785K7E0OszW1EOlzqspkJDh/7XI0G/gDIfD3aCSzkXrcJkzo2M6XCx9
hu/A0McPXSPaawuwCdazB0VFQFP6krgA/Fs/N/l0ux9IuVvIv5tUqp4tFnIh
MNy75vZAZDIDP2O1zUUWmzKX8fsDk6f7ahf5vLk68OSgsvFYTBB0eXTFlgS/
PNc96TKdOLDVJ1Zr0qv+rQLxrMZPNx4B4nfADOdeYLAwYFVjeB+HI14PTFII
ghExgvSgUikWc/HFDxyofqrAbmdZAWDAEXwAfToVUpjXpIaCl753xs+caOmK
apCa7k7ZJKecq9grzGsI2C9KLpUfA5yuEDZOA6OmN2bkSR3FbNFnDId2Fa6S
zBVCpW0+uEtJ6G/BUQNCx/BVND0ESzSj0a/pYTEUIlTR+tT0umeU1y0xHnlw
AIvpVZCy/iFB0EJdd+6iWGpc6M+zNyBEsfuA99tpBFCEkKW5fQ7JSijo+Ps2
4tJS8SNjNWqPqvADBzfx5Asu2cL0mlN9QiOvI19kYgFTtfZIoWAW0nGrxYYT
QqFV0mnD4ZvGkjYfpGwBuJ57eioXCt6+QwCGTZZmefsafBRquxM2f0mhaWxi
QitLd7qT72/U4kBT47ZRZOiUC/11Jm07mSepXpFsU7aqQ1Q/HUZPf6WbI7hD
A/an+DprTb3jRVikIOvhI5ttd8GvWNCNI1zyjPgP2JgNYCPSasHDialbX4cG
FcEKmtF5usnE28eUG6xzySsohwAA2v++yBYDabJfj2y+FrCvTTf5eZFlVuvv
KUd5ncCP3AOMyytRbRskgmjE0+3D7J5GssYjTqNqtJysCzNu4iWtg0Go7dl+
/8DkhsV5hr2QsHOwxSbj258etuTpqLSb7sXeC0T38WqDjaJxjvp+gqzkkbYJ
viGxcOj+9U5b1pbJGVZf3F5VohlAA2HCE2qWkEVvGo00j0FazVQ0CZQHB2YO
bCYheGdtm5D+aCel6KxbICr+sYp1B/fys6NQVe97Y5Pz9tX8oPoeICLQBU1w
ewirJ1T8hdR55xnqseJ0JTyNp1ESWeJMw4hg26P+wSfPlsiBPZzjwFzbD6Je
H9euvmI3qxhsoghePp6teHwk3HHFiaYyj1C3K1vmogxWwRUVWfRUhpPBsxC3
vm5/txHDJdJgsl7AUtOOVg3gWndzcWS5erONNcC0xcNVzr2n1lHt2Cqn7s5b
0r4ID4yaFaM3IaAV8PWab5uc+fUo2e0Rdts1PzsSaP7/fSPzZN5elKJRqbKZ
rYKA2tWJEVaZdji0jRPx5Ta5eCahcIGdQBxlXy9NV6YrieKvgL7nbFiSTGvb
/BFVG3mpVvIySoBU14bZum4XK4wj0/OvhfjxzHFjZssX7BiXRx3Isq1k+TCJ
5iMbiNHNdKoK9w6si6/y4X07TlubOV6sIayUsHaM4F51nyB0Em4yRRn23QGR
mplHhz+YBSvHQXb5dVoTNLe5CSYKYZaeSg1nYsjFW1kbEoHLge/8QNkDyVca
E8X33zn55be/+w+y7He8Mb+4Z86PMUWjj45CTFXFmVFanKEIV2OMaCQY23tP
86cGFdLbDRZVfKW8X12giyMJOlf/d4jVaVUdCOPzd5qBgak/+1kPrhtkZF29
F5bzhMtqmvlcVZ21kz2htFRwJkC5nReJ7uoE/N6hH98CuRBhTicJLtYrfJ+F
gA9IGwrAKF6yo0cShdL03uj4LnfkfbSG8utNvxK7IzhJRO+hvBg+YWFs8PBx
ETr6GgYJ81UEr1ntDcCoW1Cfpqz14at9MEbRPkRyuZZntuxUyMLcEyWXr8SS
GdOdU3NspFwAatKp1a47s89796e+kLClqI4QZ8aEbjU+s8m5hNvXO/evgx6a
DDXk9b/TwYddPBM2UJT4pqGGNeXP+68zTy1pfqlYni5/Cvp/tUSh3VE6ifmp
+3h1uizil6+Ie6tuqJht80iE/naWEF+UHxnRmXv8jXK//UOmNKhIHU9jnhj9
FQ02TUwP1FSdeBLmNbWaRPZpAJJYCSKUtJgmGzDU7yOnUazL38qnIt74XUcI
gMtRigYk9j71oJs3jO66TET4rTTkYY1TOjH+eFsDByw+xtutN93Y4JLlOhcW
WeJPJHk7krLF7884EPfdrYGrDzk6nO588CsXCaKpA9WmaQyPOD3CdqrCzx7n
VvqfgiZQK+qewyC5N/LNBS0xeU4ymYadTK5Bo0UvXIbRbl1242lxBh7v6vpo
PVkgMvDqFM2xe3+8j4QSjUSUir0K9nJHk1hZLLmUSV2i8diwQoh17qZoCZhY
AoxXYT6PcVWf9a1n9R6mjSSD3t5Qwfb6sM0DufNnmnti9wDYoFkPRsH5rT/I
b7KJC9ZW1QabOaVQTGkRY5lcY32amk7WeUbUb0Ovfe9V6ncsbXo7YKgsXqN0
8673KLd8T7n4/LkMyRfVQQ2COhWkrx5kjgJsfAnEBuidUHkFzHQeOj4FvYT8
rxRgGjrHlbJMHdOYpq8gx5Q5IxWLvKQCNUIcxZB9fujiG1SpQ0XV20UTFDxi
s+5//aL9qoecBdd/WiXPrfDzh1+FHHt0Cd+O9aqlW+gf3xik+izXczu62jJ1
GXABs33I1zH32L4ouXflMVV3LRM8VpM+rM+pcyidJOK3rDBXrX16apH8aUF0
OWQkFlpBrUi9ybB2gS29Hhva9Z1abxfSDSUjH3FXJ4uamXbZOF2YmSQsemEu
6lQOKOO/VO09A4u8ukz/DzoNAViuLl9lMThvqK3UeMPuQb5V/Ou8juwmUKe/
nfDpIMhPP2jxkimbmBtEXlOCSA/kLq64y4O1MFPx/Ecq0NaigmPSmXIDK1k6
+5JnL8aC079Hc61sz8Wyl0Eb0FLHCmrH7g31qEY4js8zSNCINL03NRt4tkq4
hM7iLM5GB3Ji2dDD/ZojXjuU9qxvtF5p8XgF50Us6CpVjizoMzUtcot00z4U
M6OiOgXERnwIwTdX81HoipxOO0HZ0VFAuxEJg2XQAB0T2ksDj4gVNAbpXbmZ
6BToD15UuFfDeXFSjthZ+uLUO5wvTnx8FSupx8QDiyycjG5b3rksC2vFZ4s/
1/PmgEfkMRTy7EsoyVXipKMC47OkRrYsS/uTMPp4ZZT5uW+aevS0sctRWPw1
GJGVZlGk+M3IQum+F1ccTU0BYWFNzCNloJh2Smwb4TeVZ2ghqhU+uHk9fOMS
IarqzkvYgDFk0l2zCCgGifsmP8QivYBt9QBc/gIu8UyAGiD8htvAOKJIT9Ce
/gR3c04Pp4TYEtlbN49RRw8ny98nFY2+44MINLMWN1eAigtdiuDF+6w5hqfL
cLgQX3PBGaHPb+wNOUohDtTV16V0GSXfyPxE7BCfof+7OE02lJKPhJMrORlo
cWdH2eSnY5IoIZgS/XE0YIBBtiXLt7h9UIk8WSj39769/Nq0vYbpiECfIaPF
uBLgiVi75Vbyb/9AVI2R9qhUuHO0Hw2JR/iOMgu2mU44fwKOJl853zXq16C8
3Kmj3vQN2VDm6VHJ1t7D+1Mh7K4Wc38hsYFVuIzPY50KF6YpFKAJEp8jgx8B
tKdwof+VvgY7uwtASbQoQsNPdrlfg0u8vczApwicDtmJWre8mm9NH/jX+8sK
g2LeGu4JxVYCA4shItEFbgF2ZjDU8g/CpbSj5f0mDiE79pyYk2i+lf09vv3v
qFbbSkmu/F35LLMgVUwTLZJ8rswRizNFMjjy8k7nuBbvd9q3rkufRugs6eCG
UlWaioHKpqIyb9Mq7pf1UXj8AojaNc1K6iEc4dlm/rOG0912//jEnrgHHG5O
2zz3jyx9DtU8fwLdYg1ADfBssG1on/JPXSfUW0FAQ+wlPrX+v+7yvxNPMzch
EKD5BqaqKan9aAH+hUZjtwDPPM7i8x34nfcTod8AyA+Lw9bRJQ6vG89KSUbn
+07iSrGbsOJ7vdHMfUR5PrOBNPi589WLK96/y1teez4h4gXzaS7RoSM+y9VL
YYPv/Xh6fhafYJidmjsuQ7VORTMwqgmEi8Ieig+AO9mvLNngVoOFRiOxmNMr
u9mC03aOt3d1Wo2dZ6ZuW8pRDZQgRzrqcvBT6CivjuYQx6yIzaq70RfS6UBp
YqMBjBTnjTAyjv2Q4FM3FvpVeimrecYwDgAshKD5INdPxKigp6W9XEQ8tQN8
/ai/YR7t/CZBtkktCXFAa5glz+tTqq0H4hED/3AKxmNZ9lnsjNZ1JNpq3sIL
NNb0zHRhsz5Kew9wwExZPmP4Pl5CCfNYFRzhvCinJn49llpvgebhUaZ2Tg9/
5C01NzitKqUUH4RdvxX9TMUi4XWnm/ledZ1NxIK6lscLfs/OFMF6swoHgKXf
zmdwRickmVlVGzJ+dxunAcMWy9yO8yCs24HsorFrixmI5hbE14pmJziLbJBL
MeF7e1VNxh3/h+eBhfHjZ09jfpT5SLus/Z8prMOjlydSeZssmu01Pwqck17a
OIfzYrTn0KG6d+dfkar56o3nHSXwy6ust6gaJWtEin6Zl9DMf/Iat1BjpCv4
LJ5D2ZhlxH0QNiAAgiSU0GQuGEd90U8bO3QamvczuNhYWhBugZXz7TITUHpZ
gH6ckkggMyJ9gpOyCJaTjOIHwlcI4fk2Jze2qZytwzN5LQfP7WLGyqP/PVsX
iSHkpxMVPc/ri3PLIdiRygYcbcovoZITYVa0flKQcPcAe42Z16FJCACTY3at
YVIpgu0S+QAbDN7GR35zULEnmmCpVGYjLDUShjxAyKhqoU1ui3QmBVrQOov3
n2Yi4XpvJyyWnBVMMURpVC4Is0yjn0qDd6QwNzQq0AmnOczMtdgBasL6sZla
w/eTBHRY3xUwcdg8wN5ciCt78SnxMKDANHt347wshjUeZwEraBDHwR/ripic
q9eG61pkZYBk7UtUlpHdxSoPL85vqBuNSY4EzdIRkHF8dRbcXGueWgmoLvbn
JATW1auuOblwnjNVxkx5lZfyMoGOhe0A1svf7rAoXI91q/qVXt+sr+7BDSSN
KTxkYlL64l4eUAvxI4qEOqr+RqoT4tJAQG960nndNlH8qiFP+EWvSS5QYcXD
NmIFb5YGw8yxTeYykWUXMyTQS5tegI0XIRxDQjCkOc57L115pi4lV/RhoOSE
2PoEG+JYaXG4Nt6FRX2+mTpqJa3/WWtZGslNQLUHEPE2Of2nSSm8IPV6/vT0
TZmCC95gqCRyWNRxDY4DVtdnz3biPemsvLieESDnCYAxsl9Qz+gprLb86pAp
rXGCP91Axt+IIE8aPfVxrxr+PSuR3pzJ4rrjKoUaNnunPMD2IzNLPRpgE5qR
qPA2q2Ulv7bd5/LYl8gSF/gCOTZDvjvBLnO5HrljAVpCDXqAoAEjOfTB128Q
LwQBoTUT4EUzl2MPhIC7vZaoKggnj5MUDMjuQW7UgCEF2ygmn8u1EkGoIarb
uzNZIxUNqQGax/NaxtrNiDDe+q+UhJ7ZPsjI2xMZE2v9BC+bh1KKiLzJjqd1
0ns+/BvrzOtVHWwh+xkIf7ZvSFexHs2cjivGPy1MNWkef8ojiOfq20DjT4uA
Zl5/2WnI89U43Br7+OkFeiMP7Oz66uqjvt5IqO0k7iTA2Ew9WMCT9unpptVW
UOmKnaSMKO+mlXO75gyTEpN0DAGNXMuXGzn4bC1AaLUEgbpiur/v0GasKxrb
uWjNLxiigc16LUt0VJ/r1xTIZZ18yvfAepQuUPFjV3LZ/MGbAEfjSrFhBNLb
+LtuLFoJHgDTWkooDlmzNjNQynvtVbIN/VWQMqVWCYMQn6N2k/5DnmAAnGeH
PoIGBiaJDiw8Q1/VMtqlhRWcPvS+KsUHdTcHh/IzzPl5xraUkJ7Yr50qG53Y
PCg93BbpO70Qctqhv+HddbqzyuoFfK2Q/bXaA3ejxAgdXG9WX7+Tid/L2XJB
pv7OZilJ8ngRwQDfiiePOb/wA2vh4pJCvMJhCONU5rL1BRAvMDk4ityTsXV9
9Crih3sToLRHUN0r1h5D9I+CAM3H03Krn7RSswlvvniNAnvqVbvbtPN/yPd4
h7hLS36nyq+00eVD3rxsgEHBp0Ub+X1j2og1OwyGl0uDfNsqAI5rth9vxwzi
8vLqXxkkVQsStkJA5Kr1WRZszOyTqG+wFdglpKCDhfYbsNko+Xk3haoqSP3g
TqZ1PQwndeJZcKr4E0a5qHLNnj4ibsYsoeUa3yODrVZvz8BCJnNauSc5POls
N5rV2CAF4f3V83tSRR8VlrKhukmHKGmYBpd5VjfoQcA/voZUSYJBMR279t0B
bb+He8XB8YKvcTlLWQu5KZSA2z1PBD1WrRvf3jKzWhK5Jj+BkNdYo3iInZH+
qzPCB6kgm0/0hR4j7oD8pNmbM/Me4v7sbbso2u1oBxxwP82bHqOGubrbmETj
KiCYqZdRxIgtBSxW5W3FqSlL8UsYF+s2n4wVKDRE3z6KwbkcCTfDF40FzUuC
WEZcikDnWxkXihlimPeBPT6Ne+GDvN2CxJXCgCKohDTGkhykFRK9h9+eHO41
RAM7x9tFzJLw2EcsrtlVpmuHA0GHI/N51MRzMgSjrsPCjd0R4vsfvCBOvwCX
GSHZ6sM9+zXSOWSUCW51CUuAquBxYDD1UiB1V3Y2nOayoF/UtNvXmUULGV7u
eEqybwBOJeIYJQL42oC+D7jcquC/cLUm6a1zZMyYq5Otyp96AI+1ApBOgUO4
mfTPdz8BdKBFdh5VObvFnuJDIaBqgj2quB4l0PHnmBBCT/t5BoeBMPlAnBGN
HekLtxPAHc/+9hh2+z5Mr36y9nd4x3Vgw01MfhGfe6W2Z9+zm08D/oV3cYJ1
grmTeNRxyrq9CE71+pwk4RWRUNnjF+3jUakYN2364sAAZB12VnXu+KKNMlKa
ZpXFxJ52I+hxvQaxDyGYDWw7t1tUbYHzGuvsNwcVo8RPvvoIuB7PsWwNVbyu
ev4zBvQ3Ijrl2blaVNQXYRVXI9eX++Zef4jfcaeV6gdWdrgYalCEQOILbmmy
HR00gLW93Yjx6DJDC2WxVztZffDZ8veke1J++2KFC4PE4eyRj8+A+4wHvuj8
eK07VpAwEev2TbdTLvGx/8sk2T7OZqPxmcBi5t/Q/NyUltApVQD1KWPcxzJN
x6b/Y3eboSmnj1Rqe3XuF1xjiiO9ds3H9mZLCJ2qAlYhvuYXH4xfkDEc1zM6
2pNrCUpVYhTu65mneXtHXBznXgy1coB9xIM4k3IcypyHIR5PjlIX1di62qwv
YqyLeQAGfFu8l3MJSz/q6w7jloz+gIY79F6PbEpU6fcl4oK6kavYZIda1Cyy
2OLk7I+ohHvO3COGR3ViHTlV+iTDbZuieYGrNz4leKZBpjI7o7SWXiQVlCWs
rUBihxo5QDOG0JmvspLaLL99EUehtmOtzK9VxAsSOzrKcCyueAdIJpzoHX/B
0a+ARC55YjqNsMNFFxV9qVdlA/nRg4JufnRP3xVIX93Yg316QOC16ylt9Hi1
nAU5OzXYjHwNVuJM6CqqyLl5omfTYRjg3BtKIfiWg59UTQMNm2Yixf0buOyX
zk/6/TMfUyYVXWQMj+XFObGw7y/DyD9n2deJYci9lgDrnEnWs9EEC/Hn1NMB
2pSRYjFZmNQGPLQY92+Mo2aD8ODiwSybvv6N9Bm9gGqJoqCUKYecKjxRuyvc
i1CY0SBxiVd3DmihK82Rta3U8xoTVbB6hYQ4KOt/4AURMwpXdm11KiWPKzBJ
ArSNooGqv2e+rvD/2Qg2Iju06D/7kJ3Fa2lESALclj0nCPqxgdxruncYkEdf
+lyfIQYCakWB4///z8JmsccsScmdXoTuym6xxnDyon8QMi2oYSLBVcCN5JPu
MWwO25TWs52L4UVNJ1O7GWtlPXOGFkPDPzXqvSi7BEwgf8Nn0tfenq0wNuDO
oRXDmjS2Fzk9OaXyH4SdzcIEeUYkLv3+34zZunvGYe6vFKUt/tio1dCFryg1
KkMNqc0s7LE2vm82d+gK7qeGnCjF1JrjYr+hGh/1Ir9m44ltMRQS5+opJBtU
fBShsPLmAJ4Unm8Iu8N8jySaIFcnimQO0vceF6K/8RVzBooBrqvJvRn0JvYP
Juxt6dVF6af1CUTw8hjRDxWLyhtdHqGos5jtCKIztrh0N6BcPKnxR2Nr6+w3
aq4wh28exkwmwDliJgF+MMS8PmmqvLNNM7cjiwLnVskoJYDZf3shP76Sykp5
7njUxkkz9i+M61AHlOhVdWPq8ZpuCoY+OCIYgPboXd0t+/MWs5i8XwArvbXj
/HhyJUd6HbvVc4WfteXYAPvia03icbg3KvrN/VmTfnJKnUrAwK4Al7++dvYM
ohTGQ9INsGV92TD3XFJfl+0ZH+QUpRmDqTZurLJklUiDiBhCy3MosPVoNLVv
4a2YJp1jRgupAPv67wlOsCyi7NcfHDSI/CsSiLah9dqhFCPASOXSJdyzry+Z
2Vs6ZSeqtisPYGtdoP695+RCSlfJq0PyODXMD1cIpJlMveRC7hGmTCIWKBex
ISy3AqZEcuoxBV+dSPxMs/MPWqb0dvqmhHnrCLUa9eM48Tpu3NSv0wdjtvCe
5m7loqurF7rmExWX2R2qA6JNG/tQL3hpBX/f0AMv2ElsWbgcYmNcTimEUZqA
NBYbpJH3Hf87YosBB1yDkwVZcOwzycq6Sd6v5lE7xi+qDfQKP+oC52ymwEgS
Me7oFf/viJRrnCwO021+iCEYuCvZBkjheHsMKNv7w1iaTp7j0bF5eGu4uxzl
kM0Uc/1BgpRAFL9HXdFm3eAd6FStO5lbklII1gFc5xnlRt/T9H5bKBSpGCZQ
LfRg42g2iVrZgHT7xiaMiy3lKhdBPRNbu9St7GFfnUin8cS7eohCwQlKsroj
/N5CeUvRxoqu/u8DIrft9Te6WQoohyE9SGfLMQEG6T2UPxcubPJi0ztD1f45
+JTsGdsr0K6vKQEFvLwQ3Otm70fP77khghtVrPwG9dXBtDGt+YsLJaqU+KDH
nYpbsDvyAB3x9/QICYRvKiW9AzWa6Gjm1/f3e3OkfA7i7NDaU1xsILzgJk/H
rpyxLWwkU/TCt0xyLJCvg5iCGO2nAmr2XS4h4BKu8XUX6ho5WfSfYFOtXy6b
MvdeKOejaFdLwiB/7D0CKUZAn8QPdPGcLzbJNmRJKWOkuM1crWJe+fmCw1/E
qO65opwCcyOBGCArM9rhX2YaMpQRt+F5iwup80OujJegfLfG/ZLbQ0obP+dN
WfKkhFbnr5sr4r0zk5HnueZCbXECr3FsOMbkryGBiVWKikRBQmIsG/EbFrjz
l0CYWE8G3f2DqMxGwgA/px6a72wnCteML1169sW+IauIPSlAFNtxzkKJ4V4b
TT7jEgOuxH9mSUHB522dcG2QeagHSBRdqu9UNS5hBrFoUODiPWpo0d7tLmhx
oCeARj1CS9tVYuXD8QsF8n4Uqc9fHSykQ/6e9mz/YV55zFo0itbq4sdcfSDn
x/1wSHMcIa27r9b9jn6vuB2fXaWYuC5cvuRqzEXghj8YCxiJDktnZdMVNHaU
vAzAbn/t7JfVHUTKCvzDjAxVlLlz7Jtps5THBBnRm5v6AcbblQimpvLotA71
eusaGLmNS3uAhtTRoZdOd6jmcuUW6rx9utw5DNVGgjcYmfRaD40rEN5UEVK6
1n/lzMUYBnO+48fko53L3b5jcWE7k9KWM70jF3IpyfdyGkVE4ZBp0hsn6ofX
CgQQUFuORqp+oFSNt9DDr4DOu5cmskrPwdDoJ9ZOO/C1Xm/7l85medLEBNbO
eMdPneUfVKvKVPgbwd5JWKIZRhR0CbFANtzRhmGNGPRCmHIgiDxbikLRP6FP
NdHITj/KVuYlL5jrwjO+j+gTDxC5yfhQbhDf9XCr/6Rta+4Jyov3tK/HpUaZ
1odJj8BMJ7dUm95JnH7t5AndfPTzNz84admiphqcqI30pDFe+4W3R/Ckm4xP
2XextbuQOVF47IK4zVlQ0wptme9L69YQlDq3dwgsnRk3W6FOXFrULeP2akdA
/czfuwDQ0Aiem0iPh8pc4UdZbfEsA6gt9GnozVM3mXfZLFRbyg69+7A/rg8Z
0OcXrxvFlWpVoAqf6WMzLOnQUkp7lWgaPmfm1CRk3YMLfqLB/U+FBRJmLcxK
zFeemJmLFTLDauv2Lg56uTqGjJHRDJoCMtnvG3XBibeQLNX0VxZG0N1+ErEZ
Za4uKQa4qnx4Mm287+ChBLivTgQxxS89lmFm9tqiizdswyWdfFm5Zu+OPYaR
V20xEvVBkrhr1J/bPohjbTXCYM12eaMsJVeou6pGtLIKgvbD2RO0wN8H9xSm
xxaphz8hVyckDPPkKEbGyuLUo7VNp3FtEKwnO15vLmKVHp3Hc6n4e2uOvB7R
I83Zk8RLxVuXffgK2jPW6UOHNevyck6b0At9QVDDt15BNBY3WA7gLMnEZuE8
cNZKVPrTNAoQMQTtPP2KzEOGDPEyWF/Hi3gJi0Y7HtSDyV4IKxul69e8QvgA
Uttkhf0kmgBQy2wAwu3rSEt+kUxnRDETHJGkME38GzLnt3Zr7ZkGmmwnbkgh
tfIBcFnoFVQos2WGAuT67goQa4PaWZx3UvClI9AcOTAF22ocwIuvBlkpBl6X
KlCxbNj0DKQMttK1Ru62pKfDzcGYr1eLA3G0WlPfpp58rNByTDqLrY7WFLHV
gBjqlTAQq3nUMvMxPT3icVMInXkbE4NvTx8Ek0oQ6VlP0ABJ8hjGNr7Ijfkf
AIMA7vp6DmS6xzDAGfL7Y4dT0jLWXn3Gr5M5aVqd/yhpMPv5vJFt75JdUmr7
IXytRc2mIn6CT5ye30iHvkbDeHXC9Yd9QGrUwiqcLCH2q1Wh7KMsJwJ02WdP
0iE/PPqo8FLFKIjWMhmNMSdTkma9ebPOwu5Qa8VSDiPII8qMvDbZVCizUCPu
BMhKzBc5y8aMYr4gvWzmkPUdOykqjP5SA9QfmepMWIk5aV8LfoGIflZM0LsP
GB8RBopqQEj2ul1OfHHI6cCEu2WrVgbqF94SUQCTGY+q+OfzfDW1I5kXjhYw
i3QTY5mg1jYs33OmaNoF/rKMHIQkOQQDMAalK8vPBNUotOUR8uSa5Pq58vlA
PvAumj0pcyHwpVlm3OflcfsUTH94pTptrKP5db0AJ/IvYLyfLh9U0eok8DEF
o4lDGhYZNQg2tN1ThrgB8TMpoj/SV+uGJG1TRKNlIJgskDUvdBjOWfH8jdFS
J3ppS3TFQtITgntfecG7cPww++Bi3qTBmlEb9XNQjeeSMogRa8f12EyDr2jz
2ZkTZ7MafmhCAg0cinNqg7F39Oeh5glVORI9WMmOAoO4vgJZN3UcQibs1IvT
8PzaSr+4HRAHYE2fxzA+BS2viPt//FYHkRt/JKutYtFks3q6pCBeoKUpruF+
Ap5uTxtzLc9jY+I+yS+WHSSNwVI1NgXQDBukhqYu3uFmEjraT4KsFcqD5LGo
qgKhBIR2dnqGwoFYPQTrnu/9yfQ1K/91xT2O5g6QwypXg43yHfvtCELtOYRc
XKZC8AjgcPvTtbsxQCfL0u3VAfXF7zRL408faevkiq+QD5S49Cm0LzK7nq3N
axqNZnQFNk8tL5VoSZFyl3gKHeXwo1ZWj+fSY2p9g9sxXOJ49ex1brjBwaKC
+hytAw0rQZ/61GQo7UPCQHsLE+59Xa6I+nJgXl/URMma0x6dqBENGEKsqkOe
h1S2a6bof38rBeWzCk5qyRkNX44BVN4uLI8hXzBb/htF/RNOE/qNYJlo1EBA
TaPuJ8h/t1OBlKny86L+Ofa6ViA0AJey5jgY2NwwgdW7gDsUYceqw8sRFWfS
9TgqvJFIyXmu9u9h0o7BHpUJqhRqABY3iQzdV/W+z4TdCSudEX6phX6dsO4E
2C5gIzcyYxXC6cf6lAf5OWm0elvVEmQBrtriUK5E2uizfONGjUkP8kYdNBh/
6rHoQWn403zIAldet3/yXvhLsSv+7g8lJ8rTr3vrpRHSnOqtDwpWSQUZIzdR
99AHtOwB6IjmGEJIW3rqjRLPmSU6TXnM//lDLCUjQ37VkapMvEM9FsJY592f
4jsF7dpnBCv6+vCmiG3lz7yJZYcdHWsR9MeKDgSxTOJ0YjmcYOuCmaO830vB
UeMbSdqxtRdR199gcJCDG2eupL/fz0p7n8Op/SvxMR3ESzJuTRrmri/XpI0g
BtL/2rBLrljGEzVwR8BmlExtFw4aeQdUt9QJvUPrpya6r6ibYcbofvHpWH7/
50dzfpoil+udXEwcYSD/4zp0D41DaQ1aYkc195Mj4IkoLejmt0y6t5/4UDBp
NQMqVWk+sArr3B0JnaETlr3LhEZYximsFcXQPfQuK6Z0ix2CJIU+iWeEsNfg
G+Z/7i/O5UWdSCpDWh/S90Kuhp0f+gRJE6kxzHCKNWXq4IeMNmx52mK/rvbL
2Eou54oxRU2ipGGwodjKU0kim8lps5rOEsp4fZGpisr4brTBhf2bKizv6ot3
IbXyz7UwenEBuEB08Gp4uGc/EvJ6GVKH5e68Geta0au10RE3UdWX4xelWQmK
p+qq7kKbvXYM/By4/SpdiVuFYjq6Ll4Rqem/BXF4UvlMmZ/VRAgXBUDUGl34
xowFnXRdF0sqiuFYXiRs8Sd3WuI2lG6EG1hnP6knguS2ljeXdKdMCBuvgD77
+NfL92PU4RRYP95/9aZNtlaZVyG9tC1OKIJrgtFl6aIdSw+IFZGdye33EJiX
69GEi9VwqGk0UBlG5n6WVmhHtCYjcabeyvHctdlweXXKYSPWFlJshwXSCCcq
tgTOY4UVEdJGso75Mp+gZ91B+st8H29FLwKFRL0rykMbohIhPAL33GNmDg0u
RLFw08ZxgI8tO42iQUgpVmsntTGm+S8xzMh1S4zKwW4B4wvBmFQZmdjkQoXK
GlRHGxw6jhbgLsiPgzagqFKRyxUGT2xE7oo3v9JVM6gobcAxrMGkQwGAO27x
+6Bfu/itHUabcwjRG8Qial8/mm6WjEQwShfpdzToA7/kotmOMsWR/UDsUYLO
gvVsoDewH6Lh0v82iIxkpo943w/wieBowoHit+N4WVMaclc9ogAJtTYaQlwf
70jIjwZkAN+rBDyZ7i3u6uH8x4CCBWZ3Ftg2OC9Nay5feUNljAhhIjglIJTH
Ul8pgDDMtRWylhxq+4LyHUqQzEnVEdgQ/jKQ7eWrAXtZVqP2jUzOBbAL6eZF
M1r97oltloN4GzWRPlBXpbxeu/EaxtMfuoq7facdzl1PbmkQhd3gGP3nZ2M9
/VmyJq91ddryDYlhZttfxDwX0xsHHCjaW+7Z4vgJENjXJKv4AKY1tLIftKyd
13XEEjvbRMxIireIlLdhIFocb0y6fLNNwI7uhKAxnLtju96cP+ds4KtrADhK
B1QZvNAxu/WGX6t6ZULXasMU+rKo2VcNfNB8Fy3zwHgkPVwxC1KJ3xC25HLC
7I8igpNI7sz+ho0IVyW20qArZu/0tNYQcuWtK2ESIa//fZTmmp8KQWQ7g0KW
xinTLZDIulJptMR14bXqWA9KUZnW1xWz5ISK8GAqX2JRAjKeJ8u1qA71w6tJ
eQMRqGbobv2YWCF8oYfsf0cs9TZPptp2W7XTiNcEP4BvmmMvn0rX6GHb7vrM
UjFB+cmOxDln9IRYVV/S/lNaoeBFwi4UXEYNZzVBYbQm2az0ihpgGrpdJNjh
AcKpqvQG0SG6a0w9CLfglOef29d4DwCHJ5UpfM62xajCvKwrAoooK4relkTL
1kKfxL1+J7476aKyBxsYQsJX6h2dFgpFplNJ+lVGFgZ+5mZG8rJdySd0igkJ
Tm4xHkGBvBbAUd8QLRhpLXs/k5lWu6SLfjErfUfwZ00QJs3AyZ1M6ptaXNr4
fuWNg/sX8Wk9QNG6s8gnLtfjSGw870SfAHoAKPxt4bQhZ42CFsrLNe4GRRgJ
AKocRNW6lK19AJAldHEpZU16n6xN8csmtC0ptXHR8Qm+QuZWaDVbAc53HQAz
D3nSCzbemwOf5oMY7wEe09HNFncVY596ECWYSFhpFAk4y7IIF8P8ojzLkm2X
O/TCjm42v7bnxRqyCF7ZLaK8jIC7fUNn5hv/L7ivPnHF57akQ35rZaNLG4sc
AwWCjwfuMQPBY+SqLZrKdLaNBpKCEFYPAHlg63IKKIodhHCKnRth1QBvO38J
jmdH7eoUYaiYPYIqiP4/emF/mxyBWm+jDur9p5mItyiPtHEeyw6yY2DFWCQn
h4t5iH9u4f37UdZhaxewyy1SjpnR/rCO6xcGbEeq8qj5XEumIeyzWkTLsXDA
6yGRoyPpCYsDd7sj+LmwAZ/uSE5TifDw5QsmrENzX8ZTDsHaY+rNXSNXzIEi
TqNz6NE70FsOfcNcMqJQKd9TO6ugODRtuc3Fbl5m1v8HPJ9MHp6rT8FcC8bA
XI3c0+CiaJk58CLjzXaLIINTaY2Vyk6I+UDawMP0Q7rPJQCA76RXVludSgyu
0nsGaTnMlQR4TIsuyFObDSKda8BC4zISrxiN0ZxSNDws107+2cPzq/EL3tRB
TWgHajEw2+4mTVJ8Zvv/UecTclWG63O8ErIwGaKqS5s1/HZ2F6k7OBnBfmMS
G6V3RausYmcosmVdnJHImJ1oPtozG27frdTLCFeM6T21Z2VMip/pw0HQfXAW
f8HKxbNS1OgvsUMb0XCmlXrN4lc9TmUmIfuimrbJtG3pXPke+k2BhIHo1cYE
rKKB39sl6Y0yw2FvTYD5XST3SpDADpIpj1JauJ8Y5nIfseWp3jgBmPq0jbBu
X+NbwVQQxTrSzdKHO1/dQx1LoobnnGLcbi2IOGtvfD+EE2JosoXl5rCD0Twh
fcnjUmWxuxMD9r92hmJXT5vVofhOuHHGt9KCl20957KI26vpisbk7A+RFRWr
ryT2l5EuM4N6kObnW5+Pn76YMnQnueS8ssrW1UizopT0oCACxETPnkzwPaqc
LyHkeuStH0YBU0neBCeS67TrdEVFpn6f5llmHl02NbzgKleOZwV6vfv2WrlM
9L/t2a1LiZzZNH+Cgr2KPX89iSsEYn68BA8O5j6KstAMKYie9CRbLSMyGjY9
Lmc/00xQzE5kqpL1ZW+k1Pua2LZGvgBLAXVkW+6b6e+Eo89a66QSQrfFTgop
MKNSgt/nJu9gfYMzhbJ+c0fWk3g1x8cDWuz7sx9gFA6DDhJhXId5iVeXKtkl
Ppj9AGlc4JaQnSdBEdTqpw/i9W4Lfh/1KYSobQyPHaDFQsT7Fv/tZBOzASM2
5R/EorvEKlFjde9FT+EQo2K2At/QU5c0UE/Sp9YrqoigVLcbLBVOymaa6P6C
aeXGEWOayRbx9iyqdJWS7Lpc5uRxyzbBQoSPWEqTt+TOXPgpSRscS3aj8sJO
YYo4nEZs4QXfrkdCnRZMmWkzVxGABuR13gN82OAQHvIvXoY4qGXWGLjA4Wbb
LRIF9l4t/ZQ6J8/AsaePC08BvNGUfGD8vZJELeqe7onQMjWceld6OmIBknn2
/M6khSI/876Y61spcRQIf6W54Prw9hCFkZz6EUcJ8fvxfnwx0jV030OikK2C
pL26C+Cc5vCSatevmbFdwq/ugaif3EJnIriD/nRv3L3Ix5Bgq82mZ2d19ox4
Qamlg1yaycuOjh2yIYZi+fH291e5hNoeYmE+EeSf80Ueb4Gkb0h3FIq7gnb6
5Ddb2PlI+o4ACsG7Ehuyqt8JGzpORhSYJ3yw5HpU0zPpYYmKe1ME4W706KU0
5dGICMMXM/SoCMfxhCfzBHLozV9LKmlQYoifZgo+g0tkkJuZYdvBH8hjt4Kg
INlvCxwvymUNabEW+FSlZvqLR7SpOOnj8zCfd4Kj9/AuDOtNVj+ZtsnYQa5m
oyixo2lAfiOFC1pgG7n8/M9VUIEyar5Mz0fXCROglttDse/uCLBQHe79ClY0
b4NwKPvN+3L2TqPmE6m33XgoLhC/nCKzsBzlY/rGu51KUuItbE7N41mu62aL
pSpEyuxZ6UDceKGkyj9IJsi8gpPG/FtK40AYwvPyM/qEUsuZkkK0bJxrlAKm
Lq707DenTNOtlaoRTLNQbgb92m5bQUCaq49WTFtZ7Pa9KUxGqHUnpdr3+m1V
1TpzNpyP5ke7jSL4ZChcSn0AAQ6mLl1Q//ei6JZ0n7WbCBe2hkKlpP11DUvG
MV4EAHfre5Sm51oQPxlGaKxi+tDfRGifZtoF2knBd9fHWO0NC07O9o/M9fUv
bFiHl0Alop4STiX/W5S8MD8763Fp8jTZEd5QnkSfyJKjRuh85EAjLec1bRbm
9W3R0a5rimcbZq+abyBhvWZGzzpXecUnUJMG5PeFDPua+cnh7NPYyB+awxfo
ZRnifcnE7Gq6Zwhaquc9teEQBl1iojgEPEUNCsnB8Ca0PWlZALvSWhGsPywH
twbItKKMyL2YlM6vMcYvhX9r51PUU6cidn2hyUfeQ1rmTPyRMX6ckImYOkUh
G1Q/dkRH/QIsXMpP7Y4aDSAEr4bmiUnfGQCZBmViOFuOdO9FYul/6WLa9h/k
4e/6GXAYonD5f6OaG0i1O2u/MUe9EatduRSzkiBA3POCLH7NHUiykO64tiuc
tYA6iH1zO5Jvh2fvEmj4G2d4Wh1ma44JtTLvjvtbi809ihSG2mDJuH/ptFui
0XWzLZmbYATKlgV+xt9n0foW/TEHOzSvVCPjLPP96C8+7ERrpY2BJ1SLCSf7
hXR7R/TU+kq4OwuczYxNj0XPCZHQdsg4op1517nsKnSwEXQGKavTWuieWQls
tlH7TOST1gd0X1pJ8VPbobWkdmhMhUkd7CZwnq3XMVTA6UjvYpyUzy2KS/PH
aPuSGGCBo9mbwwPNhRhSM81R6QOn1fnSdWu6VZhMqt/nkPqDlRYJa5UK9VzH
3V/h6CEZyl+yYlF7g5COaZSxMv897DczJeL4CXzBbldVzdbWX2ItTaN2al2N
xZrccFAR4heBo+Df+2jtlxibeudgKT5v6767l8zwGLsAJ6cTQBWR2uCZeCx9
FyauXanIdW61tLVGHV/Fzr+Q2uxlLkL3xNUJSqbO/IEPxESj6CM2J8zjKyDZ
JZPWgAA5/ypbm4VCXIzyLhpw30/FspWC43zrMHhQ2PgNaYnp3Logj/cVVFXt
CdqbsKwF2PDHrvFgM9q7NSbhHuHaGyemcZZXGzT89+oVYNTOF8afROQRX6sE
0x02m8+p+DSevsGDvfYvsG3CEboG6OxDuwc9vp6nTX90aCNSRrt1Vuib75HZ
AwXhcuKlbFIxBZy0R3D8AJ8hFDxjd5YmuLPbOzY8IdHPQKt0Ex2uEXR/qXyw
AEkmrCl9R4BlU76TsywePs57ZxoA3PA8td1nMKf9UVrd65hccRmuBaXttCr1
75WNq8x92cHhQQi8NOCLFnWNK3rmwlXEzgTajo7rjGLQXlhU7BhZzcRNoPEc
kQCFqXfkmVnuY7dVcEp/iGAzwCd7ssHUBkwjEpDZ10VdRcgkbuYCNrW4OAZf
aSBy6v9F4OMfy33erMRVRnReFFICwW7AmaLrZ1GD4phcnJuZW0dwVWXn/f0/
DLOLscD29yFKPmn90MqrsasfWuS+EMQQvxKi6pJ5taS5merEL9U7rsn65Vih
qLWC6xOuw+MF6d940Xn/TtQTzp7RWK0x40n2/DWvXOxxhvbRqOL4dT5cjEk0
eWpSGqBv5lbKQ6tKVluhM9mwf5MsgT0/Pux/qaWwBrAPL/A2xk3tfV7/YAgj
UlUPIvBuuYATQSiJtt9TP0LuTCqdOa6XTcwCYjsyDkyB1flzjR5rQ8QXIx6M
FyMtG13oV1FiKm5dlh5L/WoR2RriQrJfpSgDwWFgxnI5YmIZCnYKlotBN+Nz
Bn3RTnHS+6m1fzamCq8MR1CiF6mKwmUE2MYqqGMtN6nOuow//G/Yr0V3IjkN
4zCBpwD4xD8tulkE/mN23QcfybD68d8riy/706vVJZwXQJIMVXYc+NWbto+e
v9rP+wWN0q7IqtCZJ6W7gznU6MUB/BMo9HtbiXurJq4ZaNNweRKDmvfFgxkQ
/agMzhsEc8giWgM4NJhlVVwQGSS2xlHwCLFcFplnWu7gRPX29G2DjDXwnejV
BdsV5sFdNqgeTUnBfqT4rIs73fKNXrt8RMxfQTSOVE880jWa/rqgPWKT2LkF
0vGpczR3ZNdcUXqWRaFrSrbp0z3mguyF8YmwdgiqfCgd7pv+Ukvp6d8NCmUn
CHvqWCFXzsYFZmomDdpPZUU2gPg23Zwq39OpMTNgmCe14uygh3Dm82ju5YXb
i7Gprg9Mcve7ain4DWgqfOpLxV37JK3JImeekVqqFbtekHEoe4+73mU3qn3q
AmBA3r3IaIP2K3C4kvtJWrxr6V5IOT5QjPfTYlc0SfqClNb5DYA48bCrESj3
b2sqM2ApBgcVky/WNukibyZ1cR0U2u/vwvRHoAhRajBC/ymwubv7xZOwKWjb
iNM0498xFFfHTa3ia9A5AGZnqdXZaiuKkMwFsCMjRWC2MbWEISJ95SpCMBG3
jmsRpTCXwN5TzUN4+YQJ4I1cybP+6CPyMjC57pWKJO3vGGvVL6TwEwzg06ep
fdP6yzU/z7lRddG0Kj/mWIrx7P+aH31zMSq7YF/dRVIhjw3Fc6MIjeLpb1It
QXHtkugqGsGQcWjs14g9uazNBwKDB3iZQzxmbDdo1f0k0P/e21B/Y9C3P+Eq
/wUx8WMIuzvKh0RRLVjsfCEvmpcOKuUtFG3PCHRgTrvV2EZc1JQq56GiKtRS
4cAFi6tznbEqGN9LEcHz5RT51gPEmET/Vdc1wptaPOnicoTOl5I3/cbo8qkY
gwwRrz5j6enbMB+/7uJUF5HHxphxe2GiW53Aqs8gSOu1nLFHftXnwzAjmJMh
ykas3PBtapIA3xGxQej2CPTd1TjkiG2hWF1rEDlZZxjSn0c6W6lGoo/l0ZBH
oQkZbQA2jaqndGFSWHWQGRprGs/ZUgzrZulJe8OiPVngBriMONdrclmNLsTc
NPG7+GdeEKzYOJAO7+uQWo8UTYsxIlufCFhtGY7NtgeGhBkZtyRpjzX/DGd8
qB4T325+9ZS7Hgv3VISV5MzOVPRBGBa5KUzngKwl/MIDz7kqAx7KdBpm9+6w
8tDBYpLGaB7kg+jqazhCdhAdBZ8wlvhLdEgUubM3JIMf8NdhUq8sovhRwGTI
iHVvhagUeHLOHYtqbQu8w7qFhQRfBFtzSbpxfrlQ8q10Z96u/jBH4y27ssg9
taC9cZTJDcRnYmUPm/m8VDgtr6Q6kX9F3Cs4SeRgKkxCKVT0OpTDC63DhBMw
QSuT8t1Pr2h32xAiPSA9OUZw44q3gTJwyHTp/Z7sAPEdBmMnMyoLsU/ouY0J
IKqNIWJEKGcOhrTMrAAY9HPR3Uy241PJDMVZsrEu5x2F2m7VgVb/cQpa+RCz
QDraON8PsGHk2lEqZymrQvq2iorKl55f/PNrQhFaHRTmuPXJy5BOqJqicngC
b0cnxQsarU85/AB4hWyhTqSvEXgMhFTxKxH0paHgusMh52i9gq4PKoM2ctld
Md0Ka/OhqH8sBnCSl74O4cbygVxBl6rl4TXcjru73XpqF2zfl3tAdPWSlIls
bEq9783ZvwZx5k9yp4nSkipHeqfoX/k0pLcjNmKcWo1Jp9bY/m3pjunMrCK4
28E43FhtD3mowjDmoGns/44IInQCMZSnIqn0OgOH1+3a8LbE9A6Co+XHdzJ9
+Xe/IR1abInCRVXlE/Y1cvWapm8C7VLVxHki/DKmNYyLZ8g550Pi6Wb1pCQQ
00l5qRW1MY1keukF3bJDx3zxFv329Kl6dZ7oa+TPi0pe0XMDHygep24Gtsn4
HR0LMt3xExuP6dliVSE3arlg8/uF4Jtm8BJzX2nDArFZZx1Azl91SZON7StN
3HOMRyrsQt/LL+LRwLX5Yfvd5Izq/SqWasfI9JNYT+4ATLN9A0XEoQraJlLM
mOAEaXm+j8LUtYpGKyOa/26CYd4aggQbOLWPPZ0gVmrpx/QZXhvN2CepFsRR
xzVJDz57vLfaqShG2zkRE8eZ/CooUa/BZnpII14hOpF84gTfsPC5xkWdS/U2
cr4tKEHSs5QnV61ECB11uS4g7EUH164AxMZ/6Jsdukanoxwr0Uy8CN/9yzZJ
g1acV2L4ButL5Xz2dKJAsERYWo1nJgx8JYqHfG+OIcocZd/RjsWnblohuU+W
rYd+BDDO+lzPy2fMDMlVdsFIdEGSGx/vHLZ5sPWF4nzV/AydIV/shDLUG+OX
/yAiTtwjBq6/kvMaD7DbPHl0u+LQzgmnZ/tDDmpAvzpGV4MhvnFs4R9anaam
8K29Drpcdxwho7Uvt+JAkzZbjyXkuabbv8EPHLUt4FC+viSYTrKM6MX53ySS
B7UFUT03/yU/hsSa2XbRNCPAQGDSNuX14FLiHaSYY4LkeqyxjCsQFdT32lGP
MRpbnt8Le61jc6i05pcnMtFtS/wifaJk9Qo+0IU7VvFlL44f7G7h+z9ulubp
IAspeObpbrPk37FdUmIb57spJLrkcdnpqa2MwMwclrl39lravGHsXnjb5jtm
O7N3qlHwt/dV4DZe667N65mpEGxEK1uwDAqRlCs/U9pUPloRRnzkDflHpj6d
9rjwvhbsT2j0k+Xav/CwN70CfcnHIbgNZBDu7j3fxrMwJlmd+96ADWr6QkUg
QYr3YcDOpdEp0s/7/GotpbUS0lRqoHCS9PEEuGJ2I6KS4RD/WnFf3r327ljk
jtSjHyzTPgiGdZwwiG5pX4A1yANvcsHHNEcLfJb+CEcidcK/KuMDKv4If4xQ
4E+2ZplfcHfeLXEcsrSNoyULZZCWNGHnHwZtHUJeD+cRR4AK8gZp948Myjfl
sz+vrMs88p48SPQIV8GxOOSqs6PIwIqyYcPV8D2MLESQvN15ZLQBVbh4sPQ6
oNkFW6F4Tm2sdhgd8sZVbSJ1BoXGahA/it4iF8e5Han5BNl1tkc6vEvLw7fO
ZCKzw+kUU+KrGr8ZMavpyFqpQYss5AZCcNh5pvqnll1vj9sftRjcWEKqWzgp
Jifi3Py65d6wQOoWXEOx/QbD6jzPbwNmpl7bNAwenhqfhyINdsnU1dL25kzu
v1HIGnni7PLil+lq8Yy/amNYRrexyYNHdncFwda0TfP/82aTK6aL2uHMC6LD
PCOEMPEORrp6hWem0YUUjrW/KPfMw04PF8nWk3/0VI+gy+RRIkeii4NSqJDo
0RIleibab5JmpskSoMamrYNYxe3C5GKZlFANSA9x168OujjFQ6rHjYVjC8on
eR3dvC40ejwX7QOD4m4o/UGTRkayj3a3zRKo5AVaZXdAnktCp7Msa55W78AE
EvIlDGLRjqHmnEzJXDDRqAm5RjX/2iOo6ry6oWcZhBl8ddmEb7RXKbVULtY3
DriQ/07Qlo8scATZfEgQsTeSVqOLKG551xVdDDGwlo5EG0eLH3L68EfH0Bpz
ZkMUW7/fIswFELNwTvX+Kf7zrUZTLwABZN/3Upzm5ZJaFPlR2NUaon2rHLuU
w3ZmFEj+KTVmtZ29t1FUU/7V7YW5P/+VioykhfINgIaopbB7zzwGYEwTyVMT
ZiULcGFqttzDMdIkpY3ynPSQ9dV93uA2IVIM2MEbcUa7GPXG557MamSXQ+w4
ciIMwgwKBAqbuQvDPRDiLAydINDb6Wt/9obB1aNR0nRKDFR2Lp06p4FtxHPN
+bXO/PkLLdiIR/lrZHJcMWqF9uH/PSpIyhb9IKYJ9vx0hlnyk/+ZCq7ndCXg
gltkE6ZKNYKwMqRoHrPD4HQTRX/Gff/nwqevH9cvrHOFJwpBxgtay5Bof1UP
6Pk93RTf971j3Jsrt3PSOxdMPo5gF53tWL9k0WW/ZzmmsAh3KfHMUqB3lAdI
NoqjxNKGNta/7qerjpKqXieynz4hs341opArtPmd2T8Ddc9C7By8j3pQ0ST8
6HuNexNUx2wmidojxqs9xcaUmdFnj07+lRJnS6UvPyXOWjIf6ESJoOCUJj/i
B8IJRDpL1ixMS17S3UiKhZSP0riMiEYUHuKP2QmFUWR9sotj3mzJmVb8/uac
nhL+QQPkNwKLRFUx+uYTf5OY9nyatuHkgbdcKOFUcvacEJis+9on/gQ8Kkbs
cv6b8qWG/5KLAtlwbSnO11w/ngv31FOieBEWPs1uOgMq6Nxa9QiFueHxSX9/
5Q8SN3yATeyWFE5EofHQf2zLvP62wEHhaC0q5Pr2DsKTJ1Z/6MGB9nlHKigS
ngBLzD+4J0qusI19G9D7a8aFK09FE1NlmHfa1XNS+Y5pNVYYnD1HBEAvInn3
nm43uVsid0Rot3s/PdDfrVqBV2q3+Zm4gdkWhR/x6U26rL2wojyPTt7qkGdS
EEN90vVOAHD9AawaSyqnIkm/aWz4MtiGkTNj31Y79bVkTFwL4dTwt4UIYf2o
bLxePyYAZJiNs4sVZALMd7l/5Rlh/F4usUzP+/127+j9ikM9vQH46MW+XPKl
Bs36y1AOQzTpvIZRYRNjpqoy2gAIxM3TLzFaPnbFRcHKpetQH6yo4QAYsi6Y
+DK6Q96j/Jz2OUwV6c/Bm9MLPAjp+yBdu+e+CuGDBOqoWcV32l6t4cjt2Y2J
7qjQSQkar7pW/SKHQ/aUAn4Rs0WfuBB1gG6BvoSmcdmbcxLqVif1QMJ4PukH
zY1GQGWI5l8F4AfOxvvamaGvRDzbUWMaHAKtmg+2E67X10mblV6/uyj8rkGd
kCu7IeqEGeOUncO8VpSJYKGoCXt2W4aOTE+DHY1i86Zi1LYp8+rKFBv89vj+
jOaDpu4tHZyCi6t4ZqceNoxA54p9LxE020F8aKo4B/SF9rSprjKPz/u7ONr3
ikbzJLMB1xT/0WKkJKcGAMI42+vS4lby+KDhL/DY5vAIwA/6YgNRUnEkxFmA
5klj4wyLR7tGsBqaRcDmsKo/HMHpTQmY8nl+HGCZ9yqm0zmuxvQzoA4VaR2Z
GLOWQndT+Xilo/sJMYrU7oGQ4HXO9vt6Jg3y6ibDPcuZ0V5hDWzNSeixQtWP
rsVHgdhjmhTiLLiHprLkc5Q6JpT8ot8NlRmFySmfgvYajbVIAWGCCHvqe0pE
ZdP4CXD5IoUzO/nKmGds8sXNw39CWTJUs6jrhk0aIQ/8DWn2B2vboXdabZVR
J8rksFP0Jzm/Gdpn8IzuKoai3Ly+bIpWmuQ65y+JdslL8Spjodt4qOvK8ufP
1enAevfHgzYURYQGGixD2J0GEg4Yawh+gU5CjEuKlE7lC7F+haE3DbWaMJnS
700AU2mytDHtnIAXKJVwEKN5jSxU7gacSWQKrLtq+haDZU3OYowYD5XTofI9
txJW+xEpqkCJnlShHH7JTSzvGgA9Xsx2XHfbKFWeo5vnQRLQUOVts6SqetXk
gdyTlwIAs1ozV5+jpxT8ASMCcs4egDmquha1ZN6udWneVmpHrzoTZAeTH18L
o2gpjUjfdgD3fpXvtBP5fNqz+f9d8/DaqsbKMzlU7CWjm7h+6u+LuO6cRBrN
zx0jl4Td3KstWUdcribH0igR9KAeCsEN+L8+T4tQ0fDdFMMoQ8urGOXaPCZP
Exzdf0J1600CDk2J3yqbdFa2eMhQGww9G+sSb7VvKd+oaYGY2RwDHKDzwFyf
fqf0FKjzIlFcMujDYd2qLukSia+qkoCrY01oeDfkW3/vd773x5mQpA0ZJh3u
mBByAyntW1ABHkCum7p7vt4i2UmPoly/ouuVX6yO1A9l8PXmbYFmvGBLsQt5
aY0q0M3mSVtqfveSURDNJSBsgA41bxlXzhw7Igm3+yxfp/c3ByDll0hje/Vb
mJB+MdLx0cD2OGtAJAtjbDDCMJI4FdRAR9pek3Dbq9vbOu8MLd7vLEtaSmYh
G30juEzDXNaxPizFslAdxFIR+p7kHtvw5P+6AeyqOQq14DwpqVHeLzh6PbSL
O/7PB3dL2kuTJ4IqiiBifXnbmLmrY9CtbgsemrLaVVMP0wDPK0HXXPlerxWR
WZOZLoVOkZ/TrexsLX74sU85pEpA8YnsTSOPeeiA7uHQXK/Z8wH6sMZ6UvQX
e4a+uiCb3Fg2QmD/o5GusCxD9XUoZ+RIbPGsSHnfeyvr1yFp0xlCNmFjXzFv
jn60CAZzkRXPjrX62Wpq9Q+f7Nku9n2ILkT1cmtneI2isjRPqCTd3MOkiMZ+
vGuGMIH2ZJD2rJ9YkL16xZ3oiOwtEqVc//L7BZD/D5oMNhMI+PO+XNavz4O1
Htg/735QaYxBXLVQiZT6ZXMQArDoDAGfLdConAj68RWGXzT0M74a5RdgAKQx
+F8wdVlgBFTTuaO0fihce4BKBQgHLBW8IeV9Aainzcrv3B+wa2FCA5TjLJFn
eM/WbXXgQoMVHfP9hcUGQu6hmOoEfR+oqAF+DFTibKNvZL5qcIQQk5Pll1La
NeK6q90c7nqIW65PSrrDIQXB4tbl5pGM8Qey5//dbBpKu3CSJTcpfzZSxfdE
7a9XjkA6gBC/qm/lPiArAD15Tj1ugNur8YWs0U3KWjwT/7LgC7yY3R+wQNWh
fwkk8/ZHWAs3JMjaI5htZ16UOHSjJAoiKVIzb+PysdjEYhudqlXyxJwPzbOO
b/kEhCl+zmMMy2lxTECOD2HIk3w2E8YQJXkuEPKWD5UI7VDuOxeOa88WKAdR
pPHGPbsjezwN8pgmDOXplVg4UoAxZL62BOO6muAt4VGlXUpppikB/ctmoSAE
sQ+mfX6+v35gF45s1x6GbDKoM3vpGtSZ8QFlpcKSpeFuBX0dnRrAXztAS7a3
heqFKlfeIJEj0ZumSqWu1Em6ddp78IBA065+sEZUl8tLk/dpMWtsv4L8DuVb
g1io4+2KWCy4dmBj6SstMwLalDfOczTfiX52IwukwyoKnzkOwRAHv5GAqerK
Qv6xTnnfyzYxWPHbAfhjGFHF6Xbw9rrGdSaZ1Ngem7x2gZVu9CfNRC79TqY+
uWXAW71OxTw/3EpN6h56nxEtB6kV9fWsgecjb+n3r/wF9LjPbpSsBb6b3QBi
1VeR0gV9xEyc2aNo5u+7q+ISMsx0MI+gVjZJ4Ej0r/su0knbB0wSArEQupjh
SPmxG7pdJRsmjdz1ISRLkKINASn5ktPQ/p7vmQg83F1pVr+87auelN2SnlNQ
aUrjzRCfCNfsFm574g8hx2zhOQ7G3JPMxPo0GG78647pVACAQsfbWVX28V/c
z7c5/vKe5GJujKU7ORapTLv+uLrGRWdJtC18iWRqwtTR7IWjmkwxfc1Hbozf
9ZM2EbpZxon9b2GmRdryf4ZYxbzcPjd9wPsvqDke2XG49nEmFGBwm2gI3dVO
lfU0rcyMG5xvPwSIQ/lsd7fGkbVLW3hIDrhsYghoK863Mzwsi3iusrJQi8HB
BkTpqA47qM5oPtPttzNpdsE249IKWb8a85CO8sVdWNbnbzt/XhQAtsKEo2fx
tIsduwjv+UD9x9KOClfGzS+3QExbDqQsMkdvte/nAbNxvkO8k2Hy2zSZKld7
85Lc9WJJH7zZVM2v6QFDuidNP8bGy0LRjYeOOgHRoR+rBOiL2QhCddXjPmtK
4BDkdQzgOPUkyYIXBwdSni226os3B7wFMMiEu8r6RQ1guMMMM2kyJG5I+BfY
EMDaY3HiYvCan/Cp3L8OruVQ8SYayHw3ZV57BgGYpjiE1giDeRX5AMoLAauo
bnHZLpKTnDXxIUh+NmeaO3A44BbAPudwbsD/0DtTmOFCaeCmYOCd7iy3c+vZ
7pRB9Raruy6J+86TYJkbeL6uOEFpWl1gdhcgC2I8HT6j7mpaP2Q6py/iJDRP
99nA+SOPKa+wB9AnfJjy8PGwjN42rXvLRVqpXfrO5sMbN7zWRZ9MYp8QpOtD
2XnpiVV2fH3Jq9QK+WOtvnvOOox49V12LhCeqvUim449Q3XKdxu5N1QQg7nw
RFM4yijfTYc10oMRD7IQsiMloJwJVRqwvbIdaZizXUeC+UIybgSimZBZKAbf
WFoZPUlnSw+luR8mttNU17W1zNGgX+49MCRpFJjAcYTZxPsLS0mDhAXbzBHo
RTtC7Z9X6cU6CiK/ImjNRrLvmiay+JqVpf0Tj7qzdD3teE8iScbVxF9NRlly
eOo5NWnzactsNyAKKVdGW45OYsxegxBh5vL7y3ksQDbO+EWRPiDeleX53QPc
OIt1pHz0KCI04mjAaBNviiA3KOWz2gcVdYTvI1zk5soJy3wt5OG/3Km0Kk1I
aKK594wY2TPgzIJ77X8IxPB9PbfaEh3GhqJ2jGyxYtzt63XgKs/tJvtiaTM9
A24E31UU7TvwIZhTl4KDfpWmJrTdptr4LRCCVwA+v8rc0hzxHl3ZSsNncgkQ
pDkLCG16EApr+iode7rPBeDUMCk9elqZxSdswL9xU8X4YjbWQIaJJhUu6WNW
47lkufyVTiGLpm5t8fJYo3P1/Wa7qXG19cLiYcNZlzBvTU8nznTnJj9QyxZU
NcFiy0rMOB02qY5JmwyfbiCcEPAvGybUPirYul/3fZafsZVU3+HwYdlzNISp
vTo/T5vbSep69BlLEigDAC8TZLQ9/l3TvkD1r5QyiuaQv1D1qnMEOWjWx+pk
sw+vQef/j4eVCJSjvNgTIxYd1hx6+0/RMKcCOX49cUwOfr16J32hqaMu1VBk
0k3oFDT5Tqdmouzjv0GDGE4PxlnLspZDD+u6Zhku0Dra4oJxQnO09NqxwGUE
5tagD2Y4LyMssYoSbfFV9b5GQT/TnzeI8isaNp8RuZedRFTwIk5cjPlyt7xQ
bn8H9tP3Oy4rgg0204oteDqp+AZ7Her5VkZ1k19Sv6RzOqdYNs46n18InogJ
y1WjOhfGBW4JHUd9kc8s1A9MIAKHbcRUAMxVXipsto342wxPCOyN/dBkXU0f
nhH507PxejudhMXpSrGrTtmX+rVHjMX8JmOYcZTSavxBzTaRz3vYXh5cm73a
M2/S2EUjsGOGJRTbTzV3LCRE/Nf/47NctSLimEKULaQ+m0wukrx6RML4FmD3
9rXCEhamBC22SJ8fSntbmEL2MPTrUgsbYj9qp+5v+uaTr+AdwXahaPBivKVE
idCGBiD5uPF13nE3TainWE8NBoMNHvIfbWpqz916nIfy9JuWHGeyjxmEeQ6V
LEJ+jRnA6IwJccO9CiG12JSLc7GPT2DfOligG3rMz9gygsuKpcmzazYbtQ0k
DC/OuccVUDoRkG6EinYqSNj+3KWmV08kClBFEKZxc38dWqQTFByWU0FZhNRR
SY17x0MA2tlUsUFZ/M3mn9698ibRznlPTCCgcBiwPUcKFx9vTwOBcw+aQqM5
CKjydEGQ9gMNwDaA3WBANPGRfeS8ZtS8232reCPkFsd6yN7WvaUK5Y6yGysr
Y15sVvrQUINB07IGtFHix2qvviBlXbRskNp98om0NCt4pEEYF3nL7Stc0KE/
NWq731Z3moTycmmm+gS7iPjncuzsYK7ArT3E85ZlzYyX2zxOLCjyfUZTNhym
i/VaK5zC0lMHGkSj2A5ShMyT6+4BiHkKgxSPqlG+pB9Qv4PlDdCO7+Mgk3TO
ptaoJfb+2bOy0f8gZ/kAN94QTvxIeSh1nxjPGWqwTJZtHJZNm4IPXsI7pX/D
nyI8GvWfKAw1MxWRNZDYz4TqzW/KFs+NHFPy5/y9UWYvvagKs/qp1VXQKcL3
Nf0v+l+xjZfBDNvoy4dwhbZFWTPKn47V2NudMKUWcHGv5P4pMM7qc6YDrVui
bXgD1NLzpgnQU2nTvMaNhSZjZAD2zdfZ+v+qgd1Mk9gn6/XEccHBqu7QNdTp
ii4II5eUJi5kpo33XFCGLjws9EyOnIggebmy6SZZ+VdAGj2Tnkg+5XRaWL0v
472/Ev6igQodZJykMp3o1rXNybvtqegSMeoBx9x79zHr52Ug9h2VhkiqJR02
Vq8F4Nr3EBTW0JZbhPX57SKCgwdohB7ebmb/5ECDVnnqbtAfhXBJO+fjvoaQ
fTUE+RqEIBNsQXxndzEJhXvlHVpY+pDJ0yeUslJUlyOxcMmFts6nX5djJdZr
7jX8T3tB5WKkkzQlPC4NjR3YmB/JqqCgjjz5irneyI9eIIrS5E8u1ox7gM5h
B/M/Oc15iz30obAfi+jiO/S2aoSPkINTCreYvB60w4TRdtNOoot3c0oKjEWo
VNJID5aKc3tDeK/qbuPaUFVjrm9fMl2y6yoKRooRALnb6/SWAHQ0DB0QE8fP
Z1pT/PBUXBWK9mvxwoj3VGTtyZRbFET1cVxCzx85Az/1j2Scm87lfFOB/2JW
fjzvxlZ9juA/JtIMFnz6CUtf8XLUJh6CjkddX4ymSCCfAe/yNS7cG63iFdB2
MdsTZBR2S1CJjwOAjeREHGNfNwvC0+g45edjBGCkVbrxQlJfjUAbyFeAo4vD
KppUDKjAjOmpDksVCrQx5l2Jf27CM5Y3EaXvWDARVRjiITCpw6ZTLPUcU9Uz
FNDTzmlfQcB8CEDYTIcvSvZmJGjCJ0z60M+DMG7uubNLMY2AsJVXSQLrc+TV
GHiK3OZD9Chb1Gu7v3nIlef+I2SAFzvKWlBiWcoypKX9tyNYQjlFNNlArzVe
lBv1ZbuMKE0FDcFe+RBRys+oOjruKqI2tPzT+mjcmeQPOk9XwmbZTAvF1UlJ
+WIu0HxMo5e4iUvJqpcb8lDF5QXui0rUzF+WAeOQarCrs01Sz7gPAQmjBaZA
+9mN/dujRigRjr4A3bZUhrZCNfCwJGeezfwqaqb5A/Uo6ZWaZyolE0KG7J4/
4hnuWET7xQ2Ob71GlC1BiKJtzXaKcWQ2mzx+XFG/Ho+38YHyd4iM6Lqkb8gE
tF+kEbq5go0evWQ3O4HEa8w4NForSO8v4aFsD2oMyeJlBx/WuyZm0rq1X4qH
riNHo1mI4XYh2iB2rzbbyLDnfgpU1Hi8yF3tlZlT4RI7wuzTGfDKx6AljmFB
4EaOO4jJSYkIMCxLoNAu2Eg/qwReqFeCs4+ulpYkhPIal8GD7WISlJ98kCpf
KH3hGeQh1Sw0A8SVCq4zaG43xlvGvUWhGuhQHxFk6bugS2OvTigISDfNIT0z
qkoMmJUuJC1wRdp4hcWyCcbhU1FlrRRZJ1hyvbqXJK17+P8LDih31ojMimYX
YVQ+X9oTDC88Sy0HEsd50lk0jmla1OEFrjCcO9oyg1PHnqeeLehB/ymTkBcO
wzFEJVJqQ4mRxLJ1lGM2Kucj3cWWBKGjLbQDY1DTg8XXC6qN2tLNc974HujA
Skivj0uJA+sH7oKH/VXdT4zSNc7HSq0LNfsLe4y7elX9JcrLMBezQ2MxdZWy
mcGvIHAQa9dcf6i586VavzFyf3G7VLSHQq/OkrqHw41CJ3jJaNWFGKxTq6+V
rjkd34wwpwVVqmBxtgaj0BfKeBHl8V4NuY/CSiXyMMs0qfTjnRwpNR32IOtk
2JFLzaqxriHffYCESQwNjUAWbd9rWA8j57nAQphqB9T2YDGzLVRfwMqkpI1W
T5xbgM29PJyiBbBBjIkenbK/kUmgNJUBXtImY0jPTYIPOGUeRN5EeYFigAMq
le369Icudy13s2MXuberyu4tJ5+3CN2yDfdOMCaJOdMO/YUq1c7raAoJr9cY
QuPspMYeNc7yhQZtgoNd5TPT9BOl6PcL4QAh2uzeOtHrp8Y+HjfzfXXEbAex
ZJFWVt+miYJPY3n1MzqcPA332hdE5KSktLhbME6EHlpZZQdNerETqGtyicaG
Ei8bc3yNec9HdHPA8ai5k3mvuyRx4Y8JsZpGW4xL9SNfQItSa+V09OxTMOVc
HZy00TLL38payTiRpHL6qPUvCk8OktrKWOas2knhkFm5UQXEkMnpoUzuBa6c
D0C7vZSO8NsfNfn1lQ39JUVIbrJq44ZhLtFigM3ueps2DyqH7BYHybY4EO9n
87sTfke98WtTUQ+fSvn32ZmennCVoGsw9bQZNEx32/9ItvLJx3oqnKVXCwZR
MN6hnRZEeWHGaGgAVcGLutrj3W/5mfAsu9cEyF6pXH2QK9YG0RgAY1OFPtCk
z5d9yJGi0QLM2DBhxtp9AfYRS+tZzPTCTIvdz0EPOUZpa5drTI7thrI9NSbx
UZfpiYU7UbmnbtgWwDQBmzWFtGmmVaNIQ4w6iKdyW+l+6tnI7z837y4NJ7R6
3LnrDVh2diD2IbhKvH6sLOe6Bpe9h3Rb0ExYWrTyTYFurxCO5cyKDcxAGzql
2XnhWAnQqwpOZP4Hy09CXNRkhK7UWKL/eX1/yl7Ivu/ijcbrhRnlBDF6eeLp
V+IHVhSXd38vUFLQljMbdV9H0giV3C9BUZEpk4B//TNHFWaluDxT/4W/Ag4A
56fo+N6bLxXSMIvFCG6vCQTVE0ankpbgPy+beLfzbnfagN4ZdJ4zdpuG/RsP
pyOR9QqXY35ZSRZLUnrKbuPG3TBNKNHtzccsd1mRlLYe4Wz8YbmDWgjyK/Gm
vNOwmvhqsCs1aH0IQckmWkOggtuFj4qWzOpJla/XkieQ5K5h4oFT1LKBWaDf
wyb2xpnbt1NLUXSwQbLTmwT5PE46MAIviH6fuVTBsRfFg95cAPH4nlegJ7mJ
9oQdGDsqqqnvtv28LuWQ4zPFKz7YGViwRT3bBA1/4Ga9uGfhs1qrqP7tDBoA
Oxt9FIW+bHEMjiT+ycxVf+Xp3RO1ZrPItaDD9O+nTZ7iM4jKlSFuNFeMB0Gw
8wdn2GzSsLSdSE5fAWaFBSQmJU3WSEmGPc5tkr2U4qRP6FqWYafCPZBua4eW
7gekIhHfwF0lT5JEDFFVz0sk+iaC9gN5C+O1Dw0i/8u1uKWrN+Xpf+PJ9tD0
UmWgMeQ8T90//JrY7BC1Uz/8L9yhYHF6jBDPC9/dd3KglsBfcQGfRuBubSvU
yfuh8vImlacgKmnyFjbyv9BzLwmzqR4eSu4GA2Df5AfiQqTN2XjmKczektKG
r9UUfKw1YJKI0JDLE2fpsc7TVQS1t5jO1CQ9xZfktvvrvqv+MAPzzgBfwopS
5SMJ9rKajUffrUZzDz3mY5zizspqsaYNTG339U+B4d0Mcn0IZnia2iFMqcSh
LCajWVBMzFahPM3IBa7kBg8SJ+ersswv21lBnycvkA2r1V9hTCy4lxaIQOHX
g+hKt7U8HWD2+Vq/DsdFKUcSZZ4Ao7bDKC3uzwBVqcMy3v5yHDk/yJ0IDZmw
aKVPSUQ3HH67HOE8GoapsiUYi8/L3sN+d3h52+VPw4B3IPpnRHbVUtZ66oKv
IQUkUbFre8sY4dw3AI4/TjImq4MfQywPvtcuG80rIL/IIn/HFa1rFRi/OW3y
6GfxRcOY6j7Sl7MguAKPVHLvgdwjUCZyMkF8PAp9DRH/TX2+V/5I20f0PTED
gXHUBwahJ2qV1Z29XVUZLNerl131ls7cX6xoE6xr4keeWKyBSrj6XcrRoViu
2Sg4YTxvOGsc8k1pkgJua1a1UUXc4jTavdEQWCKSrN3AnaQqCpcgdESYquM7
8TLjmFmNXg6Q4uSxdY3VOT7vFs2JEAws7KhzQC9usGL8+cL1HIQIxEdjl93/
wC4a+Uj1VztyqVD1rk4VZMX1t1kfDvqgwKjbSFhBed2qVC3pWmz6TuXHk8cL
z/Z1n/8m+fzSiGyqC35GEdF5Pmmu9CiAOH/LGKSDAieqtYk7N2Q8PaqKQhC5
2wzHx3OhiB2YTg5FYDi6Om0a7ZuKcLTdSLrX+uEx7jBEryXIZkA9S4dyCqZg
XNdM31CHtF54tDhT3ISqr0qslEbRXGp79xAlwJsds4fkE7SgJAhyXOtz54qO
me8AJIXf4APoATRL1VupD7pgywdj9bWPwtXAcLMnyerFiPqawOWNsTDCcdkl
bh9rj0f0aiEnYC7PFpnRhbc5P4DDw3WixnFuI1bWSrVnqB43ktqwj5RxpTFA
9G7KaoMF8IlXGsO/a5qYmJ25OTE17IURZ0+L6SPEtimrDOGvhNenxog4yop0
bMsEwoZFXYfz5gy4z4b5kMSTy35ztXCeZgATRX0c7FKurSFSpGbq6ct5dZ5k
w3yF7SiaR8iL2gwkdwXCTQoboiTRL54qZ2oNslM8nJJ7oEZug7u+66jVhCDS
SO7U05R6VWSguCdVh0oZ4RsNuHOiXC7Z56mjRIEyyLmDJC/PSGc6UweXHZJB
XoyiyAjUofBuu8n4NXw661kAy+qa+seLAdgZT7p3+THCmFmn+S4cI2daA002
QdWin20780sEz9xvKUuqwKafdh18yHK9qxPVX3d3Vn4tHob5A9oQ4VD2csJQ
9GxXlMDsPy5RyeQE6t06SGy4kIxHFVgxACVS/z3HeYq3wSdp3gtRZG5bPCdm
yFf2E7zm7W/zGeY8TKpW3K+NYMoNoqyUL9k2eD76/+ijbb3sEUyUBHAbkDVL
oilAFvRlvWm3xPZYtdGhVaWnKeRBBfUl9NNBxB98H/oAPXbAFx7l0GJPel0P
5RhKe0GtdWIu2GdmTiYsbV+h7qGZNjkpNcRJU9dFUUAuDSXYU/9lzZGKn+wm
nkLVB4B5NoqDC/WmDVsyaH3Nos7WF/HkklV+wA1+ooHeM7Pu1viRzrVHCwk2
PASjNt1mnSCewAOm/POisPOeqXzDmfa9heXkg3yid1VdwRVVv9mXhbcsTIAZ
NPUjMriOLCpnIXU5ELMU1EwchtLQLslMMRvNYOt7KOqJsS0l/ytYxeFGtPZu
ZFnJSwXHHFNu0iOg8WORd5JCmPMHT+SHJ/hq6U50/ZVVM/gHCF/VNQo+ulmf
ZN3WHj8qnNe5FwPmH1Ij1P7bOwWN2phDouElfJZXCWviUEdYppYJ/4cYtPW8
ZSCbJvIC19uAkmET9UPONivv+JyBDx9UFsRkYq3LnLYsw87uWHmCVKZrxNiI
NwIpR2vGEgb4ZClg5Lz/oRCRd+sdjuZC/FMibEblxSpiFFlR7cgmM+c3Jqc+
q5G5R2YJNTeV0GqaHgI7mDzUI/KF4sptzi7r5cDcNEMai+A6IzzgMOUJRO/6
56D/YqryGqbvzAWbNAEQ46nnm6uzMFE9NbrUPGfWRmuCEGSPWUMVXzdXtgit
m7HQ50CV1hd38OagJZEXwHNnL61CSq4cm4L6QQUw+bsTku4bahRWzf4JsApL
VukJItyrMWzEOOZuJUgvfqchc1CrDRIDPHabVpDf2iZ4eTnyAGKyXzjQ53Vk
tSLVS0xFnOV3DIukqKpB6ax+cYG8748lPaSyolg9spB/CyVn8NIwpYhttpsB
nxCrBrxwNADnwMRNykwCKAPKZrNHeNqGKvQRjrmNIIjMwnvTuuthpzxAButp
2yoOSOX8IPVn4+EWD5Itwb4aCVjQ1QgY61fgHOfJ8RIYpDMMCgJHFLwcYfju
ba/NN2fDT2UbTXUTPlZrLDY2Amh0SpndzlEzs7DJeZBW1f2MZ2QTbP4LDcCr
+6tDu+AkYGQyBdrEpN9ZUnJ/CpeKw6y0ZpIqB3/RLpfP+cSbDhWViC/wE0dC
Of7BUEkPFxE52C/mDnN6BngAUqx+sRov7aQzrXLBi4BafpQpzBmv8hT2wx0x
ImDlFhAbpX2DEJLOlvr29IwXtWXhrggaejvZBnQ9M7GNB8cCr8Nskp15JeGU
I3sSQyRq43sEdCQYs7kwiHOSiz+Uf8/qQjpoSATlGA6KBPi4csu90QaF9vHo
UNkyyenjvhbCBqpVTUceSEYr5kKJEmtsAa6VOuTwIZmVVMdM9puBVdGQmgI4
QPNi38FqEzhjkAgfNh/7QKqdEejG+diow8xyFKUrT8MUQKYGeOJnlcztfDYW
g1GdKGWYQ20qFlbCEowlla3rj2AoJTWjQz8/DUK7A/kLKRCMojZx1b//mL1J
YX6FMi+Qi/KbvAN9YU7RZJGTxX1E4ln9sSK1JbzuQQgnB8UYlmTMP+wVzQ+g
drCVxfhF9JUWXx2oCehOczoZOZ7ARRcpXizhujDq//YNBmLQZDOl9bD33X+J
QOkLOBhedCLoNymoJbt4YXO9bp3RBrwj5NRVHwftBNQfcEUQZ0LZT8ZQ8Y32
YCWsmjncqjGDipvWreRYB6sb3RKq72Y2oa99EPJauUKQHkMBJxQA6QzHWURw
GX8YPaDmw6E6oKMkqL4S5i9pG7v/U4IeF1YRW/2nav5Nt7QK7/PxKMTnUUj7
1oOSuB2jxN8C9+uuOCEg58zMeFp8sADI6RgXnrkdeZ7dTcQukMwyntvKQxNX
TCPr9tV7eYtKk5Z6zsxk4p9C0MHFNnTwgEyWY7qTrarPRmVJE6+QGcmm6YrX
mTU/XrYWYSegg5R6IiQyLhdI58oKtS7Xzyd/YzOxmzY2QUHfldtKU4b1EiwB
wum0JzZ+3xHYZ81G066SjJOfxopI8511LkprjxKr49RaC7mWgDDy5zR1ff8w
dM8YJtpB+GdoOuPapDBsgxSR0PyjfbDsQatrDnEU7KU8qthK9caa1gskkbvn
W6WMzeOY8jgv7HwqQufI5SEA7NA0SkfJtpVdqdHq1Vclxtvpef2tU5ap/z4u
q2IHFHysTCtZmuN/E+vfKEYSvNNd0ty6x2vn8dLxBUJ62rAYJy+HuR2s1hAZ
cPJfrDHUPjbKB1cWdB2kjdEILChq6lEMuOZKuTgow8bz1pjcIBwERj3cQWJZ
t7tKt59V89VED9wMeTcWL+hGm7yAorKIPvHcad2OQQnh+r9LULp/8EGnRoI6
W8+Bd0LsIMpT9SDGgU3W6SAjoC2890NBw+uR+wvQ/nFCAB7dEcXBoSR+Qqqc
lcz8zeU/S1fS81z0VSZa2ee5857+i9OhfTY4UY45mDRVzQfp+cMjhSmeHlrs
qhFBuJKuMot3up1QLfpaJ0udd2heo6LNr/WjMwYTo0OQzwB/CuGEYFFspcxm
nGPmq52NSHGCmdYht/gxc7TX/2QMaU2Es6kiiT8tszadBkcIGZuJJ4lkt8ZW
PaCgmzXo42lCKTjIo+DsKhH7h2M1gN7Cy3kZ4iLKElymmIQZZhzV5Q8PNZm8
oyqGgN+Ke+issHVPYciWGHFvRqnB+DL2XLRBPb6pdtNB7gBC+QOSJAmh+6kh
jaNKfgeXBkH/Jx6SpfEtRTjVK0yM698wmtCa4EMkZBNOUur6V7Can/v1wMV/
LMcTg/eUNsgD4g6ttoM4fomAoZJAMmCsGOZ29i/nICrfaAJ7SxsHuej1KZDR
LAJyVhv0Dqhfn7IlzMX9Q23T8PQcnVzKyeesWQrg1OWoaskRLOePBdDWhWTO
IAklSyBuyzo0o9shYWs9Cz/+v2565xObsS8PIyekg/eTC0pHo87xB5fV8ciA
/ddV1vOo414C+ha1xjFET4NJ6gZZ145Nw6/TDd+3wVc4eVBubje9niC/tQjc
x3h6PmWDFqNoQXIdz/21fFEnEUJM6+3WpQmdoPahonJApaP4oE72qKd0tntx
5Xc0qF0yMXZGQ6Vk0/9xMCVJ4d/L4fPyDMkNt6SFRKXMh/P5J7nwCWRhMqAt
pjyLzY9OyI9UYFRhWDDLmazKveFvGBWBejGaOxftJlFo1THPn4VyYi8IpW/a
IQidvKJMo8fcij633to9XusPf8n//nscLWZAwjlU2l4b2U38Bl6eAnKg98TL
R0ecLXtw94B5cCxMMw0y18q90kidYUG9c+AA4aaQNdxC4Tzv1YgdSvj4kWPe
m/ucuBzxa40SSq4o14WES9ezeGfozJ5OeSv2JLeOq+E6ThS9JlpkEZ7InCvB
ebDSrqivLo6uWbVhOtpWV1Hf3mbt+G4D8Lwuif5tkSi5t2DUc5bH3PVNDGXm
V9Tl0Kk1VdzlJxhCIZuh/RfkYi8NYj2HrfFT5TYm8wn4umLIQAnc94LtupAO
4i1dvmCKxFPqCqfYow9ZVSDzmFsqR+rVynnP96RIAijEOS+MALDNaYJ9gSWX
3jqy7CsaZ19GkQLRFnvkC7nAHVeQUa1v87du7hUAjz3TKtL2kaksNKjGg/P+
xVkUjIz7m1cpbRCtLNENEL/Fl4l03TTbYAIzJZ1eunj3ZmUC2EAMlGtD14Sw
TGI8M2bXMRa3zCfzuG2WSlpLHYnut7iEoZaxEiFqT/5Iz3iGG63ovB7bvesl
19RXCyiXWhXPYB2mMVt5f60VzeFRvbtfEuZo4P8QgcWdGFuqXoQQvYnlpjUz
RE8dne/IPnWbQ69OwwGqGPRoB6z+Wr7gF/EmyHtOWDiuMmmP32az7TVjWFMv
ZDmU3cKeCqSxliPhF5bLtOzi/rRfknskNzCIxAkfDH27c2jL2AzBW5zyqpfv
USobxbSqrARa6mPWlxOkI73QygfXTlYiHgJrQi8llbCfraV4+lvfGvDQ+Qyb
BR97cUtVXYgeXpd8Qv2RIR6ZrWTAODkgnqhJsJ5QsT2yI43O68e17KjN1iBx
STt7k9OOmAE8G+N46QOw9MKOFFCDRxRxii1YPoV7IxzT0iDmtpFAqXXUOMcg
n4IbXqwTTzTUwIMt+MNr9dntlxmiuFXepmDA1lvIGdFYNocqLh/hl+2Lx+2u
VUmMiapSici+OGYjbW2od6TSHq6dImeeG5zBzyxtm/zE5/J+Sh65BWdKeuZu
AAYsYp0S3x5HXlxAB+8tBDhhY0kIMMWPQzHUHewnRyfbV3lcKXEqiavKwGu8
u6C324awxoDiXc8zlpcWmtkLjqZe9seQXiZdfvD3UWCtFOTZssztaxfq5uOm
swu4T6VYV8GgCxWIdVDeeDhr/kwLa/qrTG/hgJ0dBU5QXRYLktnJgsmJ2KLz
mxNWBtpEeAgmzf8EApTScJAtY5nmu7eBgrRTtug2EjOKglD1mrLXXJ8/BC82
7Pw/SWxRLoSnTubexfyl9TqHYULaotH6mAIA1uYSbRqZO8RPVGXJ1LkvsrfJ
f8eqjJNjClK/a3uSlxc56rsutoFs8dU2zCLQta5K5ATH8HvhZ57rJWoTqT1s
UC+HS90hUj1x5UISHfVcze9l7gIsQF3zb90QpZ2qZSIcTrTwb4mI8Hhs+93i
qTwzRN/vZnwuMq7SfNTSPw/EdmPEyO87dNCHRrQSDcqYHM7NNyLVV5hVXLb5
bQza2FixIRtiWak3xXzk+Zi1gMSmyBFe4//bPB4LSkumrMYmRT7Ez8YnHs/J
MUnB8DTBQk682z1tZu9ky/rX6Ya2UgOBRmC6ndWcxXpmPuJdz53XT3ptYxS3
JMlkPPpUA0qIOwsCc5zAjPJCDFMhUpq5ojoDOhFodbKT7lY1aAwZsdkW6xth
l3ouz4k0UBLb1JLEOBRsCbZCMCE989N7DWTceaFfDiORKl3apB9ggLcarLHL
5knAmxe9qP8h01Zw+8WbhDTXlFTwuJ71mbZFJRZ+6UWdJTkzRgm4ynfHdx+s
MaP4JVPSL6rnfp6pS1kkfb2HNCmTxWuS4+2M1I/O3dmVdYobewp6EVAqaNqC
OTaD2iL5f7ra3vtw48v/KRKUg6sJE7fP14F9xbiM7j+q8hcyDnS4kboR6g3B
e7LYdK5kb6GEuT/EboNmckKAV/AIyahBo8UIu5xtzlmVXGkFx2k+ilY18LCf
Vr/1F1QbuBkcZ9J65y8Vhz1rW0fePIIwSDDHcXcXPZ5UV/dh/tukIxoFNKhq
EKy5IjaIiq7EN6r0nlb4df3fYmhBlOL5unhucGlBqXmDp1Ujidh1i+2QOW23
ueJgn9j7GqcZ0VmovKCqp8niuuV6uBVvJzWKDwg+3xdupZ2BUSpZHwMLe6jy
cgxnVWd9UG+5LeFtgm3yukv4iFBpvYpjPQG5XPLgkHfR+v5MTcrywd8KFFmF
7exPs/+foKzGIU94y5HVqP3HTP8/NWRwlPpjkhyNtaiOmc2oH1WJmOhoIAdq
tQ2/x2tL5VYx8EJx3ed44OFE078LwST6JHXJwL/YiYo92e0IBT0K4AcWZlKP
6IsSJkNQeVFrHkPoExB/sQ1py/IoiNKA2sLPigxylzOr+8/UXi6nfIieXmC8
Boy/MSdpq43abOTvXSY/okLuD+Ijd+EXL2gNZu+qhEf8aXkjxWs5nTsEAWHK
h5iwZgZmk4+RRzOJJEmOlbhfL1TEyljJRQ5iSzLAwxkNW0/9RkM64W1zVNOs
t+sAp+LILWiEAHgHjMgqYz3P7bfRVkooRXdnz/zFjyTnAa8th2NXNiy6SGPM
q+iWXlbpENr5am10XEt/1h/JAw56/RTFyQ3pr0SnF3CjgYk177/AdyIET6pg
siQ72SCVS43oVUcDAlmw06aESqyQRi2Gz5cbRqz9tIojLG/8lKYMOxgthr5x
PRrqATS1TbL5Z/M4jGKqsuK/G6KpyEc1TK77exIfjwP9PzfH5kvW+qhe/N9O
qcuEXpGO5bYu8mfC7jPkFKGAToj6kW4nJO5i4I7CU99je6UWjgbNGWeb+TCi
/UgC/fYLG4NSobJC6Zczb7rwdku/yTUyg9kXwHiThVp4kMQ/9YTFVvR0VZ+2
ntt2AYhJXQOdz1lQ0nWrFsLQYURLmiTQH3RZOM6sHm9hkzI0bcZYUZxWVXtQ
ZGx7pSV80y7UHPcIPuazeRFws7ka7nniP3wZnKVcdFfTrqDAxZfJRKU78Hpb
Ye4NUfFGuMHqNQ4Hcbq5UYyESMjIcgzALqIvEcate7m1OyF5/RY53BxkoDU7
UaE/QMNROx/p6V1suvHn/8+oOaq5dIWxHMqk9OM+q/uJ2tU0P1xkarsE8mOs
nVQIjn5jFs+asppl99O5nzl4+QjvF9b/WF8QOVaJIrCJ06yBCn91pAnq61H9
drr6ZTf9VMXr8UG93AxB7lB7DuMxWbgWaSFIrw34MrBsurPBo1/e5F7wxq+q
5aHiqPcB3W59XhzToc0naHlZEeAO7ONhgtQJ3cEBnEfduviAvAepVh5D4FJu
oAzfIbHMa+evrJcceAgTS2uc5gI1/NxwhLvzE5D2vWj6dB+3+I6YcWK8HwIV
FDjgGulOEw195qD5HXplfnAjBZdBJV0jqL/gjz9YXOhRgiRuuBtgd86pMicH
suz/3vbsbAvJFhiCHYETFPvrTuS9/my+5Wl2Qt0rBxuEKk4SRfF9Zjs9f30r
bokJvYtkiVIgqsT7O+n9cTuLOCpevYGCykHWSmYT4v6sB+I/BOYPHO6NqxHp
VT/4p9IOec9gfDDJU9rh3FGpLXytCUWwN8JShkFN/WHOs6GBMyActP7l4Y0k
Fim8gEVS4La3SXSIsW/nYS7SxWK0yrqPRletxbwAtGI2meKcH8Yqu4T+ej5o
e0a1F2iQca1LqEnsKNEAVjV2FnoPkSVZmznt0GAhfbChlerjeWXvboqrhmIR
KFt1Js4l0QJIePyzheUI9CDT8rvC9XqKwDyFZLd51I/8pQZj/Qli8ybPM+SF
YM56abO0yjgukZX2oHxhuhrvXkYOzxCS6CP+rlgiCf3HLxVWy4tc/f3Jemdb
0U97fIz8fP+BVv51Md08aqIzQznT9cB2BWX6+gKc2gpgKccdzaFx1s+uBtxg
5FI4sZChU/y6wteaCicwvrZU+RVpBjiYGn9d9Zapd7Yvx2/GIAXikfR/SsGa
E98L/0ElLqJgzsXr2JSdrooZglkU0zMV+9cCkPjQXWS+JPuI+0fwNenCKTGp
Q/ixC+Qg2cAwPVhHKJ1oTA+5Jw99sQpT/llLny6oG4MYy7qg7q6YwIKKagdp
k8tsOJDuvxbBxf8lvgJp8lCP9eU8mn7DSi2v+t3QoiVMRfQktyJpA0qtLtD8
NORaZ8EXh5m/n5MiXXY+pg/c2f4Dv6zDhiALRYQmGGhCwIH+cFh5ptFMUZIo
8Zz9QPzuX0PjsWiuaSbw+OBondxTiPsix2z7t08YFnz2z4BPBQ3yiO2aKfoc
7z3rXEak0Ryu5HD90Av8xUWhx5PoHTe8Ik4TCCbXhr/n2fSF2mdeQXG+YULc
impchow2tYMRz2FOa1VY//tByAwrZhOBUdWKRQh/LtXbarAv/gparR45r73d
CV7DpyRJ1JxtaSgRpfxePgpNLqV5akEABjBsN0RyIm0rffCEPKFmIfme6sc7
uLBwcd6R1kUWvhRsQJ3V3qbbFlefP9CPn5k0sgm/f6m0WoPqKEX6ZklA14iB
eW+psUe72vvIs7ZyD1OmCIy+1Ni3+Tzz6qsKdXs56OOIJp3BQ5e6lvN7jN0f
T+aBgYVywD7eFpDqhrcbxDorUwNFQ5czdwGhyU8YSsXnYKWgXlh4XXP6Eavc
uudayJ0Phzs6F2V0sKXaOvE5S76rtBDmrFfhtwLuUYLKEIQY9cJZAdCYQGvh
4NhlIWpOs6LejChEvoAK2vxalOj02GMcD50bU38NtvQZeN7tErgATyOJHpaz
ubY5OR7be2YTSgK9jh0tq/eThot4vzFZzbcl/qT/w+TW7RsTe4Z7dEKcNvnp
2DlD+1tBqTS4UeHZZDse0pA7OKwprOEVMlVnFis3WsDfyR1jsZTciF2d6av/
22+BgvuQqiq9IDFxvCOxOChuFhTHI+2TA97VfEVvKOx8KMGtOUXBrTLC3Rjs
TLt7KlKR0rowk7N5iZkvu9LH9JhxkLzppSEhj5GYrR2o0w2IdK+OuKvsuVdF
5QnM3BMjVr3N/CoeLkRoMBdljKe+1Fd4701a3VIHd8bUTukMmFlGV90XeEIb
Pn0Poic1SRwL0q50LHSZdBBU8pHga68M2tjRlCnTF0Xq6ga0AmHzYp01d9v/
Fp33uSv35s4I38EP/Qt5pSBZ5DNRMei566ToUPzGoK0oXQv/qpE+rH5aSGEk
0ex96mp9qg7ZA+uvSWoo+2tq9HnEmE3x01QpYT1fO8LNz5u0Jo61azQ2n8jH
n6WSUCpEr9zrdH5G5Y3HmPQy2RopN7/Gniksxf+lDcMKbw80U9X8bxOToq67
n8rJeNnopy/tzTmliVj75bgCMRsZQ3XSWKqZWdnxiWbVQqxQKysgLMoB8Ghr
AX+GLPYt9iEKAIT/H4mE3rg9aMoo2V8ohuiCGLgbD5siTc+Qv4quF+oHEi4X
T7HPPVva2n5ddINBjFj8+iTfJ0xJUlYuzhHijowTSe2Gr78hjDLuOOmRN4OH
+Q0t6fb8USk/S1GlHIcTLF/LDfRWT9QgNn0D8wG/qY/sMmVhXCF75wpGVnEE
SpLD30PDczIsMsVgcpW1O4VwfCOj8LzvaF3/W6OGvNgsyO3qz0NWI2p3fI2v
blK9e2GtTdoQLkzguFKddBlVfs30MPqjKvXwpduF7fuoXSyVJH8r4p7DAouM
qQrwvM9L8DEMIsypI3jTMAZSCm6aXnd5TgzYe61A0jJ3xnVvb1auwC7Mx5EV
Hc+e8r1acePOfD51tIKDK2MQLI5CMUlji/aeehLFU5o4lpXyAbRGpIin/tGF
Zk7QtZ5THnV54RX6cTor3tQq8dOCAeFRGv+NuQFszfNbSSfQoY1TZMK+Y9xb
Z2+GzTJ8Qp36mn/Ag2tLbzvTarC7sA3VvxPbTajuRhhm9i6eVfZTEeZf/Dzl
b3Bu1D04wx5nIB9MzPIjWR8bFSAi/e7uqrnM0N5hw6EU1q1t6EGGXnMikY/7
7tIMKNPaWx/cRvKYSX7fPax/r28v03b784YNAN+kUOnpCxOLdQs6/HY9S00k
r0NcdGmMCasDf+AbpDb9A4GvL4u9IWIpFzks1e2XZEVaJedrwSUdyLg7cwxh
sKTKaKzQvPVZtT4fI54/KpNcww+ZiN0augeLl+zU8ciVcdkmzXipNT6Rhodz
8pRNFvt+YjDRd4v83uFUOqHaP2Ew+mAq8qf0EEXx4Zm8pXDsdDEtkEDODFaB
uqeyX+zdukt9d7QxRTUIADeu1WdWJDIt53CrvWGd4bdcWEoJqYIg+FZcm/u0
L9/k1M5J9myQKXBaAGid7wYb80wt828CugAr4rQ9KCvYiwy9UAyFLZAc0WWN
syfazYUSORhKmc00TMjeIYUOU+/XHticpfFw4N/Fr7aw8Ql8bNnDtWAnaRDG
h0ZFBZNzwX6NlVO8KA+/C585pGA6hz4Q7ixol2JvPI/BAhP90zT8eRN9govH
o1wKYNoSYoT0zO3tGS57+RcPoR3Y6NZgmvAygntigieExcwaTydyQltsD1gB
Donr+/ImJJl2G5uRke3EAukTrv/lVJJNDlpE976WfvZ33If3TT3IF6pqcWuN
uI/wh9nktLYZVf7UU65Pfo8UO+CD5hvh+yMY3OHJiNzS+da7T7oTEmyIubFe
u3xJHT9QvPA3LBti75KLRnlE0ipVTTl1HNYp4naaapuIVAKHt1FUSM+mWXst
pJKagheUuN1DwMm4KNb8PLefqRwLq75jzdIcHS52bTunK0+HcGgg9HFm3/ed
eqsxgOtLid6ApbwG4DJ8BreOq560KYqBHAIVmNBf0ohEPD+rR2Lm9leG2uSK
Fw0xlga8vBK0zgFWTSqtYQD5VRE64+9JR9GZDbIV218YHRlHwC7GBVM1LH5m
sOLS/ESIlCcO+fU7W2SwVoPCYE6EmYQG5m1catlhoTP04qAMcAeoH9rT+yzj
zXFpnjWwFpHSBq1gQzMMvttNvwLNqq3gg9D8oDZNNvwoD2IoLyO/EE/TGMZP
/6h6OOTwuKOL8JkcoH7b7a7HZo7kGAW7R6kEwKHFCvarqoXweqUnY4/+O/yD
kPX3xLZvrxc/riA5sstiCT2QgdC+tPN182RTq7IIHmZCbR9tXn1pLy5/7wrM
CrgrPIKOZ78An/Vse2ifUZwiyt+MFMGL0sL6XEx3VXDIPvsy6aJIZ9u/b6a5
Zwyh9CngmWCCoc1JUFfK3JRu0mLiV+nchkcd+QfiIqMpX2fja6Ib/3g5hn+p
FvfIMaE9f2Yds15uCznIOKMShMp/mGUxh/bJH7W1L8FN3O2huEBHSd66hjJi
T4YHEtg2fXG8Dyxi3f2G/ZZVfG9ZK1LmRc6/+8AnYq4NE9AeSvCf2DhSnADq
Y8aa9SbJdhVJO52b/mVBIEIQGdZXbrQbV0IG+bkSO9d5AbC2mDlpEsX/1KA9
nAIjG7mDU9/p0FHl+cIyvVRhgC9gKuPors6bFo0eNX9ZbW7IgHfPGZWfumnF
1kiro+wBXNXhd85HCYQy/pWW6XKWgJCDMFdpF/J0FJz+Dn0hAgmW1+LCPJqT
hcjGJScZcBBnpq43xJyHu2excNSx7VQ6cvIw3OtAcPsMVXkTg/c/kghg6ANQ
EfXaVx7iZ0lXiA+f3Diy+7pGCG66lscctApGOywTedykC5vv+oHpZpJ6wRBd
VSz6FXphSyaEP60oUXpoSIuy8q7FOzJvUIg0BG9MLKFkfPI6VO1PPU3doifb
8Q1KLMur0dY67cJ0yxEpvCOYmQB24XVR4hnM91t7W1TQ6/gMrkiiAxtU0/ly
jPNmfUji3LekRwegvPgJ5OsPG43Cj/dJ8cfCcZl+KN5usY5YPJd15w/jTWa4
XXvpm04ekFCWShBG9SPOPKMkjfJnlqmHFki53EC/n2vNj0DCKu+SawSav9nz
AWOOQrwNPraSJzc8nVy95qb6NgHHhONyzOKUaiomSAYNH6OXPJH0pl4D2T42
JDttIzdLMsPjt3QBfj7z7kEplK4Y65oJZpjdDpA7ErZfMjdTA4yIZSLHwI3m
+rCBgYetSOkZ9JfBIvzOSKX22Qhe9oyVo63SAeHXGB35DNYsAg1PjQS/Dxd0
BgOt27LR/9jSV3opgjwhOsYtcElWLz9TFg957NupYvQrbtQOAUtmph7Fs9m1
cY8VBFIDBndjinXOt999l0hdNg9yE/1XYXLECmjLa4vXepmg4McRpoSdnf7g
Xjf3+fTadoKJlxRdjtmarNlL3ubTP6BQz9kgTK1GUu5IkP3X7UblngYqtsja
P9u22G/o7ewO0HoUIWs/agEyqkXQbx3dgggmfMZkX1pUBstS2O9D6IwFHoBV
qS80WhuHGLTd9DB1RQr/WX4875SDP2uH6d3eB+322U0y1pMzkQtEzue2VHNF
DGY4g8MS05XK2jV3jzjjzxNzhReV0Qy1HJ8cJ0tHzRl/2ecdfBctM0J9LjT6
Q6dfA3Py+rtsuBZNppnzhzS4dmEUhW2/B+Vk0scbHHm+t6ZRMl+qFkmEA7WR
hoSSg1QeqYclu7XRHFdOKKOa9X5zlpRsejipbYZ/AOVW2dECCGm2t0eiPunM
GOpu+Boh2YrXscDwDXCD7405Cjv8xpoqCFnfezwP2ojFV3d40FoN4EirjsHD
Qx5KpEg3rTOVgSrE63DKRumjo47OgrUFDcZavziLBWkSl5nMgV+w+P5jVo2v
gWNJH1jJszI3z/PU3G2AKUFTRsIeuOXHg2c+9Ho4gGVlxmqOrSAbyC0zyck8
caDSjggNr6z7zsfxmyTWJ3haRfNTWW1AJWlh0wRPLYmMKaiAEwg6+9dFZgTg
F5fTNn6XVGPtJ/P0NqfpNel/r/zjeJMCeWf+ulIFlQpobgNB7RFuDSFR+zCm
j44Ww1iNMiLsxoAUofRhXFb7rBYXs7utW2dNV9rP9i8zp25vIcQcwc7VOuTK
RWj2i95a/A11CakCdIrz9pf7hEhUro5z/TKZcLTtigP3gBfbfzd1kDygb2yq
ENBnbJ7i5+cQXHGv61X1G0nraKXb+N+osQpCNIbrob8qnvWqpVR0EVvUaNjk
rOmvZxcmqkx1x5AWRpgERG45o+hbtrFdP1nkwSTTsSZsyegqWx7EdLcWcslY
ldnTmHH9HcKLFX60mQjvHvTcf/zgpL/UM/+h5IFx7267Su17S9swVNZxzYUI
JsuyG4WBGAvfP5tF/n5ee9kbnTmGiBziIbdmT4RtR1ZRQBT3xZFTUgF55k53
qGXEpHiCQmpLj3ouMDiAxZ2oAW4hHs5vMe2s72z/zFe0091Lk1LClGF1T0a2
j1lZkKXBzk2uo8lqYJJbfZ+mOa2/Few78OhcM/nLmKauafl5TRr4nrmZJc44
s2VirngocDZvSB6nN68T1VT96G/IOpjgXLTEfqOojaJQepcrIa+evfLSd44B
LUS6H2NfaaUljz3rqD/vH4jUTVyFTOGXQsxmi7kfeaVp5rkeBMYdaM5plONg
sdaI5x6yG9zn0mfYGC56We/bropUt+FchTM7AoZnCimnOTSgw9lPNws9QtHC
162R2y4pfE+RAg0cPk/aPQh1cyXAZD4MqGU6tiv5kN+OX0MUazo4pjmVzG9V
/MkW4gjAA8EN3Mt9k8Qe3CZOohuCbVt7ppFGVpwO3sBwkelizUxOuvOuesyZ
L7xEF34mGT3li8a8V+X76s0U5UiGfcLFrlRGZaZVMLLYYohmaV+2GIbZgzf0
iah07c+/gD8mdv4gUIp9q0dAZfBkjnlcyrIXBW/ofe9+TRcjnEB8sUfk1TYN
e0Gg+bHlv6AApOwkU5QW9nGYkJCvRd5uHhZPqgA0gY93gbOipMT+uxBhT3lO
RiRNq+wPnswsol1Mq5R7gwAzTOZNQfDb9Ed3S7YKbuSFC64cT4LB1TaRU5Cg
M+S3WBhaY3BsYEOwnk8NLfsBlEOiAlLcTjsPLIILD8YLJfVnE8xbeAJELVxt
MGntvvbjottG+zKcqAKeMqEKIo0UWXR2vXxFm6XXlLCJoKmXQmuKJG50ot7n
mTNMXiQSz71Q4Bu+lXT74Uo/5F7jOsVyh3Syy1wzYp0gLSj26D3/UYbq+wh4
m1IWtaose5zSTbqPoFmZZ1gk9QxlKY97CgbN+5hNZWfIz9q4BxSKgEp+r+gf
6NDk8nGvbsC2VCGw+wW0VPKvj4eScJn2XLt+qvyk9V7G83igL4ZEtqOe7im3
bPkj3J1ewd9FKFkEzN9bcNrJvBj/yDvADjAyOJvcrhuaV0U/TSV8AbSnq3bR
q3D3RGwOM6lp4KgezLW7T2bRpszr269Ao2ZISacXb8d45F1im34R2CB/kNVg
VNVrYS44WYwmXmKOghQ55tAvBl/wQQ9b3zi51b7id9F4cb9gBg+Ba1t1rcrO
Vf95aBCb6x9cu7Yk1jtcSNVnJNiCrPbzwblL8p8JHh+ouZ946ADNRGN/lKXr
NiaxXKTkEoc7iddPUKbdbKZlylkH3qQDjzts/AlnQd1dfKIcZF3upRhWQjHj
NehtFjGt1Rh1gONyhG/qS9aOKg3T+wddKkvTOBXl0/LJBYBp/pfdjtXixiDL
N+zEP+zlItiD+XsXmJRVxqklqHSTQcWJ2ncQFv+jitIHYHUXzQQ7UEKSFxOM
UFlBRsIHhIRppROAD4EgqKXt87E7LvUexHKnUPUPeTFih/lq0lVHVi/cmhSc
Wx3ZVz9m4inJvDrj0gClJrPpMvanMuDbtzlQehBYkj5kkbBxXMawQlftxJJd
2ms8CIDe9lgHAVyIUzkNRqt5uEcxPozqNQ+3A8/+GiJh5u921ThYhd5FNj/h
UuRUfkJkEsB08NtW1oLVkWv45bJcdwq3L8YFSK28FMHQZ/vp31bw0z4cm0jI
1Fl8eYLc+LdIWj3Nj0jgTXG3KZ+KUpOaH/bemTM0d51Gb1i/L17xelEfCiVU
w+I1hR6rzMfI9YPoNFFtY/sMAcUNB2Vjhhv5wGyeXKGEYNnbvqfrjVFqCIR5
8ypJ8TzpDUkAWMVkXwpqANs/Ydjenry6EN8NzqZ5g/5qAYCl0mFmcKUQSAMt
rNcwIVzX4mFlRX2v9THG9o5fnfDX0geJzxu2+GBbSnaBQyXkRYW/9N9ueWpJ
PeauEj+zQJfQl8T8k2rJ9A7acEZQUXXx9qZVy02dKke/7CdDVr2LHN6WvKgy
37jebzr5DBUvUwi/cMDwYgKcFHwWoSUvpFQPz3tOA/xoKkFEYCeOgYZO1SRb
d9oAtE2qlaB9sC/NJv0WSCCpSj0VMHyKRz6ShlfsmtExwx4iuYIEfQZcL9Gx
hBlFPN43NMwr0fCAiwOAn1G7hraKeEePNwDae1qbHSwRuGmV23M5cVflBYJm
SRrzz8N63xxO2B9fQ+G38VxXatIZkLMgaP+ubtVkVuFFS3U3CUQv9pmbTfF9
1fPnajvmGCwSaV8rCQc0O2dDdkO9rsDsdelFOEEkBNisWj3VWfLIscQzCitv
4yyQNl2lW8MdVufPHnTcXEYg5Syrjl3CxJp4Y26MvPuPRbBbMFJ2EbKUoPzU
TAB5niMR8h5rTEcNKiexOmVyviUzEk3ud9mJAfKrqPvLiHP0ae1f/6IiUylX
rhAWYWVrWsSp/R2mlp3DhcjC2KaAal32KGIIIikqmA89f86IMlWkbIzgIcYM
p4R4/K7zKZNRMNM9cC36hRYJKg5HzuTiRDvsZhEaEiC5PVa8YJAhuJnAuka/
79D/GvpBD0YALfRPFvSZqoBuHA7M/uuXHCkfobs33cACGc2nWIl9MsfDN2Ij
y80iTedi9RYVcmaFKZGGKBBc0utixt/Z5UX5f2T5pak6WSIPaUHvVBrZJL3Q
L/K3z5v4K3XdLukMlwx02WL0sbUTV/CNpiCMMXkjjiSg4LjchxruLFErgkgD
R4V0shAcF55Cvwlh+D1uZP8EIqRS7ntge+5SVF99+5kdc+PxxTGZrs2G22XI
rzHEOQGJ3VQq6P8BQ+Mzv2IrV1vi+pQjFWdyLms7r/kqzMtY68UZqRBzMTxT
TEMEFQ4oPeWbqRyN3oIA2Wu51OyK4LQ7XlQajvM09zdGvHRldgOb3Vu32zqO
h0vvFOiFXebBKShmqcSQIFOIzqJyqKibYYbCiUZL00Tnj6nvWzLaiZM2fCQr
BMn1kLbceVX/DvIeQcp1z6eGEKkog4x3POWXDBqVy5mftRvs3SGeIkTZj00m
75LtE6yymJHAbFiUvnCTOC9Wbu/iuC+gim0UyU6WD+9LYe8Gi3oXZEhgmMCY
viqwNKb2YKUtfzVi+lbv+8WREhvWRycvrBu/rn4jgGrCmvMS6vt9iuSblY8t
JkNDjLWVkasyHARd0wIf6FwtE1d5kxjb5/u6whjNhsQfFK0ribKlKSMRRera
RJk6p0gzG7yqiIeD9K8vJBHCsqNYD2kFE0vLv3vIkEpVFkK6iyFXybUln5LB
cfmOCJXSQ067zml6g7N8XbVF1JieRozIgitt0Ssr8nYWUpH7z7cIGVSz/tD0
Wkp5GAW3WBWkNgJla9BLq1fg2DndGBM5e+LrStFZu9Wj/1XyLiqecv3uPfR+
EDqjQdTF/10LroWMlqe8M3bITa86JXHary3t6MTnwDuoEcN6cT0TCRTK37+0
637D4dAmxvflhWSOw0pPSPfMwy7ih3E4DABHcpEDVdONeH2T5KY9U+wbnq39
5PSR67Pcwg+lJntbnLDAv6vHGjuxUBab+bgxhB2Udz9wWu8Wp1tycFdLNpph
clY6G6rFSDEK3QNOIj93sIxOFRmFj/i7uJEW3JtQ9HLlBpFrnvXTJKdhoUgy
vye11KXsS0smoO+Mkb6Q6OJ71EIMuFjVWCozlYBuSTrKavpavN/CFYZHr2lk
W7KEM4Df2jCJjHzZspfpA5tKfzdDdx+XjuP4ocPMCJc7qlM40HKHoOYisQv2
42JnZ7NCiI3H57qlNLp8H9LI4Wdx+Rl6ifoZI/CgYgqdvR5etRbzB4akX9Qw
D9cdbWr+miKV0kpvhCtSPxH28sihmvKMrCNpcfxH8pU/EyypJ2lfE2dfrFe+
GZpmKx2fgoZP4hQ2YuOqgRHi18Qw/TO67W3uRXWmPW8LeQGyt5QT5Z2dTIb0
EXkqKcypROxkiF+lsZjrKaD960XKvCQdkCDhzpzJdvEQb0nC6tQGl2FZreNU
oCtfSnhc6gxtnL/Fo95e7MR9oWtZuRCLkBSmDbkcbMSA3MNqekRqRiPtjEOZ
S0bCxa53EThiYaETqKoqx5wutj7csWRVvxCYYUC9fNnMXCtC9wYK7pkQKJiU
+6Ng2ClHbzPs7HZeo9/FGRk0FaAOsW7P5dSP0gay5nhFd/FmN/yzRhW4Lq4r
K7N0o3ADW36oWaCevOMRJO2bRXyigwl02hEVIs4mvWayU59NdaAWLfnM/FSK
+EsgmTtPJmyZ8sbZnrWOU2kTgWfKQD0/vGEKx4NFmnXqXhG1edyDUqguy9mw
z89HihJi4TIEU3S+6yPFsGJmoG4WWEDR93nV0+Z00qkg906zaZzXRjQmYGMs
wgoomGRBBSTty1WCjll/ZvIPlKuSSJs3Ro5+CfahAR0pTlln7q+0wz63wgWG
oCVsM9porL16q5l6uKog8EEEjnbnqj/RtB7cP/vRU5rhJ/uSLQVirOUWoQ6S
JH7Cc5tnY8wMGZOlyH51Z+J+TyPatzmqSD54HxD10CueLG+Vvd8VANpdopoo
rjoD4lWPkWvbnaewgIjDW2EbixMQzbKfEV4MY9QBRsChzYtgWMj72km1K17X
JxgpqLS31ulwKRy06kaYv5bMuQfXlEDMRbIL5PkApiypWN1b9wYSu5uNI6oK
HTjB2xr86yVQJNvhABv46+ZjpWQxLgiL1LLwOVGLPbtw8993RQ1U0o1ssXA4
U/ZImf8v5QCyz2LfloFN55bdHvKUs0EOfwNMULRYFpA+qWlW1iom5IDXasDS
uciobWfXuRC3AdMnPBFDG3XFGSsSex4JpzVBWx9zRyEwWh+JMiURxobDKYKe
wol3SaqiOjoOXMPE7PeeSiAOXIIIZOsevqnoEIjygjWafTRoS+GoF7Ry/zSc
dLI2rtnYhM0Fh4be6fJ3m3nwlMwuzW8bvG37OHQPnif1TnHIV5Yu6JOV4XFm
RIsCtc37SKd06KeV3JxcDF4iKU7yZW4XiAjLTIohw0CVUmYc5TdJ28WPI9Ko
nrsGZsdKguPoGlqaIWXj1xN5K+qn5lPs5O1nqdidMDz41iLL6p6ibU/YobIO
GNUlIf4PGKhXf1s5zvHFhPprx05rj7KhEWfF+AE3kIhehSgqAqpAqSKirYsu
TArrsxgPIpFR+/fouBQjgoW8f4lyE8C9PDkSI6t0HtspzNl+4De6f52VdEjm
alz4VNxX6pnLSnadHsMj3FuudKGvjHMZPI+T35+aYqBkQCJf3TEH6nTbbEHm
4dmToQvicfsBmahDKuV2G6NPNBrBCy2vsKwKlOyV41oDgjXhAN4G84H3hdQa
HFo7QG4MwK0zBeLf5PZLZZN69WUlg25PlYshbjSKUosSdIn6oufjsOUsU6O6
kBUz7DtlhbBe/DiXs044DW9NE3lCuv3pfrzBEqKLx6kzmCRZRH0b2Mzw5Eaf
QhIAVG3Yq7UXY03tzxrBAON7Gm3Lbb/8NONFZKFDmT8q12Is/m63eJ76Ua9f
ugc4CohHSezpj94MVPjHPHETkstyL5gzx5XAHBcNO2rVNqJluHLIX96yqWuX
3gurCxlgw7vQI3mCa/q6UssLH9Q1CJeIHTKgD3LzTgyxgDTHv9SXfGFsCjvL
x08Yy1ITdNu5RSlOSl55u0aLwHJK0PJrc09FxwmqZdkE2coQ4fwdHxBAFPgq
3Tnd979fGR/NNB+fGt3SjxFPftdprmvfe8mgdeW/iMQYQTXHcMGi8ex1XQV8
XPjBsdeBGnZBZPtECXnwgF9SOZ4LS+FMRi4z5/Jj+P1NrAttPjsU/79BZuX4
TaOWQHGurNQGTekTjGONtGKRfGRt9DtekjIHJYa7KcyQFYIbYAhr5Yufv8OC
Z7pPtGei9sLxvsAYcEk4iax5rb4bxibKXc0oKGCJN+zjqILIRI/In+BxQXON
pU1OxWWvcw8O3dzKmrDW2eTJpuY7lPC8ySg6uHSekYuyX6sSP/vTTFmppfnw
63wumVIfbKmT4w8lWJMILkgDKtr8SIkui9AV8gFWX0iDEYzPq6cXM2hEldrH
n9avYbW9pnEyYQazsuObDwyhOPyXXFtHiO9EQ25qjbu6qPvf6WzD6GXR/mLD
ohw0UXcwpI7crSthK9g68kYuJf+SJgNH3/cliJ7sPJ8E1A4YM3LJqlMh3fYk
PykGAnWatfaE71YbR6+a2nY3zXqAiZ+1LXbXExmaiob3FEmCanxiLV3+a/A6
nrnSda6rS4uurpOBvTmJX8LPKQV6mTJoJXV1ufUg3/bsJRwTFijUvSjEeuwM
eDO+DvL9j9uPfjWdE4rQ2zTczFj5deKFS0uY+Kqwd3QMUvwd8D9SeI5/HxxM
VxIMsE8XaFLeWUsRjBHRK8HUuBpeo/MaSnNg5HzVS3M2dYq1BaSImmb/cDly
ptrd+XPV+MOBYcb5GLboQYNuApvzN7P2l9fDpOjsUa/cNWOADxCwAXMvHx8/
ORqZdqdH3oYhEhFCtn9yHugKi0qiRnceVk3gkhDL1l8UAyIGcWDxdtE1B/pb
XKAinhRkHZ3ZbqH/kJxd4HKLC3sYSb4ukqD5zD8vlEEPV7k70SaVyeT380xE
pmnyXApQB+89+8zRyEN0pYRpRtCc164lhlDV4MtyXVbDNj6aB4eF1ex2t3hM
hlHl4FWn14A6rqxOktjothGG94YuT3gIntQSUpmAco+i3xCIfAKdFWyquKnX
Gzw8ae27Gx7jAypCeXtXCLmRsN6Snc8aOhiYdKfGa4vw/+2dQROUw4wNgZtA
4+X1/Pkisqg3bdsMpkRZgQpK665fL0Ez14H14iML0lalQdnlYZqkETnWkaFG
lETfLvGV4w5gD9aA+9KhveOE8ALJPqRNhJb4+PsKagC6TjZS1rvls8sZdnFb
TKZ12Q9QpIWhnjWzJKAnYvnRiqlf32KUB8JsloZPph1WXy47gnkjjcdwJ1In
sImb/LrA0foAA6+wbAcd3IcxpEHowE8miBBfCkjQ14nPcphmmYruHgZjoAnP
Xzx3c3QyFNfuu0bY+tqbYEW0WC72C4FgSFLSWXbBqO7sjkVtMcl6oY8ZPqM2
m8Ycbg6v6EsxlkaOa9vaseGg8sZwmAhbiS3OKNVtiBv3j8Bs3VDsHTxKpf/K
4uE+eGmXrRptfqhfmfNDNNWvyzRCPMDwrHs63WouXhySVpLuvM6+EStejz+u
Fv/amzOJjEYkDzcfZlj2Zlds0quXbcTwSaPkuQkETr7bSgE3AABZCsmJUm/S
lssCgUVs/QwlnqoFpE/531kUcTx9on2Xvxx1R26/oxSd4slO5/oT4R9+0mxh
S1tMhggJLSfjxmOUOcrDEBySiXjJsuhexEiwPgdYQQ80GDSES6p/M7daAzIm
3JrnxTm/RWICM6IRL9aw6Q3BQfI0SWRKTAktrQluA1t+LrZgE2tg9QIPRxrM
YXH5yyh9rsr/DHP0oYE2xvGJ+Li2A0Bnf8jfGcUu4IUd2n3O62m0iTQzZNaS
mrxoX1tqnehRI1pbAqgiYSC8gRC2qsYnaNhCIO4J6Kf6W09Y1Nx6B4uAUGs0
W2VVhCSpDzRuJFsCzsGBvUJ4Sq0gi++xEQ445KU/lSdSQ4rMTpnPlbrUXeCH
ZxPAX9VmlG1QGAxgoSCQHI8y2HNOEWCFZYoXpWtMZf3Q1DcASrZLc0oVQ+KV
PfyDCMs9LybmXHSSiQiqsCfRiy7UNSUQRAJXCvPAeDWiYQ7wKu2q/K4ox1u7
hygnGTuu8iFcCWWoWsA+88mWbOcMns32oGoHdg1Dg/wvScrx+lS0bBCigY8g
CdJ4vi9xmZMxe1GhsA5wp28ffgvhKLRLpCLaUNtdlsZfs1S4E46+pYt5VG7K
cmiP9Dd9JKUaAgBy3erKSGqXNkSqz3pLu4VziUR1c2FXwyT41kLsFiW8QwD+
kbb7nCdzrvTII6vYBJQ3LebnzKcpAtX4HEEZskMOeYuOwveEoVH4dTAnk/Ll
BAXKWDO+oTAnkeQTXy/qATbceF44I8+Em3Ugv2l2tVjQNJgDABV3o6yOwCdS
/FkQ1PJ2Z7Tl9vJCoBju03Eifpj4BdU6iFx9RhyXLZ3W4fyKZSM27zK0Kcd/
+CQPM1gNB/NK4o1AZ1uuZ9aCaMSKVAKGBSDVLnD7XQg3NYORPLhUbr5hyZQj
O8P6GhwflcHS/0rbz5Ifp2XsqhXAwSxyTnq3kfneJt/UxZS9yCTpv3j9LpnO
a2Gm0oIPih2qN/fWrnDq2HL2O5+yu6b/fwYJL8xrhV3d7s6JUtQzu3BT11Tp
BnGkqcv/+ZPqW+wQLtfimhnEd0NDHSb6NryBFlR5PZ5fbsn5ru5rAaMYJZYj
Sp2ZXxYYZ8Pcp/nPWqbPD+DsKafWR4/FnXSx3WauAP7TgGeoavlUMGsh84ve
dFkhSANvdpi+nsl8KY3gAeYD4gKGxd2A2//zW7mgklds5o4VQO9VYzLLcPcW
zWt7m9G0yeFrVLUIumjc3TYav97BW60Od9tyvh1er6eu9EovJU96j07eH5wv
s5x3+JgKfoWEo8B6fkbCrmMtH10VBa+l8fkJ7L2/Jk3kNxDzujpn+MUppy1f
GdehmQGGHfhbK8jL5Z6QABZnZraT7KVS/oh+9s9WGsyLMlag40yn1ywIEqYs
ZEpuxFkwFwMdBp6tMSM00TSKfBRLK6k23FwJ4bdOchyWqeRtHluxS3k+47E2
ziQwuZysk0eCK1UK3B8bv09EoowSudNvcdZHxU/TahYWcMCtWLpnABOOfKy0
ABqwiftK1VYaGWhTZ93F8icAMXDYvX1nP2Zo3E3StjJoYA5df0VoP82yKUxf
Hvv5ObTR+oL9lW+q5u8ewwXlu7OJf8YJ5Vq+R5z56TzG6fE3OMqHPCIu8QXS
8vL2L22BqId84y3friBI9/VumJH8ep2xlJs0jrFTt4Cu+0OXUKVODhUv3Sl8
zxtpd+4MJCpiKUyyOxq3qmYsOEteHUqyxiqA725aT1CRyUs/Uy2OFEZqlT2u
8wkKlWXjjz5u3VFoVJbDO621jhPo8YAq/2IGyBFTErC9or2vRz7+zblsrINl
STaRe4xdmnq0TesQ3mHrgxgz5xV7vfOAacf+aQx7o5hWV1tZcB6FYSHvI0UH
0vZSxOyRQZy1Z4BaRJHJhcLgrJ81oroBuVTgN2celYlTKpTtYkruzBdWi/mw
wTeD7GlfXjJjSVn/ktBuO7p3dqwlHmbA4wDrCLWMqyvPnSSSJX2pyv8FmdsK
RbFby0/1yP/3NsHopxsRzizelaNw46aX0uX4a4fOxghV9uT+7hUMOVC4BR4Z
867pCQbGuIXaKMO5WL/KDBkbmYwG1N9FH4fh/sStHW8sIQu20PzVznSYmKaA
8oKI9+j1gDPE+Wu0tI4Ch/TfP47/rDX+YBOAAfd3KHEptCM+t9vR46f2GjM9
ukDX8q30l3Xrh6jFblAovFGC8z+SKMha5pDH3dAu+kRzdEIYDYwxrfU+8d0s
iRWhN176BlFUOIN7Nxk5loEXkDdO24gz5XmTaTJCXF5hQa3GnSTM5IoS+/pl
jYG9W+NMaBOJJmiWPptf7kEiqdeFJPkbG1k0uaBl2PVlGO2wi7uxLh8Y9cWg
keDVPRAm/FXKLZe6O2msogFScR+tMBXLcTe4VB78gZaOrCMb74jnR6BYy1Ye
HMjjvouGgK16LofzRFd2ITANpW/G7vQRn5t0Bby9mdjx3juPrgy3RojViij0
csOxBjDHN1ZDx9udzzi6k6yiOJZrrNfnHeC737sucKDZSfgvI8fYsoYYA6O+
QjK8zAcp0Yj0PTV7mJqZBhBLtCKgWIVNwi/st61JY59eLNrJHC8tunnwiG+H
Uyk6EoBMvpDbh25nPq6GbxbVcZVCVubm066IjBlQ6IMAM6pn5laYktIzSERA
pjBxbRciH+F+BJt44lkLHlxJgm3LRkXmOKaP7DjpjQaYo45XTPUemHdoWdLe
mtUQCTig73KNsu6S6Rhhd/rkrxw0Y0SZGJBC6svaMgjJn9Y68W3L3cehh77v
8yS84SgBK/BefsMiwB8+KhBV+IO8QWuVQ8B7Dcp4rni+zv873wYv96bZc2+4
ejPLVkY8vXmd/UTd1eUfFHnVr8AGO3eQJYgSURITJmgim1poLEvA1BG6vTed
pFi/cm49yzTh33Iv5yZmV6ew1vGris+02A1R0PMDysndZVvaFvNIynI1hpYF
KxYFGinIT0jHxdMyEvJ57tTowNzLX1ZIRGdDwIUjGuKCeGAJ8bZoxkBXYarF
mvpqMlN0FxoeXjGn3eB9iHfPxHrW4z1omXoil0Nz/RvSK8gH+OZxiY2gyiKa
iNp1FtzNrDJ2G56qKORM6lGz5/JpPhk4OIl5VVGPxbXXgzQnv6IFqivl/m9l
MW63kH5XN0JN95b7Jr3BHxGz5mkbb7WSHKAn21gVjGWHOFxIg0CIo5ekuyhN
S3l/uNPYlJhGas2qFJUlr7V1UhhOrRq80QmZKxRcSYFvVLkSHP4E2EtL4sap
HOLUTLObfK1gW1fGQUnn6mDs1e6CWZGOl7+G2oFDucqplIIvhFg5h9ygIA6h
MCOE6WUInHDMfUktOXoYcEaMwvucJQlOCWRb+67yiEgb4IGXzdm/Yy3s8pLg
+cpXn/+SgpY7M5O64nBc/kRx8CsyAB4nA6o3UiVD6XrYDcYTZEz8FPrU/Ftn
iYc98IRlIG6nTYMKWaAA+L75dvLrX7SPbUUXCTyDx9fSUiKjAhUnskuLEZZC
hk/koQzq0KHED/ynUqWIUiC3aRISTCDUmUkYWZVF1ervAWCIb1v2rf2g7Vu9
2KHVZ9w/VkJWkTp1TCq8H8m1E11tH4WsPppq9bzAjUnp1XBzVx/BEOEw+oON
ZUjeaLYiBP94o9Cjx9NAlJy3rlwwt/TkpQ30qiouqTzMD0nDFPEYQJavze1S
gFCvCXv8rne74rnBDX51Hirv13yY9O/tPvwAVhX/7tuGvZ3uObV3Um9O6Q5f
tA+BnKkPHiXV/6sK+jwEk97UIyOz8/pGFAnN1JokIueQyVO2uEN28k7W/DS2
w8gcnxvN/C40DVHyA5rGmNR9poP2MjA0c5G939/W2gPf3PGmu1la0rcftn/g
sDX2W5jW0HB8L5dS5ikEr9Ur8R9+CMVhpUQXWQaYvBuS95oxR0UXULO83PxS
8iYh4cSfrURg3ZbHxAAaCf9exmTCJ8of7fvebB6SanWUErUpt0vWvZV0vrW3
im3KIN9Q/87WkkySyOFqfeIYpD9Gq09xNIjNEf3Pj+8PtTJjgYSloMbCLnfM
iALmt63H5wIWmaalNClsD60+2kuTxjGHLgxhd+YUzJpqPx6oxl8J8/bWSxsz
0XhYwhyAmjwIXANoRBM6Q1PvZzAzQUOcMWkqnWIhUV/JUzNV6stne/jOJzES
6X5a4aOreOP/eoRkVVr86G2sXUDdDfOBYTOoHC41Q/8+R6eVYeP5mtOMXU8o
hv8KSqjzeeZ/7DfNGWJdY6AUiv9oqeuoGJ/o/5bXPrV/x8Qjz6dNNhrGbyGN
jE9MzssypMP1F3uWVJZT7Drk4MzFlXEQyu9SCg4uVT5cLSHbqjFDLSRcMq/5
kwomJL48TZfuCHgCBPsOlxlM2adiF74fZQJ8U4tpINO/KKUH45akwWXJN4Ph
Aj7RBSk+uufRmsfmUelAkbTDoHylCEIUu+wofTKX5dmwaR0bjTtInza3L4aq
q//plxKZt7yMLZm/RtOpp6ERNnWP8scWHU7O2+9PCXupVLXbfP5MIHA8tzoG
EkHS/YFllwthIFyLS4PCQqFuTv4oKeybT5GlCZvF8TAjZoG44Vuosj3M2A+d
gO9A2kxTAAHfCbvjNRlfmKAa5PtwvLBHy3CICrQ/PZHawmwsDi6rx6vKN0KA
wTS1gvY+3chHZnK14P5qmr+nCGL++pZ+XbGmSL5P2jv4ImIH9dXw34A48CMN
YMbhJc+hf4Ej8iqm4ORxZShmLJNIX838RPR59aXD9m71YB6ouY572bMD2Gtd
iCSt5xjRdasfx0Bwvc73roRDW0BZ2OKWRXBHbLCSiijXLFJCjL8RQt7cz7pS
mEyJcx8fKRS3dWyCqypK6QsHSoi61gB5NktMcyWfGfPa/a8fB2xhGpshcnm5
77YaFBWzq29rmpYPGlj8XL4GX813W7MDJP+85aIJezLWzRXQytHm6praRPWH
KDwSUz5tv6lpFrhwcNVEfUgKfPjwYKICFXqEKjqTf3Aqce7yVXVl5mgTQm2P
SJ04XyrLhW4epmCw4osvbA3EvOl59rBghw+ZNcxb771RJGiWH5vjq8cG/Xj0
nwL696/qKQDQ53N5JxiOid66hTexRKoSVq8ce4sCMdXBxW2yo411Oja6UJB9
GpODc8g25oYXzuTxzkDrRqIapgoJvMXxjwo6pcfOu3G5ejEZk6ssbsdyem3w
Vlimeb/XrcztTKaEFafNXS/GLSCCPiFXnUu9gChCSN0+536fn7l8rNa6JFaQ
cWMje2pIKWAGuWyDh1oCPCRuW8LaDtheqCo4X919xrbfY0M+yA0Wyjy8Y8Ke
YRN+JBpmU9VqaFte/QlNt74cnDu0XnaLat08bMfBq4/+tcmKTIh8xSNHoofK
oiN0QBKsxVwMrsLKHSC/F/jDiBT0PkCMZxT3MEk5O6lvFRMBixvDNDdVak2T
iMXVv0yaOdMD2u1gozBEYo4Ex8rIoaY2i95gJJcoru2zmu8xpu1H12zVeE1E
PC5LSLgq+5xTbb0j/Dp+JmJ5ZCEEL2uuBs3IQRpAzRSceglRJFlPP1sxiQY6
bh9iW9ayAuiwKx555k/Rv0dG7Zb2Kj8ZFK22/kQcQ4XjHmCHht21YLwou7+L
XAlRE4V5FMzGRb/BLheXuK9brOKmX0fsNtNszjCjwTGNJnpBVrFInoNRzyNn
3YZA06SF06wjx+SShCx5711k49EagSy4ClL0ikSLY2DpoC9SCsvVRYkcDGHu
lxKv2VVJSq0cS89PXjG/4B0h65wAwR2GdH5KL9b7UEF7pWuY3v48jDPOasEP
qdrKrEYjqch1BEFEV0WvEKTPqBjNDJvKVAS/He92pmMB75WQxdu8ngKDPhdM
1x4U666YOoVngyVR8Cusl3FQYqzl8pvXxDBYPp7WbhY6PXod4IOuojYYMtcV
1BruodzXaJNGEmzXRNyrDjFsq516CAA5lOaGyCOPWuOl+eCllMv79Gz6O02C
szXr5NiDV7Wws8Sb5DMm7ahC48s4CupSKBh90FA9L70Hn2Vw/mjqctUQbTs2
iSIcP5iIwt3xwAk9xcAkw3tjAlNmGTxD5MqJb89N1w/25Ib6eBaILCewMj1H
kbcJd5QO6UnjpnA75SrHtoARyNfAUqxyL/rDXV0/1KcgaMgeAOUE92UraaBB
/99Y4f7WVE1fsGQNiO8E4ibtAWQQ+WN4hkHsB0CFi1auZguFvLYat+VjjqFk
WnudblEvCbKDZxmqmXb2rwH9arOj256y0Fu9O92hTyQH0daS6nEnR1hmYVbm
nlWYyhzBcmeAR2gDbhpUBONUMsmBK4wwqD2KWpHPQfe5qqJAgUiVKaZ6RfIf
DDn7MK1O1RIQem6nyotqbxyAaZ/LdH4yw6CYlZgX4w78xQelznfWCEJtsTfD
O/0wxbtjj5Hv9YiFAHgw5lThsqnAmmdNCclbtLY0eg0SoQ+clB8NHBSDVGqS
ICXx5ZxGTpz09KF/zdu6xCiCPiFV0DUV82cSbwx05lY5LTCbbQ7dBZeKp7GC
rQOXa/DXI47Me4qE7fWIDW2CSWp7X9irSfite43zP6iHkSP6Pj2fWKupV817
YWPcZZuYCfgo0Xd0kvBZj+tzzPDWeZyphTOMHBdhg1Qs8GL59O271GPfoZJE
qJ/K/VEpz6I2XT4qMvmnPUUAiiKtOMeCXWYzduql7utQYeipid+Qz3fZD+jL
Zfo23Ll4xWXvI/fX5srzQ9JiiI/sev+R8KdNruIt24P70dZrULpZ/AZXDB0m
9uxcXlvs0/R1jjt/JFNRLigjc71pmRUOudaxTQBgHd1i5tGY/KiM8o7UPptb
uOxmroa+WcJOJ9esbJhqC2RoJFSqLydGGBUV0YLfTiz8Hqm3lzM9jIGq0oVr
aML9UE5IyXfL4Tuv8+UpehnbP3WigeCAJUQDacUUVVKkVrv51QOtxp57G5EA
Nbn5JhBtDLkLgy2GDGoe9821TXpEsq7wqnn75ULEsIEUy81faK3ZvOqb6I8a
9jfhGWf6X8JxTitFK+JEITSZ44KTe9CMRR6EroaG8W2JybMdgs8bY/BeLM1B
GnuNQSZCshIvBqkpYdsaFpZK/cNxUoKJhNOPEmSK/o+JLiYmnNPLwX+cWAiF
RSVUtWEoBosF8XEyVUVI7ZUaSG5opIG5AxSQ5r3yBx8wr1MYhlrFeHzub0Nx
KSWMdvj0FzCR231HvodK+nCveJjmYqpM/4gNID2HHkYTbFzzayYprg5LjTj9
0EL29pVtvYH1UmyqsruLt8+VVFBVlQe7mqoJV0pihnR/VFFRqZDzGIE8AZyi
DcgPdOMyN6uT+KaKRoEgTjWIDAaxBIJx15fFZCQZqAMGI6PTd4IQTO7yjkOA
xtP2g/MuE0cJlfL2mvPODeuhyyhGxdmc94Nh/IjU3oyGQtFBlcDPN/iOgnPx
SmmXG6bwgiN7DLtK2mg4uG+FJfmP3NAcuhnewHmCDpnUZqexJlXGsLw2aBxO
qgDysPutRu58SHOu5JSPgC7i+AVnXZUdWgJdqc9R3NF32dn5BCxnguEVb4Wg
GTBIZVjkdNHe5ia9ZreXIivWIh4Dk74njW4gpWWUbc0H2/ppElkrLPhMz+4r
HdvuJvy9ybM6gRSkcEgzDfzzIiCdBtGG5eb213RLABq2X8WaVH6q4vLaGaKU
Tk5yVhR6npkT1FjohssbG+vMYMuSOUahhheazyaB6r1o/hUy8Euu7sXrjtLL
5mlie0H6uGZNLMENev4nBU8XGTUYtNRApcpeREO0APfu/Rmk5PdjlYwUkV4a
fLv9oSchjSFrvuw3kJ9sSIuUDIan+jpG3HKNJZ0e5mMZrzUt48QHIVlLRs1n
0MKU7fosbMigJEALau/oX96JqvZxYJqekmvVHGXZYCi4GdINJ0+ByWyiK4vF
H2U9ry+jHP0Gp3X/hrF5yijqKpLeM2xwgYpSUqKvjuZ2/nmgNET5Muh8fCkc
kzd68bwaTxW0UjFazo1NmDN4eKBrGlpTsTNMV5ZozSbO3hqo/0XQitc7+J+A
4m5dlB+J/4aJKgGtoaTbe7MqtG/9ON7XonNYmcQGZ/G7A3CUjjbsR7RSemgu
IVf4L9PKKUFxvOw6kiKxpAYh7PT4/FQqfyzd34TJfxwMSqdyrPtQ6b9E5/uh
fJLMcieFxEl6uPF59JKy13aenIvgMYKk4Zr+sRAIks0aBIGjqBJ126RiipJK
TTESYxtDrkzH4C0KHuVEzZ1vCFBJ/Ybxffvd32Uto6RkopQmu9lbXf5S6h5H
0WKgJyjOqoDKCXCXvtKSmvtbGzxvTu2UNoqpS0CWbxv9sG+GxlL84s4Ds4Di
dC5ErmUqyxrj/tdD1gG34eZMny/8Fk0F83HaZuY+xkUeGuwRisyramG0Th8Z
E/fU4plSFdla4LREtN2W4m1XeMCFHceCVppF1BglOk2HYVmS8vrHlL4DgJKa
eFNzGjGUBAyZKfWycUuI4bjnjAQP6M9ENnby2xzQGkuPdIn/ss5j8nGlw+bY
grdFpkIYNZ2csw6oaRZY6ci2MSxcyDqRrnk5Dsio8/x3u/P4X23L5G8VLH1v
4F7i8aM1z8uZWJnlpSaYmCg3wNnYEpaTTRMwGgDr1gSybzcsa48qZw6VcBNW
LjhgruCGCsRrwo5fykqCfwcit/Xrz01Ig6nKC6pCHdXJkrBgq/6DD4r33v8O
dDlRWPeBjq5gJXNuVrDdr6+OWxPB7E4119nL0+csshoVBZkXmgo+Ww9ezyls
250VJST19i8LBsvY74iCl4ONhR0cwiSqbi74KyZHHI5upSS1Ppj0Mdwypz9M
naPAYVECjCmeW91Hy4llKwBi5OowqzPvR8SGrMlUTjko2HdXEBIiwTEDDvgr
gzoenDD9kIIi8VGJmMJV3PWLcD7ZoM7KJCfjy1RTwlCXBOycFF+04ofmSDML
otI+b1r38N2TOYtF467MHTiWkY4eDj9E7Cizw+JfECrQQoGzxPMes+WqGKBG
h46PpOSyVjF0mkNzmR0PsBjdGSh3BYfHnao9Kbbw/TJne85xUTqBnMuXABtm
c7DtRBasq8iWEEnqKWLxvh06AzZdmdmoGnaJrYBjAZwtkLcJtYXRTYE4ghJl
sraAysUco4qy6Et/jKmsVLkrhFZQ7rgDhGFuzbDwlkNsh8SYYSajQ1fcg3WT
fnVrB7toDXrirVcue6SVWRtRQp1Qlj1gBeiqA11n2wiAD+r/y0/9I5iARU8f
Hs8iftnmbS315rCOKla8qkCXU8XMVuPUGztMRdxnNiec9aXBFdqoPb04NOPG
AB3T9qMvw/nIy2NyObBTdB1yCsX+CbK1/U2Xi+QXum5rM/KYlmtqjO2iEZmV
RlgSusZM1UDtQEICSQiS9wN7fP7midnwnU99kGI2XIu3mGQBcuDnrCkQ4ycR
l3BhvuI+hJgRfvPvWbdLNTxN3H8+fkCO+RbV1FHknPZPXPxUmwWazfJS/eED
eNPmN9n0WjpCDnj/swo36oqgoxayJ5yb8Pg9LNxWnDZIkWfe+koIQLttK+YA
jSTl4UXt5HRKmE8wWXtNGWlSg0P3f3MEs2CKQdbdiPKZRekN/hK6SS1Mc6EG
o/XadBLf1AU0NuHwfLCS99vFYrirGQx4M9C0rSr9Afi0gSJV8K0rIfMMCscf
wEqahCEbT4nXPTjDtvAL2D9bh/qPoY4Z5FNo7f+zDke3II2MAy2KEd59XWUP
qiDddrh4wCf63zB5aM3FNcnvzpO8Xe/pTReloDLNeilZMClVK8KHWxkEUS8R
OxH1NtfidEWLIWhd6hEij9fbbqTmJeXszb+8VW+QWxBAF1hz/fGqQdvvEI9E
BkOwlKYOofmVKuympRtGZXT3QFkAtq0ANDUoNYjPASNaldTOanCAea6TjJjz
ZObBmBP3ljMUHTjCQD4OeAbw8Cltg/sEmcAG1ZQxYx4+XVeMmXbI+2VsE2U5
0WgBP5pLZyauuIGG9gf/YyaHWsnGVr3l1jVE70yCotIh2I89h+klulXnLQ4p
1RSDlFUhIRmeo3lwlpwcKbvFMp6nt/GFX64N3nq/uOCrrkFoVJE5Ip6sIDkC
sHj0+3ucb+LWPL9kFRxQEqM4Q77oPbHPULxbmvSj+CPMHmVd/RDisevj83bM
g7yv29Vv99TpGcWHGRwkJGQzOEGWiGrkGJNqYDS2clB+gr+QobSzEKeZo9KA
G5sE4CC3PmIMVNvjDDzK12vITYmFLHK8RZHmbBWB4nZvM3clgeA0gLD8ie+N
k0ktu+/L4iUe1EnGCnyX08UWIRtNAxGdPlVwqjMjVZkLkZQ6MS3Uo/xJJpMT
7Mh2v6CqSdUTelZcEJXToDA2JayYV8eaEgSGUSmfJTCFKdZ7KPs++Xl3VstJ
7REUGDLzlqdi1IOd1ojYAsPAarMJNYbvTowjTh9Jht6Eexwg2w4ENMp7UBt6
bXWpISY9zb54bPW+LT+l09tTSnH+4M/Sl7r0S/0NuHqpn7Lbv8zES+4+Ey5P
+gcyO7e0v0/68dyaEye5itdFTu36x40bWXVFPhB/ZwhVGkH/jJWHzvzwePmB
zeZkoNodWaahGfC6VUQKyzBfNMpbx4aL/62ZsVf04CQyhYkdRXki8Ua0vRJb
31gFmzn/LW7+cYLB13BWRFeM0IdkSFkavIqJ6APvjsw5KLIqVqU2TKck58sB
pzjZAeRSpq5+zHMP4NU+sWP/P9u5vmJtVuIQwGa8yYF4BSThyAMQCju2JGLJ
8EvRWuK5WUv6JumZlJpSOmGBFNgZfUONYkqzTTwMYlxMOxeHrufYuD5JgZr7
RIbHVYZCcBiVc2SqQEW8QyOB0fKL6FEX3GuOj9cgxLLT07VKfc/4Ffgzec27
e30yI58pBhSgdelPF0IhBHuIeQ1ujDpFVAoguwujzVDBjk/fUq/rHruAx/mW
H0uR0fyqbSxqymkQfJjPwcQ1VFgNyNEEWzQPILxAr3KtPLTeX89Y0miEVhMP
5q8NG1KzG7dJnpBWebH4QhKpIxngjjy9PWarpESZ3VRiO5pPq8lYdXltV8Vd
gBiDgQkaArlqedQv8548OibeqcvEUa6/VzDiDD4InC9i6njPUYjamP1YRm7+
xZyP/MEzPvH45oKCjWu7NUJ4PoyIj7QnWvSbxQYOTFWXNRKaMnSHVhfFHLBl
vbt3ztGsVCmNra/0/n86DlkzODN2kzDsrO2iinyDSP2Au/Z/yVLCfOttxBie
EHjmQIR7yq64r4it29vihdVaJRxA6CDjvypl4ykj1UV5QOdEvlHNntcL5YtI
BBQFaTOeDibLz6WVv2PfyapDOsvKimIV4UcdRN93CA9B4/sKMTX+Up3rzG/+
d0aEcyAxB9gzBaAaWX04zJGw9p+KB2IvHMNAL0RRATbaN0150BSNg8Q/PSlZ
RcBwl65pZqjeTWtRk7f9yhuXhR4aTmomrTyql+0M12eTekga4TpdY9WjweLR
cptKJbn3VTn1XLvnnd034TzgpY7Jd+x4Ae2GbRDCYyCRiE74NHGFOnbw8DSu
RG97kc33jgseyIluWzVL+/gl8izNiCAoyoPANQSmm6/A2o9Lp2rVpqBLBqdO
MVK0eFk9AhbICIccGM9z6S+oicHE/KvvHhmppICYstBzGbs5R8zYRkXPqXLl
C2a4CVWWszEZ4df6wTxUY6fnN5r3llDbH/BDKTkGpoy2jC6bo8b4hcp+xdJp
M1ffwvP7Gexx30tdu9ypfj0oPL1h/ediMfxH/VvzZ1FkEUPXDZBMc0eMJEvn
KSaKVcyT9TYyGmN71sXR98CsF/S/tJ13YxRmUY5AcQOcq0thhkTbxbax45Jo
eZaxvnllSqMAbapwA3wr7CXWVoDoBDEiXPZ/xPKFhVGAN/Sx6KE2woGCLwHD
VFVwl4HTYS0xFJI+e+MQcE7LIQxf1md31ybvRc8sCCH/GrpP7WXKVyI7WuCu
oRorfGW2VXw05hMI9tKFwVy5PnvuvPmyTSf7c4ONDetEi5cWIM66MyQGLHs6
kBDjmjgiPpcO1JaYAbiquxcHHlnrW7qvNCqFF58ai2ESY0bzQdT7H+rbRDUk
AvQhGl+bhr+AuK5vcLxRK+xcWFnFBPYDZsd1UiQ2FRbLa7pgD9CPoDwQLCbE
7a3DoJaSMRYDYcM7iKCNE6KdLlcHRep+zDqdLuY6Q24rZnnslzr4UKcpBl+o
rC0tAdVgcd/obDA5Mbl0ZDGb9mr60zm32RSjxcm2eKHgXrYf5vbfDg1YWsm2
G0hhMyOYyQcL0GEPvqzUK5EwV6oicbXL6peLp4wAvMbFqG837zfEhicCfACK
KeM2/6gBVAn05ia8N11AXTCPliFKP+5b4R2/TGKzag3wgeyWw3EmABJJ9CCc
Jo/IfzxK+Q4ykmWO6nTxqegQO+UJSZu3uLSaROeC1nukxK5VTS3sxQTP9vem
dL6sLtXuDntJuxf5Mhtb2Mr5FJTA0WkfhmdhqmURGB9tib0MLNGW1eL4y1if
xOZqCpP1WWoOn/ylDkI3qu3jbJKNgasSoE8KfOH4++zIoIvE/jOTF5Nk4qhd
iOKOPF+i1MkS2/c2Lh6tNYAvopDkyD/oX75kByMoLNfg4pwn+aT/p337rop/
4bLFGehK2p+fSs6zsIgXLnF6u0cPmDLlSlVfSKSfAK1rY5gEW+8MIV2sofK1
tgE/eZABgN5ikDyf7K92fqA5SsTq9H9hRNvhmbin7lBhw3sX51u/IN4NXPwG
lN82FqnNVb+rPkwRpEVdximjmgPfAOFX+dX0YV7oWQn9n5vMlEXOZt9Ow7+S
27PgCqb4KiTTeUVMAFL/ThM9c66N9BVmXPve2IPkqu6MgS248u+y0dMa8OAb
S17GO8LiYyIPnD62Ej1I+F8Hf4ROQuHRIZQkKvp1ZTGNqSeOXc/uBSYqAC1B
mNXJrtBvTj7tW+hoqeQYFRWmAncirWp/3DQvotx5FTaMGo87A9hhr1i7UaHi
tW7S/BtD0xbCzZUmSgkyzWf28TNc4vI25oAKzeJM/yYMB42iz6CyTal7SLjb
HoEm3q6DQbOMSGVc4zB0uh7OoyKqE/2SAYcP+EfDHttmGIfO37Fgkgaz7M3h
x5+WS/sEuRj1tHvDighsAFAKr6QBerTzaRA7pfj6N4aWzwg8csDISmBPx1CB
ILsmoKCrcPmXXeBLUrYB1dBX9ao1E6POsqlBba9/ftF0zYxQbDFfwI1Sms+p
qK4iC4D1altVngY+G9NW/GJtLUTBQlwNa6kvaRk+nu/4t5RrG9SOtTc//hwb
5x8Ko0HkAhILOgWPic9wUlD3uzbzJNG2fyqeqSCRClWC+RQVpwF2y3UwEO4v
KW/vbwcT4CD1QuYVXMHPo7v1kNaKh6C5qUmDskJZCREwQMo5k2+LUG1i1Kki
4QGajaf4Qt4jYB+d2GHuhc9mObs1S7fVww07hzW5YVrZvDLhNBAyKeH3djLu
Ou4aeRGaP5Gdu38aSy1VOiWjxYsAYeS9OnFQerWwnTg+yYJ74M3UpeVQhiPd
hpzJQjuF32w4A7Zlaro80dUO1bCNoyEqa3W2o92LWhp5xHJeORivhFsN/PPN
gGt7ssOGlL0k/De9cD4K3uh5t/fJpOI2YttkSleju5tKzOLtdrIitkdq1qdm
tRBkxki85BvdYXXCoI0VUu3zjDm13duSGLEn/VHW0e7n8cxg4QIsT0zsvyWF
04Gf9gak9U5axYiqTad0Tx8g4zCJ1gfcjJa1cH85BrBvhQH3OVK93rFZE4za
XHeTDizJn7BDArw+F1rE4E8zX6q7qelSJmnoSNhIt++19kPT2UwXZrnZTrTF
EYyxIOXp2t6nvCLc1Yjxn49ZAozhOkHIGLa3vHrf0Q5SJWeJsJxN2PysqZrS
auu0QfS/BK91Lnel2ESL9TxUe9oRVnRoeaAIoVmutD9AW1b5h/3sVnFkEale
zRsP7tMqeD5wvzVOmRDwz4/TUHQPMIMFRAQKwkem0KY2Y7xDP0+8WdZdYLZJ
RhmVD4F4AJkOSfcm9x5ql9dTRFkvRIPyEJb0npJXqJkB7qHq/Mpj5/MIgT2f
nX6pMiAt5Ks2dpMB3uwFTEyGkr3Ari7MU2PKTgu8YLZ1gxVnc7jiKLCj58If
kaHZnCMzVinH3gVXsmMczFw85cfl9pv4NDTYKucREGqZrMINOPQdVkVobxdk
5A+uoHTmFZQY6LcLt5tG8ePQqwiOP2p+ftUqTEdP3mrXLYv/FHUFOjFhjfDv
CgDfLjWNJ85rndSIVYAP8LXX91V5NbT4OKbwS0OdhPRnGMj8MCwREzTHBaXd
5csViDGN7P9GrKvk9jaQ+C5HXFES/YMS5bc9Dbzb1Mid1QRglpUUOY62BeBL
N353QNiF37dVXiIYi1zY5xBF+CUsINEdfuCOI5gXTi9uhouLEa1EfZ2/jDBi
zIQj2rjtXqrt2zlBoYzgNpjMFhk3kE+WeDqDc9G9aPur/fJAP493pLlB3WN9
h9JmEtl2feqbwP/mySBt4XuPF3HSsA+IxpjOPJ+MlguZHrfJroSUqbNbSbx1
bCbCQojHtjQRAn0/nulK+r749bIVNpGgzLW3Hyie35v9Z4+IW30Mx3sdATJJ
cpOku1imY5n3pd29x5wpkxP/kKMaA+r8aSJqqbtzQQS2ZQSp9xJfR6TXymS1
uXkeIQ/wIOeRzjU+196d7pLbmO+mn6Rt3GMXcH3qvHwMfRs5XcIAjpL8rvWf
ReYTfKNWU3RdVGwDhQR80LtvY4pJy35MuDyFjKjFYPC+xu0zwgwqh9Oq2Tol
If12a3WsNXzt/6vgROQthWRnQ5G8gDCxa56R1c+ZDNNqXFOUVBsibDMi5SWX
6qNBnO3DotiwSZHc+QoWFEpFE78Wmrd1x6Pgar9BdWUerdl8AebE3YF0zUIJ
RLHVTFz36Yc94xaQ0A9fjre+gsFg7Q/AUtsQBD7sQNjpSXvIaorPbzPZwhRD
KuBv+ZZsj6CcdeMifa3zx6A7KVr41bzKGT+vwSvKJCGttiM/3L7hx9byHYQX
HszHGfz17sFQScAwiQEuHaaXPVv3nyWJd8Q1LFgafhZI86ikFN4ycL+CZE/Z
gF35027BB0VC8T4zEwfdjxY7h44cAZS3zZNI9FOPzzdNw/qLbfjQ+8wqOK66
xfVP+ZIQBhYOiZTiMQTTredPCBCzBVB/hLVfrkKc4ppkc+KX1oC0o6kdbly6
HaAz2g/PBBWyM5V5o7OBo/gBdKwpe602Z5hp5jJDDOJqZrtJis+qVtrZjENX
1QjyJ0Lbp7dzZYB/BAzOpIHnOI5tw+krI1zKVzNIJSzMkBvCjS36mNvlUzQR
p6CXNuTAIe1ioyCt3Yd10sLVngyEX3Wnl5dOA9iyQVtwEerWDZdkKC1t6RbG
lxZQihw3VTSSFUI3ZCxRFKD8yWM9xVMNcYbIekc3QuxXjARQkEM2gUAoPcpt
u7xMwrZn6NQ3mvuFOWXI5dJYRy3kpJ9aMAmrBnoHc40Am8IjrO/Gr5kV28Cw
clMG+Of2dhuhu2rjORb+WVnoNMqlTsAHdHxN7rQQ+35WqMfc+OjVn57sRU+3
QGWWHuV+K8hJe/XAsIuQBXdPfmLeFHHSdqDoIuWfKzC9UfhOCRheR/SV22T9
b6Pf55OEgg12A3PReCteGWMzff+iZAM/QhyktRKEgPoZvrBBVCi/A06wyKQD
65zPfEQMxdhRfZU4iI7vTN0JP7tZUtQykQiK3h09aO8SibLYberm4cKt48vk
S88UjZkYEUOry6sLgokm8gQrE2U69hHXIPzpZsN4E0gZuJhw4UW41CwKiP+m
bA1P0Q3GVJKAQ643RxmvGJymzHpH5MuBi7MMmt281VigCGaIYjJHhE9F1eAP
xjGYU9fLE6mEUpMWjuYa/BMU+FEhT04618L1ViV7bPxKqRllTciFqUDY8uQO
gAkhXB7paX269G+lKnSJOMJcNFTXVk6bk2dHAozPwq9ClKZaR6OiWiQWyPdM
YWCLdmAQBg7wmwSIRbIy8++cfrZVucV0ThsillVV3/H0/jAjdOceDpQ/4Xe0
DAhUIHIwMQ+tg/Jun4k5tfdhs3Yy3LpQxxvBn7UxDbnQbJxeMTMikfIZkc+v
eCIp4P84N28EdSz2oDMpgnCOxhGgApdG3Z4quP+D1fOqKutG4hwF9MwIPnFc
/p8wGM1UiKSnvuni0wcItGBficooIJRblwpEu6hWuO7v5qCU1nWCtCzvSjmo
8dvUTifL/7Yfvy642SBELdFpn1voj39XJ6OeuNm+P5yFwSGQ4w5+xpjzP4Fk
PIfoxEXcF/mk/tK04IJNsc/yi07IW52HuHaLIxSGLaRiiHx9PoHvSG1cX6sj
l9h1SwfvusbVRJ/uRyC5ov+PNJ9MkOwH/ouQkWgZFdWH15JSeN6RGfeRDaMv
oVsbbr5USmbnhJD5rcVvm9I49HsOUZLVKjjZz8OuzyuCEXPxZwSy2RZ/Sna8
2wnDoTTezJOcBh9/GspWXWLLrG4b5LVzPeZT/attKIzIjZKPYZ0xK7xIF+v/
MTCcZUK1dNPs6/fTruoRlOh8IhpAQEwR6cjCdrU+p20dOkAe6pMF4ZH1ZJpz
M6m2weZToT9mjYzwJRi8x19LxIc/5jK/6C7xDy/Z2LyM5B0/AUyRKH5ecTjW
H9Huq7PYRjdwXggEYa9euW0rFhcmIF7Cf0LY8CWhyY9McILCNM2Z3HdExOVQ
re0cTiZKkEHUqMNGPA19NQL6+ldmKqaPFyhka98Gr4kvxIWKC0Yuy52Fo6LA
6pGImFshWRHD0IhzDZxWgzMuT/H5K7FwV5kVbhvl+B666e8wsp7LFjHE8WtH
gy1xLK6a29QFbLK5EauaKeN+QwYQTBIsqIKSr1qntaEBYmt8IZr7GCYxqzYO
8ejo0JKbq7lCCUJB1P7PGnDKss7ZYBkNB3D2b1S9ywVipJ8OUVDa+QZH0b7I
ubzvCxCA0J6cPbUzm0xug38cq4e68JYSmNN0zq8GzOv1ygVRqvC1SAnbtrtP
/m/hOZYkEzere/j3M7o35DLsW7osZQc8wiBAVCeQAzKDx1WopUpdVna9/Ofd
0w+FIMRdQjuU/GxJ7+OlHxI7PPPRTnk/f7PQX7WCH8dJJZbxsUv8YLvX9KKu
W+h943WlvKYthaQsBHjK7Ga9BQN8ElvNU8Bmj53dUfVZeR1wIYFflcxY5QT0
ZXCtCjEBr8/mrWqf8UlBjnN7AH7SczoPboMdEDw8p+SDbmWYEWNWdfP/rIK1
ts0rv41E33HLWQMXZ4Prf7JSIIMbxbeeDvrI3Gf4KrqEaCZR9RZKdHPGl9wC
oqebSelkN1uniMbVVh0/dIpKlpVGoL/aDgxwpID2GP4XlOk8XW2seM2UFMMM
uqiIUMLmPI0tljtqOyGonbEwyhffiPm0ImUcEqOnlmzgMS5+vEZooRdlquAa
7TyDp3SwP9yRynlugtVw3CHfX0Go5SasWPs7T3088BznE2bbAHNH8Tu5mnWE
4DMezy3FUZ65M5LSvAo2QZawFP2iY99y6ndILq4SXiIrQ+mYiaYmj3pg54p0
IbHuPYDgbgKAtVjg8ElKz/w6Si29nr8aGlsGQvocH0rZcPOD0nifo69pihoC
pdtjkc78OAg+D+E1cfsbPcFAFpklsTDa1gkjycXQbRK7XbRXK76GfJgr2IaB
qk9llPF2pWnPBq4gNLj7xIwOGGhcb+3Rlb6zvcZ/19EWkFW0tGiwf//Najk3
X3Zi6zktBAG5IDkiBs/NtiiC1jGUBdWrYxJBbx2b0acIqNNkj68se//gUewl
t7YdTjMpBwCxq1NSPxUHe2mJhQo7vmdk1xN219aAHM0f1cyi6ppwwwrCjFQv
suPXVxUhI0ye1KxFJBvR8QupX4KbiksUuTe0CroSDXdjWO/12F6P+6P9lQk3
dbDYa4ZD73Nfoa2T0FdIdV+rdXXXWzPvZxQcDwJHRJzA2nFKmfLN3qpSq/cw
3qYwBDJcvTlpmM0a3GCUumR/U3j3jBQ6Qdw6Lj4/xV2puCEgIy3jqSQgcJN3
EN+hQWDVwhUsP1fSI/fPw0OUkZkPTXC7ytbMyUUE/eOqy2XlbbqfOPWxY1MC
z7lmAMGtmwljHJxF7TG/K3a1BkOG81Pk+HxgjefkoAKmpqrBDb9isMC2bUTG
s3kn5cU1KkcBkAih41YzE7nHryKA1j2oAxuNRRNajIigH89yAkI3dDgbZiM3
wFAOILCxX2UNs4wC1r7qKVyWVNiJ7Lt7vfmQZVpIGj+TxDBnKQjIHM26A0ku
BcBvPjcoEkg4R+hQ/tQ/E1xnFeV3CA4QDMhEmEJm0Pjxwu2NIPQ90zvAyFhP
sE8qcdcc3yDDcAw+3Pt3+TecDOCQHMf7ihpHF4frA+/NJ5swiLmkfjN79z+h
JryyJtKWfaIOeO7+6mp/1LNRFsdP0s2mRRmaMSXKTgNS01uFotoG1Oon+lVR
UNRCry+Veqc9kOsrXP2tFXY5cjH82SM0zwkk/l0WAx7+9y1yRGWynCPpubiq
fz7EmxIcyVGxsAh7CHndVDZbeXAAEtc8rouDpfDJCkVaebAL8Xhrz9oy+zO3
fLkxDcQ86SAIWNyjoLpAvepQDH7K3Q1grrQpuMhFjLZwO9kslMutbfZuADQY
2dF82fM3OVSwJhLEbKP0vkx+mTTzq5V5o4Me2klAJJ2d/JIvvowI24QTNrpK
gMLp/Cx+DAnX08OyNKTtNGIF6xVDUDqeHGITqq0VDALONXYfx9p6p4o4dsE1
BI5VO1ShvRXkLFwVQ6gCj16boiCLoptO2Xg/SY+vW8FDkObt2M1d/FGqo7fz
T50H44NDUue3VFxrviYLTK1HDy93ZttMlQW9ajSxnU8k0scn9sczPKv13bn/
lvAKBVxTOf1WzUJp0GAaGBcLKJo3b4Wa5q2DMUSl14ThPuLLjDLjj7QHYDs+
0ulOCBh0vC4i9K/WFXbG5YJ6Ecl5B9B+MH5HxK1yxMoRA/3hFWPGnAD2F9iU
dDMtDFkmoaGeV28JWjeeMWogK4SVMuNjaJ1aKDiShQSMAhEv0GYMtlt6gz4T
9yYQqHhzDW4BzENMfUNx/dPxa+1S3KYujUN9wPAuMme9XP8VDMrnGDXec3yP
ZlVBV++mM4eh2DMcJNjehvkiV0Rbqb22l4KfCSZ9GXHw7Ob2wDNCsdhDdkbQ
X4cwsQhPQ9n1/tYWwEBGbbWifi2XRbUD0jBWgZguS8R/yR9kbuQCTMOVeEUp
cILg6rqQv++i07RMyA7fKTFCuUKCnlqfA/wpILtIJdmrLSIesU0+d+zHYUFw
eofKIPA2ZZM7GpzNncNb2dSeSJ3d9KIgku72SKRX4lEVwh4Lb3iwDlhIUK98
fxZ15S8K8n63mqb3SQSaY1//LYTHY4kyIAbQlo3L1nH4B6LlKxSegWgZgnpL
X2EwFxf7/Ej9RacsdEAygRtBG0V6pH/jqVQy9f3laASpKgkXPBApwHdaJzMg
+UfvwCCXL+wIhaazVckw4efQd2JuEeiSvlRmDquviIIlNrwM0f8hp/N67Kp2
UgIdZSLDTgNB0xGalKdD15HGOw+5wQewqY5dPvnSbPzScV7ZmcMYgn3GgYit
sJhgFXuaAuz//E3tPBk5048EJz/anVtt+8uvBfrUMcmIspsWKppRZrzblC5W
J2WBI5iejclNqlrbqbgRFyKwxZjwmH6K8fOTEAQD2JZRaFtep/5VriNIKC/R
yNIAiopiEmpgAi6f3BrvgncqrTlO0esFR5kOT5vmc/vuMFmtpy2E2EcUcnex
1P3TJQMsR3DlMf/Xl7ODOfStk8YJEt4XjvqzCqJPeW4E0rrXsgx/vUSssiPR
dua5qrWoMtWmXttv4xlI8e10j7xDo1GsrI348wiWHuDLP4lSaHZ1yN3T6M+7
qZx1q8iEyfBNJBlG4Hx6YWowy4XoFmq7TIFYFEYrzOLDh2eHl1c4fmYIejeB
vUw0cUiOAt5X0OTZsYpL5zSa2RmlH7oHmaIdljf55rGUE4RgGTPYXurdN4Xm
yH3tUuK0Ws7p18d3YTD8WR8L5NEVXZiCkMAw12co/8nxlwVgoJH0/v9M3cIz
/oyhUWPBGIEJFR2Z0MH/9YhvelAroDE7R29z9zf0SSNI3YP3WMyb6yqNYPZP
+gTOowi2Q2u6YIXogdSyAz3ot1BPr2A+vBlEqQOuqzRnNLRZh+2WYgitSB1+
2HcmVMtKxFP9SwSpd/DpaeKg9N+x33Tkp4ESg5gXo7uTh7GW+PHGLTyTzEM8
/kKVuoHZJ6hUjtgi4aqqnbFu7zqA2HdpsgQgWZd6x3FdHlNdnzpuwMJ0n9kY
gIdtn9U70zRoINv5IwIQS3y10qIVw6zzuFlPVl6ELG4lI4i5rUlXEfdHQnZ/
XGzuJayDdHelZy+lDe4NVj7Ho8/G5UpxR7BLigzGFvPqKaFSQqTW26p8vDz1
4CNHwlbHwAGAD2Rq922ulYbG1zc2wTJQGltKntomlzH7Nojt465PoQ2Usstt
HUMm736u0N5ZPxFfHKZX3ybYsl+1jl1a77L3IuevWs9K46YZ2BfKD9xKpJLO
JcZhYKDehXSWIX/x2pnGsmWhPyhaYHj7p6WgnRmiC3Ub2TunfwLrno9G1i5e
6Th4s1fOsAiHIBB9mFMGrRJjP5f1Q7/jSThOmDo8TvvvDkkP7V07PC035ota
3e+J9xKDW1xhjg/FXYpkC9RU8TvykcTfczc9jEdDSzh3YkyOxDANlatOXFnY
dRibJt1j1sAOmD2/qjVLutTwpedRLmQi18H2wv5OKA22Sf433Wzioy5PAIEY
9UmyltVruHuO0niZqlisJg4w4geJnxGCbF67b2kr7OQX7JSiAZfXvKDwm6ry
QDmgSRWl5Dyo+s/P+diYAhOmukl2x4eENTXh6Bdd1KKRu7onY1eOYsxscdcj
rwtaUdOsDZ2mREbdwtLdTYqtZQvop+Co5pxC7ukP7dh4iEDz3LLlkYkYWaaC
M6DYHO6/lZ3xKzlDBgkfIs5T7VnT4gkvxAkwpYI0htmQ8bMAknMo1uworfRb
J9/OClcD+GffyFC1UuoN6z7kUV8DruMah2P9YNM2CmzbUOM7dmnquC0l4fEh
PjcTZi+bcBn32HmBAVKb8+wwj11g82TDU2Q7QEYOpecbXuDoZhphknUxepD4
cyy39HieWMctd8CfBwt962/GmwzbZ19mGMbA5O3MMBjnTiUYs2wNt8Bm/Nu7
IFuWZLWMl/EjfBKVJ7wfKdT7SFjRTKduTpjcv0Ag1D1OplbssomepH9pUyeu
y7dHt+8AWY7BihGKYlKIDxr6julbsbqviebRE81txoAFiVOKknikFmxaeDa+
IdsWUlutiKvvPR78os5bA0RhsklPKaAHJ19d5jScWkwnW+X/9dmzgrem+eWe
VYgSWX2MRKOCddlmpjII+RcgxKmNnEqc4NFbTen8KeMBgPkdJLUYoWaakmNa
5AQxnPH/Foi8TJWlRJqfLMRqbu+1itVM3IL3Y9q1zyXr2x6F2YZKzS9uIGGE
JyNua2VL+/OHL6+elbz+azdRbXSKWWT5g2crNGwrqDUJi5r/UC6Cgh06369x
NqIifXClBrEcsxziaWmRAD05IqeOgJpv05NIU1nXE8wGPFgFnQG3Gl6HIzZM
Ju1JEmxzdPw6A4T/8NxHRtreR09NmAPQIo1u7n2a46y6aO7dkp1z4O/0rl8o
eRcrtdW9kcPMvsUoUl9i4Rp25umrfXVsVD3F22CSpWzScq3T8fykynqrteFQ
/TuyEpIApNzqzYS2fAgnpqy1cOSPlJqDwFMhOM/z0Gt/IOBHKg32q7+hTUmx
OL0nvQOs4lhxhghZdZTelO7RR9FtmxN+6QI6b0ZeuoB9IwwSm1QZ5PgjTXjt
Ts32N9Oa9kWxbUSjlA5IngzXNvAZuRn2phYXiEMQOQHnAPAw+zv7PSGQ/R+Z
CXD7phQIJP0cWR5fjfbKzYA4IujXjUy8ATlp0GjpIxl1E4S9GnpfmGCGSUTP
dsXIB/TaMmQbMzqtaLwjkiT8gkmuheDR3/+dPnGzJCer+WtpxlFweq3W8u3U
rHSpTtvusoV+TKPz3Lx4CXNkBVsutOlgVaIazjB4XU86s8o2CxYWL440BAIf
PlG62OfA4y+B+VcRR2IdmlvftaXRBAXaQJg+mNpIeUE+zxeWtWqo+Xzqn+3h
Q/wEr4Dpsn5oe+yW/DPZ25Pdapv5kVV8Ms9XOSrQ3ZtSHmgbPWywq61+DNiD
mPEGeHhea/yuWLFLKs5mHt1sBVKLAkeMNqi2NVQ3ZT/fZWeUC1uZ9jb4JIuT
Qd8CAofBmQT8mgqYmZks3Lse+vzFtZgPXT44LpDS3C3aPkkaR4mNwvVrvD5F
/wpNKQSAKUmwHpGaU2RHOzekth1egsJPiGkhkt7x86xsVOclvJpfDtMfE0ro
sPbGgocQ5jgxK8FMPRAhTtkVV67oY9ofsR8If/FkjsUqV6poKnBSVv8J5s8c
2q+xY3W2+nAIntWUvgcTf6ycq64wAR8YYFdJDC3XGkVYia69tyiXSagFwvoo
DfdAgY4lsC2x/TEnF/tX1bz4IHK1X1U7jZSGfMfrB8h/qFBRoXamJhPzfXFG
pyfnZHZwciKYbuHhlnciZgAkitVElijxnGPO2rh8H0sNSrJwkAK8QJlGjw59
jcLJmvqWeSWGfYCG1rYGmku8EXYP3FAxaceULNiRibm0VfCx3T3pIENqPyQR
ty9wDD7Gzkq9VLXVa8vT4uKHV4NvmOjLVQEovATbHqomRYqCj8o67jz5Btq0
A1m7uh7aBml5jK8Fhv65ehRme5PJvlOlIm6CKtoXHb/awYQPq35gTXqdzQYv
xYYwTffUcU1gYJeliifYun3Zmd2PvXv9117zr+UuzBwpt+dONwpVyp1bPSP7
5hEzlvEv8MpHAVj6Q+tF50CSLHi5832vI26Rtw5zw4iL7ZUhKRmHC0+Los4b
NhCX3W2Sd6cCGkRXtIEoLTOEzYYwRD1HJE5K+792z4SX9IsWqpQRl+WGPMv8
c4zraY21E1Pb8Sifjb2YRMVI7CZxssKv4nOpM+NYKdSaMmZ8j6ET4UaidfaX
7RLH4MH6HXwt0ymJMStv5HwCVFXJKkDakj78K0sa/kQcPeMam5iyOW06fMat
tzv5RteP7xFxMnf+3V3pYYBMKaJa42ywETmFdznl02bYk8okHbxabqC6uu+3
pmxS5T1lAKwlmXCsPA+j+LOtXhKOd/Rr9FyseqDLTaOQC2xSVyMSzzeFEyPY
yaZ1KvBBEFMqKmVI7yDpE5kGrrZEoq0bQFQf339hXVGHtN4PMBuanKFnHCOG
5QqxcD7tnGtuYm2vYKitj04Ih5/XYQB28Yz1vW3P8+MOXT1h5y6B6RU33UXf
qryE3L/V7I1JvdeSRB8ZynOkJ2gFeDp/J/+jTxI21H9erv72Pak/KsZX24LH
u58yFunI3z7mUuYoKN69l54sWAHhwJ7+b49K/br4UomvbWUydZOWLjRSMDRC
LTblybU+YdI0xwgBsQ7rwiSX/ZGhy6l3ClAGvAxoCnvVpC0JLCW7skdvE/SD
0X28yrLzrcJwRKOp9nlNCo3B3QWV2yqXtBw6Uli8hbQjjwjGEx5/MOD5hY7S
ReIpQDup6svKL/fBDERIbJIZLBdn9HEwVc0r+D5C6D8HQDo9U9CxGeVoTl9a
sZ3DjXjPiqqLdMuHudXNGfSnezdTbnkTjuciheJMLvTOvEK0Yfi1BOD7u8UQ
moRqNcxIz7sQuajS/MqKc+Y6Pfs4sdj19nk5cTqXy2C+zaPgnim1PB6DuuaE
kKc3ms4OjFoJWmr9XimQBRDC1ohGsFRhDsmxuiu0kG083imf8iXmdq6SrJzd
TznEl7QlfsdzOVKTl9GjveoKJUhejpHJOanswbtBa8CqBVHS/8zi4ry0ahDF
qSq94EB+wO1RFNK/bMP58MDr5JC9ofr9r5OnkI8ZNdh4XQl0a52Sa6zFY4JW
+snYzRd3seh/6NDIq/xwAITuNO8ULXCo/c4kQ/2z2EYqmIHF+/7G4bThD3Eu
WG5ZVeW+m+O6deSpAmv3NtiPnc6ZN/VwxE95YnbZ6CNvaUA/KpRBVhXRp/dX
lcwV/V5eSiNjScuIr1G/c2d4lgKZDjpUeXqLbmSjtUyNNTiTMc9qJVrfe7A3
HXH6ggVYiM5DbtG7JI0n8ZLAP55nAM1wrws2csQT/LSObvU/YDcv3dG/j35q
VMaqV8DSPxpoxQnXjsf3sJJrnYqdnZ56b9RQ33c0b7QeXxZHnH5HOm34Qkg5
nuR0o3ACnSzpXKpKCPCmPGE633sU/nZsfIeH4tmHrQrcwBRi9p2SyypG1qsp
wCHOS8/qcnZGwDbTVy1EtpC1wI/cWxg/wxzeWbBBzpYRwv7OMLYCjeBqiUol
COUfQHfgIeOvJ1cw/3NHbH8TsmeTH5NOFu4JZUSpfQFh6rMBRdVHxx/YFZ6j
U7pxOb5GPKbm2uEGjGruSeaeBU2Wx02RzTm355tv0DKJOfq/TlsvrYmEWRZO
Qbfu+aEKZTP32wXzndOrUu7VFlFw5/tLZfm168lJkbnEPtbORg1tK4+9/w64
N9xzkBnoVgPSRvWCsyAEC6ix3rohHq7Irf5UInWRLOGrjZzlRdLksdvHc9JH
kK2r8+Lg1PZorpvUC9H4fPi6AMd2HLlgUpK1HBXLBtbBykCZlS2kKB62jtMn
Zppt7kiElZfJOGmJvAWzbRuBsJzNF/VTSUXDxisXBihxnqnwpACeKooJWw+Z
KdJ6k8mlhdBRb9CNa4MNW++ZegRaqlfZI9Zsie7GOZjOxMeOBSnbSZWpVw2p
vE5JMxdU6H4B/I69FE4kwxt/zZz4jbDP+M3QUsxLpwM54WaZTN7wlgHREhCr
kDAxhI/mDzOTn/7oJtdgVTm7/NasS7R4Kcp04lxbtMNRHcpRO6TCeluop8l+
mL81MemQWcL/lnh+Vuy3sJguwUDKhCK3PqU4XqPt/9Hjm5C+U6wApxACUZ8w
q69422OQlBw8ADhDPrl0uQffPk3byb0V9D/zD1zCe32PUwQp3PAK/J7PmxWH
At6+y6g+MpmmL/KhGgJJQ55VcxbIDhOm40+VRVK9PODGjYK7qcxu4XhFnzVF
2b3snjdsiWVPrS4gCb7Yx3oLF5Lrznbjw/jg/2BybLBwYaUBW4/mnKO9zc4o
uu2z0el3ms7ZvJn0CUEE19pj1N+6nC5nuofetn6DX13LFNqaQPlrH/t77eQ8
bdqM1GR8AAqILHzMXCelIVKLJRKTrSRrxf8utg4p/MBydOvYbFfLjTAC8Jow
Se4ysSmi3xvaobMItolrUI6X31f2vq/74cwbmUj9R7htd4NmOqthnpxfNtFA
iZL8Wi4s14bIiwOS1T6DhjQKOwKj0yRUG+zyeh97BKrsUmk1Ex+uA3S4zFZp
Hta0RLzjMt6JDTV6FZriyy43TxXodWpHFPuyrEQxgu1JbnPVeS5P8J5n1+S4
2MY2Y4RwFQGngRLqUTQNyG0F/aCJBZMiJv0rfNr1NYvKPzXnyBY2XIATPdT1
sGRZ2GWkmALdL/kxLAboI+CBV3Y1bpsmhF1ChnMI0jzkNMLj60jO9NeZtKPp
16GF2UUnm2UN0FhrzhbIJ1IFBRldPbDzbBCLXJuZQATjGDgQ79Pf7ie42BCC
EwhSa71q41HRlZbS1qwbcNlD3EW7a3VuPXQAh6dPTrPGAu/OkFq9A2nLq3ve
254hFNE0xT/pr/1Ja+GLVrbpIJAK+iULnI2k54DVodXxKVgbBs1QZo2BUR+B
vmJMzf9xs97tJAEttjqvKs6YjgQEn0WnnpkRH4GVsXEiL6ollveXUnv+PaUr
FuRQj0eGGFUH8/FfDJo+mzNQTIUgLpYvWaeM/ECztCwX4nYcimdlFBI0tr1O
D4DYX2YNtIP3ZC7zLao3wp0jR7bmdYYZdKL7s2Uj+z9uuuxSSYtDAEcGrk8l
i2+4mG2abmPVn+ZjP0TIyvsaQfUsZdCDVYtCFGOttab2PT0P6Txm+IeBocrY
sONrUAIfIHS7x9kv0f9GIfXPFKrPn47sBnqiz2OO+j4F1cyPnKyWtsz7Uf6n
PUc6YdfKVvdTobDpuXAhLiVgBD76PgkfzpA7QCF2sqRWE+ibI2xMLoSTlVlM
DKOBbYaRtpj+92fKMbEWibJUq3QFxjylwIC+K/4oKY0xFA5R7PCkIx74oTns
W2zQ1U3IY3OCvLP4wYaEb3YUtvGgkaxKJkZHtQcjdH27voWLaGdsl2r6CZ+2
MKckEvXxNc8shCdTJse4xdsLmwu2jnaje291hHrP5UlqWhWmNZFPTfrAWz0o
DLXYKMlQ/0a9s9mHknAuD2SNqEDwbHSq1rSdfAr5eGDCIn7Qjkmqmv4+32gZ
q99Xo3he/K/di+Pg8sEcmFIfF3BdYzAA257NBdadVnVT8BToAZgd0SJfyW9Y
FcJtEwKZceq+1bZbRf45MTZIM90FfkYdf5DimUO7ARQbj9idEh9BlP/GRfrS
UEqaBrtijOMJ5zlHimmnKl080Txp0RNuDDdXjGIFZBPU1Bi+mxQUBupYwlBl
clofzxqyVMbH1ofshR2jMhxOMEHdOg5mqq2d3cU87p2t6+ouJQ37cFbeWZSW
86BCeLJKw4rKIm1aFl4JhjWmcRkj6sTcDnumofmV84j4j2G1mzfZk+BjIVkK
OCoeVK9IOMPbyST0jVwfZZqqxkJ172UPu0xwmQIBuWpCdwMOGtbC89sCBbu9
eSsTwbqJRp1V3OBSR4qAAF2PbH3wSEwLMEVAwExrT0/Agmw9WP/wZ43p7i1g
/fBc5GbeQz01okrrPrDjGDBPLCN3dUxUfkDp5HAJJgv5AlhvjT71PfN7v/Sb
67yKsx/PP0NxbZPgCxjQo+KYBqrM7MKgtqSwQO0k5Rag8m3FQkRh1IsZyGn9
AhoahDE16qJ3UpmevT0D9v9fEUvVvqFnEkMvc87qIxep24wm7FCHT91F7W/n
6GWGT6GpGK5X94qqfgG5NooXPgbcY3huKMT3eNscxGXYJ8mxV9mtORhgSSIn
r1bNsWx5jLDMXnuA8NQSFhOZqAdKvS9X/ALGS0IgEINfqoAv6+hNQC5aM4QN
02iEa5QsYwPE4OpR8JA1SBwKguUnR3RcpfiT1czWOqdyeF3RS0YUtTg4d5ar
wIhPcHtvkHmg4njDlxZbVd6+a4iDK6oyrw+D3FYWLlZSr4tQugeVNDOX2Ss2
WF/cyKdri2JoE8y5jfiB6WlWIO/0zrNnQnVpbRIVf7WbXkUursFkMGCdNTd/
ETGeOig7sN0EWmHb9TWmQGDN+bikgQFpYMlTuj3HMhOexUYW1WsBRt2Hbx2u
4bRZHXdTToyRQJMWeSb0o0wKWDOijUl2IlbKCEQMKMyGfQvrIyE6X7bWbTrf
E9p8tHOz3K5ezAaq8r2evaJIS/zgfSIxBFHYJYEOdhIeAL5k4ai8zdjKvd94
547U0odSIp50fk3YzbVSNJRXiofVPX5zfotGRwqg5CBwXLXSwoN8uWkAHa0f
kTqNB1Gof/g4vQzU2AWPxRbmYcct5w45mwEbgCpm3mZM95F7e+MV/SYj1omK
wV1kRoBj9yMO+ZiKqE8wdml3fv6uuTuYFoSc+keqcguOoCw3O5kFGNW0hnd5
SVqcfZQVUw/XlGHXl2JF4RCDNLIdfyYqeTeRiHDE7PHX/pv4x6hImLeUmups
bZ45t+NLB3c9e0EWGVEsfDT5sMUmyPCUVDVEcdoHzntJ/MnfM+lR4CYaWtzT
eFxQC1XusdfK643nnGCqNfttGCVwC+aHtqcwO5OstiuT2jabqj1xlO77jkR2
T/vGzE0H5VXjMSOl85OYOhdgl/c8Td57r9RF1+Q2IkmUgE3wf9bkieB3j1fi
VVkkXGicLFHdlcD6wN4dK/p0RDg8DLoFQADnBMwnNy/rcd8J8OVlZQRt7qoY
3YfVZ7pwhx7Tg6FEhPP/o2whcyDOuKUG0JJvtTn6ikAigelzJsry25n/OCsf
e7nAuzQrZMUyZT8uUsQ3fZdKIMbGvdaiPq5tfnonJ1QyZvHN0IG+tSWDbxsM
Hh3+WNqYwgrHMvWZ1sPvdCrf9KFvDHHeGBr/jYOJ05C4Bp5FnWK1iBqnyAHN
3CMHWtGwQXYl74yhe4OLWmI/yFCyDbcgNL9lJEVlLTa5aUp+0HIvDEYgsuqN
MDi0XIO7MEnqSuKeelq+amOvTlhDHIOzFut1a1aAq/81PscqYrCy2g2tErsW
uVEsrJvzX+EzXkWt/cJzVYFMt7EJQIGqIiBym/zsen1W20ILhKzEy3k3GxCl
oSooH2pwiTVuiBAEoP5rxlA7jwPCR4wx3G7eAFBK4XtUSKMZowNt/fi8An0Y
4gQMG09DAAA0WcIeVRabsXEkZDAKQ8GmfIVJQMg4qWga7sDKgp9V6VDlGmT4
f53oWPjpqhuVsNBH9vAGwpXCynsUYbBS/ZYow9T7h4G6Upnvls3lOBENiPx6
V2a7eNIgr60aFIOBSMZoJjowU+f0M3cVtnTPTAroifrbC2BcNmLDhBzlrLJD
MGg9cpSQUc3TpUHbG+gdw6Xbo7dUXX2Gr0eyHtr+ZUFz+tx2FPeqeNjx30EH
MwPPtJae3x9GgDo1I4EbyIO1niBQL4v6KyQYpq/vZfGyWdj9iqaZfdabWNqB
ix1e/nLp0JgskD8HZoj/psLCXU3PNyEkXqC3mI3iEd/cbwCaj393+kG5kmlG
1fh2c1W9aiql1xrrCGZzc62X/MfexTPTsPf7FXCnFJ0cmLbWnl3xUBvFhOh2
x8kR+HCFBouCR4rEcjn1I/8Jl2G6Eb9KLC/CC3ZNnpbAPD4SQjLSnapZyKKl
GUd/tEVLFezVgSk6bmVFp177g37ExNRRg8WANZi529jwcf0w+koCJ6VZs4EW
N1LDC9kkv4BreibhRvzU8gZFG0Mo/KpcKlAxeXz9bpQISC2U4qa0fwklkaDA
zwTgtzUDyoyC+TRzSgZHc1S16pKgwuGDv2IUvDabWqY4BPcHntCgxtoUgNOp
W1dDPmrZaFxXCi7m3g/M/h9lndb0BjkwvoBJPI9NW5bse2BB1cGoV78FxdFL
1VULxqM5B7TCB0HweSQ+p20jX51vxT5DAhQfPgOfcL+1IVsULtglRDDU6sM9
tqb2welFVvkLuLnQceZx2sF9ZAt9iikSVz/sz/jTimOeQcSrOALYeKwTvcTc
0m4ig4l+Kx9IEoTkV3ar71olai6RDtoJJfWkP6M74PTpC4OR6aTcck5wXRNE
EZXtCZWGpPpqDkmoe0YzWHaIcylaKfD6jnVPzbw+sjtQ5kLjbJBkRPTUu+mG
oMHgQCNWuuGzriBAjQ33/zk82iDDWBANxB/+vCYNSi50vv2byelB3aOEF+c8
n8arbE9Sa/r4oF7Gp3XXDtor+yO1cbziCWkK8yHmUpAf1plXxWko7oMrFyIR
ISBKhER/mkAf8Wv27FRDkR5o30tBMNfrdrU6KU3uE3d1IeXPrtOkyvMBoLlB
+9PwovTgJ9GlM3Av5U5eLAQmzEMd5RT1pzsTOHKCEPdAi8nYLwWUj0qp3rXB
cc14G/RRFwl6R4Tcxvb8Ye4dRJZ4NGXIc62D8u5P/F/TWSfFQ1QQNIBuDAwq
yEZ+N5a2u5RhUNjLLdR0SOqmfPeUe4mCMrNaIkYPM6kwkavTwxKusrPzY1Mg
xaoHS/GskN00SB9f3FTfe6V5BZowUg0GqGliiDZ5EfoidSKRqkWkWB09EmMe
Ar6amwKn7/kVD7zlH8LOSYksIctAQn66TsVn+ovwN//raLEP0mPDRL+IVKeO
GxIYIcdwr80ycvO/ghbmDTQj92UZ0eNuKtEl4KYxGdQmh8a5VOykXNm3sUP4
p22pbk8Y2e2G1NHukNddln6uvxQ0jJn1VwRFJWAR9SSHdVq/XGrgh3YaYgw0
K8gYkmG6V7MZBxZPBtBqyXAICubXjD+Yt9+89NsEly1onjmDt+pbZYx1nb/G
FK3hFTe+aehe57PnRYW+bVn5G57cdGj7HBKHk/zO6OXre5lxPRWc2zKj8N7Z
KqsdGdWPomUBhOg6FCLjTqeGTjT6U3aw8WvdIXVYW10hCRIRNuBUfhOv9lVy
WOfxXr1Wc+SIy660Ap9BIMR5Mq+QxBWkSBG3F3h5Kx8Iqb9ypr8hdWlhIbMZ
bSp1jIF0YFbR+B3vW00Nr8YxGa02bE5c2Zn6rAr4YY+8BkGUOZYCi6LrdZbl
NF7V43A/q4DLyMPu1C1kZccdWgR7oEcK9bsyiztNT9ePi1hVJgbsulnzPUGN
WRcgSNAVmNKALjvU2fuVo1Yl9MYLFd7uPo8ovyt0+H07J7DsCH+iI6S7lEZf
3mQt7vSCmJLjPIvcVcNSmpnIMW2/W8um+rVnfnVCFUBXH7UMgrIGp80xMOTH
SzKertaBjCSNuyyQSdn6dpyqhVqhhNv9z18f6IPSZB7tADYSuvjiyPkueAoa
Gwt886iEXBVmA3zVdUypnCH/l8sxAtqvefyLvpXBhe50LWO4laGjff5veXQA
MSP4C3WjydPd/jNsOb4E1tZPiKHXvNJu0Yyxjc6eIekozwJrR/WKBRymM3vW
1Ft+P9h/g41qJh1BZszWYvjKyXLdmdko2qMeOIlpB2uTR4IRRqHlpN8SWLBz
wBZdXzTJySa8LtzRHIWC3IrTFnYJG78cozo8zrCmnn3Fdt6/I9KV16BvzuiP
7Z5bTwVdMfsIEtlWW6EzP8OeQgMLDeJd1d5R9nrfB2NX02DW9bhW3XjiJ/2g
b8foknvgavgTk9KVk4Q6/C+bhlLcwjQn0/fUhKmE7UOIOSFSm6mTHJQaEXYy
qT+PyKdmzOqQ23FrguvOQ3qOIq04VMHyqR67Ti/aYDvRhnSPTUy6IUrJ3/B6
BjVvMaMQNbQAdjD5cc2oyWvzc0TPR1P7s2DGG7tyiyvmsit6TPz0DeMZ8qKF
lwsjP0A/iavvq/RhlJm2diP3QmkeEPfAvmyRakWrKY70ghcbmJaqxRqUtNgi
5W1XeLrMS7ZXr5UZXc/esQzQSaW5xB/auajsmwg+74Xnr3HC6HcKWhMEfTeq
CCL47xyqAuuacVxmc9jSlOEkbK5Jw0sFt18hilTgvDHYq2ctuqsfSy9XDIHk
qg59m1ljf1JThaOHFUpt/2J+47PFt/a/s7W45HPoJC9+MlDAL0epckrSliEi
KOPQvv4iyakekxzAAc0aOq3Q47E3fpc+SCcuyKIA9Im4gpOln0fxTBPZLvoG
uDgkf8jYHoRnkVt6m1D+JQmHzxwFIs667rjykN3rMBzgXP0ZofUUMfRPmfk/
w7gE5F5yMhS49TaiQv2ehq3P0qpQutJOZHykAg7cQe+JG2FaxXSW3Hr4b1o4
OzeahAHxIpPpAy7dnUbGbcNqhkXCJmupT1ehjtzkdSeiN3YBsm/7zIOUrhnP
VoDMjJ+ueaKQnB2dfLW7cQfvYs4IJvI8tm6M3wZtheorGYpvIubPvymjdLDe
ikMseRuRyOCPEL1yVq8M+W42Vt0kva7DqqUuseDqlQbjEc8aGns0WSr8Uoja
p/A6rHT270HqKfhH28RhMkIWtTedfC3Szdah4HRQc4aIkfacmQCN5Es10Otp
co2vyPvjyNfDdnJQQ6KwsH0imkv6KWyQxaRxWjoYgTbfNYnTjpvrzQbMPjD7
kV8K9IwENTNeOhkn5O3k/GapGYD83q5Nu/M7IO+GSpVUFfksWsWL6vYFNgYl
dikiZfxgj4ApeMZObj/otB/agqWXyG17oV9zK3s8scVWyFjajZeZiINe83+1
tuNGI7TYZOeSqGfpBUoK9H4ITVf3EceiiglcTVLVnrL+SJZCG0tR7juu0RL2
wvkxGL66xeyyEZ08xnvETJeUtijafeqo3lsZ2Vv7GbIhbb9t86gLEXGTxNNm
9zBG3HD1+n9DDQoXuh2nkh0kSCQKWTUGrVFFBw2S69QSAVvkwPY1XuJXTc6Q
TZAIQiA5/yM97ePMvaPpgKkxXXvG4koHnASPY3M84iGDNaqPq+EPkdp52cUr
2Fr75mVYqkO/ZYONg0n26FgmdRYQ5UICNcHIiWR52T3uKiYKYICOI6WWeka2
jYZfn9pZPp5Q3plG9kTBWxarY6jCGXa3Weh7u8pkr32PPS6gjZ99pU4LzBSY
ioCgGj3z/MK2LXyEgi2gtzKPtVcdekjA58w1YanYU6fDmTNZpiKcn7F3xXoB
CSSH1bkTQ6vijnnBNNMCnnVBYmbQxuveqIKF8B6UFEqwP5fpqfoRLYaRN8Yf
IdIxBaprRMnT6HOJJqtqV7amEPl4S9nyEC5A7lKhciUnfweUw/+rVkUtIgym
yvfxr4LATNTZED5pQod+4OIaaKDlmEAXsTVQloZ7tM/0ZCcwjNiddQSTnE4K
db1HOc/Q6X5Xy1MziAbCk9FOTIutkY1znNZy7LIBpjff1V/m+S6lb2qXloDC
x5lu9oEmr3u31yUgEst4HR7XT9IKEev1fJ7nDCDdjeBUaawhCIgtTkTO4bH1
4NizfkNI9bBPPfzuQ7YAljYrGxcFqcp9lIqO1Hz0/2t6xNEC8VsMKR+A3vV+
b87HBXmrhyd9iWkPYhVsoRqBwEqDzysI0qQlbuC1qz5qp5bCQPU4Udr4y/xM
VoqtwEh+MaZvJcaoHsnXYWxPbCewtTur9saA28Q7XArUltlNSSqF/rPHcRGf
euBtptAHd6Q4mkw6/h0vWvrdC6SO654eL2XcMhzFjifNpvULEWr3eTBx6CgC
Sx+PBBjP5lxhkOa2NJreaGdk4JDvDn7iksGkRoi7pclAZ1ORdtcMrEBYPF1f
9iQZerCc/R5/yFhX6c7VXAiJ2jtNqN3UfWsg56eFwSN5szbe4y2d6C+OrTK0
OU9oqy59deIfV7bl/pYu0xvJmSI7RDU3YdC5cmqUoKV5WfSNU1vEs+TkymKs
OzlwNx/2RI7l7OJUKHF/OJA69yYX7QsWGnmOj3e9123zrigU4JCJq/t3NT70
zSdAT87Rep9o8UXT1vvC+OnMMqgE7HWeYDZyMDPIoqRTQq3VzoUO3phpnLsI
kE7j9fJ2iAeXm6t4LJE3HnhhzeSCni8ntyREEE0bhxfIWoRSKgWPNYotkoNc
ITg9lwbph2gVhQsTwFfQH0Or5Zbhs8DQyrqU3yhfdYz6zeupLMDvFO+9WyzW
KBhZiJ6liGJgAwntUAIzm2zVX10jWI57HoCDOHsw8+77OnwcfC1caiKRjlH1
2DhIOtQgBtyAktmcBoh4UGC8+iqfcDQKYfU3zK149kKgUGBY01KVtJzJ6gmI
IX7duZejqAfaLXpw1wZ6lnMwtsfuQUe4JZoJfjJPEao52KvGhHCzaAZ6ilB6
j9v//yN2BGcdSQWLsuhGUdf7aj06mhT6xUJAcS5BbcTDHGHLPHfY0CB5w35U
RboU5xfWvMup73lK3WnJGOmtEFvFaFAX4SQNk6ZB7R1bQ46/uJNoJpNvP3mp
70UBh4PW2BGCdDxL4HIYOsOj7e59YqIrLsgb2nC2icLVhjl3/D3yMx+IUJLp
3b+MGdKY1DEVnEanNKu6H5d0J4QTdOJygvoHBp9iOHG8TQ7deZL8QRyDK8l8
CvJA8+5FuZYidxKQuwkL8Vq44+oiYndFL9nINB0iIrOxMyo+cW/3GCbZOmvA
4Qaxc8ijVbCzpnBAydSTv1wQbxZTqkg5dGWQ7HZanp90sTBgjs9Ax2PRjjJq
MfzvV4nGrEuy+31tgADbD3gqfXRW2LsVOTNzIAMq6WCucMHW7Dcfs3wIrJq/
K0keOOa26HUindnInjX7uEsE5QrEIKR9pxvwoZoZu5hV7Jt0cTqp7TGYSjPP
8ioYdyle3PGsxgBrbmWqXwHFc2dz6Q//VqcWmUTzp59wS30yJ25aPI7Z7tow
g0y0icIv0/nhfwra7346qWges578R09O/L6Ue0ua+pyW+XQx63/A0PnC+/lP
5xFx6CiOurpukycecCozNQ5Z/JyGN56DlzThMoZpj+abFieRrcrcyA4lAM8P
HWUAJ4cUpHt9xM3v+E1HHrUYXk2TRjoOtyv84C2WgeV4FhOcyRyWDnFQD7l+
AmHeSDN251nPOuPB2Q0EQkmLfGgP4bPV27nDGI8pMdrAMfc75ZbHyISNqPBM
mx45K52nL/U8HnFVoj8e+2pGMr6EYZjO0zyiXXT8jk5OHUFHTdNg39nbDkua
CSv8yxFcCT8oDAoxXYQv4JMduaS2BjU+WJnzCRh2YlpRjEotJEMrYPw5yt4g
cG1wY1G5aMpkUSCKmIzYkxByurhzRgj0ycostMhcn3PaxrpMYSKv7I//Xmjh
Vv63DYq5mI9Qf7bsc4/fyooMPM6zQevZ4QGhOxN7CUXFb/fV3j4w/Q9G6tJ0
YbMhfo0DJU7UoyUZQrrHwc7qMNxahtm5oQuo/QhnZxjuZw3lX5F4QRpCFv7T
uWFszTYzxHRf8PZ+acPygKuwDlDDVY+MgijgXbDB7vqx7l9sj7txQvp9+uNU
KPT0+5A5J4eB2XFy8AcV9cuSVciVJZ3ZUf/6lc8P9LskkptIMSxuL6mKWiFc
4qDuBG6Kxx/CUCdoYTKSDGXfp3il9uHZ2294W5BJVHxVCl5i2RO5VnLoNsA5
tz1WNw1ewD7EPOAH+H+zH9Vph6fWANh7Q+SwWj7v3C9T5dSGnGaf8Iq7pQMb
6FwOC5Kg2U9+1zRNL1kouc2kZhmVpr9qH+/GzRYceslD5Gxw3dNuld+3fI4t
WhWmnw7RBs/WXG/yFUXi5WQ+mYFqLbihY/2j3Sb5qPc2ys1JrJDjFgf6ojoZ
gKQRsVhCWO06pGyxaVLc0/Hf8aEL/qzMpqKKobavQoHTllZvlb5P3aea7Ad3
WHYSmkjYaQKi2AeSFBFcNNsthWeEw1zNItacKSeOLyaep7z8CGnGzd6DknUX
NZ2CxjrcBRas5+fRL7sugKRQgWGc+1Dl8BaJQN4vw02nK+A3eji1vHLYAhae
PKnMzx7dnRbTrm3G/nK3LB07lkqPXvywxAxnIHQ8nBhrn/yxbtGoUM4P2NIj
55BxatroXhaj7ZwZExqZGRxrou791ONYCIMExPOh39dq73FmUhzjIqX89Qd3
SOMZhFBPFP20b4Z5TGs0ITJ8tUSd3CVXX9cHlp0ZOEbRb4Al6X3JZM0sO5z7
Dx8XZunG6Eej9fmBEnMGmqrposBL6/bOUEWDGiGNeE80+J5R/ArVARWRXcrN
cDVWYjesKOo/+cX3Fl/J2iCO4gwJ6b5DhHlVmWuFD5qmyYOgYoPMvoRdSYQZ
cSOtXfxwVSO+NXTFe5KnfVPgNpO9J7vIvipNrElejLxVKXgdJaRe+5K9spHo
7K1iNZtfvMRwoZEB/rP3iW20fIWQhT1SQloYhm1+51HW4pXbx1NgzQtuBbLn
8J1NB64dC0p4WKRVNXq8ilISqB2iGVzGhyO4kvADf/aidBmF7pDjkcSKuFLm
HPIWntyY94VJPT7k+5K5j7kjSNNb8KXChuK+RiCaHUXwlob/rhzIa6hw7BQ4
koQhnXi1cTds5cFI0pByf6139AkbmRh/eNE9ikh6bqFwqbVv8lHvObl+47Bd
04eGcaFHwfpmGw5CRrq7toG8/bHwizm23Snwn2mk01jRjK7U/Lgbgy7BJbds
lWIQwtoZtrK9wFp2Xj0QI3X8jI6O/NmZHMehkTJXSiGM/1Qt0TllP9mjVjEl
RdnVCKgoc2tTDPf8t3364Jqlul5fiAXvOvCfm8/GglbzmjeMT//RmGLJOPh4
sqzPmuIWAleoXrMYettTtVOKjkHc0zyn3tpkJnZ7/zTCJgEbG1SGKtRKQuhi
wGsJ9QQXljbCzSSuWZmX1nO6XF8lR7F0JHJcPcKrW0HEnHsMTytS/WPgByA4
4eh+teYzAvhcDIeZwdGVKUuaJt9gSnvShJBwVJzAWx0OdhXpCy4w0KkORMRK
f1kWMi5BLnfM2mYktc/qo/jnORJr4rTwbqiK1YS+ZromHCCVgWV8B97iZCF+
XkYHgWcvCttje+IjFIfSnKXONOkZkD08qBmWMQrB3RtbZYhWOWX4HZ2B7svY
CAohE4VP33Bj/p3F4o6zDAm0UnNf9LfMgcXJuXIHmwnIQjX0wslDU1ozJ87N
C++dXUKwRs5nTbe16yg7UgaOo3rl0m8mEvRKxJX1lyHfEyqMKEEiQiqFJ48u
khiOn08o/fYi6Re4Fhd1M8eInN0XnEIa3/B9L1MWsjRpqOhq03ht75e/a6SY
qO8MKhEuKBVq20UReujFKx3DsE9SVE8adBLL/8luV21wmpcqImi1MJwwptvf
DcPmLWqBq4fiHQQNLUWMYDysv0MAOjs64nhU0QsLwK1RJiJfiN9PYfotj//n
OeFJWVD+JEl8iTSEz5koQkRw+u77MKXJ7zRfqNBbUv1oeF8fI6V1kexgzv+S
jMoEPtPa96NvOcbLjkERRH1uUgzaNvY/euNH20Dz4oF+uNdeURz/+aUtuyQ+
ANkMNFQXPhCDe69ok4gOwVdEQpmOKqKX+mQvzRZsi+ayN6yXTtTUBqeFAO/a
GbaI65LOunTkluWhG1PqYkj4G4XepFfH7bt1+KgVhvFaeYXFifa6kWiEqjLp
pcLCux+FGz9XwvZMlbiMbtZpq3WFyEPD3wSTvgspqobh5z4SO0+O6E+mXXAX
oCeEYgLxeYevyjlxBL6xQG9JhyQzgGGi2GQgbZWMEogLQg71oNAOTI+vCZVn
jJ+X3An/nYzm5V5OqbVvfdH5VnUm1GqSrfCxW3m7PKx5+m1q+er1VbYgjHzl
6+3TENOS4MhYpV9O7+Mm0uktkTnnawE37wg8M/nRJEh0u549PoIWzX+sr53k
VwEPVBq6r/OSIbQnuN8Z/Kb6wQfDWy9WJPOhv+E3O4662bvN1PhEGyRdto8+
wjcDgMoeurKR2Qkk41W7mqJNZKlQfegHMftJkNYjwxBhhnXjQtMu12xJqtw1
/aq7K7n/nEMOi6EJrAW/9YSMTfHnkQJJ/18FHy5nlqSeJAVdfzo9xugZ33Wz
8xR2tLxKAE8B2xFR2aF1/XJdAgeUsx7/Lm6AIYQZ1jwY7/qVfX/CSkLV8CzK
TzBsF6I3byFM0LEBhIW0Ba6+/oEMXr/RCZ9RIXCaViVxz3v0o+RFTWUv7ijd
xGtftEIjsJ3uZWBf2kDmjUMNHmmzUSw7sa6QKLsNBpMjwkQGBDgCQ4LH/PuV
qvHLtlr3cYw5j5x0Kg6PotSLd9S0IEODgcK6YkZLHS1FAtITpyXj9kpLCSqb
uSKUD9ls63KkuAx90adyLvoTvo7ndx9a0mKChNosDwZ+PmJCdL/sCVWn37r5
hxKEnzjPdKzbmyfY5LKcbP8nGewwXH+0x0W57pGl5xEp6t8zv0h3iPyaHHt4
xXFQKzqo6+IjdPnqqiyckFi/90b0iYTMS4lv3ax0KcKgd3cIykFoC1vST08/
UImMZtk774oGmWWpctxXkHmW1Nw92KeYWbyPfnq/7D6L4sENvIeLx9mtogE+
yM8RQGaj+XFa8rVrE9uNysomlkt5iwi0q7KwY4FyqlDPbRpbpCeoaQ0sRNHD
OpMfeuGTNRLxKVXIZMPFcRFAttwpXbmljZ6H7QI44oOFPwR/owqOeCT809c/
UOQ7KpjRtcnvPmEap7gIRMh4QvixrinDjOBxKRuTmP6GlKqFErnu2bGvvOZB
CjOeoerbfvHXhozAoY9UUytytiZ9aMktnd6N9PUIdl1zD5DEjz8MvJpDr0iF
hSEVp2uwPO4hplWO8oDJg9216l/kBCtt3CbkS6RY4fbTyhFY6ndQmEwATxzf
h/j7VRYEL1bcIGbzdk4ua5zNhJHbWxHA7p7j82a/9QW5nIr/9zzpj/d6KrhL
OOAkOOOzO/itJwNY6h8DWFjNJEJrYyR6BY4SYGMaCIjgw4VUKJ5Eiihq85k2
Yyse86Wh3Izejjvx2G/DikX6uLfVZpCF5lWpORpKD9hRm0QTQQNlWlpLafWj
Gizpja294SE/g/+cx4JxHJYIpN8Q7NfySZufDbwZWQg1eS/CNRHTkxaGYKLV
OpNiFbDVsm/XrFvLArNmSLHLJ9w6qUQ3VBoMxNWkAuAWvKEEO28m2sob2dhS
na6uLSplHOc11iYRVwc5+YjuCVfTzW0p3k88i12OGlJ27HXWA3N1Se39/6l5
lz+7ru3hw1EK7p1Q3ehp5Cs7t8hfTHOUitQ2PjW+aIks31SM8J86jBUREncC
t0fCTrxVyF9nJvD4jVonn5OrJ0E4Mci5c0y27GZBBHHDqVmgGblBQelVxUgy
13end6ur3YCJ/Gm52d47meXophPmJGu0vZPNTycy0dk24gg0Eluva6dzIBXd
ifX66JzDxoDENZZ++PS6z5jDtrvAr+dGx4vFbnWWKWf1mt9EGWUNe7x3uApl
38Rta4pxlkLNAr+BqVaa5AS51p/Ivu2HRmju5EvSSCqhxGu4Ya1qr0F8JCHy
/1rMwafwyjivrk/qAbLQVINjdN/YjGYzXpo4MnD8+isByHz9IcfDht1xzAhM
U472BCfUQQR122xhIfBuBju6uhAKv53c3mbY75h9VGVlT6ehKGVs9hnopKOJ
vAmmPZANW4/LFcBTdcj6UR9Pbcgj2PJwYH16Ok5f/I1XnEUSDlxmnumGxhHS
PvNLrYUY+1B6PF6+Jl10EatsT7XYbRFXgBPCoBYK/P3i8bqlk6UaUdDwgq9N
1rqwd0GSgpk1SGMw6ryOndynJzzARAJRxGnhJ2Ft8JaG5psvf+hQROM9btgY
VtFJFgLDIgI6CaogEy8mxtP5USINx1wwRt3PXcGUyi2RmTzO03432j79NAxp
wV2tWRfjZYz2fbvKNsf/Y7gI5O6F/GTgGKz3IRJzC2m1cm9IHTY89HIZ5sgS
dKz8DqMTEWvi/jQz3bsLGpUxZLA1j+4aFTat6ttArQ4jgnhfLon14KIEHK7w
JpmS0N5JcNvSaEVBJWuIW9Vkhd+J+iVZOBlK9pXC2hbJafBx2TpVxXzS3ByZ
hHWfbvg+2Zs5cdYfmARr1lEQ50Nh1iih2ZrQYYHs4hS+pcgf+mlByTB8nQop
wHae+EcDuPH/qdMe1/EiUnAVjVSg6fwD0nhP40ma9SfgWeZGvjkAeRI4JpgO
VI7VBuMXydcmZSenw3LnSV0egjzSsv5uIj9VrOoMNffs6F4ZvMVOLIBmQiZc
gTtBD9Z7osD2BBOim//cn7oYB+ixu8zfEup/0GgDs7R506nt1PaHqVq/kbbw
gZ/8DRkPjgdbzTAJpFTs4HTlGI0YNCeVQhqoCcz4x8kJ1XP91QKOzWK4aN5E
Zn/vvA3aJBHz+dAyfc0Wlw3CEK9CR+0i/PEe5qGvHvZZPyOWhPzq3mBF1WEp
uz5M1qoBiAog6YQ3J/st6heT1Bxo9+mAVehikrH/ZeNsq9ZncZ8cNBBnxpkG
J+J0W638FmeQR+P0DBsGHF3KIalxEHugQPhlwIeiAFS1IAikwlQiQwQdhdgl
4mMV6v2eOPsBwlAAIcrHhbjO0l2H44Bt0JgG0HrNZD2fiB4miXcnxn1t7uWn
bnyYQ2cOtNynsl/JXLXs/+ghUCgcsYatgAO9RIZ5z95WxqL2STv4Yf7esyR2
z8rRQgGy4oFI6YneIINUKiLdGSTUTmTgziaynhuBMe7IGY8MS7ECdvgLQnhY
BZTAsjdnSiRMYZ6+EbI2WprjaXj3LVWplqNhCKXd7TKIA9Ub2djGvF+dRiqe
Ib1N2aMOF85wZO1q+fzJfbdNEHfswMmYo0YRVXjjrlY2CwIvzWqVZz4WnYTI
A8Qkt5d7QNusR4rYebny674AT6/h07W+AHqayA3nvG3IXcNSkbouCticqpeh
4YEw0jbMRsP6zLwUqq9lzGTWc7j9L7g6wQEnP0aqViF/IJbl1NMxuoFindyV
jtPR0IOTUAX/H2WLUBFxR8hVsUKwiF1Ixra3Nk9pq6vG9L5zKbNtIkdCmT6h
YXgjSwsROv5c0DR1xlf09WRmPygjhnBAuCGSxV1V2o2DthvVKnMs21HLe7sZ
+2YGAXNQTzT7I/0SpGS5qT7FR1XQneWAtC7KWsYh8HudQnjSRZFxJiaL2Q8g
7i/zBzYrD0fj/ONgZNugrOVdjXNlYRoEkAeV4yCvR5qz4rKtOJWqYYwk0qVy
7PkkrBKCtlhc4Ru505Q7oYpJ8UOSRROxP6fEALa1i3raG4CFxQ0tgq+5FgDY
oBFEjVw8JYgxlBu6cyo3IO8MPOQhhNpVV2QQEuMw1FfCzZ3rtAeHt3XiGkzd
FSfmELAPK+95q0Z5/q0MPoh7fVXO1FRmB3cMkUs3EmvsHbhzPxEXxY3AYHra
FL8gwqlPAkve7XAQCmU0a4ecfdHKyq25HMRovztC799cROKJ/KsBM8O/E82N
HGa6ro2NcerSZx0OW7gMeAQUQ9tgwwqp/8Zhp0y0oKYfk56YA8Ez7UEr8v7T
/JKiTixb7UEhtdwVzMRSuEWfyeyYEawNRhnPubnIQ4R072c1+xTnUF40bB+S
wha8sKfy5vdMnwFTlw9vJk8l7/ZfDMjDdmSsNtnpd64QQWGgjRFYhM0Xl8y0
d3KAboZFnsYIwzFw/NtVZ8wjXudM27NX5VNMKX/yiovEWC+L5zvrvezCy71U
smqZaDO7WmuvqOv2lSoQsOa1KNUTpd8oe0rKYIYzT66jXnEHL4eqZAIXiXnJ
P63M31D+CXI6jmxvouAv309nWt5Pu+PU0wnl15UO6sPj+05OVIFTj2lxxMNx
2LiUZM7j7eE/nC0oncoL4Xz1tr1Isuf580qh6z3OnNOoBv9IhxbAKISpFOJg
fhHxmcnumYNMQn6rMB/1YXsO7dpHL+7j7jyC16LNF0sC/XdeL/ElAvYhQVwk
vzygyvMP3bvnI3Wu368Uzo47Jkr//d+cT9ZxA7PmGEHADCAJ/BX1zVE7z5eb
bTy+XSmK9z5cELjnofTq7O4tpoIfE+xuYGvRi2+C3S5dMDGdKDt/c7C870vZ
k7V3nmDKT1GY31iaf7atN1K4p94lBdZtSz4k5y2EQVReS2DID9AtloHoksqv
++MVNDERgi+r06lQ1SuWOFn3ps7BFDQp545y/oIZZ3OQWElWc49gBBdEG0Xc
hxhKywemCoipSzckwFjDjkAbgc99G452eoy46goTv+UP6ZYe01PUbVljbLfy
pCMxF5qdYr22qWhSVc03h4iWMnYst/p+ky3S82Uu5/RLBO1TH3ld+psdDBf7
6se2nHdsZ3o1OhHOYmDGqzIqrheSWFNT62ky6vOAlmCYE4Y1yXzRSfiN/ymX
+5EwLGA46xAK9AxYlg8v3jlK5NIjNGz4vkCokJ1L9gtI27dVq075nAxbzLjK
JHdk5gsyziVBcyMHXL7Ltp70ZSQ4TR1Rgj5eX9Xt3bWyDesko+d4Y5AWA5te
KUePMJzFjIPiXNedV3lQ8SH0RW0bynq16hH1aeLyQxZirs9BX30jYJIeC24z
DmO7YPXccCrGQQwcG+47rFIKrlDyA7xi9XS77nZRBEsiKxo1Y6kpfKl2ASHj
norNelqqkhidscsz5BxXc5R+9ETMTDMABcHULX5S/4dzDA2QIgNblH8iDSZ4
dc0rANMjgTtlhkucsRke9cihGKvSe+HQXQwtno9wkAz19ulXKL5yj9fHAzks
HgbOLBufDvZu7MOGzOoqU/ujV5KDW948YwluVhXFsS+6o5yK1RM2jdYsRRNO
mw95GvYvOCVgLdgyeRAvCJVWyK6o3HjCworkH5/SIpzgTqZKpw1ts+/3jOqt
9Q1DR8XnjIUZvDgrqmdj2ss/oexTPh7/yK/+JrhYP66JeQc5nzZ6r3PGWQVH
okNVJgsSh4AIwypw5bf2dKTt/kUtJr7Q2uDW8iBMesYw/ccagPxQlrC3vhsG
g54wXfpiS8e2s2PZbUqe9SM8CGjpHfqwvko6tfwr9ueNNrskgCSaEBXHUuT5
YuJirk/lAlwE7Sk7I6kyzAC58YUcvCV29Vwd7Sta3Idyr0tQnYHfe3ulkMeL
ZRMUzcd9Hfrr6ThHMrCk5EYnyHvi/wcy7ID0MxWV1SLbEPN626oXcdn4bWV3
TPiSxNVHKXtzlNejRonhKZ51TGlHSFYjWx3KDzo94JI+3ZaYCkpViSNCQdAd
cd8G+qCXLBAdTWu9NhgR/h/48jctTszJSE0oL3mruT/gaut93MQ8zO+In81o
Hy6zxkmwIaBmhAiKztBJJfqA//9EZFQW+9dCpkiftEAO1Ny4C/8pZy2jCo2U
8xgeGToC6WNvM4ssKn1ImNiJcLBwxrESCXKtr4cS7iFFCOnxsiy3OVreaBQu
5Trt1D4SPf94XcMWFX0WePSkK541U0jaWm6lDFApULOQ/uczjBWk5n2hMmbO
VzRFXDdJkvDVLbByLce+USGbt1aP8AFW7kptx8MwBl/tUAecXpOYIf4LoFGz
pwnh7Zsr+kCbSgcvXSkRXzUXhDgcuJMtfYkw6qp2u3waedkotpkxu3MQrgeQ
i6mbb6Ns3+elO8mzznZ9XkyjLn6afgchMgFHFU8Ofeemb2/sPrc0/m70FTty
+uzDgWx9QgwynYr2nilg/3I7XX4Uni2t16C/SAxouuC0YfWPim4X24FherYm
xK9Y6Qx5yryYgcJXCVzszRSp5UUGTDjJqYEgNrQ84I3reenmvDV2l//qoHAS
Ceb09nUZjajs3RFnXb2S7BKp+ulGa75txhuYX+te2dLmuhjyGFCEsOOHAfOT
Aavv8pe+s1DBW+NpBDpV1lU+y1/G/Lqu910DzOEPt6gs0Vnhf5h00jVJ+96e
KwzbxRkoCBzF+SRn8Xr+qNmiP8E5uFS1V1vZk0dPaexmQFyBcDa2z0BMjqNq
4n2gaEJq/ZgXcegFDIjVvqfQMIyx3q7jw85ip6dhTfmGpHvSaf7RvKBWOs9s
DDp8FHgE98Kku/10l4pxJriZI5Yf1AX/brztK7mkIoI/6N4PDJIRvLloSh8j
+nqVdHRuRX3RqbqRNJjW/YMllBbDRMn8nLIyZfslSt7LsUzuzp52BXtNJ6db
NByAdXDtVYLS+vgt/L4LXfSCZh3Mb4BO0Ucsam8p7/YUkWKhRYN88cTB9nSk
RqudU8waq13kO66D2So0dfuHcTPe8g4ymK2LiyAlOrOc4TeHNofk9yTIZ6OP
LOVsqo2vGtCFCBLMGC0UpI3TEkZSb19GC706B8FfdEdcJ08JIzS0kFhmcvD3
mErDMr8iMS/jP4bHF36mvMQidXQKU3pSHuAsURKBlpr83KuHv2dQzm0DXFHF
hdiis73GeUt09Yertpd1ZaTuah8TWpSgXW0puFqSZETXJTSQl18aW0rajJqg
b+oobkb9eNJZPvOHmIcV0O9T+tFJmEr7mDJlQ9hOjBEra0BE83vthTxfeKsG
P5zKJroayf1FtudYH0CFX1e8gRjaAe+TdtXuv+tgDr7K5+4AQidr+Zo0IFr0
A1vPK7AIc0eHZhlOIivAO4lHDKJL/2GRV1kUeM7xZ/sKKd7ODMy73POw7Osg
pypfvBjNFF9BIiJMsyksJP2Jid1rK/IIwWjRYPyGQh6CjQCXh8LpRypRuO9V
ChMBDnDCq9NhObvspkP7ZHBDl2NeeazB+HLham4OX1qvGJp9HPv4oXmUu31B
Rm1Gfznu5oozpYWK+L3nk+f06by+trsg0xj6bjb2kGIHkktZsfBAqogTv5SQ
xpeVaztb7UEBhTrelIFSS71j6+KAd6wdg6EFVGryGtJw2fWhNV0ej09Elqq+
SUmrvqUIGExFzKVQgOlRXbqk/fw4kpIEdKTIDuH1Gx4ZIYBRMrNcRY2bldPr
A3fKAi71M7dS10HgGBZ+sqIK2jzUXe68JSnykzE6UTSFvzICm4j/6L41XfQA
3SSfoi5OVhHLbwPdkEoXbI7WN7l2Yn8Z89o7Be1AhI6jAO6TX5tTUbM8rnxl
xpEdPCpKX+NRAY0bszuXftPdsCN/zAnq1Hdn2sJQId8LAkS9StUoq4NnPw97
ODnm+rdg0ZDrbOM1V35zo/9sw38seAKizwpJotTAMjYSFkdXtyFCW/PbNBko
Pni8Lhc5Pr/YTi1i4j65RcLowpUn2WwGB7idI7ynrRxbDiXVx9Pm+TCWhU8L
kePN8SiNxxzTGWzVf/2zV+HTqzEj3oZ8kqJ+GVDR9JXK9AvrFAynkDGz0NxY
IWI6woJX9xWRwnEMmjJsDU1f7JkoUmQ9UCQmDbVCW9IrzPFxN7/NUxt0eER1
RvhAHEtNfy0dQZRVoFwWb5FUBaz01lgGBU2z+SOKYjuCsOsIgGXdFZDZqxeD
Zpee+zKDdao3YhUMpmloO/vYYPHI2S5EzaNswLYSjN0zBEn430NjSqQVVxDl
zUgsJ9mjxF2P4N2xo16h3a0clQekjhSIZgqkugR/5+mK+NgzuWaVcWvPMnqJ
RdCnGino4YNohgAPuHwbBeLgQ52dloOw/VExU1nAAO93+K3f+GnzSmna++ci
RXXk7yajfS5BiKWgrPuqygX+y3WUrC6kL3oL1GwUTnILcvI+26szCbM52/bY
Tj4aZ8kWCAa0JotsCzbdE3B/qnuhM0HpD6qsSdBD9Pl93UU8v5lxF+6BtkeM
we3EaA4ak99ImlfT42kXe6xldKhPUbPT9R1UzD2R8q8ShfkEdapHhDXYK2uM
MuIYuxnR2swrl8xvgGAUa1dMbMzAsao2uY1a8JGd7gQDUCKKeO/HQyYHdQAM
2f46A5yuvojrb24BkE1Juxwulz7Zme/WMdVtVQ+sKx0fqhiRT8V8HoPnuZQ7
HGfQsNOr3W88LXoBh3j61Tmmjcog7llyA/+Bnco0++63ORb1anI2wRYVPiOA
3HQZUq2DBIAOilqkDb75JB9Fcbh8OAiN+1/VY4C4MWawVYPEaftjgCiPu0MH
oM4s6V9rENdWKtLBFHjLffmbpDRFqpI0N+UX+NOL5VHaDm/DfxdEhSxgjX3f
wzSD1+Ek41g2p86fp+y5AjHUWg1/Iol4l4McG4vxDGq0tGD3F/m2DCzmrGjo
C5F8GrGAV93BCeoIqoVwVPz+/kyxHLiNEFXvL79bskHkigudbSYj9ATrrHOO
m6iu1Xd1ZMRqIjRuARuIZ0fZoUOgolCbHMfmB13VCyn5dQwjtoGt3zN6aJTo
o2MaRZK/lD1uZcv3UR2FEO32pwGdfIu1a8DTRIm2FiKgcbCuvKxbbgUsUl+z
YtmrQvJka6hBOpP0dklwUxzoKfccLWjkOGyTtsER86OTDVTtJq2x0XO7a0BK
bVfUkfikZKMSJCkqtvQLDGVnO5N012hki/eyPM4hDrxHhx0WM7LisW4Iim7y
oU/UZQkqzwbZkbPpgJoJ9gaxsJbv7vUVYuyK9g2NjR6qUdZ5pPfj5uwQyNTH
nZczmVzwmSI4lyIL44NVmitJj72ApVhaC4L6tsw1svHGt9oonalRYTH/tDB8
6fsYM+4YUd95QA/RcmbH2FKhRkbpiGQtw8pQeLgXdmUGq3EbvFmeiRPINMBm
/wnG0oHrgN2ZmSUwMVKI/HmuLIcupkMPWfzBkPBFoH9NPyrGJTDdRgQRKMfq
GgS+IKyiG9hIJOraSQHxaDQjAKLvIVJsdnD7qi/icic8RYUIlzk9N8R7CwAt
YfQZL6mvAqc3TDzzjfvnmC/8hDRiUHlilGAA5RCu1yMQpp7GUaPVie6/o+eL
3+yJjbz7bm6MPB9yf3AF2G5j4Li2oewkGOwj7hRYd2VEuzXu6hUZp6NZ2dMj
Bf221aUlS5CaWypDvwRIZWQVFgQttn2jd75Li4B4oLc+yRRF3a1DjmdNVpvX
rT6ZcjtyCInqrCdehwGwZsu2hv14pF6agJJ6UNtVrjSp/YKCTu4AhIyz+AA5
duRXWfrvrFax9RZr8ftdzPH7O1s9mh7uX/F5R0fvfhBkZy035t/kvmXYaDU0
bI19/hoVXKfZ3iQWbVva2EXAdaSPabMnYFUhFx0mvfvOmQNMlrjTU1I1NFLF
y226lMUgeV0wxHD+9Jb4A36HwSN7C08jE1b5dMJgpyIvI1+4vpkXTif5449E
E31ZeeRxlyQj2uy7MZNXHsWvCk8wfRC3S97BCvXBJ7oCix5Q4cJC0a4+zWPw
WAstdt70cMdzTbscX10vnSS1ETna5nnTw0Nw6hQcGYlbZ/rnREvTxW6icnPe
i1xcqzof+qe4WlY9zb9X9yXR2V0vHd1dnYLLyYIOUCehoIv5oCPxUYmbtUlt
Ne7w84S3NDwxvq9CbpzejEgeOn00YA5H7KLDmRS6ojIzmago4TPnU1NuqEY1
Tx/Zijtn5HVi5yOiaBE3G170Mn+VdU9MeP33oBqoZnFLMfD4DMoG0MdvpvE3
9Zi8y3PirrXX1sBkT9KtoTUsj/rTqZndyd4vB3r/vqZ3hpieFxe0kzIDK09J
j/8IVcKPgY2Z7CrJZvhjrA/Td1QC7GLcxAMd/1w2PgtuODgXH4AWkweDV0R1
Jj9aPoJjdgVRIa6/42SOlMqaYbPrfWclMAnRTBUGvrscVlX8aQe2Xr+usbQk
/sTVGe0TwaL3Fg3BiWiVAnyKS6qrRWtBTL8Q7k4Lp0P5YopHFAqmATQI/Kn8
FtTqiPFwoJTXnmY5jcpDgtLiGZ55teJoKOGYSa6MVMD5/rJFBzuPuYQ41cCd
qBjhK18Z2M5ND3ucSit4y1gQiLzi9MrTXcwvYLCITgyiMhBs6Nc2iQbGux6a
gWbu9ee8r5K6I8BaVlVXrh/8RCKaQAANLyLPQwqbztJvLwnfWEp4cvPlD6eY
+bt6qaQJZgDMx/CxvvxDSbFkuH/n4SNtGe4Qq1P4AiwB4QC/3upAoDkPGIUX
jNmA/qrzqqnptyGqB2PRONuLOMfqTZa+PaqM9XDgz3pZQ+n8OxdJS17a5doR
yBVbFyjDFI5JOa79Oc2LnxHqBe9d4Fc1WeeiNx0HzNCwCLxnpCrAUAQexyyN
wKmstteQkkINdagVKWNKGWOOOkR0yvTGydLCsEV0W8y4dnuhhmZs+a/8v186
1qVUXm0lsCZlPkeruRnmhRAm3mcTNWqlAyXKlxTsfN/pKC3vIOT1bFQM1aoI
2GVxv8W8hiZyfzLLQ1sL3t7ZQfbszUi5Oo3/dEfDNApJ6sSKK+5pyVFNfN7e
TuIttNlXol8g/zZWiNmLIxAdnaA9ZG+3hSMvxROCCyhvSmvkyKFAU0/6adSO
jrvTjYuMtvGYXuNx7qGfySaKvs0AfVNBEoDzQMKCtS6N6bE+TmCkVYS77Jbi
SJlqxx/ocGfyV8bzOfXrbxpL44TNU0ix5HX24HTroDJCU+EPAZkr7RPd70QM
NXTqAKkaKYYBrJqqsvdCYq1jTspqtYG3TuxtI1d7iJDYFmP1HAvzPUCD6DGx
4l4NV5zmZiB1BZ9hoWOgDinusWgxP5zUuGfIQCtQOezDO1QMGcoJdy3VUs6D
waWpsOcgUvNv24lZ0osrJX4x7G/rqmh+aFzlj4xAMCCs+hzGXXJAje5h7oHN
MrJ2ECGOck41i5hFeQjYnxU+z4XFmooea6cfBBCmvJLU4kZjHjc73PLCuDQv
dpLI4c950teFmK5GQg+RI3p7k4JGyPpJaW9+E+HdAyhXSOu0bVp4TOYi5ovU
E7HlegD4VB8KCBGbWML479wZkdQb6M8eQhoYy/bfnProuJ2Fzx7s94Owl1G4
j8a8mx54A9z1DfQytPIxE+XsUm0Naw2wKN593WX/azWKIpbaluRAMx0FSjMp
KszMiAPTMX596yvQ2p/BgvBYgpMJGKDtYJJRNmNBhgp0cGsp+PsmYq5ovqlS
+1kiIzZCS3qEoorz/Mj32eUiPnkaRzOzwoZ1EByfjva3gM6thCh5pm2P8KVp
E7TlDjZhAmJj98aNygaFA3UTyeri6cbnpx6YgL3wKBlTyPfFKYkl0L9Zra0A
PJkruc4JCnS8ydUIW4jL5ilrIjCUtNy83okarqdPrWqv8QdS+sc1jIl6SeI6
FD3H5FC85wcIReJmRA1mO7wTsfRsfmS6g5yZcT1ZrvvrbRMhc53reJ93pcnP
aREXzMfaYKz/moeANUkuGNsQDmhVSUWnYrDjQRK0RrLoVRhAVR+wuDe5YSR6
pTt0WsaOQ7JHCg0pQnCPeR6GYGMappx3vn4NLDxm+txp1X3WRRSExJP71Egl
OSbKISCOIGjWEe9NhNCiZMgiSfum7OUxPN5kpxs61d1odU5Q+br8WRGZS7aq
6h9/Xp7+intNAiLQfGGn2hS7+8Azp6hqca+oZD9ADuAQbNtpXrA+se4sZZ5I
JWOnLoWXcymhYZVwyzkuDXmW21kx4hv71oFIRhVdsyLAqKiQ4ge0LExwjcw3
t2nK+L1gSLlwcIJ9jcFgOMouGJArZFuOOZ+24Vl+WmCh9kmBJWQEGVIkAKIU
BhTur0fZoHwqIOj9KPWEuOn+ED5ZDcFhXZPYDr468FvCFUh8qPOZQRet9wOd
kcvqw3fuEMJyaLItk5nQI1fEb5+qhbwmJnwHUs49ZWi1YhY0mqYnCUry5jVg
oD39Nl80Nr50cqMK4zVYIdpMldmX4zsq6hEVh3g0DfJefn44qdpKEBXQXbNy
Os7A5BEZsuV68icXV0NfB9+D6CRbzscH/ibpZBiILU+jjYGyHStq8vAPGkBS
/ztv03JCu2A35FPx1u2BUxZJsb1LWrwprR2Wh+aJhky73zOf+9Nn3s2XK8CF
7V5SVPjXaNVfrQw93LDl/gdvb4zb4ER6LHPgua5F6jRw/c5MHDLi7mL5sSTH
VdVQl18FdypcIQwPrtAy1bj2GNb7/+QWoUyqehtGRFnHyFBUnfiB3EMUFyeC
uSIuE2odvJ/kzFqO/P2NpSDNOKk0j6tuRfpYnOBA3qRTlXIZiafahIXVDJRr
/FyPIqv6l48IGD3bvFUAIWJH/Mc5HiXctk29MiktHp1c2U7jAndi97jQBmbt
WwfaljVrAJ6dvEUH/ZajulROT174NJlWph29zW2zP7PsPQtJeoHnF+AXpwLD
b7EvGiHoxoX7UYIyuALEHqxqlnfeMTOA3iQgd6CckZb234AumAXrNKof9Fuv
5/CRZ063MXGiLlsYYvn6ICOIp72qA6u0eqBufEBiomzA00AeM0YlJv8MdgwI
ZBrXSGyM/XJcM4RK/FGVDiOMWjBUNP/l4Ti9mqXfcN7q+4eklwn1cN4BqYIy
FMlMt8gK6oS/hzOX9nL5ehQriAuSVWPqkZC5aPYzwqj8j9V8R27nWASbxN+Y
9tH+PfcFN88cemUNX25gt6z8ZHqrqSyRdpAQ2gQenyAQF1wxiEJdjuwyz+Hm
3npWIbTlu3W5GKzc5+TC1F2qPoQwfURmwY27NVQp3yNwPkcgRziUtPFMSbr2
ZsD+v1RfKWQoqI3EId2aBS+GNPO70TkVyZ3Bt1K6WJWTk6sJl1rdr+0IumRx
WXmgs1UGS3lpqvc4ibgBrvEXba3JQ7CCzgaumMu1SgaaX8Tp1PItC7C2cGOm
7bEqMyVhnM/HRJOr6syU98RbtrELthdFwsrra1FaPxe8HDKAWDZ3h6BHd7zA
79FHauS2907NZkCCHXTfhd0iHjH5SE/HkTg3DN8oIak3jd7F5zE9l64UuO+w
WwRmUdtG2uoho6W1oC7rC3KEAkUL99/J/Xu+CEg7rFvRIeMDv8qdHnUYRKKW
4FbSBXzKXgTVyzrqnpH8FTPDQqUJEj9ghejwZpS3bJbLvUxt/9AxLQvu/7EG
5dUgIsL71kMJubhUXIUDA9UI4nCe0Je6pFHOxqAiBeVMu7ulMAuiJcWLK50a
M4mqTl69N7kc3B1ucOTHnskcVbhJ0xZW0yYQb6r8temaUHBmdgX+GxiXZSbC
lfFaSXLC1M+rlbuBxDxiSfPp/VBo+bG9TkwL9lj8DNH0SvrFgn3D1AviHIjc
Qrpdi9q/BgH87pYXWy54qFbqh0sBofmMbzi+w29Py7yrhwRRBqDaKb6/YrqU
iQlvtgNEwrO/T6K2eum5OvzakmjGFF2y9r9fGY9SarRSn6d+kAU7GP5j1378
ZcZ0IZ7LCL2kBp0xMoHX8GU04rb8jd2RYqqU791nufEQN1jLuRKQsSU0Fh1P
dLVe46CJ+c/NIsq4n8YB6efNOyvbZ3YWMEkU/bIruTwjGOHy240PPko7vV9r
bt48kWnSn+hxvr/lmViYtxEWh7pUvghi1tOE8tCtYUwZ5v6rAGDhkEY7KAtk
WfsiRX+qzb9k3VKAHS/2gRfmVfuSzameFYj+c/Qpml4yA8Pz1QshE+tPY2mO
d1CYZ1qttyvljQP0h1QA6kvWQUYWGfTS0pB72CnttrZZvSsgTh5np4gaiYL2
CB4ga2FRMLKPej49mDcvzvrIE+Ghkgoiq/9y0/NEnySOqx29WNSVM++2c2uo
kT/aVEv0a3EzLFm0VT1TediP4fi2Nen7D9DCCo4te4CwwJHQIiNRaErb526m
oDxxuzICC5T4Q/KW04VWSRfb6jqr9Ncn7z4rZP4MarX9eHb7w5d/FxETNMwD
yhRsCq6jwj+YWFKGLd6kD+hhNr+dI0DPWsG36gGJUh+cazGnWwdQVupb5SNb
lZIJSsW1oegMI/tBEWAiQ9De/lvxSrc3Jb1U8mY+agmMN4IOUbeB5WbREvOD
VR0beKKbzTvLKEEfKlMoXpiEOMCIWN9vKxwAoww+s1YmUvv9Jt9x80bRJIIs
z0VXT0g83XJmhfrIFqqy/LwBR16benj/0BG8kYW/oem28sqJpbzbFG8ASUXv
Q37m7NW9ldZAoGAbBG8lh7QXA70LWLfvr0xfATRPmTWjioQMfrroThoQxoPu
3Zk0PDgNjY9xp+4NyJv9/RnbVaqKRo475curMVzaydVO2ro0UZGNsLQzqHDx
ehAxNfKRVhsiNpQ4GRVajOZR+9nLN6/Uvkxrap9L6ud4yZ8bcj6/MZVeG1Dy
7p0Fz3x33ciH3RUKF5SDW6zbgj7KtdHQUY7NV/j4eVSFKlVYc/EwHgihVDiY
TIdNrZQTYWteoVIvqsCFtl8Jhoj8vZXRpZJKeGUnar2rXeVrfhzlDUBAN/Dc
bXIQKuCFLtF3EtFh3wNXygVUP3xvg8RxHsbMQl4lmqFeOzYG3f9W7AKNalPu
gZerHudTa/GrO2B2ok65vQ/leAnqsva+dufr1dKNptSGaelNKGTu71u2QIzz
/Ckymxbk+dFGIsbXv6jSrEi2AOHEhnQIOZ8yo32zzn9aLFj8PQwXSAxQ9ZsB
iqVRqyqUaWPX3FwFMGlnmj46RHFU6aTpAi8gKfBFE+hRPRGrDzPHMK4uDVOL
AnhjkLvFhdA1SiSIwKLHJ55+P7MN7h9rMo8/HV3knyLMPHu/7Z/ctqBckEPF
EcwIcLqg7RKfOgK2SvVjXPHr+5QV4y0woGJwZE/lBAfZySjmkBkQNhLNTgVl
LS5RT+NCp2KD2cBs9n/wMEGvEBerSYN8mwneuN7waN8K+5j99POEVALad3HF
ZMdPr+ryVyfQ+xWfoGVRk3dU1VlYKPyX+JZ4ZmQPIt6R3B+ThLOxMIjvIW+t
B+UY34Dj/pWpmqpEAeaESJgrM1xR5qZyKGo6Ajujm2toDCcXed8O3pSknRRf
NbHLBD941SWlgyDGL8Sz4DNMm97AuWONJW5NCLLyPHQ6yvcWYCVgVehj689S
J/u/TwNIz0Mk4+u8tM1fd4ffspl80Vhof5W4YFD89j5ayTGwFd9o58VdiPQA
7Gx7fOeO8ofKt9wmzfmtF/TQ/RcyAoOKThgxTJc2THc1C7aTHVoarfoVycjy
tchE7vQJCSUXTVKdC+4whoSHD2dGz8JhJKGQbJNcrOQhIvGv9yBK0/XQBXPO
K1KJNIvF1xgkdSMlmMgmFoSHYZesa8yEWWYp1YwhwkF7+AFDK0VyV9z2gfqw
ZmiYYQQKfq30+AMkavsYQjOBtOdAoTLqhuHaGd9Gz9Yal3Utm+fKsWVuMZGJ
n02cnvkyfWau6geTMBHvsa1aDd5xLP+v0BRvUOJwLu2mXK5Gk9NIeIcEPLyq
8+Jx7q/7n9KRgFURcKLN6tytdXYL5Y5+tySiwsZgTs48H9n6un4DGsqz592K
jKYYG7l7KPmluGScfRufC8oKZBX7PFixUZfy6eYJL+jszYdTwqJMaXVZWvAN
pg3SaQxD6Ie4PcHC/yIHAGPaMfflwx9CrxGdE8Hico+DSx0SGmkxHO3PFZpO
adNlWh/Xc94/DeItUzbd4qww34pCegOAW3zuIriqDCyKqIL6SkkzHDG16own
13MptWD9E3FIb/y4AJycXO4VJRWi3050g+IhpAXvu/Uzu9f++nMbRLfZCmi3
4hQzSRm6k8o5eVsc1aHSZlxIPg4bEWAqKEmygwciPhGqHhPi2NeJM8utoJXL
wzBPhi2G+pxIQZqw/ZCfMO+cah/04tHKRxJeqy14ow6e7ltxbZMEs/817yrU
a7Z8STioL7Un85fMjqfyP0nwlgKPUPef+YztlsYaPaD7KvY7V6ZTO/yGMC4U
JiH5Um3PdORJnPSpnF42cI4UMgxZcHL1vARTjSB8K9McDs43Wu5ygpxD6Dch
J8aUUvN1Vvp4gMy0QmZtg3onlKpE6ZkDi3dXZBcwTDU0BnqGtOQ1WJoLbBLw
tBg1a9RLCc2qLxKQONp/qNmKMFQDHmCgo1upK9W0WDrAwxVymVwzJ2qK33iF
Us68aVEpNWkls5fKfa92czbr+qJjbkvxVJnsGfusbQ9HW3SWw5fn3SGJSmqZ
BLEbPfwdM40mnxg7UAVhlSPvidG0hbnNI5BtY7jLynaW+16tm4S0HudX/e1y
bOXVYXI5qAKHGFb6WuSx4xAcuh2/4lLe0ONMRETl0+6JXAa6lboBxyryiWB2
IaJHITyU09MrzxMLAY9AcxBOX0iRxf2rn09an8KSVlXooTlBzkXys2OECmDN
xCX7vjCTtST2xse9voSoKFTNTcHLz/PzcenbOaqdFx0tRZPDAzex4qyHpYzm
teGvG6XLMSU+W3SnxBSaULfbGJdM8A3D3wI43LcWAREgxsFzXAdJueJQKl5v
7MikimUVHXQK1sh1J0PYdb2pKbjD9RxkPdZbfn6iRGXf1XWBaTGsEecE8CsU
tSdmn55TUE2aNSemjjZR6rGCtgVePBSElGHEbPXDRoylxLNhWsdIsASUVhSg
ie81EoNVX8WmXlec3xh/7R2O6UVrJdPQlQUCN9NI54lWfzwka+pKgBnnW+LI
CKPbt4WROWTaP/8scJPtwD8aJW0YeJGYMf0AA+5s3044v7rMawMQtf/3IikQ
nM9jY1jv/ioKXMeIc1TCpNSV05t7WAKwAbLu2PD0rMVrLT8xtMaLcqkt/ks3
ziGuNf8oEQp2rvwUfzAPtFsrAa3/nP5p9AGgb2xZQ/lP/B6eHzIfHb0nZ8fO
Asbu0Kr2sQjrG+iWbYCTUi1OdVAXjV4wzIRVgRjYEIriOWm+TH89kA7HrM44
316HFYllcKU8s/ogPXgVQqEVTbM+s8HyUf9jmKZhBzTVhhI4lydsQ2r2XW83
rukIX2ar6mMrl1z6KcLkrpx2/2X8ec8nuMme/qd/l3QYRnhUgShhOJVACVkC
//SOAHRUhig7BoD5wqoQT0LX12IOhLTTj8nEscHC07iHuM3PK84dq6kfRm9s
rgFhKsvytIU0TL63Y6XXAWpLNrhAJNX3KenTsZ9uoerg16udvDcJ7fMsAXwa
s6PLCYFrQEhUEwALoTWH1ic/v/7bee4dcsvQuYJUARYpx17dYFdqcVsntTPl
IZPobeDwJnlCfigDZt4zB6h8yLk+nSuRwEKT/QIGHDKVTE+3AT5fX2A/Pwfh
m6rBqYpckoSGXiwhTYXA8BEla2t+4DeCH+rIoLxCoiz1hStelTcqK5zeC9V6
k5CA60KZqBl1WeWJWM0o3PgzXNwUQRSkDGjir9znoVG6qgdA8szSVuniE+RU
1udcN5gSz1V4axtu2u/Fs/gsGDbu6eOnUdBk2rq2yA1Zt4uG25BYLF5OdX9p
HKK0CxwMRPSFxumXt2O7rzSSGdnE6SsIbJpEVL4vXE2PCadTt/mL0qT6IuBF
HRj5V1pueSzE2MWY9ZGKVGcaCc62594MXD0UOtbapxXs+yiyvk0CP+xZw3j/
qUdGgR818sKffSRvDEFzDuf8/XW+BLO/l7niSpoJcyfbHYT9DXKFqSF0Gmg6
3lw5oKqngrSWH5Tw8vJ3nAtUhL01Bxy8dOSWs6ZN2lhjfmjj4wvnTvZvJov5
ZxmeYiyoshGuv3ip/Vyib8Q748VQf4EQl544g0hX+cxVQJyKWkM7ZniCypsd
f3p0Yz+okNv+znmR9oBvaI1MuKo9fjIR1xVb1+kIeob9Sb6iAVsxW/TnRmKB
3qAdBqappMBJ9n00StY0EiEgHtokN1MdzphbRqJ6GP5w4wR0Nm4gCf9GHFX1
OedJ6Yc0W6SWuOdXSZlVsQt5k9aY0P6ANts99uO3+U403dhm1QGiTuYSvUsd
2XSwSTqcsDRcF+GrCMZH6cgWVqV2vXarvqHXJLrCT/7AKzbfhAaTBx6txKhe
Ubb2E8wQwrfxenqsvolkPg+2N5NU8OB82kw9j/C/JEt/tvpfuYyM3Z7drdrC
8RyMgcwOyOSpkmNRPNo1l/mYmGltoUg+f1wx1Aqajj0FVFjT2RcII33feygQ
3YDx2gufB62xhhdWBuugDgI3wyjRANefqt+L739W/Z3+JBJiBFBRH6PHPnb5
/vIXcZxviuHu8fjZ7RliAMXm0O1M/gZ+QDcy3UsOxMVfeTYReUqFFGYfRJRb
CGpGyZSXx0zkXRRQHTzk7VYQwCINvr1yrTJEUgn4bwwHH3G9PXlRDPPIssFK
f+Mr+SqHLyazMhKohj842vlpBE6MOEA555kz8Ib4wCWL+bZi1gT4OlbA2awf
t97O2wIizTqRZzSf3GFj8DzfKKhvkU/3P5D+n+Y9FqrKtzMC6soc5gPT4otg
jl2pv6E5WMLXthv2lPwKKNMyjpxwr7kSxfva0KChUsGYPn52dfY+cnO6BeJ4
gTaMPf6ubJ3DJzcbXWfGvh11AT2lLsSrYjHHmbxvJpfk1Ac/oi4Qgdv+LWav
axmQhdraTrFPkcaXCwMZQVrmYNBX78gVqlPVa/0aXtzJjWIkqfaipUAEK1XF
5XHbT0VkSonJkjkxQFZFbwPWQBpzzT6AtwvXEbJbvpeotEHSRL3+Os0sY5cl
dHKlu1SB48gZEerw8IfTKuMUmaqFOxqYU1osiMoLYWHstpt0oVGz9uuQBMCV
k+ChLnauGW300lV/JxCPFo1Zt4tcDZczdGqi13DPJT5dw8gjDg2ZiVpLOEab
ywPg5aI8esBV8M8qolZfzaufr5ey61OXh7iDMYJcfbsFuNKyFYzVoQqkBM5G
XBJOImb1fhwThURH/ttbCW2gO1y5ZUfq9j2beNplPQVZik3kxzay0NBBMMVT
jqwBvhMbxvC4PF+myloRhThxjxEpbPGMk7DdT+bBWBOocPrcdgA8JES3Ea31
yMkXYSMRepxpKwmeMIPJBHDz+8lqbNbBX1vgqzd4pFt1FANyNlqYGtTDKCFW
zjqZ4Cuw9+XqzvQUoLpTQ3iFAD2bTYYgzVnor8aRNSFxaEE5N4kfGfeQIIeE
hQPD2iGU/qaLXsrFWQczhC6wEDsoiymsVBskvmJLNKCWUmvr/aCJbeTSqeF4
zpM29FL0X0AiQII2zXgQbhDsMQHg61V5NWfPbs4vCwK7rVftS76BhG5bw+5m
9fwF6K8rd4VDDWqJ/7fWbLi/dzVcmRcs69A34h2I+VOdaIHaN+EKB95gKfhH
dSVxozGWlK5QiKvul4+gdragckuFZIatPAABWkKR0GnjNJEyQHFskz020r4C
psALkz7/CtxI7KIKvthHodOVjyVgf6tEyPESqIyNf46K68196TLC0TRQg+X0
+oTlKFar0tiJlRwiaLhMkZGN2ESnPSKqQmyFEiCHn1v6xYcOpKADuadjZvjK
TDWSHCpCMHph13aNTQ4BdN3BM3I6K7laEKLDbkaMdryq5Ybsb/C+/Npznbqg
pGexYHRgVdUhbb1vhWj1JsQvhzTln6FUXhjrRay13o14v92SEYNDUPBs4t3n
8uBJ85BBXu108bL2Zw/8lbhDofFGFNhA8beeQXIMJJMqsRNQOqGYh7POd4uZ
LFogFRDVaZ01wbzGmMiXe9lmy4YTOm1UPxBHuuN0FQlSGWHSoxo5ys48SDmH
nkSz2UWDsMi3FxTxYileQySHjOCjPUumx+GEv7u+JISXhZRzD4fy/OefYRS7
kvlPJrGCCAatMH8+vJG4GWwvoEFSwRFJjXYu1bJ/Q+pg2q4O7zyheWtg11O/
wzexzYjdoNc7M+neBXjEr4AxXkdesw4UrSjorIFYA//UIA8C65z+IyM2XTlG
Gk1O6y7+5MCNY+wzLz+0Z/ES5eVy4qOl4CC8c/9vxixFW3MGI9qyrZzJauAQ
aJ+M8LlK8xUrZ2K0iHw0KZAkowMOaBCnnxmvwAZBEHa+qIzHOeS3dJQ5t8yS
OMZoblonnVvHXDmMPaNqv//76dmPX7MaZOLWTFDQgAS3PpIGxDN8Ss/QXZno
zxwtQxhFuk4kVbYDsthHhKDW9m/rG1O72sl8JvppJjCyRmUp5T3Qpx0YzWmo
+vUnIpVi30gC34DuJE9NlmjnITtQ9/gvqZn1PdN7FzlnMvaKkBQGH3LQPaue
cLJEmoy5VBtreYEDi1qbMofvllLTwllzBAY8mHADmM3+RPXUh+ehnL4JaB7U
ZP7SK26Vl32BCDe+TlNEvF7kd9Pf0jy51R4v+sdquuHDnhNxHL2edtFeWBUa
KzF7Y7Vs2uIG5ItVECmvMxnHKIdzMleytvJ+7qggD35ft4lBSyrI2tCET1ja
sH0dpoEHPuWMcSRNcldxRvSEHVeJ4HY87cl66K9BrsVz3jwOV3WWc9zsCHfX
uITJIMUU0FQUQ2jUb5Sv0m1Kb2d+rEOAwng9yd5OtabSW6bczYlZnmoFurEU
Q9gD/4WrYuArdgY5LAJQyg2FiMJrYhPidmP8ltiL7diaGx2a/qvD+kEmqryX
Klz2IjNtxr34ZiSksfbwBXs0Ce2AOpMG9YTyELSPxl/MUFxo2kMJvDQBHUxW
G061k92M5CERHOs5j65la/YKKoz8YdGtzMnCJRM+G8G6vW28rLaV9PhUqSL4
9fQKzY2o6bHKje9NjVQy5Alkpm35bHTRKOtoyVOkdhwI7PDSavyNwWGfvkaG
2cKOvNmtaQMtEb4ZLTnaxUv3WvE0pbvRJbeUGoYd5q7Vxqoi7sqmSWyV0PYS
P4y3hIDfIbFv+WYWsKV8hyBjIh0RjwTjiWl2G8f+avrH+4+jCkaYcT9eOAJ3
NodUdaWUO7FX4Tgs0v1vIdDBVtOXqPh3cV/u0wA2Kh2j94KdifVTLN9+QH7A
EAbhYVQEvP3f89IF+17lqOYe4xrNOGHzNdvuKG2YAsLDwGlHlr3ziC0gqK29
NpZoTyHR8oklMMy15KFyOJfbmfHIa0xzkJ8hYytDP0pP6thAx8I/K+OETHqp
JVC5lCx9qT/VbYtnGqCgfS8xFqEnfSllkmrPWn6c+HCBxOvx559n0Lw2ZY2S
JatG7puKYJ8TdZ933X7Oi2zrEG7Q5sRnv+Woul96UxkBo0BzAIc356iglCkZ
J4XXdfZBFS5D2hJGzva87KByiHmgzYz2AJ38pajnmwAVTsvx5JQ0gBqX8CZQ
r+QCxMCXsOJ9IxA6mFwtmWlTRGL1VRuXI2QZdHKUFJw9eHi4Cf9PC2fC3AMX
wk4jxmuQiKGsUIFoaEzUzmR3LcJRXOQTtOflOE8Du7NWpQ9xn4vbEOLDDZe4
bFBZh5VE9rNafcK4m+WKgRTckA6gWc0QjmXLw2Mk/1heG4vhf1DAFVRykX7y
nCbM+ToUX+WYJ0Z+H6bx+Wsgx4wbBicfkayixfSzh/AyTB+VWEQQkb1oHNh6
6Jw+7C6mfs3zFwJIplqUOcIQPgWoxzF2pnaJ6uBucECS+o3yL8lyvtE4MHbn
sfmJ4ovBBqnbfQ0uxolCzp8RoimX5XNwVK9lzg9wiN5EkNxJE9lgJvyV5kKr
BR2srrbwJK3gphIR8sd0dck7Ix1cAhCOvLFqIRmvKMa5Ou0cvSN9fD3sGooe
yNqHy7RGDS/lNvK83CFOYZF3l7BQWOpx1OaeFctqyxLHIjN5zzy/8yJHjFok
2jJbiktGTm6h68tGHtQgCdg4I097kztUQ9GFSnj/KwAzxls7qr3OM3LHWg2b
9JQVHNaOvfvNcwIx/eX0vv9OBvamv6tgnDgIZ7M8YVcKRBDGlMTBjbBjodod
qQRL2xrkTZASei7swHTYshrudH0s4PS1Xfg520WHGHB4r+CrzYb+lrnAFkId
OMHVl15N/bgncPwPn5HSWS94ZaKFwOFN8mYvQ8JC6S9OjFi/7yyx1djDojE8
o9BAs5QQgj8P+pGxiw8rIcBxsmivPKho7+6Sf/GhffwlI/nLWPrsqLAQsg+b
iLDXuQCnzgXQxnusDZoo+21LhCt+3ABfhmIXmVQftnknISJmWW8kK4g8T97w
xFPQQGB0QeBsAbNUdcieCZXAFpipaXa+2wXJZy3rxB+L4AYmYXQjGhmdjacu
eXAxSd3Pa9aCcBBJj7aMzQV03n37AN44QCVZBUZdjN0lRgEq+DD/TA5uUFA1
Qt2PFMlahk9MS+uIkYO0Nsiz4ACbt/WtY5mEEkOhedEiadE3Pkdc16CXbD9M
iNQKjVOwWoIjgR4CDbC3bwhbJdzPuZIBUeDQzJrr9DOPVtWdPJTEm8KyHmq0
NEBU6X1fjZz1vXzxq+ZKcoCMIjfXe30lwaK/NLz/PnKJ6zBcArsFj049t39T
lKSIWCIc62D/mphItTOfDFRXCSGerADTYOMK08two1LMlT3fmQtgAsho6Wjo
m4p1bxnJh5aDplvLSJe+CjA7ho1xTxmlDuLCGP8KfKIazpZ3Cf2npd4PCGkn
u/jALQ+3ZancX7Y/Kqt1yEwGpClOKzYtgVQRey0zDTP/L33CqEk0BCuA/esM
3zmjPFLRcUHSojsHSKfDhfpm+Yw4TLXhVmivCd9Y3EvNHx89ZkVfg287fmGV
EqfgKQt6tdGWbxXFrSqcbXH8htUXS15ooB3e/lGfHL+gJsXEmqB9l9VYvtbh
NzS5SosT4QyM/MMc6KjpaflMLEXQa/URRh9S9LBSC261lNhWeOK6/Qw/TKMb
Bew1fqp9yKterjeH/gVyN1ZeOG9D4jaPl5hhR7GIiQAgFnt5PURv4T1c2EZy
IZycRWKQF1zLyR+x3+qKGPpuOklLerOeML804Kj/34gANRaILXOzV9V82WXO
UOn0GatSi0AQxOSw+F2iFfmxDM+/62kdGCnkyYwVICh0qU+ulMse1Ypqm3ps
tGVv1bgnabFjzEf3aVXin5UoEKDy9WUZXeJrij//Th2+JEigIiD3zemr305V
rLEXMsvMP5g2Aod78Efc8OsQ7x/hDAhgGR3lKNlqU5Ez9Tvirz4mmrgWL9VJ
hjr5gWlMB32j8spUD+QMT6OHXQ32WYXk+TVwcOMRYACg5zN2717/Ei960tvm
nPvk2WYOW1phhYoF0jDeTuEHXlnO9iAwYrzvvRK0rWMOadf63TF3CJGPLRm8
9pJTaAOSXXbhDLDPHDlEqqVWn7VkeCYbI9Pg0XtSR5GWwqaeI2RG7K17lnug
NOAVSiuFAuVz6KkzYc140dHlBw5ouyniK4gk+Vh0Q72wHjeFX1i7SudFLdj4
T1upsT/gFCyIIzue2mNdnax5mLajG+IW09Vxfl4/FANxzGikqT2rZAQvFkYM
Kg7Nv0jxXxL1j1lbKd9v55ZiG1iqRv1t2qlLmpvRorAjBWN0rMbSjqBh9rVo
13wExYf19e5tHrsPp3UiHS6eDoUrhEfkyINUur59xp0Dpygt1l6x1sydOu2z
sI3/2YiYxNNm5I95RYn7HQs3ygI84ex4USZxIbjl9Vtu22fmUoEZsE0Eq4sA
sZRwMDUi78e5joMy366Ib163GqiY87okK/h6LFTiBpxhAELrByzp2vmpXigE
w6Fc6599GRlgCOAjN8H6KNlwA2S7TRLHfvbyAH1uJOoO7bDXZ8lEfV9t7MVX
0+GwuacUeWHlxtrwfsroQk7JutuoUaq/FdaKGz8RuaVt7RtrOXK4LjrI7iDs
76p3J5rxNmPJXiqqKVuM/fI1n42/dcCvw5zpHb81orvgT2bdinE/Y9C+nIpf
uPubAJ6ItF675CI+5tmD8rhb5mXwLPVik6mS5izeC9hzbC5SAau/6dJ1cXYv
gWcULeuQLbYF8NJjVSNSBpLglYDM7lILduZdQAl4Hp8FvV5wVrfkhkgd9efJ
fjHzIqKzp66amMkRFP5qdlKABIBKEII0fqg6VFTxf5JgmQEOqBToeM0qa1ZL
WI6P054imwYl/4yBuQWvzC8KNGVILOO8iU5xmuW/4ARceB+671NYkUC9rNTu
iYngPKFDruhJFGlI9di6SEB74eBj0Z/EzgGUa2yPSoX/edW/aBYLCQkfNC10
vqtiQhlkGxVG0u6jImE1qcDvag3HgMF122gKW5BMUByFmJscNe8z8tgivmLz
FChn6YVHkYyEXlxjYDCieM2/R3Ml25HS/pqjKR7+5Bmyh+eJjOiT7+ybvMJ4
awIf8GoT2NKHoit/hqqSGBfxJyAPQwVk/G4jPgZa9VRYDTf3jzVt69j6ovmT
dIi9zIjhqtD+wXNivkoYRnQKuBT0C0WSQYEWCckiXIUkM91OkX7L2qvBIX0S
0NYt+wPfPk5iyNPz0Wig9CscuOMoujjGlMqw7hyv6Mccg6gORHuO+8OYwZOa
u+mkHHx2boCAXFsn5iCN+Bf6T4BovPLDKgBdM/LiYM+Q2B/PgpPJ1aiycpBb
FMg4J12nTFeUKJj8ajWHXUs2+l6eT7ZB5UwMV9WUirXc7K4h9gIzRL7TIMg2
AfYrjaNf4EO35VuMXc+iQuWzSn4XROuwHirodrK+cL6vfUf7KEqfv0nLMpRt
7HdnmpAY5FEkETYq26w+McH56JIKJ7+E9JqNuQVj2trJ3O2ScxTS5wvf9/Bl
5z/zFEwj7HIApGff2xyZ61I7Hn5J/LIh48OzY+4XW6o0xYrFlQHDl0qBadEO
79wICMUCjbsRKTYqMbI+HBg3SVMoXkwUdWNa7/Td8QuweqEQGbot4rXuWm02
eYTCKj/dAK7/eQd13hWb3ahrdUNzDD+PtRouONrFTjydPZa48ZdBtVHN0d1H
7ILF2AW/0gk48eTibMkdExOH0NGfLzcqHgTroJUZJAv/6JvMDD/bqr3B4hk4
9JgcL31xGMtMPQypxtXtvA2tk9fPQFsaf54b/KXJuGDLqvCi99UmHejYkAgW
IIK00XgKVxKRMBBzq9NZzCNGAtAdSXGz2MwoxOFssSuxnVZkx10kCGUQZvw6
SOOYJI4zGvt0dh7rje7nTCaEKFhHpsFn28DZQvoUlG23q/vMdsIo86dEYLsC
SKk5kTJiC0jSAZRlb7B5LSfwW9giTQ4GJi1JbjQaOssP3BAOak4LwWxNPpyN
dEhVl/TW/e0T3KP9DR1ALAWvT2EJEMORenC397EofrkO0IK0/1ofRZL6vWoi
WAhOVVzA6pAPgERZ0EjjmtdVt4mIDCiAyh4etqSNrQfRa9zlGLJo1pBih5jS
LsKdFQdMoHAE35k5G8rRuKlVmng3q7FogU0yRy38+e6MQNISIr9GWvMs8LLn
8jfU2VDlH4WgxDSpkVfy7Om38/f4yAlSuDnXKJPKWcIkjuBwFow06Uad+oia
VV22VCbQGWJ/d1wFeVmdDL9xyKK7Fg17p1kF9y99D2zja26EwHSJ28BbV1ul
IDWZepyj768KFSKOthVaOS2rFvknNuRlFm0AdF3S68xclXyincQzIs3SDfqa
fWuTChpTq9gL7UNg5AZNaz2TCITx3sNbaJ8kDaykEfgd0t49Dz/ConTUR4bp
mBCkQJgjQjaVHfYRzIFojBNRpac71qz3s7jt6+ccfI7GQqYpz4LVW9xZMt3Y
tTA9AtefUA8hNMB9+zXokQWTZYkvyT5ewiMdJcFFIbqZWMUiZDI4o298ea/e
5XYx0Tmj9ffMOuWFlFxOLZqUWx6yO9DDdkP847O29DMBzca/QEpftg9JASxU
Gy8m1XxeElfmO5gSMRG0D0yYPVXZtq/7WDiGRB7pHp6wHkwljvCsA8glLdiQ
h3mAU57WYUwafhtRI8UkjDNRPfA1hg/nmqnfzC9WmdSSrhg9UlZ/Bu/6Ozro
kQUuGzoW4H82YbxEh8oGJDrhYK7SOl+CHYeFhP7FvlY7sALQDhjhDB9lqGhC
rRDdEAOw6FoQ1+ZEAPOCDeyYe0uaIiLEjSbJ29zeU/1Ql/hyDTDQFosGFHu4
4f2dWp5G+ykle4tnrUpEEmrcEY5CePqD0k+QXLp3hzcAU+3DQFDgtVZJmaos
FU1MJPeXcq4GBVfFzGbWkTamcoS8LRNl3YWoGl8EVtGmaGx6HNbx7huEjDLZ
hDMoaJx9vNcb0ScL8RpwZakU9D0Zw59xskr4I160daCv9X+c3a8uE3hmD3y7
hWVd8q1QL/RPgenXMj4o3I+rp/MUQYf7uKh64P/HO4oD/Ooi34p0Vymdp5Tb
fShurXZei1DH4P50Vb/3mtmKzufQJ6CyO/6Xz23tPK13ynhsOW2oYE9k+HRL
Hc8oBNZAkn8NSn+zSgMtpqFirhWCvGiTqxWLl0+ss9hg4nfTEdcNPweFnvJY
rnl46lEx9pFgXGVzuoFgLWCDXZK2E9hCRkq8aKE52XUyt5zKHOf9uU1G7ktX
PmwRhuJVkeMAvYNNEAevVqaAsFOUkDM7j9j9thcYRpZllKvRlvZz5UhdBXSN
jBBvBKKK31DX+9YYv3zXzhaPD3x1gcHjY+UWZqKBOMagyzwfdpn74BZGUxZ8
zWTQpOPG7G1AZPCTuJeYOw3a8ai4arEIAg9BHeSCKdcaWjCfPjEVYVJEmwzD
4eadhHr1rO1kCj35nvIzUtV1+3qr4JXvEh4AOJ0ywayi2KWEkivYmw2DfJRQ
+Qu1I+mGoxrCOeBtysT+UJsnvBqkr0hoGr8nmNHK4E0YBu8DdxZAJJO2ff7M
vdb4cqK/7+2NToQUoo15gYIeMIgP3qRwpFjNN1pDOxXBZSO9I7/RYxI87NFp
Sr9MaQBKhr3HxbEQML+SpKFzHHPn6k3H9bo+TbWk2fVmw0NgRXqa48vZE9gI
C0D15achwFxBUQWV5bnj5x8C1cTvsSGfakGSMvqSSl1delpw3ImTK90kylaG
c/H7S+6f2P6BxpQF6UlnMCJGrEJAgerD+mTMxVP2vDZZTV5T1YJLigxYEd20
ibY4vuGxt0P2xB7lHbC+Mk4rgz9MS0xr9XS3fOZon3NYHBK1NzHz2WZf0WiB
nmY+lB6wCQ4RWN0QF/qnrBS9W+Z03+b34Bd6lDgFuF6QmQPYPPs3XWLf97Iy
2fGSzyI1Lr+yL8uXwNDK2HbyJeay5HosUPQkLchg2NKzjwcFBfLK+DZjw4Dv
WkvO0c5uxdshq+Fy+TbN/UVH78rwunHLa1RVvB2OWQWD7h8NI6ReO+dEJOHr
FzL7xilc2Dlw9OuMH898n/pyo4SMK+jxvssxE9rQmkco5CZSrFX/t5jwHeSF
seOaCSGr2KHiIg3q+0wgH+6qkj37fOdIZomQe4EdIQetIjFQLu11DH0Zv0yk
IF+BnhyKOHLfOjF9yaKfg2y/AsiBKEEIl8N1aHDpTNr0sr8mTU4K+6oOJibR
qAHSITNWKozLGTy/m9688P4FFD7XApL88OHoovWH5V75kP5AUH6mSvTBJcWi
YeNB2S9EGRoXTEDyRo5nI9wqX7QqG1LUHe5nxnudAjlDvbroOIbMKXF2eLRm
28hNr64amxRKGZHK5orjZhTikQllGEbS4vFtEkZlaxuxccIct2NfgF7YhHYW
J/inLxuITYgaqVWqc1iRDBqmP8E8OYUihecJ+mYnNw1FVDEy2JK8zYClSWes
1bWdvxgUQY9SmMlbNG8FegGRjws7RosRUM864mu7kwRVo9z841OtlXrP5MmI
2hZHEkymgqK4i4LgAtR5+gEjGUQfFwh/hltmEozLvzHL6+Xx9G643ZL1+kJr
jkSgJl6MP9Ub/WNq3k2fPtMb8vwHsBIbkxuh7BzgqLFfk5QWC9vhPMdAlPSU
tEruxApy8f9ELpvbh5iATxa+7ITvXobHxGI0n8qPaNhZn8WG2fLVPv57Gs/k
P6/mNLy/XQnWEps4fx3Hl04zSr2lokI3F7n5l6G1SnsDUc52GZM3nvErvJee
RmaNrex0zUPAVz6ozTHBfyg6jue1/J+rOMRK5zmTfKUcuzWxSDViz62XIQpJ
JSQ0gpZg89gdag2VgRvtyAqwSxftxpkBy/ff25M7WupDlLbyASGI3kApGi/G
azOaFr9DY3IujCYZ81H3R9HG54snjzLZ8qLV326AtQm3eOfJX/FFE5eVWatR
7ro2UlXoyrt39lrCjUpFYee9sf9sYtEi+5Q542Jxb/7hBaDq9LqEAoO6as/8
zmMKtNEZMP/iXObexrXrj6KH7NSAgGAYp052unP8+b/GoFkbf+OFI1S5uxTJ
827JTZZbYTlck6ZB64cbFaVTk/1IlaFHIkJvpKkXnEkdE4j6LxUOGdye9Cms
i9IZSX+OnGA3pu2gmuEE4LS0pbopgd4V5r2+aFdCqna4hv2RHtTT76g/oflb
X19SygRyqkewh/KygyEf/fcHuwaRpaVHEOeERCkaFKbT08YPLwAAAJ4njs7q
Xvl/h0hmUpnTIyOf4mHtqVdZ5NdhIDUXoasCobYTIHizFOVfV83TxZgGvNqg
FoNM1IwZNxbP7cAK4FglxLNUDFQTyrqGWdBzEucspY1mcD2eKZNhe49zDDV1
HrYr5Q+sNfQrrrSDsP8Tz/A181m1hfVHwqkplCftTyz0yScqIVmOm8+ZSd+q
YzaamTl0Iv2I2PMOR++dHxvTnCkAQzPNSnZBjLfOLNmwSI0eVBmOhK9QbRlP
rjcbbCQGtkxzYntP/xq4anXsvrQ3PBNR0WHZsi612hGM93He6ZsRYVK+Spga
INpWXa7ODNrmc+CrzusRCgZenoDh8pVUVuVybpMoUu01JFykhp/Ump8aPfmG
/vZ2wxPF7gtcGEJ4ncGj8gXD/PceqDKyQshd+Ts6dNxwpjgnvaKipK5amEAd
N076Enol/54UI0q9cFgpce2WajJkQzZWvXZV9veAxcZDAT+w8VrIWj7ywLF4
5Jj2c7KqL/+D1SvPLdGnCkRj39WwD2LE8cHReFt68Es2d2G2YNq6q5smhrCb
gb//nU4NGFKssEjXZU4QhyWWgvmBaiAhQaBLVDgqff041EwMEhy222pjcz3+
CNEOfcOss4n9dfzVnT06qdB1Lq2Bn/FClODNir0JXNen1DWs/sbKG2VU+70Y
tPfWwtJ/G/fbufrxhETDb4iFWAyRiq2dYtYAMcmemMcIH23nZoWaQgcToSGm
nt1BnVbXgBPocKzHuF+yRuew0ZE33E1+KQoBmacrrBaowqB9Oz5GdUyAZGaB
w4IiihK9ycxpGifOuhsSaVi0eHSjMFBxRwViV0F8+4BTNH+NMnGW1I7ZodtC
/xyj0tiF6Vz2QoIADa9x1+ifUpGnyEq6JaP4JT0C8b7+tJCIIODZRIB2v/OJ
qEDgfVFH84myo2D1x+qVVvnElLCjOmjt9x4bYtfTtGQL/w5CUMqtTkNeF+/H
Fks+OvzJEM8ZJqEP0eoVL43vkvg+Zg7/fgP1bbjwiANENueO3cgJ6L6xSdEy
TP/c2XaEMzXMh13dct7JFlBiAWm93a3Kajqy1bJs0AC6G/YF6skiPI9O/rDv
4eKR0qAHLBz2osZCijghMdR//djXk9PD6cHjYQjLQxLjQfQoPVxAABXbQA1D
Ta1g442I/zoG3ZlJB/1vhLNzO81rt+DGP6bIJpUj7Ij5n/FF+bT48Kuqevdc
x3F0Aknh01Sy8lSKxgY57+C7cCHFDavbhU53Qb3SRMdqWKsT+M2l7jtomxzx
UYvTntV5a+kUOtpNxXo9OPuW5K59R/5emO1eAIH+uk4AogtH1ObunBXlf8r4
rZf8hrUUtTk4zljOzVO8VRf5VEWVPzmEtAMovnCAHY+Rs6uCYw3CNK9JWImX
pBxQJ369p06RAkhex46NsnhLlXKdNbP/kAhfQj0Fuy4yqq2RXm5ZoKAEA+Qe
zzvHRK+2Fmas8aq4kNIGyG/BxQQrmqMDH2MUbfG5E0tDH2Xvf9g6nDS6DZ2O
Gdd8fqinrF2bUJZeCG3ItMFjofJpkwHFsc7/RSNST/VVmis7EiSpa2uX1taD
OFUJHkyK3fqq24oWknVlKtmHm6mjzr68e46t989sDTVnkEnrSiRsUKyCr+z1
9r0nxASBTaDB8v/E7UbVX9Z02OUvCq6q2pfVmglyMyZvEuUor0KeRor3qQM5
9Kyf8v6AyZ+GW9YCBUBTof7ugCqZdB2IdYYY3BHC8593n5NyZZ2U776Tc28d
3o5A3L4Saakm9XOOP1ynxRp1hUncVr6kDuKiFj/YIvaJn1GEtsbQVf84QKnV
dLPA/DKKNG8bKhiC2se/TCjRy6lHHu9ahtAzYX7hrdQPlZzbWJNshZ/gAQUW
ArtFGydE9h49gYv3Skh7a0c/ccbVn77lbEDEDiyUGZIdUFcKcUS967SRT9V0
uCxErs249QNY+8DbZYI65RnZWvmmcyeF58v5nsWpvvS0dDOJ8WRDYzlTH5Ko
dtCUZHk2+2bzSAi8DD+Dlx/24ePbnSTAJ6e7py0QSwYO2j9plFRcwdR4oaGB
9tWvvs9/HlUT/NbYDPbV4rLN1qMlMjaPZbOS9Ivo6COehMmM0ZHwAxoFczQU
oSaHcbNkjFUipz2jU1oEE4zbgVIzKntXRVCO9LgETJhiRc9cDm34guombRtJ
6zY02tEhNDXTn4SrPTIjm+KQYxgzCGFwFmpDJ6xoSu3VXNaV5hhuXOht4/TI
xbE5NJjMWxx08TFTGV9hzeCqQ2/IZEbpF2LeDPUwJbj49M9Y6/F1J8ez4z3C
U9ShC8Z3K6AF2pp9U5p1G1Lvbnqz4t8Iw0/Jsm5eUbpwxtDlUv3aYHl59bHP
ki+CjddD8UqhOf84XH0o2SzyPTdzDCiS2FXBu89QGjNOYFdRmaKsSMJwSH0/
AzR1lhS8+oRihivl5yxV43r+APyfywAaE+zDEoaCdhkayPAm+OjPtk1H6Mbt
2DPufd8fJgp2XjzN0/usSyf38m6nWF6ne9J2AVuXop169ShZ+GFaNkorg8S2
jFKJaFVLyfUs9U0BZXmQswq6HkTpd3h6nI6+5waWhMqxCA23xugC5D6NVpFN
P0m4261CVfi9Kj8OmZZurfWsjR8xlb0aR0Ee34CekS9LXVlIlEiYvElQpONR
8A6vbvwsatT/JuYdPnfGBsOYQMqctL2gDtxzUtKnMhM5kKTWzGwCFDSsXOkY
qdLxXFymHeNX4afJXyLcfy/aSvmCg2zd3RgVxIE3poYuCO1t6D/kMOPK3qCV
8rHs8o4JxV1LG3N5cj7S4DKhLxboDfMZ6/hOtpTSs7SqK6e7VvoRrCUT/kXE
/aJeRJWWMgu3QMRr5OU10fJ9X4ZNbWS5FIdxg7bbKQS5pYe2D6JdEP4RSqgM
zSStkqpAx515/oGai6eWtj0PmQ0QugaNC7tG6wWB9I8VbPcupP0sTM9yivRg
aTdaS27Y39GnJWMwpgndeZvZ8IfvHxrBC7YtrPllOhGcH/D5CHmqEb8jrhyc
sygdRvEWESXm+2KXklXcQRWGWUEQr1ZsF3b3NGy35jI6RcJ/VdTtrtetwIaV
3M4jV+zEzSKjWgSkcuJljtDvPd7K6nBa3CEP6lq+j5a8nalcqhCoNeEyEx9j
L+wptga422d349GFMX1vZD7fP0qJTE5RdKqTbAATLp+fM1Qx62tdm4S/TUwh
jOON42Oct043YgrG65Tb/t1J7oayiI+KgmDgOs9p1UB7A/8n9ACCvEyoZLAc
2xF1L6XvTMgRLJL9fR1JnAw/KOm8cA3KoEEYHu2OwEAxfuyid3MjzEkRz+2h
TttnqxEl5Kr6oegKwF21wF4ljzK4PXA5fSpKgvzDW7cP/Hp/trg3zLfXL+1y
0BstTdK41Za0uQsVgSwD47cyW7qFrLjKnui/XZg/hTH83J5YDfG056+3kA4D
Uf3vmQmXlf12jUeETWiJIYugC8qcDKX2eMDBFAl43BEyO6PNTGgQGi8/Kk9Y
2Ge6kahf8Mrf9DUtg6CQMdp9fjpqTUl62fOPkTWfCozajMuY6f40R19blYIz
bjhIfZVgh+09H+DTUC66luo5zNKbYrZE7JsVL3gGzi+SNRLDd0NL3rO1SbYZ
ShHYgUyVXF/QUDCIOQNxT8ll4JYxRpzcoIQPQLt3ILrGiRmN1ufwJBosnfni
0vOGNr0UNfnj+hHoxjLMiPW77v1SVWoD93p1BK8CaMifTNiO1UK2VFcKkZSH
s5XeWb6oVNVXBEgqNnHveKZXN6Hf3mOtOPR9HhiamPo6nFO9qAd+hlp1Ykry
sln72YckVLqZH6SmS1r/THVzWhM0r6Emr0ICmhCbUjq+0Gt/wVyEf9k8EE+4
0BHE52Z1i1V5cWWyTrdBQ8baTQ0zx8Z5JJloPYYWezfV4k/h+dPTatDmrjsn
xF/Br106Mg3MwLMpb5rIrsdHDzahSlQrEC6s70TJEIERKJg5WB4Ov1ei/wWi
zvmn2mwFQzcNouK4ExVAYn9YzFb5SY0fizOJbCryQJI3/QxwDfXHt4kjBg5y
iU27nn8LM+I8UXQ2WwKe+p1Cj/8pfOWLoR5qXlwiyv7mSZlmAyaMkwAZjuOI
gaEzNW4sowpGx15/3F9pyFmSNLXgj/zO5H2TaZE7LeZPjhhdIFoJk5k+rHSB
OBReR+/z4ieklMuYW1L0ZJHzG+DymxPWWb8CPja+EePtyh/NSvL4BlQ1FHOb
70fA+xyxeeV7z/10FxyRZKtjyzm50pBlY9DoorhgEgjEaoKEWRApkCBTW3N/
EMkrmjvGPUNpu/wO/LG6UMJkRI5qQZfvxpJQ7WdRWVmlb0xhbnO6qKPLKp6X
B5seeobrbYM7Z0C5uNlXGreKz3L2N2kw87A7VQTyT+1eiah5NKu+03HXaX/r
DhCeUBSLqyzEqLfyvbOk3p8xBVjbckqpnR89Tzft1T4mMiobA80aBd893qvL
dmaPmCAMWdxXaAhlhUsl1PI6cEuvKAY2E1baQEtoptG3TCUh56qGJWYyPHvs
fpBSNRg+1ceQxNamKiJQAgL+rmtrAQConbp6sf/NhFMaaYhJ2WsyXfYN4cVU
x5d9J42OxO4frakaXBaXvUg3GXMkyryLZGda9fF6FAB4vcD3foz7JbOELlN+
Alx3zzbpyvsrWsv462T1Lcq3Nu/AU/8zp114nrb3Bx0x49EwzB3zG9BVggSE
hwjZ7ZK09yxRA31JDdan1kK69ylRTlCU8YxVASJZ/aaHrSCgxbx6j0BShB4n
Xzx1rBNGAvuNOs5OEKyU4jtYrRMdcPrluotNSetoYjP3y0AuGZxfJxBUE48b
rIYPwSr/6+ltL533pnupr43z8L8OmF1evCWHqeAeOI6hxrwxt/V1I0BPPyNN
xHC9DHWAl438q4aDIkMQO/BIVwU+GgF0OulPFni63GnGLM6ga+577MwdTwP7
NnQiqMZqxoN6qi2g0q4UnOJ/zDaud6MCK96zhJLB+M5MmYQoG8cFc3R0JZqm
Tq/bO2MG0sd+eS8lbIfTAs6fqSgvpGT0tVJXZprYBjskO+P/ixGy6jUdH8Al
rdxt5w3XHfa6m1hWi82V1eH5AjA2D2IsG98FU7aAgymR226C465JZ/33Jt72
TJSnHJR6JGngXEy4VAzikiEz5ITyvdc7/n0gBNR8RppuOgdK6t/C6anyBVcz
rJiOxBFjqYCX/bWsLCVs58l0AG1t2XLgF9p8KgOydARycJf9AzAqvZjBALoK
1tTBIjlN3/c0Rw1D4D2jaIaolNgmZZ+PiRGmHqnozMozzRiojl5S7QFm+aJi
eE/eWdioD5CXTHk505qy43cWx+5hND95deM9G7Z9lXlLZO7VGJoN/1g/hA7k
6+D8f85QCr9chg8/D1fI3IFh2jf6343kWB1lh0XWfPU5SY/jVFROhnFGR5UC
xbcUjvl0d3xtr8k7CqkE3dSUsgOkP+qklVAfb04W2jrycR5mENYR2mVOiQLs
sOq5jPu1EKe+r3gZ7zSbpzGUkdr/XI+URrE6fPCWdzoXbZ7yWOyUvmiErXmG
qRBMgQglIgqtbf0EPHQiIRjPHXJDvOsQoHOEWO0n2oEzelh/8c/HmZi5YLNf
rNoi/LeR+x5b7RSjWc9fPPKiEIbSoKFOu4mTt3ANsaeEY+ZOhivugq2mblDK
Quh3sBZFeaV5PBrt+aP8VmviuRbswDkzejlEVAqrQ4tg/WDhOVXYDXsaDpQT
f+32R6Z1+fd2X02fZvwCIox+i44T7r56puAOl7r0bgpEx+m72sMunOSplYF5
Q2/SeBGIDkm6ruU9u/Edwjiuwyx93nv7/UvMwFRMZq0G4fGpC3apWuTvUTuV
MRedUqTbQ6nIwddb65G9+LVkn/ybWHGPfqt8kbKlKzVP/iudTitNwd1GKtWs
V3LdxLJ/ZEqhNpWEBV/jrcb0/XSlvivgzng7xT1I03fBPZYKTTRLMdZNVA6Z
X5aUXwHms72PGZoXUCcrlah4cYQO2fIHl0o7jRJVu9MwEe3pO/EukcZGJuun
sHi4r0w2Uoqu6G+sOwvuhFN+HhvmgRgui+Dde2ui5VI8lvJSQJ18b+QTtSld
/C/6vzkOiQChqpxEMPc/oHDjmxdXGfWSCsEN4apIFyiK7mxk96iSYXTrO9iJ
kyWaxUpMkfPCkKS8+RBTrzQqilBcziZfrD6mR15F3d5+7D/pUWXJIaaFRxgA
DdajReb739sfa4rH19FVLOqLBi9G2qq3eRBezzVd7SCuBKEjZpvc2sqTG3kx
DUPA80kcF/60ZUe1xPFYLl5SqgmMDlLOFfEmVYn5axL36cewNhZ4WjejRF/F
i4CSPbFhK9kkQsm8/HKBMbTspVXmnFAFPhaTbj6xLDuanGTEcYMomxvK2hkt
sQxdlzWXPeKugfP0DkIJINanqZfPcS0c7+yWgmrAtJuaC3NRgV226TP+5BiE
xLHdjNRru/e9OcBGJ6UjoQDVTSJCmX9Kvj4cGQSWn+UPQ1NBpOTK4xkIzDbb
2l0/eJ/Yv+tunqyVHcro7Y90p3z008aBu8GuXeahZERKC5obq1d2e2r8u2DE
4q89m06rnSaCbdhebIdPtO3xjMo/OgUdRzDa4fJ9jgZaZ7+jUOXUNlnplch3
AkME9nUzfCPQx6gsrRz4WB3Mxm1y7NvkZZIwJ7SI49NvYLP1yq9iWeQJmfoX
KSfpmfnC1sbQhmZa1Yxw2+XeuhsN2PcI8KYE0SbmJ6Mso+B+abPWOHMDe8WK
r2ghiqUfhXUUOBHVcqbUcFWP3/nx4Fz27JgmsTn3jbPlpXUDs/slS+6tMA0R
pWRb1Okj6rTBkZE1DwijkyEEzuksDOR26SYJDZTOXLvBVOxYk91I/Q3FeLaD
KsEgZJrZKF02WPhH3tdEeNggRCjMDweU6UPjbh5vn7agNzz2l5OSi7hZfMfa
aI9dh2jTdqyVwbo5SOVQDax0fLnFjCZl5w9SJAF45wud21KqKvINnd5NsGoY
PquFzcRgr1+Z97dtsz1nBFzFkd7CsxtPE4xjo4oeXC4KNSx2PY4ab4lzd/Bq
Di9Tbtn9bA09XObV/ieySmWnZrkrklzqqodOSpV/PWa2r97umrXcmY+P9U7R
scbliOO0FOq46Yw8ttseihY7cY+naQhVfSbMj/E1vA6Yupy+6K2hwdV4/bZP
ohdXgvccTUQv2YqWzplW33nXLAyIbX+RIdr+LNvZCfTIhY8MIkgpWaopINeu
xunVv1detu4FqaB9diZr/1BeA8xS6g3i/3ZBDok1mazcdU/sBCOX/4Yk5vXl
aahwvLzk4J55rGEDW1wr8x4sjS4zsKkMaloEgR9XSK2/yJkTibT37P4iPOsO
kiqS8pl/tJmsUglOJ5iVW+XfT/3SZQe8jo9+WFOhEA74rWGZhRWaNW/R+v75
vB2SrUQzDJPJ6juHX2hfkye34cTsZPlfX09slIi5ab8milzYRO1pJ0zWtlEX
9lcmDOUrIoWWYP3ZJKX/1H5rHq67c23QTCINqCcUyLM7bYzDSksSGDvLwSls
hqlvyqzTZZvhJlh2f9cWBtPzPfWEsoYaV2O8mEeKvxjwLsQPyKYv+hkoOUPN
76m5Ucai0/kdAb+b7NMU9dvIzzwsbg2nJErkYweSXEDP28CspR+ZdQVsYIVs
mK40SFCuJWgS227xBTruwNl52ohVYd7b0rirRXrcKt/a0LfGf4wLQ33gowHU
PxU6pbZZO6bHB8iVRjP5Dsz0jLmiIar+/4aQ6kK0YRcbc4xAmmy3ktEjF1sr
rmQ2KFGPYVWuFdJWOZQBQkrt6lZDegOosaQ8uwpIGoxqsFDQIvWhVWS9MCRF
urRvhzCFMUmifWIAjDQoEzuuhRPEU6yQntjvcuhXzmq74sqOGaKfjwkvbEH5
IR2Dz5zjzi1eHqUeLNKww7vC4STy+hpPVC4lloyOBihjyzrwTADYmUqg0QS2
WGKAKImhKdebMGJRvM4QgpXIHIzd3fgiQM10c1sjwNYD3ZnFIy+N2Ih6FFmu
aAOE8PaXifPVdPA7Ccp4Ni/xTP1v67V9U8B2zzEnN4R2r6hs1vqwvePyWbFb
MtSK9/AOzp9/nYyu1E32mRcV19yPHBbpLacF3uNKg4+4tlXE56WQ3ZtFH1dw
jyoepl13iPf8jova4DpzIi6rjTKuZri08/4Mqx58gldRGI0lLRHIXRBNhFVw
Ix1wRiuo6A+1LPyXLlAnO+nN7q+L3M2pVM/L9UXZnk/RXWtECZCE2i5kof1q
1JLzpP55TctnuSRScpOOQvmnIlY57Gmhc5mozVsPg7d6RD1JzeiqgQZJVn/m
n30QC92fE7MfgdYLv7esS9dbJYHRs89JiH9SsHAmkuTi7TwKq47L9q1xc15t
v18Ei0/0U15HKN0SvdZBXR5wqHKsNzxmgV0Tzv61CZ5oh5HI8V+UUhVfNi5G
v1Pg/V41i/plFuUOqh+j0erz+Io5QUGLf/Tq0BcpdYSJtjYH1+IOP0q4aMKb
4ElGP0Pt1xMQ8FlMerxufs421/GYDCqVk/9ClWvcDlg1QQurOrX82Io0Zkfk
a2YV8Ogp5VACGK7Pa2GezF+q5O1MRA+UZ6lBnfXtFcpC4/PF6Ugu8awcm1sf
/XgdgmYGHUbZoKxISzjgS52wKpa7K8WHOLzH0lskQVOe+s/5rFETTvuzb0+K
NwJgpu0uUAF4IeBNEFOozzvaMy/+onh1Ge0okk817wRaARSPQM//qktlZkrY
C1xlocZjkbBX7uYO0Q3kQPnvAVwB9tfLYuhPIlvTCG6li+wlYTxp9walHfaM
+jhQ9vA+i2+f/EsdQQAKA72H4+VyK8C+gWjRenKV8MuX1PEvFYohtsfqk5ZY
rwrKUnOCmRhj3HrPSbruqded1cBtv5SBVrsg6+g3OyIftTkdh+iU5VoNVo4e
28JwAH2nnd96wmb/xSbZ68DTaZnLG0716Jdyy+5SHeIE/B48HuCuT9g6t8pB
gYrpgZLmgqH9A7YA7LqaoLTXS5vWtMRl/B+Q62zmneqi9O+nDzbXfHZ/5rMy
DLzedRRFHFxlsXmqkvpXwKcZ5JHHxNXzjpt5d6s7y5v8UqbAI0ytZCYbvg0c
u0xSHuVPlfHVhazggCpxyWcRCLUOXJ2eqR5nLFsVnSF4u9Sc0DIDNuJxzrGM
5NZg4fomJtzUzVyq5Chz0Cs4wK1Yuk/OZym3YEU1e81CGKjew8I7DM3ploG2
NapnWghIQkh7+1IzCXhlGATrJ2a3i7TCZIpgWpVn7Esu2toAx8vwbrYOjEEB
gL3Fxq2Xiovt4BSERTmPBfM3S+vCh6ESH0LhcDtbwCkxziE+mP0RWNzVYZQs
zkUFoSMQwldHtjZpOwvIY0YecD9WheXiCPhgGBtg7TWlBlS5kDh64YjWYBfU
p4YQGpmJvyG5Ye6SI31l1QCeNc/sro5Pq5RcQfSNFhN5tyRUtC/Y/5cQTCPz
y6+o7XI7M8gZbsMGFmwokvMSEFXPhgkkhNgOKtl085mvqfMzt2QkGE3dYW4M
agPbtHX89qh9F7wYmAHVPFO9hEZCvrvDpMCzDu2OX0TFG29KCDLkUR3NwqGg
L2y/yaXXGwfzx+fjG3XoZh923wyrRAgl+LWuYzqALxTnAkUQt7hYlGfCVnBm
Z47aVpnmkt1unFafu0+vD8O6SvCjzNWTYUh1Lbjsnw0s3X2o2fAx7lbhpw+R
zvrkC1Bi05gLPqnE98MNCGvex5+3fKpVK1TrLy7PJHzP4NPG8xx3VSx3o+IQ
YZU8eGfvG97Y1WSizcYiez1qLeXF4xvV6U9PBIVcXWZB4jbV+makYZmdL5Q3
EFegYDMArOgEc9eMKE19WZomIbQwGX1VAVHOnMh6/J8udVqSTgr9/ugkYe9y
xv8xEOdIZGAII8cQB4AtqXSvHPU4mzVLx3sCKEXeG2Opfd2y+VZZcOIGwDD0
FFmESicxBVditLKoQPieeryh5780pH9YXXFY+kKyxOA5MAKu0iWeQIpUsWjH
MnhGsCpssH+h5ZvDJeCsJV4Os/LGcJpozMnMt5ogKkeXykFwYnEAEXyoBJ27
7jbO46DOu9aUjIK8odARNx0fMqKsTUpoOW6K5cdvq1kJMSc4qRAU8geU8fMO
JZDV63nj2+Oy1K3M0AvMiv3ZiWppygjyeW+MbzFIxpIz1IkdC7araxJtph7N
pCxkXx50JTsGgi1IEuNqsdpIW1brPzsJgYoq6Jv9KnMksj8lkWDx8/UHw1rH
/t41FRJAw4s8N0X9dNnN2I64Np3cMd/pD/q2Kewdamm7FzHAl4oA2WiC3HW9
EXAqGahY5huHCwsbwUSHM7zhRF9+KPqZ2pgSZON9T1Vt3JW/+W1ToDbtBCP4
/7NRmTnE9TMN2GpfwWnU+V6VvPFIQfYqaIjD7CH9VkbNvbhNfnr3OqeyTj5g
CvTO8V1ym1WQFCd1SiRfwAxOR7etgXD5B7omVBX9nWJTdg5RE3hDf8T1OVim
ytzLkfxSUlUEhahZKuW9yFP635q0fueKW9ohxlklbLWJUAMqP7PymEsFNd/p
sMhatlae4OnQlJUq1THC21huEAqNxmqgbkFMUeKg7F0IZfpke6uf6MdJop5+
w0rc1g1FI2yOh4VCxJ0JqWIR4+gbrL0hwAf/o+DljzhW4J0+6JVr3UQiwg/h
LIfIPpNdZZU3aZrbss7bnv5TMkdytFeNXAFM23MprWG+/UY/duc2Xu4XG8ZR
lHWlu6ZSyjNaU7MR1Fbi672uhOTNB6efIs/MNhfj4zvPZ81h+VN9QEX2JB+R
Y4yzbIllTsfEnsihEqg4NA2eweHTOehXJANOUD3jszhSTzKG77njutvZwIHw
68J58GwnefcvMpHMVLSOr2jdG8I+70OcJrE9v8aAldnQBCndLLdj0XTbuln2
9g20Z5ZP8LYRDVIpizfNTEREtnLPbWOiYpK5qxcGA+FQjYkEL3JneEnQPp3M
SMgirxT0fXeB11djH0X9hoyPLxXnhrZ/vb1Lh90LwGH3x2ysclv5qlJL7p4M
TKGfJzSTyntfFLdWDy8pImkN0fgzGcMOXYAt8z85ELrA/yGJSK4k5ZhcCoWr
2Ifl+amow1AiIoph7hcJbAA91PThPH7UB/2lcCHVtfg8/2QKKyRj6hVQILCF
7x/CQe/J0gRUu+eVMUXJhYGiV//MrGz6j2KOeVi1h9wXbWG9L3eQwzFPgbAG
2U8LYueYxZs9S+BHVCYpyOwVL559d5n0yT+tYTr5Te+Dl7uVLpty3oNwCVlX
vbvcqZ1GkSxXHKDzn/wrj1yHva+CsVs+kUEcME9wBk7ydHh/rHKZLiXa81gY
Qh+53XmKaC1tjL72sg3/DJJsOa3+ljn5CNsciuDrUiaiojAGZ0x7ZuyVNZio
sST6mQGVBwr8qYyJTV6wtoQ2neMfnEDivSOMy4uKUuSnHC/qpVNm2UZnLxHV
sU+zQgR5WJdUEioGxtrGZP9B4+pzihRIxcGLh32f2EVi/anVtcAByLCK93BI
1JzOnPQ58xqzyUF0TZXPoHyJzUMjgXLIyeEAeSRaoj+GyXZXLHG5HbK2tZCu
KXKLq035+UhNGk50iW4pScza2Z1dpuirJsJKqwqwo779UEMmrne4loMzi245
PVrSGlxkcbtzzh0MNwQCOLOkIdhIeGUOOqho566tq/NAQO8YdzcOgVr7+7ir
GBtxMjFjuFLxUABmYpzHoFLKO6b5xX7GXkDdIdrNeemup1GC3rabG61pZBBl
ymxNvDtF8W18gZNSpsb6eJP9MGNaagtr0KsL3QeBJlZkv7ioRKlMfcye/V36
VQW621OnJSpq9zF4fgwNwxWSdu6WO5PdUsG1gByDWXtZBgbPRsym7Z9m1DUN
VmeJA9o15QC9XdBj4cKMay7wYWHgXiliW2eoaNg7+TlJYVw1yKb73MbngAb1
/FbLFyKChkcn5jTrqpYNpZdnMxTpNVeDKZLEirMkYTnDHXY/qEKZtfP10m/W
gyMsuI86IlAltUc5QO/lNid/mvcQTEhahb4yBDop/Le4HKjlWsch1xTvC2Ok
Au4HXg/5d2zaKxDQyb+aGT9o6x1wNYKrGsinHHb9chLKqdO2ICQcC5dEhprL
rYUwyl+njOBNfcNKzro5PCf+RY9shY+/RXTtHSBo8fABZE8U/ndoTuNI6WcF
I0m9vy/QJa6M4trGOYk2UYOuWK8pi5OwJxn0GsSQP3k3E1+fB9dflkJ9oqob
tSWK1duT690b6GuJ2WhxzZs35112LC1lma/lFiZPBQ2/EBpl2LVCS0XSCFBM
YvaoHEgz2X2II5lENpZFDKIlpH5b6Jk46nL9gbpo7jD2Cz8BMrGXRJNqC5Zv
WHeFKltqNpyLnrmJhNrwSJq3yjGTBEqbICQV38Vu0hHkTMMaH96hwiPT5mVn
3zdYs8+15Fr4euQ/njyNJUpfuiXJtdrN+K3/HhbCZQozKsTGkkUo7hY/0vfe
FL8A+hPAZq+1QC8Stxg/GWLOa9wivsIHTpxqRAIxhfQl6qRxpaqbGenchh6c
WwJuOiu5kA2LGvkrsUq3+Rr2+RzjyqxgfeaXi4QoTk9a5wvdRO3nSC6dn7mB
gPV5RlxA3z21gUawN3SsVavjWXV4Jf6B2siRGAch+vrcFbfVM2qZ+zibrdIi
zVnxROsHAghapigYE4lQJ6R+nsUw0rfOOYUgInwTqVuoHr0MiBXP+hxIuAn1
C414NtbGT7VFXw+tf4vOiikrMv3IhV+/prPMxZPptz15b2PHcqjzCSz3UBd4
oM4DwGK+DcZtEInNDpn1y97XQAq4XSjgT1b38fPep/gu55NrjgowZqvNb6ng
mg2s8ZNtzg6npj2jZoiclHGL5aHnJsKp1844nnrhvjJEnzHJXcMlJlWwk2Q2
I8T7vGR7Gue6gUxtWeer4KTHBGhIytJonE9G3GmnxVveqA8EYq2HS8wq8Ufy
9pyql2NLQ8e4qWUpZtl9m3CO2krOuOoIguIGkX4AQbDurPS4K78vNhIZi0zR
vasbDUoTvZqd03d9rOnhEG7ozoWijslRI8ikyqBvFzeP0I5osYgoJCwDjRaL
UAadkj/vL867bny5/8fgDCkPQ0mKwy9wc9AKZGcmEbffzfFHIIbob28Quoev
KA38QyF/jwSlTghA1MHDc1JWFlaCkSXbDAvq/sWKWkG8qyMKJo2snzfas5mE
6Rf4N3O5lOnzwebmKVz3iLlwwHM2//SgxbV8WiFBDs6zKRYl6cjf+hfKSuhc
ldT0iEjY6UqnyLjGDZEuRphUjxzORCo+cpv0MCSEYjO/ndtFIKzC+mrbWF8/
w/YKMyFTVr8VQ70rujVSbL77h0rrvhDtFDLTxfx3VRQUgZNe97jwd4TR0lZS
JN5go1XxnHvrj0SlbCFJSJQkK5TfVQl2eecUYWI/p097XVySfrYOk/thBQBt
GQNaoxtwDFmeWDIZgnpTrvdEQEqULbXt1+bWdaPVtg+2W0nbscGoMjJ6HUiy
xkNu+4TDPl1/16UGKk8Q9q15W2m+P5v3qvz+JKU/jFuLwku5T0pAEtDgwaYP
aP4eac8E3CSvR+/qMPlKV87X8PLsPDiw23P71LHIc7e53YCXfOJ6rrWt4J3g
42JcVejUSTy5Fu9TGVKXJUKDaT//I0cUHVRvDj2/ivs4+ZqsrHkgu5I6dU4F
PPKd0lvgyZKNmGEv0kJ8X5ZJV2EL2JlKAsgib76VEqhXplGXqTho2Y+X5s6R
VcMRAcV/DbNLGFr3/XgynXZn0qm80a+PsGQBeWbadr+noB405QSmkfLSq863
rNPjEyx7Sz4tlm+UkyixZrYG0XuRIxJcT6Wa30HjTHzUq/bcBw7xurzSELqM
IXMDpISRqWVwDnWEQ0lkkm3elGMBoT7zBde0h9fM+cGpmkHunpvD2ZQaqFJ0
dSOQhv+qGcgPqUs+Xf9esoykODuJ4FzXIaxz3mISdncDQvCSRyjFaOdPE9bW
3al77xI4XA03ltiJuxOViyL40Yh62Xp7Lj7x3LoWCADzfNDP5eLm0rj9uifD
RQTnPLntbU/92EsySr8Lv9B3JfYjugf3rolrOS13nhTshhX2EwndZtCVxbMh
Hx+jAL1GwrhZaCd8Id1xHOKdupYVCA/CFZydJqCTJ7jfyh/Av2M64SouT4xz
bwEVkvIlTQtDDbRXMsv5YNS90McAdfP4qrX4FIBOAzdO6e/4Tf7698P4Vwhv
7dXxWVxpgwiJfwYg2cGqW8O98fQMgMAExWW04ePXp+GFdSkJoSZNh8H+Y0NB
lnHefMVPNx2Em0+Wb9DTU/3+ryXX79KcLA8nzjyKtzoxrxm277kEkXpFrmE0
ROyDdEwwCQkga0A3f9SSsNzS+2A82iWVGFFhxSzrEcBmaSqiKYndb/gPorGz
agpxelzmTYXfjLcvZh36Z30wrym/yeEvz07et7RKZF8tIqPZUksWs5xC6dGI
w7yeh5aQrdPEFWHY7o6otyEkuVQgKIRK/IH6zKtvVRji5VH4DUJjWgZ9LWs5
y4rZZ+QiYBx2kX25gbMu2T6xMooXkWw0O/znfOtYgnZM41AySxvAroX9B2l5
e/JYAnop0TWCCgs/Cq7KSa0ZoMw8JfJEr7AJKv+QgYu4XT6c85FtHXN9s/WQ
s3gIiS6zlp9Dw/HLJeDZ+WE42ccA10zEF4E1w+hHyg5jhMrK22HfeV5JX2Wk
XNe/eeQaOfoM3npdVvn4Kc0vm0UjKiUxb6S/8W/7IV7ldCUZhAopblikZoIT
8cU6/YXakLNNijvLs6Uz/1NjFx+3mWzZAPnxbnOikuP0FEWZlWnG11+tgJnz
+H2WsD3bfG04ab6SWWOAid6TTlosr0x4JIhDSinWP88dkpRmU97pALXWJIqc
UELdm2yvVRsiFpUgpurScSzo9vcYR0R8YIdHNQVX4jova0CxIbS6nR5KneQC
T/saW9HzOogN97bBt+i8xvFV/njgkKLMGwlanSC2E6QVZhinrRuJFKFIh7Cu
QKQHpiOHsGi/zCCuLHQlRT9hBDc8J5rrnIdM0ndxaeb6QoQ/RzpCUKZEbLub
yuWcEyhN0jGvBO6k0JTQXn/cknrkz6ZfMoVcTWj0Ot2WF35M1Fl0i00zQB8I
5x3O9dwZnJoIIO/LgqcEPtgTuA+Eb/R2PWwm1XCMJQj28uSQovBCXR8Nn5/b
+6yrHmoKdF4wxpf04YcrwOMHCgWfuyKLDJC4bCEbKgOiTUzBR8N26kgJxEAC
WKfKG/wTkaSFXjOINtLzCTOOeC415FO4yBUENNzk5wv/BHhTdJoV55rxdoPg
kXr8qonMot6xaFdr4Xf//BZIKHUIzDcJI7Qrs9LfSQYIpG8gAN1FnV0hYbnF
/LuBY11yKCzgI+nuZPlsdkgP6cGtNBrQPZw5Q2xcG8n7Gi2FAXLSjDWW9z3I
qR7IOsiSYFQ3TdSsJ1lXQSvE4URgWO8+RufhSwOrQ4GeFFyFmWhRolv9CleM
6cZOJNKRSZsDllqZEoguwt5QLS38NIKKBbKkxVnBccFad3wXOZHXO2S4xLQ/
nhHVdhI3oARtGLv5HKG6QtysLsZYyosY1UlfucsuB5ye4oUqKQkMKV4EAOoF
ixkbfQl6eXH/sAbCYvJoI7aieZWVVhkiG2UFXRhZCnXER0nST+AiwPKNz1YN
425GKLP8e8VWp6Klnse4qn+h3RGbLjFXRVfLU0nmxVcCDdjNmK0+nqf5I3w3
4U3jA65IIlQ+Mk1TmvvxAA/OCTss/ZKZkxHM4NCBwQQozxmIVlK//y2d2wzJ
YyCvR+N3iZl/z0IHGWzddaDNURaEICaYtog5X3v4uqPJqL2xLohZKAhZgZcq
4ZwFiJYbEojKPdcsJ39LlRmFEMmsO+v0f2161vJcAQEVm3L9Gc/lGi3JEhNz
qZGtTuS+GtR+5N2Z0gqpddio7elrY6z1VQRX4XuLuc1V4P1R6b8y0PqZp5VQ
CxySn2gl+84edUiR0E34fDRvjkxjKAWI/Kqx8B/5jBp5FG14CvjQAbAlCRL0
K/T7Gb7AnFcyY/ahoWrsfs3sjF7+YiL+AXKI3lmehJyYl1ezCHNdk9Cq4Auu
eCedSqg/WXiEsrMq/zr+bs/VeHh/Y/soyEci7Y/y8lrb6s8iZjRF2fd1r8i1
m8gGQDbhLv+CpAjD4H/qKUCIO+fEoxUX9AOCaj4OgfViX/MM3NOb9zNWibL3
EnyvX+ZliT3cnJORtb3GG9tyPYl88zA69N5ryFFYMm5h7WRz29uWEip5Npad
rfRrV2Cv7aZT2eXv9e/V/EX75uzclhahCTXmapyIuMd7dzICU72XTPhSXeua
AE5DmMd6Nrt0KOBU5r8RQgun96egc5irLIqu5fibiFObdZt1IbBmQtxm81pl
P1ZWINfqgEMrBT5ypy7Fo5VEsQn6+wLbZZa671iFRsdxlzZ6Vaqu2l5+f7Yi
U6mdHTcFdGMYYpGukBfLFN6LcZ2S0aH8782Ng8bDcBTCJlDsNLX4+MBtEQ8I
kTeUxDcBeIX3rhzSCgXYBJ+k0ap8pwyLHZbHoGffxg2toj3Vao4+q+XVyKPH
rtTIxH8A5KTHcSxFKipoixdLkktRHgSTeYPkuy0UCBPXUgMdq7i/33Qn2QQJ
msr1re2hR+kWQRkPiocGJNaaG874rhJwBG5HU3Pf1nFqdkCXtz5Iy8HfgMU+
LtToYYWtcpvGnCa662g/bv+U5PKb2yyhwN6fB31Mul6QSzho02J4drNCqRP8
K/E6vyZ1BiV5ZdIoPxqwZ5gF4KoKMzQn6S2YRvL6NuOeVK2BxsDQcT/xRh0O
NltjAMKDkmK2jTOVP+cF5DXqw9qValkY4r/5m+PJiv6QpwIgAG3mCM1rIBQM
yq2/QCFcNMummcKUtMC6YcQfZC7wyCCJEBt1AQ+T2mdKAMaOlzPponT4B+7q
el6tLOI0BIaQd0f7bDwGqLGLb2V+wVjSAcbyuLTIQ4lF6oTJeZnrhHS2Cicw
5zSk7L/W/w7w7S0Jd3pj/6ttNOE1LOm2Fcp9HAFtURQE4m5emnFUX2TEwYwf
k6bw7yjOFDFB90TgDT8JuxRWxO8fEivAtWUidw7UEl+sHvFzkxJjcUs8YKwa
ZkYf29ovK2QjDFK/IOCqB4xEl9OnuNPOFCsLgak4JuHWRMjMAv+ntc7vlu/X
X5NdTJwkq5Myk8VZhV8Xd2AAZixI2JP/BvA2NeSLmj+TlyLtN5Cr5PsZSHof
I9IeYdVlxOruk7VX772n4NoG+ljrZZUhlFyRFJ2Ny7wmVD8MikTYYp+3vVFG
VBnXp5+wsJcV6VkpWvaDJMkF/arDaprZRqeUBWUvtofX/LOf4iLmNnO2KzF7
9j1CxR+9Vk+8FGyEw1UQQF+E9htxQ156MW2CyuMWjAt2JFgoe2Wz9hPJMFr2
Fy3yhkvMjWRDQR52qvDGwzGM/ZMrRAVGd+EaTQp++mcCsayXV/mNYDqi1MIq
CwMaCZ8ed+65C4NWVkvOD6pXdS411vLwMPv9ObwVSusXMsqkSP64df6PuaQJ
ABnNS2jsc3cGZA6roNe8j8518Np72xtJLI/AlsvegC5qKhexIGqVytp1YFu0
7a44Jl3DzzZz4xYHJ3HupFAB47o5B67YFgz/eCAnukT7n2b4W4I5OehGD2ZC
yaqp69X1pa2oXMcliQ9RY+uquNkkNAa/wmxX2D1ZLQcQuilMJH+b0fWsuRLA
06fhkUdVQM1nlu56q26m7nTpigWw02Dcw8Rkr805l11XCSntjpjOBisHDW4d
geFWst98grmo7aC9ypYQOdkHYX6qO1FwwtuZOXEd5G69Qm53ljE467z5ISBP
kAmOJmxGMp4h7rfN6AEcPS6k7iV55xfxGf81E3Jz/j8ZBnJrF8zJjSUOaLdX
CghVcabfch1LlxJSFnid9ixcDdcxOm0VW2E/WlQCb7cQWvod6YZwaE/zCdRa
bcNzEADByX1AYQcN+Jpt9AQfOe7N3HSd78thf+4oB41K1zI8g++Wgd8MeqPE
XgLbTOlvx8zBaJvMTszUjCAousJMHIJR8x/A6q7k0xJV1N64rDLACWBzrEeg
19xrW6hS5HlBM8R+jaFRKd4zdVgoXEXoUCpe9vF/zprVEIuEzpna8/PP4nW/
b7jwmdZm35qMB73tAT1QYscpmX/dqQEBdKXz9tg0RMq2FhS1KgD5mwLJQ8tD
k52YpgC+pdwTFf6mAUXVJMqtW9V/jJcVS7vE8t4cy8HQ/GA82td3IL4gY6kc
16F2xfXxfgk+2GZjXReSJdkde2ou/WdE1wKqEG6nSo0jII/cubm2O/Hg9Kxz
/U/IoLuEk3g43Jun0Nnv8t/l5c3q9xaV8gAD3VILABijRP1Y7xh6CCznkQkM
fvtNuPlalASch/hmULsQLU40oK/l2DHVuZDbULJE/nzyRfV8U24ELfN9K5mz
Lo1P5Dh8i+5QRLx77Q6iqyZsAC4hKePLglFQPppabjSTPTrmtqLRvjVIfy4C
UJwj+0oWl3FsCjRsJuEeTeXohkdiCVzYPCUbwHPiXZ7JwtUkUr4OpHWZL/t5
VlqbTEpEmITqgSwkkcuBQk9sjGb6n94lSxOFzFkwGAZ7Y6cpz3ItjJYvFGSF
xWIBgkKmNJcCTbxflYqvpwjQBD83+A907OECPbP4R+hu0cL3fmrMU9fRlrKN
C8OXMxooKRAxbnZR4jsJV7jw7Nb9sYeJuOR8daNpFdTRughOVdXcB4/uIDJT
ts9xa+j7l/h0hka9H4maeC48I3QsmXgHO1ogqyjrTulSGuQPdTIFyi7+8nnO
uNWiV+etS27b8svOsCW0X/zMZ44oaZOlMl2dYRompBzZxnKxocCbCbIcQIAd
T9fF/wtJshwjoPoZ9LpWfjv7ZX+x3rWA+YdiyANouCsi89GAnhUu9sACPejV
PvNVubEIMHn2twelrHTS+1q992xKzuuzgiB9MfT8Geqc/TkXL1gOBIZqzN1b
yggs8FaowG/+FS7w5YcoHyyAHY3JZ3b29r92Eia1Sx3LXsnVhHYKHlD+WvVq
9O6Lsnfu9j7x1EveEcqOGPXubsfRe7V7N7k2dRZQRpnGr98uJAA2C1qhu1zr
KtIERC9tH+BIDBCnxZC80BQvTVVn+Ocm7o6OF+qdWvGg7vCwHIhHolnz2H40
EIYv5UTGyJgJtfI42Wt4QX1DSdGGH5hHtpFGKY+5zvNV23lGMaLcwz5Y6Mqs
96DzJe06ZSLgN7PC469S6djZFRcIhfWDxmIQUfw+X7mrlLD25SplikPUDPWb
NRHHRmhYFSZQ9oaLp7WBNxlhIjZQFtu3x1a2g7jvYrjOn2poTeErZaJ8kYgJ
jbkGmd72RKDIeB/Vqni629pWVLmeOhe+beYIxISIa4sVQpsnsgp2VYX5oMXo
GLZTtA6/S9bHAOW31j3tCMJXqibISKGWxmvqPrVNOQz3FSqh3Mi7hC4Wnm1d
RSAJzpH1MoNkeQApi+vlYOzj1EZPwYmRAppWPfDFbIw/dpcbYozxnrqYQi9+
IwRdS2iFjGkNATsY5HwHnvfjGdgBIz+jo0UgMSkrOVAf0B1kd6d99dJ4TZt9
4q9SEiWcqvZDqMNpxwQuBQvTdNonXG4vatmD4WUzrPoJ0zLIqjv5lq/iRUBo
GFG73hAPdYQtEn/Pg3XTtKtrWssb1IBNRyPFZLs3kzOanCJrnjL3czsKx0F9
RbuEIQ8qJWRRmftDaFQ9bpkcm1R7GulIoIR5KQe16yQ6pqcUo6pLEqDSaBS+
xx1m8ODvPkytn6d8yQ4G284Jh8d0SOlPNha3LkU3Zf4cihMaj8N550N1p21W
HyqwDTMHg82czitdo7ZVn2+3RiCTjiT4egwAVsdpp4HMFo/lvLvJQXqD06QD
BMt50+NS0O86gGFl5iSaCH/4j3Jgv4WROhVMvfLsVe4aw6kWfZs3/3tEktwN
fjjUcHdnv9Pa6QqG8jNPouDiMA9rA2Ov/E9LFgxXq67iLAreuo/ts8G1VkCN
+6NRmw1Iudexd7xtD8uxS0JgQnTK4y6Ffnxjcc0LFGLzeu6q7eB+dweDFyas
VMZVzFStGDtMBMTrBcS5QuG6ruAF9ytohEUXcr514cS4BKhPbimerxlTwPxK
n8pAGBcgsYMi6t4klYbxlqVDY6B8BpJj9UcHD/3xS2Ru58txcC5EEY9rlf4x
sg5RBqgFfiLPNKt8C0650CkC0GFbkHYhR59Z26EyMsMrc0Pwl6P2hWMfkUsS
UM5rJOsBI/dvDolJSqmrLn/GK8gib+hv97rxhs85k4AcwBvbwIh+M1wDr4nF
B+jziRL/c4USo3rQnRoXlYxHr24AvbQZbJpkXE46h9j57jgLgDdmD5chqTh2
SSRXbc8NODmlkL3YU7cq2xK6aiJOR9LK9sNuWQgwPqMpXeKTegVSuXYWy5gG
Ee8ukD3PCiLEigBdNA3YUeYNyXCw9n8otB1n29rv+F6B0JDfA1txRkL5j85/
XnrN2C2uYppa55ZMkl17BLPnfRuj7efU3ISnzccMjzXJbvgUXjiLRjbAHROZ
so0eKoUYZg1FVnuZHRzK9Qiyqx2k07l0UgwKD+srqwX763ZOyPl3pE256H3C
DUOONIQ4q8q1e6BTN7du2v4msYSThRTkmMtH9rx3UYIBQOeyAAsGw0vK/g3X
mK3kHvv8miIuJmLZc7sDgGBaD/3MREOz6Dr029CqPx0cDEDWMfz77OeTTnIb
xWR+rO0/afMF0c48yEj+Sba+mCtjpEkD4DuqU8OmmOSpm1rmE5RiMt++m9SE
7dwOv2tn41fB+4Gc6z3u25srsLEj+GQMsUeOFVrsLn5EKsJ6gS3Pjt+NU92h
I+eT47DBAJJo9De6/KsR4j/50Lm8tQLUosV8K5HZTSFnHzlH4WWIsJ8UP3/n
teietxbb48M9TxF/1M2s3nME4wxxFDF9QmjPb7i4ySKs++3DsBgPpkyYI5a0
yub0noiDYR5EbuNWiZ7HUFYAe7kMwvmQRwxHvaiLUz4bTIHZLjh2wSicj34P
aRwJeoAPiNWCcWTo82Ms6/wO8Ue1iGpzS4zJ0zfcfGPpt6uzTNkcHXGMrItO
pSWU3Kj/1KQdupHDhuzhkwuZeAC74J2yYRq8W9KFZUEtOFHTApfj/sfDJTHF
HYLdpzSEEjnVRU7xxeShL4YH2Do+wQtb6IIJjSZ5m4gPELo3ebRzWq8PxWE9
ZAFW+Kn0nlyyZHqHpke7c4CZsVtuhHF/ofBNakUlPhAOKkqZTLt5tDZqaG4x
qWYzn0qY1yIqbZ/uRGlI+ix+H+pzDcrCQyqvQNtX0tMcaFX9qJabiKFmPsMN
nooYWQbltHTY+LraX5/NPpjVwrn2VkHcqxWQUue99ohlqo6mtzNvv5MGVU4U
Llhu0mPBAGCI0KzPIBvJA1Rj/892SqQCofFj+DgpIUzq/wb1UiaRVWy/fi6B
ndIoVuSUAS5pYF0r6Enq/eljldMAaTprY34qT6YHRzCm7fmrqxoTmgCc3sxP
R/Dkpq2W5OiVk0bjXwxhSvj13ZfPl3pPGYuRzcpNezjplcoxWEJb2+11iFrb
y6PXB8avph7CjbsEmG0MjzFppa/CXnxPcCEPKif59Hs5ER/3Sv5z5Ugjl5ML
CE1gcLMZbvwSx4Tn5FotgaV4saBqViHod2WcDqDprpASGFCU3KcZ9HUFaojv
wMofVCNJktoYTOGmPA+j6nWrOK2b1VenSAaxqXr3eKMiSrixt+xu9KMkBqQX
7D5KyrWs7eU/afxPKQiOaka8HvsuvEkVdvFG0+A1rz3LRBVkxIv/gwDVkIiH
WdxYKX9VWqEAAKLE2SWoPx60rsBqBUQF8zmAvq/OFHf+GKvL1ZHbsmYx7lBg
sKBOwIYYUY4Dl7GL2QOcZZtDlTPFObBIPG98TK+S6yXDFC/Yh5gYwtKgU+Nn
bL1y7uKgE+uLrJpqJrytZ0HgjNXH16YzgPp9b8U3s8RlL1N0e/WwCYKRx1MW
EwVLUSuE0X6vJyFCJob24I5cR4K/L9q3dxgmgLaUH1jAdD0a5gomSO1hBBvN
9tgDu4+60NR4+6guuu0Sz98Mxf5vyl26npQFQCINZaBjGRoUu+6L99/DbDDQ
HTfTTkk4yqaELiwhbWbwU3Qfc6pOa6gnkvx9vQ3d8RxTC71nvQ8mosgW15p/
osyZANlOwroq+Jzrw68ngs7KU/6CVXJvSUirggJN9p7aHMA+ex5nkLBKq6bb
2ZRJnPDhJDWnPwQucHgBETDky47pe/6YjHd0bfxXEZNb+hNV8zL4Acf/uCh1
csWw7VzgP5qZCUgLue8gytba971qtpg8mRus2BXKsUQsDT13pJom5qZek0nK
p68xszOEqGz2kxyOamT054elc2iC2Z7idJDGW9GrQRv2wz3qqZTOtZWefoqT
ShuSevlu/GI0uYJR1EX0YGi9crDiwt2hcMhCFeFw35HrcAxGfC+W6wC/lBCe
8VILUMlqvFQhjTFE2etd5/GFdG4KZVzIBBoqR+2MDQEuziLbALwfXJzoYM/P
CL7Z0IDaicc9yKHnsJHH8l4rOSXj34kfpowVN7MUT7CX4gssfouzUJrhGWAI
myjslAWp7sgcEil6cZD6/3EWa4n5KcIlclVx6fzAul2Dy6QAnb6UkdVsyaIU
kF6e4g5iYeeDKLrHd13V/s90CadJkNaB6WGdx1Ob5Wjeo3/cnY/QbKjqMxVc
zP2Zp3kFQRYvI3raLSCPkhFkJcPJtAuEVzU8OosMl1GC+zwP3cfToD70nh8S
CqpxtBBRaukKrJTtx8wxKPBRDr9HGSrKn7EToUpYW9XcVfNRcB/TobT0Qv0b
ABqn8E2VnRM9xcHRqiQDDGSZgIlny2wb+vDMBXvorrx99lJE6if2SOHY9pkf
db7QYIj/UXtI/Ia9ME04z10j1WZ1oaoNNB/6m4Oo2Ym/tr/N93ehyCta1ygm
nD4M8y/BII7VdX1ASq3WV2h/JJv1YD8HJrAD20cDcazFa1hHDSJ2xBMdWo8L
3gZyclE7Y0v9+ddE5yNTpG+8qlsOhGy/aXRuihtyxC0pjvQ4FQ/CcPsfjiBi
Zrq00+P9Prz/ZBE/ZkuJ5sHARwVHWjXv6NXJldh8J1SsieqZwhxsvRbZEEZV
KLQHFjq2CuTl3gk5mbqKF6pf3fEz9G+7iZOUIzEVlZHSn5SMVXxBxJ5iX00W
tHKguB7vw7s0zSdKie7FK4BgPtWzMtYPQhPtFbv+Al9AHl9tsXQkEgdnmmTW
uCZYaeRGTAbrrYsGIKLtuEP7RUZlDaO34Dt9+scivFEOyf8qZzX+XyBWLmu8
aYUCiCVjgMUbQV2MkgSXkS1M75Lv9eMOBh4NQoZNqoDcItcxesiaJKRewRNO
Nuv4esaQuphy1/6onJCdjr0XDv5exdCiPazUIYRMEhDTXi22p9gTBBya7gy2
g37k5XbkNrLyuZf99T4iTy5NWFuKTZ4IFh6yCQYa4w0DtipcTlXDNu32/cVD
mkUWi857uillvdUPjKcRxnGk0dKRPe8fcY9ns/v0LBDYhkk2BLUjPhU3I1iA
PSs7swyo8ziKkmelcKosuizoC/M080ra5KL+a6rTdJyvbsGOYlMrgrbKER3N
mrbKWSiY28nfxWS2kfgGIEy5mTO+zN6+MCdBl2u4O12b4Xh83UnF4KuZpFNs
etYKeCh/NhhFKKNkSaXFqncSSP0OwSAL+3QBhRHTbzrApjIuGH4soDoyMY8L
mmssGqGkztsqvMejURmUgHK6Lms044UDZETYJOYLpDtuk1J4taYBDXqsa2vI
udsE52IRcOWLLCCarY9TgU2cCxinynG5ZcBMBiUF6AjpE8VB/hNqEwpPXe4w
iZBmykVQF53HWotkCQ57DNYbSQl1/B34O21e3+AnzJa/vSJdrbakOCbFkIR3
4tJucF/QAfqzu6XEiq7q8RRriDFPSRM/jvWvaA7A3FUtGLBir/ks++Ofq13S
PDIGIa1tCY/kHe8L2dskqoCeJpaMvvB+7TN2hqz32qQGb10PmvRbeVA4x3Up
fupZ2HlfYGmZwpN2LAGJkziAbE4ZuaGsEkVmz0eQFFvrwJbjmeL075n3T2U6
DDZE5WojdkhODNY+VICTKStAmPd8bB4ACrJ+FzbltUFckXXoBNu97FncI0Nu
mafi9NKbrEA4UrMqWR1+YopLSYInzlM2UmPT+j4RY1zaRklM4uM1sISDmfUK
WAJ9oUf2QwnmIiNXCeBAUlGINNRbkkJPf/VCJp1ERWzhbhByWjNde6f/vZuB
w/otDVOvHA4bhka3Q2KXI8SgZh1hRK0u+TEoA04zcOiqq0Fm4H7cbIL0oeqC
yWy07pozqbZ6N+0B8TADyoiTUe2P5cif9gfjlAkw2EpfS/7HpsVV+XSExFZa
lsF/p5G7ofPcp2EG8VoRf+1ppOsmeDIfrjkYBuh+uvAYw5T51la+CMCB5Q87
smieiZE1QnV4510b9kYNLVglnnCmpmEuVgICZwzVbRePo4sCSc0+J6Izs3DS
caWJyRS+BzWtF2AIoug4pZZ3Gt0L/1fsrQHkM/7qYbTjU+HByiIW+Am1PP5H
zX7HqTR5VLBZVOy9DxMt9E2yXFH0ucrxOzwfrW05N84yO7UBALtlunMA0OHi
MiIfRDxlqNk76IgP+sD04LXxzMhjCMA1fO4xC4N2ceyPgmtv6LR2q4y1+9qY
HtsBffsL4c3Nm2hVB2aNB8UKVKqHaygCLSZO8AfTchyNeihAgESsCvCGcVNA
HsoBY4NVPPcaaM9N/lUqxbM9Gls4VQ9X+J6TNA7Dd/gQ4Ylx1c+l/9SWhmvK
JvoeUo8XWSZ+yrpT3oOadBRwXTLNXx9D2SJ60b1lvwFVFwnstAefGVHw8zcH
d834qg5HUgF67GFbkbWqElaK6Zldukzgjo319H+rNahV/uLLhEky7hqQdAnI
66+8gQ6PHuUdFns0u6EChubIwORazeTwO7Ms8baobsp93tSeChWERyf6QQAW
7jd/xqBoUJmPjMaddvZ4HwJfgbCmf5egDWLBNA32MVXKHDz31LP33UStHyrd
harFnMtbNxPM9X6MBUmwrQzE6F9NhCdha0rLHevbIpwyKtPmv56IlNoKkOik
xeMz9TznCivCos/tagvUKdyGX/h8h5/pzyLfM2IOwwzRhwclbHKpvdybdNlY
0N/foKzcYEO+1BbbGWIgVpS3u0inNE48p96129tz6lHS3usQ78IL0ouRrpZ9
Mfe4ki/xCZeWNgGFHRxIlLNKPawVWzVvVjqEzb3BPd+GPobsVsLJ8cyOG1Ry
21To+DU6xPtDhCfhSg/8OYacLmJCVzo3JvP+NF6sauqIWNZquXrVkeNaDdrH
f2x9DZtgoP44nsqvgJxmlxCIijeY2QPIeVqMCYvIeYgT9T6Ixq9c9pJEEgdo
n9xgh8VKdLSDWH8v5DiOJ5GeRjZDa6ocnY7DKG+GEheXAORuJSXd4RSw8i2O
/MvjoFaxAmWMZPmdqfjNWPsoDgilO4LlTnGzKiiY1UCYYgxOIn3/x9RUG2SF
6PWVWWb6LQqYBW7A8C/9ldIPmc5/AyujKWbDxny5y56vHv0H+2exjf//igY7
2+paFDlu7/1OJaGfsgkc3R7iGDGu6PW+Kpey3a0MKH6wQvwYMUfDZM8Cx4I1
xreJIsahG8BDcITGqQNTSydEfqOR7fl8HGLyg+zqZ3Kv3jopHP+xuzkfz2it
8Xzq9bB7Y+IP5lNu7h/PoefpP+n65UXzVxJ+P/42Ol9P5wW0q8r6I/h2iu23
rrmbPd/QqOFNVIFN7eUOQWyszUuSe9IGWWukpw/cUBmjWOylTmujt0iHPNe8
s6V5FUcgaUDw1m5eZDpsUwKjmq61zGjNKvJS9KHFRRcDdZSyZMlWVJ1QGRYF
06aFTHP1vbp0gDU666C4usr1dyfoewm1/w3SEjC/Re2pkeclyO8x6w4nDgbT
pCxWy6GSVoRWC8sEiN4pTlhnpSbAS+93SGfrayIEI91sRJak9pjri8E/cCnO
PsC53cKsQNTKXTqMpDvICSpHsEO3sZfUWPqgu32IyhF6Ue4ZcZQLtK9rMTqX
i1Td80keEyv3pow5RdQcqtIaA85PpqoYi9enfFsEXnrpS5y5c+peI/ppLnP+
PED8lifMStwT+i2Byvda9RsXkmMQTUQA6c2GGA1TMPMcqs0fpnM60ASTUGfE
q+fgIa/Am71Bn3Zy7yHuII8xXG+hKey1axgmC9oFy3KsgG/pwoStDTEun+sm
p1hHOn4eQ9GQh21b22my09Zyoj/JBkmmeJChYWIxAkbbKO5/a8HPMRuqlB/z
PaPR+gOHK9CcHRL2qDf11Zk0L5R2ae5KAyF5c2a5s1CpXoN/Vo0eHMxIBH4f
JVlJZYa2GXpvVhY/Tq5mEXby69L4OBAJKOVySUfVTPLy5p8xG7zl3vNGYW8y
7lJsqrxiXd6qWvt+1DOs/8slX8LAddgpeVgIkfKPD0+lSEIDdkhzwSsbPLH2
FOxUTE7+dS0WQy2oeenihmW2YcVMApbut6YJep9UMGGjxIdY8pXduuGSrSZb
u8cxAJkQSCfsChVdwx9WllCx5dJ9KdGRGnb1lpBbQfEU88xxmacQ9PkBBj0R
WU3CS7uNwBEsMtJ0sSsnbOZaFsqsmMvRl4DZKbfCTPy44F9nVfI7nsPvK7BF
gwMHEP5UTiNBEBjVTG0y0qzN9VPU2+Pbuu+ZECNi+3xeCF9sJ46IXRrfyQDx
FxJVU3S5YZrdjSyHgh2ZNKggjxtTHNGJWt3pQWnVjPN9BsaBXU+f0ICU/SW8
icD47j3+dZmPc/LLIb65lWzESC0gyyAlLUI63niD/PljloHsxOSYI954Ck9H
Xq7jyb2VZylSH3VDcKDC9n2vKLKh1iKGptVp185nLWKtjeQ+JjE1YhqC7kBa
kdsMGkebB7E8ZfZ9/5Fq0GPc3lex4sCRx5T624iRVZPX4SnY8u2HponTI+OB
9tOUKITLZSaKfOd6iWFL8HutZk3sHs/cQA9Q3qeObdv/FT8uidxAeB4drYeL
SFU1P/v7pcZ+6NPOkmyn3HjmarhufkkCc5j0vSHesgHXqlkCUlTJ6x5noO/R
wD+RQB4RcJXyHfDn/mLt+hJl8g2ERMGxlp1EqhQB8SyFDK+a4DOqACzGiWkW
BBCdf6yxEEgIwBCs8djyMTZ3B2SS0/VIzqzmcwprtbZlUQOdriKFVuopp3Ad
f/uJuyKtSpUes+qOHtwMJmdy4U55O9YSW9UztpU3s+PcfxnqYQ1SSXWDTUK6
nNw2R1tiRZBgJmA0dMYbD5qqP6qumJp2Z1iwVb3Txx/aBKPGNY5kaECse7+r
WHYxR5eShQ7D7N64DNTupYkyw0AAvsNoeZIr03PYQZes2vFqt7MSLHOO/NSa
LcuhxsuCTrNYEc07wEeF4lW1XBJmYIq4HRsLeYNS48F1hfcV4kHg9YLSR/M4
WO6T2YJMNdF+hZaIJygtDtNNdYwzKDufORL2/CFOGAFnMF2KpggZ3pPZwuxo
td9+NAL0FQWN+L4HQuU9HpbYPh4oqnLHuE2ckh/kQ8aBEU7Ptz51Fgs1ey9a
sycOzdvFWq1urEYDDbmMB6XuW3Nq03h6DKGZIlk35JDAMeCn14iNHwxObB+b
MK/QGrZgf0golSBan3GevJq3ZNkmLHLEugrKWA4f09Zgpd/T0CtTLkENJosm
QZjlLHuRRtQmFbw1k+B4JPZJLnAZxKGF70dsZDKF28PzQzAd9AcOjJhPF6h9
/UIKcjWcC8gci25Y0FscszYRWqmvLIcOxkiLpwKRIBmfla+iZu7rBBdInHPX
HgbeQyL4XLaTuQNRhp8p/hR1UbdfV1F3+3xZVpB4cGEbSb9cDmdeCLxkNy3V
BUBh47whveBHzVmEbgSbFow7wwOXF2r4OEs0+mYTRBDy5CbdIVXiSj52izHN
46qStupBRDiPL7m9VasvvWwkWldf9CYzdGDaHxhkXlzLJ7N+UxDhKld7lwqH
6TEketFzZP/CNFqreSOgHgHS3gLlWIx3Ts9db9L8lHSYFOqwKVMjkJx3mPY+
jy3/8UC+1oGZucxwawigDOnbcQIpfO0qexVWpKwnl9jBOYLbTZopqHmrYtGe
RzlRmZRiiwLqoCxgz/c357h1RsKberClCj8QI7lRThJ8NHaSO4ZYwM2yPyZf
UU+m8B6rkwzMjJfTdkPXWViSi6J6Y2WnevGNxsNDcufdfvINJIfswQUjQcPy
7bQ1G0avCNZPgHCCRFSZq6Nsk8nd8eTlbwOcSXt4OISftv+qYG2yOnq8ctJO
QgL/vedb+yoEWrZuG4fxbLrdeX+KZ0e8pfuSnNcg+SvF+r7fgVL989EFaLiE
wAOWzX5Yd2YGbmBbhk+AbadEvReITeKGzIaeYN9YbK+yLRV51QJrIlLXVaVh
YadGe5OCs+N2c0I3B/kLH8K2tSOcwjIo1M7qZXa2Lsu5lhhXUJxh02x7Oti5
zXcd+k+6dYoXY2VK+iinTOq22AlyZVwLRwFMBtnWJikOT+C3QJ8SAVs9x7nG
xBw4Hz51Xlkrf0XtVjdrgI9C/JQQBtEvfqsFZes1EYLNcuL/0r6WKQwObhyD
1I5vaDV4OcZWcu/INa3aP/Xfu88wmMzYuu7sH7THs2YJSn4LzCl6e/g2O7ai
K+JWIfWvgAMiz/7w3eByT4eKdgmp4plZR0AvMks+IIvUjqYOij9aCMtsHXGS
+9V1STwFbHBejl0co6A4sEMJZwaFGQDYWLaZxOEp4DltfL2pv8mGWDckDw3O
ImxZUhzsZP8Gr5SpusgGAbKv2UnFxiCmgCczans++fSPWRCI9ySs5nkQjfWa
SifJxEs+yDoGTuPIpBe8W7L0Pi/3lkAsPkOMyhWtybaz51TBSA/7sKYTFEJZ
19jAe1a+wyXKwU4TLkPXryMGhIDOT+/lLs9FYkTbLsTSeTIzjOE/JtJZUU3J
caJd043kuxti4qeIUbTiJWD0t8j2qyHSFzAKc3zuuqngegRMaY4qUMcgKHiQ
sP7I03El5zKNYIrusLm+zyD0B3Tah8UsvpIgejEpv7kjxnUYbZdTP2pL8GAu
f7J38/wA/qThQP7U2PJ6ZSaNOwWHinCz2zmoUuaSji1DNBET0w0N52Yr+ev4
lS4JnVJWB/UlXver9cXHH08BbDz7YKLHduclI+2jKqbpMeN53UvQT4geyu8z
pOLU8re5IlMhYsklcbWXkvzuZZ4wLXks54v9JWwk7riTyzFa9kSRux82Sf46
Ef3XzNNW6FM65518I8te6Slo2r6cNhR4F+jDR1+M55uFjdbI8mV15kN8Cmbs
m/PG74dhvQSBp+LOYAPa2xA9o0UKVq5iRu0STPaXBHkU65L43eL2JZz9uDGe
uUSyK62EQEzyufJv5SdjhMU155J7TjduCqBBXS2/CLSPcuexGtDQE8qgFIBu
YaUaWrUZjYQoSaPZz9JmW77/b5fqnOsw0+erm6lYs+XMcb10+FGwqFPk/i7t
9Fh0UrpcEoqvcQINnUBj2urZIAOwI+O855lqVImRa12Tx2LlKY9kr0tPCI/q
BH6rVCx4bFWPnQ14XC9Cz2RMagHyXP5G9a9Lnocu5UE794bPM1iEf1kbD7MG
pINhTG6XlJrFkJIizx+l9YzSRvxINoUDol/XiMoHgHfrbihCZcYILuib+LRH
y+mZ+gjCjWLzCNurYND0vRusYOuo2xMtucHT/EJ8i3DbQY9/hFXQst5lTETx
HIg7E2WS6WzZntU1sC+BBg3/fQej0cKG16VWaO0c6aaduS9ZezV7gkVUSPCH
BEWxYvr/laO/lcV8lVMMkbvapSak3kQsHFq6BviQnFIWlq2YrM9/u1Nwp3OB
9KrkO/8wnzb+cEg3hcUepMca0lBi8at0f8WSWdt2DJ0kLdhtJ1Ndqf1s4kgf
Zf4UO1cFF0N2Znsyfelky7isBy3HmRJfGhTWeqv3hOxfDMljQUcBJt0hTtCh
zkf0bf+ZDS2geDpMVdMcrrjfKUb4C7i6PZ37puPUYJmdCPflt8+gnd/f4nyJ
5XLYrOH0NB9YLoebGCn0GzCt2wZBDsjvwSHHLcFxJLgcuZNGj5Kg2XfVCS+S
fwmdZ5qcwi/VzdSs2PFCg2pkeqbKikcJL87Bt13YNmMLOnII5hZ+T/Ty6Rv1
b0U/Q1UqGyQxqlUqqk0WeR80stazgW9d6H2HS2KDGf9JeGY3CuqdyMyBvv6Z
B85zzG7m/TiXUfXy8ocsAAu/vrI1PNnSv8udiQe6iKKZIbqImnh8mTwVI0CF
xtwSSqfT/CszHAmWnnZpClULxvAe3M7zWqAh9CKxXK9z88qY71PMowiCgpcS
06NzPraN5JlFqeMfCcEXDVe6EbC38BkCUYAIcp/GjhGpc+znx1mUzU+iT5d3
hPMkeOVxIoASwMNhhUUQe97f0mbI3lNjRvWyt8r2AkJhpBWAfR08+4C5lEc+
JyMAEh6stitsLwuqNCVjiPDjZweL3F6MvurBn5ZDTtpL6eMFXjN52lOH9nQL
BQjgxMKcF8dMjzbIgyVh4wn/E8Wvzv/tVIn8Ns3l1oq7sDQbmQNOasVv4nfU
uKQXzwAwF0Nqa5EIcjglFAIuYl2o+CMxDVuTXgKjqEmn3VcwVIqfHSuJ+S+o
ODHOC21fjRIuRBIhg2jgoP2KecVFZRI2hiEupQIqSNY8zfXfc7Grp105BGh1
9ZJDQicH87XM4Nsvirke1h3VdUZZQVqMM0cguzRKPMLGIKTwW1He6pw1JGIl
O4K/V82EznpaSZKoSy/lcq2qmIwPavA5J+UdD7L191T2M48W2zhHH1f5TS2d
roWb/baW+DeGeoU6Oa0XrNTwawd6MSW63QLQiVTjFSCm7ixAJovT0ZtYG36S
NUpW9y9tIgRc5LmOBaBoq4PIuTNgDBkuLFjxp1ZzI3ybDGdC0QBmZrpD3FoR
KMPVRjbPRgVKmtmubgS+xAjRlX6qGAdGG/HefZN/TUPEa+ZcbR8UficA49+w
7HUQ1hL9/1OjFQHuYMJAZPY+LcuOYhxNy1Jy5fXL3UF0bF2N1NKSeLdbTlj0
ypRD5Q2GOFyA0oYhqXZ8udFPfPsCvYwSpTW7FFBouZywkKJBScornEeRuyGt
3RjTIwwpvoXRot2FV55weiwjZq8QTibqKCNBekxKdWJZs/IEPt8R7X4j9pPO
GcTHU0jOT/UQNN7mBrLRmrCc/xT11tNIY8JLFpDv+aoJABnMNLNS8kXYhSul
IbSVdPMQtKVdZRUA69fAegx9Rvrwhai3eBmgJlD/BsP0bFCmRlRL9Oc6fJJN
H1Tr4XdRYNp/xTwl/hkiw8JniuDQ8BqH7nSPGLl6S7msFtW/0pGLtWiiEiOh
j8YAyYi3dmIB8kkU07XlFSQ/SmmzMPdOw+632JHpBNoigmMxEw07JWG2DxZq
xAJu06OWpVreA5QCSOck1lKgwiPTTH9bTWAa2LWQk8eGy8nNWB/ioivquGz5
XRmBF8aHApcyMCthsi53N3ywrnVTgLRSOulVJPW1lr9Xp2BvAIvLQo6q4+d7
TQh5CEpcAQHCfNzHQ8usIxksKhGATPDDyQK1Q6Mm06CqJkgiTN/V93ba56QT
deybgGH2DzOtn7yb5ucUHyLAtYTp0dbE/ecWBGA01kiGCeZThZNBUjTwDBRU
steW4nEBLktFbHIc+aa42ho8qfcl8J3QGbEHhlOz5lgoZuRLX3kKsAazMee5
206lKrwIzp9n/Ikct89L7yb9RFnrINZzwOI5/MnHrlJzoaQ10AZdJKcS1yiP
nJHlvcY8SNmIp7WmshcOU8SIbpD++hF+ON7QiFMy2VSjxWzHY0qI8gl8IP3/
6WEAUnaeb3dnL+dJK8B0NFTMGDsB7hcpa0eN1gwI6Lwjb+ksDX2CbyS/3Llz
DeCONHIrCSkwLYE3Aa0wyqqqiUanupQ0YI/3avOyeSt3ygw220vtNxbXCCIJ
vMd2dtdyG2J0J/rWKHMMIn+7OMr2+2/MUtlG2kxL6hxw75BaFcOCO9UQU2nm
L7xp5Xi8Wl4N8g4OOeB9gWIzDESFOSzwOvXGO/HstoHJrC0Tq/kUlgioksRZ
MqPlAYGqkJ1AAkpqceYL8W7gM//y/qMysFwiBt3izUmiCqheEI7PLoMmwx28
UePslPWrg9Uz5I3euaiTgxy2sIJ+Dl35W3ZTk+HWYVUGpW4Z3iOK9VzcyY5h
1xYrVfLemHC6CaSadIywJZir0t9bXMIUjB9Gk4/FHnEK3//fYgyXiGOBIEm8
gWQRdnL4z9mcWqBuNQOWr1Crky1RyRlLFZql/UYEKHWM9Z6UKhuIrTTgMvIi
jQQm2QA0QZWwEeicno6mQVNQGtKfaw3ADuOUSuoA+34TyO9dRzfaasSNzni0
AVA4xCZDRYaDd2V2djOpL+BRmkC1HyTee81w6rhyIhps6e72d17WOg7X6oVx
p93oVISbbBkzNtwz7+h3dlr8oASdiiZyDhqARkelW0Xky2nxia5wCzNNc2nJ
KFZxuFwP+KOgsjd4w8CtnHxijO79yKwRGlQS9rMbBhILANDF375RtoLw3Y7j
OwVlHxKLP1wJB+Zb9tAaDBWNKXo5ocwqZniWKSUHllfxNm8Jab8cP4TMONu6
YHvVc3ROR3zBcoWxUjOF9Iivwr901BeOfdqBG/pz9hhzRkCBhM4KeglDDE2Y
+zakGBHSh8BMIu1Jj/99qx7QaFMKBijGRzKolMLQcpm4WuRZqJLHrYzweNDw
HUOrcxJSLkbmaQAtDgp6X9gcfOCImzlTdCr5awiF+W6xwLqBeK0V1reDxJWy
rxZ+9DGMPiAE8M1a4VVr4Nz2j0UMHEHCJ1TABILa/pMA1cL3TMDXRiOIB/7o
RzLSMIc5fdSOa9ceZ8m0OD2LG5c4HXnQ4E5TtbWMzlMCdquESMMF/lN+M8Fm
ciq8grmFgd+aRI8pQMEukf0wgK0MAB5PqHqCoperJ0b8u48NRHifT9xlxU+e
F/WYR7EFqh8RUWmRIA7jP/+Nr56ZHNg+Emx60pnz0k5UHowhHGdneyQqxM+5
PZ+OgriHS+bfEtWRO3VOg1dQuLTeoNhfqJPVN/TrKb02KSrGAndBjCUcYB4M
CsLVtK3TiVcM6LIVyV8BOHciUZTRRBwbnflqzIOqcgwaUc4+PTpqm16BaLwf
XUTv+XxOJO7dM8Bgkcg3/tlhGlJyNBV4wIf4RJjt81GqPWdZ2xNBr0q02qex
jB3lsPW9XgRyyMbXSt6g5/PO9g+/yx46okhUjTlLmZEu00kO2Te62SiOwUao
nkEc3CXfnef1cKfDFhjmuV5Hq6FLgX6wfEQj356ug+A57AWM60tjpX4298By
BdRL2VPc4Q4Lq+Tds3QtW/YLZOv/M4sSJviPyVnJZkPAFPNWTtjcLiR8QelU
v/eaZf5q69qGis7s5rKJD9x7a7tghHOhDkt6GyNgkVNa8Axhyi35vvwz9YF8
ATuIOoFAk+czsmv3Zf1TBUYjujDzPHpQj2iJuSDOWdS7CQk+Nxo876H1XSJ0
ZY6fdYTGbVG6FrcsUWccwn3hejUrSh1An0o11E1R/T+lFkwEjo3ZZ9nQLkRr
x07y4aryhqWrQsu5+5LDZsGMY/2MZYZqFiofjBTPDgpzjXIaCnj4bNuTIq0l
70IWCDvc8q6UUa9gFW0Ux9XLgYUP3ADxIAossxhQ6diCqszcjXdkWhNfOf/f
OfQBzk9x2XVOOXbCiolQpPyL2g45gCMxMip1uRYp0pCu3fa83DNJgf/wbcE9
oCkZgU3hFiJugZfRkRg/pfV0xpLAA7dLRyQ2+tNWoZxht47eQMGu6SQu9P3N
sWnnv5y/nnfrcXuhnxOhSKcHTevwX68Rl2Fx4wDcSTc6jWPGB65BDwGPdLCo
xUYavwpLq2QJ9j5Qe5WstLkrtKKco+sKF4MmeHt9hjMDv2KmGvFfXoIkraX6
Rf5blzjH8ftzE5zNx2oKAtwHI3cATkpae2/2msWXf/4bNw3XT5o6qnrYXTz9
ryQJBKNekFGkWh1Qyl2D44VC/Gz9rQggvJPO74ys4sxNOywe8KMIZZfBoXdT
8vRknQO3a0lhDm+nQ5J9p/aYQe/Cz8G35yLN8Z4GfLPk3Xz7BiTCZGCUV1K0
Q0Jtu8QaK6GstfdGHANk5n4Rireq0ZPr2sA0O1Yz5K2cPfyV3raNyNrV9ZYH
mEmgyVrK+V2cGRCjBlA4n7iy630a9BdKdrXz51XOQbpSsnbwlTGBFx3/rYxH
8lB1Uwu80It+4z5RosR1gpMAumHWc3fCuBKErOaCzaU2hEYXtIPVLTpaV3Mt
WsHMqyso6f3+F29Q4mVkMKb4OLlPpUFn3YGQGBssqPff3vpUc4P4nbbD6QR8
Y83QnnMS75FUZMo2R0lagWqPC+FAm42u3O31wv6F0QOBmiWWUG5CiE8QSL4q
2GKb2FmoRzRAzZhp46MUTfZbiQgxTj5XA5mt8H4iBREADegQi1hhfR8YU1DD
U8Z80lWIFg91jArbydK2NUKW/3LHTBPgDdxEc9oINL+4M3TtyW5JjBT2ifpx
cdFOiferc9T8Kz7iaBLfTgf90mQKW1nKd8CjqhhJqorwUe4t2VYTJq2dUakB
EdGXaCnK8+bu7Wsh4+bqzOngN4DL1IhCs82yAvtXqVsV7nufw1F0Jl8oZ/KE
kzpiS6KaeRQTaDxw4LLcfVTPf+KhpfJus4fkyIY56QE6/Y8tbtbPeKOSODrL
NlLMf/YThTmVfEC6CxVVUP9J8zkCo3Y3zIaVvvmkqM/Xv9xD+mR81UKRRpYM
zTqwBM1ThnB83ST4Ds+3r52eOTgvpT6cURTaLVE2G40SfWIsSp7nfSU192Ud
w6/U8hO2TIDEITps1WKERSncwCpabyE1g60u7UDT61+Vgb/MkQR/J15UMjeM
c0zCcN5IXx4+8qBatAjxSxx9r17DEbHjEHM/m6M8l0YuBZMxCdr1wTaJmOG7
hncpenydTIPBjPmYtfZiTqx4YHQ8hiz/aetwVrz9MzRcdNMDXNW5NaFFxU31
t1flHZIn9Js67H3EzptpebMi1CGd8VxzdPZdfjIzFkJtbMqjbYFXE4Z0qzL7
+t1ZxSAPTgOQWzmtk7OvC6UyVgLlgOnk1bLNGYKG1pSK6P+iavk3j6suW1h1
gDSU8p5jYguN8wIj48JW39PRZqcbYybh72BwUH9Tw48m9/+wz2hbftWk6yNX
s0xG7MXUNlqTSSlarf3DPRd0p96Ca0BlVXrqegtYe8lhgOLybsszDLNN2yEp
PPBeiUsDzRVXXsafVJqU6VBBhNffnRvuiJhtXZR5xlTXuo5nskboOs+5HFxq
pBXEd73+1PJpd29xW7vr1Obr8IhM9bdy5m2BVvL/CK7SJJdxeqlIb4YAodiW
mg//kVmZOg7Aw96PDAp91YSI2ELS4oXTI3qZKNalTyot/ojLw7OmUt8ygqZu
PDZJTb4sNqo30/x+5ViE21qX75Xiwz9ov6p93lGPcgDif8YPAx9XPme5QCEI
HtW1bbOL+VpZgNZfYcb+Hj4HLcyX3s6JB8/kxR4HwcMu2FbIP/i0skki17wc
amugDVHjH2fOK7w/9My8gVt6qeuiqsUGm7/s+CcWrVlbvBoO9f4PgaHDnW8N
Hs0VDm3DQEK+EI0tOA/fexHANrY0wcCTGMXAoeL1WIajYoXuEclBfCwVYCDt
X1w2MAEtKL1PbA6rI4Mw3pnbe09gTJqlGquZwi9j/TNAUC9VIkRrvcAOAWGe
6b9zSqw6Eq4ofq8QakRs0mLjf+W7bhe41zpooN5lQxzOWzC+Av2AiAGh1Gfe
SMulXGShjf/XaN22ibgW3eZsPSbKpeL3g07qibqx5HFzlIOZ8LSONp/kZajH
uORW+jP3FHggnhXda3XjvRvuemMMQWHSmZ2B/oWh3oGonAueNJ3AIn/Hn4t1
cweTVZelTZmPiCa82OFmhDPrEs0t2ZXzrixYPpGW+0Id/mgqZpE6b4Bg4TaM
aBt6rkBKgyYVKECsNqrNB3FBi7GAc2sIIR7FPtOzMSjJC+/VW/AtVbFTaUF8
qgduw0feI/atz+LpUjcQ9SKMkPg0n4QsJPe/4j6jZZMOTbipzfqPoLDaFqv+
BjvD98sz+ay7zHcyeJpTaDNM5DS3C6mpnsM4B+d/+AawyXIKKFnEGZguH8tf
wm+7mNJeYYHrk6LA0ZfPkVEJC7rBDBbSjNfFf3c7RRVD8RXCWxL1oeKi6zkP
9N7Iyqiy5wTe4nq/xwB8A6cE5W/gUqFCGwfZ9UNlAoFQjzbTQ32kvqR0oLDB
1GI8f6jiKBs8jdL742R4lVVHa3w1xFhMhpIh7tckQssMkaaa1x/IeORRWXqL
HzbET51pRskUEE4M0V0sz438gMPpfZr602brsmUm0AfdpLjFZWTPYiPzFWjt
tCZBTcYKPrLM3UQITTAO09p7nbykhK0W5JTJWy/gsbLIWEFv8V7j26DS/+4E
5VJhzl96FYg+JZbJTBXpcdH/cs14cx67Wp5nKRi1FedOb9U1qeVKXoVvmtlL
gFFxDQZ0T7UxwBkmhZu9jYPfI4/9AjH7zdJU2tN7ah6G4I3zAZ6HPqT/AJaw
GBTZipd+vA/cYNvLa55kq7tMeAIaFp+Rk1CQ9Glgcouq8/hHE2rtCQv3WOYB
RcaITfbRIdpQ+1Vfl+aawWZZJMWURDj0Kbo8cHotn+dG/LdVcEQqn8XMqiWd
1bCcVLlSdxDLqhXzdCyRxR+lZ2Dv34LNGVO4a+tr/qiohB6ONV7mmpnuuI9q
yY7VIM2VpiDQULMMmKQrwYW0SpGmaQYzAV4+zjDAn9OxcZCSro+e7gesG4iB
UUeX7aanlK+ECCgOz7Mg5iqWnur1WF/heqzq+f2Kt4HkgGaINjeFu2MoBZGg
4ucp1Ck58yMW+pdMpcWIhzNIan4AXOYi7oIxNHKI6isD9WyfRNqtFncQZ6B4
ZNxGkiBZw1pd2QTEDK13SITkkCunK/Mc2tSU3v0zUhE7XmliVzDDfyZYKJfp
UkrpF/qH5ctjjLMtDb0m+6wgf01lRszM4nGbxu7zw5UFpbVjpAXvWenb8RtX
QnuqtaLNTV9yknv/OsubesZlGiors5fVVF9K8AC8/AHWKHWyhBSSr7dbdXwx
5afLxmAXfJg0qm5lOGiZZo03785gI7+iL/+UcrMxKXSqGO/WbPAyhzzhcR43
gA22cwWjsbTq88FuKUM7JySY283ZBxJeYYPHrZFBrXWT/QijBFEu44qG0sIq
I3QLyV48McwzG5s5GJgXkKu2ZZEr4Avovb3LR6rol6WXMmPWSp+s2hZPTeXJ
t+KMoWcdtwW5qUG2m368ue9Vgtcx92Igsk4/onn+uY6NJE9z9JxFZoIrdp2u
gd2N4TRMaDpikzwQrEmxUgIxvWFgZs2bdaD6kMgelm1Hucx9Zb8B61GNwJh1
HNLeOQlO938wsgfJB+4w57/wDaSZf/bHc1H0nOQUvPEedD0LqnMjv4sBtjyQ
+m7hIY+EVQSaHY33p6RnN4Dva/Skz+NLiOKh1BZzvzEZxW7iWfGZaotYrFmY
3Fh3KhCRevxjM38HrelYOxwAVj/zaWVWI6buKHGiuLHLojxmGNy1CLwAgb4t
MlNTm56tirOAuOE3k4ccDG+NRxp07yfz1CR6FZ1k8QzQVZVcGFDshGOLHYiq
fik27zz0E35sM2Tf3H51m8/ZJFCeDaLBYxK4UbdlkPtasUl8WBE13mDj8zg8
g1KEetoiIu7FEcow2IoamMP9aoog1easMwN7mJ6aT4EFMMl0jM/r0Toyuer3
6YKd+JhOjf32LkVTE/g2Z0Q82AP3n2nmqFMCGhQmfqJphz0uRK2xvmMGJGzW
BcM4M9PcSWPogsXSu7vTSi11rTaouU+yuRYImv/Ta+h7IbTNE8/gUxde/KB2
im+HQ8652l4qVDJnnFweRfiOL5qgKcRimcOaLrdlTe+7+aPVnl71kadyK5ce
673H4Wdh9HnYAEkP3KF4twxSdfSJZOdMqUKvG7gof02tLCHdhixJM6khhc5Q
JuALUVDEHBVdmO38U5vetyqgMDNU7+1ByfYCdhSDRM6hP7URt2bXEdbiNp+q
s7UR97zdKyoDiAdK51uUJbT1J/UJZ3Vta9HDkJ/TtdjkYoMdpSxtzBLRgCcn
psjI5cCVEOxp0IWyQo2OjIvhU8CCQ9gF6GayThFX8P9yclyN+jq8fgpTxIYy
iFiAuW7tJbdMJTNyg+EKzIH4HXg9VFarjMUR3iB0WcffDoMdd6/fyxnvgZ86
AtNl+SmEZc29vIQNG3BnPdW42tq72BvyML1NnbOLcb9vZScod/F3NGMC4CSs
+Gw5Wiv7N8Wn5XrSrPcNRcbqwmCT6pA+A4FLD2nnB51p/1GQwPui55Nhx2Ob
EYcivAwtoY42c+4z7fabb02F6rta2+VvMvWhQ0cTgvpkrfDV8hhOFitCj2Ig
7xc2oNbre3Ea58KI9ooOlr88TzLVLbjtAKAkNWVzq/j4+xo2357d7QCYxp2L
Q73D1HF288GDD/DaR6hlv7aC8Cp/FJcN4ptNxTUhLC93TBLEYTL64XtCKREY
9DEaLCy5s027p92DeHMwnqfGN1+aiHGX6lR8NHmOWaXNsH+nquLcvuwUezmB
ewEZWYylxEVl+yAjDaToufRgMf3CScwCJ32o/fo3VG/Okb3BaTuGnvM+xkvp
FipmU2pAZO4BSbsCm9uQWx48a8pHQJHE2YwSmTJribi+Q1J2fiu+7pJ/E2JS
cDV2TWMFweNs4j74NI+0XIKJLEaFReEEmmjj8Dx7ACZysiuFV3OQ06uv/Kwb
YRYVMT6hJemUxVey+edT3UliAvOBEbSuoSx6hEHka5zpb4Vpwg0Pcc9x+NQ3
uiA4OlesmvCRcO747ZsJsWVIw++/POfbOEk63qDd4pBa+9/NlGMij37s7ph1
c5s+c+idTyKVRuS1COkLsTJTyQRywU00LLqNYXl9pI4XQ1TfQXglwjU1L5cw
qr2O6EKawPhq9HLwf9d4R34vORSuaQdFvQ3fYEDqGeNXrasHn+MlIBlYngvW
fBJeoxYrCpedBIJ/Vooan1CMyK/gz6n8B0MF/9D9SlNPW3ur+MWDur0eT797
/dlp5YaHp/0LGGx4Y3J/Dgde8B+JVNfMFZuBt8eqPB1TACysjhpdgU5ws7uB
0gQrggvS5T55c5/rv1JJ2/ESUVdSkHvPf6Hx1DMUjr3YIaK7TL2EHjAB+QfM
lfcDNlcFDHcd+AZWYsSqcWVzKC2fMSYbeihDDRJcxfh68HTR/x3zq2MFsDPf
d4bRZTT2G9nNlg94BqWa5Vh2Lvr1NZ4fz77HZOAtoxbnZcfyiezkTu3JzrSS
OUQLdyv2jkZobQ0kGPk73ualgki7DPRbgGeZMe9Yame9T/IerDAn5RPf3QPM
KxO570sk3zwB5Yq9wLslN3HDMQ3Q5ZbaWP0I2UMjC8l26LOPBm8dQpfPCrmJ
dB1eHHupluL6N5j0SZweJgluVBEeL84Vq6pNNzxtBmnQn3FZeneRa4NcyECD
mHUn2tKfug/kj64zch4q63vdQ/ShXb42C6vIlMXqYfpg+eoZnz4/jgsyx0Yy
UVwHcrkYYsGpbCZv+mWRdCwbMq9OT26vGd6lWsRxNmWXY0JajSBvX6FDKRhV
4LfVbw7deNeNVLojP1rf9p+w767w5durw52j0l3/FXGpWb6eQltdQVCtXcPE
egh694ebhQ9DafCKdKGg9/Yjj2+bcfuffdTDN+Tu/iCUAqxjPzxqbjp5RERj
iRiqBZmtHvPRRBDlz/gcjxo2BjLY0XG+TplsbEq+NlYCfY/kQkiJGALY+WTz
mosvWUbAXb9JPXbGeLVsWI6rxFBdRVHP316KeLFApGogKH05fSbeBwJyRizC
Nv9rpOcqIgiZGexLx/8DzuV5RSt22hxiyEwWF4EEh8SYmgIuvrDHAs4E2J1G
p3x3Ho4m/U3Luys6aalaEiXlQrRnOOccHmj6VEMZS6fElO2ct96s+5VqLPoI
vVb3f0nB74CLf6cu3h4wMxiEnDjpdPonvM5SuJZ5Q/FHIt5icschdypclAfr
LLeRGPuI6UlIuLMOFJAtVpAWhN4EwotkxAEW2SRT+YV68uJKWRTNrtIW+uFL
jmSQEDx+n2ZSgUvg8B+UY95HCjbQpgatx84aDdofhJBjjoT1bvTGJOKGIbqa
340m7XmGgZQkpjXuRE4cfIerybFo6L7icBfcbYyrRxBdQfto1pv5TZ/2E9rX
41px2hdJEXE+tmffds9OrGNp02yenlY0BT0R29MFSgUtIMC8N9QJUo6zXgiK
VqM4cg3Ev3+xZq18sshNkOCbY0rDTapv0K2GzBoH278OdsYMrFEaecvJX1XQ
yVtThw8dQ0DlL26gyJ6iUVvXs29Xi0Gyw/LKWguHX5Rp+Wc7oQS7LxKRazHX
1MsnZ5+l4LaxZrhoRDhDu+K9ShTfyERLH706Qt06G/qliwW48u+2r+02bJTl
GgkYbtEXh9+V+rfWD4k3CjAgjShbPpd6BUOXbbm+elI3npC1RebetDk06vH3
AbYgNk5BjMfbQor3NrFN6qIdOIET2GXNUUFmn5WBF55aSxz7pR/rr0TqJQf3
AC6lWee8Mluz8+TMonaLHh90Npqzse++eBHey3jxrDwBfa8ODYjQR7nK0pro
CNf/nHRPaEqseCaIaTgqmdo6TTNOM0g3oNt75DTtsbz3eSKHaVsWqHjOwtF8
AYTeNjt+0CwO+1wtrt8PFjEUd6Xjvv+4QV4PHEa/G4ydQY/P8VB+X/2d9o9F
XlZydntyee7DthOj27cGG9Srr6FyTA4to4QXUIhAzs293myWtOjVFK/uaVYY
C4fP1qTJTW5ISId5ZY+hmQrfOLhDWuLaKXol/hBQtYGLiIaN/zOBM028KXfl
4KCuVWHOoFM9RKdbkNFNsHiQu+kcgKNTFtM6SLGoVYhV2aGFJt1ERuIcZjJE
c2iqQiSF+v3HcuAw++LiZmadLi0UB5BbgNQNBtj8UV3l4aIjtRR6DpbPbIir
J/V0RhDC+LYQoggb4YafLP3Pw1NDMkToyuAAVRB7QLKbwtvtrBR18UkyS3ZQ
C2swgpUGPP7NJOrNFSt/+/mv40nsQcx0YslTpnjrSELfRxz0YTvdgbMfJFIE
o79/0aB2mCs9Iwx8qPF7SX5/gFAU/YJmtoVRl3yrQmF9+j4Y28zGH3tph6ZD
TeN6FzCrWQoZ+7aOq0QUplsAnggSkZbsls3nCC3KSCOY5PaGUq+IabB9Abkb
woRZXXdVIkhL1+5KoDZ0rQzvxQdto9ZEVLS75+VaYYSHdKTqV3Y8fpuQN6xJ
qPUDnpGRR0Ys096IAPa3JcbJ9Wt0HVLWV41uPSMDVOGzVAioROT9dR3sRF2F
ertjIFKsfGNXKkdkJSysM8tJb3Nus/s5XrWOKW5ntzaE09z/xxgjByk/TrO2
f0yvt0eL6Ha1Sh+0p7+kZziF4qErLp7TjFhVd68WRyIwQluUpuIrnUoLk0ac
GPxBTF/opxsSbp7HOdFNvDsQv+DuOHKug0OY1nBLPtYg2jqwwhHB/+iEXrG5
febeUjxjp1E9lfnxxN9wt9cznsICGG+Wvkpv89V8Vplc7cGwYqtISwR9ln30
/6tZndFnANWv7UC77FoaWEEjWmfkiuoO1sSSCSExNEZEzExw/OWARtJ/JEDa
UpOb7UI2dHM3fyQr2AmM4KhB9mZ3U99gytUqpWA9ZVF3vVQzXTCshhet0+uK
TEnokqNrnEtR4U709iqivfbKiCXb4MxXOx12Ii7fNAcWerM3J9bt2DcAhTz6
QqZca3I79SDQzSmKxxKFvpkxYz1biEJCB1qvwp3u6Dftzq4BjQgvpaD8zBW9
mmKA+xWPNypptoBmnWRSaVH9LWJXMTAzlGEelhKRUvI4YLo4/uzeddD4woEk
93wcvN67Uf71N+XgDE/ZVj3sOLx1Z75fxu5Gf4ngL0gqIBZNksxd6P4gmE1W
RLFX1BYy2hBJYquWWNMLNdhFIlw6iKjn1/ywkjgzj5sz9f8M4fLuxRukcezA
QFBAH+eMlWOE73BlbgGXZ7unw/6h5AVCZ/39p6h/oeuDRgRSXAbUYSSV+egf
yKecwQWPyLx7+h3v5KEqeTCip6gv/W9yCmafQa0XPz5kyBDhDqzGCK86Rrce
dll7cThWlgWedlGXCDfieLZ1lCgViNVnU9RA6iyp0Q70/nu0aQCFoGOAzs+z
kgzdhmj7aV8eUBcv2wtLknEXnAJo53AB7rfzIGe7/p64IcOuDhaWm69PlaHK
6O+7g1QFFs0D/zcpxt2wJWgwOrH8uiPOQkkKzPo4UYrJ+M1hfAj96CvnOAcC
7UWf8k6Lb5dX+R76KrFS0tWzRc69KioL3SJdoZsE9pY3Jz+RBGwhL/tYsLsM
7mzkt9vlDvr6gTkx9Aj2lsdEjVzA8UW5w/0u+XmtQ8YHTs4om7wCdBLYk54D
+ayBqkfJVln67wSFPCfycipg/bnDQmx7W5ycoPo9tCHn1j2QKnTAeo8ADTrD
K+a4ekzm7VwoXeypdWveRVvdZe6CJWx2K9hbfpmOUwo68DbhBRY6S8YffoGL
QaY0MO7mRW2haAQd4FkAP3GZ7+sjbcGM+RuPUv+oC8rHW96zFcAp+KI3mE6T
ieHyk9095JXTa7UMdrld8G+XngFLUaVb4CVU6j+bxgqVKiQhKEmR0wKW7jiG
chGdkgVSVNvUVNtmtr9akPbEGgI6wIi8+8vHknP6yE4ma20JqOmiibhvG7NS
wtwQ/mr4VlmsNs8YZxjsmMxdhnIjRhgzgA+GgmLw7m1pv+iCgF7CabmBF65k
eA/ezWHqmbn3agPDEVlNXti37X5eomadtbMfFneTovJMfp2Q697X7zqvCgyv
72MIOKAeaaApAOB/uTPZlAqKI24JMbc7i4h3tTUSZlVZthoZpTN46j8IghLc
s6bs5T+gVGtzLPptQ9zfj133lGisJpdqHaFy+MXP9KbBbauvKTOji2e6v6of
DfOXJxhTsN20netJzLoHQE172TyaE689sZJcMU0wQ5PCJf/iprocAIIRa0yI
ArQpq2VyA4VSirHZ3Ufl3SM2suwrF4e8BQd4Y9Fi1SmnzhmLzZ9v5C52zWnX
Ykud88GnTNOrzSpAhA3T/yqlBKvOoN1F+yXlUtMr1Pehw1N81yKu5+nOkxHZ
Cag5FYL8ymsmKaHMZyiG60no0Szqhs2ZcnHRm9YeWlCUTjXLcxpecjgQC/PX
u2X029Hh2G3zeB5oPFFs0/7y8u/upNn2qOwgdjIHGwrpHuEAzDbPgPayA6RB
+yEQH7b5LGNQn6k8DNtcXzY24amYeVJ35oTZ5/lPbnP5zKzwuSrnR//C2ceM
AohQHB095ZmgHprE/iClr6SAGzaxtWOLu31Q+UwuaMv+NzTISAgSuVYkUQu3
bqJI1sqVWmLN+Bv96rETXtDQPZFgEWuJwZN2EgEIJc/21FyUlA+5DWf4yr+N
4TddVkwYRMDNMNV26PvsPLTOZg+oATH9otDxgUR3LX3X/cmfZIxqoAzchq7h
I79Qj6XfFCqTqz/G9oMMFPC/QCd4RcVe6gkD3U1RPnvuu6xIqlQ/g9AzWk0F
22EJyX8crJN623zS6BFRkcezeUKChw4vgCCMF2V3zDVUWBRvrrceVaKI99aR
q3IcpdGH1nWfZlN8V1cyQnEhrP6dWtHHAUDVfX9KAhQdxNz3To3TzGBYveBM
DblkYzjWuBhG3RfhIsKRNItFbqVzfJm0ALyzXmvkLOIllH43xqsLOcgbgJZq
55EJROS2uS7ZdtALSn8brGv/hG09X8x06nyvktQTqsEXaZG56hxfHfrrpU/c
UhN7s63vtpxqGI8PIKK24rmGPW2I9KY3BqzKzk1toclMENxEQr0fdtx2R75o
AnU5TmawhsMA7mdmt8xelczqXwKMcgRU8n0rvxRp/vUdB9j46PP9Mu8AA9Xf
D1wsNfLE1y+vjoYXbiAC+HaFOiN1gnOp3sZdldczQrxUIXC61l0sP0W31Lfr
nqvmbtjZ526L8gywA4bLblS2vdYGB+sGu2Lbav/4rpRUo+7rZH61wU1eueI3
ENOeyu+4mFiBPZZK08djzCHppoWDsAJYAo03rXWpcjg/+7hgzdSAlwI3Prk8
33LpJv4gy0AINMNtP+u5kIzh8ZwTPplBFn+HOHY3HM4EWrhJC4qq8/qy1l/r
DNUcYMQJk4DSXP1FzVQtjN7fXAbLrPGyyHfDB2moqLH9VJReN7B1sWUmLwfY
0RPJ9ydX1EcJ4zWWqY83tMwfPCwV8xxnqwvWS4jxOQ+uxMGxh8LMF8EI1VbR
Qe16OFAhEPoyYSP8knq+x4U7BXpEwLSzPstqxM3dHeyplRWZSicClO6X4ci8
NTYzLsLVWUxT6jBT7NdDhmt5SfUk8UNBOHgRUg57nF/k4RjPbEMA1QqcniIK
wTqKqpjmG7s0fq6ENDHMdTIfzOY4qCnTYuNyaQudYQZakeNnsLhdXv8Y6kAJ
oVgQXr85WV46jYoPJHydWwFpTBpYjbv7JF7ATz3/E2qPwXnC17Bh2SXUByiq
5+ip8/ZQ4zznRxEZu39AJCod7zW+s5vKJ3nN0BASuu4M6lCLS4HgrVg15PY/
plj3ubEFH6nMMa18cktpWm1qP6TnavJyqm2FSd8/MuZOaEYvbpMWHWxVuHJg
WAcK3cZFit+O4ktOkdLUi4Rufo23mDSwXFBNIxTb0ZWToYrPJjp8Y2oKU7zd
tX5j+DQE02e/v/EBUnlzw3Vx4Iit/hfbQajhfIevufaisAP2IEw3JrfrcyHd
SZW2KhPOESWupKbd2yVGGqjJEbIrnEaIcvXCdlgIYaOzbRZuYBuscj/56cUq
IKQ9bGmQ/3EdSF5Q8FpIsMZ8JVz0ZZk//3bkFajcawlQ27hKdka7pxDgNCe9
FY1JKYQM7W/+dLGCtcbk2iei3lIT/PvyuZaAo3sVHP6mZ5D2/aTere7KZ8KY
yDT5EPc/czScQsQILB0IlvzqbgX191Ccswwg6Y0IHgM4dXT6IRYIxdGoi4vi
oHFuJ5q2n0zSol5Bfakh/j6khrztCwIuVpBqLYPQX1Y9NyMBWvJFEQoMDenq
m0/GMUYMTEHi6BZHezC73ZnFEcjVtIhgGuWp2Hsq0taKMh4Cue0ozPG/yBuc
tHrv8CMeyXG2VXY5UtOghu5crOXlgBWk/eOSPxa2WgUZEy98SN854/c6Qspt
bKVqYUkZjojWVFZyDDFGkzT4jHYGmuzk3OP3EsT0ZQPrCXeHemvAT/NwYmVs
jcmWkSalaTHqSPatUHl0YnnSfOYM4aOlHI1sRIaCZv0BvKrS0xZZsajw48Gu
IP1qM4vRHANGouFINgYXhowmkMnFDxTrYw/Mwz++Ds6dpcYGjpJ6SyZcp5LN
GdjNdLt6yoXnMxMbRQLwvryHvPqXre469/uryYh6wbhUS95FoB6Zgw8RlolM
Ql+D/SHB/GAac/NeT0SH4b4rdQND3TH7TV5kx91Lc8UTLZAEaviO14lURB4t
BrN+4EEpqvDpWECSd7btZvfnstPDMTxGJZv3PB860MbxqwULW8OW3f75T05z
DguZQI4llijiq3QRlnlmcSyEF6Vri9jrJsl0mDAH6+9AdUPQ2ohgeaTgisoy
rtROGXjwdZ7354fH7zncwyL3j5hLyRbnSu+Cu01DfmCo5kxHesKPZM+wlnfq
pzNjFifVpfHciZqQsVVc7MHbd+yh9kxJkYCBXnsP7axOeaeZnMyavimD1f2t
0wL0LYLYopDoD5gz0J+DZ4gQDYRnEFpiBFhd02+bhHJbho32pqRniX2rcNe6
lQOulO6fS1fd9TZey/MQ60UUj0isThZBYQxYM/+bsmRpN3giiV4EKoqVpZ+R
HjuazW3bjiZed1rXHCB5PwJJLb34WDkEF5oCSXSk40KRpV2p7HjMIOcP0PMq
v1YTidef0A8t4Q7ydbHe9nrZleguBgfdsxaOvHufjDw3RCx+mvGqGOXrtKlx
PyXTbqUokT8/FITNfeZeiRdWx/fMFxV35LzlT9XH6jZcLuB4I4Ay3T5Zga0B
/R/PwbNx22E0DvK/pjcBgJlG0J0oWHRhBZYhLywFxm7fzeSK0P0hPoqwKhHN
NmzEQhUuqPxc1am8BV6PNOWgvMqhDlxVFn2H97/HlXmMzcGav4i8k/qdEX3Z
maWWyHlAPuR5vNW4tPMk/6ft25FeCDm9UN9pYDLCGro5IimKyW3GtbC2d0t8
6AsLcJ6Xm3G1HSsx6CSQaAzmMeyLxHUXVATKiM5nS81PJiNVGr1n4kOoNkM2
7/USRb2gZMFwBBkUS2ZPyszx5GMED/1/Flvotxe0wAX9Ot9SseXdAZ0R0oDx
WF8R90mjrsY7dkCjxIL6XpcBFG/H/Eh0LZj+K2677SZMwA2LGlXjt6GaFhc+
zQn7TTAer+oDVs4WNvOsUdJHlihGKnueNZJn4jqSbwzeLIXEaHRywEpAJ8Ck
Q7OSoWiPJDxeh3YhT9ONDn7lsrOl4efxJ9c3N8wgLihMNBFPKs8/BgiNO1Rs
D7HaVLPsfVeEP8sWmE+PCa+Udoq2zABRoaTjV0/QeLJJjMlpg6Px1brM9dqM
Alo1Xb0MXhVpaslW9+NcwNwROlVtjpxxxOrtSiBLqL05XIPMNYhwCXvsUSxJ
RREsDsHYIe2Sqw1ujTowhHNVSZzsXuYu3ff2oIgiciVxrzmLDyWKd/1iBZfk
/FWzXtVl/rxPveqXZ0Ceg/KFzSEVb1M/F5lR4MwLJwwP/o/KfUPZP7gYucHf
9CK/+MI/47FyNkKK7UY1Khtn4QCvdSwjg7sYoZr8Wjx/j2Zn2G11m2MGLLid
5aU1Z3V1hZD8K2p7Ir5iTSlD2bzcdT+rDL+V41VKVzXIBdXViApMFJrq32n5
dfbv9y9eE2gOay33JHfLHJLyM/aIri90b1d1OaOyFtuOp3ZI9/8Q+58CvAb/
ZrQ59gudHPHeekUs/7R/AQTa648qe2i+aIGX7yMMzbetEn/D9h1CWLCJ8Vxv
fdAUF5uoGN+UAK2fkyYAmvCV2m097s7zTG64SAS/yEgphejLhM+KAmhZ91wl
mZ/qfkUAHVuFSfbGUpinKd8Lq3y80MKUC5wrZFwkFddmkM8YoNsFSsV3DdgB
YTZP6w+TePxj1rv0DpxkNJ2cQDxjfoUJQVYB+aGPqrXD9lvzxKVzArUNks8r
ydQSzVkMMePc9PwNqyf8/wAzJO9gf/JNdPz5Fj+XJnqDF6VsUbBkWHVCFCyh
qUb5Iir6Iy2J8QjROhcSkFfWPyZ4DBpkXyXVwPj93Y2spM+ChClrxxqn5/jU
mRLjXdxlbO2j1LTDdfl7EPshcEx+gIP748Q6FGs+GF6a0NyKFM+SgDxvuCVN
kO+YxDM2PBDDVY00i+qWbjjKhKv38PQUEmMZun7EzL0Kj4db7Y7ywOJ7vAV4
RY02noCuCJ1yJ6bkWG/im1Bb2aeWLcO5cVz/tC3f8B90On/cfeYmnxmODF3c
ZPQ3ukqqdt+gvrX7L9ofL3XwVProC11wTz70UiB/TnkG5ud0TH2QUohx3+Yh
c5FvfvVqQTfnhECKMWhr9i5iqSftZabdOZ5u0pXpom0aaWArhZjKjtY1gI9R
pvlzKua+AHfqnu1RgaK/SYj4IUGgPuMkZvNc9wHrVtWjUC4/pZFLs/jZDdul
VN3PsVWmn9dK9tWA1PRnOVnneX1rQgrg5iiaibezHEOGYmtvcMlCcswcHE5q
ZE5ovOZ1Yqt385bLYITyJjuthuuUoezaM3moFJSJjWpVOVzC60tbozQfMuci
YCnyRCNaFkBgnR6o7YjAQ6GI9Wah6S0PgkTgA9O0rPjv9Eb8hPzLZnYz9UX0
V85WlYWkwnDlCBJu9KIF2u2uepTu3SMRbjstPj57mlTPNn1NZXPS3BsONwCx
1UYUpQQpo3zOLJ2SxibMdne+j7iwBOp/mjp3PTJ4Rms4rLH9auScNci3P/rT
XRFBMcpZ17SVEAOlRNchWDrTHvv8hvEryH4b5JEQPOPQUzmfZfR9WyjEgkfp
3nMMbWNwUPmPuE8u/YS2+1ptOwvGCKsUCTCcjoj9pk6e9g7ENYEn07iM+V+C
9wTXU4Sb/qeZ9wm4XUOOeaLJ1LzRW/Ad7c4FsUtFLdziJOy+NmDI421f9PGi
j4j7n6IG7HKHtP73AdASFCfsykWAicaBkIzEjsZVdMQxICaXqBaUgCEB1y4E
GHm9X0xDHH08vJeZ5N2GnbSMFmjjKKZ1iwD5byfyq4C+CQWjwPmISSWSPLLg
npM0DL60Uuy/7Y73Vm+c4qejd0fbIn9ktFfu0GKW6gZfZbH9RjTkQGKsab+R
lZpaDhbU3Xbsg5GXQXXEotHROFXXelteGqp4ok/+l3QOkcWR6ggx+QjEnlJx
kqu94uVD/fKKf/HjKn6tS8/q8Tfzjt3VnCdIv8ShkHwxB7XPDBe+QqUQjdPV
hySDfYolIII+M3Ayh3AAHgNvS0oM5eb18by/41gzt7NA7AxtIWx5wwAlMOQB
7dG+yT1bAuUXURTd83hrQgu1QxGizClG5NnBKbKxuWUMvSaZeAzQK7kSLtd8
puXgdVb4eXrLxfs6Z3pIFKGb0ngLTETHnCo1ylGk9jQZhwpDBumHIpFOtf4s
6PJyrh4tMEj71on2J2OyVNZPiLhJ0PL03aPV+5oyxDdVF/jh6uv4qBTkr/yJ
Bk8KN1LDcjJ0ylNhaiyZTu0jhHD7vk83zrY2J5xV+k4ET29GFzYPHQZaNyBr
QOrFTxsuTz4UBMes3vc9XfqHj+qOs8XSTKWGQBfWeLpZSyGP7c2HDQZj+Fxn
q4jE9bLiD1lxvIvyj+tJJcuEheKwQ9vUTNyjvhpM6FDE02v4GhC0gEXAHS2E
IRhV1YDqF7GR0RhPsSKw6w7b5d2t3YRF3LPt3iSw0zPL8UVnJZMOrHuEisGk
zRysrBr5KMfa5yB0T7m5NBZ9eofr8Cl1ZB6A554puswscAMCEfln8bpyQe3I
VaZmmf9vTKsa29I89DRNUbELZ4tahfX3KInVvmzX8C0luA5/gGUIEWOnt1CR
nrKBgq2HOsyG10x2XdtghZXPZYABX++tN7NgLZ1FL/jOueo0TBfKOMlax2ru
wtRyam4nhwo7ucB9rU1pNc9MG4Q/I8JB798BW8yMFJApLACFLEOJROcQ/9rc
2Lo7cjsFffl+OWlOsf7JqLSbB7pQQzt9aLpBfyxil2dvKsnGhO038gWCnghm
n2NwOAxSgrsnPcri7F52+wHsQApWzRC6BycycEJhD68HhpYG4cweyzjjk/EY
MlJ8zkRl8Hp0T9Ts00+DuVWX0hgBCfi8FXcR/2e4/Gk/6o2aoLgAOdhCAvnA
RiTaxSBFpXQ7auO/1026fm09XpB3LqTAN0rsLIRm/63mBwmEgS8YGyzKz0Da
oOmueGGUMH/yha+5MW0SHUWEqO+KvTyOsLkZVJQVvjyLjNctPFH6KydPsjZp
1H3h1yA4JW9PLB4aaMJfJp49nrHE6GsyXBkBGusTRDuzRTQygCW14TCszD3b
FWwu6ZQd4AsKas0lJWvzXFT3j8QRAX95t3ptOYVqqigY/nXfBuRSRcxSFsG4
VqBMJ+vrOiFyPrWEWENmoL/fRI95aFtcC0ZxJmXAWuqgpzrX0MXKU8fmRe4m
5yvQA0LbgGBRTuu9k2BSeUvqYiWWTlSWgeboRNiVhXCgY5sBNkVovoweY2Bw
uAEXYD+GUnFR7HJ00Wv4BPLeeackXAojMChAKKJQvMIZvTSW/krGEUPZEb/I
pEXdD1WMbwbuh83n72k4u/m/oUbnZC6uiTXMNQg45UvDXol4H5P0Xu2KltF7
WUZdBR/18Ac2hMtCC3pjy7utp4nJSvLsHEwuE4kR7fN0Y9DH8eFCmcmSuHQf
CnojC5raqw83utJP5Vc8k4s9zc1kRP0uMhclh+eFlCbBSe2vLkvy+vgAT/+f
IvKhYTG9rr3Af6eq7QKRZqoqy4lzztzyzqxQjm7zVYeplM9t/wWwm3e8BoEv
Hp7Tv0b4clVdAFqK5YU5b5ida07I3qrEwBkwVxDFqbhg6YV/YsHObSkHzebl
6Za4jBItYz3K7nn5Ne/UcZR6nzds25JnbQPogWoFfosDUJJ9uR55/DdH94hf
t177kNqIscV7CTadZZi37R0Os/tzBqawEu+hyuFSN9MUTGLGuooLprV5h93U
Q/LmGC6Jhr21g0cmUVKuIEiB+81hCVXHEu9dPYdbcn2LjErgdgMvfxg0k+EY
muHjO46F8BQ0j43QIDBdUis7SGnv51tPrUDyBgWJeXEIeFSn8Ira6SLXI9sY
gB0e9UenvCV/j6AOvT4kixKXDN4pZUF4A/zIiFwoEuul/6w3OaSfeWGdOEpT
T8A9uSrYcJaMs1IQuEzH4GmZuUcGl+PnMgSVnvH1PqRr3Wwd5X19QfLFp7ZB
x5GjwcCwU4HVw7mEma++R1IQ2q/UPA7FaF3iWC2fd3aVaD689Q+HYqPq17jM
Kq+1w7t/cLUJlQ80CJESHstttRNCDtShOwt1eS58PgAY6/jEeupSgfkrnMr0
9ChFpAGg0koo1eRuhxjUqPa150d1zF+3MTdso0usneJVFHIfkm8NmxQ8aENO
AxjSLeVlvBRE+OxrSwrvM+TfnfJhC/Ip4qiTMNNGFT8IwIr2B6cmkW9cnkVh
sbynak/p24jDOsMeZZ3tgjkZMj5JG9//JSri6NH7jLv3tOKmSNgDM2BCY3qt
FiiK/43gjeHdVXUYDLQMN9bDrrYaMQfJANN8Kfllt5xzfaOcOKyI0XrPAlyH
klNJWmwmgGngnxUrbJ5aVP6N8swwRhKUWKn6QOLITDejBZG0nooZ9a0DJdyp
/BbEflIYuFHiVwlJ3fBmP7o9uuHZXufxYq1W27PdM62FXkQHXKyXLbApVeND
PzSmOCBpKQm9eiIHtN3C6xT/iAOD0SZX+9gIUzxjRTn039YD7D4l1u3rh6Ud
KfTK1oNwWSNL1v7ezi1ska+6YDdK2IN9o7jY9QEyVgy8b2j0kyC4tDfWAEtA
Cdx8aCKd5yGa97HM7AMehzheKUipImFyEQZGDlv12cPdGEadCD/cBbnyWMN3
j2RzvGiPZsva4zNrn+dt9Xde6zkSjOspbnkPZO5xTDmcKyj+0sIgHxP232EM
G2J91yKH7t6MCRh1qnLaISngkc2oeSHvcRy2opfp+2bQvpoCMNVbA4u7FKEb
ScNsFB9qD4vTIyaOFL2hghmX4F4YaBRab0E+ZnDtbFCOVwaV4lhnCUKUJYwG
qSEBrYyuy7oF4AcKLbXg8/d2Bke8Ta+FQ0A9PGTGMohCI9G00Gq9Cy9XI06G
qIGYsjDp9ZiPA32XN2HRtDfjI2/tsJdg6VvdIxxkezWHcxWRzIwmwL/NGV+a
c7iRUTTj2z8SMc+//WeCH24o8jpHyNFZiH1iuMcbretdRC3AxAn1rHKQeDkI
yYp3rt8NzksCbE67CKBJ6Y5mVchdTuEW6o6nNKYAVshk4fEsihZA1StBE+la
XJGb7VjvAfPbQdHfj1q6JRAzBSSbVGBS+8iAEeVlKSEZkldiAyZkahNTRCRi
sjMyoR4wC0HnIfW/rMp7qAZ99r/Xz2TZQO/BuHE5Zgw0B25l+T/oLS9SsoWJ
r/lw73XKiBx0KtSimguIUzI16LTViIP3v7Uwpnmws9LKCe8EddVMx2hKJ+d3
0BxQzxy46PS16OZgCt0/u3wL4tmmx6Rz3axIJqy9kAydoZAtp03QAXsAzuu9
2iavh/uPE4pXOmGSyv2ZBemqx4L0vY4jj3CB6feeW57NF97JXijoDrbhtO7a
LGzjmwfsWX552kYN7/cHtMfcNW3KB1E0/FiygE2BQr6fk8y6vCLv0MhYs/63
/IKtqa4i9172B4NeaeSVp/ZHK1mb3YeywHXDYWHF6ZTW9CjzLjpRJuzpRK9h
DSUyr2O+q6UGxTMNi5200TMnCMAAbD39VCjsXxSEiXc6hJfMRcCnjzQm7lPE
+wbghRFanj79F4nqqxaBEqYu7Zs5NE3m4xzKmez6gwtLqewsyS/pvCC9f2Y8
dnMKvXYa2nzzwfkupQm6FVveN6xAJSnvNZ6uSdu2DGrYidhp/gyzEEm0mj68
Ha9jHzJ9kJN7n2nFntEfP5+L4cBDCuBUxkvic2z9fYsz6mtoJ4P6hXMVHBzL
F2+Al18gut38yqpgqgamD80SYn6iDa+FwSiUVfbP4AK67rtoCkN3DmX40UGM
em9/y0vP2ubDeQY5x/EQL6LnQKweqNXn0+2c0Xpy+DF37oQau+0GtXjq8NHQ
IdcJyTv0aSAHVDjmYCyHtjMPuQl0p2j5XN87Uc84ac70dfZhh0OLiVb9trMI
f6KqiCWOF+nvZQYyC5HSkcx9dos+G0VlBH3BXuWDBPJLxtGVp6t+9pUXKniZ
X7negvpZ/Y9/lGqtAqN9xreWpl1p3dhcP0MQsPh+OUkJHwv4amrU/jVfB38E
SR6S04xXACiw/305j7gwqjKO8LIKVwIJwiw/IZz19CChgqT6zLk7TFUuHJC5
AKPHNqFgT0RKCl2Mn3SdYxVu3GVzRiOKMDVPM3dLftnjU55Y3IEJgBhaeCbj
1jJ5rPb889+Ui/2q4r8g3mqU0/LprXNR39b+N68F6mtRJlmGW9U48nUAU5C2
qdJAwsLPrOVzYB+rUuZnSdJ/uwb8kkiiqeQkZs71kCkCQN1IUn95GkvV2g5f
Xc8GTsEMb89U4vD+QVEB+3pAgfeMod7d/3ckriUg7A7tkWaIL5Jkau/BlEbj
dTc4eMM83LC+GzSD9YDdaO8DSqR+V0yY42GGLrwqQjyLLwNWEmbIgtHBvjl2
v0tUpJ9x/n8yQB0gnyqwMyJXLL8FOtwWjjz3PYorMNMr51U13Na0oNpommF3
KMitOr+QFWkmd+d2yay1btwPDHQWCMEhK/d800PH+26RFTWlJdLU0lBQXpQM
R8h7rXTlVW+uYsCOJhi+X3mnIIDi06gN33fPj12AZebDcU+2p9lR2Mx1yFqn
yn1HZMG691mzKORvl/eMl+uwryQ/PfYG2Mgnlj0+NQj7y8KCLq18LyshgYJJ
d5oiYXTXvKaToyCspGX3yAR2nVoErgP1T+SJgoNSEOk38q/CpxbB1+YfdbqT
V+yNNRtmQnNCpMHPmaIleZ6c4gKe+Mmt1rJ17LLlv5yQua2/bZ1jirguRihp
VQhpF0O7b4P8CmuXta361fM7bzUGJwo8f1oEQeDxjw4Y0VMvMfw40UPjN1U0
9t2Onmrucv4LtqzanlmioE2M3FSioe2DxSZFnEDlUgx0rrdKPeIKDVjz4TVA
sPaE0swd75x7c9YzixhWMDjU8zgx6EPB1dQWJm7Ov2fnYgCnvl7VfhVj8fuH
6lcSaqGOUtxFnPuVnA2dDnYUigrcMXbRdep+UqPHDxpkwyEjOFZREQxmijlX
451F3nCOMYJ3ETjOc8iygkP+K2dWi+3PgoMflh394QtTFrgYaPM9194/iQa7
+ePvOW2XzHQNzKqzqKGMoYEOFJ0TmOWyFNBh/s4Cxek4dOnLxK8k2hBikn8R
FevtWIUwtHHlVrhkc+YpC2iLgyVeTCBSTn2gF0b/5mL+IQDBpxEoLBZ3qM+v
e+F8u/YrkhT7cc1f4aH6sI2ZvmAe34zvUMqOqi68Ak2f8VM2f+vrU609Ftly
MBJu/H1X/GhyRLFpbRkTXHRv+arW4TCJjatHT4QZYbid+qxqkIE1fhx2UGXG
AzGJ5xH7rnS6PXzZ0vWcbjEfVS1TOEpsJAZlS9sVYhhTgPEkYRKIFsX/W2Kr
+fBUndAYuEYaMd1iQkd6PX+8xVCsaUZ7R/ArAHjnQjw0ZL0qTaBC4jmC3ESv
Z+s9UI7HiP/cb5dn59Ux7udmNxSUpYhNe2qc0YkdzPr75UIvmzNhnhGvTQp7
QkBrdJeP0I7ZqnL1blHqALU8o+2pWYEXEVpZXB5ARo+U0r3dTyUGz92Th+d7
j0zGdwvFkczzuIfu/H27AMMhwb1/YJjlCXy+CuwHDOi4sXj1MAiTKHVqBt6W
9bamg8+gmXqE/gQzstQnKm88N5CxfkiO4U4z46ihqRLz75yT+XtGLLXUkko2
Gy8x0tqrkT5Ko+AvapwiAqUkCcGeWn9K8qH7KNtOx+cb40KXpNtEDTQMPDub
eem1Gfj5Jil4Uq3yFBLsdMnEw5YbgV6Lp0N4kyPxUY4P4vXFI2VuirB2SXIA
CJamPgem7p+Tf+jh9xBOpFZVzDnVtKf3CFjjDCg/1d+drs63KANzlkmgmtI8
jqueUqnE66TUP9+XJbNArKTeB4dRTppSuqjgUo1dmWxQDuei02QuAu7zMkaK
xQl9qHLYUvAf05kEv5NyfuXvtY+W11wwaUJ6grII8/lcu4aF0da76PNNv0Ac
tgEFLd9A442H4hrEWSSUFQ4Zhha72xZKJdoMHNT1wQcJBcqurRSGCKhF88w4
2FucCYEr3JGHGtmbxcpvqDZpWz9+hZEg5z/fWxWBGHqYSvVmhCy+IvXNY9Xr
DTPzRocHvJGiIYGloQ5SLQEU2GJ9s5V70HcdM3zv0QFDjH9LCUwq/vYhZbQH
lXKuWNZIClm09zITt1sJnunAU3lMmmT0uygX7IRJogoWLaG4ifzkxMFVyLL+
+LvkSVxd358GyTpbsXeAVWRT9pQcr6fhopsrqwYF7i7cuQxpe165qroI8U1U
F4tKvF58QcjAvyVl+0b4f5PYusJZEsyepmy63rhza0erKZsfOVPmdS2nF5fA
VXWcvMqbiD44A1vWGZtC4QW/80ERQbi1AMGKeaRMww3/Qs79AjIeXHRWAlxb
fuh1G2sToFGH6XGBpJF27BP3d1CAwOIEJs2PvYhC/IuRBibPm7aBOf6lPcBw
ShOdCQW37qS01zF3YVzj/0DysuEGZvzzABKK7v7ZWdESTXXAtoxR6Qyfbfux
AJ1O14KQSZNnfdqPXTsk0T5MYnDQIkvoCCPAihSMLto/ZmdSZEWXVx/2VPYc
O6oPyV+MOG3af2wo8vWtGaDCeCQ/n67PicR5I+9RVLsUBzC6C/Dr+fXFne3U
pNszsZK7TtnEMRL4DYhov/E1Feh4+t4tXX9q/lCrm5Fd4D8uf9WiHkHi+tPL
EGyLqHxj2hnL+uaFdUeWwcNzubgwS+VJXwF5V2ezRwN36JGSOoyLcihkQYWW
cuQYs16rKyCmG1SMd5GY/TPT18uPakIWhOxL/YiZin8GZSM8NcoUe4KsrNNi
UrLIJpX3DoSWGRCizKr0EXxYAt+xjO042fqI88yMMKRrjJ/lWaGiRZfbDIDD
k12M7VBYH1C16EIwNI8/l9mWCpEtMD3TuZAo1CRY89x2QO4EHAoUY1KBg15Y
B3/X3buhid6mXofY6rHJedGwU1eJKXLXv3SVWLrWaoDo5QBp93nIw6h/rd/Q
hyzxOWszI7ZU0gTd0sFli1cuomxGZ9L9Aju/xS6fKdAfpQSD4GKMw9SPSMB1
psadZ4ZzpKH9tiyfsCrgMm6lFbpcZ6XwY+xNgd73h5uTTb2/wf2z3d07ORFn
cIga2FLzxa/xepetaTV0h6NVyTMzp90Ruc2MoatJgajpmz3n0ZxrNn7mEtaV
IvqlKBzPCVlsArZLHb9iZDoG86Y3nyfxeBPvd9VRoLo0YgLyjvwd2YLayhT5
oTd8VaG2djjpJTV9ys4+FTDIxqHGXEn7IfLFxvU+uL1eIgsDLaKwQAcUA966
MSPbPC92xiyJ5kDECaKhnrLa3VNN3CoMojYAgcToPibxJ0OjO8FJGBpRnnne
YrItxTRHov3ETHOC5sdEXAXmIlf1eLkYBZXuqOJsHBTsrTbvg6OhiqH3Ab3C
aJeN9YNrDN/Uyqv20vTfnuj7evw90QpJ9k/y3ZTdkHNNxpYzb8efhYJKepKO
0HVutooD70uC6d9dzZePpZOlLnCYOmZJLEPGFel0KNS93QaTpTs5sWhwhpuB
WMsqeV6hm7O+DdvUpjWtKw1eRxG5c8Y1zw0Y+fIQJMVaUdnv0zqpJ9IyiRPk
vmNDTCbxORT7wUijIxXVGWht+GGAuprdbcBLEfaZYbNE3aeAl+D2nWd6CmvZ
jE6O+hSsMR+TAE9fg4IowAdjOGfgqv7Yn7p0ZPQUFVQiqekcyKfONxJtHgvW
hrRsTFLMzUfM9FBdTWicJ3f1p3Wt7N2JZd7Si/FSK+hZv/YnRSZ+fh8M4Xfm
WrKCNxS0oIM/LmgPjxRtzJHBEydSe6092JiJnGv1gFTc50hsUZviLdxAOzip
AqH6Ok6USlqLdtvncWSH17ZUGe1CCtvaAbW+aiDllS4vFh+OUVkAzweV4COW
SAcHB+mZ4Hyxn/bSha/xeucu6jvT9IrbiyZZUkY5XNXXmrhJiHqoaliMEXKb
QZPbB9Sp6I9H59s+i5AsQV00RQRXEGdi22sRgQz0M+NSIdkorVWJ1fKWSZSi
wvAL9oQ7A+l9RSxcwYsmZDUILAQzXvHqID1M/WpzGi8KT1kWgxR0m/yCfAsB
U+uaM0D89REGcr2cv4qXQCoCJd8n4v3btno3kWDqRK+8Efy9O1iah7BYSYre
qB/mbtdgO/jKeDnj3m1ZElHUEZd7aWdrK6GoOmluDbZMN4ws0DVyHjyc73j5
DzcCZ1ylbHsyNrjHaHs1CKpVgAsOmLPImQbf9Fqkvcded22RXNAup1unz9iT
vHElpBRoj+2HctAjiU0OnkoYtheucHbV9bAq1hohTDKlflhZgsNa7Bs4Tgob
M7l0DYuXBkb2jA87uB5ax0cZ3dJFwa/3+dxMS+9NrHEvYNi1hRpqJasV1+mX
rPk3QIE/8qy7rDyRD971VDlgCZyvxZBAqYItadG24oGWIa32DnxeFBEQ07kd
CpYPtb4mLAoHJPyE6mIHTWDw3bJbHWKC8suYx5pkyjecKzve0HEbGisUC2ZI
zB0du3HiKwjIoN+ksKSzwRnXgfOQ2pNiloIOwwnj7ho1XAnGEGqJp8VOF51i
PYXsfaGqmxulJRqZXzsAOOKvR7D9zcf56135TduRZB3TTzmujTjn08ozsR1v
EGDUwmGIGxGDvuDBKhq1VnT4AA7coXoO7jYEuBHAycaq02o2mZYPnVat9U5J
0KxBIkSQcEaUXcakoitWeg4oU5dX3DJXzaoAcKoY7NDAE8ASLncT9L/BeJae
8oae7uO/5wt6eyvdmGUiZ7UgWChQ7K2zw9kqRNHg6ZyTL7OuAggkw72bspC9
N6nv0NNVYXsMqFnq/hNvfoAXJufDcSyy59bVwAD/DZy4FrDV6ILTQVWPvkso
56xisZNjPhkL3VxtsbSt2wcQK5iaSe8Xa1uNazh8e0uRnCm1iilRMpWiqkfu
lwTPoPuuMAFmHn7suRqCteD85VIiQK5hqZ77369AIuWgeYW5aV5ba1Mwnf9I
Ow9Ex+R2oDuFhXG5O+T8Q1l9p9OBORXF3XjxJUuOvgYJ6MvY6kxH84otvxk5
T6cwTpb1YUUFjpw5QHM+ur9PA7CCGL/qV1/CEK/pVt53EfTpnwhakotxyaTy
ayyDapdphSIIX7+sXUPoakp2kH478E+O2BZQhg5P1SPHX1IfXG7AgfFBWhhi
LZHwt1eyUT1DURe5SobXcKq9zL46RAYUfDLgRstr5ZKszs/NgZVXGAXmWHMa
6WUxmats4iz1Y1WBW/k4JEcuI1MInuvOSYkGDTzpBDx++21z0bDeJA3wZIqR
V960mZdE9E42tU5Yt5OEJWCjiC73VXmLCzuzz6BklYhgTs9pIslY8K+2fiR4
GEeKjgWWRqU8lb/sDFhfQlMofjjCJZuj8rrLyptevGox4S52tXW2ibAr6DG5
iQlYt5hn2VwiWmNH+Xi57eAvvfwhGQifoT04vGK7ef5/2qly1tj1GpxL0msn
94B0gWJMC3FlCMfaXUkEsNrucQWkI1PgNmfZh2fdbEkmBK5Q8n0UZIbtej4Y
STle1LvT87hHH6SQMuwxXxx1HBXCAGzK+OS1ogQpx2COSBclyLBXwlYMdPsH
gpnAaLFDlFUzGctqvaE8a5pqo4O5jQMJc0d3C//iST6nURjOIGi694KDLjua
QuYtjzrLX6qb88eirj7sPx1wPleZ2tM9XDgYF19ymQ49wRJ4VxiNeiF2bH1W
jQfLd+Il+Y3CnIdbbMtZWQ09MH8J9OW93hKYPkUtbbgOcqggSNeGEhMbT2hn
usp8Np63GuNb8WHEgm2L35If/gDcQdS0sYBQJ7aHZq4jxidT2lnZTq+rpGgq
ZTV1zjO90Ibg6IaV6NbA8sd0AXjY2vxUl2bNUTU9pgkMAEHsgOJ0/oTQwpe3
DsH0IBSl1V0E5Rzl+zLOcUz7mL/KMNYCU2hkgytRHzziVaikaisgHFBjB1YZ
TZZIax7/vgaTTwi1CYx4MU4aE72KOPW71nOoxxDL9KmccLEbzhRYLKkqvVGp
h7+auX12Z/FGS1Pvf1cymqRjexWvx2Dd0UOX+mUbhnH583JRX2XkQcCrIxK2
8cw1rGfx6Sdiz4Zk00FHDJOqNfDW7M89kixYUSc/K+putFiLV/NLx2ManXZr
DLBH6xSFMEriALCr0dwTL578L7hN3GQHy4yCoOgscO16nSghmA0OlhEp051O
vNDfdMI3Y1GUmGV85ekwD0sJZTFBJrVlAOuv3I1anLYN2pb1PYU5+plufacT
cRyAyKt3drhO7uoY5cYuW9V5cGqaMWsBbcjhqIwAJOIMVveiYsNl0v3Oq7d1
JQMLy5+gXw1kL7rEHWEsN3TVVu5i/kEhvoSEEmEgGcV/SLSZ0MTrNaq17hmu
HqbZ0CNkF5Hn4uUQ+/vNQs3RdZyhw17a+uOa42Xs/C7YkT91yl13E7Im3eu/
cZMPWggTncIH5LrOstSoY6OhufVoQuEgURsCk2HGBrbWw9YjOjEDq5dg6aXU
uH3+jqmTjBkJWsqLNwW3Ah4RLmJxTZYGWk8evWqt0+0YRHCzefFW/9go+yQn
Xgf28EA9oWG4V3ae3Wwsn+/nb+ldWKRVoWOc3+i3amwQMi+GWF22ayAIZyXZ
3RnFZOCSb6qirP4l2AiagDmWroyxzM/IvGvAw1azEKt3jzE/FsXDJAQw4i7l
0VFjz8lWOHpnXmeSLSEgE04QevZjfiN0iT6oB2ZAxnsApZo2YPp80+6dGt/6
mTiUTKSmdNITYKHisLoIv/+Dyu9WOJje9N8isB1RW5PesjTuLcIYehnp7N8V
MwW3EHID4Ihbz+c3au2AttRjjCzuuWPRV25qu9SmOZVtUSDw9uZGI7/nLedR
2UF86eNAUhTeJYP4bWwYCXtFXxcXZVnHt0ayTIjiXiejXfp29i/xfR/FfjRv
xr9WmJgM7d+3/IXDZBlXDzOh45b9bDQw+mGAswBUP1qBhs7GnXHMJkvlfUSa
xIXB2awaD3AO+U5PSP1odNzvNVVNmDljXXWjddJxCW4XHMtvGmHwaGX+zHQO
fOLCKSnDfqAlXbWHzeAkqr+LtdiRkiRji4VUoPHEOIBsfDtxPx/KTpISgeGj
3UFCe9TBva6NOHWk3zO8GanuPp/HhZGoiSE6Cj6HHtVMevG9vBFIb+LL5+Ti
/4XadFyPYJFKrql8SFrE/YxLkhmnzwp91Iosc6s0Axc76lun3ZT1SWLFSsF6
63Y3T4IW5s+2G3G7alnh/n88+y0YdY4Qk2amFuKeieq7QsNeJxYy41qBKyP7
xiF2A3KHLz7n49BpGqMfT6rU2Cxnbs+9cu8z0kxsZISsBjd3fwV4tOTjzCGE
S9YVkGkv5ln5R70kvoK0kaTQH3TeOIt7XJm7UTjSfIWcYdufISfLp4xeunlU
LeEjpX4sbY5P0h8TuqYExEFAn9svM0PaJ7dXh4YZs+e2Di3uFFK90hUpOxed
t5WIkaEc4QdRK/XNwOLo7WoX6sHGxNDprUu+3RG9YHE0KgkDHmhON23w37Zu
4k0PmvMcK4/3S89G4IxFyT8vAF/h0BsX9Fy+8ORIGQBeGKIHnMcCUCq4yPzk
cVHFtntfj3J6kEbLiqI8z24wWnttc6Ll5OaDiUPhcDVcwtUm+nnhoxjNWmwY
+qp17QEJoPc1YgyLQvk+tKkuKqSe2vMyGK/vWIBuXlIz8gCVjy0TBsQAxDO4
B9N7Ie0f6clxtCM6Ei0qrQpW1O9z104XiC5yWNqy56nYY4Hd5/nN2suvfieK
YIx/NDpiVrZmoG9y9jSl+NKPTIYN3CupVOsJG2+fNSo+S+XCGN7vbysibwI1
5KlemRdVatWMETcfFFt1jwtcXmjEep5ux+z0y/v9WJIrXI3yyoJR5WnFX/NO
PNCbyWKlstvSPRC+J5gj6oiasuPd1HZ5f+71IFfhvc6M5sFmu7hIwNKhzz+X
k+QxR6ME11ygFmWyhiFxbg4L/XyZ2EbFZ0ZHzuP3nr0u3K2Xqt5hVHERP/9j
074EsJvj8tuQX8iZb1M8JD6c+dW4cr2Ep7oq/+8w4QoLnoCGFeCsp1HImsrF
CxRDpL7DuAIapLRWFOiY4AJgwGllbLNFzrLNV0WxtTVgu1hJIowODAmFupSp
qOQOw39yamtpiueKAW/oKR43tDTkYOHgZmznciL6JNAq61JUDZFlEBmb4OPy
ISUSsEq53u2qxLXGEo5dsIoCoIAgFmwcRYil0OL7B9EkNQhf5JmMidEjlKc4
XkmGDzcfiKaciDaNhW2jDrXjw/Jf8r4tkNRIv+5mRy+tcrm2RT3y+LH2oRKF
l2Ol3ly3HjTDCptcZYUb2h0xcRtO/02/1GK1/wWJLfC3m2mBP9X2htCf6eSo
U/D7UuAgI9PWax+vLMirh2nzVjJ0obpESBDf72q03vt0omxFru+eqD6K5wVP
98xVf3aXCykLa/CiOHMda/r78qmyb6VYZYEyN+cbj0AJpYsd3JVxZaV6qd9N
mWrYfUVbCqPQFyCAv0eVoKpE31UE/9vx1U79RVdvM/qU3On33EEwWq4QGAmP
TRFUKihbcJy1QPoC1/RUR34fXZRSLTokqHq0NqVnEd24vaEKAUIEDgjQAin6
ltdGleuNAxdXsNqJIeIyyWF2WOxEuGFlvanyScIYmPisGP2O4VNsxLhKVS40
NjtKYlOf4wwEEmCJme3d2DHdyV7woBzpKBHkkDlSRvwjfzIvHYXAwFgornE6
Y15ZtxPvZUDnSfNRY4tq0oJRlB3TpytzCuvy0xndqfLNQcP7wXqx3VYLwM9g
A8NtUyLKyAhP/PYnvOjJWrosKEll76ONGwTkar2QhdtbEndeWT03sIi0AWx0
xPLGmDvFu27wajs5WmhQ6U97upxH0aHdP/tKaltSJrm8M9u23TpoKfXJSe50
kB57Kd/CbTOiLreZl2RDwF9QSdqU6NcM7N6urBbL9wBVqN7++sm1KBtNia0f
u7Z3/m5HEFfwzZvmiGnUTwjU1VmkTalBf9/4AvFFL1uTqlSlKvOgfP8Pkqkr
lUECkRi4CYeIvWIbmOgI7MoXvQd33i5F6cOytjJLbSM8tqCBHbt0qwbQVz+t
ZruaC17y65JL6QDxNi3rOmc5aR0LnsLhCHt5oMSLqB3a0yKFHwBcV8pIFG/Y
15GN3ful5A4GZcw2uDkKYKXgDBB5WlfqewV83q/2XREC7IdXIeQ46kfAo8jo
AkKNDvuRJEXklbCvybaXUdLkOiBjBM4jx5DvsG/3KjbKS8XpulVRmYZL1Q1X
Bj0Ls0cNFPWox+0nQO31EdWX8EmOUmJ8RK+tAqgUyVYTcqwz5lQ4UyineD2n
hqxtJU05m9Umm1oJCko/8wqm8dLkivA1lDZxL3dY1NdIT51YgTzTgqszAryJ
UZXtQDrsHmC+5ZQbiZ6uafk8VHEA4eIK34EPDmCFeRW2eBYJvwLZoZXmCwUM
OR1gR4dUZ0qO4hd2KTtKbPOCwe/bjS0c25q90NBJ7vw49E50o0ZaBxngTga5
mrWqTIHw+gbyKB0HXLXEAoz/jzHh8rUORa41acC+WcRcqd+9Mx7/Hnws1Xuo
LqpBPQ4MRN2bWZ4xMNqbtoEGM31k2L7Eqa1CGOnMdFY1A9J6FydtlR5Js124
RyDH4H4nPDH2rwIfz0lgt3Qo2kFabk0NxBlN3y7ylS2vJIUNLDhstzmeQTvY
ljay0kbe47NhqtQPmInV8jLiHVSMaWZluxxfGpUI/iiRBQXRkPlcyIS+G8kT
zqWJcXho1byQD6Jx8jdBr1j+rQQMMbA28GB3e/pfZ4zXPzs0YQgmkMrPzWrt
VvVofDKx6rSllAm0c4ZExLi3M3hc9FJgaey+tQ7bz6yoB+sl4Z21m3kdwux1
1biBX6GXSDMq6uwMh9mFp6uPUc8xlb8SCMnGmlXxVtf/2fpcBoM1/KZKeLEG
wSJ0+6kaxST/7SBrLINH6b5/doz2/sVBgrv8abS3FAuDCxJBQ4H543uAeNcD
8IyQ3CLh3EdOdzJcoiqRL7/hEjWKw9aSAf4/x+sh7zglMD3av9WwSykz1YbW
WP3d2QD9glzRk4aQ7Bvj/MxSnSlNhgDGU1AxLf9D4dAyVugc5xRwUS//YDO4
L15knvcY06UmltJ69NG1aW6LopQsIAbxPKAs1GZnSmNEV0x6md4S4KLNw00z
n4shsXk1U/NkCiGmLRddbL4c8mBNib9RbaYj7vLJfLokZUlXDbxdHa/wfUzP
PP/+ffKikHgryqRtCUsZPq68Si9DADqbxKpwtpQOQh+2zfF6hYQrT2up1MXi
0Txfqd+sbNjm3fmOMUyDnVPbdPkU05NjNbF1AF3eOAvVZvcHb0uRrbXmxp9i
3005h252UyrvcAxD/git3s9pnqrIW16tVyO8xCm7nifi4fXjb5xB8XFVCroh
emdVmyVaIKlUXzPpfxSEjfysfB4CV/Q5Z6TlPj9QMP1mFZOzjPZRvP7z8KBU
nVnfnM4LLlkEUcfYatPNoa9PcaAzGu2DtxtJtGDjgNbdkF9VOiNDdmYSLiYO
yT7f+uBT8c2baAWdq7l3/PSSG1qAsRuwx3bPeVtzKL3s7kSLFjnZX/GMHyNW
CmJoSwwlj/xpWie+TU6mHAJFzy5sAkzls5Z31ibjqXFqkHnTnB6x3/9mqGoX
q3NXJluEGaipOryU0K+Lo+igom164QrO4qE7o1iWyByMYSMOpqNKL8v/x3xO
n5uDieO6bvhLmt82jnKJUNmPM5tE+ZCzHQZnIFFaBM+tkAxhH24RqOTOfPTh
SMkOkDeDKVZb0nDbAZImEkjcsv0tIOn/U/XWOBO995UsQ36tDlWR9f/2IqQs
/kmqLeLsnLLeIxtDv8QYRzFNcqfjcR/7+whM/IKBxBR379oFV8OvmjA0Klle
Qybp6BU/7yIt7KROgAnq9EwLLpsRixzuIzoDHFyzzUeZfBEXv+rm2FSZjJP2
FtioWEzitoOTtcmj5ne6qPveXdkEuuzNm57CqGzNR5yL6XWlIO4w2aaU/IYt
C5WtWSdxqQMJ8HSaeiL/wTqVrjY/eEwf4DD6DlVn13zbl7hfDLRdg2kwKgXi
zjbGUSyd2wAXhygeIhJZBzvIvd2LGuDlg3wje6R18a2N9qTpk/gtyiet64Pz
18og7hIXke38lgXUe0WlIAZeNcqPAsAA67FpSEEq35YYPZgR3VP+WIrd9QRa
NttRrZMXuKq5PzJynll1gXTlgrxxxHSRPAN7QFe+yIe+AuCoI9BmSxm1JHAB
PdzSZbcrKPUfSoaTlvb60QVwlzb8APTSAoi+wC/J7+1w6jXtah9UJsGqMSYU
0TATVyZUOZaQv062uYFIuT/knTRdccwJf8sRr6zcaO560EosYE3ICZIhJ5DL
TlV/Os81MZONpansWhbC+YazC3wNgZGWgicZ2TI6VC/Lu00c0lbIJ4l8/N1K
uS4W8wZHK+iXIMGdkgyaIOwXJS33vNB5DZj80xrAp4a2WoH3rjeIEenUUull
AobNBm1x3ctyugRWWK1LRWFsAXymtk/Mr4i4VFAzjgblDSvUU/PI8n7MYvdJ
fyLaFwYtcy4RgwpstYZhxdH3ODJg1RunHpn1jFNflLGfAhMhcP1gKN9B0+bD
oJbrDUsXiN/5ZDQxKSe2Uafx9JkkCyyP3T/0lCDpJRnsLAvGXqC65VADxt7E
7ehAAmxU/YXg5lw3xjpmkmQtK8HQRmu43j6SrpjvUqfhiKDGQHIxnnS1iz67
UjBqsOrfNoktAoGBJTDl2eL+naGX05x5JpOnEuaqI5BNXtL/OK4KFitWUwbx
XXeYvHkb8PjpYyQzwzvaqvaIVMbkLuuT15aAGca8gdESzMvi7MLk7JI5zo6d
SJYfs6eCLYygLisqSzE8oBN5R/Tg3TDMH9nWT2acJOLLbSlyYsfO7mZT/cZK
k5PUY9plo5g0dr4nF+KrRR26cuqhnVuWARKPHU1kZJKi2+bCZPgmZt2HcXYh
cfHCNsaj6l3k7t5z+VPJVgN6by9RNJEoV1f9d6dMHzb0I3URH1bfjFc/VhWs
/OUmIH/C+Ndg+s2X1LVzk3zh38KlXTZ6R39liZrQbxxVxAqKIEyqxorOTeAX
0TwRbG78eh800a1jHCOiKhIInh7M87prymxgSOOGMVjrPV7a5/37mJes51wM
Lj5z/zH0EbWREPDgzxz9s+tzDjS16LymMxAAjCy3L6ZPaOrq5WIocywJXlH0
Zv5x+I5vCyDpFPerGXZjxLPmvwHL8NSMfyhXKgcpA5bqNGr/BCSfdSZ3JiBf
DFZ+L2A/pt3dUSEzLyPapRwebwt9UptXeA9rIfhlXqFzzGUaXGHjw/pqFHsb
/ZSTdlOEaTQ0GgV5DvWn4z2Wd/FP7xFhn9a/tqP+2Swa2qQtaVDZU7wfkxCl
aeidRh+w6VwS8Qzq6OlBwke+oQsuzNYZTrc8Hl41ygBuYqjAjsbjyj7L+1E/
/nn62ZX/gEjLai+pHZG1a6qk6lkkLp+ifZU8s6zAbX7yFjoqKgzdY+MIM1m3
kk4HWmY7ldfXy/Vr2OlrxD8JJcxPWYDuHnDzW7Mq18bsJSoEpETf9uE1N71P
ncB5Xglddz2MVwieMkQF14/uwuciZa1nZ3KzBjQcbjYcxHjv4JIAvChCEOUx
Marc+teuub0Um7f5Ui9WEYgq1Dppd0U09CMnta6UFeoFMDcn2NJvVnm2quqC
HXa8v81pBZZzXk0CXhbbeaVtu+0mUZlBu5uF9m/8/tCyxkvqy49nYO3ZNz6L
Ie+Dl1Z/xexVPXlzMgASMkIzeyQYxkktYy6OF0PR/PbpVQG/RFhM7YAMa9Zi
0cpURfDQX6e8+TUBYo8BS4wo+tRBPwT9eztfgx5qghT8CO9jHRVa7GtaN+HJ
1hanq8sLvcwjG/tLkjdZcXYOkpmEnwJKZiZ5+4OM1zdB8WRZdbSpR9PLZN+B
diKyn7dxZyPN9RHxHjRIWKhG0GUE0IjH/+qfpDMY9xZBurbSAZfJaNJL8EJe
z2aIoUOWxOg14gVRWEUTW5SI8E8FUp9EEyWf0mNFPy43cqTN9bNLVTJKCmKc
yytFSa826BE7qxIkRKGGR4CM152RQSdWtJly0RuEZx2vM4XLLFbYiqNBtlTe
vjUJ/xBB4Ws0c3qJ7vmb9lWm5JhvVs9vDsjIJvIswLJhgLdMWjuSHR5O57ec
ZmLw+3xCpKwEzVKo3CV2PdN5m4asDxo1Hrg9+siimCoZfkBKsKnT5eOqIOgM
Ez47Ri59sNzAs9D30QNVvxyKbbN7LjMn+GQupUDPVeAqEjfkRo5XfkT7m3OL
z20p1/wBaApTveB8MIb9PYCCI0K0YR0wFxKl3mekmj19WzBeFlDI/d27R6dX
EPTe95KmO//39zT/uQxMWXUKmKHoZYVwZHi4xyJCTMTaCip2T350eWihsGtW
dYdmiNgdzz4+MDUYpK5exnDekouLLbJcgP4os9qlqUZhmZprCvSutBXDUZhZ
ECktudaISaDY8J+iJLeq4vSm0ZI0dh1RRZZXglt5natiKt4jkdZV49GP10uw
z6lCZnVX5jUT+a/CDVXfOWWx+Q3q2YwKntPaAn3z8mJ0MlIFnpa2noseaZPO
PkvwoRt+2kAjrcL+R5F2jM81mFY8XhAsDvZeg8bXJ4n47jVHzm7hvsOsXNEV
FkvTvPchxXzQkoUKgA4HwTj17O+HlH8NG/Yz4HJfLiXfmHhNxaOOYdKINyVB
qq1ZtUz7nC8uAzEyT6ul+uUBVanmjNdiCXbG5XPgPypz7ri4VKa41xyBc3pW
NF4jWwylE2M60Co4IHk6eUTmFf120vUYM6UoNy4H4KoPmyATjOLfNZDfPwSA
8Gtbcj+2b3C8qt/5pqK7xqyfLBIzfOJNxl6xrxoW2JC6sM71haVfWMoRqTUp
J+bwBS44dHxXSOZISgUY2nF7rKdSKOkeuErCyIi5X4qOA6iMasYGPETxWuAZ
1Rg2Y0okb8wS1Hr281UX7VrTS/kRM17z9Nf6Gdnrdw1IX2IgtLU/REtDhyH4
SGUijWUojGUAkpjb9OQJ9hVgKfeatzIdVKgtQyxScVhJpciG3BMu2NAMHCs3
7fQmV+SvIdFO73+Pzd/pSgscCDLritNohX5yZ9Ew6yVAX1FWjFaY440ed6a7
8l2Pve4XEKPX5Ke8WwiXl42QFPHr6jq3dZkObLSp6rud+q38S15B88ai52r/
D6eczkrfFfmtqxiu3Bg0ioLKL7C7rYBPNOTi71ZAHIL/LTsKweQCwM9ehGNe
U3s+Y+uGr2gAtB/foSbJOUyUbQza7I9fg9QTQWcNiIFX5QrnneP6Q9svmLko
+UTRZ/OQITMmu05l3V2kMTxS1ZPvjq7IRToXHk1f1jcZwgWVdv/LUYIi6MNM
NK8f4BpUrO/33VNPkQJf3XwbTRZA3SWQWYQAIyM1C7b1hyphWUMYQw0q5EUA
8ztQ5DcMbSza8Sdp/RIdbRmouD+bX5OcysAspCBgrJo4n9sjV9BWczmXH6Pu
xMO1cAzz4WzmEGVGmP/tgAGaZBftjHzvSXs4goRkHlTlD3XS9Bze8/q3EYXL
RU7Wbkx8WMEpQECYH+X0KOTid2ux/Gd8iw/YQroAprd3fRZQME3IXMOG0GB8
yZ7HOKwAZGFHq8ijwG77KrTfVxhuCIhI6QtvaUOvIzCi7i4oz6lORWZ1OUPo
LZvkKkIsQyypCTWygWi9UMGamKbczpuJrXdouxcdrhIRx4mnXbijK8SWjL8B
oWN+CbtxnbbjSLqxXr0zMxNx2xjeLItJAz4dbqKj/6uw+7E0vR5pqK136XPN
uHQnyWRsiBzHazhz885VDMKjmyJ2RfmTUxwCo/OKSafOqRIzEDdJ2XcbGhfV
0LmCfUCorqn71DmUvMXDMzWfmB64s9dcewwzA5DoFGdng3A6zJHWtkWbs35J
5Ej+LEmA8tLyTf4YjnRG85cqdCWzP7WGekJKoR/+0dzEwYKEN3DyQQ4qEo0C
M4wZk1EBLUhURv81RLl8hyjq2SANRWzYJX1YyMU4DTJ3OUybs11YrAWhhsVo
7fFpCWzxWoHBUrSJSXNgzXWNyrsB0IjM3b1a2YTmWb4RYXTXFMC33o5nz0ux
qo6ZfRVE6s8XS+1aMBVR6h4vNtz1Aka/OPktgzS+eWfrEQG+LrGHb/XUNC8C
huGw3aQ1zQdagp2yEUSAS40lxrnRikVXwnZ//Ueb5+AIF56ivqfwgTGXCeN7
OUa6roppgWiYXi7u1PHamkGTpLCexRHdPH9GHJA0za/+czS85z1naE0yE/Sj
xRPJ3NxjLhv+/+DXaeueglH8hS0xjJuPb6mdV/OvJT8T2K/SqumzI45Ri6zb
K/BvMhUc4HhlcJxsapt03TxU+PMsJ7/1pOqZQoyeo+gHL+WcS8NCgeWDwmYF
LdfdrNrD8sMlkKHzQmHKouvRElRghKp6qIgAdJjvsi2GBnV0q1u4I8Gkf9wE
FDv2McPqOjHe2nYFehMDWraKZJyrZXvZyYq1eJ4kPrJ4f8uFBEi8yUUw0dGf
CSs7/ayKpJUJDGXsGVXEpL7doQ1isxvta+Z9SBUcnrS52nbMXaMrRRhMhT6C
843O3kapsBpYn6nB1ipqjbkSIRb9jCjuVheZ1sXhnjYHwFTasEGh4PO5qLqo
eYqSDFwjKEaIs//kEyd4NGudnpYS8YjLrruKag45LgxeE9m7XTuq4qNNm0rk
QaIqn3RZDnrAgHpFCd/EdKN2FwNvoYQPveKNOeyBJFZJfX4A/fPV6LGmrHwQ
tnEcezum8h4daxpumMdSk8sz+b99kA0aU3UFM3B4y6WFe5XG4apIgzJBiY+a
Mw5bp33xrP+CI49uknunbhHLJIcLGjrAvOhWFeqU8QF2YLrT+DWZlZGl2u4z
cuHbd9DomG3mYg2CHhBhpJpH3V1z0Q2dkC1OWh7X+9IHtkCtnPLym9uGLvoF
nXTF6Q6nA+2zFgH258yf0nvkVInAOPMpuGltxxiaKlMI79fdDVesojML4JJk
VWv+M6mszjoQA7P2km+cgRi5YTU9nbrcVlE0ZopcS+sQB+2Yg+9Tw4j/oShN
dWNmygq96kC5ecJiC0BSPdvSPvxh0sE56nyHw5vzL1NNsT/IzBbO/DHoeOLg
YGy9m3se7+459nqyYW7pql3VCP0wjQ9j2zDawKfZSOQqxvGVGI9AwwmmDPxR
/YLhVTFCozeqO/biiq6KcT1GeGyVLDp8EKpiC9OrokBiyK0xevf6sHgDNMnQ
ALiGzEcaaUMTT4FvKjKHTA416GuN+xagGGcb/Ihn9bISzeeKc+B4xoksXsjh
j37bYuL9exF+ntMW2eLW3NGqQTRKG9b6XjFOAS9dWuaiHe32bFHt+q662juQ
qfMGkP3b+8XT0fbk+jqlQmbXJXhC/dEm7Mx9rJebDuz7kdwBK7yyPwP4tXAL
OUzH74NZwuem6lMSi6dkSq13tYGoAf6x3Ixk7hD02KXO/cG0KI1OKXQaJqgd
l1ICjT4yDkFvOKW1UVV9Y2JuEWQUMJIrxbDAOab2IeNgf3mBLdLPPn0Kc6/5
pcPkhVYDOqzTOtzWhu3BiXxp939iYUCtDjiXvTQ3OzT6rI3AEhGiskV1Fl+N
eedtxA1V48f9Rx8WdPDUHUJGndW3aqvsyeVm+5tCVXn5hKmaU54nW0bYe5J6
VxTvOi9zgoEo46Ffbuk44WBStHv0bP7IwtpG2k37F5JKv3kREIxgENoAJYFG
nBRpR1gZsL1RTq8G+gwtGtCwHq7PeGoZlsIr5z6OdIu15JxpP6LgyS8aPOFw
loRnqI/vzpcspOv6gkdde/Pa3qVXg7SGGTFmFMRCzp3yUIHCZDiTgA/xfkCt
S9x3ArphrlHw9hldmAyBa5i6Z7tV+On37gA/xHo4cJ6Zl3bF88Idfu7DoyUA
UBTfovIW3Y2kYAVHugiuO/1Q50+6tQMWUjJ/7lDeY4HdJV2Wb3KPA8Z9uPvg
3waAYbjtxS2hin9s8lbwrGHqfun6xNBooDc386C7pvyavZsshqWlLzLCzlsx
9XSeEyt+/fZc1DZA956mbuw1QbaztglzpHIa9jVpxc0d39ozEB3JxEm/PeVf
n1sO4+NkuNRZ0g+UmyrE1ktJmuhMa8/ocsnhuaLU2XtkqBY5Dr71R55ISe5m
RkelKQFzRwQvK9XPhf1NZZKztQUFsSnO6v8tPGQwxcC8vJN6iI1GcwG+kiq9
b+tPoy/GT+4S58bajT1djr99s8Mp8AIXtFeD8zrrbBUZ9iT42zW46yUoPyaX
AKrA8cz7DGequJSlFJN1rnOkZM0NmkUGnUf+qf/koX9tLXmhsymOXXAKYu8J
ywHsCo3ZhnM6yJBRqyUhitnMfWW6rvhCnTxIKJT1vJ+v/3tXgw+KbfCdRZw7
aE8qcBuQhK+yCAMgMQtiiNTuBrXiKYn2gjUC7vjM9u759zA+gIONlAkBz6Zu
L/09iAzLyosx5dSVqm7q16hwNeAJBsOvYNsSorwnF8MO0F2H2a+0rftEqDM5
z3owp6nICuPN50VxyEpVYHIidqx2A/+IvW9mt2GoDMjBTibHh4IioSILln4u
d4KXQCylT9DDfpO9Qm24zSeUbepceuCV912wFj/ayQsIt3ZmmatisqDz0A+y
XohpQhJrUqQLqquU4fAbnWkozmG+SGeHrYw0V42rziD0Q5qwMQ2BfHrjyxZN
w8hKxBfllCdtD0zbQx7MBNS3J6ZCi/VMxq0jecISiQmo5poA+NcmbcNT2JAA
ou4OXkmBcMI/g7u+6WX5l/iCSSRCglx3T8wZmRJOJjGeXI2NNJZWJ72eq6Nd
pppJDOXcGyYuuqjaWm2eS4k22wsMpmTOeAeo93WbC2xWYARS/al8/GNRLQJP
sXv0N5s9nJFvFYoyuCvsWKI6ov7ufZKb9I8BA3V+OJqzKf8N7aIc3puouwBG
Yb9JlQ9q6ay4oE/Ei1F5eJJ6NMHKJhifJD43XD3/a1FMazTf+IZE7G0UjYo4
xVf6ms8odVMJYGIjFzKWeWCvy2GwRDA2hNsTjxiQdjnmvW9gnpoRY+HxXEBj
rVUh1/Ml/7Y7dJGlThK5M+dKhGCJugaXqN3t+YZtbLJpbXBOSZU995ki7i/O
LAwc11PQnWnUcB/dEGaHMcIQBHVSnv86ZRGqXtpePSLP9LDAfohDKdgcvNcP
Rp7Q41ZUCXqUJG1z76RLmRDxuG97AyplR2hnbxMaMFScmt7Dlu4PflM7c7Ay
Oxz2BHk8r+zV9Yp1k7UO93pQ1wkNIThH+snbb5zOQcMaxqC9sdFi+M7SAL8d
y60DpT6CR5y6dvh0sdtu7h600uj2/8XVe63md0I68VdErZUPRdcxGRZ94Qp1
K/sYDoxWMKTey1vkeFzePUj9R3n/02SI+vtbet9S0EGDIoyadTj9svN6fXPj
zvisuIM7xDw5Z5s/vKqVC59x1dPWzvT1d55K8ZXrdaLargAK9UZDDu9QIW/A
7sMwFhof6mXh4n+eOdc7F/XNhKeqQ5cchILLUOce7cpv3bg9Gkv7hortDEcQ
EOWp2XFBCqHPiDJAl67f4irF7FaX+9au5zMKvObbjGMWYj6k9T6qAyCUlzSy
CNJ4tXNj46YvkZFLhOWWpSwMtjIJyvvSx3Y+ILFL+Qo03SSb9gl0zKuFU8iU
IXJ+CsHeeTdFyOHMeXudL99BRbVggITMKpIY32PM2UmuHb/A/hn7TYBtDFoN
wsVx/135nmKSC4sa6SAqduSPJmKVHvpWvuEdNGRoPvvcdKrb0payG0tBR1Uv
9ztjz1Y2NJNciR3OYUJwbYKzvMmleHNnlejNzKL652uuSv5S/uzaeQ1ynp4t
oec7mmJ4ppp98nqjIJmteyCQffLRlDsdbaQZJslM2CnqAZUbCfn8MfttJ99Y
hywGhFYowszssEVclMrvC0hr4auOiAYke+SwIxRyYrCawAz5XlSXEV6JFdnz
lR3+zZVPJH6oCReSBbgmZmE9QiSvGtfDnLWvr0qYoGz5MfWaof96VuTZqSpQ
wFvfirDCDPtDzIKbuq9kgnp6NVCtkSGL1ZdSgGSE7ANLgbTYM/PCWRdRpF+H
geHjZIZH5/hNQPfW6DzqmvemmyTwBroLR+FncC5YCvLHbWiZRBf298ueJBgO
W46HJN22v9ArMSWbpbP5Gvz0kWsCSUBYxA4zk1V+BPe3SjgCihEzCGEj5uMM
Jh88Gs7jlItM7NLtkOG+MRSC1rC2vxPWRIoRM/thHyzgljJ15F7HDaAWn4WP
RkJGVf8289YjJmD9wnf84WWR6YopWWf7DowL4lfaF8SZ5LT3sGIQv1eDgB1Q
3SZxEK5mgxAG6N/cyyq+3HNKRnlFcEwXeqjorhjqin1sTbSxv8P8FeLUUjIY
5Q6EcaR3UZs6H8cE/NYHazODraAECaRkVA+9UChl8SuL5bSwlnHrckSefPVq
68XDO94U9xtBk1DvdQADy7w//m8RQaXGQ6wlQFBCrNR1lN2afeODiGyQ7cda
hIsS6GURxJLVJ9xOHFhW4EFmHiIbl3ONl8ZqgMxPG7fo74TFyhJYMqs0edPf
0hVTySaoZCgkrfWYD5xwzG/JyfQVlwU+fTf/Oqf03mA/I1uIWFlEQiUwTu7v
obn4Y8IHeyXPF2l9DyEteDd+LaubER/tJ3hlpNaiqiemRhm9SKTAwzrKQQT4
fsawRcnfPWObzGPROvp1oeIU6XLarpwDvTpb4AG+Z25LAexncdYj7rC9R7rR
sw+0oGoNXd8RyqTg6ufLYLylsowk4zcdTfwNky7EkgGyheR3UW5JBKxU5T0b
n2pFoP1sRJD3Td2K8XAbI3LTBuy4HyVGaAhoFnwXB5XEd9zWcrBrCZ2eQEAl
mZUWg6qcz8ROnYLS6ShPPl/h5wiu/BRLqMLzKoJ7of/+0flDYaKX54lkToxw
CbnzR7+SQebXDIOPrTJiDgeCVE7NLbO1hky+XQRVx91kRPL7r6590HyvQpO0
MoYqsxCsdmZ4nkwoWsJzExlxMr7vzCa0RSPBBvkAVKL6npQANIij9hDXBDsk
Dm1ve3/eJD47DVWlwEdccgl1p5MMt6XGRBxKUgOFevA3UfvNlqeZdF3OeMRq
M395rLXSKsKMmkaYNvbyBYJIXucfBCeNfT6INLC3ymQl1JYekUp7uSJz9CPr
pL/Wta2WzSqy9v16Hja25HjLVSXF3yv01T7LeS6dL07BCiGxSEpC/TXxlXmN
RcPmUMGyiyUim4/HYfvFBlj8lQMdFN4fXCJ0mUmwL8y0HdfWwntuG3hp8lgd
yu8+b7h7+HHtVFNfBCGsvQ9TxeETuN92hjIuYoPYc/kZAN5CHt9ZnjnOsIq9
EFFcqcEAIBsnLlTfhztI2PFpiN3++wMPkabxjbhN9CCi/KzcEjKQr8MYc9Fk
cdCuMw9AqRtkA9L8un070cVAHfK9oBVlUornC3OTI5fntYRotqrSSb/24Lof
Zpv0fashyqjL34ayFoGxD+R2P92StqzyHf98T3DBAdtkynSVI7W6m57HD0Au
jxpi9uCQ198t+tsYsvsfMp48VNZE60Kxihp6wGl3Bc7uVit5jVS0u0ZO6B90
f33vzSRiM0eKJCAPMxZqg0r2JacvyLSlX2swnfuXTrgkzzmGqSRzPtPZMiSE
h+/JMWBY1RL1c2S1Gi9pmyZAag4FM3d1CMmfAHpNVpCSIlSJeLyCg3oNPEU8
YrmI8yNf599ACbKW3V6gpl4hgLoUdOkLm9jMPXIUrVF73e3KdWc1H8Ux3pKC
ujjgJwMjoSIEyjkY2R8A/7X7Z3zqTqxwxEd64B91zYrmglyhDR21lXDEriqX
pSQKN45ECnsJcEQ3OaiwfeifMLND3xNiLPurAYk1DC6wsS8+EVEUSjfaTj/l
wDZWex1TscC9+TTyasHnTL0nvoIliysM2VNfBkc73P4RsZ7rngrn/HOYUXjI
9v9Hx+mqH7Ds7m+tidurPE5X/D26F99oG5sF4uEgE06YHvAS94iKS6/Ls08N
9jll3vsfJZjvyUtIQk/heA85EdXEvDbYebvUF4ZJML3DGy/fv/OUD/EaurOT
fKzUkdT0ISx0+b8/X9ainXnO03SSPz+pX+kuivJIw3f98qzgyR6Lw3sgOeT5
SgN4wJEoNxO7ERAymsMFH7hTFntCk8kl4AS0izKAJtW5oYtgndOydEtLMHKO
8SFVzsLpk0q2JZHk8unvkPrEgdTfT+h/EXTNSkNOE7cg0fLzAF9tDaCetvvF
rCNdfafRYPVu2FlRPvQpFhwRWHoojxKpjCseukjdiM06GJ5If8kg1qj0tToo
Qz1i8q8adQbCPnbETYemAfJtCY6IWakZ8lcG1FihhDH37XKqszWBrWLiLouX
twgbKX9/NyH5MrYRbUYE2SacL6M+DYt4i4VgaYCObUmDJnNVFxIs92MuyAV9
hd9LGrv6TWn/HwVEwrp8yGeI7n9EqeJnoOvbpkcs2dg94/R0lv9e/PZcciFe
72aKbBx3PArAiHk3ftRkG7qkPP1BoBRzk72pbGspluEH7w17G2WJ5GlZqqrJ
jOB6APOSISoF8pDZMGiHrSmWD5fT+h+kn/2CNM6HGqqyWRdxYEpBvoaQ31x4
CyL+8FiITdksGHAnZ+7MVNP0KP2EM+WPB+HadMESIKPW0mHXozhTKe20PXQL
zSdQXHmrfjtlrZUn4kkArNtp+NN7srd7K5WAbUdRmQ0XSwUXl4g7NdltIcjY
dieSv4A0kquWfW3MdD+HQT+kNoCXTCOvNfOz5Ua5jWdYxI48kcZwgIzOI6Zk
5dYRYx5Q5WFCGgeZbiNpzor8HcvK7vDvqFxWCSa088eKBIU+q3Z+Dli6YraJ
THBYXr9tmwC3c5hvTq+U916QRoHgti0duhih6XnSqlQUIqNoltRt2acOhetw
RSPIwZ5LVW5kbQD8IgzcYbwVujjjpcdTIuZGftdE4GE4uomF+ifFfcPytXUb
voAurbGQxHiMO/1ZJzqRN8wB6r9qvBVkakpwCIOqxkWhuQz4rnkOOpvbRb+F
Hg7WnCOIY9w13X+IS7ZdpK3ZXklUqShf2o5pG9HgMOEmGng4P6CjPY4QJACk
lE6MxiWBV8g94SnDnUXKCGeqGfpkruf4OX0jk6Y65Mtkk/U/1XhAqx/wOhWR
6PoRxZXNEcGPfnvpaJdg3NyoQE+gRsBgK0sKqtUZEmrj+Flz7vX2O/xTpuc9
NEb15wOljxbh0IThSNkbN6T82Ul7INvL7QHZmX2KAnBmLR/Tcaqphb3d12+2
EBl4Agn6AbXE8HkhNfOFobgCtezjtpW4TeQuSmOdYGuFicIlTkpsDfmcHzhU
0dSE3MI1vdeC331YYx3qHmsPZ1MxunnEXy91apxhGoXu+5e0ub0kOVRAuTAv
s4LQmw340oSbWJeX+kMncMRSUkHUk66Ihi5PZzvPO3a/pU9sCUx9tu8Suw+a
gBvYapVYVY9Vtb1f1JeQuU/Mh1v5b8rRoJThX14hxA14IZy1dEOnpXUUjWO+
6StD9tdM4NWfpNxvtuyQyP/adqvBdW/tz/vKfwEmigah+jkzUMP3uPR1frM4
wKqrJpMmUuGd0nD3UEpIGu4u9yPR4LSM3AJBq9SWqIdVLQyRC/uVc6n6qeqo
/1HpXL7KpkxZY4xYj6I9tSzL+yuYpf6m3xfS9fpB7zqN7/q5B8M5n7cr8XIu
YYg+DDvKXCzA5OOsmDH2O5ZLeuTMslUc8bzpHXPUiyt8Wr3egFkwLC8KiIjT
Fy9j3xQcSAsQFs6guZALk1TUxfeRtSCJMkQWr8K7KPmTC6dDbYez9qLciHyE
VWbXbgrM2Vos202Us3U+wfiFa4wKFneYblkj8dHy3vyCaTyYWbHqfI+p4knx
Gg6QCKpJOEWeXyu9KklpYuWyMKtxupLaxw4DMttRuq7uetZ+/wrSPwycwfZl
XN5sGt0GYc0fFD+UnE1faFPUTZAUNFyNbC5Gu7BqXiSDAKhi1yVHDZ6Icyd9
sZMG1YvogDKAsuboA6HDMFPhaokrGErZ8nU4BW8nKY25Pee29DNW7xTZ/oFw
08czGUqWr+cbzjSWCQD/IMfQFG9DmS895jKhRuPr6xRy3uR4DfNejSlqptMD
yvfISSk+KTYWWLpX2Dizu6AnaC3FlVL6MEY4CzGGMC8WgHhVbGxut/9dzQPX
xSOvnDJCrzJNg+CkJgQWf/74LUzFvvxCVkH4TPKukshEagUadJNsrgv0/P45
HF206EokelbqYjJ818XcD79chXXNBxHsxsfb9QU31jEx7f/yX559VVvqiui9
1PMBAtxyk7inSDOYtqmtOJ8HHCMQG9SH9DMO9upL3BGkSBvJ3drlDZDmGgD1
0/+Fz3CXUxlJZKjvj5FqvoSt0ui8RVQXmyVFwKvhBCMyon9xa4TNBQZm5M7F
G55iNWjTrSj7aAVFe3DnER2FJ6OvwcYvrAUWUCUFR7+8HFxPTV2apIOA2Zbz
hccbSjPK3b7sdAWGdoDkZASjkPCV6HjQD31nJX4ZWj62SnlyofzT/PmruWzy
9cFW5E0iFs8EtZ6U0pdVBq1Ky6O5Em8nlDtLrtNslAGkSFXENdSRK8hWTPVr
7v08Xn4t2m5YMYugcSV5T+gjCdWFzccgfOfayoAika5ZadUXr8zLuxBC60bO
Twak1gN1ofk8fVCRQ7J/bPjDJg8Bmq07QXKKeYAwPmZp7rucr+9hEntLVv3i
z9XY65yFxrizNBoaJMle+N52gXYFMjo4q0ytXjOsYf+ieFeibJ5jbyoFjBhN
ougiTHhMMHJeZOS21lOHRPIK+dCRPD0GuikoTQZiRuKhxKA+Jtxe7/bWrJqw
CopVl8U59P58s7BJAbpl5Gr+CqPeOQIOFxAWiQbGoUmRNdX+LDK3i3rsi+IW
/S0kEbS998Y3FTdGNIHhiUGur5eqpy9N6+hoCfayMgmzKTeAvZVy9chH2N0H
PjAO/+jDzc8zEQyEq4a4v4lEIkjjuyV8svpFFhpvG6mvBJpi4AUfU8slGrv9
qxuTXZbAe8ER0ARjp4hrFTCQR/H7rxpmsYmyTUAIWxFMRxl+k/ByuQN93cAo
l8M54tPZcXVI7TYfIfOW09VEmwYi2Ndfdi7DwdiAnfGaj2m7omPftUyTVlNJ
p/kj3vKXUUesGRH1JDmWdzPQg6nYEN688OMHDXky7a5hF+Q0YFOg8WQayAUQ
QutCc1PFCDoqEadvBRlWT4wSaOJRIdezPvnuIKSrJYPCrAbq23FzqioiydpD
cwrhUuw5eMkuxBavA2uhStH77rU5IzhSqFz8EKFV9a719sXP4yRl5uBcIX3K
TKFLP5/Xd49tfrGDEbrsG4m0T40K7rcsL06cTB4Uw1ryIg7BTrx0N8MEqPV6
oQxc0n23yZgSI54jypF2hURHox7trpsMurxg87Ys7h2urSeyG2N36u9Hs3ia
GqCgCN1780GLAIr++cc5ezqtMjf8ik8Vtuv18VqrctnesQxXcfe2r0JnLE1A
D7xMYtecVjKA56l2E93r+CucIRjoq+fWmNJN6Duy3i5/69otWIJ7xj3ppr3C
UikjxomHj9JJtosBGE9tjHYnpn24CdoYjlTAUbXzEQvJ5KtMKhcRjz74WSq3
RVvrMXTcf9eQl6q1ym1b6T3nTN0x81wfxFOE4mHNxWAQlqRV+4emR1ywB6cS
u+QQZodFhmeItTV9jkfp25rg3fmiMCs6KHPxHXV4vBHYGxau3rO5/wEAZ18w
/qKmNtC155Eo5D1LSlw0H0apJ9gjvcTVb4RZhQ199NqQ2uujH4Z+GukQ8lZ3
LXfxIu/VJdpm2xynrmPcZTCBBM5gaPZoIwGQOn0sQoua1Nin1aNSFfn0AEL9
tZPye5V2775foEzQnPRNUS7U1hyID5xZMonpdYYN7qaP1Xo0zj/pQaOpgHbp
UWMcts2rqt9vdcThtwUHV5rMeU1DcW4P21GZSeL+Zb3LfcWHxSSmaQPxHGOg
xdFnkIkoWsArIaKlcQlwVxpiiDp1M7Rt+t572Qwa8vxRJmE2snjUY55M9vjL
ACmz+4fBBV4O2J1EFwZ1G5TbqRTmbjD6qIaftL4OJYb74T93uQXnVja1iTwG
6bJkTpLep3KS5Rjs91DZRsXFP5g4wdtz7XMiDcB/pGXOOcmuQfVy5ggfoIs8
EgpyO430/UPar8NJ8dGaLDRU8KmUXA3ll5wEehiqt6fI+tKCWGDgicT1qiVR
8dZnuwcfqWAAs6bufuWxaL7wQKuT4VJ2o0jjfi6obQ+fSbAyIG/WvRsNB2ah
wdbxukghs3D5KumoLfyd61yjvfZhQ0e3fXHn2SjwxYel83v+uTFcz00N9Khx
3ZIyo7VyYGN3kAM67Xj36eyJ1XSQn8kMzUWLcVKVTrCDIicmfjMXnSRWT+se
FFDXcXnynEfl66B1XDIyIVcMWcHcR2dxD65/ieHJAzN0jhY1wxEaT+K1vWRw
dmZJp+j4btR/BUiy0sldwK3TIV1RlsguDAaFIRmQ47AdSCnIroEiuHIVON1n
BzXGIOH+9+KXmKj1MysV5wZaZCIkbHVvsmMLCV1ma+nG+rHnAjQALGPeO/FI
e+rdi3ahr/qAxjizl5EwYneiL0DoHPHkOKGiqWsDQmt2M9r4eMRKqi9Y1f7S
iotX+nZJ992gUDegcSXTqrIbedGdHUFJq0GNgpCjLHi5B4cWtt50jwZMn0iE
TKEapsb4TwnXgHUNW7uCGYeVFA3efsAUHDvAPkZez5wb0lrFNQMEydvZlMY6
WkRO7K1yRS+oz0nozWg3aQE7OpRtcKXWtPlX3tbYZmfobDBoxY6y/JEYGzKa
084K+jAQTiQvTrrzVLOzEjMYtM+i9omrvMePxsTwN+mjnH6IUPz19AIdB0vN
l8oFENZUcFMSmuViCt4fFMg8Oq+O/QZbI1CQcUOGjRpHDCRaZwgI6AKban71
On7P8Xibl4e/FyjE7sLPVESdktcot40HQiQK5PFEXKG1tdEITYC24+X2GNOi
3Vr8RLkqvo1G8fNFrjo9UIvUaoDYKQMjqEqTGP2okToshcXliBw4TSHdjik3
HfmYvfxSdMDDnA6CXkNyBCD6GdEbkuxIF86DhJm0DsmSSPJIDPiGJQJtvR45
1+pbKfN7qXW5mWexP9Mne1FbZfVI2J71Zt1alOt8EKUlb3p3qXL0akvf8cvx
SGl3uJ2wTwXzjPNp69/TVIYmzIeZqtnxiU1akP+Cyaq/IvYYKAyLlXRaSPOe
HtFg9mW/EAwJHAdvs+DaV55IZfHforlZZx8UD2TsKTZc2t2iI0gxeaMFhhKs
5NB+Std5ishp73yqCk5wjA549eFhXDlarVeObrc9uh8Yf1UXkZxusWQ1uXs3
FE+c9LwDN1ACsYuYDshZ/DL7Z1VpY26H6E5wWk6fOzLSbuO3Fy0kh4Pb1CKl
+zdbmdAGrsvghMOZH5tcg8ctTTWh+28sb97F7eznTdusuzcutUK/hQNk/le2
PUVFC9QHQLOCu8mYWjD7OVzJTekL3v0kS682fRRR7rYwMbOaK9Ub346CweQq
2nv2hCKzI4OLXHVee1x0z9IqBRq7iNPHzYY6ky6sVUaogxH0aHM8zePVSJ2L
R1PVF+v1uOn+yFcHAtf46OhLLv/OQfHtk6l2fZK0W6RbeJgaLRI5yyaCEdT1
gFSP8AsvhKLh0B9IbcchFIBH2RH++iMqORwOTB9Lum8Cc/998Y56WEsbNK7u
uPs8+QlaF4uvUqNXg0oJU9zJStgk4lIwRLRvmqyM9KjMKAn1MonTrCF6cdKV
iDIJtvvBboZKBjOl6mkUe4I91HXWtDJ+kchhGxC3qlvHUmSjvAVv4HE95dUz
sULCtTQOuFuNpK7tSDVlgLXZ3lJzFiIT1MaPePVpjdJe17+lUIxlDCAmrCW6
DnDl2n+PsTrjnMPl+KEh7OY0BXVO1lQCTTyYB+NR80AOoisEK0VAGms6ByL3
JH/QDEmeZllIrBxtVslccNFXOIWyM9mX47TLEaeREcYvjseXwApbKUXFBKJ4
2fOAP0DdSd6iGBBbDjXg8UE48yJZ80LgjYDXj2NcOZz4q83JkTa7KmuaTQXb
iFPiQSlbP2Ca4jmSwSGVTh/K3gOEPJM4KjNDtIon/7lhFwNqORwd7PKr99ES
MYu6pM/Fl0N0IpETIj1nb/T/IB1KP/IcK3ODPbi3Bo5TPxLfY78xn1bxE4f9
AHtFNpTCBMLFumuWx+GXqoWSx/0Ldx2knTYXlIMKsSmCIwOxY4/8T1frDY6l
PvnJDLQLP6g+8jx/CK2J3oH0a89DD51wtVDY3abkfjnyT6DHvI8Kb8YNikLZ
WZJXUag2VMdMFoQwOZoVh5lu1dpoCuFLBaHnIUanGBsXOXqljYbvAw9KiZBg
7Myjr6AQnWqC/cZXT00G2qY8wBvXaN4t3dxZADYGe0lEZEBTP5rZyGKcuLVi
TurcFQIEp6lIhKfUM1iMRbtODAO3zrSROxiP4s++mEC0SLcEHj3lBJnXAMYl
CtZMr+YcKP5HnuHetBw0PfY9tVrqDb0+w54xJNw93FoldUD8qjCA4bmmKx1U
/uZRBeszPMKxZV7rpl/LFSLAlN7Kg/zvpJU13ecQKuoDDlKLsRfBAbw/CM0/
DqqpbHcAZ1qW6Y/mX32hf7EetmZxGR5MeS58PaMJ8v29d58kaugvXagXtEBC
DwkzEvASYExSFogb9ozC7l8OjKqv6Hooe2o1h9B8WGZsq8WNRh6j0StOImx5
LVDYV5eE45Hp87hXgDEoVmFVeTTpqDjWmWKSPoGzFv4HkSEFS0s7T7gqzQKw
FFCTv4BHAKpzncAUMUvvUawN6cttK/aZgMLw3X2DwB5HqkpuF7Rl8nzj9mCO
eRLpVpuWJtNml8RpVFXckopJPw0JroZEFf0Sw+7/Oa/HtaxKeGZRCKW4Bn3W
O9NmoA8U6qlqsV5j3RXHEAmqGKdRD7B6uSkeVUM7+7tDKfgTuc2sjpWeyd6v
pvcreMP9Rfun+muNl7XTvNOlueB7RktR/ZWIpyWIRdzElCSaw4792Yca4Lle
fC1M75Av0Lf3LUoY9FSVf3B4jHLgl8yO+rKw6VqoGRTWdDS+pHptnT4+rhYT
qJtaP1OP1HaHbm9EOmmmGfGY1Y9wvl+B+NY0lCsXTv6U96VEsLgz7MT9sMQR
yILca5F9jl8FPDQ/0EuPwv/xnya2+UqNw8MvDFYhyD9wiztlrgP6lBfOV8TX
RIEXi6Ly9oemDeKanJK/mNCDALX3MlJTi+KdeCoHC5E1F30DTI8KDCI8FXKS
VFh9JCx+UqyWe6V0eDFycFnq7dFMJbRa8XKk+2awubQWiLMu+0zf05VPr9gt
DwdTBd0tvlmv1nhivGxnpOyBaflFTBn7vSkt2R7UMK7o9EL62RWdJw3lHh5j
NIWvZfqa922mlhAruuRVk17divUTOSPe3VwwdmnY+9z1diVRwpAJ8bzWjG8l
GR5b77ZachnOq1yr6RmCZZXH2ahTEsaHGnq2dcQvv7OGvKTGPJbMCN8JiTZh
4JNPDpBQ/OjmIgZpQZTcjlgOcR3ynuKrwOQCg0+Kt2G/0R9zkg0zuBL6j32J
2kmaSc3AVNU/SJfS09qWC+bCTQ3ACeh1q2VodGdceFmPBNri2MEQ3s+ZiObM
BkNAsEPi6asZBbRS/h88iPJXNSaHjc6CqYNepD+nZCXXOeV2GRXsqXYmpB9u
mNOgdIxOGeUET3C+MGjEFxarwupVqWZLXzND0u8wD/mnye8i5Rxs9JiGQ2Ac
A21JtQArjEslT77/TaMXWORerH6ZcBE/HlxUfrEa4yIhy8ZJubnou4Fk5H1J
zUq/OXabJMpZ1xl8sJHo2i3tO6Nj0pFyoDvRMKTavjNEtMrimFavB2YKVni6
gIBV+oVVkYMHebdsELDlTgv0HQZ6p0QirqWi/W4XHyMIT6C/YTV+sRpPN8AR
BGxKrtYzkIJm12K/+BJujwhY7st9lrMl/rMHnou3ee/Hc5xmxLiFPLI7Hgrw
MH/+EgOOE8rw5Y0JeQJmBUHu8k7LfR6P7tZkByHfzTg5+wV/ilbEiqL/bWxG
bTmSWaHeFNpAQx92rfZjaTi7BpiO8FfKZR2Ocvy9T8uveDaSiYAKtmkoWs85
7DiEuDJsjf0Gi5YtQDj6932kRgPGl7MQhIb22jmex8ZmHM9nTOVsG6bIWd8D
hiJ8wx1vzVL+moG33QpzFmEll7yzTFKs58TMGu68WYCIgXuYMgSFbWzLrc0D
2rcK4vg0X9nWBqTs62veYR8QqUP0A+B5h4ctOaKQgACPEOCqvNkFJ/OB3SXM
FjJsvY6u4TMZANxwIX3r4SXhvw45fOWv6Rt44lnRoFgocaY0+8c+QOZBAadZ
dzbAJciTZf1DUBUmAoHhx02EF97pmRsyS8ArEpL6eHR5OJGB72z+ZhkAd7gh
cR127FWM8omgbgiqN/xUn0PeGEdjaSzm8GZ+eH9IA3eegx3jPpOskiIRyMC3
5cRVC8E7bUdJBg2qPWy0tVXbOny11N8Clo72SO+DAVgz1Egs1SbSEvEJZBBu
kMeLlgkmqkfRR62dORQjf6zGWkOMRhmzaeC/h9/xELB6fkQDGYoMTTeFO4zD
hEDAoNN0GJVaSQEW4VGNAAfxFTa54/vGdc6UWO8zAxLtbU9L8W6lOLi81HUI
g6hBBwrmYaX3JndB0G8VioxMlX4j04/fD0RBozCTjOBDNXJ+kD5/L7DRuuQr
jVkKnCW29kpyGYJxPtPYV6KEZ2/wsWk7Sk8nz5rPXPDR+C33YiV1M/xNrXHB
CWPSbsZUpU3D6EEn0lo177mdMLo3gxvRYj0GUH5H50oClkjD6O7etUkK3kAI
sAKIAuchiOBxmjgsP6iWbUcHcnuhEXqwuaMf7liLWVSirh1lrRepJznTedDv
t4gtpxYCKvfSDIFMPf1JakoJvLrtJyuVL2W5WsbSyOMUi8v0Afaxq3MI6iU3
aIszIjmyEFeJZlNI2KmA5oGyJIHdkpF+xKtg3hUo3vd53hOLz9k3neYwWPyv
DZZXPp8PhE4tkLoL+AAy9rvagOn62PIZPvFJcjnaxNvvaWoCTiAQEHsX6al6
MxmYiOLwthgY+ecl0qMSAl1g7AUSH6x+YE7wPJwLR2Qa/OT7ZLp0u2btB0JR
BTYH4kOyhducg7anWV58KQdKBaPI3xTI3iipgs0CLN8tI9ZmcKTQw0rcSRPb
vZ7jni07qOFKq6rhWy2OS0eBxjvt1U2ahN6iAjFeElimHSy7vSbhAKhoDbRN
VRBjhooNhHAlWKlSG36VsSJAJeCvuSzDOgk4zcJUlhwmTX5erKvbF/frYzVE
LLCt5ZzWEw5sAFHatjyKo+uNwZVEsjd+okMLDLu1ZDh5Sr6Stbnq6VHqyjb6
VxoDx8J6nhZAULqBf3oJi1fhhKZfLYNsi6+ryHvOBMv+aOiGcNdz3vLpSsWP
zDOSJNtvuuLByLoSzEIrqmUpRJsQPrMldgGc6j6V9amkyJ+hkhI1ZNrqocf0
IsIJtIo/OL1k38yvHcnVB/yy8KQH+IfJtmweh4OuZCZxBxBOjs96jtg+tbMH
cpLLWTvp7EJKlIj3WOPtvjdNZ06Kyjge850cMYyXFDb9YtfmCw+e7vDaSAM+
d51aB9FAv5Lz2z5wv60iJI3Qjpyg/XSMEn4S1EwwZaWsvBdSvLI4Pzud0Dl9
vcLFy0gbl/gxlTXIpdX/YOWhCqcAnalmahQ2xVvSdES3IaM5RyapKDSboonj
6pkHp75++43Y4vxorhbC9qW9b5NoVjL3ZjEdaSEgN9JyR3PnHQqktr5a0IV5
u3jFLxBtEzn+OLrKPk0LjZ7aIW5L+bI3hlWnNOtxwNBE4tYErgDs0KVgP7ls
gOMPCy6b0R3vKGO5NUG6pTGnVN9sldw6kBjNclrsFQGNK+5RzT9wG/L3zhW7
GTc0NEcMDmO9/AbHzb5SZNCnDBytgn7o+SoB/vklDe74wl1MSBW7gMya5jRF
7pP/Ni1BPqj5nacUfMwAucBL2l+dPiIjcvvHdWAlsAvcngqQvRLQQurCXJYY
GRWK054u1TQLY9oXKcOJWsUcAsziNaXbUJEMEj77FKRfE2B9ERpDJp60IUaR
yJB0rWwBKj4v/FYqEtVdpvAYrMWMXY8QdjnaVyRT0VP79QITNWNiII8YX4Oq
jV0uHG0PIhYzJM4JzaOETjS3YySgUYq9pUOOlgk4KMEY/paT6IQPthvDucGC
Zj8Djd/OED5VWWvf5l21PLL4Q9/9+B2bBRVwdFDbKVMFT1NXxxNRVarephnU
50LA7hHPejmKqWrvOC2RfGrNXsOlpGMfB34Ke6rfXwZQWJYz/ARgmQhf380R
1t/VA3+JwQpbEwFSSCLADRuq3BIo01l9Bt9G5iS4hH24RhIQo+I7K7sMCxbo
S+ym4Ry/hTUlWJUGwMNVtNp3gO15Ux3qUGT+gBk7a9UoyNElIKmXedwZRlFE
wZYX5xQJ4VMypXCfT/GpU7jHHQSBIos1xYMcHoSzKdO4v64va6NtNJHNowI4
poQ5DFQg8Kn9ShToAGsrXueaI8STGRvainQPQfI3lNhRBSLsHEQK8xZSWnmh
UEccX7vFFEqcgo1I0sacNajgVTbn16zZ2SOtf2kz0PtwVHizVZ+w9st+edB/
o/0ufz3C37m1h2WVU2IjXkMhPhw3n5yAXcdz7naqmeU/s/cPN2+mGFUaDjvX
gShW524jqsNwxjJRPm4qBWoalAC/FvENm62WuEUp6Lw5KejrGf6X85fAIY5+
II/3ZnZo3qmoDU9i2tGUbLzebqkwdeXQ0bNzvgtBhxXvbZftGNx2m7oWrjee
Ju9E/LV35AREWeDjPkXEgAXYJ/CEHW+cx0u/gAvInZZ4zsdhCdfeHVc20tdF
wtf/Yijmd0U+AdskEQyjHSyIjhVJDCDuYsWpWfkg2Zr9anlfBv4Z3g0c/zJm
7CFHk1CsJ8JANFYSPXSdqeLXCYXmSEIlaGGzhPN1au+9Ipn23GluWA27FUGG
sTK+Y2hXnHqEIrYqalXPQu4PHhOdqMubh/Y5Mr5OALfDE7iVKJLPlmxyT8xt
as8wY5ol1/wpXlV6QH5nSyMRMKAOSejF5KvXJhzvBuyKyqWp+U/jpuv6ZLva
mTttDKvzUlGceSMFGUzQMNX8yFRXduozyugamy+pOt3shQOKbTdFkSobO+eh
C66Ptb7H4F05VsFrh2uSLmthc5fEuuyZ60C45ynUO8Bt9qJ7LQJ4pjAoZUeN
sZBzyMbAFAHW8UCR02P/OO2H+rMRfuZnN2qGjfWsbxojMEeVkfsLYY/BCm8i
UrDPt5yolCCIxAFHc1bf+ZXuaB01NEq6bNLH4ddhc202oMulBRJUNnMFmxvN
bdfA1NuYyjRcJAVDmWVmAnrNZ64ps5yxybOfRDmkPdkdXgLBKbzopJFTsbBl
t5wvEB+ysfeOsZ+k3rewio/3UajjQj5Zvd43qN3BiPxn9ZfQd7SVmuN7LpR1
9R4z5uvuvmPb8tM2QBLG/XsapcDNHi2Wo0rHhva1uEMUeDdN9YzIc70BgtDE
uCtM9UiyGS/6BzWX22dx7/ZYueo+b2L+NedRPPCGrZwAFl4A1y9GnwF4dclM
52urZklkqm+FNBO2xOuk+J6ibHAWfZey6QerFK/qf/zAI69hCsNJazXsyvGk
LooYqKgrRNv+pN9SQYa3mo7xOSjdxBNwgDnPInW+YM2sbBIOsAxHb+xlJuGZ
D84Wji+umPVKFVoTkDDJ9eXKd8BewQYYV4JZLH1Q6+3UzREN1IVA3Djwn8aD
xZ67zWOhV2W15WfZk/n0M+BZQbbbLegv37R6nU+IzXiTQRc1JwOrSavfnaAs
0sn8ziZgc/QxT+cdK4Z95wXrZ9wpOinrwVozyG/GumgZJAuXIo3dKbxmAab6
eiyAztbY0uJbzkPdzc2rXBX27TU8pJsAuPLTsxY7HfXej24ZJwe0haOS4pYu
O3D2u26sOmW1XbzIvYHeBNaL9s7AQ8dJcMg5EJMHcXXH1r2uo1d3tDheqmPR
9n2i4LqqrIEYjLKH7qYA73E+82I7cBc6kdEDZCbJBNLaEkTJvyJ2D39mGqfg
Awh2JmgvRamM/Sjd2YA5XUuDHF/fOG/PQgEye52qtBI1tUmYHX1mOnQckJ9v
77nbKDYPQ3aBtokcIFDcTnxgu2X4nsIqXCFs55TSrfvB7ET92AwDMDVuWFVz
JVqkw58uZcaTGZGE2ar5NcXRxqYvMU1agOjxQViz18nTrzmkX3xcDoQkMsDx
fqHHm9nhuoRX0xmr55IZuoiBuYVK1zW5m4JZlraHS9ud+SY82478cxWJTCg2
K5zQ/oWGOhENAD+G0Y4wDB86F07Kry8/NWo7lcLSudvZJifocj/HaqD9rPIE
ljvhdt7JwyxL2/KvQGghLIgzXYlm+vNu2EIdqpnETFkzSUH2gPsM8htMYkUL
+zNSfSyi6Qoaeai/I6om4P17VhZLmr6/hvD3+/OVzW7YnjnE3wHz0IxqvMdi
rOk6uZq2tMp2e8Ze8j5rw5vwLwhNky7CzwO/5TuQODrKCoV003OyJ4vYk35t
mPeF8/d+7Uh5pCDEsIvFxQNMSAsOLNZ0Cr1r21W4vddDvZDqKXK91w9H2kQz
j+J0QDLnryb53HQMCqVSogCW+xgNGhQkyZ84Ww16YfDNnaSU/7RHcH4adWu2
wejf6v9lJC551/ZMVyaIxfhOpQmT8+7ZywVFzpyC6sHAND74UfCraFASRKvM
RkWz1Cn4ikAcMCnhbuCRFzfgekudoIKN+LTRtmPp7TPI+oABujQin1wmWGLQ
OYPdWruxta6NzQq4AQwWzdMJ29qiT0eYMbFKq78GT41ht14wH0prmkkHwtPR
Uu32x9Go8pPzQOuRRHsojK1eOxN7mcD9va/1Zfm7YhOnNf2jOwzy7X7yL9UV
H7qXAvw+fLYu4Tohg6/+nPZdy7Kkvvw4tVKpmkwCZI+HwWSoMNTBscXR0iKN
wc0nsHCu+NnjhVxOcj7nckfx897QmE6JHfFDZM1H+FnGHouVMkGXqThRfJeu
Lx+KgjVu0XqhHEBVQyKExLu3g/jZ2K7JcSq3JcE3IDcTn3gGvI4tQ6sQogRO
TUp5ZYAbNmqUawKihFGzH4JPFQO4UYW6yTBlfAvWi9Cxs6m23sh0q3E6HT0M
xYSjfjVtZeJDTAA0gzgX9T9Hg+90yOZWvoeQ52CsY5zsD+rPQQkfmKAiXxAq
YuMVCTeqAL0H9nbctsTtrfW3EaJr5/xCXiRJRn4Qf+myEN6LZ2L+f+Ikt8mv
yX5J6VcqA7KUbcHJy8SMlGmb16gVbOM8fzZSZfppYDZclp8xaTMMhuUNjHLd
4q540N7h6cvzHS0rMrXxfebV7q0Iiu7XKWGFWL1Vgz/ZFeD5y+MHVWWZKi76
Oyvo4euJrIHS2C18pvS13YUBssovgiGyAPnVNsjtHYXjbGnQrK6Nw2/5tQm5
VEpujMEOa7HK+GNeIvQzdBiXG7bVBlKPbcCVASAN7f0+Au5Elm6Sm6/2kvxH
fa2N2qqtLCvH3fvqAgUFovbObwZdKmCyZ2PJyyEDQEcABiXNvhaEFDXA6i7u
rKXjRdZ2EuRvCbLB6H4v43N7GeGA0vx7nIaQMoL5x8cD+5SbRBTycdKsZKS5
nPbY9JWy+J4mzHra1R9yuDiqp7H3wKCP4ikZewGtf69V3b7mvx6aJtqq6x6j
eWVzhaN/Kg7ppwgpq25gRPvZdfP0Ei/YHDa3qYL1YADx7hIVBnluGSE9zUKO
Z0ncWWDT4Q/nYr+B+qiN/72kXfYkcSgR1nUWN2+k6hE0bnAL0AvIqXLucqoM
MD63jNJc1G8ZtdwkDYdc4jgv+ReJ9X3vBI3PHdK0pK/2RoYW89t3QD6SfZwK
lPWxIL38+G1OuBVyMMHezX7QOnJhmbBFY2gmmMTLcWgrWNA6/o4WAcaPkVXf
tIkugpl9+gtNoaJZZyVqzgxziwXDKWDt790biw2NNhrsbnSH7ngEu1TpFcp9
V1jk4JU4DUFpJMauA+fcPHNSdYapyGiXGZqrrS+Ef8YYP0WdkKtJZplARRFg
MsuiRNTLww65Lc1qSysd9mGQcamV0bt7Y1kgJJHLS3lQcKsJsFFhYwNMu3cX
zBgtwCnIHA/TCj81UyeWJQ9Nn0JKDYi0P/MxE9hbrlNbaxrz8IpT9E6tldFY
eXK9s1001F5+e0j48v3eh1Arya40oQ7g7LzKWZZTCoqjFBfjIae0OIDYyFGo
Bu0yO/2jA8S+RwiybLeqz3UEEn0qNyPMIs6tDR6b5GcJJPj0J0mkji1gbbPd
3emjXISyyyi4SntXClnow9ufgjGOUc0Pv6T4pn1jCeTPRJU7xGFkUQL+BshW
Y5vNTSCdGTPjjoW7/xj1Xu5qkUYrLYA9B+GvyyEjcjCdMuOmu3Rf0fihY0cW
73V+FlfQx5EaPFsijtd4AQdbOKIMlAhh9QuUeWS6BwpCF6/ncvqej88fN11C
4Rt3IirM5D8nL4LH6NptKA5BN0qI6uDEHrsWUyBF7m1vAYRYMv5Hmtd750XW
uA8PkzaCdZiN03Sm84EHTcC3wfh5d1nNyGm49EgabzzAXSnYKcwnc6zz4mbu
B5qzTD+NKR7T1Fko5iqYiCRwR779JpS154KTYpllbEdPIooAe1XC41kBq6Hs
q9ZrDBm8L+zwEuql2hfjGxspZ7Z3legbyhRbiMfQ7pjcnwahPS6O+SlBNg28
cBkM72zgP5HeMLyglC2R7k/kgvctGZyiHa0fKlGvs4S+a0jmBnQa/upnKNem
TYdwqkw5CBbqgnboptKpRlyc9AhRytSyomiahWxgTakip3dATrtXqDP8S62N
WBL0oWO+9yNFdCEfrA3IA2puS3bzXrGofF9L3f7L6uGZQCw100g8yXUXKFMN
L8zc1oX3EDm7bW8fF8XgWWbJ93oqXlbRYJUIwsM0LEgu2EdtgLzhXLdEYReG
JAc51+x6udR4oyf2ntJsjkYN8BPPdEGrDucKvbTJwKcGh/VMLMevt7F4RuBJ
sTknRSGInkMW/oiBx0RQsv0aserp9VBsJosL/IE7ozNJQTBFBGAZJ6RVq5lY
7SqrOe98SNqPJA8+IT3oPMVa9h+bhOvHP8/vf0vhs7Jydb2iPq/43oQKtVo4
pc8TN7x84Yj6eQspZf/TLsWHCIFt0yRByJiMw2JCXpWQibes2rRKO5fL/015
JIzEeyye3oRrqaCFQTKQtlh+NPxsPhgfmkilPkk+XnFs2wDIN49i81YN9Z3O
aSuk2RVOIxWtjthjZrDyI3H2vxd9NvKURfpfcrCf9e5rFeCCx5QoAUOZ98Sx
EY/KTz/Unwlf7QfVh3epjgvT6aGDNis4x+gPVABDGhVATFw16C4yrhbweYnW
rM5i5bs4agxecU0vTYdtMv5dtvSzHuCxUo9bl7ATV/xc1GkhP5DaFIrL+tmo
6/9CGIQhAoM4H6S6DuyJ0rnECDofIW2FnlxMaCh+YdyU7zDzIqRAKSjWMPWb
ac6bHQpXG5P7WjJwkdyL41wvacEVhLRNpikgo+IFdSpvur5BFe49Am/qjPrB
4NWARkBh0hRXGBPdBfpTOfEGRaGzRiifuqazxOD5+ov24suboPmTFaPTtvvw
75aBa/FutJaWMk9JLfTnsGU8uF2ofivJFCL5PxHjB8DadR1kFKjOWv22z/IM
X8knYV14qkf4ogG+tL0yCHD+4OR4XuWRAfsDOx0nHZOLin+aWVWRE8ZpGQ3r
NlXSCNKlu+Fi5EtMuDSOt58Bnn5oNEfBGM1h+Rybgmkdzy3nE72+1ZzuUhwq
L5F/30ezgTiOG8UWXMZ9l5HCPbpEGJoyOo4ntm1FiVT19rdSaTwD8udoHRLU
onMpMq9p70wUXlGuNDuo3LUONEPQIwAjXk1v1HpkiVGo+RhjOnPT2swDOW9m
T8EPVbL7umw/I10WroS1+bmVsdBuBHvf1aVaJJTjVmiBGZzLR1+t1RUX6r+H
4TK9KHOce8N47hs353Bh04savIqrHJymtj5876ESTg7qxO1FrU7Kh6VQsCFN
Y4hgfvkS+g36luazg0zo5AWMUGq0uLbHZ9o592cknw50s6+ccQ1A4uco7+gv
bL1bmBdF+5RpzlZkMRxYX94XyMqIv8kGKvt0ccvA2zRQ7p/YdgOp1nq+82XV
bhe4GUw4QriwwasyiV4d6I6PzlQrjalrQBZvmbo8tRrcNm1ySoPVynZuOeCP
+5PwqCnyJlsccFj1PM8ZULZyOILQvJ1GZwZIprrJYjMGaE4SU7VAIXNYLCuT
MC/gHzHjn4bAc+5TKOxTcm+rHLJAq5QA2Mn6oKRvtPWCcFkQGFLJNVGiqwpN
nexHFSnz8zSS/ms1Wauooq8b2hwOmx3m9F5X8NgDoPQSdvA/vIZAEUWjqo2K
t/h96S/RxeHVq1q25yAzDK4ZYgmhtLfqtUgox24qLdwbTTlNyP9/nDaUezJ2
977S0vinVjxWCQr6IV5qLQf7zmjzvujKXuPBpGPasUusmT60uns4DkwTxd6U
b7P/1Di64fQIGNAjDe8MfiLM8adlMSgnQzr1l0Abzcb+b7ppRZd4YmHB8iw5
XdpbxTwo0XT3L8KukuF36n9rAXrQV5rQUgO5RMsZvBSXKij+DMyYzt5kiShZ
aZ5PWCAgluEpo54FKdKrvyDwAFjof4ZOnAtyCOXEfmgn3Kn5xmgRztEPhvwG
OQj0t4yPVxxJ4G3JQY3X+sciesyshZS3jAHEfc+ptVwBTtazOYPAuvrDEQFB
e7MmcdE63zEHVGE5mjYiUd0bmy8D+0G2L9UKvxbkySZcd2M1PdKVz+GSXcqK
w7Ys6oBtlJ/af7pDpqT9g74T2mXdCjLfC3+a7Plqe3CoKo55J4Cq/5pSES9M
tE4mDlD7jc2HGwHpu9rR6p9pCMmI+lt3f31Q2D/8C44SQlD/OpvbnK0QWlc6
K/DyFh6MTcMu9A7G3FDyqfC+kF1zrRuAX4Ai4RWV5avX4vqSsLmvEbX4+8vd
afhGQZGwlpUXpw0Dhqk2PSxyTuNhHkeICrZPuHJzSVcDgH9YxjS21GnpKBmc
8mdycuB9kK84et1qhypaBGv/HL+nLvM6P7wR32evy/o/wpTTKGC+6i+WNlAs
7o0jU8QlrY3MiOuLtmK+VU9K8sQA+3Iyc4jjO2hV82VeK3FOgZofDJHmGVzc
GV90Canwq5+UMIkHeG+CpXioS0NnKcytIUhXNpNyi9IAAYYonMM65x4778PN
dM8jwT1oqnvmndFxp6LNqBKJgHaAJpqx2w6gPk506gvTAmjI2X3C4AcR/4fB
YdA2nFNQtDc0PxTtU5Z+iTVcq6TEyNP90SkPSv8uZJ4+QlVJO5qygSTKag4m
3yB7CH5OHK0TB6zxDz70Z6foUpI08tlr1+Fzs63Gj3ATPC/59uSlGc19Cm4F
u8nJdXzybzlTwDTi9GEDPzyIfiZ6DZaAL+Fo/m5cwdl0FbqclGKR5q9T9jJg
8+mtYbyvmZEph5GmTZUFFIddp7c2TaXtLyv7uNbiymN2xYhHN064WYq33jDH
yPZQ6KKSI5t7LAi5Fgw7i2/ogAHtP1BiGUerAp8cbKJxC1Rj+rnI0ilch/5p
N30+lb8dfnx/YmIE042XguzUwpRuMYj0zTlvgTyexPs63T3jq8PRzAPe2qqS
9zFPxhpArsKuG63QUVtP/qxyLzVP1THpDfONlygXc47Omgm8XPsRWYGrHNXU
EI0AY/yvvTsYJsvRNaxRq/b2FJ/4s+RHld4NccjPCNScUCSlKkziX3t2eikm
CloKrD2SUY5VZOYhAxTjSBEJWaTCOqEEZHntQan02He+sSvVBFIvf4NwvSPn
nrvbrAMpAmjwNXBqk0FEW1rgk92vv2mpJvlUuFo+UgantANeXHXl5y2m0wws
T+UjJVQeEFS6Xzw64MPHkV51uKNw8WxZ7DhIONItiN5NtPFfgW3lcW5rrZ1G
4sQ3CRXr4tVwGQo3RZPxLBO6IOrtNfR4R4wsQVzCvDop+M46UnEURh75O6UR
qRrzD0i7a3ZTSaadAtj0jGOV9C2Dtg/M0sv6B3RHvo+T0kWmahASlaChfTPk
EHyvq2jfp+33rwpN0+Hi9rAuMjbWOyOe1AIZmPfYGNdBOLQMYYMrETncCCO5
hiWT9HrmfWE5kqyH5flLsPNaYyhwNOJ7VD4Hw6sxq3NazWXjJIasYAATnuUf
9n3pnzNZM9AnArUkVbezpbkYLwjUodVIDB0ZrlI+6m5OHhI1IxcsuTLqMOo0
UTmsq3mcal8BvULxo8qAxP1SDgGiSRex4HnDb8Q72yDmADfdpMrYoN0mYC/5
srVHXU4NRIExg/M7Px+VLP8Yz78ma+KzTgKHPP3sudu/r6/u45ccLeh4CiTK
8WblUwS1w8kfx6pRh6wAvxMH8qxbVc+kn1Q0NUoa4nGTcm5tSkxjWNf9TYWy
0DtzEmDuyvvjA4T304pSq8f4/2785suvHsXYEFO/99FJ4NB0g6pyLxeOLgXP
YLAF4I+THSYOveNkQhJaX6f8v4wmOux4bwKbjbHRl/IPrbIduCgDiA7tvbJL
RduZzsMJc2wkTG6smodLt0UZT2OgQjezPINwCOAdbhQOpiqvlcvC58qMa2ug
ZYD1qUu3SGtp4XMe7MlJ6mNAzHbTOXbJexRtyYUuQPT+lj6FrkQOaNhS2CSd
ZyXHDHXSQPYruhsQhNr6/WkYQZ5JotmKE0QqscrJQ5mKtl/9uM8xBtn64ZD6
fY9MC/4Bg0/eHYmM/lvLek2Tq6fBMNXrIxgcPOuNVc1wPAyu6ITFPVAA0Xvs
bYZfg40tCTwx3yec5BP8OXCyubLytiI5dbhfg19BIUZL8rAaVeeuvfOLmvO4
XKkLCZOnpcpfWKn4VlDSsQPWKSs1A+JEnBzMsIvyAifp4rBakbS46SeqWJ4d
o8NDUsnmbxM4lqKDGrx5EGU+qfoKb4jSBRqSQgf8QKJChaSTNcUmgte8DEQ1
cIdLMftIB4mnFXrCut38nVRjbGCxPvPMJ3G3Bm83kOG5heTb7iXU7Sh6b/Iw
wclnxNY9vdzFZk9RcGERKZOiyMmA+OG0rlzcbgjx5OsCrLN+yZPGgMzS4pr3
LIivyvTB9PKXDztgHsxda0WPNr3yf0LGZsDmItfhikNTUTGCfRhSoaiCuGCy
SaLOxNmH2T4meIXYoHHbUGxPnI6owgETWN1FoZy3jyMSO+kZxBJHl+1WNlN0
gEMVwa1jbj7P3Mbt6abbrYFQJmr2eLVWJs4/7OlHw16e6BgZlDG/c1xd7/9d
jLNyOP4zS/jIy50FFI+TUSruXwuR2rjPq58Uaq5G+c5eT6Xg4DgyaHT4XA9H
f31lLYxXxBx2e+D/KeWw8s0qZ52rOFAyW3ChSpsMK5WExzMMxvkTbSJT7jQB
LP7/m6x8qP+0u7O8lfYDQGojIJJ2tlzvkrIYeA/uJ4ncVEY+7CEOF2aW2qZG
oWH1S7reIEOGh/NoEh62f7KIGZAvSIfmRDu1ry87UWgP7lkGW8GzmEFYdZOR
bBJy6pl8fB96CVVVZa7K8euerTM337WW29SQX09wtxjC7oUa5MeLCJsCsD2B
umV8kH1puv6K3fP55XSTFjeDl9YvJZQgzXpyYQnZNZZzABeoxDykc/DHCF0w
Tp7W2n8HympFEKviAatm36ZXP+fGlenb4sPlBnq0Jtd+aEyirOR0/xLwX4r2
hqrEz6YnDvF5oj4piT8EnF471YpB9uU9ekQpjA0hzk5GIXLnGrctguzPKRC8
FsE+s+1RalbmWXmnHeEpijhwt2xFXxp9vnCMmA9o+8RmYA4eZezLosgUrwbp
XFdY3A4LF39KkrfHeHRJ6gaPExy4zWvFWE0jbIdgJQ59WOag7mUjomqvEe+A
/h6y53F2XCMQE/F8ETNX63XT5F0wXcQ63ATRjXVqHQVnLgFJtNqT9oNvu+Ug
C4VUDIMksUcQkaAJeFcmz/wOzUg/zBzx+JVwupTZ3UOT9QbDL4eEx4wiMjPy
PskT2Y4qN4B02HajE6FkCzclp83Lso1nAwhenGCd6/ubhoJFbjeSeygLAsDk
wpdExD2ZxYmDvY+H6PilL3DEfJ9nr1h46z/v+JN6Ye9KK0tzpjbzlPXFP6F2
Ug5T8KZkKh50Bxm/dClUyVCrhYQEvMpzVEdnZP6/vLRKwE0IAmOq8ECwCWNM
WrG3Yn6srROWkHSpImHblNKbRqF13ucCxpvwgiM5f3IAtN4RZaTR1+9hWEu4
WiZyXmKqlqTB269jnAObzSQ63fLcjXMOSTPV2xpwHw9ZSalbt/2SiAO/oJJX
TGD18r2wSLRYbilj6NrqGMcwO3KnNhR7xxJpSvuKQJFq8876t54lXJhwnn29
Teg1IMYzqNXdpQ47LX3k17ann3fKksLUj3Cp+NNmK59LqsjPwyBwA1yPyk2L
D66yvhxmGxxqRNfQUsyYug3OsnBO5A4MbS9JjogT9BrIismOTP3X1yG56NSF
x7SKJLYaiOJUqaaqoYA7PrebrXJtUBMqIuowb/0bpi+xgic5W4tmZ959lxPU
S5MZzgUndCoaJcVfNx5C91wdxMYogHUGrF9CGBpoLSdw6UvP8z+R43VhC0gQ
ujtMgEItduyeKWd3YGYLRH/QFEgVYYMpoJPEDD+9p5yDd3ZdXq6oDFOgiYLO
mgDcYQ/EVGw7a4Vn7sdLFjG/ebDh6GGigOqEnhLXclAbhft8OP6d3faVgmrP
Ycm1nlzfaQMCdhFHkyfJLId1VykFe27ZpLfwlttwZTVNr2D5i3M9MD9gK/oQ
a4TlcmVSKEWM10FYn1JbnJvYyxiAeyjuqztyIT9+wemiH1YVpuWKBmN7KYN6
EEKTgRdb2EX2/A/HrNoTc2thGRr2Ez0Vi0qNJHMpPiQ6qd0aJ0kenS+6TTe6
9hznBRoamjTP6vZ4yxSDXwJsCb4k4/xXSsWfNn4NteEoXGrsTu0QXEplyARi
BDgO9qZE6Vus6Oj0GvXD6fdDjD7UzQmX7Tkc2F1qkayasiVNQb3aclYbIk+e
zhxeH4yEkf2jROcYfiE60NbokdkdYsXzkYY4ryBBwwjgV0r4JzG9pLyj77M5
4ser+jejlK/pnFlknY5/dCup+soXp4QQhBmjwIHIOMdw5JDsVOJPMkfEC7nR
u7pp0Umg2MmccL+8satS4TZtEa/1iZVKBnfGlL4RFDSW+wo+2xglv8wYN2XA
5JIeQIE+edAcQH1+NqbLpuVSkAf4twnOZG09PlMbtoG6VHZED2YI/kpr4eX4
q6gwJ+Ov7uJyYK/m8KHCyCEv/PvhhVl0GoxGGJWVtfVcnmORNkdXCT5oH7S/
BfQrI264k3v4TgQyExTY/n49FQj5T5BedTs9wA2Ci7plrtSDRxu1h8ohxT7P
4igauTqSuy8lB+qOzUqvoQSC7oR8erpS8tiXfmVhLZAT6186CJj6Wc1afM3Y
rL2FwL3XYBslhWRLVlN8SaDMkvVznfS1TNqp3DVzbc00KkIGcx76DOKbgmYc
OijckaTU0YNh/Ko+CjcnB8+FL9iIgFSpONcCsp03zr7HYRYB8ymxvsXhE++F
UHp5hiWjTeBmTexEsJ4QfB/GR1BwmpAMCb7FelYIQMB9AMILRTLjAacD7rju
ITSlPtmRTpSDGPf31yTrzO5PzytQ4KF3RMD09UpSaClFRDHaOeKX8YPU6Jfx
4IRyX4HT6fgkS3pBCBs2iAZ4iZqKZfi3u/svoyI0x7Cq4UHVJhljldJG4lQb
NqK6376FL47/gboH5qxLTuR/9Ct4STYMDvo4GawUyAZJHewf0rilHEmsvD6A
Kf8d+RpqYZeHObToOUdK8N/bUU4J+XV1B7aw2CoWE9xa11hBAHAHEricRmdM
Zv3DNSe99AWH/qOdeVg2YJtKlmPBdLzmz49Ph56DozxU2IUMBroyd8RiZnUY
OWXuNeVHXB8HIGMXSWq4dGRB3fBpli6OCk/IkxhbXqW+n4LV3QSzGho8G1F0
weezOvFnUL2ISnJp7w6mRNwAgKFMKvMv9gCEpJ4Jf+pQLk7G6dSC155jgF47
LujfBBQTdP2sanOmgVXqCG4zbFr1xUIz/9s0z1mfuEQmR448Go6JVUEGnIZl
GzQ4bJdXdDotYHjfzVaizWkqPQR1MEy8DtO5e6F5YLXgFBk8QnH/KbtSnnni
nsL9/e0oN4wa7vHyTCbPMvU0PojECpr22M+Qmw0Gf5hTMeTqqt6jgjpQTpNr
xjqU/rOqeqprYi7XSSEn+lUwRqdHGCu4JqcNDGltmSgK0ylBSgVbmNJgOX59
M1CxBZsh74hnH6WXzaaqIbrcq5Ilh251e+gMKKKAml3j6De8tIRmG7MOpuvS
yZ8gOcyCt+x2RxUUsX/m9FB0XG+WgAYVZbFteNdO0/ltSeX8RZAu0wpLhwwk
+5FuDAOwMVkqENJp8Tcga7S5ZaFmgdFSdc3fxH9KxP2zHd05oJ/F3rv9X1xK
uZMUTA8Stt3qddmAxFEKXmOrjKS1gUuDI48PwmCftOAZpREqL1pgeqJnbftZ
T1fCDxmtrOc/Pa7adOlUMtEFbV1cgeq0qFthIcqaDXp4tILI7PZxlOIQ4k4n
UgDH6EXuGKhJpersQrIduPt6Sw8nfbjQtWOryiMXBmLpd7YL4NBCfm/P086X
qg7uI53Fq9aDOnIURDIvx+lxBMbpHnJVfK0fYGfu62seyRfv3HeT7AKJVCRr
pq5JunTKHH/OzG1iIWwKcJtzTMymfxxtTRi3fCj6jOFLQXdTAdTjhzg+sBUe
KZkp4doDH2/qfTi99lY2s8FZWr5K3WzHd3nlXXLqYPstquK9NAFg6ojz5c0U
UxtG0w/ffy57EyllJS/yJWSBCAo009lW7BzYzmI4cjV8xZVUdKIGcybVhDDi
qxhrIxvHrUNFi7qgCEOt12me/hpSh7bmrU8C7WRre/bM7q4AXZRDIARiymZX
b8afJiZHTQPgb+zU7Ta4CGSymaTmkbBZ3SsM2R8SMZtx42gdS+eCCG0fwYcz
LVR5L8kVkhDpODET2Wd/z3lUToHHb7h7lRZSjVNOCu/SvYCZoqyDEEHJO6pL
IDQu2JyQe2nyDYdFyjo69kvyFZmBY/iWy5vf8TcNIKXeIDqXRC2D1Ss+QArd
6g5OAFqrlKLiAAxsNRh9WKHpYmkbKKg/OYwC/wqsRLWCVCI+dyfp2TgklzSK
oUylivhRCgUyDfiNDfy2PcQdHVR0zndNoDIMH905b1WZPGOrDcp0iKALP4ca
oEVDTMDNG6nJKpBC76WLnYNCJ1O47Sm8Tb5Uu6Xvg2bkDiVzCIAs/gAqknKS
HF3FyK7bX3GWwY1mweXj7YOblWCuJt58wtkn8OSySxXuF3urg3AU1ObPxAMl
Mz38PwVS6FisPhGYmrz5tcWCy9JqJ5dofHKjxjcGxbPwfdIvQjHj66HYLys6
cbguVF2dVPM186Erg4TQjZHTcOnHFshsK0mKGNs6Pp9Q1ECWmfD8+o3vtOo8
Jl/eTMMN1S6ZW+bMNc0TQtZOYjQlWIkVgqhEo5lKzA6J093GrX8GXhI1fgH2
j3SzppRxoQw2j536QIbGWvAV826j18uC3NQLKAmMdscHT+sqzctkP3TDJYhx
QVXej5ly/5og5pWWngtICgtOyo2Qqz8lCdBRcuo/1Pk5LbRweREQrPRwJg1F
DhrZK1Kv7mX//CvJbvrClYMjnAHEdhMYVIAWDhF/bJ9cyBlNKV5bzk1LP4A/
Veg7gnGF5bPiD6GFr6+shBNjngHmaJJypKfh1ihIvRIPUtzIfn8kK04lyCHy
qqSHIzxQOPxB3jrCQaHtpSG5zQxke7hoQpjqZLInGONCZEnwunjRVk9ErcUc
qGZ658/Kk7Meai0iztSyKBKwJf01HEEgpoddsqInkbdL5oPhHiuuG9gILkzN
VO7m6N2yOB0MSHj/mQHnoFFSm2/NGP3teasly1fVj+ztZzJg9/9xz30Bw785
rkuYE/lyJbrleEiPRD03W38V5e5HngloSvTuwjEBmnCwjhUOJiHMdYgO4WtO
ajSVA9zyV9lfvsgxMIje2d0PapZ02cnXiIG8VBc2M9bISMCo/ul4iduPHFv6
G2XZIWtyyB8iWsIDq47/URR5Of6s/kCfU8Yrl2c00dy978sXQ87ASHWS4SWl
E1qQ3sw6+ryJJ9+EuTP7sUNresT183uoRMXnS9ZjvYAz5G3SVNdqC58HqLOq
90pjFzZfE4Br1FcB1wpqa9bP+sVTbcnZk3SdcxGMFG90ITz46SM3jvOuD2rt
vOBFYBEbJAa0BEeq8vRbgQSdayih2Oh7V6NWRsD+w8dA7TIJ/9bKTaj46XVv
YEop4M69e5QMGpfnEkVTZDRZvVkso2gfo2P9H2NC568L62t0GbM/Agv4hndE
qi5bsHwnaYjMmbc/n7NLQiEGfKDw/63Pik9g84y8N0Uwz3xp8Eug0OVOOmhU
PD9qWxTgUYeMVh/WdhfkhEhC6q/JlkAC13oD0QJ4XppGIhLs0TkxtyjrqEfX
oG6FdwLUhgN0pNbbmUPAndYQ8KsEsnI4hpj3+b62FB30ygUPElq4l3mbUNl7
o+PhLVLHINu2R8oSnX6QyvhHGqU1vqA0J4vymlowwOtWNDOBnCcac14gjgMV
iUVfnajDaSP9nVeSL0wewtpJnfgY+F2P1DFmpfCDfW68OmLtOMCgzi1bogaU
6Q30E4A33CyxmJmQLh05OKT+ida8cZ6V/PtoTFWk8IxlYVAjNS5dF5x2hHC4
uMR0MMVmeEdGzBEutr79luHcg6crX4G/CeZ/7rJFFwshm5NfLhLkhyx0Ws6s
+6skRcl3qwTdE2feri4pUXMztqZ65yX8b1hpT2RhoA0f57Rg/naMMooCza2f
bK+eUSg7XCzq58GR+FGm/QygAXma20JOKx7ahq444u2NXSfAgM6L/DWBKnyg
h0zsQfDLm4u2DmJxg6VDMVl++4+FXETwCHMbPOUIEWHrMPi2OtfjYifCYoON
+NmYL4CNddAMJypp2Pkhno1fT0YvScWYl3gYGTvAeST9U05Kqu1AiGwlha+k
cYGbJ6pDHmky/9y7+gGXbC8CNrIYxdK/TDPqmCli2n098XutGwIjtpUuc2q7
uzHgOUYx9T3bZYjdMPVdvFMqdi7wMf7DNGjGTNPUlU5DC8tBqxbGJ7/kZ+Zg
Rf9enAwOO18GSj6+5w9iQTQs3HfAUPIWLTxt8+Jqs6orWwQFnknZddRqtZi3
Xwz8jv5VBUc4PAFIUIxvCSNYAWwPi3N9eHycPsfWCz7/exo42xMS13WU+En8
y3ncrizj0yMe4vgg/JOgYn3iDx0TD33ugjRXhac65QStO0enNSoKC1jn2+wd
KTz6NUfhJBI3o/lAZ99AePMbrvkxEJBKBhU5+vc/p5wI0Ov29vwHRhbm5Ih1
SBa9a+KeUmNFJsiY5BzFyFH3KMNL9I0UA8xBXrg+MusDU0MZsigDCguqx2h8
A81+eQUDA1IVmj9zt/Fyl1qNjZZe1x89NWIWDAeZoqdA3bUW5nv18ixmfMOr
rVhvH+pSQP4k97c6LlP26aB1oJwnRVT3/T4y+bTiT3HtCS4MhGld2uQLIWWj
e5tmc+O/49Up5LhTi6uGK4k5FASbdeMuQBnxOYan6KQYzmuT9fgv++7+9X2j
Q5oRQItjWV9HPTdTh//qtRhfJHWSCXUvd8tMRa8oQybduzPdvbKcdBrGK42B
GZUaOcXi1SsyNfXGFKykhGqNVeCy2kxqsm0mQ/8Rh8CIRcU0KyWooP6MlVI/
GPvNbXmGOCHCXDR3Qcw4XM9/wsODj4/CjHGlbnTC+OBJutpd9JPPz+3OhiM3
sVXABlBLR1q3gNxTU0nAvUPYm4swau3XwcI9MV269BT773rW6zwWCWbXuc1j
/NlaaMuwg5OOxOzDgGVoTlAXZp5u1CngnVOLPG2PnwII3jztXqa8LXtLO0j1
cCCZMMZWD//fuNHsB+5sVohsge05yVvEoH6hk0S76iQm3QU8ZVDZAFBwLmf6
xobTTlyzIGKt5kV/c5Yvz1kN4iuKKY2JwaWVXJNEU4Td6EQ80v5/1YAhiIsp
9ES6KXDD4uk45UmcbWMP4+eZTYZg71hkG8nVP4Cwvj8dAJ6TZk83k/ZxzpXX
m3JZURCbdb0uqFccJ4Wg07r14DeD+1Fx77qFCTtRmp84dtNMZjaSOSAsoSWq
hwjK50aZNcs2G8xVAi0BcNNo8Mkb9Gmc8n4nz04s0QPAXj2GlWobx7GGfrS7
05ieCWZzsRntd0amxRA349pLErKArA8YaeHmtbc6opDep+MK+GoIez91Nipd
b0f5Gkdf93rphBGsgv+/xD37idyYxF1s4mhLicdJgWqSjYQRObKzDS+Kfhf3
wGVvVAiT/r42wXmoeXR1jt9LmSaNY7aHsFZifQBVfBo8MSoW1RS0GXFikQwM
SmTiW2ik9hJoCxOAmL37wzs3QlUCRXPE5SOhCVMe3PyPAa5KV6KC9ZFA9uDq
21G6GNGqSmltppsBGu+L+y065Twnd1f39DKSv90KtUjAbYLtH4bAwIrLqZv0
PPraieWPpxjL6pIFvOpBzJx3Ef3gp+3zgpGupTfpRl7f1hLbaKH3XWoMaALR
lcvaXhrB9yPK/IZeJPsW5S9rD4+0I/Q88BqWe5g6vajj/hrLrX8BdSYm3q7D
TnLutvBXLb+oMVvEjH1u3ZHGX8MvQSWCLizoYQFK5emnURxSVUDfkaqpAoWJ
SJbOJXQ+hbNBLB8+CLG8V9/Kgov9XuJPCFkUpaCWZpmbDcokFT+zGlX2rG89
iJRhIgTB+kJ6vDVtsDvexilAlDd/YtdDLu6YPmcf4OSN4Ql4MwfVZFrEz7zq
+O1o4VlNlZy1IOeXXDxEe0+nGxWsc9qW7mYpcxnMTJ5lTzYeEKxenryykDtc
0N79mD6uw8Sam1Qh2J0wz1YbNgub+ouX5qo56xx+FeBmtwp1uqgWcijd8oN1
gCox3ydmseZQ0FEARptKeuvfEl1mhJWNh488oaJJnS2EnJXeRAS+K0AJEyE+
EwJi+LXJTPM9Ras1ES6xjM6u4fkOP7F37kHfV02V+POW8guPdzFng2VAdTyZ
nbu1k1BXM89TvzujOdRth7lU4URHpJlRo0SystmB1rdd45TuUCPrhPMuYSBM
Y54Wuuw/3z8xUFNaoBZeIyEAFKvkTs04gZ8+TuJM1dvsD8Tno23GbB77hVQ5
jSLzfgQpsoGUmrVCfxh82JN8qUnOkVVsIAqDzLrLuHSHnCb5ono8T9XF5WGd
1qx1S5mADXwUxNzjo6Y2DDEFD7fYKXq+3p54SPUU+GsfdDSNi9Xxkpe2VHbl
0jooylDbJveSOlKXlqm/GP+zv+1wfM2rHt2Jv5uZb7aT4g0RsidfIoOfkBD4
tQMPZauKmeeFy48Z+ZTCBkMUhqAUjmHZm6V5gc7rhdIDWvxinrOCiEwJFXGZ
jO0zZzQJYSx0vWEld4fBNkfY8H7PfCPWRybjw0rsC03W6edeksFkcSqL/Uva
3ReYx6PEobn4Xq5TPdAzJiFO/Mx/VJZngVz9TMXu7K4J9pa+8juDEMg6UtbP
eeDUMPPS5vZIr6MPqKkV6olWHDpU6cErb0a/mBzDYyVOiRYwDjE1BHBgQG8F
UpHhF82JORsa5XAgfSqzeIp6r/Y+B99abmAB0L1XS7y+vnG3CHkGo8wkL3Cd
cYbpVA0U3W+X/BFWWXOyoaBkzfgOfZl5uxQDWBCwXWkoqrCOUGGXiaKBhT1b
rs3fGifVlR0GsO8JprBcH7Nj0HZbmDzYoItcw7s1bPsT7uxxmDnKvRpYmUoB
E9SS4GO1IOT/HdZBZsYnyvjTuOT49N0ggdf23VfnheX2neFNHm2zPrDQK6MG
cB8sXTjXAh5wI/ad9P1nAr6Q8ANgFcyJ2hAZin/YR9gFyt+xdjz7xK7kOwhJ
bs/3FazQZp4THBIbKT6QVy6P4WY82KrWghswDHVpXNFyGVHe8m0qcb/1WUj/
tBBMH8WRMlTAiyeZp1wHeyQ2ASmVA0mFHAPSO/zXG7IVt+jhQoqHQDUHw8Rj
3R4++Bumjt6RiJ7Pg6Q7Bhndwuaxh5li9disPZca7o5auWeqsWqLCGh+VObW
2Tha8eWnI9/Yg4VZa1WZZtPO/9Y3G+NfJhQcQNoiF+eG0cVSH/lbNi+xLwxl
9fbJ0Ap/bRQJ+Otoq3VRMcRC2t03xA1TCtH16Mf+MGgVq/1bNKGhi0Xv+zd9
GpomFNjzWcRCCFWRmbincHhv9FvfTnU+6CdiSy/6aBupjbLPcGjwjiHbNdVx
PeZusxtWjmNKCzbhsxD/snxCi8wRouza9J+egs9DNMTrQjcBGA8IWYjFPQ12
tl0wM0uOjgrAaYNxpXlS+ZzLwGy30xYf4vJmluPiPYlzZqH8uYCuOpcCV0uj
1YGF4bZD49gRM+kKKQgX4l5eu4jpLIIrqgj6/D26JLOo5ZAm0wvStLIDMm4O
LIN45hXOl78BrM2e4OZ+vJwREgBE89wFNb/AvDrgql2kYbe6Xb3LSp942i+D
6oktVsj0MYO7FceH3OpIKTAo2xs/2xizyR4nOdTgIC6bS/0gBJ+XqiPGeS2D
eaxTvRzcwLjkAOeEk8qJ2HeKxNoHE6LlVlvza+oV26CXJw7KJ6t9oacmHKnW
+dklG/LBec8O7SOpBMWxjMH/bbl/E3QmVPUiVPCuxeQQnzL7st9/mbcfqh9f
5+xI4t7mEl2rfzQZHXRH/eV6MgSJMNZEQXd10wSLIU8i8/3FJE8yBknyZcqG
23xPwNd8cEtdv9Fv/UK0+C/XwLZ8JS8HeIDCjSP69oEoQMx7fMga2SPpoWQC
NI+SRBHeUgQRFSjowPVnrijYCcsdFWfeRU7nIFVWDBHNARA9VrMnV4Bag7uR
ODaFJey7dGK8wEdi1UsNArnjix1laoYDcPtEn1VpqZTwAyYgXkrNUKidw5ss
5PcikOyvXgvq86DYLMDb8QHUmGeFqmNRZSBfT9WUPP4oBcBDVJwJLvrnK3az
5WFGIdkmYB/BaBigWZDGgqNDZegINbtgbV36dar1h8wrf7QuwzMRUCTYOsrM
GiOPQ+rWeEKfu5ZO3tGU0dGLd3Wi9mevzI2DrSf6fL384mLfDr4clScweQ6I
cU5bI0IppR5TyCL2io66WMis9znVUHCgOCogYwQtC8R3uN/KmnZK9jqsSaT2
S45A/vOcFmTPGOKrUx8hV1/V8pFdBcZnKXN/MSoNLLzj0U7o6OtA7crz/Cvr
ydHiu1D6gAe2akwkVUATviEk+wLJccQr6JOhlYRsUo3H1N5NiNRlo68hxGWT
C7y+nFlAP00vY6uy1MsTWh15Glej6Yv9wFQbXNqq5uOkFS+gpbHQ/BC0Zi9b
Nl/EesQ8oSeNdDyCQb+me9FTZbDaoOBB/yBLp3OIJfv3ccXMDg9RIVq9K7n4
XvIcL3wx1rPnvSSN1IZs22/qbjwK2BwHqrSHJhKnmbAsB7nvQ2+N68V47taX
YAu8LYJBmINm/9on8nB5OvsuSioQqDQBZI55Dvr8ndaZUCIEbUdgRK5G059t
EId1EFj/84iY6jnKNSn+rpPdKPnwIthmPHeFUeIVnO9CCvpeeV3ANtZaxEje
9iBFxPqKtBn6CC1Lt2IF7sBNrHpmYSGy1E+aIh/eovIrl+cPrW7wwHUvH8By
231/43rivjmJGRSYCav3xNwp97NsCZ53ghI/OeDuNPvKcfijIM1eod0nHd94
0ex6r2lBADEGxclX0ZXwWkIV8LVZwqrdY/2h+bkMPdhtciwukJV+7aBq5pfD
zMFadeleG7hj6OK/lPbOUa1s8+O5F+1w3tePBaNSUziCHnPoOW9bZm8dM/i/
5GBBA1x8BKZbkbjZ5XpxT4Ptlp1WnTl0jTA0GFsz6AD0pdEU3eaxq8OgOCVH
nsepj44wl838DPtXbjxEIrI0bXm8ww8jA42NBvxsa57Jt1w3yPMKrNfvihfE
A0pgUFNxsACQ7ru7+pxam4qMykpdizEs7zTZa8nSC1QGvxeyEgEZRJIyphG+
UsG8Mojx4GXwwIKEfqx5FRU1krc3ui3h5UuSDlcCYXn0k2Tk2VBixfuCebXT
ry223xDdulXtTmfMxHmOwbHoKuPzOACaS43g0DL9306JqbbEXDKU247ig+eY
U8CP2bMzIiEixYaf44wMXo39e9AtrbcUrBlOLQ4B8hb9xKnzNf6YzP2W/FVc
cm0qs4+YTTAXMJZPUMpDsqeOGYg6VE8nanZL/kecForzGPSlp9jalQjJ6LJE
dZbh9xkCXf0XEr8GNYaHmMKxF+kvmrX09kqYA+JbaZ+Nim2ajXICYV+yhb4q
25n5Y8sWXv0QW522pBd0bp4Hsh0WhfizFWXWAKfHr6c0KKthUiyawh2TdV2R
KRcOzSoGoU+5dJ25BIidZOgDIgltxEB2XHGVtQXQNKmRwe1t/G/xBdjTTaB4
nzomZOD0vxNvR6RohMrOmzPfXAghNjym8muCzNd0Qv8TH/NDf2ZUCqvT4Ux5
+c94hOjM8ByS8BXNlOsDJwV60xtSuLUBy6GCXKkxC8EqDfOBH4M83nMGTyM/
psDxbYD3Tkq7dBRbDgkL/CxEBR3FUA7bqsJzKtWnHUzM62rYXcM4Ff8vLNva
wqSbp55EgF7ZsxeQFon1JJFyTGBx91Cn0S8cFowBXZNTkxi/k5tJoHQOeQhu
Sezp9/F1KCBuaPyXrnVOUuc6h7Cl8lE+bV15yHM9xo1VVx6XzddWVJ+MS0Rw
rmWkoGPhEcLCklwX9rKo69UrDlVhjUb4vwYOwdXUB1astbYW+Ztg3B/TAgCC
QWZpWGt5PLVsslISkKzDq1CJqKh6saiWwO8NcslD2J0HQzO5hW/+PkSVfJzP
pbiA+0+uoS6ei599nNyr1iK21Y775ggyHnRImL0kBJ/kI/2yDBZIWrPEJ510
9R6lYDwcoNXEOa3eS81Wppzel7y3wFmxVB6TzfJRIejgAgkGNeTHgmYPNJFa
rQ9wilOOOGTi2pcsP1gwnyS2Ag3zJifG4eEMzDX4spasBEFTtPD/QjCIakJ1
N4oZEnEvcaQTtAuHEPWV3W3NVR8zrFnc7mWkIlKUWv8J2/lm0QJTtgW4sReU
i+PJPScyeNCgbyjotY9TvP4FVXvL42jG3NCKM0PijTrRo6wBhplFvYe8H7lP
+h7j5+A3hcb3c6vWnmCaN4pP/cvs9QurGGasN1ynDOhAMZvPtfPTFcBfgoLt
dhiE1D0G1YmZrBTrJ2CKDiJiafeusDh8kSuDAxLJeZq6RYV9VFuWuVSM1V09
TVKZPMYBm3ifZVSH37R08MFuWJMJN3Rc5bzJZzd84P7vG3gFiPlbZuafWqUu
CyTIJQc+9VZUtFNrwDEzLAir5xOsEsMwMn5RJofKS1dt+hMPMvfcOb9J1vi4
kQCo3Iz9ZByxUfhLBeCQOw/4tILiIGu+qcsoVTTR0TWohP7f3A5LDBog7zRX
9LK4cQL0G03nNyipZ4649RDhH7fnx7bp66L4oBUO6uZJNURbAhWgarrKJAN/
x6fFH/0S6CALM5T6UNgKUZlPJFeHkgVIrdqtFOvofcL6ftXMIobn5vIvhGj8
VV2+AbbX8g6B7+/MTE9IV372nDLj84mkEbVmOiW78gR+xvFScrL4zvLLo0x9
Vn3poDtaHniHdiIVqcXdIGvNrTMb2F2WYT9uI32sX/dI/xcEowA3HLagEmGe
sKkXwDju9+m8sDnLRuymskRpat5+8FnI2vhuRxtLVGOzdl8EmxCtfodP2jDT
AwEYukH+4xCCDARuYeqKlDrgckxZd/onmBKpTYwdrhuvovzvsUfmPK+JfBju
ggNVBYUw4im8U7TZvSCno5lCv7aBMFBrVsr/Y+3teHFFcpw7tqLaiSzeaqpS
q/dPo8+SnTh6rwP/1GX7b3xXfg1HwEPHvoSHG7yVzus81o5lO60sBteK18oG
GCd1VvbcDPU33FB+AlChyRMO7HdReh4Vep2MO6+bTJlI5FCuq1xbGaD9HOgS
aMEtCiIOCr7v8N9xURgaQWFhU9Xu3uKuNWQ5klbBG7TjxEDajKNWcDsfZ1t9
uNNoQeGljrIf61HKECssYlOH0NbZAX8b3CqGEgh1gPtiwKfBCtHh2l0ixj5H
xU7KZXgWLQzqPGYJY0uE414AQxYrQW8uAdFT4APvU4jrl9SwhJEc2IX+6yqS
j886uTGDCxX36KzoZm6iHdUWB7NpLu/CdWVEeWlDTTbcmrDIuPLyHDNr4XII
NsHFBtT06xEzCAI/c+1P1MvMAaOBnTqTMFyZEjB7wgIMJ9YGxmeGTEIVH2vF
pSlZdcpF47dWoCZv4i9925hj/TVMXuyQUvVjngM9wf8xNYnKi7Ctq+ofnFMb
iXILU/Lw4LhoXqLZWze0slOdYj8LXwbrVeqTRAQg2JIGle5ghwaTxiBmnRMG
4ifKcHhI1RpHLN7FYENJMxN7djjsL309qkJ5lXRqEp99hyw2T+U7h0KkypCc
KQ6T6N8O0x3iZcyVic5N8MFmZUt5yGzmww6gQipysTqMZDey0nnbxBfmueMY
oAj56m8qVMkB8E4QJRsPs9Z+Aa/YHE8qr0Eu7gPBNBE4W2EslNKvLjXuYnra
esXvFvh7XrzP0cdBlbgbbMWFj0QxMpgR5GiHLiT3chQ5Jtj8EILCAgq6rZFq
tRAtODrq0CS9y+S+VUr3Lf3Pkl9cqOmoX9gTQQnby+t9LW2Bcp4MN/WbfXfX
9SXc66VXWEiLPw/fd2momodqHxMg4T+xBMW3TJz0mZKDv+7b+iw0bB9ONyST
pS6fBb+HiTHrF9l3h829Ln1vSvNUNygkTA0HgVzeBmxjdtKGie0K24wuwj81
m2hy1SNoExvf8hsITpVZlmfMdzNJKZ8Gfs6VEr51E/49ffacZMkCpFR/IUY1
oeZiSyl2BOr4vjTyL2aH3MC/Z15AnFCPrKwKfrHbtqY16w8de7wVxod+s3QW
q4abvvEJaFxhurjC5a8sjAbpzC5FCcyuNuoSSDjx6KLgSf+wI4TF6q8pUBfZ
Nrpdr8hNlG8irbq4YOG1b839zNvSx7t4H/p+WIGm/4KV4JAUQXYJjASvpBt9
4YaU573v0W4nUJYB3jBJ5wWhgNQ/Wt1gWaU3dzI3d5ihMDOe1Odd3QZipdQx
+RL8e/9fgeJf2WV2phbUGjNgGLvjCDCdWHhYcCuFGmBrE/6VVnm2+UZqO5ez
QAJOUKu4Li3oyEki9QdYZ849Rp64TQv7wWuP07+hR8x8NAOvQns0go/1hZbk
Ul3+pGbQYGtqz5OmAWjuW0DmqgJMHjDjAU2oBpjDOAnY3FgBCe6lMmXxkvV/
IAzcxizKyLdC6wznmoSkJDAWYKPeSE1ROb2zqN4xUqKHk2/Oz5B6iyoauYP1
W3YXUcdDJgHtatuNkW4Y3X7tao/1+k9Sc3HK2rXE73ZNJviUih6GzUYbQhvP
Q1pW7QBC8dgteg9xfDuFPHhLl2Vvp6ZN8Iv+fjsMGvSEhOtu5NmsOU7doGlY
1J48Nquo0sLN+0uIveDjZXRH6ap9m8qkfqYhlUJFoa/l3k8f6UNuC8O3xClO
XImOtWrwMM5iIYWhIrexuYUcA2sHsMRP6E+AqP6YwaKJu75qjwKEAzvgfMw6
G+/4hdZ36tlh2a1LgHZU0EltRFws/dhomeBVntDLw3hVGyRxdvum5ojGoCHr
PE5IZDNAWxDZHMTziKS9MOiiHNpL8kCIqVueXCqV2gB+S+mEJmFrSq5++4cm
KaUkE4xN/RDI6gfU8YdJAFKQo4EIRrFKqSRdWptfNHjzy6/QqfcAMmR42Ivb
Ub9ok7g8I+n8r3VfpKXoU+tqU/6LDaJQWPG0SepYtyHt13KXF9nRc30GmAVf
+AlfVYfuyHH+xJHIVTZAy8EfhJHiIZaU7Daqgrr6SNpSM+NbWz1Od6DNGC73
92UYPG05zJ2Cz0SFQri0DGFVN8xeMWPryQaZsaPaAUkttiJh+rICM8vwbz/T
9ot9+eTKnhXarbLLgDVBvZ+GW3y+s5llOrtZkHi+9Xc3h50FuZ6kv4XZnxyn
Ds263RNPnWo5ak2GmZsjuI2g6x8xhKfCpgQMWIYy2JGqdDAWv55Ba2d+YvVs
eCqi9T08alyBs7Z8b8NHyk2TtMeuBwtkFN7WjUae6yEmTY2nFCev7zVqkRF+
2mXwLVeJa0CHRhKfGDSWfzXNBaCLBOZggMqvjnpjCrVNZv/fA3F32Z/Yac7D
4oIQ20ZnjrsRbJJwtTsMm6jF/rQPCQ4Crardo+hxYV9T3lIz47XnN0QQyrT4
ASKX82nPdi6JS5q8Va/6E7PNVkowI40qEdwQ6vMaf+lMJsxEtsZv45cVoKJO
YES0UR3euObhbCkQ/9XdSxXAryaq39/ibmMoSRD4a5rnOlcAfjjaYSqLDfwS
X7X/cKqjJLYfVUQUYi8xkHrbrYhLYu3uSf382dPdu112ob70BcxiW/3NlegB
XbA53yHEix6Akbo9kHNi460ZB+6q/aQ4d3wXNE1HaqY9m7/qws2HpR+0wU1A
LPcarwBbjhHD32R9ijo1UPYqTRG5ACGBQScSdwE6TWXPQ0nQzMBgyBMPsMeJ
P5IMg7mkUv72fHxk2m54tN4p/BfBowvxUfP2KecYWi5C69qtleHraslGF6OQ
W1u972PJNbe3uCK18GlZtEe63E/z2SZ2RqdYx6FZtgJcFdf12HNGfd1n9brL
40FrvT3DAPIXDTDauIE8wAi6tc7FdGHxB12IExLtgb9N64sz04O+SCa9oVip
R2PjCS+FgDoH5QEi58TKHw52uBC77Of+HLIlqa0GDHfI1d6wedZxN5WujY3k
2aeW59PZehwCOWbTiQJWJPlPzCvrRtt9dI6XbqEJv87ZAo/mfovHottoX9bt
HbEG2Sph3PL74WowobRIeprg+8uUT/N7juKLx9oWHn/pXazs8LO8sC1pX0Vp
EUPjFIGffd6PH5OiXwW6hri7HTxv79be0nam47i6vJ7QSTCPQyJNHyDBrCWF
IOmBW70tPf8XyYMH5/zuqmluCP2TZabhuFpFuInaK8lSC8+PvcHKmih+qTn+
xS+C2S31oO9mZNbMP5MgYSrvH0jiom3asCFZGPOguz7XxhxTjeMLe9NMIGNR
oDMecyH+PgAgVg/au9KgPpm7Q5bOH1RC09LZAfNUt8aEl3Z4XjU/09tJwMjs
ea9PCPcCDgJdgX5XmnzRe2uQy8rQdWmSdb1hjPdYGa3LjMqaLhiSbvgP7jRd
yMTHf6ROsRdni51iOF3lwbPRlN+4//qrLNHW+8Y4w2X0LDcGZUFEBFqVvFJ6
7su9NVr7dxMlUARPJ/11XTtsAX3URvXK0x4tgdHqZx+0uZ5cnnjzEgI7z6qV
5VAiIMqT4jbhT4viwX4Rtj/PL38FQxgV/ub5oQY86wmfgvq50h8OetYY6llT
coSDpSDx3HKRfzKjiOYR99PHtHREA6BsCPN9LZyJRlVPGQa1eUjFLEP3CvTu
7xB9kRg50C4hJKVR6mXzFm7hCuznWwHehGr0P3t5bGdhNTnFTRn6rFyEENt7
ZPvCqNQ1Jnf6AJDNSG+EOoOGB/MtO1erW2vQ8r0+EjSZlwlzT7n4XH/eMzdn
kqSdktLXPk7S1DdA/IrP6j1EffNwJk5a4gGikN0UhBJJIxNzei21DkPYuYla
7gdfD2MjVl/YjurKAH6TKfAvpppDbuDkwHP3eUbrLeDFMBQWsPIkNoqFTc3+
+mFihhnWQFICw0NITgTzENXb9ysrDXjFoPofXv/p4AZeWmQqOOUVDgI7G4aa
G7YSUlimaeL4JLw2Xh0Ap4Yx7ceo8lkcb6UYOH/TrSO4L6hawnhruYj8VyGl
tcekInVErqx3VBXZFPuKpq5Xw/e8jdXiCBboPq/lStcuQlJQ0mMZ5kF1WKXt
a02kMflFIbIloXb6m/qWqssfyRvN36shnvxA9yTp+JVRpPeebNI77WROMlwT
XeUXB/EQWBHohAoM3JEU9NcUbpdzL08lTdx1L/LopgtQ4AekWgLhHhTOMm1B
894iECHFVOvXDfadHnXWDXrLJtUAnaWEPycGlVPk+gwroBdAftgAIC1T90gG
Qn9A88f0lSEurv9m+NET93WSIhBXIHx28xbJO0KAezLV+dRE5wq/ifwzY4qO
GXdLsx+kmianTPbHMJnoOPNbpFPQVDHi4cOx1lFKOEN23sPGh18vu1PltKe3
aK5cPDXSeWPazoIUpfOthrc+xxyKld7NAuqtnGgkMyrN4rQqcXWZFuydC8lz
UqRdotPzsWT1qRI76R6yqNPaZIWoRXhsX/W6iujud0LjwzMqLhBoTwWZjFcr
JhWTSnvHSLAK7uKCuzSgLZs7gljxpjhN9B3N6B8buBRvnhK9fd6etba+b+Xo
r3S/U3m2lsTJsYVnCIXcIT+naKhbz2FebGNzl+lomk20VqnBdvJTJ4I+b+WR
hv3amCJwGkkcb3fP7V3zXmNiQG6aOxIUlImlHpplITd7qpju8pJA+wA8AxKg
82l48Zgd9ZtN0kxJTCR6F0mhUSXLmpCmCkxZbJ3vc8uWkxi9oJk4rQ/wCFvL
shQUP7rzJQ4OnqfMh43wMdSvimTupny7joWh+T5NkH/39oY2LPP95Blh+RVp
UX0aOhQAW3LDmk5731U88A9wP0ivUASAGFgFMmAMCTQG1PiGZ2u4yDZebdiz
ZldI09aMS5DFVD0sXFYZWQW4gU5uZ86LepVXKp0z5UbCkHI+jTR7u8Dm+z6F
S47i1vN2udXo4mL3jxFqYhcv5Hb+/NgrtJ8nrfrFmmOB05pt05+LgPck90hm
sVHfRDiw3mTeSO09XEcDbC27iPqNDqyHlRFeNuVnSVR/UunJsx28ACXQVF0m
dhNa4RGeHiv7LdwVaGde+3zISkqqrV4N0CVP/je/WTLiCtRFLoUa7ZhQ7uis
XNMfJmwuU4dFgJpW9pHTASsIwfcZXtewvokBf5vwC+FxdM4p+mLt4avqryaa
PFUmy1RMVZPTDg3IBO5wwAsA4ersoHXLOWPonmMhIy2cb1ej2nKaZxm33iO4
FHBm5CR+7wStUkdNpzXcfTVwsyk7xv+ouAAKYtzgagQuCwCrsfr7RdKBiTUW
FL2/1p5bGXuYgPUlvXwYjZBBhweMNXapZa0bmA0xDZFs0X3UQOp9lNumnSdt
2OTDGs3jkvyIchw3YEXOpUyUSRIqIWT/596kbROsdXafwEyEmICXxERIaoHH
4AYQXQYydrwKXMpclB0oHFDTDHEzCLmRWFn7/4GWAsWLEUOa3QjO1qyYx2YH
DcDSzWq3fQJDd0NXyTbsBb7Vzyn7Ehb2ksjIYqDnARMhhgLdPwd29tVBJepn
i7ncs0tE53o1cHJCijatqCtHLpr5tmpcpVli3QrlVSTvZscTI40PpcFMaXOQ
1Uh8nUcNm4aHr1y/sPgkvq1vpRLucamXomuRyFOCl5cG0uvIxh989hIi6QAz
AhqSq/VrZbSrDXOZpkCQPQM57hhjuspKwSZdzuFq7aIroHT5b9vVwcMbCR1V
7BbHW80uxKyV2z0uAmWk/rsj3+1WP0RyrPc+WKOuRBzBpywrn5OFyLPTFMN0
PUCuz5dYkyfcyNufHvRWDq4ee/0ppVBsbkQd12e3Wq9mCBUMxQd7H0cNd8OU
lEW/y53Y8oQiW2y3WFVvk3QxBBueDmokejJsD1wa4XrgKth0pJv5L4D4geV8
HHyHucyW2NWA6zhSYfP2EztyEbBOYKjU9kMPfi6pkQ5OKAaPf2o1qZ9PmhvY
PywQcOeFhYM9HVHMkZ7m0VJtbEPxAzQenTMgVzBvxVat4Nwt+91hUp+ivaqE
bm98A94ZtvOHHmatqn8j0d/NtI85ZlJIEqAC/43fIEcWFP22mABXG8PYn4V3
Wrc4GoA3CoPx8ctF51CMF1b8QVJrA0fqDQm3KvYIr4wgHYRMHaLPhOFTX4d+
rB2P/sSi39ixF8kpc2065KxMgDy6m0O0sO3SVk/txyyZya1aZeNuyLl3lNT7
XmtIxi7HSsE+YQ8CDarb9Z/qmofus3U2JF6jI7IePlDMRLvhJd/U46BRp/0J
SBk3Ie4E1bJ+yVSJP9tulDT0QJlfAfKXK/8nWc0DUJbD0FWqe3CqCczihekl
A/1RY3oY2shtMHl2v75oai/HuYIKCnWAW5BA+VYptdvf9qPFLu3c6xB8liLj
797CmSnOBOVGnu6CqF1TMgmH0a+UJxJF03EelMwsKkYCIVYD2C/2uGCN6RHt
0/VHEsajAwbF3DuiD/cKsdRcBauGcc8wDAvZU7qDZji5zotMfWXrPTz31uWp
c0oLlgrL3sqNal/NKeQiWjiTyI/ydBOnZjqCNswDCRqLo8iZcjcolUACKtjE
kBiKJCEtePHekpqiTSfZCOZL4itdN0mczd5TgMPBOKEBYdaGyDM947UoTleQ
kg4aDvWXhQDQnvW7b8TgJNQumei39SryBKY8MJsu82cSj2jrRuysVibg3oTx
Aim5PpV50YeO1RmFOkDcELqi+d01Gb0Qjzf9K7U/xeYD96YqkkX2ufH4QZUE
eG5lYw+BuCUdINHpipbh9ZsehK1RGITsZZgSbOG0RZcyczLW7yEaAq0xIXKY
uoo8kPyrdMWiMaOWu9EsU5dfsvejHA2g1rrHylMwapqYlrNMP8x2dL9IqCV6
J1hox5KnjdoJEiJ/KiWvjM52YGojoeKyhLhnSYDfF0wHx1c7VNHOwezsbMm8
VzYgAvatuZLfIvb3wOY6WQI0jN69xpURfsmhWW9cTV5nCwmqzY8ZBIkyEhch
aBqlmVlgrnsG3eAK6FOamu79bPamrjnA121VmIX/Ui+F1Hl9dTO3mt5/zUWs
sgnxaBquIzgvyZ2RUcsjVhFqFlhMVQN61dAsYdK6aB38cnvZN1x12iWEIHb5
ABxZGIpp96fZy7NFrxJHYBDu18Fw0UoYHouJSbNc+xF/0Zd2WA1VG4O+byCl
2pLhjteuD/TRQdlVfL2Wk819nlqLNZCNTgCOEaLCeltRUtjOKw5uoOHLrheo
QA7Zv2OnfIceWE/fQRrwf4mNyLnhOerUtgfJKJGo8ShaNpqIlAev+staPKWw
hnXF2d8b/bNk4aBfeH7q3cU6VRmiArYtCTGQ94TMZH/D/0LdnqOmkLD5GLM4
w5p/cgDCjxOqFQ4eGxDOZS6nCZJtdtS3XI+K/rdACyb6aSx9pLWCH/Rx0IsZ
M2HoEShsNgsO6laqLNw+8AR8gOW/oNFQzUrT6Vh+kREJoTP9QhxyNOn3XINJ
WQnHC6a/8G9LownDXipqJMUqzkvcvHfOJMAdkbY6LI7rZ2VnfJaulFY8zK0Q
5kt3aoD7iWGkACGjc9RvhBtbnk4Dc6AcdKb/NSmJt8CoTJLjXr8m/0MVda5j
TEOBo8BEExzLr7kJOSstEGy+gcwUkwkx7OurSVQ4ru6XpdhPVXE1OqhFXRRf
oFdSe+UK+wl4W1i448ySTqvBXrhqPKvYzIDpBXnJ8ArA2fOpTQtAR36lO1tN
GyEDe/e4UG49x0B5B5k4wqpv6caIWH+B6OdSqsc7SDJB15sE7mZ2MmOFlyW0
RdkV7zZFc8L6jWeZBdoEUqMVQh2bjFcpxMovi2GhLxVsIFC9nOv0x2V4ydso
FivI4Brk2pS1aqPZh275lC2cS+qAuucn/Et47hF+Tm1UP9vKkJvPXWlzu1nr
BKGVeMcOUIEApKezmHXb4vBQlZECK/I/NxIlMmdFDnr3wsvA27MrUtxrDVQP
Fg9VUP47rnr3VyUNPiC+a+n86YIiEsQwURu6nMbylLbmNYG3aVaoMj+gyhUt
gldmNojMOExqGJ/wwswFjtRjYZbgSJX2OcsMtbOuSnu+6e5Z0uZl4wpn6G3W
NZvRYKb2+80ZyED11EfcFE/bjqFpyP3eJ+cg/TpR3vGAMYl20bM3KWwl0KUG
W5bEwTusC6E8jzsFQrKkKyFG0yNBt0u4TEqlpjZIWAnoIjjzMg6+0r5Erg+6
hrkSSqw/oFWvAKGZz8u896KpV8JzLua1STtEi2NBzU8WvuQBV9ILpgTEW1tu
NB0G9/iLC1ZcZ04eX9nHZH4C5/kKvSB6tk5JFB8VY4bFKaIVBJao5PSlV7ly
8ThYipFIr7crEbAQ49/T+gJHNXoRmJPL5A03hZsAkcVPzDf2jGq38DTT7CtD
Fo7dY4JRM0J9NgkuIvxSjfRIqXOj8nScn4MgH0B+F5rJUaX9/CbPKifiS9iF
lHFzq4PdIrQ6MmZ3UrCxqeh0NoGqTQA058ZK7VCyHK8T845xJxB35C70kClb
teoRD0y57ScuKYw5LNWwpKHrlDpGIuQcazFwJehpjc1tdbUZRTFIGQq1Y4D8
1XCISH6DXmj+54YA5TvkYXSHQbgflIGeeEXdamBUMdBTyAgnhX+T2ZrWnxdl
hL52M5oex4ZdiA6Zm1kmZLwHZwEQYIQhg4TEq36/atmrapk++i96AS0f/Iqq
oUQaqRhIDtoqNAxU+XSLq9xIkJJVNQt9wu2T4CSHeDSAwaDMBUidqCI5Wf6D
BQcdt0y46ly/B03IdBFYQ9EUgyMkcRAvGuVgqq5+2xOG92SOkNQyuSto7Ypu
oB04C6HJIHAWTHRy7WkaycdOQPbPM3qs8xuIqhd2tbZoLSrMNV4opkjZsI0I
qBQQSoV6z1d+JYCN447chfkTBUKUcUQGA8c6ep9g/nBqnFHs41NeZaD5ebJr
4fGNQnrnyi70MRFBf4PaG2P67ifr3cnZ7WFNMwb3DNgOWGFnns1yb7l1Ia+1
aIWgRmokRL17AwDl9AxHB0G5fk69ilV7fhxZGzdCchYhQB4Lq6OB4cMUzX53
e9Ed2o+FtY3XdplX30yt78r5mlEv5n/kbKoP1NXpJEEt5hT8798iCuWlZc2x
dAh4FVb3vIS0rCs06hKMTNAiqmf4RpRjy+rgrQZ0EJthfBKtki02EF5ILjxp
QcrY+1gcuzk9hB0f4RzoMc9HPgbawwnYDVc+8Bjql9aQ7dRGWJ4cTTHpcidA
b8FMLuwBLv8/b27fY9QTPh3CKr5HdLtSrkESQrrfXONohfx6+CIZQFqgDaPF
VOGe7BTluH37uCnOi8Qv678DIauFaJzoQhlQo8F32f7m29P3gKxuA2xGohpn
20X1adPr0qAjB0aZfa+5rNM5oSL3MYpXcMIU66n+Bcs+MQHY7d1FEV2dtF5B
d0BZmBhAF2KYsxtT7jXE675BfKngg4Q44/WFa0swcmRyfloec/+ZOWy/ROin
E+eqyxB5s2shJDFpqk/whyGnyeVpNFIm81oy8rUt8ZYIZoIrcBQC/v8hsGhL
JLqyN8u+knNLVzimmsWCkBUPc6d8t3xAngSG8UOF+Aj56oO4Z8RCSX+MffTK
oyQG2zhaQi9yRT1UEC3BWUv/9VHHDjEhDDbAhP+53Aik4QOFWJTFf4p9/VcJ
x/dIcvAI3ijU4U2tDqonBjubgsOdlShqciqPSgeth3BYKoEqNQpyOQIUx4e+
BWghaUQ5Tx6aJq1z6fNTmG+EXM/sVUjcjXUTtAvl7ILkIilwcLbGpSErQk8C
+7iSe/bka1ot9N6Z+jMvYN4AKhqfBwBzqsN4CzKBG+Bu6oSh+l1q5I4fMSyw
8IZVGSpO+966jYJ7eUOlKgFgT/ZAir2uvgI0li2G5Cv+2dcZIJuTsdaPhTa3
ZevhQmvMiuQO+8RK+W9OX04+HixCjxACPiMvTmYJPkshlWHZg4gxvpDN9GeG
bB4uk44Hqc0Xaon+VJ67JEfs54H3JZvt5a8TO3DFdbnRj6MGnkUoPPtkipIH
VJ0v7KuCT0WKos8VxtCY3ZhamDpRG0T+6DSqrGoxlYRRuk0cwNhfMWLQ7OWb
HxBb1REsIZp7otX82/X4NL+YlG00ak1Yu7BIRTm7VIRxH2zo6Ep9/pgDSUXB
9gWFewW3q3thbYPCsflmdCcqOuJJHATzKCRw6Cek4gsK82U0BnAmcB6i0o8A
YRcOf7U8WkefHDweG7uOejxACqrAAOn34V76cKfS2SypkbXmWfyjrhH0GYS2
E7DP3NWRGwpWuVRA5opcfhNkorFtya11wSZIEcZlhCnWu28wlJVHiv2O2MBQ
fAb8F5Xmh9/m/K8e8FEEfB9TJII2pf93XwKoHNqQLZXxMzAObpHCEeX1Oy6R
pM9iIcNtQFy6anM9muTjrVMMMcpgsBoJP8R6/lsr0d19DDjhrswjJEED0ziI
qesUsToT7VaP4lx4Khq8ftTKqr0c1sgsWa8hCTxVkHlQOf1jizWKJWt1wa1g
oh8rOc+vkjMNrRQTj9s8H83YbZ0ZSmX8ODMh6UJKmDIJ5U6NYFUzLdKP7KP7
EKuu3Xkh+yCZmFPScYrbV6b5yew7Pfvju1mrTli3vCTySCnDFA3ZdN4Au8Pe
6pSUswN7KgPED4QSzJBBJaCqkYBKEpaUa72oju22Kyw4zz4tTo0A930pDRMG
jGV+aDZPMpzmAQslL2N8+ql//L8iX1K0t2JPY4l19m2i7Nvy/43IZrbyp6sE
35wdTVFkrdRAtYG2v4QFe2lryfAv4+cPXREtBeEjM37dVObbpxlUFUt3ihH0
C6KTS+XPprYh6VTis4wD8kNVDFUYwUiycLgnunhOOPqANBQ8XsaHB0WG/EW0
xPKQwuyEIi9yynq2aFlUWVt5PHQAEHroh1SQamzkp0FXlDcbaoy94eCXXa+d
ULgdzR4Mqad/IuCTDxKsS8MXGjH/nzaNx2POpstEM/EAIzJkkjwyKOfGSjZo
JIZylt6bSeoLa4NssEy6SQT7Ym6PpXStFE6oJa2CZmx4wivWUVA1k88NQm2e
s63grk2Fe9EVxxhOJh5FBO4rVcfoh2tDvmHhw/AfGxC7EvoTZ9+4XOqS8emx
FYfPSJBd2W0VjZgwUfWGTbkoRCRmXEnqiTRzQP0REKGNEOueg3QkubgEwQK1
MvJpyp+xnfSekWfYnlz/QfhyTJ3C+1cYRu+x6Rg9MNJY9WP8a/AwopA/BtR+
IWXSteCaamdqTyrJ1wu+6m7Tum585hQiuMd72Hk6jbOzZrAZ4EJXRE72M2SY
lfbd4mh7m/Axr6KdowHPtfA7GcQ3FWgX5k8Ij9hd04trp5Ie8NtN87ScyNNH
GdrL82QXnZR6emccvJ0FyKb9pMiTL7smyYy4INQNhEvw8MBi4jR+lIUWUmn1
czKT3SnqJCYO13GTzMsYaILDDnEw1SGeLc0v/gqL/EjoZ5HC0lSJ1qTARBuq
9jjN2Bec0lKrnD5CYLd97RlRv9xTnoQXfyqVe/LzeaBjP6lSyIZfE8tL+Tcn
9mpc3p70KvcH5ViUg6ooFY6W5lOmO1AXX/cUkbxhxkRovnhln4ShrdxJ3fJu
lkl8FX6mheV+IbJ8C07MGYz0XKVFxO38QwwlLiBI+6FAI+XrktGqAlR/N/wj
CifXn3gB6Z6gD7kRk1G2GrkfLIz3yQDCaxPbnkZHUI5u7ojdB2oEx49LLjFD
xT6sX8RcxcKhTI43HoZyHW9JqGgrIttfz4nfbge5cwx0nQkw1L70yIsPl3QS
0DcI7xA0cjg/G7y2TkynckHsSLAmXU+6T//GtlrFhnji1fk4NWxGHNAD2OH3
bIn9zevmk1UMX9TfghUxkvrsUzxfSO073hLM2NyFcE+32MP8X07jKeZsJiUU
kA0n6Iwcc7OWM7Q+/C5p91LHu8i84Ba7GKWvDesnWxA8cWRRWapr/q3S2Dw5
7lLakJi5yGaVlMulp3oyJV8z98Bd14LuuUdf3651jU7Nct4kO/8SLCWfbLI4
BYGQk35EX8EwGAhOGyWizBg/5bdCzNKwAn+zVqQYiUSLiG/On5MsNeASYUmS
WXBU9CgCYP0cyLgJPtxP3edxqyNDtQB5gKsKKy5qM3ZqkAHFUbU12x4+M9cc
cJrbL8bYGqK5n92sy65j/t1ydEDJsot0rOzv+QyZA5oq6OxocrNU2ONaWEzh
DLRZ9C0rCC6BbdNoUoXZzZDRhpL2SqI6mwXBJqJYgToqc0QgzTGjs6R3sYXL
7ANlGihrumYhbBjapklpBKfY/Dqta3U+XMUzURg3yYrNIHbHP4hrAzoHtXFA
pQqrvuqL/eG4hXdi23f3SRb1oREs0Cr2OEmEgy7DEoFtnSZM0CzUCZjHC/hB
u90GOvbVzc6HWA99g/yL54UgiWBrABPzTJ3P3rWDJgJanvqY7kXnkXJj5tzM
L0MBJRHxocZHbb45VP3tyigTh26hFELi8WVp7gMXS8Z/YT6WkJr7nS6HW1bS
d1WMWnoXcl0qq+q4XjW8yD/ZLUTHw0Zsm8DfLAEWDFpLg4uZu/B3QsPeYjQl
m9pEAVufwC8nnuDa3DvHlUxEWhz2ERSroWRq5RLuQ6J1fR73vjJQEJ/T3Ixu
TYkI6MYb3udc0nwytGnnPQq3q+dnDWwe0Y4sAG7Ti+RKqAP1ZqWa+PSQeRqT
G7KlgsvCXHr7i8tFhSy0FypPKrqx/ka60qbqQ2MFhHmZRneyNFxttK0a2jRP
addtzIwbRrAAidQhqRKYdynHf3oOW6kUmbvRfO8UUGIxjP9j0Ij5kBSqTFd3
qxugmQS67qrXSHYI66WVY74x9RPRq6kQ2jG1Q9fl+7WR4zQtG25Qdi6nuFCB
Q+5hwJBf4JvaneTtKi54AVOpm9iaNso1w4Oj2yeAyPs5/JEvXYXXGepMzdyx
KbgsCa6eucarSRojR0b9UYbG+4/bhOjfSn+IlWfJUWN124xSDZbIuDAVKx5Y
q6NqaVDnq9TD6EyvTyTPbQb4IULFyz48C3rc1Oz4qFTyslLTcjb1lhGiOZTI
7yZISy/2tToR3wq0UEu3tuTDAXs7dm3THuibXn2X0IwFysNWiP2rTIJuvw/A
iKkInjrzKUMOOuWHITRHSVJgM7gjZAaT5uqsu3PhdNkbd8aFEWCCiPNHDdg5
R3XwPHuZewxDUih6hHOzHY+Wt4L/W2KfHw/g3sXwbXJvg1M53M/quqifxdY3
0Y5MhTTXaDPRAw+SG32s9plTBN7F2Vw8+b4/RsYeZYFHf7gLJLfSAsUrylpC
uo/zIZBPLbSDOMHfzIbc/WkdIEMkiSZkpyDXxOayYOY8DuskiT5ZL1euoC5f
y7oMoNQPekezrDshbxC+Zeel1FuZvTLUtOxAMFUmzoc8et6hZWZIp3khKMfh
KiWNDyx1BGWWx9Avaqajue237/510WU0BsqbejVEuCHACaZv1aPTYBZGDOTR
5LowwYs1ZZzh+Rf2cIsnQsZdFazFgPJE4aO7jcHWW/fJm5k92oXcjrMAftev
uISDp5rFKG72UBCReYwESu7NPp6HKjy61JxVoRtPeWOgysy5rLGsFj721KbY
NL0NccdP1BdjXS1og+kaNALj5guU6hS+EoJ4yPjc5TRNSNaBkrjoh7b826zh
IAyQAGjOzmnN9XBYI0M5py1oa7Zmogw9/t5e0Lx5DBfZzoZnAtHopJFFLxsL
Vg9kDzx+B3AFo3dFQ1ozVV5Thtl0t3cv+JTSlGeo9i5RIHo7mShtpxrNAwR4
AjX8NKzmq4H8/R9T2+MPIFK3TZ/uE+Or4bH0ncOq6iPI2joUr0lXG094Fmu1
lCLQZZPwD7AS7MvP5vcpXgFmuUDPC3YUrkJMdoeRFI4LWW3DR0ua+cjPNEQP
V8gAqmU9LNPuP1IxMxsUIcJA7NyAAHKOIsLTAQx0ZuuX+eGJ00b52wl+uci5
N2YDjUxVIMBhDbn5eGbX0Sbwx0S218AxOWTwpXOKZ0GD4gjXdRsAtQD9pOqn
0yu2q3VSyUdASej9HPD4iJDO6YvSeAYBqRj3iXpuWHd0WTLWlIUirrzWhXKF
fGoCP4Qcmofid66cqnU5X4T5O/L0FhxA59fbcbLfJDQzfqtoOfWJ74xgNzdI
SoJR6KQ6evjvAz/UOP165QXNJs4LEd1AIOvFqL5iMcbJXgEzDmEXBkJGQfk4
IQGm9YhGZn4uwfGXYbLdTmnNvaRwf+Pwwy233XitYbRmlSIioVE+UqXAwNGw
MDu7KghCePy8QWhooNl3y+LzvQKzJGHb5LwYzmT/uXWGX+14zXZD1jE5UJ2Z
+lssU3wNCKt+0+29dbIyllvgTvxBIciYAUbDhWHgBQBH1489Kux6XlgXgeBy
kGixdH3bFE+rMV9gva5LNWWDfigoJgO34KpEniEdmpZJ3yGwgegweq7Hb13R
nZLgpdgZYkhtcHnwPHtC6Z6dmJ0aY4xFaWi7hBG1OYLpKnxulQZw8f/59JjS
sX47v/7VzkopJErKPyoEUcXbLo2+Q1G0T1obP0G+HbL5+UWzC6YKQ+Pso3Jt
1nPPAbXVjwdHBbP8VCOqCcCCo3cokamXfKha3qxvrmvQqiy4lP6ipSYYFh11
ISnQs+fSQ834vjRsEwUJWxnjcguVJRMhIzV5aUE7oxFnoXAJ4QflOkGJjuY9
jZ53vHWuHuhY/+aCX0umTh1MAU4GoS6I2+lC8vuBz8ajXKlYldlU4AJ9BCNt
PrXLc/lukKmpfhXDN1gGO8KXAgEUN2CIVA8V8ESv3HcDBddm6T+ppmyLf/q6
p2JMxBJkZH0Nh+XFWqX/qdtyits+A4XF1ZWKKOLK1nE+DqqOGjl1JGtHhzHM
0L+st73OM+2FVz8Bm2FqE1K2iL5ZKrV1QoY9hohx/Y3q3WAy+2FAoNsTYan1
6JFC04GqJCYxkuA44YzZuyp8SL9VQZfV99AwuOXgq9HGN4EYiHYSRNVLGse/
OwZQBhqfE5ysn1qXjBeYhcXpq9oBsLPTaR7OpwMSXzvqp6fHZU7MloGXSBJO
op3jJzuqH47HPy6NNj95wBJcBKCietTqG60KN20nXHGdVyCveopFLVatefVD
RyCLUe6E+7fdLSNYybdRFr0s0em0Pp5b+Jy8IGY3M/VpakSwxHsEjl4tUzoL
q24cyO4iAUvvdrnA12AlmffRklNSZl10rkDk904tOEqi/E1vz+5wvu2SN3Vi
o2XaT3fXXNaWT6HSHZflXxvEBzDYels1JBM5Y0baLgNPBWfzlePJ27QR/Nhr
mAOcwwFs0BgZjCgqzckpU7JjcU2/py+gFBEbdnc5Ru0uoNKhoRjBUF5Jye6q
DZ/w0fjdosl2DQLVVJXIKReot68zwve29vabl5XjhnVMnhf0yaDKQy/J6BxP
wvU9/Y6RtV4JOOjJknGEICcSRoqRTGAtvMZbuZYti4LSsYz1Q3Lv2YmGa8a0
7s02AwP5FC3XJ4voaBleVLiMp0PddiWnMWvPfTMsgEa1/zBRENYOfRuo1TY5
E4yg6vYFXggxnsxDWA1BiCvLM/yMvOn4qONAJ//CVSg72iNUwoBu5d82hZNq
OcaCKQN2a94E+TcXLoj70Sdufa5t65o4Uz7YAAKani6pq1p/2izQ2PWEf18Z
8tq+4iSwu0IFSMCWXX+0fENuCRwtYKhTyyknXvK+7UZ7HBwmlD0oLm6nTOGE
+F8ruYQJLx6paZdD3WJOb2n4lceWVjdO9dxnM7WncsymS1Vf7VWiVyRJ9+TL
bZVMad5soxvrC0KRSr8zpqJRdQskcVyCndfAfHnE1hCz3tigTgHc27gh7aKY
DD4wVBAANHJhIp2BNjfQbHqMrihIdBGhvsIFJ28tqjPzI4erPgD3wnCQtZSz
LqaKNaSOQWEWh+oVlA2QSDUwvCra3j5NQIiRJkcLovuqS5kkUcapnaP/4wld
F+6LUp2Nzcy218uAjKt2zDcVPV0FJ06MVDCgB8c9v1rEjid/rHIV36lp1sgx
xfgzgZnYJVRlsPXD30Pz5/MbEI+UNsxceIr76mM9svifkFnOlmkn5CfCZV0s
f2FQDCe9rePd11dodu/3IIKPongWzMU2QLbMe32hLmaJv/7n8uP0jgF2ZOTm
6BU5GghXOJUxTQ/N07hu86oTPZ3KePFI13MTZa13hobty/zybeq3AsWIk6XA
DEJStpONwvd+6fQIZ+gzFQ0AF5OfBXgtDoAeXAAuyQM7VhWByoX5URFOBqTU
k2BQeD9D89a7fquTWBdsKfrZzRTlVWb9s5FAi/EjtNQmDaZkXYmrM6l/evqr
wCAeME4jacRIngvw36r3k//HAdavie1XCXOeebsuFKg6qNlAlVQK0ejcC9VC
sFar4fjBKiQb8ykmCB8Q8Aweqps+djSdeOPDeIIFvqDDUbtCE6/l1uKuMcSx
mB7wl07WDmZqhBy6Rc13ElWOcJxz1o6b3yp8cdg6FF565yZhBguCBA3Uh0w3
VUuY/GeqJ/9PsqKQ5kUbZi/qPH0HWuorZb2H7l/thVEFMNfB9xLg16VrEQH5
hty3H0jDQZNVq4nbluGiRVC07kXiJxWa744y9EAGI7V4ccfCXLd1ssqdsTNe
A+wosmkTen3RNMKIaqxbvxlTxMrJcw4ohVCui7sb3+6KGobdIdz3nHgX8ahX
syCnrgDJFOW9WfdeXRfDbv1t+TboNnYwC3n8RpEFTBc3UGhhiEOcYC9LY6I7
fPW4d/Rcsij7OTvQYiGt+Uu38HDUxeUokiAlM7vLc7YoLDh8NqJpReVqMRmm
A9lLFZxQF3G+sBDBzm6kymAgjgSGD8kqzmZiTHyzcD9byYQo2eAKwKnShKYM
X0pshIpmsQBN7aQ6qLEYn/X/vBH5VT+XsfIwV+fJWK/4MsZLDmLVCCl/6dF1
SbRqM5FYbM/7IiOeznANKBBcaACSFze+3RmKGo7K0lGL7rc4Zp3nMKRsge1D
mkmF5eOllsUZ2tcCCNnvDrzAnfim70UGrmCRC8QpWC4h40TAEriRvPvpRxKq
iZvw33Ho08ZNL4fFmKOYarpHrHAVkEtXVgHcXhCQHjUq0WEQzk1WQRmvykSI
lVVshZBqPxKM34BTtKcXqW60IVfCfvzB8yqSlnjGaOrCuLDkJwVZhamrzfMo
sKoSDVlmJjvTD0NHd+UHEmDs/bsiVDIdsC5Qan5aZgfRIVQEzUn+wl9WoFZd
/k1iSL4DRXlfb0ObxmAV0QTSA4tlJCNgu3x4h4pRzZ7TuzQvW045rAmjqGDq
4CA1i5ja7KWYlfX4RZWcdzNCPVDdD3S8U4pCGXs4H9pMbIcITYQy3zemF21C
Z9qGRcpoajq8h8fAU4HIfrY7NPwiyTYgvX4IrL1mFI8h/cpllbR7Ab8Yj6o1
kFAoak+2w4mdG9P/3OvGQoJhcUnRqRvkVGkznILQuE/W0vnGi/DO0nQKOjKH
YWGP3PrkiPrMu1S9RM/oTmUxDOjcgsz0lwQ5TvRMB+4RWN6etKdOXAmb0QNY
p/oCjD2H1E8gsvUIs4+CvQKjQ6tkl0HJDGJfoPMDPQwjRsJW8PveUinSn31E
D3yjb33tZaNwa83jMG2YjMEvcnSKBPTz8D+xwuzZ7NQgmeOMptw5J09h7Aek
eTLxLrOCg/+rwdOuuJWENoR/Xmn2l6SIeiMDx4Ud+X8qYUo8waxScLtRciGy
vqpfLESU4dG54VleKkxAXu11Zk9DkJIk/ANsX+hx45VWjndibZFT6Kpe8NoQ
BScEokj5zjyxSasLaNLp1FzxFxI7aJPxfZOtLJWvLIiho+mCdV6N/fuquxQW
rZ3hTF8JELJBtqKjTdoBedr7tyk5XM34CZ+unnuXhm4u3BoGRAxOvnjKRCVZ
b2fkEAB/xYFt3bGCY5ObfsvrVX5VpyWZnpZkbqZa8wXPjs1Qne6SMLi+aolD
+hiZgAMbsIOHA9w+HQXmmW6wDs3RofBEKJ/NX6IswF8PErY2GqFhYQB6f5oj
JAYFjGlM3OwUxXogaOvTxgpHNqk2kr8dTnwNbNLSgTFhGjiWzyA6mh8SitrL
L8kvEBAWWn+jeA3djChpZWY2n5lzj90qu2U04kf7o5UsMqKm1e4lvmcQzWvY
UxrTvAR7eY4xVHq7VwfcHXoY3QOT9LQOr+qMeLAziBFGEiFxoD3zcTAKkref
vuTkk3ypGWCokKzPUVjkxzhhUYJ7LaCDzOFdYMsFk5Nuoxe/e8p3jLmhqQZ+
i2ucz4Tz4ce8krN4lu2bcetrMsjY+3Y8oaLGtH64ISmXptG2uWxGle9SpVTV
ocw7oUgyDaQ72ieBXlxhXTPKcQQQq6a1Kkjix+INp8cha/TcLujmYWwy3nTp
w/n9YGR2zp30nyv4mEdWa8lyV1YPqEYxbtJxVP3e/jHMKNet38G2+vf6nSXi
ptJX3Vf5vi2LA5FTyhatOcm8jFYxsEJMBBMLEOy805X09m3YtnlH2zDv9TQe
voVOalOqTpkLqp5VYmkpc3H2ysp1FnwLl2c83siGpl+udLwWx0l5Y1qOJ1NM
WSQPAbcCp3zxKYLCsmR4yj0ZcDXLcNpDHcWYGMjBbaIAYeVX8IVyowTUZj2/
C6fTH98h8wvocA8KSQlWqpEte1eG/pJjyumWnzL8fKy7aj1958Gwe4XM64Jx
OfkXlKATLADyN1RNXpNdtrkXTKmALwcTFI5ck2Wc38YItqW8UV6F+NvLQOl5
fQYWCt7CJH8uQTi46wnjFQmXaQxPrhCqLhPaXmtJX/EOaDoXsVFvvmOtQEQB
xImtkknu106I1MD7fpONjPg3SxuVlsvcJv5naNpDoY7/q55BL3VnwUpqDp06
xDz6ggdb4KzheBv193KEBXY/roQPetruOwNOvE9rG2ivwkM5HVJ4gcIxLvSf
b6diZq3xSEg2tVPmYKjoXUzH9EEDN8ouVD3ly0iXt55WCBBSgJoQMaIu5edF
WAlvVZQBOjV2CG07IdxiBvHvPhMEWTrusrxCLyCTKlyw/37UqxQ+KhxX6Vid
VO6Fw/t4tDLdtulN1pfhv76HCnz0DS6u2aUDIlR3DzEDZlrHGnXAZ55Jk47Z
JT9nZl3jEf8IbCrDJ3iLRgNhNu21bRkQt7tZxZxle+ooryWnyV/JRiRGvi5u
TrpT55EVMhdv4FtDwvZJJ5NqQhgmMckjqS2q/tMZEGbbhnYnNAMb56Kg199O
6PYWY5WWWkj5IPO0AUCcfR/9h+V9rj8Bretk6AMmBAnB01KfbT1SSQ9T0HQk
S+F58fu7ali9CPoWgeWQEOQsSyH6VTFPIDRXOK/yykFnHj4egAMt1t15mtMz
qocM+u6DpmdjP4iSiFKB/OVgHKvDo/lUzHUq9R2PXR1VcOS0Pl5RzNL2Q+5W
jxbQw+fVJppgbNnaLmM7Rb6BDYYok5w3kY+gxRMk6lYnYbQjJNPv8Q0FDmrw
Py1jODcJQXhzDvuh/p4H4Gs2j1H10FrudMVvsEWkF6IkXdT7IIrXP1f8Bmz+
HRgRMziEsAdlrQDw90ieeIrQm2ZFG7NN3PpfEWE371j+FSejXWKUOVM/Ynxd
nMZdfIm/zhGLS/tN4l1hOdU8zaS9nzJAAS7+rS5ug0insPwa0Uh3HuOMGtbU
yvFYf2aWLQxvtU1KKs5+WOxA8utMAEuAWhPc5gkw6HYjyvwAuQby3pRa/KN6
w2Bsz09NR39CtHxw7dg7Z1FbDreXhFYbb/cxJLrRBJqi6hvXa7MeOvvTzxDj
8x7BXcNulpFCG6ZudS6hY8pVshxQETyiTT4Ce1e6GRMUA6nu0tmsy2+gWv4L
fp2V00BAJ1qWi/RdDT51u1CdFl4I3ux4a92RHzYomDRx6GIyegrYkzRg9Av3
akQvbCCUtYj5irtJVR0U/BUX8SVRo4/82uAoctumFOFSGTaxiZ45ndDf1YEW
yDZUnxay/0TFZeHEgCzh0WpkiiI8XYwI5vpeU9kDzmQufqhnPOGuJo91YRdj
rEKCn2gH789hvq52dfFrV+sfiUSVnCd8h9t66tURu1NpKU8TYezV4PBRxU3M
jaTbAUWn5JJXv7O5gT4oXfi+DCgyPjrF0ykiTximVehtVc0aox7kwtMFCpK8
Ne2Fxuvgzb/EyJwySMkH98cKWCdvOpZdLY2vtR94tWTVqxzbB0XkxlH9Mt5Y
lBOAbre+7TlBskvYTx+T8rGhdIHcLQK7VS3egczlJkEUvIp23gxDt/oRVy8W
5DKbzMGS9qnge9+26Bd+6VS/AZhoIBagjm7LaHurUgN7cqC5yst0f2V9ELY5
zKGjo6OpT3Wrd0ZHiFOuRBuR4QW/ENEKrSSEzhlUZq8CfYJ/vLWGMsso39as
6byS4LTUQ9n/ZiOJrGOl63tYquvNfhLPWvmrLBJW8WlBZ0XLYZaOgVZJo+YW
0nGeg4JOWfMDi4/C58MqgA2qu56LQELPNfmIp9fZnB0PAqL+4ksnbZ1CBLfF
CnPoyVPIigdVnZCzQQNpsd4NeythrSLOcRGoNjGFHBtTYOpOeJjOgXDDpK6m
9LQYZN+LiwrwwIMn14/FaZsBJ8kl4uFTOfNydB0vWcKcuHr0sJtJq77QhmOO
5lRAZRcitBWSARM2dwzYONJnKy5/527TSsq+9Iv2i3fpq3iZJpWfErVL2Gl9
cncIP2P4n7NELV0I6oznuKpIgCRg4UtCG+31YkpWXhNIwZN+aJgDVDOMRSyn
JqzHf3whZFFA2AiMCGoLUrGUI92D2mog8VQSNCPCxsdv7F6ls3hRkKKui0Vl
2/wQ/8250750aoWrUuZHjlDSmn67ih0yGRUDIKEqs4cSptLvLcMqyXBmM6y3
Pue9SNKkeMOzdEqBBRuk/CRUEKJ4jh+9NdM+kNFxVl4uOs/yr+nzOotLOebS
VoUevmLIjeJnSatTBDr/1mvqUGHwFe04Kd+H3HNXAXivAFSMohqedzUXNkkC
SAaquAoxj/sYpsrDlR3hO/JlT+tCNvsu6rEcAHUU2cxyguY8W5u4JrTETSd+
w3bk5VDKav2IdRQ4eskZqS79LiSciUI65GF9HHi5u6l/iSSea8FZQkqgiShO
f74XCY80NQdNfXuCB3yB2wL3PfFbVrGO6ZX3/77o2Eufje2LllDtK1+Ztobw
/RgprEYZnIxFpxGS+V6kaeISTWQtRsM+s7q5+ADqfLxNik5sn+vMDSvDHP3p
HWy6CD9TnBBHXvtgBw1L6JrLTBPNMRUBn2rkwS0GFJmqZ8Z8hzw4g2esi+k+
ga3Fad5NPxCWX09VeJfTn+JlEm6aUwPpC8L/SrezPf9CdA2nlQqojxwlGWIF
5P74UIjl1TTKXNGV3dLa7121xadqKLVLvh9WxvO2fZNtKl7forInKUNQcuJC
k+vVsfaQCJehzG1LnNklRTyXwAm5B4kIY5lrR6O9VKHX77siCjtrxdElbAkE
+t/G1HYXWHTfL1mqn4qFI8lSSTMqMXnH6NSwSW36DPJ+3G+BQKszwBzPKYKN
W0loGmG4Kcww6OfD9MPw24Qd2QfXBJjjALIBYP75QPTwnikHm/82+GuF2HWe
tK0B1pNyhRYRxZMVOvnRd+MpcE+HbUArqOG3r6SczGm+y2PbwFxaxanLBmrw
qyKyDSfzLVHq7C1Z1h2/2E+NY4sLkoBc7VJRDYIjBPD4EWzBoRWse0G+9lR6
baiSuCQuo6N1mSQRsNHqIj2i9yDwLtKWshX0LWjMRAvO0pBdj8r1BOj/jvtV
wo/9KIl588FxJxYN7hYsHH1589NAatQ7B8qojCm+A5QclZaJoURdYV/BgV2+
GrMFzpZdmYQvmCvxMczmBU1SuQoJds3rZvBNmvbHPs3kxg2fRtgfc1R4ezuk
Bjvk5j4VkJlyW9vVugHjSrwklZgmHH5RDQjONfrfQE/CIiQJ8aOF0aXFVkwn
DlqYseTFhnVE5aLypnlfMuxDDsCb+zjNPfJxcBeplCTE22bWzwJUMabVc0sY
/32wOlKHRRowESgLOptMfjK4zJVTYT2pS9WyY0/Rv4E+PY7X/1Mb7fLVTUKC
L+jnpU5Pss8CCv3PozyePWI5ewCK7jvZckxcE5skeKhgsBJDfTH89aoT5Ed1
MrYVJD49HQoPmnNPCl93VyJM0KQr4PhAQYEmtF+AjW8DWO910kMSprwaBUA0
Og+MU1hdAZzkTRhgfGjP3KYu5rRU8I+6SOcX1+m10JbinsgQIB4xXv99TIsa
q+CRfkd6ke/S7l75UP/Dh9I7whVp8sF0qHIAoI4xh+pGyUNxNBMQbtb88nBO
kF7rAAv1uHyC1ScmE3TNkeMHcOKz0oiJylJNe5o61PCputWipDxAUEJzRBMV
PQuWfP+B8B4a8HTwoBiu7jMOOfQ4VKMCtOx58I+BMzBjSD7Qcwhth+HTE4f/
fr9ugjMwvSj0O2vgKswjv5QueT2k+dCNYhyOuGX1YqFFT0fv1Su8K3KK/voG
ZNf/ocHicZykvOIZfuWGJC2HaJNSAxHna8i2zWe9tGRyNEkF2s85xxjGVebU
xdr9mw34LtD/ok33/2Dq3gMPbTtjMA/QliuXgMdI5bkUHg1RV4N4Wd2FJmpS
S3J1LwsiDTq3LDXTpu8GXEJfMKS3w7kBQKr4FHY19G/USHLQe+/FwxiRftmn
xl7JPdY0+rFu7+68THb01YIh9yQM4yZalZeuVXmrYXYlwY1cyehV73SAl87N
ut2EHaoOhsz1VNdp4bteMf+8ATqeaYBUB2PPPyBtudr/lpYTqPrMmic8WTjW
FhHMqVInmJhkdaEELn3uidFPIJEvlNAvGCGCoi9jkrZxjg3YEV8HU4qTwFU4
CALOAo4UtIo40lNg2lkhYKwXAMGCS8NHYlb4PuSzQZ5Le3yJCuqtm9vh5/sR
akJx/7hU7B6qWD1XBqvq2S1AQ45L7AkQFy5bQ/yLP99CxDY81MOYN/GqvUZ9
+xVwdv+EE6tKrvnYU/L/FO1Qej9TGXZlL2XSqN/jGczRgb6FqpHBUUUu9eUm
S+pwWVlUWgURvyqCWSm8bNhySvCwaVvWSPPclIlS6KXjoY8j5c2hU3Trwfsy
ezal+M48NyUAXxDgkuEa9McR4zNcRXGCjXx9i/ceg+HEnJmBqDMcqqJ8WP77
X3/O9rdAxK6qOp8GlyYymf80vcj/k3dJmBpdbYMoAi5qoStrlxXXggyF14TC
SYyWJwzIA9ydCSh5X2Pmma+ebPlnHnlN2kdh6trR8UswVb7AA5M7GIJqu9iZ
q5ish7Bvn4gVDr/fY1uxbepZf+4mkTIqQPW1jw/z28bdbUIbtrO25iVDTNbV
RLJySH7prLrlexoYjumbW7u4LmD6JaIYGfTyh1pQbzZzhpwXd9a+oSdtWudD
msMlFVuf4AbbfrG/cjK7/e0Jh369NHN43yJHR0vkypegpWIYn2UlUyKDqwQ4
s2+7BqrMV8oiukNODZ31WFOJaQkVoIiGpVuSOsbJjBDjIGQZph9d4+nC9Tkv
X77rd01QI7v4qgs77q5X9AdmHuQSWnEzTQSX5RtWyETCSmc2NpiYeh/kh0HZ
qH6+ho7h523hA5cdbBq5P1xt2OiNTSBKUSs545PBalY851PFM+uezczkf8Z/
soGycWfFJLuQPxRYKrmaEl6+E5N9SGraWVl6BU02xRPFPiDrgZUoKnS9xM7t
4tDdbDt3SM/F0e/iRMfDMQ/+5aDnhvT8NnvW8CNFOpiLOzZb0jjAi1Eh6JKL
BNRzEZa1FGMKwgHyTBe5w787rI5Myw54VjtX8aIcZvsuyHWnwgETE2Vmb4Ph
lzfPg9Ql6NqPmbrxdRWG/f+PEhEPlyDN6U5UfFm6XtGGZ88f/4A3TCm6I9IB
f21KjSmvix+kgFOe13tj1c2pe3qoGCVUPUcQMKrlJhLdepy69L4mOC+z3AaI
sCQE/mEys1OZUp5tGJi0IKKy7k/WCkVPmdFVILSw7EM9uMHjILq4AInIKrcN
3zZAxNiLodLrpbJ3vXbanPD8AVex0YVb/47+804lnwEvjE5XJqY950ESS96p
J+vKqVJeNkOUxcBAdS3QIF7XQvcg7T9PjrurlTQBYIw2pL9neruatXz8vseM
EwsOC6ljTlHYpADJyC59h1gEz53lZU3/RGopkolvTb+BEWJ6Wo8OfulNIRBx
W5hV/55wR4PhpPPlONYgw1fAjux6SrdQIUhiA9LTzqVH2XFs0/UU9Q3gawl9
cGN33H8AGwKFVMp1HvxnfOkyQQNC/33yxNjEuFZpnHy4BQ3nEo2m7StN6wuD
j+RESVYM4Uko0/UJK8aMQvfv2Q3FcFJr6jqr/5+nfgFKE//i6EfvooUHYkWH
roJvJj9JlXCdZgw8x0UneqsOW5etXUgILirAKqInrYvHrPlbU4PeK2O/VlDw
ZQ2D6VKXa29miKrheqLv4+hzKqwlchSOQB2jEGHpF43GAdQ5HYJcf+rQZCnn
BaFwqCksDmihZkofBcvVO117SciYYWbYsv751DyfLnhKMr8wY8qvC+mb4RZj
YelXbpoMEPxI69k8rYy0n7lE8Jg3isJhH+1ni664t2x14A93tVr5A7XZiiCA
aj4q1P17Bqx+tCj+ag9pY3uJoQbbtGaBdyoIqOCeuJLuKLoyNYZTH46ma3oe
07l+EZagPC6fgOqEftYMPZgaRBl5MLFzuTIH5QTuKM1U/vtuoksyMkPYb7Vt
CodGOuMQ+0LyPTbRDAAP+X/lz/miLCVIk5n9jIy9+rp+cy9QSkDsENu03mts
bDGL64wiwJOtUe23jjHaNlKfVzU5zncaKrIJGzopPQdhGEsv8hPcXkmgTt69
cKL1ewCBo2m8W/aZF2fFTR+aipyx5Op1Va+uLEW3t71EnuGOAKIL5Zc9kam7
/aZ836ytqbuuAOQSM3w+EG4TlxvFF8XYCuWBoNdEYnJ4n963rXBrocFAuzR3
HgPfhKfyRfICnBctOLYtJjnwgckU6qtmmUpNC4SbJpodnGSbzShGlCjBhN4Q
4aU4iy9tXRvIujn++DZgTI3MaELi3N3JCYH3bY9sVDHe5PmJ/HZjl3CWXdzU
oKcm51cUf1E30fkMr/ParQKVjusqUKiOkQ9AhcwVwWadEqGJnGiz9n/jju1+
hp43oYlfjNo3HZtIZVIBc5aulxWRCb/igQZVvxB1Y7LYIXKw4zK/mGlIhowH
95F/NN8wphZY5pPMGUPINw1L1uAVPhZOo37nus/WJ4k17ssduKUt7ho0E6Rx
NlHt5d6c2d4fzT/fWhhHLkB0/J3WYCpWSN05JPll63uIeAfPtNqJIaVWO5sQ
ncP+sMD+0UshG6dblWfHKJIP5aM71DJ8bCKvnhteSWDLP59tPlI53QbV3XEC
coPyLzdN67PgDDDql5wVWgDcXI70twM8YhlOxE3PXGpZ1KMiuWPFkS3bKhIM
eUp/2ppRr8ihkkYZyZOXI2fV8YkwI6toNzN+F1BLygC/0zPVsDzZMqBXK8Fd
aQnKjR53yYRuHoGI3tra/XmRjaugI8cutBuj/RRmKV8mcElhaONBSpsLiSOC
JwiyfD2jfJqvOrBBNaAt8bHnJnxbkp3ar/3R30tp1Qo8iIvm3q9SVI0yctaH
N3bmN4J2GYXabbXqCy2k0C+8fB6c85zx0KLgMh8/VqNCezMH+Ey9cfU8Ae5/
MalWjaM2E+aEXRlOMp+Kk/kRtvHYCcf5hftH8dmaGMPKx1w2zHKBPlAUXzXO
vPex8ed89QP4q60DiK7nxZ/RIIyFk75e7N5Cq5mYlrTCcXGQqEjWikVHS36O
eMJRxm8figJRutCGIrPTEejaTNWnXuhI43otrI4KbsoQxuC2lKyS05N2zCpC
dbQzijKIuHsFpQGJIovpDnpZI05XSYNbb1D3Drem6y+BdQ+WZuoKsobkpt5k
qJ07ziS9nWvmRYsDD+t57RjjKlviDufT2jlztMvXQAmF3GAGs6gSE5meKCHk
DuPf7G/EEfYn1/GQt9zpxpSHHctA5rU/UWC/Awc9h8dVyYcFAgB/4s5Y7fvQ
axajSJ8+wOMg903qFpBuajdy+XUBfEImKNYGuOUxTiLFjuBLcX6f1BcRfR0G
ImfUJuH8fmQLkIJKrIHDg9CnJsdxGFDuWsZ8KVJJJybPxmzm8iSwpdsuK+FJ
9030Yz1RTq9mGXAmQEGU3GeIVfidCNxriQYtMPYujnP/ZfpCKkyT9+U+RqgE
kJ4dnlpx1zhRIV38TkJeJm5Vscq9rNy19xRk6YjZ2AGEx4z0MuW+lTkXwQhV
76t9B7YdRkPYsOmuJIFzH1efKEUthKFXjP9lQk3Q83y0Dc67K6vbfHCwUG8i
zTABqZSOdzqa9AVsAlhtHWV7Cdswf8Z+6cpG2F6ZVz5X+WA0F2qe0VfAjWPO
1CP6609SgednfOHUCLtYcKGY64ZdIT8ElrZZqZ1eEQc9zUx8fxRP9O9pE8ut
kmMNQWL5s4321XWYS3kiqJMjKNLgiQ4+A4B3UPbQRJcGneFxATIyWfYK7KYb
TP2x9FitZ0w9SCljUVrxXoCMw0GLlqKYjJmdu1+eY3jxZO71c8bQWmh39F/C
9GfVn8T9zhemeoTALl8f0ZZLPfTMvzaCZtBjBd2GetV4JeEAMAfpVRA377ju
x9c72QHDQ/mXAwGKzLTpQubVrZp3CFPm56NkWB/GO2BJG8SQVwiiZekAdc9H
1FPZ1wX+CA1CwqRsNP0jzA1O4dWw3NH/0xHaeXtgvjfIXpxqfP2f7t+91st+
u38qGlJjbD8bfrSyT8cfo9C9PtLM2CDDnGkFBuyBr+yAaNt5nkvOOM1fR7AU
54yiZPwobl7tsFlteywhwx9faGVMpr0UCgoZnCIJ1eNh1EWrmyqvLB9bOGyK
+fa/1BjzHihW8cGA49bBtw/0cNKSDuv5OGEaBXf+GGO6K8ktetU2CpUqwijL
kInkpIPiiI3OWcPgSCb7r3cKvsXsvUcAGtwNogpWrgcTXpKvQulEou1IifcJ
qTjMYm/RaLdLSe4ASBnG4/sKwb+/bXmdcNdUyZRiRR+qZRSfQppK9IX4ovzz
lC+mm3u1TkrwFuZAqbUirQrW7tc59Idd77u+gKTJxIWyunHrOvX5t2gYQ1Bp
31bpslYkE1nQeEeAQ97J0ZOb7BwezR3wyuL0j2F88iKVypl1qcN9BFSE741w
aWs0XjflDmK+582EeXpCYTdG+fuMdGzdXCl4jk9t7l6rSB2J1xQ0OLaOFHW3
37pKPUdpMxAzyYsCnRCNoEN3rXfQepf82+MsBUVTFZ1/cj+EhW3mEeqGTdF4
BrsLy23B5O8vu86yqVBJwB9+4/iUq3SXBOhVXA0YW3uf/4H1oP0BKwis0w7H
uRZI5ZJF59SO1sOdgenzSiVuOuarOdDGdvIizhgNTlKj+7q2d56Gn7v6QBBe
+tW8FWw7M1efZZUs6r7g9kkKZR9ZLlj00bTIT23QccQt/ZURCsePBeHCtW36
w5ow3oUdkwTqYwS7xPcxwOjp93AVHEPrurQBWoAJw/4shjsG5Pcs9FwlmCeq
96MU2svmCbFJzeEKKcQ2vknZiqVUG1BrkivLYOL37w0CdHctUej8HXf25pIA
AjXNXQHalJVytyGvfhouqrbiHypqrudjyPsFUJw97UzkEEq5BUstxh88PdaI
E59QD63tz3xrBs8gNWXklc9Ef7aH8cc0wAMRl15+tfNmI95HEvXSrfuqQ5Rt
EQOfLIXzoxLWnOE+U457egL86NUVh8Y6EwAI+qZeMmrHkCqzyYGg92uCQafQ
Oc70vlhlliNpG8c55cUGFflUMIP61wLG7YCHG62fpQTM++CdZRCmXB98AK1b
jMITurXhhXHwi1VCZEGdpKvB9RBivK9NV+aE6BktjjSz7qPNe+DCxezAcpuc
1F+VvNqdBVlxBzrXcsce0ntDVBm/9gNfGf5/EZC9hv7WxpOWwdTm1dAaQTy7
ZxOvWhrQN9QwTY7oxA0g+THy0zZ1PLwPZlYixyb5JsUPxaDHOwIcPYXDs1JT
eG1lZZf3T/BdJ3f3kmElhRuSaas6XWcpbX7YiPK0TPe2C0j1YxR6IcHMhlsP
m5CyyaqEnco6cSGePkdVjD7T/NHjtsiTiT3wOF83HLAi02qarRwwfijLgDcC
NfJ0uvxNNaK8MM4Bv8/U0HM/9Mh/zf8eBL/2mSg763m026uRTL6CtKgCyfbI
tSJ7BPz5GtEeUlMORbtTg83KJlHtNr/8m+1K9l9k3OCdLjl1fsOMr5tOg9xx
V0tgx4uSwSwj8KNhLAJ0d6fAsa2k2eAzX8FT5jOykIvLdj/RkgsfcqDqSFcI
5GW3DT5hdDTgWlUdvNcDpIPeoMrTkA3tB4Wp3ZFzHSXLT1vLnhw/ApFNQXCI
etPpmCjG7j2x4Dyw5frE/m9PP5JqlrXi/+Ji8hp/8V9hbWZG4UPkBVyEavdi
sj+NAEEsGhTqgKmEIdw9JKSDLjQwWZbtrZ6X9kG9er+Bxg1O6SA7hZDfWB3G
TRvaL8fSCCDDmm1X5yx2/Z7bBU9RsnamDCmjhfvmYv5T78sU/iNuj6u69FYU
T0IL6r22WWfsTxQNVbxRyyPyWBOHAsyloEDs2JtXTvnHivJOWWkwFN2RXCLY
mZsDGbgkpRD6K512iqLReBvmiiNf2xvnOtTOX8aEOKBCXt5+AD7fWG6L+0Si
ON9k9nY9QFsAV9WXLMOsEOcO8eLv9gSvY1FxG/igI0DODZwy+Q2q3fPGF8vJ
EB1yjRPtNNkkQuQs9t0u2+/C7vl7Sy3q4KNIEOCLsgbEPK3m75iLo2iz28b5
aXPHN5wfDOCtemOAr6LzhXYiTDQ36XEe9vGOttunDovHrYKgOplS5eo+2TJs
AuHXX/F3vRClb2K1Zf/bLamq7pYTPt43pVhGW5YlYSKNZeYeFriLpHW57kng
U3wIYSWxUPGcUHGhyULjlTfd0nHAyQFq5vlk8DfMBfnXox1PWoi1pwDo3Dup
Tz/m1dAILHGD6+BOJT1/rr8CyevHtlOGaifqCWMPbjKdh5rjqMWiJi1b5ZN6
mUxkgI9gXwoQNbdIPvt6KvYy1UBkuOTRchphIZnzrmKWLwLovusbtRsi5cR+
Ynbnk1HnlsqK3Ci3pL8Aa4JNZwSOe90HSLOrtHsho2yYblSAjd3l2DyrRl15
ZMB06VtPlIuXS4L9ZXuIZWc7KMHCCXCXYMpglZMAIuuVDuSI9wj8gtzwI5Fs
OoUAOJBkgzIAlmJqXAvVjTIe4cylJLJZtPHhVVCKRNpZd9BLt/+1hrDuDt6h
VC4gk10MNB8YiCZ2YC4g4w2Tzq+mgwVipYEDq76ef0Gntye/Q5RKTO9ElQmv
VWXiDcaclJSxwf6y9y7bh0IVBOZujASTd5+yANDwJYGUX0JqteOQd8q7g6qJ
zfGCiuvirRUp/6PkCgVkFQ67J51qvi20Ahe/caKmRTyNzEJrtKdMvsxN9CZ+
8pzym3kuOXuMyL8MEdvDyUZi+9zLI5ooUI5cFeqLbUDaC9/IM4PTRqXhiTma
4W2N3o01kX6cru6WVE082JY7Ov7lZIelWv6dTYiYwgfUjAMNfrlpdzzE9poF
F8SQOnsHo6krhhHIjMHWBlu2onm72a2DyLzg0FpbYGuO+SSigSk/Q8Fvi1nM
YnhGCgNuW491NHQk7sjmW4IpZgyFOoqUjcD7U+ufIs4KGYHhv+D4k8fvnHTC
UOGvYujEm9MfNhfW92/AdcIt4VLKuEtIQH0G0rytpLc7bhmuwacK3miiAtL6
BDSgu4C0xXlHKEVvGG3Vj+vSEeqHSheNsGWZwpgdTpzUlzdwJxAG4GZjhJBx
drDjAjgJUMr4jhnGvsNnnES5RwdtmbTFoLx3LQVqX5/ge9oYN3Q9MgX+yrSl
/Wuhiyb5vSk5FymQrfojMUH+/n1KU6m2rcoiG3+2YfZaxWZIRkJA6w5ijebJ
a15I1o8i+Uub0/zOzf9ZVjQzfHk/HjJD2c+lSLDjc/fBvx9/nVSy0KoxvqxO
2gkCGF+I3GgcHbM9cNlS7PHRDYKAHHHXNJREOsBoWRP1cKuy8JvdYWVQUDls
MTv5qDH/pOjMAMzmoslWYy7u+nxq7LoZ6zxdS683J3DrYS4exWwk8eDcvWeR
EE69MMqM7NtBCH9HOxAskxILPStc0/3AyXHK7tPic/vRPAhKGbkH7F39ouuT
sfULdfDtIwWWnGcnIFx8tYt4TOG+gJi44EdD2XEN0V8tsUTAfxxFY77tAqBs
+N2v3S9B0UXezFQbeBIwwsDhKzFcKzLubYf7HpJuFYV7MZekuvcGg5x2Kkmj
C2NRO8DjJ2Nakgfu//Fu6xeBMlgM6QwHyVAN3/XTV/kiCAkz4eRngKW1dnBD
PW8ow1ND07H4CVCzxD8jMTC1C7IgB68KYqMwYsHO5rroCswZG3jnhLhA+c9u
0udVadu0S8AcXammthAeXUhM+sCMqgRSOaCUd0G04BHmr+0RUBRTHQire+aj
y4MU7cHDZpFCPiOYq+lTP0kmoTYWwqy85ZvdZg6GXBl1yl9eZI3kdxVj25BR
ooMVz9Hhguw97u/a/3Ax/q+prnul8ocp8Dj9Z8xvUFNNQFDJfbZrBPAXLXX2
sT0+bfrR8F4g6P99J/VoGhxaU7jAZELvUPa1Wmb6gWHTTAsTRuVdbZQEcf8F
nvX8/1vWAhbaM4iRhHumgfoEYu9yHQl51FttE0G52JLDXSnwFraqFzR5eDg8
6sTdmUt5UfWpVtnjNJpgTwD3XDLWlfTcv8Ra/HwXb7pFzCAPNfganNFY9/RH
KgfbjD2rNaWfi6FJRPdWIY2pg9SUOFRcjAJ2WXBejXD+dIc9BpCO/JNTjKdf
GFHnzxb3M5iZNcCdKugLQ40Wy54cHwdj0KQSYQAavIQGZ290EgIis3TEWvq5
RPKnsuLlv2DLB+eL6ifRWpcf9zmALhUuqIOmsMACHK659XPnXER7/r/vWsdc
AVh2JWU1+Y5SS2vGZKs5T+btCvJ/UUVPg5+hmXu2r6OZkFtePAwGfPbDwLNC
SMW0mAclXilFJkr6Epeilgks/nPDh4QCLUyeBSzeOUwLTZOh5X30RJ2MaI0V
lkPhH4vdrbWz3Jkg/S1OQ8eLdKVuaXuQMWwOlBG/PANGTuO6cRQj3vapUvUl
DnOFvyeqLBdMJXOllAYjwNHH5mBVSiwBXvQdOM1Ru6Zc8/6hMrFR5NAVKLlk
8qlyRCQL3uuZM5g+eu9yq6IO70fqQlQFl7+1Y43qEMveMhAfowp2c6X9gZNw
aL0KAKZYMdV7B4+rX29RCHOxmD3PI1fDWAplnVEnKYDfXvKirmKKqAy7Y1AP
lUHmKSyZlXszyOYxlIrCufmVtVsutYFSzbKbAiRq7NOCUhOoHYxrMNMFFbuQ
aVouSXn9nXnoJK0EbKuaS0Sbx+/Fqd5jxR4lRJqtb5i+UGUH+gKjNMZd3edU
54i0wB5R5PWZu4ZFetICjhuWHvgoHES7or5WgOCRhdT0fa8EZujJgHO+V/g0
nTH0ptq1CZ3VAKnGA7YqP18mTeuin+2wlR4vP8b8SkShc3wgJ/MnsS63aDub
dKukihBnNoey/rfGVW549t4mX5IhfDEp0Tjc6Ksr425hiI3a32DkhGHJ440R
tFfzTBRcpk+E186ofwxyor1NwDYWwqy89qrCS+L8kSY7PwLs+asQh/ppQFOX
rXHgS5noVWnjamKdVbrmFeMEIQehDSmHRkxqJX+3RgFGARHf80vqRieTMiU9
LZ5Li07ze9BawgnMA9b0+SDJS4VVnxyiCLsN1Md9NqFcAfc499omI1MymTy9
Cnx+6v6kLK7JUoWIE/RjZOCCWRFepFb2JMCLun1W0i+dNIOrPDvxkfaDG06w
u3m3rZljF3aBEOaoMdEe7Fm4uZPOyAHzUEHqP9BBRZfiy+u3X7hcncidNuaW
LM0lqftCJu92npstwElYlWEnta8N93JRPfyNzGXs6EWCerx6dP/eVHVKnAVd
gvvv6QlWyo+wSs/eB0UYqKrg3wXHxWCNCYCELZWCNHO/a5H42IAD4bKAi+ed
Gxxbz73n2WNtUmmIjmCQWpZfaaDcOQ/3yqupU4VkwaPcMOc5hs79P6Fq0K3Q
9zI6gtiX0VAlEOrzwfMwouHjllvRrdr/RD3wcP+ynr29LX/keELaiCUPbPie
B3d4tCnq2sHLqEl+jtEkd06qeNdWatsBH027jRIsRKZezg4omdGWr/KcrM3D
x5oe/LHZTtAx9b9lhptrJReyFTcsc2ZoIrUrcJRche1PM9t/mD+MQECtwd6x
cUq6SRgKDWaoKoTewB5oazb1+O8Cj2QSMKOwn/++gqERMmrNP3aZz9YYNqff
aW3s4XboiqBOw47smkQqubkTVIxRu5kxiAcBdzz0fI24MYS1WUdlPMRCwC4y
omNZTzrPdHO7Y+QFe8teDBy1GM1wfihOyt0iMnfUCIyLTME3IfrhrbWm+fJk
SX9nGVK03QzHAaeukaaOeeH+FsJjKsjYULni+KVODPLw+VoPll9p0Kwqe/5d
eMujXNHWfUsK8wPfisZRy/c4qKd8jow63Luy9Kzi+EupXfnQNQFYzJ0BACMW
r2noNSAitsFuJ/VEEEKYgA0TnIsNjsafmPmB2i92e2DgjWynD9zsI5HaSHOi
326MTKOghggDk9+FxvNFuYyyilI0hEpWP2iiSc7+EQzbL06FzgMU7dLze9AU
RIq5z/RY+ta8P0f8FFPOPOdtvd+k+qFsQQgWHX95vvxIf/wSld5FcJxtDzO1
zkjZSRqkHMenqupQ4Lp1XQ1xhzICeO26hwiHWU4eHMOlM+fYHQmPjIBra4tb
tY4qUvGS5Orbf3LvkwsKRKZNC1Q2XHBckp7uwxklYtJjjWDTKx/7n+ltffGV
p0QEGrO7ZTdo/jUnm36cRNdlVwHGBx3tZZkU/SVSIT7P4nIYD5H/JXvqLepu
JJJGNqDOeyNZDhS9eH/u69hsLsFzZ66tBqXcUhZN3g1wQbYVsrnlc52/8J19
Z07JNuJ+TE9NnrYkPhpCbrZDeSCe97hDcMxIcc4dhWblmiTP1SbJpeLHe5lU
WKLluZ1JsTmovE0Eb1EuZXTkyEv6beFvUgPYn7VV7WZPSjv4n0QeQ0r9piYc
Vrbc/b28uMsD/BRTk0a7OpKZVMEc4xxqjJlRD33GEK8q00vIYFLdVEgiaLHA
KrrXA1X7ACSSjXKebGitG1rn4M2Q8IIqG9j7RTmts6s4VKyaFe5gpHfKcZ6r
6LDUXYWBWOV33cq6S+5p830XmAU1MT9oWIzACqgoFv8xx6El9rFlqm8TZ1fA
hFsfSUoWkp4Z2+9RL9KagTu31kPlHYPRyYzAsbrGUVZrR34HLk2xMaoPzwUA
OqTggskP1E5w0QsMPxdamCTJ+Yf7BT6LcKwJ2VNGYZxwDkAuiUX7c/Mh5YXf
TDm5+Q9uBCSjIH+1h09xjcfB25aLfrQvTKfqusY7PAoJOxEZmGuVaUDvAYuL
ilTpOgprpCWFE+/vkTBibB9Ed5q4xVgPaHCVVig03cn7J2lPWRFAQ7x7fDCE
jN7yM6kaBevqLKitcqpPF55SWYZZGsi0G89uWuzvjbir4KWlCnmdLcHPU8EI
InHN2qp7UBcLGr0idqKmIb0tdyhxGWCFJQ53p0I/W9BM+lcVgN2xEOSsUQ3H
dDoUhVKfhzKK0KK6f4Hf7+JjeJ0hObidZLEw4hGAQrxV1UIJvo+BaLtbVB5b
N3ebv7FDQNL4Jr7vIaKyb1oUyyIjnLrzRCY6pCLfCMSGd4APqFbvo51RxooU
u2GuxmG7YX8wQ6h0e3Ib1D176CbPfzS2y/2IhI/loOor0vCwkEtLEASAidS3
4vaGhTYDO6uPfv0wNebJhNsQeWJDeB6vPMdwrmKpSdEGwQnnBWbcndaEVdeG
5fSGHwD9AXkFh6MaMpJEI6YpzApabLzfM4HWi8DcP/r7BCHVhSoWevjDI+5x
buLfvjH4EfZEYF6mQoSEkI5YQnk93jMrk2tdHrCs+iMhNicYWvKcinuuZNjz
HntC7ART1QJrbqOZHTaDKmf5iUdM9Y72dRSkraKAfUMGFVWUaIZm0O9CZPGE
r1RZORamRJ3gttxMMnNLjGW8vm/RI+CkbaL6VS3+2Me8l0x4L4l/a0aIO4z9
LBHZgbrWeo338WBWACvT30/LVbMuD0xZx1z2fR0rRoK/l+F00emtUP+P+/9z
lOVhXFjEOOm4+oLifBcLlGQFQthmxn64QAhjBKJ9nuKoR+MOQULQKMT7wNs9
5mC24XJU7UEBsqnLbdUvFDhFb80KVX8pdDsuI+GhplQJDSsOjt3oEGdyDSlV
Q/RydvpglCvPgimtKrgDUrqYdL/wnonPaO4+YKUU9TqEteOjliKfy8kyrJRX
DHF9lfrqEkTrRnuMjAfD4oL5J/zmxqBkZQmQjnCeEBTCHdujRhhoiHNY3rJW
Ynb63MAywdCSCNX+XcwVlPX39Ps1BS4BNbUOjKENmqlrOXd0CI4qugOirRCP
LeartF9ZYj0i6EExBBalnBXDgFIhsiSJnwfGyvBJyyiwo3HN+NuRRHHyqqoS
fbFvth52XDbPXmQaZv3mYYG+zTPNs2BI6nIvepDV3dG7Z8ftm/ueXm2H2fZp
8EbgKuzQaDCFpptH1aQm0lNHnPttvXThceUJog2PdP1apz4gAGXMQNKYGMpM
QPvgXJUzr31PW7Q21s6Ky+XbKvJ9cEsRdJ/Y5WU7HT+6aZiArzapxOxlD8Va
nb2RCxIQFQT1Wjt0J45Q+qVcD+JWb16P/bxdbvSfC0ri4iqzQ8CGOvcT87sC
bQSERFSImNcDaFtl3eaVey49Fna+l9nuiyL9JeBt1XOzOTCkL81M9M88q4+a
nEbuVcLTq1VKGyNDPxI2k/rKsZyPSGpwryS9FmrUq34+yar8rQFrNsnCSFoz
jOeIreZcowuJLZ0HOO0sLfl6s4CzAYgDqEoCw9yNl/ZGlqurmWRkqGX1zaEq
Eq2yZq563ZZicxUn4UXuWCdyOJQdnSdUDtglGpTy6XSxziWzIDsuBLH6KMeQ
v/S52iMllXLq4i1QN3GuregzGS90hvGt5GdE4YX6JJ5khoBuLW6xEFNw0xgZ
A8xAGpj/1+o3dg8uOGsGGTtB8w60VY/jHHYbmuGq67ri6Lvg/mgb5BX8OwII
ZNrObskBjbWsKJWu0ItuWZINsYLBocs9WYfcTbXjuRWiZCwt6FLn0spUe3xf
rbzAjSU7qnwCFpmqjjeAvhblWBMl8tGyCD9KxgjCQI2eni0+1yx3nzhLdc2d
/EpW7vOTnIf1YNLewywP5LfmMQrJH55w6x0PSlDZreCDbNs/EDiH/njP1cTd
/0701E2Qn7N1pcro88f2h105a048DrPC7b5by4LSIFTVN3a6/M22SxndKC6k
cVn4Wotw36+wUDju64R5DlYITZaqUGiPwMQTN5vILSovyvURG2cM54scOdEV
NGOAq1kHgpW5rUYx2plC9QoEkC2/xBDqHvA3zaRz7KkXKUcEYkn/k464a+Xh
+mLHVAA6FHQjTwVLFUqoE33Rkg2h5jt2KPYW8Hjvct0ppE+KFNVKcniORLnV
mi4N0m+UGfxAwmRSHLUS8nDmdbDLKRry90y1pg6JsfdgA63U9uYD+KVv07Q+
PEJ3XBYniCHnXuupKgJEtNH0/Rlhwm9j5ztm8sTF5nkeQ7g09vEtJRJGpa3A
QEJ811Pm1Ly0SeAK37gPyXGHCFTLObskyCf7FL/+qvgBRnept7wiZvTj6R+I
JkgOyNUX7BVx2C94CfZYuEfIEp2smpNkxhxL9U/3H8iYQso26BwQamjlsLpI
UD+L30YhUMuIPiYEVqUrZtcWIhhnbYuTwV+ZH2IrQXDsNoFGxCZh8um3HuBN
UUmo5EyCI/yiORwUm/ppv72vA3piuIK7kkR+9g4vIjkHXVp+r+cruAu6UyzD
KMOsIyPuxe9LJYrtdtTMeE8MHKJg+fxM+l4hlfoMv+5PzpqGcbRZQ6YqGnmm
zhg+8MJxLsXg57Kz1Pw1ReXVKjOmOUEvcC+r5fq5gUoK8YvmuuvDJzw6fNBf
I98aE5KY5hTgEHVAACFnf1u//TLgqQagxqDVu2IBTDb5SOqGoKwvV/XoTN/J
jIHyorYQMbohQnqsOdQ9dVvGfSbqFP0GrvsYBCj9YXH6AHlCkwloSz/VYMSC
DUrs9ea+WHL2uU5tF9JF/8PgdPwlTW8cRZ2psqAuzdHOw+imWO4mCnFukf3L
olfMJ9xcz0Dn6SGv9dyaQvtZD5T8RNjSJio72Y4+/pmGoKDXN+u0XUk9StAP
18EDBDdAZtT6tNqRsaAi0dao3yifmlZgzT45HjGcl6Tg/2D/fCgx+adWhwmE
ZyXD1ToqUj/TKfaID+bs4nghawzaccjFuo+5FWrnSNwAEOQVMIoRAPdIIGmv
V4Z2jrs5VKlIl+j9dKakCVA+N0gUIsVrEdQre0THtqa0LqKp/r+MioXAH8Pf
35qSXYg+2b1+Bx72jaEjynQR8XA/WhQ1iUvUvAnUWi/ybGu3YcgkyFegjeK0
vjNy4Ra2gvwdcbwvVUoUYvrQaa4q7UXmeoCR2e+loGSopRVTWC5fzZsodfEn
VBHMeAmQp9noi5leD6l3sgI0+YVrU9eirPEnpHv+d4YjPsjAMAnlsogvo+aZ
O8XrDWahbtOeqYaZukVH7cTpEzhsS7FG+bWM/rVZ+t8DQ+CLPASCCH4Fm12d
iHSqrNbfGi8c7l9T5W3z7s9dEUOBuzBbez6iCV8WRBhDK3jkCzzU35iJUDPs
vVWUiYNx1G/zvd81DGWObgJP19bSqcmdW4+qqBjdH5fpG3VyPwOZ8duGHhHA
S5CSIH5dLiB+hhNLYzZV3zfy1DiTUzu5z+fK4QBJ9iFdTyYl0R9Lne96f68x
tQorfhEaOwWIHCKRtULGnVQ9nUoe7iAqIK5mYHxfrGfW5Iip4eTmE+b7V69S
pH0+9475QMBrfePnOYYsGvx+RpRHcqwTEi/sYAlLx9+Jx1mhfHuZDmigkeFr
KCsVefywg5+x1WzB68om4KSQd6leimIN18NloOHq5sZ8LMDkwxKdegaclbh/
JkQPmRY+3sVnjyJKp8wAmFVdjXdEgksXxxs20wchWcePpqQHREusxJMyeAc2
p5Fe4OzOUlHARtE2M1edYuxJgy1r5UG6MwJE4Tf9/Q+mTtujZ0+4MF4jlzBc
u5DKIDn9HgAHvUEdjsitwp7QmW070b3jeZGipHZziBW1axp/c5pFAuBW9LzM
z5OUWsoj39ZEeY0DNiTyUarWV9LPHWvHPPa+AOdTSzHFTpwrEHunWP07zRQx
+Fini9mqTpgD4DzcnLJHHzN/1nDi/g4sg5GaDPX+r4gSL4qJlqdyqn7qLH1I
fEOibPT2l8bZOJzm8s0FDXotwLmmvyo3CTrtKfT7XMK0PwpZ3D1yvSXhhVJZ
s7lcAeN35EvdQyDGuAwt4I2ERZh0QXGd5jgrCXFQIidNAp3PziPRftGt56+3
s3H2tzoZaxlLoBW8+IKJr78rL3EhAWDkHiWjaWhhTIf0pfi62yDqI/Ki4TD+
VDtVhMn6N4j/hhELK/qjjyvslMP8D7Mbw7MX5rFaPf4pJ0y6mZdf9C17oqDQ
fvBnqZs7ZmH0GWHDtIJULCsJjk/clujQSv78nsHFhxKXSsZ4IV7lwhEVrfB/
gwpdXEqAnjOft5sQHqaCjId6pXPmY8idkRE7hG2LW9fk7QBihGwwIIgb6ntl
h7jUh+Jm0jJK0mvZJBg68YOWksqXg6ooxo9AveTGUy+/8B6K9Wo2k6GS/cnf
LGwGnVQt2vasUynYCuHtXbOPoc9LBkkfxgnnndbBqydx7SZJeR7pCdNfAPiS
HLWeifIIsglPyvsA9VjdQju8gTWoEgtZ2xvgLyQcFSi/B3Iy0PTYcyXLgiO/
Cs3gbwvTidj+C1XLYy2w8uIjQUF6UlmVcSdDNXB815WXiMKtuTbZLG0L5TjL
jX49oL8EhyjezqdzMjxnaQN+W5vO8ud/v7ColPQ3Kou5tWPAZIlqWn04IXyH
82ZqQk0iySZd/tDDHRfcs2ozps9+xvQfNfV2FESiUIDauQOGFitsXU2k9mmM
Kqu7W4xJXJSgjbLb8fC6XrpDSyxjPamjEj8bVqp9VrgtoeciTuPwQIgO9mKS
MCz5ta+C53kg9SJ2f7F6j6clHrWNQ2pqAThsQKSSm6I7LBL+XWXOsTwwmDoo
Va51zYj0gsLMOSjvgG+C36UxQJ/XHTIcaQd4RvmuZaC/eJxpTQUTRXvauRUb
UneVf7GZW5DHkVsutN5E4lK2PUBFXDMtfc80wyiMrl27KqRtRYUqUPRdX2Uy
3AtxrXkp41v6aLKJStbARcCYx9O9tvwTDWXoK5WUJcpeSUnUtaLRLDDLvCVS
fenMUelopNd7dMErorF9Cpc+52UyfMSA1Q4WjjsX042CiE6GWcu5vm0XYkU5
JlkCLt0i9uYHaPVsEK3/UPBt7Mycy2bnJlVV/ZiSNJm8H2VpBaJkJ/QfEpGY
Zdi8PXNUnR+YcLeZh3Zvw37IbRarejteZLqWIvpF/l/Aoe2dhKnUoTs94wU0
lzkcSgXXk54WGmr42XjB4zgMl4Jq6ilxp29AAQG9uZzvLbMb+pZmr2uFR4Sp
HjmnvO7+IuuRLYuLsI244WuH9Lzvd2/laFwGXI2ScM5a9VWESjgI5Dod38fa
TKIUAVkAXPbAZxaVGYUVkOtItZylhGm1BgdzuqHM5cynEC56sRo8hgqLKeDL
gvgmrLORlIU44PImqEfVE1TBK70v22/e/FEHzs6Wj1eEU7mcOCIHxXqqdMFi
itgavaZ5PX1x4zKWRnv23OiLo7oy7M2JN5AetManLzX/MomTcJFyCy1VOaWj
OnqUANAC9yECmFbiVBTVWmhwAOqoY1Rr3o+YgBHzyEAGUVbacNcx8brN9rEB
15AdaaIQm+4ESet3Qa68/PdavIwjdWoi7dTQRL2gFzT0PUOSey6FU5izWLsY
GNHcTKnfsTLhF22OtwbAdpNtKhMDo5tWyICmDhNxeN6SRzWrlYKe1PHIgpvM
5/71IRv2deLEsNTAdm94kjS/filrvLxr0XpK8OwE0zpm3SZomoeyobLeG5Au
S2lgPRPGnFhaoDk36ExFY1Vgvbc/FZzuBHdLj/xF8ej5WvW1FwXIDjSF1vuo
YCwM3W1usuYo56chiTeUaui5LEWUsDjVGk8Ktq2ICxeqS+9jdVdOuJCAmQkx
vuGTeVVeRpI4pCgTQ/zsR0Zs9muUl/d1azXhlcL1ToyqdhUeaEQYpSjnCbnC
9wXTjUgDe9kHdxS6cpu4L+XJkGy5mUbJ0uqtEBFVw0VZHEiZ11bblRH8htm/
S+eQlCJv+DVrNchIjUK85L1z7k9GuTEpv4qkc2A71nwdfMklUOpqrVZpTJDL
YJmd5MTUs2jNiC6ih2rxh2VmA5yXmPkAvhI/WDb+v99yMCTKAF5bT6IXG2qS
pqu83gBMzS1ywLdxNB9CXB2W9bQHzsNZgC6hFj8+9X4ngUo0OEY5snDbb11T
se7CFVdRQK3rbZxyUvczIoKwmya5z28wIdFDu+MbpYRKJqX16lfuTkn6Xuhq
6rlB1swKKhtLU+mhsLr5J+NfFlEBlOUOvDdhJKRX6+RQMdSXty4naKjZklpS
AL1zYrVcM8+a9TPzdaezKtJ0bZG5rSpyvLIoMhZqZ3zIYbZiUOxyzSKP1fgp
Wi+Q7REIs0fvi8QlkoWjz/PitgJUpZssSYGectPOZmdSlgJQJrtHMBgTxb1k
Vt52QtEawDGwldg1n/9upo6LWV/hJi+kQy8IeeRtR5b/jN/rB+WngWFgCnIi
i/r4Q++Yrw+pU5xi+msNxBYnlCdTKqOuR0VZOxpxGWL8A3xf77yfqLeqkp1g
AEaY5kFVYYjGjIVcrX/r81bdYZVYWHJUoziqp0MvzkCAa2STHvrDfTKOU9pB
e16kTnMZJm+7ZO2/MCyrpnH86aF32FPiidDAfqYTBKJjSG3SiBjOjxetDmaD
cDNm/QBxUi/uwvEBjL5jvb089s0lcSrjzNbz/6A/Vf3v/TADNvIn+CwTEKRm
81+3drexE5z2tABcdDXj9koA3A1lbVtFW7JjbI2D8jXeODDXY0boMICGq6Vp
IJCweqm2EI2yRuJd5cIxEA4aZWJHBs/1bf/xyqN2MM3AS/VY4ynuPW+XNSkt
XOV2AsqbJl299PLs9RvuTLvKDHNsr5u7NlrA0yVBrpTT3VuLstqeKU4QLE1A
56mXOFbjHG7Dhq+QWgcTOoOCTe9GZQGvY8SmaKAH+D8mf/6C1ueHU9CQ8ZS7
aSPNo/FI1bUz6IWfH1YtUqPAFmZb47ZWlO4WEBPw36a5TWhf+IbV52UQnT/U
Fz2L6201EYRF4QsM7U69cBeFzDwk9Dy5iAaDXR1RsR/UDZ5pDt5EBc+J4urs
gxTDaRx9f1fJJ/E6CnB1Z9R5yirmaPVruopy+MErCzCGt9UuRJQHLvtAi1+a
E1tBxq0j+B0SzwL9d66m6PfOgULUdNWqZgFlg9o5z89oGE7ZxZvO48qlMX00
t3+FnUw2gYV699fCIt1ZuQVKyBmGJ44IO7gmLu1/Y2XiEIMzIMhuukCQAS++
t4qmBp27QHr+GJER2rTUu7XxJJERS5Pyacrg9Sj6owNmx1OAl8AXgLwnnRvM
Dkxzw38C+yQ5c0m8SNAVyUmqp8iOkLW659rqqXxto4tsDvUEfWmlyyjt7hbM
zmH5obn+8gGeRAIs6aI6jdb7J7+VmdUcUkNRDYfQDXzCCUikdtn5IjWxWte5
/SJvi0CH3pwFtvliwnZYDfWsB3tk+kvzWtXc4qWez6eQrPfYbFmVk4Gh82Xn
9qHV+U3SmM9TWNGBonJs9NAKavc15axa+QFQ0ccVbBMg1u/F1ybXxv7xcvSu
1CcyoGrFiV1kmmI1JIO+0Jp+7ih87fyW2HR/XlyoWlAWtuI9FjSVEn3ViSS6
q4BdReZPbQkDRtuDVKryV2OLO05KyRCPlsEr+RrVYqBl1pQ41wvtKcS1Zfcy
oYoA298ln1JqaDkwN1LxTfD7p6s3UlqlJMznwXeJuUROQTRX/r50pf1cZkpg
WBrYMopZ8eONZqI9mg9oBN/aCUk6cTwGOzHnUhNCdwbMAvCrPlNpVYrQbm8e
ZPOriX1itiwNdKytkmvX3tzry3PUVyPE55BezKbXlpYE5im/2KE/JEtVjH9U
y0hX/3v5yfzsDO3e5vtN/8AlUsucShQ80zUCzCy1k7O1wVH1WIkfrSYAk2Bx
EJ4l3sdvYdH3xlq/AJYq8ub/g0QK6lOw3NVw9MbJf7MJd6hjDakvTfXIP7Gd
VHvRqVqFyG1yN6ktJxGfm65ZM7K0kl567d/J3C6KfE9l6fCexOEMEqI9DjBL
Msesq9zyd0vDcGm7bcTNHRbPmAUjLHQEAPaXj5P8ciaTxPTevvtkC1OnvFTX
Pju8JEEHn9OswiibmuqcHAr9XFaYG8lVX3ro/r4GZ531REcTueMowOl40HJu
M8k3mX+MNgeXny91EZwycEpgpXW0WLqZUy9mofJ2bPxzqp8orhrOX+nLEDvZ
ZYDSybClFtruSuSQVlVJDj7nTJ7J2gmlSuCHmyYSafeYcyJoTNn9HRAkrxpb
Rae78KH5vbi5rpHWMljBcRRszX3pvvSqnA0KWwegpfyB4XzOZAdsP79Wr6S6
By9PjB2VwsaPyDQ4KSARiCS9WHhHolS6ACwjE/RXs4fUlhwJaHN5sztL5QiW
DXGH18BA5HMSlf820YiVYj6rP+ouaSXDGhMzp+7v/KeZ36rp4uCJ1KmYJVkf
H8RTO8jbhqIkRK1vUiRQJat+2NZXUeiveX9uCTwyVi1I7sCtFENonqFTIPwE
fNgO8LwazPQp0sRcC+Hp/IXhA/bTS1HYI6C3V/0fDdQp1ep2EnzmxdxH27ZS
dQsvYaJnL0c7LoJ3ab+u79i/QG3m6ALPJHm/uW1x8otEaOlyxioxPTja7Qqe
YUHqg58sNiNMCTwkz/zDMBHO5mtZ8J8+TAD5XjmBGBUCvHbhkOSXitKWJy+L
PLpgbHobz8+kmoqZpCavpuShndYRMem4gZHrJheKoLavHz9lQbl2P4OdPerg
Wk6VRGISnkn6oHK75qMY5jsNHYDhsdf2PbQw1labJ5m2J4DR3AfjKoaMvF7e
5Dv2uNiGw0whneEkmArIVJMAmlxlw/wdOP3E1YEoYh4YiALWl+xdbgPzly2E
WCsSFOZfkT3CVG6Lf+cFywBIULJW2Ki5zpMdTFBRbPzkRtnZBFdC5BEyCzNJ
8Mxno4NKTUYN71EcfEzykQmt6xWTAgaMDqeVpISfKyL6QB3M1n8wFkkUJ1jb
JWuO1cmZqJUHpPkMQOoTYHhiKAnzqb+GS6HEIe8cWeo/ryqbaJmInlFglZyh
a7imm1Ah0mGNBW7wo1ouSPCZVq0fR01UMRsJDlV4fbbzRCFQ6gM2al+3UuPk
h8jDClJyGajHqOw0K6xDdHQ/WVMsqdcVv7XIiF8YlL0TByYOQouzM6smEILh
KI4OXh7MIYRPhhFs43e5Hs8lhPXax9E0TfPjmUbVlnEIIrTACsUKhKmq4cCu
+9K1Sm7z8nHWcrBwvwWnzKrWpTbJGrl7r5hayOoRlnEAWED6U6GsLIdeLvwD
8XzxOhgjkoC5Z9ZYvEKIMVZRIZPCdu/qYd78xGU2VZLH3wSVBRhP1caqoSdj
6VVvTx1Qs61x6eudGnyCDadX6QLqsbPhGycTvKJ1zL2/XVzk60E5/Pjcmi8h
Wu2PI/bFM3nU0iRY0er+xOvb2sUP+/f44y8+3Roekor+Pnp930w7ZOWCR29Z
p/2w+64enGMPRA62FXqf5KqCPuoKssFHXOYHaqVZwR1j0Ef5WIp7l1jWvx74
zST11OOWloZCUWikDf1w/detSP2xRByY+HNLQMgd8R+MWmJVsB7R2JP/tHUk
GPVtsShs+ab240MW7pJxAb28v6HoAycRUvoO+3eWwonjtv8jQA7T9S2D86ZZ
Dx44DvrnoKy8vu6d614NfAkN5CuglxKRAB7FwZwCYMwIhmBRA+Mvlp844Mf5
pBzF1zJ0xWPwbdLFYHmkRLk3md9vrJYEXH5rjall4D+S7Htm/zmmr2shCoXU
uV1hYiaIm8KgrDz9hZHDip9dY8VlbsM8mpBrMEYVQsfzWqiH7LIjo/xkr4uu
QIVMfCLX3+w9J8ifnbR0ypryHNsH/kYPAHjgaAR+vaT3w4mC2EzSL/CdTZVc
FSX27Q/kGAetdcaPQZWpgPWxhIJgLG97qUfawP3rz+0tWjena7L6TKNJq5WG
mI29V+ezaY5G7UpLT/iL28h4pKp2/0rMZTaBBvvTVt37WEfDP7nfjeTZpt2D
Sk4PUHM2/B/rm2f27wu4jwccYh/cTpMJb9/pSWBmobQMOrfKIDnj1Pz+mPNg
1bXyBoZ9fq1vXSj0/pbf8r9nCUvors909e96n1CZv4Nr9fpuX0YQGm1GXU8N
olHqwGIlflhyYScDKJi3K0Li3WAOaoZq4/JrjlGaAuI8C9b9stnW3TNbIdI/
cunrDaCCEcWFrn61MXDnLF6X9ax0bdOMdkSXqQ7ntdf/yrYmxz+2s1HsaN1N
xEhRkCGC9enTcgnbRC364FqPhaRmlcEAFUPOtEELNhTMsL63uix772UcFPeA
9udDSN8Q5LFj/BED9swlpHUf09qXzK0xXm3eOYQxzfTUbR6W8vjqRLrz0ODZ
MLvgLJiXVKl3GTlqhpLMjmMZVT9TURNdSjzdSDxtpIhYsWlKnSACbfvHt5sC
6ACvMiYnrLxPlnN9yLd+2/gRPOd5aZiKAaNNmIyYwrzTutDuG0JV3FOow7nw
io1X5TnQwiZ0lFyIomudFjWZO9uGcecjxLXxFULksmtv/qbHAlgZ1we3/905
BcB6Mo6QYN2KCS5aauX1JXXNICSkprXImzOPYi8t6rAyLvg4Z3dsAmt9WEwG
V6v4Egbin2qbfuimqpUZ+3cD94D4XTI4ar+gEcajHwiyTXL0mzb87aerBNAT
P5w00tEuAE4X7qQxc2m+GkQRjdY9NfSh8uCPtHrovDSiPYK1o3HO41SvaOza
gZmedG0eaVLOA4qzIMalPiwLqe9QfQ4fbXtfS979XCi1/VxZ3UQQ8PVNUFPB
teXRjzuVe+irTR6PdShkv7yoFm4ShahUunklndk90nz3nzJSwS2a/dupi0/A
pHW0toxyb9Rtq+PLYxX0WfrKy4ssnDm3me6MCI3vaK505C5I6ZC5z/wT13Pa
c4ZkveEvF4VuCkfOawxG7u4rbpHDtdCrnjbRAsFKgO4bylYxeFuhGLJPN814
szMmE1vhuxOHa7in+0TJQAJWTwxqVQRNNtMdz7w+H/8lC4vRhU51Zlfo5PA+
F/B+aaupSoJttbMESK6bHZpcHbLXUNJP3r71A/z2AREfQ2g08AJ5K3QQIC71
JuKBFKOisuwrRx4V7aE5jRKOOTQEqJYz7ja3CzHnLifb9dA6WoGSx51PmE//
ZavL1v4rFjtdNdhiuHlWdQNWldo+yPbDO7sMrCu8f70GiuHXQyPZSyXm/Pp6
JR8/AV4F9FblkhC6fyMhkndQHq9UVWsaKDPJrRI3IPhqLjWQstKsNOLxqsr/
tJBrioTKkaDDHEbrDxONPEDzSveTX/u9FRky3uQOIuOuJnRteD+vO1vrHtIa
OjaBNCec19MvanvSTONlvZImN4ybZXFGDx0+eDcKkyI8nSaq8t7Oq3TBwC9g
lZsHOxta0XrT16LjZXD0AKjdny50DYdRiWvRAow9pHr6JhDD1lbSoaygHjtt
zZ2UxX7aPD1vlewcPgKjDUG/1SNkwERGgrb/sglKQs97M3gFmFgjMwJpt5V6
TN29q0H5mDG/tKyL/QZBhrJTw7a0ksLn1VSbTAChWxk6QCbaiN+0/yIn16ZQ
5ueeDs5Ks0yRDMtaTm5EUNxpXQD3kQ8sLv8jAffkmgPnq8jgOsakHJDIkKRe
evrJYL50+LK9aFHPZ6aNvuMEDk4qscqt+2KAJ0yG0OQsfQG1uwRf9V0PTYTR
9yxhY16zkK82iJXnaSJsPgOBBF+3BLs1CKVFHrfK112FdqIN0ngEgr6cZAvX
3yesaIwvf5vf6d0uBXJ1MTV7AdgdUTL4QaUJ5O7Txhb2+WBsV2CJS+KE3q+Y
lmgq1w0wB7XDrwd6cob/vYbQWUiF69KCcQvsKKqJy+1QWLSXwTXuLsCMjHoI
eBuo1Fjz55IHoIxyzZun3of63oi2136IfLpc/gcVKpL8d94RpCYVtKpt1DN8
2KyJQIsahmPrLZU6XgFSnR03knL38Pqi5cQdfw21KQDzR5EjRtuaYkucHwnW
YfYM2P+fZ8x6ddJ+Ysgp2AeyMiVD/q+cc02EQk4PUrx78eOQ8AF9lB6n4yrE
TCRmbt1D2WKPmbTj7ub4RiBoD3qmMYXZUfDVd+yWxmxWeWZ0oU1kfsU1TL4C
ipvc63isEw56W4L76GSmcD7KuxG+cGP/kCO4H8gaqYVEmBTojFPzCWCm/oYJ
03BExwLBco8itDjMWufWiqtpNkWbAiS75m+37uBjRYyTF8rA+YVxjWSZyylr
nrhcURDYJ9wZT2ty4upDDKjKMYetzabvGAy1k8ESfu2ARIqB1KOiq3KZ1pbB
cHYyes6r7h7ioKaIkvKVYGdw6bYJzK4T2Z5DauIdALlOe8vQsvi0xBIG3X4D
jIB0TWxKOn9FwvfbdlXgkZ/dWQT1iELU04RXz9Q4R/pDflTtciz+TSLGGT3z
TZr6qhsNDP0TcVhgd51hkm/ySZ9+wCfiiea/EpShyjrsM1AQzluHXwJGWS/F
DUnynLh88Tx40cHLqIRMw/X5jhw187dYDCdZS7IJlCFJM0w29igMhjSFZuHD
M+XEp9U3EpenZVdaZwfSikfcoMmrIefup6uV9WD0jPX9UtbMQmDrPDPL6GdJ
qyg2jIHOF1y1pFJ6EP7V3ch/n1T8cirXat/PYXPKiyt2w5GGcD/EmHZ9gDpQ
U+XHOc6rKUEoiP81P53+mw6VZDiElc8JaAzSObQ+MZD4lZLi5zLzWaTDKqGg
qjSIhCaXR7oh/XWKELTZo5LA9LBLET1jnWO7/RcCilFtwTrdDraj/RykIdOF
50H62wJ2ytMbO+ovZw07anNDi38HV46BJc1IB8dm4r0gzbKhbxuv7tmblG0t
QWd2TsESlOgqW6H7PUT7RXJZnzyUKSBsgjuQ7+yBSeZMPxGvoHN/HYFirG3O
OVqIZ+kBh+M4ufRBKCujYSKsge+0DKO/jYHFas3pBcRb4FQYs8KPF3n6PWgj
z87rudQ36Z9DoZAuwL1chkbKuKiptLj5Kid6roikHVNf89hh85hQ+PnC2tdM
mIrpgUkW1CodUCosvyi2qmaY7012jxfr5moalm15lvLYJ47cKaL3ppKqgrd1
xRRJ1RcRQTt/RfALsFdyZ36QhZ/AJAnGxwsc9c0Xv8ge6Sg1pj0dAVALxaG7
wueA/uXbVTEh70GpCGYvRzoPkfEkHYCRRsN2Nj3FDkyzCuqC7ouZW1ybktQC
W9qjSMNv/EG/tYrOcmU7bsKIil7WVvsuHGuBY7l8fpA/v/HtWCwHA2xtUHIi
iL7mFIbtHZOt1mNurGB/f01tLaknUCW7gvaVwF/pzKzL6zRMbYLMWV1gXH0p
lWF8yJRb8CGn1dqFHQ3t1Vu4dMrdgO7QOSAlX50PldWhS4B/cLC74N39X9/5
XnzbChXCh00IpU8aAy6TE6nV8i4uY1SpXk9r96tM24JrUn1Dz+lwcQFm2CMg
dqhvueMXWBTZevpei5XaO1NxM1lED7n2MLkW+48dw1+kOJ3STb7OU0aKmfKT
kLFgXvXA+P7AoxFkM1FtEVUAIXWjg0tQIgfYSp3Wyrsqbsrx3ajkRyaFNda8
xthI+ahRowxPCQVRuVOaOqV5Wq5DnQFEbnnFWz8jHxOzd/3HpFHtCZN2d1ou
4JjBrp3LII9csP+R4+PPrwbADAUHfqXvcdTfE15UROGZk1tNcWRUYpk8HjxY
ll+Wc3eD1fJvunKnLvRq1h9DQvVgBBZ6/KqY+0sZKlCVtR6PAYsjrIIIFzf1
O6d6yCic97xbz3RUVHrnYCE9LlwAIZTsv/WG+0xuXN7xu8glANoKBtlmTOb9
X3gt59tiplT1t5uhybAkzZ0lxgXf28ALw0ze+/HWiDFO9ZYrG1LZC1SwqjCC
vu3v79nuID9ZCSQ3TKNtzpjPlyYwNApESoknvSkgV8UFrti19KRD11AmlcHF
cpwOT7F9VP/iRvlxiGqkOVM8XY8gpvkE9BW/ccsLCQkUlQWVJghBiUO1Npp5
mx9FifjCUau4UJ13Xwwx0srrgIB7L6XZuUZz3YLsIlZH2ZyCq3mLbck5ESDY
tbJTdiQvsdZZDKXm0NgtX8WwxvEwpWI8PDD4LMGBwUnw/OZkHBf+AvPpvUE7
hJdfLOek1tW3Y4Ec3K4YeKMRr+6hpbZtdz2d8azcy5v9noj3r4ZsOmsEEOh7
9UbpU7XhpB2d74WAok7dhfjlRCxVKZqEk0ANBNSeMcaIzWiZmJPk5HRrSVNu
hYJx6crva++71tnQShpSf4cysZM6EWjKcqUsnPJVMIYU1FJixIBmJDCQ4gC1
JQS7xTNhgf6f+T9Dc5XilS2gblOw7EX1mW1StXwkB0a0KIDBo8uE23y2Nk3r
uP9h09QORvwLGjQNsWxnfX3ZzVrI2TH9xIseEVLolGRjIz3f7b1HIbZbl/18
Bs4SopipV7yC90B1wDHAYjYOkW+6Xq8klas8l7UbERTvhmPnyebrdYa4Xq4+
5G/jkcZgSZvuCfoVdKp1xPGKvuSTSoBnyGl9u/+Ew+pI2Y8HIKR37ONq52MP
P1LMvNT5ZHnXf5jUTzukj3VUwbF0PwCN8VdlIoGR1XLP6N9/b8ntOq4Qx/cZ
ZnHozpTjD9qU3KbaLPX2XztTthr2dRqZcJXOi/UJN5BWMXIJpw9nuxGwDVUT
+2vXCxQmc1mhNRF1z2bkmug/g/IAEf8JXPFm+k2fJysz/Bzz2gRTJCR1piMA
bYehlcgawYV7TGeneX2oUOuZtOV4m0hTF0aNl7yj9/zWOuMp/XFos8yX9GNX
CKlQsqj3xjwpzTz/XmJOO7gCS6+QObvDKqgZkvIiqFicXp3jhdSEdkYutLOY
ElRUhkxNWuG+YCTzVODOLl//O9zktejJpVvTGkhUM5wB8kdV2tlawZIO+waY
X62AnvI+/gVYEluaQcvDR3boj4ih+Dw0j2nRyOhBvN770LAxfKuSzeeOkFBP
raSpskZym9UPFOPL5dvG8J0NOH5QgY0jW4tdOJIBIszG15F1ynIttjHO2YE6
WHJ82i3OmGLm8v9MM9AwQhNFudiYLuy2asPkbstaiORQqSAlRJIooSxHQLNT
V37elleQgTZ4YT2aJkwqKxN1GVMAKtL30nxBi7OZvUA5Td/bplxe/C3eSo6z
tkI2o0FSgqjJyPVGIZXbVyXa24JvilXk9B40YHa0FzIn8eX7sM0Gwko2mbmO
GzRlnlwXVOwwba5nUR3VTazEm0IOZnoQQWuyfBiPs5chjkPB9f62JYZsd+D5
pRDymhdFD7T6m51W3jJh894EYE6wZ394Zm5aHt8rstc8NCFHDqYF73GA1W54
ijXDp02XYBBoK1+1B8ToT6U2yGpR9LYhYxV7RO0O/bIxwYGkEuiBsbjj08iy
avm1UvgeqH156qgNigAuTyOIgx0eDVBqoagYAz2U05iggJEIMYgx8DRSBx4v
EINd49KKgcTTo3VK7uq4HMqSOXwOvHAZhe/t4IZ1L/YaNhQUDNJLBOuNqI4M
H7CDgW+iBeRyEBFMD6tIf842jhvv/PcKNUglcQdg90bSNcSYgpGfyJxobloU
0Qntuwaf2ufd5DvniLdtiYZaGzZ0vWU7WBn9sfqpW+W2AFAiq7SxCF5rgqZ8
pgq34u4orsWNZqikFikOL2/6B+uNQV+5whiNqiRR0qs6XVv7E5O7Z9yb4Z+v
7645vMJdbza6+osDJZOmFfdv1hnIfoG4p+UvXIepTogf9M1z9ObkOhceu+HU
hJEq3edJcKJPnIlSZJWYwh2IhVFMUB7DAyomVEqLH7csIWkpVBxhuiuheENs
773S8Ca5ngzYqRRJ7PWxNR03VcIXVarCgrKMXKrnskWA8sc2Dof38p3VTdoe
IR8HyUC18uGZWsxgecHJhikPsRJ03mNqhQvjgjkQiRw/vcX57zk6vDwlEfAY
8By2gINhkwPqqMcZwK2gW+E6QCKnwzYBBezhKUMiyOcJ7Y9EJ/MBqb2FY1tm
irk5fKIr9O5u6GiUIhiP0ftZIZ3LsF1d0iyTtd+b7kw5ZMX9B+xLmL2zeAm6
pvPB7ldjIap5ippNKThJ42bL3er1NRaFa0uPLaUYkh2RdHo6lT+DahSU6Zeg
5XJsE9+HvJzmN+gR+XkDoFVCIfjjQzlVGTvcTRi19oQw+mfeDBQt2+K4Dgj7
rwMf9OFlRRMBKsDVCX3LrELfaQY/QVoqJ5+aUsmRZg+TfQGpRI91r2RXof/G
tN2PwqGGcluK5xfguDZO9rV4rS4DMN1SQoiOSQbblB1aG5I34YnTzeSY5pph
tTceLSnP0NHodMLubddtwFrHOni/t9Grrc3bGYaHF2IwBm5IlZ0cYygUK7vW
f+Bo0fqT1wYbvgdCcLD4+/zxmFwj6tlN9WSx0eoRTjcKhRsod6xQvANrFtLt
knIAY3Pgj/6F84qkkf8lsDs9LJhK8Tz7JR3jdxXFrhkQoiTQajZPQQV37f0M
7Zglj5x5vXBXzomukxkmamUT94d9ZOdu31Wej+/bbdlO2atsuYzbpezHR+KX
X1FH/eXXPd3JikOYMkNBnp6stCyuEShvMfDvs3ifzuNmEkY8Hufu5pTaHIRZ
0WrrBI2iW/pgtb8zuoRerzlPc5oismKJ+cfDE6EhUfVuobc0VuQ37tuTfdTm
0v5Gp0z0kcKRYAajjaJWj3PRCYgkpO/uMfv82yH3sepcSDZbnvaa7GdfnOCl
aBFchsFtdOECC6WXkJXBFf4+R4KUVJzMSOkKlcR4Pe2a/RZS5+JXyrEC0bE3
jUxBjpgwHLR7Hyw7li5QE+bNwaNKMcBjHbdu3GwQ5mug+7ay1ik8Qtib5klH
+y/f5sqlah9g36OKQ2z92ic3zBYnfEBHGWNKEz1KaupPRuBBUampk0b2jLI8
tnhDu647SKlV+D1tTn6wqWmyBat7f7AhKO7dDL3ZNtdgpnKkENvHBQwZaE6f
wZEXL/oVe3IOGrgZG8gxmNcm5zyT14S7w0WLNC1o0O1NLUbnzGOA5ttbbK+6
U4ReuHKfzjYEQTQ8N7xX/hphrJ46xBODlfoKYZar2GgIniILU2zLQHNv2PuN
sTamzC7Phh5ajUlh0XWbS/ixV457G1LURd7LUVZYUd7MrY+9W1lNdRRCp9WP
DMEe972x04pSQluF7RqslwXXsQmpW90qBJEzw9E1kbXEP+5P5i7wZ09fEOpL
dQoNroukHGAq4rmj0d1GUglJNkZ+ZVagBefAaHzyczCNtXn92PLkWFKbVDFm
Br3NeY1FtDzlRIiUw/yFn5wGWQMuogtwXUxvsjgZKrg5gyTvif3HzcgchSPX
nQ2IX+3p4dizrA5pu8/MfzTQyCXR6WgTcpMAb+M5OQA3GacG6wfYv7UvDTn2
7VxDmeEYBmUdJDezT6PF6syN4gIRV9ZFc25DFOqw1wNcR9u6fMcnjmVu943n
XFhAidgHiEFvuZ61aK6ek/HvvcqdiuWCY67kM77pNGw/dWbPSY3Llz1m95ae
JHDtbayQKBja/BGgvGx1f8ZONtyZwgPOtFSs51nTxvRsKV1XzIHWdggw3E5a
9cZHfp9fOSr+x09aRnJIhk+GgmYVYoyeYJdz9U3PDTq05Z0OzG86+FPZvVTH
1CdSJOZXhhpj5DBtLy+fTbm6IVBfIsxHyoqyTDnzec6hB2JPsH2Gvnjv7EXr
FSuHlC+T0clgfhCIkFhV/Pa9y+abw3LmP9581tGQ40sTTsq68kFzx8wZ1E7k
L1+Khu3XRQzzKFkTKnu8JtckvaKMfJN50Sr8wdcuPOKN5CYnBg7DxUxtZ/s8
RndxTyF8ECxqHBkQYwS6V45LT55CcHcQIumx7jMlKeJuKLwS+s4tT1dYzjdB
NhdYAdZGlCkr2hJTuNyvRyOCE3oM3yJDAyNKXTVUVwPZ7LOVTmn1O2W6aqvP
H6pQn3VYvOPCwCfrqqu+nHPFut7m/EfMER8lu0wNmdhiFVZ8OSdb/R0oo+ni
pVcwjXIWNsrHlDGnNOWBEdeNni1j4ZJu2nR9/pfIT7Nsyb4Bbm4C0eRrePqu
1ZXqOUh+2tCM1W3GbyDTMzyEfiyb7qgdlNtKKrtZaC+p6mLd1Agzs2U0kN1O
E9JiPG88/jislhJfKBYzfssPaOPSeyBpYAO0CZtY3/k+FWqCa4EeSuvI8Qjg
xz502Q2gTrkpIVrcaGhDGxKOmNe94/4IaiFYCt/sOSdhWVcBP9pdFyUJVf2i
G0GX8k5is5CyrHOshUdAkHz+H2nxEvqwWS1Qd5S/FVx6J5/tyXbjpz+Rc4wt
ObJfvJ0OQLDyLyR8qvSW420pqhMlBwhUWgiPORhbAG6N+EY4n8raGqn3jACv
kUgSRRDk4XBTRG0My4REqok7WtboxoQdZEFjS73MGlXI81n/RgCLqyNYASIW
4Ch4xFm5FN5Zd35q7GPHBSuu4Bk5dZfdnIYsUDRfaL+mCFFObwwzF9u0EEUc
ACMcixYUJhdCspwIocotbpvEB9/BpoXZjhvkJjKVJjl+sS0KAheQcuI7okiy
fQuHo4aKLo1qKPEI8c8dr/JtVGQCXgaet6LwtmhtF6S2wDyRURYTFwQMFL5O
Q+0v8ch1tN6L9bOW/3eQcDJUm2NFyuD7o3TrjnYaLtqN7u8X3I/9xMmrO+QQ
V73+Qeqdk2ftirLmCrBUq7ZQjOaxQlbkP8aie8UHBwL0FbnWEm9KzOVdvI5X
wSbw5Gw1RsJMYe78u/zU0r3Xt0OzfLUPDUy2K1HXIdcxvNk5ADdy/yFea0z+
aOeuu9D5evQ0lCRYtoeAjfNPNMZp0OptsAH/+J/hK0wF3azoTW/70q6Y90Bv
VEkASO4m4Fzr3s2HP4IGuZmP79Tuo79f4NmESF3V33OVsR+WJqCohxb4/inW
hb6Wft8gYf/kW/cNB3dablR+Ywl4lNvVhobURetZXNn9/HFm0ZmeIvyHguYL
6e0wJhHrD3OXH6iNHdkDDAvMiwvv7QniRcWZf7R0yJh7LgARz4erltI/1SSa
1R3c0rHQJ//lgdSaJqnchxmocVTQ61p3CKYah6wE4u5Q2CC2Olv9g4KdreVl
RtJ3/AzvZD9qB7wU5GZcWko5gHQHnmoxlvjn3xyUwYXJ2uiP9UB1Rw0ArNk4
+fsyfsUO5LbEVIaF0rtuadgxwnASaplM/LopcAtBnpm83RnQHLt4wjTPT0WI
GWXwCU01arlda+0VIvJk6eeCyQfLlyuwOyUpn416TJMXyGNf74ykQjJcNfJ9
0ZWkCTqwnVz1g2t+jet3hw87OsaprGwkOZa6Of4jKWBVxy9JFtVYjUP046k5
iVyu5IslrefFHqvaAMz8SVo0dJ6l8cxlpCqz+p5USW1oUkwZb4C9f3RNDgTa
VCsEs9K5zVTG/7kjQcYI2puKW1LdW957uUnG76IjS56F4rSzx/qJZZB/1c/H
Vk3MOHkn8obg3FoH2tveyCdFQvBmkfVraBM1UyS/Q96M3zgyyDlqasX0o8dt
o0HmsmjYEpaQ1WQTJDnQqn25blWcfMEBsGvDI+fbuVxyWNu9Fb45CmZpj9qT
bQfrWQqQO0UI+ncZb7hXenkp5omVYrvtiSrWKguMwAE31lyqHKmksTM6FerW
kXJMeGljAnK1zrjoQAY/GkWVDjOuoAHaxoaG4vxLmtUkIqZytawrXF/HsDye
Zj7hqLUFC3THrtC59UUB9Ph++Eq3jLc5B0ZP/WEK5T1sxXtqM2FvDuGTVuHj
0z2ESxVrDu86hSycTWVxs8YCFZNguLhAnzNDrxHfn7jJD0qdpj88ZC/TuSwW
TFYLKHRV0wvJMMvNIiI5Tp61n9IkVPEyG9qLTNHb1sFr8CEKtaSLNsDPhRaM
MQeROUp8jvYbrNjZgSIUfOgckjcYAK28nYt2NxfbSqL0pOnZ7103DZEKKzqX
kaak1vCPnUEr/TpM9JoydAsf8PObUqDXlFHhO8nHeuXpgp/K1JcR2wHhIByH
VRxch7VY5320bv3HQOzUIVLhpCmdt1zBybGlMVnt4ssM7I0gB1GnnpEAGHln
v0Bo1ODMFFtpSJY5+o2KTA+fEZon3k5+5yqqIgy0C75cZOKw/kaSTLAudHNh
mHZc12x5VdpNVV4MLuspO/i8flrGMmkbLhMLFMHrLM++Ryn7DlKMU0JT2fDf
lYXPmfFKgzRYdfen+zlZxkrD4bymvx66TwB5AddPW/oQs4xHDtD6u8/h5kuW
AYMZMXHz54DLfWR+ahlAcMLOysRR3Xw+wJuwHFJ2mvw4vpCvxYgG2jII5v40
MxJsrvzgUOzUW0F0zU8ioe2Z3HsGOSaPWXRkXSEiocIHItAhj5+lXhQhXAs9
4iNkyQtccF/er9HKBRTkm2vQyrblWKlSQ2MywRaOoTESDI9W8YpWBz9CFFbY
VSTVkiQkgR7h9S3MFVQw3HKAPS+oK2ayc1zvI7+zJ/yxDFUWBFZhodzrcKzH
+aUu6UT02NmRdIWyUePYUErSsJ4yqYksqfgARyDUycYgXEPy3xxQNQHbot/y
bzvLkHFPaVYVBQXI3+1gxhI9bBBFbOuvoovMr+Lx1ho7hsWO3MMbnWFDcZjg
v6iEQS1oMIJCzUpSbtdsijGCLG0Oh3uU3hMM9gFNe1FExSSQx9dkGfkfuajR
CHQnkW/btjed4BixTyL5RF1TBy1Ejn5zDle2kjX2aIvHRWjAfsQB+lut/TJ4
xnmNaolQpiqbYxN0TOMfCFApck6uxWEnfSwjbSeNjGhggX79SA8pqbddKQlq
MSKKgKO32uOGbohWECga2/2Q+ql/k7i4TD3BN4uWH6Pb1Xd1RpU3opL6PeK0
7u63at8iDZWpcSLfyyTFPhSbGrmvAo4ZUO8jaJ9DOrPY9LqM7tiTrOmdaC9t
7qMIRweXKE04BWS+fhYmMhJSLjOgFSP2aP72KNff/yB617kQWh8cTON43xT2
2JY4zsD9m7eG9J7JRBxfB8O54FororR8tVmjRncibmeKmUF421XwI2SHvNLW
89j8i53wsxAIvqbZ8tYCA1ZzvUuSIC3v6VGxJVXH7aZfJt0QEEOhVWUa3ORy
XfDwt1bTRv2nnfarz4wA9NxLvOqxzPhtZu6ohLgnSlwoQKBbHJhDAHD/whzC
gyNcntuFlKLvJ7dpTj2cJ38sD5YTEpR9oxcdIhoYZocIt7lqQQpSR/L9DN25
8GlwaNpLUUFv4zeBDpBAAQSdaPvfcDq2Niw0os5KCwCyUIfRCfNhyEcMCPZa
uOLNL2/k79tGnv7m3rtK6AYfz5y57x30xFAgLwwNHhl2QeDr0OntDaa1oY1Z
TUBFNLGRwx/nRKTBpKBKM7ofeZQJlNPfNBGNf/JiPKVV0RuWx1glOWI8s88R
xXsSw5dVOis0UtLO9Ix9nTjcllo50ZyDuyBfWwWIb8NgloLaW6E1OXeRLDoC
fwMALZdPzR0aW05RWSWafUEXzZcLxWDLOJ52X2+0fS+hfs2UCNySvHRZ1yH4
T8gM+4wO6sTQKW/2TKjfCSFtNPa7yppsY4jTnXS1cNLE+ybo95e3A5vUWi+r
6ahU4V6Mc3I9Vt0P+2fxkqNd5OX0hQ7tqo5iISjnsdKdGx8GJw5eeDnUW0qA
jHtq2BwsDDreckTjFzbidnyUJyWjVSK4g83zWkUPjdFdt7/nM7v+ovvk0ipv
I2xFfxnksFmmJ1he3CONiqym9NLnwWXOxJauVTnDGQ2ya1pBSfIicWJbbEXX
+A6YShydXBzJoEL3nrJKM8d7uhw68lCVSA9xyqKjQqSK2dexvm4KHNQQRbdG
LNy9jfdLhK/yKLuvo9XfaWOLSSWTrXkIA3u0xux+c0cpMN9FR4bksayRSPy4
wQUWdSTrxwUxAph/IgO0LRY5S05wVWxf9TLDKrMxoZubAMWnK2ApHweubvkK
bnnqpWHn9h1Ttd16fGwuhUkiZQS6WUGM0NbRlLScT/2TeO3FdqJABhq+VMw5
HIIBUJPfb6c9+FIqCnI1NaV5wxKWrA785Ufoys8yuX8mPvobstDS1Pgz0UZM
iulbGjJM4U2SVHu7W7lYfNrP7XfNWh5DZlOhrqj0gQKv/rSk27conNN+LGF9
UdbfVjg9pK6iYQGWNc8s4FXZM3Q1idQ7DdwUFqJj9GZw73MiIGKmHCfdsXVp
h/OhC6+V02CLpQ9jgIHpJxr1HIPT56PmiDnTcKZvH/Qw0G/ozRGRJWS2HrXj
+UNyFQMlzcaMy6mgTE72vaTGndQaWN4zftJZ4EqHE7eg7mXVlGIhGv0Ql5sF
aaQrKJH5ZnquwPOKmromjsVhX9DfNBG7qb6hL20x6saK1nPxLZ32VnZ6nEY1
gP0RcjeALVLM4tgM6UXT1Zeto8p5wI8KtZqabVqVo5CyOi7hRbRnKa2VrNkm
3ioQGZlB69IgK1LwiCZKTq/fDTbl378ObNsK3wkY7FwqexkYUyr9axtpDQQa
b7xroLbIac0d99O1j5UdzS1HGvYeaUa55XZdOMr9N7aF1BI548+OS3LkcZxC
5f1j0Md4VVEEj7niNa4v6m8i880va/O2EC3MvJ5n0dxk7TxQJmAp1e5Z6z5Y
w7/RULl+jEov50144SBTsVieOFt5iJR5M671UjHWp269Q9BcC7cEQMgovCFf
aLhPQ8RSsXQ4zcDvO2tPCj5cDvCKt2daLfkyqDBschDdeI3pP6VqNi7kWTbs
AbPTzZeNCelXiVUh97O+Rvv4Z8F+5q6qyM2v+n74ZVkPzAq3T93mhZV26a+E
7Y5mcLHV41XrErWiB9Qptg4x2nHT+5LlQabV8B50YP2n3IkwPsEkh1g1746y
8FJqCByaJ/Gvae3izwazcBCeTeiG0sV3kyZGsKYnXNjiQ+EOu3Zu3TCbDMyz
9wP8kqbuNZdcIiWvzYNSOtqiYasMz/VVjPt6FN3C3Rvk/BKoGyYZ9vYApl4U
KNHFhIRhroMspAtPPt00l4xIXHT3b2EOQ4r+yUeL3rYbwqZ2TC+pGIFu6L0G
y1SRfK1g6685RRiPMO09JSBNbbs0TD74SjCK78QkJm3rdDPn5XWEpYK02tu5
Ao9AeahJxLi4tWcIYkdqgwhC3s92iWRiQkd8N18zD8u9iSK2jxOLiI/hleQH
Len66JXagp3vCcR62lplfTto7f14Ihn85m5hADrrXdHVqiwzgJqzo19lATIV
6skybuyAM6/DXaj7CFs2K2DmEKMTGj/q2EgRo1VKwiNkC8feQqQ/y7lO4vJ1
0kL1zZ8mhyvDSE8aNwEM38Vqe22oaqvC2pOE8zhXwzkjT5utHiwQ076iOHRo
kibebTbVV3g6DWKN0kaNGomTH6N9AKLM5Nih1SNMHlBC1omdCsJ6G0fWcqVs
N4qOWD1Pd12x6RwKDkfR0NDNAHpEyUTSEjOdTEm/AGofvBFLRw+Fvr6odaWy
4e3em91x2y1zzY2Vbe5lKSBqToCH4Q/t8kv3dBPVgVSfjtVXQg4eunXN59eB
Fsagcx78AaICn+4XBaBV+XsG4+2JGpDmTlh3wWaVu8Zj+i+ptb+UjfW+eKYk
0Ux3/knuyBBHZUilg18vsmRx+FiiOEaCQhdMVk4CXodXQBGmEF9FojNnwQ1Q
/aMbys2lzcOQoSAz6Z0ogaZKLJXCTFy1iqXe8Y3Coe7JAHYMetzKXfzhh/8T
A7fJE8IJL6BZYk80nUxX8IQkwTAM8F+PeA9WJNVh+JuJ9mEIt6adJbXWFasD
pBaFK14ZFZQ2o0foxVSiEQyqPP+niH+RnBEd0/46UGDdmBYtj2lUluOyLR1+
Qrkixc/rE5LGQHdPAJNWrdVAs0GhboC5tvg+yZ3ZO9v+BJ2w+yClIDbJuC7S
EhBxsbivfMwY8KM6bWL0xJ03MAGMbMJr1v3xaqDJbxIqfCp2qHIoOOyB0p3U
PIBd/919hFMdXATW61asSMZtV+jlZwSvpcyYYHgFNJwfEK9JG7O7oUWGk9sV
2h8V5fwsyupSn6IfczQkma+vb1PCtb5gr8ErteffbZu3q2k8Uy1bWOxWmAvv
zJdOBz8xDrY1SD2d4nBIQgifOew7zTW4a+0djb5c0yIvfG0azPeBcCVA8Y43
BWnSrq+vpT7ok2YJzw5fEz6KRCqrNJeieh2bHSsor+2bQZJUd4ABeY3U9yF+
F5sKUUlZydZejM0nT+kOlA1aHLyCmLzRn8LkNEFyJv59XY+kiVI/E9j7g0kQ
wcwLHyb0uLX1gqndUYkB0BQRyCDmtFSgnd69GPNvsaijJoG/Td+6MQd8+RGE
TqUalZswabW7a3sFDL3QYDbm/zNuWqpvuS+U0e+jzfpPLKnKVherxO3CQ7Yu
qvhZUgMeTAA3BNISLGFu4p8qe9KyhCStfpNmXiuvuIBkFsz4cavszX0qkUdq
uqeVcIPuzx16pVjpUKhAEquvSUiuy4wg1U7VuxKoVJ2haKJ9KmiF3/GVLYwq
oYiCZqMPx6UWL8WTWKfPVILEQstFrlzoqcnFNSXG94M0ySFkksrWaHw9r94C
GU9leCERK45Ea+jQP2n+X3mu7MjfWp/rvVcEBLp99vA4t2Ckbgn5HYIjx16X
XR2YvJVM63fcB8Po6KHXA8omWYFmM5RBu8RhYKZ5nsDtGrVjITJIXNLCVW3N
LrG7dXmNsJ/67mLbH7uiB290LvYURg5hmI+z8kwENKa2C39cwSwlA93MJ0Qe
orwL79OwlKxmFoUXvd8UE0gw8yKA+pvu6wdzSwBMA6WtkIgZ/JzrdZVPd15m
wnq/iWl23tUGbxHGG+JP2CCIBZNFuReH+nF+i6FJcp6CQWc/svKkWwm2RHKR
LBcS99xiNCcm9iOYgtYQp13CtmVHP/geM+2o0z4w+Pfqfl2NY3leLcFTTrCw
RM/EgtqquXp6g5qdK+Yucz+XVB0gFFDitRZFrCCqRj8UmeSf+bO5eyfSnbsp
2Wwh9WZ82hThpy+P4yivTlLaqR76oMo++Nn+kwS4ce0BDo2vCV9tXO4hELIe
DM7A+enkkBc/pYVZeIp/P+UsEFu1IrImbO2C7e4nOvkRnB6lyBcTKrnsnlu6
84f0baPHYwHgRJAn/mnmdbyoLREvrp2V9TgobnmqIovPqWqs3aRR8BNlHkK9
I/DCx0EjZKW/cwAiiZh/rZ0k6CnE7S/PQVo5zv7QL4ReIXdfzeaLLtKcvZoH
Zf6dHxElY+5nQN+v7ZPsnJaRy9zXdKO9OjrLAfV/enQFzJDk7H1+nYPhPAdo
UgLItJY/39NcDkpCi3A1pF+H6R532vnGZKa7LlmR+OGwYH87eFgIBeaQmSq0
96P5iOFfKQ3vBIhYuGOJurdfcQ7nYXYlW4w1N0JeejLgCM3creRF7ioVCce+
XtJ0jOvx5fo2iwsyetnTxnpAE+K75QKnEK7UOBYy4/8H+Pi5aFMBbIZbwFg/
sdgxG8ZnYxngR/3fCoyIG2QguEiwXHgSQMD9Ad+glDDSh1nBjC/N6rUIyae2
lkdNgO87Q45U/WKcdUOPWTqSR4D8NhklG5Uci3vMdJlGen94znVdf2iVC6CX
PO19+KpRguTgVHSvLlj7hkLqtPLQ+Id9gYYxyoQsMYceWy3L8LYojvOnhelD
xdr9R/6iHrAUAUZ8h1g4YfxBPVLnFGeMX8e/VBZAUCuwft3er2WCcU+a7XcK
zhtTgnnXbj3TTLFxK+4Ss+HSjCjabLsNYQjdZzPUTyDwzfL41OmVLwm9YbvJ
Zu+rm2KqbViQXFHmDo8iq2v/9SCe0LoJs+lC25ifBN3A9lJiGfa0+9giNQeq
IpPkU9Xpmq8Ax2gZHjWh/nJLGsW4ldDQWRPFSQbCZ4LikScrUaRWeSU8ise7
H4NSntZ9+kHraok0Cnss9+FjFsaixn8WrvHqq8OkduGSOVb0lMIr7UmGLQco
z7/krElFWp8s+FX7yVEdxMcCi2DNusz3bGwFXhvOhmlXwDSDlVjFksLFd3JB
KHJtrrPyYMUVyat39XPCnvl7WVwdxVdM2q3/L9NDZXCDhEiAOYh9GDc5cDb/
dzqJrdUDD538RkTgA1lU+twvYPkIq6JuvxdFb23bHtYH2GazOfBBpgwxRKHi
yloFKjtu/bkn8/l3XMF9gGRk79QV8t9m6aH5lWdQ3y8LkUPG69U09fO921aB
VGKejSpDX10/DcQYXbc3/rbUElmlBnN2CebqqyGCTd21iyaLsfJELBHCcR6N
07sbZ2E08PGzSXqND2E2PRqRZNaMKxGBnFZKYGq+XNzCCAGX+j7m7KxFfmg2
N9Pm0WsKq97U5VdANRwLJw85BrpO89yzaQPlIgYavnuGDPg5vVJP1xiG00pl
zLb09kyfcHxewOj2Zpny4TSVaHYebRhjaF/ED0SzhfmVrj1VPs5DvgjDwZ86
yTNcOs9oQEddq4q8AIOxqSKKOfAqz9gqIGPEII7WY0+itRzrIiyFriRmJvEH
8wwuE4mUsPvHrXCqSCoeVxPbBIkUh61+iCiNUufb3fioJz4BM3WBewuQ/9F5
bjGrLif117ciUXCMMrRINZVu+F+K2VRXHLPuHbgxm2Xa4QQOI/TcCfgeEf3u
IC+1silJb+8fTpIaoKGXENt83AEt5ThbqEQ4jn/Gw4XZyn92uv2biNiDzb7C
d8Vhn6aeKklhZlcyT9q+NxVYzzJsfBUZlwURuZLpjmMPPsFd63hwobnaLz+7
e+tOuHQ3td38QlFmMUsdHvbdGhkmTLA28jLxubgrFjWKq9K4BjlrlaFyZ7oQ
jowkaTknU9RRkhwpMVQLlo3rn1MuKOwwdISRa3bHUeYCDTBiGopOphnFhdYL
PsDyZTlRiINoza8qT+8bbuTxQJY5wXDYi3NPTX43CBUTXYPmKu/kzt2aaE1T
6FoNeJdlh0OL8g1soGTAWs4VupKiVlRrgRBmifvgumwIAHoaRVm9nk719rV4
jyZ7Lg60XfF8N5+6x7X28D/pKPkBwKNm0mditMDyy4o+pDhWzaH8eYYF7mYk
TI1t7riNUl0s0PKur3i7EL38SjzfL6MucPDulePoki78QvHB7cPgSSJFmmj9
SSTVELYzIhHouhGTv5H0+P8CuopPguVw6hRAe+hmQzfFYeJlShnqxBa/ma/O
+1+5RvVeGv0xlejFkXnBj1MumjPUXXjaKGAKBwGzQID9jbTgUHF/E2IXhQVV
L+qv/LKylBHtAhZO0aFPdAz1Zpe2fc31aFMhQnZSSF3JhuyYTP6uNH0pillR
PM1FGMEk90Yy602RsGIzXyl6NJedJsAmjr0Bd8WeaV/Pg9crurxhMDIjSyzN
HJGGEtDyxcJDGMWDOPDzTxFlcD47gsD0MEKEi7+2MIhgGPtbgPPa5UolC9AL
XpG+Sv+4e4vpQXDsflqRtJ5MqBXRtfjliafZfdHSDLuTbmoFA1GTalhH4aTU
ft4MhmJW0JwTVHC3ViUDjtfynq8tU1sQ5APbCKOM/IFHHEz1YgRucn6X/8+K
ik7rKfz0JXSb7eNHuYumbj4vkFfO/Dl7VPvIMEoNdrzNhD8G9sOyWPL4jETy
sGx5chT9zq73hN/bjE6G5Vij2lcLUl2jhETmYARc946Gzz7Ky/MNyUWOD8hS
/Jd5Pg/6CccAINvKBcw0eqBS5yVze4s6/i2JiszlQz965ERg7iB83E2x+oBN
bXmvMLNVpp37uFGoscUAyveWHqwClpRmj3b8ogwk7+vj8sDU0oYiVReT/J2v
g56X7SsCs+JAroymxUZ+nu93FmIPFc0VNdSZ/VLiISUBk/QxUTOXeHr62TKz
RnH4Jnhi7f6lzCN5OE8BVjyZmccRI2p2NhycdCRJv3nSfbgGaKGqEvCaA9Op
le/7qNkbSEwyCQJc/r6eP7gt0uDG/WzrgCzHfYmu9hX1mdSZujXJSy+Q/S7Z
UT/uAbqAjAxXujWwGagGPJ9yVudRj8ggc+C94mTPlsOfShBo2EuBIdL46Nyx
M7sF3/uZk5pGJUARcTIyIkHBIRd+PI0H7/UJlPulS2nPeNO3hSvEMvjMfkek
5qSqw2qEDlB4sOMhqKimo3oz5OZE1dJNGYx2UZT2xs1gEx6S/bM5CckgXkhu
us6o6ZKhqF0tU3QJNGkwrLmUKKI9E4dqCeh1WysFcwqcpA/FOIy13QOptwCR
D84OcqBaJ7cQBpEMclfusqgJ5aWbQZ2HRrSj5FGJcSmCsBjuQJCdPxb2MVE7
tYkQsHQtQ5LMl1WdTsySXQAkZlVb1CaZR2l4jDndyeRfbKZz8YVpnK14qjYe
UUZf1eElujsPIQADUl3ppZS2cBDMyezfofEmaSW0rPDLnz+KSJCvaZpxQbZc
njfL4KhpPKDTRa6Qmu25Vtw5aB+R02ztGkIs62iD3NP+7uunnylOk0q/bztQ
JSMUz5Ojvz1jeQUfraJbkR9gzzseO8vp/24LyEXc9X2DvRgiyPqn1xNLo754
+malMHIE6kuLJPIouVMdcsW/WFmKd1n+ytyOEmAvnIyhnrIQzcFwqlKl29Ft
Da4oIy/alA/i+yNqjDlRNqujCqaecgQQDgiR+JszFsm5L/AIkndLdINvNPJ8
5geeb4/w5/hasK1yn7jfIfOD/rWQY3RPB5R4GtfwHAvGR8S5Dsu5181py9NN
2znXXc1l1hTDxW0wBAjaISvzYHaPvUwBvxm6mXO8yEJTdh9pHvn5SHXBqrAU
p2QavHBzaIcZUNhc7jR5ZJx5XvLLqZWfnaNPhWV6KSqsWIbH3TFqEY1v5aa3
BpN66eA8xbaY1DCg4ebzcqpV35rLY1l8oKyBlLa7MFDQNlbf1TdXYqjkKtkI
+eJFHUZ42EREHQKkP7FNuWIRxD8kZgF/9X6QGRi0U0rmmy/FinUB3fRNj2Cy
kurfRF7yGeBDnr7cRc1uKGukXqg/ZTW+wZ01E7EfMRZKA/2xGJKpCE0jIoZR
IUm4n/27NXfj+FNNpc8gfbJex2q78Vs0q0EExL1K2lugplPSwy/l65MaIeDr
SRjuO9XHUPOz8g3nVP+jNxiZ6yocWSKQQV2nLoyn7wN2ZdMcJHdSOqoKB1QC
+IyZgZec3LAouDtBary2aEXqyJBnA/j1Pv0qMQksjLTVjrXE06gu/fL6mQhT
LVHm2cXVuGARBGLZkc7kMVkGGBXNy6EQk4rjc/Z5b1IDqqtqrhEIt22D+q7a
pCDDJrDtKlzF0Pi5N33ZsWkbb2qW3JkysMX9UeGujAKlRb9Re5vmkZkZuIw1
LePy8mFXEQx7jf2fI+tinDpqVoJ/MhhPx/gQ9MzpCNqs7vUfBLnbqiRLoUrp
1/NjD6QJwq2bxiOwgN4T8SXD90Ux3t6cQYMJki3lx5kGlAAWUNo52jSHrCQv
wePlOqgrfLoUWAt3kzfCeNwA+O5aj4HTPJ3hkN8+pBHNYIPkuXknHxK002qz
9P91yF1OO1e7Kil4A8GEex1t+A46n1wA9oyK97rKNK8Fcs2l+8kEFeEpZK4W
jnh5cif80nix9qooDyGKlEg0vfCvcvb1i0MWGLaY+SydQsRWRIG03uK3NKj4
4NGOTOjs6Jt1OrQQZ9+KRt7lSxMyWZgBBc8wGJNflkEgDsfYYtdzNWxKDaei
zkuARVTTJYG+lYR4Vzlfr6NCMzz/ADgt7bKDxqLSWzRdLqSSkd31Fjdk0wQ1
lsDXUgvUHopQ5ViXrZf+ahhcLUxwE9PR7zYgqvlfHKspV41VUH7hvKvm5Tcr
U71kemrbT7jhLADRo4yB+Gq/hbLxcRbUs1MagCrAOE0s/+MgUr+y6ePK7TU/
E9P7xfa7Zle5JSDr5Rlquid08H+vhBeHCchgqxwzpDYZtyy+MUCgOT1Es9z2
zjHns6lQisRlPZ9kb7xgYkhQDd1K/Lf4IVY1V9Bv7v7U7IkmyRGe0QgMGbv1
9cOT24NP7DitF7fwbXuEKfYrcBpvbGMK7e4ljfORMd5Mz9SfUqUsngJNp1dI
RGfLECDVA4JJcEHnItCPCajzVo3qUj+9QZIG50Y/8GK6aaSTfj6t5bxNHE1o
KvFwMfCzsw5vaqKAAIx+8z0oA5p28c85mL9nUz47+jLgstoDWXV0fkiXWNeI
WCn/wne5vwO3TtojCcHlpX59OXfzs+uQSnkkFtG08yiDRO/eWbABe4D1WQ0j
zAIrXzFpF0BeJgi8wdHQAhpex6Y1Vhz0yAkNE8BgeHU9U3SB6h4PIk3FVhai
aLs37M7YBc2abUNGw/G/llVdm8Ro0SxqldJGZPmt/mQJTDvD0zWHHP773BQZ
aHQ5KlfHyPwC4o62EngaggILl2LCAQrtb8h2BupXdt5KJTMUGGq40imm+Mi1
Cow6w5SuuEvWW17+qnZqMi00H57YBel5V9DnSGGO39hDA83A1NVD2eUsEn8X
t7CL1ZG/eWalIpTP8wdKclWGuEPeAN94U8bKCJJUrgkrBNvXjt9Kz8H60BRZ
KfJfnrPhlUrRP8WxHRtUhYmUs9hNlTV0ENNQXHIRorLtO/EwCxIWMPis8Odm
HVFsgryoUk/4g+0wa13+bT/VTKVODM3aLT5kje0ARvxqUkahM+oU/PX+wTA4
8/HkauPxJgsd7wTAvItq5ENi0avo0ASNvIRtbX9GVdPdhKubVvOmyn1SqeG4
0ZnSQltfvJCq4STNI5s3gIWGzjwEo53mynw1JYsjN59dGldTEcy631IqlkMo
WpVOjVSJPtElS8g14XHKGurrPTP7PtN0/z03fJlEYJdkTDZRFDh9sCiCB0OD
Ri1L3PNkhsUkfY3CagbWDKkVWNt0XoI+gyDi504BD4lQBnbx3fToF0oNhj0z
R7y17ufOZ3n/87FzJxDFEJ2dQKVoK6vTX2QBzrMSp8kfDMMpk+r0m+PEOk2j
vtKhsqYGgWE2tPvCv58BOpP50Zr9JwlIqVXdcOUA7yskkp8lPGL0olGZ8PVA
G0kukKeas6UqVn11/LHDYY16sqeKW3oBnxqf9kCaqtO7uAkm5TTDPdPAaEp9
BzQWaHqA153RerdCQMwaXMMWOWNXXt5rP704jgvgiLbgiYLx567Ck3U488i1
6HEheRpgdFqpmzmaVH6+AAG9bSs9EGmsK/Yeuj1eWOrr6IXSflcePJGM3uHA
iyj3XltQxSLZOLBVxuApuDDVdvrsTBGn7LesQtL1jMUlVclWIAU69ilOqg6W
XO/d8Pq8CrGjcTVBMH4O181jUsTnfFCyA8py7863J8YsAHz/igHIY4kCtCV1
arSMUz6+GoV+335bnn5v+G0LeMCFtl9bRm4emIhJEs/QuuX1QjDguhTfh+Ad
wJpZ5OaM5oGIASo/jADCbb0hN67ELtaGi9vsYxXy2W6Kpmj5HOSPV5SvKJFb
Mxyp3EvA8XXeADKEd7fjCnjZzmMpF24ETTObZ7Id2FGnk2eiZv3JJbauchEe
2gsid/EDdNoJot0ZdkwsmFwZ6OuDxguBh4pemO6ii3RAJ/sZVyotd7eSGSop
LuXmQdZC20E4t4E59xyQGTCnu5zOzqS9kV4roPR3DdpZmbzTrsDyg3sYFRsM
jffCuQ+sRnK/PZ9XFOs8pX9vd7qyBwaj/bYg9uGjwiP1iEIbVOEp+Lg1yVkw
wbPsQKCn58DXR8Dx3NYrwW/RykT8eOhZ9si0xNyACGILgzILenWwEi9oZMDU
FZ+9t0G+vrFbg/eDstLJAMqqOva3Eki1sjah+cXwFy/fzpyGrXMWyD8sQ5mW
oru9A9m4w0MEsLRWIyiqhk5/5CVSi2gYLkHPmGNhNG1XOLvTluTjU7p2yc46
K8nh1xuQGiCGJgz3j3eWUXqYYtVI0Fv7RRdYuX8iwylmeSeN5r5b+6LNkzmW
ELDTeSHiOKx4kqb9tbDiUaC5DW8I0D1NXrQy+UBXtoxdccRRbHqiaSxRSCSS
r28xypHEstYcsG8KV0gAKsLECqHCwH2IB/vHDWDYqNYnMdhkcLEzgwmoCTkA
8DmF8PvDhoPRKLdNjygN1Z/jEfsQJjYkm4cKXI/3OR5ud1nB5P1Hr8rjTcE+
5tigm7fQDvo8qK/uX9btXSi5wD28VSLli0ijdtgjbGqmqcX3CIyBPJgo1Ypw
8KEJ5b+LV9iGbOE0GQ9j6RIZdD4z+lVhnzHPYqlTpnrEr/Sf1+onrdtn/I2r
hl03ldH6o5Uvmhxn0VcleFKDdMceWHxaZlinPmz+QEB1DS5PhymOvCWIBjDq
EUsKbe9ewpRbfw7j5nnFoZ3rL3I5JfQy7wTS/td5FkBsj3OsgwhatCo+K9J0
wGorPWs+qFmWVrfthioYd+fkHW9RwUhCwFrIIthC11+SL2W1/inIt2nyFCZX
bO5fdaoKVwyl2zTLsy6MfWD80f+6Rc2Tb9wEmzpPyMFNxTIQ86KhppXPDI0c
isPDnRz/qa1SVj6Tvz9pFyBh6SFkasCXD4BYldEzohsEuUGVVXncIP03ekNi
+XUO7wnPFhq3GxyDRAAW7tT4ryXhg2SWVaoTtE3ODDas1wJEwgHQXliY/CxH
ni13X6vtWSkmAK3ZkcMwk7OXGrL0+wVHcHAaR9dWB1l16dDD6lH3sVxGD3fN
jScq9MXxX/nce59jbGylBxiNgq+FJVstJpToJE24jc/Ont4fHCy8Fgpi4nog
dc/upfhdQKyqo/TLCeJSxWEEPKI3Saq04WHtmmxJN44rA3jEA8EljOQJUsFz
Q6Hgc8wsLLXezVmhxHQzDBKU60koCHyVt35EpoO1BO+sEBGktBSzMkW2HVYS
fjea0wEbzqnlhCB4seJJbLr5+tqCXK90iAbc3fCWybezWQpc2n8LE5FJCo1i
qloHOY8rN769dY1/IOxDrmblQNqkR5NsAf9vw5oxiEpIaK0yLSHihHj4a2+O
GyLKeSD4XqshEZYib9YMcuKkNRLbHal6CznezBn7hq2I1ZgG+f6sN/m7e4Mt
9tEm0+wZxfg5pGqxTgJsXzEBT1VPSCzLUJhRSQEgewfOJywt3FMqkWvIiBLT
7+FgzdSo942C/KQC8vhYZMz1c3/11P43+Pjw1CvsOxYNVc8XXoYL6PRosZqZ
UJzd9O6E4lLWgbd5zQRfdnifJsWrZAmL+UCNqkBYOvrVIztV1BkQJEVbuhHH
cWhSHrxOpkPFAtGQpsH/mCjjc7efbzxwPhXJ6/S5Oivkc3BB6S5dZKnymq/Z
X9SxrHUzvVxI/2d5yqxN+DeuMh3tgZWYaTHQ4dBgBE/Bop4oTv71V+mc9s2z
maQLvKtlStDwjV6xPAtEO4HeHPvkS7EaXQ5kURBhHtDk0pbEFui9Ld2x9yCB
Bp3eugZQvbxlbiEv/9gz+TdmqalDmEB2SKaNogy1Q4/UVDCXvv07iT9PbDvv
KW2FsssFTAQx7coqg6Fk0ZL0ztJp0p1dtpeapZbSRfEgF3B2vaimlK2q/ymH
TZ8z50uP/CwNuq1IMC6JT6Asy/7VmdGFJxMqOdoCT+Xten2fot2hDdcrB1kO
+qCkdOHuoRWzlYcNjGGQMTyB0KDplQRhR5tXHh/dz3ny60OA5g/3YDwuf6Cg
P0nwAw0aMhZKBLZVp/iiMfrblEY+CuwOAl3UU+Fhnghnfnp9CWtSrETUgihQ
JYIRDJBIFGKZOAhIE/gm8ju5rFJCoGjWdEa5ul8i6APnIIeX0op/HH3oonDH
tpOabZWFmqvYFh6TZiy4LVkxFW/ws8/2g23sqckv1Vp8qC+T0A+FGx/rpTuw
iTR5xf2JARZ2fZGUeJnNoOdOvwoeyQ9u0IH25t/ReqVktAHdxjM8xOJAo1y4
MFrzIZ6Rqh6N+EhFMfM2CqgKCik/Kfj9Pykxpe/nvTZPXIGugZ5SI+rAwu/Q
Ph8e5/j9jdLcgPmfSw4pjLzdkcUIFjVglL8GtJ8IQR6LHVJMn7WhKD3TaUNP
n6dv+aCx55VZxCNPfgyT4uKtPe2GD2BQMu311wrp8Hu39fxx0z7ASEkDhBiG
LNkvw2UtsN4asPQacPRwsmkJTCAaFogsFqMRER+7aB08MOFUe8IZVfGwSZYg
/BTK4nv5iWmLJm2ZXYnRRzKaKuzjcUaec/4X7R43WA0SDhMyJkD7IiREIbf4
EQtBu1p+4O2edY6B5KWyYE4r7xU9qM2pBT65PahibXNpt6ulq43es9zXN29q
N4sYGKIPZzTzwrHtUZSvYxu01sOLa4yxzPt5UZ96Qtx0L8YyPQwIqMRzn5rb
xpxCx+ZRwx7IIwdn37t87x/Q6jefPKlzIworU/gYU0rS3/67qwyTQ49NoBSG
B9t28vXeuoyKeqwYy5Rg3scFhxHj7LTcIQ0gGiIDRbU0B/a5xVaSbZG7Vx7Y
peQvhd6xtooVi4wJsGclXicltj/is+Qnt2QXgJgx2bg00XXNHs/HndmwroFi
8qNpkL/HnQCjbCrKA4fGlZDo5su0ZI9qHaYl1APvYTc8WC+OegJS3w5d70o8
E8ow2ctMH6jg7Yf/oXHivvnnQeEM28uKa9kMp0mhCFPExrQcUfiex9++WmHB
i3hRwLaAtkYWxKabEsZ/q/NCTOlf8+/AIYG+TXG9VG1FEK1MapS/JYEsV465
tZZmbbqNgq8DCkJa419jX/OkWPe+CAG1uhc6PScGvPis2uaDkNQN/kRwccfe
gehl6/wbrYLmeHYJtkdvR6WEB7ryXTo6LXZaHaY1gbXWrYWRRfAisTqddVvK
0ufYRSheDOxjSbYlx90/xDbUdNamTj6cfl9gj1+Dzed/o7T63oNnTTyJgvYG
z4k+wWA0UWWarfUmFwwkb6k4XAtLIYyMemI9VkCEH48m/6VNJ2H7PpweK6gu
eLdgOmGVA/3U/WjqiRfNNH52iPKM2a1JuXxV4bkiWMEpFoOY7VM15KdDkC+6
whg9IqXqKGneBLdUT7wHng7jfT+QnoeHV409J0QQoWbMGvUcaAwyUB+ydqbn
WEKNNuS6WfHmb+jmA6rdXdFZrw/MmHKG7qvAngtTGfDstNmTtc4G0l7h4ISZ
CuC+70tzjRlpix4AG7OVXgol5k3mKyug12DuWrZ4FySN155SjtR93AAbgo20
o83IO2krc6Sxd9mBFJIOeag8T2+N2cvUw08B0l0Yy3qxVSOIlBqSFu1TE2lH
GkyEAzdwuBuDwk+qIWlf5kCOHSJX8edt/WWC5MXGeQtd9QXbWKxXzuLbKnrP
K6htwdlBLLfA+mO/g0F2uj3UbsSmAKMq2lWwizq5zZyUHqWJSzQIg3iKktxs
HDRx0OlMh94XdkrjgTXOxOwRU5QmjnOfn6RWn62/5YVixekqgYukZo4h3YfW
x3pw7dox0dR1DDhsrAQXdb6ZEpj3De1HwcTfBTZr840C2+9dCZ0pbgiIGkpN
nVPsLDisMzm8z8h8OjNIfcC6aIF+r2/3CC3khUSQBlepK0rX6pinOqwxGjXi
TjfMt2DuwfxuYTGln81ryzH/i4bPiwgAI3C5Xdto2J6gvO9jnp1S0zrvksTL
j8kcR0HMu3fbCTH6UaSemBoQ5SFRdHmVNBm2Rj/3z7gGI2JaLsAoBfJ80GtK
WI4V/VwTnY8pCTLjTkRx70KD5eUyX+5FyWSXdgJSEHWNz1Zkmz8tWe6CPRdB
7YSNq3smouJezW0QnheJFmFVog16m55z735Z4+JrhdVyk9ZniyTgSiuG72pA
4+YwFbwaX++EutxYzJwFbLW6XZpfITAQMtcCPf/QkP8rNkDENiLi2gfSY2lz
ypMWXMXmVBVNlS4WFtxJ9Ii72V+fHAZ2OD72jkxvt4lxSNjln3xkNhDAYnRO
/dvC1XMKllp0I5SelfzJXIS6ej7RgRFZ60rxXuUyROA4k7O1GnOQXCV21CeB
ukS6wuxEE6F1mjnSLxa8jWHnBadkNJ0CRV4pHBrqE0g/PkcDJEe/grgskwBJ
8YYdVn9estc6fj0Q2vAfv2BizLb1dvS81Ih5HHwkRpiDKKCogPgePCKa+E+x
v97Ha5Vzp4yikyScMyVJfnD7uSi/zQ+G6/0DpB2BYC+rJuw2OZRYn9XXaizQ
UAHpL3WQb00DKkFQHRL/CsrMleDXPeNIxXGYNzOwZh3lfCkVlTFcIxrsX4kX
AOD68D8O7WseD6exo4VNrLnV+Dd9BvirmEIczK5SyzXCEw5T6vVMfS5+tCdA
Nt5mrK+xnOXoPWyHHLvwweWlQ5u4tSRVPtf5D9GIyI4FkgYyoV+NvahOZGDz
MDkVXHL3Utvryy8zKsLbhrfizQylMkhhvS8rkcWEF4uIrkjYaR3wxfLZk45h
+Ruel76L2CtI2UPUHGEl3aME5fn8aYU3KcmTd34vTrrg1tqlrFSZIUyKQABn
qU5/KurtRegv+dVbylWrTne5FfBgXJMQ7mn3IQ2SLVq7Z3T7rja1idfa70Nz
ZBjUy/Rk1e4gtdxV8B1juQ/LWd6fbzyNdd43vVhjbFbP+lZrQG2CkHJs5imF
TezcazK/p3SXXpqIqn6eEQY1+BQFZ8FxPWm1Le4GUh1kErohxMDVmSIH1Z6e
MR8gwoo4oUoCYkaVNZVFuEVJK/i35V9ASoO8gAyDs79X4yVAVvB2uJXTaXB6
7KDs4KRzFVGgFXkdpCi2npR1UNGa5xjMklCdkz3rCcTur78DrnhWtHMdO6CN
IfJX+5ggghW+vc5XAeB8YnBKRnfwrxHg38FHECwgT/s+4XVtLX9dsyemGHHZ
BkV19h7mrKsqbzJTrc3HljT3cc1DOK+I3Zo9mViqBqBIJs/fxt3xiLJGr9du
AFBaCuZavrR2jhoLXMVtOBcNb7Nf+CArnuBOYj1r3cMSOAbwZwzUimBYzW/F
RlajK2I/GxjQ7Qec8suNWgHayKpawyYd9GlP8Gz05pXU0vzT8Gl41hKzlbQM
G0vfeT8XkjROcAQi22in8OHxGP/bRRla7TmGaYO0bWqaFUpUXTBNoK6FN4/C
PNEEMOLoM7L2rKUddqkO/0ILf3RxMjW6e9fDtBviO4B1CzBpSm6RFXecbIi6
SJApkNyjKASzCUwCDVVUZs3bNtlE3LGeGCs2Rz573oH4jgZD8bWNSfjdF6iR
MqS5YBevrHaiHfLwx+IldVCCwTv/TV5TMvrrHaQ9F1Vz3ZVpWmxS13AqmoqL
XbbplAvMJNgXjzaayJVw8xkN5O+5W4d40IpAqkNMOZ82CGpmI4IvDHWyCs8n
ZjT0a0DVYsgYDpvwRE4n9Sf89NcWtJvr1YW7woT/aRUHEBFdmFHS1hCU50pO
T2LGQrd59Sjb+eypapbeEvBREacWoz2nEhZp6akgRSHB4jWdReF9cEVfB6mF
Lg8g5xJ1WkK5E39iJ0qdCRsedtGhSPQ5x6Aai1dzePqU6mWr+hKMH8rV+iyd
q79BF4JBX7qpn2WwzWZEKt16JqqMa5jKXN7fqMvah4tkdQ50EUsQfwTeig9s
/PBQmfI7A/jEVFgUsCoKuW+k1j3VbJ98t7nh76icORYoIG637p7KVv1M9ROJ
pBkncTieRmpe1KE3iBfO9xd+CST0sJXGfOHffLzZOO0c7YNffEEhQ0Ck/+jt
9LHI6qf+UyixFFYsCUebK3fzjyk1x20NRbz/a0bRp0+4u7YN6sjXp7sjXYqa
fDs+JfkT/ZP4daAG31wxgQvnfqLzXHqowxGrqSaXMTuAY5YzG9jDENcY/AM9
EwAPj29UEH1XMQsSSW6l//1C3ER6v+EZnZywObplYWsCcGZAtMwo6yFTMOzt
QWElGbwJ25bVvDTr2ai3flIf+aM6v/g19+H+jo8Cf21WGCE9yLiug2XoMHz7
4EpvdkTwkqZ93Bj4a0qa1nCOS8boP3aq07Rx850Ie7L4BOmM1orcLD6xtfZT
Dhtbk3pu62U1pauVvMR4ikR9YS8FkMUFHPJDoUGz4fwwMX+cSkLktLPWx/mR
bhSZSUcEBc82mihNBAyiHnc9Wggie7iCmpueKOUj1Go/aETWqTbCVaFGF2yZ
QDJoS46ReoiNgPXl1KYEebqr5f9KxC75tsHc93vKlZ9eBstDVKyjUqpX5Os0
oXt2Fu0h4bAZYHEZ+G7JtKQR4uTREfARdygMIFX1AnNOiCvg7T4TxOI6Oj5o
yji5yYTF/9fvTisC3t8IAJEeJW9tdrgpTYC6MVh+kt3VXBNnRL6TBSCliyWE
8pQL/IAK/7RvWVmJ90Lr7ZUxOY2pRND6FeQct1reoAsMSmZ78SoqLfLrUx4b
fPlqrhYyAfkmKZL2HLeGVn1x4nBPWItXlqi/vQwjYMlcaBxOeoxaV46BWrnA
HrBilcPbO10wCLmfO4n0ghxJwhi0T+oHlyAzAZvAvRRVq9+9M0Q7gioEWNdc
woyJDxuUarUES1AdfUdQwISz1ASRnW9oj4F4aUnpfmkVZ4JQzwz0RFjgv1TR
7QbI3xCbh/Ix/TvgAGpEuwtmLH3PNkFVCWdBp1IXoi7rNRuwDnS+nRamHMOW
iAx+15blaA33tvyOu1yLQjNQsI+T/BGJ4tYJXFijntv4IUUnqkQQ6hNh7LxJ
4A0TtW1To3H/JefK5HXGmwxx1Qd5P8PfSpGpIoPpnUOzG3KXKsUq7vHD/LEF
ZckPczPuG66QWKiiFXkRcGQRRnyG1APneFFHLfsS/Dj7pWFDgl7RwvEQrvWY
I1KhFj0NUqbUek03r6iOxPZiba45mR1/bs38deRp1p25wSD/HiqCjwawsFtz
/BNEZbQXNwHGLvhEw2ulThD8qFt/gX5Lmqdhs64MawHM/myiUIC5NIIfd5PG
pnBxkr2jvCE9ePHUXCRbJykTxgfxUrebAKZOypfj+G7RF++3zHuOmmy2kJs3
izhdB/MsDh9CL0KtkymIDng2UrPPMcRTz9K8sia9vl4x8oZxKcLRWfoCDT+i
1jJerQHMB0auY2j0mKGEOoazK9om8VBg3fO42wp86weAEptII+E+yP1KOx88
pD82WuSv5iYtYCIYMx6AnfOnOZlXyjaiuN0oetMNqz++O1LAk7JzmjZ/mCpX
ONgn6268sWKXSCiqvCHJJI2GaeTTpDy+bd0hprszZTBUdvNcNkE3uK0NaBLh
npEzLUAQh9a3e6PpjlbnwPf5XLGmnB64HLBu9U7X4hGLpIlaU8gw3TVDjlta
WJbqGrRcTxhziF9XaDU03Kk12ztX7m3fLNyKOyD5gIees9kAJCdsdCbAJq7J
Nn5avUrgkNWGZjU1puvucs/YUiWo24M4gx/HedZFDyqVXzB+scd/UJc4Tnul
QcoP49IY50DgNZSZYKYLcemh8/NYbxm3tcYvHERMd02Mv3sVoSqjh9jgKDTL
Bw/wNh6tKUoHjLCYKDAvn9uSyxiPRS9efwmWnp5ox1m6c1DOOPonNJ6zzHnN
6hdur3005nRHkV/UYJykHRjbqnHJ204/V0/b0kkSglFIp64P0OQ0tjcV1k7O
lm6o68tmpIeyQrDIRD3/tgSvE9mEt+gZvm0qmZ7I3jouySf+8tYPG43sQNS5
7L/uiyNeY9Z8g5tVgcYl8ot/1/Gh/+/Jn/2YYYmhWtBWbNaO+PvSmOR6eu4m
7KWBG6PLNkRXIPZvRlZgJGhTSZF8BROxZasKJB7OMI8jBVu99XM4cSzUILIq
WvO0Xi5wwiur8T41yJVh+JpybNmKDMfuPHCcRD3RUtMH5UvtdaDEUIfp/kaG
musOAsHdeZBV/ahxTKAuCN42VWxXhE6wIUKOA9qZ855ktcNjQL/XVC+O9v4K
L9jjPRYR0jrk/+UWY8txs/526uHc7f9Clia7/b+6n1Px+EeQli2wpf0iN1Jn
RaeaXeD5jgCVn3CzXsbowAFn5OhQ88xA9Fa35kdcNZE7/pxc141zkQgOCDJn
DnCx4aiTehAJsk4FN8sVzzJgm56wAkr6bAHiELxkITWt/5iuNnRFHg2N++Fv
FrKdIxgL5STSEMAr7XEZW3I+ELZ8JOC27tK0qbG6R0DUcAVcvt8gpIEO/pNe
yU1tbXTVChRIxh2MwZMJ/jpZmzzBkJBOblndPJka7+eVceKWmWuyLFPqfiJw
QiK4DUelPCZnDgm5WODsc1BaUf5CjmaVnBnoakMpvc4Umui4YmdJuqCrzJdj
kURB5XqRkzpphPX0ckXS59zKwf1/9lFizsoE0juM88QM2kLodWq0me38jfwq
3rCOqMULofUTlDYbTE4y6VhSPZr41rQSnBxoafgpFqPnAsVQv0KOR61o99Fu
UEuq8czq8N2106fCJ4MMwnXtASbHOuJJ+EmEngen0r0e9/7ynBZ8lUWrF+39
DsHD86KPluan97QOMKi4SWWt+m2UsJN9M2rquRg5+RGt8DL6nDTTw9oAEaKN
vPvu6fNpW3x8MRH2/Vy5PAB4zcnFvGaHQZbmmFo+G2xF4T9AgzlmKTTo6aVW
86cgmHhl/NBs2IhG/ofXmc1dn/o7u1K4l+ulOBmsKSsQvODTn5vKcp67+plj
yIOS/+cNxBlGRbi0JgKGiNnhnUV5lS3+ViUFPrFHBK4rkEuOKI4vFEV8wdiQ
0Bb+w+rDot52hklCgRndaWlCuZc5UDv9YkjcP+wCkpCy+6JNEMxkyiAmznk2
NBWMjusydEuHM1jS/NmVupALHLz/pk3SRSxnh++HxnJ48za9K1wvimPqsY9g
WvCqVf8kjAoJnerZswcsMhOBGkX9yaJO3KP/N4eMQIweTY+vZcXmWEnzYwNk
xgZowtpkWjJ3ymKO8kCREBOHs+AYrztk2o2NACikFEDQsCJNYI+xHF3S4a2E
91uefCo+JkOmTcKVrHbsrAL7vTRRBIri5PSzLWrhVfVXJvgnAE0D9nDRpbko
nlL854bXIWCAfQ5rDKGHdxqwuRxXaY3JIVbwIzrZg3v3gmpklwt6zzffwZQG
sgMkXpj996n5InD3Z4wegh4h2M6hrfe5WPxOqyUvO7eGobG4RUqy4UWYajkF
jWk2OgLSd4Z+Xo/GRJBCMbcc01L4+gTAvQwWvmB29ruaz4V4mv5i+qe61LEe
yClFd1hQ6OuWctzZODRC8CeBcOt5+Zlnx+AeRQ+Fm3DMjnB1ZAAZYhluwozO
T3c2hAIowbh54rbgQWclL4UPfIvJL9Tte5s3pr4uf5K24D3G7TY/cdnnmbNM
NViEQWNA13zd1KEpG0LU1dxNjDz0tKe0TZ299h/F8McHkim0sKaBU4sf4qvF
FHsPoH2CWCGsyY0Qm1XwpP+upiVmoFV0jfUjiEuuMl5Werd9PsdenZIMgKfZ
UvVoG1Z9+1RzWdVy9XVJxjSBzZpE1Z5EmC5yv4jO0GXCW3msEvc1ttpsDhw+
JfctUOAl09InkK256/n2AYq+dU/bBaszWJ2RZbj69sGcygLT3KPnyJv9/ohQ
V/MwDwTPbMwlCb7gvidIKG/C7QLlrpvmm0UoDLbQgSh1NTNsF5wQMN4lu5vs
ZWa+0Md9BwhPNd2pHSh9864KqLsDkceeGfRpSvDqq9Xl0t9G1FYkAytqhUj4
VR7O2OFsz0bTtbQLn/tH48IuOxghwroOhnuc8Luu5mMc6Hvp269QoTW51J3Z
oVSP/t2KLdvAA9lDNKNfImqms+iUKua81EVtTEmPzJ6v+eXLRahlmkIqeKjT
2AKJ6B3prFbovuMd6LqFFYcrmqxm8m7JYxWqp7xYr48u1+/5w/g57MFh9soC
WRcYQG8MPPtZ2ZNVMM4zZHFQjmppQHayFRXGlNws3dqoNFXCPpcw8huiaJov
uV1YADrH0AjgzWAyBnp0CgCuz0hR7+ho7i57vS7bITDF6Mfmd5mhbdRMHqFa
wAvTpSKvMW6cwdFJkCMt72XMabH15gItAkP5NWfUIyCn2EqMfeZcE66Bciup
ts/nUUT8TJ0tHuZqmLeePs88cEXpTl07gZ4hRKV0jqbZW2z6AJLUDpp/iSGC
wCypI92QpMJmDbntDrErmODcD8FraRD9d8GErg8z5wVkKXQJgwq12hVKOq97
NAUigfz5sexyZlq8TmF/T17Aow6ICLPNKAPh31GTTBhNLLLG3Fw7Gwki4kPR
9x6cVC9173rHuyo9FKWxDUoY/P4EGB4f5tdtGeaia7C8EUx7AIQnYSLGUSpR
O0RirSVryMzhoFRmwP+usYqq0VEVHak2TNYJ0gZde1540DASRa00O4OB1QDe
HEWWJqVwSSMMJ9QCm/Cjgke8c6GaWHrkLguwPoSrtBoBNassfCBiA96ae53f
+FpKF4Ci4T4/Bu1VIIl55xkmFRdhQ0/bDpwDj4zFMH4aGIe+lusP9DkrPtrm
E0eTjfVoBtqQgHY+J4KWTQRmu567y1kmfHPrKX6qTba/DwlmZhdsVKwck05T
dlS6je11/f+49Lyl77nTEJ9TFgJ5aM6bxZvVhfF7tFT1un79KHxP5wy51qWI
uiv5a9jANPm5xD3UgiJeToShAXXbHTvpG5Q8AMRveTt4jzIl+d02Gjv8qLRx
RTsNvz9Fcef9Lrc3QI9PP39/h+qOJ5iAPtZAfOlaAF6qaEeuGPtdXabxjspf
sGQbTEd/7yNfrWkJDuEXWfBuF570TllrH1y/ddZhMqjQisBxS4gxmZp6rgbY
oGRK4JAQh21pTB55PTjSOJuuRhPRBATABGnpSo973wV2B3Cp1eEynvoAiw8B
8Dp0Y6peCvdFceRqEzH+ErKpsSzGYiOf9oubR6cjsBApSEhEHXJZJU82zwEu
7DhbLoBT6o+JgxhYCr2jEU+ugH/1vJ8r8NxMoy/dklNc8o/ZBfevHRLMzYkt
7VQgdhDB6KMSzVkeoEZfAWIlZS1xJguOOR5MmPGwuYafB7DLDLll6eRDEq7X
/EiGgfdBsSWQIfFZLzykFE+VGZn9viNTK3zfZN7z0bJQFxAbFguQz/g4lr8J
1nQeowG5Yj+TEVnjSWUGEfe+GHJuX090t7BGc2NSkcgGtu4yp279y6R5Hn5m
2OuWVkYL0fPaOP/4eTWV0EkaAMAvSSsMXQ/YuFq9UpXv047VF4UNOA6ulLwx
fgPb8sH2VtyXTisnuH2LhCpb2/YY24a0w8lRlPHs/ywLOUCsrsluOTGIMVT8
XHIcKgxw0I5MBQ4jV9bfSRtuImbbslhLM0DLjydeGMmxvPgF9qvlwWZ/yiAT
oo8bI1LPHanjG9UVmIF0dy7uz/y+DZCmgEXrGKAYeXlvkdMybMJOtcv65KAz
z5J1WpFdWLIZp+tdyDdfnHMSZWXhgJPQfIXVXalWxadZRn9JmaZ0E+C7nFRj
qVI+tin0eeb69fKTfwU3bw+uyy5/U+3OK5L8EJqx00OqvD0CuEv4l3K1Badp
9Fi6NI/MVUby+wGII45QUdhBhcx8CRoLJrNKdh69uvrxAWBk0zI7lhku9Q81
AOM4Osb/yYFZXjGyPN+gUGAq1jb1kbzBruDAzHsrzj1XFQQC+pgl33eDQlZa
dy9Oc0dZxFRCezlsmoi/rPD01k9LJyFHSv1ySNqwwakegxfFdTkbpomJitgH
jL/T533ZAoFPeBu1yGB4mWvnJwV2gCrTyKyvir0/C9eqioV9X5XNLzmn826o
RXNE3yvdHOKd/WEcH/SEdRpfmcd+unATVg0CxO6vD5faDtsaUgHYqI5tioxv
PHj4lDamJACwZtbhhZGr/41iUMdll0x2Dx7h9KaZEsm1HdM7zIksBLre7DV+
Dkbq8+v49OCBSuodXXuMPD9JmlhIDbB0A5wCUOE+1vN9kYB1qCGt4/97jAAO
O3gmznvyd1L8w4umm5ROf65aIcFY0qqyCv8oGPV2SSkaJT+xw1E19EkcOsDf
TwY+0AmYVgb6xRfU2tiMRJMN9D2z253fcICAFOpExs1qkcYztaNdhd+FRVIl
e1IViNxusHUsojwE7u54ViERVWazD9QphW7KXzfVX1chUy5eWw4pfvG+nNoA
RwioW5xf/vZGSTt5t9tH8UuhuEIOgHwRZ5FHIU+nvPe20CztJhk5WnxdM8Sb
JraRjH27A96JbR+TobiGehcqr4BRIWz8Qu1uBxO3HHGz4asfIQ8OUW7RNahb
XHkqt5XJAxIqlK97Ikc4+JN+6TYySyQeW3hl/hMPdBZSdY8WafBysZEQxXCm
PBSc/QtE8u6FAitmnb1osiNavkkyFJ5x+0AtQNS9KVwH3WVjbmknKii1bQVv
HbCagv2svCW0yDDWrYpTzE5sSxRKzZAEAcaLd5oFrxJjfCaUzfqgoGmZGbAZ
fO9FCYfV1HvuS0rXxl5pF5/R08fNz3K0suK/hN9Q7BEOo25IpLWFIMLP2jc1
FhridPTUjvSQL6TYJ3ofDr8u2Oeie4dPXY760OcbcsuAT8DLUZsBEQzWUtHP
Sy7P+qZ5QlYygh3qiOwJnajMrdwf+UEFZwA+EI+tJKWUzgPKMiCCMhBnWXcM
mG6dGuok5G/MdgcH2W8rFHngCApTj0UzKAPGibIzEb0geALckzwhUaPl27e3
f2jLvbPGTBeKF3aQu/IUe/sjgtYbfL64fjNxO/ZSChmPHJ/aOd/8ypu6d+zb
bW1Kz1KPo4nkxccY9iX5H3Mo6Q+u1BXH25RYJkjJSwyRNyNgldHHjpQaGyFQ
4pk1XeN5B6XtT9GYhrNm9azar1l64YHheMfvL7X0HmSQCmIcA6r8AvSrUUyh
K8qcf0TyHuSxrSWUlTrnt9xLC3vIYVjwvTqjYufc7+dQvH9idqtpa4Fb+EEv
grXjLmTGqOFtGXLkeQKL9Z5Dalsa0Gaa9xOfuWgizvlogt/IzoGnT3XSzerX
RGGNxA6zbK8VE41ZJyK4lvXametcD8LzuQdZ0jtE1K4d9eZ0PBqxfG8A1Uee
kV1nUqiFWxqiEhkPYHSffQpAoklEvkeGn1k1PbjTJNYBu/W0bn/HfbGcFU6o
JrJJVuZOjRR5JmECcoTxauXFZsWdO3GnBqWeE8oJ+2dzSA0a6vJpOVaJkj33
aFFujE59ScJ9BJwxrJeLmbadOggnXxZtl1nr7UDuHjreTnLVtSvBPLo2t2m8
dTxKb6YtjXC7Kj0d+6LhUa8Qo+SGheOpqSzL+XwImOUCRoqecw9APFdwIkZz
B8ZWA6oGBu7HvhFKRU7k3p2lEONB0E4XmmnA+ZeDm25ogQWChdNpfzBPKGQr
a3k4FmNELmUqWV7pk1v/KqJhUUiFEPZBp3TS6U+d6qjzj/bzwOzN1xGB3qUZ
v/tO9aVVA8DJHl9QeHXWH1ckOta3sOf3orfNQ68qzJsatOmlCWOHQTUGQFNB
EOgZLegoxfbCqIx4FS/01+qmOIQgf4PL1Qy0g8xDZ6LOnY70SreOJA2FdO0C
LHTMMl73I8nF/Q/u3gMRcZDmlr9dioM4qNCjXEdEUcIwZoQ0EuccPD89AyMe
SaqPMlqo8Etfa7FWhgOxJUV3T8BxZ/YFEQyhtG5PAlcXmfk5hNnQsQnm6LxT
4b1glrWRshd0QT6YpAo7o35b3Jh8Y794YQoWNwvf4+QjQKrVtWwbFqdJvlGH
rMv1QlHiwHPFOSlVOvQxuvYuUhBppGBa+FVp5XC6N7d+8riHe5W+u/nCgiul
B1lIpLOodq211TK40fwfEtlfFiXQtruNlbyCfgi1rjWikhQUMWa8NQkiopvC
LpDPzWZQIzPCKXhfBtZ7jytde0OGjLMWJA4mOOo9LSVB7HvtwdQFhcW/CVhv
gQYJWfZrbIa7datg6aydFRExDE9MFXEngScchUOwjQC8tF4VinzOUlzRwZbT
7VgUxyvoVNjgaO8F2L6SXVxm7r+AkQ6js7xDBsaBcD85uvsj3DkEqjn53+hl
HHw+A8FapZvub1bP+96d4qU+wz6n654wbq16rFYX8zjkf942vwpb/5mwm0fA
EFyatxeM3KXgnfK2cSeXf88xSwxmVMj9BbD/exB3V9Wu142oJTNO5yt+vn26
0MNRegFejuee3ljm6/vczuOl3HAdc5i3wkiV5xaPINW+3brsh2eOvEnG97eC
knChPLPultsX6Y9b9BTJFXg1/BKPKKT4z4pNQFOaAcM/RfJ3rsnpDOHBLCSx
8LJF2OOlUh9y6M8nO4wy9BW/+909DmL0kGuHjtqaH4TT1CVHT0Zk4FuSeCwB
a8ChOKdDT3Hlgz4p9eccQC7dP9eU5i0w1fZmFrGuYu/7rIZP06V4cXZk9/x0
oO36P++/ViSePfLvIx+1AX3ORB1gT6nz1b2Zp4Fcwdwl4MPsQcGXOWPQUaFR
/maRNzfj1S70tUkLgq/WSTw0n5RhjTpX0jOYao6OV7iaEPGc8FslcM5ZHBei
fEbtwMG0+F8ChGC9CuGLZDioESckB+iNdZf9c+wvSy0PHb6YDc30S0/CiQj9
KVFoM/j+j+L+m9Bhqu2sR4jTN25QYFnvbUka/ggM602uOiKS9JBud5oLdHTW
rPb15SVzpWgDZ4kG/aQpervkAPMZdXiyGgTgNk8bjvuRZS81utr8tKmFdmnP
CN3k1cFtuYLaXkif7+Es2Duw1p3AfMUdArzVgjs5EeUOQbGnRy8On0Skj3oc
J2y58doLCvzOMPXM6Jh99SoAT6bZvaEXkx+AyXJxeJ6FF9wcNTiE7YHtPoqj
IK/Uv2rRI6o2KfZ9J3ooAGAJ75bK/QZtrXwpcaRQSBLUjfykfKgF20pd7clL
UbbbC6wfwy8RzITgProU9WatpTMskLXT1VansBvbvdF6paOb4Poo6ESqTDWd
gYBxs7zBMKNr8lOsX/URcE0R+AMj2075cnOHhmy0BLNYocfeDkISAkBQYCj0
StYqB+TIt2CpBSyxtpkHOkPPsF6/0U2fJqPLE7J7S8qFZt1Y2GRjgtXkqgP0
z5EAb+MH1J/Oph7OHybD2I7pNsWXJGRvrfiFbK8b1aVtxJSwkU3vcOE3+oDt
hvVjMNqXjVuo8iQu/BPskGAeXwin+ds8U5kvZ8ES+x930idjIMzcu9jJKdbZ
Qa3Gn2Mn7BSy+kEDWyHp8oMv61aLTN5uxYGECWppJWnYRzLrT2fW88Kwqg1R
3pPdomJZFvcAsVBah3SxrqofYKzPEOM5wFTKArwYcdtJAm1z60oWVbWZ2ZdS
cUuDVhaUZ/2mMHaG5C5Sg5N9EcXAmv4Dn88frOfrmYhByCCmRrDvmuc6yIym
mE9kL4wQBP1R2hE7Cz9H07FceL02bNIi7dH+Y0ynO2QCw+45qFQyWN7KkeYy
WY1j85lcxqITooZYUrXS/ZkqF4PbRkT7BaLew+1l0vx/rqAXvJO/IGUAMmOw
Y5EAOsVF8CmqBUgz3oeQsMD7eEHOTeD8UEAEo31lEr8OMLT7JFF5ie4IwJRd
NlG7cyrK/xlRHot3hDNT1EPpjT4uyfSfNDVQXoy7+ILaeMx3dXFBHeoIti6N
XaUvEAvRv6S3pT64csequsy6q9U6xYHMyGJKMDng+4aviRAsuL366YtCu/Hs
fJKOJUmm0Zq22IULqtDwMbMevCKRa7IYpgVIIY8gYaczVYc30b/NXQBtSnZv
sKPP0EU1R0M1TBFle8iyqK+8DdlO4oaQ+OwPU1IBMEm+61D8+iEp/URbj6OP
08Z3pLRlEBrcbYK6k0nB0PBMn3advJ5OcGDkpBELUORkzqqCsobE7fo9++2I
Ax0vctINW3rl5QH3rwj0NI/Zfgh4iTVavdofgENCgWTlYVxG94NOmYrlxs0/
BDoMJEj81X4qwDLh0gZTHe8UtK93ZPgYGtvqANi3FBD2Ag+Pw6gx6atLCpxv
hZwJDn/6JZjtwwVZ2x4nAPf6Kg4B89ApoImq2YRSdgdyTEkUYNoCI0VYqq1C
xQKVJ0423gQukmxcjTQpmlvg/hWmmN0rE/GfqR3MpvN0yBqp6E43U1W11BSk
EoSDBbeCUqYedZ0gKYg0nwTAQqEmtX8OKGbBPeyNNtmtAypyoSnQ7DymD5DA
TQbLFkBXTPxhs1h9szpLAxDPzGxWb8hIFbq/kRpK9UfL2kKnK6mw+LS/Iolm
9mjecKVEcw3w/ZWaejYQDsvYHo42ayZDGGFuJtdARUkEb0g9D70rskg4/GSQ
15OMNWTe0Z3DZm1lIB9ccC0CO5ypoDEKInfThWT83Jee2hBjlT42LKPXs3gZ
bIPkvQk29nj8wdxgYGswr7pZnPbHk6KPRXlltTfhH37V2Uw5Gv0VZBnkzA9n
jGDOnEStLPQBKWrlX4ifk737C9jtdrIjKmCXQ2F1/f3B21Lrf7msr+3SVO0N
TriFjns8zOI9v02OpwmsVpFMPyi8GUtGSJS4ao+bTzPxAP1TzihrkXQHx2s/
WduGiPD38gfwOetmb+hfYM5GHIDFw3lRKbOcwCzPaVBh9vCwjz7lR2UgLWgW
EiKRyG2vUS8QpcZjcJd06QzKrPRo/3TpczAZmZjlTHQ0yazdhn0FEBTQHCpP
eA6qYIGOPG7dx6A5JOutW+hjxcIr92XI+jF4iLeYOviLcEH2S4pSHyIbRHEO
pVo0wmI/j73J+KfzHyKPuFv+/a1YkOxSM+GE5efwp9Gv47Q3MYuF0vP0rriH
gJrf4fZ1wmiQvpScc4BLiflyJOz4o64DeaegaEsgdsDLWXJFAabK6MDAz1ZD
SLt97tB+fYccu7lodUl910Bp8BjYfPlK4q7cFjBWo5J1sFsrjdSfsyPUl7FS
P5ve/to0sO72zXntl+Wa0FtpWc4qOkiUugwE4sz/rQY/WLkgYydVmF9OfkaX
BV5uIbzzLVF7cRT8uBW5ZWZAquFm0PIbHndMIuudBcDJ+MjHK+OqiZjWfEbc
HsPJKDaGbj7a5f3NPDQLp82u59habGSL5ZImesaT94+j4f/6xY3+BIv2Jey4
JEKtmoTfXuRo2afgPnEIkdjmglmJsiVnpnlU1ETlsel52NP+JtYHtxC9W9kQ
e0mpnsoIVJmUYUbJLAb6CeqZU1zLok7mPVX1Gw6lCYLlXRM6bOOLLqZ45qcV
xja7Qer7LJey+6ybQFd6slu34G7VrM/PtZOJcrAjncBL1cpOFplwX6q+pzk+
jSbQrGTLP+iWSzexEJn9HqRbMdSUtj7BB+u15zBOVhxL1JHaZz1IfrLFj12Z
5YJM3VKQ3vPCQiz3pi6FL6FGBObvMGlBkLbonpOtGTzX7xglUGVUcvFkJIQm
fVDCJ7JJQ7+qdRxKZ/7BM9Zi96ZRp1/STYz7JARK/jtaCDtStpjF82LBEMw/
/4c+33yazFlspDVFjPUwehYLDPDR6L3Z3qja83/rO7kepx80dkrT9J+HMu42
DaLH+ogGl1o1AxoGxRQdGgJffIk/IAEM09pWljBrfM70OEZrhQGyFFXJK7xo
1dHGWM8199X4GX86P2+wkIyZVADZIfCTPLXU/4Jl6jHW7oC1lOBOr/Oqcqic
8ZmCdoxfTc26fZcmGB7+/puAXnLwSuQtlRHNTbw9WBPwWAet8Q+JIvaZHWq/
suM8+TCy5ZWrwhaFNLv+YulPIQQ+1QzykcAcXOv9j6uB+6xCK6qlswI8m4nr
+Ue2zEmeWdkIyo7/8kRyKmZx0OZdT8y/Nrrwa0nLRQKrVL3bUL+MIZ7jZjWg
BgX9GU0R79oYDzFbSxdRrcIOXsvj45urGvWkSFzXZMvJsmORwkgktCMKBbEo
4SxBH2HFQL3HldL1f5A6koSOqOlgSL4q5u4oUi0NsNeAaQxkX6fIMAwkT8qa
9NaOxfpHyn5rAxkeaiqWMkXVkNkbqgG18Oo9rQ59Cf8pouMOjwyHjpU+XjYF
G07kMe3jrdpcwPUlLsCqKJ+9Flsf0GVUZL1I6fTxvehANVGM+kqOJqsSYi7a
6aszCxofBXW8e5D5LdbISgtFzwfSzDsDZmkvOCw9oRxMZtd1ibHtsuzKHa9l
7XQ7QdCBquVW6vVcmtxfFFYCV5aSoWuZ9LoFc9eMfOk/zYXsjezWYPCmRENm
U/XMr7btMpel42LiYUfPF0GSFE3BGQg5Iw26SJV5XnTw4wujkDaQ13OJTwHg
1ROI/dYnOXzqRT8VYjbhoH3PUVkgz9LUy1pVa88+52KOKw+Z5nP2auLInWp2
jAKHMYvCeAFop1cgIgUHDH9ovEOY1IuuUyBUt7pljvuGLrYDGoeKMsozdUky
4jB8KLchxOS7VdDZz3vxjCMvo/OjWiEreWOVvTdgAMXrUKVYA3IeXZ4IiE4M
nbgDOdTV6WhsMeWjKIdvu04PEDaK7jxHQMZYAM11jd7XIh2RhrxgrdRc4UAQ
Qp+ZmWyZ3by0J6NFKJxg/xVR++50iUe4s7d72xt5Nw/p1xluBCyUfJ/94h6S
Q4HkViW72DR7xf+ownrEsdJqIqg1RMByiAFfZkfxlpv1QTHTpEIYd3gZUexl
WgXluntV6k+dkDFschbOVNGiX588lhKHvnlfxO3HL0C/0TjTxaOdGHidJ3uQ
emNbIk0O7UGBR6ByYqIs7RwZdSYrcOW6q064CS9FNt+PU/yMEA5Yh7S7HuCu
Usvy4iHmNCpnrTaZzwSdKFYcdK5FSsUSB7x1VbAFcauSppd++acX1ygc9Dz4
11BX9cE8cgODJrp+1qKTfIXEAL4TYO3MDklMbk7FbnbzMBs+Xh9HfF4VLvhL
vFnvWlSW2SzcykvDbvecTeeXX7rJfD+QDqupOGomgtiw1TEpO4ntCtsU14ze
r8fCJQz14XwqRxbh/YOi7vey0jaUIl/99typsBXBoOOHrVkF7b4ncVZNrKB8
P0evAyEt8JvokAcs8Q7Aj6Za+AA1Dz6fLfiTodMwmKtpAvcc9nTYKEFUWcn9
+u1apyPHDRx+pFeGQrMDJOSLbgZWlLfMnhwGCXP0Bj6jSU9Bs78zbGJGsOZT
BnWhWnJFZkO85PWq5OWpss5WQZBuiFKRF+uhlrlP9rj+jonhFGRfbWE6nb2m
BDT2yGoNdxYoKbOsAb8j4bwS3Vdv07wcN1F2rtmVvTZvpUeCHOJIgJeaPZw3
EpRPDEWio+vu715b1ivWmUpnNdjhMfEXmaItF2afzq/s88Hv1kMr5TYLQeVR
wYzxFZXD59sfcd+IjhCuiS+xcxVWt7U2D07A+NjVMV13LlX+WpwpSNumFm+C
+LVz2nTIz87kRFfcHhkkduz1+t/gzAvrDislbVQ0rByduD5JbJxrlXER+tQN
LKb4TW4KBJffQmYVdanrVXDPKoLpJ++UyXBY4NfvLDLwFm6mJSchXyhhaC9W
5u1IM2aqW1jmScgo3e1/PDLwSMlc0EnoWcu+WfQ/FQsapBjL1aCdPp9d3e8B
JiB0nIhmOGRXrrTF2cucH45VjZqV4Jc4QRjwKErV+4OAHc/rIpkCUEh57HwY
1EGtpIF9Ho3NbVCvd7z/i7PAiP6AzyeCbOVcMCt5IQOrlaXozMJhBQffdfk/
Wi1wBIIHlHSluAKLojJmI0l4ctokjd3congoLq6tDO212uGVNjvIuQC7+ZNo
yoWCsMyTEnmgQZMWWipg40+2Vnx2dIQN2pVpehpgJjOIJkpabg9LUr5tTSqA
PfO89CFypJQJXocKAcX8dJyoApfttnJcU9M6VilE/Mmqo5OQAfKY2IrtjXJl
EVrFaw2hCJeGAvox6rloBndgY0xKz9BLx9OYGPqqvrzspnF1u6VHbXJLIRJf
wJeWIwzLG1rZzIYzKFin25m8a81KIXlm0yr1pU96JmayTtukWdKjmb/ckMn/
SMmTukDHPV4BBuMey+YBkV93WtxUyybCCboOWAdxQD9InQU75Xew0wpcOSRK
srL0BN1TElfBJO8zXiVQ8tzC4ZC9eBEykVWN+mD1WznE4zSVIhYLGFTlJvlW
YxKVkaT23mVCRwle2mwDHpOJFnsoOvYvpZNHynk4w0ZUifcevBJLh/mU2If+
D+XnT95rKWIl40MCbldODTTImBnZapuc0ONCShbYhOcnkd1IyFsZUQvL19e/
rD48fr5zCnDz5ybN5Y1miDCXRL9ODYqujfhYBG+7KFxwuZnCYWhsT1BQsWNl
SWWdGXiy8zQZJbTh3J/+3G1KDDh0GkIPlYVq1xNk1NTk5fulvBnqDFhjgZZD
aaRfgQnHDhboS5jb7o2RXXbqTTPAiSA/cHJ9Zp+Rj/31PSl2wwPT+EpcFzfR
7/x0r3AWtwZvJo3WI/BMGYzV0K02dx/76tgX3e8seFeS9DPyrxsb+NLX8sJt
lkHqw0SO7SGzUSBAegTWU9tEsE2KfZKobZktgex+Va+CeHkPpoU9I6bMiSVg
fPV2wwI+9NnG/gTrenX/rClK54a1Q9QDLKLzMJSq6XB3bqrWGSTEYoRfQj8x
QF9cr3s1O7USPoSfYV8GhkcfN88SINFet9zFTc4LCRqxPglgDzJ4MpGFN5hb
Aq9IzjaOKPtfzrkRGVN9WJoXh0+gpbO8gQx0iDDvYzyGDBeQcBrkxLyD97+0
TPPhsm/97JFLbWfD6jzQNcFe2ofqGiuMvsk6X1lLx6QnvTfhJ7Flh3/pAIgv
81xnfN1nKZqx4LDDqH4+QJGuiJZsuZw68BQJ2EAujft3LL7p/s0XDIXGd4Jv
GpTFhWuzgAJo5PTo16qnhu0CwGHnHCZYKNiRbAQ2P431OdQTdRiYDr8eYEYu
4j4O5G7KkZmYI+BfbzcUrAhruwb1ItTycI+g2hMrRLFzMo9V582gDtwhYM6e
qdJ9Xaz9Je7O4jmfJGZTVEsw3YbMEQ5zn/IW/mkSDGrzpSHXcC3YFRt4IvHA
AZpgB4nohn6QByNa7sKMQMG4PkuDGRulqoIHoaJKsCuBEPI0CyAUrPmZ90gn
v60gDqqp092w3k12qllCNOEfHtKoeS7TCWzyULGmyzuO08Zhv65Hw2yzJ7sT
3eIzK1oeKYYC+SseS3W5w6fYHrRnZ52sqa/o4v5F7mZWgwvc/8HB6bhsVmPi
ymczi0E0Bf67G3v0FEifJHwTX953M/r/tEdjNw0E2y0drnKGr1o345IYJUoN
Yhaw7aOueqMaFDWUzijA4VW/6Ikmqn+qs8YPBjjU7E5gbnit+tqgIVtIeM3B
gcLp92QiodhXNx0amTp5Nt+CToFCYM85KdAtSF9nxObhpR51TpjdsoZSNEuw
/UBd7xK7O/suql7ZbWpXunp95QGOQLdCjor4Rr6yxwRN9Fk+wAnbDty59+JF
nMQx8mqotchaXP3O8Ojs2fkeI2rX/uG7Df/U2trtUzKXXQjJu+11Wy9s+okz
0a3gbHbC94KniFOhemJWo+fk1t5Gdlzdk95hnOsls98HEi74deGif8IlRtJE
+VXoz03WzJ+4SiD4zY4cE1VQ7czbE2nCP00xVntjFmljZZm3L8ggahKTCLMQ
XZ/yCxNubWgqLKsfjE8hpNcacf0miPoDzWS7B5UIMppshBZAxR3Hv8gjE3zn
TMmnpCXeieVMx/3g960w57HZLZE0HgJMgkombE/ioy5oTRz3YCQnPkc9DOjQ
AGPOgyTjpxfmpjO5uFAHT4NbNeY4BQ2Vf298HiWFaCrnysNoeugTh2oW0xgL
FblS0LGMo8zGJ6tvDTPa+EOF43EOZ3xU2h0H2MRhVQdmuyvutgosRFIeemQ4
HVJkEudXYpVKU1AD0gIJlxjVJ2x21SV+g8fcAa3RqvdFnzOyVSbcSVGaUnTk
bJeOo9Br/5XjlYe3m0GnsJVrFslzmghp+erxwrdgrQ4PvgFGopWwQzZtMmAI
NKHMXLWVrsVwS3l5R54xO4RC1FADvZyeqnkwaAg0jCn0M1htaC/oywBNGFqj
3YFXXTZG1i1XKdeFuzCIXoPKn4je2D2Ri1V7uCvc4vubs3UmRc4QRqzvAxk8
InOU//OdTOF2tOe9TSyLi4T/RQdg8kjke4+L8UwIxzLaAocrB6uva3g4Ggu4
iN/EIafmwIYKP4fkip4r2b9tHbfsL+olgqJAHfJlUmASIcZhKbYNZ3V5zwFC
b3qyJdRXAOqrLF+R8clmBm9Kv5dZu0yDFDuqCJTw2M2wovGBq6pivEHPrIbM
LPdAJ8I54wUg7UlJfgXpZ8JAweLKt0TDOxsP9jXmK5/+X9JuHVT8IrGdmzzB
ScH4V6ke0RJkSf02og5Jmrvcf2DFSLMEzEVwqJ7ADQt9a1J4+3WVeaapsMK1
kxbkOncEPlbrHKKv617Nnh6Uv3j+H1imrmlgmOmpbZ9W8Lb49en4qNquDl9x
QBKAyFaexhlQoMlJL1EdJFS5llDIrsB6J/zJ460s83SYVSVURNfkj7JhXQk4
q9c8beBo3BI4M6SKxmS4+aIFUJ5hiAOCDXl0dWaOQ549KpZHDuBs88Wy//D5
zggDqEHpN3W9avneO+3ys/kckIhLz+dGa8RCorm2j4xpKHtuX83u4Uc8zEkB
3FgrQQfH6cpJ+VaU7wzvbeCpz1/Ee7Yr9MDsluxN0EcOmNZNOwdmEgtmalZ1
7X7E2IIUMAhlfApScE1pmjSGzL6sj5jrUMSneyrTFmWbIzLj5aU2dPVkiTfw
QOb9QY4F4eHFPJz44u59rZ131avycM2uCOsxz46gbz4xVvkIKnc2XQgZYUfT
/mEGgCmDpaDoubOZkklrwh0tzYPHr4VBD7esGWj5iKxHPqQjWSkJVK5eM4mj
aqN6gzCQ5K7sUjw2vWWyxNlTyhSTOtg1fV+jIhqejdUZx6Wz1DlL3uMQLRSb
Z3VyXbvoMB5xgAoIn6nSSrkC68eNE5FvUUntrhoYvDKTZihTa0LMvLF47QHt
RaiT4w42N1onuSBb3RN+9Es6xnA1SYQsX5ZzR5BJ4goeUv+e/Xw0QoMFCErJ
BB9mDrfJNP6BUazHLGeThtFY1K4LyXfNYoorUXXDJJ0MDbCGwWveMneal4tx
ui4MKCLGQi/xkrEx00YcgcsOmmEGtbgz3lzurSl1sOkaGYtps2sNNORdVtjf
Ijp/7CN6djPguHo30BzNOwJw278iimcenmsBLoOcZkuZKKDLzxrlZL8Vw3A7
Mz009YpCTV0lPTwE7RJEa5malOdIOuMd3yB0JZPHkEvWx24xKMkwTcGYOHZy
A4TCIq1Hs5sVOlo5aCpnZQBpcVgX7vRTlspZyuW05kgLyYGxxadrRQDhjQCN
eiPfqBqEZksQqFdFWkZo6TtO/eFBq8sZfVGUu/X5lXGmgwj32rlRNfrNIW3j
HS7Kd1vgFA6/RFyRdJkmXDWPibyg3bN7g6Mtst/OuCN6LwhrYIFDfwMAsyK5
Mk+1aCBN4xGeQdtvLj4poNubrftDXnEOZ/pS3Ek+5zclWHd5SkPCtWbhNfhU
ZBXf+/GpRTOJv4FPtNqyE3sSWcu+nStV7Qgl5QbxnJsgndz6PCAsCNzU2Faz
z0iQKsGmbfzpZACCrCF3zC6GFxaZavApF5xaYtyEoyuwplfs7ei4HRSoMx2x
qJRw/tLXMqvwhpTKO4sqeMsiqFFIC1aZ+v72hq3OPtDTDb59vnCwHZeMKyLc
09+xKuPdfhXcqV91eDBiFzM47xCfh1w5b8Sq6Z+ov6FPtEI05sFkPV/yVsCG
PACJWHzTRG8mbBIPENr4ojq35ydvK7HmHBC6YeL07OQXw7+fQvRvxPey0CoR
R0TU9VGYia/CxZ64m6jkF21uQekyBBR19lQqorpmlSW/GPqRO9I8M3zuf1RG
oLog5DJWZ9VHxz97QuTTKP/OP9uCSopsgMxndS8+4EWe+A2i3OrHU0YWqPaw
/8uRVW3yA4yy9VZp1Tf5RgH6EqVoY+4l2L2xNS7pMaNkweC7m1R7DOniiqXn
1SUfLfJdMbczePPIo7NsnRfO1zuVeau+hpUsT80voUrlHaxuuAqR395tq+4B
awf6dDvb2Yzkb3ZPW0610JGK3TFamdVySu+836awU4GzdmcJ2FAxrHeJcB8r
vWAPIHyB07JzizLSoGA80PceeMCsZ0s5gLIEgWVBsH3DZozUmyeFxiqBEZVV
4jQ2ul26nfxHCa/YkYnN25IJ7rrRn2Yhs6e/dSi+Vyhj3OeAfkdAIckOLsrn
TP7Wr4kkqUxmbP8JyB+rWP5SeSidg95nvBz7oFutV0Wg1XF42iguLsyY7Dcp
jemVM01g8CBkJcNS03YSNoXGuY4IUjaWKUkUotKYtPJISJn3rLgmjVHFbLJp
DomRJHoejwA99HhW9DEtutPtaxewUHDVdEVSwZveEs01rZFdU3/ulQip9P/f
8tmob/0IoWt4iVpqNzUbze9pS6Q0keifQkC83T7i2tSEv2qlxcQBtdTRyB3N
0X2XjIbGDT8M7UNI3RqfEPyqjR2qzYwv6XmHXxNAAnMxloogDMkk3IVEbl7p
oex2UBIi/y4jnSsS44DVTYpWCm41DtpIc9pjNzHlsSow4fIXTvJHkD1IQ8ii
E3fQShWOhR1mWqdhmFB46SwQYs+n5gmow0MKDwmYJ+GRwRWnR02RLOtT5/kn
0prYEiwwLDhUm+UtiaOX3dvmQKQ559fMoQUEKlFoaAwaa4DYd3PdMEsgxxXY
wKllTxrrHrlqedjbOXEm4/SH2oKSv/z06bMC2nQ7qJADbDhLkrG0H/mdAAZK
QtQFuXiKwmTIgoaXZm4habHyXu4baHKYgIFUS75d/ozkXX1JBsTdGo6T6wJA
mTb8KhBwsup1SCtN4lQYeZx0Su+NWtZtwADyS8c5Zeb4DxaduVCXp8BS69+2
TB1I9WUi38gOjeL4KaROyEg9F/qhxiIR30EEGygckW41XIlnSun729jBuYKh
T/fFcP+hxaZ4KvGSepO4igQVD6zYZ+z+Ij1QXbF7hfgd1HVcFapQSdn8JLx6
M6JopB+zAbsnO+1uICclJfx37VaxyEbMcnGNOvbzFSJwKtsxvZzwBIDrOF41
RXC/Kt7Jyyzx+bgD3gTRT91XMbmIx3NjXg/Rot6qur07Wm8NJGw5YWceBpOO
DFi4HZhLZ/uBZRBj36zXKDUTqbVm8wrjDmRrRyMYbJfQgX6mhvtv97k15car
eS72yVoBBY/mHkGBMOgzftkjKvq3Eo9wgeTx0gnfqBzuGSefnX7SCma0jkP5
6p5sWRWs/jkdUlsPsTp+LjYmpASn8Hktq62wBKq4f1KWS62ZORF9NS6C8HiK
7KMzXIlQ4MhNtYIEXQMfqhZErhfl2zuS0gPf0Y9IquwXE8SckNPReoskugYF
YMX1hkKebVY7oNnzcbRbnClsKWoFFKvCtk+QnNuIYJTVLMT4NzEK4CwSoGXY
1JVSBrC2kutYBPuI9YpAEMTyEK0ZGH/kniWeBpcHZ6kzTciR6Y5umUBA7IMC
F1A5lE1Nn8gv9c7TTJQqLM1FtdZ1md1UGmvEH8Q34GdyGm8uSRE4bsO4gKY4
DWWNyleJhck1C/hf/RccOIqtoR/WHTLKUOGafnVOFPwxX6g/M0EHnJk8x9aS
oFays8paKilw2nKgewM7XrJF8NRVI/cp1lkIr1DVYONHF5Omdv4He3YPXbOj
p8xsUMgfMnYe8bNeSDcTlEFLGUDzdmR812UzfKn4U8OPPFrsgNnBTRYpvaiY
jgHAg9NKL2fOa+sRE0NNa23PiIYy7PNAOd8dAjWea3bgvR4YccwYYFcj4opK
Yzoglz8+mghs4T1oIf5fa1YssONtfrY9Rry3anNqN2DkoWV9WtE9s5d2W5/1
IAS43pXwdhuxjxwxylhgTvFhzEpGz1bKgfT8OYhRqEBTnHxd6JITakV9g715
irD9TCmLr98QH9pJZzb3/oZ80vdhTtFr4mN6MZofsj3nw3uINXh6bbmysbNI
jWzZpgb8Nuc9ftkd0LysidATLwiksO4549KF0kePecEgOzVG+b6A5vT4iSSJ
AimDE0TOSmYCfVnNJG/+xBr1qs8PDTrk/KzRTxQGoqIdWZTAD/tGUm/NroVC
6QT1LMW9g2Nzj8a3a54BwR5ItU0OXGtgEgaJ2yluMYCjJkbmTlK9ISShU/Fj
sSADwFN0hAhZYHmaqYJLyBnE6CuHBKULli/Y0IcSpH0sXzsixArA/g9FD5Kv
g8Gwd6ZtuybgWkp7fQqPVkc7PhQoKEJ8vq+d2bomrG+a/4qLBiwTnG3gQoa0
XrQyrK62v8SEUztXp8z7zeUpRFm16hz3CWZn+dLwu5cmtM9aj4+zx8nH4Gqi
GpchNB8zEvd0RMt4BLDq/Pk2B/uOGQ49zdxcsvZdBazTaSdjri1RZD5bYtJs
ef2e8aa/IrqGapYGQuZXa9iMzdhvy+DoBWXEpcFnQKBfc26QWN3AEYCECfje
b0nAK2asuQkLtb3kaAJn8wDn3eMrdfEIQwtgmmbfIsxoPzQOEcg7Td2c3VJi
QLZnt6H8ytvJyL91PbH0EOIvJQoT3oEmcXP64AtOMYlOaNI8/YuRpi9JTxGg
PqlxA2utN6cE/Ms03IHG7zblMiH9fwmTXOqIveQqSJi52QtzyvtI92kAMhex
i1nsnqJXD0CugEfOhEchd7lw51oNeJt4+VgU+2l8tSF9Y9iidU0YhJtFtwgm
SWyU261KLQm2RlvR/VJriIVnHBWWQERL0VhiYgJriywuUeVVPqWAn0Sz4Yyh
r75Y9XefLZJxA+l2ktlqBsP08edU4sXV7FG2erL+9DNyLCHmKSBSuI1zgDfu
ijjR4JzJk7kiP8i+63rWtPuWoLBlBOk/IWWP2K42lPqSQLLOVtog7FPuQAfs
xIzIcdPVMRbyHWCUzFCEo1PCXvjleX2zx3ddYql+zFL/t5BzqwbA95Q58W4X
16GAjglLTBWEM44OKv3Rc4+rZgBaJVF7ffo+9h6YLvEfueyyaVfxpuZBTQCb
py5POrs+HAa6KEze5nB/SCp1uWrYfu6OFgvm4z0wSuLhLr1Vt/XZxeg7KLhM
xlc/XA/0YNvpYMgYn/EbKWSpTs3HxoUxnb3fXf2W85XwJyg9BYXMwyBWNAhz
NAorkI8y7q7+kumXx3ksgdnxKber0cKYKZsjrsQ0XF2n0LfE9/vAtKohTBzo
8kJybm/WIUguzQQRQwwj4l02tivjFQA9e3gvHW5LEutd0T26xfuk6yJXHH/p
XqNI+TKyVVdO2TipOOHSUx3TI4auEWRA9vSCmq6FY+ngkpPT14K/gYg8MOPU
FoyUTw/ggdluYWDU+KOliVJYCnzm980tPtmufN+y71RydIq39Vf3eJ2ca5hx
jl8PpZDDCKHI+4LAvbxW7eGPB7chJatcVeXB1/BgBhO+5Prp0UtAlxuyV/5m
6nJwXlBB3u5RiVj/yJXkLTc0jxTbPPqZQkhh65MCe5yHtMvVy7KFkykGaMG5
H/0bjhpHmk8Yn9HJ3wPUEEpaDW6omWEKfvCZ9EHi3ivOjwy62zpiGOLsyrOW
SNiinV9+9PK1BUqZyXMeePKLZQvYQGqrSflW+j5p6M3S6/XuQzGpl6pQpqaV
VPOShOXEr2PzP2dDLZBZ4z+xHMZjupIliUa3vHXevACH520VbhUmun7WYqP3
HQUYm092ZzJL8SfEq1vx1h+9a2rTQmEQ7aJUeH3nQ4fM4XMQsN+8ymkWUf1i
zHMrlYq8t0g7AgT2Z1NWu9YaSQaXQxSKa11vMaG+7M/fZ0wWouA5jh73nkfX
wyHz5SsAWKefzNFA+G+4Kb42hg6zO+cWoZab8/2n9b+ymERoPVVO1e6c7yNh
p9gpoBbJ+oPtMF9JBW75TVnRx9hefu6MuNc2ZLcofVeF8DB2AivEY0XBuxcc
wGmT23kzRxi7eJUVrge64HnbGw+RcaXwk70RKUl5rdtyaF8UUxQXJ9IP4Uu3
LbHKh1f8ikuL60oEbYJgWsKEqSxvhwoUgRwgpcxwptD5qbVv5jLiMGiOU0Fg
DmCLGnzJRDe4G0mQrodwoqhcQiwUxvfLe6z6BoOnFNgKOwmJ097m4TFDVMIw
jrDXF08Il2f/6kJaUZg6+3ttwrdaI+9nE9B59+rgpA+IliaaC3W3H9mpk/52
uuiUFbwSvFCPQ+NNlwkohS7374D22a5TcufzS2elfq1W9Z9LntmnKxCk3SZH
i9z13iy2/UK/Ys4K9pu5/qnV6+wK667z9GcBKsmtKKHdht3uder9g64cOTbH
UNlgFqcgsPVdiqD09taH/Lvl0uBqZuD/h0LoPOsNkr+Lat2CrK0SbJdQkTME
PvleFOiF0o6Hk7kvMdpQps86DNRBzn61VGsbySqDxByy8tEYBbVVu+4iBIfg
nVpDWMo0AbU+bWmBrR3VWojBN1Kwt96b0zmvww2j/j9ZH7J/aWT/tFA9r5JR
y7Rohtx8gFqNtFvfztMXWNlN/gqJiOFj5Q8U3dlaiEHLPGwcJfuExbxtO2OO
OweT9L2JTlbxQ8inbI6/Pk8QHBQSWnxzOcEh2dmV3Ol67K8EMAluqSMsSN/8
5T3UJnfG8UuD8FgO8VV+IkQDsF8O7IFlTAC2rj08FSLW/TZo0YJH9zZu7lS+
MXHu9DHZQi1Nh/wdR7/Yp5WiIQgBe+MjQo4GC3fZvyVEYrYInxaSXltelDY8
ANaFQ+TepCSDUWM57WkjWHYsw+JHRBARSetjL9frpOrf4R3y4ikuSsao+coQ
pax2VdLxRGmcoCFGcV4/1YJ0sTORaPvpcJqDLME1NLOLl66vZg/EvetiLMXf
otKWeplu18PAtyS7MDdH3YDmGvm02gY6c0u1Kp6RjeSdCUEuAinsa/sIAO+4
iA4TWej90vqAe3N+mJuh6jr23ErPvl+RLn/v+S+6uedv4gnPxUyBjJLK/S3U
8LMSUjutl0w7iyERZJ5WkuItaWT1KIBU6XkUghvRAwJ9pDSQrT0ViH6ODlAQ
DXHSYqNn0DDFRuk8nEhGo6AP9nJWGaXNpFdLcBS7rzdlnkXWJ+G6kvR0eGR0
d0xwZNO0x4ZjDJlLuzDkShznv4a++rcBQwXGSb7E1StsTg0Dy4dOrsFt4gic
GeL5ukQ9Nqyp+hfDJbWaFLHIy3BSvasHD8CS8px2yglYVtI2KhuoVYqql4mc
+1WiWh9OStnHfoIbhy8JOzU4IvphqfFOpMlB7C9cGye8I9A37mNp17Kn+obB
neWSrk16dt1RkZj+jFG1zPdil5JVd89pLFl3AaLWj6t56V4Ex3TppXx3J1kT
Jc/8FXCr3pMn9VMcq0yplMxJS3fTpXs6N1eGMVJPqOQqimPOrbMT5vFEHAUq
rpxQmqgFYK6GHKmBMkOI+vFGTKPgCV+ymaCm7G5qZewh6djwZ+wjV5iSTm98
VpbcRciKN2SdynoNMc0xtUbvDs060KVBZV01Ez3SgbQSypk1NigcaUleKcUX
+lIR25YHtFZ6W0Wp5O8qCD7GhbiDnKym0fJlv8byglazw2D54SW0WuuAFWsg
VUn59Gj7e3NUvcOZfNcZ9CjlaRMftheN6P+VZDf1xziHNwvTrO7xCzopSa3u
Z+WiysDuWBloOyk9Xs7idthC4/JTuL7tzi693WALeMBKNR7KoioY4kzCr5Qw
cfT8n7aGfvKgRP41H0NizBarvQ21sYLZLBebv625JMjSWDz9TUmfx9qoH6Dj
raKsXpl9fbElG0aw6EQzouTzKBE99cfehfJPPB0mgDts8e86pj6iReav6neG
CEOyU5tdnWNrf+q8mrkf+7TMpMfT/03iu5SpnQyj3C6sTeZq1Z4dBvZe+SPZ
ZfIlHKSypiACay/rE1pjKN5Bi/4LJVKM59vZuITihG/K/zrP4513DllypBFZ
xGSHwXWCsUqb/B6o/UV69S5O5wJtp/jex8OzmV7GQd2kABlzJ8pWHlEKYYap
l4e2rU4o5FRcLPtBzqkt6fvruqXIBDti78R2e50EpoeGPzKylN0mwvdvzee7
ifNzOFTn4k2U/NyxeiFk3BZ6PuHXIzyVTdbZlduV5iNF7/ZrZKjohSkR5msC
gtJxn6+enYOZKq3HQ5eYRJfrOpK2NYJQj+sf8eG1mIJSrI1Of7+YQiGb4tt1
Fo/hNvam7tnu5dYE1gH8CeN8Sn3T6AIGia3YfWdaOidNj3r6u/bXQr3loZEl
i7yPGv+NWxHcIJr89ckDDvrhu/ElMOKvofSb7DEwYpItvOBQ+Me2JpNF1nWq
pZeUiSjLaXHf7dj4PCpC+itFkApGIrNplw65hl83Pcni71l2lCTuuMXHGD5M
j63cFuIgCcJXWJp9QSyddIYqaM5mSaW4v8myFaKvkLZ9uxjsv0BVWgVwZdYJ
4Qhmk03InCOm7hDKY1W1TbM9RO2OuE3/9h+maUfdbM3FCTEEFMhoY4FP6x9z
V4nimgCTobZUgl7mYWsCmqbfiA7uHgtQdOcb7vF+ayWatkJB9QNHbKhCIy+R
TbcezTZiqmnh2f2jK6Vb8DRLNl0HxFgy5Kdr/5oxF0xmaAGxeGpQhewLz8hJ
NW7G5hEK01HYKQ01Esktf/AMRVzAfuK9WFBVyRYHjEb27soJwLHQ386HMfpU
xloKoviysxL9Uch/G1ldhzASpRn335yryk0PudvFeWPtALldK0hWdI6KzQic
f142iC9pXnsL3kGsaA8rHWPvHfiQu+Aicy1Ti0L8XwABmcHrNR9MzY6ZPARh
TfcQeNQDVXGjMtnkiRA/z/obBQyAQahAIBiCaKRAO5FZ7E11V2q0eC5A2UJK
kt/AWfirj+1ocSLRKaCjWInQGf8oWWEbYwDla4nOG8o4eQhFRNt3oRLMAvCF
rvwOhCoCpU7+YFoIrsbRhzJNcAEhb7mRjtvTZwivkmfXJ9NJqPNF5CuH0uSF
vGbeOzUK43OyTTEZ2eLX6PoHUSK337kOiy4XpNS7sImLBdYF/ZL9t9bB3dWO
mDCEkWkjyt7w9i8m/wXDkS9luyk0XGG41KxaC+Qc8yjd9AAel6C4Jic0bU+j
3U8C0i7Z0n4ytA1qwMpEicuSQXKYm8PDvIlVijL/jPmLwENXZ4bYduduYwq2
ryC+oOBcORzahQvF4d7fE/y4d2ZO1jQZyqC7NnCH8uD6bBqw+1SFJFYaLePP
V4Rjzm1WIhsEcvGkMby5ou5dEdrTJ216J0PQaeA6ITz8SlaCHDrreHA8arrg
K26eH41IP/bE337C0CLzXhcnWBhteWaRn6xpfgf9Xsq5e+TBVKsRXELJIFGY
phYWQZH38CZXOg3L5xKFOkiVQtSlctHRORcn0bmwBwjUtjL5GAVI5BUhfF0k
9m/TFfIfHCKcTiRbwYjXnCVLengkEZEdLKz2I2bxnKec8ne3saEpK7QIa2ES
xf3ctZcjdpV2cJEgB9GIq1Ek/qwGBqwiRlLXpCVQJ/KPfaJB394TE6cCxaB7
zKrtJADKhGv5+jJb0oR3+kTfMmaFfsM1cDDGk4719tXrIl5PtHQ6hUfpB4bH
wmNFrNIA5R+mDOv8+nYoiuq9vR5xGzDCHH286jSV77OV3mZ1wwDBTlr2sgBX
zZ+P34tniZYktJ4dalarmfmyAfluSKyYqd6HJ+7Bk6TXmZ34Adjam44ciqHC
vR/jPWj0HWFJdknC7H8ks+8tk97WwkZI3jVyy4FvPcsdlUkQ/6pbmhKQkQNr
6AVyJdNGfNkrvDyJ0jNhDZo0LNs3o05xMn+v/rEX4c2JW5NjaySrSMLsf9Cg
yoHNhytmEGVKe6R3Hl+34vgWIBaA3OQ1E/TlFTnBFJz1qEceuWsdFzVSN1Kr
6IFAWt3LzzI8X1HdMQ9s6Ux0gqbYcoe8R44iA1oY6KYSIWy5MR45CrfYVcEh
ZSyAQZy34EwmS70ZT/4Ot/NvYcL9qTIUyQx5NTcxvstVdAnSvW2bxVVcZGvJ
On0mROQscyQhRJJEB1F4HW+TzpHo/t3GNySVo51h36cfI3o2irQeeOdfV0an
3yke6wHBy6AojrlpAF8iFOQxLkwSfo1/OZCoz92QlbwPjttrg7V9tq2HV9rE
Y4YgVsje6WnNrbf/h+i/egj9yjIJ5xWyGmuxP8A5BY3GaarXgfuIGMhNHe/J
iuzBh9oe2fYcYdfe35O34aAGMCb9oVufriO6vUB9rcBZeFyiJCF3M+RUW29I
HJQVF/yaX6Kp3zeieNWoMf+9R9yhca0osqYYNmgHjJxG60JbTTqGT6GqryO1
nGWmtqqm3Ptc90QM7mkuGaI/yOhijLM2AsdVd8J1PQv9d2uOJCnx1/A7fiGK
TruECwPU/cfXen2pEJNyuNDCtTNZPT68hXG9C0AngTgba3guZ57iEwKqjoPH
+xB2SXsszFUMmtJMCz7WLHf6G2YFeAZvE+AKuiqSj3nEpo5AskTvZXbUIHwk
w2EkqrPZFEK/5HudO0LiMtFAx7dD+vDTsaQ4dvZWJuWqTbSKLeB4IQEUHqXD
0Ijp5a3PYkXvy03Bh9AR7905UHGDc7Ybo/sCKYEYyNi+8r2lZdTV/4EV5ceQ
5VAvqurQPtRz7xQd/P/tS0ugPGBXrOqMVjMXFIS4FbBmIiwqju+OEgigP/+X
/E3w/Mi7s386p1or1PpWW43HMu35aNFjL+O/ZZ7ggP7X7qO0T5TmGh4NDHaw
j1Vv2OArP8ZIQZfm+n12+ToW34E4CMvtVAn/HwAzsxXFgv/4JSofxrzHult8
90MMqvZY43Zs6czPQOgMaEjglOHJbMTKiHU9i8hDXWpGbqUMxMGOfcISieK9
P+vSDSKDIOTMUuTQ/QM3lzCSFV2/K2siBqgyRI9zY2V6CdqCXIGYMMTGJTqQ
6W/64pPz+ldJzBJS64MAhEgxRsLrB+p4YHrfMOadSmmqSy+OQ0FEvB4oq/gS
QIoXRnQeAuDNhYDnFtsgb5PoAFVHIXHuVgewiS5yvU5Jq5gMh9mdbpUWxdKo
9ZqbycRMkeo1sW7x1AUAHhEPF9n4FTtJ8WcatMV0HxTs6VbriQZuKXaND3n3
QfQqOkc9kFFPmDP+eOaFU1XExxIHet5aeBDDAWo/9oRMghcDz+3ALd2VfWPG
7WtfwGV3i5pGm4zLjm0pDLIGcLfQ+uyxScChHKVTf8mDb/JJK1peozpAZkao
jkIimeFaiMLgR6f4qPmBK7ErqhbGUXJzrU7pYd+0nT5yRrj0rRZNBm5TXqcq
xDuybGXPoxMllaYvOMXv4PQFRc6Qx4axrCIZBXPltHgplOHi3YUgDZ2WuCeT
aJlXRLVEdo+4dIpBWuZVbYUITyVyaz8mEj0oAjSH/IvM09Pjup6OtUQ1d7HQ
G6nOkaJdx/iso2YisSb33z8pGZ/p9t9nuoFOgWutuyP3UUGCu94ePbo1rcNn
69ZPjBKNS1FegtqYJlgekPr4m0LDGpbE4CuACxnLDDVGshAZLDHSKWuEQpQz
YwMIVEg3jTt9VYhmb4M8diVS8cjTcubLt6sqR1Z1s79Cr6XLMJnsHy22Pc75
ivZKGPiYlVcqR0/immst4jc82HMIKZesPwiji+zn1PFNUrtd3sofHkfMt5HY
qfgG0lLAQXkmzf0uuBMIKg/2Qx3NhG11GQmpo910eA2mwJuUfjVcWBKNMhqg
NAUvJHU0G1M8Bwr7uVgqgiDfp0jhbrXpf+ct96o4s2wvMN5i4mF9nrUE9Wze
ZC0480gwwpcVFZ/vIxracACjTjPiG23IwjNzDimrzIL70gG9wkkwd5hNiIYz
z/KKg0rxfXdZZkhDzsybEV7rllQXtnsB5qndIJ5lzB/8+sbUHA4ooVfqjlGW
8C0h8Dbsya/MUbBsoWKbw2lCU0/HkxJX0aRYAAM36JxVxEAnBJ++sSma2aUl
6kHH9MqfWSjw3NPREkNHYAB3s6YHA/Lfie8NapiUuwEdbPB3ECih5tyDkbXV
c9/clsHJZNdB0oIiHqDBHmt/iGgUPiiSsuRqZGoWXDuj9BNmtwDxgQL///1Y
iwbpTsry4z+QCVSwHXpuEbTQnasMrBl1WsQ79AQwfUVZJmoeU5nHUalV50Ho
Md2el5d5vilwZgxhuqFIcfUTgEncZ01mZoFnr9d7rCGvb45yYNzLMjfhSG26
zrA0XUpYYQJ2G1BAs5oe1EPfrVjXiE8NLfQEDqMe3/ztwdqMqCEIbfRuyJND
sQHTH42+1SalWnxxUOD/Y2az/Stf4XDAf44kq8GUzUBVMBm7LRu5zJjlDdy9
dk+c6nsOKsSX2udgmuhV2a0E2MnlIfiOQHjRtmci7o+O7YmRWUxv5Edqzlng
m/81KzybPKPJtsR4m/08U2qzDZ9G+n0fDSLAXL4ktGPFZnfbUJbNVLw82iPG
/RV2Y3g5iudnI99cqdKtYM5Mkw5el2B3y0ziHRiCSi12bpL4V2yrQ86GwNUo
mPmtTTbRzKR6LpyNJCqw63iAUtqlKGv2mNFOuxmt5OIyUrL/pz+6AoS+PPfE
q2M012XppbvDAUeaXOqqzOB1r9SO+XUawwV/NmIqrWc3SGYSzSoIb2gcDtm3
O1xcyV8U4/hNcNZ2jXpJAXmw7mqYyVtJ0l+6sbWxRk/trLWG+62W80cYhQOk
6NCGetLPIIfcjoSuVUhd/FTA7VG51UhxY3NpOOiqFPIF3psPkQ9HU6hry9Cz
IESWCbAFj1EQvKYWuybtfkziK99Q0eUihu8YMKf7ewMxWCsZHkh6OV5MXJVz
fDeUN7+N4P537O3MgV+VtGCD0UA1XHeXxWYLylNRDtmJd0dnvyiJ3ikSM1Gj
DX5ZioocpAiqA+NckqV6+CANof1pDpqG8gAVe6AIENJaPI3xl2kZAeRCq1ui
msTazTooq5surjBqllPMRXxeiPb/ohgwPeard4bA0uvSf8Rz9xBPh+WAfRMZ
Ovpvr2Z2Wv4DrCB3ZeLqJ8/5tMLJG+vaeojDWaraouh3E998KczCrhKjbSV9
mZo568I8fjfdq957wO5cWHf7nZDMEcefEV46R1AqD8CCxdfDM38Kf2rXWVQY
nSf3GsfiQHrh7nnHN4LEiPt74LHGmBdIY+neNpGPRBzsq2a5GpCebEH3vpG4
2ZRuejZd61nNYFzffB67sPq0heJSUmx09uhgEE5rsrTDF6QMOOQKM2sAN3Gi
RNGxoWIsu9ZBKGX1OpLxGAs/hnOUMJ89WHd0cY9TZOYmIPZnN2olB78IRmGC
bt0sk/+qpq2aV0poJCOcSLpbcxCXph4nJXQViA72TsXlnBezC4lTbzjwrFwm
bn41EZu3DfNPsro+MIsqpHt7OkRGLKTpcJXU6sFdTkTOTQrJodIJ8xXIc3Fm
bwDnmY5Pcj737AYPozYJc57eKa2e0lK0MD+LME1+hc0wJEHUaA8sPYY5oGWC
bmUXcEvx7mCdoT7Aln4seGsswolnCmQqk8qbtpBDIWDm3EKSCMPwp2YjmdvX
akA4i3lpfdspcvkBH+F+Tw0vt3Q7bh1+Sd0L04jKspsSG+C1FQ/W/4EVxinM
NisZmR16dJG19elwqpsB8AxMFZ7JCrV8lC1Xt4OPbiS+R532llHGo0HpL2xl
44ydRGMR0Nau02iOcAj4Qt99RRb3RcPQ5gWVuiwIncA0VZeipzVxu2tg2un/
SdjlT6/8axDctTaJjyqH6F3VaVHNTY0D0AOZA9T7SyqRyC5lytw+nPMcb2PA
fISTEdRIO4gi0oYXBG6APLg5Wk5HXcFfPVT4XX3SGXG0sccOfI4rhKtcxE6I
B5TeUKZlNRFu4oblqmfDXRVbbWU5IoNuqfjyIAHlF4jR26x/p1tsaDOmy3fo
H1LFHH5Mvly7g9npizqeqeDrJNeXrq57tm+nU8WBbdRYAiwgAz68iN1tOpgm
vGPQjZO6FnqLtfcnfZJOjJreGhm8DwmXpRbW/EKELA5t4vlVm6uV3XNQOgJk
oZ44vyTXmRVCZnw47YjNJuP5cAaJ5x5BewbrVyEtRMbYapOjhNPxhJLdgtVT
1jeW/9ZAb5m8Gbbkz24kzR26orYdMjra3gsOZ0XZWUWN8UEHqwM+iS9Ct0hA
mX+pO+QYqfqNM4MZ9QarMYk4Ogj9+Ny1sx+FwlJtoO6470JdGRoP9JP9zqjI
rhdXkRQhi/2cFeHlIZ5G64NzwMyzdi9UTt5ZWViEXf5b5MuQgEOZPqRI7t85
kKiDO19Rp7Wu/UHcPXovM//YFgT55ly2qEzpeBvpGLY5z1MZocK0iLT+W+sw
6F310SVVnK1qDWaxx5EzHkxfAil8HPmW/fFeOdmA73qeKZqAShNsnyyIETWh
UtpfIEG/aEvEIAAPTyGCbShW/atR+fetLR0rpifQn2neFB6qULszXrXoChq+
b9z6/rhnWogb56VB+FpDhgolpWxsKZcIQhGpCX4hBzlkI+2YbFFFLbA1igiz
YAN7W5/0vDfr831cIo8UHt3JgtYVzA5+R6qZmVwonm6/5WbKsfFtdvmlC3We
oiPNZUJowelBYNNfJYdaI+hXYq0D9zQF0slmnKgqp0HGQ2X4/QI1QdqzX9a4
x1Lw4qTudkOaOyGImxR11Hg2rmKIZleGGvVdLiPNfNthVY50y0SI/iLUa9d4
Kb98AXrREh1A4sW2aJ3Yftv0lDZRZ2JtFP/+vDKnUY347X0qncLCJzmMez2g
uk5e4nR4lke4g8k1772dw9Dh2f273kvsKIEdjVutQh3YQLft5UFohaEAuOR8
qNAe9HmajTi9pEg1AfbGiOkbj9G2x64fglPi79CogiuomIR6kzcGEv4Eb5oK
Vct7zHoWylkvB/b9Pm6Vl4OQQR4BLkB3BUZ3HzeDPZBQZO1U5SRcskKdajk3
IAyx6ZCkiZM8uU2yG8b8YZru/Sk6f4VMTQxQwRzCa0lxVwggGqtv8lD6idRd
rHkRZW/G6E3c6dILQEgZyYCTsbw8LaB8pZhQw3zE/MQH5HmNSgttS7FOee3K
bQy5hJ0YYfzF5PGFHi5c4xVilgRrv6BvP3aYmuf0tC5Tyl7a0EDGV2GApoNl
xC+j8B+BiSj9bqdP3Ak22L/T0V7FmPibzoBw/zNhxZpxkjtz5hLHrpbqrfdw
TTQTm7A+fAlw35xyNraDuey77Pw+8rNingebU9cogybe1Fe+o57XUMdoqC0G
x2sS1oXStdmbjhQmOfwAd0+U6aRf2HsjGNicq34X/Flwjc5W3VyNJdvkiC7K
gZNcGniWpdPUIOjSDpmkvaMV1wk4cPpgfGHxsX5uIwO0UZ7NAqNkyBRB/k+b
4gGRjXCsluyqKYFi4DVHPVHNFx/Kn8UGX7RLrJuQcWY8Z5SqkUVvuKTWIuXF
5YKQgAIFrGoMYu44J0idoUJmvWbgI519fPU3K19zkqQtQ4KdrHYUMxluG37P
ZVQ1uujpnlkhyMKnqEQJyiFzYFlEROImWwKXL4YXaenxcXdgKYnuKKDsKOEo
8oz15PWemDCRUeZH9Wk8hAnfW771l4cz9kXOGC1BAppWAwE0L/dXp6fb9bqs
tllXycFaJvk+ntOyef1XlHcJWIPFKWhBnErdDAVv4az+uZPZjP6SYaz3ny97
8hSThHh6TjR8Q+larzcyrOol1KfPsRaz9gulR3XbPTiNb0CgznU71PQE3jy3
7Lg5o1g0313sVjjKB2U8y71SXZxGiFYHxbEkaad0G7ETwn7z3OUFi5ccBbue
akdniZ+x1JeC1UzT2tI+6cp31lE3PAcgAc+XrLUdBtL6RkVnuPlD/O9rJ0YW
RKSJtyKM2xBSfJiZDQWHbrBk9CmFuqDeLi/N3jzEAn9V4eqaxX5FPtHZxXYJ
JKZ/xD8AKVdMEIuF1Ztvc33gR7exu2REiawwbz8qzj5s9F3GRp/zzNc3v3B2
+mEafDbshjEVQboId6Km8bqxXV2ZDNFIZMH9fA9k6TfdFA3xi+wy8vwCgTMv
ZJ4krYgqF+QiSE8kX4ApM+3Rv+7e11NM+YxuCHm2oC7EAzJIB115sFWxZu5V
OrjyJAoozkWQHql3hcxlNqW1A59NtcsLI0VQgt9efJeadxCmRfOwcjZfdeR2
zxxK5JOoZhsNMD7TI1NlLXWbtXIX4YQ9HMnEC6CN2SSc97ucMyJo/H1EA1uu
MmOdQyyHcsEsmSKlFzrfliMrsx0fzOvIsQNveJQMWgxnKUZZ80kYf66is5Rq
Hz7Y6kaedk0wolY4p1WpwMLMMyJjfe7IY6o+kasFSw9zX8SQtDNXZ10NZXGU
VpbOTIbN/3gO0vyTRBhJU7seC4nssuMCVvzp6m98yx1i6Cy1GQSgtgQdrdzb
L+V5qxZG4PFAQUWB9vsgGLWtdblSOI/eelYoxegpECVdRHuJLi6LBBHtXaCT
Ogs0MysIsT7NBiWZy9oxrrmdY+Oicmbd2/GRu5bVmQuUE4E2ee/ETKx39iiK
r4Y5nBUc4iwOG+mMzXD1FdSuWcfQYoZueXwzAWLwxZYKuhVjm6n8gvCkhfSa
QsEAF9nTxzEK36p23INYarn70cQ/mCUmU/fzvRnbzZy3t861DjG90ZbIyFC1
jL1gxyRgn/zGyJintQet8GBDqbu5jU4i4ASsMyf36UDixILqb9drbev92Tlg
os4m0y0C0w/OfN9WifuXFCbWmmHzsi/9HwiauMxc3wvXOviviCNRT01Utolr
1TEHCfcvbNAhGMdHVaUwPHhBmA17P27Nj8jcqi0K4XtsAjYyRS4dmZ02D5Eb
A7uoBFAcVHetnHMhtgoB4oOPaYAZLtUvEuhDl1BGy5c9WZx14he5nMxBnCv0
ro0gYx53rdtE8JCT+ktfHvesa00Twe1/tL+zoafN/SSvffmMFERFEflBCS/9
NXDO+FzgmIKnhwgjju/l0lTXslyALXJjyRgz2Yloc+vgVCpr6LFL41+GytRp
nWt7oVLGkzoMGHrGHF3gTmBchOoBP8Bj5DnQsTJmP5eovk3ZGYXW9rnxM7NK
fqmkpcLuOELvlddkg/tAlQmg8ZgACGDe1/mT37ImqLFzrJzUn9kzmzjbaSBT
joS3Zx/PipvWnZlFulT81EUrbWo8mhcVHyow/gPz1Af4J1cAglcJt1v1MAiR
TVamJ9EsugPqj/oyN5UVzepPrt4O4nhx5vwSHud/joJneYMnt3hAIMV08+Ux
DnlUOYyM7O05nkNRmCiDF6kUh3NgMJ0Hkgs6Opn7ZSkFnb8jUlN600Lv8xbm
Jhj1pIjWf65Rq79COWYS9QdA+nIfzBauniTx1pw/OcL+qeNtFeFHSbVVdjX0
saiW27fTMvgMq5oaLBsLw4dd5hqmHNiMoeim4MfHYZlp7+EcliW0v1W45t08
Ti8FSe/MM7iKhOC+w1wCTCVK/qfBmOSiCVrSBLxPfNTZ+aeuM9fGqRr5dlD1
HrnoRPS440fGAVDz92n+Cw/zEC8OIhtRZ73i4qjOZY0fe/aikSCudo7jtKIU
Bf+Ctc+4s/Pg5FgZKnZDjfnmi29ujiucBv/Lfq16DyZ6yFLipJ4m9XSgZ3Vk
xN5m7lfXcLS312b+85BmUT5TIbgtL9iRUdBI+m2J7XBtIs77GNkjPEWiSa+0
O3ge31CXt0Q1kLZUIuw72BOutbVTJ9NvmuAAKoMh+b0ozpSWFNubl/EmTr/e
J71FC388s9TmhsBIBzLWqm9YZEhvEJrRo4gxYgsCAqWrFgQPKZpNY1CYErBS
kqvcZFKiMzuyMx8byQnqzS2yjo0kL3GPfIsEXYsIknEfhuwcJ3uHuyjcpTIh
KnqtGtvySBreyE+QjQhquQ5sG2Pbxqz4JkPelWbYOJsdlHkx9QN2CkwysYeY
DRINhDAL7HEnFwbqOPDeqksygj7ImuO2qWfRddRqD++C4WTPCUXa+eMjbhW7
ZJVmkRn+6n3I3m5aHCLOol2ru9OLSmKeEEsDkhhArLIJBlox2+HJJFbO/MOq
tPPfQLUT7U3DdaN2yFtKTj/U3ggSKVZ6qHru+x4MvFvblagv/CRAOht72aWp
aaRu7Ly3cAGPZ92+c53x94QFyoDHWmCCw69hpH8kVA+p3Jf0kyU8m3q4npiC
7MGB0606s6vtVNltXYxb4omSlDxw15S+7j8xG9VwhH2SAdy0vJ41apdOBGqT
QJzkhvp0TGQCU/Ks15Zotc5DqMlgfLFmxA5fjLeROqi2mC7+CGVsENY/HCJ+
cbH5iiMICoWnq50le2Fqs9KYipwZvSFj8HNnt17Ett/qko3c6HLCueoIx4Yj
ClCYbDaBQfym/cuIl/hxKjRBAiAiaqLMU6bmwy5PSKTKOyO/nbNyoCHHTKF6
1tjTJB80xOC4YI8711RDpYtnBU/pHJEizv6QFDPkzqZBmGRDyjsodE7UG9mU
B/+ctFomrvrUZl9OQPoRC01t9cvJgV8i8UKJT9ToNIu01MgSEm3D6mJm8+oj
57oPmzpI/OIC1f9QzFzPmytP1N6aIi6QmylnNKdThY3rOyYLLIMpbfgOhJ6Y
3VBqOgIPt+PkXFZFp7whA/60K8Rclp4BqjrDcWGFd9MzdMum8ncZ9a8oU+H3
Ef9H8ScpbMd6GH0ngieVueuwHYmDu+qkdr4RNrDk1x5KAEGDQaOQXNJhUqU4
bfIhl9SkMSIbp0RV6d8fNVOUlsSvScFak4mLao6tCggBU1+DWpyCv4tRa8xz
1A86APfqhSDAUbpOaJ5bgS0v+KVKXiZhDzxqeHzIDC7G2jRfKZ9XKMc6aZK2
90H8Y5iEJWKkVnbzzI/aGzqm4YRtYKLgMZvJ29ROnjgbebdiyY8ICcGpfQNB
nN/3irM2mXNmEFmX028GQCaNFQklf34rdODmuqGnlox9Ofz2c/MLYqy2x66K
ZFhMaHQJbZqZL0+R+/5AtiMOifY6lHWgRjSnpw0rdITgTs0qqNm08TWyxSV2
riwCs/Ow2RS84n+Nzmr4q99c9wQup2K7eywTJELW9zxyf78CT4VN7UQ3dipp
f+tI/9164DuH1QOpLXXhTCxpKUPvvHihTckCWGRKp4foHLVCqXlVyCM9xCTO
CHJ3aoG339FsJbLtOSxP/h0vfR8FMmIM6A/p6BtULNXktrriuy9FdIIbGp2M
KDVU77ia+qgO73hq0BUdsQiYu14zB0E7vNSnEICf2u6L4YCc06/Rz7Ze0F3C
+z6PEdNHcVOKtEv/22G5e/+3a5Py4A2LhNhZfbgVTfQNf9Qwqq6wm3YFU6j7
JPRexcaE17qvyNubAo1s79ZgvWpiBuv/ZxuMSDblALUtj9etkI4OcLc1LLo/
rqE9mOSFcOlPYbI2KNjzXKMVB5JIsye9eq0ZFn4GLo0kGvvGZ4+fQHjyk6z/
ic0S7atW+t4E1IgkFah8BaSxv7VU5Jd/rGqmNSx9FVKgPooqA6YvRzu4fHR1
ylEnknk1GGkr71Rmfs602ZcjNoLH4jqu0xLwdRwXMZyhMAqMZgQcHcfVym+i
xB8XcKwHVU2qHXWBlw3HufBZP20NSjWSWGxPUEdEj3d4GitBLlQ3EAgjL35J
ymf3BqIgFP7u/ISJFA1DRU6TbEiL8zFiDhNtRBjijRwLAiJul5aZSNicIX80
hciNUmrh3EfzMvBYmzyfttwbVBCcJeEwev6HLO8E8pxALJh2uEJEL37X84Sq
uJoD90PmPjsDwV1fkzV+TliF1YRd69P5H8E1PhguHpvhF6n4sWDVsGpL4oqC
ACVuYZqxh4aHE6xyjQg2NHEL7PTACI2eM25MEecPpr2zmx/TZQPPJpTOHBH2
56BEZnhigbx9EUz2mW3q4iCN+K0OJsR5h/4Gr9pX+08XMtV8g7J/bHvkx3SI
D0dJIuOpstlx/uhjIGDx0Gaw07BiwYuyukMEDAM8tFngx3YqwM+F9JpAbrMJ
IWwFHWCmq52JQm/h1heh2lqgfjP42uEhTJ5uKqWu0XMG8hrPQbq3wz6ZO/Eo
MlPVkATMIL25D+SdYhlCvbAZJb+qmqNsJ4SsGTTcWrINzyHXXwJPGDjgf/Q/
v3cp1ZyhSbPyMycC82iW3Zn8RPTGNR64opC1eymhH7DdMPbEZuoaXqaNUqhI
DfuuBrIzKv7iprsUu/Z2tSrWRjlIjypX7Ila6RCvP4rHntu46KvMJBP6U0wo
zNHY3/Hd852X3aWsPBD7J3SCvrxo9IfWIi+ERwPg4uaHQwqYIL9De4tJczND
CN6NaXUfm/gQP7f4Zu9ZWVcqJy4g3+Hvpp8uDT4EsGL7NR894U2hAKsZjyWG
izWcYACPMxVkSWcGGtw2lAdYwSgKQ4u+JsZYNCF0z4vT0bG7wrm2CA+F1qJb
TVDVZlxqt3pIrrA0RJk1UXvHNFiPSvy++Q4YQfE5M8bCaJTyQyAU7gIMGn84
4e+Mn396Xt3+rAIQ7sjjJ2zeo9hmpd1+yM9VXEid7OWkR+IBAcBOk+75niK2
/x803BUBofUsdUIc0iFikFKpl4lVYjMhBuAeAPi+lMeVDkkwUuMlqrcDK4sp
bZV66OHHh0TmYdtlYRIpf/0kzX+/1QiIWdYTJ5mBVVj4d9F4KdjqvJD4J5DC
nQ+hZ/53gAnYK+tpuAjSNxtj/E582PgHg98aK1ltToIDEvQI+2ZjMWa6srnp
TS0XWpQSyvOOjQmhseg3Nmp9x6KMJVBTtg6gi5rYXqNa5QVb9H1tieC/Daw+
bGie2s8h6AUaqKtKSHDv5+yfK0hlb/uea4kRxoa9IMIp6yYXxyp2d6NWzWlM
dWw2G3e/q01UlrBP60WnDhxpJB/A0JeYB6DSjjkPTviMt15Au8D5qQGpIGJ5
kH9t32nS0LMMNwOP4/9JgXz0aLd5iVL+2T5+gkEAy4hvPNm7SCx2M5Tgei7i
1s8P/kMepwmGif+w0C0ESaWLwHiDAkvpgJLBlpLoxXOE6OoJGW7SUvLDVT+U
MWQnpHyqCTpgSIiis1m9mIV1kYJwiqulL+T0TnevY4yTcYIFoFkgg61LqK/f
JehbchOQHVgCaqSUT2jz3g8soGj5+1qzGXX0nF7hrrmAR00fi1zvKi8z+fTd
Q8J/OtXL4BXrjyWyCxasjKOOxusaN7kIoQUoh9nmNrjlIr4joeC/EDIM9q0k
SlIaEdeKknclt00135gw1C9mb+VB15w0Tuv06lS3voB1WFLj8s175c6Vdp/X
MUJ8TOiU/yOhjYdzEo+8k5736+kq5PWSdGRnqRT0IQ71QwoRrPTKbJ6eU5TU
XuZXDrq+OATuQ2c44/tGZtpDJKurIT7s/ahCGOjOHqrvkumj7iETN+yB+f6I
qTWVJ3zK3gkRQLFWUZrlrja1U2HyBz+ciE7YxR/KiNVCzrFAKU5ONi660yO8
ADgOaCrd5Nec670hqNmwZ7HOlcDTRO+HcWbasc+0rac21bZ6CSBsvr53jsBJ
ohxItE/RW8R+PZZYYT8kV+Tm8fvMLF3rssLJze/DODX/9IhhZxdLl/7YXuwV
ItrmXKeSR6sDKLhV2IkOgMay2Ajnk3EfnaeOJbXgHn+H7tPn218NMErDHiP/
RkYMETRSGa5ypJCn8ZynzqE/WfkqjzlVDveYOU3ZiIfJwPOxp18of7NsL7jX
y9XbbJayqVVepqzPDTCrA+y5Ck1HFsJ9Jygdh+7Nvu/k+SN6MFj7u11jdhRN
J3NGf6NZ351elKstwArcJ8rVKwrQteZkHI26FL9rKLgElknV8NtETclO8fp5
yw3LgD+H1auvy4jSc1ic91KrhN/yWWTcYXokqECtzPNFVkFhtS7RPdxcHfmQ
0njT2psMOhj1Jcen0B1da+Hb1dl98Ik6TTtLVScrWZhCKSsFBTpa2ifsqekb
/29S7pEkAJTeVy2P2+kVCyfG4DazNSKju2x+zhAYXkKytQybv/VfaQcjVJCJ
gDylgd2q5R7X9LnzhVexgumA60Wob/AVD6d0M4TnvqpyC6Btv2LrNbOiSwoY
o7r7OVguUtY8F/vEtCXF2vAtsKRfjzHXKh8g4zlYFLVv9v0BUZc+ng/r0O7k
Nwq8jEeeRVkymnLAuUIQxA9JeiGq7HT/FdTB1MAhtRDR+op2uhYulr25Yx41
H4lsc9bWQ3sk5b40hPpaYOmSxj4jcGWo/9ZnWK2GC4rjaiGoIpLA69zb3ZeE
t3XVmrF1FHOr3zT8i+afFOTtJ2MDAaJ0GEDbmiTkBh547TfDDU0JBy5w/qCa
dOjc/0oXUVKTpQxwCaauvvag7op5Yf4fqG3C26asEnoZUv7FdMP4lBc15kBd
9bDZmC+MIe/ADm4EqnjMwqhj1Ymj8iBj7WrtnohB6FxNkR6RqCEVFtz4GHUC
K7nEUDN2ACu0VjbMR/0TNSmIRKSpc/OcqJrWzSTppzw7BrSLusEV5bxbGTne
bj3K9kHSaKPj0E/u85+OLSDK7VfuitvqH5vb+eTaZXssHSz75akq8ZJWZ53Y
pIVCHi8c9qYB/GU3KAAv3ExZXGKMrPcJ2lNTZv/RN49ZANUHUJWXo0nYlq++
DsidBBFIvaak2QCcCTdpExpdbN9Y3xGlbppZEpfZweBvIQSRUpJJih9XRX8X
UeWYnQr2DNQt3+gkyKNhvM78w3fJPZdzNz213VdXSJm5OMBA5RKW6ksjhk4s
M5GHYNV5KHAoGjEQMlkm4DWNUFvbu3kCTsKo1qFffXgKL7BL5cdIrmjKYhCR
CD2y10iajF0A4GuLrQoA/x2FvFyf9ti4gMU6uPIFx1FlojLSkr0JMiEEoRS5
LJn6jS3uqN3upAZ4jWVqYfuJoe6enLahAFcS/SPgVZ2JQVCeos8TawmnGREg
wy0eWLHn9Z/a1wx7G5VhLr0rqHPI/iqqsPxwIyj7soyqPjjcTQJyKEFGTtk5
MNJHMRbCleJqd3ZKApB+Pw011+yBc0is+Nff9VGlb+RMLBo9By/pekU5jYID
YEP4pffH20+CXh+7174cA6GygHtV66nySPasV7yhi9s2+D8zENh71Wav+fwt
MlzgP3KrNXlFkNJ5SVemYYj6Pg6T1u+HVGT3fvzMkLo9XDYJOM5xP48ysJcx
6Lc7AvWM8hR5yx6zrTfKklVmXw89nFlOAtrTdvjr/QdFh/C2J4crtaxCTGfc
k8eiJFX9NLB/Xa0qzCv24Bu1Us8GnPeyPCgMo8LKX0SxRvj7GTTU5OeI7mz8
l07r48WZU8ntHr2iB6MoaKIXGlDs0e0BPwzbqw4q3SBAxhKJydJ1s8AeWmEc
P0ziqwwahf9fimww1txqxOdBupB5dGa+fc2eZD4O1bXi0iz7I5tiHSfdk90U
s08jMl8cVVv/lGDIEdcu2cJLGhQEWes6993dAUvCcI3Jglob/KZqSOiI+ZTW
IH4teREJjsz/yYs7di29wpOMK9n0WBW6DPKz8yS43Sku8v6zqoyCLnokUSk8
qOO+gdIHKB/h94Pxe59EcMahM0Wc1B3IkrQIZQzzTVXwnjkme9gl0RyS19KW
6JWPy9GkO3RF3Eosg3kbkm0s1+Loo+VA65UWAFCr+ZHn1Km0+bwc/gWwDAh/
fo/8u3YLC0XqANJXXfDaGYSJPabvettKAa55zE0/G5c967RDV/C/FCLUhlwO
UOjjoU283Mn2IzQGk9CaQSEndyDXy3Df3qxwaK9tuJXpI4ZcliDCA4stJeKQ
8AJLXPPNbrTfwUlthbKEFpWu1WtEm3dfWr6BgoEV6m4ZULN7pkales2VpGkq
yBf0Xi5ke6AGm+elo2G477WN6iippUuxgybollEtLlD7JKscG1nYnxfViu84
styYhQN6wJMdwp9cIqAsd6/7tC/fdH9qF8YMefMz9t0lMLGI8TbYHsWVt2Lz
0/XpgGBvYNmFJf3Xsovg2DGui8pu/kSiOuzx9KV4DoM6ZH39DaoU3l+G9KyQ
viXaBVDWvoRz3kTYOP7Y9rImkWUZtW2OszagxMghiK1+9u3R6REyWqhF3L2W
aBh4UmLTqg7W3PIPdT2ZWa65/3w20CCe8fcymNfhO+c1QqXR3uRNvD0NrRBn
KHxcGD+c+zomnhY2VvEKb67im/WtrjEQRQTAZyD7uSSIBIfNgVjj26EGPY1w
E88Hb247mHi00bB24q1+WLOFPGImx6E5q7n47YLGG4txSIxyEY12c3HloOcd
gZacO6QWRltOd8/rkwvVVX4sSxf+g2NhU8fP24VdgVKIp7gCHxF9UY9J1RHm
wJYSj3hvAL5bFqWmxMulIRUuP22K5046UWkYzSY3IwvkUmnn2z8AyWq0DppF
wZjzL+6yU+55YO9/KWxImjObjKvFvlcZv4pw1j11d6kRwK834rMXCw87xsNj
zzNY6vA3DCOGLlyhAHD3zrVJ6BVC/17ooRDLc/Vq9SVclYbGpDFEcS2MAZSS
6Ezz0NAC9h+mqf7fpyFH0Q2v7oLUQzkprnNVjX99ay9K8KotY6jxm++w1iJX
4gINNJq4CiML5IdCjhLRtZKBJpl2B3UKkeQb7cI/+Hrjeez1307C0bwGgvTe
sh0kRSpafO2hMrigkwWQ+gGErt5EOSAOe8cNpFTkf5u0rKwNAVoMw4JxwO69
2fLei3Ny3P2axAjAEF/Pdl3jGEeXEIs8kmL07UO+o0+Xa+RMisGLEcirgk2Q
ws1SDFiUR0/P9xh+QnoF/xYorT+srsmgvED/pHqgSRcEnWS6nYQ1s+7QsaNF
kJcSoyBjxYAXmlF2l6kI+9HNQZxYTDdvMxBHM2SfpfYYwoKYDbdlsZU/PZI6
r+37CCxNAV7CahPe66ZfsgcuG5jt4C+zKBlak3NksIFX8Sj7gDKoXeAjmrcb
wSqVAUKH3mNpthrjtYFC2mozkYc/tF3ilgXek78/cZz2vUxBplh3/euJHn6O
vwo0/mIYcTOvT0jtY6I2+Qfsro5fqmAxoDX0aCjs3c1BE0ROvDxIlHMUF5wE
79fXKIVqn80iZWP6Rl4JYc58KAaxp+aMb9D2sf6zAEfYRO2i6qG6Z/wT8XGL
W8dn/j+H80Oo6Jjrwv/ICdKT+8L/n6kFe96jQ/6JndxUHFE9At7VirSkSd1M
BPpOuxnoSX0jGAmsptlcJH46jRqkJs/gop34KOMxlk8v7lsd626Ia3LymfCC
kQ0FwuuQJ6eftxAfzcWa0DGJL+yBxeFot8XTCh+4QcbjL9WN3K5CZ0khBymx
8PA3MeFbXNp2gpLX6k0VY1Cqako/I4fiuvfB4ZzDB3aI+6mLtLBzW8vj8IKf
NTVqfwDtswxUzibnX1Vmi10KdDbyQOQCokC+eO+cwaERFKxfCDxi0L6T5dS3
ohjSuz/ZfflNsUTFco1qWvKZpRuKiCpAtpWDVzzeEBImGmZlAxRoiqTm7yMA
bCxNlqCUE5xKlTwaUW3gJ4P6YyP7RTUBNCcCOJkQuXUxaihZcYaQIM4Hidv3
L3z+OjuPEX4MQx2Use0ae46bm0QKsTE5I5Jrfe1GSdZbR7KtMf0JpCiZ+tZh
ir71PjxlDDCuy+NN3SsPlDSUMbZRubuMtHhmgfrWar4VELDwVkvmPn7/nDKq
pkKzkpOg9Cpt7LEWEw6zLr6eHphEA4Uk0MjwKFlrvUuRjMWTOUiXSdVMK4M3
dFdQRJHD1Go4h05eUKomStIhtcbcOOoxb9wFa+4S/z35muPR7Df4ecXE9rBc
iuB+vHzzJv6nC1N1QV2j+dSbIug/QLB2SnhaWUacj+2uBWu6yOMW4Zsel4y8
Cp9yuikAdp287J7wiDLEYRUKssAvhZS1QtTthvVKKWy3SijAwOZPkLo40aZZ
zzBgxlku8u1U7cojNO8bBdTRV83HzZNhInWyegnjLluxClYuyKOcniNILJZn
OQjhSOF+gqvemqmytKo48vLMrM9Ue7qfcFhbHOfhtzt1PL+8zFU2DWZtA2NB
2MDUZU2ANpIH2leuE9gN8a8rcWqUxKrPZTxQlsOwB/SUwo0cjRJKQ19F0DRn
tKl1XqE7+rXFB0e9J0nCaLkw/TDZujbMVaElQ7WebDlWnGg8EMg/LswSNt6y
Wy+SXycHICmTAZ3Ex/Qop6hGI5R6vDQ8tqB4l4S65xQnBPQiPiQCZ9hJYLXw
YtHoJ5vgnQABcllBSo+KSSGDDezrR54Zs8qOaa/jV8NGZ+g/TSjVWBAnL6ZW
JVwlaHUAV/qHk4nJrfbDDbO1u5U+5JGnkf/dno5Z0z9lhbuYtkAJ2eQlH2vP
/azSxmz2M6IEFkXi/E9HPzCaQvYqMib08FZVqDcfNjUocgD35EwBeFWuyfOO
ggCbi9eBFZK40sGCN1Y/7BOqex4RS9nDR66/h6lp/Dixrkk7Qn2NDzK6jEcM
9Yh2YgIOebY/bwwQSnY0hhAZ0mr/fko4aRAqNw2C3Jm2PlAQIcmXHvk3Zjod
KxuHKYJRDmOMC5jY84e+AsnQDsW3nXuxvAtV0Wgav4Rt8RbBSOYLR4Pxd8na
Y7Xo5D9pdN7XrfssIXXYvanCXtu/4g1c3nLKfN/3HibQ2hr4YJSy7nfabLOn
QoLcwLKxLBbTtrcomKvu6OGZJ9W/hZeIqWmkyLAObmK/WKni6QnTYyB0AOMf
pODy/kbaOD+QwfTik5r6YaH3TGDAGDvYfGv8LxinaYwCHYLqf8Z4bVIH8HTK
Z10659XDKbutwpG+Mo0o83sPKVATGUH/0yp0LHmDd0SzusK7/NNJUby+mkp8
pr9nOMNyaCyIKZmuEtdnVKy7Awl5LPxR086S0zco7wqv7erqqkZy6rqjWl2k
fg8dekWZKltZ2I8/KyiM8HhvQl/tXpjdvqPwJ2I+WGfGAG/34DYjGF/VbXbX
ttobyBJnrPlGxDHklss7M70dimVSJdtdQ2KXKK2ykcFRP4gnXzcpqq54VHPv
zQLgTITy10roCDjo38Hi+YrlyWQmSOj0wXswgWLJAB7E04AkE3RK4afnbzza
KwsZxT/POXAy7L/HK26FEBVpQZfpqSCk47rh1CkwFddTVOecbMy6YmN1FPAs
XUS7HuFtX12UqgGLFK3CU7FhzFoFi7Ovo9ANYX+PB0azZaix4WSci2W/4sgQ
rfo4WaAS4ePgwL1sZBdlsXhuWqmNkS5UmrvJUJZkejh3Y/sI75KNtw9aj/3A
AxfajT5leqNZiPSmtSz/ooPR6gig7s++ZjuPIEv2Hg88iHzQ2hj7RcYn+UG+
jOeD2dc6dAeHmjErUcRf97sDcFoTo1ni+OWoJLYdGXoqQETk+9Zrhj+tgbIt
0pseLaPrakH3FR+8LUDMKQ1d0sSRfe6SlfgqeQ6FzSutmo89oujbJ/LXa1c6
8/PawQaTjgy8m9tIuYMtHFkcfEk9NnzuZrESrykDinoaWXExhRRXIyresIky
dgyCUH4ukpfZTTGXLNRJqfUbAgl/LS1/9MyUVhXCsStzrfT6y/W/nR8tHeo0
/LAAySndM1MKKS2hoAzTTBg5qhEGv3jBDRKRfcEQcK7LNxPOSBNLs2i6OfIm
2gbVnrx3eKI6Ko4J7FjDlPDlu17aSOk+/7yvEYJDoCLj+9ns9TQYopxtwDFh
jym5L51gR8ItE0A3iJmza4YQQ6Lq8pxaMAlh7iwaKBJNtp0wdmxek9bFm3Il
o/EnacflwwaBbytwX7h3Wmb76LjHwiR/pWJ4FgFlnVMqszM2CBs2hmHBqjbM
9r+JMPmLfG9kpSSEXdgpk+wkQBZSW0uifZPk2nprRRKLIWbgnCa3WwNWnCR3
W0BHicj4g9LVUP10qj04c/z9GIV8DS3MMU82QY+a6dJXt5g94Y1zLi4VWZwv
d6q2Is9I2x3MZBwMX8Cek7vUdRbLh10312XvKGpZecB6pme4zVj4gQvzFJ0a
O/8Mfi+vJU5FfgiLOMq9raOxnyrrsS8BitMMDMxM5ULKN64DkJuAutY3Gpt1
PQWTX/53R5+jBjLZvFoZmf9is1bTEK9dACkCjrwLwW05zEbuBn23f2QVyU34
c3x2yOhmxvy96XMTQFgAIpXApHGbu60Yb5D3M12Poq7We7HGxweajn5MSc1z
ukur+mzaA4pFTfsEiJ72LdimUDrz88ctymjyz69+yKTDtloyLfcfiwipysih
/Hs79ocApfP1YaJrh5jE2h5/Ly+PnKmSdYaClZNl25HzxNMkvl/dzV/vnIFm
W8U2hwnsI0l4xoIwS4exe3KvZiASXARzxR4tCa5t+4l+HdGBQA4NLzWNmINW
lw0DfSeGtQyi5+HUzUjF2cX+fCjRcUYhzgV6veCuXR/+kIBZC/BVN6BLM0jo
mlCD+BhcIgooyStjaqD5hqKlwPqogqj+gBLIga328xCB+y+3wlkDvfGSR52O
4+QaHqROgOXXPMwygGX9XjRfi3rkbvbswwWScMzghO30q6nNvI5CFcxhdBI9
1NdCFcaQ62wpCEHS76gYdOTNgl2/cszPMlqULTfnijlg6IkKHPMss3PZkHCu
YN0QPeLmYvgTzgmZCu6pl7zdaWgpManbAru5CCHLwV1sALAEAyYC5rW8gD2j
KM+kqEWXH8gL1GLydtstdiOK9T6+VGpJ8w4GYewUpxGzr2wT4sSuerCHuzCP
pJwomQKLGaWxnNCDoCrymjuB0j6XUwwQ/2FWLKkXfZ2/A/M7IaII+cldYvra
UkYq3l/G3v1S355ShVma40KNeG4s59tnECUkEM+bucvb5FC6a6uolr2R7s0j
Im+hEDidFiFg/n1bkSnqvSDlKrbdFQWwKb18UGYEloXMgYzWxjkYK7ILP+PA
WnJcZ+LWPys+FePzqPorOQLhTKzAfCl4SCxAcHYAMkbEZIHpa8A8uZidg4o3
5bPhjFeT+8yleJ/vlqG6fGMXJ71ZcUIvrm22N5PsxHIKQw2A1ghofHo/0xgy
J1xW2GJrA23/scWujPoHJ7D8PlMrjZ4qRXAwzLd1dkwjn4iQC/qFSOVjB8QP
vffqaBWdSNgytWTeS1GVDic2fWMZvbViQ3P/GyQeOjYT8NUVi/RX+gEYZ4F7
nqY/zvp19y8j+sm3W1JZXC3xS2Y/vHkh4q/BWLXYmQzu8rmum5VWBaVKnY9W
26U866I6zGXE+uS9sugPjPLYKYoenMW1p2Q2nw0HRit2dLehy6wLX28apx29
y8c6u7jWuVF9DQPVGq0RIqo3N1p6WjqfJ0LbePgyns+vNYW9wMbKImt0KHjT
JSD3cb6pyVjqDKthuxZtl+bN4MdqQiKCi4edWHTkUtQyXvvVJwAVGC9NVTQJ
qhRno9bJK+w7A2Tl7xH0DzzQOQwrDO+EgqVYbA3/0/IPrhJkjFgeFK/XEdyj
ejBf30emXeTuq4PPzFZoeZLXMGhWz4g6qwwMB7HYbmVvJpMn5wprzraL/D6X
a2cBQrfQXf01aQnpzEkDHAePFK7YJTSuQTkIPBEKtV8s9pBlHarl5wunhM/Y
DrO7rebwwb3JKTmmCSB8HhEMLX/qb6jvz7TG/PdXhXwrVEok/EDzEfhnAVyE
MHspd/A4dz5JZ0+QdkPMkQ1HgZfilY6USoCgrafuqMsodA564thqyVF88F5/
+PZC1uG/c6QOicc64+89udL4PhFDKULRXM9FsvqzRZFV0cNY+g615OyGD0vp
soduFEnjRPvtR1PFu3n5wF14sg+6NoCEUCGkMH4bFNaPNjccU+GQ4BvkeXGz
s0eCLULf1caAfNULFqiposBIeOPCat1LUcUPTP70sutW6qq69vU8CZhEgWNW
5nk5zL0VOz5K6nC9gShnUnvjOxu1+q5qeq93EiN+e6SfiWy2Vu2HgJeCb/rO
8vas4fvB4qTlSH5D9Nd93bkiluIgZLkdq79BFNlJseU21pcNBUUbeCNdCxDU
qPyOAP25Ghb+dPEMMMnKbCLoRQTxBcy0PNmrOCD0C27cyiT7qaDxVlN7lz7M
pnsXA9pIX3fje3XnCtE6XuznMfdb0WXx8Qk+pfCzGApIVYmr2MZj+Hth/vyr
4avW04zJ8Qq1eL4ApKwXxNfxT03EMGjbtX4+oOKQHLLWJRbCPqPGbQDBWvPq
pBPu8Z4tANcbkiGUyJd5kGBvWTrks8omlyBjt3GMW0hF2lg8HQZijEuIV6cT
q5F2EFsym7Ul5f/6msiB+gVD+KQ/B5+j+rU1f0wxUOE0kP30uHo2HkSmY1it
+PQN2JaYCC/Oyyi+4EC4wfi/VcSSi0IXQSgBpnfgDyXgAkOjtqWDPzPXgdyH
6pOBOkWs4r3JgeUZ78ZMhYOs+aCYwgjs+hBFjIKRfuDUlRECj9iYXHQfWSW/
uHM/nygcp9SOndeGknwhXsjP2d91mXQWPkqwLh99CdagKZg12ToStXouvRpu
PPKgxn67/r/VrSXf6e+nDnM6dWYRfZw8G19ufBvTlgBOB2beapxrn+e9lr6W
I5kArVvl/jbf71bBppqYNghijqIHjMUvkeKRcYr5PZoU5aPKFQQ8XD/DsmMs
1Rz3OFzfGgQWX1ooSQ6JgT24EZ1TpfcTyWeB2GEfLfZFpgOPpNi7D4eDIG1o
AuoJ7dC4XNYXEvRbGELIIEnrqgvvWbOhH1zyGzAQZsRtWThu0eFk8gTCxQpl
1lYrzq0APjOjugkDSj1mEfczw5ADoXbP3HlUkdOZWFzN0Pny+GcQeqtfSPQg
Adv+89g1M04Q7bv11kQP0FSL0mq5Ge6WQE3r7H+uARocAuebRN1geTjqzVvN
LYB6OtZAm+pJrv23TWf0G5oneO2rBof5OoZ+bHzP7s+IKk9CG8Ufs+FlsKIv
A/Y6I1QHDbUTg2Y/JO1dUNaX0pwjj4Ocqf0OAO8gPUFOFz/M53hTdGAMRPw/
5dOdvt6jqj8AivupJi7/CO7sLYJoZ4JUUjoFWRuirTcUZPUubPnfLmAX5T23
kvRtbqKFbrhQCfEly5AfchHS0NlqzC3AQ86TSQhKqSjSgK0tE4l457k7Df2w
mPa0HU86utnfO2zGFkH4iL9cy8PQ52opzz1vYYySIGuYF2yNlE8vg21NeCti
xNGIWIdP9mUYz47Lt/75qCohthrKvoTCkXa9Jddhk7ThXdHP477G7x5Jz+wd
vKBwwf+MiDyF286sFvccA+onOZtTmI3pBPEzRvd3ODLSIlqvJiFWFlY4fM8C
I0BTziStV5aNSufWfZ7u7FE3JJjh5h2FN6uKGbI1HcpeeDlWdyHvDGPXGjhN
7s+1+Mv9AXz45QTPv3yXlOHSyA+ahQr8xrvuizn+OsZyO3ozsWHpdT2uxh1O
UBjOWktHpRUjYoAdXZzO4bTkeHr9mPYc14ymM3WDZ29430E2xIpc7LNXekFA
YnbxyXhQ2pnlZ8dodq3QT1Ts3wdwOcTGm9UItjLy0du6BJPziDGru7AxzhMF
yTsLZfSvahhF6jDe3YE7gw9Du7Vlkn+EwsWKi60YB7zW6PNqCcjnYg4tK862
YPsz/SgNfGd0xREhXNDAJkz3lUCjwZKirdh/T/dD5BrIRJoj7MiFQ8ID2KSc
lSTQdY8PZql1gYDY1KOcubCAqlIalTGiFjrOVpS6lg12oh5aJs9ZMn0+GLUP
sHCQwEPFd68fPdAkBPi5U7PtQSuDewAIYVDpRZV9Nsu6euj8JNOzy5vqNFEd
904FKeLjer/+7iHRZJGtwqN1f/hwf89cvhZ5oEDFrzPkUHjx5izv89QR21y7
SSWQOXvxj2zL+Z+wUq0pCE7mNM4r02e2NoViKtqWRi5bw4qXzxIX0JonChRd
Ch60xmh/uLlo4rz+DE8SF3Pk50DUO0WP5kxcIIRDIq/LYFXwSCS5y4+ulxc5
gu6gOAEJ/ho28z3QgFNwrQPSmHPOHLbRpeva+jCA0BGrqy3H7NRjjlbvAzN+
DQ9owK2XfSUJUVsFCq4hk70L9AZ2602LypDudOW+3SCXr4WyuLCmCwdS9Lop
OVB5Yt0gNqARjZPox8/i5Epy6YPPtGLPpAyBzV+nKJZ5HbHtV4wNv8xgc2pA
OwpzkQLy9LeR2f7wI8EcIHTpQbSxvkj+tOFBAUOuZPMCmnAHlIrjZhl7bn6S
0V5hXCmDg1ROg7bRM6fsdRe1Dyv7xhYge+Q+KiMp00jZTJPyB8n6fLsH9azM
Q5Lzduar/Egltk5KaVzet2qVYUjqvQ8aC9MNCZUb13Re7XO/1L9I/M9jm0bJ
bKz4eUaZtMPf2scpOsEs2W6UF06LzuPAED0we5Lz1ZCNJnMxAG84Tkd9iAKM
quc1fpH1PKb8zbCBxKgcDLojazjn7HdK+ac7Sbjuki6IQnOXpqvW9C81LuK/
3BebKEIUcUt4HHNCulnKYjKzgDQo5428G/OQprSOPc5ejU5OWGP4MxeKIHY0
Xq8PIBN3kKPTHJlfxmxItiKUg5VfoXhKXyV7JeUvlfUTh4pjX3m2GunM8AFA
miFPIMJgc88mU+ALfyP3X8CXWg7Aa8rEJlF34AYkixbvK+CMKaRGlMjp7/dA
K2kxmm+yxZukI/mYmt6oCtYkAy6AVksPsam86dqnFmuKk6BV0Lp/MEGln/Oo
3yvpStxL6xpsLFcfQG7exJsFb6Xo+EDSZtsJpkHvcVqlnwDKWJ4NVmnEZgF2
2FxmT1YjOSEMOVT8pT4kq2TJVo6J4ddgbZWzI46G7BvGzydfvWnAw7R4LqUK
okcVLtG0C6mlZlRTg082WisLCaoqRkaFW5kk+SftXKtvEk+MO/RV+92yDHEA
S1FzUWp2ACqI6iNvEnuUGOyA31ckAH6R763dcxMbSiGZVH0qCWgq1Pu1RWuJ
uTWydmAFdA0jCyNX57itLjrB5nGMmeB4oAo6skZCpdt6QDE7quGEY6EmLlNe
Snu/JCEZUCQ1VnVjPaBu89aZ/NC/FLcaA+KoF2xmjm/Y/i67a86RiZ1dvFev
dY3UagnJlZqjRXfE9KrmLGArWV4sbHVI5J6EZbX032ndZh906eFrpFhFLRbo
n+5PYfqeNlN/Tc99CPWbrDIOB6stoNHRKJHtJGY+NGyBpf8I+kUNtZYA3bMi
Tpy4taAbMvLMxz6zBqFiTf/bFf8mLvH2f4YbSAjNdQI4lAhGzbsWnNr6BJiJ
PMhhvNc6QPYFFNRIppBoRtiLlCnSjSM723AiKfEpPOlgcblhe5geYru59q0i
udETN90n+g6+I2ldPxOYJS+SjxUtqV6maf3VciVSZmIkzFaXl1HK/fbBzpJ8
CiHb6r5WZKWn1fKr9s3XB9qiT9xXxUjHlb3Uk0i4PoJ2elE8mM1M+mRPk2LS
nrDtPeHZwEtaufOJFdTCO7eOMHrw4lp3Tx8BPno2EtvbkJI/UsmbBNl7/o2o
xno2C8GjZ/l37ieof6tg9hqFA65zlet4dblbOPvz+ekYsVNKimKo1l/DLXlq
NpLUnUR2Qgu12rXHzAgoFOKjk/pEr6gXoVPwdIFmm6k/D28BsgjbKAj7nvKE
kcTDbqzJhNWXWiOFX7jEuCOjRw7M7puXYPofqsDlIYc8uuyaVxsPPNCCEuHz
VmsbYpVfHRfORH5+OjEt0K00WrP2WeaAul8BySMF43/0vh1NWHnbLQUj+581
LbXwbdOLMIQz2UK9D6GQkY343JoEHPbH8JMSj1ChjWiimZmIbIuzkQqIQJ36
379fmlZgUxFG0jh6aA+BC8U1B3BCz9ANW6see6xqnBjJqMjU0OKwFURRhQDc
m0l1b/fs8uPXLZ3ltroI4FtwoFrQ29reeuOh6c7YLk+c2NI5YjHe5kvRUOeE
Ko6eSVCjVdAQ1YScNVCR9kz5qvhushuB8eX6XAqalgHf6a3qvvWtRt3UYhUr
iZUFHuWy4zaKsqwVJKmerVIzjbLLyZFBSxcvsCb8I4aAq2BMgeiB/yaqC4k3
+Bi5y0jffPD5OlUUcJaD7SKhJHbciOB4iif7Fi498HMW9eoGq/I9j0r6kazx
tJkGq3AcxVUYh1Z2/meGCMH74uyqhkjI3HQz8wc327DyIlWnCNUfQATt61rb
6JslY5e8zIWHhCu3v1MDdvPghVT1vBXAeB2zoeEn9SnbHNhljqW1p/TyMH38
mQbwFHEpDkB90hE7W6T4d1AAiZKCaNbwvGKURJJksn4Rs/v+oQGpiqkvOD7p
bFpF4mpNk6cbwviJezCSh3/OkfwIS/h6fPAUz9Tlph+rmai90xDVQRmFYoUf
h6enmza3nEvrFeUP6YhGBivEAhMhH9xke0B1q6W8KVUb1qk787RzjyzJm2v0
jfJuDKpISnSKlEc2G2JiObvrOiQHlLT8coOWF/IXjjPTXPWG5S1GXheNGCv6
FPG7Egi4RJzWmJHOus6GcmDzkKXcd5GJWr2r6tiLW1X7MUeIzHHNfBV5GdL1
NahM8HhB4j6Px5Z6lIvXyXj5yNNhp4UDMtbS9hBpb6CgQqu6jJKzEHUZwc8r
AffWpoIdggs6V+3lSVvZkTWxqmDqpDCmK+UGSfewToUK385d/o/IxHLGGlJB
35CdaTBjesqtyzSKXhIhsr4474ZGAlKZu8Kfzbye/8zIel35mJE6sP/tItc2
vsx87tgCrSKVzpq0uRghOhEYD/7HihIo5nWSnbGVDOy2UqjUj7sfvcwN3pdW
yXiWu+xVyFSovSNBafPqPLReWfwg9hYkeQm0ndBCRFGb77BYzRXbGnX1l5dZ
E+n+p559X/y5TvLiws30lD7I0jjCq0WUON9WT93wJk1yActzUXLuC7pW+IsU
TyQBgZ5QAr2RtbolMoivDLtMqL9C9KG4KdC6cpyp4CYbclJQ3uvFxitt9KA5
BDV0q18nl0OE/k/ED1Ft6fiepqKvC7YEzqIw3fVaIbjCzXTX68pFQ7M+mh+4
+13ZwudItwRK83HRqCG0VvNcoqMGPh/wAMw75z5jnLfbKyNSpFWTYF3loxwX
7/QDcbuMPFFVILzZsamhWKAVW/zveMr29UaxM3vi+jsgXIaWAvGs0NjtI/Gc
BacJQIwekqK0V5Erxg5vXOyUclnpYYnNS4jxfETgzn+uursV8pfrgrkuDooK
AQud7i+SuRV2d99BbZeu7B/QdJSv7gJok4mZIX5Zi2X0Z0X/rkePd3Vjz5Jw
lkxKo49m79esX/QqyELp9ycejMX1Xlxc+lN3IUyBBgZht4g6ZALgBDp31wsm
kWeCDydIcj4BUHKt8X8IkbujQfTUNAGwQHLZXux9ho4hsEYxk3yQVFuaCCr7
zNk5MLxY1zJJdy6pLqWBApkc5X0SS+f/9oBXcYUwh2xMcEQdzEBu+7R/qnjH
xvHBtKMbVvXFMINdwQmQBCAgNl2Ykrx40a8yL8kqorgBdwBQBm5bAcSNMVHH
ABLUyXCXscy48c7m3vwXhrneqJzSN8tIBlDvj4TcHeFe4BZ+EnRO/myu8I/X
PgXV+F7P6Jm+dBu+xerp6b8Gq9IQTJrR0673mfP4mp2Qxy8ayuTdOj7ZFlnY
b7gE7/5jzos1o1yQMSs44cfHEuIwXCcbHYDlqmKlA4x1EzMVXhywJhWD/zHh
WQmLIAE5s5nmAEfuqE+i7sJszsl7bV0s5GD88sYyRFPK9TG6Fs5z0bzDN7qF
++nce0N9Ovj+71uBg2ZbKI1MmLzgFSkX7/mSiDtzexal19Cp2QrtW3F467wt
GvcnIhdYBrLOzLDHBoYtB3w5Q0tzwYeJzUmP/zTXy+MVfOpL22WeJ0t7Sv2p
TiKjD7MInsKDXvcgCmFhx2RWsQZeyRpwPJrwFDusybbrcG0CX9Mmg0F0K+M1
UeCclWLK/hev78DKR6OwLJsEKjB/QXIEheYeAfWcEtIXMPKHnAUPfRnhzGm3
xzKyPPEnSmvM2wMaCshaeLj4MbM/oTHbXsFfALTAhefv6Jq1kThkdRXLrI0z
J3SJe8w1MqiGEK/hlwxxMwR/bNFtF5dZtRRxEpnC2sjgHQbj0w7e4qFR38/y
t8rx82ngoGkfFzzZxh/Km6xuivaK6D1B+FJwD9WO1FgYCqSQ8HB07EIvsylc
zcYE6ESZY6vPl9HcfQQ/suElliikQ6aUa0791t55umUeiSRmsBG2WcAzPPJw
2E2UeEbSaD7UAlaXiXWlpGcPY/wUm+QWIKuAsiGSQ26UH1kHYHyAO0xCZUrI
TdWCaCmDUc9uUyDv8Nw0bGJKuZamMT7APn1PVBbibR47LyKLFGgUnt/dB/4e
wkAIkvpnpTAF9/c6iqYqaisfWOLTTgZeEgHNo0UK3Oji4g9fhGqdWBms5nAs
1m8tmfPHAGG4UAP2OHZzqGOLPNw2h9iyi2y4Nj28uC6DG0Qvpu60YyHoxzc5
rSMo2z4XG1nMMwHHxuo0/cHXevYT0Gz6/g+6ua6jVM872Ht+y9I2Bix4aT2O
VcsZZal9BY8G3TmUGxEDJMMt7npc29GuiQDOt8TplvrQl/GlAxHVTFtlQM9z
bDUkC8ig5KEFLUB82+iuPN/yr4tVw5g3NOvoQWBiaezQwMr0wWUw3pYK75B0
S2w483Qm8l0Wu4EL8keZjArEZMXDl+6iavCIAqt5NsCndwIKRpGGClMt+BdG
mpym1j+yw6zMIQnz56kaz/L2Doo0/Dgas27nQRX4VFlsUrzF5K9ICHS6ZadW
02fdQ21Dv+QDdGW4rG4Q8A+Tr5fPOnHikG1fzaoYGK4mcNLrvZ/s7Vf07l7Q
F96l08Zis2ICTg/fsbfeIhMOc4E5mEooMJOCbdTCSUrs9tbp6OuBl6nscNUV
g4DTWoG81cAZ/CWmjDwEHlDu1DRJYNEgkxHUl3fIBljeG6fhDBMqPIkDntDN
v3FKgfeTQBcAAjnfutYjjtZ41fK2n1oMvfYT0BYLXLLTnsyZ+1rNGLDRD4cw
LtpETUC4OQVZTWcd0ntGpjuYfoaCWEZxnCKOU9qHyrDh2kOduLBnAsAmDeXA
jsN3FefZauPMhw6rz/UjHFUgSXwNrJ6mXY2TZ2A1/8Uyx6MxNIKRxvHSalsi
/3AhGh4DX3dI9E077+obgAPG0kakPG238OUbTME0qqmi19h8NG5hDAaWo23c
Wnm0NM7xwraVuUizkEvfi6/N7/tWxvJsb2/i7fdnp3gX44XF+BpQ2Ks3PkUq
DIC8Y0auyHQNKdUHZ0bDfkNyyGaLpzkK+KCCRG5D0EpUJn1uXXsejmTnufWY
hZtu19SC7KB54pu/dD13PTSbXz4XE3b8Y1bopkw5+wLtC1WQRNwWKZRVoKZJ
o6QZS94NKb0nEKiDfTxD1T/2C1ty56tPy5jPIH0TNF8/DQw1VtXOaqSLAzA2
zusuEOlOsjEaIW2n5Ia5WUFLstRj2PWARbczJ94IlQR5hviPzn7402FDO9zS
qArNtZi8AeZ9d0OHhjUVclav4YOl56I9dNesF7T2wZrz/7J043MQRq6IZSKX
dw2kySL90yKVEswNYxsp42SGD8LY7I9slRFTKdc80MiXKHPxf6r0yn40M8LB
BeWJYtSwMNlJxoO9jzsFt5EXJDJVeUn+94iiM/hnE3qiHC0GJY6FlAbq4lGH
DTt1pthqOoHA7wfM3u8zr9Goo4vrwL92gS0hOMtI80M0kxP4gYgXgyWFBD0I
/4EK1kW5vP8dRSSpwN5A649FYjbED/Aa6yp2D/00mhOy5uLGZYoK0Sfn2OQg
fT4KZlzHOS/jRd4RjQwnwKE4u9w8ybOMPNaacUta/PZ58iHLui0T/aLLOj03
xDxZHgdLLfYEgzR2l7wbR1ae70ZOkBQlImxBMuJ51pjguFZKVlG0a+2Ja2A7
lBXwl9dsYB4eHNtp+GLmC6KH8NbImMEPrOu2CNXiwvvZhONXASYd6FhSu674
4d5qAxdF9L+v7J5/SyRZvzO3SrCCmvZKMMFSt+xolSnYov9Hpgw2N94IUvI7
9vSgbyj/73JDr/1qcyQkB1y/0ck/OAleEGOTxZZ7f3MRWBxw4SAYDl+Ix0TI
89XHj/0b2FCvH+qSjrbDqT0kfkFr9XU1EOdBXnXCQxiLl3BvVw5IdTWquNrO
f/8x2OngcCaBoSeKWQsa6OyA4K5Oqk/il0XSrXpjEn8W1JbeUsEbcshKwqq/
/nxOJJDRoi1C37+ztXHTdhlgWR8lr86rEq+qYG5zzoEk/H3xULV+eWPc6B20
Ub872ZnK/5seZ06lZRj0ce6HEHdvmqGBxHLR4RYGRNors170s6NsmgoUuE8+
ydXhlgC7bfJoO/kwELVv2km/u8m9KRE9Gd6HSdKLN9Vil0kTrmh8D95kPdU8
hIFtqNOqB8S56LkcBsdyl43gr5uwVH3WasZvsINWLqMjVHFxTABvI005oFcP
2C5X+Iw8z8I86R/2eq0FZRr48Qn2dwbtq/6Y7tt4f2Eh+YihPobTPrss+arE
OfuKQctOHHkJYa0dMhqqpz28ZVTP5QlE0+a82o64UmvtxPpt+ip9RyQWeAc4
+517UOoPN3PMkxrA8AEptL/vJGHjjQvYnYCHEuxqhN9YhlAu45wRvRKVklqk
Xgr8qHDAPfI//DADXeOnEspeBf4xzhnvw8TxSr5rF36LQeyvmQhHnjILvOc/
D3C+QoApmowc+v0T6W2H7eRYEGMVGa3hlh5XHsgTQ2LwVlZodY1wA4IGh9YB
CHGmDynjxC2PRg8hGorqRqnai0PwI/1lV6xvCR+x55RbMxTCqA8CgwX6Ir+p
vGJwxStIy9FdQ+N+c9Ku8xoA7yMRWg/Hu+NvFu5d4wbWsmsUqaql7DnTaVB7
BgC/5Lz+HcUqjv7VDZ25pqIzVodYH2d7hqLiCvyphcCzOGWMq8LAiKmNhyaa
j24ue1UCQfGekBKfBaQWyv372ge6ihcPZ7gDnlezBeySRkgtaCqGNw7ziojc
vNQgxcw8Cxzv++nXGtzDcuypAFU0o8ptTE8ILbbSNTg6Rdax2cG51CLy5X4u
8uUXD4HkuoEM9Ly+D95lXVLMu9KZGK7B9HX15U8TxqgtBnMndW3kx2iVQj0g
fRM0oIvoU1p4MeZ3gpgpP0ndfJImN3xShnv+PHtSOO8cH0qhudfvzFJKQL1q
Bf+8DmR5NVhGRy9NINP5kRSBhRabPAGu5wR47IkiCHV7LBBNfRu0TubYdDGn
yYYfazcIEfaXCAUa+bDECg2eeEYJSk7s0vSuvPqm1CRtNZyBQthwmbZMFo9t
irCrrK/236Xuv4yLQ/yLNXAKU0TK5obt3VtYrpe55BD824KDsYTVqEPwAqpA
kNDwazPtmwmXH6QlnX7lNxwmKJgnen0LogGG8kc/tupii17/Y//VRVOB/N8y
nsw8TXME2gv3ffBfhGFG437R5mNI9MyKJSnOFfR3600y/x4c5ebbg6zcp4xd
kPF3OvZftQnfCFEx4/cJaolqgvHxvfBAXjCon/JTvbDXPB6WUDZ4hHHmAaYu
mJFNcWT/IhjcB1lXSSqy47tf/2Z006udQdC4xBatNTbMTXQNsu+oUJp3OnXd
ZCxKJKPRou2rr2GAtFVe6s8KZX1Oo0UsVWKSG5bx+sM6TIVg1ofjufyK6hi4
o62j//bzFz8xRdqtgE9rPiB5UNKsz6SgNGh1MN+BlDgMwPlouAvEOKXm2R3E
H+JSbgWS9suV9KMu1RDTFmA+r2greADaD4IWfUw8CVuNL7HFfwnZn7BCotBD
L553udQE52H7MtuR5St+D6+Yn4lPcBZ+fdzElunP5fy90g8mKq0EqubnDE0P
ndZp1VZ092rxbmUC0ZBrUKo5dZR1WsQcfXMszekkYpgfN/SRt9/4qmR+hee4
8E23a0eRoXJTh1yfX0DnxRSNdiq6S/4QxFQPUkBA2FM3UrStD5kViqIsMY5K
78NMd+ACUTiJAyGyaMb82wC+9ZnhYQ9LG0jTLZyGtX+sOSWQF85PKvwtYiPT
TerA/Ye8ppTmj9/aRG0ivZYsvZ28otmg8onv6J870Lf6zjw2AnHJvaMg4Crh
xL3B2Hy5ebZsCRHcFDrg3znQYhNuQFFoyl2QBgyRCHab4p9nAttG+jWvNO3c
XlYbYQAmZr6ubxFNwx2XaqAwsFBH2JfWpKBpZCFkNxEy6S2m2UyKkorjBCBh
gwchzuv20f/M/DAw09HfxTZGXk/ZI2KXX/CBT+RYypwM1Z87LIb+TRwBdXUj
CxX6YHpLgkToSWQe3eLbVdbU/E9e6S5AIFab7F0DZ6iHexpodCtEUMl67pTS
WyKMrf7TDVxyEOXrTdXCZGI46HLTIdaTfrP0aVS1pCO3D2cZLhfbBk7FtHqD
KreBRm+31uylB1WxAQv2/MEym9wMLKKp5sioB+3h2AxogT/cO24cExemoq4S
Dmt0VkLoJwTLfSoFOt87kQ8OtO8qadc5xtqBhtcyidw6xfb4mHoUF/kl8JyM
UxNTrExKtaJnak79EJVoPho1ZX+2EK9soxuXG4uX3OZZ5cjYtk4hrtbUvePN
msCNMJKf5rtZznSvrF58aFGyP45aWBEtZwB8OduX2FHImj6Bf8jXyddXA0J9
io6r078InaJydEL65+OUwFIweYrexrMMZ9cEldjgGVNGKPunVNAOvCS/B0UL
vN+cAu/4/ahbSY1MzSs6JiqqrQVEz84sIn06IhfA7Wdg1fhR5RV8fdvBH5ie
zdsiKA9oPE4D6XLfQgfj1/iPQdgXh7ikj4x8QllupUIkA12hAObFSVl+Wgts
aRh1UfzQVMXulpTFLWC2CWCpqjJgWkw9KOIsi8oQ0OkJOJJpJh6FgFOeUxyo
qVETyxGO0UYQam3DSxjO21e5C8ECoiwwv4/qX7fC4LKQioWsOsPnrk0DkZTa
HMApfyfln3Slf1TmICFFt41xeO1qm5zRsBJLbMUY5bdyUQZcehvpLjiGGiTx
9JSmVNEP5z+eWoi6I4PoJ4gZS6eYW4ot/lEzOZzUsEzYK23tVFNkhLIoO67/
UWgB6alHCNp2OGeC1ENnnJtRzQgzkLYiRtFE56GAbfcyJ2X/xBfTnixVwFxv
Tll8cDkJcRPTDd60iIfypae39OKLf2+qywOJNKiGeFGuxyaiSnhGZbh6kRgl
6hTjSKYR8jedGEzJKYarFErXkjGZKaUaI/o9b/9/e8LZpP8kClznpaADlW9F
1Tzi75revV+LMUxB+1XBT8RBUV7x9n2HB5PCBaTglnrjNrn7SzVg5UAQv2gw
uufug1HMQoLIalz97WUSJcqqPkKAguhWWP/N3CHqSPsoROsDAylVza10lVx9
wnUW/8QFvwiePAjf08uMY4eGyRMCwCc3aMriodoDwYveA3NQ6+Ld/PAu+jwG
sAcaaDD5R5bJ8EjOJgZUMielIuHwTd4NSukawV0UkHwZKbjPjrDC3sEvJNiJ
scquhzK6ogNSnY4jWqiZtbXBiwieg+unUskdCHEf7j1A/XICVfQIdKE4sdo4
ThcamUrNJThPcI5VptRbpOP57QT6q3P5vz9mzPbB/N7SKESLudffW0aaBkf+
OEF/hXQOe45IQk9M5T949UnIa1g/0sxD0n0Cz8e4n0HrNo2KMeYljt7GvEHB
SfMOMWPrDOr3ZCGWFnMxdsiomYYFYeNnNg14kaEsOpHbzF6VaxIld/mWK0ls
rzMKwMb41HR9tn7ecl75/7EjN2Ps1L4b+Z00eVWiIwg6ifSgAI06DUoxQGLa
1x3VZIKSpt+gUzMMjoUz7SviDbTBtxeXADDvE+8oSkcbPKNhmGidCAvdRMJt
Wo761xufrVCCho5c2fFWkyz1QJM00LD7X/6+hzXLUsj5ufyZjNcfO1iFqQva
y5Cyf6umu3mC3HW2gqzu8o0EyJNuE0LVe3X83cog+rumX1VEHSKxfSsTcS9R
G+J+xbNyBCHtzeuz8iyahinOXW4CnPZnrEHBaHHSlgpgu8pQEJC2Fjx/xwSy
aiMynXVYtzbDm0oL910wSwM8zVZRQANPyCxLV6qXqD5cK0HttTiK4BrB86j3
uBur8LW28QIBE+as+2W+uaZfEGyDQ4C+eNg5V8uiJn2TrWIfDWMLZRG5P9BT
h1BMwmMgmL61WRLfoY4BF5Vj0Bip0Znqo9zb/6QtYMUdeY6lC9tSK2lZjZAu
oMiLUZA1MzUyFvAfMllcD9hYvdWKsQluL7rVoo8DFLElyWQAaHin2U0fuORh
d+/60Y6kKkR8qV5TjRNf89Q9IcLZVDIyx3IKVUYx2COWIr4YOufYch9E0GRu
Fus2rlnE2NeBcaxUPAtrx+smhMfOOTCF5SlT0YF9M+p9LmFaoerLEq8C8FpU
WeYXuUY8XkFtN04o41d4G4yDghe1FdmESUkulYk80z8bI4KQjIhoH9K8X48l
DFDVJx02Pvg305BWHblKT5I+uAmeSBmUkaF6TkiT3kQWsBttA2NBMJ1KfEHG
8thRE/IDskm4cJdqAJAhjchBYygbxQsxl0/KGCq0k5r1dhaJBv4NXkbrbi6s
U2MKxVLEhTgwWDReQalCbZN/ozPj5pVLDSdrz2KRhRDHEonFvDWmUdPqOAMk
fAM66IqkiQXZt9OE1kJ3HL3IHICuKrnZSBpDAq0UfZrwQYvfqRZkOLEdoT1A
UHD9IvudSlymSe9GNfZARW0/gXBt9fdkTbP6XbA5xDZ0F7HbMd9tOILiQccM
SyCG3z8qxkiU1gkj7PevRFsMC0b5RSLgeCRS7ps87tOF4Jaf3ftH1qMrkRFG
3oO3RDUjwkvlHLaFVk277XAsuUbnmoHDOfj5SL+1bUR6rrWFSIJcq6EtCDB/
n72ANwMB2Ivq0EUqFhrnYzS4Ejrck310lMQFGunhaErTGIlvYYh6L6HjFNn7
Y27Q10vExDrA7JiwB6tJFwfSVtorVoZXIgeXbsVyM9V8mT0/TNvpp/uOOzah
4imlgR88Cyl2InZxQfTnkz1okB9CG6fNE9rPIYEazie/MZPqwb/SIihedhnA
JDX1e3xI7Ah8s7Vh27M1wbU7/5isWFc/38xkwrHFOgDz3OKp3o5CDQBoP0wU
Vl3zin9raKdWpgHW0e1R/PT8n88yK4eUyHk5lnNAMo+/wNoZKPt6b0bY4/Zw
P/BWS+M4PWdM0k8C+qJhFrZihzk+RZJkFkZ/qopovhOfa2BasiUICdZ52gAQ
IMXG/tcwSSd/ZazV4FFE2mulQJs5m3EWbYdqAY1ogBYHYBtv55Lw4u4qT7Dl
g8I5AdSjNJk09u40Hi8JNUe2s5R9bbe37elrYbvTKgEqaWmy1FQSKvbfcbd8
iD1HCmgxsfqtn3g607nkHPLF8OMg+0SlaTlzlaSf2nmKQ8gy17/DLTxis7LM
llP+BjMN2tE5CcCU8MJsodY3ZqavWwWJ8MIRFW1/9ZVt1ns/b8bprmYq4h0I
hlCdJpYIgH37VVn8VP2URh07t/VfykOmY73BL4+NIbgEHn/l2C/IQa38p4Fz
nLR6fexfwXSUteAfI/kXsRzVX7iym9vj3JmPdDiTOXeVA0hBPEIsRfP49akN
APoGrL5l5dC07hb6rZlJxXdeg0VK/84uIi8LSRIKM4K/lQhMFQ8VDfmI+n0i
a61+lfNvsxydqt6juc17Q8vr8e8B4XK26a+abOctSk99LO+kutsOSdDEacHO
mn7+m0Zn7YVk6dsg8s3ze1zsZEr8nDe333m7cQPmhv4bohpfXmgyIuFNYm6E
jurDtSwWtRfJxe2BVrkuYO9wRVwAGGV+GKqYsGwDmD2o4Kf+9TREt1l9JGO6
E3NPtgwbFqIBmnB/8BpBXxyuoE2Z29rMEOEu9NtYC6HzY2h+eNYjqCWadCOy
WYHUIjwBpXLEVDoI/VN+/R3UkoP47B++Xz0EBuTS0iDpRHp5v8/DDbFKi8m2
b1HZtmBc9A188zPTaq0YzQEeHgrJV6p9Sg1ZxwEviS3zZd8fLIVjHRMTnmWu
sRRgybmWV+GUGeFN9m/2EpKqAgDY8MXLxfUYsJDh4EZ74OTP+zTAjb1+4erH
63fucjQqh+1mf4OliCer804Cr+0qosQTz2ghmbh/8FJwD2hb+MvfB8cVrZnU
E+Rj4oMHd+7+7bb6Tmr51espswc39ojaF73TQUah6aV7DdH1Iw48UHcDpimx
yI4Fy86eI1EJk7IdINfyyYHuOGtXNurgE54L31AGJwBnSfYlKiQiV/WLmWu9
AETcyUO1lCbdqNszQZoGiVwzXZ1ekZwWiHuI37sL0N8a88CiA5jSlRGKHYCZ
9sJOsONHas3L+gC/tJ1XInw7Jj7i6cVN6OYeVc3Kjpz9GB6SyoOnlf1a5M0c
ThQXDSBKoHBpFNHBzo7y4AiBxYUUaq6o1tISNubbrlWUhW5a3nV1pExYZG16
8ebJF/ougqMkTRYwGLCcqQyeJLife9DGbKsxbKwwTPKwTSeJsOkDtQnxh9v/
bvJ0nbjBlj285eHdK3ix0ZHL9I+cQ5xVOuMU33IlmR8+LUKrzio0g5eGAqsl
56kuI3S6FenwRV8T2/TBJg8UF/mTqci+b46ET/+y3L4/Si3YU3NQ8n3ddZ9y
6KMsB19vPCKyrMoiRDHtzXdjgMtwZDyWfcYy1F5xzTqElAcFTLl61t+jJu0g
BFb7eatsrHly1Cmr8ceiGd4o5miU57IZ/9h0t/a1oQsV8u+1pZD6YfabXi4o
XJQDPlQ9q1SLw3QEJnbk+p21Z61QivsNfmKtnkRSyk87jOTUiQK+ssSw17ok
0Jz7q/RdgzsgN60Bl6dtqm/pbHq6UHOgPd1bsodtFICtiSbVfCSjgAS3ov0N
BE9HXJn5kyq3ui8UEw68H+7RsYWfHnTyHO7z1JsYJnydeuK/Y9CpP6WLRpKt
RqNGXrkKuXzFfQcGm0ZQIVwgsrU/2utKcC4mZLwmYKqZmFYqEOLNS2fFSOS9
FckI7lz+uWP6dRImjV+YqOPhwRg8Ev9NXNCsxrZo4t9WP8+7GYCWCMt3Wy//
yhKQTcY/Tv5Yyy+y3ztHzy/30LMxWREtGLGjBt10/7rCME++ra0bSGbVc+ZH
VcU5Vox0V9e4cIxLncN1Bu/I6A/97OgzjxsMPQj7MIB7Rx4WUcrPhUGaImDL
mNu/vZ2mX4jPiucWENdsjDtYbxplZPCUWqMI+k2IykXJIZruHtr8pU/ewlWB
lrMGsdb8Z2Ut0iPvqMX1kihDhzLGvF+OwIgFyBNoIf34uX9UEdCChB90eZs/
mSjV8rXFmcaEjpTZcIgmwKQsYImyF4Q7Zk+DBjJxji650ELcZ8RyJHiBzPv7
1asLQ0O1CsftxpP7Mq0ZG0H1RnwyVEEccQmzdoX6IvkTopfE3RRT8YvF3mYz
hxeUuwFtxBG6W/zDM8N4uiSyavYCVlhoWvLIXH/YVUlbhAAmtEpHfa8KV6jX
ZpCvM9vO0aUHK2ij2lATpabGADgn+GhN/RCsedcSWiUjxjgFLSSuLYDAdwST
ZdgdR2M7oBToxhavIYIxb87qbJ/MQX2Inj/5lkagdSC1tjsbhlQ8CJxa+nJd
6Z9EgNbyqpu0BFSCpur6kRhnHxgRivb+R7SF1DJsHR1vBY2Vd5AgPcrjMT5M
aGfQj3379ZnG2d29c61OrBJ6lH8ma5eFeJLIt/6Exu/0zCX0GXIE2xposcMF
FYfqdZo7ZdDsdmFbj80JgWpDhFE/PZf3Si4RmFQmIIAegDD7Smt42mFy3mjm
+QegOc+HiOhptewJ3cuhlTJq9jEuVZ5Gcysenp1/eNtaQ1Pcap7pH4HdInmd
p7d9Fv2fWMqbUL+ZApTyHVN8676lrr/+58y5Ce9aEtRy4j2Qf2jJ0XtI/K1I
ygZUdiiR92ajtEOpjON83IrIryDOEZ9234EWt4maFEAWIvAazzgEo9zsmA7v
KVM+3tDehgxXS+kcJitaK1+zZW6JHVmNHuXZsCVMyWORdzFzNFXeIhhPat54
7ouvlRnj+/67CQkGSKoVLY8TblkzlK7rKvelzI5yTQdtYbEkIc2QT0pf6IB4
DozLzBjNx8yNk53i/zwlAAeTZiYFfep5za76AIWNONRFPlWgBxgadrAwdqpq
pQ4XNC/yuGEbJ07Auou+F8Pr6RZ6bfryfh9KhEIvtN4ff0OA1TpMg10yNBoL
w18XZ+5SkpJIqaZufN1MM5DxKqnkz8CkyxZQXHpc96aNLmD2gfg7t6wiH7kr
rMLUvVB2lh/ehdFAkMjC5jBk+CmgkpPgGua/JrKO9me5rVVEp1NZCzFxGGVB
KBDjX+3w23SQjmP9MyJdjLAlZKjkXthRM3XOXTEPJKuveGvHsnZeXevbTdv/
9JB1ZInVrD9FgOH1nl4EaClvARmPe8XI4zu+a8nojW4BAYagZk0hLzc0REpp
26Kxy6zHvBLKRy1wIRmMtyOT/R5sFvhROruVXKIeWrAzzRBgzBvmGQ0hC/zS
MaFqlMWjBVNJimbk7fT/2y954dfJhOKqLqLkR53UYXqBY4lxb+BUW3bsStyF
bV2BpNwM9GWq26qVwjsevKQRg2KhIaWlTyE7Od8+NUSUH8EpD5kus7Si/ORs
PTQesoCMCSuhKex7DYaHxKdvkY2nkIancpZCUpnJWFXyaaY9E1x1NkAJuDy/
/8Km0RwGUN/6Lib+AXRMM9iEsc354PRdX1vNkNiyrMBgLNOlRsuObc+pJPNJ
CkTHx2j+YX5YspLcv/9/K/bLEgmC8TJNAx/YhRXTdHn52NNgN6t7QPoR985E
enVjLsKNRJIC4K62eoXyn5fLjVaFg1f2RuV6coDGKjrK6RjHOLgmp9AZOCcL
mttb/az2Bnkw/LxhOHheo6dGiNuuWQa7SAA7A4bX2Vgn2P31PYPXSGy1SRW7
1OubSC2MkaF8SHeiO3iEKIpcytpIDJAMEikuTsCO0w9wHLkA1PPGCQ55UTCA
SdM49y9tXm6KsXKZteKucMMjv67qhGjY6inr4kP1RG9Lise+cWuUII4yO/Si
tF61SiA3B51Y5oW1LHcs0HTgUBxjl85qJDf5L+iK8cr3H+E9fZ3Z//oO4Pkj
WG2uOSFyy7VU4LVDPAtEIdHk+59r5LgQtYwqrfMZrLjpjPTOXPK4IAYjsK/1
TKmNeJqLv6NbFP14PqgzxER40TWqOaOFA1/twJNXrw6gOouIrA752oZQHdAQ
ooo4m+6LIxggrqhes/rO/ytFCDGZwV/XiWLibryRDVQpX4bz7CDpn4qbqxre
RHJIe66RY5v7wEBA+cuM/jsdqMZ2ZjtvU5hZb6O3hZsIqCCucNW9v4nu2gRJ
4VRS7H764iFD37oTlspTlfyzdnDcOTk9IdqvFuvLm2dJKHvGMCom/OcnlzNU
gN6YNiuRN5HuSUYpGKbmBVQOohllIMvmkVWA12YtvwTw23Ov6qWAytqMpABv
HLpR82xYVG1lDjYLYalCELHEdX8NwpAIG7k/+ExBZeriy5xt09FLNXumdxol
q+C0C1ktWInxl34Z3KDgeVVTustk9eyUPqMU8weiucmt5OYItdble7jv3jXc
vhVLggHVQwcIVP+rEQTajio5VmqmlOyO/y9J5xZ3pxseqnJ63JwrpDdixvmm
ukg3CVSxwRcwSEaw7AQEUBWOS1JuaKYfGXQXPRrbHYw638ziiMo28nE24Nbq
NRtmBrSCJWsh+KsoinKLnoO/7Qjh7fEiS7oJaScWF6yNzTxs4mKaamUIw5n0
ZQLVbwgLZJfLaF4XxGeXoSgO21utPXxf2WEeC14f0ilEdRNw6gXAeAoTquB5
R49luQ6tP+7CIWNF8sm25zRnlGveiODI5zlqlsn+wRrbaYaaCCIDAQS8Stx4
ixVvu59MuaqPXSkzWrV0Vyveg92bjxQLmGcHJbffiD0Otbx2fde1QReZFi2H
j4dBuS5AykjiKFghTkLGZIAPI4ugvVcQEc2SGQo+aiAp3uXPwMD1KHYtLFsy
kpGSyzxAHDc0Tgd5zxBBOlqFFkLTkRjOQoFHdsx7IWi8C7yiMoXDXucvBHoP
2syInloHWAiGA3NlOtXdFV1apjxKpeywCItAo2mCv5yVCa2tLbxtSNxxuziR
Q5TPuAwcCDY/aCrjyCQIiz2Sc8URcNe1CLiOMuxC+zdHjk7BJLsVJAKcC5fX
DdM0ymdoBFlryqz9EXDBS6caPw/q8nKWCd6icqovON9ELAFLT4zpuRQkOYVK
nku+4YN1HosAcwZgQxWFu8UWpyUqHFfDHnXChIZz9djY5doE9xWNbnAP/NaE
RvFKG+/mTFlQw7WSg1xAL2TkpVeMeA5mJxuO4thUgvMZltngK9lanXEHn9m0
IjFa9ehbYKQ3kscbnHJp5tbB1e/hfB1hdH7i4JIxqpSZ+AA40/CcQdxse261
AwGn7vMLlu7mnAoo1/ckyqF2EyqrVLD7dWECqnZJ7FEcEKh59y1ttdP87O8n
eAZwwas8DJNxlz8XuHjNVHj3iftcEl4h/U5SFFoj0ZmUoSxS4yYWaRjWwE81
fIU9X6WTZ2KOZWD7KPYpSRMxRaQWhwot6VuYf2yS1X8YZnBPGYI54jpIDoz5
nBzLCAtnIDOWHhYqbkMQXHR5aAWCMLkDCfPnlHGdnTQWEF2wBAceqZismfU5
0lcQM3ye/er8UbfJNY7rCC68ukLkiBY0c6Ae6yz0f4GVb+YZpa273dO/q1p0
1VL4BeBNhwQdfiUpSvCsu9RaJxkT0bPb+u/MypXSlU61cVA6RbvhsFTyMKxm
vS3wXqu7EQ3cSVVa0KtwqJN+ueGw3QtRAKJlilmkkwipDhwO5CHusqEuZg/o
eL4GjYD94LCvVWNlJH11a+DJjmw0wvNVopUiysL+tny7Wuadp9Eolsi/WzzH
BAz3xz+sHRVqQczf5ym3bzh2LOYGDodAI2vg3JLjc5aftMQW3/7Bwmqik5nb
lnnlJjjKhC9erdQFcEl53tc/vj1GjzH7DLJTa6G0hQ7x+OD/gkkZRESgv+r+
TKLoZGTsSEz57Xzc8lz6mbwtM4qF0zWsxUVcc1LMrkOvOu9isf0LbITujQMs
aKOuylODj11PAPoMXpkRfNGn+tNZAot5FGa/ce/ys3UFnZCXLg2sJSTK+EWf
l3iE8Dx9Tsbi0yeHUpc7Hw4G7UQQ1/KV6MTL9aoqodJvJd3bCvMoScaX+06T
XGWuZJ5MyeOySTeA3SmX4D7TUDMU9lS8UKp6RbAI5dxN1+ktG97v6xaGgbAo
XVx2kkqyoJ0RagNjkf9uBXYLo5fhEzzLJdLq5vyFhjlV6Wqv4+3P+VgINmL3
Id17G3gMEz4Rkwo8cTvgsvKGUqGDo1vZtQAknaqEpzxTgNVU1EHQkxPtYKHR
kf2E7g+ajO+2qRHHPl7SeaozqeBShthyJdoEONr/KN4Hvjq088L1L26rGri1
WjdOL6FAJkNIm6p9gpqVrc1m8bmiS26YHBmba+CVRDqA6aMU74lpSD/PC1aA
DCSTJDABYwEWBHlvfXGAjs2eFw6P+iLoeQaS2R54BDw7ufiuezlfJ2tNzUwv
kKc21pvy7sQ3QA22YRI8z6ojM1EiaYsroeH/6qqe1yAwCEdcLeIPor16HJ3h
U4svEBAwr3zjOLuw7JohS10Q9V/S84jx7NaPaLaOV8K+mF8Ph/hSmqsUSNG/
I4REwej6pyWPDz16mECPaBvHm3dM3ExOhn9l88cw8Oaa62WSSjgdpTBTGXf9
BIAbe9PQCdhUKpaXou7mQMJ8jTvEaeBDFH6iaB/8F99TY5AaqmYiJhSjK/Oh
sowUmndJ12ldSzJzc8+dhl/xA0wab4DyDCaEeHgPRkzuXwXgwCUBdfqD/w1S
hBHpBqCDR4aUOn8uu2o108zQMur/WqeUvX9THamPjrkYUBeExn7ZzE+SJK5V
8SXAfXfsX4mR9D5ZfVXU6Vxq/sYHxrtao/rt1YrYNOcgeqneLsFYYUdb8HGG
vdTprwuBYOeT4uXFSQWDO/F3RZC29KhM8GMitKoBXPbnNSG2AVX4wXzRWuhp
Anej8bt2UuLmHFUtdoOkT3xpupuyKHKEH6+r6XzJTCP4fFByQLlaBw9BA8sL
r6UerAIWCpzKHCpWTblw/zoiId/pHwKfPkE0oiw50BM0KM84R5Gma5LioWwt
zgfOfPQMjIvW/Y/BLRxkrOdOG7zaG2WXPzjBHLdEX8L43GWSoDeFPhkwJDf8
UqgiHUALLJkVX3UoMdm/H9FjPeFOW+wtFECh49mM0mIGl3gTcguneachiBEL
fbUOqavK96ryrz6hGdpag9LD9INki3maOanw+kVxN3cHSnoaslbUf0dJ2S6p
JitWV9pMZJKbITjLYAuvQzucFvoc+5UX09ClDYjPXno1qv1B5G8bH6S99PHA
QJRchNgUGcTv5auGnqzokdZbRASQiRKagWKM0FAS+ZcOkXT1fa5WwDBkJDZG
uUuFK9ja8FopvDz7G5GYhYyxZKRmRqoQRDbA5f8RF84eUq8xRcmne+sBFkgX
kzv8o7OGLiifajRcOHHR6b6kCGtzYLpWk2bpOihR2b/jkGWvljtNmQVr9EAG
kHHmW8FifHsNENzU8PARlBOzIDOWyNoV01bdTIyywonvH3DRs6+TsY0CxGgL
b9jCmW2f9o81K4Ke6UnECSLiD/nJbYvdAiRxVj3s8bMJkQoO6O70HYfIiRVu
eGKMO5eDDyV+jo3reRY2skUAjz2Zj+04TAIDT17VDNRIi2v9uJwgZi2h8mLa
wY36GqPG2CVdnh6KDloJ8PdD/kZbRQB8HajdiBliPXPDaBq44XZIv+OcDbkp
ey/+VNrs9VxTbwcf614Xf019NTbLmY047QuqO8cQoBzbPqIfnd7DrJGYdkyf
JPJ3rxyDnsyYW5HkXCXaxNr8NoPjkhDihtM0mQunKnhQG6Yyd9Jk0A+sTik6
ypB1b5zNG2Ke3toBdDf8XEiPeouTxkOnDErRy6YCZ4yBHvHz+vDig0IdqWPt
fKPcWQP1pRpfMMGFCU+KnWQOXET8qkcB5uUs2vZSQKmmY5P+5iD0PeFcVzpK
ahWB+CSrTfO9yXutuR5cX1QEFTeeYu4Gaha0xI7F0+4Hc0bltecObBuC6zyn
bJ7mvAw85ocvHJCZpQ8iYcD54TwNgVB7BphG07j/DEyEpZ6ciqEavDazH2hA
d/TgOiN2c/BrgwIWX97c+/xp0L5bmLGUDlG296BLTz3Rykap8CH8KOS7zfmF
z/nfaNPYh46X2Pw/VV5v5wZ1Wfwijcq8h/ajBhNe4dkC6c6XMtPoWHNxTOJT
ijJsmFEuUUCg2FxccW1FGFTHNcadPszlywEX3QEIt4XTjZcsRCLofbrWhzHE
At8MU+Mnx6/YcOCL6gSEaJc7u9xZOaTfFj3TFYiqYhCmkcBUYx3+CmOIHvs3
zPCkV7eIFhwfcYdcDqO/Q3gABO8N1lYI5RzY+WFl7fZo5u2CgYD3kPaLp0QX
jc7wSpPqSk5t/0BftCqoYk7FmWjxZ/Di5m0gHml/0sHrMTMmuJgzL2BhZwzA
F2dWikO1RsPvUo/mfvxZ/yw8IYSFnR+e0O+JCQFmLlHZ0ayZqHkn+CezLf2v
OUZ1BND5oGJ7CDW1ytFXxFWs2JjMOm7nuZkB3H3s35PxO9PVCFrnbemAio64
bgpNy1cjHb6aNZW9bdycB2Zgzsmux36equDCjjPbIL48CzFQgzl3yTWtcPZe
Od4X3fISnzne7mOutg1anSqNXWLFaG8CqAx5yR0jJHCzd0UwEP0VCMuF1wcQ
XDOeiAMnUOU0D8tOpo4fgNyZdoPV5t777rDR4rLCIDA/QosJ6FRPCJO7PpKq
HVb9o5VT7e0bUfvy1r0nbeHIZZbnf0anUbwSBbhfpRNvxtuzajO9DXIpKGy4
/0A1YQxXzbAAopDyhUtpCCGNtwSIIu8sUYYHrF0KoelAhkGjEOpGq5XdefPT
/UboeBptz2CpY79FzRbraMIxFeJi/JrnFOYVVXfMjLgACzg7KkRhBpLeekQb
zpAg9xaSLkdD8pB3N08c4xvxQM+hUMg5I4R4iweIkx9bpUrtpbpNJuv9snco
0D0KTQSojGUg/Pp2pKPyhpA+E6ObhFUv/btve/l2E8Ubn6DJn2yrQY0dSveY
tbkeD1u3VkEPYAGXIlHGudDhXYpzS1GjLD1qCXGZL7k2Yyi2bBQcYbVXKhph
ODy6OLCAwXtnZ6TZX/Gpq6iXZBVjOy7z/8dEaGy2bIFGMimUaLxqSkSO4Feu
pwAM66kgArVtuGNCbVaUZtkCwbkftwSFZrBhvcsNnJeaehg6HqGTYZSxqMmP
fi3CMxbWcI2o3KyZgjo00aA08NJw692DC09x8RHHQsmuE+zpIM0h26It2vTn
ZXD3aA0+6Pt52mtSxHff7f3vm3s6t6+GGQ09x16pfsjYsuQRxMcJi6i1PlEl
s29NAXnLyw+29Iy7PHwZKKj1WOTgcD5BYb3mbX/JcDXBctZ/U3Kyuub8ofDz
kE0/Gi9YdzYjitSNik5RGK8R8EgjPxlELAe6pc6wUy1OZJb2lbUR9qbZlVwo
zA4P0QVVioBmIEo29FUAh0l5BhyjFIevlKQz4HQhpUAmzRVZ1WgvltBLcDFz
B1/FvVQg5semIXjqX1p/Q7wUFgQigwvTD3BrHCFz85F7rdBGpFgLeN+eafir
0xq0i6uq9+rg6NUX5TOiKEusZ0aP5vDf4NwemV7SvhQ3LsvmijhbvCTFznlg
srjqvrDbu0iBmowC0pLviVap4OyTTcxgfmOrIkfBjlJwBRv6C6g05bjMDCNO
mm9+eRNPB3i8asz/o4OnlAosWxaeZEO9nA5T13G2tBXwJPQrGquAQ/QrBrdy
H4HiA9QIKIl15uvCHsFGI1+2qD0FQnCheW5UYcc9KayQm5lWTNPf89CAPpaH
XgE+u1nDvddKXMA3mCWLyO7DAGM6VOUluCF5rwOtcuOjYdzOarHtQpXZMQdg
m5a1eSAgmq8Ah+4Hkd2ps+cvLk3toOBJGzHnD53CWPueODGWXY0U7Wx+EBEf
EAs9Sg+oCm2eI7fxj3mmIgx8KSXTA3+Rjg+BP31b/Sn50N82cNaHgcIua2Ed
cjoGftd8xtTcmK9i5wcf/RsT1PkVDazHW81NIJcXuoJ1l8twO9nhuzUcoJgM
JSqYR3MLur1LsE7x/Qu4Ra9Aq/WNEyygu+ZoTykRYg1JoE9X83lO0bIceQXZ
dLfpT+DJsX4joZoE4W0aiUqdpRwitaoe1AKHrfqMgYDsAj5iOtLUPFZB+kBe
lVjX4Py9AxVJON6PeI9ypVwP3tj/ppFsisyRvUUH2cf2g2cHyAU/nOniluEj
X7nzWOJEA1fy8ttKvXuI3Yoo41DhQvsGn1k0AfZLf5Vcl0k4mo6DvpxYRRlZ
uA6KWTz9tkGR//4YvVx5o56EFtpkKe5hVgx4Ek1N66hodf3wx+9Z13lgrNCo
PU0uIlI4zskGfDK2sWISmF4Ej5JzOvkQCJNbYLKVo2X2lUEcvxdfUNMei6bM
jtm8p6iTciL1evjPsD5wX0jBq+AuzCSgkSJYrcnPPqUeBkp4YFnhkyM9mKA1
5ZzTIHK4HiqEc5cQRdLurZE3oBXtnSNCtIP6VgXjvuhXrEX5ZLKyD+YTfGzH
h3NNWhumNiv0LV+odZ19bKMe0FxvYavp5WT+wJEbFlepxvmjyoyatr3U88K6
BuYc/5vZQsSjyxCJe+Dux4Lt6WelvA6ejpLiyw2EGO+p/3QA8tTnA2abSvFX
UjONHE3nCl6bZBTk2HxMWokNpIwbZlHJ/JQmtUQ+h8VeNcPclD4K/0pMz+2f
D0IjreextrF16+Uo5vG0r9N/NWbjm9Zq25xPQyBQmkWCEHWlrLuVrXmZtRZJ
qOrXx22V6GQycLUPYJ8qvSFkpxJR+xJMqUJLAr6P3YU3pkWzOWgpbcRxDGOB
dDwsAwapgA1cDz/50hMlphalOrOOV9TvCH8URal3mvv8oqyva7VDuRwbkQSX
ScOx2pnJR8da5Y0cljor3ZkqGUDAbZ1VhxcIu+mWXj3TLcLWefnUN/0ECwMv
vI30NrL6ePXX3x4XHBbStNaQ9/IkqxVZ4qENIFSOqAQ2Vjcjwrmi4vpdoo5j
L1vPNa1L/9UjN5WA9B1yDsLkaDYvbrWGiNkJdEGw6rPEefGnQLatX1fihjZa
TKWl3t3aVSo5zM2HuGugqZM0mx4ab0kyjNmWGls0dqnuEEP5/iiFonEvzDRw
/vU6CqoAESmQhQVSX8r2Tf4thdGrwcwiWwwVr7JN+0MmnqiMtv8eRmAGL+oG
1zgnqa61thnkCvKXw92gTwtURvSl6hP06jmNtoUjkAPJQzFPhYAc3ea6EIYc
wTxtboWpfaD6zoBbPdTY7dhFnJr+uxV5JRqguLFIWbNQMcpcl0wrAOx8X8Sk
ljIGOdcSgw4PAEeB8Pz6GCvfH11dwIMQ6PYGcplEBUsrXXaDA/HiUOcj6Z/o
jpUVIQZ6Sq4KGHAnPEtpnGI4pOS0vEvx0dptU3VFS5LNWKDqvvHdegGwCfPU
+DbTLERdDafWRt/DX2QlLr570P3EOV0IPI7W35uHLVm1/BdHn2jT56kXOe6Q
aV0f0D0xZTVRKJeeXnJnAMkcKKk2fbx+cykC3+bHOthsn5wchnJRKW8KjYaW
599lPduBeDMJPsB+ZXSSBYKE1jpHc91/Mxsf7UavaOMDQApvg14jKHBk/t0W
S4Xw6gY9smjAPHgetLmrqlRbH1au9oXjrnsiXv27uyRFXzRmu9gI4JHsD1nr
JUpnukhRY5aB5IULWZHZcihnWyysSpp7R+NFuaetlK2DuoxSJVK7CJY02AaS
EqSNswwEv0eNvH2V8/p0xaip/pNl7R9614iSun/zgiW1vjmyU0FFDFKWgSxl
XI0YkCPaXt1b//ID4kiBMmGK6LU+JpvJaCmou6UMRaz62eR8Xh3NWfwErB+d
aToPzJ41fZAyQRAqZg2OFTdq1PiKkF0USFEcl7lKzfVuQv49zey4d7AYYPwC
QYMtykVIvgt28lbMWlKXSl11Te2OPLtsWl6x/DPonC8PQD3bLFKK7cSaroqx
6PH3mGChR3kWO0N0vcQMlV1B03p4WC85I/gPQiBVEsrWgd+7wS+RBfe1XyBV
S9MR+EwXdcnMODxMhlzXPRsNet7fxtRBNsDv+KNcveImnYKgMeUvg/N8A5s4
j1WE9OqTjWxAQxpEs4I17FOp/RFde1Z7y7EbbTWah0qznXDBCuLAivjckqB7
ZmfP32Y3jyw2x3rCTPDFlu9JvQ8mt04SsIP94tDnLQVbXckXQBOh25Oar2WZ
AaNwZWQZy/GjJFuxNmjzWkZK6rqt15qGshJPdTRIcgkCScVBXLDcFi9NXy3O
55eo/NcsaZYPTuac/WTBzs1EMx+F0Ww7lFpTu42BS2X7FPNCuPqacxJ/aBtX
3ji8IgGA6jqky3GDTwqh0X2gQxbyfpYEXHZ1gjSQ+149nibWAx3IOG+sVZtn
ayWmEEp+aBbp+ufwLLHQKzaZQyY8Nu9Zvi01I92kp9GhjWcDf1V+sFFRiPDi
ze/Wcp9Xe5TWYBL/n64Z37gL4hFulraFfLXtFj3w8cfLjd3DjseepcZAYKKm
iiJQW6lrNI+QqUKxuy/iE8UV0QOWU7SpmtlSyVtxNtss2gcGA25XUkRdOKy3
VgE1lR2NSGMbH8xRR7zST1Yr4MvoIYE6m9hqcAOUHKssaTSpX9+EGY7U/mQF
BEQrpBZUWr38lAJxND4hFHfByQ+TjKBzZeGz2rCnQ3JVoVo8n6gvSHZNmqOe
1YcEH98crh4daGkhzozHghlcTmzQhWdJNis2Wi6xW2OFimCtstntwfjmtSpX
OAviqPnl/m0MQLacmhHo5B94qCn0o3lOjMM2CW2QE0Lz2fFYQHd/C1Kdrn4m
uOS8RTFIam8iUuoWfw9jY3fXKLTSEpeVECpMJeteHW+tmeCNq69Yf4YBtbKl
7lQoCZY6vIeuMs1fXTv/cD6P0mdcq6GkSF1vnuglFGpcnY0T+wZF8EL33urP
OA+C0isDsyPidgdwrU3O/1e8XqX8XGEvxG6Y3fSsCK6WAcSLTZbQnGOLhPXq
38+PcKb2Nhjhrjzefa2gTuRheZboTmIVzoFPCP/NM5ugm31McMX2Z7Lnz54h
e9xIhct/naHPfrVkYg7Po/buYwNVVYVKTQWFqI5mzF2JnSei/iASZsfqOKPU
L/LMBDrfmi3kDJUk7NT3UV2KRkcxdISfYLyhTP06rmQLFJoVhXPYg2IG8vDY
XwBt5LeynuEzcOayKi+7/tUbPbJaUWe+EWqzR5Tgn1fprbBt1BoTOfZnl8C7
I1jcj+gHXr4sTlp0Sc8gi+3dW5sV2Is6XxBZ8Pz9cTXxbpUeSPLTk3YX2Ux+
flDKBpmYGjsOdVH9a14sISR6y/eSYv+IbbhwLZPLAU310mYl5b3uiHgQC4eV
G89z7IUXNo8KLgtRnG9lTwqA3PwSk87fmbxaS9j6zP1dhsgnRT0lTWBuiUSP
xyXJiPqivH+X/DXT+ZrIq0vOG2Fq9Y82pCY8tb6McML2YbhGyO9bCsXWtx9f
SIzPiqUt65p4B9bA5QYlpZMQ5uepy8GAtIPRip93ZJuQMNTkptHu1S/shMs/
I926+50YhDxWmH8lv6rpChXIL7Svd/ILrw8pMgnGMMLG6C0YFMGDjtqz0Jpm
3dbwPbzW0au25Rc73sdpAWF1Rgwvyki+QgNzzCX2BO8CKU0ju0mrdtaIWRFp
vae57VyOWcVqV4clz8mqKKJMDULMDFaNHNXIApYMwviKhnjKT3Tde0OuEG+q
fUcv6pRUVUfhKNRKoq/uVhNyu7dBnt+EOZavBKc5HMVMy8VzzxHD1WNZwEH9
6weG6bbNlpYyeHOW55CrFG+2o1Uk/e6z8x1l+1tkczythNSQk/whbuDDos8W
1LRT5zcZwxRy4MUjHBbCRVg47mpQT5Rv1XuiGR4VSEBU+1AEJXrQUMuOKjOU
iOfIshkug5cxKyJ4Xe0Rp35PTRKIKdnlLFEWsSZJoKC4ZoULRt8m7UtOZF0g
eGvznIDLhuQ18A+DizXfB7rrN1NHRUgq4QuLphXizNo7yHZwi0k77dXb1ian
OEsvAcxCVdoQM+wVJZzbVc+b1/5Tq2bJQA/9HVXZ4+ceI2I8FNUt0A0OBylQ
ox8ay6uqrF/Cb6cmXRZfHSe6sCo8k2e3VSbSLwKJJaDJsvVvgHLabc4eQGKq
yUbltocnEOB5B+x7W2uQq9HkSXp/zhZWpqmAX+91ylc0YfLxWVSkQhKu25DV
sYlsu1LmPaBrnc3qSz8AgtydSePd4c2cSZZ1/cCCgTcdSBcOeAq30MOYdt5b
Wb9OsBPHD2iRWc72NeW2S2Q6l+xbVX9MgZX1dClwIMNtnUMxiaWrKMZJGFBZ
IYvBqKUiipV8QmRUeHEIfyVBvBEXSmupoDrWX/GVpzdb9iofs+CJUmVUqNBb
ZcOXaIrRrAUN9clK+zcFRunOEcRSKW4NKH0dOl+vTTw1QO5ow+8rIgPY53OI
jIwbLUGTkGF7Is1ggCFUJ5FX26/U7DfbT10OcORsiFbUjZbM31oXNQmrTXWj
60PeUlis3EBVg7bbipEDeJp15e5RKeJIsKjL8El5dMwXeZ1upXUVkLdtdFYO
Q7LWGynJN+yy2YGTNA7L6kJhBw08oCe7CXLT+11W4Tlxf8aooUPYG5rzgJI1
pfeou2Ma39/IEv53e9W18tbaLvyRZrxPD9BqWkWYHOOXDlvlyTX5cuclzdn4
CCmhhept4nUjDwL+VamxcXWhlyeQbe3gmmcmyYvurr0rkmf/smDu5vnulwVh
sU5usfxtKjVPoNTon3BIfNa//TaIKE+g8GfRnEr4ArKPou02wszpLWaYeICm
F6AA9hPWaQ7IISBm5tqzur0V4KW0Iqb2DmAzvV7Wb2CBq5oVJnvfcssbhuP3
1uU9SAvcboKfucBRhYWMHOIyzXfEjbD0/6fQj6Mu4oS2C3PhpeJkYI5NhSTd
yZTunJJ2SIm7J1K3W7HY/I87p2yh/GGBSrlQSqhTpod2EZeKs3uflqIEmKu8
p6L8GOjqZV3EpF9JiXeOGiN+/TzmV6ifL9/+Hq4iPGd5kep/HWi6ng0ys+GB
KgW12fxxg0TZAu98tmsXnCQR0uNxe2QFQ2S9glMGeUBBMhj1PgzaKAhycEVL
aSvplRoOz/vQCpjXSnQ3dkfpS3QAONRZHNWEcWTS9Y1SLATtp30yAQD3bf5h
MyE3aHXqZ8HZAFF0kBe2y2JfXXxapT3wnKfI/0Wnh35vlIhm0oqKwFXSW0eT
gXuqDrtG6Vqg/W17l11PPDTuDtWQMowmBqDPwSmq7DAI5AWUN8UlRAHbSGh6
3MKp30ygJUPITIHxVOqI8HU+MzIrV705xCB3XQc/GztAFborc+i3ezASPbUd
L4YH6hSxAQ8RAKBaa1VM8XQvPBhKz8itNue56BMexfKlnd2FpXs5yHfahqVB
UqNc463lUmFKYFDCCzvfO83nBJl45NafCSWBiTDFjDqBRMQ9oc+HJL3P3DLH
7JoBfNHppyJBYEZViOPuqpFEw3icl8ufQr8NVIh06nvY2GKcdLT0tC819oWm
HWgYZlce9gM6t82kacYjZpQ34uT1DlkEZPqUEi/wNfZofZZ2Lo9CnGN2/uqv
MTUFsHRHLzIWopJgtvXzFuqqcb+Gb3jVjsMT4IWpvkFPsj0VfMt7u/PAFU4a
818XI7y4u89YgX8a5PFwh7mh6FE9DZFzND+QaIhru/0FWWyKfI8ubpznSUk9
or/He/W3V8E+FhhB+9dmQ/dJD7QbrRgm1vqLzXg+ZqGmfVWftQ0rzUbodt8M
i33UoOLBAt+2+IAOYc0Ktuku1ANUOpYHGMl2rr8CANVTDgTHN+sX3QyZAX/e
ryuD45J6hQuVGRJQJV5sA+lBCgIKLlGxENasusfI2+lLFVT58tPd7rOd1OXN
im9aDKnCjBDHN/Qdg9vQ9cKDQBc/qwCEqk4TkVJVK5hfILqFtcnRTeyscZ1F
h9MZoNkf1exyzcTCTwI17c6deFWqhgu/SLjb1G43kCgqDnYOQFUA+01wJSIW
3seiO/jge2EQ2FHtDiC4ttBrEhOg2+LfrJnqaHmtShzKFM0YBA7L9APQVGjM
91T/eWk1v8vY190ibesOiDYueN1xqJrPl7/ooz26z7t6b/ZKrPqf6XH+2RAH
MJVDi+NGCNCVvrxgXiqvxqgIm8dIeVdj4GCQ3QBODyCow+AZPwW6kO1sZSiR
sVt0TNkNTdw5xRJVLC17qN3BznFfdEZW0xdp3AAq8QI5D5LnkoNtw2crasuL
fOURGJkGyy/0yfptJNIm/9Edd6Kr/BfRvEdxfFqr9lR7Q3F676a46zhH6MLv
bIPr+4ktzFGUS76rjgg8EdrodJdvIOZPcVZvF3teqLOVmcUPcE2Tk1vgMx2I
FQWDI/gXqnW3J9zJjIegfXkXqCCtuz9jRiAy3FE5ZToLiB9VaNg6f7Bj8uCq
OoMfzNLij87W+iAwNkJoubeTlAv63meNvHKdhcCMUaa2dobyUHV6InLb05h2
NUzFKOaY4IoVm6DlXMwzwGShT+MzRK9vpLhSdXJaRFN7+iSgSsRe369g0GqD
mQ732Hm15BNQzLgef8kJakr4o7eC1uc+Y8EAhqcXC6Pme/tVtOI2Krz5aVeG
invl6y36fuOOI6KsJLWnnsQUu1AHqvBxG/IK2ZI5HiWP4iDKhl25DoH9G8CJ
pBoWDSfnjLmOChs3PU+odx8Nr1LZNCbX26+9RIa6LaLdnj84ZQ1/Bim3LFmj
npMNB9xvYJCUDDOVCY+F4ingHEK/hUnAWXG2mXL4NdcDlWZyo/YVov0aa/jo
/RFUQ2tx/WP6w4Elda+N6DLkglusyd2UXgMeKOnSrZ5YWfVnoqIJ98OhCqF/
uHiWtsrVDSEokZUs1a7IzYa5+w511PQCxwIpTyvdcBqc5jQ29BG0g5aNrGbt
InmCdPKpa1pAccXwBvvqyZeoXR3HA0FTJnW6dyC5us7XaCzNqmfBQGsiWqun
p9EmLAfh/cEGm6wamWpD5R3o1QPfCda/4CSr6wMgwop6MHqRFmx6Dosai9Bo
fq34A9WyVYWcUjS1MwCkK17kujO2r4zvoEIpGCxz44LTFdgSFS9E5RtXwxRQ
yPpVFTdA/KXkgnD93ut8nGaMuSJ9vgNGVFLiA+1fMraCgtGvf9BOnelt2jF/
Up3o2i4it41V4luRSy6VoUp4Zh/fxRBTFsR7tLvky7wveNXFF136G29Bhjcv
SHJXzZPMbkXt93MADKFbbf0aua1XTMQthF/UQ2+mnVB9MrWJaQMejHefAyql
DNcg9bDFMu1xvNTTT3Ctw9yG5N1DK5nKB1ykAxfjjXB9ZJyfx5reikIn4Njq
Q0ys3vJf3TOsdGCmahKFYKDoKaMRGFMbV4kM2+q1GrXoKNXMY6pDsDeNqedr
CcbfqvCmcrabTaVmE5xYN+YVoi8DQmYq4kIbUPiCtMC8VlOKEl116kO6Uxd+
30Eryya6zG0/1EAZvKTatKJsHePrCUAK3pHQTPcbmDIzADmKp5Xb8uQ/HvW3
LF9oOQLYZ7tpWlIdQ8U3ALm/GUmW2rHNaliitxcqUVVBJS0jRzE6EQV06msT
5SKiy7nqKZ6G5Umrm4x6PdrBI7EAhS26ch3gY4MNB2/ADJSI07xfCbCGDLX/
1rqAuDBbsckfxKQNzA209ZuHCsRAltEPrmGL0Ipe0TuvZRhGZLfrxNiplOFA
pudidzISa3v8Pvge3/3ypmLr4s1XFMwosQaS1JsEktKuoKz4sCS07LET5zhp
Q25H7F9hlE0slo3+Hc1SeeFuJ88IiLKb98aezFt/kjtbPIPqvnM6lbKu+h6Q
kVWJsY2cIb714qJ0KT2y7dpMS00y1Dyr5rzsBl1jnJw3Pk6cGqHctrhnTyqV
nEOEam1gLW9xb9zuU5hRaTlmjqlZeV6uiJveAnDVxAoA+SoQ17SsYcsD6iIx
LPRMKceQwKL3RU7ErO13wd9JWFOWg4E5f9mCZqQGbkh39yfcMOx8/1gGiKu2
OGEZSkkq45OW3ZCn7+gwnGFyqO/YKC0PUxqLl8x7NT2NvSz3slCSZfptkUOr
95h5ZgIbfL6z27hnS2zdd+kR5pWpAmseXP236JHy3AP8ReAOs24w/jGrwWeV
tbFU/C5kK69W4GCDZNTTHodAVNtjD9RF2Bm18p7vkpjzzbiHnPHALWvHfq3X
40l0F1uDi/vt1qOh7RkMsR3LU6qpjNR9gYQL8HXsM2om6NkXybDWt5YtFeJQ
qOOwsi8jnFdHpq3pBQfBirAYiIGbPfyjdv2QdMRGfSrid81gtqPMw5Fyp5kd
Oh9+eVu3WOFUrQhrYfJGwuc/VCPbnfrZWi69uCLZb0bk9Hml02bO7ZfbadXD
Zw3B/meEhH076lKQhcuw9Xd1bgcCxzrMQ+nMkQiKDvCBKXsR2ysiUoauvds9
iyay3F1QISI7BrwCbRQBDM2rEFu/0RBIoP2noC22GpAT6pweRYQRaExcs2E9
3Qy1CoSY0yvFmPap02KQUKgPJFFdaGaXqyWMWHbRKTx4Su04efSpxKPwYpm1
bl0Be9cGvxL3aMD+QrFX/2Vwlqq0Ea7qyfaRwFOP6js95mQluc5in1ffDsrR
YKf/9eSuTbQRuEwRXGeun7JgfadaWVvrHaCmREOA9oUEV+dGhEpxO3/jFj4M
gUzDcuCjatdQ0wx8rFb+qN32wsSy0FqrRM2yaxj0cvEwlYYNyTYcGoBAFDw/
v7/A0FlIBbVl1rJvuVsBNSIYetLeSBrs1WPfwoGkckIZ+FSAny0mxE5idZUK
Asmblse32JDPdxJUskD3tGppXoWhBxKtk8vYwBDpwHIDJxsEP5cfXdyr7Tgt
99gWPdY8ie5bfc+pn1pcAJ4K3cfmMEYDEAsWskUSJQT0tPmzcsRZTAOf3i68
ZeMyvoWb7Ek4geGW7jl3ts7tcPbswRJN7gVERGo8HqG4cyhhJI0uJtRPX+2V
NeVjfaWCavPuRyGLJWkqie+lGW3Y84ZZz/ODsLAujnsrenCxS+3cPCqO7FMk
3kSd6+5oJEDatX/kWSfGmln3bOfdXtNPr2l5+AH2aYSdbUIZxcxXlqloQqrz
WXF+VoB+PygzWchZAxfytBLGB4uoFHlp0MJs827do3Vi6A6A/J23Pw75XcnM
ki0VqMoH8s6EuCxOphRhCmDe4k3yFZIBirazjLoR7FqYzI5NN91cno6QsjdJ
ThoI1dMR9f+xVeOmIAAcSlvizRRvu0ns6MN9OjuTfjiRVhe4k9lHxUT0ptCN
QKpN2zO+kTW3+el+nWp7I+biyqmsbWYbWofL1CxT22uZp6A3WBJa4TN/jQZL
n1KpCLffdKDBgy+9fdDphUYEpMtfZyweJNSQYRTrN815IhiDQK9imShuycFV
jWZ7m9NwcB0iEwKO4NXnEPXDiw5SKR7Ee+v65bPBTBQPRPHSGgLQJj5Jnf9j
ns/tCYlbLkJnZ9dhC4PxDjfR86p4Eo4/zlHzdMN9unFdGDbbYPy6NN3aHRI5
mfX0ZrFSnsaw3GG4dUvNUCT9f7M+CEVIex8psDng6ziPkfB+hBlHDTgsPoP3
xQ65UEkzbZNDSPsuMM9/GTFzUd10qCLkEb5E3laL7oovgGFgqDzG5HaVzhfa
tG4prFluv1Aag96KhZOjhLBRmdib7lCoT7IQB3EA72v7A++xnxrB6OX28DhR
srVtAyAAgJNmRy1jS+hvqo+AEMRALlzKkdi8IG9Y+pGOsOqiziuFpAG2dnia
1yVSuRCAsss+0oxs6V9X5sNsY5xOmYMlpFJrwitvVXzQJmNTPEuXHwGMJrKx
9R/scPdWBNIwYYy+CsoCySHbVtsgnAPod5vx2t8ETWa2RRZTaVUjTWDY0uMk
SAIsmI0HwdVcUjLFun1xctTr4e68Lp5wYaiv7Pbmn+q97YMv0Gdp78V8/Fj+
Hl5jgjdBSKyMoSB8TqWOoX6dYwK45q0E5e8q2SSLkFkLTH/MnGRN1lw4o7AH
0eWKQwHVvbxtNcl+BcIJoPwa7JxtPDM+uLNgq/rPgUv1wJFql3MYENRhQDbA
YUGWMcxHdU9p4sPVosJSkSXnjUShR3mgTZxb/ZdmjjKSoNGomQT5cB9bUBx0
yBNskQ3YZERRG52y++bRl0WrtZtRIWAZ5Urvg9HiS66P+MAPWXuood9osu0I
+JEMssBSVpoZ0kQHmuARLD4olyJwxw9CMImdPzW61bpg326iYV6JRil7zKMM
SDDXaJ+4M2JwHUOjZyVcNGCoD+I4E1e3tewmPRa0X4+O6drOC1nezGih4uOA
4URzRrFG8XiykJfwBCPJXzSpJWZLTd4+usaHc6MDetN1fsdGa568clxSw0dX
iHHkNMQtVhffk7jloA6fBiHwJR0pj1T6tSWVXiASFYfRj2XYAsXc/LmRIXbK
vq1FK1Oal5KJeaTg2COevh0TF5PXiCUN31WbzVZhaZyLs9wQjCLtUbj8r1a2
/cCjP5FEm+5BdEyVpd5JYoyhCEWZpcuBu+AyXlqIQLwM+4lhGL6NaxBZFwOi
PUekxFqGDdUVA+/jB6w7b0JQhZO1jx4EU8a7mwg1PH1XEWcsTiWJ+fm5zweb
WA/olFLPu3EsoniaTjAYVl97iBl5YuitT1rN5DhsGSGUWJF9DBFVqjBk1MIk
OTSsCakGN9kE/+3b5VhVW7LWd/AZ2Ip13mVkFYv2ruI9kLzO33gCLrmZHOri
4SGhOCQW75ZxWlWm2HW671ZQXdyfODD6zkbwEJc13sPJeAQjV8o/qr5m6mgJ
aWLZN5P2n9cZy/w4heLkgiIKqtinjP3zdPHDAj9ObfLR7cDUeu31EOjIPFiw
1hZr25VH+RJTtkoDYRSrzI614uXimF44Hegoj8f3GfIBCdPpBMfCFJ55UJvG
t3Q0UN6kBGsu5gBt5OaAIL0JnKgi/hgisnPD89BHWIKXI1aBdCXevl3T9UBm
d2lSEq7b7IcL2bdYOayPSucxFN+h90nFL64jZU2ZcXYxqVMuj+9eSobXZfU7
svV3FHq0LTsTvUvdLrvfymgiiVIMJSxke68ejBJe3Yry2HByaFgJiAqQh5aq
kR3YFqL45A4K3L14F9Ax4bzXEjU1Yu9tUWbxd4KK+FwMWnbgSSQ2cqNFbQ9e
Wwbg0ABMULm9LftKsrr7Uc78yMao3zmhl0b9ixmJee25A6Broj1O3gZ5f0Id
87dprOkfzUpz4+P99soIep6nts30UDsYoI0O2vEVpKmDEK8wkzcfZW/dIE8U
HaybK7x1usxnjym0LhQ+Zgh0KY92qs6hWEu0Xt4y/aZzPvjAJxst4zna5aoJ
ZbAzeZVgxsxb+UGRFCEFp+gPgcVcWdxWA+8NOpmG1YD7zSgsZeTbBnf90P2F
TqYlKLKtdI0PPpmB68bsUa92Y2O94lv6sec9h+UY16qD3oba/Kl3h2eoGBlC
LszjdQ7WyAfhcnKcUGK+WFt2EdtnZsQFvaCw74nXWHJynfbLiVnONG6thj8X
ekC+o7hFNKwzErgwAxh8lXNbX2qXAac9pVw/DOCdiNCVn4LLuQUSJFXUOJRD
6WAY2XjyNmxipfDlr1Scm3MHubrrD5rfR6nXnm1pR6k44qiQlMZBmYqdhLgX
wwlRfvPl407MKi+DVl3tocRe1uqwvUBgix16SJBqEi0FFoukJnXWG7lUuulu
TuXYFklnGzoZ8D0vPWNvQl8uQkzXHYXR5kTnzmrvQu9UNJJR/yo5KXKEYrWw
jOr54MCFtPFa9paxu2Jwei1MfdqpWULNaTgsVWXDpr0d1Z+Khb8y/9H94uFy
xTl0V7QoW1FuB0tQ4uO4y7GRn19dAWqFIrZmdG5g6bAkPkTlOHhoDf7h1MB2
m0/quttRGhrFFg4ZGFBboxfBtbqT30PK9FcAzKAneRTA0xu5O9CMGAZkygRI
/hyaL3RXqEbdSWrpLi6evgf9uIrrjrpPAKTmuYNMXhFyCz9ONIIZM9NxIkBc
xl3HYR3bssnP2IgFWZ1yaFCabahFruDpGkBN7r1fxGhiBx9CVVIuflx0CZja
sDI2cbs0ODuLzo5NOZaaymARJ2XxW1CB7iZYhZCgW+KvRRDGTkE89zNEcWh+
w8HC0MqjEWrP5i7Y2TAwXgNVpup3RpOqlEw4KpcKRDjS2FEcULYqO1RW2H+S
c01U4UtdK4bAe7BmoRWxY+jLUSbeCNWK3BzA1YYe7UwqVcVEKFdLsL/hrNGO
cKnYhT99DW2SgyQUx73E0YvnGG7NKwfVSCye6iI4rZfFgThuhNR/KAgMJQId
6+mqPesFbMQHlknKGsKMEESOFF9qO3sIIgaLE9FoeSxcBfs7IXBoHa3IMJ3z
8UpRTved3mU7DKH8/si+jYmDRj28wwjU2A9KNy6HK/TASfmiEqY31i2Iwozv
BMDLhsIiRi4MNNe366V7fYMgaljjPIxruBprSYXtgDKI/GyvipoM7gu/zx3q
RgoIjkKeZVVBqnnlHWbKi8kcXsp8/sYwiuwYG/U3zt2AR/niBWIxUYrOljHn
zp+/zZQgxJXuvscTfOM5dpDA5ZeXnv1Y/ZU5qEAegG2mO5RXbjQVMjwmhBeA
XUjOgMfGGo+GA4BBvlX3S5trnlVzV8zwJPsq0jTIYZytLTIeEwemYupoy19K
dX1h5KfQ4tFoq9YzE9EvdgWt3wjsJyKqSht50C38AsFAIZUyZTntuIxJ8HoY
szy32LCSrzHwfaY6WSZFa7GJeDJi8KMqFIKaYoL2B53TgpU0+5CX+tGm4G94
BgvEGIMxhKcZR075wuLhm61qXHpQ+/1CBDKe0lD20WjwgiuHin37JZyaj1xe
BHDEgLm9a6tfbhd+qZK9y2Z/951gYhPOQSLRPwP6uqwz8GwUKfliJO11mZNP
RyQfYLmS5ik1+kkRc1T/VsBBhCtQNs9essFYpC1TQUl6Cv8FaCvEhkc53Z2Q
32I6x2NdTNTE6ARNA+qw+NNDxpHIaAvxtHxG45TbYO+3JZU2YxT45VxxrznQ
E9KOHIpsIL9utuBdjsycUPupVkCTQs2VL8Dlqjl/5HL9qpzAS1lPjmYwE13D
vy1fc96ma8iCLB4fZfG+fuFqNY+KvbQl/PZcc4cSme8N4nmwJuzeY4G01P9h
bfrAyqrORkBnwK2e1wXhBT6f1y6u0gVw7PgP/Y5nbdfCXRpA55oeDRDKTDZP
RQsaEZGiyJ432I+I47TatMHDO+wMNX6iLA54SyjdQgLKZyx8cEL86Pe8dAmm
dcW+jGex5NEfYzqW1jMDeWY+kI0sggBTMmhjgUCzbFyhbfPoIbe9Hh2FEex3
7Oamiw2efeZvj6IWTj8o+S749Hjq7sJAf68tjUCP/eafqJ1xj7y63VFq/1MW
sQma27qv/ydDsBhjP2gDxhKGwEezKsr4QDkEVkNgGYjdWl0OxdLdCFKF0J7+
isDQ0ONEEHzg2GFY+KMG8gPK71TkNDukHMH89s/67nD1kXCsFfT4QAd/+ym6
oXD9n5m8nCvh1cvkk3JUa8w/ijNC5Sc+e8pk425+VQuO8T4fqnLh/JVZHZLB
r9fttw6jZN0M0GzqHFWZajTd6K/D6v3qqOzTrE8DGMExVd36VyaC/RA97H0d
r+tZMi3VfyVFihEqS/Y8+WhcGtDkkC8lgmVbFOkSuEhHfune76PM0hSXe6JK
h9AycY4BJA3UVGpL4KgrAghhEP6m3IlNlWAPWWmmgymSC4ZAtLej0UzXmwlN
ilkyIWlGbazSsBGgF1ksel0HYgvZPCMXgAvEf07m/G60YcHvwt8cBwu4xDSn
WNOIpZajNECaTuF04f70FaYwIsm5lHOsuOtuvgoiBODZx4Sclfz+OCgiBA7T
+gPQGBZcjH+BChauuHZAlP3FRTu5IJA+p55r3yselIszdNB+E/0VMu2BJlif
1ipipk5tNN5/Rx57d5WEeQ1qk4XgCEqZtWHZHe05tzshPNoGPwFoPjvzyya4
bVlB/dlBvOY8ZYp/ZBdhXSTUrxIrNRY4X01HTTpipROa5yjZ6CSUJ3FfjjDW
0hR/jM76co4qqrUT1jXz4jTHSJcWJ4GkmAWcAhbQ3LwW2eGADGFzfF3FqDJn
7CLIo8WbgPMbqOFKM4cLYLvlj+0P9NiAh2vqeTwZ31RQTJCQpTsPx+/cN6EY
FNMOG10GVxp+WLmUNkW41hu/R79tZO+dMTvYYazPrZgxeWb2JUPT/7LGSbbU
ExBAeQFrdCnFHrMZ+Bhv/GBu1iFOuUUDMOWtwkXlr+Snwp6+2OPZzd4rMyyV
+9TgfceMBZ+MLNhbPhJa3vdrxZUjGT+tz+oP2+k//2WdO7YxPF1Hj5SHeL5B
ATcyPxvatwnL/mHfd9ZQ5lTKtCapZsIsDvGqizZE1CLQglQ1TJKN7GYBOa63
7uMfQ02KdDDwaH23bwuUoGB9NYbaO/EB0nhl1zd7We/0Fy/RvZNCb8dKdMjL
4r9I7f14QYDrCIeJadIPM3t5HUUSvd0PSXOxiMJLJmFXSg4Q09sOIprs1v3E
4aheCGyOeIBvDkgBoJrbUjzs/6Ly3mHYQIPoeuU+J7uDP2ZPqaajFN3oSE4q
IqyRIOD6lZs3/g5syHpCYLiQ3WMG7wiBx2YRume5t1J4XKFKoImd2pizf7Gx
NNC9ZSCpxpKbnspJq5AEEDmg50Z0KXVnj68/Vg9bNuKg+evTbTdRsULQG/Io
nxoIqm+nPlfe6/giGqKsRbd5WO5cYfGYfEpaD5wDGOr8hGW0CIgnc+MhVjVK
jGTISKl+VnC2d6u9xZf3Y7TKnInaufCSKDbclhyeOxPPXBAcnc3skcUDIYS5
b66oH1b6HX4WJyDzKtbhUjNIp+8IvGvxts2MeCsWK4Mwj0DAYH6wGU8GeSgd
Ur3v7naE/SXyLiSulOUfRhChKRmdlYOMEDroJGNB2q/Kc0ZpQuiBnINUN/8h
feSbvVVtFeyjGQr7sOOVwg+K7ViYR9YfO8GG0+ryRQ+fkeoMHLu2+w0Rs2Ks
bhpxVpFA4ghZzuXQTuuuFdRHu/zLH6rWacUpI2SYtBCfLGumHqxeRfaIkWb4
8Zmqs2z9icvuuCZGW3GXXx/9+TAlD7KQpenecXnM1LvLzT8Sm3dk/R+ahvl6
ur8avQxt7/5rLTDTdpVkR63vBeZ7c/wvHUvFA8E+5/Q4K4uIj0zTtwdoyHNV
uld8I4ZN6ta/Vn2s/bJaKDdSvhZ08wverQ8U6sJ3k+k+CVfdZCINa2lH8vIt
SFzWwrVrRqbMED1nXdQIcZnzQ5QNb3qFFXIWYv0wGNbw9VB2PXe9B/cIPDE3
SvAlCjJsVAoMpNVjB9rfC2opeVvZFHN/2H3sEMS2dlnjXav8SNrngP6RFPAV
2iNCag0J4633cdC1Q0znXUFMu9XiaMZAXSaMIcPbNMlwsonWSxEAMVo25Grb
BqT+4hgh9XUseuNU6DbphuBEsjScIE8VdhpqY3Z3Ua6KD5MarOo3MCJfpIFT
ebVbSkAnUgSqmNFoYF1GpqfaMJMVSXBGljxQ+qnETCmw00zgvUoGqVY9pMMu
YqA5ZQka8gXZfywAaTCaH/EfnrPcsbHKrIelJsQJs8JyiukiQn3OsCXI0nRr
kNESPOJNXbwRsl5KGuQcoLYvznu0Ik4wsrmj0pzhh8sRv2eBY1tmHv788rKg
O1Nlev53SIkHLNgjxchavick6NhF/juUfb2lWEsp+lQ6+2mzOZ4RDREGy7jb
pCJycu+AcMMUquIQ+yGC5Lu9NelsxSFRdXN8D8m+YN1tSLi19HRonU03fA2I
P3/Mo3n4+mmP+Ho2IGhggKqWAcjh4Gav6+iNO/rEgbf4wNUMPE5a6i0qH+ua
Cmm3NRHHwo/W3BC+IGyv9uw2Dyb0tlvFeMzTEBa/j+N2m+jkukhcvWng4hfM
g9ZDhgQ9DzncB++wSZrHCIn3onRC6Us5u+24BhCKMyuEk6KZ6I1HaooZTSey
vNapOlDhdNUxOTz0J9JiDYNq2b3lPaGJ8jZBz9CXaEDDS45oI1zhwyvAomr0
omRCjppNGUYK7QZjwecdFvH+zsFOnTFGeF6FRmAPJrSOTnP+s8i9w0LbEWqg
DGUKlVQN/qjagCSW40W7KD97D/nOnDG4DuPXhRHVQLIYI9K4grr2h16mZzQu
3Qu/zYttc6S9aDQ7tmpZlaZuMvmX2/f0ECSaa6yotMfWHHTce1Od4Zyf7bVh
h2+dzRcfOKH4GM2UqDag3PwztBsy9/ygDtTXSCqnQrjfmbYMMS1FmiHGgVB0
ZNd1ags16xa+sr8Bz9cMp5KLRiDw1np4ANgPb4m8ktw4HlM4u3J6tdCKMA9t
Kov94hfke9YtPHm6VZzSHy/BmsiLtIQji6WsK/CP+2Zf9F02jEuukq5nWvPC
SQygBoo8pc83u5r6tDDrnt8d4K+zWw5Eth8tfD5QOg2v+e7f1KS/yMS1m9FF
Ya4D6/xmzCsYUEWmqv/HvLnbV2NEHU9ztBdz7BrzyeFYKzMkx8hGIoLlwNQX
qQkUnHqPFEaibEPAuZzMJ/5s/I98VQFejGLaNRFdPHbQI4HsQJF/T6GRzLR7
a1HyZlDbnlUAzARHLbM+TFiu4rtoDNDCfdMcwEtiE3NEqEOBR5YXA4bd8vkk
DY+M8812DOzl/8AGUB3E2l79aTHjQ+hP/bz8MqdQFvAEFM/MJ/rVZnNPi505
jCsA4AD+/1nCiMDkdF1ioA5rib+qPdsbKBz/1VNnlgraqqDCv4VEqjewMSWb
EKFyI632ahHgnirNw+hMCz5Sz5DCdi2nmWXbO+FiPGKIprxCZwuebRlbiWXL
56SfrGoVHHpMO9mfhsjZWNX4lcImxvs9yXhzcunORtFKtU5YM11o/+/eGwI5
brJAlJ+xSo/t8HGwQsKdVTe3LklpGw89Da40ddaj9oYszsXbq8ufuDHkUnSx
BNrrBu31CkO+bAIxMMwj+Pg/+Q7WVXDCKsTQDNKsM82KiYqsuif39q0awu0/
SxvzsdkPhe7cBy6pryjLnSDHvJP+kDOUrtbvuzme07vA7RVi95DWX6uSYJYW
2ZaOR0wFbM9wxje4GogABg5Z0ncSOcDkpbsGLsrjmVFdo8LUKlEwsh/09rwm
pDB98mmbw5EudffVmroyEns0AnQgZa2Egu2952MB2NS0OYsE1ptUuqiYl+d6
6JvTzu1obscgi77SZI1HCrvoHE8KuMmwlpT1YV+SkuCsjVZYn5pIOtbpNgTN
UQGULShXB/UBUEB5GamIC33PqCoZuVTpK6w9Lkaag/H64QLbTWjRspMhY/ON
pmS6QCQc/J3WM3DV9v7s/Y8mcrtw10hm6VDJLPDFB40B/bHCpin1KUOoSZpR
B7go9fZ028WEA+HoDuv6yOyIp1zxICalA8ieyuO9i8ygnLFO/2k6pnhbT16/
KMWXW4kY4hSQeik36xWGZG9VmlKYK6mZvWaXnsCTJRmFD3DZa9BqOW+M2RZm
xPQdf4IpGnIN//xcObWQxO2E/c3BVrdPxeXudWMIszTBQqQColi3eesPuALN
M3BnpjvyUeZxdazG9UwhA3u2by8kKRjBsT8C2+hi2P3KWXThCVmZ22UOnhjQ
btVkCwOO5KSqw1XhgiUtPdwxBesLRlj3jIQoXQ9FFW+Sph8OlBcf9FcKJfSS
pGa6du+7w5LWxZXtQaUCnJrbPTSVpVVgfA+JAQXOFtTOPTPj8FpjY3GilhpY
O927J/yShIxWL3vQxA0qxBXRJz+chOzbzOfC8YtL7EQxsRBIBmeUyCoVbtq/
fNM/2bUJpuV8mbH7thYe2bBxQRIvQ5KVT4rhuI3U+IBUIVAVKuc291e6pGv3
+C5s80Eag24wOTerQaX4/jEiFu43xyrMVvdKTxXa2R2ydBsPD/El/xEK+4p9
P8p8hucVIesv5hzKuF3oRr/RoH7yrQUKf9Ak+Rf6Z+GT3c2cEstbYWTFIJpB
cXkQTPSgF6QxGGQJaDOJrHr59uTYFd8C9vcc2quDJ5dTY6M0m8sgDtMOySyI
FTaW/ndIHpT79VS2e13JOqWpgff3qYysalxJvmHKXDCA+Iln76+5tS737+25
osB1W4ioqu9I+yvzDtEq7CzbrxXmEnWPPiDqkuIFf6/o3srzTGeK4+UZIREt
6BAwvW2Fzu7DmBqfbNTBIefayV9x7ZG7O9vqq2bYhUzqWSupT6MXf6cgBFUj
6uMLMF1bTFIPM0QkS4u4NM1OXBnrENEj4XqEX3B0FbDEkLs72gLUSNmyLsTm
VGUZq7yFOUlIrE3bCuoyw/F/559PUcODkrGt9l0MODoBSyDuTfksTYS3biGH
7BqQ8K2PsoP8eVXck5r/VWjCYZloKWjcQnRNztIwWcGF6S7nzwVLTwvuMk6b
dsT7UMQSZ8GlEu9KgojNh8xJPXmlavsQIolISxY2RFP6/SH06yJKXjNB7AFq
TM7ZepkK2JaSer8B7DcJkR0/f5ruMFzocGsAcb+ktobL9Ek14Gkxd4hh+myN
vTGbifDAPqBTS2E6L6Hm59L04INlCPy+SoPJ2JevW81UV0NNfbNiflRTCqYf
lPGX739qsbONbdJAjlh3RQ/rtvv5kedoiOgVwW0gtAp4X038p8A0uK8COkQh
6RMYB5XhN+sKSgSLSOOMl/eyEJ9N/NBONCg789qYvD0nuBxRGIKmOo9lybiq
DYxvVHYzxp4jTrqZ0wm603dI60mnoXpZILl3XHF5ShPwUqbMcMZlcQ7j/CuV
SmW98vbA1w8SUqnRjDQUEKAOajj9bhLTBktL+gOkCc2Z9Zl0UUZ84ew7mh6h
EedsReT0o2eWG1n0pYYoHfIO2Y8yuMV+lLsMzUZSk76wQRINXefLZFtFo1lb
cEL1gca1pOcIkkUjxpcmDDOJxvQJiFpfIRaALQexx7nxziVM5yfh+jMfWr5C
nC0r0byU8N/Cii9pKqIfL28gaLeNFOanio1v5eHha53a/2E1kgFYHDJ8RE61
VU4Q6OOYTHnvUdmDQDXaBJpKOTc1XOWb9Q1aAwMN1CQjZmtRd0YtlDEMligg
dBYzXcFioWpt7Ud5aaEdZx3vYNH3DwS2CHmoqYrEyvz2LePOVyPPnxLXKSBb
mcRTyIPyoS4+w1GduFA7kdGpaYl8u9ZLWCkbhniI33ZsoZkRb+Bj5cvvDb5e
LXfsMSb4qjkuaCQg3bAjiy+yZUjNKHdHkDTI39oTVuHCbYaRUFxP5PTdGCyI
SH+2Mx71NCZhjRsgP0sEDL0ZV4RnHSvydVo5tqXcydWITvHFES/2d7zUFaY6
D/tC3h4xTW2j923lSYBTExWEFpKEUldtTxVhlRVReA97WsT85z6UNi555/as
forpqKtkEcObQDJusYnOT06g8eC+BUZBPHdapodL1m18r0UF5hJenzzSwUjd
x48k73T9aEeMjhit15ftRw8fW16+WaS8uaZM6MMu73V0nvwtXOYXMIsEOpQ7
9v95NTRYof/hh6+yZ4wRUZjqES+rBCzdDvoyzA7en1hWg1b4DS7Sqt8oMqjG
FiYDhQ/aGNrjA0y0aZeWH/29lbqeT5W3z3muqOje4jtKftWznbJzCrCuL7Ck
yvgZP0K4U4oEjNb/VcCvRPdL1OSywVQydWRlGHSmvmnWG3RKQR1ZljArgpWP
t8BKdBWTIP6fAJl5D7KppZ2Ne3ql9mcg4UxbTNidhin2/mWS15o7HTFQQR/8
38NdQmBxgyHrra66cgaBpXpvfe/JhAuW4/29JR12goWHhwfz5CZxv/uBW7tp
AFayn3+Opbc08TrBXo62UDm7MK5pUClNQUYlhmyqC61fq+NaKF7sNQn9sWjI
sh02hvLwYV948GoJVrLGtRJTJ7uu/Xo3AZAMJPTSZJB2SiptLLjHZqi56pJq
wAjHLqJLfL3b4PRetO5SB1a+9cvTsQgySJoOcsJ/xbUzX33PQj50fuQEtja6
Ko6ziuGt3lloUuwS+LrvbGbOIxCWXd/3Wxm+Byt+FSpOCwx6N7wEc78oWgfL
q1A1p0dw25/4AvKtonAJlAA8TVZZxBlmIuNbghAw9cYIt5ffHrRIjeBbI7k0
vSrFsbpKBGGrNOT3Yg/XTI4rU4Dam4oraYWUGtPe7HqcL+oTYhA41zDuFKth
/OsSjY6K8O4WV1EvyjXd39JInx6VXPhdKWZUnl2TtGMXmraEjFDp5OW7Nbqt
Zq2EgSjBgbjwnG9Gw5B5RtWTGnH5q+fdcugYk9OY9Vn0cYiHueiKdWsnxoOA
+NlFjUf95POeSkcwGoNVQuKbUJ0Xc2FZb/VGpUN3iZjtWLbD40vGqwa37A/L
gkS16m/xjlZglAC/6VDTsVxqqeXzHCAvHfCFTUI1aWZRYMBZQCDS0N3BP3UU
D+ZOpk+rT2JuEekJkwdvJZaf7bi3kVvXXRDtQOXq90j11VOv5v2ZomYNyriW
L+STxYDVSh6ZV29tgutFelGVCVElgtKF1qE5KO2cp49O/AQBPNpZigyj5ApK
dAn7mubs7axMMtUqoe0cOS7hLZMfAxsBMsWWNEPdMBp9j6Jwq4v6er2ruhcM
/rMXIUn/Y1+XpuDDGuMpFlpuTImVgStZrqo+sB+xt1R7NQ5aDwwsFYQ834tU
aZyVBDpBYpTRRQkCDnvM8AhCCxqClS155tJ8amTw3jvkY5Aoec7RovOe3ZBe
cJUQzcwGm2MneZdgG7lX9IuN+3cvG0PzaBEh8v9e5E2OeA9HLEvoRZsOlRVV
8dCx9K03iDvly/41Q3ExS+ikLOWriOvk8wp7a1In7IxnnScIA1zBquKbXjGF
VkYYIdoB98cFqipvdWC9wjrmN6iR8nDd9IYJ2NgDgPkB5itxsnbOpj799smX
ZM3FP0ntFYFJOd/nqdl7zsy1x/JB+8mzZ3lJ6kG7QZsX+0Q5v6z7ht6D4Dfn
U5UMI66fkmTasXn5YZQeewjYUeFKPlfEzDWrIQAtbsX9m1BukKQR6XAPDfya
e21KhQ1RDDw+iy1gGRm5mRyUcGn+RmQWokc/sTLt78JWwozVYtMUxufSm7VV
gKaAE9hnyHHIQrQRvp3mo+myeKfrP2rVAGd2N84wLSJQARupo9OkahyDmNvu
dos0t/SpN26Jn5bxqQZo6fWWfcy2Os9Hyp1bhHT6+2pwm0F+3+7oUR+VbDOa
uUTmLy3xDiiY+KsCys+m8gogKOGsPn2wp7FWrrQ4TgSTmgZ/Evwr3d+90jRy
VQl7S8iGZyevrgw1LdPqxAT3M+s/JfsohbzO47lJRpUqGQrEWbUAEs/yS4e0
zmgBmh6ak+iPXHaVBiIw0m4HHBh3ieo7gk64waFDWRdH7oeyPJHHXF7QvUnS
mxReEzNNDoFT8ex1ZJaxUnkmgt7jeuCQ2CrCloCvz6M7L1Qg5tUq+47BtDZ7
Ageau0tuJDX3s7KLnpLfws4FGpDvtUMTHoAtcoyGUruC5ldJxoJY8LdVoa/x
CKLJ5djBbe3Q2JSHFPAFcLQ+cWIhn3xOUs6dPsNrJ8B729W1z2F1BPwVmRPV
9MyMlE23ep5sGLiV7jwpTqL9uygprY0rOEOAol1SjEvsI8MTDIahcdgLrdou
8YL9fewup6O8KYKnk/DZGeUURWip6h3yOTh4P2fx81Bwd3GVfY2UEjNyE2S6
5sfBdRA42IA2vruyzr5Ml6lCIJcThppbp1jOt/ZEG1U1RdChSBjE7OHpzOhK
bWNgrY9UFxBkcPrSZ+PvVDWgbm35W+ZZdpSm4uxIuh58JWNjGwRAbE392ICh
2/ZSBXvj+kkgbyJ7JRErXKPTFwPBRo8h71U9Dv+ohBdDtUjIssNehqfnjxfc
s2LWbIMomzHSg3UysmApwQFkYm3UqLNbzAS8JizEIXI8YQmblqF1O/yB0Swx
VewdNcODaskkANv0LvxClXPnoN79tswaa3Od6X+slQp0r1ytd9PFfXtAiUwp
oPsM0tL6fmsXhfPwosQMwbKjMbgdNKKfSTsIumbGmvsrDyTlyWxnVWnXEPwV
8Ka1IFVzAALnqy9FdSfm5H8OHV+UzFpHhWLEBuPUjfE6fkaUXItzHeQAN5pV
AtomnXfyjvx1fiR1q/1852k8pzKNqbTIifaLtmrPc+eEhjOW6SoYtRk1BiUG
8AQMO8+Rfhouo7DWx4msA7TyKID2x1dph08LqcpvcZk6JN1m6KK2LzqEU/pM
CxAGIHYCvZb6hzwOkD2RmN3TwBLTUP30RdSHbG87rRphhQYmPAOgo1Yty6nN
4j07gMJgOhVM4zgcA8iOEX3GGVHTFHewwSZ8REbWVeYXabR+s8nZpiQ+PoUA
6k4RCi3JGnj5V876Nh5rt2BMzvvpqERA+fN4ypy2H6SglRoNwxwDjU+vIsAF
EepyqEMg2DrCgUOfWLuhTJR2ZVDvZLT/q66W4lNkAn0rDZ1YqjvPNTFyJS4N
1tz3U/h2lQNdIn3Ls7cjVNV2l+Vv1mVUlz9hoQTzsUbcfJkIseruN83HlYCO
N5e9wBnns/JKlJ1iot7KdPao5u5D0zNIapC7guU8LojY94vEpAY1Y/dKCYG1
ZfLX4la3WxY0KtehSc7cQnhKbi0Ab1PKNrpJJdLsi8FjzkaQU+cukhkal4aB
0mRoFVer2Dthj8Nnk6KjAmdZ9cehM9P47uW11pfP8JjMJyhAnxppYY3lHUGs
T+nOAU8GhrSLiY0wEHE/TFyf9vDwLTi+YsY/6Y4VnCMHNMTc1QfoPm9HOCcV
Dsswe08yDBH7bGFjIU3eXP9d3V1mDSj93ci5rPwZIJUncBSudBSI07NH56VQ
DH45i9Es2215s17ronfxIKVEjRKCZFMmW1ZDbQjDxoHzdHm8vo8C60Etx0GN
MGzP6N694g9vyKHA9ttfyI2+6Pm6c/OVU6JgWwoBIYDt8nDOh3TBKY+MHV8N
0bBu+4ueUuzeRGCG72BZc18MmdCkvmzcz4lggWxSoK1Vqo/m1S3twThtO8oz
SJwVCkCzL6OFwuF0LXMiNL7tRpXWu3n31RaznrEIkr81JKYQaQsmYMDR4Tay
tSN4BdFCMwtT1AMg11hNQgaqaf0HaDiDhYXnC/fMWGsL2x1nSbwQ1dZD1QTL
0cHKOv2H5Vijg4qFkEciVE0O/NDPSJ5LxHDfKwpzq7AeMoHOHBqbw9r2ylgZ
pB7fy0IqVm+VEC4SwVFAfRXNO8jojAfi+v/w9qwQM+VRk2huvGFFxJHo/ak+
b4KMYE9/9gFQf3ldlIN04OxE+a35hfjOJodnHPEUqQWozbxzXuwAiupWg7Sf
hzCm0fMydvqWGxNVEhWxg1f2Pe8YlsSQG4lV2A4/Tk92kkPkx4F5ukkMRzY1
MD0IxSnMSV9DQky3aXJ4P2rbMTqI696+6EdzZoA29VQbN9r5I4zuZFNVkbJc
toTefcpzQVGx6OBolVNDJCsCSxDvK4/rn2kvJCD+7gucfaFxc0TXPc9NQMGD
oXomqLIKGztfkZ5m3hYIzQd43heNhb9REhv1Ji3RRGeYuvNxRYVb3EsICm4z
XgjJV7A0iRqd5CAjkOIsBYonkfBsoBC9mY58XeEHZwFCIaFknvSFHm1RhUlR
YBYq7qmQLbad4AsV7w6Df3tTsqUG9jbxzN27MbGAczkcAdgKg/Vb5W9WwGDD
6q1XH2xftkcbBPV8vRTjNK9w62uL7ZxI+XjGrX6EFaUXvLEMvNJI3bRa+iS3
hwTdvb13oxI7bGdFrgrj76G1izC6RSWxXoK4tQQaVTtQl8aQTGrioiSpzPZh
OJIpqLXq0prYGxF6uHh9FqSigi+FCeQ/tA+lurAvWbuqD6LGgj3wbMAwhaFn
Hms/3/BNSTHIoZa7ZeI1I9qUXmBPiddRkTxAQCpNmMnN/hzQLTTJ6GnCKEMv
TU+jgT+Sao5FXWby2VYzr/6upTPm6HpkUd0aNHJwyXGoaunhjdat956A2eEt
7rVi0kkha90/8l3ryNDCx1FuUYNguAoYrgL+RCTIBxVu33qX4glf4XW3YLCF
uRuUGwKejenksHRxEhyxQPJsk21sMHjj/EDza3YhF3idmo8B7J9113sOdpdg
qvnsBup6P0uxguzvYeT4YYntI1Kg12ivQNPblxOo46ojrr41H+XfOY7p1kyd
0StX2vxQctPSkVfl4bNQrSbuhgH8S83UCOtw5mydau7p2DrSAaMmpnW4rBjc
7E8FOnpHLFwLNBdd3pwGLvAljKMfcTpDW5+fhPnZkKXmAZyU0eUeVD6sSHE3
7XkEujNaQsYJFCGD5va5eQ4uq4dqGzpWQRRqmrmmlr2KLwybj9j44GorX3Tg
UJDF/beKZ76Vd3/5ytKit78UCfcE/0VwyIVwM1OWhUh75EqP6i6EyZYF5jCc
7opxKQLtjGO9fkzmetSDcumCezw1HR8kern8E0vyZeO4vvxWFOwklSQA5OAc
MRBYnGSFUQuTeHYB/8x/g0GaN/WYzNvVERAnOgi7OiHKXa81EyiOmgKOixHL
/FjcYD+53UVV6dCbk3t09W+9Lfle/tKemQG8cTokLoYpsb1fLVV1eHJv4lzF
yK6uFdRO3UCcvGa/2OB/TxwHQpy7LBlwAuKF7muLs5zlZXjD5k8JikTRlffN
l6ZuSUtzZcXf9SL80tsi6SJzz1Agym1lVPaHPfzaEdMOheEd2748hfhT2wtN
8a/zHssNFdnMuh7YZiJQiTqKqiWJsN3vayCC4+8NDYAyqeiBLMMT4uwuxtDE
k8wpo3HmP6e2b+tS7bZtHO1zR41VViUKcrUcF78whCcYEiiZvTx7KZNRqP2o
88xKGFom6zjZlyynIADjPcBqdjsIeSSGdw3UGqPQJlTGr7/w0C9wmu78HlBC
NRXuoRejRKmLcY1Yd7D7qTR8zdAWwuQFo+Eipn/Fwg7ZtPeY1DnWiAkL5x4Q
Lcer+gnPSSPm1+xK7TKjrNkY4oFEWsoaer3hoggsLDh6Z1OHrdQi33V8rdAl
AfvaFiR9s/0KtiCtwvP2JRrf6jh0KkG5g4f4zehHIqISqvW1L11UgxYBoykw
myCShdm1vCZG64VL7AP90R9WkaJi2pmYdKfhv5WeB7SAbXtM3iE/UEb9UYTF
IUl9s2EzSeu/G9puiemaR1mj76zkbi2I9FG5kxo1eEDJG9RqHtFLNMhIelzT
Q8h+qny9hA5DadUDpiuvWYsX9iII6gG7srJIMXtDwUw1BBCj1um2BHyC/nHZ
g+Nqf5Tgo0IoMQhxxo9BEJPX6BARvxp4Nhp8xP408yeGcLU3w/dqoJ/nY3G5
7FIyyVtGGMp5KEI56Gz4YAUeqXUnHqQHR1iL6eOJkdF0iXb8ZjNH2ZIilFIW
msWCKrvECav5B1kXtmw9pc8gTSr/fA/FylYlLHW6p6U13Iu9lJ1bL5AZhPqp
nQvClaEjNyeZTNcUJP4fTDdo9qvbsdqOErMQoyF05Om66KtlHlfAaPrlA+c5
Xhu7tFL8uIrfotD4gcXQJq6ZDDivW8P88FkOV+xeEZyZfHTOBK103ubAETcZ
q66lMHKMTI15tX9toAQDpQ6uoLCh58/iBC4Oqh7ld3Y56SX352+5NO/pvmRD
UJAleTYAdnQetH3ncV7+fXdGigodEfLYINZluTemWi6yrkVjZHrHE1JYQwv1
HVa2srRCcjg5IREARNtraLrJKcPynVHt2jWfJblCM948wS52cfHrwmbghXWt
+rNhV7t6GqRUH9w1VhOLtuYg7arQMkPxllpBdS9VSZteqRjmamMzLkbsj7wx
By5IIfpVI0e2weaN06w3dFzDEMg76rhbtkpxoLV8jay4MU5psq5mouSU9Nu3
h35jCvRMa/+vN/4B7UGBnDSX41FMH6SXooQpEI5YqA4AsqWlA02yhfc+rEtm
9uw5rcEJI799PZryDfyUd5/TR5r9NBdaUtlHaaoeSOpuLb5Z3N6XA9YrqIEB
l6PqMJlzvr3jAvgZvkwmWSn+h3Z/Kt1ZKcwdmhtO5AEBYU/t24tdI5cLHJoS
v8OnMpsJraD9/6jfVKkTXKCJPCczaUwjNvdTN4hNIKVLabwdvih3K4eU6Try
PSq9TB416wHCdLfWeQwsYFSaFTxpBaKjdAQbFOJygGROq+uYkwNIb5F/yGsi
IL9CkVz4BQkLt8cMGFsWKzUGbzlXWEOuh5V8ZKjR+BC6NUEuhFI/3QEAmLvB
ZmJHn4gilFzNFabLlwxaBY5zLob2+taV2OCTqt1QTTmdX94aPO7C5Pavgycr
hMBgIYS4V/yYlaAnodCpzro+X0rmHl/2GdZgIaW61hZigkZkutOKq+xm6ZPt
iiKDDBnXOkZomv1GzCV1x4WyB7PS8yeG54suKPSQSkrFhvieAlQYdseUy38h
sRKbRcGukApyuswgld2xX+Ex9bg8YGOaYNF1Oipt8cnDN3MRWh59ptQjL7ZT
JdDQ+9TRIxab29OIQzkcCKkfeHALw7Uz+CGtmwu1h72i25F4MihwNkaQZR1E
tLmKZereU/dVJMkjno9hLIwBPejGjLvVfFxIlka4BjUbZjf3NApgBBcbV22O
KEEzIU53BkEKTdPNMoUu0/Vu6tU2rvl0XOUM2HSGyaXweUrI16cAdl2efDlB
IDY+xAcFKRlA/vLm/UeMyni8M+bBTZhxjfU+kO5PD72t9HkaN8wahu0dXUhs
lKdlhg8jsMk5tj7OA5YQqQN65DjiAWGv+fsBTElwpALOtA0v5a4B09dBp6Cj
8HZO0dWZ7vB02sOvVXlouJLOZbq6wTXuUnqDtLmMZNYtzHW6xZYzhSycn6FF
OXSifgMG3yemqHWK2zfGM5rD3KCkQYufGIp0+LxWO7PlaNjmaOvyrMg+nVMX
X1xEEecHLlMQ19Wc3eTCGNzcWcP86vjcc67ndIUsWn3yaJUr8YSnqWFB88Ge
Ee9ce+KURZEWJFm+NgZuxm/Nt2pVwj8mNMU7W0nrEAfGIzapKa6trUlxkSMT
8DdvjVFjVVHe+ERp+ky0xwYvR9IhcNjVnoOSZGUJhtegiRHQk1xAM/89ijgw
x+dGySh6gkndtOMt7AsKFx7geTWJvX2ljGkJZgFdyE6pALTbeO7myJy4MzDC
x6HANpx/6SYug7lxK7K9hj924VhfHTZvdLB0mDPPyr/jSUaj5LlwHkIlRBj2
ggbwi8vGxwA4SwObTOWjdsCzGtDw0KRrr4DSkUAdgDCLQc26AcUPuj9I+MXE
k4DVU2xtmn3HnhiQ95YUzJoWwC0GwX54rRVOq8xmfm+t5mmSCIb59gWRU6Vy
8erbCILO0oukii6HMb8ArZBozBcPBjV3a30BYHZ3ZFSA50zXM3zGqxcLTVwI
ISVo3AvJliaDZkkaj0gti6ZV3zuSN4p3UwwsSv0MGLRfjoSAD6EYU2i74Xw+
vQQH+spFvH7dUuUXqn29sDCXdq10emRHBzTC5LDkAHGZvNDJJ23dN72d8unL
MOrDEmeD+qd+JUoKUKnvXcTuoCxljar54P+skOCeSR+Wu33WmVY9hYdc6Srs
mcA1S0pBik6oq9ru2gD3IntDWpG/2GoDkMuf7hXMRQ9oeVoy0cRLoY6dZWNC
EzYm9Xm7LsrBy27V4BCojUd/EpidVOHYxzlbFNKCQB5C4wXUxnT510NclEbj
wM0pIj3fgwVvhOArg1PC6fWdURQyioi+fNiCzllIPM9BOCm6vWFkjwp23kGJ
rVa1DBrWhCNPzsq6HnFpLNV9uAL8EQsZxxgCRaUNYYnojFr7zX/Q2M/DiYrC
9xnWZ+zAek52Mfjw5EsHF4tH79/P3cj+MvRmK+HC6h/ZlKqMfmT04ZVLMqUA
pG/te3rezXVMqnr22CwxbdHfvHFEY7ao1wWsvp/2d6hnltUUji/760HuXh6m
AY1Rhaz8ohje04JWHtmnO96n7lkVeLllpsyUcvgIiLtTRRPEguM79LgawUMQ
1UswUG/w/EdgzOVAflXDcZHfkeJItdaHWKevSc7jqk3BNSP3hdQLuFtkUtUR
+5iH1TByWv/fJgd1KdVYDT1Iae60CvLFnbaXtc1G3Z6GAN0NUhE4An6hDYNQ
GZi3zLaFRkyGfOSGWDGKFlV24AuunSecv1FsPmXuXW5jQOJA+fEQmoFa61Ye
rCVI2rb2HKJ2jt0H6Q6K5W+23mBJl2bYp1G8dmDlipagn02/xG3FlNb+Ansu
zFEzDnV5frvfKf1ywMVW4RRYCq6yIfRDs7MITSBSQlykaOeFeKg88ZjOyKOY
1cDa3iclL+7Un3UpZOEdXydkCAeBBgBQmxDh+pjAfDb8hiwervk3yuoZmWiX
1W5410HlxhQ5yCk6sRx0qOCM4MQ7F1Z/uWCnYZZTzk68C2s6xFvyclWYsHr/
+js9IbzV24r45uodDlltAmB84gphFkj9cxCvFCVBUYEhOfOHovCzBL0wSmka
UFwi3PCQyeWUt6rIDVW9rg0tsX38Ev9ycJ25WfO/O38OK9C5gZyPd2UGCbFF
H7se5tQicY9F6V7CJqIw3583VtRdT46PBctknTPoRpr+SOVHganFKkA0a7pW
uLmc3FoyWpRDWdN4CKIzbSuCujlp/E6vBcO2s60Uz6jHHC4ly6eh5uB/fR/j
sjgW2T6jTmOYTpuMmuo8eozhdAVHqsoV/X1NS4dMQUNNBEJA8mFFMubL7f/3
sRtd3KUMRAFTwnzQEjwqjGNtGG+/GXnMXiHE5ut8QwsqM4g8PYFpM0qfDkgL
mdi020COKVEC3jp+X/t2QFgJ38gJy50mgCKGsDHTmdlyUEqfsojm9ajGmE0J
hacwE2ELKHSyHGYky2rd3ndyOYe1HIpYyezueEzFfiYB4JvcpNk85OIKxX/z
CLMOqwDkoHpyqPG9F5KXBYkVNopPe/TCUOIKrqJbgiFa3Q18TdcYyhvjInrD
i+rcsDulnihdh8ZVLkfcSU6mziyuC5VxYgG0UAVahSkf1pUmBgr1s/21bcFm
F3ZBFxEHcDQLHwehgZNkcDw7duW5rGWiO/noDB7H+AHNY+C3bft3nTiAcyvb
VjLVcsM5P90WNn/+NxF/qZJzaDYfBC7CBuU8J9cNAZpSpZnVBzdLL660HlU0
0XM0TOwbfAGPptKish21G6JZlNIpV0+Hk9NtqejVfuJBpxYXtRV4U9bN2xgZ
lr2wFfALxyp24jeLAotKd/TCzOZ6XJWTDy1su8plcML5wmuBYW+hFhJOiISp
VNLic0/YdyCvQlXrRij6oCDLs+/tncvvxdDgb+wJadqP4OBK6ykLhH4nD7RO
aJyHzo7YEUne6+kf1fdpUOPx2mMoXK9CBGvFHbUDvctOsZkKOnV37/z5uzI1
3bHAIEwfTPXl7+CpN6H1ruqFcm7XsZCLKkyMZh9Wv+TzJaaU52K9ZzDqrKbA
53LfAIIYi+oXA0kz7hOLNeABzNzfBh6+JtJjM/wQFoVsQxL1+EXEXHUM3EJf
6pCE+02qM1jNv+mJPGsMCDLQwZgdzsGZ9q3DXUY+bhsjOxnVTvZYsPmldp53
iQRv+JwhbkVs1J+CjVrx2sTlWTJT2Y8a7p9PKgrjPodNHAXUy4q366GuYP+x
U1g07iwOb+BeD06+MEDVqcVaDtfSCRrqPmif39jd+WzwHbSnK6NZb1ATRD/J
m+0L8/Lv+gquDGhjRlaXMGigcnoBw5EH+/VZmmgFsXAzRQgN9VR/qN3DYxSk
pzV36LVGFGSVhMfuJUFiFKjNjpGv1PTw8kq+nZDkZZH6EKdsAjGpwr/7taCq
yghpVcbfLB6cs+X+B3XCoGJpasQnorh2XV2eAURCkAE23k8gL8GxpQJg8OWJ
3jFreBKN2BwX4IpL/aFeUDjxcheUa74TWwarzzHD3UGpq8UWfLbnouTrETdM
h46dH6YHVdrWFluiLbr0xFd9bbrbRkrTvrabtRw2kgD6mJ2Z2kGZcUs3IcOc
CRrDeKNKGt26jL6UZtBg76ZKl2xnQi6i5laYawvysyZM/vdEPLtYegvmjfl7
/kX90jZLCqDG9pz5o/1kQQ8ZAFNdj6AClTN1tMandd9RtzSEGLSM+7I0Zlut
AG7em4vDiqm+o8t4RPIEJpoSFN5njlgJmgM4l5dZch/q2CaYPntRFyviTYSY
RCOnShHC0yTk+0icEK9g5W7nB9FUDZvUCzvvkxWkdevvXR5RN9OSwhOeeO91
/s+fOeQ3cz6PQQAwZCZFwZdjZnFy+SrHBkmbsFpowlI/vwwbLFa8XQeYGUHL
PHaoTWMJ0vLAIP6OmtBFkrs6Q8WEikwNpXtQi2MLFtZGR6fUb0sV6K64v1nk
JlgeMV4Pag4JEpddyL/pcfT/npZHJ1B5i9q800HhjSG00ABWFHFyUVkfu0Pd
rJr5gYD5qaunpnwD2+FAFMqHQrG9oLJY6FEUmPjjCHpCrz5tSImWBQEPO2Zk
iwvIzmFiF0nj00LAikEEbLmoigGVjdQ/OOtqAQbJiKcapKVYv0Iozu0yamoi
zcCwFCznkXMfDrUVK5CYkQ06tXWF1S/Oxbc9U59ukOR2J7phoMsFINpnHkFz
LpsZphWdroOAQlh2uSlY7fetf8UuXKiT5raxQULngfD/q6k7nVMcL1IAmOik
+K3abrAn9MtiX2/f4fFM9/E+rMEVvAWFc2ZFq2oqOhPeEezGgJE1WRmCKumS
D/vUIYzCV0CaceqtgJKqubq9v4fyEy6Pd9xzwUf5iEiKknsXUtKLefz3vaLh
uv4/t64wbppgsxpWxtoAFXe4M9fzFsm9CY7Gfx/ke1XuvaHcCIskROP5ubvY
AYVSqUXk9RRzpwqD7qRC4lbjCc0T6SE34sDrAatN8vKV+7ilzkCPvNdzOeIK
F0iGuL8AZCcUameuvtt4a0kF2ocKrT5+cTWcU76IeI/zUmc1odCIdwxdxUs4
psRBQMakQtk95VIMeWRoDItEy6PVR6hx90vngZDZpYoqoQVh+45AqZpPno5F
CkwiRsu6qmi4Wz8q/G2EjjEuwxzZFi62dP1zoQ+S9FqgGvx9koJU7JYfBxoN
dqRousEJ2JDmEnbdQwI1da2wlTf5vgYv5gGtrNYXi8QYJsqzKCGgzgpDuSot
g8TdK6by3Uonapv2wpF9BvActvElTbmawuC/9EZAsof3XtMupxGKQPaZ1Bav
LtNWbOCtv7OrkIZsjJMcl+jUb0BOGRieTFrI6AT17HDed7a/AMXvJGKJ4ICX
okAmeX5kKovkjOlEiLEJ7E5eMHiIQDJCdbnVWxNzWYhY+JiN6eUjHsUZitZE
XqhXOrO6/oxA3qqLL1SXZ74sQatQq5QQOCRvYsysskDS1R3dK1V2ZuhIPlQP
23SZEvSmVrooOv8GOke1ngtqdocs/QGg1w2tXDtz8/2k0S971CUqx1FxhSkD
2TmBB0KW3cFrX9rRJc+AYo2w5DnNUCajm6EtiIBW/DCLhG/yfXKAedKeb382
G3JlCGikzGrF1/x98Vu0i0OZFAquoVPQ3dvq9UBp2PCmf52Um9ZMp4IG5Oc5
50wi7erqtwWhy2RDHjLTch6qdNULlxixRPmJ2O3TMykSFu6HFDNaZ3R6mKgt
z0Gvz/fNxNhRuvKrz5XOB7NMbc6YztzLJ6WYzyMaUU992+/wZ7J1Om7LesRL
mgWDq+vHkd9MmPlaiKvIEI6Pf0gopEqbN64iHl+nx9Yme6/AjcEVT+nPICmh
nLaivth5cBGy3cQ0Rg8AjFOsNLWbelRLJc/Div2Bb0YWcDFOD8pMBvC+fE/8
nXc/lO/0eHcpSIqswV22nik3ELIvzy9o/uzKVYyjhko4mbZbjgqyeIhMhWgv
9SCZ68dYK1itArOEGi8Rt9aCPfQdFNvl5xD54D6UxxPgjdKsrsGkh43nkJ29
+Fj1LhBfRIMCb06II6EuM/EXs2a8qMEBGon6Ji0/Cw3xb/jVPe+aiJJSIs6T
2g1C1cLPBbZM3hklVFCONgnjYAeWlJ6OZwkZ1ydpAQ+osJZFGONRueroax6b
5jVOhw7xP7O+trmUbs56OOLvPq65Tgw23/aOFS1/IODFsi6yGwM8Z3U/zRc8
bTLAb7hUZfMH5mp0eS8tAGXpWhwLXxjOchn2SmrH1ripmHPRHU3CE4UtosGG
kVbDqoz2JImAl912cgUlg41c/wYkNDn0gbobziziL6RTbemIhHxoGJLgm5ZH
b5wNYbd2tLUN+VAFSRNIMDany/zZtY33X7Hja/4zTwV/JNga2sUhuDGPHkhN
mUyN0dSO7vxxXUjmvtdrKpdFJFes0Xn/+41n+UUgEkM7VvvOTIVBTqmirw4A
ZAiGc5DW3hiY0OLhSmtvhOpTML1f6kvjfd2vPRKuMvjdR0mNs63umXrLS+Ix
7hH3cfqaGRpY483iRRXlsS2xjORrskhL3A5F3zbGZsA6zVb/bI0chuSJwD6y
RZmpu+KKQkUpqB988Vfse4h2j3YUQEGWZIzmLhSWUfiaxvokEipsLNBSX3Vh
l4UOk+A4E+or6Zp3naY1jOKlC0uy4GeF3Vb/zqn/iawsLgSnqGT7zN1Fbw9c
G57qoHr54mC1sYOTyA9Y42tcc3TNzpxoUbDnHJJ++rFRc2dLjrKYPQ8X5v32
SIcVLX5JvuuiM6vxAskVsUQ6nrBoLkHnMbKUMysPXWgi9v33s0yCy7xc1BL/
eqtikpc16UAG8N01bWbOFChz6yzSVt+weM70bQYQQ7fg18Vbt7HQS3bBcUNH
RMADGLsIGgUVOZeATMDcnVOX9LRaogRO09FxzkSAMuIIUu4Yj06PHApkOcSK
nq0Ys2nHzW7SkSPNFNh+IaMx8696obUQidIvT3oACUiUCFJz5cp9zZGHXBS3
n60rmGTuUGklbcpN/Na1UD8dcG5OnlUcvfh6oB4xNry2+IMDFD2Rv9g86KRn
cnXJlUliSqOht1a5bND/uRKIqCMrQ9QaGfTIoWpRjFAMXZV5kuiO0ZDCEMSA
SAJ2PXhdWgb4l8QG7tgwv2OSBR5pgVEt7YxMYH1a/g7sT2HigoR3t4bk0WTV
yLcU2qYSWG5lC14rrEtlM+DxTadzha804HKCYlzG53Y93xZiYb5yp0KPTwyU
uJDOs6iwMWzotX+7xX9uJpA2+Fik/W/oQBA9UN8Xr6RAcmCNdxRTwZMMa9IX
1MPPEnlf64jR5vcU8JDmPmNcOLxBtHx9TnTOyjntxqFK/1PXmLV2bsIZEO80
S4URkrdAauzgdkTJSzPm63ZUgu+qBcGr/ekmJim0O6oWf8kX/WUVO6ap6Nnh
0INAj1NI2FuGQe7XOMJEXBZVA0xoRzA4WFSpip/Ddtls6qTuvfgkoaINTu5+
zJMIerA1aUZFfQU/H2CeCHg/lkfEPOJSD1VNWOnuAt6hi73UE7FN7p9p0wT3
RqffcrTKyolVxFyNEJWR51R70FQ+xkqhKNab51GlMyzONB61sSooOgR1z6Iy
vyKvg5CRBpTzna2d0w0OQpFdwXqfDxk8Abx1zgHUku593bmOWogO7uWmnvQH
hkEkSQc3XZLTAdlswVB/vfx7/hDrADLFoW2BjpFqhDvDcsWYFs67JhT9xTbQ
Cl/7TJXQXIi0yjzV6Oa7ERSAR7lgK2P95gksXtxklfNP0G5yC+9TdwHkp6QE
YytnIWVGeE1raHB2U4Ooo+Bs5LaPgFsIqm4JmptH8pVyRbONI8FkZtoebROt
IV51EgunAs5ldz/MEpH9dNkLFVfQYfp1OItL8TCdUnwgcohLb/SlWwEIoDgt
0kTngoWhHOkT+cQsnH1zF9T6cVBWD4vUF6gG3SZHJYcmgZR1DA5o1eG+sPsj
ThLl+Ag2v5oEUtfvUi/oIRO7sBU98UUGymVxAWuD6G+ln9Rl7T0MgjZEN2x0
YxZbwMnIRupNrVpPHxmt7x3e1xZkjBTLeIWQFE5+DehkP+vWf2AeHkNPNc7d
kOM70kMRyT3Fo4Ipsxg+5cVdJrEiQZKslBQqxoKXeCLiVBikCOiMBjXGt0vn
RjagYl08I1ShbskoS1E5FNCtm9KAi9ew03iYRCGQBp1YWiPIRBpqQCPLqTWf
0oHTx7vLgiDLAhHoUNh2U1vKQzwKf842QIOmoYFpamU4sXec6lkEsnyI6prh
avL15Tq8Hmr6qlKPOx0L3l2NPeeWZ44v/OEtNFq5tTJZmyYktbiZL6wbkA1m
NuhOx9P51ISMRZGliTo8oJWJdEx4y+63knj/HcUdk+ZRqSOET0gSEk0yMpLn
SejcysGc4syTnYmOkphkAZ3ETe9OfL+NWOu9eYDaTLMx4/1fvVgL+dC9SuVv
G9+yM3Ge3bs7ZyDxvUMsS5GFCnO0FJpEDC4446hmi58EwEUBYikeFKHWYpq1
f94xVqI4v8TNV4oezfRpsTeSIBfxrpJcfDhFIOvCmT8fxdQp+jLbHxE5DsBE
RLXPBqN64kBluwcRjmWWpX3Q/4hyEsBvNcnxJRu8YBWIXVgY9/RRXOhHVBht
QPwNaXzwxhXqjDLYlVPBp9lmFKEFAfJ3tgjrVQfSwgM6tlEVLlEHQ/pMi09P
3X2Ui573aBfaCxMmaEL95iPCT673CLF52IlkpI+Cjvlrfm6EJjWExYDQCAlD
rzusGkBhQ0Hb/DNfJiSsJnllO9/sKNsW2jLVIWdBCvE0Y4pZGMuP8rcHtT87
tt+u2Rr4dhiHKFKLAMkrdDUAtgS7fZWqvsvte30N/rb10ZS+M3nZkRs+xQlg
VVygu1fNu/xXVgT7o7l4vg156eBV+Eh6Zw64eY0oW79v9AnkShizlhT5W3Cr
3QVYxkJ6SWRb6FTrVj36QgdUfuCtpYawRET4o7UDWQy1RG2GL6JgSfqMweBL
6rpdjHRBTU4aEP4FZR8233Vfsv7I6Pd5OeqweOmAIjBUutyvIOV1VN4Z7Grc
i5TFSNj/fRO/stjcPMdBbfuFm6dd33RsuuxqoYu5CznQ730E36wq3oxoAAyL
0Shv+KYtJb9L+vb5p36T9OcT5TFd//0+a8KT9cbupXPXKi/Rr4cpE7wDGohk
y2rFO7QYf8SwPpPHHFLGx9gEV/UE2E8sGisxC1RsmGJzr62NqNw8VcpFSh8R
e6wtbdWfGDMGSynp/D4qvvdp9Eam5oy+yJuJ7A9yVxz1hvvee0abW6+mTlev
yw1sKN0qPOtbaoNb5wJRikiGiJyu06ltmbkFX1XbanywqV0JnBDGnSHvR4nQ
j4fet38Ihu+QWO+QlCzS/OQyGK/+3Sz7YzuW35tflwcjtEAmUih5bk+hNOst
EWUTeCteSvBzjUn7Uh5KB3MAWhOeKbKTDxmR0IODKBSLac7FHFTLYyDvt/bv
BSzyoQWqMW7Y91Dzb7haEU66nUyVlIdvBIrpeH2vYzjvfxmIaf+/lmqZ7dpq
cCEv+Do0zmKdcrCaSLauEUAU2gxH6Yy+OY6QlpY2+Rc2LsP/y/05dBlydtg8
E4jqlE5emFHTTbMsz1xtRjLdMYdCGJNIv3Yr2fc89RKHIzqEHEnZY1zAuWrm
3JgXyIKDXLdKHKV4jBFd0bDZIDWvfngCklEWQXYDImedUZnKDBlSn4XVL6MM
qwXJL8JO4yZbjxGwNixuMEvpYnnrIf8jk+R43ME48vRJOd49b+dZl1/oDrt5
+mk7UtK/N2vfwp38SeCJjvWTwcW5D2vQ49sfLkb+N7un/03F6dnbjGCqXqJ0
xFJAxYA+ebUceRmwu4ZrdB8Uja4StyQnbCQs3eF0m/UgGAoAtmeHMDAjVUpc
LTFF5E752M1daAh8VkCJw3BmGhJ6N94vXCbhmB3RS87C8ym3Yb14w262fuWU
E8Uj8u8ywHQlyuyBmzXyw2WxKr9JaeN7oJQ34xg9eyunh3nx2jUPKc7Xt0HK
7DaDqWD/sQlkF+sdg6pZp6EldQ5b5daniUb7eJbmhm6vopU67ksfbq95F+01
uynWSW6RfiT1/qLA3pBAHGmOqpO5+X/D+9hheQHACpwj2pYYjCEq1p66Gg4S
xBs1Ap/CgX85kZrQGwqMs1ifOh1XPefCQ4g1Wmo/MSFAKZ2mqg4RGlEZqG7Q
a8qZqQKxdXw2XtOfk2rlAWyd1tsGFHX5yJXDheKAt2ytLzmdLad2Y3fUyQwe
JQlGYYq+XVagPzos95pHVz8+sSJ4YjMDMnM5rKeQsuCbPBzwnw96qa/sbJhp
aPd1H1seuOL9zNaIuZn0r3Qsup/6o65sVBQdIvivDfxToLyP/iFjZ744AnoK
bElwh/ysrSU6HzShNrkOBzIjkS1X/shFnlzpO/zQFy+Ml5btwUltEi3LJJMj
IDVr2yoLd4QuNq51P5FwoC8U6Xq6eIEqg5TAPDM6golx4cqMFmS1+YwuR3cm
NDgp35ecxjY9QtQRngDRxdLrkXWe7t4vCgZ4ZuAdTTaJcGXQbUZcgR1bsukM
WadzTSA8tZ4xLHBnutdgPQtzPygR/lnhRblMUssdqGmHUiLQChdnHUFWY6e5
7NQcHFTWMrQQwZ6MEpJAAyniEYPfAURTz35JSBgn2oPtlxxZuIZs8gkBHPXD
Bz2/15DHg5b5szKfEgncGgGaDgnywK6y4m6AtKSf4EWzPLSaSDhsYhJ1GxDZ
HifAABvrQ3XXeL393onk6WjUzbwcpQSgFg/lFEM/sakpq6tH9WhANNM5LHfI
dgdaxZXk+cWk2QPrXjkQ2q1Jq5Ks8Tm1iikhXPBjRPtxHn5fPY8MWYepnqlF
c6vrHg6ZwyIb0PBrRBxufNWHVnBz9ptgURc6e14c5boGpzn/2fgqcNQwrNdE
F8B69ve0UbbSdqGp+jyll8VInO4N3oKGYKZnNhHZZYVZ4qUv7uHNjGGWIqjN
oWE+BEEVBo8puaxi0u9M2uqE/rPxgpjNOJyXPCfk+Ku+aFjFqJwryGoZUJFF
0kXykqN4IaOCDWMMbDjQZIy0CFJVQvEWrXFnOZYbanM4BCIBNWQp84VV0fg0
EyU+0w0djW9VVdA5vJ0qe4bfcfYEwU/CrmzpIz4VMpwx9a2QZ6X38pU2MAGl
9KoTPJCQx0mbCBxnahJ6s7PQEzh5HmdDZPp4If+3Ictdop26p1dNRMF2GCX7
d/r9ufiVlcs5VHxvoiWdRaLkaGJCm7GnOu7BO8skRP4spiR89ZYl2XWcb3bc
43S6CY22DyfXtFhd4QS2/PT42qgUQ3udX84GbYMUdB/IQZYR8RLsz2Asu2Hk
tPFIvTPGw0cDXB0bGyxvBVdtHVYEHKnRsJx42zxWbWtcoFPJ9+oTvboLGOke
EwwI+BwTAeKymS83hw/B27Z9iNWRWqTDrr5W2bnKhkq3QbViTrvmUrtYi8Be
UeBbnEZs+u2mFGu6wKQiMZbfcaNLAggCYLSXSkVe5KUDmT43l2OpMnFrPjzT
mSid5xhwkgGe72GhaXyyUjH6fUA7RDB/Bd6u00nPnznKwLt79L4UARMBSZBu
sVs1N11YJJVeXbNVushGx+YkySbrzv+KA/bhzdZadThf0wwLRrGW19ewnzPb
qxK7ynoLAbBbOVfIxvlH8pt8BydsRev1335cIflt8c8Xz3WXMKXG4HVm49Os
p4eBgcuHVYKmrvCWm4aDbhNm0XG+amGizIZwPLxhztNv6MZFcIzShML7OPbz
qnzG2SiuVE1wC+P0N1V6UCBFYBQwT5g3v+YAnoNVHnmj8xD7PSTDZxIdYxZf
7OipGI20GXJHiXaWOEwBO5wuVhIYq4j0HTBZhpo7YmeXH5QN97YQ08MRLKeq
V3uIhExpqZUQHYdacLHmUpvy7VZxgQdK0EgNwaMHjHzta7hwFZy88AeZJ1pk
efRw6qzvMI6WW3rLUsGV7xEUZmD+Obp/nXFYFKtNsyBVp40couYFNgw6fEeX
a6r4f4thLtrOQRXaAGr8VVftRliRjn1rAQPjnvMoeQbApCVZehOpCNPoqREs
VSfBgJNOehA9LXHMN00uSE8VBB6xE29mNJx+32FkhHL8n55o7iQB97e+vU/p
QQGVbWzA+gXtL1bxNtc+nKMyYtlkt8kVTVvudadspEMxqUTJdskrOyzukwEe
YEJ7+adNzRUx3HrG408+0ZjPPTgmVNkUy9Z5gG5F5/M+U7mojs/4MOZgKekv
DMzgI4P2hCurozu73HcZjmd3JIxOA/EfAQ7F8ofxMvrz4dUwZYJOI+kbHGCu
8uf/A5dJJ6UKCQFSYx3QUhOaG5ADYs3li5Qbv/OvKPvvJ/hzc8PT+PZI5x5C
00vjJQ4+isUDIU/OcACN1JjX6Fv2NhaW042s1QcA3A2PGLjhp0hJiu9J+V/d
WIgLfYPlv0rODd25QnD2uY4nE03A5iXWtQiPraK8uaJ4joYEARKHslI+rKOB
p0EC3AORmuasFXyJJaBza6B4DFhI21g/69BDy7SkJrQ5LepUMRzZo5z/ly4y
h7051aQttvIY5LoZqXR2XJPxg0CDRzt2alUkNxHZzs2rvTt/4QI4nKGMRlXs
aBfs2+oyriFmxlZmPl63xvv+5f145ftBnq83P0cf/p9oY7T0O32iSwN8XkZz
NJwx6vEtH5CRji/psPG0XBuZgVZWN/5e2HjHCE9f44IcDgSW6QANLoSlCuWR
BYAsVl84sSsiwnvJ2flEzKvpL/7Vgi8J8Cp1iJVQv3MSppt0LQOiINPVuKru
QUD9CQX23TL7nCERYwuyZqDG8FJjS0cdcYi7AGjy4u4YmQAsE9YReO0O9qTI
/hDYU7GaxQ+UUPR/WQ71LIJzhnDYFqPYImpRX8istEHGxnoAD88fmyYtmkM8
wqXWfPGETG6pS8D69C7lNTtOLMIU0TMrtxd+zzApMV6ObNN9j0dEAmlIHbAP
O4Ni8ObTfIE2+hYxOiNkqNHsivdvJt3HYGv+h6huXHXUAQA3N+x+B6Jah7EG
xcn85dwikbAwPfChLdrj0XVR020usxh4U124DYW0WlzQ/gmi2zea5ydS/qs5
nBYL4OYx0tsOlatEtqnL/VKFE+WNtdenpM8BW2QSzutPGT9yrxRD2Jf4Tdyo
8PrI+jt9j6QYJeMKbyWc6Gj27CadnadHwHmLhtaOzqExW07LN+MnbQZSoLfS
KUO+hEw/jBDo0VP9bG871e5W4A+iPNOYdFPsN99ls4i08NW7yj3D3RNNsUHP
pW/PCBRtPWeM1HXwy+RRu178ZhrNiZ4FjHvVmn9k+Rdmmn4bxfz06rO6QqyK
b6/EiHZrDP7dJ1Csut5at98xJDCCqlV4zW6uCr3oJWOUh/aRqJWqVFBOuSLA
tnhhZO1sYFjT9C093mri5QC1YF1bg0kCIJHQ4b3ntoDQcy3GaeU1dcj3Q0SY
e9/uzdLhwJHyRS435ImS6P0Kj7Crkg/RBlZdvQAya4oX72UJiJhgvutCpmc2
bHljTBrQrmgefE2wMCEefBv+MKjXCCf+8WBeUs4avOa471R13E68ZuJpfqPT
IUF469tap10S2/fDca7VgLtkRVfaL2xMnM/PqMuM9+wahEGM+78mqt0qmLY/
zlNQyjIN8wS+rBsQHdcQQ0YzjG3OI1uW4IxvaECXosZbfR7j6lYf7RsB0Izj
NbjDdcL178O2X1iYtfKxEQMsY84kAMyQ6+HLHMkTJDS8Fcg7cgx6JGYXdhwd
z8XSFZI7k86AKe1y/EJaV4JtGfXuPT/t9q2DQxzAAtT5bFQt0vpxeTbDByxd
143K28JO2fZsN8UxL0vfh/3CjY1gI0jHXdhrpN9qYWIpPEpZZFm1B2AmHAhH
0hGLr9lTtLwToErfUBEkb3h/xv3pILikszDKX+QM0mhtnznEe28sdG809XnC
+NgsAHtt2VgX0WuwdPTbZFq36J8GkfaRM305kvWtUpgypmEtVg9dldsYTvPg
uv4TxhXIzYV5snYxMpV7Aj/VC0CRPpLMN1++mefyaK1cMKXxigTj2K9wTDoa
V8yXgLn21AnqfZklS5oSieGT+bamTMpqVdrdmQTL2ql8t+Ch5Jse5EGPgJz4
6/aw2UVH1qPdUqidbNyzgK8KrufR/jOdbEn/3OZKkO9Lkytv7ebpzbc/uK8Q
8uP3UJjzJEAIl3Oh9C5oofBz0EfXMPhHU/TQXoj4F17xDU53D1jl+xNz77Gc
1spECBwo7xAwjLpy+I+SpltvJzq+KlzitcCuTxiQ4DOH5VxSTMSHCIWde/3X
GfvxlT791kDGyum+JnB/zcnieMIoMM39ShFlRh/jxq8ltdpOOLS/PRKswg30
BR86vIHH+8fiiRfd65ZKANe3MBkx0YEXDmnFiQ0dCb2YfOvlC2EWT8xSMywt
FYIE3znASICnQes/Pj/Jwr3FrtFx5JpiR2cZSv9v5j7vgL35JmYdtAwms2h0
t8hC2YdawIXGwv/9TuDd+0oNoXZbF3GqdKqlFwu32pqjxG/987vihqsEdcph
SzYaC/UAQfDlVtX3jLoBs7WGiy/8Vu7GRtUosndJ3myIjYvvAlj6bk9qsphi
+BLFwsb8pq1G3XBb9TkDvTCfUta+VeCT4nN/ziltZoJsmM1hzFhQKTagDkLs
rJQYKQNbalAM4NXwZsoPz3C3LZE1jr5tOzDCe6yxsJpThcPMWO3kcYACEmHj
Sz7gjt6eLFhRIIDCA/ktWz0SsNO4x+1WJxTh8LLuCKGs6xAdol4RnLpfTtep
jYY7CQRV/hrkJoEGssiJpMY/wb7iTO7KeNspEY4lzswb345Sk/2t5pMdk/yU
RDvN1yu0SGi86zP39Tpvv49I3ZQAyNUZ6tKhKfM8laIHe+7QY0wwjl5Ddzuh
ooDoNRkCwmVOJxQdlXtkFHPwALohCfVh/7V5mO/egm+pY0fEuWhKOqoxiHsS
iF9INwdflaTfCLMhPp4WSSc+vsBE9b08GgmDh6oEOkbJKiPgUdMZNcSzuXiW
o2PvZ5OcOEfWbMUNYAAcjZFw/rK1kR8jR5wIIq/BdozEcvIacSq158ozNBvV
r0FIzvcOto7vvDk4jNzIJF4QL5sK36nwXTFR5CR26EOEN4KULsjo+SdL1x3D
VOJ5Dw0Jv/AJZWdIgr7RtbBwH/u1LQGuCFny2igipzX3AD/duKalt/B7rkfK
11Wb2YelVbbE2f9HJm7QF3kEiDp+UbYuQzkmCmQ06G/S7us/r5M1MeFoxwBL
ku4BwIR0/mVdoAIy3Odwkf0/pb0wi4CsO15lEz8Y13oGi5aTxirsyXV8dV75
sJ34c3q8Sr9dw7860uITyJOsbI/+i9vN+wn5NjRfGGNg4YlfZutWbftjwBr7
R3UfqgWvUwbuIl0J6uSwPpLozRZoRbFU3Xns0PCPwbw5shcZ5kS0vN79mQlH
+P3g7Pe0OVwBQ2EGYsX4TF61nDVE9H2QQZzWxmhySMpg0kfMPEezIv5OPfg6
VLB92yroKR167hRutWhHW7HKU7FV6RHjsdOzgn/5ws0juwheKU3dtik9gBqG
5zAqN+8hppII4mStpP+idEbpBKX/hrVb62Nj1NyhPPQ55gvO9GuAcDajNnGS
KQ7BG4Fr8fK94/4U1RfQj461fmMdUfccrcdwK4Fg0c3pxo2apmwt/B87ziz9
5bWOjNCP80sdawToibyU67mIGGBeDFnfDGYD1LFfvBgiWcpgM+C+iIdivWSr
jac7l4g/La5B2GU0rIJ0AIOWuIAKfRgans9gKpJuHwctwuGEq7kT6jiJD/QB
xL/HdJ1OSjN9D7NK/tEM1Xt5mRLfHSdkdLffHzk2ryGB5HSwhs7okscMVYDS
QaNx0KjQHXSxnVlVhL7gLaPsBys7qz+CcsA4z+ZakGxlQDtIjA4cuYwaVpSd
mnwk+/fsgudReMEp+YiJys7sXUfl8F/3GVy9MyLWxBB4DxK45ApcnXxOCI/4
GY6LBNOmpbgokYwzFs48bYkIfhSWwvgAUDUTnKBUBAQR7ZZ3vcpd8ymkprY5
5dEVowJ4CNFdpHTZMxXFvgnJ+moxsrTyU+dBqyC0jR+B3rvaKRv0z/5zQLNS
RpcFcr3D2tA1XQRl+VLGgPSlHLPu/BV/+zoUlMw2ziyqSIPsFSQ1EtjnLWyZ
vaAGtXnt9iN/YblKi9GuorHvuNDHCBYD4Iom6aLk0RDgpFoJxEak6ZCniInS
GuL7NjTvk+5+Y7/J/lgynGwdEguz3aw4oOhmQ8eA9S/MWCxi4UaAThFz045r
9NDDIXLXE8wtjomOAMa87ifvYeQRuv0OO38kYoknVbOOEbeg6LrftP7d3uHN
e269t6Ofp3kArRFtw/cgB13bddtzNTYhRAZXcXpKEnURpBPUM45NxRoWP+xV
CJwEpb804hLu9rEV3HectJbwo9HumBR2dGF/Q6DqCjn2FwaICEwgGtmJ6CRK
t1G6mqgIC1hI+/3rBVRtiXZSgY/Gf/74SHsnS1ksDl6gbe41xt3cU5F2y/jg
VPNrCz1rHfbkAbmaC7xS/CjEbpu+GEriiWxCjO6d2BzuerWmk7qs56V9JLYI
U5K2uioJDREBy1/Hwis5OQwlL7R9pZeyvwqN/PCC4vBVRn19UcnyePsxbCTy
TdJtZ5uXhHQL/6FYkS4eWr3kqjtlH7VFjyLz5ykkA3G5Wdt/Je86fL9TYi5m
7WdTVS/OkjWC4xfL9Nd3qPDKPdR1NnuNk8A7Nh2b3rNu/BEWw1hyHytrUEGH
Fg2+SwVQRkDX1SHv7EYSghYqmeHFcuZTdb+A57WNK6qwf+BPJoJRNKsS7H2F
5LeGJKf16A0bASuLO0xg2wOqh7/wC2U/Z68VxB9FqQdCmm5ENm9J+rmVWA86
b3W8VZ3p7LMP45G+q1Pm1o+zespRl2fcmMzVtqPUcFgdQ435iv8Xa05lZVEu
fTs3hkp6kO/HWGSJna90jHFTczWCKwmZ5vf9O39v3TUo9QrpI/3DK6Fj9f0q
OY6tN7DncEzxivflTvoe32amAnXGl2aNGeF+NzjsjE8S/Re8jHkBqkZH2k5o
ZznZQQ+oedz6f5y79SSt+1cx13FPtyENGi55cKe1JqiInSrGYBEjmO5If8SI
5pB7VtkPG8AgnF1dE75uztHHz4tzLZ3lHFmSKq6EOf/RT6g6E/8nIyQtoswU
PPtE6iHyXhdnDstgXgT5yX9GODGCLpU5ciPXodmhQeqMtCvNH6jhtem41kRJ
rDBAfl/KBuMwydVJksbDK+igBVR4jOeuxwzfFfnRI9NNubCzZGufQhXDjOxn
I/Qvp6o7Y0uqrE2BidY/leAStcFfhijOa/+KciUc3SefHkhnLZcZMnTbMMwR
h+G8SDvNYpzwgJX98tsTL8F8/77wWcVdInuMODJArJhRDXzRuiC/pgaiLkaA
njulAcGyP3bUPX20IzMhTuc4WRZIJT6Ky33zVKuAKsIqaxCA4ter8Zf9p3SQ
rC3BXqdcnArZv6vUKBSuG6X8GKy9XArOVuWYfNYaECe50rsLu4L+JbnFCFpc
GIsVyoMKNageUmqPQCnAzr9F86AKvBA4ZQKGAGbkSWuPNnTEVoZidbfu7yk8
W/+I87Pb5Bz5IUKKYWRbQ1qXygzOSuJZuzjMw/GQIigMBO4evao0VH0z4z1k
ZhUHVqFEssd8u5xbiQV3GKmJd5ChVXfeLGk4Pi2AXULNGayd7Ah51Ory8uie
i2J/6J3Lr3/PBULKqDsEjn8VJfkoDewRLaJ7NIp9L1H1KrVWXSvBTROgL+Sd
pO12YVv/CqCY3PCLvhJvHPv9thlbTB25OGH7Ct2Zg7EeHK30nWV+fy/hEVNm
GNLOS9lmaq4YffV71oB6JsniwBdKwdEua9aBtWFhK9OjYF3w16nWlXVlYHAk
Mw1SQ10YnB0H2JNukxltt7LKv5vgCx7cNLvI9GzoZcwhG0uLw55FF7sr+koy
RoVfmkJa8ilazSmI1fCtUh/AFaWwAZrLI80gLV3uzEydnDYMR2fOqrFH7XyG
CK09bOwHzXzq7HR8fZj3xEMMNzuP4L2dpIxvtJk4L3YoPXkKE2DldP6YgYxD
diN+qRV9vI/EuScLJq1/ljC6S2gqahffjq919WbGT3+zcGTcUbBHYu7gfN+8
SQeoPSMLl+QU7Fht2PKzNwKr3OVs+j+PPEnIj8bd38ijOzWSC6DCWAX4ITdd
1eL1w0lDZnInOkybOx8V5EOxA/NZuwkWSwAtafgxJrcr0dDqpiJ/0R832/z7
WIUVekL7fgbRa8/We3FaikW620/P0t5LclzoSfBzVJ0d2Xzu+VcmDMrXuZ72
8mp+VGGo1pejoIPXfhZcsWlBBA3qgX9EOkQjkdN/YMVSNYcpylqPevkNIgsf
g9jQCejSQkeopvI00EzAZDYmV5fYQuCQoRTmde3ivbSTS1MZqxH46z9540JU
J5MdIxnmglyXoZZ4UMTBBYDSZATyaNjqsNxy3QXjP6ahWIjRJN1PI8w7Hnpu
9iRnL24dNv5od3sxuvyAe7NngivMB+tMEtXZKqZqE3Ww3ykZB4R58PceCxBq
/rLjYPcBiYVMev8unYF5jBSEewjSY1f5goCTzKpSB3jbSj1tsYeyYvPCA6HF
K6tvnJquWcndqa4Z3fX04g6vVDbUOs7pEHau5VNUzFYhcZwjRxQXt2ayon1a
B7QbWG6qhOTqboDOEbtFI6YzFKfbTyu7RiV08bxTk1NrlclboYQ0obSanamk
Na3JmbVNJL8kULUJI2rLA/R5LCpBUOcBew7XwlDhkrNwb7RpO5W4dbwiqxmT
veOkQv/rCu65dOxKuaP1tl6TT7dlXLmjL/Z35kxw1uHxz8ut7l9djOge0Vu4
bYxw0380FMJXTVCESkLKtbbFBO9XQHq0xsQdkcjpFaqKjsEhMRp9LivXJ/64
Bu8dD9XZcj8ztyptGQVzqVhswKvWl9nyLda2/Xb9mlem+EOtZdggr9l18eP/
Vw6PuSi4LmOsVKlg1N2/n+roWATTRpKBOEWM0NEp+EbRq5m/P7iN3ZIAHZCM
8lYL8TPfJ7OrBdlX2cbNbJtg02fuAMJpX+VSl8IUI0vpiaKZar04Gw8fZr78
xudNcu+cNBsgNTcxowJFToLBmjrCJhFlasJDDl1SspP0z8iiTNWdkbCI7LJl
rfpIzqQyPNso8PzpYvp6jH6lFl45JlHqim9vpkBD09Vaug2FSxcswCZbA9KB
O0cUBOasUjHoNRLfrNnslarFw8k3C8hrltRbaLlJsCc+TP3vrGZ9eu5+C+YJ
EUO4fPZJLRORDnih8k2G9y4NLu1Z1liMHQTyP0v+Nqav61zYwXPPOuRX9zoL
tKqu2FKp+TCIsZSYiClbYRZWLi4E5bkGM7BdhzS8daWUjvkHn+D2yt4jDNwU
pjMFxkM05ZEUnj2ujB25gI/CKhppAUPUVXUkyXugviTm6i9U2JQHEHvEzomT
ZPK3a/eJVeGvrGxN2O4vkCoHCBUkt4gIA/kqvekTfY3vBcN2A1wBiTrs43kQ
Bn6HTs1lO1d9rGQrykegwjR3kYWA+2DSilDo0SoJxeiYjqQcDTwIK4IeJBrk
er8TvAVbEAdI9ssDH6X2ffz8FC/Jai+oeXD3DPyvQmrbJ7G+Mn4/86VUE5LM
SMIx5ye3AuqhBs9hzzGsBwNvFo6gX75RhhCiowqZbdsP70iPXsiF8XBtDBWK
OqM95J/gni5fs5t8pzCiC0/8QHjkUhmSqL3oEBg8It0iKjjnfcBn0cC+fECv
bddm4K8n/B2sz4458uvkiSDxnHgecU/lkO+ANGjrFodTAlb2dWT3ywCIki9X
zvo4/6c3vLks5XQuYCH248LPlSuVf8P28/qzOGaFJBz9mDteQeS5EgCJpSqx
jEGvs3kWAdQKBVokHqIRUKmFq5RW2rKsdeGDHlyUIFdGo5jk2I+B2wT4kDxM
2/G472O75kp1VeAJ/jNPZnCFKzFW3tfgKCtQIUAJUK+slLfe3EPGm+rkwB4l
jSUZUjag+vF8XL8UVQCMNE8oF6eroz1d8M6lCMCD7Vv/vVNFRTYW6KoeTTH9
S7uVLupvvRy8ZxrMxdXrr6FDdnjz2jgTH6n5v5JqCyHkr3QZzl0rZP0blfUy
TyalmI0Xm+/wV/xlJbDwgSfNB+JM7oJECvkTXYPRAa/Lv1YJ3W3Z9UirgNJf
K7qnsoSop5hPie6+NlBpZTzu/aD7FdmN0z8TIneseY/QVNFUbhFlUY/d2HR5
fjnqUnIQuCNJNjd6IkP2uI+5qSkPknC/42uTIRbdYgZ1IeGGm9b+yNOXiYeO
vCneGQADI1TkubyoVrnLKbvgtEnPWYgcIlW0dKZoxDC0tCvsM5evaiFvrAJk
/zqgTsADdyBRgos7Aqb3iZ/BB3CVwn0jSU+9LK/GJ/C+vk5p8l09+Opzdj+U
OJPeZoxVDvyG292rksdLDRZMpsuRv7zztjpc+JO7TR/7Ful6wX7dP31/qMWE
QEL2DfM2cSS9SptPKGh70Qe6PFf8EPANbI/hpnQwC7xRkperXXS5yQIUQvpV
FDKqw0fkLvABu/yGs+aNXtg6gRkTyLFXAu02Df1OAMV33LZU5KZX2vTX0Swz
kn3fk8eApPGSGivGIpXOmYqsHQ3XzY9ShOnuUHAUwDKin49Hkm+OfUn14hfp
SucFczBv+Vf0yOtQbktDMHcA++yeEtoVx4sZ48pJ4ukS3DmA7eBy71C30nmR
jq1NARQTy+sMrj6CQNR8mwgvZ1BQBMYiXiprmUGQjJyEQPP8EkEsN4FmOkvX
BwJcj5os1jPW6OqolwNek3TlX8aG8hlvcCTgJ8LMkVxMazr7DWgdDeQNC4ku
2IOdRDJMxfyJwUtJ7oc1Cpkvj5FC5tPd+RGyq/AlKvTwqN4eMULPTJOLL2lo
rYsCoa9q9RV3NkvzVUyIuHlWLWf7Zx1dRGXVxwfPEwqd+fH9Y4qLhkdxnZB2
8P99diD/MCRwFWROBtFi7gg27Is/nb6Ze1pXgVHNg/V6am+YmaHOsbCHTmm6
rY/QbAG8wALgauv3Q8/tFW26KtnggvgmWQthMriLW5ryiG9n8LqUE9rLBetZ
AHlBkyuWAQo/yIIj7dGKZRuqJxUJXCMXarV/nC9iTjHqTTGlqoZljd9tLBhw
QP4bNLyatQmSyEVnbt1G04FdAJxUwaZlyYf3eo+60XDkZAFF3k9IXTbPZCS4
TeWay8TFpOsyqx3t4iupXw6pXnE7PK8cxkGjoVAV62l1EUmPTyVSFgoJPIKu
gtvN9aGUX59PkWSH1ntNibay1VuqiZl5pR+J9k10aU6H3S12ZNLYysOUYkN7
azHH3bfPV+poG9rjAwEkF9RRHhvjPhSyxP4d8UY2Oc6WhbaeZ0G3+LkO5xMy
Un9GThxHCUSgl1tT90TokIL6e10b+SoC8WMLs/sPSYbECjYzRRysSfeLdC7Z
G9NwOJe+/VzoBN/EhgdORw5gFHbHIGtZ7EgWK6Nsu9TDOt8ilGmpP7DDYXwc
rDVgh9qLYwftuiz+kt0TIvTPh75dnqHjVLOnVe/o35l+YtShv7/yglsz9h+l
EJVMx8fhbKeDVRLX7Hg7hHU2zxocRYHC5Y4QhitGbmVKTyt65xaLY0q6uEiV
NqvLGt4g89bZDlegiNLWll4lgfCnBvazkR0Y6p9FqQO9ucJA+FS+Q6F3TEeG
bT8Uer7zNUU/GsAtTiam1Y5Z6//HXzlI6Uia0EhkuKXQcoadTaLUze37xbGm
2V/zx2jEBqpcZJ1uT8cOQd52Rqrv2c2L46h3R8N8RTJ9kSmEFNCJNpApszTg
5jefugQHPud6H682A2JbGO8pbD6E5pSHOdYFrB+XFeptRTwYoefjDkQ9DJWl
5OYOoWlWpMNa5O3+Lgbi2OaHz9OQg+kqovoJ83vAg1LG+XgWpgB2rDVGWSsI
vSMyfFZE2PWHGCyNNqWcopeI/sHPuKDO2FfHzUid7Xee+6X3xLB185A9Ur7F
q2JbhavT/Cc7Fa9g0LYyudlXSdMJ0ucUauUwdNGcgLfKB2WclJvPIAtAXrct
AMFBaMt0p0gNdc33gdxSVKzqpmliV3GDdeOY5CjfxoZjjjDuka68Hb1yhAm8
rBHvJJiql/vyrKWT65xY+hCBmTqeFKFynPiaq06rzjR5KIJmO2cWxYTE+WeA
88Qik2DfYXHX4MnJgq20rtd689uR9ZvTM4CrTv2v1FAiznm39pP+z89AkDsI
MNJHw3UwdRP+E452Rz1BPmtaZN5nLau6/fgaNLsgGFB9lp1JFaJ0w0kXYRbg
5BmafdqhZLcjqjFSlcA+n1OXd0GcjFswQscdB6VJr8DoRdXNfOYGs7N/F55m
raO3XY7MfcKCtTzGDGLjdoMvIUA2gE3a+u+F/458xaAXvf2oxYHzB2AwQQ37
6xOgCV2FxfSQX12aQP0MY9Rk5fneBjSTqQC8SJ1i/9bOMTiqWfAbKc5sfW7g
OrLC/wT6G1LE0b0fn1/U9hOMwvz2D0OeNgdi3J4xyexfBdqYCgX8QRE5AhM4
SMmlmX0mpXA2bNQ4yWt090NaGGxMwN/w43WMBZqAcigYHSeryL59uCISWw6b
bLzN2vAln9eJ5JkO43I2Z4ZupQLAA1GYXyrWZmvHE6CHiZjldrSLAn0zs08f
Sqcmj4RhjYJ7PFFeeOO6rqU7gnuqqrWZeRzQbelOe08a2dmPNZh2ry5XZs5a
YYXYMdF8pG8Av4GpcjJFRNVXJyhEFjDsg9msZbT9lD+3M04WO1sHQ3tRn1tU
JTqtlQlc/ivzA4UY18bvDamyu/Pd5szkrsslefyzgVGIrPCtqHajo+61GA73
0tSKJqWyOPVbqGPKyJ1jXnGNHyClIzP5G67o7m9DuwyotcpUn+uMcoUeRQzN
EslXBKbAqAhUZBIg+FqRPdQkuikTgD7hXvdpt0nB+CZcSTbMn70Ah4jpyHIR
ngGJU4Jk0UdVwEA0Lt45DRPgHMvOEihT8jVk2PMTSsA+9zvIE8FP3uw+0K0N
61LdENkI8LmWC7oa2+B9z0txynp3z3IvxmuQvEvajjfb1jjeEXnuf+YbY+cp
8SOkGrjKYbAOJKeyqhnA3CAGh08tcQwTB0boTAUqngQnyRVLpkX/wTAdQkOL
/kAxY/NehlejioLbWaRkF2GM2scvUFRIi354ZNxOPLb2R2H3xSHKG6bihUMU
NnIyfN5M910krGzH9NiSBRGhtjSrR7yAE0GFGm7JkfnK+52XdkpqBgi+WPsN
ncio9GJ/KrDoWYI4z9oGDI2zU/6Tj14DqUlr6Vn63JGrYThTAC7xR04IMidv
+FHcsI4GIyLRp3WcjnJa8nq7xyDwmOX++IaWq5jjnrz9xea6TQLxOGZzVCDi
DY5oC9k/Yo/itaLn1DkYbX2ZnsXIOR3YsQv+1JjPWRRQpvpGzMAp3ENO36q3
c/yt/ytloV+EriyDa0IOeFvh15dtikYr2GLTM71mGby33qUY7UCU0bRes+GR
z5kcCPQ9XHYEIRkiJWgLtVTf0hd/8EbvTqlox32mVPgl+NhPB7R9hE5rBHl3
SFAm7VM3OHgsxjt78+m1nxD84wxQZswh3k3iYB50FDq9GjJQR6ojOV3CeHGA
gqvWIkxytvHA53oUVAHq3LhXcWfxQ5Tbvf/Go5Zj8qtktNgRmfCPyqgzVAef
95gjVerPmDpdcEzf06ZR5M6jHaD/xN3MrJFkBw9gyxim3iMMEiew6KLEla73
8DUrFFTZ0J5oYJaQiPB33q/apxJ3n32hM5PPhLtkZsC5dfetFMZjfGi6gy1k
aHB/vO+bQmGIdaT5limwc58CfrehBnjQXndeNnnhf0JWHwiYCTBNbYqQSnmb
bpq0ceRNDop1RFAOfxA/b6XamLw/xliYgKLFwjpTJDRQIOZ9K4KEYAy4a/N/
lWadrXt5AfSLRW3OC29bnUA2W1ttH+O+7S9ZBSjrvSpRFv/vlpEwM7xt1SIW
gYwN9+oeuccV5Bu2DuZNfaHa01BruxR0nHsgpt9qr5SU8BYtA1cRoGRG9bOX
365Y2Wc3LDEme6fjH7X7tNY1N0H1/3Est9ZddD7iCdqmZssMv5s6xLWDmnRq
fXEbqyzAS2x+qVN66GRbeVmdkHZF6V5AANc0S/QMikdKtwI7SBaXFNK+CWZx
X6qFHDHqrB4+Kj4vZG9ogNIpan6XRBzPfnp0mQX3jfWvPjncJ7/u3uPTKXuh
gIOM/gN/NrzaoPDR46CEf05xJuwbBQH/Rg9fiUOCwBvPJtsYUTiBuV43qg3a
M500vFoDN4smom9qW63Hnv7Hdq/RJ7OQiAzIvOOVzy2zcgVWDBS4E67LCOT7
KUgAgJQp1Y5keQI0Y4KFix0wIv3bNleWHBZjClQfFRqdsyoa0LWkBUQ4EuWh
3iUPA24aVy7zfA92wIwQnXYTpfJiMdXRGkZoWEtSj2IgwBerEAvhNceUilR7
AB0NmHWUoQ31QWrgjkn8xT9H6KKTSlQBJiO1yBIB/rsO1YAPX/X0YMFXEWHQ
E5hJFEhzlKjh4hUVVM5ZufPOs2c2ZGLI3ZduNk2xKUlDzEPH7lZAXVIoQrdL
YASmQHBpWP1kHfCsZGYbBNWp1axU/PglQFvVL7TKnJ1zxxNGxJ+ePd91fize
acLZnGixKm1ta8+1oN5wDcNHWwLKmeQ9ELL1+gc8dbrokhnkAozzFOhorO8A
CYd3VOx89rQWCPD0LsvUYx1qjZVEwWs22pNxRaM2fHkE/g2xEKlzMULyzEkt
sqI3zA04sKQQwvav/eZSJ9cCQj8MMETm5YWiSPLMRWVWL6dVWJorifwf41Sb
WewxldODLCgbPX6qXTWbcrPuNLwKpsNmDhYzRAY6j/5zRC4PKWQVrHAlIS3W
k6XXUDiLNu1Y3PZtEWYFtBNJ7tUowSAqY6xpIX3ieuwzzJYMxQ6IijWMsD9l
NB/6j9uenp7e5AWZOFKB4OHyOwlyHGw4qC7KkH8sBsq/UPvd4bC7N4DT/ELv
I71TNL8ZZM1fGNwRfo7iwuNhbZvBGGMPeE6Pxn2pzNvRwrviik77zdF1xQF7
hrujtHT65q0vkJ2UZUOeUz1ACo/qeizme7lLEtXU+Ano9qoo4xgwMpVzm4rs
EnABlrhuTZmti1Wnnu6TPu2xZiJ/VBo7uvIUv8QGAsBc/HHdrk4tBE5ASgAO
6i8xm1H+nuB45BTBPGLT8mmyLeZ24VBvTm32VQ6xLrBn962Q7fPEXfjlVP3K
NOjHMRfhaA6C2Ns59eMNJYArXMGcGcym+k99nLgpfD0ueZyBTd9tU8Z9ZgkP
dcFyJ4fZINxoRUsI154Sz3lVM45KUUpPMKtnM/XPzB7j95hWYDfvzbuiAvBv
TK7h3hVesvQaYEc1xXqRpAzOfHf6eDnQqrNtrsZmkbOT3JEuW5gRlF2nJW1+
Ocu+WyWiS2ETRW6mMFZDHJeOdYM1V6CHVP/eclM4LGeyeNwsne5TRpBHGdJF
JdJoHLp95Kr1Cea1BwLI04L5jLqD9w5e0pJaMWY7pMzqccfIpLBiDdw5YIjT
w0Biy8jLXwNwswCr/iVuYk/ScQofLTMjf0VXiBzYprvofV4hUVhlepK3xReg
/bUSvornSxfCtQZa+ujOj9rJcw8e3s1BYXKpcayY+BTvIg3sDfXizAcKOYPv
F+TgWjM2wJV+U9qDc/bJrlSJtOvVb6WHSaxpATlDIEdZQ7I9ZQ+q2jOcNNvv
n2SikkeSaP0SQgD73xSl7XOZ7RFiHNXclR6IUW6woXDAxsPKw4Q6Uiu2Jw++
tJycTjKuMDh+gX+mtIET/jSgXv7uT48PYtyaHEztSbsbEQ69Tx615y1dxzLi
1qJcDRZ3YoQCI+RCu1x0JL/6Nit8dak0KriO72VomZcRvoY0gq7I1rINII2M
ipdAvgif5couSt9laB1fihIPb+FFCWz+zj8CvdKQRkToSDfoM64oXt8FHxht
J9hpjpg3KhPVVzjPMG8wL6SoVfu8d30NqNhDT+6Z0RoEFQj7P8unRy48xJkR
AyQKBKcYL05t2zxqeU9PMxrfdjmUyZOr/Miuu5Otb7nCBy4AZb8YUSF1hyTd
+1lSSC3xpx4SAz6bN/MF24qvgUQOE6wRjd18qSSYVMhSFEhRaApb6ETyWkWJ
7InM6u/pldlDuHqGlieMJ6+WhfZlca24t9I60BQ241n0NOtlGPQVdKhJxx1W
fSo9n3Yhd3FjhVnK0Dnv/UMo1vKx/nnkd4+wEUJrs8+FZ1pyQe9GaCO4Xvc+
DXc+4yaOfYvKQneb+6c62XPHLDR8D6tMKgxo0/gVaua/2u0ryujW5YF4YAU7
JFSW94BGKH6Gesb+1oG5A/VCizgx0LU44dnx5Qv/qeP0TjF4Cifbg0vA0fxd
NDiP62o3Z+b3Q3ZmpQyY3lsZP10ABAYWdLN+F4/NOk/Bcp4vUZNaeeDaMcgQ
INEFbx6hmS/5DP/OSeJy3jMZNVfYH35UNSlEazkxcKaOloNIPkjT4CJDt0h1
6hRlMXJKRQQqEEa/BlsbbOMohE9v6HCOGMqHbdKAl8ug8ersqmy4+11zKSPe
J+synvulCUEQyosvzMi5PfKfwrxG8fKhIofBOs01J+JZMY6CUhljOPI9UjMf
OfbsM0uzTCD/wROyWZu1Z0CgP2W0QslKgLtEmrhg2xuJNVB7dBOBhRgFPPMi
YHluLQiIK+yoEfRLlSFxMwYyddbtDbzPPATROFKfaWxKGRKEQRFJm/AeJNU8
rCyCCn+otNX88+qQYuhN4GLooPKpeCyk00OmEOKI4Ib9Aeg+E+/2E1g9c11L
Sgp1I5FO3d8Opl8rVvMKm2LGECFKGpFMDLKx8+2H4EhSuDUAsOPIv15M9kRP
ZWvNLQHmOEx2IuBU9BjB8WNKwtreET2rqiW++dymb6QxEPU17LHQF0Ltp7Iu
rbXcSRBtBmaGzcvRH0gQlLC+NXXHGyhlRcFp2X28VxE0T7vAoFLEMCJbxVaX
dkAX3j6c7i3swH6LfsHXszjtGI8LD9ZWwqAN3nZ8OJXqxmWbLWp0ElsKs70E
8ENA9C2RON6F6EZItZ1+cxQkWxApINzFf+VxVenVnkXTt/bKUs5IjDu/vZ2L
9+Bs4pS21gQ/0munjvjrnkDS5TcoeyQ0iU/DgVKAAtKmab/aDIqZNdo+oCwd
IFOBYhSbgZZmu0Gf1Nyjj7HlzY5s1mrbEkx8Wk3WMN4NnEEkogNuvM7APW0B
v3PFLO17Du4DY71xqz3JkEdP1LH0dFhGs0Eka2SSYKdOCw+VBXO0ajUHfRU2
BSk/pxCRhoH7CqKTnx6WBVGyoCoUaa520y+iaWAiq9xcTG1esi8GRg0s3qh1
yNuaoG6s8Md3tOxq+8CuvsfI5gS0j0gWH3Nz6wfKRQWKgGu72oYJ8/FRlyN5
/TffeN8e3PU3hUD/9wxWsjIQ1cXpourcuhd57nk+r4iGxDMROcqewps5LuQr
gMgNP3m09PdNUlJtOCr8AnBwc6/aQgzexdGFsDMEuPbTPJrpn0rNpwMdQg3/
1TGNbZkX3HwFhQ6j0xK1VbCz0nsm3EFs//sttbBSbKMb/UJ1R5zYl0/9OuJM
9graTTO6LYiWIVFwo9lBZ3XE8d3KTiO3MTr+NFRsoAqSo2XWp26nOkKMNryi
0ZPpZwWU0iCBXj1eKzy+UrYGS9af/D4ruFbU1hPhvRS+lmenYCrMe0wbgtlb
y0D4padTTw/PxeX5l/MBm0HNeX78SZr8g9Rnz3s1R2pfz+hPWGOajp0pX0eb
wIbQefa6qe2xVUE0CXE/f3T+I0lqZxJSX8Z3I7VmGfo77eVW503YAQRpsCY9
i0y5NY+8xP9ZGtD8krIfMAYXrl2SA6izlN0XGd1YSFUHVT6oKs+KDpu2+Kzc
NjNLXFa8xOqEoerapv+Z8nZGSjTbv9N/jWE7+7LlJmC3+0pCGPOe8v+xEtBN
0SKCi3t9FAADMnh6Jwj19vgKpJdCgLGodGKcF/AtgaTewYTdWqZsU/WFL/5M
eL4DjSzd4J35GZ/7ek/BAnaSi7TAMD6s+HRCV3k/Tnpt12A6Ji8OfNWdv/zB
o3PkftrQaFGsxE3NAvX8jgXA4SccPNWA9DfUaA4M0CcYGrjgUAhamGyzkT0R
vzzZ3hBkT6NG+SOuLz/7CV+BAtuUY4YH6QiIh9pi5hQh9IcFyKe/5RSEF/XQ
IpatUHL287GaGI7duvvPLiF/3ZgAUMmsjJ1QTeDgSz9eOp5AJYq660XN4T4M
eCk/THr/WQMMcUf301qIDrqAKdU5LlCwmaHefuv3jsIWxNuvp6d85R9gNxQF
hWl9gGsSuKT9Jdm4lLGZ8cueQc8Q+mjySCPOJOo8yd30oHe4S/iCvLXKJgtG
8bTXRT1s2tmvLtbjp/j/GaTPxiKNAdwmAQw9NT+Tci7nnAjrYEn7L//00fRE
tmV9p4Z7jtkcyX4R4bPhVUH371ZHlFxMHIwe3Z9doqBiRYPvETWrcUWeo6UX
EbOcfR/eobh0fOXyhRQzaEY0X6tJbRGovFRLhll1O8UCEUcleX19wLC07uY/
Dn0rq8mScvPR0KKO3PMFEK6GJA+e9xGPih1WolIgGH5C7G/KIzL3ESJXHCI2
uneVlhYnQ8n9bPqI/TaBclUd9ObxndVw0gK9aWzOn4mXpAvXL91605RyGWQk
qbcyqYyOoVwBo7qlyIqcoM0+RK6VXnuXk5rjM7XVyPJ2z/SiGngeaVXSKC2v
nJM9lokZDxtZcrWoD916Wf5jBaLdVPp6MVxhRHXmUOa4DOoV0KwPGwZAVCND
0CPjweN3eUMRhgi+9JoNSaRxJfkPV2y2K/AJd6IYjk8Z3sGXW+/VMGV6YPY0
st0I0ZnVoV34tbbsWbrXlvL/tMVofCtUiZxsfQ6k+jGk0Rcu3gjq3hP/kzEN
G4Dvy5oSCk1/ps+tmJQ/2xsN0hxwouNXKRPQOngQJw8bi0wivdhvKxDXDFYY
ZTt80zbkVOb7H/bihTkdu/uWJZB+RxRoZMOlIbStV2d97o0/ztadk3a2w6aN
xl339IMLryvCxBZCYupYkUqklQm6vr+YQxGlOQA0GvMJKMxpOdDryGFLHw3D
V5pzyOuhkSRiTqT6xwZ+bQTxo1lKgSc2NVN2u6hs52/1CocvF5gSDHGBzRLB
dh+t6TmqYTJoxBAFZ2U1P0ZE1cTG6Zd5gmyNEtrlVlB5BaZzaLa6rGJHYk2B
Z8Chv0UwJLKTsKgX52RpLRApdehIBkiSIp5qfPfN4Gruzd47hmV0LqCKCRei
TCV/cn01ptQJ4qO/G2cPAq6ba079+Zijy3aV+7RIKYqzmdP9wAfKr8yoS+dw
gzPW1u72JUPFUvxeYeTI6o/JZpl26v61rAUEWLi0SOEy2dD6b2cX+W67eBWg
Fppn7AaEHamWCJEwvMdQnasd2RfOQMWloSGkyYgEXB74HvQZfP9lVPzyJEjM
bxoF9iU/JD+Q5E9WzFOQVrO9Pkfif4z0zQHA6mzZHBW8NscZpWD01xfnctJ1
/ZCu2/qTQpIPZnnxfk4hWRB7hJKKeGVWWOWddkm8lVhowu9UBO8pQRkIdLmr
sISKRULKjGe5fptF4c9cf1X5c8yey8RkVqzHf/O1BnEZcDi8Ki1KCLek40b6
p2Mn9eMG7fodH2yrO7CRCIszujSrQ7EKMT86W6tHpi57PxDqw5hNYOlSFxu9
Hd2ahlENs6SNakUMSmrPC+gPK3AAfSWdm53xEszVyQTOmdMw7fR+EpJjUn+5
ehdBuEu1EMmAbhH8+8mCdi8o4YWlYxn8cXcQ1DRe94ErqftW7VtgOtFt1dP1
nU6D1lvFf4ar4AN5dwN+GGW2flnPT/Xh3zzdXExDVMRihm/x0sLwoJgUsUMZ
DPPFEyV112gdsHUNw2iGJzLpvdUw3/N8zXV2aUs16SGFZIsKwaBuYMLjSx0D
5LiIJfr2hCbbveeQhxtN+ElJz6IVIdLiY3BZC5VC+ckulR99VtsKeYZxhoA7
dtV6D9wvO5tOmEJPJ673aizVkrGagmoggHQTdQgHnt+ARURkHwkVTgC78OOO
aJsGtjnXciQnZZiJknV6ji4yQa/7jsjeKIRLlYtVxCdboqGwwDl/JPJtNtWJ
qD6fIakMQADKPf5yVSKPvu4NkcnN0WqstCdhoTCy8YHcA+EUBwSzYymSgjgs
Iyx8P3DsPYrtYrS/TADISpfuG576XlNyc/eRnd7qNT7pNormFrxTSH/s+eLM
vYcPQIUBRcD4ndwE1x0SLyJ+xme9EHyfgWEbhT7aL567gL7+TJrnFlOgDWsr
isTgum4i/Rpc8C2dwXd+fiIgmNC0fmDM0e/LVN/loggEweRNg3LOmFEzYnbh
k1lpG+zJERJWLN2nuDpaD7ceh9ai6w57tWXL7PeatsdFhwZlf+DcBA+EvSGV
pQaLfxkMKEuRs6lOBtPkyq2pQQ/4mc0GqeOZIRMzQmFnu8KYcodtfuGvSNe1
Fq86qFQQwyBIQBDCVchWfrxvXmPh260OgUrukEnh3BMC0Uc7us9fbZs9xYl0
bbQAP40cJ+LnrXEylXzInFNxPY8Oy3TQ2KbpklIrARIBy6j9v0GdaGaMmKt7
4XCuiUgCI56xbU0RW8f4WrtF16W/Uxnqrj/ilgJGmoQqKYps2HV7L8o2FXBn
7aXf97k4r5BAH+Vqs+yESmBH4Ijo9uRYCVf1959RLBv5P6AwFJmwe8kNoCsr
efRNMY+hlRFE7Zjuq9IxpHsxcUxDW0jEwMKPvbuYR8LyQEWOswu3aFzGN0oQ
AsCepZxEhiQ6fppRubi44LH1BHBW3dqzHUps7KkJtyfQl2mZzKqO9VVrxZIX
s1QtGab7OSrljLgmWSa3tHkCEQdLvPjKwkucjvor1SCBNoHfP+FRVXBcgJGJ
naeHDLWAVHOeV9lSqvkuKsaKq8QWzLFgt7bX0xIL4fFXLEmC2YFK6drTouOS
ywHAAs8DzGqxnLMxzMnlkRcbnqrONBStR9DNhzZT0apubjk07NtoFDweGS5q
X/4XjP9uMZeJce7+mGelNpuREJMeYoQIH5r13GUx/X6Bsx974fzKcwEHMihE
K9Ll4Hr/FXbhe9Ueqo+6EN1Jii1fgEGxIEBENaQFEu/sh3BM5dWHLJiQ2BO4
6y8W4lEEmquVDyotlkHR5w3m0M9JUzq7Vd1zTfBwwnBl4pMD+gVT3/wO8aAK
r9jTM/+NkfF7RaA4uJ7gnsiJFz6kZova+HTagPd9uEAnwtnzJZjJP+i7826m
7c2GHBBFQUaZo2EyL9ZG+aFMkoUWBb+ebTfLiSVnC0XHs2dkZPSMlj8nVXKw
ndWZi4zOxL1djzZx3fNzZ/CBh/JleAKFCWb7tC97CQrk38T4UphgidCMV4ik
8p/Wqx4+OQSYS5lHPAYrfdeS6Cgua6qYSXD6Up5vk2qr9mqaSUIInAoQ3GQf
R6eS4uDh1I7cxpVmCrPhFhmMmqbdXY/8+3g5gYXFz1NCFrWDvYCmqRhzW6jV
1pQ30mWgXlGPkMVw4GJhkmZ4kWhCD+VCfY03QU0brbSslmttOZkADxeQlFQv
ZZ+WD+kwYzxFN4MJS/EkYiDjxS+fxtAJgczlxPkgkI8lbjiVeVuNBt77NCFZ
PuJmZom0FkFEzKR6m4mPkVvxV2PHC5onwJmHwF4PGqbFe5qz5YqNyOse9X+L
kY0ZFcwfkFBXPrVNxCI/1WGvxTY4SbbBKsnT2XOIkroTjp3Z0Tg6LLtYHOaH
yu3+EHy4bCIRxGpBoqmTNgIflDoFxjCPDDtnHcaTLfWCqgnenoY6CMl3nWsP
fTlzpFlcqjeipMkn0UQ6QT2PMLk5u6Bv7x1yEjsahkflfBLtdH+IdPL58rkD
jWSRg4p9ioYR/XRg24woCiynEn5MXTFwozJufGtdDCJWVGsVgp0kfMYbkrgK
18pwPC/2zX7IpQoBVO+T6r2vzjdyzjcqnrFGTG+BlOWhWA4asmVHjLOYjknZ
548TcnoRTNCikDNfkz/2l8gQqZCqwhMLjpCrjcqnqYED8ccV2NrevaaOflEr
B1grYWJlSleKaaefWfAvxm2LuK3ijdMX/5WrEQG7/eXVO4y6o8cgm7a+ASfR
WfmTkttsKx6Zh1aEaRr0SGGfkdhLCYFurh4e+zch/Cjpob8W69QeLlgUmJW4
xL1V6ANwagDNkiYNT1ko808SPzBz0YkrVJwNIPfRGyeVbKlAJszwZii7JmKF
y5Nidlu3C8DrrmyqA+R9ZWslcV0t5i4KLwdjo83GfClQYIlW7z+pjjYfW284
PrkF0f3kbPc20a77+kOsJlqU6WcxQjLP8aP+IzGoEhL0b0HIPnlYy6K6nr+F
iDppEJypS4JKRXQqXW9pEz8xaigv5oth3g0+J1y0a4F+SyrrNfsU0gDyyA+P
GAULU4AHiQkqNiU5NL6QpOOY50nRv1d2o7nRjHSHAHXCrWeglFD/DnxGX6n1
421BQVVh5pchVxRZZvmTi5dC4Z0TIjlS5LFZJe+sQ+vOWeQWh5ffSMkaXXOu
3nYffW1BHjiFTUn36sv4FVTPxKfo7sRVuo8IG/Bj3pxxD0+m2em8yAa4W0wq
mXNni5NoOOrgNF6N8WKwk/p5H7HHzcTn3Hyps/3gybpCsNiamkYqv429vh2B
PM3i06wQmBUXZbkfsOouDCd28yBE523AS7wfUUQY1AziHwLfJHaTx8GNdadt
vwdrgWZ/NSbuOcVGC8lRj8HE9a6aexB4zJskAdmeS0O1QQ6hl7kyeKLqpc6c
DzHtSJGUh8f54U9029ye151wvfQ5NGZQwnV3GMiFLNFmGuXX6ezeGP3qrr3o
lf4x/OskSE9OHNalaiPZbe74lkKVfNkrQRZr/ctLOjufKTv+X6Rs0oPPiPD7
it5HscwDm3N6jRc2skKTNBsPxrQt2McVmdhFfFGbj49cYpb1pMpLjMV7/5vU
Rx7v8XBmoNSJ4zCHN6vyMVnUBBI7GY8H6gPC2xymMfX6Z/EibHJhYy8s/3W6
wabVW+weRUmfUIAOcEN7d05mX8qDQ+mdyZZ7/0hNK/W+V45rw82udtYQOEK2
iuq1f5ki9Fvn0O+2JeORbHfvA17Y3LqMrZzLI2Hnhwm/OeSg5zhE8451u4bN
osFwusPF69pWAdh44QrIZSvZGzLHU/0p5xldlsKKNfIvmj+rKk7pnD7xljDU
uABpxEZrxfBrz0qUIhARN3akiA9sYt0438ErF/g5LGeq022YrunlVDmILe+9
sXG1A2X+jmuwaTr1r9ZhJ1Pjq3+rqVSRQQFpf/OFyFH1++77DFcJlQ8AM1/t
+6z2LKPLkwKNOY/MO8Kw1oOcvjPc3Rx2S+1Zq2x7sd+pjBNq8SHbT2CLvV62
QJdcDE4l321Lf07i8ipJ84lJKavSNrWoSf9gFHLGWW0AXmQ92yiMFuPLAYqS
gnJBKCx6E6GUr0W+t4UAjUvr5NbmPinHeMcsQYaciZ1uymNeWz6eQ1nSXB7C
f+sh0DqWzs8OLFPPu5VIbvFYTTwIvuXwG+igcL8AiLCsPV2c1wkmSqN1sB8K
xkS6hWFxnOT6odvT+seBLmO5UBPRtxe93rKGH8I/aRHbUC3Gaw9mi1ubWMNd
z7T+SV5ytavvuZU17hqRudb5gEWyMPcTmTPV/V+1p1qZwUClvmxs8wJvrZX/
ng0GLnwPW6NqaX44Wwbv+j6cYhV+ie699x2nIkAow4uPnTnV1SNUrEK1Z4RV
hM84H4dUA3G/HmC3Y842u33olGkAAvwYp0zSH9fyUzC+O3Ic/fPorQ12rsB+
LO6IUhCRNuipVuXrkcG/VfMtvCfQQVAwqkCg+GiES75sjgxAaKfzjZeCiby8
qq+QZBkJ4Ju56Fra6sZRt2lJ/cg9/0+yiJl4gAMoi+YdWshLkEROCmNlMuvy
+Hv+XizkQdSIBxZfodqIFGa2lFlMWP+tCSMxjNyE7cWnNReBODwTxU/6bv2h
JIplUUVzCWuvTFaEiztHoBaoRhIWPH0hiTMqqTTaUHmcSU7vGlTnf1wE2q2H
IIuDVL07Mq4T5FIw4e1OxJIayJNGX7tfgkBoOu9v/avkZjeX6OH+QhwBCu27
0MKgIdH6xOh8DdMiWqD2I+lnYloUUHDvV6xoERXIJyNoUJKsgE0zWwOaKj4A
OCnx3SKDmyrZ6WlR6Ove4jrY8c53dfaI3GF+yNKjK7BLv+NvPJ1hdjhl0Jgy
xQqXcrG6+cZhnEOQ35DscL9nyWdJcZtoYX9pNNeiYgs8UgLyCpQ3E7nRyvj0
kKFIT8ysAMTpuNoRsRmIEFa9dyCBowpIbsjzreDiQBWORbOfVcEdYpolJ0GP
sBsdtiu/hvaOgBycB2duiXhV9p59Q6duJVexwo1+vEG1mHBe4/TbwG2khurk
ChmHTCHJ0wXZU9BxGZpgDEFib9XNh7KPYaQU60zxwgNJC9o+z6idr30Xngl3
lNkCPFTA4WYZSfDmWWAOkua9T7RY7t6tPb1KeBpWbaacCluO4YUS6JScUfga
MIdyQOr0c910ibEWXKMXoDXv+E4ReIzB7Yn4cAEFPuhFl3XMN+Blw8JVmmBV
voJGOabqph3iCsPJxJhAaG78bt3llIeCHmJJBKL8gLuoudQiC8tMaY2yvtmQ
ADjP3KSgYYO3nz6eaYG3o0kLt9TMvoEo94k1zRz4IVXnjZCPjuCQWBdsxSud
tLbVBF41jxbK3TmNMqehXLlRY588MT+bfoF8cM627Lpmy867TYFMqgYR8UVo
g7Bp9btPM5TcNch2pFloxJfvKEXRvj2Wt1PBegzbBRfzIU02kW4ptbOCZLcc
NBKHeO7k4vGQlioZ8tO6JjebZSsToVvEzoxSwgk+G515emZdfnaCv/4lxKb8
hQ5Jb48I8FmrHNjLOtgaQ41nmkcGch4xvPqSulASPy8tSl4E2cgCoTTJQx6o
DiIvO+sdrs1N4/F+oe0l2iZ67hMf8ZvfrnGwL7CdrNs/YVjCvO6rRiznxyDI
OLsdrs8clXN8+4Prw2OefhORjjp+Xz9/2NgAFseU5/Ep27YZqxWUEWBYFXrr
A8qaKv7G23y5g1vO6pJYaBD6oojgo/dCJXV9GBHZkRNYupH+jq4XkvWFaLs8
QHiADmp5DMcDaQnPY1kwiXS97gapBpoekUBTWwo/rgWhHIwyLWyzAngGI24B
mNCKjIkZa2mDPKhU7/R4X51UUa73VY88yBkksoVlX5Z4R9sSBOrYHc7lyHWp
zkTIuUtsnhKJha3AX7bVal6KblydHUU++Il/9Kua93YPQ4PRyw0QuoEDMB4e
bOCr9kehKI4v0DbkluX+Nim5733ea7TiYSyRNxEaj6PJ2osvgho9pLtLlM//
lNXhFVno2LEjndnC0pg8qnZR9rrXZPbBuZL1L11jkxZ4J7gzJkgNSzCaolo9
xpqlbZCks693506qEHJUDnODaO/P+k9IQdP4JWP1PBPhuPFKnlVSAj3SBd7U
a52GJXR9cx8kwsWmuoG8TdvFOO2Fztw2kUAmiRz1rNIY+vWrnOqVfNBCxo8t
s40VY5oRXc+BBYZJ5UNqgHGRII6wPaZ6zqJiSowgupEMkE03v8XuN3LazlWy
0hRwzFFhrTBm0QqHVS9tFuRhz4mZdjeAhxBuSFn7T7A3imeU1+OS+qw/5vY1
Zb05StalDA9fNSy42ZZKQoz2TKL06+7UcpveoKI8xBLrP5l9TfWQCNu+EXGJ
3Y4J5ximBoyB2VmWJ8oVEeOGv4ObcObKljbRISRPqqpdxAQ6xiGcFH+PcOhF
VNz6JsRxHqbo0cL8wkmqy9iKMEYg9NhL/sDztB1O6heoQokqLn0+pIyZhwEJ
F6LSZUfeBWRe2zB24yhZjvW/aC3nlTfHfgNIYZmqN0l5zZPSnMqAKwJhjJr1
O/zL4amJLN8pdKvPUejjU0CULj+YqqtLu69OR3C6qRoP0XjQGo2WSJGsddUN
/TejPT1jJLHr4M9G4JvQDSQgQsD1teezg7LfmHO9hK3A7wY4qJJw1ADPZaU4
BqSQpjzCN0BViD0xMm6+hbgil1A9hOggtf5XnGBNkWOiQ+R4PhwbhayImpO0
KVML7it9oLq07AHeBPohqj9qh3lyZs0pt/k4hc1R9mAOxY76oWlUmyRur1Vc
eCJ2h8tPRmT74b40hD5rYNm38SJTo2dSSM6zLlJbNLg8PuugjP4x9jaJzRw+
TKGPHUFMcfXPek4fxpJHLrBKU55Kqxv28Isa8rdUEsNnZFaV3L1c5InuiB2K
mBx+efCxU30zlezZAgGOUBmrpmX4sx9sS1G7ftt705z18rz1rqi/CRBMgixf
6k2flfrhDJAWwMRclcWeZgzRyy6TQL5VoFaSeZiQPSoT0xEUOUtz9+T0WsR6
TgjCrw4TlFZqVNxKwe15QLQSkbTO67CCIDwVok6jIhvL64TbYWZxzXRGKTw0
AGGTpWFot6PSyUUIAxwU3YHz8xOQ3Lj7DrP+ee4Vt58Etc5gXUAOVdFDDqWS
QdVX4a9MXhsQ3dfP9rSHnuiqSWQbXO4xVLU4Btg3OSgQLxo8zJudmDY8vGqd
Lx5TOQz41D8iKWpY9g4HKGKpIQUXYIKktmLhRAydbo5XriKWZUsa9uUyl/Dy
bO9IAgKgAhtjPf67we8aUk/cvQaG9jnLQ5PTJVhRM2k1/CZkDdWCxn0FOdYx
NknNR+26lmViuILFTkum+CMUOZK8uydvGnfWo61vI+S5SZW0ATXhych55Rx3
wBPudZpmlsshTZRKUR28q48FM4ZyYFpCcrimPd+T5zEyBRi/wMYuxIPrN4K1
ePaBdYgcVDkIJtQWFUwdS7Lv8Ieiyas10oV99j+koMAi5dw4nbbaAFBMDOoq
SnwDcujMfmGuWO/ShgGpikE5uvwwVT+bgjZa3WMpnIWaIcdYP26rWp7xcqYu
R1LnHMDxsQ59bj/Y0Okr40QKppSyPYdhtZRH95jaWvMRDhB9MeNga1nqm5x8
IzE3qCyplFAUdUZjVxJtu7yEYXZ7tdzvlam5ppT4wB7zSBCjCatUG+0Qx3fp
36HdO8W5NZJvDJ88h/+a9iPKNsYQtwEwBnzuXY35IWS1xEja284q4iJI9pxC
7NEVHmwMekyXQFEMpkYevuChkRzwaxknzn4ekGgOraOKN0NNiyvur47Ev905
Tp2GBdEFngl8m7b7SaliQYa9rP+HmsyFTHWdbzaHWvz1sV014Lk/wkEky2fb
kvufbAf+tgsg2h0uho6uuPRmxz1pgddaGvXssvpeiNsrcDv5zFLXhF61WDLu
IG18Eo7EF45jF+esMSLhl5B2LAcrUTmbDPFXn+BI6bM1iVHFcZy+PDVQxSWg
HmRou/ovPo/26qZFJ8GQ+Lj+aluQ0IviRjfIfVN/jqZHDsetq431oslCnvxR
unB3bVfseywT3d5P+MLr+ESqz0k3m3Vv6f6O4TtFyCdiM+U8Kyp2K6PX8K/z
RCDXpclQ3TSEi4iMHeEc/LPygB95XGZtdhGovcRWL4AF7+zgc3UcxHZ8Pzmx
Q/lW9Fur0sxzPYglQttvdLoq/DkBoXN6pnglMuNUMcWFptwYjkxHz6HvkTG8
ktkmkmMq2omMaeV8wTfN3zj+CfXQY9eK3ABD8ixd5ikpRhRA5hFVQUw3rTiu
Ss+nrbCrkCJ1BtLEagyZ5pidhIKgoK5r0OG1kFtPg5cFblD5tjnTT0ccFVc5
O9vWT0qg/OS+h8tO/MBlFTEpKgTj0IwCoDYExVpnBaJBED/aJWrKp5RflaeN
AN00a4GgRd1ZXiDoeVPBsrYmuMEfGtTQEovW9OOyp1H6AkarZhavD3qu0SuN
ugw3jn2meodPWYNyR3Vda3m0aVhoRATlwssfc3guzB11toDuxfrFjDK1UMQa
GzFozXWu3EZ4va8qpwS7JOTsL6FVokvTluuMoR8bn9D+4RdzgPSy9jOuXB3D
827kgq2UW9i6t45igOZ0GEL+/PFkWlt/DZKvTT1+e8w4W5sAUV0Vq181XYaY
RnkHIFJl410GX9buMthaQYQdmXFsYXBPy9rvosx8CNFvtbkJ22MN8Ns6EER5
kCcVu0TE0wn3wvBHS7LME1Nu4d3goMpEvgcrF2D4O6ULlfT8Uy0sV+GUeayJ
VX6p6/v2tTmAycwDmGdGofNmljhHKvx3rLP95Tm4/LZovggjowyIyLNheahk
FqNRV9LqGcPMviPY5lAoGgxPwWxv0Hb+5aj8iwoPiuPR6TXIrYL/jt6LQdAX
UeLIJpS9n1DnVHvVGWWumpl0OivZHERFC9etCC7v1zlW42GoRg9bmpP6RE9Z
NQTRge/AUbzrwkqdu0lmWFcCDCeQcmBUD/G4QAOoltjUgqjz1zvlOweln4Ix
i234DAJHcvrG+yhbaA35aTzZ45SrnDxDScDSWQjG6oAe12ONPyXi5uA3oSTF
eAzsabRy1nNozs4w6YDDmTbW0z+JZAqVoo4pZnWcQDrYRo1DPGRcC0WdSqXV
9A4mQcpNksbGweWpqsy7wNsNGAt6u8q7RLwClrCF5eCJLyeUtqmiLR958e60
ke/lVP+fUXchGZDVXr8euMpaaTgB7MSdOOsuwmMmbaw8ZU6VYpJdyi8dcE++
qYmL+U+P+fuJpRl0yFA8MwIpnIBYZ23vTtb6fZapYRPtCjuWrjc/OUiD0PPy
mxIvF5ejR/EkPQcofVkUz08WNJnEK/xd/LACVJApOqwWkhuuRZj45GrV62uY
vYaIkSEOy2rTkzKAALLmVHNzIuZJFxmW7H4se/hwqdYn7c5QGtSw6/ERfOdQ
DSlcJn1p5XhFf75pWj968gidr3SixsUsD44efDjcrL7iuuHJzOmnwUrguBv/
Hts7PfU9S9fydjFirAsbFbDjgt/OFgHuUwil1Ohg2Ekqefvou5UVFpCbRPOU
VbXVnlQ3ZCD1V0egVVPACRaLxMwMVwINHMchAyf+GkTbPiLaOpDD7LKl6VMO
XsaGth/thVGPf6CV/Ghlm/PGtV1Sks+yn6vcH8sjAOLTIzt8Amo1X3d9alId
Q2i2Goh8V991A85gOrETK7Fd3Myp4y1QzXMpaBOUMF6NC2jrVn4q38qIIYNo
jM9QGvfVglKmeVIIu4qu7SZzpUpLHC/Xx18vhOpuauky59mgf3oVmlI/NCj6
bfjR6C2fXgil99P2SIwpXKNkFLouWhU1pFNGi4zbs1XIRXola0UIgl6I9+4z
w+NXPqjRFpe4uBgmTu28ArRBCjEVScF6rpZmsDoGX2V0VeejxZ0cXVUJHJnG
ya9noL4hEo3dCucMENj51avXqZ0Ffy33/17VuvXm78y8jWejSU30y975Ejm4
g4fetfEDzkoeE92TccJtlDgebd+bOpFvMX9h1o+cElk2FUMt/hW1JGLKFxe1
Sp97mUU/0vy01gkz6kE+AOo+IBLeKTwz4b6DfZXJ2+XoKAdJUaeoIt9wONEw
gizmJxwppnv3ZpI5Q2mjvjZV0ZOOM4d+DZN7rrVGFlbQMFJYF5mNetridJvo
4eKrSsit5eXrFjTdNRS4xKs+inF/CVuv6TW7/TBGlXP92hPS1SZBh0Hm7k5i
Ysb/wh8F/CU8VzAewiz/h6CweLlxzA3qeM/o3hTV18bvpYr1B4d6qypvmrfm
u92gK8zu3OqvsIY/aX5scvLGQ87cikw9SbC7kont9PPYrm3zHCX0ns0SwmNH
rAw2fYV2E1hinbbGWPz131ejqJ/YdzYfXrCbnCcUm47suykQcnPqKUCXrtib
AqmlSUn76BMnZ1TlEE3v0tj2dIJibGddExh4Ppb8oodWEHn8HkZeRMh1lkf0
66ZkjpErcRUpkJhnpoblOCjoxZt64jsWlmA81YxQC0KW6CBXdkFxuYvy3NWl
GsHtLekNWfhkelcaMTKIARVLx5nFyQ6cd1SDgEFpcDVOeS/wYhGqZ7fErtu1
8VWmOjfO6SWJ4JdWYS2jikV+dlleUBVZ4fgD6XN7XiQ5uSrRkbD6asL/qMQU
2R1DzLcqZXve2d/D0JXk3IBFDQVooDysF3Hk99rWgVoOrIblgeZHSwN3XjRI
F1wh3D7fcd5A2rDyRkb/EigSIgCaQv2/+jJ+gH6UfY8dcjl9BaRQiDzCMNir
+MUlrPW4jGOIB18+9CA+fR8KP95w/mOGe8GqO9diWzKWnVKuVqJ6Kg7TQGa+
L/FI1VegqYK+oToHAE6YriquPZhZ8UcSpMGNzckkjqjBaF+2ifjX+OjtE717
yGM5Z+U7joXWGehmtOds6qt2q+4kxs8grI82H752QT1cIjWSEGrnbYoZexlo
KrXm4T532cvG7Y0nnaTUzKCHRmqyQA5W0Cty2ThCnxxs9JcKuGueDZYWV/XG
IDsH5cGvyTp9gqg4T+hnflsiBjUoAkG6qx3ZoPekKh2OoGEE3DcBReROHoFx
rE6CFCpWDAfWKMAIHz86vuMwSyUTgLf/E5ORla1eg68O5SQJ7tqZ59Rjl+JS
UQiepL7Xc86nyToPpjezn8dYZ5kBro+quqmEwkQfWyRtvL+uKQKJLAx1MzAK
Ryt04qOQbh+xmxRpM23QfYyWc+S1B3mXaT/yMF510PpBADQa/q0s0djNKGTC
D5uqOHtCMgVQFLQG/IR6chG3DvbuMo+xdwTJjoanB/2HZ+oHb+QbfJMj4O+J
0mtmDQ9LE4v8t7pGnAFfCnLzu8rCO4+4R9O/SLKZJVSmGUaYFgtXSSKL3BX8
RW3rdg/1xSqv54RV7aEggm1jQT/+1oTx3K/MiQ5cG512cuzGVAJp4dQNBEqj
leC6rjStPxAGpnm81WuCLqUDpA9aHdsMY46IGrCwUoHSX7iLoACxum9co5ux
GrH1uL0jhvo3GBckDA3JlQ/q8hs36g9BZHifolxV/Arbaa4NeTHVTmFmCFQ8
92TS2OdVr0ryCyeRRbrn7qenat99It5O7tiarJqMHSqJCjPXo7rcF4zfFtpM
c3e46YaSxYzHNhCdMg89+C6/NxhY/3pWpbVoRHRmdW2DfRa8UofBd1HtZcyG
sqspUhBuK/2yTLTriQ/YjSMVYt3cM0CzEi6tvHl66LtJlT+V/JTUy/VOFtWU
w523xLYZYPqgA2nYGQB7opeThWY2Jo4THX6JrxfLmKObfTLctuCQe/7uoSKf
h4EWe1uwN9mv1NHF5FLCdyjs1h5yo2MdX0rpiVp+N9AfrO8BZiZRtucYTttU
F7hlwUeTExLXFwatS8cdB6PqzSc+Wvn1HzVNWpuZplEu6NrpodrTXOJHDElF
h9hnT6pXlXgF2LF/i6dttezu7q8Wb4R/GZCfjqBqdaNGD1NfypVWcDang70q
Ss7/v96OzcFhi4S8dQ0Ovgva4tWSoSW3lUV6XEjSdAM0//Il1Xg5WvKTBKg+
+NfYzBV3NhetHb3jDZp6cd61tTdOb3hwvICFm7Ri6Sdn/eWhqNu/LZfw9Li2
B2woFqQqGnAHi/zxOVmwrLilVvp8y6opdnbvCDpOUka4sd7IHu1Q3MYv1NCs
E5uS2oO7rxCskSIao4mbv7Jrh6XcFdg3MrYA/tfa1QDAOMUFGJLugbcRT0dv
5p3ELX9sp3/Vt8gDE0fk9n5fQQQEIOdK8fLEHAMsNGbzoWzSanvxBABl6kFu
xAEu7ZO7xGmtheI6R0iO1Ya09F0pjKRO19VAdT27gWnYjCOuMQe/thQCxV2b
CgBibdgJ7tFAAIpjK5yPRHQJ1O61+cEBor1cGdx34/M23Rk0gCfcmiYhI94T
nG+Wd4pvE7h9p2rzp3XOco20pmCvZtIijVS4ao4RhFIeMHJ15/I073iHucK8
OzsPdH03xSU0He4vMvO/QaMTja6k5mt3IQ6OM7gqqWC2rLvi5jCxiFFnJdaM
vm5zm9G2IHafRV0SiFGezP9Ht901YrGmkaxXRxhuych2hSBFr/IpqSGZubnl
ahHPHfC61gXnEWCzqrxWqbwPQDs3nPCISIViFnNxkhQH+xw4XIX1H9emsbmX
0T9kK3u/1rWE5hzNSbdR+FUDXW712eoEPZy+nQhdWCAt5sDoZd5BHsnKY4gW
CpiLlQ0amsEIygYug8EcAjeAxHIuuCyQR8A/gNAr1lYBAEpSwAaZHEUWmDE3
xxm5JISB/6DdhdSey0AcLOHMP3MS79OnvIR9KCLke5TSKOhrMn0eWCHyOP6z
cuVp4M4VG09mrKHSGxURlMU+z1xDxTGlHw+GLW4jifidszvc3B/kTpsjbRj3
muAZcXKz51iN8NSO0FNv5dckhO2aXTLOdWVV0HxkNH7j1fszTJI9uZPABwGh
NGbKbNgF42Jzg1aXYfkf+GvTGFp73Crc9gFH/4KB7J0Jh8PNYX3tA/w/+0ag
YVZUHVDOpBrwHpUtFMSNsvLTsz5U1yqkim4f/Re1RKK6jMM9roRN7AbP9AE3
ZvSsC37C2xudNVq5+nuLhb0OCnc6zNJxOI77fHh6UDaEIxZ1Oxl2mV2DW15g
sfAJMyj/eJKO+AYP+US7D1tJ26eBzR91U4fE3lkCiqAEKzSUlYXGIXY+3x3N
OGwuXpFrHDFI1FEjqvj/do4OZp2r5Ahb+myHCi0hKDraVylxEYktu3EV9EPq
aeGbB1FCs9kuIIagV5cEi1LWLA419Eguqvw4ZWWJ6uTA4faxpDGS769BFqSs
n5c6EDxgFXqY0ETMQdT2BhOoP1mFo44MQ1BqDp+4/k2PbKR9A9cPiuFjNQlT
vV36QLpAZFJEUZ9Q2eFQe6lH7HxPJVOHeIHqTXq9v6l+5i8OIZryGtVpTwYS
Mvk2PW2VwVaJR0j4iqAYE7t4ySN60pCClhQ3UdiAIH6h119N+7F0XrQPK6hh
hE/a+QfzazIT8nUclSOT2l+C9mb9F0E9umBY81A5iwjKb/t9taFhMZYPLfaU
RhcmQEViN9UO6GoUgpkhEAcMhJCLwjtxgyitLBS4Sxn3JTUyv/WeLXxVtwSp
jVBNwlwYytzEhqdpAfSwKda4Ie+dNdaILbyBiE9ann/VvoOqMgF0Bzjl9K4N
WsnoBMwVpRQWssdRcqXxfbMdzNeWs8dYCYBhBlqnia1+ATdEMS3ckmscRP3Y
Qjb5b/m4P1DoN71yJyBsI/+CMaQIFAIl3yqDvx7OxKGDZEhb9mWIwtaT9d/V
/cZQdckEC2amYXduu5LvZXr1IGvqHK7DKBN968pbS2DCowar98IO3VnDccFD
mIo09IQUjoMKlpuk/yPTlSDNEagnTs5iiALpZ0qwLP8YeYqvDugI1IDGTsoT
hYlzUHiAR461K7+fHyaqYakIAVSyntsU0ZGnstSHmEA8QX0PY/WSyxQuYk3R
Z7T76m8a8z+yHiNRePzGaLCYnm919mKA38GcPT/yOmE43D7RP3UaUdiSDjww
JwBWZBpO7dPam/z9Qvs9jTASebDj4XEoO7oe6dGlXyTdV18xGiIPFAejsUa7
DvULf6CLbDQxR2gkXYC89P3C0tZnLCbN+tpkR0PMxtG7H04WApeNpYRJDgLc
HllbViLNYgtO6be0L2tfgOJdbQhzareo+MuBvIM7Hm1iRyXh1dNe4AA5dlwg
PxL5k0KLGiiruTj988ABE4fHjDctdlrZLBBM468fp/1KhAEyuFWZ/hJjWVn+
ZZMzBo2WjCn9NS8pjIpEX3S/6yv9wjln+kZUmnwt/d2xLeWbg7KefXFwgCSC
zEhEQNm7M2YmddEnWqDLe1ZdTlaLleLVirymeGQqlvmUZIGNPt80CPOu48cb
Nll+IMq9dnzKCRnEIQxMFuo4Sk7pbaMS0DFoOwco9fv6F5DnxaV6pc7mVlG0
ZAjyEyg65Gv0Gz6V6pQlV9UUQTvSNfGDN6pWREQ/ZdlntCirfJBHK44k73WL
kZ04qIXaW/BAOUMlmJwOQb8/4PBWgrK+3inYUq0W8x0bQ6jh+G1tiWrotLvj
JXyAEf/dLM/dxFitYDngwM+MRzG9p5c7tThywj95JgdIvQH+eJP/3IDiEYnw
8PMMCIyhDxSNOvfuV270H9AL3LlXAYsG1As9gX4AT9CMgy1fVDJYB6caoOp2
S+nkhTWk4UesGkhChz4U2zPWAF90XfmhiB2FIFpRU+Med/3iO3Ra3ni7IvgQ
VpMG92E3nmbLRaVRL/U3l+b0Ux9aL5JmBBH2CaKWqYMcUKdwn1MzyuwLtIUD
FbFgWw7EIfLWq02J8U9o0k780DLyGWkvDAPmhYMND+Y97KY1+3b6fiaTbTa0
gRsC2N214yHecAGnpduH2SS4LfiASuog3Ro8T+R2XUoqnLLJtYGFhOQtP1Jh
gTP6+5zazGeWoA+71UKO9PIkZWrvSpEvPrfHy3ziO+X4IMJwy75GEeL8OQ2h
bg8/zfDtJT4g0LFbzABhaKtyi37mJ8iyD0VeS+I5t91ta7XEqSzn0xGcQJy1
vHnN6uQ7SAXoPttXt6GmISXLFBMDgRzY5h/geHCejwpHOKhI7RaFZlrlQFfz
ui8m3leLSd18yYor+cg1fBUCAJBGVF5Qj7A60Z8HyoY+MMi6jNeYja04uk1s
RB0avyAToYrl7GAsfJtyufzWq0kKn0uJGIz9mwckFYzMmnZw8ZmCDRgsg/Ge
yrdXfVAnOv10gWVH6XW9HLElRmxAoUB9PG23LdWmIoKlpILvXqMrPneU9GpA
rw+eCppy3KU7HsTAM0FlCC7CVXkDZgW4Wgxl/0u9gxwnU5384A64751IPgWw
sz0W8vKDmSWJEvKho+gomYSl4SaP4/mDgPR2ZvIG31M91WoryL6cW2PEWSWU
5hJmHLIPunAjdY8ekZAgfvCuvYCjRffoxW77a5lpPES3Ns5ZpMzmgT7V4h7F
aF1bPQVyaxP5IK7gI5YRIbYwllNA+vRtEqGI+Y5joYcnB8IjpFUDw7uKig0q
IrYC1ZlCj8e8xTT+Qn/H150yS39/lln6jLNP6Pa85DqCMZ7L52p9RhhDr1UN
DrpB9iFKs/ZYTAcBNygc0E8OyXm4iM0Z2HU9aqjjWqqqHh7LIET7jYEHlTbv
MKiJpPPkZP3tVrT2xXo9uwtoC39YKhc3qDemzHy4rtTD5S0tiQG/SXyVD7eA
i/A5GBLIRw31+1FViAtn+TXzubcafbQFIQgYZJtHJuMl5qyYOv+k/361P9x9
he99bSlf8ff30T5ToxkdtOsLJckVxRrxTl6VBMv/RIYl82CIZLKljeG9a5Go
qDSUys6KKQvfOcvZW6RKjlaJPqL/++w5W/59SqzlOVIPZPK9bbvNofXqpfP2
ZQrnkNH1ghC54b53LazK7KYdbgNC4cvXx4kUWGCKBRQ94dIG1sQJw1LPRlNl
qdl/ytQJ27Mr65/iVmS+6pjAw4g578tmcpsM8XQk2T9Jhk9a17NPp7c13p+e
W8CGIrKQIO3DMwq3TRaAFoWgoWy0/1CUOxzcbKEw9gMf3tYfSanbcg0Fcxvu
Q65qoYvze9DICHnit7DBXsUImoJBH4Fs5zZdod7V7jqQ+ohSPS64+So42RHV
JeCJ9YTtROs4eif9/ZKdbPzT/sMstx3EK807rtjA6lCAq+Msuu0qRTz4mZ4I
hlKO3IdFmJEe87lFrXLDMW5ZGG81L3M1ha7lClf1Hi8CJw7dEyQlG2YmKxhY
2ujI8TEdUauctEltKdAicvDqM0K+DwyhCC6s3RfOv3H5fz33v1s0vbvtmjF2
Le1cHG0lhGW+yglk0I6ktBm1RCb8Xl91G2k140v1tNcjm4ts2fsRtPMyICdV
pk3ZDHLuhCUtSD8znUeSvuwwfbDdXE7AZF/k2OHB80H4HeAnGBpSNz0eHA0Y
89ZZywK4Y1uL2gCjXdhWOONVN5ZPSAIb4q46JkI00jDu2Dh74mQB201KNjc0
o4LqQBdPvhaLO2kdnfKo0BCN5wWauDf1LN123o7QYyHdIFODa6grXYcKzuOy
A0GbmcebfehHzBV1qvlJPQF5LmGZmuyNdLttMe4RK5nJd5lA6AiHEzrgdAlh
O7BS4ROMCDEef8aPdWIoa7HgGB1y4CAPCpDTFUPnIjPmllyeHXhCGV3cbv4p
QhbmIXqe9hZv35Ia6FXYPArkJvFGseNugvZ9qWuJL+fTlQY0GDvdzJnezmvz
XBUgygHHhgT/q+XBrvpQqlT7QyOYQRqlLgx/vi45QVQgWWkIqrTb0G9ESzlC
l1bXZcLt4sg1+KLfal50ktuW7UP+fnhvaIqpy+ka3tEJgTgkwdjzNNS6GF70
7/MMMrPld0jlcLHHg9yqU9GwNGCK5TjRZ/GuhZx4FOBURxpjXNVZV+d67+9E
c7WwowYJAHHD1WiD4Z9pek7OCxzlPlbLvZ8Cgu+mm6A+MYLRqWTykNJYRkOc
pebmzHRDNPzOILNofz50VbpXAq59kUSZcjD3dJXGzY+ENMe+f+05Mam8gkFK
7nKFwC5cynlG2Zsd91+IQZKtQhoYgNoT/Z59oSCgNP7iqnJjSO4M5qsuuuYN
ZM61SmxTqLWcLpd2S6ffL7VGaOI0SH4oDcxRTsXI/XjEQ+NJoPYs30G66Ols
dD1vGnSN57WX04RvVtjsuEnDMVCDe9liKbFKi1SwJVZGu0VGlE7CwwMSk1bG
y5w151edtG1dLVmDxWHPfEuzO+ej2vqY424JG4n9sJKBJEUqdWdlmqO0pNrY
zGw6Hoe8Xq5sabtP2yaYGMYlyJYL0de2fm7/05ta2nOHLRh8COslnqbMr8xR
n2Iz3AElcdwKC731Ejunu2P3noex9o2kMAieAfnA/zxQYV+lNBp2Dm8Cx5hQ
vFVZxXk4kLTe1EukCf/8ex0GV1NDBXAMMyet+54wjweqPAOEvRR50rCwRLVH
Rq00ds00AMdC8Tvd3eCd91if3MJrcSzLKyYNCOwEHYOHZSltYxaOhXqo6MCj
pohNjvaHTJ5ARXGBSFWHr3n0252WlCvnmStazie9LBXsuT7UU9AXxZqmVd3R
pmID30wEWNwo6QupGVp0r3ikbI6GELbeLeowNslevw33N4tJAvngQXMKsOd6
73e7lCUZzod3VBjYeqyKrr78AuJGC9UDNKbipjfcyN89kv9v7U/sX5qzEUMc
RwumSInjeYBAnPPC56Q8jeJBa7FWqtXxHQP7o0dm6quIwEt7qZQCNf17oVm4
vhl+C34C9jWXNqqq5y+gRiOLkr7ALrxJdYNaJ+r0g7xNm6JJ7p38AMpCSiJ6
2Z/xDQqRhneA32GwvlEdEnb3uw1jOXoCuBMYFmvcInlx7BBmBDGvNYU7sU24
zm2DyyfiI8PsYL6izg4OtSoa8y2XMIlicxjyj76PqsaZQ/c/xOunUkDDi5sH
0dIfCGYqk2pyH7n7sU36KqesoEcASJs+/T8eNCeloX1CFWCu+GAk+O2bGJwg
I6BiegjtL3lA7KcpVxvG74Fe7yg6zREaysqoyOGxHzVMVTRBs6Nw+ql9egDH
/hcl1+Tw2MIvLKy26Nc3GYFZrquYFzcaEjxGtg9gxxAREPfmvQJP4gjaQjrO
iDeH/sKMw/Hlldh7Q6xP+6IFgUmtL4JaD7BZy0c6/rLpaax4dlKfz9gDvPSp
clsVmXHhbmjyJqISVieptm5czw3xAOu6/3TPXdRYqRf/i3tqmFXLgmerzyMY
O1LaKamev/7QIC4bez82WkWvWv7ZfurdbiOZAqxS9svSmEuSn+zepJvIL5pq
O1BYECYqtjCZoOcwGZNCWhBrjvNyfMhdo9qJXlThZnFQD3+CV7NkuB24HVIL
uPGxR4kgraag1mZ2O1ksTS69rp0zKDZqas2NuGsl9SsRfoh5NuO53PoBLyZ2
1SiGZQ6ZIGTSoUZgv9gSrmcZvbX/DIivJI3t0+y71p4aQiRjA8fdu0tWYkGA
1WvWG3NA1/Aw4TYR2b0hZFvwVUiZ8JfDCdYMsvKi1Yu6PkpJl6BNsiPqyprS
91fYtxkBsdUVMj6OioaxTGwpZw92TuwT3JJMRK7S+UBbaaBQaq5Ro/719jgn
DJ0CkMkW43wPfQ0/c5tCiRIZFsLHB6+NwT3Fal3pAixp3VeKrFydqD2jA1yP
WlljuCJAhAaB7KbDhZl67AmIQpFabl2N7VZk+JE1BP1vcl/qT5EslVEJnAwJ
m6X8o2BvPQApazJX1vjdnVswctwiGWN5JUkt0s2bSUXiZdu7llD2sRJhOrfr
Y26g4pSMftkvzpLzrBTv3WlgejaSuo9WoqgAVzSZAoazfcAKdlmB1mGCXzTn
WLtJedjETWJBWU6yM8ddvxfur/eaueaJm4JN2pAOLXUIiEhKCYVutvcOcPLx
e+wMUJHgP8LRfkvcBx3LPgDoC2rAqPPIweECGPs9YkkhdpRCACA9dUhhlEq+
Znz3i3dC0f649bakPtVjppN5D//uabBqREW2x95ANCi/rKD0QA4SiAVHdTTG
pSc+jpwSUXSzJQ5i3YRp+mnyC08JQ91oa8fU3se0awyTO/2dMKVt9Lx0QCxy
yBcckEwb6+dPTU8ufehn03armvCDJWN6jojhsKXpBNwNiLoY4iQIowmXQEco
oMgFI1YUfBp3AMH5n+lc1ekr+oVFoq9mudhNHMTfSyPlVhEpMFuQbhCyyCKT
JSa7M9Bw9/2JMcaMZTDH5NTEpULDfinzU4EV4w31WVZ7knIMXBztOxPywXpb
EPxUDfNfIgr8EIck/8L8socnybKIX99ki1RB0itJu1qSxBBbcUXdhmY7hClT
YnWXUmMj2kSlaWYyvnxYQZtEE75ALG3X44WTmWjNiTYn18TQQwugzFq5kFcP
XD9XA4c/XOJjKGCnKmkNt73PKoJqzh+B+w3goYVI1QfT1IohYDu0vLwlWDxJ
+YKFbno0B+x11Rb8UB4vxxEGN9tpMoRZieXKPsYOLLEfQZBe/3bMkKTG/XAJ
KgDrvLV37aNF7ADV0WzhrWs/hHKstXkk/6pYEjvLHdd9ld9LRZowGsyqxi0o
dSN4cvCZX630L/8ZslkvJkyhmVzKiFT2gvilIKGxQBaMk5D1EkqjyeIP6YdF
zMrxyG3XzPklvgchBvoOWFXZSnS4nrjdWwpVLwUgCpOE7AWSoWk0HoP6Gkq8
v9sB3UV/dZUpmISXCrUy+HHIChZHWmOzOzN4znP/0V/SWiagA24YLN6WIsIj
yceE9K2ow+hcyE9b9M4jpLu/vn67XCn3e37IJutKDnxLuHc5Wy3gruajt6IX
KOKuejCxcX//MSwyea6nh4SaHz6AvCS6uI3bfXIDnjfxLqeM2lhq7scVog2h
fAAdOofO6j4STxwxgrB/uXgLQb8mi2dgtFoYS8qZX5yO7Xf+y24qoejRWu43
ZLza7fHBgQQ7+5qXgsRn35HDSJN6n02YCDBPLN4w96ZF8MXeW+oTpzxRSAUp
QwZhoRl7AxYrTVGju6fo1EHBdYIHq7koOAQ29Ylr72sD3z5lazsw5b1Ys0kB
eLinkF8/5sJkFYGBAcgjbZPmgxp/gqM/0OVELxmQ1gcWMCBrCfm5v0xd9m9R
c1dmIQQILnPDzR+MPTz5iq3xkWM2dAf6yyd8v5y5AIFv7tFWJuZ4nTh8lPJr
r9vvQ2XhdoPREZ2/FG0LldmVh/4Rm2nV53QoW0RVLfLoYSvO282udD/+GbE/
wHP3W0H4DGVSBCY0MtiPBJI4N/72iGzLBm8s+cd1t2+p7Nr/tUF768i75VEl
xxKYZd/VuN80lrVtCu79QESjd757t71cvObCYSoRWsCxOi8DgI54ioQ5SmAh
sfDNKOxiBlxRd64lM42QxGNYhpeEMsBa98kobZDXZt+Y2Fy/xRamnOJazlNw
dF8FmMxRZoxQQZMJ8bsWFVYM5mrU+NvdmlpKDd9oai9SWzZkXsu/k4zd98wO
mnc9rKSyVO02CDkAm083uQDDnmQFLDjA/LOQ0jWpdLHpQzkMoB1UZt4fTpR+
HccwCuA0M2Jye4IFFdiL77X808IS2V9L4H8HQA6ihAkI1bF5DjTy5riJWqYE
UobU2AmI+GbGmq5pr1JmNqUneeH97LFr86apqKPqY95P/ZL9j+GzeuNr3sCl
rub7+hhtRdEk5YFMa42xaeauBBazGiuP1/aeaQQbB3CuhGpNBtkaYyt/4BMh
aOqt9KP9XYhQTJLKrp5blY7vzQfqqloirB+oTXRSnOMYSqyrn8vdxorwhWut
l8vHbmL/tu4Z8hJb24421PPLCM1u2exbxbF0uEFB6tYnW8VDm7lZ97EkZHpX
mbDURX3hKPNZP8acCdd2n9urgwsvznkYVjY5wzWdrbJsLR6KP8lqBAkoijJL
5HqsjQAN/SefhasRrg3lrkZwdt0MAY0zqsaheK75+Rdwy9lRfUZG+KM/vXnq
38aJgD57ySXlpbPrTPlIusFN9JGw6PBi2ubroWDXQGX/hfKXtUimoJyUC95x
gRH49owaiLbt58LrR4PtQAr5pTq4/zfUVV+D+jc+s/XeML7f7xkZkexFr/F4
Hlf5GZf/dBaJwdekIAfNYMIPvka7FJPZTYR5k2P6ZLZzDae6Dab+SjRNFlGo
nCkr5sC4RQGW7CCKbnV2r+zv7cvus5lqmsOIb7nMKXdTgk25H5UK8+NtZ+Od
BrcMrbGhPUHN4ZdXJu4sy1mpG8ZKk+vwDDkSxA83PSS2fPVHV6ckwjhlhPKk
loJ7NgtHnzPExmtJLhxOfjzeYc8AYX8urdiQflCzz/N5Lphjo7SQ947R6PZi
EF0AiA2Li5JNYmbTgh9QUDZjCjaE05ZTeQ9RywHETwe4B9MO1XbOGAhjP1vK
bjZjFOMCu6ZT+6OfUJskqWstyn2FpFv1DVUcs49H+NRUwjDU2fRJAXJ5ABSw
4+gozmMtyqejEGjNZhvd1wGZPIXcl30DOl0DB47PgHdgD9PGY2lLJ901G7w2
u4lo+R3AMjIDx5oGgdSlbQKQ/ko0GQN1T976a9jgCl6OyAfU43P6gEhEDU0y
r0HA/C660NajX9mi7RQcg8nuLo5/HeqFOvP/6+OlgHtxQdnXL0F6L5g7WN4c
eW3+7SEoarvtxVADaGkFXprguH96ZBLCqVmoziC62OyCJK77VpWVUerFDvkw
6q/pzExXvzG5z1sgSlssXe3w9K6s5ifVhD9PD8iDx+laJ/hH2HFE5nInzV0E
Mt/uxwcKloKldsVpSdphjiac2bNw66wK1mdlj+FukuCxzsrCHM2PomXmfUh9
R9wqQhP4u1zs8KIDWfEDvRbp+A9zV3DxXZjkdu0O0GMAxmDexG0ui6Cypum3
7PlYVp9H/gB9k3LyLaDbduX9f1GSI6qHYnqSfnePu8UEG+uHOHVr/mlQr37L
TRYA5P6wHnhFFnRn8QcNHf32n6QL5glMFsvbRTnpngPaDykS5Qw5RSo8z8RF
AjWUXZilHlzCqXW2eUPH+AIjZt46qQEfGuSB7ZvloK880xpZ3az21xdcYJ9+
R3HBjYUmpLoH7E+YK6jP71g+9Ar1UPfJuw0aXknWLvTVb+A/I6VvSI/yvLbK
2eo1geJBuDUhbBjMqBNXRITGQQuWcBZ6JbYMDu4ci+SffZyu195n8oVmaIgn
Q0QAI9arTNoPZS4us047d8pROuvL2z0sGOJGwHr93tc585+Tpjr5/h3ZdPIl
Hods6PDTNAdNrK1UdZfovT43mBXznwlsiVq74eTo5QcnCIEKW73VpN4IBjld
wqaQdrPKkx5QhXd0mWdUcoAhXLvkux3Eq0VyCvSqnULS8R3V7V6HGGSBDgLW
lQSINlmZCA7X1oBuSI3QluyabSzQhhQ0XNGkC+zUgA48lpdPhpJuZQKIhciD
TkwVurkASGdS8zcLataaV7YCkLHh5zc76hSKVK5y+L3K5N2N4QCJvQ5wQlwu
EnXCWrPTDxrWtInSURrWys+fC0xMVPjKMO/KhRp+O/ULGE+G5Dy72irRbXM2
MAJ3Sh4f3mVx3ZxBm36UeyKSWR/J7HkgbZ7AnxoW2ioX4zNmGHdod4B0+28H
6jYPwM3w3Tv8haPIGikY1wtpb5xYvtqshCUYxOoqWirjFb6tUlTYdYEN9FxQ
jZw8qonEFRJG9fmBBdzbeAvVwcd0BnfvcV2/UYxLZ9G/Qe+LHEKsvDJkM0s3
AydwDUBoKECPRAJYsKrne2neAA6mEloc4Mz3O9qQYh2tz77d0oP9IIgQ9EOY
mHa1Z6b7PS1h90QwauOZzdd6dN8pu7JRBzBYKvAKhEvLKjJJdsOzscKVR4kf
t3cqLanPO3YNmzJSxt0PjblI3W+LBsxpojNDe1PuHfK8/oDObtRODzPw/WV5
Cn38NRfTwjad/D35qAFTFRYCmzasMq7Qj3xec7i/CU+bgqFAi3RZbQVBnbcd
V/Zv2NBiUb2xEYjYDAIkzt29s1XRrafiCNpWXLoefRkQ/nermTFkI/dxjSkd
EK+pWDcmA189hQYWlHC92RtZeNlsDH3EDvMZV+E3oFPYEbir9SZe7NEsflq+
lSNYVaq9pSBj40Jx7th8wq5QJKjP9It3+U80n0XByKWCynAHyyY/znoBbqGM
2RyPWt6mDwa1hxH3fz2uFwbABWKSpuQM5HWCXYfHralUYz7ReoYFH31EO4ka
qTXp7RPD/qf3Hfb0vRDwmiRN8aF1alAHOYvCPZhr7b2hOA4JEHSgLJIsU5qm
bTZnms2NUbqUTUY8G/Ffwox0bJ4Z5FWIwBx9KyRfdl5d0ySn82xxXkJ+gFNY
dX5ff072vyS1VKVxIlVpQFAbw+5aJU5a8IOMClBqkAuOST6QfrgqAj7eQ9JK
WdLwP3yCD3lTpBEgulL4c+VZH3cNin4bdaFNLweLrERyJ+N6y1lDMORmtz7X
NySq7VjmSUTPwZnpLgD5oJxeTLO/T8i2M+NlFNYiga449HQhuOwsmfflzcAh
38I2Tys4qMYssfLjS5dcs7xPyCwxf0LhIHOPXjxa7DZbKS69oWcbFv2d1cmo
cXqJ4tUO8cXPPpTqHzHCO/65qgum4UWlHoAmDKmIQoWPD+arbK54InxQkgbj
SzPyvuwJknr6DYVDRmU3PI1YmmjcAGxbatT76oDGL4sXQ6CJEx9SESgolj+l
iMhQ5s3um8KkK0GfiGpstApF0+GUwKC66tfbC+tkVA1Vxwq1n6P9MRW127uK
pMYc2KdEmuvzkvcOSEh32lwgQSG1Gnn2/yQuDhblyDeaEfOmA0+ajKsucmaE
RlRd+vyqM62JM8qBkxExrj09vNp9aqjReefdjS4xONnJoorTWPML0gc+53hR
VrN5jtXXdBlc+6BEMGzBOUsVkcaHojTE3zE5r9HsCsNgmdVAOIfb2dWEDYBf
hFj7jHlhvL3RtfyZzeI6S+r/VmSatsqNvw9Ea0SuOLyU2FNz+d0/Ty/ub3+2
PqXVevqrP9QEPK1QShTN81R+EeI7UtUBvQjK2uWpjN81T2sYEftvaMYsl88c
ahqrC7NJc5/ccIjvfZlwogp5ARHxzgSSzk6nvLMhxULB2s0qkANGhXIYIg9t
djioL3KfwI2GLLO58GdmReIDpygj/JWZeeNL8aVjFLueOTkxI9qFeClwOW0K
0uQH3fvmrPEeLp8D6lk0alWRBKuCJdY5lj+DX6Bboqdj/FD1YoDnsoI6dkVb
acC248AokxnqGrFSHbpCjHlkWOXhvY2AWoy+/8gf9bTAUwR/h79ZgveOh97v
uK+/XIFiuFhQczQfo5vdDtGLba9FAPcNnGDF5nZ/5zyyxqS+nL4pbmlUyrZE
V5nOSsuzA4mR+5JJd+rVKwiuabKnOoNdyczLcWz1Y6nPaP1KM20H78OAO859
sGIYlfJtr4EPhZF9nGi4L8OyKBETb+ZDOzhBHZTzsT3A5WZ0igDHrAWDOdk0
IDmeYEb5sLPJQYCoSRD/ORkFzLpu0M+WixU0LypgB0+f56ps0NOzcx+nCjE8
YALlJbj6Dlx1gS9gAmw1O2tlodSPboMXmNRpE8qu7Fr2QyF6f4xh0MT9W/Hz
pP+PCvKyn3NS/wyDEUW3ta6Na2jMga9mQs67LHNaIA1f3GTySVcCX6JvVrfe
uljTffJN/yB7noyx1fv1eHuVmggnTRzalvMxNIVrAWkaTDpETL+AGS4P4wgt
CUvkfsPjh800t+bFgt5ruxIYtp9UVTie5w01+kYWwuq3ELrp/WZEEE6QL+GZ
R9q2+ODI0NSVtKjXdXSqvLIwGem8V8gtNFmMhKMEyP6JmP+zeEMdrfo/RTY8
efZj8ZxdI8UfzlkBwuWoLZh+poloV8ZQa/sqO6I4iFDu+FVQtCLTKznTbXko
/zQboOgP/l5ofI3KqYhpGPlExjdB5fsCEisyw2CE9JyiIM0qM9bleKACdZ85
3rb7Gtacmi2fEyJ7cL/bJYxVjS+WrEGIggTTCl20G8SRJsjFbX3Ne3/AULje
JUd5VfEgxk1sRkuQ1R547LNvvyY/vPUO8NplwAsbn3ED5qYuJnTmAbvTmpiH
u08HT9vb+s2uOVGEcDyefZS/KwU3PkOJ72zgbfVjZILA6TjpDQz8kSDy/TQe
1dyHPt0y1t6QkQdMxfPX9fbR6nNio41yHWiJ/yqxtvKP0tYQc+ExUJj9Jb6Y
+oo01vBs47LIBrM8kgeCWXxDf6ZyUODgN52jKYjrT++Hs71DsUVzSwGf1Zt7
QP2nJj1/vJHetu0ALXbu7fiMoWUj9VfdEBxwBo4dfFm1D5g9E4yaEk26/vKN
4bF4LS4XUsFLNHR0Y50cZj9d9UWiKjTVfh3rjDENBURj/b0Ih/AcFZJ1Z+Rw
kCLpGD9JotZuYreZUDKMkUyK5gRE8ICUlFpzXTFFNEuxrh7JPIzh8jxlPeSz
0mQS5MwXZh7lt1aKul3tQzeZWkJbOo86O71FKEyQulZInZs09mCwGEkbhLMr
9ay6KoGPj8p8prCXlUY4vkArn7/FzixADVrdlUbzBadtUxCiOEC8mSw9b+j1
kVzkZtPhtzL8rGEqrSnqSE/WG2llBaofrTnYtM/GHdm6G+Ume7Z9J8WCGvU/
3MRPoJl3Jvpf9iiagWsj8wgUhoRoQC0WT6O5paugQaSSqyjZ7URbXQ27te05
A2d18Jy5V7tDh3u3VgSoiwT9JtdSBUrgMUEkry82toLKZiIPnL8GkQ8g7dYI
ZYLh2mJ9I+X4aMkc9737B/v9L4AjYB0t66IW/OgmJy95xlcsS/RgmoLyFU9h
okJfP5f6i4ba1/nPoGJQjTPsxzBr/7Y9oNDJQ8kOdG44nMhJ9+OkcPY9wk7k
cPTBD6S6k+lHMkgmOE60Jos4b0ftcAPJhp83jX4PYZCtmhSc/0A488cY1vGG
1HO7PcUvBEXAZN35sBiYOjIRQC26QcRm0E6Nq745oG/eOPqJmOkayKyWfR/R
SDsyrr7qV3dHFVpSM6o+ASa0Uy/OufITMYKXOLP8DddRaPd0bNQ27d2eULNk
CFw29bwFSLU12gF+DH15hyoKQouLIp/l1QYchKl1QsgnhDf2ukCYyrXL7Hdi
KNd/U7WXB1QOGzwKcgsSkT9qM4liLMGij36TWHtOD1osSGl94vTHMC/F4Ky6
pEBBlJboIKh7XVkj5l9eQYIk9yb0kOL2FC61pabgSGUHYHFjdoT4Lb7ptsk3
E+nlgeAnGQsn3FSsf2/bqBUZ6iV8l8RYVeSxyo4hNfx6RhTs84FV+oDv21OQ
l/JkCBNIbriMyXQcH3PqiztzlvrAcJXrSVMxsTWFZ5hS+E5xodMDU1RTS0vr
GCkQ4bPaI4TD5QPruaUI+5sRh2DJtoNcTG2OIUkyESPQQyoh+ako2+Dz0Meb
tDJAxb9lxAJ3ElJblXNwHjbg4sAGav5roLmZreJ0eh1yn67yD1jYgGrFS0ss
Yt+fCK/2N0YS+GzTU5n4vRLDfYrrmCYAtQsWBY3qfTlPUpQhbBLRh+lMJaf0
1LYO7zYoLjzKmZrzxPLGyT4EAizxUx/cZeQm641eOWpnJlW3b8cIOINxCIXs
TThyZ4/aCPz5Lw/ti1UMEXdXvyFJ2MyYLxGwfTqbioQamf7vFGldcYt0tYce
VKnQneMjMzqrDQVo2VUnjQpuc1vVqPa+/ASR/TAOxtK0ol4eLSqLBKBeJKEJ
T28Pm9sX/00VSoTsGrfdK4T66a/rORBZRSlASdqaOiz8Uaj8oZi6EFsl/pN4
OpJaLUKeDYzOz4uL3yIGkoKFTTAZasaiomQoyKumfvkwcFQLqK95Nnt8XrYy
L4TuaJ/ufKZ0YMETYqLXLTJH/X9ai9VT8dO+OwzcoI/0zOrdc+3kTRZcdcV0
w/pLZe1dWnfubUveEGuRdxKF2NHF+8VEu4Dzo8ucBkmi1inN5IAn3tSvy76N
x2hBDIe8Eu72SPsOdEPIU1BZTeiLR1Fj0oSkskKrgWOYebVN0MqpOYI7emHC
98r0shzehxKDnBLdt/jkqNE69fX+dFYpU2QhKUyU7f+7mcn/3bIEnSZFwaVr
nTNE3nJLUN5KsedlQoZ9BLMmpledO9s2/RumZbDgHCYkQIjdydX9jTjJTX+U
vljk5ljs5c7hZy8OGQp8N2sMCRv8n2yD1VIRTQjwqjjwgQdAP9fYF7mXplCM
SGKSf4H2/ZJkfcEfjvAcYbS9tpFYngb2BvRpAFi1DRzm6Y41nwifV7E49vAY
h/qjudk910rLxv6fpzDW4Y4tLBuZvQZftEuM/1glSa8h5eFMGpDqJ04O3BZt
Qm21WoubG3a/8+NzSBlQ34we+mN/Xnxof4KorgB6JTRrZFAE8WAeFJrenacf
zdacoqMP8YVmL3VcXhUUetVH0nWAWMhraRssJqEmF3EdnwiCdjOdESxxWfIL
RSexA9+nc6wKRWSAD6Qr/vHjphcslX86hmIrDLxE7eQ60D3mEHgmXMFpOeM2
vf4Bkq9p9wG1porAyGQKmYbj1jAdIkdHY7mOySuJgnPMrBTpJu1LF4qO/83d
raY1Z8OtVeJbI0LQcNN0aUfxbqEtpXbx7+e1AJD1aVa8ofAevJvFnrDIsy33
GXw/3D1VWz7+QAKh3cTQCk7kFiwW4lxK2pUF8tQIn0UnGCdtgjRIQF1jFngh
A9A0AXKFF78rFISpu7R6awpFmAANWx/nFP0urKZLXHFawgDy607SToq+Xalg
kyT67yunFgWSwCqMkJhC/obk5gZwf3ydhl3lCecZ+rdxIKJ0OoZexuITdi3M
Krw3K9jw0UWmkvIOo1jXIxOo1Sf4VUhpU2/bb0hnq5Nie/xZm7mgYsjY5K95
kMD7UwALeKyvFm1D1yMuWnNOdffWGWmyHeb627RX1DDxsMW1Q05/qGf+I4GX
EQXph6Mr+r9fnbkfylsSczPFcD80iUhJPjnX/Og6ian/Af06Rve+rpVGwEnj
HLElbzpc5X5+imE1KGoUhqzVyKlQdf9Dq/uhbOVD/y4WXELgBrwKXcgVgtJM
x27rbNN2QcvXLPLiTxOvLlRpuAvywEKnG4HO35F6nqs60pNr/oFmmBkN7Dsm
oXRUwxVKcPdlMwabC8Pi79ZU63/qWbWxFyuyrbnkUw3cV36ewRD9eNJNkTw7
/He/TtgwE/KisAET3kAQ2RoYhiQ7VTKHDoeYvhoueNcDeNNHbSgdweZXyJz1
sg8PcRpjQ62piryjL33oVT7gcsXRGQmu+aK0VNMdb7wHud6scK1Hr7UGCTOf
StGvZpvqlOJrAC1RkiyR8EEzGCQK+z4jAjYk5PN6UCepjoAYSfWA9NhRYVew
OarT3u/GEBV73pId93J+NdbUcbV3bmPIMs0BA4FEWSt+dpKgspYsLzHS9QMM
BEH1XGsyPhSerJ1jRd2VFeWhNnZQsw98F+A1oBpX5ZJd0YdAr+t4hjdXLdqf
JD1cYq9O1n4gxYe7zsNqFWJbuP6qPwSmsPA8xi/kb1iYANgkZQWugwGjS98A
AuIF4baX2VHN1F93+7zflpWbKBDrAj6l3jjzZmG6TwJ0nHbOReYiddy8jU90
yTSPA9aFQXBjpe95lPMl5yRYnXclYML1aK61rzF+Kq8D3dTAnufUIvq+7lnD
vpghaM1CFjXbguCm7/UrzPYVIquofd41RljWHTyWySytLPzHAjztP+qDtUrK
6SxlmTY7jqBOyOA7kHApIGlDWSQpS4j8WAniRLDfd+Z+CqSSvZCmrxfuClYd
cs0tpuvw/gGzORGmuM05plfYHZBK+d4G684py6IxV+oWilxWbaM5WjIIdw7H
2RVHO3v9E1lzNrkl1JEzusnFRI/QYgQVay5Fw19n98FVmzmSwOd1WQ8ylGVQ
5traxeKz5bXXnoFz6GXfHgSpm132+IZzriqskqusxqu28IaPOFeI2OOr18l4
ms0fcmSI4ma5aHAVkgqkKg7yAjyxac6KsGj9GtfQrPKaWzK+TpmBp1Qrwguv
zGLJcjVJwEj/aGhEhfGEcO+YsDE1ZvgkTpU4X2uwHigDOioMXZVn2OxLotmi
09HY3KpwMusXzD3CJzTktIIWPXuj5vY77eSKalI3CC1jhuQHgtgswBAiYxe+
V2/qUvb/0qwpq+gqsZ5OvZSrsTHwh739QWlST5j2le1HM2a6JPq6SbEuaYt6
2/yTi508UcJme/Atk1Obo1/qZOittesuFUGpZnADKdxuhXFBWbMpCsQIkrnC
u88iHd5z8Ipm1xV1GciXobMKoOUk3OrLMWh8N9uiCsM25vhgDAeS+VB2MuLc
vylAZxVMcATp6lWXzljaIjr33GJC8KwZvoQjwW+JUuQkuwOa3VEYLBz52h41
ksOxac1WezBpPz0BiUF5ZraIDeHLoS4AONM4HBxKPcMz/8HJZtnuZkUkPc1d
eD2WfU8aStAcXYNK6QgJxcnTATWn7orVW6+R0gm/RfnX3WPqNACR2malOAce
k58NCPN6RzTotVVXatMCuwuYq8HbpNA9A6d5WopJQNTeU6Tk2VeIJcYmaDJY
dyTJzAcfd9JH7uErMLSL04Q2OGB2ya0/7EzWPqSd95Ol1WJVEWDvP7tFl1jP
G3CDcp1A6AmMJc1uFpjAKMJBgJUg1/HA+eXCSgcpmBMcbqFjGxmpUZpZjReG
IYPPoZr/VQsKAFB50CxJw+ycjPn3+aSs28EWj7xBo28XyB7uTB+66VdJqE9J
Lxz7g709/9Z923J9mn++h+8spqH97mGPQ+tBb03MLv94lz7ghia9DYVnCP6S
7KQvalyF0oVNSfKpMz0QlzyKVPGhBRpEAlXHHrV3mTfNzXHdMvtvr9UFzexh
roxdKj+T07vkQ9be+1VLAlGw5bN/ZLj7faBxGq22ze6aEmtFnyF871q8ydOy
kj9DD0qpWZ0HTx6DVu2m6NwO9QyMMdAF6+m1OQ8Z3pSQnSOIC2/T+7ZV09Yh
I9vR5C3k0qavcdCOMNreDt7WApESMHOXE03glSff+wjO7Amduk/WjTJakjOr
kmgaO8nKgu4U+DUWROGkvG0hHD0Who1YcutzbdQ+NUu8WnXRjbA+5bKOT+4R
b8TvYb2IJcle/xFWv0DV9HrHz6lUhDHRxNyMzPvMeFzzdVSAQzgqrVxbLi8+
yE4rDcuMP3cXWcCHOB9Uj5Hq5qiUXXBiFCX27t/INuTW6rNowtWgrqswPOcD
7yRbiXQHp/yNBkM/hCNjBcvBtOcq/OwP+k2zHa+Ya0E2osOg8frrx/bZBvVn
m5PpPLb6Yy/pVsxntdxMmCms4HVB5YhH890MapJqpxXaI/btlpOnKpztEcVS
Wr07fZY6X6moKfU76fANf23ImbfTKyPWVh/2RhoZ+RO+7wPrYiPJyZNqDNVJ
A6vFTJMvxsuRld0GirWVfPoAUjoHKEm0aSXgWnn4R7rKu88spsmkAjbGQNea
DzzRO6mDAcncqaImo/5+U3h1kcGc+lklxtEJIyTfwCPaFsT9TPAN+NNvQBhg
aZSh8jinjQl/tHBjYR8QMjqXCdI6tfrzTWBHNC417daWvIVxtHmGUtj3AapY
dUPeIyEM/n4FGkgxoWHDMbrAe6VRn2pmSIkljTQSEGq1++9NFFYJvlYHTzIl
gFX3yl602Q8IuDTC5WeLrPxzHOntShbPB+fOshfE1wzW0dkvKpi4QT/O+Cja
NRiQBuu3kedQsGnrQ2wsx9C4U3m4BS4IlATwmdhq/wMUevfKp31U+w0tqqbj
wFAZt/yKhLnMSVhBnwy9KjZURdiFUpfTFE8pe6yirG/kY/qMvMer6oUPxHnT
wKxpNAHHoef/BcgUjto+tqM8xJfWSxhUJHUzlMf9A0S3oQrtf9xxSE74enmd
5VcZXWA2jn81tUi/RMvN1w4GPO+jLCXk7mjB0zGnGWtFOkGbEpuWvwxBba45
yv5iN9M1la8H6gP3+GZbIeZrgRSywQU/qmWijun22Q7kVDFXd8Og9GfyeBg7
5KOcIEBWBz/WGyJNEvXB4jQNPgzqJcE8a55ZcTk9KYub2bI+ehEACcke75Fj
yIeMmGNg83+l/URa1Kv5MrZBPWKd24B2NPBO7C5OsuPPIxtkkORFbp69CoLB
CznLOoifCVduwy6FIPDRSLHNnx879tTC42+SI5ARhZpB+fsbQWwhAb4UvBV9
hB33UdMySC7AQqdfAL4NN0fSzf2QSUjMQHuRXb/ttzKBFVcBQDZby73ZtYED
tAGrZv0uTKobcz5iMj55TkRsiXPl1CIr3fvnlQQUfVU91Xwpm/e0uhYNxTlU
ihnYAneo19LEgKwLIS6mIzxhAmVEypNeBGFq+I9oaAlxHo9nHkMS7RO3GRXN
owk2CrxroTlJyUXG1sLR1O8C8I0wQ6bdjG0uGHZyL2yb1Qnj88rphDp8ntq9
j9laBwLd684wEOMB8zaWhFqQx4NFXOkpgtaX4ogqwqsTA4El8gpEVW06Akfg
ab8rCRM5DAJSpImUV+1OsunZ26M41sQF0/41WW7yN8WjUihV7hVNyfNhVfJq
xdFJpXd+AGdeC/reAU/dg9PQh7xRyMCrmllQ1ekPo8lfm1JvJoqm5JPQP00z
m54JjLbN6p4g9EZh9en8f0Y6MWDVXdrtQuuZvTxBWJf8KhFS2AYSS7fXI9zc
WVGlm9+gOTUkG3AC+oyDBvruqsJFd3QmQLvrJVuBvGkmv4SvHbgwW4VRzcM2
5mNlziD8PnTdRhAgEO6P95UVe5LVQrYydLj6DskfFrCruuqGtlY32SH2VOnO
zD1kmjMxYtfcplTTUjTx3gPcml6R6WGqWBBVNEJ7Yoji7g6dFCU9qLWuypLC
vZckEJUGoZDII4NHkkX1wph2PxEQXe1n+FZdJiBGn6+OVNLImXhVjbC+V8dX
jeNfGQHnG1AWk3c8UQVHN3UvYsl3zpjCAhG3daz+2LXGi0C3sWSB1nU7ChtR
lk3wBdFqWwZmUHyTExDhTl2L1BzyK08eqJIpkrbJMCr0ds+Pv6MA53sQ2DQZ
F4zGD57GmIxw9sNOti0A0ZyeKMovUx7Zf5Y6pSoDwEDyzzNr9ZzXKUNdPuOi
WKMHMUZky7Gs6bMwNODcamWxX74z3K9Kl9ey43Fp6kp/gClHpUIXDgEuaz63
Wv+NcEP1ROG3lwL3eqE4UOkAcLcRNW3DrCfYWjnq4fMsPJbe/lOt2lHLmdi3
TAb6Sa4uwbmHJ7iX9dcfsQSroy87S3RvYpkdS8iEAEhza/eivEl7uoCqFtEc
YSNfGtPSsfeyn/MS+zdevR85A/4y8El/6zMmes60e5cGfnwkoqbAjtZyA/Yh
n9riH/ipJS/lD1ZbHfCJl9y9XkyCV9DDOp3zQe4eZE0yvDra8B0OPB1EfOBE
KRg4pn5jN04aEPT5bl/u73RZa6H+3HKskMHwOhvl8Rv6pi4wae5LKINSYVSj
ED2M7ZC6Hqzwceog6FRgWAwOxC4iHxTSBH5d8TFM7PTKKYy4DSo9WEqCilDj
AVzW/Ru9+wdEc+I4EtY2wQaDpkIJbfGLuKxlVsFG4QpaZyznYttEcq8MLAAs
kv/pnMZckAHdcCTzjD2xewXiRtw25fsCOZghelIZJ/XHfxY0EtmQ7pJSe41O
4niWVC2RR5eEVGlVpKkna2eYn9Fs6zMZw/Vay5/tsfLkWB1vddQQ/PDenDTt
CEbWvy+gslutqg3/0Z1490gbb9Hg1d5lc21e4+xEMnjh26g75cLsQ3hiTcux
30v1CT715jyciq5tH9EMG8fAs7mbq8gvdAN7OIlQzb77GqtYLALEjkcKefSE
jSYren8DKHjWZkCUq4+6/DtmRx0wWhshz14Vem7JRU6vVgE6CMYYjYd1cXZB
ay5s3UtpfXs6iR+7mVQ9H5fJKfo/eV6xlq+wTcr4X4wpKPJNJxauLLMYJCvN
aDgYaOzl1ZCBNd8HulsBQ2Qi7EWF0m76qlbtq5vxOD+byoZfC744bSd7KBC/
t3VvgHlGphAEco17ls7qw0Sl2B0j75gHVDXU5t6ieEqJblBM3GqLrJ5udVkY
ovxIfJPKYOgRMYHUXgbLToGevVg8gIAiUMWBt857NPEZHAg3HtB9EolyEP/W
eskWm+cYg5k6vmIdOEC+atr6lQ11g1NwXwUEPUtH6JsF+t5P5WgxFq0hzudX
ZBHu8jIFCrE0MKhPX54oTAoIiU6VVT6JYmniNM8B9G4nANrgC6dMJbolLvwe
FzMzm+bVnDxFhjGWTiAo/CTSdLNLExUP4NxCMXrWqJ9+li9AoclK7iRB/qQn
8yT1x0ccB/XK2CfVhPnWZsyt4egi0NsA8fhWHSww3VkupV6Q9D6fKKR4C+vb
BW9CqwyObTWOndgeSX8HukEJUxAirI3cMPHGFQkYmE+zIi0bGfF1fcpfWg6j
PPhsLYsfiHxP9KJTnbzBjQ7b9F7vNBE7wzSNQG4oyGUL+VG6d5g6AFFfi59g
iLU/U7LVTRhABNQs4BQDINB2RFxehl1RKhu03sjbM0p+5jRlE3TQ6BMwAl64
qzhgtzaFtFqpC8MeXW5/dJD3BWPF8msPMSvbA4JGSLhe7367UQ5CU2OQGNP8
B8L+0NeJz3sG3f1LlugRzzUbgzlcSYzo/tnpHJZ2AtcdHL89PN1wArpSpVMx
+Emu56DQdOuDRJpFPcBiVMbEEcrtB+rzqrqW6it2PfkxOkAl28RVUbUIXXmB
58T+YBGkFJx2VDKA9dB96udQNI0S3a/bxzfIP+Z7nOIvD3lP5u7XjoclL4GT
R4BC+gLcIFgNOZpI5EKEHzC1+Cdfj/TCBSdyfXDfL15zKVsWVGHEQKLyuwjp
6qwQQNYdx1kcVI16y9FUffkn1yZsHAvE0MSPQVJ4ikKTwtZXh7dd7Jxg/tlK
PBhNaKVAQgl1DU+4FPI23eQP2dJafUvXecLDBySek9K6Ir/iHLfMsgRlD9i8
BzbthtgJpp4xgy/e016YtUnc4IeGc0NCaXv8cWqD6loCRPAeXYceUjYtzgXJ
h3XF3aHtPe1TCuLIA8wCQaxYpjn7jRU/XPhIxg0/YiPYUEKhHR0JRjy1PQ7V
mQCwrc6thxuk7Quq1WrcHgqjaGZ3ZOiUx0R+F0LPJeRmE+8+3R/ONUVTgbz1
b3VYY930+plVCJuk1qJ/knu6dKngZx3/l7bf3OaRhOv88UvhJw2j+hUIoUTW
qUBj81Xopkxd7f0T/33ITCJB/SBhW8qEd9s688NnmA9Vxh5ZaaXzHxd5bG6q
VPqSqwl2rajvuEqCN3RknpyCUCO7j40N4mOpGEJL51SKMARGKMDX7G6OViE7
hkY18iTf3jwpMT3t7Vdru1RDLl41yGOpHopYE9OLK+iacEZXyPHfgrnmtGyR
eKXJuYli8Rox9PskOMICg2G8FTpnpjc8oGY7nEv1xP3VYLlfXluR7HLA8p63
H3VpmMBEo9vHtCz6GKAhxJOKNCclsXepnmUlFsgIrLbxr+kBHw2gzzk0PIZ2
Oseq5xgW6+QYRbbr6GNyrl4fzVdemfYJzoPBHh/Yf5a3Rru8vX1s6cafd1kp
4NdpgBIGcYyI+V73xJwBHiKpCD7BA3XH+So478te76cEHQbhH4lULiizUDEx
7jCQRYWnc1nXnej0pJhWvrlsGAxR58Rmzd8FMV1bysKV/Rmw7F+JGbEYsZ2p
Lt1ORnxGHoBcFCucjOAK5BOZHUMpqa5Mmd66+9aRG+5xyh8L7ACHQgnTZuZt
tg2B3MfIU/qPHCYQeFKJcoAZGTmG9OxqlIaVJwmOCLD6zUygAD152FgNK4eZ
HxrwzwlES0RM2rrpF5gKmGEVTu6Ol7ml+UJ0KDZOqScPoZaWkUYtm4VXf1yE
L++mQSSvxTti4wrDxb6IZEtt2HvSNtZvJc/G6h5WQSH/m7coF3oxm2ZSmmaa
02CwZWDalymVmKHlv8odx0v2pbXh0iwlXgTwBbFzGNyc3wTcTHn6PkHTCb/v
TJJJG60LGy5u5qqiIBpa2j4KiWC2j8uP7ZRynkbtZgcKFWKYluLCqHhY9ynh
8CAs1IdwebRDPvbp9o0Y9eEE5Mv7/VetPWwhdCeR/jLODqeHoKjPGoB/H5oQ
3Vrv1QCn14+evIKMQW45vGTEbIgImd7kkPnQl0fCMOtfBf3zIqO9dUo8gb8p
I55CRhBPgfG8QulH5Q47Ry5J/4ceQhwopV5Tqt0Yf98R8sAdVxVq73SCjHqE
+OZQfOpU1KEw9OKsQYjH6FPfelHpPObSrdu3W3sbvCnJND3+jQd4NWHzeL3/
K4gk1C0pYgQBCueMOAix1yu/5xz/TaG4pkUxiOcP+UDrZHG2bpJC5uHE9lar
K2JJES6JBs/mHZzppNvdjN38l1T1GQkiI+tQ6yvqQuhBY0vppKMkCYYrOouQ
JTBqwu7bATVd43OCZiLcz5IRw4/5Z321qe9AWtKTBZca+6U0jj0Hl0IIzkTy
l/7Ito25bOsROzdPz201v8y1BfVtAAgxiyOgo7Hqs2IbKwOXRdzMnWc//jnf
r3TfwX9Mq8o0clpF9D1JwlMY/JDXJgTqrGrmkAj5omP0fulCj/okut0X5Wur
+aIp920R0RJnAO1j8Q7cBiUBKXmZnb0yi57YJHS9xFp6klmnelT77Q6/WysW
T9KgMFEOe4Q3brzsOKFIVu7zvhpkh82ZMjJeKaDypvYzTCn14LxTiInr8vua
LSJco9s+E1q3nMgYCy8VghmI9DbHo7gL629LDej1kCPxueZ7m3s8sTiXfedI
cxcKK4Ah/yx5kMXiobmq9O9QrpvFjnfMnSSPJ4IUDqu4QFoTu5yPmaDDyqDz
cOylO+ySZ162weW/EsGhF6AO5fnLZPhXnCfP4YBdiKpoo6z2PgQ+lbMDlqJ1
9Z2sqn+DM+lDzLfHv6L2wsH+CdqhUsxGltbMljW+sXXKTc2pXArvcvWmWIg6
2AuwUn3vXuv7rZj+3UBXfwrJLz92zyYO5la6wrmyh10myXxxRE/HskqbAfHf
yl+YURidCZ/9m7FhOPZ0oLKoSuR/zx78xky+G4tA+iGmsDS8pBC8JzVz01+y
8hdLoJqtlgaZ3aQotESwBc+ofXuMmr+IKCCjWdXrdgfEUjNhVt07hH4+gxfD
ThjFyMK/tZdBYQykQRsHgLDXSgpAxtY5TDbf3HYkqUlNLcodXlqABPgjGHiL
REizScHA6IVSeJG95N0/nc0srl8/I02gLj0YV9BDl+j41m+1ioWwChPY5W1c
et+HAVXJ4An1Re6QsGRek98JGAYVxEZTgzmW0gT94TQ4jesEpYfvRE/Qv6y6
kUT/NzfShWqVC4pPt7XWMW5j3dc23TGunn8blK+yGdFAwF53NA/JKvkmwWS6
EvUh+WtF3//8qUtPwfMcA2ULYXUK7Q9QgdzSoYBv6ceW+w61bPm4IArLpJrT
GLhUWN/BxOeB+bIi/XPsoUPMVaF22/lRcXH1v+h2ReDcYgEuHVOCa27OLTtE
ul1YOnvAtxg4fklX0r56XgMPbkpXGHiK4zJaUlRh4a30u5N6CzsZZHnnE/DS
SrgjzyDky6QJfG62uIUhd90O9mWYmoXalk3A6VJFqvckmqH1aHS0bazao6ck
iLMsJxPjfzgiI9JBqxOaTkSsEdeB0EkBYuyAjokdQTryh1ZU+SV5eHb2zFZu
hEEOGv49QrX2eEVP5PHpQMmA8Vv0rBJCnApRPxq9NPJDP+OYyNRWQj8O1kGc
lkfshpOadWu4i3jIZsszU5XZ3QSKOm1Vt4JGgs8HRutjXGtrfWd1xOZHimct
Q5mQi2Rz8NAlC5vV50jtDhDT3vDFjvJOVQf+/BvVED3tOI9m1qP8HCHzFbV3
f1fIWAWToe6a1lpncxhSzIQEp4H0YM/9t7BKBb0Mf9y9Zw9Y7CLl/WLUIzCh
7XBd5gu4C9SMKlY6Pvnlh/l1iaNUA/n4u3XQ6ynQghpXTpNjrdZhBUKkuVWX
wqgkRvIM4mVMamnNvucYcI2AEJFYh0uWbnkhK5yG4LYRo2nU4uop5/kDwa2j
e38wZ4oSv9snzbPaHp7zwm8/8OZvybRojFDJcLy1Y11Wud8pDIfrfSfimiFU
qLC/CeZDBR6csgEU2jmM1gR1YWSgtDWkK6Mm1iiMvQvxMzygEHhvxQYlcNLO
6eo2B2KGDnXt+m1Rl67+QxfRAHmAMMSeRigMb0XFD+xKNLYzWebrwoB/fMme
XEgX6JP+Tj7g4krn17qV/0EssirYdF1m5wSK6SVyVYn7TcsDKwr2usq1UROv
u4gtIhBmd9k5kivaorTb9VGmxZHJYyXtFTaTAtR3niICdCk2YrmUrUlAqji5
O6FBNb1rZQQ95BrbP8pgRbyjKGB9Ld+Lh2qK7PXfCFi5a/JmkwRjn8YDgDbo
EXtyjQSC9S2ovlidXjvhsWqCi5JRFs9auwSarkHgwvdcMTSrK952lDN0jn73
D5cFiDuWoFnNQd+qE9IOFrW/p5r9rbxrr4JSj86aZB79WSuMocs6FuulyqNS
0tlPefNAaoC+OyARnXbItoCfd2I1Z/uMEJeRSbEAUIYu4GLM7q4AC3KOqo3V
JF4ExaNm9qx4w9SuUmueJ4ppBN20hXGbYR0vUN2iHNnrP3BtAU2kQns1oZAD
VaASmfWdHK+hSDMysDDD7uphyf47jbLoWqjmSzSUv+uFkJdYwt3go2C8KnYu
IzYbJbSGP0QnonfrSMVZI2rzkbrVCPzzO4loGOAv6geak103xFwtZ4A/X0q2
Jobkn5cJ8vbSGoo3gtLbpKLdTB3zQYv4DKot3zmpGQCZPrq0aIBi9quwSqGm
qMYrHR55n3mHdGv2KoZ77tCg7yaQ0sFXTQ0N0xK3uc2OPQax0whTskY7L7lp
30S2ekifMahuGMKkz74rYuRLU0xMNmOfKIjggr7t1Dm3z/Z78/HdjnhCRhkA
rFsZ4pScQhEHWhIs22res+Kgf1nHFyqVT/Q/239y9HEMaOfpZftJ5YY4r61x
HVZCwzS9+It462pdSeQIFBDpsbwl8wPEcp56njoqeLZMM1nHsXProWx2pEGG
UNvEi58xxvhINjgB3uPymjNLRoU0fRP8sSUYUT9e+TbxnbQ1IMmj0zkQrTtU
YM/hdpzGtnYGIKNpD0Ffi1eO0Bc8cWBtkL0+9GF/aFTUi8odUal4jtM4/6HX
+gPOcydFfx9wzG2+iacidW4WSDZCgv7/JCE8CvN7FWv9ZKiJXobrW96DCchJ
3JuF+3MDwzObC1Euril6rQxcmGGC64M4harVA+sF8g9wcGb/Sn9PEWJw13jU
8HnyR6+CuaedQizLIqhSf4z8nOYbxhFSayioUJXwUJTKQLFPU1Tsj+uXIo3q
qTTWAbW6aNn0+SZ57lv0EIqOjrO0P8su41w4V+TxRAdFBKSbcufyRJLkHv88
HLnOKOvfhpvtnmIHP+T5jiijT9MQkR2K0xMS845qj9cwEPBWuMEYun9I9wwq
Vaw72w1cWnwfVTJXYO83E52mtnIY/QeMQQKGpx6Q6X/vmGzbhWzyANbBs+xw
8ry/Ix0Phpbt/PQMcZgjtHgxtVw8rERDrwB+tZp36glW5gzmVXDOY2rr7c8E
oJaw+NFjp78SZ1l+zerkLtPKU4lWyWThaH5/eeFXUTqs12zW36CC3lPkH6sa
ryuGUBMMw4wq8uYWxgNotDLvwlSvpefSPrWF+cCXhavA7LxwsrQ0pfzYyRZg
nLwTjxgvKMxmt2EFgG4tAgyXwpPcz6/NPm/odp9RiYwskwtG09rj2M0JV2tx
4pT5QJCY2mxRjIpOasOMenF4shnO7lfJsTeEjyqkaQu/lp8ZBy21ngk/xqB9
5oxMypLu1LLsrsEkHEDq9x/UQ1O1sEsY1kjjHSO6R9nLtiX4YPQ0o0464pf3
DW/GzEphSX/DCzA5H1mxIRuGQq4YsycttPpXfDpSLIwOkV2QxCxfMYGd1m32
fUBE76JSfmrT8X6BmwOMSUzwNyiuGDhtJFudNXtULrUyPq01AJz0fwBT1MqW
HsxUp1R3KlLrKwCv/POL2AnLz79wsSzhRcIyBieKaqrY3KGheHcpzUsAOrcg
5azExw6YYd6TzePY3pNt61AiizftiU4HGRBAD4E3bttp+rvNotagJhSX25dK
9v4UV8+3slc2Nz2Ps7BHcpo9YpvWaRm7vV0X5DFxYQT0QRXCBqevRl30kBRM
i63sSN+tOfRUsupJoCcoML/Vj41ibTKOb9nKul8k8bk8ERqNlPPheGFX+64W
Fjc26DaqhJY9DJaf8cYQpObDEPgUK2iNnkU5OMdbfupFuDwJbX1S7FYU4n+/
OE6GIdobZONVlqDhiKkViGsedHezW9gGRdcqkzhgbpmzJoOkq8AoM3CGCSgw
pQoT39KxTTmrhzjBY/P3KUa2f1x5eRCOB3skdwH1YL7eoWo2EdAo/ey1PPtd
VaOS8qlDfuxAqWduZ2l3wc4T23MeQz3jtdZKRN0Qh8anOxedSwMYGp4w1NxC
IkXWEsA9NPLVJ4x4b60npoFa1/PSf0Nfrdd+EMt2nkBmxfNpsDBFBlBHnGZL
SjMe+z0vELRSGupbGPdE7IcG/aEuDfdHYzomP0l8IyOcbEW4W6e4fWjxyHGw
TcW9/RcusCGg1RFOa+UrSgRZlMSLPjVfEAEyV9wmXiCf83APVLpxLEJ1Ld+W
fVZR1Y8wH26qY+AzdylqeCp4f0s4QJk7sPCcHOkLxABU43xc+jTGpjW97nUO
q4acQsjuCULA890yNsbWOc8SbDjOJ/UUoewqa2PswsG7+SqAmt+mu1BMB6Bn
hEe4i8WFoZb+/4oQIvNBs6m05ys49m8x9aB2anOQrRvKcECCavgO1BnsDtIb
L1C2k2cyGwFxhoO4j2jN/yvvoxfOxFWRUAt/CFSdQCTdGALDM/I+8iK7KnL4
4RyIc5ZFEZtKa3bY3VlGoLZSRR8Q4078zqyc7f+HKciqlcs8ze+VRzosXwC7
MQpecp/jLSY2UfWVFF/Inz9LopjKwhlh0hnMMhoUJMg7jVj8Kkc+LRxmdyt5
aGl6U0Vg+uZPo5jjFqnZGED/vvrfvKuhELHq/iQuMqSkc6WBPvHmSqK6d0j6
0gumAlDiX1Uzz4By7JmOxQvb1QxTvvUyOLc7xgF2RvnkbkoahK7swmx/zt2c
vxGEVg5Mq6fVq6tiDXQFNN06iTQi5qV8cm/+H7sVjK9LZdbYUZ68snUr7pQJ
s0649Ht4yFVQhOdxmC+4IDxMLUJbRvQONUGqtVDACAVhReLORoyiwQML/Oub
DJofaSP8+dICTdOoH4bD6z8VcNfWVEpqhnclPJ379rjqOVwCDonEL0/jcSMf
QVAdNTaUQHlFDNTldCfZAo41uwYNLoPGBUE7d6m0YYGl0lJRrHn4XC0oaIp4
/aNktGu+0800TV3iOG0BTcWGMxLXVVYfO3GlcNqT2rXf39ub08pQEhbJPt8T
UtKl8jDAzUpL5Xyhl9kBh07asXMkPd2NfpTZsLgYfC1A8Vkig7ho5eGo7Ynk
kA6w57IpfhvXoPUwsKsWRHY+bmlFzOi+4TZtKl6ecHO8+02dJAXSwxZIhkIw
umlUoX9X3W1Xm/ABm4xl0WWCyx32oXukzRdleePVmiu4k8+PhIWF34b+vSJA
g43upIvVkuOgNL2hMbLLQ/7uqGFgklQbUkBJwYENpRYWBaL2xi3DH+KVFkDQ
ik3fo9kR9QpuyH9xPzXAycbGbOFgDfnRykUX5JAcTq54FAdBcZ0IwI6XVMkV
oIAd2ReRa8Z4qIaOXxb1FWGMUgyLYvvonbRFdy3Tyhzir8VCC+Q7Ndl++YOK
3u1gHTIMiQ1q5yStk4I9q1FWzQoQg40KHmoJc7UUHOJuel9PxFqQRSDhvqWC
tbIV41ey5YXH36/K4upyYfZXmn2vSWCZ9J0silheBBP8rJ+9HTmKmH4IhzKh
r6H4HUFvAcPwwpMmrYIrYZ9sP/HM0z2Z8JbrX83HwRFzhGtjXEq5KNKLOqxk
L6oXkjmME+i+LtuM5XDY4GsxAB88eM7EKacjz5tIvUDTb1ERUncg8HVbQpOB
8XP+Uh2O/+2nPVhQjOJM8g+rtkkqbAqHWA01gXhKeSUHJVLL6uScC3g0ROMX
e38RXc91/RApPVLaQQTGd65qv+w+MZK3KV9gP2A4+k9kI5phZ8Z6AyvFNgXV
NTFLzeUqfwOGCqaO/UGLadO1YA1lttLjlUgf79hwRT7KJUwKhFSpqjj/Ycuo
dm2avi0kop/k/rvUnCQPAno02u2qb6wFRCN/wiwjegId3JVTOlYrFgpH5OT3
b0YOXN4G2Mnfk+3e+k53xC2x+SmD+z2c5Hq90wWC2O2BbmJ8az9xysQ6uFPS
J9yOp+ZWSpLfh5Y2/wB5DmyDfLybK6gMuxqIzQIyaik2GBvf+7xMSOxV2JQg
D4IGQDT5Sq5kgqeJd7H6wmrwAzAfqT9eSCpjm7x2q7zSJdfuW3e8MG9HN0H5
68m50KEktNbsqHAlBKdVxEtYGSIHZ4Z/YKNDzIfRtnoRU1SzbsR3FGHlXv3u
K6lblilk08/zUv99g7eA9Xn1vwLSG2iJMhwjEN8s2gy2qckLX7E0k52SrJVT
lKTMwicPGP2m5zJNOLrJRjiA+lxCrNrAO1IzKILMfaYF0R3ZTNYh9bnPHffr
o9bqMFKOYMI6N299lOhmhT9a8ZACjUzpPpcGrzSmsk1GTloru23qXE45+Zg7
tWdatY/1RrZFi+pcmjQK757XU4QXHBu8sV++YEuAryYeIjjybqnCLTUx6WN4
zoqxfn6kGUaTBoeBX2s8VnNl1gSCPoq5Z/4BxvEv+8t2mt/3RqBFmE0fUEO0
5c2OSY3ljW0o863SZs0k/vPYd/z2e4ay9NqnkWRA1obmSXYSbLT8zYLyPfE3
dHfylt7lnYx2bt1xkOPzlHlQwh7pkSgKzU7zaXygjrs4vv7gRk6nImydf1Tw
tbmZiY2A23rn368YA1NhPSr1DPub4pmwhpsFWu2WL67QgqLgf+M0dLHiljBA
mBlmetoMsxoPplRjn+G5TzwOIf6LOLGyFCccmHE0rYfU2hurH+4jv7K/DOFb
mWy3mI9LYZD9qQxj3/ji5q94G/NsmBz3Lrvq5KhJn4T2scGMJOOsQ6kyejKW
To/ypXQMZ9muEn9g6tDyThceVXZcnLL6fv+CAdOeqFlUYGkvKhyvjdXC/51G
4n7U0K1TRz08fj/mvsxp8yGaze5mwbYEFS4mh+JATPVlMbSuWCKyWh6SvT21
MTIAtRCGPxpyUB5bfphWjIrOE+6AIl4LXt/HBLDvkiyu28qQM4xmbcSBewcV
D9ZG28lBTMmw/p7mI4FTeb6TuMmQ0UA8NOsU7SyI2G2S8bNuto+F48Oz92Pj
DbArTpCfunLdiWcdMOOfVbU8jzvWXyZgi1FIjPOMbqT9HgtHEk8A4lqk4Pk8
XVoIFC1sEhhaXzhsbME0v8n1wIca2g4f/KugqoG2/Syx0oT0WeJT5gNKwE9K
/LPAQ9nIkGu9cOu4kd/YnL0tj2DPpoTnM1N9d5nzJ0kioEZ97uhs4Xih3rOj
Ib21RVUYKIJPdG5VIqt8WIROQYOtbjtFZPIj5CmjYxlXQXUr+2vne/Esh/oo
/L90k9paEnQaHxWgYLBUYWu4AtOH66WFrELGkgo7JtBx+3bhY/Hrgl5pEls8
f8rLlQ9OzU2rAo6VaNPb8nbsCOy414hqjlTmLzYrtFaio5+1YkGL1l2BKT8i
R+MduUyG8EYzYyI75TEAp9FvyiGa5Ra19y9XOfK9+brqUXsCOc9+ElbugR8A
QKLdA4NxtHTMKw3E37r9L6C3Hx4cWwtDpq4cnLBZwQphNj4BxxuVJaRnB9ib
+T/6jXPCXD5G2OfRM635gR4P+uMtHuF3FugXCD5gBqqcEDPz/MADXHJ6iGgY
cbCzfiuZiQmrF7ftWQTlo/U0dPWIPpKWXKF8vb0Bxr6Z+q3hLFYIyU+hnI8H
1ENc7g1g6BRtE2fiepfbqohLJ9X4WNKWPknNaM0dZwqL9JvXLBkfM1yq6Qxu
SRleNdkC7kZKKh+zzb7Ccl03vgl8gkeCyCmxwwAst/VULLGnBnJrgEA09WGb
qYqFXxzfqlN+NdrYAiOhRTdCoHJND6G4i2U26Evw82JHI83Mzv8PQYv81/QO
GL0YxdluqYvvOt3CriOQteg3+Tud+WnQr5gQbPc2WjRLEtXJOw000R7/ZgAa
1e03CIs/+aKXr6YP3Zm0wRN2mJxj7UyBXAgjIzdlk04tmS7nM5C2uiCyBRKH
v8lNQP3UCmbgWxL+8NAqQqzv9CF3NKuQoDfSXZKsKQ9+t6Uy8kP89I7P6rTf
s+Av3G44+WwguQzmj6W9Ji26vDnYNFbyhqv1gWJ/3V1ZAujzVZEaApSUfzE/
Ao+TolODUQF/GfNPUXSPWTow+T5ihKuksJdSzckZQHRChya0PvkoZi2CaeSU
etAzkw6IIol5Bt8/yGTdgL1b2DEtl8BeNSqzNyKO2kmAbXApQH/BZ18usKK8
qZecezOd8giXusa0JKOx5GHxlOX1xPKA+t4slfDMJB/fJS2NvrwKeloEK5c8
3djvx8qm542vKKHYSuMTL7Jdr/CFiLe3RcwHtak0lptvUYkBqC6rxI1evv78
eEvOny0Z3prURHEiNfxbCG5YB9QgZ2EuJS9Gz++ySBHuoL4FfzkCiK/U6QXZ
J3VBUgy64gTaFSOJnDhlTzKo86UkZgHOfTLY+pg2K8BYZkM3JtkMc9Ox94Rq
E3/7adQfmJqEgIFvLyivGh+O/YME5RwrqIsG4c6MAfPEZ1tMWWePfdYY35/Z
zrxdfVKQlzGOIHtK5Tm1sVrqeifp5LUVwb2PQagraHJxVQSUJcrYj5Au4yRR
9BVUhAZ9Fwag+o5751/v6Y1UAXB0NFl1MGS+Zf0w+mIL4wU8dkodGp4ubD1d
4a+4/z4umkRy168KTK5XzfnTKap6qb+ZNy22MS7RXyVwyZ664qQLEA4NXIeM
PzhwF7y2SkjrY1r2/0wp0l7aa2SKEwTcIEL75FeAu9nMh23hDYVMLjtLxg8q
VfgWHmMKZb/1xLBV04oOTfH1ssfmImO4fOqNGf+tFzE97JUysXzwOono2rIr
d4uTcUy/tbCcLGnqisapXu8oZ7tOx4B9GMquU8Ap7nndOicVBkxju44iVEHV
G0RpsHNdTIxuzvFy3M0G/nrxQQdB69iHmVPHXYhBGpd1s2j0nXCMVRJWqvRX
qZ6Xt9WfNDEGDSD2PGjKlAYF8CZZHd8tbz5AXWfnglINx4kolxfJ76kIKsK+
mbpvTKbUxoZpRzFZAMXb2IgMkGv7hTF6tt5hoqa18e3ppOn2DGKib9gFlmUP
0jRm9hpMc4Ecu7Xyx0jJT0aUq2FNE41i7ly1oyE3StQSvdQWhc7fyrlf9oYe
nFdHrf6hov3ZaXkwU/RN8oh9xYwivmWlMvouJ2gpnDKwqjTf9lDOWq1a/PVd
nwTsYgPH26Qsblzo7YxrfIdtx8eaGOHlzlB9Pts3VMxSgjz1pf4CZcWIBpq7
yLms9TdS2yosXEJNHa0VE3+z3GiViRmlmg7DEitVxYP7I/eHzYEWpqYCq74y
sRNCznQX+jWv6l0QLCq5ZB5+2Aw9nA39zmY71pXxkZsZOgdqdC/7mXc4kMc+
cVHsBj6YSq6Mg7rOe8YoQFmFyRvC5VlhGsga54Ahp5EwCSiHOW+NUHSEVKQH
djGP6uAKTUnmweR6/lNGtdq88ts1Fff3N11EKzpuQdq5s72AaTUGXs0u+iZB
MM0XuyGTLQlyWA78mqdEoBJ/HJzyu45sW5x2ZXEH5w6IQusR3VGpyRVzeqt7
d7LvrlCzCL8GOU6EWNgLUT8dVGlh5i/PhdWRbQH9nC9KVVX30C87YiU3Zpkm
u21Re1DS0LxSepsaTL/tHYw46Onho4kx/RKZ+XWY1pgju/sGTnv/3ucLWxLX
MGAtOYa6dZlapp590GeRGSGwDnUsJ5ewEJhFVEw040rvsj9r6o5KCNtxbfub
19WPY//AG3mIOFfkNu313gzTKIFcTbbsuu4ZTJ0k+WY6gbRnVhUjXk/oOFTq
3nJToPS7YempN7oRa6Gp6aVDEXcg2b7wrqq0ZTlLUvIGvzGPlwn2sCP4Eikg
iYzqGhVauAbseh6Rl7kJI/2JerLnC8N3Pofr9Ebqhp5/UwESoHj0CH+FbFWo
yMpfIA4H1y57xiY9I4kxoi3lTRiOVSwRtnMHiuuhSwV07fO7OFC5pXbnF6ql
idarPzncKIN33LiyouGLWj9P2ljOHzK/EAkWHP2ZdHHEf9WsIBJybVnCBM0t
4TAJEE7J8PDdFEhAlLC2CAlR7re98/tpf6fzJvnPK51/nSCW5nbs6HBri6xv
4JBfgcgRK3uqiBBJe/98lyNE6YRgX7IkkthzVsH95mWXChpWj1UFlhpQvevg
bmKG+jJSfQo/5+R6aoo4oeJCyGGoec2Gc7xbAjTr3AqVoMJ5+SYLi0WrKDiP
L839aRKEBGGTf2kFwvqdP8JhD5rFge2j7qqAO+4mwfx6RGIVIN9lldVhuWrF
neF2GcdW89gjqhGjryg68XxMcUGY7HoFBoMThB79TuKvWI+8bO6vV+q2J8ST
rpKrOvX1U3BCuhs6sfE5F7LNceP4Uj/8sqtOLtOS1nfkmSGz5K9K3T6CTZVA
KXXizmKQzqU7psOvXv1UxpFneFoPwU/ofB+O2Zb2Cu5EUcjDiBe1SMr/gF0h
8avc17C9u1LROnTJZkZ5BX21aocC1B3nNzuj/gUFWfbew6I0BxDjLcV0MvFG
YDGNGTXjKLiaivAltYstvgN0m6sYtgF49jGZLXNS8VT2hsJeQojc9/LAqgnd
yxzZFrLf1f2UJlMu1wJCWZZzN83lvutv0FQZnwAifPTgbcFsZVGkNTuJN5Fd
MkEt3N2l7Lh5x4DXYBUOfDsvcF2LYGBwQ/RLhu4YhkqpK2JdQLwy9X8ciYrJ
CICu3HqgGA1Qu3R1rSYM78u9rjcGtlGVO1DVv8XAF0AgVwmJ8ZhFph3h2hSV
C3cGWST9YV+H4iVfcloq1jeyWLMCb1IDPcOGWX5DcWI+QavwXNRjax3IZPBx
xsxqsz6yxYTuSrt1XfG3CWKbdvVPXIaTL/d7D6Hgox/Zi21qWh9Dtohsuw2H
MZtW9T7ti+p8mgZCPypay1CIBUCeu+P1GJPIHrUKC48yIrAQnVqrJlF3QwSb
+wIfTbqNamopJCGMm6jFAyTzei+4S/ySzU1xgvE9J00Wyvw1ck+gS63FDEkx
P9nqFHqKeqZVA4RhafXmpGw98XRsy5GEPVuIc9jHSygXSiKC/DAlWMpa79Fi
tss/xZ+T0zpnYJ12v0XKIr+5UdEDowihppKfUM0quhMYflxmNeWNY55s1jTJ
tjaS3DDfDKlKZGHsQnC49cwK/JiKhNlP+xBwG0YU2m06gK9jIhmy/34vjdym
6I1qM+ucfK+75Z2B4pt/o+GlDvgSfMq08EHMfJAoOuPOjSB8K4p6c8AaIjPm
JsobsMNUhnzIb+wOemo6mRMKlsM1SHlnHjysN6cTM7fgi9aZPdGrMnEYTara
qJFMlf+itpYEDOTrbdAch6hmOB2bAfmxqMtnCR/ldqtY1BHw6zZyF2J6vyOe
7WoqMpwS3HKM9HkLrq+5AHpG+DT27suu5ltCDtxmD9abnZ6eHjXfUdQhEf5k
kpLU6JYYNp0YGgzQaDwtrZLDNXmHBLaCXKTYzjITMTujaBvY0Klk9xPfPJh3
3j96xXIqWSWoO3b0eaSWSTDP9pgOaxzD4D4DmIDWkHg63ysU3BuhW54uLHV9
Y/M/HN54J0dGK3Q6N73EfFqT+anxMzytv8ys4Io9egS9V4eAFk/igTx/VsHg
40iTKuXaJBKl5AL6ltByzEnXSKOFSBpsca7x+MscGhciQM5cNdO2jIY4blPU
lEtv9ZlXEgfwHKJirordpFsHunUKQU0NWLJhC41LtKyr/eNGfyuY3fLeuC6C
8UVRYX9HI87dfJpPP8qQbVIqPSE9v3XHNfxfWC6VoLjFvBipKXsH9AY7oqnr
GoKbHy4kX4L4R2XO87nCfl72st3yN7ygI+ugnSUrKv7/xVtv/H7mnkOlcMgY
KHS5avp9NICTeJ5nFHtvEftFmoISpd0wiLqcMh0bgvv3VgEV8X9LWaJaB9gg
gux/8C9k9oW+C12plFZwDgFKQrnCULV95g1AoiTVwhecXW+g3XW76AlJEHPK
z013RZ/HY6+HHnPImVk9zPSy74F2+ZVSSwlQQScwpUZCgY+sIwLt6VMQf/Ui
MjEosq+UF1hneyF4kG4UYDDYtwhUAtVLfWPn2gJMRsz14nPrM/h0TpCAyCPM
NOcJT8HhPC+f/XlyHooqI13B8pwH5nwS0RHLVvxZ4nrAm4wK7bAeJhrncYt7
ulLCPY5MadytJIoHWVi17Tgz8aq5EFtqKW8sqwi/ehmagne9h7ugDMOx4tkI
AW5jJDiWbkTo00+C9Sz4xwwMlGhdREokYCE5fUsRn3QMjtdYduLWEGVuIoZF
hlz5soaJCXwJVxo2soeZXTEh1Npcmoqo4Rm2GNplevaPx7v+YWuiXG+wjs8R
JSdJA8yqcqZdC8zEI8advlEgOLe6ZBKwPYlGtX4X2uCZMyWzMbzxX/I7qmJQ
zbZ9LdCpJdiAGwuqxFgP+4NAAQA4Yf6/dhdk2pBTuIG91bpXDm/CkjpoOPnB
XADEhb3VP6f6nLr8rjYN7MMtZwyGyxuLblYmk0uRY58HlJi9jgs004hIxce/
6ldolDsZ3Lx/N33F/K7UI2iPoKWAfFpOnvnVUKPm4LIhiMNxh7BenLmwshwe
X7EGN0ohGZnJVwFncytZwN4S/wqePf3twOdi4ekcLQG2MeOHsPSKweglHP7v
h/0EzWSgiKIjKKjrJcpChXbU5gjtipoi3EQUiKnZxIp7jRkXA9UfOxaAtcrQ
dtBsWaWeR+rLEGlYPWXc7RyUQLwxTt58tshS6MzHZA0fHvjOXbBfI5XzVITN
3+TuPsELZhGhRsnhhR6ZRusOHkAKTdzqja21frasT3SbkNlo4SDAkcJMDSFY
ehgdX7NyjGvGe1FXLIKFPvXNhxEe6wOVZDALkg+newKeG1CVqOCNq7JZRuqd
TaNFAm80o6D0nX2IITNnZai8x+BhkxXOiNVwctiC0JydOVjBjjF/9fnOs46Q
6bpJtOYTIT9ofwQbqe4YdFfIYDQvPKJWky7z7YPkPdgnGmPTHDji1gUtkpDE
CCoxzvKFljWq8hLSeoWEZ5THasFqaJPOYSOBzqEgC+fJqZhJTpU/cmp+pAm7
9xUQBPeHL9iHXBfTZrBXUPqXeX+Dw3skmGVHd9/6Wz7gEgEGi8W18RISt2/5
ggvUSTF/RrGtbOSlKVea1IaSk788DdmD8qIbQWEvNMbHQ2sQw9Y/V8U1j3CI
tnDYT+nejGA6fW5lYA7lsF6O596H+n2XVCsGMYAJLP+Lc5wKowR/0he6sx9t
MtzdXF9/jRc0oIJ22UqPkNuzJD+MRWuUOn4MuRG+9FMYh0wAAdB5tXnl/Pe2
iOIaHwtxuXFwVnPkataWBsMOuetrONOrNUEwOM1epspnEHOOnjcwomyjvx8+
EF3l4xgOI4XMyO/YaMUwQmCCjN8Soo0+ntOJCSmex6VtgkhIFUNpYOwBoLny
X9+5UosJ7EsjT9nyZUjHYvXcngSrBoeCs7ZF0Yzfmh+cehIF/G0vkTjwsS9/
76n9myaLPuR4R8z5Um3lyw10YsKEOtYiXWQIbyMEnZGmssvIeY/MS1loYMBv
O6II05rkgvnj2MmxdJFvTdXOGDxvpZARrIj6/TttzTyoSKquv8STqel6hdEO
lpfiOGGRTZzGP04BZnO8ZKNUoPqmjV0kNOsW//3e3pK1gEHeFMuValgL0m95
dLUbEkr0GgR2flILfIo55hl3UhDJfsZwpUh8ToqB7xDKjrAkVuONcbuB3/+X
sx1eTOSYvHsh49W2NSxKAy26xsf6CgPZRV0GIKSThzi2hFrxGaHEtg30EHG4
oqkK/+SMekG/l+Pg5oGURczgtUN4630sL0csS4mYoeRxH2mL0C6uizlDqJTe
+ZtOfT6Z6w6wi7KNeBzWhnPL/3BDlZpLuZq6fsGVednSocCG7Rw3mRjqRpqx
zo8qvmLvxGIaxrtE97/x1N+1GjeNoCfWG4XV9hNH+Srfa6FpaiVg09sxakRW
BiDHoaNhGNlLb/bucjnNddf7OEwaqeAmIz2dDSa7whtmKSC63oclmFIJNtyW
pIUmlleT67J1Ze0GUrWo2pXBSMG2tyYnFc7zMbv8JCwTRtXPOzjtAhQxjeMj
oZy7tk3EzmrhW1d+kLfXGdgyg3arPQk/5RfOBbwra3obD8z+++tC5vJ3McTu
E5GYePW10blZrTFK95wFcGn/KtI9m5pHURG2gQibvSdO2mljYcBCA57uyHbw
M0RKcOkN9eHPNQiKF4HImIdm2hgKkN76KAX0JNYzmy4O+CbYe5XuctmASpL6
c0KRmFt7R2g8LD4S7cFBmqgBd42uAEdbdNpnSSrikOycQRyiP2C+3qxi/TVw
7v66dCZIvPwBgkDOA1sYdrM69qEj0MSdq5Oi4jLhHu2djo0ouAcCDfisw2dH
R32rMmp1i9xBHYg5iesMUzwYtMuaKMfI4DNWomzubPqkiaSaUPq5BJEpijwm
r8tfObQantc7nkgCMUH25KQhabf47Gi1zj0Rhd+Z4N0RZmPIKwR9LkWmCQdQ
N0lq/GhR2q3lENyLpn8ERIiALAkVGRTH0TRYK5Lzwjtzlb/uZ7eS9i5d6EuA
Nv+CfbYPeva8ZYw//uway9534yC+USWSXEHX8PdWKhBU+3Yg5Pi64+WTdWx6
jSBloT1w0VflPQWtg2GaSFqr/GC3h04GXVBYTQHnH8xUJmjLov7JSBa01TPv
C565ygJcTXrPfMWcbIFoJoBi+LOZKC5SwOLlq90SS4DKhiTy6U729BsKtqpV
9KJmfec96N92SP/v0IB9kVaS1f0z1gtfjiPP8sY4hFYeY+J50qF45VO1mQBZ
vVnhj/n3Sao10lSO2LJ70HaL6WgtRPs7/FUi/jToL82e3+T4eWq68UBAiY4W
YFGxVrnARQdil1tihCnFf7Aq3f9nkTdONcwCUsgk2vWjA2yJ/BXghBXRce4V
vkWycRJUNcv7EN+Rf8r/WEpeCRSZnNP8zs7bmtT2mAcoG4nlG0NatwpgNOrt
73/byVm+6b3THre6G1EnWyTmyaUJg6CAfFELqJLnMszd20xKqRpcmRiYMMWe
iZV42MfTiZ7WcCi+mfmWgy4pcQvfg6rfjTNqzcggJRMEYGo4rIyYLnLtDka/
gQsT9xE1kSioQ2YQ+20Ahd/0pAVxu6jf9c7VQFl1FT7ujOGsnS0bzh0yikku
roRSWiMvuGFNIH19+gE3b4aCf0wbbHLq2qRQ5Uiy4X3wXNPQpagoxH1c/gge
cJ2UOH6kP4aHD2D3ZXkXulQWASQo8RaDVRVaveZLx4EM8LDn/OAZcwJvfiPx
hLoy/NMVTlDRN7DpmrWDuIid+CWtLmOnGR3QGKkOLxPQy/rvZfxfvDmtKc2S
JskgmO0D1lHrekujOd0NFpmGJr8rclWWyxG74tHujOp5v3GssiNyOe8e27nw
nkb931T3GBMM4ufHkpKAJZzx0F+2yimEV7Q87qMwoVxMiRRdQXNAmIDFscHU
13nYSsmMacYgDERxWLBlFV8o25fI71sGhUzpafZYXZ3E6pQIW537uaENyzi4
gx6RpKGCEdWCi5dw3uEdVPZpcuNjMKhUE7ukZJMjdUMcG1QuNCKw3qPNdp5v
s7DmK9/w5ZIQk/4U8w1Go2Sk3Gmod57pIQWr2z5BFZiLgzCWb0sD3N/AQzd3
tDQdVAsxd2H4iUkFXZOo+uc+H4PeE451ckxU/St8TIKdY0sFTO4O3dlYokDg
lFeSR3dzBZO5LYZ/SnW+ZW2wLGhXOxY7ruYddtx5xAE+T3arIFGRTDZXLALv
VS1FEQoBoCWmAAl5iTJ5SppuBxRVcqcuXzY6bIlQLjm0rX+Y09WwHTZnYmAJ
kENBWyW6hkll4s2l+nooogzXd7ASogI8oN++42NlWMFkLGhF3ZbxaJwihfNj
eRCQvv/dyPmvPL1hCdLk4G36MCvJeZwfajJZFdhCXSYoMj3fwCJ+gi3pZB+V
J+K5kU7ohlId+mSDju+ifwQLp456dsamtImFIQ1CcOdBt7Zu2hX+tq/mmSk+
a2I6tdmdwPt4h8FvHmFV8boaKjoAVneIrvQ+d4FUKVjHGpYW9sQwGPGJ1vWQ
vqlw79jr9M7WuzkXcHKxwLfbfnwTzbAvUbLK3I3oeta+VxH9abWE/ai/iRia
OvsVB+NNJOhSUaWrWoeTLjybdk9ueRESmMHqMqXEBPjWgGk0DRTFeP7ZYbPf
RxzBSgdpKcUOFB32kw92/uygG2T/dvXK8goSJfrl/jUQvI6+htaQkwrhPhUi
qJhnTrkSBsjTzct1TR2EARRZhbLNw9sBDTbKCFzR6jdsSmaoXN1UGLc0liW1
pNPd9I8YUXXSTv8usQrW77w8qVRs70mYQeuhH5lWlgPmwvMOazwzJ8wLt74U
xYDS/AWhZu77j23yew/mrHwYCCYqyJBd4Vo73CjvWtWnMtVhjgWbf7ungGAN
FJPCXKeVHhypn7ENa6ADXua2N7XLYNe7DfeFjnMWr2OITnqSCWPLvEvWOZJZ
zWYFGjyG7LbyFXdCKLv7EB/oKzJPWF05HUNqkK/zTTHM+Ep1yfNd1dqY93Nx
pkqiCnp2aDAUFXkaoGyovxbAclBhqQWtBDNU4Qntx2HPLXolRdkCa0i/qCmR
2gdZ5u7nXuWM0x+j2XZeJzEnjuHGq7Q8TUepXCrjPHgl2VyCtAKYsv5Fdze6
OI007QWhFEEyp2kCa5PMkwu08j6CKQ3IY3yzYP7a8jOyMq8NXnjB9ETQIe4+
McMThzv+IPIDdJFS/x4sGdHRTyhs2X9A8MA6FyxVdhU/aGXFAnYnKVnL76hd
wyQn7Zxrw9wtQGconhJquY8zgLHO42NMJ41EQI+mGMJDBKxLLgE5VB6tQxAd
QodfMBQ3os2xlNRA+uNiiSKBxFZzVxovCjO56HG2P8s6UUiwsLf2iQTnRScV
VjaMy/Cda7Y5VEkGmcklyM6ykKinTjNZmoHR/Tp6u3f010a4Sqsl/lfkpsMt
WMuL5oTVIwi94xtEGvkhGFi0Baw/D4oWvglufZuzA6oKURDRRLDku8ekjlyK
mLiaA2cJ5lZ7dg/DgK0YkdN/yK7GOguljjaUmjdtv2dB4mfgRoBfk4QirLAa
yYhQBJxPGAWlwhPma9jXipQ5KvCZIIttiH9pvdBlJXe4QwJ+K26YBJ7NBrcO
PmHhLgg9s+sHQMJ8nmPNUwGtOguGFC48aiosxPdp3EHt78DsyOeCfMa75SG7
HEi6za+suPeHtZhGL9gWqlGR3CXxoDlaZ2ekCZwUEgXd+24H1Q6OSf61lA6U
0njY9QlDW1KQndTiONZ4FdEKtSufNcpWYeQJ99ASXJMdH/qtaXsn9hxKv5iS
pcv+TkCndJg1mXily8VBgO81r3BpTRGpodJikOU6PE7XvrscgdMBDkUwM6N+
OAEdwjPceSEJG91V04VycFlas1huLiQ+s3uDmpmm0hbbsJq5ukE5X6Y408/t
8giiYoAr6OGEJAfQldy3BkOzA7DZXog7mvwB18sWezgOcyoR1M9/RC/O5bJT
HJxaBMljpZLO2M+yI0PnOjTV6txSvq1gIYsMHoqQLkb0a2WPOFQmp+ORvujv
lGQyLbnX9UoVJ14PNoYFS4oFDruzUiTqwrpQpWs4cFMSMSdGtAU9NN6t6Ziq
nKMSUJSovge5LTm2WCnWDNlbwv7rUJaK4j8PNMVDm0e7VA+B7VhUI16Au31e
YMumrkAja4OHuMjcm5n+Xw5a0TWqlO0dhXOSScOf5XdO/XRoBh0CHyecerTg
Ad6IZdIROx4xSwX06kmIWYmA8D9afHXBTBa4GWPu7D4HwvGqNnwGdrKbBo4r
lEC2duWhedGtkAKlUTJhH1c/DfKw8dVZgrypMTs0mSCAfk4yts+Fg35uPC/S
XcCuHWVPU6+GUQTu08mJXj/sjCmKP2xY1xO8ioRlCKJ5dNM5kHQsFb9dExQy
POhSI7CtZjNKyskcISjafmSCO+5rp6VmzDv/OtAAna72g6o9K1IoY7rMqczE
SRItZ0yMJiEuRGPDIg5TjoSjnUVWL9weUkmCLBNbDyHR07KKultx58sWapL9
+ibYMyDLoVmlpq1zrV/pQpivqtMC0aNiFjKd2UnPddD1htOMiko9b9rTWAxY
Fb3n47V1kzbY+kxdivBhZRKyhuzoz6S8KVwuCFTMM8+l8uZq8OHgBAqUMIf7
gFOKIlpG3GJy6WVWA+EK9XGEM8fpsup8ssg6jIYMZ44E9oatm7FWamgHJhn1
9bZL5+jrYp5G3FdUNEyfUdvwTSQvuTeokGD0Ea3/SX5kWy2vuyl1EUmrOyJL
oA5FIsS+hvXHSl9uUa4750UQbTfBKseB2nIj2iH1qrYH0p+56qbwhTi47x4Z
HqYSSO8axQCvWRMeuPfpITF3uQgIitvpfjETIsqePcLIw+RzACxzBpkSFeS1
Ze/MlRtKTY1398ot0IjFqUce8r4w+Q318T7TJAGDl5PXzugFw56EFBxSB9cY
Cry0AYSzyYOuYAaY+hBJYVyaTR22iN6M0rGoxkU4yOfpX62yuAoSqKz82Ej4
fwQ9XfJD8v6dbRros3dVEgf0cVtscm/HWojuVl321Luo/fMegpAeS0aubQ4E
9Ak9y9chr6b3w/DZZyTtwrJS7zLCaOh2RAFPXa0UljRis57B/eDW8W84q2j2
cRc3cL+TeqKcgD7emSzYINGKzuz0tBnVqw+i4cPMAfZb6SoVihlv/lniMxlo
ME+C8ZKMAcBsASOpfa/1sJiI/VBY5s1zldWTy5FBPl0/6WYpwfSxPimSDb3l
TRGo+JLs2Z4GPlYmaoWldQBjutHhb3qYCCW/7H+4uhusD97bR1mCJbkUDT05
oPPq+vmPyTvnf0cbyMIM1DF9sL7+3LSxmf/ue1DvBh9e64FGUnuq8yTCkdPP
Ne0iMtl/D6/faO14S60QMwLuIgQ6/sEe3LaHWOL6BHe0cTXmtxHhkRkB2tgS
tY0w4cl2riJQknGq82xOZS+TspiN73zj7THruNX3Jt74EGMy+EcXgRFa1VAU
mxXmQG92XvLH3jsch/tzI1rrSyZ0xudNjXom2m2iidnttgJjDgrpqLy1ZI0T
ncxmIickwx31ZDe3VcRVlEu728Vx2yB+6CD8K9RTUTL+Li9iXx19Hi4A5/vW
Ywu+BfkmzxoaMYtKzLTpBHH9eFJyQ3iX2CmD0EFuS4St3wsDFe5Sn3ai99cd
seR2t3EPMY5ulgqzowSzRLk02MmcZzHVFLdJdkvkcWjaQ8E48cvZGjPUU1Hp
qwa616mXKqL7x+N1xk586Sze2RmY/0NGA3ZgNp+zrj4ku7xDVQEEYvCKLynx
mIsGYfvU/6gxSSQiiQU5ImN8q0Dq77ulKChoykIZodRJ7E8thIHyzz47BLWk
rwp4ykDEwi5Fti+sQO+GsoX+0RiYGxAXlRR1XzHlmufNSD6JhjE1/u0wg3Hp
oL1tb4J88hdb97/+6bx/XfEZM088TYv3JjdNluguc71lFO6W+4Ab6ODULZza
t0DSvV3jXWfaiDUoLwuNoo9fG+K8gI6DKR9155sb8iBskY8x7PWrhqPFrGCt
DprlU+r+5yoMhHSg3qj+kpIcqtHutOnqWBdxiZlcm6ykz3N8M2SEuZT7Roh5
/vSCNNZtZ7+vEbJBquxe77voOGlkrY0WhxC9oYczZ2u+7YF1QK7Ow+hfxWPY
ko7J6hJdqacGinImYcEW+ugxiVdR9R5nIsTdsLy8c21gY7SSdEBc8UAETw+6
bF189Wxh42xY9g+euytC3CLf3dJC05+b8p2fP4lVuQGpRxaJdMGHzx3AZcZt
bqQmRiiUp5Y7mw+kxCGgw1lIBbbzdsGEjzMqP0UatJ69CmM8MyQP1seGDuk2
svZRYAKw7Ikg0QrVAlp474QHXOR3VKnyWxA3tVgrz52coZ5tYgpEUzSYkvJY
5Qbig9bEuvLpX3DHzZ1M7LTj9ZApCeJqa5JlsZXMP7C+UlMw6e7kmA0tDO2M
HXxYHwaGTmbgEm064+jm66rNehiBw5XGQfn00iwdfhKRqV0jujMO02xmbCOP
3VBMoRQ8RkT7HnN9t12c0ipK3lNWT/ZS9MtIfFuoOaP3CkQw24ocQD8Gei2I
4BAOS8tvysqhiAWlrTttKI1ia2fD/rpneb0elJJQ+X7MYFCd2qO0tPNgYcDX
HNeOPjBNAM2vMyHbrmAWMOLoriNDxCpf0gpA4phRMJLUtpndz4AVCUV2Zwwl
fSQgr7Hi/cP3A0W2iDvJM3TJmvBacV/181UH3kqOWyiigaB9ZhbQw0E4MRqu
TTm3LpwH9rI3+F21IG985lgAc1PLmmPiNear1337BEKJ1wkKO6MlG8z/9zbG
WuHRMMirc2viMJITYR3uKsM6jE3yJd5OuUmwiTZt5emifPPbQ5ZY2ih18B8c
dFsXkSI1ie/z6Z2ifTxNGs7ZemBBARd4PvmexC02ITI1Fiv3ahopeDOu8DWJ
6d347u0Y3relaEgPLYl172EaAgrorimVxSY0V7hwjaySkGk9oBa7Gis9JH3a
Ys4gSwVuuPmY2Rm5qI8fV94UWbqRiCeF8R6hvu+64xaQut6Wst0gLn+51sLP
NWfgWf34fvUuvZh3gQ8ERvJMe0+R3kSsV34n+WlWLBhmfwMvPVCwTdUxWhwn
U+JkXsE0I4PHrincgoH9tnQvxpTzwqyQJ/F9tKO7wNw96MYH+J0jl+Jr7/CI
7ByA6RVAqvKYP2JmHU+DnajcyRf9W5CkzIhnSrGTu5jvgCb23Ty4QAir8Vb9
YH3jEr2x6pXWjORU+Mft3RWz0z003T+zZKhaTrVCQF99+3N5K/SGVAFALMYK
mu1inCUH4hvgsY74V99Nol0ESpdT5KRO+47dikrKWOZ1ZBakj5grohMP6uD5
Mb8Rdqlr69+GPPk4oU8FhpeVx8WBxYxYpj5fFkntL2GTHWBGgmyz2XBMK05s
/nETH3WeolJC0g9mk5imtS/WfKk7C5XUTpe5D4JHwyV/tHaxQoUHELRqWOsm
aMv0h4t1OHKBdMx5T7Nn6uWDXHoYmfpogKj2augiYW6UT0AOwzU+UkShOV/T
UwUcJOnM5DF/lzDXSnTPC3cyNQ11MnSDGP4M+as9B6c+w3VFRUYSPvBuC72+
Sg+UEzG/cXtup/1g5311cFvtDIC3A+8m3FGHoE68ku6VpZ+1/+rxZD6Seaes
oK0EsrMH7zABpKZV32Ng4qq+3CjgA+59UFg8kppk8/vTZI3Y3i6CyXpvPZtV
kPZL8rk5SMDZfRw8PkJcl9hrrxwFaYa3F5DqDYjVHMsbyUtQOxFDL0A+CXjo
1Rkm5aKrz3FzFtmLzejbtQS8g4uRBkKL15gEYbb01Oo7h7O1+GA9jKS+Tv9r
CLqck/K0omHs71vdqwz2iHDv18xwP3l0sKC5SnMLzruGnSDPWWYmvIqd6E7b
V3ztYwAGxwVYLRsNaWRkZ/i9SRmYoV1xS9UY++XFWdadU+Y013AryoWmhO1I
yDUL6DoLSetmUPQIke34TajchfJMH8lz5q0AaIyifqUj65QEYVqIq02MkJrx
is842qySWP+Tt7nffbEvDcP4qrIdOfjBxrHVyILxMReqS6MKpkuyUySWr2Yy
rUVm9+tJrw9Y4ZkmqDa6DXefRSN6VenY/PSfKusfwlDiF+roQ7/93vLhtwxk
SMHBf8cpdtqFErdptE1P4k6I/wCm2ihQUzDCAHN64RxpErJoFpTLvZr/w7l6
+1kW/JeDww2hSjyujTYrtoRQZP8zZmXb1DLhZLy6Gn/DPVuVSiRNilV0uGp8
cMe2D6FwRDiTcQpbva1YhCBkliNXQAmRjPiNb0ftBf13TR7X+238uQXFiHaE
lLbGybVAhbwt/lsmUkFll7CK9/Sg1730XXqdWYNZANF/PKY7EWUmQ66/NzVT
5CoO2Nw+D77tG0tjiYYcOxxHhfwsp4fxJ9qgZcm+szuVddJXQrpg7xJHwTb1
6snmJDWgNpVd89KWTr5d8+kg4qxLq3Fm272EAmTCbQjCXVnmhwUSJT9TEJK1
jwtJHSIaHszOApzKqCM9xSGDIc8lNO73d30VEDPXjTR+gVRsiqF3qjLNBbs5
7dOdMVpzj6BYaaHyrx4f9WtbMwUu75kkR1D/J/xwfjlTcHyuL6JpgsQIXY2C
d7mSNwP+42omQ7+kFX/mnr0NcAqJn+Cg+lYvA8r3vV2vSOvGBzIIBIv90BU0
aNL/mprlXKb3V5aTWXQlJrFEYJzJZ5qXNGcOW9hF4tAixFnvzu3m3f/ZgqgO
H0J85Tcxtdy/lVDRmnhZTLgA8V7YrECj73aMRDsu+6ObQJTLVWWSNs5k5brX
I1NzFj4lRFLcWj2OVnz3GiEg4d4UF+3cgBy1niE4BWPfD8L2ixaOxj5NuyMP
5A/rC0Ak0sEZn+9qFLBkvYqt9iJy64hutoAphUD8rfcGb7LfaRvJnGWQrDoY
tZOc8YZeTzNeCntF0ECNb2kNdhWLyUfsZqAYm4zj2ausLF68IhjSZzpWrzDE
pkxyz4/D4ldMeFvCR4W973uielczfvxqSzt4LnnL6yTEMGek2BWugan3wKy3
IIBXOggd/Ievr4dGHNrf2y/sjw89yrddRxPH+ITlfqnaiDEHfmWUMkem6lxU
7EnMP9QGZYrXSNSyPkR9Ify9u4glQwsuDgKg5ofqpRIdC87Ho+lEQiqEeRJv
fM4jkyt3NCf3yCZs5A4SozU+/Haz9BSeTIhxEog4UKT8rhn9CUd8PP9Wnuyw
OgzLIZi1FfsUugZOiGug7f/fLAx0bP00eY4An5+2OkrWVFIwZZOOIEDb4m+P
rD0EKofrEps3no6vgESZT781LQ8YPOKZmhFgBHW2wp94HxIa6bo5WcFALrlW
bp4Ic5/SlVsb4SLzY8KV4wjoi59R5vdr4AZ8j4UXGKqQXeugDCywSd8ebbh/
69Qz+FwGKOiPljkAjTs1q//aBGWDZtIn5a72oBRN3/nHK08ZxFxP3a01malP
/14RELOFWUzEBj2LOWiF3t91IABY/SsCvvr0zHKjkpPM7skOBxaPaU0SXcWX
Qw6ZIpqguch2MRogEG3D0aS/qQKldO8KekcOmzoK5P+vmBsEDFdWXhVFNCUD
9R/UXlcrFchN3ttWpY6aBJj3ZhzuDaLWQFt6LbETIW09sd+1BqFmV/SomXBI
lrKscvz4o+hxveXazoVq++aq/nL4oA7CjIzI8JKLRUDyDozmfz5TdwmnIHA5
ZmbXEkwVCCX0QAHVRljzW1JJzd1BfHqHBJ/t29mh2e40w31fWZu6Pl4bkgbq
QOKJR5lONz/QyIj6YABuhgWY4v4DzGBJ+9CYD6xeichYlKsjv/AdQjgLjWfH
tIvUD6gMkLBTjgBgaxityt2TsbgVOZ4zPM8s0BXWM27uRuqzkI/V1PgnEA6V
fLZjUeHpKfnrHXU637T+WoFzX9VeXwBxIShiPq2Z8+slXiky6ivkMqwxf9KM
Xw4Ga0Wa6Y0kePENqX5WQtQnz1Q3u7Gt0ZIf8HrTIcRfvxkbS4FkIWGwrG59
qlKJ1H6FUzvukWkdfEXW89cVp37qVJg1Tp65dmSEJfjENn/fNNtbLBtFQKHq
u+2zoeqggCsqWF9vJCuUnhPfMLWzKAjs3wkbXCJpvhQYygVe0N/UUpeXV1GX
fr0tq7ItvNjnR10aocYOefIlrhMkyU2YU9N/65atNqjQuWPuMqQvR5ITQgeL
9BDQSN10tz/iyvBsWaSnk8vvjSliAijmkLD7v4dw6HzYX0Vha1JcRdFf4a00
U5t/05HRvECqLoxwISBQ47Dj5Q6V05jc1Q1zzF7Liok+FihA/OQ+LcV7wcgO
8C5uvLTzwGD54ObcRW5j2Rh+K0JDNjEJUNuPPfFcJQ9EoWrFPio16DO3ZXpw
Ex0Zm4IoIkq153QbNBPri7CY3jGoZ7ouq4XuxdjLxto5zEnW6ju/GRsFwXGi
r1DO/APMK3h9AtzEx7rSK11cFjkWthG7AJJlNMoxQcwYxVhck3lp1r0/2yth
kN9f2/bvHyO1by8ahXIs8ffYmVyPCQVwdpffLAiY5LiOB6/btKf/tMKxe5Tk
djy7A5VPGRExgIU7f7F+cmyRu/vRcr3DQF+zVCjnNQolnUbz8smoNhC5ohHl
23pRhQoW3rq9PHPy4YGasw8dJbFHE2wH9wl+D8BhxaOXDLXabde9RDexM8ql
xnIDAtjRrtWm3ePtjbOkGPhAmnV0IFi395CLOf5LuoS9zCzMbf3Xhg8gm8jF
0+Dyl9g1W8dPkr5+Qz0dNY+Z2nqmow01qmYXNffueftXDYRIXEJFsVX6rzbL
lwkehMyqOrVr5VWcBIOsFtbxN625KyOzDdlm0WAnU5EYF4JtZ128lMmKnrSs
g/RvTEYorW8tXwFu7IC+gLDCyolj0rIaETMuQR9CsbXuNmvChhZhXm60gvB/
x+BLj5oJ+xipfsI+ByGFWxjNfdSV8A8cVLeKkG+WWE8qRVr7Oxe2FYeFtoQT
dhvqkwGbur0wukvj3BeNKdCxfqFKUtquwpduYpUvf+x44TzMiNSoyL+c7KfL
Dyoqqi98AqAY/hbKCjKlf5UnUhPSdorRJU6JbzJO5g2RiDEqfXu1YYm+dGzi
IiUT2t8tBlIzB25Wn/dSTRiVqBzjbx+1K3Qu5MR39KyctT1RVvdTRN4K6fOL
/MWnS85TZGtZGutuCJpfPA3e2E2hydao4KtSSjg6iSqoNRnRNBlod0TcfA/r
qWgiTwmwaSR5YtdxfhCEKlXYMLTgyW/LCTAdyljvB/xaFX2iViwwKeVyWPAL
Ui7Lge1rpO/ElehJI5cS/8EPNUu/VmQZp4hAIXtRF/D1kFfzI8qC7IiPHU82
Off8ZB9m1P/NAo+GXUUuzNPP3U8zIZJHSN4B+ILDEEwPHjcZxV1NO4XCNmad
9+O93Q7tleWHlZZs/YQ2YNEattbmU4aIuZJ0x4Sj+DTaHJ2/1OAss2MW7kj3
aDSgS41Un88/EEo86duuaavQdDuOvCf0tVgTRS4o1gAasD18APnh77G9iYw7
XhlQafnMTCfMOmmDt20hpQVqVWLRIlqd1dVt0vPwqRHNNbqBdw5jb6WxmudX
PU6vXieEIOniTg0iw7hHT6e/IZDG2UyLHIMfeCqfGGsD0Kq3kSWNDA2SM7ZH
IciQkNrQ3CLpLQRMLvpm0TwoEfU7Sv2TdPDaR2IZfpUHtZAWf5rrxGDybiXX
xOkYvkg+Z9CpHmYtp/Ev6f/zMuMIM1oKlZyic35mkKTjqiJFPeGFG0aq89mU
LieKvf9IMZjidZ95mL4PyRScA0TITcpg+b9c3ltB1H0ycZCZIceCr2luO0aJ
mh0AVV+BGKn/5SK0rrTwn3Gx9pFkQjmUQEC/CRKGD91Rk9Wqje8z3JYYYLD4
Bu9RxNX1biBOTFXdj/i8nbPx5CfRRuINBPkER+PF9CO+eZfHBAwrArogRV2K
WvFHKLZl2CL6WwKqO57M/pWTm/JC+cr1bSj6g3PIM2Qg3GMgRwvc8+dPkUqw
vmw3kaULQe4MiQcI8BkFYVcj4XaremWVp3CjTQppbBgkTYsYaDrmhotjzQRX
qp55oVrb1d8zqo8GgRdtaNA8yaGcgyrKtYsml1JudGaBwYwMsY3L8iEeaYqJ
qzERzIu5buI5qyIX0fpYyF0w/JlyPrEfOc89pUaVJvGuPeBhf0eSSUu+dgut
NuemG4UrSr+3Ll9D5JEq5LvJSKG2ORTcxwwHPDAf3weeLghMRowXezmUmZpM
RkN1YCH/Jas+6C62AJNqpRqF93lRHYWvgugnTMjaKemLKTDoiMyHUOFGiLF/
0EYyQISKossDXFMm5PKEQdmFyBVezsbc5ck90WYSAgRyoa6xKFdrMUN8OU0j
7sryDbpajFPDvMgXeYgvCuhxBZtwaAuMIpjBmaeqrl2oJ8jQ80LzO0Nm6tnv
qNIEiG5AAQXJP0YK7kxlU9LfJ/4FGSPleyaq5c9nanomhYEpbmVl+ETuTuDu
++MPn06E5HbCQPehP9ETTBIY9TfMuL89/9fkD2OecsCmR60EyL1WcPaDfTDy
vM/rO4giGaZuzt5OcM+bEsxwD1/xqMYBT4K4mu/j9H2h7ACCDQeca21vmh0F
Iz+7IcCRobcVSkbn1dsnoTfwZ9IIYYO0dludHVuq176B/dbLSWj9NYk10PaH
0MEerDIDXLlS43JSYRN9u5h0B4O5+dZdLKrG0bL+LqEnwtwZ9tCyt/6xQdaN
Pupu/aZw3vm0VOvuCixmvcO1Iw64zhCsa3odfOqLLDn5Pj2wH/cwB/cgZY7F
s3gmfANlxU+b72PWz2IKgdhhwJd+SKwfztj+N2Nzsz/qmRTyL4AIGzui8t3Q
qGkewKQdZO8Tju4jJ0h7n7cbS1qmFxte+nJ7fr5XjokUhiKINNIvz6RVbGJR
ftRWZe07q8FJvtuRIPna8/antwW7ea5SS9rxg1uj6FMhNc36odntosmm2ZK5
s8cAr841hvYHEpifTo1s2OGQqJpIgNurJXkZ9TsYOTc0iirRmaznxrpt08mD
zk3xCuhuHxProE1wzT8zsRe8BW4lMP4u4EKJlyl1NZU8ehmnpfix0kciAkpE
JTeHOPn6aszbaj8GQFbfGYzfrn+ApIWOcPwrz5LxYjbh28l0pJ6fkVSYUunq
RR1AF9OoKmVUsMbZjtIzDMy6dHClJGOtqhnrBZTU7B2kUtLEj3yxwdfDOHwV
b9ek8DzctPEcP4rKpDG6VQ0RG/ZWX3gfig/XPu05yuPxtHp7bFzSmt/jzDwN
TwEtOK6ofFOnotb+JJqiSybO7VhyyGxHC4LDFrlZXGvVhB5FS6vonBv7mLNf
v+lrg/MHN1W64V2EHGGAJ8R+CCg1aq5u1wDeUR6xftErFxYvreOy2GrzFLxN
fhwNxWOecTKrBjDZ9U16UjTY86u3k8cd7/EP2QIlHPkJKjWbL8KI8dw80XBc
BYEaayRo8wMjQHfH4eG6nQtFRuHu18vACk3oITK89GW5G7LqAaVXU2e5aGLN
Hux8tGW9KaketkGBvJGAkF0CsZgufaCpSdR7ndAplCj6J/vraaPAem8s0ybu
6ig3XoavDOn15I2tW7dx3j2J7RUHw2Xe7uemkdYMHmemlnNFD+X8dCSbnRPx
AJOCzEJt17hLrvfSX6ofzsOMv7k61OWsR9xWJrZohvDpOk5t0laZKUe4emE6
KhuJgP5gMojNR8iP9lrErltMOBZXFJKxjOyLd4+U0K+RcFa4+aIwF6QqDYY/
o1M7AiQSN7j1IPQOsYs5L1K9KyLcZo9Xs28zZLwoJeQPYAriguKZ+RzQhge5
/bzC7dBxcr3WvZV+Uxt4PsUILgIhPXPEz3Qy7p0sbZ5LGVmQICjPP8YY/fZk
5EVZd3aWMUMr8/lCQNEtDgy3p+K7LE9kXWmmzI8EKnsy9S6dTorQQl22hgeK
ATjVlyxWXIXsXJdHHRHiSv7IPDjGHvfC8aJ+S7dvnWCMTwuCxTbqXfSOGZhp
YjLh+lkh8WCoimGPJ/yOU5tnQiiNl5zIPM301kGMeKAlQQa2z/zyxYsK56zv
US0mHAZtGE9kdmC1R9Qmx/7q5hFQe8Er24M6bp0JxZNafdO3nYtrvW8H8XSi
+7STTayG5uT1yUYS1UhqFPMEsMBDWaE+3/HaQrgUzV1x+GQHocIOHvHiFI9T
s8kjTu0qy2arvdTBkJSH81N/5jFOyZUNCfZQrA36tZ0Sb54rIfzs2Bc2yHvT
yFFLqUrrjF/h4WBthKbiznoAJecRyYP2fOnhY6yInw7cKw7DK9l8psy6sbdY
gKHRTNFU+ZaC04DksYnjzlk9NSuqoq53MHOKJPA3/GwiSKcvFnXnel4ICC/P
dNtpxmgikyZZqBcquoTFMt37BJJii43avIo2QYOgso/prNFHM5bh5ZiMjyZq
1HQA+kx1p+eaJLiYRzjLt6NPJVEcGKe2p4IOOybWxGUnBC2ZfXBAH1hn1Gdk
qxJ70SxjMs6om1fpzoklcIck8V0dkbA1lL5bQpJgf4jojl93uhpaOnhLpZQm
SmdZzmy8gMRkFgUkUswUNh68V3hKTV6AXtwGBU5vB4gNftIdrnnhHbRhHYWN
7IJ2DVs+09dIUVFvKSZ3comlEdeMwoU9Ju80XM95xgDpMmzkOwigTQ+MH9+i
9lTp3o0gQmqL92/iP4V7GvOk5GEW+9uKejG953sU44u7+jhV3f3Z9GnPKDVU
INrbrLCz5TFdlqtRZ3kYJqhuqxjqUoOEhvveQMmmtD1cCu5juZ9CX371E1/0
5JzevBbPth3W73OsjP12BXEwBRnOtAlH0RskIhZHFKUCL4jqhPQF6NZ6J1Gx
KdYKrvNKk4V/aJnauO4e+Zh+WiDZzsPGQV8gmoqx5UO3qMxzn32fOWXSssi2
tapNL0FG9jmXS3SVURjzeAmCimHXjFyYQGK2uR556f0p7yLJVDwfcxci7UNR
f6jMco3EmVrJfpN/8wBE1SaK24Nmt1EDmGkggKmo9jJiaf7CXOIC3FUKJMtG
+X/lFNL/8ujwKsgbTeDliUIVnDRR7XwzsFXJlX5SgfzOPYqluy5MfQm5rigp
6TcHzS1YySTF2q8wap7f3tG4c+BIFZVVlkI5sacCebsO9ppOxj4h3eBPKQCS
rocZmdDyJ2kbDOXuGdFm8I7j+Htl4LdM0PvbwF3TfgsvIzNf7RD2stmBDXVD
oL5Mo74xOTdm7Y2kWnyVJRMbUzdYGnZMwLhxTz8P6BjjZoHErpVUdiZfJgY8
k5ww/bHrHJ1oF6ODOQB9WcGclhd/wkUduxA1+sJV2fC9XUPBVSyqHqutNIxa
t+4QQuceR5305GGxWjs5HGmMdw2XvVKLVZOd2OevDUPH1rucpATrArCBC3A3
rvrNNNHTCGb5IxU3eeMql5cXkuYj1OgXEkFolTSb0TGUENipOUakZHtK8k9O
N8dQcjwMsCfBi6qEGh+HeC5TzcZy9FVpjwiBSuJphaPBkVAAGMxgveh5SH3g
CgBNeYJT9X/yGEwvVlItvSqYi9su6tNEeWot9ToheFJ400vfB7upAb28ILtw
y1dqZBw2Coftutenuz+FEvbPFlBqx1ZVDxO42P9ETFuMSl1Ej8Ho13gUg38V
1cKXOLtKMJ8FKbAnkAose2JZMlRyLjGJZga5dN+7LqM3n6JptfIaPcoiONZT
KmLWDcWlWRr+Zwg1ZztK2jp+lYOp7Cma3Ya+5XI2YO1As/t+vetYt+2G/+ac
MvIF3m9JcUh+fzVmWGqa7iGW0zzxYIeItpx4+Ejuia7hoIWDt9SOwjps5Xvc
EQzcAKHdoCZ7OKOX7FIpGLcRhZWta0M8oRstb+WSKjLVzcJ1hV7tJZLHzHXi
NB9x+1P+af1C1B1vCnNAwq97FYL1IMCNboJXprNg0yX+iaTC3ROiXwxqWwGd
C81SAvBn0f5dGFmouCFy/Nz4x1jI4Wov5ya0Qf/0uCcZAO7DBejbnSohypNL
Y7WwRxyq3G3nWKQ7lzPQXX+WJZug8sTW1cMORA79gbT2DbmCoVQy/pdmb1OO
M96HGSg6cmUmuFx2aNqFprlrWnralEVzUBz0JOuViZP/c8z1fk3uUwvMBQq6
PZxQkQSytdN6pT0KRD21J/Een3CUMh0tyfxpfxHNNmvILOH/GW8l4C61RRM7
NLaenxR9fnl2UG8uxQzXJOa0ylTIwgaaTDqvMSTGynz+iAzUj4hFBu1aN033
YEbC+QlrI0Wf9E8Wngvf66C1N2HHgEMckYAzvRxUpDUZbsIwdiqp2yC5/F9f
fNx5C8b1fcsDhl1T9cPW/xo8yBQXNk7oZuv0fSX8pYMb0g/OKxs4+fYTPAdH
3t4n10MYTy4h3fWk+L909dm0EemRRgmCofkUPnQGJdXtWmNoJ9o4+5H7OPpO
ZYqSOVsG+mQrq4LV3AbCAN+qZbUo4YegQbnW7h3V1umexZ9G2GrpFaFlFXrn
gyW2qHmTqMDL93Hz4CukA+aubb5+BPdTtuaAv6rPaM23L294Am/ONP9EuI60
J1AmBVYnSKkRtoQGTDeThxnba4dyC3jI/VBLlOj5nmxg8LeI13gca5nCNJrW
I5fBtlJW+Dco3yERkwyjP9+Vo5Z1aVMH9o+z3dKE4rpXd6Gc+kMpCVk78mDL
pckcysesnqMAzo9z9lQUa4/SeunlmOEnbdyC01CZ1r0kc+Gqgl79dAkxcg3l
/5pD+C2jmhgZib25nL5tJwJtnVsLTooWRCApcjqc1oeEMIf2yGjxLTaGWtij
pB8Z4mcHzEcWGXplPpkkY9NMCBwdqQ1s9F2ErOHMTHt4MYCHf0JPWdWlBD8b
P2Vf/zJujAKIbbG5QnvnDqNLw+bqsbZL3IcjCorLsuIo/kFKqaV36QcYUZl8
ZdSgYLZU+x4PHaXi4XpkHDgbubM+Ad8v3obWGI4MmlhmIVqvi3Ao95WJtFI5
Fock6MLGBz5ssvoxlnPqYoibU8NIR4BqMRSeZhxMfasOiqE8m4D+SgclV58D
dwq4ZOr9a2aVN8JXjH23Kfda66t3n6zzgtfNc2nphqrhgy+qE0Ocia7WR30y
uCJ5iPF02MGD1P4RXf4eOgYCCLv7Ab7FP8DOXE5HvL2NRypphcwTEhyrJ33I
q5/ruTwwsI15sr2oXwPgpK7ZK7+CRx8FnVzADGkIdgElbB5w7KNLPIr3oqzf
oJ8knc3o2BUcPO4DiuEsPYjDFpVoyzqKLbhBOzNfKKkji6G0UvlLFYGBvAoC
13KOs0QA5i8WEaLkg1qs8aV//SZXH4xKxojKN4A9mTAhSZdWwg3EJmq+LGlW
k9aSElYFqD/R7dvgi7yxeBDRQXYXKokCFBy0i/uPj+lEX97pY3dcs38gS56j
9pRRld/OJ1SvyEDFUOwgta1Ht5KX+PeXPq//7LVn/wfGc38j/V9FWyW+euPq
jN7CRTZ6CVQ4RBErGGsRiPUItewIr70NipuZgw3egxqmg9b7vKriayJ+nou0
u4C2vEV+wLHU4TO7NIiHJEcssQfhv7KIQ/U535GlBFt+3lgzHNS9oKbbZpNe
Vt9cyhPcBZRAM0akFRLcGwKlLRhLDQyeC9MjqcUKvqVkXixpK5rkjFb2Pks4
lcF8bKo1ykxLMv5eV2sy9s7iBNT9ld6kESp2Yi1a8Y8tmgNa43IzxGAgJ6Kk
9n+uVc4qFWIPvrz/yWGRDqPqKn0FbFEypW0+UwD6nlnD/FeTEc1nVu6cWf3D
SSSEROAR3l1ueU2AwEmNyaqEJ63W8At1fn0TEOLb/6m1s8ggPeXdw8YV+DFy
OQ17ptOw0KDYdN8IDfvWJy9yXOEXv7peMsnLqGK110lvsrBL5MQH+lvPdkga
/ReKeoWt4iSKk8Ut0mQPonDoL/Yh96SiYHKJjcFaLBifj4NgWAeYrshZV2tW
K0MDiQ2fxiusQJ9Vwp7RKMG/Fzhc8gz9+jffQIKpuUlkqUPTFH74tVPryYRR
2ceE5uTmiTjdZr78yOFfhdfqiY6MK9gaes3HohEWjbvC1gF27hJsv0vcFiYv
UL1lFzoWAddWPCgQ2Acojb1WNioY81kotrj++gg0Kwdbgxnmw0EVIwxHSe5t
OuKOMKcuWbXmnU0lw+rvB1hW6eVnqQtlBC2IiUPWYvCqxqEt8CAFYlV/+AI+
DBR7W0gjss5L+S3h69HiVyOGX18kmUbeK9ab9xnnI3/NOyAT/UucqLWfRq+5
trhq3+Voh9zSNN83AQjhDiEyqDry+Qoi4+sSTB7XBXvowpYhuD8SQJSorGyc
PWQEHu9Ds0Y9I79tpAiYShLGF4mLscoUnstVLLIzLp+mGkjcBVQVnzutPwF8
TiV62ny+Y+KNy9BpCHoPvEPuDvxhsE9SPnXAYrQUSXReaUlEhB3V1lsPhEHY
FlHU6b5T+s0SaFQ+6FqLYC4gAtlmiEAo/z+Wsu6ACZIrcnwEPu4uVQH1BQTH
hXEKUBF7u+qJ/8pMTgesgZUXK6IFOxv9TJ0Pk9Oa98euonj38pRlpwe1kOGU
Xh+emC2X9211NuUB5OMoRjlF3ePF/U6R2FPPWERtU6bi7idmEG873T99Qb/p
tJeLUdsJeeqeMSNrN4C9Afyx+Hkz9S762YXqczfaTYZ47s3htvHJDRxWmsWF
ht3AtCXd9UoTmFX6aHYPCsesyc6xY3ZUd0bvqBetmK5bLCoPgz0EL8Wwd7fI
ez7jpFxqztQ1PCm2QyEKTsV0YwEcVeLxqLaHVQUgo57bXyHRpDqcOTEm/Gp2
WmvOUZnEFhSNZuGEH8J1gV5wuHIU6Vwavp9vnyYUUXzonA1ijbzE5/r5ZdIF
4yQy5hr+0lwXF49sXFn8+y6Pyi95Xz6ax+LthrF30dCl8auF0vqYsxtffNcp
OJL/6T8bHp9mME29rGdRCU+vE/eyelRSx4E+IPAClOt9Ow66dZAhlgflXtHt
Ss0cdSbLaOxoWd6gWK8TGs6N62CPG5P0jRfvUbJKp8aU/bD2Z8+Kl3AsbZKX
rIY+qtfSJJ1GYKiZCHuh7qiiPBsBrjj6cPVytr0bjBepwoqpcZ+/Bx/ZSGnh
OsGlAT1wPGsdqtsBg7VQ/QyEVFrcYYOxPORF3/4Yt/PvgxrKm0vY8NKluQk9
zfdOtuiggnwqPtvS2uqlCVIZpVItyPArttc7BIrZFhFtjHIPWCVhXyKkhlzD
vNkRhXXVWgwpSAmUANZvIOoCB7dmHPoclw4Rdl6SzZK2CnKApO1isnF5VOvn
F8eJ0o4jJTVeR87FGOF3kulcLgB/qixqpA9fxQKh/t7B2g0e9QyDevRkmu1K
3kQJ9qkjT0SfS+W1dVy21SAM1r2z6++ki/Nt5JvQDzaHjZ98uDa5k9gV4KMa
lTABbSCWbrpJu4H0s2jhdaEjn/y25vlvLwrM6FDnx14bTeEJAR1fmdLgP70C
ciuvilfZWpxPKnuisdE3ncFxHG2BgvPvdrukqliZqBESmEzejHjJxZK1M54q
RR/mGIOqaTIHL5UHKZ0lDcoX4GxR8BH2irGHfLDTR+veJkRUGDaL0GrsYUIz
fx6B5i88PeM96NBK47NwuD7ZGhVKMRS5/7VBd0ui0KDfBXqf2eq/358508Jz
Q7vl4aUDP2PGL0gTyuzMwMPDlzyLHXJ+3sy94ubHn03HXeATdiumFi3jpVu0
4oywSAdRdtEZHcvM4lkGTyBUqQzLYCJRS4FMaQWqCSMBFlVLoHkn3gRBqVsM
2B2F+CWEk/zH28hD8JLQV5N76WLcLTp7pD86BlSNDxdqgsW+vYn2WuMkpFJq
+X0HiHyGC5uvXubzyDUo7Z9o7gcdjO8AeYe3JkVHNt8e5gs0mNbjYNGkeWif
nRbIosVjQYeSxwabANt4T5Gx+V51ZHnCvEtlDQ/y+4hb1iRoaaVdsAdR9/FX
ngMdsQTtewAEo8ExfURdRFXeodaaR02zzhpUorHilSAhzKrusghcHf3xxSy6
BXdoJRPacQQbOzJ7pgpra9Vz7zfQphJq+DI39yeIp+w29L5kePTBZsb1jEim
9RTPA5i1LJWFnKu0VymxCM0HtGfIpKXGFFpg+oZEO0lA34eSyCgFzr/k392o
K2NmOsXMmG2CIkObkIEhW7A77q+GypAXRBMgR0FmeEFu/QigmGPAmbJkVevP
EpFBzfRKdQinXEnoGHX75FRmYmOduqWkdNd+mrJfTfyWVg8d7NukL8+dilAL
XcJivguEY4IZsLViBsC6KssUHVQcaN/Yv3BsSyvEZ1u9n8FBhk2YMqZxTk0q
tbRGbsvS3OTCSQdtw43KslEsZIrUCC97rVrbxgg3IY7IiLlcdX2Nlbfdd0xo
kHoDQO+erZGEq2jukZAXv1nd4HL45xYoShDkVAxiTs3zlE6QpLqn3EDdlbjS
ChbPjFxVShPC63hgqu85U08cR7OO+6ZymetcbfO1LRloXrh5CYT3jVtY2Gn+
eD9xBLxWw55Mk3G8v817gXvywS0OX0mWG4uC1Af42OU+gdKCnt4FWuHcB3TB
bMaq/hjIXEAAvA1G1wHB0FQ3NmqltOHHzXmTvXl6h+A9yCXkHBUWvfFJ5d23
tR9t5s8b5AGENsgaPXQZY/iu5+SgtsfuBbkZf3z2Udg4ehRi7CN6RxcXUGjQ
MxAsl3o84fCHsK/BKRN308b1hvuS6DrvxjKVYd4dSC3eMvHDzzuExj00qS4m
mwyCLTo8IEJI5rC0QKACFXVBWCz/L5098hlC2UA7PHeGTrqXA5e3Wnc+FiL6
sYaXEKsa2j7p4Si/kKaEEHywp4HPf34mRuigmUiOBcKLHeDRNAY8t1u8/3F7
xnqfHM6Lfd5jxh5hp2F20md6BtS8CuNlpPa4ZuoHnrKYZQtJ+iHqjie87owE
JrZOmLeOHhqbMcDkWHll26bGwZTFkga82aYv5/vSQzXs3vHzG+Ymfz9wzDAV
XA3fOT18iyjo34KcboLCf02/dHbfXjhmitoreBwiMJejO3E0SpTIDrnm1rdL
XAlFkose0FWMOTKygtMQ07v8aTs17TqD/7CGxNUD/gN/Nym+SrnderDCohun
x5eNDJNZzS7ou9MHGNXjRqXWFrpqEZuwKXNOtBusKE5jaRqtVBMb8sFsIWim
IebbMk9i2jBxOjmK2SVX4eu+N54oIeMAFjd49TRtmgnshfpg9OD17U+FVDcb
I7yTy1/XEuvzUAMGpXRbrIjLD6c2ggETrEDafPM2W7PjkZBJzqSrMn5qEvvI
zfolcVelQvj4qI/itKBJdTuD3/+yEVigxqGvyNoMMJO2DV0C34RLeL0oAU0V
S0MFrPn2QNwqowSN1DKgw4yCa3CBvKDovEy6Q52MbzsaHPt0KN7M+rEImbXg
4NxbxNOj/e0SchoQxA2eEvOzVzqwtmD9lAwx+V1orZry1Ngh8regM6uuA8X3
ZhzXQBUn0ddrui/NaMvZSoHJujU8rCHkMiAtqdoInE1Qe/e5dnDzDWWypo1J
fjTEKbVOVi5mkFWYwyPI0G8YQF7EFMDmOBgEtA9CyyVmA6JTbKSwPWLDq/z5
VpPehOYed6iX+2wCNbHMM+uleknT5nefBxqROBkXpQB2/ZSaUe8ordTd6E7t
RNfZoqRTIWrPVSnpDuFzmjBORq3UzCiDeX3FlqBXXlfgW91L06gV7IDPUV4r
3TbRFwEiWwCaeWu25CVsW/CxVyvvNOI7m7eTrmgzooV8Fs4gWywQ8sh3nuIJ
yzi5luIrsyhMbflMCVa76HtNU2/mEqlnUhAy76snyBfpYXzw6WC/xps1LaWh
OVofGT9i2hRN3v1mDIbQhpIBh2rqzWUA9OwrQ9B37dAwQ0uvsH+6Ftgbu/1H
2+ePMdzGE1fS4sfrA737lovztzyDI4cXtAK12gKdi1ieYPK52iAOWBRw/21p
yE4e/ErhzWg9mse22Qwd6LmEAdpJu7Ow55yBc+zRWuw2035tG3hPY0W/xly7
fhNlBhO9uvD8UnSLQ4Ts1oxM99h0yymkMkB42dIMzK6P42zGCKttZQTmgQFL
1fToYUfIQPnha5SuhehWgGvb1YBfnP3+9waTd9QtASmmlpSFyhP0QLrvCC8x
Xfdv02RMA+ptREzr0Xjpqd0Ha9DBx0YEi7jrOQ1fGAcmeFfHSlvE21TdZddr
YBA87ceIpyWKoZDc0dUhBh9p608ky12MbOsNIh1GFg7MQGYnuNQ/GCfcTbU7
p96HLsotLZU/VeSWjR6ny1REgdPNx6QO258WvBPVafyYujiDMZqrHOU9S4Yi
bh5VKObkeZ0hCNCY441mWZK8aIhQItvVjPpyMSMLG6KLwEudFlHiGTkQRLl2
RAkAhL0muRUBmozRerWKY9WN1FUXtB42FtOr9N29lQU5sdwzbqIFHXhuKzsl
h4Vn9RTM4xMu7e9jg2XisRDt+smKsWPmVf3WGAjKN3lD+5nUnz28YBzZi4kc
CkazktPnDb+tJN/jV6wOQwwo4sR1B/+NIclGQZ+pEx8zDign1ZktPo+k3Ltj
ejytUUgc+Q2BfKyFumVq0FLkOzCLNPBm8i3dP/R01FGHDRzyJHaCY+i8OTEq
8vGpPXVnaqrxB3pqCdEk9+JUNZoi67BWJtk/xWi9W3vhmxD6Jm7adX3O+fHe
as4juKK3wuzllHdGZrBsEIFy55dZYSPe+Qfk4PND7nnCN6xxxn7IuxrtPUlP
KbPGARataax/QBralsvZ5LqlCm+UV3hf2dQ9fxM2SvTofu4VVlENV1T4/Ez4
p4MyGLPNxfNOldkkNcQuBIyt2+FVEdz7m/RBAtjJex2sKwZiEHmKSd4XtcIa
l22mmg7spASq6Ap4Oob+flXzz/9wCecT+uyGrQ7L6s47xJsWXK6668LkE2Lx
u8uM2byl+LS6PSNmQBCg9PbfAuh0ewVA46VybiqYC5T/n4hZ2ht56qKPyqRI
GIj7pGO0WGhNrquOylmms7JNkZKekXGLfJEdRVLQqDCvFGkJjMNUzDR3ASw4
4IQFlYrH1IC9PxWE3CnxCcT1nZA41gEHnj5N2xum0Zed2LGUMaghnGDcadXA
5Cnq5o54kVfu4ZeIzX5VULhHYN05MawWayz+uJcjBGmERG+mzasdA2BYrTVM
UhXbFo4wvgR4HZweeqmB7PpepT512DkJjLy5TqPe3qJcz7g3YwCosfRaviX4
MavpMSegHK05UkiWMACDfEgxBrKfX8vw2cdY0WO49SBwUCWjXuwneRo67DYG
UbXrsGKvHSDyMgKeetrq2dxqpahP35JRkoBGqAIuiZJzDZyDoWJu9WRnFHZj
In9/o4KOmySaKga0CD9yxWtKrprp9Oa9cmyTau2fQNb6tUC3A+EhgP3elefd
v0e8Fl5Pl5XaJoIImSjEOxqQLkSMP4QNfN99LUswIB+dxLsTyLCMV910SdZ1
0+3fPatQeJNJPUNjDBfuNY2fol4kA6u06OstsJZMQxh8NPcBfqWpNM2cxI62
URT2a0iLsf4gC5h9qFyQkBcYU1WKOZAQYOAMNRhCOziCjMKpPXmSp7uO+wCb
wsdHK3GxF+bWFfr2qJrdpzyvYy22lVJqZxaLNPEcTmy4pwjstRB5VvFcYgQ5
7VyGQkcXFHYDnaZW0dHRFu6aJpFOVrXa28vD3VB9ySMPohCLT8tk0v4Xxmh7
XdBCQXqPr2iJRCF4yeX/qgSmlN0vtUuheslcSNU3XK9tLNPkPLehQ9s7Jk5H
S4UWOLz+plg1vo0JqvE4L9VMp3qO1QiomK1W+N1L8oUB87NzDjOUc/phyghf
VZRdzLjMuO42XCyR/E2e6lElFTAj40Z4qE7c8H5q+JuET/ICLd8Zc5Q0/OhX
f0r6Fvke7HQYAGFKe92/yFi9MaDiUiJr2PUu5o1gTelzSt4xcEGCPLHleml3
3MiA8EZeHuIn71X6LUyDXUonbz6q3A0c892zGQBPzU/a0jF/S8ZIqrPLAyLI
bcUdxz1hIYMJBOkEV+PlicjIkVmqrhGrX0XGsC/9sdqU6oQAr20BTB2ORJr5
prMquEYd6TQRBckKAk9nayN1Ts8zgz0AJTuEK+wsJbsWf9tKS7tovr0ySiYf
/ZiCOHIRKdheUwXE2DeX14KVQsBRIGMoor2i01XJocfYoBOMPsksXby6SI2A
1AQRb94tkLhnjGhNuFH/rVJzXbiwVLBrMDB69tpMAw9uEY2rYS20M18o4UIf
dt62pXBSNloJ5SFee6g6n2BEHu4uk0SjSGR0EJNDucLw9t4SIzdWJE+5O5ER
hUdm/Y0cJc1HK+t0vwgRHpwxOzg0/3YPMZKqdBvznSBppuHryi9F9oBGj2tD
MZsC87ygVEgrDcP1nJY0z+eOPXy/wRnntNqmPSGld4giafmAEy8SBD3CLQmU
FFeGBmQ5CcZBTuP0C7aWmGw4GEZLAWbLhAuvk8LRKhFjcR5bTUaEAQefjxPq
rPMFNXdk8EcCuAA1aii19HWHb7vW2crHCUBCKHPePHy/agO68Rkh8e+twD51
MdSAo4BI/Z0Yx7nWH3uVGFya/jGwEMvT/3kOmIQRyQOQLvnZtocpOoHpM9MW
2v36FDmHc6Tl0b1XxuX8NX5Us7dAcqWIaJDv+ULYNaQ3Mqp90X5azU+O9ydO
cDbkOVyidpqaYUa70X/B5LBh9xYnxcTbiHABGYzWIq9II5j7URXyv4McA/4u
46bvXUe7IGrYvREnyZyB/gvaISL+8WqzqLRKCPYYy00RFZ3k8KIieeeA08cq
E599ROCpiPhJNO/3c4doH6MIv+mzV5XwvPptTa5pLtGYrltezAh/8HcGIkD2
ERJTN3aAmRkP/j8TlMpssjo0FxEkOyQ6oQk8WR5XiVCUBU30u17AljAHo+Zy
aEYrthRAZuteNZeehaVtMxALb1SFTRyd8jA7Xq3bb0Yi2sCMx0Cw1OOrfax9
6iei+pp/9JEJTaUdduZ4A1Cbh61gQABNokdcDNuczGnn8MGAukmnsWIZo6ra
IDTrErasVvvwmR7ItPyP/GWT+8634mplZz0SqvcsXaK2pIHD8vZ21wuwC1LO
pxtqLso4JHesghZeJbi1OpjVT69apJbFMI4sHgFqD3QK054L0QfCavxwiDoR
qqpUQU2OeVOdnMyFV1J+Vqq0f0+ZvE86i+mLq6P9rCNdo3TLpWTz7n1xBVHQ
H2XGH0jwyzr1ahvvnYCxa79njItDKCM5AORa2TunXcbKKRTM+BBpEfaWZPh+
wMihViE9cwCAlDM75SPWUD7diQ5gQ7ersojSw8mc9gYeBma0PVT/gOWxZY9K
kRrybAP0NyE+oisuRaGQwM2DhgKJPE2r9DdRBaviBae3+dpGKydIJyGZSHeL
ecQtdLEMfktEwGw9hzCiBp61RBv+xIbUlFqcf6rSik/FNFhOs6Tx1x/3xdnO
SADq6wzLgkeGqfgTA+RcP4r6HbJxnoawWpHLLp4SGuVxusYxNoCXeO5fCNMU
jIxfLWQP8Aj2Udcp2TKTipEUOQWsFZ3pTY5NPecm9xKJDZF/Y0rC5A0LuOcL
rdfazSexLRpsqBGv28UZCg6WSYJJ+Xxvr1p9BBHtOLO6yB0XotCLvH6NmveY
cKRk602JWH13+SHtm7P0Rq0gG61lxmbo5dCvN7YwzoL0Ekw9BszXSk+Xbwm/
RvFLomVz4qJCEFTiBHujjo/aXwZfmOztXMZtvkxMfQXitHY30Qq5bvvPSVGZ
v2gk+WveVCDYrCc0vcWfvWHi3YYaOuWB7thp40vu5L6ujyMvtfLBN30aba4p
jIhKK2dff/mfStSUONS6MMEHDm2eO2ArWrHMlh0aEEOiYVAZ9xnoIm2HJf8L
AGC1mHeqgat34dfoniJWcLHofem2mU6hEcKTVBfEjar1BY87tjFndxHi2VjC
YNWnVpPx647SWWbPH0QXQIcq5rDVN/VIluC/2sNoQRrgDkhStL3xKgmdSJru
s00r8LlBI4xNu7DyVAIpdGbokeWJJWOoM1qqYmVkvLtpxsPDdGqx/tJPOnTe
baKLjqjLyGYIYGFTE37qnbkRKU8cvebG4lGGtGMCCTyAqRD2dtS4QTq3Vth8
b2kkSJvV+QOIX8LvPK9jSkxLbigscqPtzKrcVdZMVBKJtDfn5cODEG/hePPa
psiTs43km0ixreADy1VeT2mAP3ioU4yjScauhomfjdTn4PuIu+a4hkRdFiFR
F+NtlZJDGF9/wLagveB4+76r8kAbeupmZKY7Ckr5gbALKn/raaipZOt05qiD
06pWy15vzoevP2aXt++tL7j1Zqau7vUp75Vx2j+byWjIY4FlLjORi9jmkcUu
w8+HSJUitCqe1ZTnKNTSkfW/zV3zZDR+JIexmjD6MXcmBozGcQeewZJEn9jI
6PDwCe905RpQJbJ9N2wpMKkO4wg1lfzgHG+R8/Ex3La2A+itUHl9qHwhZ7++
CxUTi5HlDLFBz7buW94yn16SYxA41V2uX5x0QGDLL87dWNT2l7zUVHVZHirG
b0SI8whoonwdTIwVUsKyjdWcCiiz8u7eHrMQL2i9opMyk7BmYY/6U+7Xhk2V
Db4qWijcOEGeQH9ahxqoboq9s+02DXaDLb2HhCyBCYy8p+UQ2Lj3fYCb8XU7
KMs8PQK1RTzZ+HHIm3Z2MaTaIFEaUBVQhGYrRCD4xFJ+JUE4oFRe4creaEkU
u1TyhmR2Wzk6O58NfN1qY9Lvm0KUSKMHy1/dHutnNZK2hclgDqE4wfmpesmH
Dl6syxwNYWIjS5GdsvW/2hkkkDh5mTnFE+tZCmtxh0Kv5JT598Tsi0LBDrvP
2Eyjl/F8m08blohAFIX8e1JYJha1fnySqTQJ8UPG4mKFwIlF1j2UxfVSTGpI
hwQ6EzDwUrS8rj8gu0Ucpp4KBQNesUEVRJxrgcJbMBGgEp4oc0fRYRO2xeYZ
Ba7wQH443vuooDFFHiGyktHX1lQ4l8/db433vxG2GzfJlVpy37xFH1e1GJWQ
6x/x/Ysm2L7s0l/jR5azugvqzrIvAQfa8/0OfSgMJ9dSIA/HLvMdjbyulYmv
q7Rx6ohva673P0XvMb8gFLIukSSvwRzT7yLTlIxhBeLr1/vM2Oo0dMhGKILF
dunIDcnpq3FHpXvI5ryBUHZcl7ySddKJwrI/Hc4JC7NqV949Dx4u5xXro+m9
3DQYPakBG+9/8ne/59TwLl+Ueq2GRDCYDFDO7Nq80QyoNoj4HyiQlUduB4v0
o/oY4MX7HkYOnCexh1y+VvWp1oNOHBRIxiV7i4QTZTGhGbr9Nlj1C398OExS
nXk7BCYoP+hf2+s0owVSb0jZA8f0WX1qw97C7JAHK+Le/rFhDxE8Q9FPgzVr
k5BYPi2saNOivtni3szWeDZfdX+XwivO/FPqPnc29RtefnHHpamK3paWXQvU
2C3jmfSXTaDpkpcnpyNf3pTKOZNIUhaAxfB0hip+9sI/R/nS5X0QONhs9U3S
JQbE/sxuA7R5VIiDhOLlTQsS6E9GjnvSZyZYYuJbqVTac+bsGTdhzZZx/DOr
2ReGFwTWrDA6+Wc4HbhqDk3nHFsxJSpKnHg3sqWFnWc4l+LmUHz5XvpDkt7c
Fx41wJWj77CQ3KOLSIsYok8XcbI0Nlqj642A4gum9JQoqvlJ08FKEgML+uer
pdMkUobSNFOLn3x+fgqlEW5ASNg1Ie0lMGHo59JFxIGiRHJfWdVhQDq8dyrv
64dyhv/AGOn1UJDxVqvu/XQWjySI4j7UPs0mNU5TrQS4v5mG3leL8Di41WRX
nNhtqWrYdUHWzt69GZ42JoCChiTq5focpSyCo4aRKuRsqRdbfjxOnnUF8QKy
nsDeQbLxtxJUYX7kCUKfP4cG5/kWxF/iOZYFIkGgB1o12c40JiG9997F7ldo
EI28pGJgfdp9ocneOEu/J9bZf9c+gP+1ArEYHKxknNbWpplpA8TD8bOWHYc3
2g8ckQM+PBf2fLP2bhbBpDsDP93wTTM4twVpDr46RblO4Kf7L7O2XUpFQLe6
sdfNQD4BBqKKGg3ZUMoo6tUryivUhxsnNo8Q/A8BtRcpc96hboW9BVrdKybX
5IYQsuisnNIveaMAun7jxeFQwaNMWwYJ7ZuPxIPZju25+dA1niN51m+TNwyq
BJKBZJcMGaeGsloPxNEd99EhpmyB+VrGYIXL3/obNauSdjLbH7jr9nfrnw1x
GqbFk8YKag0NHosEbt6LCnXN8AmX6wsQZqSiPrMyRgYlf7tqFg/mbgWSzXTC
e59XpRDCt9BaVj0oVeGtIcyDYoy5tlLsd2HoowaEG0N/vErD5dIVJ9GBkl90
lZ68Ym13STGyzDMg79h8M3Joa2eq0UR1mN/w+FCANvlCU/6XBfCGX61ALJwQ
rcVAqrBsk/eCkHuwLR67dhNJowXv4GKRkkWVnHs71hi/sQGgbgfM2iv/jY0Y
6jSJrb+J9U8Mtt/JSLKStOYKhNu5Nc3AhABSbX26VSzMTKG96tOYy9z2xqJ8
SL5tYgGlXCNQPo2luXmSOK1XM587AZEJOs81ncSy2o82jK4xZye/j2HGpR3L
KHj6gnr3v5znjhtf9lc9BEipVh3/xQgurObchMIxJ/p+S1qMA82pR/6DGfXg
pb/4nSkqCAOdNcekgQmHLo9Tf/Rm5zpJvZW29Dhqy9rVJMWOzx6vl3vwzpDB
qlkDPLk+q8hZr/TX72NuXKLfjzS5VAraxt6b1Dgem/uk+cCz1cVcZQqX7LLc
ALTQ243enN/goreRpyBsWcyvhpowJRiBuFcBoHUutqsgkg5eg2BN1t2NxpAI
AaSxhVGOOvIrLoHBELB13O4Z6is2/hutmk4nNJPSfljaRiqlitoAY3B7m4Tz
uXeI9lT6oaDZVJRSgOXZBP9FZpx74OiqQxr9dwUmTeWoN7iSi+457cDjBnEy
0cSOitGXosIl5v8uoANWf+Ts87dNQnE8PorHjMeTlXR8a2x/++LH3P/4lgML
23AyOevzOv/UFxnCGue1Rj5sapPO54ptSfOdKdbOYXURoVGm7mjiZBoocyi+
aI+lPiW5Mi1vXKXTXHOnREc/2jiQAr5JbDekztZPU3gFL998MhKh9esGtaVs
zilyDM399cMxOzA3tTseCtIlc76uPkqx4Qv+As+02Dai3efqFnnT9kjpBL6W
KJtGXr3HJykmhEBY/Yr4Y7HmnnQQuSBBiDEjCFPEghyh5WFxJhwQxh7j/O4I
o8XvmhF7PTm/cw9tIPQGCXrLZYrDwXZHSTJPRT79l6oIP5der+4cNbB49fDy
dahGsQgOYC68o19pG9OUFrpV8wrAIderbroTVCa2TvGwbJJ0v7T4lVkpaWb3
NbiUdzuMqDsWJTPT4jqkEx1WMiThnUO3Q2DXwRsNb8w4rdtwAlGBfaY1CHfT
rjLSo7SVg9eGO2uXSppwbBewOYLZXn1mdUPepBRpwdVayWQtTuBerCxxPeyd
vOirqfqaWKJfhdyiue/fWxcOt55gCN9vudRpjTOGTwFxgdq18W5U+BJtsQfq
zyiwCWlUIlqSBlQ+kxsptbZmx6kRiZ557X9AGbwffkzodiQ6qF6GKoUZO/Rc
gK8YvUuz5PWv/uxLCGsoW9AjNCZSqsx1kcO/kBchfRYH6zoOT45waFphS8vT
CSl8Bd12BVK1ATsDb5dnAsny9yyvZQ6OfyrFDbOzMrIEtYYZKHWBoP9dOyjB
OGi0XI+pc3zF5Dx4NnigdTXWDvYRJj9Qk1uNHJZl56ccKlHDBKNvGAyR/rWB
YWJlxq8RDN/Q0IaN656ihlGZfmZAh14aJcQ3heUNWNI1M+d2QeMlYdzo8q1B
5pzZzfVJRS/LGOH5Ss+qctpoeedlJgesFi9Z6mWnVHXtODGMe8TwpfHTUQfk
AKXbUKW3uJegcbBs32SspHUWZPFZf73cLvD7/cFrB6BakOkIAloaNEkHhby3
3i2jMzT8TEwgMoMw5fQ0XCHGLJabnZjSqqZT8HqRFnk4RJjL3GpC3N3GSDJI
uoTSJI3w1mntLjgHXtP3dP9GN4UHjo2fDIdvNgVf2+pjRbQgku5Z61YIdfkq
5CYEV0wTa52nopohgwd/5LTdzzLsqRBXA1UkA3ISk+d5IXFNbbiFMm143njF
ZpSd9dhJbmC/WMql2TBLitgfBsIzY0i99dyusjdkVtoTqYf4lZKwP32gxrGc
crSRsv5V32/UiqIfS5h9f9OoBv283tDBjNlWm05Pv4vSef5DmaLa9eJ8j7iL
0sQm7890mrJLZ9IpPPUoOtzEb0kO62iZP0HRj43JTJI0uac4kCGwH1SMJuyr
ocLxwkLYj2yDgqwMKWgnIsTBWZU+zmC3JmX+9faki+K1mjYkRfZLzesHplMS
BtwiYpwcOL2faQS6mfgm8IPMip+QWGDTHM2uvs6uAyHM2M/cTELJjl7e6oPZ
Bby+F1NtzlvRGzDWRry/79/ooyW56XPogeLWx6kBvkQI5ScI9kbmjI/hI5u9
s/mwL1Jafzmr38V/RjkFNFasAxF6mQYkYXhDwjPKYjz4vgpKSmnF3np4hTQ4
VFJixf16MvDzl4qTUtdS0OFwDEf1GZUU/p6LszfUW5R9x3lHdbSUnIKP15a3
xpcZe3+b0tzv7eJy62jmJnn8245up7cyqPzc8QcXjOyEN+xpGgXGgkbvhzl1
3Og8TP1EygTvnK6oV5xk9GuBZ5INmbG/GespW8GKzSCFBaXGXOMbN2aLsemt
zop14k04wnpHve8s7yNC4w++e5Knvx3kSqX+U6vaFdGIaEdmnRih/KKeFAok
tpM8reF6Ns6354oy3ekKpZi1LaKBQ3DyAQVsUhsCkaYTATYHfE0qJKAFcp9j
sOf9EAIvqdqvUmwpT9uVOjLevYH+DkkDgq4aoSbPgPikaA4j0kKRKabO0StB
3ANvrQrn8zIL4D/TvLa8bC274UgM3bX59WqX7chiz9o+xv0qJc9Mwt+Y5EZb
RSwv75EdA4/toWFkHj3VlV6tTYb+57UZ+ycNWD5RlAwkCNKBRAuevfA7/+LM
BbdC4KA2QlXtSlgiq99R7NVTo/qGm3tE+qn0Ar84VSqHc9w6csyYo7qFaJp0
P78qTIJ8Dx32ZEJA03eEEigsazPDs1TPJQP6c5yFEx+IFQ2qFpxANACOcex7
dyIWU8Qh5Ku80PsXUjn2+6pO5SLH7z+25ubusr9QKvAXU7qDZ5HYn5qJQzzd
EvVV3dU/Pd6WOx0/oAhaK3gXMNbY1e07LNmBJwBpiDCBfCbJpETsewGn1Ul3
ubF1QX3hPTZ1O4//LgfVGVXMYSEV8hZGmnu4z5Vs9L4eny/IpukpFvI9Ibmx
znpe5r4DpLH70ReESj8p4Y7/dp2lXoQrHbUy7ISdshWpxU1DhrWQIypEVV05
6qpj3XeqPzEt6oAKaOlg7aKB8hc7NNYb7CGkEqqAeI7HAv+G4oioIJ5YPZ/F
Lkzm/IqqpdVKW9DzB/ABT+xq8z1iKrDZA6J2Cy0g1JZhPu5ZQB0Wbw2x2v27
sZA56BG0JzoM3t93EmDpdTHbiGpQI+EVwhw1VADSxiB9L890/0kEEQ0Li121
n/Di1oLf3jTP9yMyAN+zuiONZC8CFnVIqjOs+4UPhyN3merz4xx52PxPAjw2
d4qvExD4OvhBos0W7eVcIGQK9itTlO+DRwiMSVsYS0oqBoQ1M3Zo/gfXjMaJ
botuKhahoXNSOzBcsZXrPbGt3Z9ZItMlqTqJVbBz4Yccx9RKM2CxHBDbP5Js
8r3udBY3twvUGNLkr1gn8ImUu5GeDla8RXJ6ctMn+CR04wu2jSgQxEiQFIGC
5p3USW2xeDWLv+R1b8TJTxRw40zx7XTPWA4Wic0O3LY62S2cHbiUot3FWdJW
c7ZrZobPxzFMlGyh7sHIGqEaNInALemdiOY9Aub4IYYqq/u3jSj837PN/b9/
mlSYyZoA/Bwj3ojeXnAuLX/zknqKhz9e5CtqMcm28/sSAs3gCzV5XXSPs3xm
lh/moov5qfhpT3pKX9tme4449hvSPlqrr4JFpnf+kugIMaTeya7AHV/ADtj+
k3IFO9IF92vvuzpvDas63ys6wk6GLp6/lu0KheIxEPDRAzPC177Yi6wvwN8/
xZHByu1C2cGVKDvxyDh75ruMuTCE+ssaP9M3AnME9hTXXd3F/DvcVaJcDz6u
3LMadr9QPtFA+yh8B6b1/OAG4FZ4t6Z3CFK+lRtMWZldTqedjjlzr5MhTKmf
T93ci0XXVCIAzA1TL7BfOZHnaBXq/GWnYX6P15mgbBRuUne/tXYLMDhkKZo9
CVMrYxUe/meu0WWQlT9QOQ3+Uwcj4iKLfyCM8pgOqOgewpp4baPR6QI+q0uW
oTgVonH133EjqNEqkCh7Pcqo3dKTegYDZ4ulv8f8zizoqw0hAgidmaRSQncd
s25pfi+b0gJ4hFQjujKUdiNx9yCXtv0ufbStOBfPFtoCGFrCQeMFemgJz2Xi
dcSMpiB2owbJ7BZMxpYoIr3dNUc98JN3GEQGuTxsNsYyhVWNHb1hsc8QtSLO
pPTPd6CXkmZpMu2I8y3dJlLBAsMxnGknEsSfcD+ijKkgPqpH3dOtDQTBQsHc
6TU+dfHrfIe2Wmum9r+9kfanTczR/Tr5Jyjl44lzMG//DtiUJYOWUZKotfGu
RJygnIwOEjM0Sx8+b0IgJz315DRsWfR0doAbcXncxDqnraO1E+poaz9HrSix
nC9yK5I8BfNBEVyAVusp0chf8W6pQT8LYpcES651qWgsZufHeRzuwGBL4vlX
PS5O8ZWS6czfh9drza8bjB4kLjZYHHKKZEVxBNdb0Yn26nYOBsOgbEpQ3509
t84PKeTt3H90PxN6jG8cKMKECgiC4Woz3/ddjP/EHEVt8gA79Ocl1ebWUAla
SOnOK/J5KOwhukUJn4W7Dv9no6qQj9qqTDKGEWsUipI5N+9YZC5jAMuFZLkn
uY1TIId24Uk9fMLbZzQ/vl9UVjYk5SpHpqgQWI7jpIdFbD4v/uM99JGvLzOK
vJGk545bJOq39tZ29OYqiuT9Zy3MObTbHbVuj7CC8PRPJ1t8crY4LGKsXvly
slbDbTwubMr3HUCFF87EZ0I69VSbo7oKXzqScPQUaxFWWu/XMu8+zweJ75lV
NrZIdKYWnYKOHi02PB+OViR3AD+Z/xGRLt+F6rzdnvmTuFkum36ekslMDr26
MBHADb0e9XsUEfJJm2jhEzZWDLP50ZEnUNWrbm6rdqgIUYSTzBIbkl23suuB
dGBsa4slWSyNL/e7Bp25lrpWDmrTxSRUPoF6/ZQ+gKCutdfrCoZTsrHyeNIE
NBZ069UfXSvd3rgfzORSpSN0KKwGku2Tr1V8x0GaolVfgITpSZOEp9Gt/GiK
vC1j2roSPv8tJfWgEZUbTCfc3WtdnMIbfc+eZz7nu9r0qc/3yeR898klSAD+
z6rJIpUqF4LtGunFhWJyibboNr5Sk13wYCCLCtrUpKd8nvB6sFYx8B2QMZks
3I5jIWsKT3sFMXB7UsGr1nbKpLh1IqzihxOoXJ5gPbP6wbbG2Ywk8xCF5T1g
rfaP0CWW24Npmbz4uk6yo+u5oqcx22qAQ1iWm75zw11UjGo2RIU9MB06jb2i
nRGIEgRaZXPERX95rWROmjdpatWaAblAHGQc/LMEyuh45X69gOY2j9rVR29s
JO0f9Q0AZRB49mDVYHbmgYhaLDnY4zMGxn0NEDHWhtHP5lXXikknW0D9X321
NhwZSHfbaj7+aPNQhjgXvUR2JRs7xRffYQ1NKg0VuNcMtnePV1v32RK8mWjj
83nsx/teoNfIm1NFrbcI3D3kcPWUX1ELBII4ZFQ3mghXI3+WuliaiHEmCuG2
fItCHjFgaVOV4A9wHtTxYqvmLYMS+tDEyJI6Tjtbu4hT8ISIJX6lm3ZPQtMk
Cb8pclyEjUUDZ6Jw/Ow+s/7gcG/NMvonJvC1CSmVYprNw741D25yMdkT3sE3
Dpr4n2AuCjzO5aoGJJEag59xpnY2NPiMqXeQB3lIPK9A12A3XGhAOPibfvBm
A1qCL/UYfcv+3jnoyk4XhWoSqN04FCbvRABuwzaHyymbZsJCsRRv914bKVRP
NDsWw90ImiSt/c9B5vZ370/hretv8RZ6+nVJfN6BxGxCUyOUjg3ecyb3xx+G
wulVKDb50zbH9csndRtCRtaRCOJsn83aCfAv1RVXcCsN3xBAzoW7T9tRFNg5
IW7t2CsGghoUl+egIYdn+J6Saw17nQ95gFpdMBiLAYqnlHJhSWLaofIdY6zc
SoQvZmY01viaHD1+HPjReYG/F00Rwbl3P1Ole6g2NabEnGDF/+UQtmCF0dFz
ueRSXwXZMvr3twM3XrZOUNhYdJ5xNNBaqVPS4g45dDPIN0A9IEK9OncswH+L
Mjxan3CdiBCys/aKLUEv2rNvnkm+eecC7/j9LmmfB+U/ymOgH2Q4Dq9lSBba
gmOAaq8fj89dw34O5JG+rFFVMzg0iRllRurambXleeuEqTJhNG7ZT/BNTr1p
/1hQUTGLIrWoZUMB4p9Rd8cGt56aqC6cHFwrIG6do4EhKrkudEr1yV4fhr9a
MmbxvfZmnzThHWCmsWXtAgIBbiEcJ4BWnHXXdVH9xlaTjNqn0vrwx7lhNoJ1
ThI1H5AEcmTJZb5mhYbWvGhKXOdHiR5rD913ohuz6mGPquO1tt3sVg/N4QjD
X6WeNmzwLyV4eEZH0uxuTWElKnPzSkqwhGKWZkDHImK4uYn8zk3qfrXzb8qa
kcxN9P8j0mGLTiPgdgHGeQLQY5oVqlFh6l4AUESSuMEQvDVGjOrfHJTZ8jEd
Dy669NW5c+poYITL7/J81U92QzM53EHwyZO7Pa9LELxESQBE+wLr0b5t3Be/
/wPMKZe0+5PuvitMwwFVwEPqo2/oj7kIYpxs/qlwbd4X5K2GdhEXvKqTg1Rx
JQfQv8tUAjZsT+U6uYfU5qjkRLK9WMHqAYB0flEraIXp8/8+ZdIEgMi/61vU
Su+Rw0mEFZFxgCeg8pbroa2LYlWYTn2C+t55dFc52fOpjFVSseG4kCPzGLFI
quPaMiW2oGQBRwtdhpAMkcOXkrDNKw2CBbIUVHUIehBwH3RV/4rUgGEaPWHS
fJv0Onj1onBNEH836BNPNjVEPV5eSSW/2y+7A0Baq2wXHXcVLHCBR3Z80dHo
4+Dn00iu2A+k+wBYfPUX0XaPTgLU+ppK0S9WuunLWitbrvJkEZU1klfalQFX
f2avIRjA7O2SYslbangsMoUzCkhsW8V9uLdeHt+4NPV21xMeRjkjoMU+Up3R
pvGP2s8K9XQKXr60Btw1cA31yonyRCCJsNQew7yYQvNGeVAl4tg9WQfpoLKZ
ExTYOMoe2RlDdDCTlFu8pdDVPwFwiwzA+Iqz7aR/UdPSIo0+4CTk+/yHoyBM
r1o29tmFx02fYyV3ECqNeWpHf6APNKrzF4ex3fYDBIyoS1XTfVFZ/hSF1WJH
LQV3VZg8yXeH2rXYP7guJtUUQ+B8FIac4EfDzVReazWHkgLJCwD8OtHze6/N
YwNLNaTL/VuKvFoe2+BdLNsMMiB61MjwwnC4HlZun203sgVZq+GsDU9BTBeU
4+fUuGa1ksOMAdGBJ9jUN70rgIyaduW1jmCVbjNLilBAuKb0yGTyQhIzjjbf
DBoXsPx1r8MORTfgTA2BKi8lwqYM3GaXcc3n3S4vbvU8xrO4Z2YHaCsd3vWK
wqErIGgmKg/mkFFgKg0eqzl4exJ6u6OJ+V5FsMc1Vl9M3soIqevmFAIa81gL
kcTHXg5GDZQLCofM/N0m8asoSffZNUQTkH4ZagJIZAXA1k52e5NxRg69UfWR
76zHwRZG/oyhJhO8pTKUkN+N1VC64XnPaJLH1ygWwLX2yMjMpG7z42rXSr0p
4P0lwf5LHX6SO3SCKFdNoSTDnMbOCDomklOIxFjU6lYD2m2znEr7o6jCuVtC
vgHXvJXW7dAFGLltKp+xQm8U6jU15/HQK46eTvmHrvXMdWdgPdARY0cLh8cL
sSiXudGMkxKPvpO6lAZPJs5qE6rLNEZuVeTJQuNzcTxKdgiUbhIlIIaz1vPB
JCCxTZz1Z+NlEZxQqNl5OCTQ28SlPTlxJzGny50SabYZbYYfJaVFs5M2IbJC
sc3ZN8KQH4QzYj3Qf5sIcouF9Lqm+fd13krN2dvXRuLaDN8axQvcVQB8ZUMR
RdodedUzdJwvyjrNZiHi4w3k0DoJWViFTxaPdA8FsUxQKI/tSYEZCXbH3PBI
iKWEbtFzqSj9nOdNXbvKwZkQm5iIrJxobZr98RtjnFCkfKZMA6AT1lRKsYwY
vId/a7aI3/Ar+0HPX+qcYL3fcSUjcFgrKiJJIcb0sj2HU7QlRMNng/9gtj6F
04H1mz7iWh1uV+Zx9VD7w4Ec2Y7aN1zBEcRgaMDN8MOIvPIHl5C2H+Cx894Z
98oPoBxMqfg5Ucymqg5wMp/auj4oZ8Y7iZbtoa15SPwWZ+LHCq2LSt5ae2bc
Zql/Iuv1it7JLH4pfBwYRda3JhcB/AjprcLWIvjJeqQX4WCHJuz4r1hOZkWF
crY31eH8BWtgwQ+3wThPfuZlV/9F+cSTnPTaNYxDFuHvvRe9nWxeVI2WhZPo
f6S4q3OMdxyaqfnQntAXwTVEuba+4sdD2dxF7e/vRASX8DZdPMIj/XzRpxXH
h+yB9EeXjUTKy9S46z1aXrDPcS/93FYZ7k4jUWcOrKEddpRz8A4E7xFXDHw/
P6QxIDQb/q6iWVO6PdamhECrAKosxKSXIyVNdCadYfiRdFzZtDvBYDgu7A9D
lx5Ni0I2f6QC1NBLlhm4noN7+7J7rQpdqKFzLcY+vO26/IA/kpYusNqyKlxn
CoWTnZLQhFEy0VYBwXL+oLzYKgOxkFK6Jjbc+N4/Iazt3CuVBFo6A/3A/lg8
6qAegUqmRaiwAEZ0qTMuL/L3JsDMtBMGBuNiIlqk7M7f7tOwzVADHunKcnQr
sn04i4xGG/wiW1Zwq9VGQL7HMIlaVrS0SFFpQucaF1dj5ITkFv0/m4wyfdp4
3u7huujwqfn3MUge3rjLb/nTTjOcdSpJmGEv4+FCD9tf0my/g+Jr77DXN7+7
d+HxMaqMTHCY6ljcTbCxfBqvYn2f0fwf7N5WnDsZswTDihj5kAeNQXEVirVT
dUVGI4Zyh5bQYG5lxiaw54q0UpwWdvRmlYVVCRvNG7IsWXS8oc5wpfwmL0Cu
Sm9yVJMvMl2ckjK3/be4Ka6EdUqxtt1quwaJxo6vtyxHU8Em5rQGvvfMIY6y
ahB2hYfcNXoqgxZYuLnmU5guxSfeij+hgal8EhSAwah2wwX5NwKBbH1DCdgc
Z4JNZNMPndLXMWvB1DGcgbEHWt+M4wi82a1J4XVzVEpDDrTDEVEfceMbhGyU
u+NbsG7LTwrocv17OUKUlYxDZPkt4jb2+smtvHSzWMmQucdpqyJXmPMZLyvu
hAixklahVuDx+CL98VwER0wCzz5UeyBvt5FPvJLsfPSEtM6bHLbY2fet9wFA
K9jiQ64xEbMT0L2F3OQj5/CEmNcj4ESLgAlzV4xw8GdHtXvRbtUU7eAuAIr1
o0z9bvG6VbOIKYgeWPcYMkCN7jYN5Z3tSMpAdpACu5yx1ZEDU03VOTyiiQrr
0ZxXalB+6hS9VUfIW0YOkdBNUbsWjsga+F2KfbcSqBw5w+Q67HDJhzGoyY0z
Ok/6LDIfwE8xo4Nk5tsELHRdd8aXrksn0ZvRgVi8erxGkFqd/o2ke+Bb21Bc
ktYjnvKjuRBRymEEzlAo+jW1tT4mKe4dtYPfey0EVJpXQ7B53ZyTAOdPjS4e
r2K4/ZYQGN8EHdL6nmGfDLWzPn93nzjApUCLQYiCO0z9k5+S1ulyz0pnKAqN
NvQddfGzsCRXN0ykK16s3b0xvV5+J/nelRGpLc1Gy4OXznEg5L7ozJdU90wU
jWXPCYlTrCBbdZVDSVSIBeWdpKoqyPfDYwh2AAKlXUWGR/56wEDqhH99rV2o
hPreHQATRrdmoF8uB1FXvHt8g3Ll6FljwI9WoU0FE20RsJNlOHwHeG9AWBhg
xIAG/aAP/xGcYQiPDzhOED/KG62mci2ZnPvu7vhgvU1Oor00BDiSGJnfzYkL
G4Rdw2LZPssK/Y+y6RaY4WbY/f+oZoXLvjTHwhE0G1tYTBpVdVKio5HLAikP
ffWX+kHWzerWZNYx1GPJejc+FZQZBwWsoCoTA/VNLlm/OBtwwCF4Js1aegcx
v7n2XDhJfLtTwa4LsNbk2e4oi7F1tVNtTV8hOc3KEhms2BEvySzAdHkQOHNJ
FK8uX0iK6rA8LoVQ2+KQCUKQU3xYiMfYBYnSWaKDq2II9NTJbgUtZPQSyG4z
LU6Ql9nTEBPg81WCOCgqNO24CNFNhQ/R9X/WNmiK7x/bmhYOqT6TRXPE875h
xanzacMZuRIWuHbL78eFsEvxIwzpT5AlxJD68Uk8reiUJZ+8/wFS9w+Gk1mV
X8/cgE+qHU9Q/7lU8DctVHZmSFEZHCbgd7pSNYcZU2mYeOn5RAqSqnHR8cit
LVj54JrxmTga3HDoSiDCafX/YUGI7c8iNmJqGJ3IxjKsv/0Ds+DOcywrTizZ
GACEnGMi5OmKKnhfFk07XBDhqrRQKxlTAJk7+JUcxkuYqHVrLRM25+hw1xxE
K8kl1ZlIhoGZYbQTk6GES2HPWtijxY82dnWTiooDlTnr6n30BOxaCoobKHRV
deAGEx0fTqA0du8x4DtJ0XHIYFn7O5wB9dcM+NBpePFCKEV9uk1vc4lSNThV
pjlxnxNONPsQYB3DmKpSYxaz+N7FmbdWvA/AGYV9mZi/+12JACEXrTYQ2zl6
6aT3jQyamv7q9JCTgOXKrW1jaCzyxgzHvrRaFfgDsIpHQtZJhDnu6rQ/SWD/
QOTG+P3yyJr5YRlp6+apb6vcaFnbh7ATBMnAAW6Ca2er/IiyMIS/wERoidlH
LkG73nMTcmuSuZCFNsC/fIy1Snk7a1LLmldJn62+4bJRdheRpfbzklnzQ3xD
V0jEqUUmOZOD+R7UNLXWrpp/DiFpJu8rZLv+m8QQkdvVryxXm40c/jOeGCDp
lFpjlD7h0N+kpDUIF4/XyJNJLQq6xZEnswKSOUnCMJoZeVU11qV8Hu0hgoRm
a3pzw84eQCAPV6k/CVGjvgIemNQjqqOi4UUqW1rRClph3ERQ7cNlxLnlyDLp
8WxOSM3qjzcDB4SwcY7fgmZN+3kh/wLL8t/Xsl9ibr2579FhTOlTn/IBbIT3
N0YLR4KkjOmgV1TOauPG5EFVqhU6WWjscA6jE69gvF9oAcDvsNJC0O0IyWx5
Y0r3mn2lpZivitTj08q3GLk4rrh9qXpGZgZ1uLrT3FFWNx1Z4MzWnX2Ld1cE
RMtYSjMyI34BufOPxx2K0GDhjFH8t4diTGCdUzWuRexyUdriBGtVez+Jc9px
vxyq+a3SGLm6L53VVsysXY4kDTBUabopVZNllFQLaNxPij0hjEIvKFjbXSXT
hp9j4ahNnP+ukfX2H13UtlSchWPTXOJC2XfHRFbe/ToMwVli4lVyGfS5SOO+
okjDg3CA4e4iWt7gSwuypa1Qu5o20uuzjYpyIdRp6p275F0ONgkD2DxADXsI
Sump1nqXd31da87ZsqguGXJul1JFTjoz/YptZYPrRGqcs5vjobTuXjhk+poa
HyFR1M3XMwhc2YybVgCI5ZI65lyo9z6D5ZlrtT+TnKwb1GfhLemSi/BUtlq5
esBsgCopXrYhIqAB0Jt4mB/Lu0spEqoXkUMp+M4kkxKm22OrEqxUsapsBckh
uz0uFBjJRPng6Ek9XT4h9i8LV+o8w/sdZJTgX/gmxcXlKoK11x2UWqGSCYTK
R0EQt0FJScU9ow2VySbjmCEWa1fnVtgWF8/pjPRl+6pZAx9OtXP/dwEncUP8
2SDSumFGwNml03vjuxBfxZwcfDYWyR5fFOhQfPmIE7VE0zDz3AD+GY4zF9Ol
lE34UdUcemkKG71+ElbSNaGzUaZug+mE7aeUxakwIWu+tMxNxtsPwy9/Tp+3
KNBT6dIyi7F+CkVU+Ic5SXZ6K/nI7KmpCADcZT1CYYPnqjSy7aBGVFfsrwVY
IQKHoP9V44VUNLNJycQ+zrTC0POp6Fkmjj5PfRYQsUBw96ZqSBNRJlEdxaVR
0O1EkB8kQLBowE7bZoidNMl7JzxS5xjm+buK9cuiAYsmp3yXcXwRCK83dH11
ZariYnarXMEy/ffeyl7pTrD3uXqckQANtC9CR1XU4/fBqy/2CP/bB9pcq5d6
mLjTevBpYkvCGmdSCAKHR7w/uK7v1HB4wOe0H38pjC8LV4cSMIXBoGDxN5Vg
jJ9JdwmtC/lhuciFloGYF8L40e/NaLQobZ0PTUCDqYYTiuH+ZUPxech/Dusa
uYZCTna2y/M/BW+gdkB7WbLDdk7M6OLi+Ii7Q8VQHLlfLBOSufLBcgjNidK1
g2B0dbpNjIguPAGZct81dfQFAMmBXRr13Y8aRLq/ag2HbbpH/eBMm+NxOqqT
1w90l6yYlqCBl7TfhNsNfVRUBebHaTM7Oo6F39cFNX3+BgJkjxJIYNPmWWyu
OwcJRpb0A9/gYUQsQRQ1u/EL5hLA2e1U2shlFwlOQdtZ+a1ZI+bhPDFP7qwc
D0YLkz9oiHBS6z6mtW7H++GUHd7Akva/zZKk3wnxPywUEF76g5iApzEb+nKv
KZhnCuSEcIiKupvWIO0hPK1KayOb83JrlzG6CvtAaoILLz4HvMxZXSuANgsT
dj6JVS2kcSPn7hfvGIp0zbvrRvC1pzyINtCK/eN1qp+vbO+4o4fcy9DUVJYQ
PjZeoNyhXFZWugOCNIusRsbZSlb4fB8xtWUBMHJadkQ3yk1ExPpVYsWcdPdI
LXtoylHmTfWEvBxEJl/3Xs/y17ordhhahYd/622oqUHpNomjCflzKpxIKlOf
vfVV3xrEvl9qgedYZ+v5fuT+frI8sz8ah2scwDWiUbNjMkdDPZvv0SqSZgJx
FXWLJ4oHmfekdubrS8nBSbPcQPPPFElWLUDOj5zCJRISfiy0JyfVPWLYgv6t
gV77n8qIBaAm9PKJTHyAGjTREnAYF8mNBLogvoB00s6wh6w+EiDfgFGieEwe
JrbIoC9Lnqv5foayh6CtgZFy56bkBcgNoVSeqL72KgYy5Y1RoEdMaNE+pv17
IloWWbnVRqvS9165tY5Bj8ByTEPy0jtoIrf95QSg3aqwrKzGHQz1/Vqqsm4d
SsDAoR36m04lP4DI0ij7hIlRDw+F+H/mBm5Lh85J/HLja5lDSbvxa+JXIJvF
9nJRSeb18y305v4HU0vuAUrpC8/4f2MFJQaJx/7i1g+v6YQOHDtgBsh0aATl
G+WrU84yZRlS5KKanpNlTQ3uqToF2i+5UJNBGcIYnZOqj6/NeeTXVIelH3Ja
oQjGeTsOVXHnn5ETZhG2JRmO/lL4qTXZOcN9UD0BOIVO8iwa88qlWwT2qtRd
s2hzyNczUeQpKPZpIhrH3KpNQXwyuvJJV/bVn29yNel1AiG2mgiccvcb9dgc
3XyhZVmqhsirBl9d7P0dVoEyw+/R0cJ3vE4AMEcsJGVNOCWMuJqQdKrpuvFs
bTBioE3gYYBLA+TR50MuCIOUy2IUvjteEJa6mq1OukN2EUKbYs8eS2NrfOyP
E266xLkzWXWlkHA96F2NQCojj/6IqkzCh/EpqpnUin7R0TdtaczKyWvaD3K9
y6FQ93vveAjmOAZedS2O9lCO9/WGcOaZsAE8PU6I2JQUTOKfICjMJxzU6Zj7
wFg60eCE5cYEZfEcJnr9SIFQ1mjKlx6xo/32rKPj0nb4tbH59Tkcf07eiH8V
DG2/RC/kXZp5qHiF32qPd8Lx8YptcAcKhEnDCz7mIwhrhzdFiOvExSPl9lI3
vr2it6oxifeI9bWDyMmdmrKLlp6n0TgoB68fltJQ378bIIE1EukBjOdHhfnJ
4JU91tzjcn21eg+I7rvivjh7khzE8Exrwkf0YjWJqdyBqdSnBdJo6BR3cuz9
El8hzVJ9bSc1HgMlhdLJRcG3WRskdVmo2oZzTJouyM511WDI0MStD7gZTY/m
WZrkgi71lLjQbsLE4vXmmV9dHmABns8T3bzNPzzSUv1KmKyVUGL8bFRWdcf8
4i1iJd0lA0qIOsRcOz4f3f2JFRzSvHvkbHcURiBE4GXSLlRUMNAlMPkbExpC
Q/fpz2f7nRT1VauYV7yM0ZWwykCDx9iXs2eue5+LTgYM/PK/JCpywIMpZrLJ
RbeAxxyd+AXSKpEedK6gdsjWl6bmXwNS7ftkIIF7Z29Py0H+UFXMlZ2Th72C
YaHTN9sXh/EAw5OhAkAWgy5SjFGzylxqagOtO3EhE8OO7jMTMEGwajx8MyOs
n0rzL0b+iXLBYL2lKr4ySx5yilWkZL3axMlNSrjgufsjQHmXThCs6Ydgb+ZR
wKzQZPm2WhEVIZAB46gtjb5ujbTNHePzKKFLkGYAElhdWqA5t78D5KBXhPNl
N9wEPICbyy3/Epzgnv04WlSVP8Vk9/1blF8xpIaxRiO8zC2ZSqSc1E2VIoJK
kgWyrrrYJZiD2KUMDxyfw3Jy6IQKttEGsGvsgZG6MzMAyiOOtpOBgObfqH2+
htSgMlMzv15/IeT8IVTAa7mB2rQXsZplxEz5SNYR6L4RlOJ/Nk79IshstU/R
ddx9+L8MdFKBQPbeIAJfeEfRPiFWYk+W1Jg4EEMj7nIGpXjzAZOCaBRU9a73
NfGi6EjHyrTUvtAnAhoRITZqZnam/Itr3tFzr+pPa7BjWjXkRTENP2bOSJR+
frEli2oBl/w6naesP8FNbybkwNxYTzb5PXJMxJKwcOjQqlZYblrGQ/hYPRVg
KgWJyBJVREcBG+RBzkHJvicHqBCT+LTHsczFM6T4bhWW+SO58m+ewjP4MeFn
Upf3dAZuTTHMwBbQrWndgliOXqOJAVb9cHgpPhh0j7QfBFAb6gpOgV/j9wO1
YOCelr78cmKuwijYGIrRwEi97GqViv5/UuxT/FZzFZhlslt3WyX0m+DFBKuP
ZfzN7JP2Z+xwDYbnuZrBAst6IhNZJ9N5VkPcyihIJuGDliMWSANtmxHEFMC3
Wt6XRqLTJn5sEOw+hmgKasghP/qEb7OxAH9GnHoV1tze2SSDF08eos6M6rgo
e7yuOrqefBNQzDdP7iL1hrIryXlaWFogR9pyl5+IpWL0kJTMuzbiQ3qeWLPK
YT+uv4qNEl8vz9r207axGuDkCffiOWVvCAMPZfQWM3mwKWzkcvXnj89+BNnb
LciKyz5xN0AXieAWZQSPG3Mg9uz7dhn8kF8hIG/csiuplRsvZK6sA32gF+zD
cDPFlsyAARzh/FGMHC0pPW65btC1ONw5Fh8XmtGNdWxO/zMJQ90+6Bfbd14S
4vzftWU145qM3SQ16PuSqMWtV4mKYMkOk7aDVNsMPIG+6EGqutAcbDvmaMc9
fVUdjy96F5nRzLApMb2NyklXrs3CFbHjpBQThPlMgzw61zk66oSXUTfs/q2J
FfdFK/NKU//SOcKfH0A/YCvO+nwwgE3gJfgX+vzfBksQDPbMAtWwxfm1lKPw
hG+rrGFJG8bMaNxzFumlcHJyXjdUMvyWyTrlfg+JvEmUwdV1oz7IW63M/t0/
94htTq5oAkyLCeZmnySTeatqJ5yN2eVUXZLD058X+z/MSM6s7bGdedp88azy
nmK3dHBX3FfAL1GlKJ6bD80SY3GHu/LwC9nRNu0hgvUTpCz+8xlfEA9qDLLK
BmsRT7DQKXAq7AQPmuALF5lfx1YijMOaPTyIeAbIFvbS3Hdo2NltxaTl3A7a
+PGOeQqKvzoOgihpQ1up8BFtN0tWiOTJLKT6Q+z9OHxZQgifmPbE0k/ahHkA
CyS+Qecd0/1Ecu7IXEQx/MP32pS6rAkW/SfioArHdO+q4N/KnPIt7V6HeNsw
B99zK6I6BP5Xyc5U3gds1ry1pkK/iv0pDfEkvQdzwylUwLfT165q9EXQV5kQ
JbjqrRKNYueGMEcYoD1gNxOLoKmDIHChD19+FzyJvUKNkPLERySf3OnMOQPK
tgUQLSAWduSsuxDvQX0F8Ir7KFt/GNZCOK1PsxyE06HpBlzea0J6r2lSGfOt
KEmAX5RX25HhqtKD4elj/5FQYNulTZqVJ85lsxeQfew4/kqNPqL0DxsBAHD6
GJraUIAzeR7YJ61Xo03/waw7NaWODddSNQKnT/fYx5mO5R5KiGE1RxkZsO3f
dAZpJkuoS3zF9rnM81nfyEX8xBrXpvCX1X83C3nFtV/BNq601CH+eFNX0yV4
oF3acWItcosW2LHFiOpOnWFzq2sSgbd4ftz5RVc6iaBCAg0aUrIMvbNDXitK
IAgHzXJWQL3q3/jrVIBQvajJuZegjQyYTdoYN5FElDcp1/Bqvc3RD2A81Nm8
P+/Hwa9JEGQZfFuPouq0CLedDR8D0bghbJYLjUUwtlqf9tGV4xPclPuyh7OT
VoJ3zjG6xg10EJPYvUUTPnR7MoeCjcsZLTwZ4m09/ZmPzbB2JqasbZkmshHm
DOyzkmOIrphXJhPVxSZY/hEaAhEC0Lvlze7f6CwpDHDS4mQUTvzUWbGuTm5h
LVsMWtouJLzd1RV7VpjpVckbjAT0BBVDY+dwlKWhlLdhDRYZ6i9ZxbGOyXE6
qaK++maDA8Ilo3Sm3DwaZ0pBY78mDm+H0qx5uauOtnkZEfipvbE+V7ZOtZMz
Nie59Sg0SqnrOXyRATLQCdohr5sgOB4MJ/kC9K8g+dA9l6jgWhBB1A/na593
cM9hBkiIMXLRkdiz763IDEzWWDCwxTbFL36RBgaQ9at4Ux3AXfW6cm5/1+dZ
0t/O8XxEfidpbBhte0++XV45ZqKdA3QYih+bEgHylxKPQ9M869HYTaOPDKuS
ZbZiHReWNxOKaPEfVTnUXgTZIY5k2S21dv8lrTjAnI9nTefnD/+SagTKRTZd
VD1+FtOY8ne9MqhoRlLWwC0OWTqCAeChzgY02j7Rn1CyyayPnqGLJJWvIYPO
z8s5K0eS02lWI4NEU24J7wW1zi6O4gyrfJQbXTy8iTr/K3i9YqMtg+I+tlrE
xKHRgnGxV/L3UWIRPXBwSR/Mn9qKd/i6jjIT9OVbv188aInRvq9Vfejna6U7
aniyT17z0Wp1+Ss4I76yrzbTBZ3b93qaVLkds0TelTROx6ZsHXBcOnTaH3H1
AD5iUWlPHdEI4KcSmCMUK9pF82Mfkkpmby/lk9aFV2FppmbW9PzoKpgULmGs
wfvx7BKxsUe7qeGmcdeSv9zWplZef+ehEuvTqgDuRowWnySu1Xyvx/jbohoG
W57/nVEXNQiYU1TosGAb65p8WQkkGTtn8cWVHefoEvTgdAOuMrh4/FUbGkqX
YBJFbOqgv1cKLkypycjEc4dyxUkE4XFecL0GhmtUsTrrexwNAMpN49IOx736
Prqp1IvXnUwtd/0xqpyjCP7hAroR6mURr9iQh2CiqNRJ42A538Uaen6Gf0TF
FGJeebWM8goS2vbfdbusnqxOhdw/9u2UrzVtISo4N+0/86TNFgvAT/E9HpqR
TULZdbJzhi55qzpycUallHTiuufKT8po9JEFMtD/f876erjfBgqoc8Qankta
nCBELcZx9Y+G2QxXbz3/hzNNlpxiR3+xDiuXES/5b7rW885Qpcho3N/0CC/o
W4ZV36772YDXtOlyDveMk5KTpb7c3T05fQGTJEUN1rB57pGX/zQ98g9goi/L
+PzaKCXLczWMHpT+ewAUkJ0h2tIOLXeYFxmiZTfLbP5jXBuQOmZIgT+litkS
I6v8hc3IYtpkn4bieh7GiNNFZ8dK6yjqieVPuDSwsnwEUcHezsyV+emoF1xU
HqrCwSfy2wsVS/9gl3RCbl0HVM84A6P2X/YbL5eNHj7ZAobwY0n3HC89bxZv
tl7tln4NixopAvg03C62xlnZLdnTbWZGExYTq6pWPSZUNZK6yN/1qXQh1Qub
fOSWQWjB5CYHL0j739ugte2MFXfQABDnrPBvPpIBBuyZKwVz4ulguMieniE6
inwi5DDa0oNWPGsGoZX7fLOFNiCF/t6qovoPgN7Ty+MXxoGSnQ5NGlcCVFao
f7L+JXStoljTglGIMuHCRK7+t5pvhy3MKeAVqKW2ZQtSj7HDzBxAmcekK8TU
M1apjke22/QjF5MpwUhgjGf2YqtZSGswX1pyzU43X8EJ0sW/C1jsa/cJgQIm
arMYMJqjXs7/+XQOnuveO1Bku2c+Y99+0bkAvaiCj05VrSOisWScAmSmtwhV
XWtxydJvDSkAG4UriUSaTYn5sxfLzhn3Fr6FnUM0I3YHreEd95sKZmVYUPbc
zX2Fc85vAwJcZiwwgarNlZeoFWAHgYpXPFQrQThb0jGgcK7nvLmDdmYX10kO
DlkhuDteXtJX2mjJ+S2b+w199rD+z3zlnuklRCWVW2LcEV3g6Iumd4VdEdpb
Ov438o2nUq5Gh7r9YU25NdkySVXXm0XNtcIMMUXJhGrPnbNWbGwC/l2DzJ5i
lr1w7xR32U5lw/9Lj9IZRFxzeBC2Ao5/NdDqloGQYmzTiDyjfWc6itwxfDzb
mO25/hehUVgtRGV/SqJjNg60HdZlgxkyNjZY6tKkVt5n1slzC28a1stMO7yp
zh7w4Ua/gfhPjjrXt78X69UxS2lhlSrimUGuAPa7RgVsSg86JDDZKR+TeVYF
jM5L6gtjuYEFtRon/5dYUC7FUtkM9V8W54At/2RvbHTJDgMS0Mbjt6lJFo7F
BCeCSG0Pgqg/aLPpJu71TkcQhRc4RDtf2ZG2Eg74Xvvb2fxBn90jZVB/qpo+
d9z4PVGzRjCIk9/d1lzk2a6tGyDgPJH9QXg6VIxQ/2KxUbfO2YPdijLz5KM7
VBBHTmR04hLrhBbpUEkDCehcBNIH76qPPra2e9gG+9TKk0IVV2pnKzMl93qh
BBaoBDn+Jd3Cxj2OjdnQL0V8NeXq0b8i5IwjiYGdtaT3xU7uQnc3HukEzxex
CAhb3JlzOmjl2z8wVAkQr7eBSJC7vQjJorT4I7iPADtFzV446ZEogdAcHm4G
2ma5yqbcR8196D/8hYV63OhueRwGFmBrIbYi3RO+JqOkKSlywyp9G5uaTrTQ
ot1yyhcKznbM6NVXhcCtz5LOedTJ6Pv0lu3yG9sQeEqJTL7A0OI5kd2J0AOo
mrgZEuSxisW53ithzHlXISRyXuxcTOxScujo6/2l7JlJ9NLW8kzmsCDmBKvm
py4g5YGB4P41Nzgf6rRr33r0wjPtgmh4wXZR3JGJpMPtWhzF1eAHyHPVI6Ab
cWT6GpqRbl11u06mQV2OLCfTBnOXngtCd3FkCq09K1Ac3Hc7KLT1hBJtmfCo
GGhH+XdHTgtL8AdRmvbKF9TXqTB2ZYlaDqDttr7iMWJ3gYkqfqVvmtadU5Th
WYnNzt/Jl5Adz6YKVM9n2RwHQsh83fR6JdEOnGhuLD97VnKKyTCUM4LHP2yI
KtIr2UDJj7FXzqjZjAw50/a5m8nKSozuhAl0fQLYb9T5InVe8jq9Ky0Z9Ecd
YWaqCR4WhTWCmcQB694SKg/8YY+4DWvRi0ps5Rrgi8wEjC8E6apJuXeTkoxy
EHNPHsm+wkB46/6EAcuRZ2xrUiKLfaL3UXDlwYIIENHpWsetgPDhoojEai8v
MMErXXpmxHaa+0S/nMUmzxM14Ez0j+oD6otBm0h6FXMkRxYakunHbJ0SvGjk
oz3b9zYXT3qfBWzcwt/1O9eoi+t4VN5m9ZdT6Z4z1dM3LeUO2WLEbYIW68/E
8/gd53VIh6WOl6S3dxHkIS4VMV10Vd5fA6G0MEc5kQ0prPyaoljxqTmBy+xG
JhpvJ0Xd8qLzg72Gy2/47BleKscBG7ybuGPdhtgAJBhL1W6oGiH0k5y0U/+3
sHmBEFXcdie+v3fXUvIoznhhWDl1QPr6rHU4lkNWcjYRIPKSgu502CN6ri3W
8M5kliOpVoUntVXVlyMLOuE8Zz7N3Cgz9p6xYqmoeWhfiTPuPe98ZUjwxcsc
vzTTfgOv+ae8nNpPyTvAA3r77tZWp4c6aZTYhTZYtJiYNIq3fdtj5gKNTsuG
gwgQ6Nqlr5BzcJtbODHd99yeYOGbbr+ykuDwdifBrybunbwJUzFhoIBd+u4v
PKhpiwV8QA6mkKXu+VANBEOO7VDVi18INRpw2nNhp73t+m7s4gOCSOOQZMhT
saiO7jjcvO47+JKEDPq3nIo/iDeElhIWnlA65+8WzYxDyjtOkG6GDJUxwoKu
eqTrX5DQ2EOudEEAdDHh0qWBCAbjFhc0/Mc2p+xbbn9NDgVAPV152tyuFpRk
DXih5zFdXQB2CoslAAZ2IzRPXvxh3ALtUtznvwXZ77sSzJz+u8/P3D2iU7gk
ZhZsfBpRRlvswqxNruglZfK4et3L49TlbfMPqATT5WlMi+aZ13Di6fkP42/X
eBIy0R4FX9lPXIosuvhrt6L0m8tkXRmVubPrHwepa9AFkj6ALFhchEjasXHA
IvWq5dWGKJ1hECX/62IQs5gdeiCWGTVTxuu+oFXpNkUbxVknp+wZY6zn62+H
LmGU1XFvEN7pX9pZ/iwuTVV75KoF5WvtYKxkaquVue7MD6sHink50+awWm/2
8VxUCUYVmHv3UdonIzAE3H+FLf1wQlO13lGEPOSUiaTAlZ6jfwPabtqJST9X
EdnOJYeelhcnBFH7zi2Eh7pljhSShz9Qo4gdKozH4HRzmbzPqgDJyyPSEsJy
kXLcDP0XFOgqnmegSKq29Otj8ipOSd8oBvhz7IBQUockoPpd/4GhnWbL3eNa
VH2BB7Z3uv82n0SrwNxHEHJp25ajDvOf4ZBZRn9HFwXU80YzvSfxfBR7xBbT
+bp1eL/mpmxRJGWnUIURGv5fzFMKSetgdX99SM1E+VG6H8S0pHeJsM2f4tKD
B53arkdWwVd+ytjyYOmFaleM7vN02eBqlIp26ih3ZrdWXktOH+wJj2gGg6h+
hzxADwSjKksf8yPeByDF8j8ErzDEQpzseSfoX2/9F1R9tiSP9PJI68Jcv0pd
zfBCHrMJOgd1BpOL9IYNz+rjsqbGv7olCd93MB+Z9W8iMU1zSlbK+0uXWW0p
2S7iRZCeHXPhpeTW+9O1hFT2+rUWGjohT01J3WvRyFylxWA2JfpNWYZd8Rjh
7NZHVFZWHHADVNuCkIpZoeB0l6OHW8d4l33ZhLp4uGpfdji4YFMjdNqccZWD
vtvmvwa44rHPK0jiEfh3Fv3HOA/yWpry09ATrATUmhk+UbywgV2CYhlrKzwt
PCuZUJupHAzTsoG6jJ2oYUOyG4yB6JWKm4ECxTBIg0f4Xj6f+w9nmm3p/LJT
L7aULalTgZSAtLz1/42xBFxpAMk/lBSp8AqB7vgR0z3WxMI1InlbafFS8dcE
z2YcQip3KXxEn5ODcq2y3rHWpK3L3o00YsZXLWkwuwGrHhDtAo7JhfbpY0nq
VN8ICOBKI9hXu+PueaTWHX49QUfpUS4/sLfd2h3pTVPtZ5wm89/ajGjdXbTi
KzOn2RbYe4BHDmVKDAk6Wk0j4rxkn2itqd6+LHJE9IEJUS334tvSy1CXpNh/
Jfxs2V7E4mqoyBJgA4+GiXUoZ6QbX0aP3z3I1Tk2+cAphIB1yTcIbAPOllrI
wrBNbRctmnZS84ONY6danWIFNZvISJenUd1sikTBOKXFeD0L+toIrMD6AmfQ
mIMxJ/km2vIOKqF+tMD3MDgzqTVh+l0uDSh8E5Yx8w41mbMdQSX6BfIFTh+R
3AXzwgiKToEccmd0Cm4zsnMCcnwMYdgv5lhw6Ris9KgciWBNPgDQG76F+Ssk
1JzQEx4rSTYgAYK5U+DfLzhv6VjaDFX6Of0dHAry44dE1LHP8AJIexP6H8wS
u9wbR5B+vCMquuyk0RLXrGD5cze1jXH/Q0nX4Te5XwIKzf8ZR0/hvPb9JWfl
nNFrJyA8Wderq5S2x3sMHHcHOHB2FIyyQ2ABX0zl/pb8ogtPimt583DbSsum
D/EIEyDuKrLjBJFYpEVa5s6bGvfX/kTKZkTujbapoyKIm+jyAasORTwrxlF8
0m2a5o27hcNRqIhjTMDKY6VnkwIHsNEhXcyp7o5/Cuk/xFogZ2lQhggoDFWZ
4XwGi+KT3g3xyA5CY6oz0bBQ524GNVQ4oSkrnFxHcaYzAzM87J2rmdzHNIPZ
7lKAVJPSM0BQiW5aEgHveCk//Z/eX4YsKR8MoqwoS+fnrzXna0OtyPXGxSGe
hfRiOxISf3wOaNRmeSf1/G4u498ixsy/BZmRZ/h7ir6TMhUHqa7LEKqgr1xk
214XPFhx9RGV8J4axh7hbgp6v734pultepCHdxId9UWiBPSASkOuxemskyqZ
HOVSA2XdhOp7j99+HWEBlP9B1rcGWNxI+1lKh7CkK+WiQ/eFgC83TfXewAQV
ZLAlha7wDFIf/4EgBSCphW6eMAAnByOwPEWxIN6NojSPbP0viFvg0Rdx5BXV
IG4csSUVtIyAAhnjnkJGgV3KdWXZ7DEbWxBqLLextrFuMBbyTGJHZzAWcpTf
3gPlbz2aAyAyzj5Et964n8RHVqI5VW0t/DvfCyfqNX6k6tSL+nYgY17PAe5Q
L65WnJjlSgSeNMzWpasy7+R0ItwYKWSQiBkLZawYqmk+Ys7HL1PmBP4P67+5
Gu+EQzraf4tHXvRPOYBVny6VzTDyFKVv5xor5XaEQkeDjT5ifZVI2Wu75ag7
hfXgGqkGmUDMkUrOU7xgjn09H8YHChLfitX09Z9mbXdTInU55CRn1Xg9zlJz
oMHC9YqYcK1MQvKwofyCGvVArTVavSZUefJVsC0OpmRBpMrIIvUYX9om/dQp
f+Ft/gQ8OLYsuAe56hKm3HekCG1IxZyufjktE7OqXd9do1iOl2FeIXpq1SHz
jRxgcFdKox5kNUvmCczbREChYXjUa16fAKGbq8NwiQgk2Huc6fFjFVJRCRcO
rBv8FmNefPBq5E85UN83AxR7AvKMM1XXtdEMhTEGmO/O7PmT85MTq5p6/Da5
ACYUnxsawgksZYk0OO79UtwKn8xgUvrX1GC5pS9C7Zz0+zEzo9sHW+aThnPX
xZty6w/IlqUx0kj8/8sGCLuZrZE0KFWEOnl5e9OWcYDJaPVVKhMI+tSSFJU8
kvzY9nLMqlJhs5OZJH/3ZLkrXkmzvT/yyVxO5Wv9aSaVltpk6+o3Nvx5/N+X
HEeNtkUSHdAaMsq7Ar4Q5IkjsMdUGTQd7NSS53JYiKACU9U0oTdU+tgg3ZJW
KGezaPJCl+YyLE00XbiTtWHJ4x1bafPFrCqFjj/HjwlLkEZCqDAG06/8/Y4/
YOSrWitogoeSv27WT9N7o9r3sZ4UkxMmIENuTtq9I21HOHKYa1cragX0NH8w
SF7/wa9AhQ6Q1XivHE0J513G0x4fEtelniMOlBc6nKuubkAGN0uXhV8MwmS+
cnFt7hqv1sgOW0OioZSVegAr2C/Njv/dMak0+TNeCQBE4sOw19hm4LQQamnm
jTEG1Edyqdpx1t+jv2PGIN7IsTzNRNibdLHP+2JrBH3RRbUdbxrzn5HLJkif
5nxuMcx0VNLaRNHkeSzQQCdFDYw+L2gTA16/ilNE5PQZ+mNF4wCuo74kK4h1
b/m5HO37kI6qaQul9Lqk7Uvfu6v0q75reUPjRCGrqki5t6OnxZ6+F05jG58r
rD++ypV4MBmQSlKb6Q9mXrlbtx3tgyI8hF3NfwrLQV0MUJbXQ41jupX0uzjr
e82iD/XT4pPKC173+03zg/NU5ExGBJ0WoLOpsxGrrZICKgqxfmPUnhpfvd07
sDhuWrU57t2Yf47FsiZVI7Gusn1z2rGtdp/NXEhGRnacpkyxYjX6FFg6Kehx
ZM3R1WQ0Wq4RRkASQs/Th2q+LpU5gCFIi1oDi7IflxNQovbxWw9Ied3tavYx
iWRsHZ9vG+qhJucsfjTiRAt/wJMfMHT18xZycSRbS30s/HwnbjLLl6nUsZqU
r3KYsVyyQt8oxlDwerkiF4XIvLwmkEqLxR4uRIy3O4plwfMYv6eBUFjgM1kI
V32guReGl0q9vHg5XAdMb/+CZ2OAu/C9WV14nxL8mqdwSasaWlztYhAQb/fR
lTPLRUcU9bR0DGXhkJagDV1PuJsV0rxliqCPb9rs0Ep4+q3iNKXlcVNY9wfl
pDAhGlT/FabnCN1i0CO5dlUR4K1pOx/miPEDHVw3NVlA05hFEO8mNtxRCmUD
VZM3YQRHae5L9rkVvlmb9xdyRaXXD0bw6DnkOkFGr5gyhVj50WVBsKNMsWEm
H2H1r/YoiEaGdJNgadXo3EpW5V4CEaptqDMW/WPQk87x/COb5aBh1e9cnIxc
v6kjN9x6fi9LMD/aESfrVhPjeQBGyZiXuuUlqWQf35gJjRBBNYsY87q6BXrJ
wq69/s+Vgdero/qHEdUZSBXMoMr4tnQAUozFe/SOQ4ZZGdGK2dEZO7EPasDp
l7bjgergGPzsruHUarfnJWNWFkUi+4hYwsDCziowqZMMZmMrRnbvFTmztt0A
LdleuVgNJKtRybN/cKpVESwJOmcLD0hNOQ3mcd/ClpEvYt0+kaC4W1Vq9EGQ
4lrQU25Co3kb1QAdN1nItOQ3mg1xx4cTTxcKqku0L62dbYsvxlqxOfkzukOz
6c6UVk/UyZsP1bs7UZCwMtgp7wW6jmui/2tYXDYdZyS/U9ie7jVMYq92ym9Y
WrKXJtvt++TVnppc8ksE0ljal2SWhv9YTpYfQ03igx4bp86Tfj/+49YY+J8n
TT3gP8V9mAUM0ixpTf49m3TVJofAYc2NvhMLxAhCxFyW96X111OZkjUSKMBd
l1CbBokoUI8TGA7RAR1MNudFXR6zJtS3zd1CwZS8Chmio4Op3MO5w9ioQN7k
iZpANeadCW0XtQVVw21mJxBYVlT7AJBE7nb5wNSFw+h4s0baDDsrFucpkRod
L4LDYiBPU3b4Xym/5fnv7bdEfqlryLX80kIY8uqPwTwtp7muqKEpBvIfhIME
RLPTp1Vd3sjaGWam5G4tjrZWHH9er1glBWVpDMkat8Mri2OIG4EyHGxLQaOa
KNFSwmIjpm2e4TrAH5B1XjfWzfSHTURnVBo/9gdoXP8w/n5x7SuEVZdo82Oc
HI3NHhThnl6i6w1Hjdv7BBzQ3Sygq5iGg3AfHARkvGU5St8t6HDKm9SSddb4
ywR3vBVP+NZ0gDVjtq+wuP9TA0TKnUJCV0ED+njvPHovSoveK6FHS4hHPoP6
0QgO2VuUUqUAu6to0itcn3O58am9tnoHJhGZyMy+h4OXoHdUPph+/HRH5jl1
O0u/bNt7MrjKImk7OWdb+YJIDk5e0GSuMrnrm7d6LFmqNCPKX3FK6yocbk0x
q4FfSwfbifMLanFmrCaUVvM64Q/hFF+2+Ds4YeNqBy1LcUd7wf+NrJ/OovPZ
AG7liSxkT6bBXpDkmJx6FuyYt9NF3WzxlSDkBfeb+wA1waSMwHT6yIpw96xo
MXTWRtJ2XmyRGyGGHHsXGl2Wd3jal0tCp+UVOsqOrHpxZW8t1u7/hjC/tBkO
o9CuTcAcgkUczK+HWnQqqgYu2LYz9o6yIt3ythTVAomuPotUedNEq9JIAVw8
mBI3aRAlenV60h7PrWpD27RmqFg7zDn8+YVIKhWNG1/P6BBg9jHwlz4rinfQ
IJ3rXoYKVLp/xuo+YG9iQO63EdAMTbxCR8YNvWllTJ90itJLeWuyKeQJYasZ
eW4GvOVQZts1qXNJBSbEvT7+39+wd24OFUBQdic0tMHicdMlyKbJ04KB+VST
pqrEZ0nUfYeIpT8PCjIuLZdEgv4uupA/X2shTuVKKRPIiLe5gASxbdWC6/lR
kiYtUFredvlxX67R1jHZ/k4LslHcfRM7y0cgnaFrlQyRHq2Gdnn9GMAWqdTA
Ksb8QUAwlFWdU3zsV3cGADdL7I9gTQ8YVpqVq40INm8lm1x3fdAhV+noG7lD
TJr3QsHeUxjQzBF6inszD6/0lCSViKJP0TcHKuPY944N2bUPNOM6Db9s6+vg
y0jUGz51HyTP1L0jzl0RBXqoYg9DGyokQC5KAfYf8BTJrk51rmYXuj5vP1uD
2rDIsGvOwIr8bTSBirHVoSPa2iPepwREg93bY6cbdJVAlVIDZgYZIXNDvGTr
dY1hYq32zKuexT5vOY+1zsK5LN9yMIaZ7QbzgCy+xtir+l7EXjeHdi1JD6hN
WTLIOPG8mNqNn1GNIqNDc5ukzHcwQ1sgZkt18ufiVXEDRNM6FEcOCiZh1U7q
1/qrG7VvSw48uNs0aV3167wSNlrYseNf335rIARkqg0MSdK7N7V7juVZMf+h
K55Wv5T7yx5DjcUECa9j3MGM88551/rm9rt0tgjYLryoKtRA/bP93z8Lzqx6
fkXHfd8sCbnVTjXnbu7DV9lVzuX9dP3sDYis1iWP9sjAbd1orMJzuBuL+Z1z
rb+EoREQuaXLmP0Brl95EOgGrAMwCHR2yoNdrvlPKcMasQMVFCzQ3EjlySJq
8XBX1Dx2JVw3JvfPYp3aqgkfTMFmv01cjYlY/8M/X4yUtUrB6cWeL2HuQ071
O54tF3Ss8D1RHgLSQaHC2vm4g7d9ydgaFI3J79Yc0Fih65TW7TH0C3OUyRD/
/dM4MU3CYGCyPqQnt+utaQMH2Mdk+iySzr2vx9/YQC7MiWItp605T8ULO/86
7J7RbzpmQ3yjQXx5p1wbWjgJLrfe9XgqL3pac1DND7XI2nikdBkp0bvEfFFT
iisLMKEzgMzVBmzV/7ADr/Yy+kNmaC8MomIM4difAv95OEUYcGMH8ouWbsso
J3VIy4N2tQemRZY6JtS/cwpnY9YQhd4FANSk6vJrzyooQnHjhQFE6rlFH+j8
rPVHVvWaeRXELYd0ENuEAHL3P+RQEFE/owaWpd3Vrb44MYDCGs9h2IoApXNe
DlX66/LXobAEfodOb7Fx5jtqw+03IbHdBs5Nw4bXnICQH6vYxMIWTycOVUPr
XTpFjvid0u1CJ2Y2VOVWP66hXeCgf+M8X0bjBJGo+PxIK6W7nRfe91SHD2ZI
HKocGK6xHsWL7XDV3eCRmltYRfE4pXQ92rOuzd6toyNCDUH1YbEKYHl5xLh8
aQLQHNSyl71QRsj6Lhyp7YJCd/Aq4cZHrYeGnrux5aBYtmrci0n4mxz5Rgny
kcU4htaDle3O7bRz9G5oFN/gTD3mnAUYVyaFSts5ufqi+bjQqdnxKnIjV2rh
8AiinqjxZs1KZ2p1s85i1mW/GU0Qt+i8imDjLOZeh3BfZ+ZTrFqrOsXVOumD
snLhXIRcPdLyVAg8IwboAOCrqCCE6XZjEYErg6vB0lJw3fy1WVA1p14NvpvB
5Qwyr/js6tZ8VWy9d7k/0Nja72p0vPWF1+o+57AUCOL1wzteF2BOxTaghIq/
KbHrVphqTUwefDXYQNbZzNnWLYD+eTHOayquS40RiosXwE0cLGokTZX9Kx/b
lZCwwqZUDCpkC5zDSLmpa7wvwjaHAnQD4H4dBDNfCFL+n5vWoMmhDH95eDB5
7QrSAIkFRRF2tx0Tpfv2DnT8RweLfawU2bAb51xau/7NAOUGV+GT/O/YJZD3
nU8UiosyMwTLFQRU3M5MfyYw33Ce8Un6Ck3ngp/GSG0Fru5lMyS2JGdanrVY
Do+olUU0iZhQm7qNGWCalYRtamOl6WtFhb6ktlmX2trrW939xcehPde7iruc
mR5rCwhgGM1tEevw9wdq+danMJPoa+OJzMjn3J5zhsj3FoLKoSji8TunZpNK
PNN5X9/6MG1Bhe93ZEhY5vVrhMInlgP7VovqeguvcWljCcV0BBWKOMl2noh5
jhNLULCOoZ9AYEzBTTlllhd4pvv+2EdLYdDSc+Zsa/oRmY4voVfqvpSyXl6c
IgcMtAh5QoI1oU6SUM1bl7cuVnNxcOoz5JdKoy20WjCzU4pgIwJ5y1/j7gtP
G2USgfT5fSTeSpOZ7ySaHQzOc5j1+A10FMFYcbxv03830zCBhNnauH+qnOBG
trEmHwXFndTWlOg1PWy9vzdE6Pv84uWH9sPrL6K84Bb96SNe6CYqHtJTRSkQ
AaosuGZV1jLjjyU+Eb+9EseshpmjW/iVnZFUJUNnreEfbaPFexEjCSvFa3Mx
dwYCMj5jsHEGeBsdlHs/Zl4vx/QBBHc/NTCX00TscquiFQlkx9+oJ2fjQ2fg
BZHr5Fui3bhtgCkee5x9wnSqkC5CpM88aTuCpQjP1ECq8ZFMz4UmkpMrbAzB
A3/clFAjJ5ljlJlB6kysYVxbU+ZQ1iPkdYfjC7IaC51ZY8s8izBmb+GzkB1p
kPg/q18YOwec4/sYcCMtiXso4eZLb4IRSQ8DpOre1XU5N6+1dPuzrP45XluB
6W1NSN6tWKToQdfVoavTjx291P1bKTm1gb3wg4i6fKsC87r8aWQ5fMNMHXY4
+wwpYkoSjbASMb+acREvA6jpwY/gE9LojfeXvdLXX/c0V1jSkSVap6t8mQBZ
YjgSR/w2WpqVL2TDvcWWdM288kOC2MkHNVhSTpMBkKBnOJzpIk5tzSe0yyTU
UwQ03JmO0XfuO1gpZH5EQG97AGCNPxHTh5wCjyMCUcsGv/Bkd2aBOTO+zmVj
hsj/1m/yEwT+a2Bc0wk+DzUJR20MClD4KVtNJqQmQB7U4CvWzz8zdLyafFcM
j3/OZbnOyAa3Zz81iOo9QN57xEghWoSbfH90KRicsHwoUyL5UQnxNdubu7Du
IdEx0+iR/V/xmL5GUWhxpFpidkun+FbiOJtu4Msldb6yJJ0OlhxxsE/Er1km
ze/LUNl2iltURNu2dxYQ2ud96Du45qr6LYHnzc6zzNx7uSoGwzWKNJmqzyOu
ElaYTEgssQfFuo7X8CqI3jNYs2ovJN3rPZtKFPwbjFACA4+xRLjrBk5W4xeQ
cFWaH6YIB/bn+PKB4dFqFNR0SzoSxP/P7L871Oy9S6wSGO6zoIDQjUBn+7my
YzMKtjMVQvlIg5YvfobykURNIPyACvH16meE10nGzuwBj/bmOw67/q88gl3b
zYFu+LmoacKZGXIElfPzl7O4UwGcHXUPR2RUb4WY2zWD6fvYdj72M/r3y+rR
5MQLndZYQ7SwH6JiOL3RabPWRdmfGk8MYPK/EPeO0CgNJ29FFAYyMH0FQkRJ
Gsx3/H+wfXG7GR++MOIC8lCzHTlqycMR2XNANTk5kTiA+m+4JtfZhuSOtYIm
9ZF1BzUkfvP0H99RyHSKCoqF1fHH7g4WEs+hve8yWc8VsT1AAYbmxNd0VF2K
8tG2F0FnNn/kjHEX+afU15kxT1iJXCKa1Qm/ol67XbLuR7usf9ylmXXGl7ad
+DFOODEkXr+cH58RBBMmPiQZdz18MWwmXoYXtYc8llis/tIIHOZNRmNyp2tv
gNC029WS97iPnp7fT72OHne82R+yjsGtCKOE4fsBCvsYVufGMPjP/jaqbYUk
+0zUVarDVa2z01hnCXxo8I89/saclW6cMDTtEKkHh2dbZtuYwkndnx89UhYW
/FxlIhEsFldqXpVqaAAoI+hcIvWWvuckHFt3fZ+IfduLm5X46+HCdffDTvoa
pg6nwIiX/op/yFKhbko+5zHYJlGizctQpfhTbcIaT+a+J/0yBGFE+4q90/H2
u6C5p/o4HYkUEFQMrhWf362vNMLmb1MUesQsbe3hcC7bF90ywNZ5UWbxocOG
JmHteP4+cf8vs5vllYB2uk6wYdGZ/fMu97Cc84am6B0gDTH0360rfaRt5I1v
8VrPf9RDcJj7yOsMqV7oQYRHBd1y5MXDlb/U+CTBadcVoqyUuUAAFafKnGv7
xXdlm2ksfrjO/1p1PWL2EE4AU+aLvK51DYgOVpLf01CunjkyWu1URRIPw8rk
wa71+ZgTSZnLAyUD9vkI7NKtp/KCq8Ae+FxKUzjL3bOSw0bjxpCEkz1W83Z5
snMdJJGafvLkhvF10j9EaEy/g/Gv6JykYAXVcCqNSxmV77J6ZuMSC75FPAvg
7kkPvnqcUGlX1tidHByK/L8QLtka39QVCw0eZ8oMikKOfOYta3kbKdL9CQAJ
QIUPngDYww1bdbWycy/kWtKAtG9SJnFxmeqn0iJmGnU5Op7p2O2zERYkN4A0
rcBXntnEybS1iOcMUsWvqaUvV6yMdwqWJPNgfc/6GSNKRNBEU6U+7EigXGOO
zZSmb0xj0BAWg/agBr+l4Xvw22S1nt/LOTQVeejMP8rhwRSbvRp6+ZpMN4Qg
irFgiTvY4Fpqng0/SSiVmbgMrC5CZL0UIcHCmtSpre88CXfYe7Lm6emQbh0v
XQVUq019s31Jp003eyAXObT9iV6mObD41V2ooesyvA1MZcHWmjFd2LXDoWXI
gACvXveNKTTyqVlaIgHasBAULJPHyVAHdpSwyNlJ5yq/IoY6j6SePAxdyk4g
igEl9X8kmkbM46fO7ht+1l0tkqdMbNfDJApSKlAmmgP/QQt/Vf3HwEFA+o6w
LAQhH/3AiwBgTR8gmE76P81rKGMxPmzdIblPQvUoIuNZXTERN5JqTz5MgAXA
gZVEDlW4913Tjil5m6A97Vk0gmfDdmD7N9oMY5ImWOrfmgyyRPOQn9T2L2Gt
aEXX2xZTgEi9Yf8ubA+tRKBF0Fq2RH8l8XMLuum3Q/nmjVDWSzaB0RZk+rLB
Ez4ZTiuZheKAcus8Gx1Twu8SgC4o4djiVdutHPlR2yXd/yUzMMZMmCgKUlU0
NVZKK3r3PmxR8OtsvhkFz5vkcmyaoxYRRBzQQKwY1+loeKylttSECvPKHhXL
u8TdmjCVdHfi8WQKASGWCrHECcp84HOboPKKQMH8aXYz74tWP508i8r8H1Eh
Ir1WmfsOjLjUKF0tecG0XDAQOKYrPRfAG+LAG0bjdiVWOE8T8z96qHsQA7yM
eKYQuhSyMEHwTunDFjKqVZcGJ2MD68iLew30zcNJUtmdRarSdkb8v1ZDmAkd
cCp95PwMX9zoaQRE1y+tXfGOutI+mMKVEO+7grrkWLepj8Cu+l48DHhXHgG/
LSEi57cjRp9pvoejJQhozH1pajKw0WXRkqtn+IKloJE7nxX11mX2ufWVWXvg
m5Eyn9j76hGWhZ6Uy/0fUg1ubHRSnBdDKc9iFUXa1qwONA3FVY6BgYf/HJ+o
LzFWpxQg7tzVm2OXaFtOimWgLW9MkmMgmamNsIa+l8P5N8gIpByD9qwUMFPG
cJQyujsxeYMWsK4ZmaflgcBgJLoGQbTenrd7j+rQjWMTiIG+m+ZEGbtXxdD2
OQEjJgzUUeouwxgGKi/S6LDe8YRsRE15gvDs13CHWc99AIJ0XcC0TPuJNu0Z
8ijeh9pyB+nDQh+ZdQwF+IU9esbO3CWU7oSzZz4CAE9ML2Aw/H4Ke+nmQzHi
VwJ64vupkbuGqAZuv04wGVswLWmoO7cjk6fCtjPrNH9r9LnneoVPfNvTXJsf
YEgIn0+aImXqyD+ANeir4ZpNfNW6l3XfgGFd5I8jwRd9PFgQd3MsjDNXxUVF
i1xtcEJKv6Sb+nyAD8r7O1pArgI/O+MRMHqQksD5rypyRLXRPN4G+pzOvBFb
ZwL/IhGKnJys5x7iCmBDF+JoheYrdsdfEx5N/vBuZpvc9DbiYlREokwENr5g
BkheVHrgsevnhNDolOyGRuO27XFzEIBDVNK6DbmXa+yqWFVtm+7DZuEjvgUK
B72rMGypEhBSn/6Mn1leV58m0moe9Gs9OC3yt4HQJkBv20eKFFQiT8BDiRe6
AzXa/Qrs14pgKhbUef23VQAq8PUfvgFbH+1nk+YW6jHAoxXI/oLYp7Z1OGTG
oEtaTNVzcaoJE7V52kZEy7WMq6SA/SF0lRWpp2bq7KfrKNPN74/6Fbu+8Vsj
Wdd3pxFTb7OQovOyVv0T6fKRN8iDHs858lWTSKJKeto/oroZRFzYshh1CkDW
t2QXPHnSNt+iIRVd3WvLO1tRzBGaWrDzEqzSOt9FzEXiTyPZI35HvsCH1tcT
1t+uBjcYAO324UUqH9XeTw0UVJftGvTGStCuOVm1NqSxJ4IGmU6vXuKwi3wc
+3fHE8RB3Vnj4bQGn7jUluXr5GKs6oNnQywUobXfNpytuZO7uaJN4U5xBTLg
8Y1QxB6Np7T7SO6x6LK+dFCsGVkRrFuRFg2H50SYnoWgb1nZsJ/GeTjEbMda
DBRD9p/PCWkgVeVudIvIVj0Vc+l8yXmVEQvNtT6P9b3OSk1fgdrU8MGQniBR
Oga6Uy7YAWLTXCWIyhYMHgF5hudSLHX2EXcD9JY8lc++oBk213V+DpquYnIx
gmHfT2cyqhXqqrGUrxRmz4lrbmRuGC1fLqkuay7ajIkCx8ldKISOcu0ANdfH
9eDzXB2fOQuTgP4jIpYQx7tO9O9HGIadm84a/oOJnySDEyzLN0wgAVByEVev
Jqjt2GqdmS0JDjpe1Oc7J2OKPrAIaFFQLb2UMVqRpYryGyKiGAjqARQ1yzDI
tZF79L5CDXR55koWxn39ZCPZoGi92FDCB73RG27eutbmppLVe5oIgAycS0mU
qe0TbPPKtdQchHZZDHICpiZqo5h7hfqvCYB+6NZmpfJ+rnH1LcVn60s22nVe
7wO/XUJu0/SLNMI3E3kf4euGSl5p8zK1UGXCMao0sCMYOLFZ9vWXzvQ14mfK
ok484IfH9T+W2T2wuXANxyYg8oEJJ8uZmesQ/B1klalNfzEP3O8NMSHmh0xp
UulGMsWinBPL1nkG5XUIVcpl6fI9POk7ZN7dP8dYopjeLv9Dk6mOnJAWFKWF
WXqhBOvDXcJVuMOL37eLwhwlusVwluG6B60QvigJt+cl4XMwDzL9iWF/t5+T
RagKYix00KqIj1hgI48gq2jLLI+UYiNV+8BDEOGUez0HIONR33zJyB58uvXB
haX+bkB42BWdIviJzU7R2kZCkwvLjLBjKT6XnNz6MMSYw8zCKqHcGo+5uoBA
3LZ8kNxEBAqMCKOFRndUDZwj4zgBMUVFE4Y6qObo1x1Bkh0w17d3yb4qgOff
FVdwpF+yDFVfc6f+6ir4FunPzmvU/ekwMa1WFEcZiIojVcxY1LJ/8JfcOFa3
CuNEAXYkYtVH3F0isv4wSVvhBhnVZaI1PniiBzXqdvfRNUxClEx8T0WaNQqx
LbcLiBLDBGBl+/aeidND/VKQsazk+LNsJqSx+mFQ1YUF/Tni+SiJ/FXMCzus
YXOr7dpve3l+t1EPeHKtARZ88xt3N+mLa9SLVyOvhOT4pZS1NHTUjrgIUHWf
1X3EWVnO2lkXV/ImCag8+NoGF3RBAtTEN6S+vqFsPxvbp4J5wQZXuYnIGusj
V+nfYvmeeO1xVEJjay/9alYzOstx13AqDrwjWle7fXlpbTBKmmnpBbilkggj
6sX5ToeAjYW93KMiC1CLR6k5z1gJdZhJYK2iURnHQcYTmqee3B4XbBrSYxXN
IqQQdzyuLA6sCcYmOj7c2GXL8z5xKUHNxv2lseXowRSCm1bm0xB4Dismo2D4
TKhvXnWdkomRfYOIj2TJg1TIzoIRKyvmLQWlDHf9evHHx8tZcYUKG36a+8Zu
s9dPyEcwRyxo3zG6JXlC6vbaWU27tHIdzBjcTtI65XIyrlF3F09LfGAZiXhg
VVpOIygkme6QSOT98OI8f1Ghfb+H40ESk0jn0lvQXjCxsDRWND8bzUH+5sq7
DFqXb/fmOtWqYYRgj2aQp6/fPinllJ1oixTvhi4jLj8bYeiulWFDGfDjLm6i
MfjvJTf9Nghy2LbvlGhBldy8pUrt1wfBUt4pHBC3ltBGHdr0DOYKnz7VtXv5
nSm24GgnCkgygFBlbX3288bIpfKIGJglmvzJkTU1S8y+zubz9w0hzwOKAm5B
eNw+Y0M+H7n/2kB71dyh2FDl14F3lHUwif3+FHBqhNxrtI1A/pEjlClYRscm
QJju752gbuQxii9EBp+cA5BC8kctWRHhdnJbLr6TRcQP+ldlTVns20Cg06/F
NeMpcgMVvHMBMdaR32jBiZCq2aUqwkHl3hMy2+nbLWMmHX30rDJrWBE5EXTb
0j8pqfiEtnFKD3ZQq2M359CkN/ZCzK7KRJdn1KHhZBHoTwK4ASX6EPsCGWNl
Vjd2dWruuaEzkHsSzTHf8nVOZnOrm6dLXeL7G093TnhKBRqT1HCpMC9bi51V
6aIgOPuN9uRA7BOfKkP5+YDJ4PGFEXvfg8a2D/ewww2F2nJDsgWiDk2phFdI
T0JPFKZtuZUoJh85zg743Qy+e44f9wHq3x8qT6B8qxB4Dif8EC8TC7AaxmVp
VB3EVxl4Kb85VrLwBxShiHCoqIJ7aIFC81r8+moeFlearOz/H3NgDGVygRS9
DZgTupWaP0F+AnspWM9uHnyk3rRH1Qu87JvsiLzs+epHRym6e4IClJqk4NTc
Fd5oG1kE0g3G4i2dI21hkJkMU+xYI9+b2Bzt7BMFgxv1GtbcCO1ANwfPHEL3
quLXf/z/FA9t75nn5BEk7xPm85qimZ86LeXwz64ZeC5Wc54j6nXeFRUfTZVE
m2Jq1FlaI5Cgn9OKIPH6VPuEN3EyQEj6TbVM6Iu2+o1bAoRVi/PHVTLKSeTQ
KJdb1tE8poCi6xB68CWXerU1JbNAj70W7tQ8QqQFnh8LzClHFCF5QJ5zSHNu
SKboNMHFOiKi9ceYAEk/Rn7l6Y1i2nMu0CbXnfbbFPTEcaEI2xydej1K66Ih
IPj6ivgJd+H7oTHICR4pS+kj4a/IDvJ0s1QVH5irLFAShylhOFvEn7Wz68ga
PfNtmAdUO4dRGICA7LJzKgshiu3UPECbwanyhGI0+1W52AXZcYJ9jr6+RcCh
G70Er+DPIl6OMebG+S09cTWL9+UoUtpBozbHMGG9TZzDLYskCQPyrnXy7LSn
hkGK6x2QgYweoJfDuVPrsY2Gqsvt20NRZ3fEA3yETTIFaq4mWpvO0aD3G9m2
fomKfSNldseBEtuRSwDkPzeypXhnAgYECyBmuF4GwZplOuSqTv6fzrAvb6Ni
xiLdbtQBzmZ3aeYx24DdzQi3cp7R5Nz2JgPkaG07HrzuKZvivf8eTLvkBb+F
1G905pluD+Hl71H2+nHTH7r5qCG3OX2UU8dp/y2+hhvNQbRDbE5OBka+KUcG
ipV/IYf9PYzBtdDFTqr28+keKIJnZheTexzqNO/zSdmxZIMkB14IBUgQa0le
uMRB6sBNMAob0f1bul79jGLESHu1arcYvoXAgmzZk1p7nylbd7XWJpN2DX5g
7qEHM8Ynr7Q0mIhuk3TPNg9bPmhbjWf+FFe52Si9YmU2h7QC8u1Yg9Ssh09t
aZlZAf7/xh6a8IdQkmBb0jabqjTLj5p/GCtvkwxfqGd526AhBfPFVXp52fIv
6RKZYno2w+Nla4ZMrQ7lg1d6YkW45s+L9W86spZ0qQrOBMnaA98WB8u+yCjL
4eYx4Be7UMprDMkyEb3wWcJFWgfx/CYCs6g6ZyKUXi8e7oCHutd0Cq0vM+te
tMODVzUu0ECdzTAkRLs1A2IWdwbMHj4RaHURM4qINTN+mcybocPvHjNjvs6N
ANTcjNjisTUV91gbfv7DguMZwjtuFRmEeMVcix5Od16fQQA78up+qaund9/7
uqNyKeiIn/odz4tcE/E9a6Cyk7kuJPvOi+b+HqLDZC4r/+fSBSVvh02hJeHO
iLJGndTAEllAVKVU5VmCslpoNnadCS2+K0x3Z+RBwjpaOzl19rLxeAPP0S8+
1Rp7TxHnFLp33g5FwMYddUKXR4I9v3ilYi9Hbzo+ejsreRNCggDcLbibDnb7
AUtpHc9J99cCfU7rpKNLiiUJliAtQcE+/f4FYb4dFViEAYRj2MvoFDntD2El
TZDy6ItBmcxgCDgRxtwnrHaXLXaliof2qrtIbwBj9SMSEMoUW4q4cZVVxRbk
LflNi2mUY5O+yT2kZwJW1R0040ORriyO7C1TZbxxeQYYdAleu25PNic+/lJ8
xaN6dWr7vwzMETkx9d5+7rbsbzcBOe99PA/IBizivJW/6VFasOmvqxPP6FRX
yDaQNKR9qDTXOjNVFSO/Z9L/vKbpItYZ8Q/ILaVX6DqAjNWwIc2LiRr3gorG
VLywO6iYVytOZhparCAeazmoDTnQGCmuTbVh2mjV+iMCM11NrC4cr9/KyBtG
uuv0yMHvgDL0SPNCmhVKeDBgZcMUb4MBJUZ/e/QHVadzI0n6NgmymHFrYIxU
07cVYGnObOlsJjPnM7N4O+7lppZ4BZ4SKJxK7dsbuSi40SU2LB7MjEYvihY9
28wLKKjnmqaIsZ1dGuaQ2IJQHCjr9kOWAab/ica205JVa4QeWeCZRO6mqlkB
DfCwJzK+zbxHvSxFUgEbgZYABtM08glWDU3M1qI3pRNIZYfSff8d6ydQz3OS
6CuOdfwv0mmaafeGnHemCA0g5PWJg9rqfpS9FbZwtrWMKI5MVUpkDlmo6MGN
NwITZjO+n0KxhzNyy75UinPqwVYQtvr0AbjTjjupFsD+2fSKpgA8I5NZpeJz
qxzaE9hyR9eH1N5EZ3Wz1YQvzRnHkQYT6cx62TwMW6CXNQ5/m9mTMjs71PVg
pj1b0BFZamrVJdzeiw2iXtFV5tawXTLifnOjfGrL/LJX8GfhkwiczFheMgJk
+2+Q0UojJavBrQtyDd31igaHquS5p/e+BweCA/IsXMZ9oCAhxgoV99qOiW3l
bd02C5Fpe0rpkA/yK8XSKQ0Xdp3Ic3yEhWUCC6IjtgVsGgZHkvlFZ8Flg/1/
oSYsQloBhX237GNNLuPG3OnlVF4OYV0T0LAtZC0EGjd/ym3Cl366ueV+Z/GN
NeKQuMCiQ5sZHIeHJOLus/IIFiqktseM7gFZtLL0DXPdLqou6OnOp1nFPUUC
g4Mh2l68TH0ehM1GN47mvSpkE0EsL6Rx3BAEVuiljRJytilnpOEyE1xkPtS5
4C0zrl1vFB1Kgj9x5aQ3OLOgZUBpxjLDUetO2Zkdp0SKBC5skZQbxlWyL+Vj
Od2Lfm9I542RqcYshAlpSuea8Gf7KJxVjRE3WSPDUW51eZH512qJaNUHrtvG
A8nN679dGkTqWOR6o6/EQLgue4ihE5KdfbaeFu0ph4cvLpj7Pj2ZK6ZD/faG
HhKG48yrQKsSG4vR7OEsKDcoURr7iifF8KaXeSILYMkGYTS5Dsl5E1HPxpXG
9Bu5pqatCJ69zz64imyOmyj7Y7ZoQicwLbB6VrLkzhMksnWqK4n3hIHyPwIk
oEBxoUMPC7fgJ0pUjB23tiHC/DMDi2p6crE3/45Efg5bvulzkgABkqPjDi8w
OAASe9XnZKyrbx3640pswAOmGqrdv8/JaT1ukf9WdRyjuZwhzE+j9uzA93VU
0TTTgz6kk1E426QvTGPOPuMfkTbFriDdbO8T3Uosro4qc9KruPnuUx1R34OD
Yui/nrVwy9VA5SdvK01CTiNYALr8KQJumOHnBZX+lUmK4raV+5ErTEPteaTI
GtiyGqlvkD2R9UAElC+o/Ew13mLvmuliO3XemQE9gjuWlTSjSxKsX58W2vYM
+huAjHJixA4eGukAnW3SOg0N6Kav1AWAdjOfO63/LZv2aXQGSYkCrXVaIOOF
NkOJEBz9DbOKF9rxVIAzqg2SJfjgDFooQ2N0HXGux5/YVemrGhxgS6SQIaST
JIHs1ywSllLK3kBIQgxx4RNyjCoF4TYGQ2T0HVrdsVNn/antLbnovnFzdaLO
6aCGOeM3zN+tOmBQ6xvYPfqVOnbTwVaUFjDPppyN0YNj6JxbMHhCW7cgzfu9
rEcfoNLBgAgzvKeun/COCkMy3fXfjlS9iFzcmEcSzr3vMhjBuwPPfQLO+4Bv
ODygC2aIBNMHbql1UC1xAg/nceMSu4u7Oo20GIzV9QmeNdj9dU9O1qbDd2Br
qbh6YuYPPpsKw/6AD8HxPHUYRDeWaRfRRlyOq6LuPCrDCiFVLFTPlLA7oLAW
BvhvHlD7p89LanLWEFi4Tu0wF915rGItHsy/eFZyR8sc+H02fRvXtRHqVdpp
mK23s9utiJr/k3KzDmhfE/fpLrtvaFhYpfTMSf6qMIeM3dUZZtpekqMBeuNH
X2HOLtSPl/1J7AavbRn89opRD1GbgM7gL0BTkXzEOlO2ykH0au+scFF4Zt4H
gExKqQziN0cWjcUMw6hSZdDpcj6YduZFlDJy3l6iGuyYSgL6MjuGTFuomFcC
hkfVB/JVEgC+eMgDSErb3yDt/mIyFUMFecdJtHKi012CcJVnwqcup93ga8bc
8tT+dqsOrEyvHctf9b7mPFnkAtvCND9ff1t0CDqb7NQ1kVYl3D1KOh4TXPVK
nPtekKxkSIxkzCb3RJJYMx5o1bWWqI3BIKjkruX5ae96JqOxuaNl0Ur+OrLY
dwzGvunc/4CjGC4jLfZ0rLwIPC/SUXwkZUMOsWqQvUkm7Z6iPCvTFIME9r04
tvckrBMZ6RffzIUi8ggNiqZSBtshQLcPvGI7dSmZhI60rUI6f7pmsGGn2RQk
PdSQNXvbf/5LOTwhpXvDZHCG9TUPW+zQHh0FNLjry9vlTpnpBVzorz67BmN4
QX2ZvHH81bkZP8LjxJI+quunzjoF6Drp3o9jU5FmuWiEux97JMhRMjD+8RSI
ySaaEJKKwl01gRQa66SXN7Rz0VucQkfzsf/5W/cSf2RzjdRib/SkEC+4Gs1y
HkyN0zsWF12nzX54LcXAyNQckY6tasMH/7unXOmefzu+93K+upT6SszUfwKb
8jfY+9hMryv1u0dcyQMWU2WuFbebkFErtr5Gblrv3yex3l7W8abXePawnV6h
t0ZG1pbzqt3Lxt6PH5OpoVQHGsnOInvMkW+lMB5lIQL2AYnSO0gfQY+FRjUh
/b4o5J3glhzlb65iWXk5kLt1RdvTR7WqrHIbpIQXsJeUKTd31MAWsbha+q4f
XfjMVXvU/uqh4hil1M2CVoeCzlyiUkKfsNhs2K+Y+tYbpNAtMUne9mOQuNNL
GnRub3b6RVRd5YEkmXQF2djZ1cHE+UngAm6iRi34ah4mmYm8QPxmojolFkzM
LCn/9rUPgob1v5zXtS8cODusdpdPfY0DpIwh6TlVW40neez8AIA/9M4+/rSt
anm5/w5ICxacan8QKYnCzEkyuKub408vzOyd1FVOQegFRooeI2yPlStvR2oc
ItJFrsd47Q7BHQChE+xVG2Gh8nzaHYbF1DNE1Wc0olbPYHg6gJ3evkuqv4C4
01w6TGs1r6MBxEy0z3ToU7TPG3DiwZ67mEMNr6jR9CZs/nEywGG/+TXflw2g
d3BKSx3xmSbjXQflrzeOsR5hUXGnZDTFV1Exv0n+j8zN0FcYbrhlAyjz4isv
1fivBklnazHGDQy3Dk7g8pdA2kfvLcnA1uUvvyyjTQyEYvWKnmsp/qJrLJtF
J9nZ0qeawwXaF5G4cWFY/QXs9Mvrfl97bfmCIhxd+V1UXc96QfQWRXnb4Vlf
aTMJ7pVr1BX94j22Kqi8u0htQsakJ9n25WlKR9Th6JSpJfPKBoSlUbMI+g04
Qav1j0/icfB1EHXyBIu4xbs+UdOAWVbLCf8JKZ8/Afl67gHMCfUh+8a7imjr
XFSu3NoWPnTnYcZeRBiUNrpmz69NlxC7ZXUiSELxjU6H8F/AgQX41eJuGybm
a3/rFVuqFj5ZP50GzhaBdksbeWJDT5NxHmtScfHJR8gJaYOJSWv33hCV6JwQ
N5lfn3J8q33kTVR7GeCy4I+s2PW0504sXoCbTej7ojHwOa4lZedhsyDK12gL
PZR1rzMMpL4eoVsiS63ZfKW3Mz35IpnRNSPH9kCPXD1YPqNTcHADeJG7+UXl
Mwg6vNY5RwLpAUkutU+i55iKZmCGaxtaFsOhYa5yLP25JAL1e1ID8uOGQf7u
bss+toDoCMF3OaZRKmN0b7v8ShLVAn/ghBfQ83cF4v5zjjlkkVEMJt23prcX
ddddvGSyA5OdzjRjJlHRGF0w/Uv9EYce5tqvrSR+Rqmr8KW/0zrxGG8cUQnX
EjeOVHzTELcON22RrYHyl7oeCHILv8U+ICaWASMRRMLCiMNRndEEUrLVL81d
BwvZ86qds4E1kzPtY3lp+7RmYWxzYFaCyUoYjr0FwgvUaJn1Z5wa4UqxdiCw
BWuFZzW1HZZMjUf7HcmM6ys9k/MPcURFbLo8rDlBjni3eFK0zD47gk4MW216
ApbSm71OMVmDdTTIYSWLFB/84mb0Ma91V/z0e9w249Rw1W/+5He1M/sX9F25
xPxn/EP2SWW8KXN7D29xIUXoKA22yuPVD7vU6Onm9m5PPxKDKuwqmDNl2u9A
NK02nxtoGLY9gHzMucD2OOGtlY27XKm0LJ9CnxV1WMcLqDdE7CqPyyDIW9nM
CHrzAd1rHcVVkkmycJLFK3gNSf+pLUxM+odfIumbej1EdPOfVPuCqpHSP8Ub
e3B4QF97BOU8LNiZ1RlCZk1GdD4b6LlzqDWb0hqOufzScKzwfsuG1zB1jRSM
ynndEuSoUzLsjJ0al6N/KRnqEnwUQabq0tsG/DSuwYxPuAwu1IEpCibSniZu
gG91PBv0+O2AhWYEDEKcQw2jjAmzpQ2n4a0dDjfy6RYpnqu7iN8Y7Sed6KH6
vLiPkE+kFcNIfEGkujx38vVeF2ziYICOFhCjpFI47wgwHlxCuuUR5Gk2lXEa
vXNiiOWEyQHYsSOj+9Q9WfrnPS+fBo6v7jdqUj/jLoD9hatNGkhoqGeO7ezM
efT9tcXpHnV3ZyrAXepgsaxSLm6i2pZ1oJYGejvfUSM8GhByofM0mlhX30pp
LfPgpK3KVjKm+u0fGWQzg3+0o3rQnmT6fWhrGRZXyiAxqBx3R03ICChfJ6Tk
LutgKnieXZQkpSMtMYn+R5gu5h4h7RqLSGhYViYqQIE7N0L5ixN3VTLNWjIM
JQHOs8abVw0R2L+DyvKzxrz/NS9NIT+3lGhJqE/OVvud5bFZjOHlbd2nsZnN
S+tEyruQcYDJ79NosWMX4WNKtyOPkYP9u4SJoBA/Lxetu5o5EaTV8rRkXcHm
dLQxD0mGB7ZMkcM7bkhnySNh5e+xSJIKj8470wpgwjp6ntwMSX2aJXk/OpAb
hRLtWprKIj34lEu930dvn/9Q0YxCKUCevyGvrEAUC9vsF2SrHouQp+eLDMCL
zbOtvWHfynpxFb06QoBYItcNsX5UOek3ZaVDZ1bntdeyvQ61vANkIDaIot//
Y44+rgbBgNdU/VC2+TGtqvqZmgvRl5GWvhAS8LEaEvP7Bd8Bd9xDO3CR4Heh
BfxYZdy9I6+KpWKVE24OQxS7Lor6oHydkdsEYNCwUl70E+jOfyJZF/KvZSpx
apVuah3G8G29266TLmOGMgROYkzkytFW+L7CJ3Wj1duz38PNygXFjptNU1B8
QAMGiwbHEWE1BzuH7JyxP0Z6mfOvD0nl/WJw3DosDut7zBrEODZeXj0pr800
G2th0jw5gPfSF2FSlVzBYAVQj3heDtLU8BysY47ounE4c9CqK37Oqmzkt/ba
k1Bo8rO+MB0+wgje9w4lRd4NUfMyuHVaozPmprNgKVpChmpYy4FDqrU+N39C
/6p7yb2MFNjrtXzB97rxURr2+LyKMi2rB+XypaeoimSTEwlylRxeDHXn4BaI
p03EmQNdoK4tPpnBJzs14d+K0x1shUl3rV0hQc5n3qWaicuJsEpGdSMYUglm
QNrp5I6Yye9rfX8Mrwg+MQngP1fmvc0R5PUIl6Yujoiz3QFM2LcNm1IxyNn1
hRovuIa0nnuKL8omSxu0aG44b/kav5LIBbCeMmUEt7lYyUAvxSCltlWknjTZ
AHHZsVlKc3QhIfluY9PedIrf1l7UKaItZdVIqvmQTcDOtNQgGrPljO6lt2zT
nucpRLl5JzH6PUZhAfKwpV2c9EFBZ5Kseas4XvZyK/+0Rh4/+l7kspDHBsBr
bCZpb1sp5vKGvZTPaDwcIAtodTBjtOpnR4ee+Y/reH+Q7/6ZJYQCt8ZaE0jZ
wDhZLh4egzlc5f+R3io1cSqLgMkUGICVEhPPN/IhgDTtRGnW0Xpvg1wxRf9Z
HsZJaD7bQ59D936jpnHkqzLs8BMpyuZIvE33Iu4Nr0fpCGEdADuZQpHPNaUq
pWTjXUEBfSfQnr10SIXiMdS24wXH9UsLPfDsc7tmSD6rGK8kb1EjRI3VB02M
18eFA/aQkxviQ2PA1IR0puZIoVwilETpkJHJ0jMV3JFW9LVid3TLnusjZTqH
Zz7my8egbLwUhmDMt0voxXtf0PpnbHMc12Y4Z8fJ9kmWNsq6yt3VjunhjqeT
Hsue/NqTl6Zor65NKETW/sRFWVDM/K/cPMdorbBa+zJ7v932rpvZdrrjgRYT
E20GAH7qypdxVjcGob/rYjhj1aJwp9uua2UMbE1Ivai1u7sy+uT1iWt5Uf0A
BzJ3/T/onDblAQF3rNNe1m8Q/V36Eta0YSy30EvO+Jzj1pbSp+6cN7I57wbE
bx/+W1LZ1XZKpeBDLsrm/AHL72gOmvpN2zUIu5oCbYvKCtb3w1xWvULs76LP
LaYQ9djjoTLp8E1E2pp8dUO9XjQc087njHZIvMVtZ22HV5fTHJhiEMjsDVs6
1Tz1cO01LReIpzo4D81x3pUJihPtPfqUo/Nf3Ft6b8swYQz/EM2nmWN13q4i
Ty4V3p+R8E2xtZYEUkZbhtnsyrHUgq6CU0dTEUeD9GdTzn0eV/hMcXU5qfZc
PtivrjVc689xE4zgDrLd/GyB6muHqcL+2NYKZ0EvxlBZPdFlC/Cq3f0BHLbR
0+Q4puR93bXv18VL7unDkMs3sBOCPOpiIJ8P3zch2H1gHCZ2p4/YIv+p1PpL
cD7wouL/grokyUypqOs2y9KXg9bqQN3+CPPWLrB/b3cUUiGeaMskz/V9oRxp
rc+jiC4lrIRTfhydxzOEFXyo7CpW0lE285SfAPUX1cec8lOPz4I67UkvJREe
nxIenak4J4O2OLEYvwyMHnOPD+hZWE295yQFdrYq+ty9cdmBLLBJLetDC9cI
GGO30F3eR4CKuD5tDvzWA/BTaZsbALa59oHxeqpteVkCl3lgmc3CHY9KzeRx
vMcSmTTcN9YCAXEuKFd7aN8wWkIRUmTW+dUw9m2uyjB6O0Mx2nAork/ZIEFX
oA/Ld6ljp9sUMwwSb7E1QwhoIadBbHZ4L/RhubvzvjS7CdsTxtE8UaBSPUiz
HPjk2COfWx0Gg8PpqtUx6qP/hvm1ZXQhmxBnx6ZQC5p2fEATTfECjSb3hNsj
hR7vQaOC8C/M2qmo6SmzOgm+2NoY2F683arzwsul15zP4c7O/On2HHLWypyG
9u8zGtq7zRaV8USU/vUsfFfYZe2UhjKLq5NqikSACRyyK9yObG0NY0yl93/M
Ao+nCGodqbm7PiVSWnudomAjmv9mjaosmlqJz0UmSuJwaywzGzn0cqpmIG+g
c41JzW1pNmVgDG+pYfaW38/md0Ww+UB0+dWH7Xvhdd1DAw8WrlaY0VViOWzS
bb3THJkGV7cxvaVJc3qTrez2NmQfPhI0RReEp1TmLWSweeELnWYEmSDNn8Xb
Zlaxye+PdZgqYY0TCBfa7YF7lHp90ix9NHcTnrI+LhlbnQ/Cwwo2c4ZJ1n9W
sAnBycFVDuxe4MCafO5Q74MQtk2PD9A5pjkPR5jXYJ1mOHXPJjBGRBXx1hVh
TGNUAoZX2HW+2kGQCr4/V0FG1R4OHXy3/677EC1XbPQP7McihWF3vvyziGzN
XO09PWo8wObdp+i+SGN/AQCqvJyI6Qidec1/RePSYSEwU79yzFCWj4QVx55h
dFBh5PAj/jt2NziyYHYOrXuP7GhCwieMS3dy5DxDNjwkgteNBINYZp4bHAUU
FKiJ3MOWeLr58wimseGK+INxvI5Hn/zE68vUY3L8iszgs5tfP4zoQBaQhsrO
kMCD8Tl2Ukyo8dKVGcSQ383fno4P/UtBU/OxokH+bihG/gxs8pWz+YZNh75d
wnuQtprkdfkSnzJevg5B+ZAo8aAhDJC59SNXzTtVf08WNylXjtpJ4nf34/ZY
6c50kenEXDOyfk5cjqB6zpy+Kd690nYJg0WxmrQ14EL7eCWiu+q1xxNv8aMl
pq6vKkvDes+r1BRR4PTjMGs9QnxPDxZECwHTE4SRoboz9hf06UEZylxQPzdO
dLzCW8eVNFNahaSXR9/MrOL6t5Y8RXnADPd2D+G1X3buuSJQV+C2fb9WH93v
/08jpgZLjknayohHtir4p6mzC6BKSZuzendhWvvlr/iUzeuuL8jLkCP7PPaX
q4Mx+Z4xlSzoDNfEPxJav44ZW7ZFn3aw1oWI7YnyEvIr/f/h4eIw9dpTFf1w
MufnGMoruBRcc13OiH31W6WrmeaTPnCWCV3IzrFs5BAdt2SP3eE+NqWswfQY
hFdRYNYdNdnZkOVYenx40plFT+b+kiyn/DZyQepj3wKwbsNbGPoSFSHldqjC
tobnFkqdyCuRyDVoeiH8J65MRR2tRaF1eeCXaPOGQfcP1w5nh5qyMYnPREWp
d8/UQ9LD0yIm+rxhMEuUAnNpowPtcxONBYUB88DtM/+2YH5cb4N+/1FPfm6e
6zQ4QHzKwFVVmBJWlRcej/5MCGLjWprLDKts37cL0bZrNjkBT1nSZAjwXYok
0ofvSwIsz9J+tCg7cvon/pD0UA4gB99RaQ2nu+xVExurh0VP/xkUCgPsZS/0
2kMg3ckno0n1s3+woa9nM5Y8NhEfTflE5zWW2PvwemKqBTV1qgjNrUVHUNjE
xklof6HwFC4Kp7gzX57G76AzHL7zsZPardth0kVrd7Y7V8ekmognGUVpv1CI
3PjWY7rgQs85ljpn3gpvJnQwz1FrM9W/LpV3fWjK9v1N92a5leRwkgXI5S+M
d5VqVxZ7vQz3yS7W1vP+0KZ8gD27ZlzCZx/Lr9Ba3QE8qgXsMJdHrGOnlJqD
Do666EqvRUvdlPc5/a342+WnxajeT9ISvoO1zxzSa0f9Zp/TOUHbyR58JLrA
HvcwgY/JFSiBwCiWKBWwYDs3uIfjcIn1HMyveWs5+lXqTHPv5bVQGvVwOp7o
GBAJGWV7Fzg5nIn1ZAJ1ClGIH3jElbfAg6dNyJC9agiYFtwrHBBu+Y68JI2R
vrC9bf+a2vrmwmnCsOf8cgLMSyc1/6gIuLS26c5pf/EpYLblm4eM28RYLBkh
GlPDLjo9G5PooY8y4pny4zod/K8mbFmQ1fczqTSV+Ao9wONNpgZOw1LYaIlK
g/O12Fgrv+UT3ouduL/Dlxi4JA8FuSLmpyDUSZSHjO015ru48asl/ecy/+zu
peVR33s/4KRgDg0xbEF+3jHg4iigsD7aHjRjz7IlwU5aN7V+RdLxJxPZ+enU
eA2DO/8mO9dTfRgXl7u6zajq60PVcbfv2n/s3BQy5+ySBu96eeafUn7qL4RU
yXx98n5A5ZGlddq246MqJLJ9V+HgMzeIq5omgK8p6LqIudckliDlTtBSaYFy
vkexymuzv8N+FBhKJPjcMKArDLUbHQissf0h80IxL8lPOcKV9xqCy2umGzAV
PlELeGRvnAZh38MWIh2Mr+25vJGBh3elV4IZv/fEcig5bQ3mpFH7YdQZI906
bkLvT+yOAgOg/dMoKNenHMBh7JTbhMPNn01k/Hm1CoBK71EgZCdtD0sZ5+I/
E12d+wV0zy7q17Lk+P/Bme57bbIZj4vH/h2ayoOk+uHESyETG3pJCy1MKM1q
t5quKuoa0WKmXwPtSHKyv9w95BEp9nGugQxgJcU6b1+HXXaEWZ7WELG+QnJ0
BAehlpGAfo/VWGX8QdNLBCiLgDTqFvFQ1AX/cljfSCuok0wD+yuUDO6ysgqV
fy/YOodGY9BX4Z4UFpXJmtpIHi6xI3TYew+3Q7CIQMmxgaKtJbl8TTdtNmLk
5ovAm6Z8U+OuIIktdacl51awGveCQ7syOx189dyGJBktaEXzJOu9HLDbtz9o
ReHQB/H/jsMjfBVn25tU74UMOwC+EU1aPkax9qkmxsXAjzovkujUBga/H5Ng
PTc/mGXrpl6cy8mM9v5Lw7VX4c/b7dLoOxgbPa/7+L7NfqmFWQPCj1bmqogN
ZuRhWhv72VRP9SI0o6Ha8hRjDogl2z+RrRk4pr3IkRAy1KzvGRlodXdN7I1f
qkRmvnaLyNkc1TIuti4nnPM87GoH9VwfRvb7+L3ZMLi8iMEix/BKfzmaVK/E
KCliQF/h8p8jtw4FEzfubjYOnNnyNkhQ7cLEUIRNHvXfl6wXHG0oHmjcpwIS
vNZtFRoR5PxdvtbqqIEAqajQVoW1Jbs5BRhUih4wwim4rA1YqTzcXbn55Mw5
jUgOPCifB8zR5+eMHhsXZuT966QlhHZ+dKHxRvaXbbAYi25M5EYeJ+l8HGCk
epBAKawn/Ya7AI6oBGEyrzwE0f1KkRotYrgMIuP+rJjbLvJXXpo1wruiJYGn
lxJs0vJT+YqKEL9/UcQQqyboW2fjcm8GmKFkSlxcnVfT6KMspkzyGoXYkX2C
gSD60hSn3Uf/e6/SiyyMSWW8rSNS45X+NHvl5fg+g9aZTsK8/laCspNK0GdS
bDWRKG+bszUPWL5qBter27dKv3TERR758rxUwZlCNU2YcahClCi6z1yb6STT
Qtj8ASKw55s2YiY8i3Sq3d2ZmKfp1ImhbvpLhWk7LQeibNJBPeETGILR7sqh
UXEtbsOETxMJxD7UOi2YyEXZaOtL6gH+uxphq5G+dvtLJlDsZTVMhR9jvlvX
LnpK5zYCuE3lBwTxBYRBZWxIoKQqq7R5KEYYPRnwP8+V2Tj1v7Xd0l2eX525
H+Oo9dTbE3/EqU4AMmWF38Nr20YUQUW2FwUgc6fqHkb3RNfbDrKAXa7n7hAV
vZdHlbCq0RcZHcKo9Y9HgG4bOt2LnN7NVVBD4Ufd0qmPtLIHjEZ/9ONTQU1w
EzznzoCE8EXqtklekL1tfhy34TFEcQkhyVpeXsgBqvMLu8IMRthc2AnO8qjK
/BV0noVj/kTthlRtvbKOlKiY92AWcCwGtBFpKBoCmOmBvI39fs2X8SkPLCkc
CfjFhQrO4Qp44QIbyBlon/efPi13r0TwiDvI6tzhFEn9HUFx9ynwO0d+oX8a
y9ecEzRRsA/qKu4v0bUsh/bbHd92bwZzzdi+Sb0PZgP+vjCV4mgljuhcipOh
ZzwoP6mzIcXGNhA35t4k3bbc97DYzw6wc/vReV+S//DixB7lH/1z6GXKt68s
CHW2InQSyjEISwuoKPgzIx3z8qwbO/+IlaadiIsce5XZa637FzKWhXlxRvZH
ZQfIBonKfTHiKBNqxQP8Q6iWA4IME5b0Y1uvTGYoF2oSUvyHZG9dBa45Vxvu
B3WDXxD192zS/VK+Cij122Ttv/HNf5Lk7GEm2vnEQjXQAw1C7taSQGew5OqZ
JoO6b8n9OtMnuvjFW0iZDtfK7yZ4ZXwyj4K+Iu8BhbVQmhifpIBLfqCTOUhc
fbX6IcKblk+l2QNQDNhsaA+rk+PCDhlrqsduoJ/0na/Us//9yue/P0B0n/nb
Ht7UtfeEQPujIbUhhv+2GBCxvBHAGjCuWnEmhNM1n2gPubQqkmeZttI5q93f
mQ5YDNkqwvkscGTd919yp5CMzdTfUEY45A18tJ1HXCbYpUIX7QevBgj/nWaM
LU+XbcZRFPKBQ3Vms9JIzLE+po91zxdjDmQC+yg8O981GRYPSz3INT+1XkPm
gZsvEQluKAPqZ7JuPTIwpzcPqoFbT/kYiKKaUeUWys2Pzb1MLoBFFCerei60
RILMaxEXEfFkKpUPB1mBPxiBnfC69RYvTHH1vlFHiX0SO/cAV/oe5F4wC6wY
uqGNEwRm2pe/3huEqCBjAvmHDpfYtRYIHEubpqxU4wLwEiv5sSvaUcnGFMw4
9ukpDRWfvZ23QgGAkDp52ZRHa4VTSmcALF3H+3VFAzPc6xPZuS8rYdInJzAn
FCBBP4/ZBB/0V/N6xeTSSY/BRGVZulbnID/l8rf/5d1Ziy1RW4SURDkERCDg
QjDGLm/lR/Jk7RtBE1yFyedYZn2KxkIFZJtYmnucKsKa6HAkG0weVFba9+BZ
ZwF+Ip2n5gKctNuDQ8FOtonO2HrizdS6wOks7kJQ/TQJhIemKjBuz4p8J/wp
KW5DRgKuWdXjyH8KHR7yNNjEwZFiVit7cMrMgxqOrlAa4UvEdAq5WXvwHNOF
0QkRLskEhEl1EGbljfjfSVumvT8QgJ1zjNY+HwIrv2zP2aDibQhS6NlGgmDe
9Ndyow96AUxW/0qRAGsov5WoKy5axvyN+50IFNUPVdb3R+kCAOZQFfN6MWa1
RfbJ+DJBAP2bADmaboqyYav0suMgQ09WSDoporsDBQFHABlGBZ135S+iFXKd
Qek5T8Lm8HFlwbNceU41W2bAk+FtPzHY42IiLYO+nJQnfvY3hPnI4gi8UGal
DB1h4uLFv4wpdn/dCCfvI6jvTBfgjbv63cLWb2JwGqeqnQzHlhw3WaCfd0Yu
T+dHVNTSKWMVDYbTsS8WnbNjoxRG9HOaWlEzKUQPMtfsd9rON1jJytuu70B2
g/Yxhebufs6Vb2v8jFYIZrLXGDbovZfyYGWv8V1pMhTlEvX4S4WmkWA+yhnq
372EbtR6xTnrPFOCDbzVfwcbDSO1SG/kgsSTEg4oisNY41Z5A36GyU94pfGa
Hsbtwk8NHxqfh2O+W4Qu9XYP/zRZi8eQ4QrRPy0LBpwj89WViEYKDUvrIaQu
bXeHx+m5elJp3tAMbl+gAtPodjEw/csdr2Q/fZsift5wBo9xnSmOd7ItRIZl
mKlpTz2dg0x3U0GLzrewa0YuPCqEmz/xe5m843ynJ537M/RLreGaXbxdH537
TS93qCRYMOksWApH+niXp0ammNmC2iekE0f9KUsvg0ASJ4oTe0E1RWOgxrK8
ztG7lS7twtY44jnohD3Vp7Ta2mlA/AoLfNgLOEh1QV4dL5SpZqFBGLgj1KHc
wTstFDV5AxhV7QLVO1+mWpdvuyolRzUK1qXNi3OECZjwqlepqJJLXxoU1yEY
Daq12Ezt9fYAT6B4BM1HwkceRe19RgnpCWzmA8PuBbIpHal+jhlybuPmcM0s
L/0V34XBVUJeyJBW6w6yE/i0rX6ZNu4yxkxpBHE6dviPSJCeqIhaDyVOQi3X
kW4BeA8yfpXeqacGsmChWWI1/EDgl8RZy/JMqjZyS6el/xXP5yVwPwDG5lmo
gSXByokNVHWDJCYUAJ0Lp981s5OqqXj/Ie5eAKcllo4AckE09deIVilu0f8U
KkxuXmYZcryAt2Jy98euokS5AVZ8oY/SNXmA0BUGb/2omOK9MplB5LRm1yYp
D/gO6keTWWo66+QCXxhi60PAnPIG199lK72rcWKH83QpQVKw5fzsS1lQ1xy9
SMHPfM81QJIpZxR//RGtZkW8iZnHCvuzEGIt1dgPuMAUjwVEBU7T1+T4I5aZ
SHC/4C+mT77D8snaKoGsQhPVQIKtsdo8YyBo/iRMvQfLDSBqaOEkC1WS8LHk
pVK8lEoDalzfULrc6R7mcQhnQ7VYAk8fGfSbHVZlZeImsljdXLMAndce72Xo
W1g9SqgNaGO2ebh2CZotSMeoh5wGYw4xjymUnecfBzbwaY5xkgKBMj5LdADv
S0Z7YR8uJEi6MMfKbvU1fqVEnhJXlelnRcbeQAYQ9BfS/20f2KioiP3y3H8c
dOwx38pEM1dVEdOaH8vqPCktYqlxt1POyRi5D87+jekT/z9yaTJ41c8GHSPa
sX5ZKm9d6oA784k4VWK2My+2Yt8wfQG6wf2qD3lZwx3xwv2g7kY7U0uQCX1d
KV34vkrUNz2aRSV9xaHBw23wkJGIKsElsejFohQz0a/kKDcVNelvM5N9Dlcc
0utx/NMGpgO0/Ja9Wx18J6KquU1Z8tbygL3iyPpWJ3mOLMJBOK5juRu/ZWGJ
sB5dqkWaW7VkoynbGLxm82yC7/N36dF3EQNgDUuDhU6BWD5Wd2SmWfp/DUMr
7o+SnP326vOCH61U5JyjlngKZyolFTi/nAka5hSfJ7l7Ek5NAxGM8lUwRiSY
ZWJkJ6Jh45FRmZdZRhC7/JGkY1hVyLipXIfW8366I0qIPRvSbgzKwDI4gPvh
S8/xNyG0b5MVKUricb/9+YSTpYEyz84wZX2ami78sxcsBa6+KLcwTMkjLUZ3
e5xReY9nHO9Wl8x9BC13tBXWY1kLjNceRRoxWbiTtmz1vNX8RVRhvDY3J7fx
BzRR9g4ZoEVBIeKNpKK4tJ3+Gb+CAPuOXqvGBVXE8GYwJ0yhhONLfZ45nDQG
c6Ye3lMNt0FDlVwbzVglr0uz+9r+MOBidqs6tJmqiK+tUfBBIerSuKJKJ81x
iAC7OqsbvoZLaXZExMM0bTbwem4km7zk/z4/Vemzrja0jM2JOPqcsr41ggYB
YDogiZ04E858K6kaVMnyfZZinn6eepeNlGLN+b/e2X5yIyjNNc7D19Q5ZhjZ
VeOjFOImm/7Glk6J7HIxFxQX3cHylqgtyIMIgdlPIeQiShcQKYZu1SxjpUtt
9Hnz85puWTVeuP1ka74A1qSgTHYcqVFQYnJb14irliFB5oZMD6+iGQLtjDIX
MpKG+vO5x/K7Az5f82wo5HOEHQfDlIAzUw7w/RVXyGmIu2O7PxfBPUi2MFC7
0m4/J7rmjC1OgJS0SvJOWAxDFKeHvyl0jFGImtKlnhklDBDOiRjAeoohNtHS
rEXkqEniQ2wo2sPPZZyTS1sbFRR9xMupzpOUUq0WyQH1Vj1lEYzQsMtMGLn6
w6xltKfMpIfyTrmEBaMO41WU2vR5HGXgRYnHHVZMv+hfYN5SHdaebygj4fl1
E1fN6dQwVYrv8i+ZZ4LPxmckRk3VIME2ycEETrwMn1zs2o/V2OO1bwbpd6bc
9LWnY6l0yyE8jD42ziqzQSyS/bveCAYmJkuTjLvsGfoLxXna0KbFwou3w72D
kufOSlBQbCMDAiyC20S5qTIc4dfYctSLAG+eZdaObuj9/dct6iZ8MoXbvOkK
Kp8XJZ3XZfWt2ljZINJjroadEkb3NbeXiCtZ5jHh85bM7Q3VXTKA6wG1vtRJ
BwZCqCmWL5bLJvt3gMA2h8s1f5JbZVV7qzwwpNPYDZxH7hDVRhEiao7vf7mD
+IFWqYb7djdUs1VReicHNTiJeOUYFVfDrS5zy8GZZNWJJxkQAcBFvm4HUxn7
e2ofn3nsyFVpvlLnD0trz3bA0+J56yaQyBHKU5hZEpH8T7MA5SbDp28MJI9t
utKltSRdZtZhVB0Avh7djbTLepC2lOsdzepYCj6X3g2uiBRobaunudoJdSt4
ZuClj08gusyWy7uqtLH016dBwS4pNO5v0zKj9OZv1F7Gby8T1sBLdm3IFgMp
7Y9Dp7s3Qgl3fuRY0a92LYm7RvMAzs+T3jDZpTQql3ZLe5hz4TveaJ4x3v2b
FhfJXHMXVCeGaSmvTo18JcnAi8A8QWDJQgyrG8KLVxRqmcQTfiTD/C13v5NG
kSaAOpbpPFX5MtuS9ukkyTtrkxApa1SoFwa7JBVm8drPJ5kidIHA7DOjcNql
9sIUPL/80+0m0tydJh2eWHXeUaEwSD4d8Dy93kcodJE7x8FaCWotLLozILi7
U2zEhzUaTtTdidHFbcAacBQWg0Am60KAWxMU5Q/veaKfTyEL0yNTdYpehbPm
YQaqoZ387g7YA9Arb/ou3eOi7LvDK4UKUENRG8lnF2HrsRjpiz6dxXUwwacf
7JG9P5awNRQhHm5PW679EftA79cJf4hq0QH+A2K1HVoPa4O210cznNEBdlDS
hFHt9YiTDY3qCMxLNG8Okm2WLiiPdkSw6I0c060/zefFAXFpudwwPnACrw8w
ZBPq+ja1FOQvuvW98pUsljY1nmHrglq3ACJgHq7z+lMtQEBEplXl8mJkHSf9
+TgPX4KOCDm2BsjH3F0f95KbzWDFub4rN6JNp3p+f+UJDHTrAC//LV8LSjtn
G6ZwSV8p8x0WRbJWI3fTis5X+hegEyLSUrAMCZSQyvaf3S51aXcZdSaRgJmb
zb3Y2PPho1XGTzhbDF2TtAIxUq9d1VkSGiJMUP6qCrpcMAUBIG0gNe5afujb
9v5jm+cDepKLBjuD9C7jPd9Guz4BHg0E0yj1In2/8momYMKjHD6u93QJWUHH
jHa7iVCget1ZsXstXU21e1+XZGPztMgTUVEwkxrlVcID8qbp6DsvLjTzLKy0
LkxIA9QKcIyBxgSifXJlHRe2HyUWz+azCRYQCX6u8XbVSQmFYNdUsXSmKoFD
r8CTSSb9YiNgDSAAgmtcaUYNJIcMgZvMdPnDBOew0FtvOuq+aMa/tB4IpSuE
Llh49SjHhqdTZrW1ZAiE+DYU32N2U86E9Ko8WPeF3uD7+rBmeOoIX7S20Ujf
XHwZKFdTJkOEWWGft1o2Lwcv+odiSVRlUcQTfeUv8YzkoM75W+QI4Dw+9aAj
hprQG8yzpVrp75mSoEEPuBWb1wa7eMLKiq6sRri4SL9kRIJqw4NSjypjzt/1
vRgA3yQ0U9AFiiMJI07dxiyx3N6sDjdo0QtlIHwoNVl1pb4b1tEJDVxJJZZd
N/DIVg3Ah9J6SmxzlxO25gLGX89QiG/VY2V0gkXWw2o833S/IyxP8zPUdr7Y
mm+8TTmbtXQapfZTDLKw9AIseuA5ED6+QG0rWhh6PDdGyhZETjBOD+BB87uV
bkEh0RYNoig0GQAGG4haHYdGPJIteA/OYHwiljyS+B0OnGzmpm/qfyorGLs0
ggYFrEt2St9wY0GN8ENS/ayDOXX+sOs4EwYrDGqBUytK6KfgGME+C8SkX5wc
Tqi1+XIzrnbAOvY/n7VuxN625CkPRTip2P7z9bjIOU2fncRbfA3Bgv0AdBjb
D51NKM+dmeyQOzkpDSRPnRmMJuiPOuJRu6BKzEjB8R15FbZKaU+sNpgYmz4l
5PwQ61wCOmi2mgN81d3MPGxXeKKjRQnGU1mBnhhsQU7++F3nQhpIahYFuzGa
UhNZhs51H+z0cZCqIJe5C1l0WQ0ey/7G1Wa9IuJXjKHeRmANRXTgvzFk7c3h
hR1H20A1hMVTqRLELfkYsYm3ecMRbKW/CMF/Cy6OxXgt7LlBtew2LVf21sJn
Z1hNweO31VwkITdElUX6msYVYS7wFKIsxtUy+fvi2NNLmvvqHQGk9SkeM2xw
YvKIhni50flyVdFTuZjBay7K1FvzzOhyKn7jP/ESMFd5uZ+TCeLqTPJgmP+T
f6IkpkC/fV36ZqNeMlVggI0SHnCP1DEyAnFE/q+08N2TaLSaleqz0zcg0llQ
PAhrgVCBgiTvrAsxXwNQ20jQBK1AMZnasa8iZF2leMyEkhthHavilCN3pQAj
+No6NgXl8pqivOH8LOLZz+K0T96pWbemSsMQRNKKa2yj0/KPUMWM9N7s5Bmi
qNA+8ePARqM41rqn/Dg9swvMdQfUDhRxBIv0Dk0Wj/XSXXGZeJuQj35oeLer
1SGzPeJ4BPS20ujauO1I6R7FkvYaH7jg2APKwhtQ/7fh3jTjFyuUZNy4nlBD
Ck/Pi/syA/z90ADDUIgQ0jgXB/9K5B1QHI0Upccb/+BI24jRrwkyJcwdfTkx
792d07WWBQl/BLCeFUC0jfm2LmwZd6LX35vUYaA+eE7HLDHXXGEo5CPl0aFl
dNpYRdAbH3VynSjDqje3XOdpR5zoINv8ax9PuoZiC4r9kxGMd1QoWKoJxooq
Vu7oJfwexB5QQIjvrkGV0RSpwcMmEJefvI43dProyoJBhwQvKTKTLJbeyi1p
G2emKKyxkhhbwWcWuZo/9Hx6qK17E1I+vKXCukOYQoBjbl7CEL1f36qL1oCy
DIszuxLkCsgTIl38FzdFTJv4EIHEMeD3I+OlmVSzHrEbI86lUY4jeGXuBNWq
T6tYp5irMs/V36JgYQSt1UIvPzfY+yCBGj746Lfpbd/E/hIhEh1MZSHq68jb
RDVzI2eHm+N07pZ7rvvcs8bftNl5jHw/LMNQKb+kCMK8vuKXWeQv8ctajfgl
NeZZSaW9J2KUubjADCMhNm+Mi8Uq6XjCr5fkzQXw+3JjMYwVAyQXOfv7lnd7
siZX7JxmMGVhJ1cYo1pLbzg70hQnwgTqyYk2E8V6LPaOOcbZ1UJU1SCUU5oR
eBSP7DSLpN2IXVjAjrOjW7ng0Z27QAoqx1h5sdQ2pR3WfO1sb6jCtfEvaFfY
7HzXxtd+vW+xX7CXoa+/LRrkexMN05FznAkZ2QsVQFDNADsMdWRBAtU86d2s
/M0/BvSjwg5sMmt1i3PeUR0fpdgEhKn+QFi2lp5nvGsXUA1Oqw1aLdSjvVfW
lOiIZYYB0ylo3hpeYgeLoYsl4NSD8LnsUwr+RaIH9ZZNskS0/XVPGH4VNmWR
3pddhza4vRSI+0yPZKVqhCozl39eid9L3FTuTyNBMv7xpDHmhK/x/e21tWoU
X40yTHTgDPxubh5wZmVoXlDRRa9H3rr7ckiensqnp3ycyCAZADJ8fXzYB1yz
sA+/3Beq1aEZCxEN4rb2gAeatkWhLDHQjUXvnUbH1Wpt9sSN7klNW/p0t1jx
el3ubQ73lkUShUdRyDwrBj0NJ6IFJuqBqPXJdLHjUA+PDnhE/HLNVzZWSlJT
bqqtEPcAXGv9xWXDX/qDQnEImQYRT3Pf6QScuwI97xG5QbuGcogtBDHM/qYY
3z7hDiDe3jaKRSVIcYA7azP9vV9DmAtozn4dw8LoCR+nXnRuOSIWoOLMbC6S
Jd6Eb5zoBaUuv6LS61mLsRgNrIaAC4hX9ICb9TXWzeaTvjrLtkIDS+Xh7LzZ
swu4H24fFxhbI0rTTArnkm/KUQvrDqTRft8NmApzRmiTl/+2mHDY/8fDA0kX
Q0EjpLgq9Ujbn6f8ZkmEuufvz141MRqk50AcZJuJ600617nhwPijst6CLptQ
oN2biP6IPYMCaKE9oAJ1fTDWBpnImU4KCAD/rJuD7iYEdjmSQxeUU+RK2nIP
NjUOBRWI6RPJkdiua8N+AHKXE/AGteMTLYeN4LGpCqoHAYElYnRYaRfb9Dpc
eOVnpdqhl2mQ1PXNFAhGX9kcs84iFq1tzM+PypvxOSSv76m7zpLS9cP2LGBP
qUViXYIHZtDVFg/4y1Yx30F2nL+NJRCcvVskxYswVOUCQsF7Bs6wHZdETAZR
tPCxDYOLNyCaXaS6MFc/oG0Emrw4B6c1Qbl3jht24lRNXpdzYjzSTpXho5zA
OaNPxuZ+sWOW4tf1tuoDPbgn4EAiyQin+G97QVF7fiO5Vt9/HHjhDce+5Yx1
D2h4+KdHRa8Fa6XzkSuBope1UZWDJOX6I3cm0CAvbosLY2gT4YOOw3NNZeIC
w83jPVxue5YtXpQgXaH+astTXMcTgtGRF3uI4KKh6zia+n2UuVZQEpnib1yk
EBrx3m6VOTa/dJN5b5IWcg3vm5xkLHGrb6xDRjKg612y3DuRzmsAqqo5HVlo
AhKROLT0gei+gEaFStx2PPUx0cyBo4RvzuQ3UxAAnTAK8HB3T9F0vqFR2v60
wiBkvYa0BJp5aimb/thqSgm0ILXfjo3zBZ9HePJd3dU9rnXlRSrjiLWtFrST
K/i5iY/cUNuBvG/T73G+FlC5ZtG45trGlNrz0OtIz8kMq4ueUpZCfu47gN23
buBEPtEQ5sqFDTvvvzXLMJKFYggnPvSKlGLtf0G7/fVQnxZWrkB9ppMbeTmu
7/dGdPlgPWvs1SugVYR1+g+xXOJ3OAKzbt75yCB4MqU8rf2+K76DvgJBIaLw
lK87yjRGDs5rfwlF6EmS9h6tUy64QmAxCgl9V9yUZNwPdS5J58EcVswU/WZb
sP4JakzD7n8NSwC/kGCE+jcQkpZX39Zaeuk5Q3CImEW8J0PRbfr77otIC02k
nMH1j+YwgfqGgop4cRYb4Tk4/otS+IF8CnU+UOazin1HjAn3MPGsNNqgoG1E
2KXIscRHBzEHMP+KFSxbg1HBQ44q3GAsSdeBF5MKqUflUIFzkJXWPu4K9OV3
9F/Az13yXpFVzeIEu+T+i+LpPGCxWx/fgS4JkIYvGhG3biTHizdQ4Z8ovl5c
No+Z5OM1t2+7Va8EIGCQOYyUn6s6Rdqo7vJtv+Tdgo8xSN+YrOAD0VDQroeh
hf+4R9Tv9GNhrHu6lgfZOt4apORj0fv2MUMviMMD3MskO+HfrmsPkAcQZexw
nxBVDMyi7sF5ci2qD8DCqfOYBTdafUcgTamL3biJcO3ZvKUQAFQmFT6p2GD0
RWitVPuwfa9HfSCOwORYPqN6VFVGfopBekvV6si1X80fpLGEObgxZAaaz4oP
98YbHtW5ISwfhRqekFvw9cscxT3arINb13e97IwKIHwghSvl6gwsbEAFnAhV
HtxwQ2KP8hwTBpDcm6epa7dLmX0VdFh0wF3Q6leXj9ShMu1TvtAcs5Dlk4Ac
4tN38+h/YJt2jIxZkHXfmW8iqaH6Msh83vDq7li1kJPQUWSarkzkzrJmFdjY
bkV30gDqMGM6h0a4W3U0dX9Y8YVKH2ZU5ie5nvyCKbW+I4SF3LZi9w0ooDzv
PHMG1t6T+QxOWYMcuXnxM2GgwoyQAv/SbLHR+2toTem+BedyT1ays80A3uuo
a+ihdIp/AUy7B0EIvJSk2YrPkup1t4eicaYkS4L+f9tDWu9JuRbu4g8+DFyH
moJCFCzNFrT0buED18O784y3EKEwjVaUY7DIa3zQCX9O3NlE3qFTOUImCOsM
kgFWe6KsZ5veaJmxxEUzdFsJdV2AB0x2/Jg5JmsLJ4EhdheWllvFuqIevwoi
e/KHstpXRuKN8SP/Bxxy0kMTttbEzu7mhkNzQgvylDB/K23RxC0tA5EEhni9
5SbqANmi7boZSQJYsGhQL2uUr0ba9i3j4AgNoyfHShZ/6mGDAn5qcewn3R9f
k010hVGOSyny9asF/z5dsam02RCU7rCRzrW6hcBaLEdcPjgRDjL1gnch1SmF
U0lhtRmui4RvdGE1LQP9tztsBZltD9qh0szSd51MfJ7prBY+stPATQfMoTqj
T1/WHQOk4/RMobpoTQNDZPdl3UVwrUjirlW2N2wsLHs5zq/BzmMmgbr6gsTd
diYIJJTpERAKI43NLwSYEPMLWs2R2/WzcUkDyALlIHhW0IAlQaN409a3fgym
BxC+h/8ka8aZ9BnGldogbxNm2qjKzhTbUedSVVFMsmq+nCKOwLGEdUrnTPyL
NjLh/FkcRy25Cn/r7qfRgBcQnT/S/rnXJNoPeOTw84B2/LPC0LjURgZ1dg+G
FXOTb4FrWKjhU+eXvki3LQVu6LZBwkw122LiUvg9q1FhlCrm6joYxx/K4esO
NRnY//u1D3AEkFbCfk9RhbaogFyQ98r+dqZmAuG0OkT0tXTiRGy9mkk31LkZ
sgJSgHnV3E62ho8BsisCiHBEot+xV2d+MV1hE05HMnuIardmGsnQKFrAhpfP
eKvwPa5xZxh8tD7q4YEAacwmRocoo2YDiO+rFZKAEvxytFoA4rdBttgMY+Vl
YOP5LuXj/0nwrWjfN7DRoA3hllLlSx1IIoDdJ+lc6NteHwQhiJCmjUFfFOk+
k3tJusEfk7v4ei0w8iVvNdVgCjCQQtIsHv9KGW2UHAvNdwuJBfsZY+x6DUgS
AqpSOx3d8lr58TpWBLLyWEYcB1kr0HsbSzLeAuRHwzX0fxpPTdGMGucL80Ib
oSoNBN9TgVNhAlL5rgngXTYlrR4jFJ37j1haasYIXuV20ESu4Xh84GBGx99K
LEW6bj6MX+3P6dQ1PoxfCT8VW3zrxFQIi0fGimse0uRz2lKaYB1nb9xsWY9b
Y8tuRSOeorpEc0FcGE2O1rhDIosZxCKOIOIrnnpMVw1netlg5vgBJopfBcOo
/9U+5SG1bltti4fcaBw8mTpXRobptRstRi/8QARBjQRSchyIlhj4Z9d5wgq7
Tfho230PHQaJXKRQ1BQXTUjPyp3UMKvMesYOozaAOK+cZGbBOsemN6YNeIWj
KsDu/PutbZKGHXAuQ9czVhwI9pjvsjscwgOyz07bTvgPT9P17/SKOWD/cnTz
GTXIfNFpO/6UIn2rYaTptH5FhbtdTBZNfEYOnsr269pWwPRIDjv/7FnoYOf6
7CyZWl5O/arYtlPuCRYo9f3O10MM6MII6SSCDV+sBp2L3zVyJVb0dZLvR/8q
kn6QvaSaYQUDjglkEAhi0jI0hXWe2VUHKd04FX1/DM5DSqw9zbxWuKATBa7w
eE6mG6/ism8EECPaYN2bBdAUked95pWOUpUIUC1HqdfPlV8XHAyJFJnnqWye
WbMOYtDJYv54n28AforYj1JfW8i9sTUYOSi7I1HkV364mZCS1Q07ON0JK1bh
oNcBC2Dv+IeaTfUyerPCybOunxBJca2uLkMUWI93gILc6rTo4PXT4ZiO1Jyq
kGa43Se5TmQnqGFiW0rSrDp8556iVUpxe2Ug5zzzVspxDmYMWSBL5lRUUz1y
uqwfQM+wOqJQT+U8h7GkhPfRoTurOSKpKKvKtHazZhTOe1mw0eS03am/t4ee
HYmbyIh84wQ/CHLD/jTYoXUSoKNmE5h0PSWjrQRUtR8BIMNWHMP9dy2aASto
JMxxSJIl5POyhF4w1oVh17SxpJv9sxq90vpj0wDtlzS5H49nN0sgxY/DHBN3
YBHt70GX4bbpQv1CJn16zzEl+g+0oKeZpXYP3P26ajPEtce5xDYvldC8hTZJ
Ubpfjowohz8ARQupfKtAiH5+KUN6rUKsIz8UJ+mCMKto8upGPbO63lQ7wWoc
2oBsZRKywyCAjm3llezI8UJwEKXu0YP3JxAhXDt/QkRu0+l4esLVydhLcaZ6
TcLbLnSVT5Noabqmnd6GYHDOl37oqhkfW0a81Es+iCedvafxWeK+K0s0VRGz
AhSN43kP7HblnKB6Wi1isYtFUcwQenxVxYhvhnLYS2QSOllrEuda/G/QmwQb
jEAACx+8xvousJNbuG8ToRNMS7OWOq5HI6rNc0nHbhmd908QNwJ0yze1jTne
scU2EcUNfMHxCrEudHrib9Faw0X+tK70S/IdbTc3ljiikdzuStjA/cKheIDk
prqr7VwJ4EpMD4Bu5Xk1m3oc6Uucu30w4a8OJA/CHagNtdpqU8slVgDAWohp
Az+NQYuVBsgsXMg8PGwAMLDm9z9HNwwweYUs44Xi+7lsxqdT6LAUBaJbWmFV
KDSias/9hRHyxTg3YRBNDHcGteH4dyKCgEK3BG5/6BYlvMFS0bAkJ+eb4wKv
sX5EI+LdYhLADa6VmQcU+u8XHxSexH6E2Ik/J7kEQLDYpzfp4ylkNRRccWdh
3LmVEBFE5uriurNwonws/DLtjSJLPh7/HFEv8nIuGvFdFB84w6oYgS7YW5B9
UN496kDiKZR0aFWpHoQTSE4qJZtaHG/T/gkUeyw37JYtfsA3ipwGTJ7rMiBi
s14JMzkV66xHR9ypSgMOWhPkC96MKqgINUS2wb3/XZShmQ9k0htfT7b8+EmR
n/QrwMJ7caubE2FTDHd4vKftLYiiIFqZQ03xOzwo57lcZqvROwPKqGrkXMjw
ZVR5+06GO4VUlVrfQ6XQ6Ig2UiWwBAcvSVCwQUFDx51/TqQmoS7cmAEUIJog
RxnD1C1vyCc2s1K3Wd7k7qv2yR4x2yyZ6kGUplgSgwLCxJ0sLlJOfpXTCv7B
851CuMRS6UVgRaPiwauVpgO5aQ7lwbqbqizkP2TatPIt1rA7+jfpyYrYKVQe
WtynwJp4nPY/Ctv12SWfUqbjP2Pz4nAY6z2L8PXneVnPyINiVImzVLyVlo37
y9IG8xvY69NVk+wWWM3wmlC8wWCNGeumU+1Vd8UQcGEA+nJ8DYo5+IO2/gZ3
th3ga4IMKEvihT84qFrXtOuOWA+ghfZfOmG2NnQuezTvEGanBWlwkDalcana
J1o/oWjy5/H6elSpbDV+z/dMci1ux58n9+NLc2OLpwhqkKbHdg4QMiQcakXy
bYKpYSpI3fJy+KTKsWBAi2FhoAn2AQTdVpMty13kBRVuE0brHqtbxvjiY6rL
OXaLf69oK+TvtxNVkD7ZPwWWA6ezCQ9hS7JTULMCwW7g6a+e+crRbBViw3XT
7xPfgNUyMMgC8JzkO9XCHQCNoN0VTlspjZu9sFbHme2zgVYmnhsGGBhD3X13
+3kGO/B8Y14D6l3VzwFjJFi/VCpvIOSAYDC87AquTqSbTiEsWYlC+0l8DmMW
FDzuIUALaFuXCc1ZqY1eMbNCGV1keY8RdI4HIqbJIe5FxcvZc+RLkTsv6fSP
gWgwchT9nn+dWTPk9K7Q3aVVV+xiATlwo+z87KhZjp29pHjKKT6MgY4qwQN2
25jsf36h7O80YrP/Mc4LL5cgIAqVdYpoEnc1iSNObs3PU0Cl2kLYKTq/PtCi
5OxEzQoJi2Ae1ipHbCWboZm/w+0TiRobdAkbCoFTLlaNCaqp5/vFZy8cALd1
BEW50vFdqrnAVbzZxK9WnPmeVOnbjqlZmKjr+JO5vDmHo4Ywm6iHn9p0nMDi
J09hLnlb0QcmBBeYfkBRi6GsfFPpdGrs8OJpf4mC2jHonihBExGk4XwbKeKU
o2Lk1CC19jzsQsBLFhfjKSVr9uxSk/K+BlivJb5s1TEqn4lZKF4M5BT8p3Ni
KOgtm0W0QQO9QxM46gub7KyZWqIAzzRBvk+T1YTlyu/nE5s6fo2ImvpPojNO
qn5pKaluRRcjzl+7fqURHIBYn5csn9T5CtfXkDrxIWuIa6JUODCr1ILCcnkv
zfS9rOnaDPcjOCa4l0DtQTeaXsFhQ23LWsPHZAXoHVi3ZB138Pliimlgmljv
N41/N+k2j5C7+ZKSgX9Wpim3z2o03DI1Tyutiy9VfbIBgXd06IfmFOl4aYFS
PtrSQjAdQYCJ214NSfnV7sr/aBvahPkeBWKu6C3gKZucKOTw+AYSzYA8mJ2d
JE58GFdOwnFjQmcionXlEwuDr7UeUpc/EuaxZm4YZ0WXuq6+cGA60WEcEg9s
c85Arose0GRffTrUchLHp15rLVTyn17gifqlFCKgPR9Hnce9Hte9pGsZ5d6I
ssKdoWRYe3Du10MzmyzIVaafZ/+QGl8KY+snVj4yEII8wvytCCOXpjZ5QpOf
C0YQXRZt45cusk0ucxOoaPNeZuwAqo59zq2ItT2ZEGb+QRv3r6bIF8ApdWoZ
zUpAddzhKPOQmJlEWHHnjZmx4lSShBlJtfxqqH1gjZqm+Y4GylFlA4yIjYH+
uIZLrlWCwWSESnuj6BT47HgQTak2LG2p9r2K7ZjZ/xZa0omMkCQeNBfhZRp4
Ik1LIFqMjvQB3474PQLG5Ybl2kbFehYFP7Vr9nw1kI64RH8bsa4caC/099Jv
GBeeIW2FMeCM/cWB8bssfMunb8ADpfVK6tGuny2QaEkNbbrPTFZUTjnlveVD
OAaV8+1TLyWvTbG8bhZuHTsNQch3eN7QaIoPHRioV/pYgMt+IcCqB/LOGtK/
de7MRJ+14OPABmcYovRIXUcKI+usz/TLHPX8SZQc7k6Osr85qeWRITzSxbrh
t745VQBoHtGkf1/lTz2/Y2gI/2dIvm/d9XBQnx2O77MDGKikXVnzgD8s4HlP
iBVONXcGH/QcWFRXHd4toL8DjN81lGDgSY/woVBfUy2lEN2z17eXW272SyhB
qNEstHBZmOlZJQQK01gWBS6tiGfSZzeZaRwax8GN88RLSkJbEFSyNaIirG5t
XnGRT6mD0wFyMP600eKQtjyuBY+vOVxCT1rQ6PiNpKuIXTMHunaTeqFDJ25Z
dUAvTbG0KzZjVvsjKCtgyZ0XQELwV7kDuA3Q4ZQcrriadGEJuN5b2GGwNYCi
9qwUard0mzLnp7NeGsa3YCXAMz5BRk+5L0nZgVe8l27bcidzjE1bH/IJa1pe
qBpt7Rk0humpij5VCGuYsteG7DOA6nseFRGA93YEN9ziEqqg3Fzf/VfHIpxP
IKwbNYESsRNDh8HOhj8unUIVlxxyNK8Dc/9CcnSHq9qG1CBr30q0qCWHT+/y
rAgZylerCgJKEIFAN26s0TdpO18jm8LYK1COYaIHTZ4MS4y/rpFxi+FmzNsD
fGCs9qDEi6niA742I4oWfvSf5stePhhDSu1k1a5AV1ko1gus67EHw23CEgl2
ZAqfflsed62nMt1/z3yAJv5hnQ+VslqZrBrn2Xd0A3lA7og+B3KpRnkdL78G
OS6/J4MVGAxhjidpG6f+bKZnHjcosSpPW6ifWC3/nYgvOEW8aorvTbvyw2fr
H7vwWzUObwAkpXIFvhgSyaRkDbg1oO2IHAcRdYKNZMGQVumuV2vYnAkEchNE
3DeZRo3T6a8RsGatEqKv3ypwhJk9c3gEL//n9X77SeHrGLSOuP3W360hEzmg
wVhW4Uey5bVYHzwTC1ZK2RoWJU8CQvhxoxt8O/ktWqpFeJteDbpWz3TFic8P
fTghyvkpod03XmAQ0b6cAw8Cv3Xj31WNryOGHSPKyofKXVq9nAfUMb3IptID
VhrhpQe0oUZKIJfQf4syH68ldgqydLy0Nn7BiQWJoebrMNb3JgJhJAQCVQVa
IDY2RKvV5NK9ct5/uQKWx9cwAdr8BRT37Oxh0F8IzikEJxt6g4lj8kDHCBEn
aGwYJqC09Y/lbuvWPMMBGrPRGlSbTv+yxWLr8FkeijRPTi7qsCMNa6yh1Ni7
ea5FimOf95FcB9DhG8hzA0tCtWopjlEo4ypMvMGh2SHB3sQZo1HxTQ3CbfRf
V6uHP1HTG6fsK3tmLuE0JXNAZElc8JWDeDu6RVciRitNeYsGAN95hRRDWCvr
h+KPmJkCuPjVLz2ti13Oj/ac9C5f82bJfWJpbzpaAyLPvI7LE0nvwsHO/rGu
61VYu8AvbLLuC3dHuJ3s5s+YjGTV5K9uZIaVIaL38FB9i9B9TeijW1AyFG0+
5ec5utj0x9pQVVcIQerWtzqynittUehRnM1IboV/lwnr9K77AcfeNupm0FU2
tRsT+nXJVLP6ZPMhXw20Xu/90DfBIElJ2QurGbBSndO+uDKjEvqXFn0JawZW
H2x1DJwzbuihpYysbupLhVrT/hSDBFs3YL1pTG/a/nlcisiC7ffXSFd7rUx6
wHiCbGzPlAvUf/FsKGNsRvrNVyASap6wfBSE7cNZ6WesHArLhWfh1pL1FZU9
AMdS9+3XBbjvpJweo8oyllEES0bKsRM2BZQc9uZvR+/L2a1vdTVEfnZgktFz
o70qRDR0hjaTu3acrfEM7+2Dh8ke2Dl1SLIFAOSJZikHQrR67poSE90nT7A8
+2cMYKO82RpbaFqw7k4UG1kKQe9whFEqM/lVamjKG6NbNIbtesk3zMba0fXY
DlQTju/8YEtVh7bvZmBld2TtYzS2XxoZ+tizO6OH7W6k+BOvQcbLAKjpRGLS
wo7nlEWqdp5ymcNuUnMgByU6vN0vghfqXnWXonw77JTE5Iv16AqVhMnaL3x+
P1e3cOJExMGgCth19LnXXEYNnLdCkTEE5OK8VVcM0s8PUcX1p0Ng6VFVhTpB
bCFoKo6vZ3LJjcbu4J6qoGBLVi7pu7qRDxnsABJYN/DfwNAgzfgIG7hsKHCj
8h77LjwY2Yr7j6cS+wcuWXEuPUFYyfHponAnR4ZPNH2rDDUzbCEsTWX3lCrd
xManOsup7uVI3qUtIMwz3cVqFglDi/oVH42RE1rw0I1CgSLPkOTAdOTQlt/N
ugWO79dmcPaNq+0E+MNzwLNztHeCq5U8XD/AX3rGMVeEssAQc/p+ZkWDwkzP
x2ypQJ6JDsNptpBQavtI4/SgM2HsVQ3GjtT9zxgoxLnU3I0jdlwOdOFTQV84
jhaBAd3vpGcI5sP4O5n9JjuqLpRbtlYdicoTOozXzlD9DqTnuWK/0LqFU8U2
gCWQ8vpj85fvJafUhG1NoiwZkF88pC+6s3YyrVcGpLtMsmfxmrAsBhqr0XW5
5sJJ3x7ilZmC1+l6U7q1aB8LkQNcG6CUx7EyZq7Fd7jSbdbkR4G2AbMZHMOO
9LmDrC12NRzAnsOmDTw973AFBAwtUK2V1ZJN45xRzF/xqlEWA4Z1YwXGSyuU
k3nN51t8WPmmZUdIE6IgRyE2eOA2qJjSr7tErp6CLJLrstEaFftfrxzauzL9
BcW1UYvRTFVwIk8/V8OX9X984DqI/JQKzYtUD9siQt0hU7fDczl9iiBWej0I
sLWAhAZsSlftCMdkOHPJEW0xg+iLOAFXfx6UBQYkg8J7GSz3YQnFEx4shBGK
oPr6Gs0rvuTjrlSjRkg5NfTZcyr1UcMFerOBs4eqrc8W8W+3o/NGkK2dbqsb
TsgBuYvM7lE5cX2X/di2WSL+lV0+DXifn+to57UmKLRfCHxTluuf15wNp66Z
2XPl+1VM3peFLz6fj2SLIhv70uZS2rH8CJYiqD+QNoz6tZqZbBbd3/5IiEQo
8LUpLUjlF3grL1dRH8CIcWPOpv15rxTkqq/cTFLRF1eWqeVVAqo56muiSjZb
j6o4tkrY8LI4k5sa4istcHQL37T3EM9XlRzzMiwQLZ/OHjpNbPwR0bvsRiGD
A/PirXQqbglwLJgVAZrfJZ2d6BCIQurXPu5bbclJwiq2Il1USM8xSvsqCetk
fxC312luhvTGZNoKKc9dG261ziCZkHDDrhNDT3CtYVaFAHtziQyAIgH4sICw
LFrWpo39IUp+VHg2iqFEmXRvVAyKs9OOmYr+P8b7sY3TtTo5+hH/VFKXFoXM
Y3JB2DWW0miH/myImRl0yAOYZNNrZr2ubJipr8QceZTc6bAM/LawvRjOzEEQ
epOCISkNBL0QbJrGRSsDCEryEAdA3aEvBVDTcxRXKF+wTuuMUhMqp11gzqh8
2OARMX7IqAaaU08zykB200tVRPpxxKqUwqLV20mMkF+b7cc15dR89jqVdtDK
IBRRYDybRZPP8JZlAEcGr28XGvYGnOP7gzofYXlIdW6HxJXY03ZiQYI5AU6r
mn4ICd46Wo2zdVy1nXBuh58d1Zj+vUlQsqSJ63Yb+jbOB5AVWAF7Y4rhnmFP
/3mgDuvuHJlb5rxoSkhR5E/6tHA30ZFZUnj6bZzGdnasMp0ka2Y1VxrbDBnh
vqqkOO7h/YLzTbYbeYp0tRJDl9GoF40I1ROc6D94UTBKpP0QnAYG1lXArg+h
nPN11sUO8av90rDcK8nCFt5hiJX9MJoeHkmxo6q7cTZniMQfETsdOTsti/Fh
gcKIT0Dzlw6QjX8qR+DOGLmtGHWqifkColjoOCS/pWVrWaMlO4OkCKTcrfF6
vgdC9rF7+x3wATQajqkCSQVl6rbxF57HDbekCvx1ywvXj9v1rsvwvf2Zr7Ed
T0WARR6GpqX/PxWkzJWDYIlRsVqzDsSWfIGyVnTc3kMxYPTZ6nN5aQyOfOfm
qFXkHxKV7Q/QVB0juxsKs8HHhDm50BnvaYHf+fk8Evlyl00k/ubP+9kkym0O
peEa/YcRW20eJjX53knDWP2OS45i4ftVc54X0q0I+stL6GEpSGtOHsoqxYRH
TFsU15zxdVW3IqIqrxdoQsPvk9qUZkfvPwxyz9f5Y17PguI9YK6jaZdL+maj
HAKa3AfDwuvLqwkesX1YOb09ZL0Nk6U1Yj6T9mCQh8iWbAwNR9XB5m5I8Q15
7RAq7MRherAyJoFp5tRr9dJln7R9a+JCWZ2XXgPD98GQ7lOzbjXXjAhxh+ct
7AJD/BOo5UiC++hqjpAaUQe6p4LxYtqJx9TSFmsmb0GWpqjxG/o0O0uuGg/t
vwYd+fqWYT2wS82Rf6gZoS1TBehxEZejKBu/GMCDduKCiLXwpueCoFGawNhs
5Sb+xf8e9YZf6SivnPF8gir30eYnNea34nskM9EAe3rFXfZGX6dixWSacz7t
FceCGuhoQZ6YPI8Xz6t/IGnKS/FwcuTEeIuEP/bDRsENPUYyoDuawCPURMXo
AIMwBhdhgZ97iuwCDc5uzC/7tJx5iCuYsvp3wyfx1koKpw3aff7RgJA39nnC
zosjK3wQ+PtA8Lvz+ApJarjvwGtopL/NYwJ3Khv2TTbM7+phCM4Bhqpoj/71
nqK/+qqN+FyfJSNgj4jBxJiV0FKaCJe5EcUtcYct42hXHZxx5/XjFu0vE1NK
K/+kW9NStW/K9wVzLJtiG69ss8L6U9N5cAVQkG3+i3P121v7UevcCTAUqbJi
tKtBaECub73W8Tmew7tkhw5VPOvguGu3jCb4MJ+7vGrnYs/VufGm8nZdM+rl
BEE03SyIkaQ3K9u/vhIdf/2YQWAti0RN92fbjDwjHdWR6SwpSt8zdBt8VGsB
3ShyiByBP0hGzz/vjK7Q9nI7ms0Gb8Eab2/SK7MmtfGEyx2sjLAPmGPVRTzW
pTo4Zp+HcC34WkOeqnBMhTxwMI2TJvtaH7+wQ7mj+jh4+/BFW+rx4Rz4QCjj
ccQuWHwDy/1t4KA4yOP9m6/3OwzUJ5XsT9oszcuPenByUI/n6zlPPSlJJTKU
VQe53rLsOvkhrtGIThMr08xHQGKIiqkch5VVEP7I3BPel4Im5f+YZ2wxVkx8
zq/fnNAk3A2T8t9rsV7b4Cs2t5+Ikn4cE7cjrCwwrNnWaNR8OkxwggUYMAV2
5eUFrUYE1haH1D4NaOj0aTOEKRSbXZ8+zUpN4boQkZGpZkcSGRo9JQOUFXLF
mV8Qk35OyWckl57lGTdInmZMo1vFOwNz0+UPcD34wo5KF7Ti+9RvU47BIfzg
3Ts8qsdtnPXDWvv/XBeRBQhvLtSbKpEGimA4QjxERk9DdNkQ71HC9o2BekVz
oZb146sJnlokz/kJqHmgVPNB2x1TSeV7+4eEcUXJOGuWzpqm+Rw3b4RlXGG+
pR9Q6SaM5Su1U9+02xJ8XN34C/SNKCGuImWX7Iu1cY7V77aEK41GX3aIQaSX
atiQIMgLjn2MQKM3BZiY57Hhl706rFjjvy2dSl0zNXNLmVWCi9+aUsnVqXAc
94V7P37X+2blguczs9OL0iU24uH2yRG5tX8FyXsIpNoHoWrK5cGiyKkUzb+D
2BCLPGlxJQf+R5L3m+9KanrXq82mVyrRbbUIVh3mhwNY8+q7Lnt7n6miXBoW
sKB5aEGrTBJFvgUzDJ266oqGTZ519WV0r5N77tFA7aVmS/mSMTyGAdRj0dLj
2MbNFhXscx5suXMg/qgP9OeB4qYfL1BkPbr9rAphUTiF1ixB3KajA+PgoE9x
bv1x9snjucWGpf8uBJ6eQ0KDUCnRotnQeML+GM+GZPkg0HWl3n2W+tCCMfWQ
T7vnV2YsKbKXECXdrp8K0QM3TnYVQjN1RHBnZYahjomfjWyvxUkf7PfU3vjT
rON++d5SWFq+h9kxyKc/PN6bl6uCUr6WtXan5/DkvV85QIame+26YqkyQu+m
Aiwouc64H8gdBtcjudnAH+4fXsNQgLm9l24yTgfCbdm+rdNfVLgLu2Pum1gk
PcEBFtyXBq7y0lMsrnELdObzDR3Jrqk5DXyTvqsoC9r0eKcvQg/WkNb5j5SE
vg3sY2u0cupVsFLctyiTOLnf/qwT2Zm7magxxoWayZKi31uyW8oti7EwY2qH
MXxv3FiX9/RIFyNKyEbWXcv+iLsVzdNt/rAhJNFzZ28KXt5i/6gkT++65vPu
6FGAE1gTA0BhOCryKxacrVsopqDhZwep0Vl2B9rJZoauZVir+IF2/3hkIJy+
AAecvr8lVb1zQ27BjR/S0d3C5jG9pM3nNfU5BjXkhVmCMloRDwTunN+zLKXP
9tHffkHsjT63j8cQt34Snb3+GiB683oXt5+bJF1jCqAHPkD2XQn3EkqotsnK
G37zTbVbU4EEnwcK9KWqzTRcAAv3jsvAHmS5KySzjfMAn6/ePTHHBSxJ4zZw
sQV5b8bYQb4mI9RXIvgNGhoZ7JFGxNsb2B4rPkNrQvWVIF0A+OrWKPoFV9LK
kXz7sTCds2poBYY/7mf1QZgEKCyHFf1n2FIe1aJFQm0PFM4p8wZLnHK1U/1A
YHGa+xITG3cCOljBJLwnKvils/MhpSF8hhkYfrfs+Jn1+7StSJq28FkP/SDl
LYVzCXTZtR3COzhbyIrFRtjtZXxP44ElmwnY7Jac1qJ68gSv0xkex7zyMZW5
nVvZCXXniSXIg48kkxUGLe/EB4aI9iqyI34Nz+j49J3LXqetQD983uCT4rXk
hM8mQrauRmFbHNKQbRzyynbf75iqwNuqjGFykyKhRj5ioObhdcXBHB6gu+o6
mL1KtPP7u89G0M/+1EenF1c8eB2OBveoKlTUlFSdNzI97qAMAMWOsbKUjGHi
du4Ts+95dX78k4FUqyBWgl1tlwuIl4nFl8twVxFztPSCT3ZGOhG0aP1j81Iw
RDF6elfOv90q4zqyGkeHFF+IoanOf0sNs8YdPHeNxKNMtOXia5oph3OO8muI
gJ2YT8gKfVfTWG5U0VzZz5YCUIK7AcqrUr5/6wsqEkjH6KwHXli2Yh3Lw9Vw
aPVflOgv+HZETCX5VUVG+M5QqwA3J2hNH2XpoN6HnQEZzzdz+mzc4htvRM8c
aBGvjnupHc6fHSCHIzHWdROEYuiwm/BCxR5buVbGNsa2bnp6oXqMqJzeXjgQ
nRTQTXv/egTAKfaI0zeVVCS4fKbYaTsFHoGrv7e/7zi+5zaaVqTtMUo4u3fN
Pab0HyiwJhg47I4u+/mUw/C55V8sLcArkj4/1UiR9xX6sLtEUkbizj5LxLw1
B6kqgRseyJTFVwiWdX+rIqhW9kcYfq1e3YIM5UWHOvaTh2pBcxNDuSLTdrCJ
a/m9waXUsklxnfEUoHiEFuXG0SK6rvb9rSBBhlYQsiMlM+NLWjEy7oHrNmCX
uCdt/BvTzsnazgVPONL1Z8Yh33/XEUvIhjC9l82L+k4DUxnjMH3JO2un3qA6
P3mep1LsnbqqmPGJhopArbzraLDhI5FkIFkdSxSSwCsmVESjc4rSIoL3YAnC
6ltdmv7TGFIyyHC9t1fLeKwqAii0qzKd62gitIfrt7oX0W3beZK38vM7m9tE
iuR2IFOuzny3iBehf9+8JFmA++o2SEfJka9RN/v30Kp9cwcrbqe8PQAxknXo
L6xCYmnxjbicIlFhAmT6N8zVqs13tvpg+1qhr4mPRw/10Cy3xF31AiGud0VO
CLbWzTYcs3RnOKYLSgyBWmCaGDCd6MZk21HvJmjFo4AtNftVmu1xHMt4DKoj
MDTksTHsQjPxNgn14YILbnV9+1uIBOvIja0DrZR8sjSeFtRyxWSjzGGFJWWr
l2/zaQHilcBnRxznYY4AsxEtY4aEeBNRogasd7PsfBD/jaRwGkr0e1JKBbT2
BWNOSJuo1ximQxlJ1sro5JPngTgfI1QJrbeUPcjZLFxqzCdxxUhlXOkTkwPc
TEqT1hwBYM0M2WE8UQCJyJtszXlo39bgxL32wP7jFAEBThqQyMLKknWxwgDb
d2Yg0Lb0r/C+6KMaVGLCx7i2TWCVh8Sohelzcgir/m/k5R7IFKgKDTSINHDg
9+1nlee5wcHfzCez2DXZpQRMNCFt+mn+FbhrZtjfx4QGWJekeB58mR9ZOKDb
5LbBxIBEzgo8qLa9W+p//o9172bL9AEBbRqRCHTA/hXfm/rm611+0UWO2RKA
gqudtYSf6hhxUqoGzlFA/xWq6bTUzg8/a+NzHB5w/wgPSh5u06r1V3D9iGMO
MDZt2KLnsMqyC80Eo7Tmp016P2uCFtkNk/ODLgH6Ii08L8/tQlC1BT2QgAs7
/Zui/atYuj+mmCzwSaLh0B+L6+3dZuvWu+4E3xmKxPp8OzZmQHD4WV4AopDC
55OsTlGF/QsfmSirHYK3zDCjRmDh08hbh1k/rRHy4iHOthugZCDZpaSznKD1
RIppGTHyYFajtewT/PUUHTIPLstynbHlWDAxblJsWVQ9gLzUT7Zc6wNIvqAi
tCgmXN7xbqTpxfdHyauPIZuhzJbMpSq3QRTP9qcIx2oCeLOhmFOBIOV1dmgi
FlVZMMXgOtaR6emn21RwkKy5vzTHE4VBoSetYuoMrhK+xw4nQEmXJ9HSXoGR
q9AYaOuW0fQhfgO8FfHDQnbnz6M8OJ4x5p+WS1HBEFvEYd1pFb2ftQwRABNE
E+62beAWKORX63m+kbpY1oZhPe2/hKBMU96Ix5MhCe5Tr5z5eyKklyMFrIwQ
1nGxRhOmSQQ56apByJZ6mJpT3wXdoCv8HSYjhpQKco6i2SdLULCpKaruwFor
f9K+SjUWRkawvcVuhii7TA4lf/pnlQkTYOH1FlfNhkTUSHBajC5wl1kWwllU
MyGnxGveF2ZZkAc28rPlc+c0tuy8OUyNELiBYV7WERVfgzL+UAkyfUtTW/Ip
Ulz27K2D5f7YavSl/sdrrQRwV10pih9bgih29e3Vrd2nJ4FZS6b3+V4H/zyc
35xVRUafNOMUlG8XrBY0Yo57PD6N6xcYy6eqzAorCbVGAuGad135k6wboUmG
tppwom7WHv/RB3PId5xt0hc1eVxNB2VldnEyIllqWFBGDoaIA2depxATXI9i
V5J+gaG25xrI/7S2B9O+IXBerdxEDrAv5ZtDuJOdiEYup5Bd9fFm8SWwLnIS
cV+K2UAIPhQHC8NgXWUYNi4E3JM4frzOt1bdyyd7SCNGJlQT75Ta3IJVOaxP
WWvyHnGFNQSKHZTI0OzQFQ3V24jJ6pBu5Ydo9SJ+rWLnTWL9w+c2iN+AC2E4
YIGjFl//kzbpe3ukbHvkyInliPafUkCSs6SLNW7u0MuOhlQ6/7w9vV/nmkwz
/It70T5GkcWp8mZPnEOlFaWmqQaVZkOs6YPJdBs6FA5ezawrZkh9RDIkpKCJ
xFN8ytJ2+qzdm94OXfT9YQ/ewdvcYVyrkiSL08gJmBR+arq3cyTh0JAs2RsN
b3bJnvdD5ONbm9948hhYCOecQQtnLSlvqlHuh5gpTsObHtF5PjkSi5opTfjj
oKUrRjYDfTf1lJaswZGTJVZ3fffJ9Dt2O6pifcKeIzgDKb4rILefiBHh8H9V
osrnKXb/s7Xrk9UhAiuXNAh/11WYOW4nSu5mClN3nKKjPLDp2XGsw7W3gO2s
l51Nz8p6Y7IcMkXemkpEWjFdXAxtNeAME7KcGme68JBBVc7OdQwDy1MAzfI3
AfP5IfWosR0j4otTJGRURTS6BQS2yPWNrZnDjeC7P6zfHUO7eOuty72xL3Xv
0vD2dt9AUpIZaBT1tyc1WKuvKEA1i5cmjzhO1t4sqgxKnBF7Nj0OJSJS+PsZ
reoTf0rsVy1pVkn5L6plK+p3b4klP0y2dj4y86R/Vvs6hi5IqykhtUyctX/l
Xdy4ODJcVKcJUEaJ10mBxNEgoToEGZ043dMlQgP2v63mg07zHSQzQ/ANi/9C
cEo2ClLH+30gNpfXIZrcgeStUEbvw7JIXy3O2j9Tkga9gokBYiC3ToIBkD5+
mK5724NT0qHheGP3BJ3CPaNV+BvP0BALikLyfbe/lAUFKPbLHi+kbamJUcNh
2/PiFBLntnOiJjrSSrsZvaxQACjasCxs7VLT7ffbGS2Q53fntsP4K4WFryy3
BaSTCJENpLUHIrQH6rjTU0R7zATHHyZb1Pt2CJbWM0FmWneYxmEA5VA33Ycz
tjjJR4FOKQQKvpxSmHVfdEIionmt8BWTKOzQ+7JKZS9mI/sOxJQX2TXPJSFd
cabdB8QQGO8VnW1r1VVardb2korTSHCJDV1aCziRxn0L1/sXa085rSnr7wlD
Y2CEfKgszGHtQue/ReoCcf7dvdbFFEKhcmXKroZBN1obm0YDbABvgW8RYUDv
V3pUJcNjvb3uJEiSmKLjCe0mKQu8f34qFwUpvHop3iMDV89h2C3sxCVaOedY
y2LFj/pZ5VqICPhXA5hnFmLUWTehUWB+am3cIbdejcAkO8nivGUGMiTwt6KF
TNUhvBAu3/M3XOXuADozsg0retTKoPyyVzsbf9P8zcn1ESdcYEVSaGrKLGMR
xrV6fQaysQarRrX2tCWkGimMytkfqeSS+YvYB9agIcIS9hm7jz2p8Bbpo0Uq
YL1Kf3gQJXY7eSsLzMHM0xf5Tac+Oq+ouMP4I5X1J6OQrkiVe13N9WwOZQuV
0wa1fiNr8vmQx0xX6TGAp02vQaaNBMvxOsPsmJp9znlWOoGUVg2nJ/m1n4iw
++vUnyq+EemtGTjfj+3ySzB47a7XZvHnIEKEPueoDhCAoae0GXRht03fHgNv
i5glEEi7O0mjQHu+r/ch4HtG4rXw0QUZaJzihCVXhmdMfk1ZcUWtG27u3wb4
AMigCO5ai79vmJxzpFbIyLqwRLdwmM/S+urBlSi0Ubw8+dwl4ZvHUI8fVOw2
HyM9uBXi3ciJoTdbhzh8ZQRdVcOk1qn0FAsVnJLOsqF7fXyMpviYD3mIlHCR
J/lRQoXjOSIuv61H0GFM/KrGALbyOs1lQKEgI3RhMFvceeUYpobOdfukUYWZ
TnwM3uFSqGat5FAINgk153mKs54de4X1gaHKcl6MTHlB5gR/E4Wj4/nll+vo
9iNNUEYadyE6iQgfEWlDqlZ8ZX63EyIRvZfCh/5yZL6NBxyQDeAoP6ufuArx
3hqH/SH6c7ZgS72xMA6lP0x/jGBMY39f27Ps4y/6WAcJfzRBp7vtA5k71Sb4
4u/ImofwnUolBFK2enohR3rHbTwyyN1eFb1ReaRd7JVz94SvDb6iZyUw/PfC
JgimfXioZboxBdFBqIkOfIz0zFDqO+aXPgJ1QdNjKpoT9K51mGr1obW+Or5z
pzOMH5MJo07yYOWkXlDeYDmn173j7u6zVpQ6K/mPpu3cCyPRFGrBDf/qLZoz
LD7ONoVzgiFdcGwv+PfDIxei2sNDuRWwd8F2xBqfG4nC78BMmHILciG9s1Hu
0V5yRsLbbIeuGsd351AGYs5MRRZVm2uC4sEtdXdOd4JA+feZ/bDGihGgM4bg
xpYSRgHqNhtcW/BN4C86tbg1b7RfVmiYpoO0ENYMNh0hKwfwO4tMdG/FTKwS
QhlxFHvze2YURRjnozm6sOQhY2yynUs5S4aC+AKIu8nQGtN5MyCgj4472hiD
7j3j0uvZu+B6PwUZBf8jc6APu2/Tvqeq/sjMvMGzGNuEsHG6WDKzbXSkvRzH
VygVhXJRGERB8anFrBNgqgWM5G2uomatsF2UZqLNynCIBB/xp0A6d9uk+K9q
IL+fv923s3FEzD5DxNgcblHi2hU59xE1ueJ0gxdLzkyhAR9TSZftQ2xRZWXi
1kfPrKfPER5vNC74Oq1EvrodpXMuUtel7NrHeCb5rrn5AiKVg5jw6dQs1dOL
29PG8Nc8PiJmTKKuTMT/cuArLYI9vY31xpcwEYZE7GK4QJX9djUMgGXx4n+U
jKiP58fZM3ZqrP+fjC9BZdCeTOKZRZY6iR+jH7hwyCHeoqXaaAN8qk+nh3f5
QR2f0YwP8TXonLDNMQwdsvmEIJCvgSP42gHZPPqzkd1XZAfphjniUEk0D6rJ
vlA/paliRdwdkD/6q7U5c5yx6lXWO44mOewBkwv+ZFtAzHYmX8jYx0JqN9ki
Bxpu5MjqYwcJouu9wJZDWRYvKUvY8E07PLBwFDoG61BDXk+eD8oDRmM6utW/
v/TggXEh2sS6PLFvBWak44cA5lzC4pw7V9R9dKoxwG/fKoZE7unJIRff8OPT
2r5+Zn+diEdFoRvu3stGY8Zind3H4sxHJVXr1xo215qeTJw44Z+E/4wzlBgS
KctNwHuZfOo9LL8mSLgsCr1CL+YzXIUkgKo1e+ivEIaVylvmV2NmKUy1+1M/
NFnYh+aQQVIldk3ltxefPqnDAVFO71bEY8+o9UBdymtXo646rqzXNKLCLNBy
BffUg4cgRARyWu+YFwMaHgP9IJW/CAc5OyIE3dBybrL/lxRgDmooszEV4LAx
HfT9zNtZz3E593egQO5Zwm+HpEfJ4hH7MhdRUmge9jalC4lLQK6GJ4zncNJ1
yWIKwlroNF9xgD0EeKl/W6ZTcoiJt2gmh/6K7Q+xRP6e3q1VtYkRQDQRKoio
wyZRMskxKrlqAPM+23vC2cz+aFDneVc473jxN0DcRVrdaRCK9teyFLltVRMC
aO1LAEiowYLTuVwk3MDZeqsmNZ9UqwrxoSw6ewZmJm6Z2onGRflAuPBspc4g
DyPMaaEAIT31dbak1AW49nl14lVaqXM2dBARVHhb/PgbBKsCLJqKKsNjlD0S
5yrLlhAVIttxiG5nkB41z5bFueG+jgETeSsz5O3tdBYyQehF8jTEVEtigXLp
wup3P0AzDs7JkTSyIUbymiNxWahDiN312iWLVDSB8XyWCgD8hG4u3cX3ARAe
nKuXf3BO6GwgP4yIgPPzgJvofGhyCWoZY4pDpaKxwI6staI2M1MXiKekoEw1
cYYY/U13QpZYrzf5DygcwwZ2zz4gmmRWXj+XIXkoQtn4d/5cepvXaZl1L6u+
rn502T0fk89zIN8SyDOMmrPtCZwe7kaxdTYqhAVVir/HVwmugWW2tbwnEKK0
yl1CACPH7H1Aw+L54tSqvbkdilcD1XfuMEGoC9tZTqVW/gYuIiB110qjG6Rj
O7BTVhoF/EUxIW2tHJmMJ99n1ZnwOx/8vjfEHRIwe9AxW+CJez2vF2dLsDVb
5jugMaEmz/7lm5WVD5hr0ZqZ51PnfP9QhnWChGAr9VEftbxFJ4H3TLzQPlne
WWPSmizr5IE68+JroMCdOtXXUYVsadGiWul9wwvfuXpXrSFnoNrGVUY2n7JD
9x/HlcAvSvs4Yyw2U8X2hSE2ZRUkGmkXOaYcTejzcWbbgbGvl+2wlKeeTGu/
E7QjCIPomwkuiOSDde2CJouVhD/n04ciJ3kU7HrTs2XYsLGrSIJPVImMuDa+
p7dMYg2EoQggWxy1aRTDp3GgM2aeJhCSWD4Dz0Q3S8ENyCIZxhMmeNw/mZeV
N/NELE8WuSHyeSaBum4k/mAUs2fCAHkMLZ1QBYvNtcNWstg99sFo62/ZtxVs
iGFtXkOTf49fAkQxwnIaX9+97/wRfw5Pt0D/6nKSYpwnNmW80l59Vld+ZlnO
R72lma4mqOkfGbAR3GWtON87FGGZCVz135lLwfo7lHlMEPW3CUGAV8ryjn9I
DUBuA+f+jC/5IeKZxT5IeebOuiRYNTbx2np+fcIjZuHwpRqyQzncMP0WzqLu
bH4U6F3CnZk2sKIVcfF56yE0ebAnZxo2zypemYXRXsD03RVIAxO0+PPjkfJW
UjocW6ARhLir6uFkIidz7SJDOaWRUwWbLLfKKQwdcRpPpZY5RGvkPfPvJ2ij
spJbX8+iHJfjInb9NOL58K1X0Mq1pCHSoavHzHAYUaV8CQxhogAjb/95MxEV
MrieNIhxGOF3B9w6iQ7Ewffe7BSLVEfZmOaErHpqdSrDhvU6zijqH8MQ1zLn
2zIKe7KOYABK/s5HCv0An4O7dRK8Ry/wDOskhA9LlJxKib+HUAX5C2v1/j5z
/PCbYfmyQQdLFcQ/xpk9OF3oRQVL+nmo57LutK7ro+YDEyHQ3+l43rBdMojH
Omt/hQ5hBhRtzIq21UDWoSKpSztCn4Q5dcu07waEycct7ydd8CA8YAZF1z5U
GZa9MSOWXnI4QceG1frezi+iOK2+CC1Gkx4AQBfpGoAX3N9pC1Le7TppmEHN
0zi/bBmtVIkF07+8g1LqJn6WntZYURUdOoDveE10mcocjd71pbN4G6uR+kX6
ckLSSxUQq6yyZabr08vrQ3d1iOquGc/Nup/v321cmmjrePn3zd7f+22EeWLb
aFOL3yYPga52wRkEIXlTEcgshy5XF1k9el+vvKDpbAONc4ddnJsneHCAU8+H
8C3qkFX5eD/d9f4OVFS8YYrrcG7HQuLO+dboyJekxlhvOtG4MMpdzO52zF91
Ol3hqxnO/Mk7rAKGhC2JXKCJ+mPCkDjrlWMJTXKlstzciLMRnymkQtzqdLMe
l5yzgELM2ntuM8XvJg/UkNt5ZwW3bQmtLgrtoBilcelozWpx7iiJqiLvL/bO
zfuhw6QOFYUMXdb7wqE3w7OedCK1jufvwQHPS/wz/56L+7ABgTLTJBtRCHFA
iNPNfZZXytWG/DiKl0wkknVfyYWoOOLnzQiKwRlvAYKUjZOXsjYKc9y+AaBa
wupUBb0ENMPRwrW85nvZ+dLLPz2188VHJD2KxOhhRofRewIzFxdji/Wcq69w
REy2IGlLFLPCGLUs6AXv3536QnMBYytkyrYr5mbU5h6EYCv3e/9oCQlIhOOy
/QeULuDJG0lBDGJ32dgTjkAtEEm6/KK7P7mR1f38x3j3CNqXQxiHwEvNEm2c
fPOOaquUJ/5/rFC9sjjrXeHHBh0CfG3kY14mguGaCDoGGfZt2WFp4SdDaOY6
pZbnC3ry3UI2RaBnSiUDskKSnDyDd28WgYrdLZWn9ip+k4MdCDuBkq8eRDjA
F0K9eLwRJclLYjgKKtzLphSDnW1uov+45bzsJxEGrmMCJnNJUbtzePqKW9F4
1spSR9iN/Yq8I0K6Eu8R9/BrnbDF/TFbjYPcgrVKHpxjQ3B6AEXallIJnNcD
Td35gNSRFFcQHsbLncfzgBnveqPS4EnDN/AHTTKUj/vUqi+15YqrTF9JAg9C
8c7Mh9VFFoXMrZpAhDkO1hWh6wfsgmSmBqmXIT7hoxhpOQdK9qQpUX3TLm7k
e9Hv2GncBx4inC6u8mGFuXXVYR9Y/O/8CLIoc2GzVUYV3UfVGgwkUn4230DL
Hbheq3Pf/5lC0Z9eOXnyc/ER/rMzGVQEDQRaWMT7qkHGMZikX1Tp/QcZVVim
mV7wlxmnkZFczTF5IuVVizezkWOoz2GNKtp9sfzzYOnbpFq/mEPwykIdRHRn
OrNlKu++1zI5W4YZlgWfoem41JncT8ZydRiUyfsW5/BV5mHzm/L+yvKk+HEF
/F8w8PGoSjgwv0vrOTIHSuHknvkRFkNY+9GfuglU0UP3mpzFHgvO/TcKBcXy
yu/SeKGt3ey2ZOC/4UhTwD2ps3hWneizioeBNJIz2tEX1a984LXVrzK87GX6
0hgVo2aHkr43+I2I6aOxlwJxOgfP092pj8zRQQKmjuePkFi1Ln/DdLPxlVzz
sepv8RjiKmxvUNYyF/U0uKJ5uDYMUnAYxCkmfB5ucM7ofi7fGIvARIcIFCLV
jTOM66nwwMgaF461JtWoaZJgF5CED+Z3jw/vs7EIOLedYlx+jiB7vF07+p+w
uZ5hSKlvmxUt3Msx2m6z8s7y51DGEBZ1Ci8m8nEw0d3VhVmeENnilrgyJECU
y0A2wZjAszTD73KdDakGe6CMivLDWidFwSrCe4WqfiA7vyTdIz+6p5nqVGZ/
KvdzrVetKNlkyMp+SrGa229mfcKdPZw/mTOAX6nmJoUx7z7TVOt9r5r3p1ix
1zJmXQATsuMBW5nmixROyXqfDSsoAkl+b2bmj/vLK5TGhSRkkC96fJY8RjzB
KeVY6E2TGHroHuYbFaSTdz+YwHwptS7+Ixe/79v2M6+Q13tetPlVVU5QCHOG
j+62TuWDuf+fJ21XeWPC3ybNYYqDC/UEGtuJOvqIttC4hayjVzAaO+93Cn3B
Een6V5exQlXuQTChrkD3y0B0m6HyPfwA7TWK6fUPQLvDlf2jrTtXBYEPRWdJ
I6DB8VD5FIrQegZsSyZrHux+hI+CNLqm/PX5LtikF1XqrOm+Q3gJ1uynuL9T
PlzsBArJbD++az0NNWJI+pWl5ONtY7C2N/yo0n+xrQQtZgwtRFPbgDkunivZ
uTDnd8E0zM+92w8txASDPhJi4WrovsEydRT27LwBjTyP2OVqjPIkVDPbTiqU
mU+99CtR33h7QQpEPEwAGUj5wgWpU9TuFbm9dncyIvaBDC0/MRmnVwT1r6N8
kHfZ2Gpt6FlnAu3oqVtKqzIEI4yMAkPl2Vb6dmjoJDtSOXLZeFlHjgZTBAJO
SC+dWK9AZWl0Z57H1OysSu/I0kpfwB6rtBSkLtTdGV95wVIawJTGbEhvWkJ6
tUafwUtxA8KMuD81pAg+K1qGlHUchdT6gI5tyg5zV2oZIP4Wj+fX0GNcrOQU
P9FI0AT/U98ncPnjZFdOmrlCUt/NrI1bqJ2L4CDdMVHLRS7NIJSmRpToVKpz
RDBWUAcalMxpFi8xHHuwiZmNYO9kHZhpwTqV8y6yr90UGGBW3Tj/ZevX6pL0
cMbli+aiGThUQoeefFeKH+S/tzaJPVbA3J09oq4xPWry1Mf7J3qG347NKA06
2rNmSD+mPikP24DmjT327f6uB43eHHM3l6w+PDEBm+H+U+seS45/TBcNg4xF
taNHknWubhbcUqm5+DOgBJ7GV7VMfMxaQ3VlLfbqXHrJuohIS4yhHt9z5KC2
lu1QwLy+BlFczLTBPBkr5zpmbKzFLwrBS2fmDZ2jImkPeYgKgDXSN0uREbFd
BqrPt74sSanLMRR/1hH7cbI4gt6e0eJywTUJ3ItTNP8PSgADq71Dl+qo4Puv
CkA/lxceJzz/KQKljUm1k1+Fw7b8MTU5MoKx6PGvQK9fbLxi4X0oWbzqMLyj
AW2QpWpe78swr27zfF2YdEelo1lXyNz3kSzzoScP1l2fU4py4QH4E2/JK0CF
rvumHSin7CRdaTfDPTLczFmOp5eU4VngjSdt1H5GnxLS/xJDP1uvf3lRUkSC
HdXBA8B+7L8m5965tB47Ne//D6QAYFXyWChLFZ4+NCX0GDrVUfwlo127ehCX
3UWCvHv2wjES6FoB/hWBSorEhPhbCBELg4xBzyNCiL/U3a3fjtwDluVA6qGk
R9zo5H333qH3STEEHdaCDSHwpsVBKYh36e5NwLVsRPTyk3nZ/4Jq9ugQL+SP
7SV4xgyw2uAhm/LDnfLS9lhjHJoNZ8e2YJNLBLpxNiedkhwpvJu1GNsD6yEO
9dhphcd0UIlfWx1zeX7hY+6YNVYogqfTMBdVb0pvOas1DwqjB2HHFiKJsDQ/
oQmQaoIxweer6smzgul6Sh+vJDJjF3IlYTgudaf3f9l75LiP8CWjH71GybiO
NKL2YpWACR+qb7JetzJLaMAWuXBdRivZKyYjh3b3j6f3pfb3GuoMPIC30f5F
oxIvEUaRndhhwFbR8QhSPPjngmtfbmLAd5+yYgVLBKnd1eZgTyd6viusdkmH
H23Vwnl8DDp9K4rHFWXb+GwUoadRqTx3UCiB2bZgZ8gYLWLxtPKlar+J1JSD
7bAyWovMaHw8Lm5W4rp11oTCfN/+mZTs2P1eWdKPFp/BGJFV8PhuxNmKTcfL
2RffSe9jjt+3XLxHBgQtRoG0EtgJKB9/638JmgYEh1K2CHYP5QTg0nPfmzRw
AKIelh7W5lZ/7yTG7F+KK97y9x1657SCrQ2KtWctmIDVBaLtkrhwKQAxQWta
TGawBkGy7YXboNr4WBdCHMSWkBO8FPGKGiuUQgzH/jfksDXnW9JwVlpvHwHD
cZQXqAHmIcHvqwZGBAqRFu0Xn4YRKzCR8U2N1Lt6g3sarJQSV3UPmcCPA5GM
iX9OliPGHDhtwikgsFKQjp/2GpP8Qwx1rYSy4RgZ9snV144e7eyc938oBBCQ
VEuUUlI9IJEbfDzZ+6XAG7rjqYsyX/YI8XWfXZbgQEA6EzbebEW9Mwn+Svco
VSfzh8QILMIDCVtv11VtHxLYxYRE+qvRKeAn5vKn9Cbwpzax3KEFCIhAzhy+
7euks/xH9QOSSUNKpQjfr2LMXU+ZeTGGlX7BVpaaYA6FIv4JK6a0hZL53T3D
bswieEF3n4dYDiSFMfd8GSNgGVW4qnpJ+bycVr/8FJNGdjvx8olFGV4CqL9D
p+VxD+cuF+h2j0O7KOtGwwABDPyDjZ86X2xtpnuiLnCDgVVdXL2/VD87rgKJ
kBQEoJaaJ0u99W6XqqZS8E+B+ZsbE91UQTb2pHS3rLWc9rVHFywiXjbPZWYw
r+TfgLP7VmlLzcwB4g2SnZ88tEIksQYGhTqN1a0K2WSVz94o2gJYnIQND71B
lYb3TZyQi+5c4jY7N8SxorvL3YnKKJMMOfZ5BYoVcF6oDgr1hWUTPLpWEqEb
0QrauL52zUg9HhkyZIc73tZ01SfpcGjvHxUfxCYpBuEp+WHfsSr+mrHYjdtf
xezKkKEiUd4IjtFb2WibLWWlZnFdjf6DnGl4OlHgYFaSuoFVoKFTurTF2AEJ
f/NYzGH0eqmMgia32Pvo7N3M65ud3VNah/iasxGh8FSg2/lSXVJxxB/0dzno
TUpiyR2yKs518W6XRjoyvy9G6hw+My1jU1lZorIiWRosvl1torH/qqcvgZfV
nyzqhj4cqqqUHcav+Qb8gzNUFObqk/1IL+BMtG6qZP5fq8j+9F8aXcUk8M2k
7s/g1chB+VHX4ZtYyXCKRwAiBJOjCVrkuU8EJBvc+IhrCTtEFxcjC9FRafLo
UIIy+pH0ZIOoF1H+IsFTM9s7GgKjXNbd14dz3fJDp+g1RYHthVzYs8VouAVi
D1pX4BAV7s/u2cBnV/g2y9ST8HQv7YajF0DHa3GK5qMY9vcspsvRj+L6XnRq
1XwO95O5Sh74+5JgMq0cgBXbfdyfl8wAUAH31WGRVxMFPPqTZnl9RT8hMGKw
xX1jWtiYBmaw2sSnHm9dn7RtUjMQxnOvpEpIU1YndnAjWE+p3f0kmmlNIOK0
dXMTyRt5lFvXchN+tJoVPphncpBvPoWIe7oV4QJ7hi6PjiEBdO6oWEbvpXDE
yeqcFD8/PUCOI7aIgPbvwf57U0/qCXqDLHzHIUZBCkI3N+Yqy2zJ3AyEPldZ
18XY+2UuWPda4jMXDtH3hgRTLkgXRm0EF41iVprIk0y4rDvSYjUrdJbAkgt7
PVXLMQkKFHHVn6gQIPl8bmrCdVTQ/VqwDBIZsM6OwlY/CDzAaofWChVr+0iw
z8/xPUcB9wOHoyjUNxHTAqaeDHSaQlqPf0SuLvxckuaYTXs4wPMVhIjEwPJ0
AIHB/Du1mS9C2vG7dg0brgMl/ySfN8elOSyvf4cO+gYFwJ4fU0+K+uUmGMrJ
eFvIY249KCGNfaKaR7a4GhNtR90wn8wgfKm2NXN4F87Qc7OEj6fk5+bIXNCP
g81xDIy/VLij5Bw0p15gb2VuVjXUr8dry8Qf05tUqOTyKBRH4G1QcAudxsXD
DKKeC7MQRwc2c0rB+SY6CLvDyQzTpbxYIBgO6Brs2PBlNw4I8SsmGf2RMk2q
Vebuysf6XYG479oSHkb0HaVp8bfp5dg9VegsAu/liq9RrjOK6nbr2ZuVezG/
+T9gO99XvCJJWKFlg+pUwTbaCmpaOmxTaOqRD98vZN0wveY1HGI5jQXsuBWC
aXWbYVEpXEGnJeMJIGJRZJ9x4C2nQ+U7Xl1XnhO7+3z833Nw74qa0y1XVLkO
W8NdH5U7E+P2BXExbSKGWQiAVMRnl94n8eBb4aA2JTh9KMhm71UdqfhFugx/
tto6tUxtJiYMx3Lgv1Veqt27Zs5e8ToJLnD5gZnnzZHwKyAg5GnRpvCZ3eXM
GdwV8C9wIS4FCyQMrd4rRMAygaoDSW4kWqSerM/lbe0Qhx42pvRnjK1HjWyW
pEdrRID4qaAgFiehLHxRfd7hqb9berxkE7SDQ3P/Xw1N+nDs1NQISMmy2DtG
QgynBEsogaCZMju5DEoJ6xwybx5C8PkT7TuUG+4uZipVJlcqLSKQF32SEMFn
lxdlBOXDP8lmRD5t/5D8cxz9WzTro8TCGq6fViKUxeV7pdnINmh7XwYpMwvy
9+/wZ0mvq3g0yqaQ5wsoK/z7TKiYy2kIcBPOTgGFuyjCfRkJ2PVnRR62J8vI
QD5jGortKBrpVyecIfRKGBB3Zky3hlosN7k7KqoBNV+ag45q5PCnXhR+M3tF
WunKAfNr24FVdTGH9531UN1Bwi3QS0T1K6eF6h2nmmlWAxPMaaFAxk197RR8
YIZJKSDO2M/0vwRdghXEhwBBMl5S6IlzjJsqdopGuaTvg3dy917PlwMD59sG
euLds9kS1iqf4QsXrh7K7Dsaj5i0SdUCAnpzxBihDMzWlAhKHtgUOUXa3IXf
3MqpiaVOHyM45gJdhmT0FtJz/eAylvzo5K9A2lgw7Dvxusap9jInkY0E1rIj
AW2LNBEfUDfMib0w6Ju0gkRSDQTZJ1/H0xL9jkon+HQEiWAznIg8kjLt3XKt
uwNhTycAdEIdK54D2vtRpfoDFGrKDmcBBeGfQi0hkdWlMMtq1P1eYH+6H2Sn
jBXWEeJ6gyhgcGsKw96WMHwWDstlvnEmrvTLZzKB0TPJPrJdhBVuGK9d6T63
fuEnkTiF8F+fZ4+38ESwvUMpy9pKAiB5kr0gQrCoXqHroMVQ7L1qwd5QVgMm
OuAgMxMC+fYhecPSDQrAy0q24k+CF5d9jGZDeHJ0HCPyZyHuyTyQatiPhGu5
89zHUnhCJUJf4ir1WKVtgP8AlLsIho+oesv2tCjj2HfeEmTTp6DY+NeP/5pT
HppwCyixGtU5+g3m5HC8f6/Lw+pxzIVADaFHBOpQWq4GaIDxCYQkTqtuRQbY
s1yqADUR71XRdeK2SqoqTnaMBMY2dg8Ce6OCSf/q+Eh7hyFfD7LIFQ1M0tdP
BDT8B+p/EbPW2ymUVgkj0Y3Hx6nMGSL77yNlhbRdfssfiUeLblMlvE4DLcSF
0HQxW390tJnpZWnT4VJ8HQf4SE/gdmndjaHoRyKAiHffQdDBnwhEexZZ8I9G
Y8Ktsbb9gBMCerIld2oDsXud+707CfxR0d3VTF+gjRX9waTYNr5yAVvzEUai
kFd6xa+XwOFQX+61pfe7/CP75AfXl89bJ+0Fc09KypCEVVSLyuTJqYX046k1
abD4l0i1SoIlGEPeDrma96rnbfMeA7fqhp7Jkd+Wgi++2nk8lzJ4sI/2a0et
bZMwHunZiv05m0MlFrK1szPmx0TVZ+ba+AGHBZT1sDPCifArsnEb/Y69KcCf
+GBVBgn5EGt1bKMrlXZISV/FQeyAW8pdSguINqNG1tVbYXzI4/JcWi6+WlWB
lxC+SscCHOy7uheyTmg0Casm8MIKZ740+6G3upC1ctnCwX5osjBrdIhA6OUn
biKfjrQZiJMSHsCtDFPEMT6x/D72+tuD/aGeAUDb/Fjuprcp0cSDsngoe4mH
X/hrgv/m1+KvQJNeT4bU5sxCinQwB5Zx0EiyHuHJwSMzaMF37K5pfkSHduZx
Wc6f7mpe9XRVUymrb/DGC2vdKQJAR4fA+iP4i9kEecI66fvYYXRwj1QJY7tt
HhtTvF5T6pIqnw57YJY9axZp6eIQ3Bm+JMnbPtIpWsdKtrid5toRTNdFO2yB
1JmW05AAsza212MhZr2ClUZpFsceKgJ7wbomEkVoStYEYcSJAdmI04WfSypO
82VB3fIB3B8DpGBSq45De+ANf2IWPY6V1mZg1LryqgWSijLB3dVbESp84ahX
hHrHv3q5uimWTK6O3PhjUe8rlO0mPIJRJv735lrDSDruCHfA8yzq36ijnsR/
EusGVdMpL1jTwJMG6WlKK1KH/woDtW/J9LdPp5mkt36tc4hmlsoHqKWIS50j
brNaD2gWl6lXIMiutpT3JA/GmXF7Iwhqc8DLgxHI9ZOO9kl0+XHpysLbB2/S
NVH/EzLCV4EvrzFExEtENbutzUctM6z7OMcWwS0y2JzcS2qtv5OjM2geIsN8
FKyvRb58H/TxagRJEJr4siPzLj6cNL2bIeKW7rXw2o04FiWObiqmPQ5cqdrp
w6BS4wjpyGe1pvG1ex/5UZlvo4rWTmVNb304pzx5WuzJFbMihwlQV+dv/Wn7
EgPjbWJC5M3gwCuKidFNATLLAPclprRqPFBgbQLZ7nj36GAnL0yT57PbGfr8
JA+IA6tymwPuMKkYnYrgMZgDZhl11JyAWsOXStbrcJVZQTIW54YLzTbxoflv
7Cp+wkQdZoMYV6rpZEgEQ6guN24aHgN+Zy/IxFBJPvs8DWrft2WGY8sEUcF8
k7lMI43prbd/z0UQiidOmImUDBiDze8UI2SxYe5ThaXRxdLLey/3OcArgV8n
Zi0+So0KpVwuCzoDs08frqfzcxTtKPp8IthNKd64UazypcqWb0P+BeSWSgmb
zSrbrgD3KO7K26gJJG7Am/pnXI1j7uhw2YeSoumWl7klDoh157aYZA4+EzBB
00hFNQjmWPcd9krF79kuDxYRyKyTJMwQmw6b9ht3RM4ebw3ZD2HQOHEdhVdW
zelQ1mB9CaqGzixT3Zps/0Sp4+i3stnlNWc/HsD5CmF14s6xN5rM+NhV46o8
Evu0nJYfwGWNE5yWfMRb3NGNcHlnRuCUGaxCkGERLNxuMb6T0Z0G8O8wtCZV
juMyHAcARJDGzrWkstcqlWMhAnlX4b3E4k7t4VQ4X3sS9EN4GgblL04GYZG3
dFDADidf7KFkFO5eoX1RVA7OrSUYF2Z9qska59RRPk2yH4BNms9oxWuz79qd
b75vjit1tMJTTiUVc1vWj/rL25YEt9C9IfyzuNmhkEySmdJw6cjcUR4fWdAJ
6QH19pWfendDMPv2Wk0L+G/ahPGZx2wbLufgfRtbEKB515ApdGiQe3QTmRnv
+zeaSbRunMKsuqYwMphXE5i33m7Im3qbZdj6qOOarFt1QmSxVdC8AN1jxwVa
QV4zXpQ+Pa+7W+U8Hw9zJHrFi4l13Ns4+8xciFlcymuAO463P7Rz4r4ePnbc
krw20Vh+z5EfRlhb8VKJSXm1STUQ6npUwyvFmmiRA/NE7ZEaNNonFXWmk685
VigS0gpvt98Lx/+w2F59jZXNqUT5SmRgVgvMeYUTGbgzTFfmE81SO0ggyBoG
HyrlA6Q4/xP35GNs9rhc8F2T0FRutDB+fd97O6hdwqzcWyh6dqcOnUqPMNyT
KAOwForThrPijXduTTsi/3xqID/NTx9oIGD5NBSjy0pr7dHkx3QSJMXKQRSt
HWVd+v3VR6FxVjODKcuOah0cyY4A6OOjhk3j8sliRBiLkCVpTZlSjuS5f+s3
aeiOAfaIqTwYUWHve9mUFFzdIoM4n28zMxWvIUEKXAIacDn0xwsOVvMQNdmO
hGwhSbBJLYRmvhSMnLVbsraLP13mIKhmFZZ3x8jnbXL5/v82RH3s6N8NJfBY
xqgXge5LZbHp70xTz92PyaXiW6O2+AFb9PQ1dTP7rx6rn0gytFSuEfbz93It
qs/w+TRvtBGigyDmsYAu8ZrSIG1tkcVKwJ+Hn4mZ3CWOGxWiJwrOB6QOjUDt
F+vx1R0mtp9sPkKKPeENE4QwL8d5ymdAKX5FnyDxnVRsjnyFg5BE1sF+98ZL
dYCYwwsq1WJgGqM2zrUFVhExlgiYGjNyvo4jtVSve+JPN8szs1uYN92XaA9v
bOkZtVbRo72dC7kgOwXp9AZ4XrUE0LCcU/nIUNRzgC7hd9Ef886ZFm+++kaW
JU1Q1BfPXDclPipEUmpW4yYZ7vwPAYp8W6h/u9KywWs4zMazIHpDopba2Srh
tDN0Lq64vxPFBfxHzEuNNzbPH137q08w7Wtk8oHbUC+yEfXK+4U8lgk97B5V
iDQ1i7ja6yRIVhmBabpjqzmPUv8CTrE5WlcL/odfazPvuojdnMs5YL2Hxk65
eZmqt+5J3ciEKGmUxGYC42QaanhufZG7Vi46ZJnZHfvKzAiqYu2blh2dP1+K
I01aPNIjF+AD9tuJ6+K4jtwX4w7npZbpB95NKXP5BYXejKzDQtTKLqgR8SKi
/vpYu7sBEtq8DlwMGmUUom66MOCwIU3AnTSIeoJ4P/14yl91HXVlEth6P7P+
od9qMmiWgzzTwdwk2VJId6HtxrqIFRg018MqrC6QqQkr/gVwwRRFaph/3NaX
PuvZ/tn9ehmFUFml374p1vJv34lQ0w2Vs4cM5L8ZQGX6DRrkc/Un2tFlAPcP
KpNU3fwHloOzanPfZy1RZyQ5niffGik8GpPokc8K8ujVnJWQOBQG2qCp0Ae5
HIxKMXH1pvColgXUEdZhc6k7Ir/heUZb8vnq3pwMwUV4cVzB50hqOAK69B+5
Zddsq9cGT59c2WMxxRxOdu05FpsqUO5cl7zwEqPsfoCN4Xes5C8uXL3QNM5m
0KmLaa1oq3MYyxihcON+XMTiWs+3elLcFaZKAI+PuGpPymgtP8fOU0YhZ0Yy
aMPM64oXCzjLMXyAjfyZwGOtALw4CmwDeNaXiMu9nBVv/J8YLTsZFnkwlu4W
rV8DpURZD8kk8PJU46JP81LSQLKuYnnaAl6x2/jmOdhfOqFA/NWj/XEDLeb8
YmDfM99UDgJvLj2E9RQUHwftZS06Dd1IT49ezMC9CBgsCk6dpy7eHIEt/2OG
DQq46E3ytaSWYisliwBtWJ2vX6T2cv4dWJbC2O2bMkMI1L8pi6xeyFK+Nvle
lYkY4ZYEd0+URGbKb2ghmUWvYxbCV+Nz6VmL/7u2g7Zsm1wigX//GSeLf4GO
a/5PgktzpdCqSvA6ODKjuLCT39CbiEMD3Xt7SIxhrIJSD39h7phVzufWRCR/
S9YfMNjHPtqKaDw8qXpIDuAzb0MdrXdtx/2epUJjLgh7CrvRZCIinDtAVtgH
iDuuxCB9Barp1CYjR0ZUwUzqHjNeB61LXjgiRuGK8mFgm8dlcVmrgR0f5I3Z
MiJ4ItIa1EkwPUqs6qU/ad/OrAksMtR7cYKsi3Tk80S9wPYQ3+/tZ57m2Gn4
kXitbqILMnlK+4zOQ6n4jkydlhi4eIx4ymRGwghvd2mbTlTWI9bHKaYlGng8
njVJTBaQTmVfH9xsi7T2pUXl/ijUFgTV9inLAwA7zGLoCUzRiBsT+Rcn5g68
L4nLq9uvhwNILxJFLHBy7paARTXgMhY7WxjGJpH9MuRDC+rxyTv/72u2mQoo
6h0pkfWeVNYW131hMmwoHjYIoEw661qKySYQp6xg+Pvf96qpkAb+ZpfYtDwd
F1OoQJ8HiJkhXe2yAqZourvR2TX+sQQBY9q3FLdtAISWGxGZtdNHXjYreAYT
8rGP7fMPe+dxNHeuhsU7tiR0a0OUwxEhUR+sMaJZAAq7pHUnSKMt75KiQ/QL
y+uzauPvLSlPA/sd+HofS/7/ucOXlvxQgEA4L3NsEKDOd5N6kZ+oXoVmSOlB
4VvuyX4rC+IbY+rvVX2+Tb0Uv/lcXSC5Fp15wThG76ikzhG2rAtRFD/sR7D7
UAQj/+pQaNB47qJsTVBpf4EKtssZgxqyj+BRkkOeP+QiUnr3G26FOgHHPB1w
Ut4JEnH60xhECf7M/D/a8iy02+H+j0V635U4Sis8eAXJHmHPMPQ9d1l8ezOl
EYtDauXBHfFzV4GBT3fwHnoNC/xzeeTce5sH9O21ziowb6nHfIKv8B/asE2j
6mgPLv0S7OVoA2h4UWTKdeoPy8O9z11Dv8Bj7UJkpJ8sQ41Q/tIBsN/iqKQf
z2hGtncqsi92X/ijLmWkKES7P7Tl+gwJKF1jfQdqJ0KOqEMUe9mOG4jbEGRt
xpm+3CPJPxW5Vdvbf8k9YuH6Kt8/+j3NEvxA4cjatvhlABN379JyqKgMaxOo
vw2enpr2xfkmbS6CPxqyAZuEFXnHZiYJ+wdfXUv9mYJMOA3TM8nghltucGXk
rH8PbZaxim+TjPTzJzKBK6I6FolbS11MOeVEj3K/+R18jhcWY5vp3qUwOz0T
TmeyXzI61ZRySUaJfcQxS9yL0PwBv4XMJuMOD6BMAisifvbSIulVkHuqoM/r
XTLg8GDbdyNvGZ3ncrg7QCDyfwz9ppCHnnboDL4vDNbSsm99qzmcc5LgpG9G
WIhS+DiK7vge8+iQWBqLjNQfGiXcGqRc0If7r2f8Eqi9JSYaixJUzwxgFBQm
z+s7I0wFXu6oIYt48H0oA9TOD5tlsrJy0qmLqMsMUfYJjHBycHZGSoVtars7
WGUxJh8x+9KmCWe9/qtphFshHT/PSe4z2CPN11AVaiBeAHaZXV0MtkupiPC3
PNIvHN0TLfHgPTZefMQDFtsAmdMb1rRmuKamn0uYC7c6VM6jNzYZNHVC6EQe
ppsZoxwrz6chyiV4K5rqKqWXoOcU7rrDsNdK0goRcoGrm69+l/287S5QY4pH
uYl8aTRJCxALF0UTKDYCEuGpQ6GzRRFI7OvUU27QNzqBiu9lyF7oqXmzsr/f
jcnj8Z/aEFJvSNujQE0YW3cmAaUpb5j7uzM+SS05winHVn5qZJUI7Za4OmAi
vPDW30edIYwDDu5X3+C8fcGw3dp49hXjrD/C+MWIOWlHPSnvNmf4yzajsEfo
Sr6LSqkYha4XdYCTw57gWExZ/MQziDHyw8k/txOYxGxeGJZxYLqpYpP7wAJf
bDcuJabYAQeJBlni8JdP8LSfO0iJTtGKHqT33W1G8JDzccTJSgpFnTZdwXwO
tMOWt3UF32zp/X/i5aonFfHrmF1q8G5HPuon78iCIwHMn4w6ico9p0JnCkhE
HNicDmli/XfU8AyWOi2y7DIJXi6E3dyGxCniLwCeOcSdhS7K+s9EJdlETdMd
YkJ1gfvpsytQg6h2hzEFq2DHFS9k5ic2L8rJy0DxHKs1PWnlMMozsLQJm2yU
nGnUPAOH18I2AT1oOyBAUCCuw1pQxSJ4n/qQu9eYYQEfuoquytHZLxcfkQ32
SbxeXV9Q6xufg9N/9JvW+kt9P9tq2UhsTb2AmrIGB/Ms9nb07OXDXKETT67y
ss1aNrpEnPOj2d2djbAFcfikgpNzrFj01zXoqGbObIIw9B3vN+gMSXnWyv8n
eIWccgxopDXlaoS/chVvqqce6fZVVNN5HGfc9w5OJJSj/gJCjyc5paC0SOQV
nsS7RidQShDtFP5qWhD+Srcf9omfDGK1MVoWqi4sqhN2hCTbHcRlgLTKV2FL
JN+2ukmAvz5N/tiQi4gIcYUlLQqCff4ib5Mw6fGcLxyTjnIaXFecxtPVFk2K
GJQyRQzlT9ynnRA3ssJTDz0TGz8G3Ob5nnyPmxjY0x6wgfbGi1hXoISVt5Bw
+lTbxtHj9lLBxI8RtnM/GEUqmma+EloXb4p1gGM+ZAlZ00tSGnTJMX/XKM9W
HTkmVDxvdgL/LP6qalUlPEqFroLrg4rrMl5MQW4+3ESEpEV73ESAGdiekb+S
vekQqRBiNtyUUOHtI6i4gF2n/Yx8JQzujjSbhimDwmPRsJKpgj6hI3bSR/uR
2Idk5nS4P+uxWW+M0KISpxGm1h9hvuvIvXfftJ8rayCqllkNOXnnogIUq4Mw
gl9u/k8Ais7UqMWAqcl3UNCZJI4Ps9/zIHZiyXpctFMld1VsBXRzw5u8AShN
OBVCyGf+unJIozGeITEoHIZjWqDkJt0pxp8RIjsDZgQrAOP0PHGhW66ni86V
GjYkhrCKyaCs+kGV3yaskosBF3dXar3GnF4p7tmh/TeSZXp3PuQFAMy1h5ZX
/CEt7yeW8a3ZBjwik67k8UhYLm4apixfsppdsgtn3oYB+kEcIbYxsijOU6Pu
vgEIOVWp5FiDqi4VmPXjJnb2FBor0Gm820vEHV3MgK+QVxFixnfp2HNKblqc
Dc9ElzNsdtiGhflExeZ3IvQITjFbxGddjur9eTQTB8TGAjV/qWaFpQrjRXR6
QWlhAbp59PklMNmVAJJOge1SmxhEYuLU9KLoArnG00s5UbeZstWGYU4SDrku
7fF+tBKab4SNTUJ72EFidixjYHdImaFtw0kQvKbjPjhSR6w2J+wNlqqFv8N0
b0XymGuAtqL17kai1C2GPl8fgM0UwACTaEbYrl7R6WfVmUNiK2B4AGS4/08l
k0AbSvyUslg46J8qKZ706BEQ8ueBSsrT3TEwVdSIIMBWOZxk6U+KI7mX+tOX
ip2E+DCiZUkP/IgS5eW4PsGZaFkNizED/Xi8ES+D3qpwJM8UlNNfJvcd+xcT
m7JlsNwy3UhTWp6Kic/BcuYEL6soqoHRZHCLdIrDIbfsMdiZn8JgjtJCqqwu
ae5fzJs6byrvzsEidmbRuG5Vtl0NArcEP1JkLdtQ28L3ZWTtdgPE6nqvjIPp
m8Bp/A0AjGuUwPloe3OeeX+zcWDM/Zdwc4MOP9BW2wSiRtJUMDNkS2yQRA4k
PBtk0OemW0ppvQvlhXIVzpEyHRLHFOydV+V13ETzvHKi8LN9oZnd6BkLa7K6
epLku6Rj80+bdx0qJ6ouQEAzJGTQd3Ot/QY0Ytp9O4nTyD5XlvB288Go1n9o
gbeaIujjB6/NefbNGUHHnLk3KZ7ofbaQsNNzB+SJngKvFuoQKEkTpazIdhMh
FWEF5Ql6uBcQCemlDdyg5Hx7L9VNBs/8SHzpZ/L62MD5Lhu9Yp1gBhaHVEFN
/3iP851X0v7gHCtYtYQ2Dr68ztWbl6288ME1ZSiAKwPFFGUy+8MabfYK/3M1
4OZMz9ntcNmMO8jHvow8tjUT6yHF8Rqmtj80iah/S1aABkQhK3S91y+aUaii
aqj9DpMROU0HJq8A+wbJWufZuW3HM2SkmmC01xdBOjBPDgy/mvrGf0KVtfcA
rVbS0/wgZdsyc5chBbXSIGEaCkbbNR7w7ZA1gIY+Y91QQ3CP5w8X6Tr1NPZm
ru35rXGhs/sUjQYF4ncJP0UI7lgQBVh7cjwUEekKfWN4gjabqWL4JX73cm9W
QjxKB40mZK2VjhdoPOsQKNe8kSjVkKds+VldUM9acBTQ7PHco7qOgfmpZAHn
jjIKZVLF944D2vFAI4BE5LA5pICiYs1DptTO/6GoImp9fJeMISrSIo+otHNo
p9OamoTMAWif/iWQPk1q1KfXxEk6nMRdwTLbcHrCl6UG4PthL2S+rCF5LjAl
lgJM2HktLy6zph5mg06L7JUKgr0+86MbBDZooCNZWpD//hQT9UYXXHsPq69P
6mWEXsx9fT3Cus6ZDiQkQMyn7zC8MGheBG2J4xEXYzn8SjRNpeD1T+g5n17c
VoXGmiwbI5eYVrLi013MqhPKi2jXdwpVcFZxu2BswfFYWXVjqOyx0P8L57rf
TP5mtpk2KR5yPF3tcNHvyGbh1rODVSHTx/gWHe0JcvqHQ2Co78kC7WMbpu3z
W8A0sugr4lYQWxS/zXL8hUTIR0zEFARK+tGhwOc4pFU5XCWh1q04GsMbMR7R
WLki0Ino5ZWHQZIBwKsOnyUYDDl+Kk5wXNOum1r2ni8NNZNyV5Tpyxwbt5rn
2Zs6tgP6UaN0MG0S8H0QMDyIUIwWhiqsIx3VSvdcbiDGajOEiPUKhxubJwoo
DDFhOyTuLjBzIL40UcFQGDgEtky0eJUOVmlDY08164fjtxQyhvYQ8G12ycjI
CTBVfCOWVyy04KZfEB+Atd4U0auXLZFV8QHWrFH7i2/Hrw7/vQ09F3ntVerj
kSYbbW+j5SCdFq6zX8wT3HGKDcRr8QmvenzUJ0qn2y5ZWO8EDUZhSPMO5pDF
Zbi7uhuA/8CGRqk0VQc8sxkRaRnI2W6Jp8k0TGK54zgldI5G0cOBIpUZcx1O
gbhGymLFGLMNtygxPiBFMNVZkfnn+AXO7blXFaLKmGwvzqqtRrU3pM15qSDH
3POP+sI+vFlPLSRItsZF4hMSaPdE0HarPlyXwef8CVoOI5NhrIy/vKZIaKC8
HBOo9Igo4ptOTI1OliDb9pZpHKYu5CDEe0dTXpDaRTZLqpgf3bhjRgZ1Uhxt
upbUGkSYMGyvmfGiy55plO04yNOEzi9ml7SCEDvWubYSIug4LQwXRZY2BOgy
hlhWqEkCKbo/W3Sh8JgA1yiQ+MpNhDvziIaZmby0BlyHzYtZmZmklr4RfZYG
yrEnH6wHKkB3/xtQDt9sdGSC4A4sFL16RBmgpogZuZMZ4OyTQPtrBxiYTk3E
mdBbZQvT+TWqzVJq6szIBs3MZlunoGsTdggw//ruuuzqQJXaIu9/Y3taWQnE
ncVY7HOXbwi416QfxZjmJb+DMLww9f8wNq6r5ldheSU173SoNeiRaSmVEAQ8
3DRofqOCCAUZCUBi41TAu/N7t0LqVsX5T5wNSx+naKoOv33/1fL06SGjDaSN
pymwvUVASqUCB3sVib6pdYKfGF26y4fJApPpMBaaMkhHQ0F87N/OmUON2HJn
xg0LY3TCpUgY73IcX1OtEhv954VM1Y4pGi5af4gFP3LLHfzqk8ij8knGLCQT
oOpoVzNk+2a/NBEworXv5yq2l5OqYj7GzcpEIGCOAiZ0uH0th882mnM4fa46
9dSO4XumMm+gmzbmevO0hio+gyrl8bygYXHtoznpuftvQsCZpRBY7f1XIRdR
WjiVjrAj6t50gqDCwu11RdETHPnD8UjsqE04HUQKP6EjBHqNJrCJhjIlqsS0
+g1D51P20fppcsQThm9rtcjVtwfLjWK6CeK3qV9uD6fr65qDIxJEOYRRCnLY
cAd6pgJi2gbvKhjeSEb4BQ6ESpD5LlAjfXjJIBh2O3Xqf3ba8Ia+1e2VPzIK
7RhtMVC89VppY57Kb9TirYa4FnB2FjlZ43FrYYsF3gy9mhcI0EceJHh1F0eJ
xfgAQVJdVd+s2OvZ01OqoGuY3KHnsoQI2Lyzl5iS1qSlB2QpzdF9e/MQVFjA
ZY8N/u8jqIO2pdhPpZrrQX0ExKa9Rh1ZSDh4PeCJB8RMrTktFLEOeGX1IFNs
jf/aqopVp8ozHk2nMgcXyY7gGiWtdh9HqEHrGRJ8mruV0N+/+JgEjvW7qFOH
Yd5x8qzWMPPHwvCU7okOvXl+IFMZKdePCbjvU1XpgjXF2Rgrc8YQFPb65JK3
MTxL4aZzNWDx4miS2TMzLkdv6t8uTl1SLoqyCbjKrzFwWTQ1+/EU4wevL96P
MjP2Cv0+WPDwFQYpbhzZDs6/gFpcv/7+YWmd207ZiCrrCZA3qOl2eQpTAsvL
qtI24+iu8VTx6WMPmUqWwTRjRyZSWa0/B2P/RSZ4/iXuMVJ/t2Dw1iMel6wS
EqV93y27DdRVxM8P021FEqyR/bvVVXgK/rfsD634zdYs7SCGn75pPnwPCT87
wEzwe/orLUQafQCg1gWG8esZY8D0pxSbT74llgIT6mUWayFCYA8i0jTTpKPU
ieJ1MAz+JND9B9z1nQlNg3/8KtAYyRWpY8S/CAWiobRAiaPOeoMZgUwGh6kt
54xl2QXucBQlV4PUfYcTju6G8s0BBcv4SYtXvYnSmqaTqoKKPk927MgPDGQQ
aNyrWYR056ReBKYwqyJQKR00PHomNN2p00wYyfpawa5QCtytvkG3rt/HoLvt
r5oEWxAjRg00ivp3iRviXn3TFIJIiBOwE2zlLDI1CpGULZ3N6Ma3UzFUK+m+
wSUQJSzvFmD4afsQfXUpgiTPTKasTSKZVzlEL+X0nYVbO/qLkZOEEXIWAVkn
c6HfkAEumR6oxZcjNlHCCZzLR8J7F0cOfjgquVteUIPnYyZCMszLPaTo9sJ7
IEcBpzUVwDObe5UHSM2PyY7tTSwuKNYhLJj52u7WcXfH28Uwhhea+KcbHnUF
iLoNVNeK9M7aUuD3do1nLrHiEItIDkKhNF18V5UdKj/snacbKpXRBIiXoWv0
/g7pnym1GRfWC8KuGZGoLZ0bmo1JAkhwVhtveR635y4HIlyI3M5NR6dg8QPM
gpzabBBSfx/W8mikrthkz7LHyqhy2c+veBwL87JjYdeifRFjwz3ClszjJDOK
BSToRMBm4d8zX5uFzUSbeuNf183+jbCxvwNFaGLAzkvG6zd2wK7OkWYfCc/h
KJ2fpJ4ahupZpEEIyL44dXtBebFy2KZ080l8yAEj+kyMhWW1k5FIZC7S8gBF
XM/BErvxMwtFt0sZN3RsvbhOuJHWhChsoNVA8aTlcDKNCqUjuPkiF4yKMiPy
1hm8fqWKGjzPuLFaVE8sdiKqkq3FLeEXn9aDAqiu0jI3mhxqXVxVYPB5ngQT
HPFyT/iqlk99n4wPWYma4cstPTxND0Wm/1rYfZAR0vsqpoZn37lJixrAoBFo
az6vtByfGYrx2BVskdWJXKi4a1qrWJlFgFz+2tId9qhRdGXkJgKjfoBgCgOY
UdSJs30mKZjaj7Q1wkTQQeGuYEADoSJN/QpKKWtMy+e1C6/JsjaMr1v6hYWP
Rkje9mkSUDRTv5yI+tlzqKr5lGHDj75h3/o2+ssKq52s6Oas+HFZS+c629wx
coXgcz+m+fbt1LEc0OIk7CZXC+MfZr9iIFWbAVUTYIv5ZEPt8Po+RyVmweCK
6B6Clk5xzAK3u4Lg8Q57TJm84EDE7hOuFpOK9l6EYPPFgf/CugXVA9FXdszQ
DyfNjgT66Nelsii0/P409VpSciKvHRVjES0Fq8J9FuN1WUmW5ijUhgtKU1pZ
HzUQEDD4kpB2zU0oLAAGW1xrebPiqX34/4gsT3UYsQqtyfIvDxCw/jVmjNhM
pgmpJ0F3nCZX6rcNaa3Tne8EH5gxCJMQheq8AQWwAKzl4FeZpR9Vqh63G2wp
IrKMP/a9UaiODFUcFH43lC7g1Tn3vUm8J0U7wj68cmhVX+THK3w1YWvqCSLh
sDyRKG2i4r9zIv3wRo+Uv2Q8qF/d7HqmlazF6803DzNIYlVQBzDcByOVaajG
cJDg4eVqn8B+mtt8gb8sIfMFGLoANaQy1EQqi+rug6EQExe+0eFCEbCiSfwv
Bo5ztTekg4P69loZdNGz9vHjAiZv94RjLBC2ssJ5TScpgvfKp0GQ7U/c87Ys
yIh06KZtDs2oPJsT0pbJZ2gmFDiPLxNQsGQ25HBjtRj1FLT1QeYiB/9bXgpI
unUUpv6h6cZZzAMW2UfPxWHQ36cTh8ShYhynlICJHBM8L+H+hy2ZIL37APwa
eXazgIvuULZYmYdAHv/BytXhy0LeSHeyBVoSOilhUXD0dTCaLVyZ7D3QBHX9
DB4P18m7w54sUrwTytMPY/m7dWL6P0kiFxGz1IcWpbxaiOjhdNTzIn0o03ya
K37LP3WXkvpgpozOp5EWr0APZlrmgl9NiLSVs71p6YB5QJZgA/ajpE/v+HwJ
HhguKxfKJGxxYCifaSvqIjcYupBtyvvfMfUI/WqTBQSirst0W76iF4rmyhtT
dEydBsIRLbBD9GAO/pPSp6lInmc/OTvEZm5iuHJvS1QkAFuhHJlXGsbvW+L8
qyFyJRJmsupl+nfxyZfNi409GveTyvqMPQqSv8/6AcLroUaVuD+HEqqSvfVm
P5cGvzoclWoD9KCkcJG2kwvhhPSf0Kwfuph8rlP68ZHziFy2+hTjIn54Bffh
R9zEteJMO8tFfqC/WbkzbnMJs7jciB3+fimcHQLIUmdFsN5S0lLSeWLBuQkR
+aU/gIzrn2bSeTEVvtnzgXvujI/C+g+tGTzhDThidK7Jaj/MIfMRAIsjAmxf
VnDAuBYdFbf8/rMKHVCihrIgrYVST+vAu12bVivcNsbN4NlTJnw9Wus67lIs
XSE88acSp9GT+PjPVwYPfQwsSPr2tCTS5YJtxle6FlifaNuEAzT8pQ0LxX8z
2tX7USfojosjNsztlMf+n4qWULg6bAKQsrIsA9p7tVoB1B0F/kX/gGF7g/Vz
VvdPZcKj7hMCIi/pLPRjRnrUuB8UwANRL8RhNOGe5znHvQhrHzDO68CQKHPX
uh3E1nnvHOd6Zc3uqhah0HYnLNpitso81FJ8wf6FF8aebMAKc61yvY+8Qu9U
c3/0AwWM5wZVWhKv4dUKrNE8LYamw4LX1lhqeDtLTl4X9QYQpzUcMhVuM8la
Kj0HKvh7A1CgA+IIkhsjWUkCyhb5oJRPvQ5TAYrWuMG0wzo2DnI54w5DabdV
ufv4PkC9nxudRqUBRXZ2yOkVXR9F4el3E7qEQN33sz889sw6xkvCB+rnJnIb
DSMQhvDk7iWiAdQva51BlhNTvqZneWAyraxApWcT+qcUO8EkRDnyZodh/YNx
KPFxNOil1hsCkF5RHYokmPIbIWEpvOOaKj+GaCvx0K9i87Ys+j+m6MXHwd/I
QzSu+pQ/2nJymBektQktTscCCgsVGIG6hXG7tKCLqyg6aI5++a3YM8NluT0l
zEvYUOMK41FsnexR7mmqdKq1a/L/5snvFy8TRZaEZX29V7BJevP9ImX+E/zg
IQlsllyc/N4EfV6AuJDvgZMICRzV2FLP5IT9QfvUOzl/r8Xhx/3VID69V+X7
sjSdZbqH7AvA2hM9Ve78LDCfHV63s1fJyruZWd4xgw+bX2jzHtMON3Fp0iff
OkXXpiBZ6VefWDupH3R6COhOkil9mPmGlDUPgqKW0N4BkWMOiAL68k7EWiw3
GUpWWK0ltXxIbYmrkauc/UJHclDF2TQGCrldM3i6hz7Rg4FBCT4bLwsMvviT
bBtHcnjrUj3mz/q3AufOMMBi5i6dTrz6osZ/xt6fYyft92TetMH6zd5ipzUR
ZP5G6U1PkVAE3GxIkio7QYtmBA1tHH4J84Hz9YzGTBFQ6ePw6xgkFj91M0mD
opwyPFftFovq7tL7db6u4mTy9qF8v3OB1CUWhcWnm0ao8EONAsFaLtXTk1Xp
UWbUodTm9XgYI8Toe0rrUlCRLiV96lRX2EBKtYuQMb22mahwMkulgKZzFwMq
ofWlyVBJji2or0qBJbmthjDFxhhpzuE7p/IgrfwhkrtGC4Waz/fBp066VAY1
Ws8C2u75A/+3+B1BwIIR1aR6DHN9S0tBtUnMQfQ+VkqYKKrGSzPjuiS9EkIg
qs11fF/EpHahBPlbSvL2WSjyzMUR1ZnBBb2UwR70oNOM1Z5AJCmaPJHddcE6
nSjXP2o7Dy5iII196mkiopfeesaV5ZLcdUPluSYAQURZJV2EJf9fgFi6jwts
USwwhXMeNgkHyr73d1z9BlyG4y8973WXQfzZu2QFTL3Mu+F8v/iEXWlj0Mkv
COlJui+sksa2p+zGD0S/oFBajRJU2ZptRKW7las1yrKCtrLxtYt0MAYkrmnR
YG9h+NP/UpjM7yF2+e2apVUcO/95MdcgZZeQhB5C8NfwcjMz+a+mz8WqBwh7
SQjLCSbd+/jRjyBWUM6RddQL+wKqXEG282TGwwhweMCk5x2FjOjbzBP30qw/
Wre9RUh1xlUFv9uSIfz9D3mX7Skbjj6PYftqtuCQz+atVgytFw45gTVffhbr
jflImlD4GPO88H/5EJjOig/S0pNWpFR05iEqU+P0CJr04i4KdK7iqH2kzXyP
QIQbcmxuo83FuO2gDSoiXGEFlR4j5n8W6A/zRa8XFyCFwKjxffc5h6bLy7ZL
DoA2P3I9Y7/NOaPIBsPsEDeZ43Ba1U19UjzpUkIOjCbLVjbgUaXkTS8Ctsb6
bG6tmmrxJ8DEsxq+VLBrRSjGKts5HTk8kzTgWfzS4CLYTSItfprBvLcaC2b5
5YkPkczKo4iVSSuaM2H2NaHJlv7VUWrWnVcwtBvkDjrMgpRHTCez3l3kLBMN
zaNYLlmjCxmfC5IHWGjU+eZUU5+LhZ22SHFlDkWO9e/9Ghe0rs+ztxB5rwx3
sgFZ7RI2kH9d+1tGndSaPlQwmocefdf3CRH8UrIJuD+7O3KK4x2wNtwvzDva
La0LrNvIVlMWHSvaU2gVJ6cWKs1jRasxyKcixePt4jRMPSTzs6PfZBTFEiGO
kDXjBjMhsvFbixFILNwxk0DcqkG5o9urt1rUjnOOdpMRN43Vf3Sv/dRaaCXq
2RD94FAEHUx0eOzSUHSxOqC9Z/8aN1sX/jB8uGhO7TV8LA+paFtOZmc0hxcW
A77yPkwlHwZ4cn3TMNnfEHFKialmku5EM89tQTdHy3Dc0GvcTLCV/OmARqPY
jyFZq16JZ30bpJf8sAndLoLAbXpTg7vyJn/HdxlULmNBD9EXUXyE8cTpRF3J
tPx0iFmxaWrIz4r8sIQtyuyOiWmiLtSQd59T7Z2wcvwFEwvM69RlDZ3QhYEZ
drcqrQzvfi7WzVYho5FCYoCQr4n9gIgxbxzmuFVW5uY5uIgYZwcdknrTgS+B
u2QEGunCidqy1xbTXo92KalnZVzSzRtBTve2woX/2KQ2bedhAwmZi6hrDT9I
hZkq/E3dfcC5tfFG9u/EvOw/Qn0oqioxHUHQLcRFF306r//0qxMOTunD6xt2
MtvtykVrs+15xGJNcI6LtEOZMuVPuXUyVmjCURHzIAZzEg+KJ+0dR4Q4LeWg
KyGQniS4ES2TbITl0jNioB0Pyv2WuqRdxQNoK9VYhiuxiLg8ItN/FO0OSFHL
158FBBD1exWaHiNqqVbiE2j7Xyb3yow6B5ZyL+gY/pS8RoR1dHuuvfQ5nTxi
sRc2T1RBJXpXhVjd5J/Gj5FLhiagWNjRUAbgs79Gn/3tahoHeNdRPClorNJX
o7RKelk3+JetmLhyMKv5EBbBHCtDEud8sceg2vqcM72TWBsSUkp59qJTbZ70
bCSpNfFRgbTEf3mBGNk9AuYqvImEIbrbeEctk6CdJnPXVQy0BiYeQw7bFspI
iHu39ayzsCFUBmrOZHAPzbth4B/CehJpFBpzoKrUs8Bfm6roOUjABpVc6hXu
TzmIiiBpFFzsl2YYLo2UxHZ3MIWCDlW19oWOAyxlhvY635LA+UK22d4UqQnU
HJVYeZGKhoBvecBzFyncvI1um6zHC+FrD1kxTW0Snk6l1Z3Vvue2Vi4CtMkr
E4TZ3LxEmfe04NbcHlcRkTqULPkT3y/XTdKVZrTtR4k2TMZ1WQ2A591k4Uh4
ZlHd/QqLVDbZmQRFCPX6QrkEbi8IH0nEsIEYmH7W8y+Hz2U9MYerTAUkkhZ3
3z9EcRuGAXN0qQO7LaeX8Eo7PYu9WDJOX7eqFt+Af7wNz0D4jLhnd+Xve1NO
/ww0p9Btgl7vHOLYwa5lYnUtbGCmCET9c/agi5H6S7TRhbDLVlNvA5oHQ++Q
rRUAoz4JcY4abmIolLVDsnwCyfLnV0Fny6FHvwyruZJonDpXqOPRyqXAeg6L
obNuzPg46zDcP/O1LyiyGsMlSrNUhPKAT/VUgBsUOh0muHYtoswdo+pEBSes
+2LbPSb3tIP0tDW63iydwd4spTiQLAIRqeQ/1EFNx/DDKrNT9eJZseUdFlpg
SAPFJwiW0oRiDFPuvxEJkjGpdu/+Tdq+QL45O303/+NxzoR0ARJ2Kt+HOMp0
uT3D/wwO+NMO0DQI5sZfyV319UUhGnqddWiNFag8YEwPmX69jbCgoNTJZVH+
ibxk7HHVeUmh+Db4xoQr/2s4OhEDSUj75vm0p1pKHn1A1KnlD6JDTVhia5WN
VXzw4UYe9XoUYTYYVEjyjguV7e5ebVJ/CograYklo/LUamgHZzi8CNp6EOBx
7Yi8IcpvK80JC2GEKj9fJwiS8FkeSuU2TQUpWFzbkiXKQsD2KlwMdrPwGvPC
fSd9HtbTRs1tTBLLjeGvtfT3DBWZOGV/E1PAFyxhzwRfdlcSizA1odnzIg6n
iET6NHd3xxkFVmcr6s/NeOe4uC8oaSa18qXKf5WTawAzzGTljkxDEkcXA9yG
kHn6/iDOGsR5Ww8APDfmmdTMYRrg8UEj1FJ+fSt6prDBmIh9HykHTRrYT3l6
1GBCuLQGUiWySNr7qX8HZzZb7TtcCcDfuGQL2NDgz3z0rG/ZjNAARcZYHrDQ
dpX7pZhAyuk5HrFrcPYDNZUmx2HZokYyUtTwz/3iLmzbYpXaHo/Pbqvj2WdE
UIdA2AZZ4EE0W6qFRY7xiqw105HIrp0kzcdH0ETWXtww5msD1gCuvJ9AKB+4
IU70JYbsEudUs9aLwwYJeNghZHY+PV3qOeCgWNc1+VhHb113PJeFBhM4H7/Q
e2cIMliJwMuyshxREUC8953awdautiFI3BOd31CMEkIBdG5Obop2HIVKjTXe
ZKPR6RmvZhNlHyDmE8zgt8gdiw/t+OnM1pF+h1VzBM0Wt1c+Vf5src5NZyeY
bmrJH+FIIV4LTXntt4W5isvGfu/lad7WvXAuaQ54HR5cyAOgoczm+vWLdUw3
C2n0ja/vfz4LrZLsJMiC03vgWe/R7cHT3LavhOxKdNr/KCX5TiafPNSuUcMi
pLf7fQ+p0My7nkipVyO2/Jxf9mJtjvDp9KYFGV50J8+0DNamw31qcc5Rwhtc
b2XslHTpov9A/9S0o9e0gzd3elooqOC/YFPvO5Eroct1bdE6eNgqpFqS45fh
Hms/huLldxjnDlciY4Cyd8YZN9FkJNZCmj2SVbtSsBPjxs8g9u7fgV07CZBs
GHbRU2Bkzb969LheNqBlKTjojAbihhIe+mGWXR97i2eydxgDukdNEAhvvMEl
1ilfNEKfDLJtVe018FP3mlhPYf4C26VWgSe5+aoeOPAA7pcK+xU5sygvAgWI
kTpnXr3etAPyEuVlNRyHh58KcjXVm8axYJFDg3FwL3Q+PzihnwaHbgwu+wOa
XOMGVNYmt4BH6ix5SAxoN33IYpRbE+ND5WQHouJip8yDIwLx/tH/EHcLY/m+
lrlehnP1BxCKHqmBlFaof+D2PhaytlkWFEy8ORV6N+r/6+LwC+HiIfCpsEj5
LW6wROGsyA/4DtlrMgvhtPxbTc61XlZcgWtRBCm8p7GDVurjEDIbOOln13OT
+nFg2zLrF2QqyhUGVM56pUonBFy17bvL6MtatQOUrvdXX6GuXj8tE7ya30zU
Tg96HjUP4BADRTbWHpm9ycgcN+eboS6xR6Zz8PqdRXmjOBaT3P2w4SGtPz2E
zg/wv4prd0/yy5GX0dA3IUntALtuDTeXOJzwnH4QitGvG+ZY7FAObGY+eHkm
/g4ODZI/07FmykTJ2txqcp2ekNgN3UYlY3SZZr9LQGwcd+u+RMHjI0fgYkMj
DTJRdn03KLKTfCbg3S5wWzTT+BosTVk7j4F2Nl65h1pxj97dn8010StUvbvS
ZiQH7Fz2SKNfTkRZFFikIJl5w3VEUrIu5bupJ2iUtuI5dsMN7usMY1J1ASJl
sFA4rXy9iueJeo/31zsJud0TEZzNfXC/4Py9ihMb8jvjdfzx8HeRHKNpUpHK
PD1faMyjZ7UN76cwEAqeba4trha2S+820+GN9lnmn7OGa+HnVPwDSQpMSDnu
UKkkeTmm/ijAsGsMW9evdItvL1Ub9IH2zM1zl5nNIK6R7idkqKfrc7RxHN8d
Hc0e4ul3gt2rCVr486JVIQzaEXftunIHYocAL6uctxJnZK25rJpOwsy83AxD
j+NX9SxvAV0HQaPAa6uGoeTLmTseGcQsLEI0t+VabkSneNd2qm2XCjD0onPZ
YyJMRTWHGPoUSQWiIrP8og8veta41l+H8k7bdNIltGyWQJxxYqBnZSgnP4M8
etpLfx3i2eF9XYAsi4IALlj1CaeJHO3DGjqNtdD2frI4SyvKPBV7MLsuJE8C
R0R82CnUmyATg74QobTUzLUVLDthXXobN6BF17WzAR8HSuGMEhr7iMop5U0/
gknc70k+vSLA9GGMEN8YCJ1sVKR5yOCpWxo+cBz/6bp4DXR2kCKQUGzfK7az
vMttwRBzW+Z7AaBz8lQqQfuE3kDmRUVgnb+X30Ve6ie2HYnymbRCYD9j6/Ik
kA/l5VRKSPXcf464mSA2C9icc4E/glMpM93vPHCPTkt/qbsP+VpqLsGnbL3e
cAv2elEsxeik/DqXWzlhGZJRWhdC9oBfIkB6A5PxnYe6WXb0XHtcGsEpptfM
sh/PSd+62ki0PCIvP8ZZpG0T5/RHWk6qjnEEIg7z5cqZrv5jR8C8ApP8xAjO
IsZaC42kWrakzX51YtA3hp0gVaNN8fSjpPKXj3p6O+Yc0Fv6RK0ftXJiIq0o
EHEfas1UaIbvK4ZNFoBoz8/JUHZWL2yVwegTZPbQZ6q9yW4dJ79tZKI8RbvO
Zcu+TN7KkcvV5jKNOQ83zwT3bVCMCUr5KShb7QFEnglaVQenZkoNNKzSrS4N
l8mgDELRtch1NOe5cr7pzZhQjwXN3OIz73gI8X//H2U73L2znghDhyf5YSYH
JUru1g3OnIuh6kPRkIZlCWdicdClCzDNKJYJEjyjLiDDAQciA7hhpvNfEspU
OU09dqsrXXMd2TvKdF/3w7xa0sMOeJg4MShZhZ9bBWdBb7WUghO6sfNSAF/P
gl0K2OTBZDa3ArcdxL/81l/a2iy34THhf6Tn8My293cnf0RnEBNrQBQmBCFK
g6j3ESGIrmT8MqTfKEiKB7Cj9/OGaiM7iEakX9gS4JEJvpNYfgS1GeGk8rhI
xU41DmZkDLI/6izW9IhiITwLIplRX/Ra680CxgOmhDKofwugzimRHRB2IhCF
hOu5yl5tJR9SbnInlDeddEzLAVMO5YWjiXrJpIKIApz0aogj54ugh4nKH+bV
YVWgqRjwHGwHPtTInEqDsg/7dNN01ScXfmvhe7NmtGSpShHGHQYjQf3CPy/S
TDmHXVN1exBXnlP2XoUurVak3YTTfGUuJYFH3I8+rMtxQuYZ4LoTx9wkySQ0
mlc+tBSuVtIqhLNQCu342WHjxP8DcvTjz9uWEdvZos7aIsNzhzlBJKNP5JjN
f5FTn665DY18eo4anopQIcvE0GZDrDPQwoP/EcU87iyNonlDqT1FTFFCf/fr
OpKVIq+rFrYNhNND7W7yUAOL/YlnOJ/xxfHsHigbdzA8XCVVPs+RWtvOAoLA
nyM8r9MB+K7O8Slodth+F/rFq6SX35wpBK8iqx6Yw/CaQL7JNDHhp8rlXyV4
I7APppCCeBNh9zThvCIlS9XGIG/ma8QPYagwj7AG3i9zdi9Xo8GlwFfglv16
tRG4tNEL2T8StQw21f/GdlAxI/PUdNbmcWyYkusNp0eOWaDd6x8zm/K/+9TP
cL8tclQq/V+E+W6pnaqxT5Qk5cD1YG5BU5Z5TMthqYQ952tzV81iisv+IfHc
OHyVYS2zWljt5YeqcG2Fe5I1e8CQ4K6S3Bi8/9NAqY0f9N7Aai4KaIb4c5H0
8y5Vt7EgbTBY7zzbQ7BDF5VbKwZZ6Vrtdyk2DaeDfCOXzGc4l+Kkb7fUFH3Z
H4ePtcbCQwzep4JULPZjhtc7SdczSDapatLUtlJ/9G4v8mCoI41w9Kc+ntz0
FPs0+Gu1aADnLIFq7AzZMybXHksV5NkU+wKmoP7A2kuhc8dLBZ3WAcZm6gbX
QppUG1/I0Sf6sldS0MCRDwvaPQKcB8PwyrnclMmLwJs5Uoe2pqlerD67S9a3
78e8xi3JuDLHjvS0i150WeySoLfl/aq1Xcykmwl9qYqbSTuBBm1hFfpDH+Gf
ZabhvgWaFnAHL8fo5ya4qcI7o0wfZXDxRHBaIKI+SRt78Aoyj6LgGPvnsO5o
WT1R8imi64DbnADoGh5PoP8GMvsTJyxr3ZVvwDNu5pLP384atx4f5WemoXhS
nJVq5eKfev0DpP/jLfaLEwQNnyU7qRS7T4BhW6BVOHAW4P6aeyzVuaNbf9fw
hEw7RW8esTnMYH8xJdC3BWJgcHgSSWzJjswukQFsnwNNIfuv/1+lFFl7ImnT
fnfV5PzlDgXlAHrG8uandMX29UB0MHf+nNR+MKmtAA6Cia35Hljbh0plbfEt
rvqVNSWQ9jvkEw7r9nY6D2NaZ5K3yxCftQMj5EG8aj3s5JJtDID4aTq8xFc+
sOKi22ieTJ7beSSpO844LFshBlY55GZoPKrfbuLpLXYIyUwnOPq75Ack6hjC
tFJ+YYPmiptUmF7LuDjvQ0Zx3j2h5wxde7G1ibTivRo15Lq8+tZFZzT74zgI
MhJbftEZudlYZmpnlo60qNVFrEoBEvsvZ28UQ36CEPFwx0B9j6RdoPOklhVt
Gqa9gvNiD6pIHlizzCkd5793vuhAH8Wb2lrrAFuaDU6g69EFyaHXxv+31mf3
X0OIj51N3QH/5yIyIE35jW3s8h2tfZtWi1aGqS1kNihW4XntW/lMboB1R8/o
4QCfCYOPCmOGRmOC4pkiaUkjFO3Pi8D5XYG+gTSmmz5W1sI8g6Cus0kDhguQ
1jyR1CtPypbKQ2dSCm6AVm2RQ83/fM6qtgm8NRQqftlrPqpm0DwgZr39XG9d
otrP0BmNhIAP/G03cN5l038fZ/5GYe4VK6B2FrZi9gXTo38xsFZgBSAo71Vg
5phSZgXFF4WQFC5EC2W7OWUv7dxZUHldBWDr+SS2WBDUhWeLJPYvgL6SW0GW
TsMAsm+HKSEboAc/de0tkc9urTv1Hs1CnHcUqLkOV7Iw0IxMkBaxcEMYhETt
+jFLqLIWUPxg2Q5lkwlcqK5c5RLDywCI8XGRcPH1iz7cfJBSgo4AoATQfCiD
VGqpcV2DHGXwTJk/BKizCnrqWxM2POM937g6RGC94J7nzSykfbvjvTAL18vo
oOZsxlm9wOCPmOsri2BO19F8TyNLIQ7xeXc5nb7EBrnsP6tzaMop7Kd4vDis
mNgLDem+OvPVmKpdx99iVHWzgkCWWYhr0MQ4WjM4nUBwhjvKbEeizeu36u/Q
1gKr7FCbqdBRieCum7nzc+E+aRtE2H3EMeAYGSLScpEeru3dqbdKq5m9tu4+
dDrPp6YYh8wKWonfXmoTDMQGnWeD3notN0glD1q9bA18MjBpJJuPGZ9cZWnM
IzWlyNYmxDQlepNC2Rex0z5WVfbppHj4VTzewsr6oeg+rfJahoN0M9pzH4e+
I+man1A86LESg1DNKuaExAYW1maYHoCjkudteZSmcDZ9xMnvBUpyN7Vh6rq4
MFZFd5ggpi9srxNpa1rtq1rwYXUVMW+d3Jgm10wV9W+aQQdjYkIcDrjaTimz
0u/R3fBul5XfydOyPpuoIOUBf7j2oxkJ+f1J3z4n/jbs3F8D+CIInuSAS1bP
7hjd65b+xbgQwEJoOSN1x/dy1QROYHZ8uHjsk9UVSdgElMaP3c6SFpf9O/U9
1bEP0oYkhe+fPSfyHfktLmHu2cBTMpu1mmUKDOh0tNggi4/geDhg6wISIGar
3M5ul2yZA3AGMKga2pQDyi8xXCi/eYVO9Q7y98KA82+80SKX6iGtfhfPRtAq
0VZaAqas66y40O/VKr7qWKa1wIk+sCP9wJQOHEHU217PZO9pMRSHBd+zFCeW
DOLRd8j1IpOl9oY58nKe+riO7C5JlQwzziVgg2C3cUFBC1MbE71hhOC20yT3
LnhTbhj1IRH5yQPP5DCIG4ToxdojcuU+civutfGGj9sMwwZK/S0aJw9xfna2
15zaGC4G3JJKyIft4dXdxxK0jphlAgsCzyKB3WgsDBV7OSgZW/j6EJSIrnQJ
h8ZuaXZ+Z6fRrTwfZbvkCsiHURZsMKhYdEWjco0hX8h8m1lAgSHcTCCz6rBn
6mKw1tsAfAdH1w0FFdswLdXPYnM5eMEj9uliprEV4t0fvzIdHg2AO6Nne4I3
DI0H5/X5sDa0XLi+0YKwvtg25JUqoxY7MY6+pQUZ5SImX8HnnirDldVptiMc
wZGlWq/+U0gNVHFloMnrCSGJOBZClK9HVMa/PYHlNfj6MYXpGe5ONJxg8gQm
KmcewDS3NjxyV31MPT1PbPUH8ycDSELHc9GE5tDAO73IwI+zGuJhztkteMaM
lJSaGcxAZF7hjX1yUyZEx8IGcCT2B4QhVY8G/PF04Ldu8VYlgo0CRNPaCrDa
/ppeNiHpgfMi6R/jj1xqL1Bg1wwSM3QW2UiPsVjBPb2stdkg53byZ5f1QpfN
pCsr9LoqK71CleRIOXVe/F68FPt/BUE9CAJe7XcFYrqAId3g8ZJ7ZvysEIpV
h3Ja5oZczy0+Nt0Q/egU05bks/wVDVm1bU8qnAb1dMX23dd28lWz2f8Hjbji
GBi17c+227LH2Fqs9wfHJ5nmw3MPzPVr/juzFsyicPXtk961XaqAn0OYoxcy
5eL7r7AyfjcEgK5CNtM/j8B4zQ+ZE1o/HrQySTaHVo8v+n6cFnCjF9ccCHiF
WHFgmmt30hXOZGw4yOe0WR7BTNA9j/rzAU8uY0fghTI30UxVfjKsX3Y7qRa9
os+diqF6+ijW6Ovpj4mW/ZgVlPTZTyknajUmUatTcFQTQMUclq0oQsG5NyVA
kpsxooWSlmKa+rEWZJL5rnTPDjXQXHoCJMob11c9ySzDHbOHMEQ0rYvvEpLi
oo1aNyCdzC/ypsilkQ+OemBBInXT+ixOuBoDDlIeyU9CPGHnC8rL/osL6S8a
7a1b78/vxYLeBtEhIDWI13AvZFRvyX9UXsZX2ur3p22wPJhUu/EUvjKNcacv
Cp191K4WNnKPd+p+Tt5EpnmS+d2A/G8CGmTskbcO/ythWgdIVTJYROMnRtZw
OBLJu8WKEMrlZCEwT7ehY7YDEtwRk04yjIq39MhW1ThA0VQX5L9aa4C8ei/z
H5x4xzR5P0noT05CzERAwIz4cMZoLAT+SnRipfojVQRNi/okYQ8cCKjyMnmd
SBPpUj5BS3mq5T8rMXBP3Is5LNbnoYXsXBGd00fkLfqA5pLVDvaK9tANBMUq
gBdWKtYpGaejfxZQd8Ywklzxpr8oppqTjurVEGxL6hDPC5mVA/YLJ+dyQpux
iZw83FhAeNqqp9OPHRXY4OiYHlt+pYsJw7iW8HzoCD7LjY7iXg7IdjCMg6kH
peWOO9jrNFvmHrOS5RYNPmGoDLYKKqBegRHQ4UFyY34aJAHX3vbDMQJqE4PU
QLPfK9STDO0RRkS7lr9LCcxLfuPA4Q4w8khEkJyHO6PXH/1XfUHWauPyOuWH
OCHk/5nlSidr5zEKsL4Iy+aBgx9XlmLGiqJ5rKhxCwU6dOAQYcjyMgtyKrkN
DkLfSn+a193Wbad3lDy7P4yGq6yMz+jUR/+fMAe9BrOouREb8G2sC3X4w+fK
EZABH3p93kVyokxhSgzyHyg6jxx5zgwW6BJuSF0s1UGclc5ACOSdKoZ1pl3C
OsBQDrYUONzK5JYTvKaQFhkcJ3GmJtvIdirgN+OzvmaSVf/VMb4d7CkHly4S
YjYJ+ieO94nfrnIk3zNHgmseWbGTkxwWgER1RpM4OLU6OufhVDeUTBl55m2L
sJivOKyt7JpXN9omtoPSxSDwwpw+HbXUafUKgPHiBLcwjjzVNwjpJektOPLh
R1xNWYkj8l4k/BEV+tHiHrw/Pi5b5jdUkE0WkdX44ljApURMI7mAWjnrRylH
oL0sGqkdJ6LifdB2Gs6OVxQwsWqEakErzCE5tYeBdUVAJynz9+CuVDdNTFJN
91x35Sqmek577ChOZ+z09uBwKAQwPfKsnvuKl0YisVxi7xPLqIB+TG6kQkY7
v8pDMLSX/9H9bKsevTGENpFPDu8rrQ1Fz6yVLRtRGuSMkZ5/OoKsz4iFhvIw
GLUadgad7RGN68kqNs8NzXWDW1ualA9iB9wh1ckB2ydi2roon6KtyJRSMEVw
UP1XazxvG2Lpx0en485GQEtIzhUczp+8ebwecLHBa/4kKcJcqBUajFGbOma1
R27qkuusQfFfiB9sfma7ndjsLEXahS8DNd077lmNE4uKgD0X49MACTk3cPAX
5obUywugHuV6deSDFD2pouAnp8wxVms2NtI6K5EN1Q4LsfhLjmLOTjUhcZ0Y
p/w8hS0v6giDXhw3qAITvCAGDmhaIhi6uUEWAYg70GNBIzqvk/tTUKOaEc+r
+DS6sVjlX30/Z8Nn+MAgi1poLDy+S+awl+UVmMjJjkd+VvzGP83JuodoqO7U
Ub6ol8N5KyqA9eYTtr2HgrLWeDolXcCN/BvDDBJ4rdU9APulK/QfF95uKZND
RymtTwn6x4QRsRf4cI3fhJLTuceuI75G7KbX0hWD/WSfb+3fr5cLMZjJpKBW
XkG9lhAnMLnKgTcvaG8sBfombgBhYbYV6czXW4HiBn/leKfFpVZQgqygQAdt
RbBmx576dIJ1tb6enTuKj9AynMlzooe9vE0tmhlnU3u4c2MhfEZ+yzmG2Jmx
R+W7ZofZoQXuXGbYct9VB1sbwoTkeDfRVmtPSfEczxHK7oLxzgkWN2k6a1lG
whQFztYrLnR9AnkGIpk/34MjI30hA9ZEOLCSpahvJwwwGXGSJT/3x+jh+Zpj
wqNfrCO3M/PLQhXFTPFK+ilcXExub+00pyV5ywqT5Wgk+2VWlzJj+798TW1U
qOAZRKVJ42PTsNt9PFASnGBKmIReXKJdyNMkDqHnY+mW9T6BnBeh90z+N1NZ
sZdlLTrivh6H14qL0j/s4iNvNNSOWrn8yzpDIQqROawgCGn8NOHUjrnko9Bi
WCuNgJ27/PLMMPXJ0FOCIu75zKZgnbsz2NwC5akY7BQpNLvNjcjh+FPMgILs
iK7VJ90/8czNtiMSI+yKoX+esSvarr0dpmW5KQ9CtkcFWIJ0SagC6izZN2HI
kyUGVOnO+/1BWFZrZqwMpcLOG3CtM1dCOoRi1o21SzvGholAgdbhulN0XYYy
i6ox8WhK/kCd3a4/DqwcbKcgv4jlwtDEIix3/ITaOm3O/r+o/IThKaouTAcN
Szl2z7maerZNUjhzKHyeR9YUDaan3SFr4zczPPjxY9dMIGup3KOIp+OJVpcw
e1rAGpGbZR8jRY92tijTxew2xRxsJjk293mqtEDTd13tyOMYUx65v5lLbLzJ
R7zGILSuQolhTEReUQrlsPiRVJr4eu/fJPnkm/zowFTX4QktZGDX3htnCK5B
jkSM2CEZLkvENzK3HfdDktPRr9xC/FIVDXBCtNdugoUAz7JCs2xK9c9nkACO
c+9FHAFW5B1OSRLbVoUC/EhcWscRCAZbHvRnzJeOCxb5+/YwEGECW7MbH0us
xJ2K86W2TvK+raa7ScmlqyerNWpydfcxYBlxolED9730p2+D2SuDqpr82Cm1
/igqIvco0dOKOgPR5k6Te70UX2nCVjrWh1lYaIxCqmJdVKYGPQDLZlKEemPU
18oB0UDAKgf7/3X4U4JTlk7mKv/ewuOuOxNUg1E1+aFuRN/5WP0SgVV9sUY5
JpJDrfm1IoXwN1Ept8k49LUy6VADZcc1BqT85d1mqzH9boZpbhf7bXmLOE/I
XXcAV1VW3Lcyc22Bz3rDIrnLl1EwSaWuZQ2ClyruX2W87zT0aDV7kVRO0BkN
MMVuNINiSLEDNSwQ7RxJk1BVNk2buK3HBLj8W+TiQsC4bHt80YnSXKSnZ6zI
l9caieB6kOia5D7rPm113fy56F+UiKMzsVDGMZOxHLS9dIKyw+WP5nLYb/7p
HuKm4j0QrMp8LgI8HhW/Rf//N39meDQxD01mpKRMSrdNgk8Yg7YTDuqzq6rI
gjCvJ5NqgRDuh6AsrxNNHcpchzOZROu/b+k/JBie5dW7Lc+6LLmG1ydrSxvF
uj89HBz/d7dSU2l6+ju+l8r6lKu+6CbLNDH1kMOtU0BvFUN127BTE7s/pD+3
a8jmtLpkVdKbXTMJbFZI+7lmC5/KXSYNuqQ20IZ229nsRQrffnUDyMjh5ZtH
AzfKY1C3a0ecyYWDzJd/KugguJLrbSRcsIuLz5y+vP54JemD5jokHG7tKcZB
HIvcjRvA8uG7d9IDtEGPjPMpKUjXAnzKE9EpjO89Srqt2daG5V6VZfE6XNDf
hh0RNMG0qzwmaMSrpwIkqUaRlx58tBbBWVo6C8TOqE/ydHA5Wj7QCYToA+4Q
Icorcyl34fWNFWKLJKVWvuwOBzJlAfC8bVK8ecK+DufOeGuA8gFgOOAaShAM
m1nK+hXyn5Ey/6MPg6FmooMSP5HWFqHjBIoB+D49QIXeplF2IIKkl7CV2DAr
0KR6/kBylvARtyW+6fJSY1lbq0lHnNCsiX1jyazEg6kJ0CN6runLf9c1FvsX
wl+0hKNRAAyZvz6tdsCAiihrMN8FKUYl9P+tNBSzrnQ1ur4rBmLkpCLuyneK
VNsWUnpwGDs63qqmZRpGoXojxXH1ksPvY+ZRvSN+iJf6NyDLs7MsloIbY7wp
iazGcEKlWDb+VcnqJDX8R4BtxIWNxLD2b6z4okcEZaf55mU8s7gjX5znXw20
h9qNtK9pD/vhL9+ljCcKA9B3P19T80XlL/n4G7rCKdbth4DbpDlRXabWK8IH
79goNc8p+o+BUj0n16iwxWrl0Qf1hNTBCL1a3uve73a6g6t5en7IT3PhvTa0
QCKeTrzAMNTbQrW1co++OotHXeRlsstsUbTGE2EEXZj4ezS0P1PS7HIi0v3w
pIiAZULI7s9Es5LD1/h4jj6djoIFBJQrCIDxTX+wz06ht1JUWv7/B+D+yz3I
gZ+hpY0V0yqysPxxM7GBCz76WzSOTAn9q2MCI1XlEJAgYnWUVd03u+u8Berm
3DG2iEWie8D3cvyLe/0WTXr318U6Zv1QjEE125RZ+bFAtLifXqVeAhfVJ1Ik
Nigd4q/xSQLLGTQlYn9bqlyj/nBbUVFDpansbpUJdPSbA2TIV/A2zMGV2mmB
rweSq4DjRDqmlWyCUk8JjA9PD0UkycyUIa7COeNaL7HU1NGI5yw/vqGqHf0e
AM4OcQt92HTe1dWtWRvftBX108Rpufa6wtZknBjrS+uwuUj7iAWIUSxBm3XP
EcdmGepj2iV5hUVo4iSofUBPEGg4ql6KJaVzSLlP31yDhqAjyzWYV8iinYm0
U6ZhsmgJ4DoPcVxK/PmzAgj5+ru62GxyKSo3tPmQxfDg7jCIhGLG7n+DkO/u
5CZ01XEW0xfH/xUVSoazkQzz+WZ+RDqdwc298OsBPK2Q4v4Cz677H9o6Jg+9
swGVYd35tLr12sReqj69CCJicgCbFESJJZzx6nUQEOcfC3vHQttqdEpThiPq
RW/u9D36ImRXI3ykQcssiU3iGMKMGH4v3fnnFKkE+6u1YQ3yzK0QCzuvksKj
f+aK5tYc+6i0gLcqcGyVGKxVTkcWwJ2M5U7kk9xZ4Y4r3/2Cp2dvy+k032IC
ajSGxZqTULDVWHogs7q19BH+Cth7yQ1uLWrcBrQ+ui+Up8VYDliqFKmpoU4K
gryAsYBQfwBEetT5F6jJMeMIBlPX0r90RemPsExTg8nck3aKr8o/YPCSl6FA
4ZoEXpJtDhkBXyuQMSqobjQZujuj4WAntKk6uS96oGRiEIBlhXDaJCSvIcg/
RtURYZ+UBwISCSw4zXKHUmz2t5wVUVC6kDLxDc4UvXs7a2Z2qUUKNLCPq7vC
tz/lOhE4VVa6wNvIRkjBNIL0Dqce3XL52Ef7xy5ED2kCpx5LOUTJTMr/7B01
zZRX39NYrqmTZY/gCeBrEvNCd8+btM6ck+A2NJiJKqAuPI/ORP9/dp7FUrcH
22js7Y+0VKk6liSnXI9uZojaLeKHHbJF+PLyduClJApTqC/IV7J7sWdTf87m
8ftD2yHo/jErCrltNkobYASMMTqqb/lGZy+4bZs2aVBKLncd3aTOW0W+O85K
CABYjV8z4x9G2v8bHPr330nULUZ+dLwabbHnRunrE70ng7nkSkU8tG4L0RaJ
HJ/xXaZShb+l9DIuhSG1B4GhgXLydF+5Phclovcj90xD9Tdp2FpcNDw5eIz4
XyhvexTho813AcL2MJd9yH0ITApbsZG8J/mNY+BPYWSycJvIyPDaiVcNA1TA
HYoSa+3X/YbG+ehoGUhJRsAphxabwgXm4Y9SAdfqLpUTbfuiUg+X+mRLhRTP
lkjrj0SIi+etH9XC6aLXYjo/EhF3cuU69XKDsOWGWYGSbNUqheVa9sVjnU7Y
GvlvCKO2RLuhGOrVNhOdvXlimNMRiKQkHFMRX8VEyUvRnsedeP+sslnJNzWa
jDVYZhjpGHjoKHEpU11vgupxKDPUQCpAmMJejRO80lV4L6jutemaSaaLC9HF
LaVU/nLcIDgDXzKHej3ji5/iB6lL5kNwA6SCIuyVV4DCrBvV/Z/lIUmviz5y
ZLrTjjsb9DWXf8dXRqyDjZgaMjVFz7cQZizanP/kPCnBTMfHuYLwH3dgVwCu
NknCpHcI4lYhYhqzuV7ZYKM0gG7gg+a8RERdBayJ2l0MYSf73P9EalOEOC+6
WDT3MKpypc46Z3f+6RineSVaT0ihahp16DctQn9s9Ss8pLYdCuJEbRxyqMJi
hXje2z+7ZCqWy660dIqtPj8YsCba/Y9JUhSRlOfVfVrlR7NKPox6hjKQgc8N
zMWIUsxK0hn0hwWyQ3R4EELoU2rBczJ5u32Z6O/QFwaKO7TVHjg6rlJ92O9x
pSEzMPS9feNZOxeQXYRV+QJxWHewyNngNaIbWCQFlyhfhKVeLTQpvAZX5Lxu
yE/PyGbnWYS9YXBLcpn8ZHhg+bPEoXWKKmAdHluWiFEIFOqD7jBUdraCdgWC
drrYd9oppjSXBZeUcv2yasWX1JvVnYHqyzepPpfHjy/6dIUrh2a4ncHqdvO7
IkKtWyzdURYq+T//KxAqL06wctPd97qOC9Ode6chcbytpHGr7vgdrHaNSiLG
1WuKz9RUQr6jsa8Tx6OucRq1pNFhDeyocGoap6Vqi7Vunye6RVyVEz6nhTWG
XUUgokvfk0Hzg3n75If6pf1N4hImA/KYtcc30fYcgiNGG/hsDNDwwTKEzElt
pPTCyWYOMSmryivAyCnQ8FHbA5puOdEukjaq61stySlDY7qfvDF2xvVZ/Vqt
a9PDmXvAYMnc8DeRcCUgVOaUfZrl/WD+3Ht2jNNX1ti+2oH90yjhQwJiYMbr
+bFRCS4iJ74sp5jiIyORILGTSoyvZM9DR3lerHSXo9Ae3clVdE17dFc+CUmB
Oceq48EflQ5BDpSa3ZuJMk4Sk6V04mxg+rFfPATYzDKDEWjnIPDtmtnuIhQr
f4HvEsyKFoFqE2xYAONo3WXY8QoIF1x+IBz2zQUriHofak0mptY3b2zNGfaG
0lcSr4qClMaqFJSNalO06V/+lfmQr0pbQZMQ4EpwiWKvxJxtSwUgs5d2XTqL
EVMcZM6oidM4OiJl2MGRg26q5jhT/ECF1LCBMp/SqZb5bv4OKRVwqdsE3WaY
fuTTepvks7925cId1mPHVNXs6LJotMc5i9VwXzyCxTEgyJObYeEZ0VtB+XwT
kjnpHa85ANltamT2XafLCIOiNWh4AWEpD1VrkFzrO4bdP80l0znT+OrU5YgN
CgetYgm24KJgiiI9/tJ85MYat3pypSdLKzLx8t+h6gEVZWjKuwAdc+VYU2yq
kK6GDrOfAhURWOp9c5omFVbHX4OTnjuYKyg0b0csX3ejXuJnrtRyXcy1kt5w
oPLMA3kzZWk7DoyGQoMumlP2qLy95+GAa6Abx72jqt8DcyaBJQl1jQAoQSA8
SiatlAAw8dhcrW4ZDEjTkvLJ3UvQ/VgrjQGalsmhWv2ezNmhztCJmM6MGq+Z
npAuRhHZLOnW/klqVfYUhpZ8OuKxkp28kphNxsR3V5Im+A6gsjOeYJO4Lopu
CxiA2LrEODF5aFGA3rmLEjCs4MEVeEqW1H/rV/DNfvFTHjNuY9xVPKKHUglF
PeeYAcTkIwiu7KToHC9sWyiU+j7zeP1RXknJdv2VGoqQWSeAtAZUe/ziCD8W
md+hWgsMcLPeDhHa1NH7OEf7uH4NLe8N2LOTRucolkb9c2fdUygbZfRAADMX
VaER/6++MYpYS3TYpUUyV5gO2Vt9tG5mASSmbonn0/YDMhm2kbEyfHRhS3wk
KTf2BhKjDJ533cZbOvE6jB6Ux9n6ZcS2bRDc82PxRBZY3U0FQWAKq6a8kW+1
R+Z64KO1dr8Hl4/qoWohDh8rYAuAgat18C7Qfe36EAjAqfHKHz2NIvK2YnJR
UKmmCFrpj33sylhOIcmcALQnmupcZADx2yuEgJiY8M3Skzk2C1bvf1lJHnkA
5sk233Scn357cMZxa3N9C8M4Ct83klsMbeb9SbiHOZZN45a8XPZIiu18EiYT
Cg4KDmS9W/O4t2E2pXSDMijaBlHGB11W3rZGrcCMtbYRoBDRG0r9Luaa5f+4
Aipg7l2eMOwNhP4whEnjfWADGy17WYZ8oA8REkZwFM/SMU+c5zs4movTrQm/
CspnDsD5v5Kay/TnaN5lV7qSNOyrO95Cis0M2Vp7RgfLoBIVnTyNuAtijp1o
AjsWRl0nPNDSGeEt1HBKZSr8rupOsYtpgnTgHpqXomYi3xKy9Zwo3+9oo34y
XFjQbgyQhzLBNZYoLzDXmw8B7vWq1tFFijQNexAC4GKjpUcc5B411EMsG3g9
5xnoJ0bgzdcgFCkly22OmkzhZ5u9GLiUSX3pjvg3AQSGFshKjZrDGlR5jHFb
neC5CIGkAOXRuJ8rG/U8AlyqutO4rnLaA8UQkcxZ+NKYichwAL4I/1jYiFgs
ojJSUAg1RhXF3Pu4/1EFTZkdb40AO8gY3zM+GoLFN0asmkQGvhEEeQAbbiM4
H/j9/cWGw2bZI8t1G4JG+1WqoQtqIx5emjqAZtmdFMziYPh8JArDrAvpsSI3
M+5eWHATZz+DSh1UqSUbqlOULPyDPtbRwtv6a2ykc2TRdQ/xj+V+LrJ8o1M9
JObxoTw3qelOuLYuyQU7ckaevMkjMtrfXFUNGFpllJ7s3Ltwt69BCRtJr+bN
Sq+ssxIMrI3T0lOAL5P+eV2/LdbJ3MLw9DUCfe9y9DFhlDM0fjnMt/FSReIR
pgQjWIHtGgxTK/pt369aljV1JLgj65v6UNFPO0jXr49dCDpFVbxNONRiH3La
LNtx/mbYmxic1hUIiHOsG5FhTxlDvmESXi3jdx/NBkVBeDDvKaAZgw8wt7UR
a7Ws/7ViuFHbkuS6iEdATjwvG90pj/Db2CXvgGTAzuQ1u+f3hazfHlRUyfb2
WK9c21BLBq/az2d6Ei64MQzT5ecA631J3HA2U7cbdjvPHWMFHnp/SlMOZwvp
hxiGHZWt5Y2KwXzUR5V721fqmHUNGj/CT53DW5Hed5h4vCU7BGUt0o3PMT8Z
5dwLkrBIKkXVNxw8nqIabDMNhW90NcDCN0RfKeScUdO7rY0/AIKM7Sqvi8wY
yOS54QMlnMkk2/txI8zTwoXJsQbDOLqvUJHNAr6Wx+rtu5nkYOm8yPfjPDFh
utu5k6PsG3ObIAl4gpIHJQFzG/JUgAmMGAisRooHYIpCJCZJJs32N4dE4SBh
BQxRFKSwG1k4nSDpWVIwNsYlG8RWOo80OMyFblUzoIVWD5OGYvQM7lHrHWY3
pAliRtbD0Ha5XdEFEC9DXhN/Ilk+/kLnuTJAUDON55GmrGdGbkIQRN8t2Wid
HwR4mKHSRcU9rm2y3LRk3fee3agdodQ1FjZICVeLt9NX1Oqh+MyIT/3R1nXn
n39GbIwZ4yT4IpgN8i9KiUlclXdCh5I7r0ryN7ptBfNP9BWJXuldZ2DmKIyV
sy4GShJEOS7KHro4YSZq2+j3Yv6E0hp/4+PTwdmBGxv37/cZF1jG2Z4WlZ1u
hE5zqcEbmEFZ5faaQxJBuIqwsZSPf2IQCcNAEfSbKvPno+JxFth3es+kHeL0
NUafvxRhXFpuyAsKtGx7zTIRgV5aNJrgDnlWlpfc6pDQk0JDhCyvix188TYm
GZUjIyBegPD7le0ot96DSxwKcrSJwhj7t/W5PUnXD5eGlaZMue1yv6BagWM9
7pQsbhyNljeN0REucOZgD3sJhmIvrR3jTYH2cxa8Bu49lBTYodq3dI/2P0UY
/0MTqhcl+0qon3U+A0IqXopAaQK8v1aDd+RTB4zg/m3B91XUPSPKAD8Md50r
xYok/0dF76uUcvo/6+B8K94stEB4KlqH7cn+HTbuBCztDkG2Hqdu8d01K5ir
slNWR5jHzh1Cg0AiuAK0jRs7I+sc6n23t9MBIXOiVTha4DAuK9ooSB+OxUU/
W77FzvPKSG5ZzGK0fFngyfG9E12I+Kv3t6gBIHijY+acENKmk71bfCb/bPCz
rg1yNscZqCKq7G/OtIDq6W0xe+rzYN6MCWMUBRovD5np38Ad+xtHURbctdUT
A2PK4GhSIAnbGo9KFmXWLx2VmhyeTQizATN6lpMuDzKXRxCnYOmSnmHBqG/L
WOOqyOxRJRtvPrYrBprRJJ/6sZxTjUu5RBCEMTl6CpGDkfyaOuopHXk99YbY
7k+DeJGkTZFMOY8964LTqcxSgnNR4d98S5iF4BQrOMU5k/CNm0snAYoDqohI
DVFOZVgdzFL3GHJbYa+y+iiFngPVC3HA2CDP1pENqyh+3RVZ9Jjin7hvMmDY
e9UhiVh6UaYvsUzi4qMTYqmoEDNiIe5WbMDfAa6scVnhPMA3XOq0bebCd/PG
zZSNPp0e4rL/goqF3rEDzMh5oBsHnBnhzZz+7N5mjM8/2wc1sTipQD6mzqhp
Z4YcyoOzB8fxqc12Q6hH2vLIdPZ+HyVl3dV1p8cePjwzJMVlqMzYq+IZCuf6
9yCL+FbyfV8DqS0ozUlPF8KxM4ZfDd/sHBfDLbjsk0VbTL8Zq+gA3zZNgiQm
cthLkADLFmmFsMAhduqVP4VbtD4nuxXnHzaBF1QoHO9kBL0BvKjG18/aMpFR
lcVuzMcj9p+rsx3ZWe3YXAXT3wwoEJaHRQEGQP82pHcMiZB7VqlNFj/mtJYP
I2uOVC0PYZx13OYG4OWZfVrFqlvCUVAmRvk7GiaEnTMjfx6lDt7FIuNdvQ10
eBag9WyLIL7aNhBYgDsb6Cs2jHXhCGRKkOZ5k8lIu9EAT2eyXodAJKbHWhH/
K8cwaSYts7DKLMRg1wTNiq1ehK7qYRrX/Ds+UeYkrN8vZfa5GC/7ytu62WLZ
gpewNG1Bc6bE7HxKcznE9gF2uVFcfl4jeps461eZ3nnqidWntbKiBPaKCSQb
xlsqvx7F2HXIsL1+zMQOwfb9R0RVoZIP7rSksgq8NpHIv4w9m67GnfcY8vs4
JZtyMT8CIMj3/xwG4qx1mgxOxMJJykVvfLFyvxPEDpRHqMbbsee1c9d4EI7Z
Z9+bcA4tC7sWndcYLznwM8xqxCIweJOCfLqiRFkse7722DJmEaN595BW0ZQT
OX50CZF1pYKjscydjhQ03W5efRHnZG7EGevpaMqAIFCMlWUGbfbROoTO3tKl
O182UO+OlwE1WDSz37o5BR6V0dbebC3WKnorW5HkPdeKr8/i4zzrdKT+PYUF
IFmUke6GBS3qwRD/O0OTbQBFX5M3l5LLAze61DCR9ascohLReRtVjiuAi9jg
pCAZF/QBZAU1YT43yRQI4Odp4djgxkGENPOv3O3OJk4E/qZ7U1HJ8XlniGQZ
vGWHjvqoS1uf1TB0N5x3brCrCIxE+qFiu5E2XxXh4HflwHvSlW6V3oUOP5d1
2nMVwmGfaWPCPXPJb9NYU2Qe6vXRduaNwVnf2Qvd5Xh9PPpAo+2uraPf1GOd
ZTsg0d2WDtCNQStaYcYqhQ+j4BBehIvERHtDaTzWuK9fYCgfB5aku38NvCbQ
0RCbL4uP+cZJ5eJ6cq4LIRPUiwpaRSNapOhsDKjBg7/APLt/scI16aaBkikO
wl7HUq3VCGfspgSKJJLh0yf6ATeel0zi19jf9BcEj8oBhqn/fg+RVQI/CQ6x
pZCayPxIgOizlcheqw2MAASwdtu3W93MgWkJk5LZywE2LHVlbl6DDFQW4Pr1
vETAoF/Tk4T2TY46qzDDq1PQTXeHhSCNsq2rOdhaNZQ0SmqZAHyzjM+dGv+y
QJ4xHg777lxFELvVtqtIrx8gUZpYWW3hdZisBC8xD5CmiUF+Ot7KEcf7sxVA
XRakh10l9DsS1MJaUnDUsNFXiDpgA5nz1suQnNBgP/bG76P7iQ7Q61rOkjVF
EtRCh8Cjj9wrqIlwxq9ovWxBksn0ub2XubSgZMtN6WPMYrigXgPC8ALKMTzS
3dKQqXicbhKLQhFhyO0+ybMmBvF84AiX7dexLOpNzLiEkz5g9DTgD67zzu4U
MOeIwMaQNdA15EKfIKPe9L9qBN8gNpWVjwUkOAHoopHW0SNnXZF0a7rS03CU
sltvJpIqGT0+9zfMRX564V9sGj24Zvtfl6qSMrOjD74Pfq23gAhR5ySEC3Oc
WWZE1XyZz72tVsifh2+/IZAmCfaxGAyRWPU/nD/T0nJhEw0ir+sW9Abu1mHV
jQEmcu++RSrMRf0XmfcwG9WDEHRCuvCxcitH8S+etkaR/uMX30fjoKkIHDOk
8oi4Mysk/idJ3bbf04ttTlm+/YJKtyna+Zp+E4RTmP4p+lHkVVKcsc84hOM1
fSO8N4Yj51X5W5m5H7k8+GRdN1Q870CPuandhEx0gsm42nQ3qTF3RntnfFck
Vo32cRc1nppUV0lUziFpjRV+C6I4XcUYACfjiZGVHOX7llPT9bfh62bV8gR+
ltEv8VewnIUcsYt5s1okEHSI7sxJi9XUUVwkRmRfRxEd3bny8AP1fQRIDbnm
M+lFEU8OIv41zmEs8MFoxOTQwQP8szN74kHxDsbTjM+JoA6ZjbDDONBV+EyI
DtKUtQUF8REOIqVjw3NaQiaAVopKE3UHhZpW2tL8aM/Kkw/8Vwb+3fxb+BVY
b8Q3HsO6ZDDM9n0pSZlwCMy6IjBGuYoiFF1B84oyBncPy8e/Q0WHNxxEjPnI
waXW33NGvNM+Rb+rOovyFaXftxfviOXpobllMAY6dpj1g6I7t+8iduh91MU0
QJHKvSSXGNTUxTLYvvVZoarhW+qv12g7wPRku2Pehdu2ygbMC0+rwA3ASOU1
1kMlGdTCgqyQbnH1ma+bzPXqtuhBfFSoDnBdmwrDk+0PlkqMtZsqYXIDZB6m
IL2TWzP8p+iv6yuRaDxnWiZP/7AHAUk3rZ51QwDGquOQ3G09Pz8dCOiic68d
zGKwdzHPKr4rRJQJANSZ3f7yzR9yS9ovOT6P4gNYogH+Lk7q05ufNs0jooML
5YGF0RLej+wS+7xG7nKAR0V2TZbA6d2KDPD416uogrovVyEY3A35v6qrIhMv
k43w5AAYeCA7SkQO9Fo6pxtvh43FLT4rR7YJKw7g6lMcnJTn6RhkdMaR+6VJ
VRCjLzP3XLTkYxlsx4o3ayjkppcKMEHZB8U3sKIUd3IP5gGL+9A1RFqFuJ/k
T2z6gvlLzCtvGCkic0ZAev0MZz/sc36cOouxOxTEVsxUepCgOBstQCdd6MxX
usfuQWbh7jqn3D6wOMGzYglyBwgwBDQLWg9maN5ovpUyQ44OLePesZyrRTNm
rNK3etYCn1bbW84w+c77apFaOYDYhqH3FYxBW7BUGuTAtH3TRXnSQpClzpJn
4kfD4pdlBmsDzG9fMFwYA4y6lqcCjlth7V5S6DyBQ6pVus9BT8xMR4AxQAOm
FwJog72Ab/InyEy/89DN3SY/9SnsTy6XQxB3WtxG9sHTi1FMvXwOPkiBosuy
+CHS5xoT0uCd2vlkhgfRq98xOiHOwD3B1cEXIdh0C9Ek5pi2qSr44cPFbaPr
wBnwNQrW3QPZTesW+Pme+GP4NrPLyr1tLYvuHrs11a6bUgp5ZzK3nsdQQOf5
DkL3FqUw5gZ7JArdqyfEgw/9hOOV7bItt8Dz3p7XvKLYqvLei7BqYZCbt/9A
c8/40n66QM7hSe6fbsDCrDrlmWtM94Uoqu8iDviYzExRMEoXDGYflBYrt4xZ
+ChRTx2OkJnV++AwJVmJMwdfL2HBGAkDzYYZjouQUuAyFv0JDVJzzs6lzWcs
VtjS7PrhhBp4xxXrtNw+1fWXjEnw6acbRvrM/C361/L0U6SsYSsnRaKtNfg6
k6cJScK6o5DJ6H4eaOQ0zvrflHcnFrt2ylJ/12DlYy9dmTcnF1+pMt2gXaaF
r1XS3l9GKLN2D1HD3XW7o9kKT7zmMB3r2ob4XEc5jvxBujNlIVJ5r0BQo6Wz
fbz3miLH6qvbD6AYkSDsUSxnFBtb1UwQVkFPqeHQT0j8bOAqzzQtUNBvzjb0
77NwjDCz2tBnvOgoa/J5cHM0VnTBqUkIjKKP2PRoWfda1ZNMEUjO8O8KzUkQ
fCn2f/F/vkZiPXP7p1p15xQgXPT/crSFVwyYgi9sXIGkkI999XBvX7vge2Na
3Uz1NEUO60sV+r67ENvQQPdK9+GPUaTRE3TTFhoO1ORkIau/587U4eVojfEi
rLsjdzI23OA9Vb3i1eHz9WKzzSaj0Z6yP9CJn0J4gdgVXNncCwzBahZtPJuk
0BV7P8khBLqFAljzGPb/lBf+VnjqHWgFn3FokxUrrOhonq1bO5Jgfkv1HB02
Nry8l8OHUJ5VzQlfbXBhFoGsIspFE2Iqr2NlL961vVHnVIUgslU4vlrGBoV4
8+AvfzWbw+ZexhJxc1AqjThYYiZHurncgJfV7jcbLgwrKbb4ePVVGXzW4qAL
iExZ26JJIwDhdOWawLhoH2vZzOyPdw7qOYzH+Nwbh4c8MQA+wajfO2roOKn3
4i6wKjOwDp7AQrab//oVzxY0vR3V6AoRtCPNcaWR8aZSaDT1XzPgNLJkM/SK
p+FLAKj//sxLTXhvcKNUIgBYynkum5LryChOL+WttVslrIDVT3MlklqhUOUJ
fXTxwLAeUs5GHLdaLOS06XEF5X1lcwfMsFXfvZyh10dEZ9PPHt5TspbikMe0
f7Kj4OUP1K11tE72LMbGE/lOMbQ7guuHh3/t0T2jnA3haalsZNy/RlOVkmGy
L8XMpxv+tFwN8pfOpW/h6nYdZfPu1f/E9bGzmNICzpQBEDUHaT05KzeRSRMS
pfeqEwdx95SUPjAhknQdNO5j0AgbRZM3pOwonfyW7rPqeP0PS1eBcSMjH59Y
IpGdLAFu9dj7+CHdzY2R8aAtuSUYwp3RdtbBFqjq6d+LRyDN+67K8tKhaN/w
F3KtJbqTn7LMDuPkOJ0e0UfZvFqGzOlAqEx7A7jHZgaHCxD58IuY/6N5C5HF
4rRSbDrS9eHn+vDFSzkab6PV5fSuM+s55tLhPtamYF4K8gSRWDs9fFhLkDdy
aeNvxKKDl91SIyMuoaieYJ9guWsYMmMCTf66Z0kDjtBGGtkcluSP/bap9ljK
fBriUVvvUdUuwJWKLWc9BcbZHA1MLnSoiXFMriJ7Aux26Ku3G7OsdLoUjG6U
3bIR9cHYewCFvqa8w2y844PY8VlRcrXKs+cUuspuLYWLnx4bfm8IEiqFEQRz
R0Oex2V1EfU4d1jxXamV4U1dckAfPQWFIJqWf/ALIXS0/SZXyr06rl01oYoE
yjzc5jY+6WqmQCZb+Dc8ONc16F3SrabHv+Y9NqlZXvc3KMpuvW/HIKRmjoQa
mNsm6qDefU2c91S5qXvctIKkwS0+3fB0sxnfmqz/WgSyXkeIQFrZ4/JOUVj3
Y77S3tiipUL3IpVGseqNyO6zppkk0L1yaSM+3pD5xWSMOeG2MlhYg06yaifc
azeJ60ruYipcMcyWCH0bN6QOjTLIc7X7jq88n63frVmxMtGzfwfw80sCYrlt
an9o17AHPMzKA+r2t3QlesiO3jB5taBSlQLWjHuyTCT6H9R8tK6GOidS91ax
PjZyTrvGAJdFnpyapNJw/lw/7YaOZs4ZbZwCasg3hc2Y4G0ktM+L13pXhbhJ
P33gi52ZVoV3siphfjC98MWKevwWEjqHaGdBTOhrvO7Mo/5KCUIMMRm00FgP
2wybTR/SCHqZ/pKxpMJ38zcxHdNiQ2vL/dNoVVsGf9H6iYbGdQJ4Up9aPrmr
/SJcLXIi9DuKdVi3IlvCH8KV42UDlD7xPf1AaO+rPM8mBiJc1YmJq9nTN6Mx
2/klBh0vuvgie3RyDVUlU7BOnGsVIIHdXJ5SR8f5ZpmXPyVjjxTjsLKhbf2N
aZ8qQJL8p0G9rAZhGwgqsvP8xi6BCeDYRzgJ7xuncaRghqkRuVjoZQl5I9JD
OtnQQ60386nwJ5wwHxB+RA2Kz1Mra7ELQjrs8swPJKqb4bcHjLW6KjamKz8C
Vr6atAPB8tk0ah/aiTJq/e6l0vSlZrP5v7Y62oZ2VTfJIkj315bKnVCroTV6
066JMHcUsJOdest/6ugeSdrGTHopS10Y/gmEIXJF9x72MybKBEn+rsjQTTQh
EQpMEbbzueGIocF0AOpDs20WU5DFYK+6P/gYCnTxeBNgxqY/XuumJhegHzGU
cD2wLjV9ri0ovsUbTvgYqnZ1i5cm4Js5HsrhAqx3tKT1EixCXzKk5ByDyMoN
uP9wZafItC8BNR7yj+WGf5VyU313eFKYObv+HMGeeu1NWVIHRGutWHfr+HaB
VVjijJojgoCp2rQRCQ2BcABj5il7FsBwkV29/sVq02MFCJvw3lxRNqpkMVGF
GpezAcqw4cyzFOGKrIRUdypzIae4VRxFunAPBWAo+7cqWJNwO6vBv9wpJEfO
AqUM243GUNDEyJq0m4eshfDZMolImEWihmhbTWUs+X33hvyXb9a0F2gtOmW3
fYWDPq4KkNW+WbpfDV9SzOVjmbET+Rp0sGHG2phX6QFMlCTqlCAmau9Nx6Zv
dF3te44H2XrNO8l8nXi8/aAFM9JR/jopsy6HWaPTuXZrh8MFzpUNGWpowpa7
n2GZ2xZl+g6WQRnBE8ICOj86hKFI3HSUKXPraWivP92hlzEcp5IN3YdF0nw5
7xza6xfFLTZf/+HRdrZJE0BYIwEHV+pnLC67SxuvL3c2ocbc4jcyRDqrND87
ygIMQTmpSIla5yDOapuYajhroZntbnPmbBZrj3tpDA3mD8EesLptKhLiBJnK
gqK2gdBai9CAWDjQSZeu+nMpYd8D3FW7pCYo7yz66Cwopms9nI6+2rxMzNV8
o6td1dVwL3OvDuhv+KyKIKpTPKspEeQl2hg7CAFvZD/hohfaigADS3cELv56
F6f/D1MCUct/GbCo+vDW5c6bQUTiViWecpIjF0Lhqv3jsz+bSJtFtep3hxjV
5jMqVTm/9AcnwDN3LQgmiPp9KlvF9UD9NfpLR+nERU7ZH8u81dSuluiENovD
Ev8LYFOmC4RZE8ERTXJ0bNc5KGGEpQOi4oKCCF3g7Iqb5dAe6DjjtzpkV9RW
6YKjfSWV2ETfktZlhB4bcUUmhcmkUEt+ZF/3DzeC0vaLvT8z2l6XSs8hMVtK
eiQein2qrv3m2XGMoIOyDWGNmxzXsrrdP0AxO4ngNpChFhWHBrNovYUnn8mU
a7irVlYq+HI5ariYOwL4WWCtOyQdya7BGhWmC9KBDP8IIJwc7exfnlPIrZ2Y
T6UvJnKH9gKG3dNEGlRvXZuB6bpo/nj+O0awY9Yw3VcRgWYOa6TZp9sr2sUP
8adGvPYUfwbysfEeoKYVDHUjvP9jVU0O1wBmn7DS2U9vxuC/YkyVQmyumH6a
G0yKxKWxkBlKojlc8Ha5h2ibmSBQZP/elekWvcu2vNdWAUuGxgoVVpNweiUm
L8naKcqOUzNaao3W6V5K9MAUUwhZnbEMjBLcDFba1XAfLB0h45VI/2F9n3bJ
kcWAqdHj//Yz2AkKW5OuKUAOVwxRba8oKWVtn+dEicnLI2+sSUYW4Fdwzn7c
S7a8HTLQs0i5Gc96qYoMg/fGRgvMl8ptD5TscPc8pdWHVarr/6c+2giX57vb
SKhAZlTznKs9fNfsW9j2v/c9W2cSjsKIKJvCf1GkR6B5tx5MAdZxIS+35frE
/TC4PEuiTiyX1qI+wfNrji4ditucOjIz2LqzmhvREMHD+l4U0hOQI2CbDlJo
xMT+gaGq5wMAjTm5yJlKiBDthzcjVo1MOkrBgc00qw7fGPUBnqwce4AqxxJ/
oF6hhhH+230Do25v6sRfXYfrmQmuVQCf9FAhhcOLAlzNrsIa54BeATRcgVAp
mjkkRiyKAlWuh7KuWOQMDfCsF9XjpeX5FMgpbE734ly99Ou3YcUzVJiEbbAP
L1OAl+uOxjRZ6Uolumm+oQdXCW8wB2UOq3elbNQzzmywja2kgTV/yyv2RAHB
PIGCQHNSyXJ3Tz6Fu6aQSVIAMw6UTlEGxyJuBki+t+A7LSwHtFTAzGWY9ysn
+Mkacq5IXb+ParNXtYdzBK5y/kTI6E4jsB+T5+a9nRuZu9pTEpu8qKhxvpPx
Ko0DVpRIRDxx2yoAvk2FpSTnWqrp4zju9jhysQnQ090G+wUgOp00zbzwxfxa
zSaxtAYnZbD5HSVbjBN6wL2o6kTKTsVUihVP88f8Y0xbaLBXW2kchWFtpnDh
VrhccE0yuGFhbb8C2FDZJ4QHHm2U2S3/ZZE2UX4jLvmxDO/oq8eM2zDWAl/K
iKmyCjYJU+ciZy6Z1r5XN2zCoxNyBhZwTPHv08tLaPJfEezVlCxsEfBTjCIp
mZVhyOhXNrrBiksJnT8CxSmFR/k6PI0p284tRCU8IBUydvWmul7DHt/MMrEy
SVkmcTeqZ4GDzu/nf4M1MZYIPTtFQ5M20x3dWHOpEcNiComz52P6lsNGd8fa
40rpttRrZysO5C6PbsHmOAg3qGaGsN/ba1QNOjaWnpWpE51O+dEtYxlz8Pvq
WyKjoWNAlYClyn90KDxQuKAevM23UgshTAP3oLZgRAdJS4k6Z+FNDneZOYgt
JX/C6tF2qmqdTla5A/kuz5dXM1oL1EvUTFEmrB+Oiz0ZBaspUYf0imLTpqn5
OAvYPyUjxTDLMdkPaoZO5PG8JaI5H+tC5aRVpQ5DfhWxiXqEZE0H20hKsrbd
dH4jkQrnciMUSK/Yar4a3/MP/5C5kwOpBgUHa+Dh5VZobzC0T1xLVqsUhIvW
wuPC5WLioS0ZiBdQhTWBHIGp5xpu5My1tLrOD7HvJ+ZSc1Tc4IAUXITJ9CfC
6W+ZIMT5LWLN0LIQAG7MPQ6ltqklHN+ksLOxy0RohF5V5re+QVtgTi/Se0of
angZXXy+3nhf8zXsLUsWgbwp/20qTO+OA8OAbXEtMJntEa5Xpz+AIGblTIWA
5fjEEh++kJMB0y2znYyrjgAK9xvYL0172YkF/1sraPgxlkinxd2XHThHFgab
2azAhQWh1NrhzovJC5XGt0Sqhw7oqcRgTxCyic4PQ947vW3+BDgVcZdCIYVw
DuXydmAeMpJLRnrGAhw6rUUsYRyN/QpH8vCjMw31RzjHIBrQSEkOuteQCmcV
3rC9zKl4AkXm9RKyX2kazQBXUgOBHu4PR+khEotpxG1AYmRHhgJlJtJF87G3
KtOniPJ21E3QEQqOELcoYXvDo1c9FphAkKYuIfDL8vsEs14dExdq90feFIDF
2sI2HmrNVrKy8+VEHd0GxfT1zs+caUDqt4K+ZXG1XKS/2hvetxmwa/Yy3evY
HVkXlWrKQmDXvQmCvB9kJtwXFxu58/dhrSeA/QM9gDajl0Hdvqnacvp4LwWy
r0/W0b7gdSj54hIuCLMX+jcuoRtcF/wqSZnS1/+v446F9wh4AXxgux4O0QF6
lRl5m2aPGACNePDwSYhJySq5vviSmC8OgdiERciQxZXyWsmVS96hucAPz+ut
K97XFjb1CcLZAfhPqsDvOd9Fy5IrBp6+VpNzaC5surNfRafy9kvUFROySVaQ
+3/gBqgvYQ27yEkUAe22g6NoDf/d/UR6cTwOOBe8v53eU7HE3MwYN+36J/EN
ANXJ9rlSrWrieqhLaLipqJjO20o3pOG934iyKW4lGz9rAFaiEYVu4xqo/5JS
CPGqXmyea2euLu+/Y9eDFxQzVArAErHexr6q5bx+U2N69FLFwEA/YsQLsJHw
oDLzKVrz1ht33dDsTMDB63WZOnaiIc8OKIJMFu3mWILXjidgZSuww8FNBa8A
1T8kn3sFaYIJ6PK33Iw3yFF9s5aC8oXQsev4yOrobuzZqem3Rx/XLCt7G4A/
kkvT4T6uFcSUIkxxZX8TWdtJFvNp3BN+ZoeulAGgHcxsrvP5syKV54B+sYCo
TF5ABETrMrqPJ/qBmlQLg3i0kwMEzoAVwqdO9d3CdXQRwdFw8h6dqE02atlU
UnNKfKc1NcpvW5uI2e3XsYKOn4AeK/kxzYLQ8/1FtXQP54x/GhA5Fe38D3Cj
1m9yc//tdENDc6oPDVro6lk91ZbQe0iPsreuGSV+buq2l0sXvoOENI4gHrcD
qcFxe61ENTqZoCBu2B0695p6J5PP2cUyt/iN7Z/Mu+LbFwJhdBlmWfUCmX8C
wTKAz/4hvdj0Ry8xRU9T5T6VmrqEXYiFPoWGQrBf50Iq4hOXSkBKY1b5b1uM
AUYm0REnixibEirGGdrYrxC1lyp7Wwyeqdwsy2DNEHUkPEGA/5vLR+9+hRal
3x0dzzAiitHNrXvQX5KoNGmKmUbP8FkOoVEqxH2QY3qJ6zKwi/hGJTZyGSAt
G0j2j9Ym9wglqOt8gzivaXQD42zWKqyDGhgVMyH3qJeGpYJKLYyYQArjf0hx
RGH3XmbzR2h4HwUJlw6DyWk0XSDgmHJ3/LlRyg1dgiwSjWx7aUfI19DqvzeV
q1AUi4iZvOpQmVAjfP08y+Msklw6DItDQRwnUOHYdF7a7WwsMhVdCps2Yh/q
dyUKlGwQtsH96JUvWp9ZODWDe0DCoWZepmN3duZoRo+FfFajS91KmQ/s0l0C
hbkZ8z0A+ainUf+wpUeVWd6tvM00RRROK1B0YgCTBPknaPnsQGrTTz9LvgtJ
B16I5EllmNPM44HxhKMGADIW9EQ5UCAtNLKtMvby1eoJBmGjNb3Ul+zH6yAC
KhY3LWZXjtRL8ZPDzMTd6OaBS8q0809a7zTfku9VgZ3ubQHVDNeFUL5qgTim
fULOb9KkzjBt7hi3t1YLiEyeA24F2pXifIKNK4EjOQZ/COp6Fe+rENVGVRhR
LaiPXphzysm+rJkPKI4KylKrziYZ3KvtphccqaIhmi/jttLktQ2sbXtzZtL3
ftJeKAZ04/LHYHdfheZ8w94gRMl8/JLcI2g3ow4kg08WEB7S4aBZRQAF6lUS
81m8wiZh8294avdoieZ3PTPENZ5CZ8tkNQdIG1Xuc2yVO3rKMEAQjyxqi95i
msliEFPPTrJ8eqSEOtXcnVga75HuEz9SB1WTXpR8qZjiC8s/95NhBMZxxvFt
BoWbXXiKIseTnRQb2QEVJUY9FSiqLVkhKL2NPw6idW6j1d3CltbgGhV1a/k7
ZsszVTN0QW0p6SjuKzektsPf4/ju7UMePhEzZ2EvcuwET70f9mdV3EuSyFUr
zyVYf6JEUw0gdZsshlyQMux28cj6hVxo5uTtVJ2tCuIqtow2uhoOAg9cNhCC
2/bU2ON6Ut8BaxOByrxQq4W5zJVyP7F0mpx+8v1mmI8nzyDf+920rcJ7SxIw
tKBofBzUdqYZAy3UELf7Qli0PSEHx4ANJZmdnHVhuMNlQXUbNx1CG5mNqux8
q+rbisTMF+IjxxdzFRU2UA/PTWueaoXbk3w8hShLfB5Hw65zT3I0Ct8MFfTH
GIcnaPX/bpdAJgENRAAWweDIV5Q9m8BhJNgKO4Nl3FL7+4wvQu7pVzbAxW4R
L9u29jlInILMyKan6STLBlOwIVUfB72onPlokK/H3ZPYhRmk2n8wHdxsnjsg
B5b98lvr/S9PB/jvbyLTrtn2jnaDCj3wQC0skuzVUqTdLOOFr8wch/Gwto1t
CSQMTX5umdryTO03f/jZF8KWF7KYCqSSsbb3ATXjdPc+HivF03dENwNat2dX
UUgPjYKFiQXNSJ33LPqXfBeDhkZcO9jLkg/sZrHRdqdJ9NfUyTEE5d1lelaX
11DGd/a0A0Z9ed84Gz3CxS7YfmNJzawMxHIlnfZw732RM/wF50K9GYk/aJrQ
I2lYKK6aU74f0F37NOOlOn2YUUgQgrAnkbS3DPtUZFB1n05PDOngzyppWu/1
Uyqla6Gc8Bp2QC25nkXi9SLA9bJKIrWcuwaJk8KX32o13nln+Cd6iK5Myjyr
Sx3CsLEoFXp11N5t/QCMld6RaQTjajiuHeBeI2ADSi5fe7d3yasGHdYE7M+Y
2e9oHe98XEFLBzF7SRSLIXPJWHc0H7zdOIYU2VtkQojA77xxq3jcYcXMVGYz
9/ctTLOG2J0PUhLmebPpQRKgWyBVlNuLtJVjww8hCPg+F8cXoxOPP7lVCpMo
C6Q9GoXPGIyGAtO5tcn8paWdBez5skhO8x34QIERfa1TeVtRemGO3dkdsvvp
0cUQez86VP3FLHcFFJowXuQsbrAtUSfvlEbkTtqABBfIRXFsl4v2t8nwRomi
9jZPSgBJLubJlBJxcoFBI5T+w+gN5rIj8hbNkUfTk2H6dZRxZ9hgTBXtXUeQ
I9L3kg1IrGsRsUelmshOzK9MUonOh4b+US69SJmQmEVnaoyZ2soHkGMo1wsO
Xbg1gZlPMyxmu2abCAetfgdWxSn0okIvvbp6CsXuVfU/RuLGAvRu9v0nzhIG
3sM5dAGc3rHUxvxx6sbAD5OpD+NtMlorSxZlzIDV1MM1BJlp17kR9bOOyKgO
fOVK/7vn43OBPpvkn0lLr+OstDx/78JosDjKQZzrhMxk6T9BpxtFdpZLo56q
eSIMX6ly5MczMQuF/HuXqz1nhNQLsm1+Wvk5wmL7IkDIkyX+s7WslwhdY9oA
D7Jw+KS4ML+WdzgZjFHQyyv9iAgB1/tRCw/Z4RyFTcqCbH84eFIb62LCqPwG
adze9NyHsyUiFjvKozf+LPQRZNPWkzFpfh91SsnmnL3XKvpW4YHZygbHLq/D
OpzQhBldY+n9+GsQ3I556qshKOPYoFJJXAZf379Tbcv8xTmzY632WkeXchTQ
aFxx6goF2ZrWixbXWeHgvEx3nUU20MFrtE+CI9iH0QfG2v3zgN0XGZcif6Xd
RY2RVDIcbJCetq+0j3a7tH1Z/9SRt59LW886BitFH/qQDhWaeqvwFqDiu4/E
ZG6t2Rt9m4b9LOPSIWGfXG0AtDKArSljCkRHOkDBwfgSm0Hip7JpOYgFrfSI
iAoavYOI89+BjT02PuFq5meDU2Avvje3N1AmPVepcxIaiT1Mr5tcTkW7a/bE
hC+lw86IJWKO3b/hNgqc1n999SRUn1C5dX+Jy6zXF+82AYuqy5LdmoC7Cm6I
8JXypUymF8ngEtXuGt1IQXbAQ7w0jfg5IpH2WDfrdKd9vJKeZyOz2Bvk3pHN
tEq+4iBzJc0S2K9lY/QHp5A1fvS378hVEbS755P5+Wi4j5QQadGSHgIeHi0S
lGNyG+B1MRHCQObJAViQ3byUM2u2iAfdEj2fYszIkzQdSkKYnOeE1JY+b4zz
Z8JUNDKQIoIrtv8Db7j9C5fiVggoIUm7h8xZRKc0ZYZT1U1uTextG3e5Yspp
ENYjQc42VlVOf8VbXz2CDNyisBSPhLoUJTih4eVfQv+Ga9Qgp5XeF/qBA9AU
p39ST2/Fr8fBa5yyR6Zv4fz5aed6H6jR08+k6YyB32kxzXn9ShNgPfl0XiKU
oMpAbKen6ponaHC8gRt1ClrYS73bEOy6hh059AlBOeGW+bxpvraTtsxUrK3G
yCbdVVVdEai04gdor30KPDxE4cU8b5lCM9aFX2NxlYuJ/w0/F7EK9TPYwVo6
ARFBGtquS7DynqH2JjTjQGXaPpnRC54+PH0Y0hSjfb9x9onzllujk9zIJgn9
ggm7WJoYLn1zKkFmk9QSXkdTlWRWqqAJdF5/ar7FI+v8+iEP/cNwxLu1uKMG
Xd4A2mZx0LiFqCB46MrWh4vZNTXRAO6WZ3TIZrGH6hf2np43eIQWS/OzmFs7
GGT0uBuzC2ceKreYZzn1iBasq+sA2m8TPBP4DrJz/BTwR5W4F3Mx4fBcPOPE
Z5JzzW8thluzun0jHQUXV8zu6vFDcVsyP6UZu3IXG5B/Cz24LaRMyRBBj198
P0uF5OhDKzJbI/oND71yRRnCASOuwloNLc83eig5njrPU/B6JaB4V0rftAiV
vjIIOHGzBMrCvTevbFeAvMBcUcxA9Nh0Lv9gRk7nVbijpVrG9M+4JlxYLo4O
+IHE44hZLWNoiViqx1Zcr825KLGeYLWCYGgaRjkMj5pMWWP9CCq6q6sWCNLH
ztLLBJ0tRSfkFY702ekaY2abUB3sj1jaEFxvhCQFzkuiQdQ8jqNkgkMUN9UZ
semx/abzijHK1mQo21ZPcK7U35lXd/a5e5A5xV44T02xc55e3fSIqelatoZy
1UlL0ypCHOiCbXxPXTEm1pLDDkdSSwqJsh75JknH53KTC725Rx7t70tpeEPF
t/HYHWFvoW62YkRd2HrJWdI/Vs3drl/7vwrWkFFengWx+7OA4W1rJmat4gvQ
2zS0DoCLCzbxAaXc/VSFJbFdpKlyn594SIMIfgT3lqcZHapQ13UoDud3+sNO
R9/MSql6Q2mTJGipbvThYAoABobanGJDeQgrhBXkKIhAMFnONF8NMd6GOISf
V5aa+KxZlGmIlGiu7v3VRAl/dohzmgK/Oht/PVKo9sOR3MnhtLOaRehebpf4
d9XTfvE1XP4Zd05FzhPCjPVhuwiPMIULjrSWDpPKcJHQH1O1QoO4fFD2tdpS
qtTk5cFae9j3uD8yhxIsTClqHdyiBA6aAW5crtg16R/YAEayWgE7Y9PvUSg2
9cE1Jw2FEevg+j65QTQpYRBdQel/uxrfeW96zKF9lH98FE4yvtFZ/AgAEPXt
xkfdF2oFlpYfgQy9Xrk7tOUIImArCplJRgFo6jcRfZUdR6ofWkCAgVqHNHJg
pw7qxKzY5T+2S1tqNFUQRVZcdi9G8LAGSwQ7/+nt12qRMZknVDa9t6wrG41l
CbFCJFnOXBIcqHwQjf2BaeYxHxNLAJ0soSEQ1pOcO+WPklVnrj+88I1r1n/H
h4K6CahAJCVZzlR6MS8kAQQmWlfaWmzMkHhnlDxRwdzsByh3pwAXGVukdaIl
/g+eZWhr19IJt+q95ibiU7mQ/ty4LuMLiFQ1/KPdscTDeGbs1C/cRZ6pCrAR
0W/dO0M5MHzJrgXTQOGVGJYkyH0JCpkhABCm6M6l5q2zKxTddAQM/f1iY8/0
uOMrd6z3MPiWOx3M55fzLb3/cKJWsrznHtj1r6+9QL5pUXrnIwgWPj11PGq3
7nqEH19v069ePtFgSaNLJGxg7W6edC7pjkTha3OMkqJ7Oeijeh1e40viQRr+
zFQA+nusT9M1ItLzpQpFHOl7zHJiaTs6HNf83ZYZybS4ijoT/lsD9on+1CDI
xpEGtdGP9DvlM0R/l7QUHJEeJ3ouMFDspU2K6OrMTEOYO6Qu/d1YqCd8CAaF
CEUua5Ro0fKqHXzUW/GEa7XWI89G+0YsxFpeh8BkljyCDelpKBphzoggRZI2
UIrEfzHwG16bqXP/3LAh+6cZiyHpNO7cQTaqFLSgAjQvm0gjEFVGsI05FD5Y
tF5l7CjYb6dtxAPc8vEU6QYq4L90kmsPN4n5m59Agnecb8ghhCpuZ2c+Ahl1
gEnU5t+Y9sqzqH7lD4C556oH59Gcp9FljJJodjcINEhwvyZOBFqS0TcklVde
DvuR5//l9zsJDv/Da1iIBeWSDV8HuJpyD3VlaPmuxSWa9Yf6tCNQObDxCh3J
YMgJXHsr3Owv6GKaca0ePbDKjFlel1XcJSEV+mfCg7ntUd8f44+/euHoce+B
AnPqc/CsZrp2PnN7K3KxDBVhZz5azlpS5VbNWFwF8JDQrCBYvv2dCv5fm1pi
KpsZDCr/9UcVS1Y3cZ2p030IVt7eS2ajKNaS8e78FPmdgJRPS1fd+3U2ijix
SvhzmC+xOsXftkAfuKiCSz2Ztjuse4G0uFh3SDAZBZpzAQMQ2xY9XCigvmZp
Ul4T3iva8jm0rHr6j+v/Sj+CHUYdLuK5FZ9KcYn1WJ/L4YS/pBQr4PBIMYEU
VlM/cX9neXOL7aEbK0SDKzD28SbsJT180ry4i8rBN2Bjry2MdcLOvocUh86d
ML8mYdAkGJ62JgDxyQ+6svYIsc+biM5M4vrKzcsgy+HdL4UKQrCVfjwN0RHE
/u8vnxeqbBp+RbILmyCPp+qf2iKyrfb/89h6PnRh54koYJYypIsBcmDbjGbc
26EABLDJCOMWvpBg8gsaOjmTQIBdS3A2PH28EvdagHY5gjna0MQ2ky1kGCtf
po+m7y0R6iau4QsFYYU2jOrARQSYVw/fDw4MbBq2mP7SiAlYeSWtaSHXTI6U
RiweshGT1BuKsWOM5mc0MVCqFUCYa79Q9QBaUK1IC0pPrsSBgwpwevVFlVm/
Q1I28OEXHXuJQlwVSN20DkRWtgYA3Zzqs9p04SgBX+hOzeLgApbkWQUnB4kx
hRYRlcq2IE/KyY2oMuRbfWQosr9bdJEc/t7CoDDurdYdCdX+RZPLmHjMK2IN
g3HhJ3UnDyo1kU5jN86MmaaS1JemaVtZQkymF3/DVR9F3mqaNvwuMKIB+rc3
tdx5JlAlInsZ/3ZNavlAcYRsJMzZR7rbgjAvYngPpcT8824biHFmCXQlfuO3
JyHNPuu+i3VbrjFOLRgjmwByajDbBRRabU3da6rSq/MpTur5rmyOn/y/MFYz
ye6Py8Q1wwk1ZyfNQzOsG1rKEbmzN1cSnZf//OukKSi3y1yraEXuipndm0QO
mOshMucz3AVF5IR+PJRaWySdn6y30xmt7Ib0qtPMq10nl/IC3M17QfTo34vh
Ubb7WCNSeov5SG4hNAUGvF9rBDWi18vvcNsRB36xseI+N3Hdratmumhi2L88
RcccVf8Mnu11jgBF1DPUbJ76M7EDUbUG9MGi8yaQm4yvEWpCjVv8Vb9QhJPu
LXRypZ5Y6lqaJVTN0ez7k9JYi7r7LGbAcyqZaZ70cruqDrxxhI/C5u/3EqMP
8qufg+glVfCU8/dwyIeLcZhj7tsbmuDZyi7X6mDtqZWliayN7RbdEQrV6TuM
3ZQRrKvxM0nydH4Zf2mr67o9NGrwWAljFHclRBNbGkBsat59rEYMUSe8HSSj
Zau+UQp0y5sp+1EyvQSbtHwoath6zaxr4lFlfPUmzRKSmIsbibVkXr8Ziwx+
bdJsSfwSA5qDe8IiHdLc4aWfwmeSEILKDnbLo4DKo+WLOl8+SO0L8IrnxHJs
fTrJ72rK8g/feZwg3OTOPX/XV6eu8V8JhATHDs+244C3vGuF2fUiKZW+It04
GIoLUgrfZcVSMBltQEd1xq/cGs0kBJx+39AmSywFzYp1sAZl4MfPpBl/Z1/y
YsAlwmkTIkwQgQ+B2tZOmSrpvOmoV+EL7bMcAdmMUoQO0nvjGux64pQFYJP2
W7s3oHbLCYlh3ey1jxOqgg0jWALtwSQOj+OYFZWC/HhUN2OgJumFZ3Jl054n
xq7E6dBaFBZqTjadAGjmGbTrSzt2vdQD99OZRTWRo8huWwIeI8+SHHAstO8h
sQRsRHPHzYobSS7SjELP0SnQzf61noERtCVFtCAKaQa80enUq7iOjDNpYaD5
pJuLpWXRK8IHxHyvlrbu2biQhKB+b3SVFbabB7mrwA5x2Dun9qOouhDCrZql
hIHUsc7ReHv7cvgDnS7IRIOndWnuHP+C6IJTgbVFGqshUKcdOVSx1rqMvaGD
jhQCQPZnLQTcz2jl61VL7uJ8QcRU9A7/ILOON5xJsOMcWhluXIE+jAaj9CMk
yVlN/9f1VFIP6R1gIpR76WntewpC1mnbOI0RrhPco2HdKZFIcX9eKmlKiT2a
+rHBdlOAFlvT+ydTmBvrrp1+1vgWjDvnxqkspxBG3wDG/LtcBSd/qCC/Uz0o
LD/u51i2mweYFi96GJUPI/NGkJ+ghZG+dJ2YWkFXR3+u2TkEhopv/1cOXiJz
1wkb7Qqg6D/wOopZOCT8D/NEykZqgKL1HjWocwrfd9ExH+ZnKMcgJD+kmMXu
I+w4Zv1L7gl9zffKMUh5YFEQo/twzj/beW3kYxmaWlQWLaqHKxbKaBCwlKd+
mFvvQRZYGQ2PwqF4PUl3Gab+5tPgIl+CLG2yxq/XsBnngr/dEhcDXLW7V19o
4nJuZ0bPvHsDOQg6w4eVrEY7C/9L1MfARcBE2PN/uJWtydCfa8BEq2V2Dyy0
JwTI6EGdY4mUIfXhL5mFBGjrpoVGh/UO1BXPpxmgh/dAuyEdZDnqIHjyaIFP
srsnXS3vtuvWQpujwhGlItyc26Yqri9aZPXbz/XRL4cTVshpTSbi4Uw3yP4I
IpxnnMsdfK7VfkfpTSpMG2vnnA+Se4bbCQSc/6Zg3Z6cTWhkBGk2HK8RMqTW
HnwxtZxgkPxLa1h3tfJMfBuzMkAw0n3gd4lQd2d4fnzBWvAEw4lBTUm/lMCR
i4/MrmjP1ciE+egFOJaLt7ZCDrzS9FJlCnmrTp6d9iKr+2uP9JNyRc70c/J0
Pftvu6c7Hra9iK5RsczUX13Pq3zMDcRZuit/nmxenp/hGODAQPqLvlxF8M1E
kC2Axd5iPwtq5u8UGZKYcJKkatfJXPTqg9Etj7Y41aeHk9eopBwSr9CGUUd8
xB0agcIVaWVcnU+RCJLaAixUV1ZaLHufRoDnad0nddt3gpU3XUHl5LLZHqKA
PA0s+XwRRWXKuJFrOLcBX1oxtOexral2FfahopEYFkdPtnBszMJ40xly7huu
suLn+H+kN5rWy2HgbXPEMqstLDYjwgV46lDQaIBiLWQ5w4Zl/2hmPhkZ/Bho
+E7kSujjVnL8BFP3wA0/uRB689tMqk9Co1kqJPkeX4rr6fuRj6RNBh5onY9+
6an+CI4Ch17BZI1ukWU5NB8PEOfWb9XS1huM53j/41oTBeBD4bViMObRzxvO
zl8DM+UmGhAtx7D7+ON298bpxv5c+z5aAJJW8Cp70VxAju6hdNmxyxNfCmx2
HLNz/X+wq0TOk0Zm0/uSJxMKvVntWzCK7+W8I1b0JMV/ZF2ayTj9vBqrIADX
q3EswW7bFc6lAy3Ie3nSltjrbqlkulNK3XtoTm2J1oAw60vpiNXDGlb8EpBI
uIuzThKQa1OY9QQOdTQbirVqVGyoCD/OS29WF4Clfzqyol1F+BvETbNxUdzA
Ea6VfDORzK2v1NRgHy7PP2dkHLGhoPCTOpE1K6Ej5VW4T2pi0494XUBKOgIu
OMFVSvIO0h0ao+Iv5eSa9juoj0wy0tjfAMr+GpfpTsL+5YzF5EuP3hInoPc9
W9P7GsOc5RcVIliswc1T+uLpa3xuZchlPA4LA8LmT6WPMch49wLk4TgcY+Vo
Vy0smFw9MQbo8JESsGqCJZgt5FEjhLShoxk/z0q0c7k3n07Kx4Bca7Ppbmlk
DdSJI4WvL93+Q8zIklAtIorZd3vKdMFOE8WHJctxNLyJZTJ27pl4ZAas8D9Z
XvnFNJXZl9hrInCP1MbH29W6m/kAanqCF/FG/AzuFjF8yESi6SOK7AFMpF2z
uzJcvVqx2B59v3HYlgWTHTEpR8UbJd/EO4JEXyo701d/eHJlF5aiq1K2S/mx
7sL7OdNBxr7VG4l6qze00lkW/81w2rRVEm008YI50DaFlVGQcOxrx78Szm+4
RGULptpGjqssL+50+itGYioGXMjRT+e42JgNljPlO4Z30kH/ciRDTgoI/fFL
aU4Dnz8o/BA9XQSW5fe1JfaPVYTvnyRT7kaEUgQtD5WKoqTyQI74q5DA8Pr1
nCf+LFePdkTZV0Am4dQARZ64jsqURUBNQBuIMm9iYMZiVI8k7S0ULS0bbh4q
ClXN+nJ596aY+LfvCuC2Lsny6T4njz9v7+iY3oalZPD2S7papDp6Bw2M2Nh4
G+A8VA+iHGWyHC4vVliWczzfpQFu4HQ9P7vJ3w6lfvt4WDj9PRdwd8Ct+UIK
+fRWQCA/P2+S/W0DUc4fdVqkzMbZ2TqoP4fYk4jqx1AtSfHUDs8VBhs0EIee
IV9hlknbnb+aDhOdVodmLwYFRXA5VY3bw0KSdeR8AATyYR1qxFL0pUwzupDQ
7CkG0r0Pv6Pvv8DgX19F/vKGV+pnMi4BxtsqOgy2VfY3mqGK7Q2RMvB+Cuo9
vfYbnMmOMF4fECxokvzCODxIc54sU+eRw/LWdMeThHdpP/GuxmBLQPIaupyc
kH8dyO/3liw97cJFHEIR1tAK7jlc6COfSj24rxAGJ8tEh1giuB+/p65xOvXP
+5dONR0xS6HOIrhTZAMgXXea1QAEA22EeXJ+Hfg+l80N9y7gcJut7kQ+Itfc
zJ6FrUtmhMKf6MXg5Sd7BnJt3nt2byMR4iNydm8x0JbYT+gRhWIWCAKgwjYW
SztMEKf2PJ82g0fRe3tneMxYgQj7GB/eF1T5SRWDjrLHWEhqrVzYi6A1rv0N
g90csqQUq/a5D3XafJglm7N61MgLVmNbcwEWmUZj3gKhEyBabeknGG7N0IDd
CaMHg2S44ua+Rhib5HP7KCEiSJHE9WKQoqNWCNTDTPTHn3pN+J6cc2NDC94G
TqwwLl+17aowq2DM1QMJ05IMNVxfbItBZ8JAxGXPjGuxtSGfa02P/YfeuIEH
/kOsqU/4FjaGD8NS9LJ7gUyhNaPMDHSzK9SGR/MKX9srsUBMeqPx32w+6/+Q
uWoKiBWrmikzdL0KvFG6eIFFHeRl9xATidZu/zZmF5a/kxyW+G7b79maLHl1
HGRVffQLk/FVVzd9zcYtZNSxgygJD5lfqdN9Q6mTFM54QrgeDFtnr/D/4Y7B
NcO3wELidQVxv+RFTI6Be/4ZHBV46j4ZeiqxxEAKCj1Wc6HfcHVVk3QxCMpu
pU1EwG6+xLMQ5Jf7tO9tgDew6plmTDzGOX7RpqgnHrl8nowC4F97mnPM7re+
1GsVCkVde61pHVIp0+DgaZDJ/dhO0gTJdjDajg6SQMKvvZvg38h41E0l0XMU
SMIfqQ6twIRg/6zECjEeFod45LeWUR1gtA1Ewi314ssSN4OL+z9oHGKNbz2b
F16PfwzAsacSA0oQfbaZpgJvA4RRdPbTqGOyeK+32wPAWgi8ABIakced+5Kq
IS9C/YbSeheLvfNl++ok5Hs/GikfossAj0CQioEJMDixAcUCykon+oWTEh44
8238xX6E9CHFXJZz1q6peMyQW5eHGmNm6kKZYij9OtaKQqtsreLPZa9oT5Vs
D/en10gW2eqbTCYy6DJfEooSEN9wlCePha82U6gm6dd3YLA8bBfwzkst54nh
Y+2gOvS75BOFyIOHPbeUDTcRY8GM3yQLfFMuzEwk4NOXSY02PikBKVx5dhKp
pl2y8wGc6fTunfwn32+PPa/73x+amovkXh4KbySQKL9UYkZlEhmQRGEerKDb
WoNU6C7aAQezi7XRkBi+UObLlYJGfngmgBfCgTflZA8ab80PPhyAS2c5bAzA
F1bEjTkSWbTZa1sxB27o9mJGg9kJ2J+cTrhrvGJDpqhBZhic0EWaTO6H+hxq
iSYnnDjLCrnxA3Wo+FoZNSN/bXrrGVfpjMtiFHISUokazfvL6rrZX7cS3EZ/
f1llvfhZwAR6u9xQPQXnC4Er6OaR6QkFPG36Vkq+0bwGJvGHAFWaUc/54R4x
QcT2M/K3hfQ2M7jnG29qCaKtSQ46hB+mGiA5Wvlcw7H1zgPHvQOfMrKSUSq6
AkXHv0wLp3UAu3IXsfdNxCzvxnWdD8t5ZOmUCRv3u8M7SiMN3Y/6NugeqMK8
9i1oT8LJq3n83TE9j44TzewPGYrLC5YkYYjV6M/DzysBu29JoRn0B1b0MA6S
kcLnxZL8G3+F2g/WtLK9FmQYr/gXSiowwsgBcGOBAG0rNkk6xO1R02wuegh5
CZ91ZeP6zgCgTYIlWfXJvlFuy234cy1uPypKAivsEBZMDvrEe7VRBopyjnf/
TFf+oiMf83L7QNnck1wZJ7mrrUvOr3kB4GN36zsQ4tjKukvwHZrFExrp6e/3
PTPZlaiRdDCCFkUmKGMW6m6kG6RM0NtJcTFNfwAPE5blkin8ZrnkOJ6k85ZQ
hkktSpTQU9o3sEWLNIq7dZBBzGX0MOfzMn7j2O+QuuyOXNzSS5EDLqQmg/Ee
QmphAB+EoAnxTRU1Oyh1OGPEpMPDKP/k+HVJmEMa+iUFNmAgpTk56nLMaMFX
/F4Ms/oX8z1pMzRYQOQTf6fVA8FFB0DLpQRlf5D+RrF91gkKmXRiwKgNQwDK
Hy1n/uxODh78qTNpJ7ZO9EIhwrB3aoDvnjQmD2GR+bxDj/O5JmLFx/Eeyjqu
J5D87NljgpLWJjKZ2vTPiihAReS4UmvXyq7LBEQ8Lh+6kcdcek7avoobH6Jx
Fz6XfXuEvI+R6EelFyYGsxpDtl/4joaE6DJ9cWLyrFePvRj3Wjo3glTl3qC9
nFQ6q1pqwXI27wQyJTV3BTXfekxs+mR8qkWIXpBEZDWvab39z+ov64VC9jb2
j0muFZQ6b5LHl8WAUqLtibqLP5m+qPZOCOJ/4/vU73m4i3xBHmfl7QrwwDhR
1u6/MVVk2qRpMcYA1xiVKAV+H5ysEJW0AFBeB47UYvs5Rdxufs0CJOgcobhW
PkZu68Y0b/EcB1rpvbLA1mwyPwa9BTGcvgDDbfd7a0FKgPqXL8Audubf0yaz
APONATHGKsJG0omtEPU62GNUuB1Gx3dKaluXkWuCOpBtxhEpMQllIUjVWcJS
TeRjS38l10IvSPojSl90Vfal70O4zRmhldgv+imfiLUQVCXTAFefkC53yeBi
jKByMQE6pJv00kWKh/bUUUJxpTDzwe33lzd4NeWQVNg9qv2rDJWzncigRgCo
dlY/gJswtGYtNWZbNZgt4wLTPwcdN7wm8ZkUEmXpE9gsx6aO0uSTkc78NIcN
JL52tRHZSsqEWay3tpv0UfgGTlPEc3H5Kvl2VDxI/ogr6PpsSkuvBaeaTEY7
JuAv8i3OXcZAtiXmIPFaW1Bg5qgLLHcOke59c29B2q9gOY4OT7gkdUE4O4MG
fqYJlwm84NEBsZKH+uT96XhXM/wkV9oIHte3gHZmhiZXE3z+rjnrY7majTsI
R8LNO1e8TtF5HZU+RHyQ4Uh0QdQ3Q18WB5F395Vi+44o5qUmi4hwBUGOXElL
PU9ZIZZz9xUdi9CjdxLFoQcCT39WPVT180HM5rngRGF0kEgIVvd84/c2HHR0
onAUjdzER0nNTq0uEH4AgleaAm1ncZh3orZCjrsX5E5tlvncpR6unQAjnkKA
AaDquvvBI/uEy+jcnWjR35ujH4Mpn7fwCshnjID4b+oaRQavp5PBHcNNy7Co
T01daYakgiNPPbEvSI24n0khbvyazQFcPhxhPH+e3PCo04rUa+bCK89ygS7b
sSvRftLuEx0NxrVB+EeTGREmnCYSacUJe+VzSE6ai93zj4Po2dw/MyhsbM4+
MumwnPPLFOJhwXhZTOFc9Jj2uFSxnZiszhA9bfhNF49G3aQ2L9OK6k74qd07
ULkAMIrVdluDxfQ90j++WTWuIp9b3DD3nE1OpJcGnhmHxRcwlByKZj6gED7g
zX+3EtaJyx8HFWUTBAJk9/YWaIKMHctdRN3GbSbPMkjZLnEhOgQNVovncsjk
Nhh1uSXp7uCsasL4+Hs2AjEgacyynBkjXGtCuEAwEtVhmuaXoHJK2kF28ogk
emknvUOlYO7LO3ovppoGRUoRktt5prljevRqPOX1ezPRDLEX+ablu0piJ0Ya
pm72zvxEp6nnU+rmzRfsmkk8OF6ImUMhP8UjbfMK3PDMS9dHSmxZZ3nNweAK
4sU4KaHaS7W0837Q+VcEu9R6GQ61XZNgUb6+GjKs6+9qxWx1NgZJkaqAn0vU
s8NczVljVf/I24ItPrH5Eq/fjLsFRSVp3WL47KsSG4mwoAktFQpMBRO3rbZI
YQG+BXVSDXhMs8z3Y/R5l2tKU7EQVWh1YNgVlP7S8El916g6uz9hZyYlSn/v
kposeE7SCUq9gdgR86erI+d/jSuCHtuEda7POUvESpPg9PIHu29vkxMFTpw7
vFn3EFigEgjdPLQ4Qwl0u2iwneRtHgtdp8z/cB6hNuflp2cDabUxCekH4Y5c
Zk07xtCClXQBg9uGreWolC6NXk8VfpJpHUBNys4SqDJ1VoDnkGcY7Cds4kIz
BAK1Xaivmb1pOcX0+1mmE/5YBdtmlcZZ3ay5CYOqLB564SD/0GeYAlUq/Je+
M7jUglYxldYhRetUmwZ1LAGTPvPM3RK65KzX8YgEvfPk9WF27nBzaEQW4Gtr
PjqGJR/0vO1Fp42r+F2C7V3ee4TYYlsZ0DtYBeBNV9yOfv4bPPExSIG78k6W
N2dIwzU/I+malPkfyoI3/XjEIao1or3JNf26XhiGXKfImcwiHxmjCBNYxQ2/
ciZfKqa6lXsvLLeiTiZ/Y7qzheZLUQf3rcd8ng9gAdB6zp6g1l9Ir9R6mAvU
IiXRHQwAc9rbE2iWK2th0/1ApUyRrB8/Pn9ArNVwb+wzqYB3REZlP815a4fQ
PaePuOLjGYUG0G1YHuIhEMdN+ZS1hAsaCV83qDSILB4qltnR7p+NipG2XzbH
sDcYQeuacuk7Bs7YpHHBbJKeu1QkTJy4OPIzWk2wPbAvXT12FoORE7uPmHKE
6TLMhn9fASlqFhkSf/hIAQvZWoKjxH8GUK3RMrV6P83m4DkB1iOiXBHMbd0+
z9tKVue9lnoFuOiJw9k/KwGOUR8eIQHhWifkXKozAYJcaTiFtqQo+Js7g5O1
P7E2JKC/V+Rcoe/otNhr5wWyljVPY1ePqGaIxSJXxtuuIPMsggN1+QL9MSRQ
l0Y1JgCMB8lzpAQwyRCWtKYYB3H7qRXASIyZTLLnVPdraZYqu/9KH9bBp1hr
GAf1kSBmvHqfH0O4maZIGDOt2HjLcPlp/DDFtCCvneHEBlz9q3d5lKB+T4lt
3smksiyHc1kK9SzzyDr/kh62h4Dw8alPBcZ26yrVSUGbiEnhr04gHFvUDRS7
0NDq3KukI0MTOJvZvtyu3aKhs34C6yHyamF63AJU5HER+YHf/MfwsBwsLpk1
kLr6QkbtO6LP54bR5Lm6B2WuXhgZ02EGyeYXOyZQQ4V7l0a+d9Mp3riwDUNh
DRWe+MBz+qUFQuLbTPnr3YK9My8azgwCtAT6uJF8W20geiWsmM6Q1NxNBA+P
Obun7Brg/3KHSTJ1iZHaZ2pZlIImNJ31CRLBSMW8CMhk0Gt7dI/2ju8Fef1d
97vNJRsE0FcO2AoWCsRQ6YWXnS2i1Jco7uaTwyxQdTzua5Ckz4JR4gDa8Zem
WoQuZaJJrdVkUo9665v0v0HkKFQO8Y2l73epbyOUMJafcnGIvEC8cz9PHCVJ
HYlcuTS0LE/aarLEBjgWiKjkgAd0ZtYt6IWknnRwbz7DhjDC2wMDYTNW6ysW
nf12YXXF/bRjSGnFxhnFFHSyKpGAJC86z6uEK8pvg06fgD208zprsMeI9Kae
llYyk0uf70I4zKMLKqRYlWVdFTS6TxWxvtfN33Wa6RFHvnmoO3skr3y3VZFE
xeBcFDzxGTPTOhfO5PmlVZnkJPl8TlKKXoFEfMRuKIcIMHUafaeWlio8B12k
P5Nd5N/WsKLtnI2IwEJ0BKfGjuK6m7UhjfYkJ3hGbT/xvYm5Kqzc/i+vO1gM
RNeV3zA3vl56/ZZthyNzRFWfWMsTGmvqWqpORLkFvaDnSBJliA9wAadfXYjl
BqPXW6NeSt/kWnKYjLlHJVZG6HuwG8Kxx/AwD/pDVF0d2AcTtFGfQgsMys6j
b+e4Om6KBCaySPbwMDdk8YRZRKrA2viyyEuFkXwb4tE8qB5nrgKUTDulGSt1
QjqTaRbEM0gjRLDiqV+3NTiJl8b9NQoAxbfnxp6cmOZPKRigvuFgESSaL7dp
YY2Iiz3+ysjGVI1Py7o1yICQChz0QI/VctCQT9Bub2wAikY5XP/piDA7nFIS
PrGzuzL4hT2N0BR4Qku9n7fvTHtk4Bf6INd+lGNlw/GiFHubZ7CK6GRXBXgA
o4YvDdzfy8S9S8il1Xa5NljD0xGpsXLxdDvmEM0kZ7Zeb8UvTrwZg/DeFJxr
goAq7a/vPnwovjgkeaviVPJvkOuMkH9tn4u7TQIMtXgTy4bjxWdyOuJ5mthk
nlMkauVOayKORUv/yZffMJ7qSKDm9j8dk3gMtGLta1jZpzd7h5/x4mMU9Uzw
dN3SPX8gdawX51Ngbt54ZagWyU1bBe021LR81/nB/i3oYfrxUnprc+ZkKNE+
L+Wi1zeCKM5tqISNXhmRntHIjjCjoI6m169KYrpIhJRwSEk6mZ+6skfq/PO1
CWXJ4vEMviWVQ6+kMkGh8CMPnP7Ap2FhyFaWtPbwSdwgQ+0EzLGOBM1F1lCk
ApfEU4ni3ANCLH/83ekpNdr3/K2qFsQG20eA5A0+6jM3g0pEdQ4NxmY8G8RJ
tMt46bXKQHOO3mPyEVh73GbQzAGsC2uqifQp9gmEDSTaJomy+BBFIAGNTRO5
OXKQgw57Rrv3UBw8fSpOJ3UnW9TDaYWmh+gJaO7U4KV0z7cabqW4NrdbSubt
Eo/RI7DmfCmHKctd5ArhXVGMFiJXyAOcPghOBcflk7uHPzITuPEyK+AyALdn
IbSDXjCPYbedhW4+UYKN0ogbRuhE1IXzNNZPjEGh9VguMdBTNZVg9GXjUzLp
9vc5o6UTmFZJY4Y4LncAQAW+5Ie+evh9qogL5T11ejUZD9xyTNVcTfD8P2xa
mlwwDbaYeS9EfJ9PSMQUFQvqe8XgrnmgOhySWCmW2aatnvWjbAm66MCxvE8e
2eCJSoRuZJaog8qPk1P3JzfXoMfHV+BSe4YjRRvIutxjfuPoeOf8ZyGW2Xyl
BaKcaRyqPzaI96yns8ZJXbEAbB5GUefYXNxAGO6NlMVCjsKvllZq9qBgfRZy
DxbDKss+TCI0SImfoby9BEhVcbrzYLFzTONDNFnbZbJ91wRHGCJVUH0Wz20g
4+tCOoTSHOdsp6M1bCRqLN33Y9tji5MAXKRgBbgfwT8P83y5ACx+r5Rv/WQf
S3mqk0xs1HZGdK3XZVSSpoOzA/Ar/YnBwxxHquqNEwbPhRad/P7Xle6GAYVu
Hr5kUxTCWUGavf1Cvx3Nt4YNs9M3CZEPraK+O0ZFTkSH83a4WQi75/8aD55V
tddh2W/WWAtYnah9IILLHgUMpu/l0sBnSo5DbzHuBaIYh6OxQnBdItiboumB
xVFf0L0471BeRbn7e4921HK/kyr+2dbxK/d8PPBUe1vXWyYffEc//cBzaZ1q
I3ouNfMsB5f1qEgp8mE6IaQJch21SJNTrMyPGKmVipdEu3zqvaFVaRWGxnPa
HZGPhp5lrB54GSHZrJZyGKtU6bhrDIh4REbm6oZ03wmfY6BIiuGc1v3Oikl9
Eo4eCSKzBC3yxB7hQBZwXC8dETdfT6GIzqL4F3bWxUVWWFZZOskFZdvCs7GB
0aY3gPgeavRNCGKRNsqMTjB6INJDuzEOYCrKBv+k/Ghn6zzf9OVzuZjgokqk
srgaep+bok+Rs0dnJtPHJAoHjk2GNfVWaLh5uM6OQEOWQ/GscejGj5fmnTjs
kcj93gq9ny0px9sVuXgX/2GjvyMJC3MvkiuXuULhgz63nz6PzqgD53QgbWBB
tLC4/c81fY1TUsfwOG7HrbHnEi0K+mm7Wg5aAHHOFH6TMMZc7y5iYJnZMX7E
3KZ2+h/6PmVuszdixsBLDcIRvgKAO6ZfYcMJ23aW6k9XHpHBBynvXHIal9Fv
GFVS4A/KMCzjh+Rs/OXqn7UTecVwJPR1AH2OyRt9B9GI1dkrSmr0xEZ+tc8c
55teOj0VfHYCw1sc6r0j+fwunw810DdJwNrXkE7AWaob+Z09BKYSnLyGWoQ2
9xj+Os2Pw7Yp0gFtvfFSns4Qv/IXt/vY0Yee6veBH6nR0vxinECa5ZbXRuP6
5OQSgBy0Z29GY2I3BZuo6FCmmitq6Js0zngEPTZA2cW8GMLlWgojyUaqU02g
KiFGJnWvLgaj74D4u8D9xBaJyZispIYztlSrLruXc6WtnKFOvbrVJtEEQxcR
glKuLjJLGVUCjrxfHIqy+jmVPtdHZpomBvlMkxZw7c8uJF1BN8ZXA4motkD2
67B3JY0mtOU5cKaTH9CM0IxQELz8JzETcVbDz8q4/6/PjeL8LVp7xM+ewQ9o
9M/ROR+luT1AMBXf2cTWsuWBCzXz8RNq+f5ONpthE8kvy3ic3oneTDsXpwco
j0MuwY0+zVl8DEcT2t75Y06u1ZabBRF2lzoDz3blDPNyYi5RRnOD6TYM7E9g
RU1tf3w/wFhu/89thdsHxvgkQrdadT/sfUP0vklmt09JrnW5DuW7oifSqHH4
Gtcut4T/l4WG0qmRXYtweRb4yRtjWB1x3Kb9HqMlXH0suYSDkcVe+4BWcyDQ
t+DGtcQez1l3fyfKNiuWsmzoAXpMMklt7AuQPY/bRPDPOIbE7DPMLN00Rxs6
6VpO27+Mgg2ZMlNo69tcr6hQA8TOaDDV36x1M+c/yT/dGkh7Vrk5tH+/NGcU
hQs0K63qjFUVp6GZWEmosZ0z/xXFHkWyR+SHyFAwSA4vjVv99314tOwhZF1S
KarIEE3H4Sqsvc3zytxZHQYTyM8sIKgvo8moglIBKE8wsFoibl2H+YBU1KCs
81ictBkki/gS01TyTwzErMBwTZEiimVrte7CEOPlnW/rRCOzqN445X3eyiGp
FuoulTS++SBCd+GBDdzs1HJvMxd97+G/yAt5Cli/ttFq2WFmTdHqa1WF7TEr
5Z5YAsho2Ub927BEADidwMCiF8/z+n8h8HPQ/Jo0jlFLk43JeCjukezVPm3f
yZdW2G5PHAkkSa7G5dNudh3Ij6IW4VSnm38ydnVnIihuc4SYDSU/JMKKS8o/
TU0KlbVYfhbUP/Qyr9vy1TCwWjbiHEdUn6w55Qhe00DIjUHfN6DYujWwf7ze
L+ElxZf2XH9U5l/4lASOKUvaBoTFyd1t4XIJCMsfo59SPKX2IiD13ZGmF+KB
N6EiLzwCav1/j8SvsdmZC4ASyvfySOY+PND388MarDDtW1fwhvgKsvr0XGEU
t/jANO1EKg0rynzBNC31IvI7+nKDxX05IzUlOHTH13pPucPzilL2/1TRq1jq
A7cvvD+KBtsIm3RkleeGqydS+lmWbAVt+SHATbNXsKb2ZpHd3VwOY/ILWWYY
dj0xcAPnVlWprbw/BnvOxqE70wqm6Ju5CTcG/xrHAPATgGEf0a++J0/a4JYM
iWOD3ou68nox5JuuXshnnTGjvTRTcJwehln2EobQ/THBLjHqrNMkNKuAo+pq
iHyeCDX+ZObyhmPsrs9z81EOvwEBpo2ZeFo3fN3rCGL4J4PkeN+FFRsa5g5v
scc72p+oDTRSnOK86gJyde0N5RVk05uNgEdt2FdegY0KoMvo9zxS/f65qEqo
jOZhU3yMXxxVk8eEsWbHvxco6KNnQukrjS0mYTkN1VAwgmuDeLcsegbeWeqW
3EKxBsF1ZqqxNJYxQoHd8OWggjs0110P+RXJfSWsDTVxHdAtlg5QCI1E4jqZ
lirl2U2wa5cXf3+9xcQfCIyOh7lK8Zr17Jr9OcTuS1VMroq2MHuyic930NW/
NX4Z//BzqHS6VEt9v+DeE6clCavljYPANrmLa54598JvMvfcLDLasIG/e4bn
9COBswym/H2Eoh6eJIgTJaaSs0WKiGnQPLacDcgMcY+wueGPi3iNWV0S/QMz
sfIRohTx7pmGWaJdEJGoGMOXAbhnRySyX87vxfplka+sOKXuFe4nv3H3Uj6P
6ctCdrtc2olsq3szcvdCHdZ4klVYbPcOcZDjAULLss/IekuSOC4fM5tq38JT
0gGWavNUNIlfo9BQYHWZwgFtslkQO6C60ss3ODnCKdOaLy0TMhp+Bh3RHtBs
mR1m2KCLYPRJaW7+cD7UybOg6g4fkAmd90eTjz5baEyTuVaH8ktDKnSJNodf
B6qS6lmSwtbIJZ/VUg2ihzk+VPx4vP53PkMocEqiCgPRN9DhHPQ5mN871k20
l+WBsw4sHCFEOazG2gUlO9dWFu1XzEWlGw0iDCQEl3YRES5PCaUDPJrK5yIC
vSewtxeBwoYawosgrmnAXGE54Dnmp/YxcDiR9sMQMmbisNFtZPhPuy/46AsC
KLxs329aapRCYhCwAjJS+rYjqtbx9NSwXx7WWNW/uoPRG9oB+IiwHNoXsptL
YVFFFMZk6g2FviFp9C/7GwRkXEE45P+b9AV9IWKr/orDU9WdCOQtKFruWJLg
L6Dgx7JoyasVQNNkeor/y+n9EYsBHqBft3dF88Fd9zU9VBh2pP3pKLTjs/2m
4R1WcZ8aZ2nkAO+bn+RgfJqan0/11RW0rl/7moxwL2JPx+7+tcqUYTz4UUP6
oNXarmiYIABGIeSEoktvWwEP1eG6WizImFRqacxdj/tIHKve2b83K9OLMiTy
g2LRWqmjOIIY39Swg1GTl5o/qvlQR7L5Fvanp50cERFV51tYZEUhN9SQycIp
TeQ7b53mBEz8Kp9RG8RwzWPYkegtemKhzF5jP+1EZnXLzD6Cd7Sgs0IRNKDk
mwiY4/+tSth587utBN12JIzsAZg1aZ/20oOqOjY9NxpiwM/DtCgERiyHBTE7
19Dwuv1qynNl8jkedk0M+TNHTWF+CajDTpvoDm9eT4I1epnH1TAUMAR5gGNe
h5oQvoWunbPj94bzVk/xxBKx0jv/tCt8KmFV2J5hQbnfWab7khOS9GFZt2cs
lTUav+/YXNN6OAUrdelT0azX5jaCXpRlkoZSIul3dy5ToKt4etMJRzwm3Yeq
J3Jq7T2fHcpAiGSsQofu4scUDR3lSVExfcF5BYjc9seUterJ6m/gKeNxuxh8
fXkP7oM9tK747REwBvjJrf9oVOP/EzxCmOXqC45zM/SU5BQNdmGm+3VVdsuw
YiLLS5XvjnXnCOLID0cRPfTUYqwkpokUNFFAN6ecv32YrrqI56Rhq6F9xyrq
G1GK9P1XoSBo+mEoLo0OS/qvEcXppvICxjYfqWMqhJkfhsqc9k+PXLWlXebB
rFH3xS3zZwXdveBDwaj/Jp73dm/aE2YOhpq+/H1pXEYXTmCMqa+apYdYeOBv
bBr/fJV5L2AfWkObwxFyP8QJe81//pKzS9999TpYIAuhh4w5YPVtau+2RnvZ
gdPF/luIwbxjSBKUMRN0Ms45Qy2MyigrR+wRn0cAkmxpDOUMCr6yV/ieA+WX
uh0FpS8ggEJ8ok0kSXm/c3iwWdWa8PIyleTVS2ZqRL5T69rulfaw28v1rwrK
uj5sjaZAE0DZAe9FTwlTgruGwd8KNVH/CGIGzl+jcgB3X19wLyaGOaqLGrmq
bVgG7h918NlowkJOsBguArik4pTMWi9WRGRgKvEFz/pXVZ34op/oSs+UfuGD
s0+338BQzj0oBayAKTN7JziDLvJZDAZCx+njog2EPaHkm+4OHyPwfZPGB+rt
OaxYPZpLwUtwc0++SuAKTKBXg8XH39/Piry6iZ1xvqrXZn7TgryysmdWRckj
FDhik+0wM5uTiUXLE+45E/DR5tzwD9DRMDekXiJ12aUIJ2x1uXvUIWWA5Iat
KCGhW2d3HsYHgGzU4DobqP3TxjGOxrzys72o4ype26sorR3/nkhwHuckwado
olGKClRxdcIT+IWI9Ew0xvUMjr7Qd51SaGBUEP2XblBFT6O+orBcJiwt5YH4
HqHs67ip8HJzT9JCbrEXnKyA2ViMeXaEOdlfr4rmDwQBHeJAi9IrIT1+DxQ+
fAPA6C7QSZamqpl/AuSN3Fe1zUyQ8Zj0dFD7fKE9bVA57oZP1znfYJskkexH
FPLM0CROjfyBGelecs8Gn/gZN8adKLZy8vpl6klNTHK1kUBrWuy3G4T0nHKJ
CtWmU4vdiBehOs51WH4RixhKV/mXoUl/K17QbXxfhV5UcIH50tUF32n4aeGm
t6ueO92PgpxpCztvkKCfCuzGyvZPTQC+/Y5Wcv8PkuYribxJIUxdye2bXDbI
fnH5jYRrDsy/P3sz3UfcDLkNxEG7BG3Cy/x2m3NXOOQUz4Fm+tTjmv/EHHAQ
YoYUY8CIywJjrCv8TMaqqQEYg+X0TDfI9nBA6+xc2YYJzsWJ66ja7oZ5q6Cn
Lp+H22+X1mjf+qeKai03p62Tqgzv6yrw9bTRNyVj2hrUHRZBeoHeh5DSmWs/
4ssJLldrD7EXlhuc54STquKqh+irhxSZI0qOf8qRrCFu357ohWWODYCnaoUN
z8lVOOXYwNx3B94mKv7JnaIuTxUoQj0ehKDBKsI4uB5eeFh/I5Dag3fLWwxa
En9TUNyDqDGFZSh4WgOby1FT2OtXxtuz/a1HzQBzyRZZbfNl648lbTeBaHWY
YKgX6PxOXq3wskj5oWJbPtA/4gY2wA4GS8HG9JR5x/JpPZy5k9z0Oz95SvAq
ka6isUJA20PoVg/46P4qLPvmwj+yAf7b+c4e4nYsUDDbHMPmuV1AjhpVuGpl
lUOEqpwpqA2hEDHUlnpTvFysk1wKM4rG8P9H1B6T9lbrInlLykZsjCQ1rAx+
51bH0NrFRUmrZ6Z3QIKn5gvB4TjqEacpI2gMWUICpB3niS/ZciOiXy7GJrYh
2kBwzWy+n17DoBN3g8HfkKKXJy4Krem2Y6AB9nhBerqsqaRMOfdV1GFBduQB
S1Sizc4iQ2ckqIvxI49/glPzD4RZ+i5q/x7plmdKCtjtWmBWmzQdcEbL4+Po
C40imcA0ViPZ61qNn+UK3pTYOiHANlJk7ik47YFeKJljLoGyzO2NSHbzPGvl
oPScBRWnGKVYVQaWC2XSCKi7aIBCKD2isDVs1RbYfVsNQDMcQhQtMqeUR7aU
4RPpMu109nx5X9i3wqR4bi4UU/Z0+0yFqSEBZGmPMKUiyCCRDvqForb8M4GT
HumqmkD/8Y4hYyaIgFkIukvIGJi/PxA2cjGlNWOEMpMjFpKaYZJlRBBS8uro
vSYlxxwx9Wp9C5Vfi5sQaaC1cEcJMvioAvUVLIC5iF0HJXuTShKfHdyjp5vF
K46jcct3r0JVIgnBmPqDmRlb2KrIaFUfOyOkzQs/EP7FHVHluABJxvKGmfBX
Mu+Fqm2TMzuVAQUmD/LnLqIJCB6aZETXbqpI6jSAHuAyU7z7As/ge+oH3V4D
dW9+RB0fFUtO/IKObXUjmcWKGtuvcwovMTiJ5PHoRKVLcOU4eNmEGB6fa2mN
j9yWiOv3jXJ84oGJiSpd0EUGzVw8js8AFaK7m+JPHHTCY2CWObGUbmWRoA56
GDX2YqFuhlGhxNWvi7hu9gqTR6h7ugDhmpGZFLnzluMwlUdxOUIOGhIPC7lq
yQEkgWyzNPL+XJp4iuiVxz2Y+8UJkpKcToKgKu/vYKyYs6TQoRPiG9qKHBP+
QItVhrhP7L9AXsSQWCxOVHvayk3VqcUGLedTkSqF+yBPw4lOdEZeYwrdkx6x
I+ebq+nqZeA93JCNbCD4j+nAdVXygtBA0BjX4d9k6URGDObmENzPkOwRkXFJ
5geMXAD+Yg2mhEobuNUFUleCHxjQEzDABFf6kx3KNNN8mpcasJuOFHRhKmNs
FnsPUAJRoN4nyFoVVDJOAFRNicqZ7FUkZ5hivzMuInSWjCkRvNX282rgcmtc
oOEgsLRQFFNeuXWG5ZuxEKi6VsE7hP/Ru4TIi91mxadVykQLLmRAyW/h3Dq0
ngPo/uC/gY6NAHh59WJuVKMOndi1CLa0Cz/RlY/AjxXg2vsrXO8X5wADVhmh
w8K/EK2gGoc3yukkDdnHTIR7trDF8CZe9aNAjkaQCp/gmRXfwu+S/DXUQk4p
DE4Dj+HQzVYGmt0YKTQL/qH8HSjVrC2gu3TCZTEs3f0vgu5p3ErehqF1Trnl
2Rf8Tpu5+L1IevUA9nJTxD64uvtp78MObFtQf1pC1oey55rXQNpXxeNAXOnl
dWBKzNqFjumhpGXLPTRgojzHQroHRPI+zK0qJ+4oi29Elrkub/gGMyfuRp4o
JkUly73cGuDU5MMBBDZRE8orFpkGcFRhStK7QrX3NK2ivJhxYiB5ZbWiPvVw
llw/poRqm35bNAFMPHLmIUyxq/c8Om1/ARJ8+3qjIaq0lqr3bmYgR8o5Ugou
GS2GKNiz0tjYlm2nCNB32hAHCNrLd0WKuf+1w2o67TpBiRMYpgLZ9MWcjlvs
Yj26Ojg2qjB+W4vkuqKzyG6A64dCNd3Ixj/mGhG72qwzop8BdC4CE9KWtBt8
ZNraqIqwUkwhOnkhuR25Mfs8cihAEgi8bs1ou2XJNNMp6A5C//UQURo/x98+
KpNVGY6KFoJ1HPG8fdaQMDDhZV7gjCrqDQ8ji2rlnfcM0lM9kAHaffNp+uys
XTuM8icgt5Ehk7vO2aZkX2x9grRu1v7U+DJWkwoVngiiWpjV+miEmCLllSjw
wSTvkkdThmJPCdr3QChQQMVHUQXLpm+KHtj5VoMmqGM8selhOWcSKqEhMRlJ
IfSmPHGYdelqULELRva/Ta8OR+Yvnkh/E5DJvC1sY+GVhqxRWAsP3qV4ri1X
NVsfEyjj/AASu10ZGUscPwC5z4S+xFteaIQfTLwOrA3KxmVWzJe20KWb4irS
a35q9ky/gmAgj7H3A6GosYjVXZgOUzDNM5TcnapXlV2cJiZYnlFrCuFIWgbl
T5HQwywBkx5noStfNQUch4pLFLSNBkDLNTDP8+lcxSgwWwwjkoAySmpApQjY
/sir4WiDtoIUWefcSYSzviXFj/3LRgbHx+d/aBQ8TI5uWM18H+od8N2gVp0J
8OGfIgZ2FmUYuFTkl39luXVCFOEocAraGGxlJSiEfysZ+jl3AlQLtWFRXmYA
RwbPRsc71kXQbiZNLrBARrlyoibmLp7tYyzxQjiEHZ/88Xtfkpb+l1MdJEFO
tmaGTOqFWNXiIET3OatIHruJQWA6CfZl7YmrWiUz0jKOxH3BY7qaW71fCdw2
wI8nBxBufCQc/6IIE07W40E5gakb2HR3KiAiTv6lvbEHi0jMDdkCNWawvhKp
dU05fO9/OJsg1Erlad2RRvTK75Osi7WXKti9gCsnQmw1JznmgBHlwYCRL9Ds
Cvg5k4WZ8vxwXFkFWmRSNbuAdQFt0IZLXqVmMSN/hskUvotpBssSUdYq09sP
6dzV+wKsYY2YRp5IFtEfWAFD5Rycf3dI/q3MR0Jq/zJ3ayakW3IadpmjObew
lk8+8WCsJGH1thjA6+N69DEHK/pR76mtS9j9wzYJs2mk6G0E6ZsjZB+PC+5M
oxkbtMmRUNMeG6kH4xO8ZvuH6lrqJWfrw4UoTiw+SFlbAqqaAUyEVu70Clzm
RwNzAa+Yv/kTNhGhm6zPWzrSfVh6PX8vt57GGXlBFWSK73HkjT2oLhLZ4O17
SiufJWzK7/3O5T1F/U+Bzi1k4gmZ23F1VIdyFOnwKtjKHzCHHTwUIpAQnteA
ix7UogBEo5M6/cOhBVmOuaeQQzPcWAe1VvtIv6YL3CbAE3vIphDm/XpjUW31
4319/C+v67lcJ9PvAWPzCFMXRErRNYWnY2U/IWZC3OhXvp7ae4YpThbnHK+Z
XkIXEyifAVtbPIX3wIOBEJcZbdjaYEtwrWQ8rg977LZlDOfQCE6bE6KeOugZ
yQ+aXpBmznKnfecJ/nuxNSrA2I38R5Fi3BioDVM6WfSE2ovulwK3Q+oM32Dv
isoDOblIpBWviLjyoMPW0OEsImZjaDSorKZxtMleC9f9NjQvN8dUEM+mteVz
gyXN/12xjL18gl3zcRxQFawfYYmr5cIPAmXcx0jVBnGXbK0k51OgQ9KUXYLW
rLNNfGSImootyj0diTRL9SpBk9VJpzCgV5VgG1bGdDmU7pEnnqJ34ExkAou5
AO2Y2SimpyQlBRiJRzNHJz3IxllXHZTzosZyyA17vxnPcLxO5sculc9XSPln
3ghtu3MYjwDkkc80uFT+8o69/k2mxjVd3tt4xPxbuTCGYw3tWkXMwiXvFfeE
enllJxdQuY2cqPSpC7pbV4aj/D1/jmTBpsRoIGWHNFwc6YUKYvZpmoiUKM4I
WTyBIei9bE53J7orFoCKAelMRPM5QjVSn0udh2t+dVLg1AYOCoWVnoJsOLVX
Q8P2eYKKzUxlEo69kkC6nZ0ImPg4oSFTrTQDQj/F+ytY+9xdV3g5JVQpwpKd
C9O+7/2quAu4LgtHOamN84YNRXJbq3tAnpJEqhPdhpAR/A2ymlVfP5pFnNiv
rlmiXzB6YytRmzaAqCuT4DdJ57sZzVHAZcc9U52pwl5keMjSG53bGDZwe7il
L13zHvr0aTM5zICEMCqOOquvFVgbKcqPNN9akQRK+yUrjSK10a8oEYJrW9WM
+TK7ZSVdioE3ag6v8tTzB5L6RJ8Tz1nA0ZDX5ORpHXLaWaWFw9gol075WsUQ
eht2khGrdbTemTFdkcLUREZouhZxDFuTV+VCs5Rs24ebjigjlQlOp8Vo8FIj
pAWjOqdLHGJrEc47EytAseuPK2RnEAIfjODGWVTWndhKO14pH0vJ/rKwVQoA
Eedq/vdpmoSh7g2OhTFIOFREyOU5tDeQwrl0fTl6S0qTJ45Isa68LDaIKjaE
F100gjPTpYysA+fzxEOYqJS5PTUvJh1kl3S3avQvJ/pdm38dVJ1m/0D+ix3u
AViNIh/O0R46FRd5BIEwi0Hp4xQDCr/o6DGU6Mh3yw7XZhcDcE77sxbWtHt3
QnsyZkchoU9sZMjceAPR5xDXchSnANBRoTAdmTljAwUrClyOO1juORjqlkpm
nAR4ZwI2TAsM/LPIScI1sOUCr5dpL2+OZeW9u73jByciByNzEZP5v8cWyhjo
ZDP6R0XkFLn3+hCeUS5i8tNVXJnVpEb6MzGV1aay/ZXnqBkAB265v4rQHx+c
THNvn8gWQXFUacG/+DdOH1lr1fuqSeOIzYcmHugj7dmStlwjFVvrXupCmi42
c3Al2wMY2JMnBpm1TNXfaCRAHigRRoIcfcLrR8sl/OErjloBwIYvhdbPiHE4
3tiwyYIPXJk/6xRY65xPi6GpdNyrAjsBMGM9+QdNECYKfue9fTAYpI6b2A7W
R5IObLawmkWOFpBkdozFm1VE8YfQ+wu0NLbgDqNXBY4q1nmVVDrfkzwkmRcT
/91P+tUJpvsyD0aApeh5Jpho6/VFkGnNz2NrUKr/LR6QtgTfqsZKqVabKydD
4INAqaMqNlfRBN1bJxKzjjsoAWmYNKhZb3ELiBOernWTVTwsZ234oRVmsh2B
0q1+pFXkMS0uM87LbE+e9WLU6su3Dski6qyzS4/i9cxah76DDghSKt4BbRry
0jLLsab7LgS0MzdxHmXO9+ynNIRR6WYUkNoYMvsQt+DNzf1oBRawz7v1Sx1u
34jx86OXrTzsZ5jQWVm5WacCXXP1ivXFd/F/vRsg4W/C8Xwm/ZtLTZd1v9P2
rdyakzAQ7QX2fy/0FLJmA9c0BvRboFDunQ1hGDseZpV1+5JXq8I9zJgbw3fb
8+sDLkBC73dMWfLrpa7uMv6kcQKFE9956Tc3uhF+0B4tmpJp5OkgcZhWl6g4
Xybk6HsKEmOc4i37jEIfhsgt2SsCtfOOAwZdXVS+ZHG1KW8VnI68xlfYSULe
ukksOd7O3KYWPq49nAVIPqfr9/dyjSAAd+Ea6iTySEzt8wN2AS0NriTHfb+h
NtuXfZ8TYnQvgokoJ+4ElO0EIPUDAnqiZGSHr6EchBVX+6IG3CcE8I/WFyHo
w3SU78A2S6sG0Q/wpENQXgXsxd56VsaSRpaPQPb6l02PA4IAGs6JKHjfa62t
63ly+VRN7AYcna7XxvnFQX9A1PmBh4RwhOe4GQQPgb/ghtKMwpszuiR66sUT
KhihevGpdp2HOnXvi0/KppC6ZkqykUGpIRUWmcbMt9CnZNSCqG2MFhY5or4O
Bmr5LiX47LyrPUf9ou03xnSORUDsyJq1Uw8Y3QneKlcXLFE0D4h4VX24GGUA
D7PDCQfyogJkL9Iiobz36VjP7+mUIHM/yQoX1XckuJD7gUukapsogfjGlUhX
fKTnciEV1+PKAwx+PYh1MFl1qu6j+1Ai3mOrSSILJ7au0+44Mp+Ltmr9ROrh
FAFYcZKIXduqENY3gWTG9XIQhgremSmLSIbZmB+pOhqMNaZUVYLIiymO9ZAo
URgkV70jjg+OzDCuLiEKE1EheBRTvKMqVw95f8NCCp7dIjWAsItIrIeNf0cX
EHqY1039RY2Efh/BtCkWehUkIPsLlHjZ28eDa2c4Xr4O760lncNooFouRPDd
7Cl35uky/NbAXsvcEXfjlu3lhAg4on2ML69dak7ckuXD7LEtppY5DAEdAoHt
gAhETfxF5ol0Nu+AsDeyX1d2aJUlQp4FbMR5LkAtKtCD/lK1DWTzOqLUDfsU
MA+NvUc8Ahd8AJiDW1onXapgKmUTA9PhAsgSQqC69IIX3PPcE394ern3AT6e
Hyw1SGxJY/3Am0d1c/zf2KZQ1aDDBCGnrg+6hbC0g2FIFw1N1nXiwFgJKNjl
NzTfSqM9xMilGYzPTVtEJIkZEmg02iaR9GN5cCLWREBuDHz5SJRJmq4zlVBn
RSrhd7FnJ8jsm9aW/i4RbIGstm7bZB0t2f8dM0XQiY2flEhiLUnap9Q5/NV5
fvldmGa+A5UVrqB5Lord1OPNzq+DMhaDd+hKob9KT0FMTmIAoob6iQE5db/6
dRmQDciVhRas8m7HtR2w298NCQHpK/GEWv4hHE5u+yyP9ApoCqkxoa/6hDqF
WBzOCPLhXg2ooJIVydXAF0cB/M/SJOvJ8bhOg0gs91UP5XdSBWQYyNOgpryo
EiBo/zFwlxLNB3xw+7BVP9aZh+vnIcMx/bjcK5JEhZaqMe3T6ESdUuthicYK
EdO9iuZiuDlNJ5N9ZiZ9B7YfPkBkXUS40Y6g1kgAZbGtR4OppRo4dzToMtNi
KMY9APH6cH3MJUp/QesgVPyLhlGFtt8N3TidItg4pfDtx0FdEKJjOFyM2L3K
scilnLBR1dmcyoKnWAIfQgYZTm/Beg7Q3WToOffeNFGWKPSTTD6En8TtPjvG
0vlWhvnvxL3yVsp2nsP3OMSwZPVgnTgRnKzE0Gr+TIWa0+rwEfgMmSWGhl5Y
jgVQXQz6RN2yctOENx/86bMuAJ9R+hBvj7C+3ASRanSVL27glutO0NkR22Mp
KsbSgep+Ncj+IDyTevwuvtghk0eETvbPEUnsUZRyITZ/YulCSpO9T3wVS37q
Blza8lQPG+FrQzZVsBfLdDqcae8njk7JvZYetOO/EMxkGvq6fqZxiUeHSRIh
rh/Qm7yrqk7geFZOHZfjVlg5IxVLYwu8lbBWh2nrgbHOsFP6RFOz6V94NwID
sxe/cB3R8oXCkaAM1gVgrfananzJkB3U4SKCDH6P0iLgRdW6jzob1XiKdXOo
AodIU8i8ManxykWDc+W14rek90OFsH0jDNsGEFU5Pg7/CXijNH1QQsmGNPVh
K0lmPEgUEpdeMOA/g/I30Ecsr9MjNjuKelMN3BEeuTIGJkDsyQzBqb3uDnQb
gpc+d6zF30Yu9yR7940/GypnaO6CtKvpyTn8ZfZz/xZ1VHdk6pGlllsycp/n
FWFsIYRFEdNJEgWMbWUBDOfvfh3/09IsI17xv2s4RFJB09efs5tRohbq8y2M
bv+RaLYiex1YeN9eZJuA1jwi/yVgh9HidcU6gV9PcyOFwtgDEumwR0qkA8ru
MgAv898WOqT5r2XvpZrrPf0PkZmoDjoURQJL5/SuK5TBNmI5UrZXf2X8dUSn
9PbjH2WeSk7up6+cwFNKbZOhLYd546peBvNGaBt/nBfs1Yqol+h3MsEl6mRO
G8VchLBD1EY9Ul8nrZBwHiW2SsRJ+TZGq/sFEM3T03ty2dlUKEYSciZUOhgl
Nl9MaOsu7QxEzNXnqBPHLpRFdWapVrMi8+7vN8sOnj6/vLEYTFVEcg472+Bq
2fB0qc5AlylY7cHY8tLo3joRe7KDeifA6uAZN6PrPsFMeYbyOCNfMBIRzknF
DJUjtMyEiQzeNB3NzzGWfwiU6TArc1GxlzLiduBkdvWHqnvNGupWPY0mJPZk
AVJ6vwpy6H/sx4PYP3iusvTj/5dHD+itajHd6EqqXRwsUvVX4pgnfMDSBCBs
o5lODNJlsjfB6O8usYk+W+FWR8jKuZ5wx2wojmC+2nIB+1JBBeV658jbm8KK
5zUJKL819xFuK9++sw6SYE0kAGni5U3CmQP2IbYxQ9A0ZIuH2yxeG2yCKh1A
c4dgH4RNipurGtRG47JmB+1+4zEwG/bV0BNKwCZ2iIj4t309GRjodvChZ4qp
C3A2q9tS8G2dTl5WLzrRNfivkLuIGyugfFDnzEa9ewrt7837YKzYCl5fdcI/
GjU83r3sIrcwGBl7BFnqPgD9gZkv/Ym1np5riQe/6R5Sqo+x0UcDeo9vVkXc
VLUMc+kJMBXrnikrWUyWZIBVpc3+9+0r8JABtEaeGa6A0Erf4LNS3QnzKDb3
ZxDqBArZGOLJjU52X5mrjm2W01UQjX3qGnwHhh6JvnKwGx8fg+oQVvUMDQQm
9AXzV3KVCABfFk80HGM8SsT3rCyiONsah6jW2z83Cu5nECFpkDeuvPIRrDVJ
LxQNm57Vj5O4GV7mwC6SzQkHZV8M1smt6uRv2P7F1f8YfPqJ9Lzf0lXH7VdV
1LQ/r+5ySablDf/4EZuzRVVdyh6dwdfYlno7Q/cEP4A0YMMCP9uGqE3crbAV
QmCFVAaMyChFDsD+zd8FR2blcRHhl+wz8TZTEdqhLySPVUfYd1jsHfxZBK3r
bdgn03W8h8jkRGl6q/VCyc12LFd27CjkUW37pKi7+g8snubiquUDzKPy/KPV
79pHJpe7RQA0BYJAvnYEXsJkqz4gKQ31egVgvFtx+Bz+S05C4cKqPxsirFMf
VISCXvueqBHstKx4+1oA9YD/Gs9WuQ6f++85yL0klLLoi9tu9cU3DA9vib2m
UiqJUvPrM8qKg43iB5jEGeomW88T7cVfNh71ogpoPGtDQ6WHNy6lIkmb/00W
vM0RTgnv3bwcC7z6kGW2j9c1C9fsyioiosjbkudS/iyNN6l64CpbiNbL5nkK
jVo4O+wKnfqiHyeeBd0ikJ0fFTk0mQ+JGc0guytmxxOrOw6rg+4sBjJBVecv
uBtlS6YLI8Q1bJk3M/TFXJWqvRbXqC8xVPoC0xX98/Py1uyKaNt+lp8lxd1a
kvDluitDTwPiOYaqRLACJVJ2Ib26DwHBiNOFYa5hbYUnpEO3CTuFowIUBDCm
X6rM09vkpDklL3IFq1tRgK84Ua0AHGbr1/6XX//uWqRoDt8GxHVdlORMAL2N
P8k/6e060a4H/wLkHNYMyNNnoZZ6V9IKJAEXteLh+0lWEv3ds9rKXpNn7YmF
amYAM4IUw8udBGVTNWIn2G0WZDAZJmp3MLRlRmJ2KfT0u+Pl+MiZrT29BvhM
l0hRisNzdydFGkM2IMKkRJNQRtrtc40Z+8VP7uTeSW6aEQtnVdBv5wwo2JbD
y9+pMFBUDnt6CYKn4zNQ+xIGkDcAJc7pa5MT/5pxTVW3rc8JorELwfyWRJif
54uAvGz8xVHCaTZ0GaPWd4aWR/jIjIv5241jrOntmcCzKw4aJ1VRUvX9x8v8
BbY/urQMVMVms2d0qcD+Kl3+WUV6IMTME+bdddgc2hgg6ALlLrX5o79UP/Tr
LJa6frGi9oYXas4wXg6kjoE2vFCo6j++PlAs6NKRtsDNAzBPZB4Ngkd23Wc8
hE5nnt1Vw61GsJR2mo+cN0Qa2eUBSmQWJsfg0HVPH+Cy092OGGXRQR6U/4W6
6v8Ct0O8PEIOeSiHQw58scv+rZjS9jGNPys8u2QnrM0A9Gzpug/77Qk17Hl/
1t0XZRByQaF2ts57HS22Ww7+xBCAl7J+7mefdvmJPBYSd7gtNFh6C08pjxNT
i9g1WbTG9vs3Puf1YnCZKkoWXdcDaTJZbJ7xQNURL+TH1n2gyO58AGlComHA
zuZKASKQIrIYisjRVL/dqUrEZjjFjv+GJgJgCv4DHgGirxBqyMnCnaTTAiVc
y2zKrCS01MrnHUFBKBaq56IulrMsPtFPakEeGYHFcS9XUcMZUODv4qX+5qPM
Iy+lWWFjJDpRADFubnvTTo7ewXhNeomBwTDqQjt5OdtyNwbZgpwD8a7JTv6E
+F1w5cmUWkLWgWQT47U9aW4KsZUl3EOFDouklBZEJAyzAdcPGSpA49mJIWQl
r+wvLTn6cyi6neKXfqvhPGPAnBEEza+8iRwV9M3ID2h93iBHqOd1cNimx/2+
kkC09r1Kow2jvd2YRxYcJpxgEREDToSWSNQNw+LbZSQaggihpm9AALz4rctD
CLvCtpcpMIAM51lnrWJ7mdmUp+Bxyhl738CecrKV1H4xvwi/i1VutDe7pooB
tvvNFKCBgqphEydi3sVUS5BGCjE0U/x40q8FHWI5Hfwgzt7qY6OhKNaDaDao
LxxByTc159o4WijMdZLhrbeCHRQBDqkmA3qgJRRFRyN9bbJ1ZeeVqZfYPu1n
5lTFd6Y8FcgoldVTGOry8G5Od+5pU92dq5I/Igq2pl03EytSr/8cwxSuESCd
8TbW65CFX/5/zYwNR0/X3d41NYcd4Tvdta6TQn0bK/mFGL78cwbSsUA2KY59
2SSZ7zbRj6r8kf7DpsEH0WVn6WB642x8/4i1wGAEYdXc55s6huX0XBnD9mod
049yi2wVjkCe2TLr2VhLtLpLVGG2gP8YPVNZ2e07bnjnAbIUQUwdFx+D0iRy
c/L2P6SV6Evsc+NQ/cIehhzX4XKTMcvWC8R96lnWCXOg4Rp2MRuCe8pLGBmp
2mjVg5L+yjxZv+djzU7Zc33KUiqkauvsqF8pEtZ3Vc2IJCU1DhHFYq+QkcEI
VzbTjm2/Z9kYSw3CP16Wvi/M82fGaBjdevVShBf/zhaG4OlGZJJIdyjB/UOo
7RxlOj5bGna0iZ/5Dg7khL76VgSuyDt+vYLRvyynf+eilxnhxU3pcYvRCTzq
F6wsHz1OPHRBkh/lkRQg+MVU+5LO3n4oyMWhrD5olgrTKNwlKntterff4uws
s3EZ/T3QEjQYUThCAduKiHkHr0xVQJtrXY7YJoUIUQoIDsLc2TFALbmjcXSi
VDXtSK/qwEac1sG+R+9exgatyTBlR5hBRtwgQ/ytubLX5xGTnVER1nk/VbyA
rlnYx5uXsT/S6EnOp0wJTr7j+G7M+YFr6XvIDekjvmfQ5MldftoLgSCXBAqT
uTxp2Y+3F2MSP7EUmaC6uqy6vynp4fCW9oMVoyvSWNCnJy0SUT2TMEF6kPqM
mgAM7lUpYYc/KnxIQ8ne0UJeb31OtZ17EF+50YvJy12V1/kpmIn+VjXhS8cp
+X2/UrjFE5dYoyigUavUd5e4KMRutyYJBZnH/uEbL0VjV3JquEtT+OWk9OR9
4xAUCEbdhVPh9Z+Ax7JeH53Y9ULjPhWxTetiMv2PjfuheKIsVcxj9/lx2zHH
UKZM8fl1cOGqNuXYD2ujLM/WpJGagJST0es+Xr7XflKb8zFl4lnUQ21iS0ER
ljEdiTnc7Whd+lwr6US49YVXMcJV91C6GES2VWNgTKdyBuYdTgKzh+jTw0iL
FrlzikWuUvaTi+Uod5Mo0m2krLgvhBkco4MnpRAQFftOOHQFzFG8b9Iw0FYY
KHC9FGY8kqIa4vdSRWDuhR2OpK9vA0XTeq3MLDaIEdz/XvK0YsKRIRm/kxxc
H6MWJ8vzgmHgiZhyKQJ4dC056tI1KJw+cdDs2SwT+RCbF+LExfybW3I8wn9F
/i0iVhrNyESWCVtC7Z17Tw7W3E79rqQpILz/iR6kzTXVK34fiu8pL6jP2tY5
VxNQObHDscMy1jXwhokblFbWUcQ1VBnWJvno9uAwCUwg4Uw/WR88LYuRZOW0
Ws1BbQmGpNnHThC7RvW/5/2Joc4dNjAJ7/yr2Jx3T/qLDvjA3XpHwZGWAnp+
IJ9/sp88YWwXztYwQpEj5GYcNSY5hc8GfmqjvdfGPWGoaL2mSVcjFMuzYAU/
FfXeol8GDB+8vVwwC2UcYcqDDaJKC+bDM3BuPsi/n1agUEtaEhQcQ4v0TB+J
um0E7V7Gl8PKJgdzT76hPzP5K/vA8RsFZgxDmvdk2wMfDdgbmSYSi9sn3rhY
8/O4Ic9I4LK3JK2LxaekGMx5KWaojdiodOn6Vxo+81X/HoHTIL4T8P/G06yS
p3EDkjd1Dnbr54oTUdNaPAq+YvrihcfAl73n1EGJJfss146EYI9emiXXcrsQ
8fPBbiOXrw+6DjAWrciZeiD/Ow0y+Vzt5Ym+CCa2GNDedpbQgZbYmB/h2pu9
Nbxr9x5bm1GxnGK55zq71hAc75YG7snjrBsyxLjukx7nNQvxHJMo6KNDlMrw
uC55xYnE78B5MrHDJaGZPXZzrYc83vAihFJbe2z7eBGuZj7TmUBKORzXE6+L
Bvggw7Fq0JBWjegIFlZY+Hw8+mA0M2AcHxSsiZE8q+cp1Q3BEAU/OFB1Uv4r
6EDGB5tbHEzkz9rozOR/8aCx4To/0yyF7NfygTf+1y/jHlfcOPG2Xd5yQNh2
O7SU7XBQA39VLIKQLtQQXWfdPBOM/gDPmwdKvqgXRL3jsD6EPo67yxtfT5in
pUPriy/eyJS+yHPdSdM/u3CEa+FtPgEevYPM4ADYC9T2113SkR798VrY9Nni
FQtLnSmPxUtAXBUwOVCLWkTMspRT753oaDsTE2tyjreoJhEVD9I+QqX04jYR
8S55YdW02MmEDjIMgib+IcYfmHArd25dvEnca6t/sw6zQF+ckCEIqDgrI8on
vJpOxzrbic82ub/dz+673zrEN5nlE/XjNjjy0sAs52KmCtzp4IthPsxf4i9x
wcdoZGG7JG9gmGy4S0ohrhEkNE57oRUXN+E3jgK6XXPUG95r84p0DzGhIn2K
ESUUghkAAxIETcRiU8GsWU0znqOtXV2gPcA5bxHayhsyV+JdmhIWqKPooX0R
03FIBrAnO2tIY81Gt101koLtS/ipggOF63bqDzsdxQ6kvlf4k1vf6JUwW3R2
axWJTGl/XopAT2jbdc8idiMwfmV2LA+ZJG+TDxrImEOUSvC4YwsQoF71rSSF
njiRATirCNZ3/vIhKB/41qUQfdm62zdImYqsrboiFtoQVPThrf8fsx61H81Y
8OqjXwAH/VwgxZC69alLFmHiX+RAnZY25EIu/cnpP9fUDoqaaupg1tH9gZxE
8Rr/dJlJPtFbqk3vwiUxvlOKh1tEPz6FT37hvg63rzlO4ZsQATcLcQx0hOt+
6ROt9eujoV6bny8ez49mOHPARTJzmnMcehul16KwAfUZmeRtX0c5+KQL5+eR
dXN0umrIJp1sKgJy3SJcUHQmbJ4QnxBSsFsdVoAAS1+OedUu+fGMPIK08WGz
6pJMyvF0FkSTIRu3PN7zDSQMBeUpnPW/1khmvkkuix3+NTKVMxAlpscwLYJ7
+BlIuOSpK7hpxDYWLrwKqrjMmt+HqhruMFnRSiqHRr1mujyU0WM9FRwsSdzS
6lqN8sQbbYLAxuEP06RLzolqY8hkn157/h/ceoFGSpiHPFIfR4Dm3vtOdnjc
zOc41lPOqblHDsTqQcZSpT5j1+3HyrvZ5MiUaIb2s7lJttw9yjnxXdJP1YEl
VjgOPr8asG14BW3v5L6zM37+Rgm23apaL4F8j6A1Poo2kJum+obkou9NBAFm
T9kJoQX3XpLsZ51xbqcOSk4bsCCMKyvMEfkwhx0u0nkMYn1XX/0pMbSmEy6M
qnDDxvg9BWC3PFRp0Dnx3Tv24VIwKi0a+jT0usST/bR5ovHqVao+IXKMutKj
FMMwFmenuMR1NMLoAuB12abMyAP0v+iIWwIELfh/Sx5eMR9f1JZaPbRTRWUQ
AokiMi8Th91jMHefeBquYeskWld9eG0eYJTBkhexUBl2mdqOtXtaaySg4EAG
wriqIh52B540BJxJK4EVjnEL22/dJZHin+g2miE7vrwZJlqnyZOfUDPEEvKV
ExHdIJd8tMigL4eE/q+qXf2tfP8Q0evrth2cRVqaLXxkbP2uiTp7Y+ihw+Qv
3+Qd81DOVKNOvSoASPkMbDpnQ2GrteS2ZdNML15djsHALM/R6M5J3KEj2jfF
YfL73bk3rqYdGsGRdvww7gs10jYY1CRWUo9tfqV+Jq8uBOwAMF712x6CiVOI
EzXOi2ZMIh+/507zKVxHJUNAy97ZgF2/Xf+q+hZiZyDDwlP130MyHSr5IZ1j
g13Kgs4IzvEwi5aE1HbQ5fZ6SH7HOkDBNNPmXkBtQsRqvwHvribKDryOo1Lo
y3qZLjiW/b7AO1nZ/EhJX1S114AKW7TA+KgagQgjFIi5S1EEsNRtYg283VJ7
IdcHVwZ8A3GIyaZ14htbxs9mqJv+YwKZ4co8WCF35qxiAgICLt+GD1vtx1a/
Q8sDgXMzztRxLCLyAU9RiReW7dHSa/hORE7m8moOt38hbk0Nuf65kCJE4I6T
HZZ8yoI+30KstnVKWaUDgniyROO7/RHuFpK0FOpu+lKC1V5fWR2+JfFJTDXA
/2jBXPHt6ADUg+q18WbVdtedrpsDUfF0FM5QEgDQ7Sf1HoBMRhW8fPBCXw9C
i5pk//fdYlaKg5xtZEs9juHfOt7qEedpl8qMAiXU1Pj4a2hn4AtSc6ZnFSNT
UKAcBDUUL20P9NKcgrMlVBPrMmTOelrEYPX7YFkWyaDTX1h+5B48V5PsJXl+
3VolqWZVoNo1GqirVTCVIf4J11qYX/nqUv9kk//lR217tB1bifwr8+GGVTHr
CyhyX3ArEkBzWG77rJvRLGPtys/4AqXF41LM+r8fw2gyxHp2GkicBri0ZWnn
UvlB8SkbxjFhhRxx01lHo9R5sNt4cRzEGgJiPKyVVQaxgVT5DHa9RAl15xe2
69mHACkBaDV/Z++Z1UWqjBcCPJUAZlBus4+HRd5gF0kjh8yNYEgXIIOpWetO
sGRkl8jl4ftChkLNqr9ooOmAaDTVkdGIn3kR5xHtYpzpha/IkamxsB3w5mAd
cHTitA0bv5xf9ugkw9S2p0F6HWHnCv4gggh4zfMvrfwpJltJN8BgKoIo2GiC
cjKyGb9cikIDBkas1dwzd58oRAzO6PSQWNwwjA2lLuWt9gdliM1N6fBT0aSR
VZXhtftJAE5i9WnzVE4vg4p7ozAZScInrf8eRm3KOGaTi458qwsb5V1TEi/e
YOcSrjgQgibGGKH79Hefswru3qf+OgBFL4ZF5ovQiZAFOoh2VLswOY1ySB35
5scUlwaNcN4Ut+hHSFWuckicYiq/ZkGAWnf8zV9htjJxvThzdfpo0/swKukb
FOi4rQU/DOJ4dkOp5z+dwjgUBxDqWHYrpX0qzDLs6Nb4Ex76XJ/v4RAEw6D2
LBqmVWuRY3yLf+cVtP3Po0zQ/ZaVB21q81BolYg3mYuMtxpFS7YG/OHeJntC
c4ZS5Ljb/s7qaMHf4OOOpCjDKWMRUFzeltAIbImLIzrvdR9YR0IVN+XQHQtG
ejsoiGGmTp3FSCXZJ0a3Fqy1e9am4kuhF+7KuyuWKmJlQrjYBy3AJLTW3fCp
19pyumNiHqIDIiohYcZFprCzPPubXNNJIA2UB2QpVQcf+uqtJx53RdjvDhlu
iuUICJ1n4tvEEw6UW/mW9JrL1eXq660QQppI+ZCbsD7IMqwwKvjjeDS/J+wR
suQGZ+vcsvGILNvDhwCEOr0He+lqGM9A4ViagnqCnz7T/oPyppDGmugnYk1j
5Nken5JRcQPn7p2/PZ3Y+CAxh6iKA3jpWT0Vrfgea2q4oFtRxtvsVfsgIJ3J
4fI6cChgNpIM5qalaGBg4FsvpxrVbmXIffAgk9kyyYKVciLrF6dsKrMPy1Ei
4AQOfZnHdvcO+j2tJAF25oONxgIxIB/xglnLW4YDs7bP4A+q7pJHet1NT4K9
q0eDlJZsVI+h+B7A9BcHdh7o1c2rmbep9yVitBl1wAKmfaR/4ZMz5uVz4nGs
L16mjvQueykq31pSZDXpDHObgDxbjGqV/7S3roAKvtXMYFIZ6OGOpvQpQ5EN
U2fBEp0HYLifRG834cvXdC0oOVJ0+eGmVfTRmLeWVUhZfn9pNiyswNSMhliP
x2Rf3QDR6Y267JfOcL0zgTcT/s7tpXWnHlVrtdAk3wEQO19BbDbE8+iOhrO6
z6XQ9Bd9EbsZe67rOh5FxE5BKV8lWn+NemS8FNHnOKzJAzgW1Xz9WtwUh2FL
J08Kj5UxKU4LtMKetOpSmR/Gqz29IuX3qMVr7ELq7wix0aFPtSX8osManOR4
voAscmrtKhWFrrmB7BWMru6d5chtiBhYB1Dr549GyFE6ovMIQrdeHn5teAZA
blOu5yxmjfZfWJ6lglD5PJL8YFHaGwqO739IRhdj9ofx/UiAXg67P90U2R+k
TmULSZc1Kxqfl7jAnfxm5XvwuRr8g5KC6XA1YJ5WuHO3c/Us2HVv0Zaf8CvF
qiJk/Md+OIhwPRolecDh0a8OFND8iWTFcJQBfFLls9t5h1uui/teWbQV+beS
0Qsgg80hizcZ34BIrqIrQQFq3peFrS4P24Gr1QEpcV+S/YRVD+7/Xg6kVvhp
iXz3dZHj8szEHCrZijPvIUIYMyW0M8bAOlL1XGmvchylV+COeWHmjU5Zy4bc
cFOJ1BMCaotQFK45zJgSxbglAe+wsFyJQ/1V+YPKclF2pYIPftYmTAFIVtA0
IOeAr8Zt5SwwXX/ZUgCh6AFy+mz5g0TSfkt2mcScQrLwDELWtCDUPUVSImAo
5odKyb7NGVUKjyXVbUlEeawlX9Y3aSXr0ejzmjPn0K3Fq+ptkO2LXbe7pNSh
r4+lkiqMmnPBTFD7X2e7k8gZt0nymqEkNU809+B86M6cezStASDEYHZGE/1Y
y70ueEztcr0mlakG1lc442NUPvqtTw5dFEsosHVqema6Csrna+UkUCeSuR1z
riS/wIQ+SIExBgNobk5sCD+VY+CgmFfweEpWZmvB34a/8S5fnb3JrYdNKsQ7
coVlWN4mQermHuwb8wuRzHdmUV6SU32mIPrbbzhkOL0yBGpA+X1ZM7eL7vfq
K8XGJ2Fkug0dnvL/3vs26NlEKOJz51ic4Pztqv95j/jtJc6PZTBb14ozVbNu
q1hLNnjISSbjNOTjcMT0qiIx3aeMbCURqC5FH/1NZb7602kabI2BbaVgyKdj
PEhXVVoIoPtEBM7VYwEn/f7+qiXAUJe+s75Shyur/f1VfD45mz0QipTo0ZFs
cztl1nK6Z2oiJ2KbEpStCeNXp8ifjv3G28DOyOQGDasSu9f4Vr1bIyoFEmJw
4A0kiuDzaDb/6iGNuis3zopnfa4t4UJ9MRyDyCpyrTz2EIbgHRi23w+ezGyd
0qpj9Kx+nLbGB9papMu90H50+0mzFmxG+UrUxEAogZ1aMhy4VLLUaT+IvW1R
Tym1qF+cKRyK8AYN8qpqlGH/tSxs6HWFWlwEP6+9NGfU08Hshti+GsTqVKyY
5izKj0JJfy4H4FPFFY0MlHBInpu70XOhY7z8I7M68frCq2FfXwX0JavrPzz+
je+fE+VwDnH+sQDtrdt+dnoL/SeKWDbvdk5KOYbfUSzUYqVdVBE3kixt5yMf
h/ve0K3zNcb+859agW65RG5uDUT64UsRqk6co6/heXtaSZpc8U8KQzhnCO0C
taKBcmYQMqWbu/H/2uq6xGt8flwi64P1CbXqy+00bSLNEXaQXNDnLjPObId3
2uiss0IhVwTi8ia76CSVDtB6E8IHWPWRM0UyYqziS1hf4PWcIxRQfP14FVDR
A/eLB8nH+wsCuSbimVYqvPu2j/pk3LJvG77n9jwIDIeBknTQnli/1m4DWTee
lLtLQCvJT83OnhHwX8VW9DtG2nurCdpQ7u+Sl3LiAZmZZz0l9V3+v8PcyYOB
9jva9SxL65pdtf8Jv3d82BTS2KQZAGnwbRJOhuu5aSCSZaI6DXrcoxLfLmCq
IwHjzwD9Ps6wYBLQYEIlLJQECa2a9d15DRsr1EDPT21nHwfSygyYsi5c64h6
AHA9wgSDQ1sqM4D3I2UXWFxw10Fb6iUYB659Cs3PqKRweQ+73/uzildwOT+g
HJhPCaj9g5wFKOkH24IB3zEEQDGpb+sxWEUYuEE9DgatSMiA57xg2AUfYPZ3
lsmMN8cvy85AIqR6+a2vskTjH2UDg5pN4vvUOQi3D1GQW7FdUCOZVBoo48Wx
lE3fBNgNsDYgHrcg2qYBvQcuAT7BG6SPELCC2lBUrVzMvr2HnqaC6Uaqlp5R
aaSZmeWi+KUTWnY2+Cj/CZtoDgHqf8ZzvYbYTlvBO0OaspIoxg0g23gCTBSG
jXtu6zGaYyJzlA/Nd9sDz1rscc5xWyFg0058txcFMQ5DpUycPxBpKt+ZlZII
IuvX5XLtALF2kq8ZtC46gS4IfohEqkF3kcwWkND2fapc7jJGXL8B+PyIS7u1
WK+5ON/ic/qa30U3y22x+PhJCimYPng2nW22b2bnUXLQfmCNnH4XM8d9vXuq
0tyBtLocofil++lVz+bneGMCJrzRUSA7HbGf9CwoKV0ubfrGkIat+Mbvb8Y/
D7aSg2oekzV6RVgdCENd6uLL2oz4mo3/vl6TNb7Ps6Llv0Xw35fDWx/hWfuG
vNJN6oG7TeDikOSy3YD3/mMKp+kB2JKARHVDFiTx5rwNX5oQ+q95ALsYeZ/7
6UkFBTpzBB4x3wyeu16h6ftliZFdpZmYWkmDRNFNz8erzRAdOPTSAtyUYpiy
1cqdDFYfS06rJX1YUUr4Qhw8ctqR/7LQaEtFfpuDtXzrfk3GHidTFjQz8n/o
9htUet3yjuv0kE9Uw3Um9lZRv0ECZNCBdsNjy1dBz4Nz7xvkBGCpqL9EGFFf
3/uaD1+ejb1R61Wycd2CamAMopl9spY9fB61j+UJpgbcOrxJ+pw38SID7Xea
7/xhZG86xpyicihhH8yyw5ZxseBPFw5qV2IzdU6bSvYedmukvf23V7rgQa7A
P0z1qmpGXLYtRk+B5sAgjooyS3suoScWPQGW1JgkPYSS1dZp9RoJWnkmiyFJ
LWCKix6Rs0RdkJ+7OzW/PCbvixAd+DefmRUXNO8TmwrBcblWskYKZb3dIF/q
RUMLSNO7e0etS9GOtnOSlfHoLHXSJJckT+ArMn/YxWdZxucm4re0f4vj7ovu
tE/3iPBA5P8lt75+zjjxmorWM7wtv6JEAGDt/FSoXyzb5od6gyIyysfH0zSU
CBRiN06IL15O3g5H3EEZSlQiIIVsiv5qkbpwC/yHxp0whpzgBX27KXZH1vZ/
TZzw9JoTNe5LW2PA6dy0TDohoC1+coViXeMGevzqLaS4DKnuRXZqWzniQcuB
CHKcACJzdr/76zIb5uhTloYWEJNpELcCxesQcyAgvoeJiwSRIqjUccEGQlnI
YVwwHys0DF48Ov37j5Y9BgKedJT/ppebIyJhxhRS+34S5ZyrEVCPq5sc2PoO
hSptl24cDO2MsrVdEkpavN/+l8P0b59iZQo7rAM/gaE63AFXvsGHzEFV5nR4
10TGIZwQk/nDK74G8vciqcMFLMDQgplUjcmsg3UJF/26yvxtp164y/+iUgdz
Sme4Z85CGab7mgIZNElArmPSJjuqr6iWlk9vF1TpnCu7Eqnyi5lbikXvPcpf
6Be7gkqU9Ffsk0Z7WaxoSjvR2Znb1omf7Dzp6ZwmQn1PlVCv1yg5yVyttnyc
ya45vQ7Z30HHIMAzXrdpthORNArIRNsH/LvXCTt/h1idtrZZRed3wg59aHr1
wr0KWS18Aa895TMVxslXPFjVw5OVq2nkWfi5T9lf0SIRaYscrLdBmWnma0lN
c6lDS4qty0Entr+8jm2rHCsHk7yQ0RDcIznM0zcCZ5VQlSNSjkhhWzxRo7am
w92iR7YOlMzs3mE2SuGgs3zhGZYwZJzKjQ7czPthADE3fl/oMRpRwSN5NFuS
6oN12KHM+wFg4cPZjkEWVsYDuYssdVZYlqm3LCJKR0mNaEk9x7Q+KCmXDBrW
79EDNbKsNnC8e2fs70S9IbjEyB+lDjx67nAqmGeTKY3kau3C7+22MzfagIBD
7y1z+VS60Tv/1OUh6q0b4ymLrqMWW9LO1UJqIHDIKNsGRS0YQtVMvIZ2VqEn
nZSoanSqYv4P4Xzz3EZ1YWhZKKJk3vL+eoW6JpIMoFhMZPwcggRVwchUbUJK
f5RTpJTcoWcmMHgPXSZfYGwEXrB6d2dFg8D3+vHRrx1REFJ+/Xnnu2IvZB/V
N7S9geiTrkOcqMcGX92LQzrz9NxxTGDuVt2aMCv1OkdU8YE+I8qirff/KGT/
cTdq+SeVVwWyYGWeqmr96bs6MZQVA7PXh03skZohG7LAhiJx1MeHh/xZDhyf
EGcOf+R/2pPZCpmC3f89wS2rCpB3Bd+a1vgJg8YZAJHpnzleRI/k2OvmKmzB
nsbDjLWrjoIWzSTSyI0Ms8iugu7ZOL0O182HZ2Bn/hCpoIyxNOWZHRCG7iyf
aMTlVjVXBrZ54sk8RDvbk/AGUbobkja1pPbJKQS7nvTyMKXLMF1K6D5oucwi
ZeSD7kprmiTQKBQZDNmBUaIQsGj/585Upo40btoQceMf8d4RFzqVVi3H4yPA
MD3AZh9keHAsggxbUASEB00xV1TaHG9bMv4gNEKb1Grp+2qZNMhg+9zKjjxC
dVFPIN1Mw4npajW3X8Zu2LuMPlK0ncsYdIBsk/LCMUfOkz6ufnfQQW4LcSyh
GDCYmuGTyYrCvZYNEyyopLD7UQHyGs09F/3pFnN0wFl+JQJukSYh0CUFBkR7
rv9PeKsjl+1pG0Vk+Q/cTZ6HnDuu/lv9WLmE+/5BHSazAZfk/31Be7x2yFGS
xK1lOAHupdg4suWfflUgk6nhNFigg01KrUZ+TmEh3wez2j9bnXEOUV0gylAn
qrVF+PnMs9+vg0113YkmS1XaU3nQe3DOvUfmk0mt8HzOcugyhTPQS1v4Pw8m
PmEoHfxlK4zCzkqWpiSnsDB4pIb9hWNJKYSZlekqBwbm4mbtEnJYjs/h57PE
+zEroI58nyueZwcGQa8Mhu6lveX9/iSJ9fYeKLJIOedNcyWDjSEz3m/AHUjC
R2TfPSPNo/gQIiyX6W6LxHRYGEqYn97plZZN08UB10iff17tAlS6N7cyi55F
9yhCY1UaA+3LYcMUguaEO1vHr/Ue0LehD536UL53w+dZSGT6n+pK3UdReggF
7InI3YWDfiUVsp25m0545cvzeXls79E5kazLdcfzsM+q+CLB1Xqpzso7fTe5
F3m/OX0ZXEBR83mDsClJ+5o5gxNtyaFQLYDzKwM8/iTEurbEAgmZLOjZVNtA
7NXZtFcpX9GBwsNnIJCn0UyDV+RWxObN4woOuvRrXDqSdTfKgVTwj9400Yc5
BIBD5PqwkvrDS9pqNI3MqqT+L6NvWs4eFAAYWaxYQfMbF0yOOP0T5mlo7fDS
k6CCFMIRHJkShbNxGZR8HMXgNDD0GtD/dmr4Sjp0AqNqWJc6o7AIW4z/lMpB
5mUJeqdHbYskY19XpLNFyfOzFo6cRd3ie5e0klEvFlD/UqBjUU5m0J0smf9p
d7Nu29HdIayKehqtqRHkPaIdSQ+fd+j1bH2jBpCGwiFGvTX6s8CuURkgJKLt
HDqpKioOqslTYU+EIBVTkLeUfqbZSRbHez7Y2cu7Jr346BpI/jWnXrhQwcyA
GkNOG8q08PXDdQ4Ma8dvawYeF17xV25VKR85J5jQNWeBQ8KbYH7Ku0VwKP1S
PlPOx3FHkt5hvTId4VzNHF873ZYJG3pv4IjMGg43IVPPGRSQ+e/xhX8nWYsd
thA0MdKx2XQyD98iruNTY2m/SajykKdzleKFgGxZe7K1IHCaiYw9i079dhUD
6RC7mu/AqkhDumBRho8l2ga+Y3KdnWtt27z5Db9w6Lg2DKWxX715RysT74es
Zh6NXVHasu+aI1vCjQygo1cQvCyJ1gtOWhfriUnuHjuQFIaeiWzv1U4QSwul
wzdd4nzlf2/wnZqqhiUPKOGGNZTWqSnroTKdZnsqdZNvI9cepfGwZIBYU6nc
GpqKUB2+hjSMCkp79n0B0bAaLX16wSi9sWdRT2uVSWRX8WQ0S/lF0vu15Zre
Zpp+XvNsw2GWdsDsnecSkrE4K4zVH5Ge7otdvSS4cV6vS7NBmHb5N98hTF9S
r7Yi83Vxks8PP4JjvTo22G9J3+FqDpo/qG+f3vok9kdKs0ABA6EliYhv+b6R
cwZFr+7vlGgW2pfO/E2fNP7chWbK98N8oRRLB5GMK0dBjSdvYH5eGzGXUCd3
PymYrOsh6kG+MyPLxjiGY+3A/1zH/ogstAYY04pGS8AEkepAItjEatJQ0YXz
D9XPQqRUtAOirS9eHVbp0/GR3h5rA5dQZvEf6LDWJfYVV6l/wBkZzjPJsXF6
pIsBYDFxD3lO7kIIG/75AZe91gkhKFTEIQVEcbYAbYD81fZ+Gs7XJpuRN9Y/
H7JncqW5k9nqa9OnYARwUasUoMGQ5l67RN3MBPFnKAMjxkKq76L7/f9XiErU
RoGb0R3gdD+DSGo5RXqyb6MlZy6h2y6eWm4W39VdZxF5Bx39kabzklzjoWXW
tVDU88/kHE2wtckUAEi6GRY4FhvlSwkjZeouhOY5d+Hx2PVFYbs6rZJp9Fnb
k/EfT4MlE2T+puZ6KsE/j6P1MjpU3dv+DQQtEVM+hxvaAJocb6484dpT5ck6
VsH8AWnt5gdBEvONbwV/z0JgHUOBBIzINhXGEpJ3DYFXY1R027qiSHoGjrav
Kd1L85kBV86OHNnu+s6Fqt3+FsH8pOZ0DfRprJsDZuo6W6jEuY8hBfM3TcH+
O21zDCs0lsO37j1ObJzwyEs9/URE2AQnfwbkgO8B9z6t5DKVsIa5onkEqog6
4KCtkt+LI+RiBIAs8utp5Ocwi8qCbOisJqo905jhRvkGmXG9n3o+eOqwZwxw
Wcmk00gLDL/zu5wLhjSvFgEVJDYFe844om8VykCPP2NCkH2AgWwqGHA5Gd3Z
q9ktey2s/hDNUrsMp1aCRFV1rVykqmvePgenRxJON2tcma2YkYguYYHv71L8
VXYx1SXkT2F80qV5UKYbp0zFMInKzlgMd2jjslPLPLwO/haAlzk4WIyHJJrV
xo/2e9kdpo/vNz1vi5gZWBDDLWyJYS1rJez+w1A0ZL1OqXZP6+dF/7F44oVF
hak0jgS5/zv0Ecrf1XnQh2tp2JZPK3SbFqukvUZDdoK4+fl0pE2kw4/IdkhG
5SpDj5i0z8LqrLm9bm+k7mTEvmxRknLN0PLCTShTpJHMQrmRg8vNVYbZmClC
/LqQPf5Hgm78H6bEmyBde/8IBwSHZJblKVZ6IjvARfy+XiGoGhKDOTcQ/PL4
UIDTIYgW6akev+xCVyfyrhZ60MV1ousnYNV1AMSTbNtEU/GVzKk9aGkd8wbC
OcC5eoEDLwQ1wqnLALPhSJlmrWAeVYfoxJ/tZqGvUDriEnNIMh7KplZ0tuGp
6FsQVpuc/0P04JWT87DOLy9c2NuFfj0mZbaOXXi7wG90kY67R6mVAOapZQoc
NMUd8LylzVnE+ZZ5tX52Fodqa0q52oWY0OIr+Rf9eRmqBi1DOs8/w2PoIY9r
fhNX0LKD1caOH1iaTmmI6lKqHjh5tPDbv68EMSVKcVdK3h3QDjNglUgikxnI
rdkq1nMg0YBuPHWDDTSj+WSJZPRZDVc0xsJdBDTFRzttCVEoNLEZgRjJSgUj
nm3elcv5eLSdrxGsSuFS+j3mT9rEitIhlesTlxvkPIjVZs99JJRlLtpUksUi
xhnlWLofdzefsOvNWJEWkb/e3+Xp+Q8xudzDEyCqkF/I7Ogur//hDrLxbZOz
YJQM7ya/auOvRfvtjOG7oO4gV6mA1iSStYwCO1OJnsbQ70SzKd9tfERaLJBr
S+wqkYz1uGheFEHw1Ap6VIJrX5qgdX7HzZJBcf0QvO/6TgbTXN2sSUDu1d9V
s2ByxqtCJTAzR9JKUcUNH/vNhO8O16lRnocQocpYM/Mdx11vXZ64FBTy6sA2
RlE03Vlg/yEITr/yZLxYJK57BTAAMz+ag8gtZxLCHpNQ7SuxrTzh86BfSsrX
1pZuex+NPD2GzfAZt5/hHO37oub13bn9SfU/KWH3RZfy0IT8CaH+DRlzZ+YZ
tCGh8gDAkQu5mDs4AcVsQ9E6HGJH8lGO97wilCbnTuBDuGH0lOFS36vo1NYy
MyuzbOsUQ5jkQBmfNHbTxWMJam8jepEBp9jEI4/98vv3bTbYJUuamZzQjZy7
X9+QYEvX+19MGxbpM9Zmz4iB+6R2nyh1i98YWVSkWsVbn+LrLCDTKkgZ3r1F
bou+MylBizP115H1cgRJwH8nIHbGr3ZRfHryeCajoJ4wjg7O7UWbvDZXGoxY
Fbd9y2gkszhEUGL1lMUhFMvh+H6SVERTnvNB2or9i4mPlGLGeRjDPHrDt/7b
3DlGmhncdl6z27dFwvXcJhQMSNCfl4mc6aDo5s8KsHoiYsrYyMtTmfulEBLu
NuMgKB+Ug+Lsto48HiTl5hB5W4QexYos0a3dE0RL9lhRzgqU1OWMTfx3BaXh
PiZF3engnrm+4iVoTnIUgtNQSz3ioQgsu8JGXY0p+mjr4NcF0Z+uazxqoWGI
MLebzdiUZNOOabEyyuL/plwTAEJtS0FNDWXUtRjXTrQW2ysOlcFPcevqcTrb
Uqon80V/VIhdiFqI4p6GL/AuDf/nGGL0dHi7Fe5GRH0YBnEFwFCuoulS1y3K
FBWeHMjDgVjr9TSODHywTmeIpGFHI0u35TEG0w+1u42WT53sbIYX84iobr2G
nY2uCmvVJLXawSeqbLTJPXMbHs/vXVEulhbCS5teuK9scj5+ZuISE9Hz9yK9
cozR3TNPYt+fW4Ld5n2g5t5LiEaXqa50z5nNZ0ZnXmFuPllrgUfpovprzRif
5LqZKmvfn0UoXbS4pneMNcNHwsO/k7vDsuN0r1LsqLesAAmNNIOwQWzrC9Fz
TLRWW48qhzGos2HE7x+wchwrKL3mPMMlBBgGRxNDpeiwi7pIx0AIhiVqx+qE
3wGAtMjc5Cskw0zEmiPiwHQMmSm//MaDvOBjdBrCCfhlAvaRK4q5/aQ+Nuju
MMBlfd19CiqrbkUJwpr/lhlxbUBYjL4RVRZND+p3f/uXV+iZXt2w3xMRUKA7
jO3/meCcqTttK8Z+/qbKWYuk5ckCfz2ioE1UL/qO7ZQYkdvVzr+JL9Dsanrr
f+CHyvpleFKHrZWj00DDMye9g6mQpUMKQ4/C1+MP2rel56yimmUrZdWqyFZ0
mwvhWzvRLtPFrpOll6k0L4L5VmwuwQjBDfqQHVAsheJcX18JD7Vq0u+j17dh
G5+kr8iPPjq5IgoQPQHEYP2JUI2d945eBw4Xmew9Q5dTuLKiQW9Qruk9S/dB
aYMc/JgQZ12B88GNJqxSUGwjEEZF6AWchkizpiWvSZd7okiO20O1pvcXYd3T
KSYoO1kb3FxH6jPTGjPJZxJbGgWvW1rCAJk9Nf4hBSZNRRE/1QkHxHte6MA1
FSEgZBYCOLSFYysZB1aI54sB5hgmqPS+xzxJOPg8mWoNqEZYlhrc8Z7sFpah
i/vCu0MipFQTR52647uNK/3xBoET+EAccWQX8IhuPU6+gaon5RzfgGJVgigY
+c4i0e0Cjn7q0MBr645GHQEayzTfqkMSJwaD8OHZUvKkYh6VV9X5b3x8Y+IA
ScHDqqoQYiSFWl0RxgiWwgoTrjyBqkWypQSi2Zhde7YYz7LnfobBYd8Ji60x
EDP1yMzVeezBPVmVeHZUgadocLTMGGK0yy92EHVDPELLf3nmebjUJ3Lk1hMQ
Cejfyi567H3Gv1xZgMuymdZ765tLADXWXgWy1el152R0ZMpA4MGbJ3TbM1O5
xUwuYKCFi9KqGb+vEZHeYqgZ5QIj7W23h7cw8J6ZC+grkCYVyuIAVkTm1dyX
/F4+lHAZLwj6ZCs41NIgQw9ovrbRrGzQw1WOcOMMABWdKVomThOiowHXFhqb
maDtJPkTnIh0NS2tysBFwM3EBaS6Rh1Pv1tBr0Zfh2zR69obeDCzFIMre9we
SvJvimIx6LVUe7swhjHcqfH+KkaAwLYzW6wy7jaFFRDpTTop0adSQauwqs/s
DxAvdt2feEJLcUqSwpW6mzss7U4UBEupEL5kYABO4x0eOnjMOaZ2OoViKzIf
rpRiMcKqKLfuLg0Clo8Ce9c8FnvaRZOytUszhLHBqWZmObnlOIe8c0XACTm5
lJ24euE/hRojVHSSaOiBAihVHEGlzs75q5UuNcqlV/Et/q6xq44buXceTp8K
8Jgd97J1mcbRzhTO1yzD+yxbuWKqW8XZxrJl/Sm5761cUGXZDq7g/QEPDIcu
xovBQPMJlJhcMyOyOYrJdrDeQ6o6e21mPGTFtyTDoBLrrP0i2BiUnmVhUsjW
oFUiNXky/OtG08CEIQ6waRA1mvSuIcPYIi3HKMWU1wpQ44JGWM00dFRaZBo+
IP+I9WVr5X3yCt2YYQAVlQCRJs+Gn80yvjvQsK+qtk3++kAIZdP5DjTvdcLQ
uzDNP2EE2NwSBsyC/e4pHiUzpD9ZlTQomPJiy0oY2Kl/9ukme7rClW0aOEgY
pjzUR1Ln1jIO9clmxhbIb9/swb1X4Wyq0119milfS8cYqbUtR34hBa+eXTmS
9uq7RVbt2i/akNOrbYV7Kipw7fLGHQ4bib+ZGwBigz9MloaqYpB9qNpBMDM8
WcsZNkbvvnMUdwQAToq9M0yi5PDJ6WiRyLDCpokSL7Cr6X9PjLz5jqt5zdc+
F1bvsQbCjWQyiSJvwHo/IvYP+bIwIkG9gbTLxfIjXtcg08w+/gGC3w0lU9dP
aVyMeX9flvm7Ohy6Km2Z9l+NrAF6huIky+ytznIozWGIPR30hd9CrHqyGDCP
JNN0c8SugMm4euALB7Qu/p/ftyw1AcTq4KdY4KznlapviON7tc+ktTvVY085
0mvodC4pB4dFGZCwd01+ROomVXf/st2XVL6YGjRHH+7cJ+OiPKNuUFYVrRvE
pKhB9qQkyQVYXUxRQOQEwhjqAojNGCeC8HrHZTJtMZsu0nbJOivtYisvcQND
+TwzZBA55GFAifbPncY6ndc2/5kK+LSFIcVk9tPDtxoKUN3Dhr6wWM5Db4Hj
HnkAUPDts7GM99noX61Xl4D+lwe8sZLZpgnuEr5b38V7lTtYDulA+o/hPbiU
JtLk9mZqcXJVxwlzLEpziGipVaZrUIxm0cTC4jWJ7sJ41u0rNoUOuwvlxYFm
qhYXdXHI8pT3ARd/fQNnUAs6JkK0TAVaYO/j9CM5rurngu9i3SbOVtvumXxM
UlsNrj0m4f+067PjdAenES7HudElzBngQJX3hI8htSt/FAkAdrrmtNP9XO4q
Wc9MNvDWmYquiOGlp5ZhMmdJ0x8tXejbLgRLzBQtlgucqcPXalMcqfTUHO26
lWlpnHbtCMH4lOjFN+21g3p75OQnQKklSw2OwHmcw57POIn+LzAl/7pkYiNN
QEwzrxfGxBAdPhFUfuHXRw8rVTr7lHc2kKSsY/MR+7O+K4QmgNPSp4wbX5Sc
O9m59iJRVFWuLnPGOhB21N/Oj7o5Mh2Fu6kF221w7siNcUrxe+jLQ6MJ5On9
EvAHyIe0krhHPgX7N7vgAMZ33eBRO9QTtCux54HVVr59wjiD9CrfT711PtXT
LRdgN45fs3HwrGEsg8PespkWuq/6IyPdBMrLU2R7imHPMIFIw2eFBodJPamU
fHHB0QCejQlcqk2qx12XznBE3zqvvOYOFybzfQWgqi9QkqeoF5lQ3PRq0HHx
Cc0DDLNa18Wd7orZPy6A1eJSiUIZ1rp878n5EcfHhRV9r4JRuCzOO+Uw8uIN
T487StPTBxN1I5BVfArbt7lCl9q27ULk01KzOenN3H0GBa4SkQHDaa34EfkM
U9M/ZzHfV1D7k8x9K6/Ilg3sLevfLD46oH+kaxk+50pLu1bhTRM62sqk7wup
o/FIN2nuaHdxYs90EeS+Z9puKzmiCen4LzsUdpjXBnYnttGDA5jmPSlnpt5/
RDf6sXK6qVXTC/8QZPqpoiIuiJlEoZRIDP5XVOGBkK7yFJqtdfCLm8XwG66t
8U0t+xPFRdhF0kz24MAZ0eGamcHqaUZ/w9pPBdTvEG282YqjF2yvwYGPUqVZ
lKSw3MOkb/9arIudsIAckKFlFiltMLN9drz8GG2Hu+zPEcnaDsU6ah5Bo7Du
eW8R3mzPJtIQlHInNvfyA3/HqaHhSZv4tZwbiIQHPKmtE1Gl1AL8L8NPGgu8
xG54NUphXmm+vK19rn7jBD7fKsxYfO40JQLzlH7CdCj6fsqARg+G+Mt9sRyq
c6vjhd/YGp7zYrcR+uQ8FwuAjqVTBS8lhvrfHYo87gPvgHeWEWV88yI3d89y
GRZ/SssKv0Ey5jycYkZ2u5/lQkoRzuhpqZus6h8uyzPIJGXndhAlr9+jmZhx
sUBKJM/NcshC6Tvr17U6B3CsdM89ReYXP2co3+qibdxPDwOl8UXxuS1muOUU
1b1znzDpd4UbIytIz+WZW0TmS3jFBR/DYpGfRunheUcxkkcuS5jxgWLOvZnG
5c5ryS8DUvbtN9XQhGLwNGRiA11Ppx5+CxOpv4CAKmhrSd/b9ex39B797EBg
l1y0lY+/X7BVipxhPrJLfgoOJcrl3PZL2+85PAPJ49Bqclatx/HhmYe+tdKU
qZ5pP96dbMnF76iZCT+htgOh+gFVfkSRQyp0gKEUo53x9vGjN0RqB+CeVKef
GmzxDIS24Qu1U1m+Na/f+8sgFEjhm/sQ7uqm+WtUvxspL8cUsPBkl3B4JiQr
Ye1361AEiszl+uev7cexzIGSfkVIejLx38/pZ+zYW31arPOU9ULtgzGMKwto
aN5eexc9xN4w8ve21IeLVzpVuB1ZZgFhKlKWQPhJFZB2V/2M49AMaEfA89nq
A7Lo5IGrbsoaNHzN74yfMViJKqDjiqyUqwP4FBbjxQp4DKHVbXaR/n+f5gBG
B9YhnfMg/vbXtPNkNOgiPZqmvTAe+irInEHeie8QTTqAH221t1a6dhUNNV/5
nBcBuwDu0ng5nXG9Nm2cC8fdoC+L2SinxZePaGxjnkjE8nOcLGJkdBdQGcy2
z5E7Ya/p2SBkXzjEVn5hrwHsgM2MA7C3sYtEXBIFJojcM+9/aoHz1F6vPzEd
pgS+Jhz/U0EfM89CYeQq9um4RRk47MH7rQXSszzlpeUbkPpDccqpX0X4P2j9
FVV9xwyZGRN8eBbklWSjSn/oT1qFCbH+BqYYQHUnEG+9pjju3OebEe/cDeyf
6MNbHaHBas4EzOu1MgEyvbLQ8482Fri1/Y7MsAi2DQ9VUXOLBLwLiYheoz1R
XcmVeS6SZqe365ljmyIyencJYyInKLcu6L7XQpSr1JccQngbFkn9LXpTi75a
P3tfaTwQozZoQnErYJAHX99uoRmpZAat/aTNvT31YhObwmWGk0AMXGrUAehP
22XWOv5JJoQfNuhKHEgpQ23jv1SJgY1yZ4EIDHGjJivK2cC9KWxpjVGyhIJu
UR9cz23f5hADTqOF0wssOv5xaFTYiFVHJtDVcTna9rYcdb0gQWPLwQp0nGPN
XSJJbTvEYxO/YMrWNALN7EZnKUy5kL1zS2PBzDP5rwJGE3JstjUNYBqcLPDR
q+XXoMsCx3t70P2XvkDRNd3PqcY+hMxTT8nRFHTHzK9NKKlq0P2LQBBBY90b
3la2VbSmQIOuRLwg3BX48J7otSev1izoCFt7zppKbWf9L86BKkz00MHDzYsn
scLLOxx8Es+tiMn39Q8hvZh4IC/z7lMvY0N0x2SUt3vLax4cFu5jEa/CFX2P
hieshrjDmA+p/uC77B2lNGxdT65UHtdy9Ar+UsWc7BL5FlbQku1RZ0TQsjNT
owjpw6DVWYsaRHF8Me0LhQXpOxUJCdXtaRvCJ7qAjBy/yIA0OjNXyY/rUuPf
OaqmTACQMvdrfp0WBmnZJc15PrjN2IB2eICUefnXNSUo0SLemNjaP2DyNT8l
zN9fpS7mBAjs3hg+AkrSqveaRBhJIFgpD++s+6cIDVRvkrNRtTeoFbWfbzy7
kpn22ccC9UByASFdquJB1pW0mHuXrjt9/Pbijtbw5QZ+zaJ7KCccbuTLHe5b
IB4SRAIgPN5efs7ea/O1750Ha5VnPSEZFtuW1HFtiM2C1z9GqQuZyoo63f48
gd6dVzF4FTgp7W65d9/P5HHWtwNcaWWGwq6C0gerhUqM4szamH5vx1nc+nFe
M9jt8JUZGwiQ7cUKxYIkQPo0u4zSIWQD22X4x6JSedF1OnYVNCJMbS/rfMU6
xSLKYXWRnQEyLIe+nCFFW3L/+IB3SDL2/TbuW0QU+FcXiu7wBEA0IMFwb+B1
B4EdOiOSnK7TpOZQ1m2+UQ4wRD4iNwBucqSJla/hRoofXr2rbSJCs7Pcuo53
XLkvH6cHvYHsENhFrWFJWMF1VpcaRjkOpNDTCXT+uzAt7SgfSx/6PvDmhSXF
Bbuyf7CgCukS4CZX4uyqDmSfal+OhF9OvomRXk8K8pyHe2EqJc1rjKFVyUsB
gapBWFnscJggZW6spPIIB0JUfmHfq1lLztSnI9MGIvKHcZ+Yf5Ij/rSOzsf4
WYERybdfVFMPFy16AQvfwQM+/P0j43Fs3VnM9PmOSSw3YKDXsPG/qV9gL2mj
wITWZGq8wckb76NzW9cfkm9m0johOay9wUHHhOZxL4JuYEVhoN0pVTIOFW1P
dv1p4gH+WTrfAR2Yz4wPNQsBrQK3s5W6k2fHCPM/c0KCe0xy3WLCtDOUlDyB
QLDCOccEOHBkwaKoFCZHsRhI12ij4JUE2lh2v2rOtfNYxxA+vpMeNgnb6lyr
K0zIGTqGkv1QEUf7GEyo+zPuGGV6HMA2RT7B3A3PDTuCZaF5pKvkowSVjuIs
Eys5m0vb7U7MUwfwBAmjysZUqHE9Lg2/JXMUu9F+Av/3wEUijvv0qrZW7ceN
0LiG/lY/7TQsxd4bl7dYw6vxKrPW/jKjmPKsw3w557LGmPllS4XB1rZWSL0r
Cja3/+ePugCQR3KaiBUdPFR02lDdHDG34t8V2HhP8ixqzJ6kfIEv2Lsoohp6
y4ihaMMbRloXItSnsCPuNEQjXe1ellbk32SQQhRaQH5ovBVAWmCwX1TEQb87
WdiMAUnjhXuWxUo6anD8F6MRLXg5VL38FSK/h9r2+DkKI1uJkPKv/uO+IlPi
H9Fta5i/DhlVgVnpyA0SKcvefpjqlPeA1pph/EuSskOpRLzTnrtrrkjrjV9g
ghEYLf38B5ih50G22zMSBaK2a5OU/iGX++PbFYN9EGUcaLCsb4SGatUJiu9q
JkjujQUZaBv2jqnEPsCb6TxCqya8ChBAO2FWCMjxN5sq0/vI1t5zEmTiL+vt
ZVIXJr9ckIi4vwj0uz9k1IYBqgoDt0Mh59HsRsSIp9kmIPuo1S+K2QwQ9mmy
Dc8x0tqV6CtZbCHkyMHtAnRwNPs+ZGXZgir6mit+QrCEWEKBWnyBlVCwTEhr
vON6xK/XKWj+FQH/j1bR6+eIZxe+119CvqT13gzLm6g7/uL1kSrrCeJN4D8h
hGnm7tIMp0MCb4IwnJ0jJrTZaNUe4f+Ab43k3aaqvad51zdBf6lJeHujG83S
Cd9vuabN2zmbwqX4AEmHyRnq4/TjUa/61qYI3iAw0cwpCHgw0GeGM7Nkc8ql
U3J7Yph4atqDswM2q40c0fvXdRaqnlLqffbTZi87Bl6UW3JyOPxTsTjWwPpg
Am8zR6AMMndVyDKwHfi5DKQKKjesebVjWlQb4jXzh3xbU2rlKz8VFFhbB7P1
XuaABgwezBV6fVgFKV7ICDY5lhaaqFOBtW73Yaovl++ixNIYEm08Ax2FoFSG
/G8eBTZjwSlVa24yH3SeuwMmo60g+0pyte0Y3qH+n3NujzqLd/t7GWx8noPn
PYM4WDpIHiqjjiZPhAeeqPKEgC2SyZVFAE2TmmJuNVUo8rj/rlxDv705Bt15
I0+WbruyGrUFiqW+eO+c2JDZLkqbd9Rp/6u6cvWcF1FY7l02w/W/1mxFGkA/
tSoTyN2pDPNKttR+C0Nsu9500XMIANApzySChO/L2lxH1Z1dwyb0jp8AQYc2
ohXd15LhZlDQ8PbfEhCRqrDphEXZlOxYcd9JTgLaqPR5fDqLFmpJ8yURbUr9
2ik77wkYncoRGy8uDx036iZyr1CietzTSZVvbhYaRgUwW0tXNGoZvlbwoZ5s
wvmwmt0KOB8u2RMLTbf0Sxb6icSjCBP1h6gmtgCK2awHx1snH23l5ZOq5Ww8
7V8mlq3bPkOPq6f0G5vApCqT7inTwDLxthk5hRR/v4BJYjl4D+fejIXlNMI4
5C+szr9QhgKYNCIYVMpgaonb70+kUkRV9yZk3MF2scL0oXMS6FMlvUUYjFG/
my5XXKqS3QtrEt91K9ufIRczoxTDFoTFwDv/d4vzrff3+c12VWjSr6OyrvoF
r9FmCOP+cw0OAbJoH3mamn/Vz/Gl78Q5l3bPVl51sTCtcgCHw1OMZEgUeOS9
LKU8oFTkgdzdG3xZS3X+fYJXcjrv7fV7K3JYg5sF1ug7yIYRfYCaqRGNOhZI
XXCPlMQmZqDtTwYhINMOp30VQbLFKznP5dAoyBHArxdswO6M/t3gtjxckhsz
/yLKqGW7nlseTbkCP41h6PafQx9lofmnbkQQ+SKODSYibPNDdk2adBQwabij
wtWegbHj6qLBmKLR+k6hn55CZ57P+fMjuO1vHWenBC1wxCdZ34hnrXviQAzM
Rfy2judWXwt+LF9QPi7OXneC9jKCxLqCJLDT6ahWfeM88T7cS4jA+zjGNStY
EIAOrxMAnf6IFn9NAH+68tnqbo6kJbyEmDzjNyMIiksU4FyuOBAo386i4wTj
aR4oLYpod/pSEJ/rktkG8vOd+slv2dKEn9rUoPy/sbnULAAotEWhS16IH0xh
iXrXGqCIREaTx/mRJH14sGHh1FzFZLvrYV1rz1bSWF8REBhfv1MkTFmxr0O4
HOQhAt68op53QC69mMuaEoviQmBEfJpveTEoZqfeeBHR9CJcXIzbYZBXm57v
RPZWSta1YfXhsUJEqRMqzvpmi0Jj3jfzSW3RlaCudMfXGXZy/sprGJ0WB0CP
eweFmAT//j/RwxZcfb2boeVy66nhkcRMGzvdvRHoC35SuYq/2Eghfl6ucyXK
6HsmemKPj0+sQWscAzieuiHwXujUDg8H75qqWfHBRMWLI5DIGvd6J/ZonJfI
57QRQjiXYQEcw6mb5CKJUwR9xFDW53bkslYoB7YGHxiVLASlGFKlK96zwyjo
5oWqYjxxjFmOlvaEL3pXTEOj0fZrDdODqbutKsZ9vUAV7mLvZvU7R4jB7QuR
XelC83BxwDPKo2tlJxoTn0/FskYbHMoKQoAtJFLDllz7LUChmW5qUnBZydSx
DFDEuaEFnS0OnI+CiQR9TdXzcGa0w3ws321o+47xDGyO8lY8n0dAsjNlrkqK
6ZgfBgjqs+UW+4dGwa1zPghqhtJCWQsACPr0fC8A3+R+i2BLvxNHMzc8vgaY
4aFMKWFdAR992o2qIxrN9jXbCL/9vSNVH9F6/DaA7jnKcxHmS7CCcJDkcc6L
PHYVyJT+ks/YIdZZW2O7okMCZhYkOXDekxlvltFzRNK+ybQFJyv8DPAJ6J6A
sKcretjZgHpw2ilFVGp4wiWkwSl7DJac4F6qln8W5dcgKTsh0Acj/BMCGs3m
23h3P2xk2b7tGb/j7kGcTnEwSK8pqmHbKqe7NwAOqpBJnxlebMoqjdkD380n
TEiUJu7UH/UT3uG4DTULTYgdD+M9sShwNxfyvAZ0MjA1WVxI/oAv30cCSxjw
mqOA9l9sS9neMLoZcD4QjwM8VaZoMmtm2HxCS4jARg0kgoFzvE+rM5CGviOB
aBj7I9ZayJzwQQZDyCsCsoU2c00/uOAK7wU0YQ8+sK30kOuUxjR/Zim3t+o/
kIPqANzOX2ICUn0m305RQTb85vr7gABysmIFnBT3JuxUykDy3/KWU43r5tQ6
Oj9c/GJKO736+NqbbYboqsuGyvE41oJ61XOtVY0FUXScyYjKrNaNzhQqb0NP
h8p0n/Ve0493cAJO3jA8hn9OMCvA6mCtWGozXRKe/OZDHHMYzLb4dRZAWuZM
mIltafl8nqrWhfaruZkKr2/ITTUM7YglgEyXYbXsevcpuBxCkhCkG7+jiIlb
aH5pBnYq/TUuS7nvV6BHSdMleNH9vuQZGJWeteD3U0j1s5VPBY0oveAu9bbu
P2h2OEg4M7rIBiEG4rDV3qgJGtPS60B9ZGrfyvBDSyQuou0eV5e0BGDZKp+B
RtsZJeg0E1xvLdQi0MBlzb5GomStuYv1QOxQJC3bx2p2zCsvt7NG+jXMq49c
UHe3+LrxgZupQ1dbU7t10NpeBnLtNxWE0ktk3SUTtL/ZfvtTOqafFpc/rRxM
Q6dz628TGDzf7Yfhsv/NrgtfLmR20UsrL/sNQPjpT5SWNWP3d0YMLOxSI7eh
dgQK7vP9baQM6sZevr7g7ooxMbmYLhwQLfHxSZCDhh04UQci1H/TR5nVBrjf
bVEt6dBsQc01R0ai2AuNOyO/wPk6imDX3R1HXucCuU7zr2d0b3X48ogm/0gk
6I3SZtRjT+6XzfK3IKfm6Uc9+njgUK5RViF2Wbw6gs+24LNXPVFjO4EOa3qq
QgV2f3WNAowEg5nZwxL59W3O6bbbEq3Q4d6qnUNvAl0w1XJZmsqNcqjgj0Hi
nOrFF+LBmmW+lcTpwP/7l27BIkQZHTkOWIsAsO/wRTPrD0KwlkFtHLFd3onv
8QFAVT46CnTNhIqKzdjdtUGAfFcs2+spBNjV8JvO6yQ6DlKHrkc6MgxVPZRm
5EWWfE66u4yKBpZteA4XGsuUXMPmVi8DSDrlEqmDIOeQNJwqWLwa8AaopPjB
aiarTiIATRdgiuNwwH4Ivd+zltzYlJg94fx0QNKsO3+vT9nDTElkowi2hnep
kS4xF83w5LR1x5W2ByIl3fmn/fgg9LmHzH1zsuGB1DOXYG4oo2dy+Vjh4JjJ
0m0iUsXzhas28lvh53vFN1pDWtGX+ST05+dEB3INtXsA1p0L6zUfi8KK5sPN
3bizh4pIzCOJmRWjifgDSgYMXrWRIcZWWWipQDErGvq0XOs4mWru7yoJMvFZ
ZY6SlxG6/lBxb7ybXs5ie3VUEm0cz7YJ6XUsfKi6egvWqy5CQ4IDB9GxxyvU
na1g513NLGlpvoHhT6s92jvQ6GNVk3R80KbhPzSqkPJFgcf+Xk+L4w05nrg9
fA5Fn46PNeEbeJpDJzJxzKAFUyZae4UptehqKfjzNB4WL2ugVLw8FwCxXwda
pRmxO7vhkNrheIYx4Td70nvo2cT/xVw0JSlvQlsvFliWHzcjLTNFgNApAwJI
ZfLbAPuYu7jCgQN66GT2hp2tfNOOcRFZHRi4FlCyykKLjQvl8aXcNMS/Sc/K
0aL8F21Gs1AxAROOXEDl9HuSmXr5rA6VRYhccUYxv+kjVC3yDRC765Fi6jdX
oKxOXo59oGS+zEntsyAPid+5Yacm8vok4OJwK7iraeR/Tzgv8lqLJsMKTEQQ
3j9fg2OnrV59zRtYmsrlPhp6Wzx1BH1Ke+ZCnUkTmRNaNWR0gmNBOJ9FyMQH
9uhhrdRWEFw4+X33kbu7wBbM57kURc3qkHo8tBHnZbc/uR77w8KO8Pz83q7p
IXhmC1VYY8jCh9VIwEE3QAdyeYPXuGiLPh5SPuT2KwH/UITWA3XKnlnirtLj
LpiaovtITA3wfip2nc41Pr2fyoyZxSFUT7tBbZjLy4idKKHvbOjJ5XeTmyB5
KBY3WupR+YmsqJKsjeqPJ0RoM+T9Vtb9fln13iotoVoOnz3Scnw3jfucYq8M
B2zBdt/FVwjQizD2G9TdbzRh86QZKcbDbMB4km3HN3XEwBur+RVvnL9RnWiT
5XmYzzKfsqA5sB5vh4RWwEHDMjYF69xaE52m+EEDaPpC7oReaEZMT44/m+ZK
DL7icxi3AcdRzOePRFeCCZHE1J9CRZbB6WIvF4chfrzRXJLmpxs1NRfpu96m
G0Cz/OAsVd0zLyG9n33+2BhPLiMZFTZ4CUAD445SkfB6g51scGHKfD1tOGSf
O1iUZBpAy4A0rAeafwxXb4rZbMkaKgi8R5nOBIGjoSFyzbMAHI0+O76PgGjo
MKl/f2SvPNJ2R/zyPRIaSVFBGrBcD3iEVOc9ueXmlEhmvjAm0wnHOm11zCkW
3QP43BiWGwzN1VfWfiTGiHvVfTf6NyePyfA43LzEv6E6AMxGQXde+QexrwuO
kRr4RSCtfL+vLyYO+QVKZfRQ8/u43HNr7qWt84AFbktFMT/bf1xCd+QoCGSx
BCfOGTBIyY8zTpPIpJVis5Pxv22m7D/XZUbvO5mudqObFJpy3EuJ9aTLoB11
OUQnn6rJDyUgcIFcyxuJ9hiKsS46uK7QYVOHuY8w0esEq6wI/Dlc+tIoxaqn
lT99s/iCBKeVuP2FPeMVz7W0QbEnOTOARKVhSdt77pWNoTaj2PLOuepQvHR3
3Bj5TK9veqREXRDykjhhGrOy2pOiUE74z7WvGXMUxxUOe6yecoXWrbTo7eqx
hfKiv/GmoM4tolO4Ft1aN4ZSYVgrCISzsX3erAh2buPTVKSRCtyqykFLQNRh
FpSIM7FuvmI9gohZwb5Yvk5AXfH4rWwyH/yaEM5z+UXlB0PsV5qMpEiZz9Pw
vq1YfFVYXd/OvNVy+5/crpQURydvwKeR7Fhz+U/re5AeOp2onbmcPd38Tjxy
GVX16kwxyPHqbvrqMg0W9ordlxH3ulVDsI0bCqkCQvHnJTKW0/goYTVSwaeQ
Q6k4clYRpd7jljv6ouTDMPcc25mJeFdDMnKgMurOA3IEvxLlJCVswgiB/tVm
DUNFOKszZMA4IGAZGh6/JeAgt3/L+NAeT/2KzDB5pfJzBP56dXLgIiXS+ghZ
p7xizUbTYJofx7uUwNzoRi4AC5P7mmhcgrQNw1I8a5o/oO0ty3AmKytu9qj0
NkKVHzdn5QowUKHXrEwirQ6RfOG64MWkmn7aonHSDgvjiYIT9I9LIWJ/+jOg
BtRCfxy2I9GEGjtvFVIjzE59/RWiXFJMhor8++y0plhIe8LJlUHNwm6P6N2B
X34duOxAPJUPr2Q+ee3C4NYCzPvcj/Ay0Y9e8+Y/YfHARa/UHQMzJM19nyeZ
lugvcNJn41PeyfsEtVKfmj8m9lQi3GLgqWU3ixmA9IVxuFS4S0O3RB8YByTw
uMgRmyWx187OqEfXY+M7woIrJWId1O64fNl2N0y71we4q01cyvk7XtVsGOUr
l9AgaQMX4e88UKwIicaVRXele28nlmSLqP2LSdXqvonNjztnLisSaWUjZ3cN
AXDLjcXsnnS3Ahi8N85rku/lwMwAAPXoLREPqSRy22EakqnA1x4UO8Oj6N8s
HiwFC8jB/qubZGQwJ2LYIYFlx2FwxsCh4fceZhk0emeuv4E0DgsczDrn1LLS
tc8gijEeRKYteO627CXvxXrTt7emlb2dPeMWqmFdifC6fMEgal2h5SIbZchn
23IX9FaF2k7ok0ctF/1pXJh6igZw356OYXr7ckEZRDDg8xphEozD30GCBfvc
fdR/FJTl1dWI4wm81QhYgPeqH1zmLjuAFvcgEjtJZGPoSskg7GGd62ByZVwU
BdLJdRMEet9+UoTHJyO/6nxp0oRA79pXsiw460y65rBkodnjNCXp6uXnBHa9
0/f8YmdGC63GCXwNNAxSAxrpA7XfDbpdeQ8v7KhV6kya70qdY/JjAY5znU8B
uknKYczBAm165FhIGihTNiq5TSXb97tB7cCAPgfnuq3XGpRX0wr+jncsSrDD
MAeWDG3AZsrjafiomJtGcGJf8O5Jr5M9hc2QSh1QswBzlDiJf5yoQ9Wk5+/1
yxpWx/SXCemhor4aeMvL5woP5y1mbrpcuPzHsro0EvNU+uY5YmPyG7Hjodel
6ZKLFTHS5qU4rMmoIbpUksFjI4NIk3fDGJFwrTabqk0N+mOFSpzXPU2JYBhW
83X9XHXaI+PvPxx+Rsxox3+V6Ogqdiqk3U98YKcKJ1N2FM010WDXE0/zml5c
GcIlNBaQnkgcxBgzl4XslbOQw2k+2M7ntYiqs6GX4JiJAehgeScJHk7dN9RA
FZYrRjkulo8ZiQg4bGcbPg6CeTWJSHfM3fMKgcf9s3M0WrlPn2An94xyxPxG
9IcC0gWV1Ooirj/n6AxQfeig5WGXR7e8aADo2707JQ/kIKR8BDEVHw9YTUqG
zg3hApqfKVzgYjTmNOR0WQNX1ib2/qQXRf2mg8dZDha6cnfAiEply/kLKbDx
ptFqTFvGrGfRpcAgPNHBTKWUad0ZeZKj6cQjD2Y+7bFZPV5UBeLpRMJBWYFU
/3Tr4ekwfr5hrRFfJZHujanHmHpxqLCB+/zgAgtAGjvZ4oWa5YamScEVud1f
x8p5gbIiAp6dcndZCuI1593IaJ9nvt4vANnDGwzICCRZZHi70dFUtrzZHc58
vBvDY4jxb3VAqEuTeEqKIb9f8OmRlJ+erZjvJlX460w9ULUxrE5wXx5hjlsi
I56dnlY7Yd/26FDsPCowfuXnpKG8rUtlorQXaafny9ytAms7ne+L0nRB7sr2
dow8uZGGgdq5aJXefsoDRzQVs/zt5lRjmN5uXW9drhZRU5iZq0/K78k+qGz1
z/5nzlndJQk7ft2p0MYnjThgsDBCa818sjftKqDkOYRtugqcoII/jKt3m5Y9
hdUNxsiJ93Z27tBLDryjTf9fQQux9SObzN55+RR/ubj6xGxcpljn2nujN/+D
fOqsiccGtG/58FyjO3Kvoaqg2om+pqqXcNESSbiluRwS0uNL6pUHkEcp46uP
TqmZpyXA4o1Vm/V/kWPtlF71vKW1T/KOTCpaTRm3BeE+VnPgZBeUEJA6cVx0
sNXZ/ehawBLgyznXVb3GFjCZ/ZKSFY4BurPPqoxJFM8g0ig1JWLg0MYnvkta
SMAN8fkwtqVSnZ1PehaFcjGJxVRN03Dtgq9pb0r1Hm/XUFMb5jkPgDlQNKaG
3U4F9bfzwRDov8vCRs3RKjbMDy9PbnEJ5KQDiJCuo4Lywci3OGqfOa7MwfC7
7L9JJiJsLXKs+Jn62NhZNG5m5tLGppRn1WGM1jFWqTldyd/Yz6ZrtKVDDIC7
KLANqKVBTIc6UFi/q0CdtwAXds4TR0qNte2/qkr8/hIjxtwYFo5TlaLRzqpS
7oyZWAriIFWzOQiwekMsnS5A+Icif6+QWJb8S7fUwEyc3+3qac338AfdaFxd
XvH+7pFK9MzahxM5WopxmcNFTsLZ2HPHvw4bgTSDThht1OFx0VEEe+81BSB3
Bq0nfElwj1jWSw7NgcfWgGbUbsJl99m6T0kGNq8TuTsLNPG6u9i/gwDzYctB
Vkwdb5vMoedUGh7yMQZehn7PlNbnHlrD6uyHSEk7a8W5IwmWfLeHVHhegv4Y
ynUpeWJjej6nG6cu4B3jClWAThwIg/ZN0jn33OcA5rP8h5BLUTYPLZmdRrNK
Y8MSYX98Mgnk6jm69MYrtsQP+c1FlpHXKvEuCiE/oC26BOIrhnyYLA2TawyV
/PozfJWkUa70Bh936sfMwlaQVOgTTeP5I4qC2btnkQumMfrKH/oF/KuqNHYG
EiHB4nuecJCZ6DenCZYMTny30eRXxRcM83FjU3sJQIircm6Tw/ALsACcSWRI
hUfmMFep4BgSWqxbkcu5BxuPPSa5xoCOc70dJ3Il9Z2kuRK7Txo2w49XJjNv
YL6mq0JER8Cz8gvZDyVMPajPD0s4Oq+AszozrVESYm8orFFXxrOusvIoFTjW
49/t9lXkGp+s+O5gH7qPK7bzjt9b9lQfcL9KApwhirlc2gKhxKWw0KdZuNmd
60rSqM1PAbBuXwPnE7+x1xFGsO/ciyJnSk/I3KeCOwr4qxddFAx54tkkKBBM
b8kXHbF75fhL/h+M7KncjnYhDg3fRCHNudFxAFVGnLWpk6RdNgBs4g19N0EQ
hLPrydmYWv3TDB6D3ZOta/M8oCRVnWyXYklPoYkPgscIhNc1y6f1243aRL27
pRpLPzIEOR6oDCrt/44G4aLD7BHp7wJGM42Ar3NBJm9vOtpGRDln3slkkbof
X36dIBH1ZS8AIVHOw27sA+m2ynhQfbaSpZKzIIPpcMmZOy1ADRyWKuq2HqhT
0a3uDjLkE8n4ryurrWo6ykrKSOeUn3qAZkIWzAQT9cYIv+IAU6DFjhplB7cp
flXUvZKVn0tGEHoFaF3klIhaLJ3a56y/ZrpCe321DtY2cI70KCt2NmB5UuiU
76WtTk8A37K0jyLTGoxQXuQOzuE7+nwHqE29bFZ4WYemk/k1XnI9t7Jb9T8o
NKyakgQRf3XWjXbXbzMpbib0MkK6quGcAiysD4g06jPQJlQtA1/Kz9vZ4lh1
1fUEsHZcbUMFLDciOGG6RtoCfm0Uy8iDWMgy+/idnucAr05JVo4SxrQ7pwtN
EGC2tfpMTD57d82hUeCtdLUUXPv2L1Ve7AXC91gD3xPf/bIcoi3/OlnWYVuM
Ef54N6m7nZq/O1Daugqr7Fw/PXahnwc2V8jxlri55hgXbKVfJvtTh2aUkdsK
fZKLpGcTXxchDDYgVA0PTdF/xBXDL5pf+3/EEN/BJO/2/SGy4nMlxvv8WebW
YgA1d29gFikC/6enL39PwofJgIhK1+Dg8/5ahH9dBWGnmXrsofiRn7SOt6I/
y1aNE5Un7P4j7Jdhy5t2Kpnke7f9zFOQ+r+YaRFdsCXpES+5fNYVofzfKBfy
4lVj8xbOs31orB3I5vKTXoWJ9/0EUcMgAxIbDkOvWDqljTYBUx6GWItaa7HU
OxgcknRtu/q2UURA67wtSpFqieG5cPkVbrtbJ2YYA4VzWL2w0S5tmhNjpuxj
ljCnK8NB7wkDmb7NDhaU+qCAohd+HNIfB4dDcJE9VHdUeUb6IwbIEBZOrfo1
fiPiZ9+cxNX6tKhAu5ulq/2oMMBd5kqHQlwLoBoMinkHTeRneCO6FloGG/1s
U9Mas5uyEl8kq77zOp3MooqUp8ENSNAgAhoX23bgSAolRUV/xGYnAvcaDPku
u/r+zyuC3eIoWIy69dBcsMyICPKil1aBd5RLNrVyUhR3Y1SY5mwzr6+dimq3
s16u7sJ0wtRjtJf9RlpFdF3/H5tbm3xR1Ki5OUdX6RY6ApeBEYKOYGXbGQR/
ZXnXBKgzhDVTJjq0Qd6tcO0BfxWbV1elRW8iJ7VZocWnIdgpeNY1NINtZGRq
bDrSLX3BG63ovsJLDZ09NDovH0Dpg2HYBIeZhY4Pnwaype0U6+JsurdJrD7M
lMT7t/8iBAX54jVJb36OI07elvv4nXI23/PysV3CJ6zFtFiro6/i6K3r1T77
RDID/iiNJluX4a26mFWhBLv5LNTj4SlfeBm+d1Qz4g2zGr75hClKc5LiXtq1
KOg8iz2qFGL7nCFcF+WmvrC3teUnYZVw9ReJMQRiyXIpK0poQxaNPUvfxFAX
LU4PmAqSYu/H2C5duJvFlefuztpAftcaOiwTXBbcCakCkHKGavq+IPlwfeyJ
wHlJLYs0/LynPR68nwppfdskdMMB2DlejfVi/fFj3ualGiyHjLELIlWbIIMp
ppPYbWE1yXErSnFaiMOj+kFzh4310NKd2WeQkLepJ+SkARhRJR+5WbQozmnI
O8mNsrskT8CViBEg7ZSVYY6rnMQf2lOriCrEpt5KmfP7TuYkQniAushufgTF
of4GdhW06m59DKfcA0JSMUvJyer3sL6WaF9Z2byTExAx7YGfMy5kNgD8yL6i
g2SNpKOmh4e7+wtniLqBBxhB2dnVSL2bDarS7O0YOoX78UOvml8X3tj9akX/
UthNcb9jyLDaEOby/YRujwKi3tay+TXy9KAcLwzouHbxpFmHNkjSJo/x2ynM
kMfyse6aYu68rNBZOoQlBShl8EtBFkYgLgH9Yjvy0pW/TSxgfNLbnyZRhVtg
tHO9kgOmLGPIj7gKB1eUp9dOnQSMD+e3Yaoe1nNaJiLUiKjQbPPKRpEIfUjW
JFPOBJcEoig2tqILpLDFsU+iTvOJsRDT/OD3+/F4+5o1/bmbULKpr73qlhHa
XLI/94B47Ex7ORT3jitMOt5gKoA1SX1GBClky4HC2Hd7AH8VpQFxlFmIjFAg
sYu9xxeZtIlkzMjOIN2u+TDDouRR5qIpwWiYX8RkOI2aDB2RGJYxN6JlLOx/
e3w8A34WGTOpTJ9mHbItGQgr/nguCyY3dTv51SB7x3mqEJ5JloHZfbzqsApe
6EKmT+/IhGroWWZQTePIEHWTIjpqos3ljyEyvMfUa9YLM7isAzECRgtJSSd8
2dD9Mx+xXB7DTadDo2kknbcLcNTQ70lj76fT8id7O+opdeXNJBuwfK+bjOiO
m2lQm7T9sZtQETIvB6QRs6CgenzBS69bW/v1IIwDAH+XgO/mMR3LcN1BjG/C
X2H4ZqWhU8/C+FqaJY9js+8xXMSWxsNWuwSZsaBxT0sN7ZPLVNHXfMAA+DeA
1gz8v0EFXaMjYPLB9UctbVZFC6RW3ZxrjzNuNEBoGtWAbCIxdQRY68ec5uqr
zp66lxisTZ3U53MZJ6h03Ad3kN3TvL4e4URcoKIczANdGYmHUGOBhxI3tRBV
qL00HuvfNxGS1PD1PuIP2Vf6NAe0DC775/xOOVQA1neB7xIiLKTks842OkDZ
dc/C9a+yTE837WaqMlm+f2yh4ulrRgV6BtHggY+gEMrU3RZjvr8CD0bp1HMM
XDtH3afka23GmpqI2OoY8aEmc3j2yL+AYkzE2ag5KqG0BMV1yOyllTGbYJbc
1W998Wvv+Igdue79hYgY25Uh5zz3hb4vBbWVtDisyauMuw8+ZHeXm2gthu27
UGMGBBjkyeaedh8eOgxXx6D0tl3roHnEFVSmlTEPjWmfECEn3QL/e0obhKnM
XlGjTMlxKVKIxu1zVScGHUtYQoeDmlRUtYpEgK5n+8nHjlLtHFtZcBmVhlfp
qEoIYk3i02AScrjg0lO6azS/h1LDUaGQ4dAHf56uix4RKTQpsfFePsDleww7
utlS6BMlYOjVpoXE1LndRaewNHEjfKiOfPD6LVp4HLxQxWn5SgAcP7AS4Btb
QWBfpApmVRMIdq0MwmFi8sNocwMD5DxGZrCrqcj+GklGI3RHhcnAafORkkja
UC1ktZEjW1DoERdcRI8ggRAIx8rgbtWktRqYtdKxgCwfSpk2Vj5WZNRJH60X
clSWXOSFcA8EO0pD/UgmEQxSAxFZWRqDE0yAsNwDJQJu6xYyVDCQ7/PXLTVg
9zAP5xn/nKQvnzdz+JhEpkviJF0PIaTopY201uI1rKQBaHHK9J7qnEuaVj3K
yORVEQfx6Q37glXAtWX3uOURz2GP188Zyb3WaRJxgMyZB4vX9JJkEZL0REju
VinOjajmZyddWISrYwKcwhGcsNu3sx0E0RiQkK/hd//mht9T44dds98M8FwS
VEIfo3Lb71SOlVRn5EsxyeEZgOJ4eDbgbNSkNA2IX/8d/2lF1UjcdQAQAShC
BqtqDvQhHKjDIwmYkkdcaYH5WMBJQnAHK8Og4iRTjp39HNfVa/Nsm8fl7RQ3
6XdG8Rwlv3IQi3XDIAfXtqORzvVxr9U7MkEkOAG4b75NCNjE0PElp0zfRdbx
GhQKJvSlHr7lN5f1xZiREa1FYfjlx6cHUHpaSoxmzgtjWPF6ShkRT2c/spIC
hL6sdSZLy0axbOOaoxFtIpHLxJEiqeDILKbfIriklXObpEhz9NyzmhTMJJhf
y2YJXO0Lw2jDgEhEnOz9V1QM4vZVhd8nQwOXKr7hGKk342BSXV8CWIExP183
UPI7ip2WrRhnnhkqusHrmKIGpECfJZ03xMo5/6RFpj3zMPn/+mgz6O/A0yrx
109EHsr0hRNmsqFmc4sIFjC2DjlqB7PUWLNph+R/VvkyAev6Az9zMKLbqoOS
UEy159aqz+s0MOytLQVm9MS10iEqRfIXA5y1NgEllbaf/chvIpXHKObUOn5K
vzbt+Iw0ABjzfHskElXGdpxZYwSrbOAklaRtonf3Rm9SJPj+l9ecOPKikMYY
yRfLG6LSV/I9z6+n8NcpSuok8FLZSBLS8/wb8IRe8taVB6235IvyVMtddl1n
yWTnczbi0GjHCVjaeYywwErbwaph8xhwYosniI/v8kxf3IbHyJl8fqdQR88O
uw+rBA89E7AEA03beGTsbjKBI9f4stqVLQX42u30tn681+4l0cPK+cXFM7EO
FJhyAVcVPejFPFcdSUkaoRgD75d6OvMkVPaQh9LohGyuMBo1krhvYI81EAuu
FwLli85oZN50oSo6W/UIDLWYiDrxH/WcBjtftVnVrnsdSXA4TquMxQ95pYk0
2hJpzWfo5sUu+kgt/yNj+yKYJFGo0W+rbw7V9xz4eVcN+95/qVRnjLS7l9ju
g1/v/xyZdnBD8IAFHY0SAv6lYwU/e5fVAXj9OX8VaVk0QHrcJTBxJyaPgRia
sGt90ZnUkMbBBk542WRCQiHio00zaFFKdUAc3OCDg3mZiQSDRfo7RqmHOD43
u8gAgFJJOy+f2c1Ll/wV1U6Ao88yXtViFMETBecxnzR03jJDz3DJckXEsZXS
rhP5dliIY4HDoHLq7jhvD4/wb3XOFex/poxEedR2ois2isGbOa6UEemy8LEs
/QVbAv1AAw+w0XJ4Rhq86yzJlf78zjVPtwlfPwMR1kv6I/DO9INbfJZGeTKq
UVYBTbQlPZ0wfVKxeEovlcGnI81Uw4jgYCZZzLkXITwwQ9OhoJTeZ/ms7a6U
RJuUMdri2XPgKVCEyRueYmy2svB98x4gnpBUOR0pKJCtfTMQAxRy8sXwqTJ3
o92cDjE9vqrNsR5TLQHUqFadxzu8xPwHXjdhmdDTywVjke/KlfTsm5+XK06/
97dGkYLvHZ5sGxjSUt/bVX7jtPcTAnK3xbbCSj06ELi1wp/Fa3Q06VF9gX5Z
PYoEh2mW0VmFe9LcF4Oyr7o3+b6FJEvHDQlHMo4jeT4lLLADEdAUlCZzeZvS
3+Cs6tzQqgjSRKB89XMUkS4aNQlKOpqJSCt4F4r+pXoo4rqXLloi+prP1E8j
1IGgfFMYWRLjU68FcC1aJmBaRRMBlRi+L8wsCX4Y9Ch0fn1TUTLZibBstiU/
SmrlY9YCIZyeHDOz0ADNF6xJ/y63KtS2E22TQ1VjksWWuzNp4JXpuRlGx3eR
9odzkbrgbOWm8QUZRwnMd7fIkZZFh/gKCSHr4NCXd2h11ZKMMDPqjmWqZvHu
X0UTOPjuS5TzvrpEHfYIvkomYs7rs9Ztm/aA52xhvCzpqbFxi1a3oQmMkMnw
tA9H0rciT7eefS6TD/P2oTorhZUxbHGiCChiOR1VgGdd+bxiHz3eiac9QrEP
T0TsBNL/tjzjaOxDTgyY76sNab5ydiMrq/fcRdV5HCc4dg5rXsqSXW0rTuQT
6q3vaRp4CLsMfpbNVMHTuriczxV3JE0YoxjmpmfKZ/UNZVRuQd3BwYn19bsm
sogthI1a2HhrZrGmltZmvzEQPY4ktbS/H+1LJiXieKNU0aIZRB9MYwDjsLQX
Vj+1jaheyyXKjk6Q1tG2oK7jbSqmwFSCKE//eTr8objAUwgd8tBRt3eeTOpU
8ADx2D627AT7OTnWIlB63q+k4iX4jyRt6z+xE+IpBsQKeixaNr3QUY0dmJWi
CjQevq9R0cKu65jbXxs96ETurtHzVgEirjo8KMJKMEx+ek3TFq0q+JRHJ4qW
kheC/KiPdIKc32ZleNOZyOVG70A8JMRO8173rOjSnC3o+BQY0Zm4mjcCaWwO
kwgzwCV/HBHD9T297TnFUSaF9aZFp7K2p7VX0qzl6C33fWduIQrIw1WeiCOX
vxHseBtRp6EfH1yGrgiBnGSQv9+HGpNdjUgCxbqJZchCSa36xZRXJb4gqxOI
E3JMJ4sE8qrsfKL/yfjTy7K/GU4d33XR6ZpGPNbMP8z5kDJfuoDCf0mLsFy6
bzFYZQI3///l0AmXFn5z1hZZVgnr7cygGyPR5l4VGOsJajCqqe/VjS2abQPx
8HjVq/ZUJqjmBiv6obYpqru1o650LbaltTLbjC6NfAC9KFcNp6RRs+A8N2GV
B7T47YWNwPxpme57sp4FGP4gvZ9Q0ub5Ei5fLVWmDCSRPXon0+m+A34nZiJd
p0c+R8N9M16h3XRbJ8wu0JO4/AZpefRayVDvS9sAJa/ASdJOnk748IRiveAu
yghl8ofQTsVE4oUNWwepQAcyWN73z1vLWavXA/K3wfi+C3luunpBXdW92AeP
vVmCJB3gruRMLSsVacYx5x9ujFUNPwdzBOm3jKdyVG8J0fLwwON4xzQlQriG
4/of37jkCIqd42QGYXzq5HxXGTo1juvEt6gA9I3Vwue//31ddgYjfzbUYbRr
q5cSsiqqNt1sAhYGKTZ+/82ASQOFU+FuHW7CYd7/XOzpz9vrkbPIepQ+Gdt/
NzgH8r3Mw207P5swINawXtw1UNqH2+d24KqVwWFICCj9yJhXWfyAe0R7wWTT
H/hxDO38sAQq1vrt3z5CGwN+lRkJkHK+frfQVZpIj1zqZwh6A4pQUiu8c06z
RWFGrEQIxghv2JGhlt856mgqhAxxWiDzigBoAER2eCPI9n9XElK1EtECaOVt
A/gIOC/NdkKsVsUloYeqhdDzpYYNzrUv/QGbjaQVjJn5D7RaiJCgcM6LsG5x
wTnvXEsuduiYLYIxuNnY/yWo8NBd76ZEspME2JYjpWXabMEEh/C9iZN8lR/K
M/TRCwE1e5FKJQ5ZvcsbvAImvmNhY79g4M/cgjDCiRWdoY5AW3q2yBAlkF/o
D5pwT3XLXEArUZ2g4rz2X1RnJ86k2zK/8wuS0ODzyo2UBZB6kLRbBloHJkWo
n2B7x5sX/Wa3VwZH4adv0X6yv0q1LhdQ2xSr/y9V++fk41OpzgTEZ7zTFX6z
BnnXm1LaYkAGNmmG/G6ljaEL/oaYmQTDgn8izFCMjbvtEuwfQIguLvk2x/jO
tyBrNIevsbXQJgQfN04bI2sSw0/kUBUQxydaHLXDOSSrqfsoByJJlXirEgPR
RYDUUnI3VguREJDbM7Po6HlbCwYTlZIW/U7P7M0iWuHB9dHvK1nlgWhvC1hW
mWnMeUoJ38VIHgqr5eqXxaF36K2dif//4YI+ONlNclxCdsDD0ABuT7frgHdx
X/new3fGNuU6PR4HnGRXQUSNwTnUgA5CUkW99lWQ2XNSCdAjl7/+59ZmbStj
FzPkjfyRnZIKznJUCcllg5bsO0rgmlx0E9xnp035L7MK5+HRj4EkXn/nYo/u
5m496aYGTVB4hWFrVhyIORBxWhfpXPhjEq/cLmnCkAzcV+8sYFepPKvAJAr+
ipELshwXu5YI7nFdkBqRqeGcVohRGT/Kh4yfWc4D/zS9uEqNb6W7MFMDmnKp
Y5tq8LsrmihP75hEAJDnxSV1gr4kOsTB5pKiEJZ9/pmANlCENAvOWM+rqka6
Me19Zc+idIazX0nxGlfTTKSw09ejlmWIYEr+qFE6LQ1hH+E0JzB5FMpTMO5I
io1dw0UMpjSK5nluHArQDkRH9NIGdu1MSZMEZ/pb8xqIZEtT2NKzIAIz6Uyc
2xWKAvMr67RI4BNf6Uhr+Sh2EizmZbU2VyF6Zsvb5L6avk9jIh20UAnHJ2Rh
3tIEFeq33VvGJSkRu/yHAQhdrWw7uyL2/w71dUr1K22qJIQClUUfnG7zSEPQ
ob0jgutgVp7l2LP3M5RhUgltYnnJxyLbT/UPTKQrM3d2KSvyDM29CC79wxDg
0oEePJAM3dKNlivaHWYPgy5lLt2YODS1lFQVosMvJYLw3BDh+hHBb9rkJ0Mv
jF0uzDWwHrLTB91wkUUls+KdpIFqvvVFmnUsYlaSLWqaJASdLToMgE5ED95C
JRVzLJrerpdOOQhMRjtLSf11V7pO2COCyoqNz3hp0VNpz9qcs3Bny7mYkajF
iTn40ty6bm5hClB80rdGGYAddVSK3qqrtUiHJdXx+pUoRS/N2vwfc2hcFzcw
cfhJoksLCsbCS08SVxprtBNGQazTuZ+6Aa0YA2b1rx5XeOu5F3iO2aPFt0z4
UEb4klLX+bzcj1kiS7ezhJVGDDyKy05PlmRVcaVXwRIDHayuHm+fZICCXWPO
iUizLpOuE2/33WC2MEdyHTBT9vlHndLw46c8DvWF2Ruatp246h8kleGOmVR2
2pDsKtxqqk700Y/2R9MsJsv+1xiMf756sDSi64KfM5BQb8YF3v/nvawvOf5Z
MUHviIGRyXAYmIRE5qVX5Gdadh2vgSG4jrA2iSn//qBoJeUu5DOh/Evt0A9f
OzRLt5UeJbfUt4PgxSbofcWaKLvYUdZ7kDmWROf6rmRLv/2looMhNgLXpb1p
NKCvkaT9WD1SE1BzZHoMzgRd4VvUeEgVDDd6XhiG21SNBy73Laozadsa9AJo
pr1/RfilfIJ86qSe1FRZA5BtCiUmxQc9M3Rve50acSaBgqa8D3hXxvYxI7hh
fPSzzg5SRzqVQ9HPiI0a0Ox+ZNAyjUaGul+LFaFNznqQxUjmM0QLEoRr4z7+
At9Y5YRw4mEzM13FwO1hOIMQwmiJ0xgcM4fhi8lIrcyyoslZft670nR5pXH6
6Hhl3087wU9hVnbbCTAYMQ7HiXgbjMnY5/FmTdZoca3Ya+VbvKT87uAdOdX3
dvHnezoV+u2PcfbGvCV1knFgCWYv6m+FJlfc34SVMZH1ER5wQmuYUX3zOgWv
cxXEqsJ5fay2CNDm6O+Sww+72VOU2z4e+13sGwN5bgoM2wJrIedYd5hwFpbx
klCG6q8mXYkccLsA/VAlnngAmmQVnuCb8p8cmDmkqzu/stBlmSwGmCmspT5k
W4MLzA3zzX6JhEAxXa3ts5MOx5V6lJdrY2NNvWqwqcwOs2Mea32QijLCD8+8
tqteXrfsehSS+JwEDejHryLTBPl/45GGIasUYbQvdhTqeDTULM5jMDmaV+hE
D9ESUFfZfPqvvka8GlzPuEsTwgPAvxLn42GYdLPFZt9QA6/rPLpAyeOPMTqQ
P08MoSE95n+2RKIdvRvDVZTWvAkiW2KJuAgtnfiyrHe/24ug3PvkhP83plTZ
Hepy0Cm34mCjiYs6zj2qRyNGjtKLjK4SmIU/69wbQBGu1gEdP1d6FcZLdIce
B5dQMQt72b3wrxO6AeGP5w7Fz1pmP+f4Uk7Ly0J+5IMbB1HC7yD8J5aP7pXR
MPS6eYuCvshRkdSYLoz8dhmr6eENWIxpyVUpILYOtOZYaDkZmRHNFzak1UvX
d5XVKPG2KG4JP0pqlEDdAbKyhLuEsUEq7iFZfEsq8nzIgGU9mXDWT2SS7Hc7
xz9gv9Q1Td1VUbYwK2m4Drr1MZXswMXa3BXZO9/DmVa59xrmMzwUqAyXHBQ6
tJIQ+dgzH65HOtKfdB2jAP6/gMcO2qMpl2PpAId875BcDd2XgA4daftMqldv
raD4PyEJk2PDiKO/77+xqcYJYHu6XhtTpT/CKituBWKEm02Ul0PtFRZRbAte
o9COpt4MjdJFw3EbQ6/xODtIsGB6DNDuyAHMdwTRsg1E1jI4EDcIfVGkuN53
dSnzBTS/Q3MlP4S+QW6JWDTbZKBbqL9ZsEa3TL8vRodeBF9eszodyRU2HGGG
HWGO/Mvw2GwmGCOa9KTvKh1MOXcP1owcBsUwPRRpwJItMswLQVKFnGZ89O1c
e+hKqQW/osCuhx2jqRaVXjg6gHe8q6g1Vt3YS8fkkkaij8B9NCqauSMUIwLg
LsBrzCIojNZICuL6Ac0n8T5mt8W5JcSeVgpFlVtyBDPhpC8u2yzq8YDV0k7r
3UqObMpAf5TEGD4iQWrwDtrQzHBLTACuVSAfTx75PvG92MwNrqQlUl2gv3Rq
tBAlfdl/V3w+eY4UtOmolkKn+9HmIsvn0DujY6pfNrIiwSRR4EsPPfPUVt42
zPmIRj2WjvOYVTon8aghNjIuPWBzX3XRovDY5BvqB/Q9OBypVs2bq6tab+7k
5wimwyBwVY/CpX/3CB5G1oJFvpuvO3i3rAeLp857ZfjGDU0YzuvZPKnjt6BX
jmjhUiVNHOqSEYPxReYDiT450U7O9s6WCq0HGQdX6BJDD+ZKyYh/NtgIfK/N
N8XISCvx0HjQWQuM1xvl7d0TxWnBt7Gx1ejAkVU+wOQMuCoOn11rnF6XCgFn
Bnkdk+AWbgw/orcSH0EuvQ0vAItbuOtFKwUQBFgTDOvwZ3MHFQvRfty1fquP
QeLPzwwAjilMESs56bJ/KpCkFu3liPBZO5ipoWvEPPghl8c61E+1622I2YSO
sCKWjzABT+22uevDWD0AxsR/FtlLbyLYlTtJtO2LMvPli5lPvFcGuiiCUX+w
RiPxQHVL5H/XzNP++x1PPW1fPu9AWqAcyF+LNXfu03vuoak0Nqo0U+PfEPz8
PKEo2TJkAcI9QnNhcchd1auiKScKjhJJoRh7c4GXEkBx/7Ce9qDM3Q3jOpig
bZqCJF1OpXMXubHOCfJJFCE/YmOrZ1N8x8lD/YrrtkcWK9zZRvPGVIx+EvNI
oiByhzXeuP4KpdTEVw8GkxeLR5OmLeGJ7l4G/YnecH6DCclwWs94jOTrtM26
z2ZH/rG3SZynmlycYt4fmASzL2e5WQEsMnbRUjTDO/FmqKtyi+pNuBCCrz2H
vIgfZhQsIdT3P3SfV6JMgkZLIKnL49tJdOfZPUbQf8OxcwQj2jGncUWX2Xjy
WTPJUmbtvwETL+vuejedh2kG3dZ6/ddCYpE29YV90y66FEe9Fj2FiDzqasVc
5ij5diBeLSrvEnqDorEEL8FgUtYzw1wjV+BvUdFDIRuqBy+5qrCKn7ltyykN
W1Xu/wCyuFiDs3KqZSykWM9Vs05YFgiAwNioXscsxKllQJS3rxD/csg0q48Q
/QK0lnaexIEPtaud/UfTHgDTPtUxDRagOavO6RlMJLloaCnhyCFnaTpBmd2b
qEpqKKF/BiV97TeIvzhcdnGAgrt/F28C44tfYbGCF12Tv9bmMQi5qgWLPSaR
kInQCQ0KvhecmzOvQsAIGynpluL2Fn8sCroN03idUAWs2ZKfGXEk2GFKeyWK
+9ZoVgOmmjuKj5sPm7TKoKlIPmuF8Z9IwSQHtf0nEkwnNfP+DY/m7KAoa1/8
W0fJhfHyfYbj/6tPxTei16CtleSCRTdYS825ERetnIwCCL0P19vxMXm70Edx
PJ6fuzfI+u9INQLUxRiy8xQlgR06Kg/XC5OCQ5ALIF7HcBvERYfT9uU6Xiaf
fb9gFhRqOWiO6SEdZDg2ntGRg/D1keDnHPExM4j2mphBhV29yX+T3hvnsRxM
keRPfOVVR1X2mzsApf4k79nCzp/PORGGtjEaKTZsirQmYaLNyZWicPraI0J2
lfMmJtTPAUmkkg9rg0r6j50Q2FRUcA9zYAs9C8wPobeiKvJz+9xEAMGZzXyo
SBMDkb14sex/SJu06u9Ua7C7t5C+2QBn6bohFqAM1QUxlvDnOtll6GWveZww
9AI227TThal/z48zN04eLqHRL9LUCBpIhegqCJUHRMxbXQ0i5aSKCkH4D3Sj
zWemn0SddwLiDmiV3Dc40KqhP4+2OLmIcHP9AwaIIHSxhPpx/WSltDV6mofD
eTgRNCK6x+uPrQ9vhnVHUF5AV/sugn7W7+XBMH7J2jJ+4m5JDogIFoBD7oJJ
rMIf8IclHIfra5KxWD0Gd/p4I3pt6NzMsH6WaYAyVOlr1ZJpTTXyFn87rtOW
RvK9ZgaPgv1m4i1fkb0bmwNvdyHcXpmcCy3sFNr0PztkZgg+BhOALdcWFYK3
49mqxWeunKqMClszrzTUHIETJ+u/4ugMeDfybKbVkdqX0COUno+xK6qwqGMY
TfAWwgVSEKtDqfpD6tXVqr78QLKJ2dYovMAoLN94VZLvJXouH/AZM+jWVw2t
7qH+CDCvnAa07Ri9gIKUEulUpNGxTZKt4C/k8tKjFiKsyqu91XmhZhdfmj9Z
WeK08qZYDL5tXrLmaNiAR8W3mgmOHmrbl9lQc0gFajex4IvfDenya+X+ufGC
+YjYsTdDte5aUAvAYOK4n4j5GOuQba5RxTsLbyS47nHj+QBRQUp0acFUkswa
lx/dg22NEz7KhOpfsOqoMPPAvm5HMCVYK0GO7/lxHqwO8MNFxlZ+EU1Ax7Kt
ETjlPyI15Uo25oGM/njnL3HQ4YlnA1DLvEjQuDaa83vlcYH9kW1Ulls2gemG
z/ma3rotTmVk17fNLXSxDZ8EcYWF1v3dpAvA2Ksu7eHVzdJP6dSTqiqua9NJ
nn1twJFwqpk5yI7gjjQPfeoszDcM5KsKr1ywHB4qSsNwsKQqf4dQlFkGDiM1
xkLe3cJc0qXv9K/V+LIM4q4OyXT1tOASm5rJyZMG0l7c9SmzgSdLL0m9QEKd
cC8YgI9DvFtEJGxeIeZSr+/PU8ciOtUf7eRh/q9yvdjR2JdkrrAkgvSNIO/O
Gg0t2yyUOE5WvhpjY4pvebOrlfzBImrGaUTSCtb5fNDLnYGFw+0m5/J/455E
LcnX6MHjy8OjMPy2YlIbPh+CmeTp43/Z9LXuCovlvIjgqweBn0b/AnncwOcP
F5DvkJqof60f4zUNy+ZlAQ0g5gi+13n7KEotkeJOYfRb/jXyl1B0Hi/ZTQ/v
oVdB4twFS060BpBpthy66thF7yokWGXDViMaXRk2XkF1RYGuHYiov+R8im1V
76RuVPhNwCRIdZJIYkM//vRl97/fhi7rGPg1pOA1Z0gdvHVi3F/Foa84I+s5
EfnezeeqE+INjVpH8Ej0nFKcr95Odba67AgqJQReJ1Ryye+P2rKAfmdk+6wN
RJRZJ91aaux1h4D1j99IBpkSnu+MOP847+30k10PVPK56Rdt/tv2QL/x0YeJ
fkV1NVdL0M9gOw9vYSmBhwD86/JVfjM9wmtL47OQhz3r5QFXBZDrezPJGqRA
F7Ddcc+VJryoG+8KuQ3q8kfojf9KQbxvZz9A0v4gGvqqHNakhAF+h6uBa6yv
mXaRgZT5csrlbfIcHGYHMaRtUmnzNhEa9jTQjpAU2Y1A1R+ILcBzhJJAuiNO
kuIQIow9hlIeaw1d7sp7+WxGGPDg/AMp1WSjE069IgfERv0RkBbKklhEXmWv
epMX2PLWyV+Lqs0GKxhyT2tLwbH927oTtHIaKMYVacHGhEMbCJxQTVJfN+p/
Ab7l3P+9wrOhyiMUVwnafjLypgDV8pf6Cn7zTNOY7dw9FxfvSgFK5NV/SinL
Gd6dCTG/SNr91vKp7bmfoFYKPS6Y6tadn6IaylBWDs9rmJFHUe+71oTCcRys
j8F45CfsLtgJx9iPujroH6eyfszJQDD92L7wjgh2KumHwOZwQUKpIQfAg+/j
9mdHst9u9cbJe7I20tzwWwFcf5y9TdmvQdDZGQ0Cz2w5mMVgwmES6mQN5l9r
pCngHbTXpKbvdTozRj3U0YcgBbb1G42KPymea12DOT5P+zOECogo1MIYOwPi
FgGxiUMssXGAoqoZgz2r/19wXZYsM7HEFZZkMPo7iqc6KAVszrpBWzgVR1cY
XRwaX4wZRWIra1hlkGsj9xD3bcGgFH/VaZIrlNymfamh4NCbnesDFKcAPSLb
QWht6w/my4qM+I9eBvsoYMg2fADvyBIAFqw69xVmkMTGrcoG4cH3KNrEqcF6
BAMH69F3zO6LCAKpfBon2ndRudoGfkvrCHJM4W0KJD+DtXGSeGAY00mDF4LW
NR2Xjl8O1QDj75q/M2rO9ZDHHBTSN5qHYnnyA+MX7/o6LVw2Ur7dbtj1S8u0
fc3k0Q0Jlho7igmf77jadIOPdr3OAh4ipgVeoY4tHnKFVuq0SI8osNA4U+q6
Z2/QzbwYk4DPOIdCrwEJIMQGsETHJuGW4htgYvm4fsqzF4TM26fe1N11cLgd
tbEyydwOsizpFPuPr2l/xdwppIihskb5cyJ2tlfDgfWghs4MWl2PPmEq0ycb
+03JzTyOh+nZki/CEektL6G4H9oZzKetLKV+Ogw105kciHDe0GgSTqJLwSDo
GL55IbZVbA3vwalTQgt2/yUjDCrelXOwwy1EDZHkfNx3BpCY7MIhpg3xrbIN
mc8//0aUQEd8iIxx4ZcTVlDEQ+8kvzoP4g41HcHwz6GBSD52LXWE+5c25nMy
Y5yaheARcWMGsBjY2BYW8T+HcpGbUYVlf+ogQwl/y3l+MCovyaHP0MmeT9Mh
8cJ5FVFJHJaBaS2lWPcxhUwhskKuYtsnhtT9uK7aRTF0r5V9b+22rkeg203p
nnBQnHrzpU+GfAf/PmSKGg/UB1YNpjuNORft6ri8Pen5BFm8bO+TDRjVRZIn
m1qSuL7EEXL9HO6EKywZUeLoU4gweeVoxFZCPS/PT877Ms0rn+3HYrGLTTrk
F4Tau0icjlL1VqxVMHp/Rv8opB0OuVfenp6n0akX4OvXyudyzvbshpFLO9vq
QxwG4sBOAsNRXu+oZStoUUyxyKGgBkmG6Cyqcan+7v3Y29VQBulZByer3k33
3V1kT5Xfxynm3bbdcH/aGhv4xnZo0wYnQqL4URxH5X+cqO2OViutx1tKnuS4
St7StlTYlxDoLjTK+bcPFaE5fpJ7NT2tHPKsgrJalYCSMrVJu4ZODrHeGPet
C72rllsL54NWNzZysv30b1Vsrfe2cfXeXMWqVXNGyxoZMz0bynqvc5Ws30j5
kh2ISDWJ3rf3iUADEuvHAABAUYWezu2sDhui19IsZUaVJUIrP9Ogit+7fzP6
3XiJcyt042X3K6o3k//k8D4llVznxkywAvx/2fIGdLJm3WVfig3wEWLIrfOy
Y9XJ0sUVFgkTzDDg39ThW5wOSc5eZNlgbHHzQyPmZSkxZygRPvJ6K9LKh7PK
1iLx4DUnPkO40AkkVDy7NbTtOoUENUOqM+fUiytir8M26l2wtMQ3PazGRXIK
AMYrfkW3Oj33DDfcjE+GHWpoeXOS4Ii0QJBOgfk7fP1bWS6pCqw7+fU9Zwul
8ffYxiApRQZ0WC1fSVNH/Ghpm67SNolplaSo9ucPg9L5Hcwb+GL4v89JGWJd
jUVdsCPU41GY0UTfkJCwUcYKgzicDwqsg3wrutNAssnEDpF7lr5Sym2phyV3
j29iioi6OhRMCPZKPrD8vivUmpSprnvHdPwFsMuAEW+2IK4VWAxdjO61X12r
pbz0r4AaksEruemTPT7hLludIZrA2s7rM7jschr6FBqda3zVuIIzwNdN9BP4
26Gg6R5lFZsWuQr1gikbOjsnumMTNeMDfy02s9Bp9bnJi73QjC//vW9DRSBs
v2NDqKiuxfgiVAihHv5R+ht0bj5NMK7AvITV6K9SARHxRqH/GhgmYHLFHWzi
Mwad+6dNnvMdYWiT/hBT2FoWAZP6Je+zSurqVtorihkosnO3UTa/9UN/q+ih
xJ5WBumU18hNtXKtqQtn7WQn8uRlspbr5zNJIihvXIN0KqFQOr9fiE3rnUIJ
bCLVgw+7XKYWKp1H3yy9N2ytk/EsetZD5FcUAFtyTIx01gQDUf85AEGvGFYx
E10TMU89GA9hChM2AZvDQ0a+zM5h+2NOLp4WisI5P9JcqzSVbzPREyTRwuXd
o10MTNgyeOa2vYvW1l3diMSAdyauJ3/qLCItspBhAkbZutXE8wGnly6H2CMo
u71nsJ8eWQnM5qk/u3bStNrS/tYl4HkFA5Wj+tiH+kEJiOSJSFpvoYbfDxFt
8LLXaOCvFtQM5vScerFss3miitAoX1gB0AyQ/WAn2caeFSf4F3l+HXuffVik
qDAYFJar0fuaS/I31qRjG+fXc9uzVmm9k+IxQrHburnn1rxezU+eVif/yumT
qe0N+ks4EpfA/y8CZM6FfvGSr2N3wCNcwqw18v3Tnmi/ROr6CJvoF2PCio1T
nzDIkA1k3Y2nporfk1o4JC12gI/nHEyj03wn2hfAvcU+7W5xe/NI0TBH5a7O
jWLQ2nPB9e3FJRCrt0LBc/eZuwDkuBtWOvxAkOO/gRdrFvlf4uXGwlVoB8Aw
16dhfw/o2wFPTtSWrtUBOQAJdQs/nuesqU64quEXSwsHoKtbWhWDI4XFWiBa
2GoN7b4hD2cGhQj7vKono2G/xLXp7+YedzjGdw5jPJJuldhrcEqnj22HEq8l
aq31kayuF6xqAh98V2j/efay4QTzyn4DZkkOkVRLyG8WtKvvNANE17drWReF
o8ET7nEaupTAyZadNTz9Qg6S5xy4V7WXguHWxBso4Lfn4j0LP7Tg33EPSwbD
5FpJOo20N+msUH3adRkHPcIu8UpPT09nPbF+rWjWjPgkFY9Kft3nr5fUdFhn
OAv54S95H51qx1GJjmV1X/19bUh1yPb7ljiUN09yXtsE2fJ7XGwaJwjCxz0w
J3cCNooBt+MKNtbmZiH1Er0OfU3CXY4sgmckki6kPDLg0Eov7YJ4zbqQ4efW
frIeqrMPEjNcIijwALh/xrD3tzFcNsdTBDWO8KRzcv0r3E+sgE6IkofjyzyB
/+gyDO3tHX1lP3EFGYdR325K8w9U6uYRqECKaJDpFQof1wieWgf8VC/JPEHw
TrRpREJlNuAK+48WKcaFh8jFTAWsPjnG1+jM7oAxZPMGxLqynMSzfIP8Ulu2
DGcAJ8rYYpNYqGa8ETsuCJGUkJtTSS9fga43zIsOYBeWTKtZG/n327/W06u7
AXtc2QSYDWFiMLF4wo3wex18cv/uHyHTSaNKLFmiUQOD1fSgBSghGoypyiyd
OYAOD6NeUHk+IlD2lXb9+7eCTEZNNuwWHhIMJvRH1NRDOzjAbYM+I9btvoy+
LsSd6kCMWdRrQJkYqIuDNtUJ4jbZPU9jT/ajHKqMtdcUHyQPMfUU23UiYpT0
0b5E9bCb2bGal60mS0mZiIQpI3R8C4UrlcB+dHy3Rw6IIDGPl7ARNtfdaY1G
t8nU2bkJ0GTVY2ihblDUOwCVTtFz6Y+ctEE3UX2/tNqGNZWWmjQi1eisClZc
pfKKAyt7JS6YMcQUy22saQRQ+TtzCsIWw8Diw6bMsWDnuFWfgA4uoIfgryzc
MZEjxwKFgUsp95j3W5y5efUCwY3zZ3L0ZoeYBb4hzip8ltwQ9iToNWCgjxPl
CXu7A9TlMlhfgLFvDOkntkwNJs5B2u2E/XXD69I/vSsezdQKiUDZYS6gc4+u
XdYZGpyFcYWG8N2jvj+IYeJVg5CKAQ0PrF7kecMv6n4mLir22cYH1+Gw0lJv
MmLNTKH4GTVjzx4JN8lNd0O2ZLnHFM3t64fqVxKxrEG/8A3dHqDUdMASoCAA
TYnjvohOBMsaKXpC66eCtpGf0RGgp+/P6n2hvSrS1Ahrr32q35UH3G+eVOPf
RmoWt/5uVbiVCvx0JsOpd/8EuSQruY7yaox9p7Et8QCqi77lxV8Jm36mGPZt
zL4ak6ib1TtnZQ9BstOGgaYdd2agfHMawW3LJFiF+IxZE6q7wwriEeobAAI1
LzZ4csiI7SUr4G8eLJw8lqY84b2buBoXq9i+5bExeSCVY0bv+t7/IpLEFPad
SkfZTD4mjXExFPf+Ksil7d4ydc0q6Rmy8CtsyHzcYtieJAwGWkZ3zebEPEKL
/V1UAGzZG8YLHxyYEwg9yW6j1kj2yoAtIlQnp8ehfJ5sM6zqmJEgKTioZMOY
t0ZVkNJ1CVa1u/6dTM7Xa0SN4pEV6ZnOz8g6XAGOdenPXS9s40uYIxRq1k8m
ZX2zuAj4jSMkSQro0W12Nar/m7tSi6BiidYb6gIAxK9Y3fyjvTpcfoLHPiYP
GlViNSwKEdYzalezck7hGsolZL+/UqKLXcamaLd/ZTO1JPh4KqDv1PZ0J3b1
2W4pOmjqrJcsGcXzKsSIp9gzrS+nTuNJwsM7UQ0kHISPXhLjBRUrbDdb49Z4
jEfvgf3W0HR1J5OnKiH2Miw38iepe8BWSbXn/KkxK6xTJXTDRv0cZIMO+T2j
bI8LVSLLm6zH+teZadHmCpl8JTgjVA35KkhJg69vGgbuHQ7zNNgjBnIdVp3o
mENxPoAxW3bDDIUEJ3cTA07R2uHqlJZ6B9tgKHjiA41dOInN2sR89rqUol8g
w49Wp3MXIjNsNTM/6LsUBfzokK2VG5sK3PeeEbFRhIpr8bMDaLIPKhWlO80U
kFHcVGow9J/toIJ7pTPyNnJvN4A2Vp+dJ5HBzcXa+LXQV2T0i4doA/qlKw4a
zgTk5XuTY40lhObWRo+Tr2+nUpFYZx2QTAIR1+d0lilvJDHJcEXGp9VvcIwT
S8lqER/8WrR7tAW1rCTgD1n6SK/QYPYUr/w1CuAbxbyCNyCD+rcHcyCk7Lo2
YhEaRgVzIiVxzyDiobo8ACbpZbw2UBZx3YKLFY6Bqy6wgQKre+qLl/+EznBU
Fc3PDrCNHCsZKq89K6ZlqynoCMBfeYr5jk7VJzu4YiXFgrcx7sf8AW9TdrnK
Clx6wAoKP4k6pcCPbhwOn6OUnwgXnBDtMSCTu4mN99zbuG7SfIxAtixfkEX6
JSev41rK3AVGzF6pCmPvTvOokWu6t8mh5zNRBJhwedBxDFqwRPGgV6cSYd9R
fsNTJ0CXDKxJsWobRA0qH/cxWpPCqlkdqrqUe8oQYuFhH7UAXGKweBAy3TtX
5N00nj6H1/cmn4xYFabaLSu8KE+t+Q0SUSax8z7mVjIdZYTK6XAdehU5OjqL
pNwIV+IsWaLzQLvXN1tC7vNHFBIab3OtvNbutQcuDaZezZRZwUinePvewmnR
tnDynRFYDwohZQvL7+0RcKZpRztS9rdqv88J45GAwndVSmmViZJdkZsLF8nr
6z0XsZKzcewhJonxlnFncvXuMt1VPyt8NNk30oHFOCqaQb+yOLG+XNJLUTJc
4TJwunzS2DjJVkkeroLIrUEwLd34ReZsH3ZoX6NVpKMn38t9xqUZW8SI+4CI
sxnVzStDT4RaMPjmfdt/zJckuMBpOfPxWjUWCHqa7lpME+jBj4JumcpJjeFn
yALxX7SKx5lMWZDEjXxBKBVyoD3Tnq97ECf6y/AmQj3ZPvtK143v+b6+/uuJ
W3IrKP5FOWXbYye7wRgfilow8HWOf4H57F1CPKoc5qTAUmUhvk25x62V25iM
qYVodh+7CxlFf3iyKW+P6ggu+FbEL+mlbHGi1c/0PdwB+Xe56xvxWFRwroVA
nsqJ1+Ju3ez0cLYorfPgMPkXjjSfPloRaY80ubXfW8WUX5XK9fChgbf/uQsp
//HO5AxGInqC89euPXI3K13rFLFVUtn8aQZLKz65TtkNA/SImK2zd76k8h3y
sM30w5syWnLv27yKkwzU+UnyS2jMOMYVcQPE5LaUHRkud5sjvKrhY0ED/iPF
6sg/ZrrhGsVmt/Mr24kf0R6My4b0aWmQOaw80KWZXVpDnzCOBvZsYX7W8T3P
vU+evxrnUGHX1M9LTJtkZ8RRE3KUL1m0tLmg9zANmz0OzMuNDzW3ERLJVqLP
j6OyUM9lORsMBLXWXs2rQ1yhHeQzO6WUJDtkU+VrfvVMSGumkttEpM8y3nHk
1Wbcd67UjSnX28H8Y4ayMuv9QDeIAyLYa/VvlIKhy+PyZV/TgMpVCPXf/cT0
fZVA3HhDf1QFOZ5+QPTiv5hInXwxhVbu8QFp4V9Yfc7pPJjpOC0hWWqMxFgx
SzjJkIItYJZAARfQkQXLcZCNTlnBUt17lTWobbrFAnCNAz6WGDC8IiMGEozi
BHCvcdK73OEAvqdeieNmkQwjIWCzAenWkmN85hq6tEoFpYnPPD2hsxqZS9Y9
6bc2Nn+5CDN5ICQye8OXXN7pD5+mwzW/9wI9df4vd5NYwzer+LX4Ru71ilFD
TZsowGLdfamrTOcZXcibBxp9MRjUec3TtlTlHLR5VDP1yJUrv+tHMuCrVBHa
hKOZDdAdZQCw0ArcU7gP1HPQNDTKF+fQ3CStSIl9LrCuyP/WEMC8b/Unv1um
LeJ+G+94MqFeIpmyQqp9RbxNB5CSo83TVzsSGX7hu10OyNDHGLBO+LgvAVn9
h6pQDRUEDNxBRTg6IDk8ZJaXz6ghxsIBPePqmpzCXmaTH1yePoDaZamqMmH6
9Wq0e1UtmNpEbe6zrFcGBxxVQIcu9lvvzK02cEriTzCXWATAuYTq515T0CTZ
wZDRhgeVqHGjhHppmTpVv0ATmpda//+d1ktfxCMnp09n/YpD9HKmW1Dwvx1G
ddB3RpDvECY/V3401WSpkHNcyg/5uapgT4CePCK0uWTRerIxGbUL4GokBwLt
4V5d8Eb5wVSNh41qiiIYTJaarrFaSG0ADWIgVAeRaSf+075Yba4u/Z84QQKy
3pIFP9KYalhqe7U5vWfzOuCOMoRo2tud6omiQay/Mt4JojxwQgUNpHc5HSGw
9d+vcNfWnDL2lrxdG+qDtRB+uyWWYY6p9H+EacdI24qyVUvCVlkvu2+jUmEJ
CP1dtdAn/V6oOhG3lB0105UcwdDkMQVRvjNXVRYB05rEwcR4GUENGXFUX+FM
u1FmBvRDJ2GFUa2q2FbhT38ezYUsBvsNjwZQqZOV6EHhP4QS7LV1ZLrQg7hA
EeANJ+xE021gdn/2dOxJ7e7PqgEKu/t14eaj2pbdTvRHIGTtld3ydQT3goA+
6A1YOcN4uqZR6aJYEdWxuZdCE2IS2rH0aTIfTusK7kie8vYA9TMhA/5iPmuP
4T6Cg8hCrn8Hb1LQ1rPla9kJRQpH88r97Tcf0VBkW3wEGZCu6cJjMmAyJCeN
kJo9cs2bqXkJeMIY8WT7KVesw6kNMdwuJgH8pLdr1kugbG33xhdNhvy+Fg6J
R5g8snksn10dVEAJvFv16R3l2mavO+Fk6rpyZ4fNkAC9uyGyVvSvgUJ6C6Cx
G27zJuVNc1/bGZ8yUVnl2nMHVnuM8l0OgbuscM1Im/nG4ABRZluPJvS0Aest
VvZyLRkD1rxJYfNAX3U2PV2eOk1zMz5P77aCKlTbjvqP8qXH4TWDZgxM2OrI
qEHoYm+htncVSydEV9ry82CdXtixQZ4JewUX0l8QBWOA/UjBEJHVYD4RtyS1
+XorJ2ScDEVgefuE07P+tuLxj1gLJ6s5viaJdvm6iY4zWc/oRXwMH9uFhNZL
Gw8LoQkidl8T+eSbWl9QW2LmGUwriM94eCUubEd+KWVzyz4RxzUGg3F8zL3e
eOhdfeBb0w0MeLTkye1AyUc+wO3TYjkWIF73X8MUhs7Z3qeNe+bFL41rLZa4
lMMK7MCc+k2xIWTCSCetY/+8yRswBqV5BRgpK8Ka0bVULNWRwuZ2dNA/6LwJ
CdrjLevnRn5sOTkzWD8fB4vomiB7tTORA9ifW6o9cudxz8HjLzoz1vuHAQQg
6nNSodEPkcUfJOOqNfI1JcZdyR1GrLB559BeAH9nZXytRKi5giKDciQ3xbdM
6y6NgkhhxDSwmSu3lQnIHO6yi5d9avuj5TLV8+s5du4VR55Q9nrHpRFJi6WX
BWbGSnMpoX5tKDi6mBEo9kYrUNfsHkwoPE+9vpslFUE5thZebKhlP1HY6sTW
N4xvMsmOYfW1jtxcPJDxNTdfoYz75M0MK7MMXPthQI5NZuJPJNz8npXm71oA
AS1Of6U0v9qxlagWo1LPhPPRqlFOzvJAJX3mnWhC/8BvBlMEv3HbhReXS8pr
BofNjMnlBGPvwLC1/ojXyqHU4n4SXc4P1bcvKhtapVvUTIrHd9+NZaski6Bp
83jJDunt7A5BzZtI2rFRU65R2Jwl76axEV7UcwNAo9wbbIWyMR/TcSQWCPrM
US5SYL5BozOR0gYJ9fG8Hh1NfyH7xByTtRy0KtK/SV6QmBb23nAqUUvLwLEd
0hEn0L0qn+4tMiGMhltHr8vp6Na05pmH8bcNCcVMzRzUTr/EkK+EEWV7e2wX
jUxkBuSef51Ek4wZKT6ZSrcM/gQgql5eIk7j7erXXjKTNgGxz3WeYAXuJu7y
sTv4aLcfBMD4VYxo5SIpPWj6I8XWYxIlKU+Dhxb1NIQnvfJ3HiwTNo7ydkb1
cESF2o62/8av/XRbql1Y3+nYRxdR6NagYy25uXu1mp0kgr9ndN8PVT9nbXZ6
vkeA2WzAWyzdKptuNevfl4DzK8yK3vgy0QO1wrwJ3OwQtWbbAPZ/teBJQkss
sHfjqNMu77U5KpYNavyTT59zAg3GO+1VVtGIWuVwDobl0yb1ZBK1OluHt4Lf
DclrA5hIq7HDscTw/Oi+v5A5wKux/9KcA9JfyjPIrBVeYrCcqnMyTa/jl48v
igsUh7P+cqciVv4cJZL3m+4eyGunzzH+raPTX5+sOmX54rhHPo98ahsx7T9P
1KanmLxyxqx/pkAkHsLPKm6EXYbpbRMZgr2jKFe9Jl7jA20qAf80yqWh9Gn2
YGL6rtrrB4W16ea3cxYTKldWoyxTJvWSTtKW/S5KnglGH10OatBL/Tmx43WA
H72DRfg1R07jT9ab75qo7XHtcS6ykmbdaNnKC6U6ciMlTTET3B4yruQAYlhw
OUWVTHQJGGMB8noJiFMRyhg9WzldW8U8KkC99do8Gt3tmuR3cYbl6kNN1XxQ
t27QawBW7pDmQOGQq18hNjpCxqQ3l2KWcXK3vQl4fgkz+1kdP9MErlRKfLt+
t27/f5LBRZ1sdhaB0ZZLrIidUCaInoCSF2Sc/NI05EGkCqFY8dNLIVuaFVG/
Z21MGuuGtTEPwANhDSAi5QyimZeoUrobiPGdrA31bgIToPcKAhcIcwFIWa1x
YD7oWghhZIpggvuR+vXqq9IdmSXnhRNJuPCuC/qWiYONfZckoFUVHqqg7+e6
JcIA2DGlZSxckqAJhEE4fl3g/YmoPh0G26FwPSu85ggWuXb41uyZ26enxc5Q
PD1Wz/oaDMCHB4b6RmP0LsV+/W/njYMBM6RNBWT5uh8du7EOEz6JM9Ny3pV5
IPvHkZefnV3gvGRP56zlQU3z6OjQ7aTSE0PDtLtQhZg7BoUPW0EyYTI9/CmV
5gvY+Ms3DnO4U/YjNTYdC+VGwfhLBVEL+7gCJcqOpGeregTl8o32WeAawf+V
RT78nu1QXOgp4x5rfcAMqEcS8jSWV+HufE6AjcHbMmhAh2PszJSOQTA1TViL
kfhikkK4LCWUp1kZnLkIDuxPk/ZQcsnI9b7MNX2WVlNl6ZVGsrHNcVaUrVVm
KTuHCFVPMwinh55528w0g7aWdYHZsn9F5dCVpRk9CTEn38pt1CKlOX6GXxUZ
N73JjmIRP5o3urL3Oia45qoAAL/kB7dU4h5wpUK9gpYoi2TVB8Eh2xuOlfVn
FzfuEasbHAhaNtbO0JEVAqeI0t+JG95Wi34NyQP+mWaVJqm3edzYtStUrNJR
mwmt4pL2au/nmwvYp5K2gKB9jYsZL5SFf24Xl6jDjlxNdCSsqunANtJ60P8S
JbonsUuv4JDibkaWOonrmZwhATAhH0Yi4cFeRn3BNpe3pjw1+cFB23xGHtcM
Mp+uT43Qq9xmqu6EJ/zDbOkATYlyffBe7nNHK3esAj3oFyy8zZAQ7yvMFCo8
GKui/TFSvs3Maa5Sl9phd9fWJaksw0maJpeZclG8EL99bAyAvhHg02U/TB6s
M3t2J3XNq87T0j8EEYoy8hHRm8l/BUnC6vU5CExTdt0S7RC81Bw8hZiktJj3
2V2RrP0i6BsSw1sFTk5IV+7YL9Uqxw12mkuI15KxJF6K2jXKucki2AvTQY9f
h3abKz7XMeoOtM5mlSWeAz21B/1hoVxnqK8VZ8fGGElRWb3QmHBr/ET26vCp
TUNY3WtHCll/U0fshrRK2YngIAUH+KqbXiD/2LbCtoCNzMtyUrWsOGt17Jkb
f527tg0CZLE5NXfj/C54vwzOw4TpDuo5M4fRaCaUtrPN3VWVw9L0pUPerEHp
26Ph8nDm5SeH37BQBt3pBljSqgXk1RZMluM7SgYaFdlOY+rzCVXaUHojxo3B
AJDMvIAdVgwaT/+oEO3oW+CfeW5Zzjn9+z0MOM5A5QJSgqk9cBE0VtyhkiHM
R3cLnKtwIy5izCKb4s7ZPsxqR/9FKHuQgef5AKvNuc6/ZF/laZPNCG7UQvIN
YQ6vZCQpSui2gjWMKAlFTU6Oi0oZ4RlzyEbUQ6O0fCArVnMF7l/KXq63/R32
vTvoR5de1775Ntw6OkS8rEidHG1c09Y/04ukbbsZV7+fAMIHqNCachpjxzmc
CDbkPbfu2rwCRR8sCYnVwlA2j/G9tWtVRkMP8FKgU7kb9aeK2GwnVvj41/NW
OCFV1G6Pk5xPORoPkg6dOG0KES3iO8AbGs5HkSnadJ3DzYAGkJXxGV8/HcB3
QJdHGvfrlk3cOSgOIG4lk5tafq1wvFiAkjRfnkzf741IBX1iIKdVpT75bVml
RXesKlQUbeqIYnrAAARMGOjoaxR3lVcyae3ore/6pYIpYyCXcNMQAyBRBo90
xX38/es2xgurNnXbleoifOrdLWCAaLdkzq41rsIaMFmt6CeJW3buqTg3a3zN
orOtSbeYhvvBGF4s2VUDwIfb5dCLXbewAf/x+guSZy+3B0vh5KDFPQCkjSDN
Nxg5QlEa6asy3O1+CzgQ1Psv8VsvyRXNn4BsWAOWAX0k7+2g93I0fNDI0QZ9
X/+U2VlBW5LZt+DL6HrtTNSAh864TPry3rpexFbOcdaTxD7Fz+BVy53swGqF
LOr4DJYevTIjzI+wYB+IMh1lb5DC5EqaaYYjIb9uAinGQeWVKvwWf+Jw0ncv
ju/MaV/PlxdqgYsuD6ym/x731rvMCRlyMtQitzifs1dpOI6wMpXGfl/ipMJd
zTREMwsAtGJPzVphVJ44NB30l6EMzxEkZriVIGOmv2vww2jDbRnVEWTCuwMy
fCxxbzL1xAoGwVUMcDB9mOEsWNK1cy2oAl4/WFPY/4FrkxThQdKomNOeqRdV
4XTVgqEdIrCSOfs8b9qxwFyZbEl87UPriViaMUOtnxEt2uu/k6E+dIfOOquW
uogIjwxoNW5GwEMg3otD3Pl+rmG+ahp2I7+GACm0FypkfFzCn5AOYseN6QQT
nHk2yUgU7gn5jUg46D6DMyRgEeKHEmtW6e9QWLsYd/PcW2JA61oB4mh662YN
X08jo4pLKnbuvE3BDN8/KuAX1MymreH+KRxFps9EzUJDgtV8hyY1Mm5ZyXau
mDvL6asLNluQn0mzQ6c/MAbqT4U5XW9rTmRRTB/6Go03uvXTUNv4hCw1yedu
tGRoINxQ2dcP7t4qwu/5/D2c8YXl2MBhizIMiHB8+SwQqkkhPSbT5JPs21nw
oVN4Mxt+ukMqzDnRX4DxDsI/Fw4lXJXf/pMbkXgQzCwQ6/tEqdaKi6hpnzp0
hs3M46Zw7ve/kc4tSKGxZpIJlJdlqu0frE6YhvKR0E+Fkzi6VV2dhy9qO7zP
X+B+fjvaCTeJCUMR/gMgip2isCZN3e4WH+tuieCUz1f3AP5dmWNvKbM9o4JH
b2Sn/594r3WHEMYkeQkGldHAr0Yk6xncg5RYcYzhhwxAdBwr3IbvTNkfqKVs
B1uVF+Q4cNpxmtlj+PRrhRML1h/dGQrLjKTv48TsqKDMPfqGjamphcI2Md/s
G1MhSCqiZbDXUaaSN37HhL9VF1TB1shibFsuw7wM6WymGeqbrLgWaZL+mYGA
cQj6HNpxldvmU6Z5yU1L2c+vD1cZzoU0g9TAUFC5w3Adow0htHt/QwOlngH6
oYLLv1G3sfL6fVBNpDqKbl35nbF66+cF3uArwnuyY0H05Bkrd4PsPtOy5Ktm
S0ty0tmHLGmeruuai5bsYnq6B4JdnjToMBlIet+XT+b7h9b/RDr28ribarvu
ohHOJjprDgmuNixYkIs04Gfs2+B8guugtfbRbezUaKvSOZW+PpJSy7P8sPN8
KoCMu3BsTeGcYKWB92KZci+YFn6bAPCzFgvQ34+Vx8mZhjfGZp8x9B6mgrk4
HX5bAKGM+UvYvhs+8cOg2wa0WvSKtxhDZOhYdcHKwl8RpHeBObUFDMPxX3In
AnkB6KqzW5ifd1lspr8CJ5I6IwgOwnnfwM6aMdTZLOLhBMdinSj0vNsxWrEu
ihNAkli4edVzL920a6kEgEDjAEQVwjlFrtmgLZS20ZSB/mDoUrEhZBYNMTC/
iL4NqE6+6Bt1nmiolU+BmMiccMOp+mMQz6pLqCzoRx595oA6aMr+XdI55yj0
vxB1b5VZpVQDr+J6bWNCt5IXBTI2pZKOXZw9n/a0A8nQ8QBs1FUn2KrX/lMI
Ic76/nbtrlXas2gXwlXshYgEvhdVDyVCZ+73OGDixnM/7ptBDJjgoOqmeYFU
UcIU1vPqFs5I+SiJ/He9REKUCz3+6aZPqCz9gpmLbAeTo5DR91VtX00Nuk+a
yuZmV0zv5opQpF85EAJIj4zi5fc0eb1PS7chMhzGdrIa/RjJTryHlOwYFB57
ww23bQxhdbGvAqTlG8tdIEJ7oxHWsAEp8qFZpeOuMgXJa6loamxnYDtLdsSY
xPaPzLA1pdlgNx8bRdNzpFXXkofOG3J6Z4wRtU/zsrQXO9E6SzlvLcYjnOlp
A9sueSUS+zUv3sleWXLo4YQCcI39ReV2vk3JKH59df1qmoH0yWyYeiavj7xD
m+Hdi2afbpttpuFC4rFBCQNoVQHX6ddf50paBNr296mM4QEi3Fw5Jtjsd9Hs
vgSDMhCoUIMXTaqGAFZqMH7IGpQsjP/xcxZZbqwijOsH8PXc73Mq1OP7lqfZ
r1PCDYZSXXsfEDnytG12WcD7JkmLcZPgikcpZJfNtUwkN9ROU7kp+xVBlBRZ
3hSY1BAeP/IXeZgr5omh6gJz2F2ZCfDFLr0X//69m+9+IG1uGNnudhW/LFAI
JedYZv2f3+gzYcet5K4iQd9/SNRvbayLfpmNOQOHkb2mxg2HlirpmCkxAWxZ
aZrhL9tMsGAawy0Sz/MOtgIpwS+sT6frSKrYCyCopZ/SbfUeh8+4Y/5NmXAf
+hrZ/Ah95pEOZjictUebB+TdVi7yciFDCBWB/flawzWjnD+OLC3u4inNmKhG
itcWrUEq/dPc1uLmWHz7eMf2rtTCNFTeFlvR2nnlpt3usIrl13jky5qpWzF0
nB4jp9UzrNl7k2bmrEdSX6l/oOMZ5uBRD3GucE8lwWAdzYJjZIuYnSt7rwmD
0G3Pdeqa5yGl2pVtZlchSJvdeJdhBZogi857z7ppiPlqA2+kGdfQ0z4p/AR1
Hp5NZpXhvyjAmg3gD9fmQ22SDBIokNf5UCKeOeZU6iDOG+JWba+4n5yI8R9p
61JnyCXdgpdzVGhWn9VslHIE6mCrS9KKhmH8V6ClI7rn/guZLw7ZTH01TM4W
b4AtNFZ7PLITjuVA77DP9gTj6eB0+M5ZhfW8u0TuSaR8wTh0VyFQpkaTrHQC
3hptHeygygcPI6xWVC8bmgL0/8Z5gxOMYBXMuqHbQbsBaiuh8q/h/hN3prkm
v3Vcx3lqCB/8Czhrso7RtDyQgF4WlmsSrXY58682OfFdDQpLiXAhf9DKAjo+
zunYwWo8QByZMnRxYZKHIBuqKWXxkHr47rm824J4DI/DnmvpJbuQEi0usi6/
OGPR38IuQTIHUaF6S2iIAUoiEBBKxZBz8bLTAqXAMcEE3g4noT/LSAUG8LZ+
2g9m3agbJY7bI3mx9lPutXz327LiERU9W1SjASwzRlhQBSi5ahaFUGOQ3Y4V
Q/ojDCObNgn0mKwW4bz6LgFDINsz5gMyD/vbSDVk1c2eK1qRNpYge8VLU1m7
wcjIkx4LZrHn17WTUAeeV2NXTSX4rwRTdtAL95XUeGDoR3XsrthAqiabsBCE
WuVm0C6cKD7WnT0RsdU1QMHT7JH5YbTPv11ItjapIAyq9EqMv74hsuCzF8b7
K+wHAqD5+paf1HJu74vD0TvSrFZI6x8IJKf7ArXkxJ+VKYiUrVF0nrMfSToS
NVBcB071+vm7071NAtbk2/OSsDKIGqSQ4LDGy95zhkxBDDYnx0JeTWXuBEJP
IZGEWRiolE56Xm5dKYA29GDjqDIKebAmohhrqf6Uxi0zFFcdHmhoiNurDrNb
90CcICzU67wbwHY03g6ztTfQRyYZS/+WVEMz72+Plle15TRgm4SMFQ3id/Uv
JAK5VYA5SkBmoMBxLp4Mk+2q/Jeii5AIoHtWbViG1xdIN8RvrfALruw/KxBr
kEzvVoNvpLaetVZIM18bu91e+8oF9fONpGWATQOvvlPpIjxZjNXx9dgF/CyI
R7z+rDc9LymHT/hhJvfEkgnMEw6rfNNgO1UhNp2Y1MSMwCnF6sz7cHmFoUfQ
jiPU74HNJa2q4tfjI5g2ZIH2ni9ooE4p3Sz0Ucj80uRVbPxp5SwlAkfwQuZ4
HiDJmL/0r1kYufUBObMsRm1HU7j6wfu1u6U4PvBEadaLQ7ZuDk/7oKObl0YW
FeIQbF/Bl5N9b7IdhWWcRxLVA683ImrqZ97dfDGsiOQRZ60Vg9FcLVm10tml
20wvF1EjtcaA5jWX3G61h+t8izIsRU2hUIkUhsssWBaKYJUBbB1JL7YoWD9C
Cwvd2yE3i2iw7T4818lLwxAbCLqJVJVOMUWswC4FKtmi2v+TCMwRgL4k2rzl
XqAPUFfgiZbfnphqrUeKDbvWlGSgeShUMcs9Gtl7KUSjCu6wdG+XSR8b1wrM
M7G2yQgvfa0Un4c3qnBJIh3wwICJ/RhnB4mMcyAD30947j6kmQBKR3MWHylR
uROk6iOueHH4mgLhKcO0qWY/fg1XYn5x7zONGxusjceyC8VQl0EHp3qW6WVM
W7hqfQLD8JuwefBBFaMTugQI/WVFhpX1247MhUFeJXSyYoT74oEPl+EmZ6xQ
RSg7qrXEc4s76d1vC01E8ZI7kO2C0w1p+PyQsIYkDT41YUdVFxU2dnujMYuZ
LVQneeFYksGtH63/NX1dmrymlFZ+29C3jfHHaluJ0GVmMX1wLSEfYiqYi5z3
CVDIkXlVDR+AmHeT6cM+DgmLWYwMUuib/I3TDcmV1acbd4sucN10DVvnmD/E
4Nulq3mloqg2+/kzBxYk7XNEfIFB59gVn9nudjgNHCUHNZmInHarxg1xWkFd
21YBmuV7GU8c5AAGPUL+Nps+SbOG9s1kUISORAA+8HGpg2YvYXQ66SAQpKJr
fb5Mifd4HdjcXylcPL/icGEyCtHmMHqJ5tgYNkzk+f0AGs2VO4W5+bVm3oMr
WA4kvjoVOUfaIJW0x0zV2qE6CwIBWHdYRSgsAaYZTnhimsm6nZ1L5lGCD00J
zggfDQeBMFZHhPOIxNBE86MkQal+lv9M5FJX4tMKUmBt1rYd7HrTejW8LlUw
Hmv7UomUnnhaUEAyF3p7YozX1fL0WyecD6EMBsNDMtnVBk43ppb4etpTMV9y
h02wRly1whJUWoVYjLAM2gaVebfFwB+b/0H/oN9dXqzPJZ1RKrbxuIN3psUx
oq9pn1I46CTJTmcFBeqTjbs576f4bkNii+Gvy7/Ag8gG+W8dTrcGNjuHytit
CNWrFSySVN4Pr3f42Ib9l1bgD3l2NBypqcjL20CwfaJM8DDl/eGQBBSPoxn4
o0/JRbYd8h0BSeWQ7x4v/Db/T8ThnUFxaJQUhIvUVxZ3cZyLzXnxtC1uPFpP
U1dGuY8088v716XaAM1Il+DoOg6BBVqMmEn3H8/Z5yZ4YFamAZn1mbcdqNCc
cLU2EMa+eXCfwMe1t+3DEKxXJANCFrM3y9cRf+64JBUYvgRjDyvcr1TjohLg
8HEYSkvKMa5UxO6OCFtOO++CGEe/bANxXWTkXktt7T/JXZJcpAic+TcyTzFr
lZ3aYdCGZP7PIsWarr/N8aeeG5sCpFTE61yZTbvfVaPxyWy8Yk3zupbOYU8S
TUxEBrIhKGtCzENmZgw+/WR3cXNdOrmZP9GHNnszuhJE+e3/uQGNjscuvnCu
ct0UzTMWy48uStHoKPfz9AjTewHzuo+l8v17YDvf7n/EcjXd4Cskc/cZm10b
9LBLyPL+Jb5Bwo7DFN2QouWASFJ04FOEKHh9nSVAYnt3g68LN1cW2VYLo5PE
tb06Io1+jS90YNMXmexTa7Z55SNeL5q3582RBbilRkJfa/DPDBsqQU8h3pws
TFet8UwEpQJ5by7OpNBk1uq33cheoH3/35tnJsSnDxHf3nANtM4Gc+3td0Hb
VUzhmeLLFMzhyr6BUFLQkHo9rMU2toM/lgCiCTLfnsxsZoqO5HkBHpOiGfJv
EYtUT8qEDRwJ3CbVxL7tzFiArIWjoJKCiqvtCEt83gchnZmWftbRCtXoF2+v
r0wLsV1EBOEUkNtmr7264IIyxypcVftGgUiXPXDPhI1+PzjGkNGbuGJhPYAK
fG9gDn+ckQNxVWPX9AU8dIugXjcCJYA871keEtiomDkWItVwbf5kNC+Bn5wR
aLSOJYhZNlJrQYsKAxMi+fPVc76HhTj7mqChUqiy6xAeZuckgzSWZnOvHqyr
DEV/txXl9XennDUua0Dpm2AaYVa438IBjJhLqSeimYDFkgCDBnPI23+OKXh2
iy2zvpV1lq9Qw2/wZNHLJNcrUr8d2yInpf+ONCDERdwaCUpUlFDqPkmTHr4g
5YRPSn0UG+OTaLIlMUTGSOWq87wgRe/CkJN5DOTFvLUnpfy+IUJaipLAFjwo
efjyVOeou/Upkf+13OGFKA44ZcnHoeJvmVA9u230BRJPXRRexl/RzwLjPPL0
u6idBdSQBmRn7YjZWZRuj9SUs3fnqJTvuBmrBDQx4JnZV3iVSKyGVX8gSd4W
K2qjpLgeJzh4u6pMw83fs57YBDqQhgB6fE/xvhffMKCq8JFDVAvIL4oQ8VpY
VROTt8t0ORaQ2sA3unY717RQ1kqMMznZKcTR/gTBhFG3vTuMsO99Cj/MWJM3
RJlGyJGclXi33t7IYwUIGA8aR7gD1aH2sQS671v/zLAvzqGlZdmuePeuP9Ec
YvO0c/i/LQSBSNCAHdtu7YMfdVbtjtsY9tr7QWUVMoMQbQ0/pX2RDcaXmnEU
EiCXU8T9zyBL8/D04aBcGfjxVubz5QE1lgKVJuYLxLUoS0b7F8KibdG/zC0S
YHxu7DWcTPMrNboGMP3SD3kzVUjQIwXIrrYoAGfSPbn6ElWXKnYnvnH7gWpf
5T8MXV0o37BQg4H4aM+XRUrqBqX8MhhTTfpy0Xl7VuB3tleDxB+nkeDC+XKa
zqTeHt2DwOtZ1/8GN3r+BmFEYID0DdqNbGOjIB5MGieOP3e1EwvsuAe8yFs3
5V3wGJeXkafYqg/wHUBgE0PS4zPs1sNzG8mSwbpVbSuGqA1kA01SmN+sOfo8
oge4pl99m6JZxGR8V/vkFlzmb03xzB5+4tvfmlYvtmI/ji+AAHytH/pPgMb9
corI9GTg7ufk3HgEWi6QoQ33s0moqpuiV87jiKvLGNb5tZLwaZ+ewvtAE+Be
TCVUpCdbS74Y/fWzFlGo2N+cWjiw2561asME5sLQEJB3Atm4qGqAAx+/izw4
2a3hMMyIbHlu3cj2P5YJz9pHBXWxrayQam5H1JtyYEjAgwOufb69o52Ocyvf
5pE5XRSQNvvfKl1wQ+qQFkI249v2g5YO9Kao6ePwtzkgG8G5k4IAX806wyYL
3O1JVdi0GtMUJP3KxYrFA29yBKxc3Y5nrScvNFmU8HZ2mWPhYQx+Zjtywa+R
4PD4Hnkzc91oA8VfebJX9RIOF4n9CoeXfZqHkP2qb3IvgS2HfbkoSnk+Gg0V
1p0eZnMHMmwoyifPzhzLeXIHT0L85HJGrXVbhDil3juFe9pdQZ2w4e+07xVT
VUKvI2VmqvorXSeFCXFtj/Gp9YUPAQWk3Fds0fbXhUvzMc0plHKoCnAKQwAx
pUJOIT7qOAXHiqHWwBoRtGiKtV/KXuVbKy8YDOpDdJBJOl6Gm/1XEgiE3btT
SAGAYb5yWy1MqsuoNuOSF84xQv1FZcoM8ZbLyHFB878PPPujGA760cdhvbon
JURkVaJoDJV3toIS9Zs2joVoMxAozDW6PFufLzsvf1LRENLYNRG44PZ59bd+
+SIT85UbhUSfDS8SKlcWxPzThSeTCJBDXiRkcVNs+uO3bAujwvr71y7o/DSv
coixiV4Fsp++2YK9B3Bi7dX00YxMV91xTDT75W5JcVGO1Lu4iweBerYnFf0+
ySbGolF7uun/b71xdXjdGyjvAUyUoIT7vD52U3lcuJeRqeBImuUVBAcIJF1n
DAgFwb4W0vUotab7J1khQDcSigJaXkfZUYOfMOkYxhIcSq6G96hAw8ZRGNqf
VXKTkwX83ljV8JNtjzdgTrN/+NbmdoS4w1sl6k2gz/iLD/TdGeb3rl+R7iEZ
1NOI6gWQ5aplp9HdBDQOgmvQ63ygaJfByXK6vWIz1sTGymNQLX2TB2rmkjVB
Lm0TWJX7RDyes7qpRInvwW1fouNxzsXkXLO2KFz0YuqcSXtAhStFHrXRIMNJ
TbNZqEzWZcoQXHil//ffXZAZXbQ65V15kOrR++yTjRzTgONm5ixcEN1o3gN6
FDXmdiUUgj069Kv3yfVroWaD6uS7TxWjJ1L/tbG+zedLLi1KV5bRfWGNewH9
Rh7LMN8e83eiFcWEIhOur17onFEJwZYGFLeqQkz2cA0Nn+1k7U16ww5zUrfx
zvHmE1RGIEUcZ2I8IwJKCMq/gxy+pfa+PISbrwxVnppATAkS8Ru+HsnpqSDI
Dw1F37HAnUSZw5+mh5ygS0XZN7dv39XfaZiIESwC+E4M2/8kSSbNE/ACDp+W
kyVU+JxyIo2q3IayS42PZgiM55E1jBtGm2k0aU/+k0uBPgJUlbAcjOR0zmrN
8RcQzbzYzHXsVAIyYi+vb167k6DTMlQrAquBuNtQjnOxe3sk1mYxSzu8gPmo
L58wvLD570vn67WRa8N//7niHUrmqNS8+9326sXhUbCYCe4vDuiFSXQBP+lJ
HLpHLNyYnmFzPBl9p2HwyZjI35YvUxJ9OAl/TeSzc23ZQq7eQ+7wbhHkuoYD
QXLGfBjYJv8IufDyKkWuIZBHm0hvHMQmfsg8Dm0K36JrN/FBKrv7ojpN9fq1
oGziospXUpx0UQ0nG1+PpIj+ZYt1swvgysr+sCJWlJMVd5WyPuSv7VWggOyK
3rnAlQW0LXlzo0Xm0U33ml/D+/y3ItnZuRqkHskozmYvXzMwCKCPryzXsEYa
5qcKyyXXKTy7DDhC7mnsTMWEXLLpxnHN9bfVl8wfsuULgSN9Xx+zFC3xJpeS
oB+UrYaAGQs2L01dmKwpeaF7swt2z7lNUzwf/uvUD/hhwBDYTg17NXibbjLW
ybC5f1+0KB3ZGUugbuD/DJ9uXb2oNgIfrfuRMmI8z3HE9415wKHtHr3orDuw
K2kvsrL5ODJXQbcc7C32h/gH/ljmhVuQ+4nDGgcdGY+bVeePAg+5Q4naxZT1
HcJ5cf2q1Scz6QzRbRqjFk7JWUu+h0VbSm50+8CN5wrCoWw+wHPEGt+CiM9k
AP4vVzrq2Ff/h34deFbkLEkPSIiIrhShxXFzMc7H/GTRTnQ66S7WCWpOwv/g
2yrimvhMo44F53dFykKqKNfRO6bK30gvXnVjx6DClrDcs1HmP2trC4hRMKfC
UpOVvQwwx1sxwD1HleWwm8XYogYzqiBdJZzzwUKg6Hkxb5y+K2HIUWMBoOfg
Z6gvkpQLV/puKIkzdiEJP0iBev7mjbTZch66rXpZ/DsNA1Gk9iX0KfWb7lvp
e0B85cx+E0M77ryYD0i80aA23OD765lqTIJImNVkztJ+dbPH3ztDU6rsRk/N
duEMrMdbM/cLhohBGkqz8pB7d4WIVj6vpukXyQfwaVwsudhJbn0M5x8GBqJK
DJJs/cMGoD+B6ogVKKQFvtBgLBbU3uCZDaJiomJU+l3WZ9loXzBC2sNo1wmI
Zc6mhdosF4b+bM58GWCOGwFoIquEse5EDfv8B34CwCPw/MqOPQUJTR/oB2/c
INXcyjiE/NzS9z0hk7JV1xioXhilLFLNzYurj+0U5NixJE+tsegdpI/+OQ1h
5TI+nXecWqdjbzfRPwa55NAaKwe2pCOI3TTYAAabsnDppSkmUlL4VvqG7xaq
UTtKgQK5d8ohCzwkDk7s1fDHFD50tjtI6FCqGxfp9pkfCa2RjuHa3qtX/etF
ZougHiuIDg41QhOuPWiDwmosbVKDeb+TKM4xiijPDaf6AgnXiBHFUh925FAj
JP+nmRTeHvog692cx+IlxmYZw/AJnZKeLiWgGfm0KsXqqL62j8nVJIVx3bfl
pq4heBsyttWo+n6W1miY0zHmYaNoPtB08RJ1BA7BjPgPNP0InR6GYGyMsGB5
wnjksPx3u9EZdmAGfTlkKO/X7FSe1XS64gs5vNvxF8dui3q1zwuOdSDMZTUV
g4tx81MdZE2S76cP6MhVM41VLRFITSTgkhsSffsbyNFq0/Y7/6o2u6liunX5
HegZeXiDC7TnIX87hXbvD9WzorO+kU3oyE8fwBNGe9ANR/bx6YR5O/8eN6b2
xoc5+zrLgdhREnE4Ra05WK9x6yXPG8JCY3lDdDIssY/JDRYaJxSIdlYhL2Ir
YiYYJntu9eGkNRJgSP3BitaTWfWhsE0ktWbVJPRl6dVWTszVriKtSv4E/aaz
ptoDkwaRg2OVbQonb+ZlSclpRdue+O+vjC0WPBbNsbkUIRwNYyoEHEdwvIN1
+8ELdgBRYZf/g+SWbpTgIMlqEGSSdLV+bhVJ7QMOIF0sQBZ74luLZ74IVKwu
mvk3Z/JQwxQv74Gex31pWwBI0cBeEcS6GDHgsB9STB4M6QUF+j3DCtSS8l71
uhR9hLPdh7Ms63tu1WFuDsWwwQyHnNSDDntJVRTNQu51X6CS2Y6Kkvfq/udu
Zc3qNrvMqAFVRgFesLcDOUxxCDshixFm7TihHQW7CnEc7FPA4ggQCrdWznD8
ISaxZqIDdf4BH82xZ4nqcRi5niDTMtxZ/uENHBof7SgYKqvReijef2EnrCRj
iQII6No7M7d8ynxKcYpFGlzeR3cl4JsSUaam7MspwBRxTYB3SlKe/EqmkhMa
KVQ3QCbrMMY/9j4FA3FLVCtYhggpgjWcpMvZ2tj/N6F1syPDn0w19MoOAY6k
Tlc3KU4sS85rjuHgQur6Hs/2yTd/jsR6NfmFX9H776MjC3UdLstU/3s/4bop
nP0O2esJ6OXWqGECgB44cWg8Wh6YYCiuPi2vDG5z51wKHwA5euzdPGlmn0eL
tlRmee7NxEGGwhM3VaVX1jrLQglfbWJXwSipVRHeI/81brkjiF8Bjy6Iu65W
sYS7Z/ZZH53G5WL5H46jpigPDqMPZ5wR2I6tgGGHauCpVVfLGfHRXYw49QKX
QCAzbWu8kIWUu15KV276At5qIyC0iA+DTmW1oc2uM2h8vP3phoJcNXRPrE92
cVY9tQW4EjffUwx5rscN/q/51lINYP057y/xBAFxqbjvMxa6Rv5QwHw3KeRD
kZaxdHtXHRTznnOFI+OVuyWWCOWTdhmBvOo0UQtvyzhNEpItMo1BCjGRtCfQ
9FKl9Koiqi5om5OoxGjFVg/au1XnesSk3v9EtjqLCmD6MguDhfO6Aq50gxFR
oQ+xYbw85G6+NG70knnZwe9VJ2yNCd8bHD911vO9tVOdst9ipMjcMj542SAn
ShKyGUXTaDO5KkMVMg8zRubRDXZ5YaJO0zSpoUyFYTXsVDMuQlESu1U1LxEn
Fo53iNfCyCWFJPtSMGn61VGANO5lmBPIDUDhMNGVLSj4XAZ6ALumot83rXDN
NYkir7tt3rUZRRbCEV2cKMvRgjtGJm5G5ITSup8gF3NPgn2i9Cgxv9GzCnBw
jG+OY5R9Q70dlU11xLCkrwT8XkSjD8x54k/raeQ5ygRmQ6FxZiM5ENNfY6II
5owvbG8gLlk0Iv7Cz0jvh5WXVNUjdhp3iSdLqp9A1UtCPIoRO69sXTDo0LWL
Q5FCV2xwpmh/g7LpnkIvQzY9enmbB0ZZkpH/WWdSnziCkvtoDHPIFJa6Oroi
rg0hJ00FoMr6GS/sMkLa+lMcpRvABIlmwudJ3Iz4zbWTmp9lgOIsHvdxQudk
jym8fVMrRxm8sW5Ex9j1oMTVYcKzxDnNxzh83vGEDIhWlBeBI5c9+diSNAeG
VcxWPD3XaRIo6ycNEnjnYvNhxaYfx8VGudXfD4qjoJn9uAMg+XUM4e1ClatY
o657n3GpMK8U9mmnDTzo+IS2pDoxOXR7q0JK0DgA4iakkr/70+oabg+IS/5l
sbjG+2WqRBia30Y9Xw3zyF4TX6/ArcNm14LI/MTgX9/uDOPCHAdelC0Phl8A
GKZDbkHXb2dNxMgn4ksBl8iE4mkldaXd6n4T/OtmNDIcU+1IcSgCRtgffXSl
aPcyrONRQh+8+VnJZYqXiOOvyGmrZxnH3/suojgxoEJwtnIqy6s2lWkzMS5m
HHtqEV05Yx3BTzlYKOo4jVKv1cOqtUKwBgS9C5qRp7vezYrnfwFYrqEStGn8
lbav6o5NBHYYUzy1WXaiZK5CMiJpuSG78pq0IYZN03Vkj9kn6HvKxhXHLGvD
hVlpLepVPP/2gJcwp8/kys+7HyQ5NvGJLNI2zyq+W22sWnNJpKToiBa5vEqM
DOdTA49rmY5ignezuzEWfrSt0T+F+KdkW2YwZJinoE9G0pa7puojcSqbd2/D
hlD+kfFcI3UVM0yl7fXAUaTgyIko9ifRWzs1qSOJWKOcaVLZRC7T7Ic4rXyt
QU2GFHBMed42Kcn4IKsUDsCXImvuKr6Ikq2HGAhuTnEIl6wNjxOFms609zvx
TzUeyNfDXA7nXk7bbr4dRmEVs0WGSw34bo6tumtDC5Gea7g8gHFvkLOLcLP8
3QNcb2W4Lal1P9HYwfZ+BNygEwAEht1sWGs/MJTvX5FZ2dM1Zwe7K0xCAVe/
Qt6VCmfXmnHYX1utNpk5lThh3fUF8tA5YTAuBcEJ9SDDw/XfXF+9FTqK7SPA
5g8nKW/JUDmSw5BztME+Tl2wy5mIDqTUOJDjzYadfmxPvEmFaMatCed28hGI
XArDLM2uZImVqBTHFknEfgdQKGr87/vcq0/wYAM4w2z7px0i55zsGqc4avKA
/P60blALHrf4dw5B4kbcaO8wy9V+nJ3T1oZPRCZklcBB5stsFJYkYLqf684m
1VpCBKnPfXuhxu+QcV9f9eecK8HQ7YnPYXaSQsxFZHDTa5SiRsCAidwfekyY
FrmRDuVViCna6rHIl4FIa4sYNLKiCNuscpLsHhG6Eih93wl6wsqlHwRPhlmH
3KYRTbzu5ls/ZSb1jN3DhJOcPMfrjWSqO3K0ASKnbiAlwEmcfSuo0eB1MMtU
cr6rJl2cnE1xUIQAr71SadKJFTB1WYLIG28VYHEK0F9s4FboINMM9ss0hMjD
uc7RestA7y6ugtRjYgBNAkk8XSgfOrtarKy3kiI4xNDcN3NcAxIHeUrO/md9
qgFA/I61aHKIsGfySopvy1nVVjwiikZYFhQufaXXJx5J1fXMtFvqD6l2VMAy
JRKJH/Dapz9Bz6uALka4PvQZjK8RpVwfxcZTOCUs3IgiyeYNUZXle9iyxcKt
ujAhjtW9xsfYHfyA129LJ8lEGtq6x9uCs7V3hjrlK0Kd/3NbPB32VrbV7g4Q
A1/yXgTjfiBBQPEwq9DkN/yUMLw/FOL+ePwcV5JSYIapEtcDmDVJvcX+P+3J
4ZxSkzTebKdJ9DUEM3FINaAaXsSO3p5zqlLYfngvFg7KCINyERUMHdJOvdF7
SbTvKPwYHOSBkrRV/Rn32Honphk34o8zUaz4kilsXM1XWdh22wNC6rgyzntG
RyRSDpqEhmUx+VeswhqayohzjTU3tPpxngg8Kg4KXX8T9+I6BnV942j5fI9B
gGPq/HC4tzTsG1zEridnj317YlFBUvq1UydHAfMdxm3XSh/NG9bRyi7Eyjr/
DgjJkBiY1UWq035cgVKFW6B/rGTGKgHTIQ5bu+wTls6zuza5Rpx1PvIehi35
FxBbi6z+TXbpAHut46CpT5YSttZ5f5rU1y5KLZQVu/XO629ZahVPZKrTjZ2B
aCpjuZPhoPZkQf4MPdUIdz2N4qScF/3Fex5qMt9f03PHq3cTXLEWRxS+XCtn
9jWLYikMZCH4VVIQPy4VjwzVyZ7BYB/77F4O/VmSP/BlmEor6DSZBIKy8C04
DjVaAvPCuWDN51GY6CTa7EuXjVkjBvjGIGIrcniOQ85Wah868XLoWKmWWPmw
nLFaunPuT/vY0UYDq2sUCvBPhbg1L4KpKcLGu9RSSdV22hz5GDmlCX0fiX7p
uAKTyT3GxhQctuMHP3x9SDB4ilLRlgWR30SgpsVp+IIOVcI/g1AUCSF+fafB
PV4r+WOElx8mvbTOubLt2xmJDo6WDOL3wNYYXfiuDS4Mdnz9FtRubVEvQhp1
qbY88B+0dFpnCxY5uIUfWiwxdLc5KYblJ7zbBNHP2O4lIqFgVWUHCCoeDb9f
eaPJqZaTXEjz39K7AsEE1cN86nD7YfMD6toK8P87ohI7MDg8BWuFdiMjasX9
8st0oRc8oEu/fJsymaAQue9GhpvAfGUnui2BiXvs6xECh7a7G2pMXsJpEREv
pPffHyT9g7gjuHb+57tjZQlcwjy1fmV9SUQIDM4HEAgKX2eR6T92wJWYafuy
0Xr1DbKFUFzqet58dfnR4ylwVCsJFMKCH5kYi7WM5Bw+f2bynBOGAXbtWzRX
tQIB+Bk1dKNWAhajPE5D1GtoEmlbJAf06hE082RseBEzzeN9JvLGTHXzwkxh
5JabQ2cKEB3qH2ggUzKHhhB5nNfbTnpLNEvx8OWIYbey2CDu26cit8I9WsII
WGLfZMJ6FrDK5GQvsMcQtFeJGyjjmu0gDigoJd4RFFWO7SjmsJR6+R8yPJrN
5eqgZqLz/nXkLaSbOd51DWirNLfPg2bKbMgYTeHwpSTKXmjHvX26hWaSUQP1
/6Yb6chxtY1Ym1z88a6ss2E3WhJk3yF6YDmJJV5JUi6MFv7g2lAujFnN0LkU
M5KDX0RpNlMf+z7aGN8l218OOQE241IYa+mWPwuVsOvTWay9en4q6/8+u9dM
pmjodHfeGZsLASt2l3kVuBOOAwZTVCGQAjoMYUvVqXlzrLO4F6slbg5tc9dp
/Z6iFIkL2Yrbmw4iKLFwxp0DGdQbMj5lAwwFtf2LkLpLqLYiuLcseuumZPdW
x9zbpo/gRCC4Dxp0Aj3d6vmAeMzDWVV4jJoa2t7Z9DzzG9df5wy1XlhVKf7N
HCIlXzktlF1pWDyxNPR8Yk7nyj3euieQBNzvpDl7+xMnNjRf4uaqa5GcIbgF
fI6ZH24BUNpQnjdvcKb4mtATq7gXsCbq1fUwf0Qq5TV7dq4vMZd0A9kQW+Cm
eYom7D+PSZNUiwhUB832KQUmCQafoMHHkxN3OtSdzh4eKcND8D9muWVms0UK
zHUL0lin2I2gmzQ8ohmU6rE1ORIS35T/CZHiORuIXOqHkMwLFSqE206fFj4t
v87cO9FpurpWLAgM6JTOn6JzKrljSKX0UHrPyFGx/pGIuJaBYrhqHmUug8LU
4tjGYJbNfT4mlNaU2lKj/0EiXJpG6aEMPpG0qrUV01tNUXJxIsed9eDOlbSl
Fw33bqMM4TUvAvc2L5eMkMVR4tdr+lOPEEsEc/A2JxgrZze9c76bEz0S+1ed
4W6+VJOBS2D7n1wMH9Tm9TIX8Yy9iIXgR3JyP1gDwVSY5hm98vjxebiLec9J
O3C6ecCV4pnviuJ3KtZKlz8D/FWB+RzifBjKzzAivDJmrnxIbMBMlcQbmoLw
TCUFJcn+azdA76IMdAODQGBHsrw23botwDQ6KGY3a4YHAjyhwxIhtHhLaflO
5iMuN+Vuokx8CFcN2HxI6ZueGbGtzLBN4skZEHlWauqLrfG3ODiNEaBRIPnv
FQ82k/GSPIg8Ob5+P6MyMD3L/Ro6Cu9kA9mA7iOW6HZ2dxl0MHSMhlgLbygP
q7LyaVOUnGraSWq4BNmo/9TL8fwkD8+aqx+anf0HXLdnKAzQZyE1QCZoBs8z
/x2bIJtViZHgPm/uuuOJBaDECkCWlpqCBPa2JW8uF9cGSQZxINdV3Qvq7olB
MT+tXB2FuVwxq4SKlyOgsIRKu29o/j5tkJo2FAnNSRF9OUlx9JFukShUiPvc
HxzMUT2CaO24T4La15nroGMOo+h7BdjAAq3Wncb0LAfOAqzBQHPrA5zOM0sI
hOe+E7bN0lhcLWTubWHW1+eVi9+MY75aSVRCAI9Ik8yoBq5yndeMWxR2fMD6
TFCMV8yFPdJzmq044WzJovXd0hEqDtK0tz3Xm8LuCKtWEh9x+b8GlDOHFvRz
NBGlMFGEYlmHDqXstP5EELP4Pylr22IFBAed1GzPPV7YxzfkmnAnlaLPGdUk
kTW/ABBxdfv5DrCKxu2nRyBdZaStkfOz4VUwS2MI7pO3OPtB5qEqKNEDrbbJ
XZOjDxZmT4W9yZVVzdt9u3FeZuNlHPYC8cmwq0V+QPqgN7IIG+6iu7vX2U+D
YctMWXhvzuGSendbKzB8XhWKmtpguQG4m6PScqn5xuPD8kbzB0sn8JCm7OxQ
QfWWGuEpOA4DzJoKfz/QnTO92WHD9d2Mi3fZksm7qHvbXxiPRajAy3/XKDG2
HpL2L6d8jtYLC+/hPtkQD+x59/p/gMGtIN7UQm2gj28zozimATh0A2bo28cp
ejqUrKJI714jQ5dLCMZaHCMNx94bfk4JXwWsD1GQaviseFUkDeTnE2k3KY5S
lT0Q9q39jFPQWlPhLDCbB8oqrLM3p/YgibA2cMK3xJ3A15OdQ8k1tTpGnYcy
iMXYNqfZUjjB2A1/flDWXA61EliqwKVw4FQcenLaiCfrke5UoGJSw/wKSYDt
YLi6RyF1W27/GNsGGG/lzZxk9f5qHy3hOqbE2HS5KpTlfBGFi4WVgRRj/gQl
lScHoOPEMBflPBpWzbccSaFvyITdD+Zb83RXwXnDz3q5Bb9kNaHmTL3oGiR8
2hmy/UZ2yHwtd9q9MLpsRBFFzwbefrvAjvzr2XPZd8CbS0oy36VoI4BrKK2u
J4plmFSJ60Rikonr3MWMmjDmsnjWCPfV4Idvuw378nmJsZbGkxMgP/M3qFt6
K7QNVWzKrJjEuuBOaEaNDoczGyomjqu7HOLZq35eIZwq9Iv07oHrWS83Wuhq
8YyvH+lEQyplQpq3qw+hOCHO/PxNT7RgqVWlc+3FPucyzpjOciWdoWtpzqs8
whcLEsENaNc6+8QrIY5Q7S+B1Yp7XJJFUhCrkwAg5SEm7tWQ19QIFdBvja9o
A2hwxcLlBiUN3CPK/wqengGRApJzrUwbgYET+y074gS+Nhc6T5L535i06Jn0
DBPq9ZEZqN2idT29ZMg3I5FgZ9PO3f2yE1Z7rNt/oqNJ0218cQFz6NySwbVO
pcKoYSlCnKnGloe/YUdC4kC9L9WhNx9+XPuSee/48KjPz5DTLA0quorHJV8l
rLoVLubsBzFjnHOmwARAfoG98MBhAEx+1TUNjXGcDjgykQmaulE5aOUn+lQB
nulHJD6JToWVkGQo26alPlPXJIfFGiTyXrJ5PPjR5tEY4BrRC72DltAbsQK6
tb9Q++mot8vVCe8JaIUWN9m9AwzEO/zPM5qo+q3hnRmEfkuZMtD2YjNQ0zgT
FZFVIxjDj79g/et2AnOepTNY8bZTjO/b3jXeEhAuCehNBSSBWMPmL/tPWCn+
0AUDLLyCSPvSRYQ03dokFW6r9fZS/jWTkq01bUxLLBfdV2ZygOt8INDOwDBU
SI+sebZqsm/Doo1tk35AVZqQ7XEkhWs3JdlfhhanfIO5J3NzpifjzPUNaK1L
SNd3IzHVPl4rJWCIe3Sx+VHqlcS/fnf7Un2b5DUES0rRewamjtYCScTk4i6k
tPSI0AmdDuWXjHWXg9fhEqZlIXq4JNZu9cpHPtCz5izYqAvcVjJugBy2OtBf
vrSr2ZuM0IZR7ajtClpnn6XUslb9uIev/wc71erqiDXCkWlrY+ToON49yO4n
ECBEDhYlfcE/UJ1gChYPiKG0R/9u6bIoF1h8HJJTSLBmGmSFhVivwgCOoUbV
nl23S5OY6MlCz3NADMaSvPXvzLN6XxcUvtfNfNjxnM8wMIMkvAiqFUhthq79
0Y2TnbVD6b4J8SzsBa9rmydaaiDkA8AioRvGRJ46352K4dTKjpTDsPKtZSkc
y+pLZcBGJYjFL7w51smCeY7rHJz/Kr20NVU/ZOtnKuzqL9cWUHAonAfK6F19
UygQ2PNm9eWr6dJ0z91sddx51TN6ib7RZBX7Bn3N+Y4J/k2p4v1Feuqpy7rN
WMo30vlz2vfl5LKCWLdpoQZ/BRKDGWnzopTEMztoM/f8m3eTjO29Vl5SZ4YW
rca0uLDJ1+3q/MQiLpNsaDA85g/rd+SgyQSqzw7ZBzqWZLAjvaGtMFgjTmhm
9fVbh1RsmhxVVorfCh6vkuXqP1RjcLDr5u8+Z+Q5BpWJH362Wv7G1+GYHkP1
KU8twDXSMClMD+xCbYDRhzkRYQeA/yeH86dXzI82xexhRAZA0HsIlNx9utv3
FWit1MJlXch4Mbvj7cko6vgx3dVKUAtBERnSQTbmrzd1n4wH6LsL7w3NZiRP
39TKDsEQDdw1BAhgPodaesEk5rSquigRMthRFfTgMVb22wIMMOM2td/Q2Mic
JvCogWMIAHkJK5HJO1kABe+xps+ykpGc9Nc6RVKxQRyCJkwsiN1nGTbWumJH
SRCGlRwTZJnHRNwxnSKMBTVvBIapVOlozSUunKoaXkYJRjCwuIJFD2bXE/3K
7MY7v4c062xhEQSn4L+TJK5nc6L8mEDHPBIGThPwcuCvaXKzHt7EGQvJxRCA
DulJL+AFSYU9CGxFuLpYqwnv4KQeNPxgKadq+D73hrNoC9dOrPyxJ9xCODPP
vu7m01XWDgZkqOPv8odgTEyVbK6/++/53DPlMCyKlVR1V4NNrTeKkH53Vc+s
66Gurj/pnjXvmL3O2E2cSg6NlKEjleEwokR6t5pnhL/LsKyketEj1+lP/k8P
7a/kEkCFuMZ0UaMAgHJTpZYKtMo94Zli+adLEfongVjE0WXxpLigq1mnvLzV
4E9bAb5N5OPJeRxFf4L27LhexefnsiGkX+YPwayaEYyv1FwkJ5TEEKOemUil
VC9jTPCDojXcQELLRmyucHvXpyoClHuoM5as2LjlGh9NoD6r7wv6pvtrIx12
Z39W+iAQHzIPn8hIpeVhigrgFpm1s8eJ+70lKB3NVG4HIPowR1d9MBRM1Zog
QD/jZi9OmzIlcpGdf5QnrYGCquccZAlGrqg1uru2BJWRqJM7YtrDcYL6JrFR
1JQeIg3oKvsnTldUSf1KvHdMvRWWeLrieklwTruscHHjHkEpwL6aji8YO6/k
EkTEYDcBhCuwcCQfhxlA/gJZuaG8FrmsQZgwdAZAc45OAqckaN63u4KHQQH+
fKOSZ0BSve2p5DDfEGGpTbtrF7gAKLw/em19K3UrsleA4rMq//Cqj70LCgCi
GWwdvcubixwNbj4oLQRK5oWStdUNSMW/s1lvPDqC3PgJQplRZTjs7T1bDwdK
iOiXqcniIAJgCutsZ/KgdqNbKAao37vsB7i+kUw6iiOevIE4KxYNIcCCh+p0
eaEYOHLAialBmLJAD1XE15Ti+fKh5pIsZYLSs8GPGL43+15NCcV8M7CfIf/0
1dFiMZb3aPx9w/wFrOyp/SEKnZJzOPv435yDDKDnC4LgvCf70q/oOTgH00im
5M5YroMCIDByo7QV1YNkavvD20GN0LCxnU7xKKgbquTNSO/zj9r4+qlg50Yz
2LTSKBqLbcWerbyf89wW1Hn1xWl99zd6r7MCCH8pND/vuSru9eR2cGcIpzwG
D7BeJ25pJ3OJkDy44Z8ZZ424w5A8Dcig4t951MByd/NbUFMrfUFlugSCPQfd
HtiQTkfd0uXL2zfUOuq3+YLJQeenC1hrH5Ic/uwb45Bct2zXtZOulzFumMTX
t+7+DHKGtM0PdJ3yMxVFpcbI+ASyWjsMXh/5ZgrTtoGlKgGeJKxvXIpL5LdV
kqCGhfBpXf/kWajoyr4oQFJL45L+MUZvYdB04jUmFXoXLgHLkIYby6z4Hvfb
q4B31Fv415SQDElbSGyGpTCwrw+Rakkq/P2Fx2WaFoGYNzQQFlgNAFh+Zb0o
pWK8SBEOfQHw40cxK9Jf8r7rBo51CgjtWL4RKGd2cWMQSbaa5f1dpeRjfepo
2R/whvJKciaAS14/L+TCS4pcoJuhI1Tn3SH0TqFi3DPGS1dRye01/NnRE6KB
LKf0D4FAU41t+SEZfSMqqu4lrMhu/vxm8BcNZptafI/bSzuCZFJOU9fKrTQR
n8G9yR34G/bNcswdJsI4grqCXDm5idwNvstF6LWn2S9mvwY6qdL0Kh7O0J4p
MjXicuhFIEi5iny4+BEN4QhnoXAy/anjgJmLxqzqUaTxoWWmHhlUOwJuczJK
WRwUNPt8dUbUFL8t7qM3OPeRthMOqu8sNN96fkExWZwZ3zXFwISvynxzWx1M
1umQDI6LuPZ/S4cjTs3JHRuOaGCiLJNCemyasvIqEviHX2IlOGgOE52XYUjt
bdYi2zkrp5ake4r/cZea1DFiaKbc4VNaCGztrAi8JjaA/iC6dFDAKD+MxLnP
pgF33B7YoOjrqZ5od7wmfkDVfBted8gm9aOnZpaQN+FEAU0Yy9Ex7+dcVglh
JV+BuhUfv32CuoMm0BboIF/VP+9q2kx/qb42HKvASTrP66mz0gEWJC8w1SuR
Upa+CifmW1svXepdUZ1UTQMZmh/nNdOkXPdVQngPy/K5AUoKdtbyZNTWG8dw
RFzkj8lXQAYjNDT33Jv6QXx3NgxqHPgdz16hsbQ2+cT2oK7566TsFjbLbGj4
mvcy3w3GG1cKB3nwA2TD/5FpGbWz3bMEDPTAiGllfL3vz9uzclTVySZ+EEzb
GaKujlcx+tAtAlsfhojjawAOHIRcpXYcCVqT5TEYJ5OwYHfy9T7JN1gul5+C
l3C43NIA+mVHlz/XanDyuQ3pxF71cdDRDHzj2FiRZYoii5yJDmm+Z5JY5AAe
wfkBslN/kD+P0anOVPbOUeizQykpKeYcMyba3Az2xL6LiB8hyX8UV5f7zcIP
c6Y+9tHFlFOyYr9vhoBmCWuymjTqs5zCy6Tt9ANb0SagaK/YyHozgAYB9s/S
Oy5ZDK/WKsXJhqtzWqcmWBELsM3npKdzoUzWLk/kguKT5gVUt4tPQiFVOsew
2I9LlwvfwiIo/Xx7Rt3VpqGdf8BvEUs/FhpGhZqannr8ew0VOouNm3iLYp2f
sIhpcBKWW8RLtrGKkIZB+YFTi7hAAoszzsKggPL/DzPXjCZ3n8TP7blAv6aw
ikiwA725BCL8Ob9KL7ooatdBUJDD99vP84+dKoVE9Hk3BDmCFgQNd9ugzot1
xv6Ik0jNGlkgcLGumcl2xNXDDuQ21HZVGqIy3J0VGP9/mqpoWNiOWk/vsMdx
RlffrZ650gEF4A8vRzEE/iDeEqxmrcC+LGrqSR68zwFF3MUYY1wo9P7KLWWT
01/8ITYLvKdfRUm1gQCgYuiLHrO6q6xm7vJVtwxACD5FsdeV6BRMy8M+RfxX
uQbfzG4tjxJ9f7Fo5FbwmEWaNqDTGqbr666V9EtGYcXXGHGISSvD43XkoKpZ
SgI9L4otArwUWnVurU5Qi0FEvIcwtNttVQ4KzHTRPt8xX8UUVxIwXitWZV6c
AORmDVVT5+pzVzFDe9PIKpQ1NPUXINWPNpAw6AbOaafaHIyuDpRMHJ/9S/Af
5Yx1ARr+z3hyZjJEVcIfjthKc3u1QwXi8aBOfgxENwJWRo5dUyn/+BxVGhNa
rszN3hsuBLzv9z2aJSMtaI+fPAJMQ3kzoYGyOofR3f4CRNpGUYPKhoAGe5Ks
VnazYxv4QbEi8THh+UID/5y1BEVMBydhW1xBOvcKJokzHl6VgCpV/rvSUuJu
FAIFhhYCIcINo2CkznkRAJSgOKiYY3dIHR34dtSArGE8ojMPJtHgVyuOV09j
po1oHSEYtkZEos1JQ1aeppRhIvQyw9WVWDxN3yTTiYjNPFme/1P292AVCvYW
qx13XN4GS8HSBHwQSkiVo38ptc/xOlAAiN+64NKFuev8Gel1DLIZB7Li4Ie+
HdaOH8N2dyn87t9C4EG1+QHcknTBlrPNgTM23j7PqyC4A3c3jiXw1DdVcYkI
J6Rfu2RjOJU0M93VLQJvCdNdgp1IMXN+I74RB2ueOcSMWiCfxdq25cILEX7q
oueNT0Jz/S/XwkQaizxi6ZrPru/dGjROKXUFQ2ISjkMLaGvHWENmVRwSlFGC
7TN3L8+VZe6xLY/kPa93zV3Bjqt6CyN0dtAZBr0IyfrzcJtuZ9/+2zuUXtU+
OvEEjuEq/oBACocAKV+wQD5U3/vVfnNLHSFyNA6vgDTNlpICF28KEvlGnRIm
qPLki/2XuUPQj35APOrrU+NOPAI8Lj9gYVfOu0nxrOVYV6I61O0UQEO7moS7
MJGppMvcy0xK8AzorL0IWEXY6bw4i4p45EhvmByMV0hIruPH8VzeUedpWqQI
r7+jlenMcMbG1AGnpylx7nuT7MMpFNg3FtXFIdNFmv9DfHfjJGn9eeqA2rsj
TINTGM9ER2MZNFyoa+ymHeygvyOvLiYGdIPZ8iCBSu0R4s+rFGhdWtA06fLG
cJkKrEhZhVaAzQHXPsp4NEUbKnwbtHBx9FZ1ygV4Bc52pNbELJM1csi2Ehrp
YYb340NFnaaWOR6HGh+rPDf0r6INrCj1Hgsu7FPNF/nNELcpM+aFQns0FX8C
73wXf12AJoYSgD5ToKQh0bfyK7l5Vd+w9N/ldX1kC++lb+YCM+GoRiQ1coWE
UZD8HMo6K2mUhuf9F60zBdgQjDg16/zSo8JCBmxJADUsldG4NK6dJCTzKbRW
C/0SKpd3+A5pe8e6YAxVWFzO8gjdtY5yPDDwmDjcDMFiW1uxKoVjnA8qwKW4
NkK9t4rOGeCo13snjutwdLTa1WCIlqAZ3SHH9s1bfLt3qW7/2pGf8I2HgIiY
1yCYfJjI1HLGVkZLNLEF2xblHNS7yTC0LkzqFqgm/uD8kMBJysVFdxZcA/xH
OCh9ssQHmLizmn7sjGRxmUiSXIDwkZ5OaKISZjOuUjuI3K8e7pxRDITBTNHl
sqkojHJ85Y8nAq8ZKcQv0YkGCZcGynIMwtmkHST58LbnNmYgvKB1YKaQ+V3L
TYP2uJWj7ywhVQrH9Xf/Y9GR1w25XzjBVAXGs4nYUlcRLPWALfXgV7QWSpRN
Uyvv8gpvhWDPrfQP9JGlmy7JlDYOWAPYPHooTkr7K09R2+pgMm9hFAgS17Eo
aJge31+M3mQOtxxDB5R7PJ6fw22w66uvplNVgphdii3z/uPlT+wWZXuY4Bp3
ANDfHRYyrrqanJ/gI9yIMoETM+jYLKB4t23DGPJKJZWk44ySEv+LjBgOuHgE
nEEXifxE0PFZyUaTbrhdENb06xBJkrq/SA9VhchSsFfwliReEXoDvAFAqsl3
Dp+SzheMaQguhvbG/wk5B+/xG51ZQ7Yn8H6ywQeDDiX+U2e2dsqtdImMTjKc
v5VWjMm4tJq0JQ8QGwWozA3uhKKxvgxZYcw348yqojUiX8pkrubj7SibO8Bl
oFf/Yr6nrNSoDa/FezTHa7ni9WY6c4SkLA+3jg/ETfC6a0hPigt/jIYwP80Y
uHmKZI7mgD9pWgeozeSs0GFhYf/cl6LIdUalfbCztLlCCRiVptn6YCXjp++4
R33LnVeQIfOceCiEGNrVXrqslkCifD8+B4tDqaPu1puf3EmhORKaEvFTDjuC
+NJwOaxgxfjSudG9OYEiSwyzyyf+QIaXA4PwyCQndiYll10InFGNiFIaROjv
frCv5+xzq0wfIWsxTHltOx9KswvmHOgV43TWxgiJ/+q6L0hXSOxrwvWrkvCu
aCeOhNNtDs2NTu8umgttu62g5+Cbkpd+2bazA74HajR46PpBSqLt53PEivII
Tshvl+Ledw8cIt2Lp+tZ1wW2yc+usTUoHnZNys57dSG6GYKrjn7jIueIE5z7
xZ7IfqAd7Fh7aNdxZzk21aHX0bT5qonc2BtNcYEpqxJEs6MzOFdCFueprYzW
uiflJdpGC2k+dMJJLWdSXUs8iEfy4/z4WLgS2Jkcg3uPnWaeih+5su5WWG7w
DnwU4/X4Gh4TkCShnP8jx/Zp2JZacoJm2scZ5CEHvH7aAh9JVIJ/62QZgQJq
Zs509T5kJYfzlJ464i9eAN//yi9AY3LMMhR96U5rgLyCYUsPHRGDQMHp9Suw
fPA6iowUuKWTfaF6C3X1CDRo1IXLgaqrt1wjhBJtVxC6oeIZlmacOyh6i6o7
psGvdI4tsXuMBzSEsZHmTo0U7yK9jE9XieZL9MklrlMTVVY+l8h2YfmdWhcf
no6Z2XLU4yYuuSmHqMeGjq4k3W9TvErSdZ2QboKfLRKxQ8zSzXwNZvZczOcI
oXkPJD0hKGQx3E8M09j5/KISkuZyqeH/FWIpa3d8i+U6HqCsUl05BlxL+qAR
hwhvITZC3yYMtg8xRi5GUtek4+yLD/sx1ZdLWaEqcUNo72nKRYI6U0Zqo21e
VQxQ5MBIZWlhLD6wooQYkpXZBcYvNB8bbaFvmqa/ejlHcV0NnBQkB/4hSDwi
G7BiUFx0MXda+VB7wwlkS7NYYsspZC+3BBqsLLwyuXokdsyD3oXYtptbNzaw
6rtTtMf0pAOd7/zdMzkUad8qjkQ2dtpyJQaSt6o+aKT9kPZdXX7qSsOnGXj1
vuw4WI1MPTIk4/4eIUXbjxMDsX+LWvI1At3HGMCg5ClP+MHK2VaVMSRSU2Zp
n7XabVfDZm0GFFPp7/Ftxlu3mb7cazWSxZlWLcbdc3I9RA0F0jEHYGD8UWM6
o5B5tJ6IvlVetehy+OWX6dFW2pamzrDp7WRQSTaaw4KWUX0jg3toRPhiYet+
tuDLSG/X2x6EuDrYO49g8L3E/kWuLvuz98XNe9Pn3joVo0mQCg+dWNwmFSUG
XYrknUCGfweyN5b5GnoTP/xoJ9c6KQN/SXytefq9sqmhQm/VIb1J+aVOJKxJ
0TaMHCMhHJuzKaD7VxIXMUlJcrBagyBkvk7eCukCrFZeMScKaE23478ycv7Z
g13JEYvyb1ce/igEnT5U5y0l3ixK+edmemKuA/Jf5t1eTSYeXmNxFjBDGpFo
uDAL2p9LH3BoWDljzYRasj9KdYlhCLFeJcQqIplGdoOuOM861rzN0/ly5mNl
VnGqNaHkmiyxeYQ6Bcpt9DsS9LsnBTt3l8GDHah0d7QBR/Hqan1YPEcO2nB8
LSgirv5wmSvavzX01z42YKRnpqoLwpYbZHyuqWUfmXDGX+A6gPppNUbOkFwh
7/7oC2LFe7nJiR3y7SQlmEDL4ZVy93+XuX/m/4NQdCOBkj0XjYWA8Md0Cz5G
WIQHIsyUASGg+yA3TBsCAkjiZSHgQU8LjVfFEz6kKRiQ6poiyXqy6BLcvikC
ERkyz1iR3pBea03G84EyHyPmZAtd+MLYHPfRnFwhbuA8nHzTz+ae3LL54VSF
BZ52PltGxeIfatQHKwfpeZMB7DQz115zCiwJbXID7Dom249qCcc6GLS0ft5T
dIPGMLD+J8xy/eRER78jKilYEdJRzSppRKC/gkTMsfWDklHLNwvGEpUXZn3y
c6ZQwaEFwzRh+tg3lTg9e5iUfwbB5X/PXHvy+a3Teq5XndAy3fpB93okRHHf
3yBzD0uEqxoZiu3uLLOIRVs8WXHxkphYb8TJFhNcv9A58o2fwxU2JYPcqv+z
hOPlxF+z52ZZrwRWNi1zg7CRiBQdrrL+cr7PgeeqWIshMqvzdBRZdp6SOGwu
M9G2th/4f9ffS7VQ1Lw68hT/D1iF9DVE+fZfMvMvF/kANSazLg0CrPysrWFV
nCtvhvDLpb6ouzoxLU/JYZJMRBqAPuM7cBjYxSjeGzR4zbuK6HxTlWwhL0PJ
5o4JyMcgRKY1QuhVXNqFGTQj5dcq/0NU437xiPkCFMO7e1Nz/0xrIdzzOR4i
2RwE5i6deEjT5ofOnBx2u/Ua0E4Fk+Zkyj1M9ZTak6B8HEgtx4kAOZs5f5Ts
723bKql4YPmAP6QFTtGVHYNzlD2btU3JxhsoZPA3bcsTEqPQuO5vWuRftWEL
LPAhct5kAR/EoAULHPE4CVEn6apUZ+DyrLXrQCqaQRDLhyZFuvWtXbCzRZt2
NlvXKOyuHLQMGmvac0KC+YUlxfm0X9LqluW6cnyiI8PNryZYsIgJIki1WK8c
Popx9A4JI6/E/8ySFYVN26mTs3nlSMGpAtAXGMF6jQ/9FgceAtpXZlAs4q5d
RMa86Mx63k4z0WbX9+iZgvCUQ9IEn0JsmrwD0Gcbi/tL1W2E478djtPzLWjC
GDjEbhY7aaeiYtlMJ+6bRPi9ABNM0rsGMxBuWfpqwkap2kGXs/BmJmSLmF9V
xdZwuEpFMbpSfJUBq987oeeDgae8QFmTMjLnSa8HZuYJRx14R3jeEUqr+Hyx
FXxTP6+iJgDy/zoFrQIny5/hoh23SFROe2UeVOa/X+w7t83mruKc5pyNHmUA
+gGRQqh56txqorRWyNHhnPX4MBnvyptT0Tsho6POnSu8L2axv/AUE4KOyWat
ckIR2PFXHyA1Bf0zVpmsr6+IddrMtwLOEOTN2IbE6GSCB0kp1Ht3/pB+sziS
lKSGradyA4u4fZuY2hBZjRvnYjnYAQOnEDd9hqNOm6jAv/xBh/wNCDFVCSA2
bA+YZhUrdnm+V5ahZzWVE4HyghhIySEQh5DLKvn1Ykew/Kgv0JIbFu4q7xtc
/uluwMDF/FJepaTKQGNYYvxWZUAbtBhFr37LqNc3OhFAFRjz8cb/DmzkvYBv
OObn9SzEqBk3sNooMrbrpB4UxZhp3yGbEb6O2uFmUIhlaj45ehlAFbFU1DF5
h/ik7cA56M88U3xAxXghdTW0BwJdjbskQMyWQuNHUnOSJqST4+FSXcrBgaek
BOuSSEA06RK72dbhcmYKaOjWdquyVqldgwBvQB3pLXMMXYYBQzAIHMFICCfy
nPLGN+0/iCM7CsJkUYLESmgJZk4X41QHoJV/+nYE/u8YqPsz0jcFJmyLohfK
bCPmKfOPYKyxMICDM//s36eHyTnH6r9hvslVjR8Gu8GYqQv4BNWzRr1Qg2yh
PWremUz6Ou2b+wRGwjFLozA7P9wtEAXTAmeW2QieNNMmtMz+ysuAiPInQu8i
BV//ZU5Uv/4pk7mzgZkzsiXMp4zzntZoNBnvRjT/8rluNzyYDPOEY11Qiqd9
fwGM6HbGjp57FJiyqUF+CcHBLXJuXx+HvJrzx4Hc5+YG0+JOpaAtZ6uoZv/G
BMPKwTsGu/f6Hq38wUZ2XeGey8sGj0iynzJ6AwxxApSIzncg8Vf6WNnTwykP
TBZcw58dUa+OdnbBSBdR7xIAs8lQGss3GSfaDNM06eBLmM+ytKWcJdZeIYI/
GdNjJNgyubDnjN4OND84JxvaUsXQEkZ0zeuk/VyaiaEwqFEKpEQEi7wV9HMA
qp0sm5mp7h/Z1ffL42ZRJ+jKhN/e4Ly2fAFNBHQ/xWeQ25uuTlA9x31qnmF1
XJLMa3QFnpArNc20ZcC+Qqq4TG0WAFQPz0+tewgo4Zod4vuyhzUxcKThcPBP
K2X98q06ILiX6hkjOd3fuQ3WMq6o0pXRogZKA7LOx47rMZmgYuSYT1Gj1NWj
fNAToFlTMfAvXYGa5E4ZFQ3h6Hx9J7dwAa5CiXyJx3NMDl0UdtSlQD8DixQJ
u9AJQCSlaupP6aw7CY6U6anpATmfkrMv6z/BlKq0+2qpaCqydt+HSVAPRtyr
wbYM8aM/TPN4Rf5k1ped39wPXJUmpL9831dFh4YohCZ7QyvJRKpYwKh+z5Ff
+T4/8cSIE2/IofVXnlx8o6nylCHujZVY399B1eXN+vUQqOAl2paoonZorI5N
usTYuqyE4Fd0w2hYDID4bwHsdUoaRJpfRe8GVxXJg6FG51dkh2wA4r0WiEtP
EXY0OiaHbndr8iEAOAvjdsK8fJ6BaQBH8XXOeXJju6ya9jHl5DSWGHANDlu3
dv7hStDtgtkgZhc5CMuMkgxcWQdxvR8sL8Wtdo0Nk4JgSIWNRG3jaZxWsb3n
Am+vXvZf0nXG89NV8ggG8ktacEJGkV3MdSiPMeR6p7R+79LW0oakanTWoOeD
xCmQDHkoCZvc7XGlJlbkEa56c61D3BQHdfENybcJsBwrZYXzVsFjQ/BGEFFZ
98kz4uiCQqz8MIp20JvcbxByxna4NOsjG6cmrH9cND9n4gwXv10OzT8N+hq9
AMshZMEJDo8u8o8jDVVx+NxQO0+9f67eeSBm3i0Z1aoY2hN1vUcV9XX4YB6G
JkXYjzZgkQC5ErA2nlZXFDp8uZR0WhUJijqI2SwcogDiDQsXOt8dZXhQqsKH
dF8di1Xh4e3m+UiNY07FSpoyRJcV7ZMTcpFWCCwpfcwD+U12ydnUjf1p54wL
MsxH0K0Q+Naouni+wZjQLIuOf4BvQK0/jf6iPqSl52jpAn4clk9SFNHqC79s
dA6k1gd5f6MIbYp91tlFbrIwGMBG7nvNs6CSi235q9ifGhA4ncyy0bGFz20m
XmZtigz3GsSbCziwVv+ub6wIfCwhHltrfULZCyLBYmVrHdg0KU3lQIr0qAx6
WAat/OvvdGW8hpbRqU3UUF7wJzzisvPYGxxCeJtV0ifzokoJODak4nUUJVWi
RcWBA0FnxY1Qpg23oo4kdpKnKObwU7Zhbub7Yn59kVhAIziRcP74nOHZS8zz
7tYcdSsskSJuE0Eg9uxExC0cWu8ZD9ua9GxrCI20laKxFkD+08prO7vw15x1
HUm/C2DrBtWXvNXNR8BZ4miF0PazzhP+XtUYupV817aVs4zhZB8VhpuIZyZM
MlD0frnM1QXltIz2rhC45HVdyxj7AC10cvJnoN1BUB8lJW6lYfhnPIB90bqW
b58e22QSzwQZ7EdfCrydZf75cXouQoSeU2UzctEtbJEUjhM9M/1dhjkTaHZI
hk4EsH3bdkq7v2zP1Yo6W9qWSqZWdwAndvrTGOTEHdfjwtlESn+LrdZH0uG7
OxN+1ahbgBsV9KfEGrjKVSanTD5rZYprRT+ltSiEqqgCJa4ObaZccNb73Yv6
3SrdvsZjMD1qrNAJQz3+BUkxfLSNB9K2ozd8K0WpNMXf91gjs6UVCZ4FTupt
wgwOleafqLrRzv1t7wULmG0nHKyNudF4Ik5VW2GAu38pmAfNl8cwHkOhCMoT
ldAdOSo1xwJ2sQvR33M58G9YdeevWPkDvoRBMyETqhrXWFWrlbbt2g4b425U
CSLPhK5Y6BygbxGjdyEHfTX/xrZfr8vXADGquOxXq1iF8xarSOX9Nh6BmPJy
w94rkPg101D0r+brCZBtVeuJ9ZuPpJhlhKOTB9OKYpg0VkozrkyILu1CLqxE
tKrHWVPiV8hRLMWl1N6vhuAe2U3YgkShRCCqJruCiaJy17kCHTxdZvkXfH4H
AnGWgw0J2ZwrjMRMDmOo23nMVM/3t0IYu/MHcOR0h2FsQPIJ+WmGk/XJR9gh
f+N7GvrYrSs9aQ2hbzt6cXZvIalPamc9FSDY1tnDSHl7630J7QtjrVgv2hM9
/zgv06rEqSc/KDfb/xGnx1ew/Wnm1pjv+k6SYn7546uwKUx7DBwk0TuXhEwa
buvRtyxn+EHNJs2LwD7GbgEO9LOAz7d3RweoF7X9TVLp7FPlqQTc3lytMF48
LK8ja4UhRuIPvV+q5l40iHUI6y2BfOGWu19ZbtV6/myG0aX38Oj30zoPzCsh
tSO49kwinHmrhwt5q6LunlWhw/JG2oH1kGycXpZnwGv2+df0cYkWtkNIfEfC
cUWpUV/GP0c2ArHPiWEH3Wf9J4Q2KbZxVFj6JkFP3aR/QcUz86c63EAemnsx
3+eSU32L/GwARo9/nwx35WFlkNmX51tdsuf+JdZru/1lMAO+zoOYqTAjV5Sj
+aJPTXo2JffIlc6MxqjD5DSlPX9FDPhchAgIbUQH8cirJHNBz6kIcnmnFL5O
awtwdUXkA8oY0WpHXL6bdU/bzK9AC2vyZ6xn9j6dnXjIC3fmLcsf5DwFPwMj
O4Wu9wva2cwINxIXURy+2dT9fdTsLOUf5SFIAuygZ2vivJ/Ma2Ri/AVBADsx
lh8Ei1cdbt8Xd5Ewe55dCZpY27V4+muHMBU0tUCqDHYxD3gWwQFGufiC8Dk+
K+kYK85aioTgcrrgnzcK4yHBKgU7wvCxSGuoAF5a8OY4MAmP5kYa2LBLI5S5
7s6x0r6yyQX9WsXjzoGEK1ZgWHaaLXyMbno8ImXFZUjHmEJenvx6s6ne/HEH
5clEHfWXHM6Io/hvXYeZH/8q6qqyRZQ5L7GVFKF457hFWOvB8Q2FNDf77tdJ
sar6ZlCXgjTgUYpRd/N7UXWmGZgGA6ZP+lVRIn4FvoCCiqWttx8fu0bUdege
ipZ0Gwmqf8up2TzaeGe1qtwYMirmCd1ILF0Z1616j8tMYXB1qQ7YV0o4lrp/
m//592czbkfzWCaVLkfL04cRcZk/ZC4bZK8u0Gnoud/ZCVTfjzhwg/BLu9N0
gE9hG8sbEHrqGwjxvyg8zqLN+O3cWOS4yxjQBR3isNirM39ovV6DXM0sGrUA
a6tVPYHvaHM7RnfK35Jo/V0y7YSe+BrkOAnYhlWZsEsus/tOP1XBgNarTb+p
uh1rVX1vBjflN1w0HsbeA+skJbSc//I4rhTxOvO1GVHilEGnaQpr81YhLD7E
L/jP3XTG7K6tQLzkp31wPSwF8eag0sZPGaR+FMFXw3ay/JWXJ42NKZV4Uyvb
pRE5IjIX6NBth3vzFuRtN/Yb89ExdInH5cMQw8iiIyrPEVjuGL9wcJzfSWoK
aN78zLI+EPCl2zjORr9D3uUodoUD0gnPSZslwACFG0T+VpzLaoiKbAwA9QwM
WC7qQknBgaBa6RA+cJx0tsnrD1Y+iO0n1+21OAXKWohKHcwBkWjGBUHZEGaK
/qJde/ok/m2coVSVIRwlipLFZXCVdP1Z+TVcObuPHayYb5Y88uJHNnD0nr2x
aiGdhhfEKlkFbnPGkaryfD//x/cxYUak2Ema4lQHDbs0KjVnMKo+VCxav3S/
qPe1CElBTbY8Nz8x//98+KTa6DwMhRHi0r0w8WzxLXWTwNuptNZM/KBDVDBZ
J6Kw/rrwSTa8rEljVD7D5JIaZkCKyjkIrIIxnIOoSYbtiDXU95tRPL/mHXIV
TQ7tYggBdgFKYPacUE1IpqZC0J80u64JSDOU7Ft8IqX8htKqXN0CRSKH0myr
cJOBWou0K+KPU8YJOrXVr3TwfAnvU1de0bfwjnM8u0aPwjm3z+0fAG1sdyI4
HsKjehf16MJhzPVhgQHpctFU1yZA7YC2YBF9bj5kmECpcJlZxpJid/t0BrGb
aBf8pRc6j95RZZDEmOyUUPgH4qtRph5BR2axEs8VW4LRE00XD1P2OTZSO70c
kQF6t4QDXK8aOMZJvtKL+Gj5tnJpRiib8G+vKunzhYguSRnmhXf+5m6rEF/i
UBoDDcDOiQdr9ViyABmdcIAaA5DdlUV8bUxs+nqOui7JyEpiDnSP3r2QtT3O
v+CZQdNUMVsjhtEEbwWsZQ0Shir/C8hlV+A7E9b9rVeYVy7ndmKVvYpbd1Gy
PI4tIPDHDhEsjVbESSgcYxALb0cR8xAywjUeocPOoGiAOGbyTSmJlNhb4gIY
Qdb88+0/IghmDnxcyvFXD908Divycv7tytxPK1Gk1YTAZSvs0s1qWwLwvJAO
ACzvu8eDHTfT9z3w59HdMyp/kgdDCF+UINlQV8L4djVmaE3gR11xL1lbiPyc
Sbce8O75S551qjogazeJ0I0XurvJ3JIEVt7hIru7pgaoCC6nqrbWQ1uuc3kd
qOasKyb8s6yRnXh1gFz3nsyScW0E9LtZgiAYgsW/5iOkRkJ1niNwQZGhipkD
pahf8XTYX1Dus/7WImFdSVxTyMcdTY2nbck/PTrhHSSg4+emBX4X2ZTNTb8I
e85bE2aLFQ30BEKY5l+1h+p2TCCSGuKUOitSMs8Kqkiwxg0ATcAk3OJgd3sT
SFw1MqMjFT0bHzXKY5zxeozf1Fi5Vwq2RA+SHpG9iBv/s7GGa1RlZSVoai/Z
qXLmfzOFpVnefpTx/IUnV/n9xQYJTzoKcF43KjGmY+/NeYRSknWVizEIUZPh
di/eS7W0L4gjtyVv/+6DJ7I6yn7jNWr3sOiE8TMeUQDjihveFU1GVqNKK6Q4
hBL7KY9qJzB+80h1m2swLAYqWVTaU+AHKZQusDFCWKP/hXslKeY+5NkvoR0+
m7YbOQctElbGcQhbuFjYO4w4BCS568VkJ5c4C9XlzEy9hCbxQhOAI2zkpEpc
jFP91Rh+xv8LYCY54uReHwAhFDsQ1uRoeNgCM2RuLWs7wbssW87uue+8lY/O
8LqSm3d6uBa7WiQHyz7Roe/mLk8bof6dGxLyxli6exIXLZyA07WVBld9Uw4A
NZeJyKtNY6tNQky2SLawJaIJaoNfMQLum5A3l7DtE8iTL49YUqnjuv+1eRzk
CZ6ql2I7coVBZAv/4F2e5OqtGncIwFIF6bkZ0V+nBZdYPHs7T1ANtRN0hJYf
Vp1cAA5PRU7mSWNt+3+vk+u8aWironN3jFcx5rzPPMQXw5rBSUTIOJSd5JIK
8UtYsudGnLAqnWQD/9j4hpcrSDpoKY7CvGnMP/q26DJqS/GOz6LohWd0LLAv
LQc9EdI39WMVvEA+79gC2LxWhbVx6nzzzlZW9xlA+Zt3aoTO9SdQUtzSf/Lp
Ez4FphjO7Q7gmt5OhB3m2qQrFR85tnHnhFJyln24O16oDxPSrARtNeLik6N7
ghec3yvs7MDb15Jg1J8idtA8JLrfscAHU6eSO71jnTFYQBtHCceuoEiUP9ps
tdCfzziI5K3b7wOisizDyrZAaMilHfksQhqwCbPAtr4hbWEmcvsYwrCp6P73
LgmsSHqbgzRQ9mNGPTkadTGTh77tma6rEG8ji8m2XfVpnlbtW5FcB4iE3UAQ
nkVHuywfYLzMZXoQZnGHprDmnHSgYQMjYW/lHCij0NxOvXqGBCCKOSm+jdUo
Y8Is61+Z5OeD5mMoxzXkcCBZyZLQfWo3SUSy5RXkGegUDE7idxSjU6HzSdM5
aW63cXeYFr6kACnZkpKbBmqlrIzoqFkecM3LyIapRY3HfEVZzs/yKGRswrfl
rkvOJTD4KKAaW4pr6k7/HFuR88XqHZ2y1gkQ86prCiGfqYZYHIWncdHhOPfL
d6EyJAy3UngZYpBQb3lXfoopmcVQV/Eobqw4B79f85nTKdEFjPQ5Cj2hP9Ap
LZLo/wd0r3mNvNKBgQ1RXCMFcl0lswGZ4W0vEQtNK30+gtSaZr6GrGdBD9Hr
EYbADe7HGFZQCRmYAO5ZVB7liazJFfQTH5zxiVEecK3Z/RGYFplu2SxWOJ6a
qWnhW9p8XI3M5Q5XgqbsSbUiXtCZugGHAfNouuIo9QkVZvcqAW/FjB6ctw5Y
r2TDH2GFVJZrUycodYQ1/wwP9Ixk7Q0vxVZlFQkbLoxesGi3b3JXVoA+5Kkf
XVT1tbgGHDt4YO1Vis1KVURz8Yrk/ZBB7G8R0+PZ7WF6xrbUEZKqzbSyaoP/
rvLYSuLV8Y37QzZMoZe6ZvSgNjIIdIFRNYJmYBbYvG0fsoMiUIbsLm20wt5u
dTgMtlE1EfIxCphIynW4JFO5Jo880MsZB88e32eIk+QFP07o+jMdHlzB/8oP
zo1fNi7a54ozTisqPKmTza+hE7mpimLsqypk1ArSJ/GOF8JAvFXGvm9ZxBol
x+xcv61vyzCI7uMLkZtknSo93hm+eZOc5qTivjLRTJVa1L+U69I7HJu8qG5u
nUUGdeW1FNYJVeRNLSgBygg0cLejzHQr2FW3GSAflkGZQ22niQSFUz+TZMmR
+rQP7jKv+vXu78JDSIA9cuwPncjZ6PDcT0XZfG+Ir+GWLsaWvgMqko0UEqGf
RntemI2i85nWQIkDbnxf6mTM/0o44qtQTJo/OxMegiGLzQNzLQzFdyiAhQCo
YJB03fT01QgPk9HDlInzFW2/yd4QSeuytSEMt2c7uTwi+MotI/Z/gM5kbIp/
WkhbfW8IpXrRTX1Zx6EgGC9/8gkEJ9xrOz8tNOid/I0VEUkc/uXjRVnf/1ht
wKwoUpy8OWkvwOaNlzd5BcPbQGMfZXzh6qDQa+nuicDuZSuw1PPwVwUa0mJ8
VYlbto8R+r/h9eqvSS1Av4r9iQ8uPTAvKr15IBQ4gjg7gn2U6vn0GCjj6duk
LmeDp8g2NIgPodt0OJaUrEaAlaFAn9L+aODPs3kzzR4njpSnv9wl+DisZeg5
8I1iEQAfetFtfOxrp328tk5j9C+SfQHaF39jJjc5eV3rsE/q75860+wSxsfV
ghXJZINM7Mbxd0X/UT4gk+Fzy1+SWIzW9q3AIc8UOz0Sk+w08N3vzgCo76Zc
4iyX9fGbbxRwah0MyZ2dNV1LuMZsvFp0NJa0LUaXURYJZbvMaYf+CGCaOLAK
6aUV2KFRaKJJwQg85rdl6tocHrNJjgDFaA77TStHrCYmhq3XnEvCwaK1g7VS
Z9LwKfR8H+EuJ02lOjKeROB2FRtMUOMtW5iTlmq3N77lM7WL8xhbzI1u+TFA
ro1IezFvClcdEP7Xg7pRNTircK8j2lggawuoXqYkHwk3So1ubUCy/xvBf8Fu
cGnl/UdYSD7THjam8OWCwSAkNXHd8fF1nS9IpnmoPl16xe9ZESMfNAAaknTD
Jbdkr7EtAoiqizwMxJZT99KQlh7fJ8bbbmP7DTXsCUwPa1ngOmubGHzajq42
l4OkaiqMscN6WWaKIMzrknUIna1DfKwFCwRpbcwlif9AadLrPdtuO1hA/coU
AIWR5hJX4hLxjuHwruuDVPymPbOcCeYY9nSa9jTdQkgu3oaHQ+YeAJwY9KmR
+rK++JG7eh9fA0lQidgOU7C0rSMbtOrtsYatDjnYYSjjuyo04xZMsrlS2qTR
pHYYsEfQgCBbuBgbGqtDgZUAMgHjBE9vo9Nm344+47+MLvbUspYN5Aw5JOPA
YYQoLMLQ6hiEU6CY9jOdbCyjzTTnXER7JACwBldmzPvPGtfy56GpwZ//xjWo
6fEX8qvPG1+Q9utGGIX34gz7yZSBmZ2rEU8nZbZ7vfm3PQpCH6c2MU9nVfJo
u/11bbTRm2nlxRZMeRKEEXqh8Wa8NQRfvIfA2/IAJ+IzELqKOAs8nKhURq4h
mBRTBbCgpEqAFSpCQJKgS9Y5E4RGO7J5Eqe7kLLk6uiyeL7+0oFPIE5Wi2FF
irwmZj2ykrUKU8ThuZkvzCMUFdtCGIJa8ARe1ZzYX6kxCL4Om5pkP0L21ZoG
FCio0nQgl0JV6/1yPN2BJv8zOWXH6dqokAKAns2OG/q29qPkry/RDVnyUULL
3zJw673cY8NFyH7dkUOsR27oZOVRYv5eHP1fF5wCI01C3v8wRquxiwvVu9zT
UEi76VUosrpUoG/US33PW6qwuiFQTbQE/jMoRYih8Wa6rEtFZcCearXPWvc+
YMW8WNn9TVdNd89RTQhKVP123xtNwyaTUQod1lrZdWDhUqgvZ07i9UQdUNKN
UvLw4FjeFvUg2BRl0ub4EjRhzzDws5ApHyyLtgrACcFA3d5+23RAeVXCydlc
at0mSFPB4D/w/Jz8nWvi/RYNtKy/SScyx+T2/64XlUtssXO3RILhmMIFF2FG
WS7m+JeLu2l3r8Tl+iV0AHPuNUD32/iqjAD+xebqafwXx4YD9jxyRkKmb9Mr
Xm6vJReERNwg5Ejv3RXG7frLv+2NaZGzGLomoqAyB4zVuS+pkjqkDU/7KkeF
SCuq95IqbYm0FBmJMVgDk+hgESM0bXS+8Nxd9BhpX7TmgWinWHRLqwry/PJl
QQCQBhwtHWHahIx7DHJPTqog19eHgmP2FjML6CZfo6C7wFUiDA2QRNQ0Oy/8
/AJlDrDsXvW/1VbFkvIvrLb8WwVKUAUagSZLPg8KhIiR5K0/bqXn8zl6JbT5
bEmYlB7aNQKB+8Jy/LQBf+v96CnraKuuLJHV+Gx58z0B205EkLaqPmIcZ+Tt
xFcYl07m5e5g6GlBjZBwiAX0RqDZ+85Jzg/uw4cVnWzDwVcXRdO+I2tc1EhH
SKcivcPN6Im1MiE4pzIxddPFGUkJQr78zTV1BR7jorpG6acg8n9sIk4wbOka
L/SEgTDniu+LojPCJo+zuBhhOAE1HANScNDdjxE/CRjZCpXl36CL6VM3Tyet
yMSjV4NfTBSRjcr1d8TnjLCc/tHBKlPq2u4A+xd2y/Ps8qO3gV1USRZkuUNB
W9a4UfemZhYLKoUbCy74iTQj20svoLinHmsNT9gyxyjYLjMnVMlFX01aypzJ
bF+J9VEVKv9KaC/mFxe4Pw0W1sJ60GJPkOVowLuntqOZj3Te9zPtkGSym4bW
ta1NlXgxs8ZNy4wHcX/p2jCWhl0JNWaizx0RVQafIHBk5GXatbCUIoh2nhXP
SDlHRA9iPS7jeaW+PEFGxqie7w1JVTVyowahxyJ4oxugn7jdvGTaKk/5i+13
vUsiHunYFuOqyyb+YCHnTK2IPnYvw+wma6hbyJ4CP8tGDiYDuM4XdaNgf3Tw
yWCDaZKZ6PLhAb7Kbvy4nFh1iWC8Ryn05X6Xw/H2FL0oAy4n2ikfZExBEFa6
LT83Cn2yIQgbFlPwVcgXvqgFpI5jNncqDaDnQeTfEpZEWKXylqrjn8Z7BhZE
5gFPqoAZcOoo4Thyt0BiXI6lfXWIquau90zbzC+BkshtRu7NYhOYLlFZbake
+THFsSd8qw4GnT+iui9UarKTX6ilFj61d8ReG0QHgdXyH+//Qnb8hH8ckRha
5FSVPlvf/Tq/lfgA/LJrFmiEkhnvGdJMBuk1wYwFZAKFPPBWlAvzQ15uu8XW
Y1lytWb2T1gPAkiUIF9b/ZFSBVSM5n57kjN3Wo7cdPoY6TrQiMiKpNicK61c
DNTCFoWyFp6NKND7PG4+7bKbIgzokxMuEVCdGBFNtsni+US57UPl4KkqLFBd
zeEt5hQ8pIDJjE+/1MWJHP4P2UMuH95i3SCsWO3pEf336MqFVVfUtZzqfosn
IisOEwPLIfyacUqBSTrS/93ugF7Ih/+8DcOZgXQNAgUNQYK0VW5PvZoURYgE
GSU57P9ASTOKXpjsDyud1LJotF75s7dMY9YFMZGcfH/xYw5WPPyNArN0SGFZ
rlbNnNHbXy7qka7wpZErtL4Iwxy1tn+RmciP00HuaPdzF5plwsKwEuRrZ2VF
SM+ZF/j2/D5/dBYTs064bKHMTFKbRJXx70hdnPAazNPMPZETK7hrwKlJ7dwz
i6FOnkpTZDcgYNnXYYfU3htw52h9Z+IMqeIQ4aF8+yEgTmPgLQ0TQnRoJyQj
854SCVnyVsjToT02XO7XKzkY0bWi4fsejv6rGcGRUaOTYNNNI3csPG8n0Zzu
g3iQChKuABQkCIS0arS6b9j41lXZPIt+PI6vr1s0bFSNQAlgIsSWXTEsL5Lu
nqhaAlS17mylKOhC7MPqSX1JO4ISmjM7E0KB1L+kdRh2e7tVQsHFqCc1QAeR
azCzZks1sHTFzAvcs2xNrooPAlqH5s+R+5d6ezWrg929GVN1UwJ34FKJolB5
KZ6MhSg1Yjn48VnvcSPLubO39tup5QUdEXaQLOCIeWlubBDXiae72bsUpo0A
k0yn/Vob/uiOjOQSoHwCLb5FnsmdfYxCK4OY+ETlwrNOnLvbS05bkOXz5EnZ
9wEYYo6B8Qr//JSGIhTMi9aQyC611tVrnaPjbKbIN/sW0befNf3C0VMilUpj
mJNk6xFBz2bNRuOpi4tVd3gnmkVRZscEcShKAOIzKD1bI6HkJhEqsqCiexBF
PnQoUO8EEuw8himV+RuzoH2KQwJtMBHTGIAI7y+DbDR8jJygpenOPCt0BbXN
tsJ5j/00zKhaNAT7ARVYmO8P4UpWWQrZPSNLZ5W9fCrvn208htHKtJfqJDbB
QxkqNkoB7F3iK8SNPBK1wSis++gwlRqJ8eGf7IwjXPEcfdkhkTeE6H2cA6cC
LnV6YVFoVt7vYOj7oqQey1V7LPRDyv0y6APgFJdz2j3IkrK4YBf1goZkurnd
DofbNxqEGGdNm4sLdCNMQra29O7ySRHooXnbt0JJ14CkuDX8VVoG9qFxTM1v
3p4uvmsH/+lVaaGY4BnoW7urUgnsh8CQvQuUwITOU4RAPMNSMVaBX2ezxcaA
XWEDFeDJ+R7ylfvg3NZ29Di5LY7eNlxvYt6V4ZuWUYpkvUkJIO/WI2sEiA19
wSQBRnTtdR36ZHkwlv9XALdMs/sU5NSxjt/1+lPXjBps3ziAc38KL5N8ZE2R
4RSaSKoOPiD6A932Sl0u6k1iScfv5vHmrgvrCRbjY64ygA/JYBBYXF4WKJjV
RLT3CPOoMedVkdzUeG3kxhVLmoIv5iAKOD6JdrKTfEiLgbb6lU9YkJnu6mFN
TMHZW8hBf4bZZpcaXmbD/tBbhSMJ/TYCg1bVRtJzBaZCFhYVyhCNveFAcw32
Fs4dRdmkAmoaOLx7cHVSv1F/Y3XHfkwNyewkPw6vBfd//dBwM3zpDcXzssHP
OymYAD0cy2S4zbJkDEE+ypzOxYfXBtF5wdqtreqpHcBzl+b0k7lvCquvqzt6
0xbKrOn8Po1AFjITxB9hP4PDNC/xm1EsxeInu5xorNeBzf7NVijON6OTcwTY
LOMWbv5sQkS165x703RF/xKvrjsj6bil63xLv5YhwTwGwNqgKtRM8GicQCAg
6LSf2X7XwuNB9NudGVZR7wBoS5vWYdEPoh8Z6GASeV5C6xbSv1Ify+MbCWe3
nIN0AYVqdRa9nnTVGx2YpA1X5S/ZXfvn0KG/YVvH+4yMnwrbUEghng6NApy/
CRjGuBT8L1p0wZ29JyIPi25YKbtkV8u5F+2a62ZD8Ud+MWT/7VYwIK+63s1a
L9uerZN1YMXYiiInInC/8kM0GtS0m0jvEUhndKj2dSnWqAyumIiGOo7UgNMa
8sUcfPLC5uKjQEk8b//VGostzRFfnfl4Mdv4GeDPXWNIhec5AGyK40Q19Jgl
0XJhCWGoXx6FahUdeN1BsMQHiVDWp/gYdKaqaYV5t4IOP2sf6nfVJDUr3o+q
UxnkTOl8/xQo10jhbWQPwcC2+kftyuZX0QyUdrjTLGnj5K1UrtTdUy+YnRdV
4HQ/i/OU5ED0gPDBfO7cWJWIU0g5WCMtviMxjxwuho4uWCIMGPMIW/e4iOr3
txLnQzvFK07F8g/LZkGlyDKePBacSaGcTAG9bUhLqlXo1Q8/8XtyABTUUmc7
VvJD7rAp/vVvxkApU7YTyGg8eeMCWK9KE+lixiRZz49EgdY/2BH7th4yjnNp
7n9l9QYKPFKhhLP76j1rjZrNoNsU8hSxPnh6KVLGapDMvHsKE6g/Fp2N/t7S
wybhriXca1zi2lPeBr91k/0rZdEa8z9ofDiEkIIbGpYPViCiyvQn8Vh8yH/W
+K5VX0vd4o0tRO6e8sjZyA8TiDQtzjn7K97izX3WNFXk+Uw+MkVNKiDDMuVN
WTJi5FmmqydR5IO8PmiTpogPrhEGp4ebmLX5YMEN16HVXx8P4AhBd9jgm+tS
WqD7KaNO807FQjIj2RXnxMbzBg+M4Rm6FFS35m5P0Wwnp4KZNGHy3bKwufAU
XMemEXA0bKUlV/XSB8PGB7Nlp7LM1WoN7zlEaMSjDCH17TXjCf19Di4rBPVk
gKozdydIrh7E1+84+bNx6NV90yekbmddjYuiPiIPOV1Dti83CNjCHA0t8WEc
GJH4bgUULC59fZyRNLepoWabjvDim7LIHhHzQ6uFOXm2bb5v804fWfOPX2G8
Dr6yAyMWPkJ1uYla3znVqJdqKls32PVdNYKI4/ly06F7IqTYCKtP+nZizKC4
TPB9LktHaHGEtpb6httTmY2qtd6A5Uv7fdRD6roWggTbJ3jHP9k/rv7Pl1CC
DPKQcWeS9SbLnS1MWERcOwKi4UYa6Cv8BE6BNtSgq4ADB0UXOs7LR3K+BegQ
DAiCMm764eDcg/VUXIs4zijm6nQclsixlvrWxawAkjdi3sPUSqSdQz+jJUoX
kzuPvEtF1DlI1Um4GwcVI7jC/o72PNnkura/2ooM9DRBIDzQ+qQFO4uf2Ul4
o8gzE0OpfqFDRXMSfs+/bJWzILwd/9A+joJeXItZK98525bhgbZ4fjBBvYrg
XgD4bSxC4sDX34qxnPSJkmmtooO6DWx8Pbc0AaJZ1GuhrbPvw1KBKtmz15Du
X+RP4UtJT6/+sVY3ZehujHbfrhy1FmKhCc5ERq2imT3LEa4/BYEoB7c02wbb
p7EEvoWYzz+yxuxe5Sal1sq++i6F0+1x2PtR5F4v5cFp/CF9Wl8reluOCGan
mVTOz8FNb5gkhcb14hZF4J5ZYgeKwrgbs3Wlqb95NY54qvPaIFCMOvlzMiBT
8Lblz8fGCTAGi3pkpx7NLbnTTZ2kXXY4hV+i1fk8ZBJKiEahKXQZQUOi8/e4
67gEU0unUffgdTVklUqRuQ/j04pkXcyEZTCv8in+z9KY3IoZx8Yn6YTF/ipn
0j+u3jhh4KBsexIg1XEKIe68ccCrOe2t7nIdc9JTNxKldWOJNCjKcrU3BMsZ
htyQw/UTzlZ2ylRetYp1MexHC/EX2ikAhXPQiU16298SKrNCNi/ACv3agsgJ
eUJ4QwIOBb9lmh+VHo2XMYN776+CI5KGXLWqwK1tehmuSts4g6Z1ePg9Z6Rv
GbcitdKst/40NToZjVYGPXJFu7tsIFk77eFn78FWpY2wz0zaeh4eOr73j/Fr
w2fhyo6IB1wo7b1xp19e7Mzclca4+ptwU/QDVkc+SgjtjWC9BdZ8AySPmT22
iQV32go7bUojUYEv3bp/bX4WhnEpxikKlWIYpnLGuiapbLrrO49QioftnWcj
ggEgx8inpaB+6O3xiW3rmx+pciO1fgsakppA0UZRdCsQJysE0zRk7G8dHYH/
7CkmBogJDPRG/nBVsAZvvFc6VZp+HkArONi6TV4Wtd20EIyNg9toLaD7K34s
5zwCCXwzfbQQ5wHXUWrlZxGN076LpWKbE3QT00VELUtV6oXR5BSd9fx78nle
85rSbZ2ME4UA8kkVW23OVpDNiqm21lpaINvjKEswXznTu9O0JyNno7VznrHm
R8DZrPhNFEaWyI6c4x8alHk3KdXChHnGjBYg1OpKti7tyg0KeeKDropEVnIw
iPDJ+qUtb0f2ZnqlDX50qhVpQzIQVAu1U4xpyN7yQ5L9HNjpRagKrFtspR7z
FWBlDoOqwow9AvrPqXph8FCwCYKTsEmTvIA7MBh9NkjEA5AlB5snhVZbYSiS
JZGCZsbZcklsXkT37IWEQUy5bafaV4JJ1v8Cts/pdoOMhiHQu+2V5l+MkJz9
Qvtn+8439QzXZrgEoMtEi+dnGuVQIFQbBwHYYjt9zroL3F37JhMlOGpFgfEz
KAi8fZRoB7AHpOkbfERghbW/UT3k+Y5eq7mrnjEAePKtUfbZZ/bKzYgtQvqf
DUDTZ76ISFmGodKVbt+qKyAgO0RInqPuI6PxyEGRR1g+sS7PGKfRjYG+F9KH
u2qsqkHZrmtta0SS4aB4gKBjqr2c7WDaPnCe/g2jCKGA1MMe44EUiQcD7433
6tZpoZMa2vjkBLb+h4ouZYgYUOY9oR6HRlCKlX5QGhPEoVn5xsuFoE5tbM+k
T3pTgmj0LgLO5XEcd30nji+oOzDhoMXDIxvPrV0sDZ2L8iKxfOGv2oOtbH7n
5BhzeS6F3veCvU3+Rm39r21YMAlPo5+6TvzkQEoY4bTm9t09cEKOvI33aKPm
O56hx4gRpxYXQmwA6oYrSTrqn28yyrM7rwFtSvlEKwBCj1yYyMjJZrFqOso/
2ZFSt9OexiEEFrX3JyH+jOykY/oS+JXu8fCjii2MZHx1m97gPaB6hDi+VX9E
mffXLvbXzknBjlndt+Et47rp5r3K5jPV8oD3F5rZ2MUihjDXypEw0cg1LstA
cR0r2XtGtvWDPPpX2ZWfOISPZK6yLeD9yHJY2/2tmhCNCE9P7ZcScDk/HMG2
6FqBWd8GwcWLb2Cy4w8mOF7O/pV0/P0MpXcLeYrG4H68lXgJZEuZWunoflnV
puFoANgEnPWUXdalmLhj70+O+2ezn1UdzJscurCawEJ+zkzuhmQueTmJeOEz
a8N1Ey2HLwa+QViI5ONxaPm/a4uQCJ6QK+AZUYx/YmH9mh6cTJhJTln2rTn7
qSPnWYo+zfjcW0W0hx0dkFzkmm1vz7qsDGHGLlXyl/SLgwQKCrEQLx6exsfW
Ke92nrfo3gaP/P/nv7DB0B7yvgbrjF90qhVfi98aFz9Wu02l3cx0M0FS2cPN
IkKv8f2zEFrhVU0r0IBGLbAGQkAI+FU08UduhjXsio2s5+xxUblcn7nPbEuE
IqxMHePQmDjRULTV96lcFOZtSOpsR7sU3ikDR0qMjIbCgLH9ElN5R/tEtDJV
UvOZ0h50zfxk4BzXVtOJVmxhg6rBKOPLCCwhwki49yhgRO0TiFXCyeQuEadp
6nE8zQblcIVGvGc4NjULVEDMa2lMLkdT5R7SZdijzLlKoG8pAvdnNjy7oXJK
l1nGeX6ZqYWV+hraMrw8Q55wIbgQvsOb1zIwYaAwR1aYVpw253IrVaSRLqiU
oa1N6/eOizhFy8Ng4uAvRepV1aZCu+uWlTP7Omy0lb++5INAwD4lzuV7o2FA
ODU5lfBZkT04OEbAhnPC//l0sqbJGuknxuySH0jKc2KwwE39ORuVnxygn3yy
G4ZlCozkPq9dW403EVUIpkESiYW1pDSuXVAbWPYUTQFCeHxhKkXppegMHvUg
k5iBs+apZfHD69Sj/RxkuEPonNtTwdyJ79t7TyjDk4bAgciOUcSYZxVLx6Be
1vgnjHr6oGTjWwaIDxLpYC6vXCHrEr0WUD6jVQEdc22C9FLetO57ekCjAoRF
5UrVpwfUiSW0fkkksdoIUF2mmWJkyPxFUWYnpEXXOHYNJhTEjvOM9nWnINtS
sAI21mTfYeUD7lExmgZXf2d/aL6/ZIpcenYf4pw5pHtZ7R5kbEfY/mVXkDYq
Fc4Ek6UvWAubE+Sh5c/hg1ZukikNMeIWK5L5l3t1DgvXEGsQ8UZ2o1fNnXbK
5/zgXUSp4eVZGfWB69DjZsr/qybzSvP8gsBUvjx1zKQiWbFBz+TwTHgamy0S
g9SHvPq5lrva0b7hToZU+a2i0pwBw/9PK5jGjt0C/UyGRIJBm5W7/tk9wz1b
z8G2u4uuHzCz0AkLQzANtHBP4ZkBB+hR+1kqd8hFiBew81Y5bv99IcSX78LL
cKLVRib0AUxGOv87S5GEscLqWHV1CL1H9zP/SokSx/mMMrQnjw/SEetSUuY/
i4lqxdayfjoT7YQgo+UkPLb70OK4d5gjSyl/LJewYWXEBXTvGAeohqNr+zCj
NJ6dKRZShGPWwbuxywKw4/uRJ8R8OoNf0LERzhQDEgjTALv47hd8bp/cMZci
nq84EivuC433vc3MJM1w5mhM0c9nDBR4DNONMzg63SvZLQqH/+BqkUZxngPv
C1OZOAWduExw1ng/9DB2dCXD3vK+bubG3KlCiYptEmB0oBakFCbN5JCQfahv
paotu1i22V7XBbakQoasW+YL3sagOA/pDyJZdGIe2b3T0wG4XzQes1yZAI88
Xt3cOsDdkYf3Dn18PSyS1MVsEk0Nkj5SZgUkWOdf30ATFy/VfW+WdHPDqTcW
sfmXg1eO7c15ZzdIdBNhJrcCPeo+0VsrcghswFbGL6JQVgHjyLRcB9JaKdgA
VdcaZHj8pFJrPrqh+pZJMNE44gEntSD/+gjkvYe9n/ZzRuEHP3IuXQbX9HMb
J8VCaccn95xiAdhTCoTkZ8yhlKmPBvKHGxWj93RWSoKKskFLnqeRjAktPiWW
Dw+2PNrWY4ETjQwZOaBAF7WCt2P4tJy5TBzleBnTf4LOunlL9a1rbcYn/59g
nymoL8CuWljEDcj8SJV147+i7JO19FCTXMncYCNKXU01ivpZwWe20Ul6oZPl
QfBxtR2ICPNZrBnlX9aU9yodC5q2+bygQTyBKViY4MsJ3B0Voywl/q+iAXXT
G0P4FHt1CBWl0QamSCa9pz97EUn/ZXpUMzcu21RxcwXo8WC/GMLRorcfMkKx
R1Kg5lJFqnGCjbP3JYr6+FEXs41xgkfVaFf65N7aRxhHd6nfZ0Gfba2BTvTZ
mNxW6g/mGVZoKubaSprlNmLyvFioDCoYJ3hwPbJOfhifQi4m8k/n03D7Lf5j
BIm9v01lkMXgtmLBJeHvWeNMPajMfptrjUEdXuhssX5iUgTQ2xF8uuC9ahTh
uTb+GfYusgu8+t7vIKm9bfTyh2MjqiIyylxqRMBN94YRZUI/8XrdWRlHrBjq
FzqNpiERqErOmlvi5DLuRWlJWS4cxyaTSpCGZdnxHyCdtJCpeAprNO9ORPeC
55cycr/y+LFN6W+dUKLV3eO9bYYWyVNLvQfyhybqRfwp0mckzWD5uB2FMESM
Ryt2sGZG+hokHbaEcRT4OmrB3exi1LwFkIgvfLg5wcA+2EYxukTiFI5H2zcW
WxoasUKpONA1F1oyHBv99i/t4hKkuxKMYOG5n7Pi+RYwZKieiJ2LLtNp4h0t
cL+Lu0aGV1iOGSqYu0xCy4WVX8lRxaBGY9kvtY8ncHsRPinKGTojyvf4b3Mn
SVIHzwZgor1wqowV3+8EYHtjRyenTtpsAFNLyYQGVUz3SSNb/qQZkXDdKpW/
JV9Cugn5dHjAKuZEzpTqwIERVd7Zs9Ul2x1jEo45GtFfnbGQ6WCc4BX3EkZ8
oVD5w0akI6hf/RxvYoJy8Ol4w+uGZUIAkezuCVwBrO3TN6O4WGUDQz4lyOnc
kwfoGUEI7oFwlAZW62QuoJNg0c4/787J95QQ1s7DC1PldFNNvtN7BdTdPyr2
87aDCzxpI2JheKlDy8IYpStO4NLf0XbOsSXrPNe8Ni6UdqwAyTUXFstWmkWq
GMXOtJQq8U1NPz20MygjYm+wSKbgnO4FkdsCZIwjDfg5VfSsgYeJCpVR13S8
3/nwrbLT+VBhazvlw6vYjyogj8vpwJs7s5CuzXp2WV53iVHYcipOtCriQaZf
oTKG/QcCP7W2MkvS295QnZ+OY0QLK2uFPWHnTKpS81sMDGBsVI12V6GC4GcI
HeqX3mCF5L1TSKOswFltXvNvMuTy7wdBUHPPkhOwonA8GSbrEg4eeiyjPSH0
B0fJIsqmWYUp2jdZWTiLmQk/IE6Iz0LT/9FoLKxh023fxsMn7rC5E2Z+uYbz
7f6xi5IXilX26IcWeVbYSsbyfeBbWlqL3yUQI4Nqdjt2siYbVlF7zBEe/0DO
cC27lzrGFx9zbKum7Y2zxZCWS228HKADfVbsorinXEFIG1kPhR6LR/Umm5Un
bs+T0ICo/bhAl87++L/rsYusiSemOe+nGrVROCE6qnpxctX4BXy1AVB41Taf
kC+nboQ520GjlhP4tSat3LWNNe+jSJHikNoFfUinIhfOwaZtjQcH0aV2ouvF
28xztvXGrX79xBjI/hPqZbYSdas7j2JmCkDQA2TfMWtvifo0pbS8getlcA5Q
rSz7AHoR7lx6Hnlx6R9f0BhIuTRPvb97C95r4Pepb0BQYlMT8UUIAHqSZiHt
952ZBZ3lUuw8AxU5VAO0A9vR5rLLa0YniAfBHbEY5gJKQLGDRhtop51XDEee
NzReiRtvhKDkEGbtxqhlUkhzv+bEx49vJlUuUNUnSv78tKJtfUEGH73YbWMA
5a9Nvr2G4gppk3y8PGRzEd45F72zpoQgz/hqUBmBXQoN5EUx7MLLON0uYx9b
gN0xuoeImu6Rvi5rjDC66GzHuSZz6cmRoIMKx4TfqtEBg9DSTe+sNM1a9qkY
8JATHJLntsPweAIkxLSMIbWjgwpuPZESG9fRYPb0XIUEXJOUSJ50CBgSAVrJ
bEuE6+dfTqYcnURuYoYIidCwjyB3INzrMANdrrLn9pJH7oG6CrWOoeDmdekQ
huwR4k/yn6QWLkdUCMrKxN2BUtP6EMuExKwSbkWvCNN2eG726O42K4oPdkga
2VdHZBuwBGROJXn43HGDCFQi7OB1li+PtdHkIHKO5Uqez21u8WX52sDUvumH
XU0OAe6goKWLufnvZZZpbnt6f5EZwpns+OK9TXKVgSfpeUGufA3YpZlj8Rnm
FxvKAPdQ5S8gbsquMrP74gJp5l9rbn+ecqsUEV/VoIVanhwDrnGjQF0idf/F
AJNiujXkErOUoq10EyQjoOHC5rcOlecR5TqFF+7rFf83gCZuLo2PN3B/ukaX
lHPbUGyZ1Y3Vatr8VERMU3im18dlvrt70cDlOxVHMSC3KndxhKDXP7iuEmhY
B4h37lkQkMCkDwr/lMbQaSbTwyssL4Nc9V03c9XY7FE7Ay578uVa8JJU12S1
fTe/KBlzdc86TACAOFY54GRun3MGVa8+sVNn2Mf374fPf3QnwUz1E+nUeTyl
aAMbdgBo1gg6EeQrWkm74u56nzOhDzVREQOv/gdCwwSs70RZNvKkQMSq+lCZ
klCtJkKDyrCAnZX6+3HW+lv8PK44jF3uqrd3S8Gal1N5p9z8owg+178/IJWr
Fo3Gf5gxwdw6ewk8rI/eiRPy9Nh/upARy74O97C6e2LHQmahVEPd9Oe0Dzgr
Ba1koiRvX4QqEkBTys6L+Hn+fE+hkljVBWJniXm1/5vSs36aG/mUAiSq7iHQ
JRlVd7vy+NZMnu3VaNiU1Fq42iNkffC/+rBk2XBCBgMTYmd4Apiw6a849gsP
qir8MGvcZ/bIP1kSXtLaKyWLiLyyQgf6g2GleMMfK+ERHdLJdMdMpvfMyW5M
anxT174BdICLVlWXKgb3pT4j7eE3ogjHwxj+WHRi63pmk87o5aL7y0WIP8wq
fe5EAEu75ZtwsFV26S8w1gzIPHPZj/l1/2B9K7WL5X3UqnmqxvQP3YRFW01u
x7t9qH/c2RKpcmVi6J+zeh6DHgBteqC7dU8YQp3f/uXSU0Z611e4R/3aQUi/
ZzMb/ySCccHdSpl3y6guF6kSoGNNv62ACpFflBy3vB1IY7ouXbV9BoGLU6sG
dLFBVIMnzLuWMXcUeaukZq0MbcKxt4skqB/NONeSk2x69K/XMJqH4iGFMvZn
xDIbGFMDuQavkVO0SVsPadu0sqAcSY911P0N6/oXg+lkukrAh9NlpsW9PYdY
CUbzqDadF/OfpEyP2lcIKGQfUOHPzoTJkV3/ad44UF0ebRpeW8NzRiac/Yow
UgsygiYPULpG/QB08lp74Y/h3NH4V9fHTPCBpPWC4ot2sj/NGag0vWgluL/Z
eM8KyJQbTy9nwn0cl6KabKBAtjRmfF/QhYpHCIoDHS23sWUCmbwqgLAfjPZW
b5KbC61/XbeOtb6X7WJO3QpvOIVgSMN7qv8+ZX8Bl7iGTDKD2zvUw1zHxUOh
iMxbhx/b8R2RTocMJygB7FVsgQkacAm8DiW9SJcPSA9F7nFyonyg7/ZItYYy
ok0Y5CNzrc4i9opfbuenusw56X0mLui+WGT2i2hkUATSKANd3sEujuHRkFAh
WrgzHYCroH84LsPxLxIzCX1sQUxOpiBxjp+kwQE98/dgRrViga1sJI9V0buw
boWeL5VFJgXQjyEYAVMGS+IhU/DXyQNU+yxSTXE6OTRjl2j2ae97H/MTQFKh
x3NzO4Gzj2zgeGLQsHkYN3RfpwkHF9+hBWI6aF7rJkrtQT2X1l/mZKDMXpwW
ctbuhhR3XDIAHRFT0a66M0f4S8WSZH3nmbITnA/qbf49WSKFS7oO/cSqhnpI
NxW42ylShqG/ZxmoJsMAJSVdP+3dBT3jrIRUquY/2L6vDaoiUXwkFntDOY7R
UxSqvqdSnI6TcRduZYsALAbVmAgPd8ZImzMPvY77xKAYAsyJYF7/TmOZjZUt
rwTc3dj0qw6c/qFKGtxDZ3PzaTijb+OfWXP6iLHGIpxreOR1YnrrMwrGub8E
zYyXN/Qvlz7wfn5tml5/fG9/DSByJwVP7rj7ko9He4tw4MwmAjM1vwZ27VIq
uq4UN6a7CVqLwnOonMS8lXuhUZPss++ZIGc+Grd2DYyjXnmqVCRyAtkAe87G
iI6SRL/BqUiuGDi+PXYg/H8Ug95hw4VHOdpAx3/ce4lsRpLTd/YdimrEfAOP
PI2P3W1h3XlCBWmJ4wzoeiKpZ0/70+rvdp2x+kZMYkk9sSm1hNja9BU7Yj5b
h2Oeppk1IzggzbHgspxEVCd9cDrCHFUooP+x/I7smZQHRozlhWUYZ2qjO6LL
kJKtvtUAoHzOhfeUhyRHD24xqmkIQytgPWHpYmgubX2EIAgQgRVRlRaYTMmw
66yOJNsW8NbtJ8S1DY0w4BcrGg06d1WJV+2Vo7O+IRpKEAPNE/U20NdB18r0
CgON/dBSrBgaKgN9sS6izDL75AB2bKtcUKxrWBmHtasb1jn4edBGTepHUHA0
YdETcAa+4MbRbvtP4OfH/V4QtF+ec4JLqXExOkCh0tV65TsOwJj9kJYFRz+X
FkKNLa2H4ko/1AiXXodG9aocbcloFKRy89vj6TElhKvpLHAjl6VmIueXhr8S
+VY5NZBVttLCw/vYHSkyCR4gn47wsWvtliJj02OZrIov06ZVlvBnGULOmOIz
Id6IBuNK4+QNixnZRObDAOpMtc2jXhKseY2eOGDpkqFKfluDzSzws3w2cj+9
jElOzATjXimjE2HXOOJnPHNXb8w3rTHZnX/QAQwHPQWEJe6mmnq9EzVV5YLz
3ra6mjBp5wyzXlUOHUjPWmWAf5O4rn3H2WOGzK0cdTb7WGtTzME5zVEf+97T
W+yTs+e+KoWdb6/pKCV+eYLW0KvTvArGHJmdQ3lzp8lBc9WqxLnMB8xbkxbG
whdQsQpoQH66uZ0hYLie/AZH5PaKzRjQl2qMArlw/iyPk+D0GkYfsxA/8RUh
yBdYjjDD+dZXdWuMVPGhuYThWfrWUMPnre+aNakocQHsi2woPsUK+XOj8E5k
mxVcFyNBqW/q0xHvclJiT+2eujhyEBeWL3THvX9OoNavZP1XQDWxjb/Us4Zg
vXf6l4S/WSZnFT8K+e+hX1ZRIlPqePueVUiFyn0hJFFVqQ74Sb6hF7kV3xgS
KZCFIyCF+fZT44t5YzpYe6X2kLCltQfKLNyynICb8exI9WrHLCeH2Z1CJwMj
vvaB6wLdwY/xHb8ogrks1Zuh+1p1gnmrKAFjZbQiB+P9zA88QpDcn1plhdTP
qmNk3WkcxNR5kflZZbydEk7Q569KltE++tJ+DD+V2EaT/WiL/SBwMDXi+OAY
00bX30PoIO6xN8WbGuKPZMjCMOu+jvd1paIrHlnhUJZIu/GKex4RV9xdE+Im
pdwzS00SBm3s7rl3oQwX62x5Ee/HSs7kNyXV+yemb9TLN0noBbUPwzD9K45v
IFgePYUHEPEs1USb8TmHgSLPpQ55mgGe/AIY15oTu0MXqs1UF357cUJf0aM/
iUP4QftgpXP3atgiAmT5Miwae87w84H4EAqgoglC5/sNFJRqah4wkNM/3ZmO
tjnbvPGzLHgXjlNEiSL3R7M9XI0ZgHsw1vb4rDQY0W+pe4pQ/hw4EiGEpqyT
fpcwN2CPdtcyBoQvxEMn100wakcwdQZkdTgPhOK8VSgkiWKyrYMeqjQk7MDC
hzQDtvCQnSZeLwPUADafcPE1Xf74SdvIseC9x/CJC09SXbLkBGlg+k/PtL3m
2U2d0fW2lkfeZtqAl6KfThqeexLIK62l4SFTOCFPKy5XsCUEM3ixl9whzHUh
VKOTE3eusqV19s7ws4Ofy2yOqQm6xXFoggT7OkIM0TK5j3srvUAYVXgdfTKg
AOclZw6BAr2Xs7lbo1GOwDF+XuShhXWBNfb9lo1/lXYTqJwxn96BM1kuvC+p
SDdLFqOMFQjZA5rHV5ixq2N/uIYSA675hVXjDfwgunFnquzbjl4Rj+YdHxCl
sis5lO9h/AED+JTSaa6/BItv8CkCNHkFuKmaEmQZ5M7rO/yPWz/8BDcRxmeO
oN3x/9/hLc+q9tT+5E9DkFDCEotqWwsUtNhlqpzEGrW2LSj0C5hIpqc2NRYg
TE+pv9FfiC4lTrJyFjjcxKNqcXqMv5DFmsNJA14dlOnb4CfNYRqwMFhozj4T
mOJo7L3/bYFEkxr5KM1S1ADXab70Y+FO1bz63cp+OKGt4t7KUT2W2+CQ+GgG
NTQ4i0s40ogVCTxlO3aYDwQksvD/2Wr8HIuvXomuUXqZIgd0INlHjBHlu31h
QhrQUeSRnNMfAUc2buQHDivveeghiEAVm7y92jk3yrmK86f+oAmJUSX56h9n
fStwjhnNszmiRg8i2n4HpwxMa/m9BIVYWKB2EvERJZSYLrgYuWi84kp2QP2n
rmKufbKtP4SkDdykR9rv+RFP0CeeNDJtPaO82jx5FPcJ8//2Q5zlDGJhv2fB
IzUUKacnN0I+US6aGDPeqS7pLtUlBZtetFCmqhR37N3O1qNCAB7ofzeOML8J
zrH1YK9yZ7uTG3A/C2BT4pwsQ0Zz6iIujlYxK2Xe6FrLxdzJR6+5AuhRbgnZ
UUbiMkZpoLJj42BPU+vTDnTadexuxQPqPoxXFvpmCD6eZdqpXRKadxP4AwYv
a72zti8XQbSCGbVJWd28AII2IqdpVVRzqVEgIi5mSJMWn39WapcAihvS6PkA
yVUxUaEaR9zcsKiU+8uP1Yhw7zB0cwsLgEzisLYqOlWh/PGlbZNjmcltHQzc
PIHnMqa8ZhjQqJEaFB/kuASPVgdmMtuHDml/79+7sy4rCN6hjhCenu/WNBPB
YNe77Hxl72orx4eSmG8jwjoVE6uXecvFUEdBiQsjMX1wVSCLt9b2VrmwiiQT
etytjeEoiDPxMPNE2nvieBKv04exYhBXG+eUQ/FySAdBS57g6HhMgOQEikTu
xxg6uf5MSP10mbnKqijhjw5oRXYXTZrURVm7vx+gB6/wnUBX2TD9ATWdboND
T87e9KzB9EA4cdjoGWhFuPSyTc9KI3GoCohr38jNYUnmNetMGnYnwQn349V8
y5OVIKRzhLC4apr0IhPIor4iu5ADay7YeFimuPhbZnRNUc0KCYNdM6f9galp
4v6/kLJSuZCWqKpdq6vkbhSsrxFs9jimWYx0nj4qLBH2vvohZ11J9yFbDjlN
RMC0DvcXwtYWPkLotpTLv0WPQyqwbrxgYqxRuL1lcLg+hyMQvmQkPm03hvVQ
NN4qe+Aj4WXpbUEyvsDiV29Pl7OrgP4FpKnKe1fJ8KkwirkgiUqjADQ4Ra35
5b4mmvw93WkUf3mPM52QvmZiLKvQVHwJL3Hx+xJQDTMR+MJmReNvU3oV3jYc
Tjc/u3BZx+F35fYGwmA0PdOoBf8YyfGzVB//0q0s7aspaQyG7qxoA5GnfyGH
Nhod520C5ft+UOhSwlGtMS5EGM0RrvbvRpz3+PLMXL4RDYxMJnvQN1GC5LYl
icrwfnAsxpTl1NmsymPT6bYx3boD8VbvTk25g1skECfICvSPTVSuVSGzYaPQ
oECqzcpnLrb+a+EZcQxt2VTECxbTQSSGYgiRj79k6g31yWmmVIDy1rUW/q5R
T7l7xgXcI8hDn2PAy2o6HRNF8CMYZfDZ7HO8Ets6CCKJHcbYHaqm62mqm34S
CMx5yv0oTWQA2RTmA7Q8TljxVQEAVta7HUO3qBzewYkIayUiV+AGRtsH3qMe
LHQaAXZsn+b8BRcuVPtM0cF7t+QdRqQBmEEOd3uWWJC9GoBdXkAtYmXRw1g4
qka9HJsjaIu/l4ufNtJ2DJ/iXxaPXl7zKA6jHtgekTcaUOiHo0jK5SrDvOFo
gasyQZXio9GucMPGKtbfYfwPcoymlMWCHwwqzyg1FfO2MV317ncSj5gBTMCU
cKzTUUvGPaJ1F6OGgYLCKBu2w+cj1OiO6bWs4TWkZw0yRC4/h04IZBOD0z8X
9W9wWFAyXb76Eoco4T8Dl5MlyuIJ+CWR6VPQoEwahbBjNfXfovZxo24eFaZk
mAgGf3g4TqXf3gjbv+DLOsJYgdTPskBa+lYfo8JEKneM3AniqpwA86GSxe1y
vWGnj9I6FHRxuyC6A0ma6Byg1P84d+CUZaUQ7IVr+uYhrYSkexFHxGe7HyXq
uTpDgHhbMgqD6xmwUqqICtnonLAoR7PSXG0bqHu2NASdgGrHbJMTQwybD0dZ
ulHvxzzELwrLjV1pO6vCOcJMUMiipQ+en0xNQwt3GcPwho3pbRLZwAZwC4Yk
e9RR0j6K+kaYFe1F7TS1UANx2fz87gO6kzzAB5SYrk55OSEtKFwfd7lUBhxR
ofvuWBFppp6oEfGBnGPYnuJpTWPTJmOBdJgVFfm8sIPc6hSvL5jad6EzIIrn
fZUZ4rdNOZPnlSXjVYijXZ8fsIKxdu+DMbDxWS9Xp4LBefLNq1jUg07zEObA
WJZ7pLZNm9eSIqg1ckD+iAGgBVx1UkpGgElO7igX5zR/X0Fc2h/4NzohmYCp
Jwc4yt2ZUSbUht2IluAtDB0yFmsQdtG+a7c93MMycYmXi29yH2rfUkTs4cAl
xUt7LeHsZeIMU3SV8Ym1KLMVcFesuRZpY3EXCUkZrjOh0+awhThTnrlLOZFa
X6i3RCkrL3OP8IjpopEHVvWo2x0ee7LDZRxWjj08uTL2Rsj7z7GINL7OhVqU
eIdctZLXFPbx7gBL8fR9/1RORtd8836zgvOBSHlXuIsbk8G5i/TIJq94Zxq9
jQh/YUL+8P4Vrn2FPo6eVGelYp7sQfehfqZ3y7L+uHBJnYt6iCxmxuVUdEBK
ZZsZLfLUxsGBA+f6xQ/8DpkTgWKxDm3kkHNv3BV/zAg1QwU/SqSaQJAbynP7
dSUW0Dx/zsv1xl8MhcOqPLm168MyVAf40p0lRHcLClEr/dywneWcdQbbV08E
9UHcig8nwl8Z/xX29QjRPBxWzPfiAMaEypykkmhEQVtOwqod2le3nE2HWrvN
ZLL6CMrHSp52J31hTALqiQzUq/A7xXXNz3crZWvDNhjOvpZxeN88JmM78LBw
DqmfcXmZUo3w8hN+epVhMa7HfbhNX3YLKg3QJYlcxHdETyCdAP02gKHMsZ6L
VYmMAMYRZgQSbR9xsD9a94ARL1pcC2DSsn9upvENJrUpvahW18e32rHfXPpK
MDccxwPHBo/OxUZbAg14yWcreHM5bOcwsAUmDARNJc+2XkXUCWgDOCpZSibS
tBGzuhi76DWnmzDLstdFFhpaHsW+PvPb+RMGnhDAe34NDLZHJF3DmsMfRpuE
Vw5h07q5iqyvAuEReQcsh0/FIhaMsBAMSH9RiMHVmFc9lfjZbS4tVTP2JwPi
lAYbkpd27EPeBQzxTGoB2C2dQtqCMru8X9l2H3lG9pjZj+Ja9i/hvA+HON7J
L5ggpe2fi4ay1OJ/Cli8u0KVsvDMa3nwEI1lnXyIR5/ldf68bgv7FgD/RLGs
C0e1yg/WA/SF/9vXqTYiefBUpLiY6Wny7XRD+Vu31y/8Wc32OTSbZn+9Z46H
wdsGfw9nA7XI75soPbEaI99IthoSx4Tz+/azInNti6M2ijyGnFMfcW+WBi7k
Abv8KKljo4uhRB0bGvQJAwHmG1xufBu8oE8UeRHxdNIm0nzLdKDXoKLkC3Ea
wJjtsxXkkVp17wRneLzk+C0//RM+GetXWPi8U6CR4Zo4FJwlHXrtFYqmPgID
12nI2m0nHIrX5ab51UXZK+WvHt4G9KprEkamR4POXjUzjhnFgmjf1/yrAPSC
GyjXaEcr63FIxKHYmK15hXjZcdh/uvhHvExkC2OJDUrw1NOEaIzLaP5VYIIu
H3SIejusEdEFJoLrcN4JEDzAt1jjG8KM475lRz5abnzaMY/dwNKD5LSgnYCz
1LHlFZAmbcXG9W9l0wrPb5zwKLjVVz51ZBvtLI0VRG3zMtUA6JmXelm/Saeo
lDawPEgegab056wj0we0GOuAbPLssj6FAHmonrxDw7xWWINNx2pAJguUPw3z
G225TB4Ge3wMl78Pyjq07yYvkxe2SpYzBnNtW29akNdcW+2VcxVmZtDbXIH5
FRicmL4bfrxafuHo/Zfk414Sr/qwKDqJCFHHpNmsfDqPJkHcz4bAa9NPIACz
UIzL9eSU5ct/OisT2+90F45U81JBJQKVBtt2KXlkfgPnWcI/EDum1Mm0iOtt
PcSP6NW7gnASjde2tnf7QYDcBsgl+HkWnFpB40POKGb7w6CshgGdzuIoWQKD
9KAxqbTZqnZS0mmCT3TlVthH8czpziIhaOi/iRiNb3/CyfGDsNFowOHbVpf4
Bjm6xPpV7VZXi4kxL0CNO6zrma2iVOaRwADNcSjy2szUI+ida6wP8XIUwU6J
aRcp0IxiQWfkMksNNiHn6va7xYTQkH51PPBBPDqhmZDDydJF4HwhsrowDRXB
N7eroCPkaTz762NBirC1svP+rzUI9bCithSZEB/c4Z0AsE70kjTZy0aRXGCc
G2Vkga5QNhqSk09IIHEEWYF0KNS2IQ/TreE65frjSZeJGZAcvyLO+iH/wXsj
jykEGxvAxxixmU7NCj9k8f4rKI4nFMFeewy2h+X54zSItfFK9nc+dwdROQ2N
aq/BML0ys/lAVYSyN6aWV+SRuAq5HAeHKmt13YridMMV7tyGA5MBeA2bsLlQ
xva8CDyX3UeDwF4l+YblSk8NSG7RaJXivMzDZvdFAjiKsvYZ2a2driD74xOk
VRScxfXHAhkJPi2l9jvFkaiDuUvaQHXp6W6MSlbAcnuNS+k4DfUaMNtMGTz8
q8Vh8TGzHM1qdY/G2z+89Dn0t3sbo3T94zQugWJjCq13JdO5adLTDDWHmFQY
MHQ3SGdfvFM6ayknxjZTpq5O3c0letW1Wjj7PHXytZ4KyTvdC9zIcS3klFZx
4ZQx7RCUy6Etjo/osYVQQ+OhGpH5UrJxpy/3m5Usk8cVoBgKCPweqra5RE/O
tJZ4a9VgvRKPjFADGzmnRvYxMhGpJBaX8/P1QTrn+BVH8tnbd7G7mDSbgck+
r6pdcmpO9pmfE+fjNTI86U12Fj2msnQNmM5mtTZOyWUve5nHgz/RDquQ3Xt3
FlsSoG79N4Ghe/t74RCYhyP7AT1XtSv2Hz++ze6fKPOQu6vJq+GhjfFXVJCH
3NOBTwY9KD5lIWN2ki2cPuHDznIP7zxpGZqFlMHPV5E3ZOQIcjtX3y8Ytsq8
wDnPAU126M3TPAoH6SF62ih6RJAOo9EZpQgQIWMVFKCOOk2qN4dg90JhVns5
4kDcYvgmliJWw0kPGA57ezeVQQEBOMfF8u6VbIM2ne417NigMChdPlxZcETW
333JII9eznzdyFxvoqnJklEOrn9uhcr1T2O8rpYA9bP7o72SkAsHbHi5G6Ny
I63ryA1W088fpJ5ya5dYmZZFZcgxYxamacDAt+j8BY1sbqhC3FlPA5L7XAqH
DSsuigybwXzPesM4+ntnm1kpeKYo0Z6Ps1HQ1hVgapG4CnB+VEllsWD96Zhq
wtayYpE2lmRWfCqVYGOsmaHq8o/fJPEYWMjif8t3qE7uqnGjyrwq0HiCVFf+
rLKHTyQle20UfQt7liG5K0nSX41VL5V7lhZ3+9pTreT8IK3lv3jhrubpaWp9
xOYQFdn3kgYEtBBkdYFPiJB6OD8Bn56AokO3F6iVIH0iMQyl2KAoBFK2X7TJ
be8OI2eE7KIqimrJKJ3cwZcO2fjq3ygOHdTGsanWKya/xKh0PuX72jGFCNA4
GsmzTTtiXCtwhuRpaTYwxWRNsl8MqF3XYXa8sOeaDcZU6w3swfLiQ4y0TUSA
6v2kvqBdbirBHwrCgr1CWepJa+ta9BK1XnNGRMMJOz5NDubuh+Tow8fMvZlz
immoDI9MPhJ8eePZIN5N/Aa1hPcwZzFuxa1+ZTl8KnY4MmRBADhZ1hU89XIU
KtOvsEJFYbsLg9gIzHiAKdjZse700sgy3TBL5H104utpt37T6ctvkXrFgs1t
tc5xg95aArJQ4luMQEV5UrPPnxrUp19cldYQ1U1LlMcuJOrrhoofHdYdz6oy
13O36x+YfLrMlXFF90xaJRP8/Aa/5brL8zhEdqPuhbLzUlMhn/8h4bZzK3cb
n0mi8KXuc/gnTUq/+ff2NCwy+VrTnRKPXRD8Vrs79HglZzBOXgquVog7jqaM
cMqsIpJKGmgd+xn2t/IO7OBE9dWmZfRt0FKEb1Rm2EwymS+9r/HjSPQkR9Ap
YpY/olKwfXUo+yIv28qnBZ9L6INZbL4EqiYEWIAY4urStRwwYyQ1zkcD6QTZ
M0m6qVvfQYGEAhOnur4Nw3QB9twsf8Qn6y3eTsmWDuai47dH/P5xgGfaK4fW
4mhaB9VFPIPZZNlWhSc5HkJfqhQAS+qTfV8iZiJa1iCtCQnLi4mehIo7XT8I
6Mtzj7TRL/e4DZHomqcAL2Avel2MGam99JBBnXKSuWWSeyohUfbHAinWyj91
FxfxNi5FDOD89JlBtS1ptan+XpA1peVSCN4Anq9Tnn/vLSw2GeTVAgGefp2K
5SylHgwCNKaWZ/M8J9pVdyRyt16oecOmNQ82sNYzuqQNvSJjD3Mtm+OLUJZs
XLLiKWddc+2xTSideQNrFemkK0IqDAUc8EBpNU5BYtuVQ/M902YHJdoYvfOb
oLBwKmEqQYYMl0E3bArInQ9XEkLJVZyFRUwxyk0wqYD4qU3WcpniIxN8ovPU
axv3QouYjbPCssiXVPxbdrKyQuVa/mYoCYePxUKh7zmObcpJJrnPiuigfhLI
qgDx7gyhsdNJH5QL+btfxYxm/xE6JnCNNO93+VVGNVQq/oA+ZVIypnZ7l94B
RQi2C65YSnkYp3ywSD8yYrz4ssYQ/GygjkJ9w/0bLOgXuBGX83NrYL7WM+zj
Z27gYXoiDSz7ECUWNQOSSGThaVPRzEnlAB7Icjm3uK3Q1Y9MAfN99Uq0/pqB
e5UfGYFII7jm7xefuaS7CDDrx/t7Ujr/sgvVEBEEHvHDmT6t9T5PSShbeGmK
UZneRbKrcmz70LCVgzskDxRgm/GCC9D+8pphgnDvkH+KW6b52gCwCpkW2OdS
8PqgaVbiT3ic6U8esnEW7vIAjWqyhDOnQSzRoyZOy1qD0ipz/D3f6k/WMoLg
SIrXm3zfFSzUjckqJkfU00DRup+Uri/boeThAOFf+WEQubAbZsrmiqVm2FRQ
1R38dWxBHeMbVIJI8sa+ASrWBlfAfjXLsnmfnqKrZTZovlw0pRixGF9fIOgt
LHtkJzEbxvl18PYKpfYW445AZaXRzeVR2z2lxbUaPS5dMQTfA/pDYjOA0BNa
9XrFNbG5lu0Xz3A5migdF9bBSy3FLf3x5iZnw9TMZLN6ZNWO2JD7nn8tfAn9
cBt6U4JNs78lSIsQuoRg723yotIa+95d/bB/okursmwTGFVvNzYC+NV2K8DF
oF3dKxiogHAvKuj+s8r7KPtn3SGkZqfHUBBsH9OMfUykXoWE2fEyuBaBY133
CuYHEzH0pWkWY8AOWsAAprnz3kUsjQ3+9p7KKMaEuXpJLnUipaCQx1+Y7ZDT
yRChOUsOvHnR3788y+Z7qP0VbrytKuUn7oR4MzBhsNk6a1K1f0nlGZBVKHo5
oljo+byqOzrprVR1e8I7x8yfm6GlnDLGEq6UEiJaHaa9v6WrUxN4d1G7sXsW
2ouU0hENB8tafcAWDu2u2fYoEUEB7DtP+zh4oWy5KcVNIbuvQrozmN9w523R
yTi7R68it8WCR1zzGGq6zYHNPDS1/hwCchbIakhf/6DmsbP3XDBnOolVIwGS
Y/3dRI5xDk0fSKks2MC2cW/4DFRNAtGstEvNs82syHYxPA4Zz/whT9dwFeUq
mwibNcTbd4X+OJ51+dhjqg694GK67/OWtzYjev+V2ebx6UzWJNey6htz5UXz
1XXIF7uTL2ag1zcI30HWds+zzFklLlIIrRvuhSq51z3PhG1pvZeOSm2zWfiu
6LlhMFHYx97Of8lcxMyPRcQTAhdMP0l6twCp24QEiN9LCAjcp27GPyNhIyzM
VSDeuL2jho9XdvCvgEO+NG1w+JSXWLYFkOcwBLP6pMeJVe9hrLz2Lws3aPbH
ffec+pNnEGD/3mRikhpgq+fRI8Z5tnbu96s+IX6eFq682EDVYKtF2AhU5ZeF
nh6hya61uwlRTX+2jZepZd6U33UK4WpI484VvRXelcGXYy6Vjz3a3KMGK3zB
3a8p7QiekjPhcYEifHfLRmofR5f9l/BTjXR29//RU81ws8YxICdpRdkvHGsL
nNjW/FGxvZowBZYjxDDlwFnkxtF0R2hNDVmGEhmJtOe9QlBNzkNeIQ721+AE
t0L50pm4M9ntfw+7Tv4DV2KeuRvThQ4oy8BmlUKW4riQBhJ0PrEZ/5UsC4gg
KdD2BV/pR+SJCIXOB/tGcrMqvAvUBXNRzTcB1y2i8QVseko6Ut8t3GDycCE6
MvLPfVce9KCEdzo7Y5L07sVsq6iO86UFQPylV02WAzGunQK8Vk6715kLzUNk
GGZ0v4esjEoi4iR1R333n2B31nLQH/XfsPvGgcZhNA5vVQE3YUKNPdgAmse6
wMHlsC3jOjLvUDKp4Rie2wSxHGcLmHlHonF9S7aSTkqva0kfxOMBpnoBujab
JfDNAhrcrQeRLZq4u8l7fcFOstfAJvDEzzSrp5Ic2WkdNOOlUaRPWl1Uwg8U
aPSFobrdfO1Du9yDZyXIBau/L1qev6eVHQN0p6DgdZIcK6n5XSaranRf9QU/
xtmmzXtZMl7D63FPMCJd2Npgmq6YEJfphNmY871sRJPml2TrI2eGbdOvEZCf
YQoUp0tYxEBXHHTQAKx+vk4PhURfCdcdgPT1sTaggTfwtiW361WoDgirE1hz
13Y3TWbtU6qGKl6eP2DtiT5WoTUZQFLMDrA8PKyX1sQ5JEkyvUW4+lmtS6X7
o2ysnqeS8bQQAEc8kcrN+juj6s92PqPul43u2vV36zQQ1jy5B8OvZAyNK88U
BipN7sxhtr8gVtgo8T4o/82aW3/rvvuFQ4UTmeDbAX5jw4pVGabBpS3x09qn
qjMqT5qNwF1G/5DWKLTyX71nwiH5ag/5D1OjxJ2KOezi71d2UexFlKI9VFA4
U5fGIqSrWLKCTHg13w6Gk15Jox9rnHcsWhRxD1GtR/wGFhd/i9eTRGUeBAdr
ySKkmdY31l1AN/h30f3C3vBjm6tNRI3i4nfmtfTSPWNVH6HZDTP3FLfdPcFD
kafudI+vFtrLUoyr/mUNUipi/HKB2KMiaScy5ICtY1Yj62KiAByTOrZa04ys
H3Gr8KuJOJ8L52I2pw+8I8inh6nmgnfasxa8nkBlSuaMKupEi/K5BLNmmKi0
ZqhXTv48nC8StnO0mg1loDIiGarrAhXZVoLPp4qoB7xgsvwj5zRDtg9IX+Mk
7su+lR2mX+YkdUbXeu1FGX3U1R97FzNnFzE/WjN5LMGbSUJZUgBuIHtWQko8
RY0qP4xPPqXmRPwG0eVHjWFQqBX60IrV09gltLTOuC7QoSfRe7m/TQQej8j9
zGT7/DLt7AC0jjU5ziZNkAR/382C03ThSFUnpFgseK9PlKWsS1QNZ82VoxNh
YuzzpOAN4TCKyO3f+QSQa2rKei4IMTNTYIUSJA2qEX5rkmJVtpCEgWEf56r4
qEnT3Q9Ozrk3SBVREtm2wFbSTaosGW5XX6sKgSKn3+Ocsy2C/7mtl3oYDaEB
+Ldmungxrra9wdeNPznpGPZiaASZZjbTRzDHAsaMIc/l20Y6KaIsD5UFVSMq
3p9u/HvzgNWaHZGzz7bRyey/kS9oirPtJjiys8D9qZ67BKn9uwEb1sO8GVQJ
gMeDmBXqjy6kqdCIs467OgrSXIQHXRcnENFf9GeAl1JOMGSrhdEMNzgvJwEu
fG9+F9LHioZpQXY79a9aUmHzjDC24lYe9jyHtfM7PkCmQxOw8/csZbu3cjMH
5dP3FvTX/Pfr65ehf2McyHSbp0p7/ZDR0H1xDmcGhnTxIhGYFvD//YWh7ETl
xNrNyemYY/FStdtVZkZOFp3ER6oNc2tUlyiTwv6iUkRsBZag7JbJYbnR1tt2
+Vv1i2K9gCXTV67Ugjcy9yAUBMHZYQZcYOsUhvqvXByzc0ayScWyAze5Av3A
lKhrSOXDu1G1OJIIuhhGciMCovE5L4QCwnLkKbRXncB3wg9hi197DkWdNKNn
x7NiFZAL1N3nZAK/gUXBMNpqZR1p1SP8ic8DMnXH+Y8RfwicOAQIiuO3JqZz
IBBfZyLBUMsysX1SFm7pKaoH349xyj+qCU0ft/PwUvSZ7ccdFzj/YNZdQWlE
4vhWpicLtMH0OJiR73/hDexYpeBCI12zLEHo268M2UnGX9BrZMtElZx45aTR
VDErEIBF/nbFS/aW8Bvlxw2MstLOI3n+9C4MvCMxmHZtnyDHM5hnUJgjylsu
rxqzFUasK6YY1S3aRUdi5yd2iPUwtpBBxn7xiAwfdMyTL+A5bAlS1azkJyb1
sdezPRHvJ4ZyLkvoAUMlEbuLm/2k1Xfu1Vrw5fC5zRzU9boi8Z2MPcZxtj7h
470t9K5jnX2E3lJWAgf/QiDx09ahtew8nSpuEiHQ0aGMRkEwBU4sJ4QuBLPJ
Cf8JmPxyh7ZY6pmnhsnZPlgRd7qkQLyZRSL0xmO8VsGlieMGKKtAM2EWH+88
uzx7CAN8/IrWCYKz01itTN56OPDIwcVccvrf1A/NUkgeWkDDD1li7kmollEi
2eUbIMgQi/j7FtbXM4E9vjlOhLdqvsXW1ihzhfldBq/td/kt2wl2F3QJ2acI
mIewJOkbEivPhWJnmmbVoigVS8i/e/vn28so6JVipim/gtBiz0FV/5Oh0U5N
i496TD1dZ/1VZLzs2uN/yV9auySWThytpnytBuBpB4WpjrOBPEIC/QYTRsNV
0MapmnMEoz/mkdGjsG1txNmCiVB6Cug/qRQgtNjp1SGgRhMuUCbfxkW8z1Cd
Fv3S3cEAiHro5icfbMHm92L7CvtsKwUVeZ7Btro4Dhw/6kQGQ++RUiJjUnPN
JBp2AveKVtMetqoU1FFWmL4JmTQFpyJ4xIwDNL802zuga7YsQIYagOfPLJV/
G7kaIcTdBSgIWdm2JffBLsFvFImmWM0T90cE1djqsEIIIJA0th8t+wNCa6Ph
grcxIUZJGQI4fS2atDHkgyndwfx5FeNQj19nKqiqA9BFF0AqTPnI7b7Zl1XA
NhsiGwfy/1PDFBDguaTEo0scLTlIffiIG9MyfxqyMYe+ipv5jV1VFF2BcQNy
dFLZISxtdOE7BJK56Mxgys2hSbRlVg262/YGdXySTLA/TLlhMoujdy/E14ye
YPOgOzyZlUymwJ9MKFXcA7KyftFAmN659vwkTzpi943jSJ029FZS7SU3GlwK
gbFLgc71xvTCjZY4usv8zx+mz0V2kE5k8yBKMwP1V2qSzEpDXogouKTgcNZr
5UqMpUSs99rmmH1LHDP2mhVJErl5NUQlQS1pVMdTiTtuvvEuPcpnPuw1yY+A
LcgwrR5F05dShnScRvp8ifI9OulUvV4mamQE44f9PtdxTiefEKwSJvnJk36K
QIq1+b5ylcZc6AoAqQf9UXtn7waADvTvNvH7fsqNgMa/AjkTuGohxRKLM3B9
CDaOzAFQp9KDVuQ7MVeSRBzFNCg3bbHZydCymzsLO1UJBmDloyIWJrGnJoDk
qIWw8PGax+rguZ1SN0W0WR+HDtyd389+jjFFUvbfq+dMIf/TMxKJYNZI4e5H
BG1H5Au/xL+dqsgpU7o/6k02yaeAmVR2Kec2EKPQsMlrzCic4MhwvANL6UIt
cpsDQDE7dPOTxpCiXA9kGxoZvjLdKGmX4szH/GUbQMsdmVTPaDUS+b3dsSeZ
CGXNsCqlMmFMZyVeRxxeCErBCT9glHfv96dSg2iT16w9eVkZGd2/ZDD74jis
JLbfmOlaVmRZI9JMGw9L4nXVMdzquS5445Vd0Lt23Ov4xtEOa6wLzO5+AEQZ
ArXktbCT4hX88TAEPBfVF9Z1OmM6lJ08H+e8MRA2EV+PD9Ne09E2FA10qvoH
LVS9bJFl5VYHdQVMUsNswZkhF4O5UOdMMBK6PdBQCvl0bZR0WScDkzJEaRxk
2s5UuwaXESObyCeKfw43OCaoQvPnfZs4OQ5RIihqWXuvvjzHTXOnAibMsw6V
2RsiMaVn4d+kCn8qlz2l0lM70GTTG3eeA1+MDiE4aCf9A5Lyvt2ZyAw4dpy6
iS+RX028vZjVi2tX7kIis6rexSLdc4TEaNq0z5h3J8W2Wkna6z2YIfh07UI2
O8j7Zkp9lQVR5rPVW23l3aj+HG6q8HIlZDpO4gghT8osDuXaKLPcDRco878z
tdOaq1ifUCDKThMGjtJ0oS1sS7xdwsz5FafvgFD5joU74Nnj5uVkV2fW15E4
Pq/uGtQKmgHpKx2vo82uCbC2jBn0DxZ3NGGZY2TWyEjEySUM735/1LyU14fi
EvKbqw7oIjf33v8eL9QQlC2YFtitJJgf28kQk6ajZTOxcpmaK3e432JRbC1m
2WLBKh7dysZX5VsbXVgqF23pnCawziF3qzW5zzm5LgIdOyaN1WSpONWxNPe4
jnkyZkXeriEwF9VJuO4rdytH+6f99tsR9QzYs52uy1DdQNjaGLBeeoqCiAPo
077dcpf3Iedg8uhi08WvlQdS3CcMXHvLElcXNIe+OOpi9KCLi902q+YpN21T
CyRut2u6aFIgFmHf03VWPrk69yIrWNb98T4yZNCyHPFc44SVDgunZvLcfigo
MfUQtVbbbHgd9KN0HuhnEd94JOsMUcSiX5qwzZsO+A5SWippXGkupcFEQPvz
wB7BebqLoYgI2IuGSVzXAJSBKBAgZ7q+5HC6WC9fWOsXMkw6PrF3FBHpSZ/L
nuFOnwuHkvXE43+k7feVdFnjPSECGhUMt7j1CA2IsgSGgq3f/7+AsIQ5NqfD
7qd9HQBEGvNZt/dQNBVd1++gr218s4B0IuoiCN5Bgg9Z8Jzcf3r7hXJ7HpUj
iPok8JMiPwkP9rKSkYDBTISfrnTZ5saAT7DPwTmq6hISMoHGgQ9Q7k8Z3prV
vxK5SHOhDLRBbUPMcXahwY/aHMII5bVh7V+NlFMPjroTFZKcxRrbfCaVU4o0
/lV6ZqE60UOP5C0FmU7icsba5BGnQsT4+s1ZrTgWClJ6oMUGi55dpjg8GjoD
MwkkiLtNJjp/XL+ZCRP5A93YXIIuDNrKAipwULgdoZewdb4vAUdSdoHijYOK
S4Sy1H1/b+WAkCGOtPREbZKt+OPQ54y520MYKFxjAxSLN404M8AsdegBFI3z
7SqfRJeNcsbfWZNq66QhW1rXB0CjqIIjRLTVwpWV+lpGnOcCPPTrB7mq5IAW
U44pbTc+DY9tCSGl+P/BDqAajEWt+oPawSuHtT4C5Yf1OUMlotx7nDGKFT3z
UXqRk055sDMxEyntGj4yUQbBbzRPtJbAApCwEssDLjl7fK2/zBODExgp2SZq
s3zjA6PuPrccKWGgbo+LOjM2ciXJCtIWN1ZQmyqr5MSKoTHepEyDmt7R6bQs
YHeGa/CM+UKXOgw1+kJGJF8ePRY1OymCo12un2AyDTQRZ0GrOvxOfTxaoAul
URpV5rOOye5yqxvZsImlvyhcKAuEpZG7jCZb8FWTJBfV451jkD7sryuM+4aW
SkaU6HUk1OFyEnyE6xW15ANTnD3JrX+QsVLoMsJR1zK8EPurn5H9T7jZo7KC
GOshMs1wAd9xVW2IPQZ34zc2xbGZThXaVEp0D1e5cK5cwV3lJmfg4HgZI7WC
usHc66hIXd2iy7btNxuRlwj9fJ/wbv3l9gSHYMqPIrYkJnxRcf11BFr7TvDw
RBMtqPVqlhTFjXEImuQWBzriospI9OMewf7tG1EOo9t2o4iSA8ccnoCM3VJZ
3XsKMGMaXKhJdB1PsrVz2ibvyKqIZvrPMzesm5GX6MhJ1tg1tUCC3Bs6gSfs
WgWA7Sxo7xEwIyXmwvihn7eYlqfySrzDKylUtwQorhxS4NSo4A9a+YV9TwvB
Va4mDwPRQSgb1ZStaXBkvNLBOf8ekNcQdE18e7k4znbIIMIfz7iNFIfuEq+6
bLZhq6BoHpMP405WuSPxv7oZvddcpgGSYBczO7EUSdUO7oca8VDeTY2AZ3Xi
t4I/zNflm2IvPvxG+fcs/yckTp04HhEypfXtaDqAcdLy3jhnPPg87VuhE9en
NkvTMSO115pkeafHvAZKy9+5FsTUxech9dT6w35gL2Sg+B68Fya4SjVm5Xhy
dC0/wWeQYjgNV4SZM0ZAj/Ks9Ox0bsLPjZgePjx40Py3lGC3fft5HGlYZJyS
aWO2uAjW3LRBpSFN/cOcwWDzAQgyOCjVxOjl86HrDkdnteqGPh4DeAHosPrU
GhWwzcpTtQio7psiD/lpNwbIL4y1gzw52ACTvecBopWVtnl/DGzNU9j6JNO6
ALSb46gG7fmbzs/owwVOA7annOdi+D8DVnarCv6HH69dGocTk6Ui60SjKJtu
mbz2ykegGAbQxqRGORXDZSrTPDAp/EDTU9DZZuYH7zcoH4HbMbF/BWPCTkRB
QYqiezpbBR0cMWzFHJ5x5FjjaXBwJObUnXe+D2NOGmZ2F2gLWbEUfNdrK7Bw
bvCnZwd2/q2Riv7KVQUfSc6pjRGaJKp/80waum+p5EY7g7knj9NvEoG0Rv2A
MP88oZybnvbDKnFEnE7RLe1nqOJKBPF1aNjJ6HsbIRqlSbjkd+MRin6SnTuX
d0SxXydwFI4bORjdew38P5kdchU6kdCkaZOfmbbIj7kAhf4yvVsfIBvkjesA
e+bWrc/N/41XF16Cg79QJrVowpBnS+Sc4mOkRalxFQukZNt7Y7RsVQT9Pp8K
kmHD+jVJn/JHvyK0mB+2cTkxOW+Uffa72Gn5qcXsn95UwKY2RrJdKzMvPJ0K
Y6L6qwogbJkomILbwt+N0TuOnW/jYFlAFkwxjBc1XBXxKftxGTlhar01pI15
YUyj3H9IJut5+sMCuSIT/Uj7bzr+um135mC7zGJ+odXhPC3mvkNevFaNZ3bx
jMpPnZwxv6udtfb+cgNSnak2vLyukLHWcENNLo5d9SA7qYA0CHCNYLtgAnXU
ojQG2CwEi7IRlgeYWhPVoXKKXZWiwkGIGoOW0KjTrEPhKZL2ZDQG42k5HB2B
SxMLVo1wlBmqyV6wpVNpaXcbsch20eADCAYKP8Md3CG5mlZW6la07oPfMV8/
t/pdk3f1v6KhQE3NAYuakN6CMXfTTZ54fp8eUxL2rPgUPAcO+k6U4+Dq/qne
CEZENYS4lGV8mVjivL4Rt9lTFoI+f9wse8WYxsuUa6/V6q5Yv4HYurow3BO6
CNH3c9I62KX7wIjthiax7/o9Y7GBg9yyFVudaOnvJf1YRet5nRfFgeipoXXz
+Ppoq4b9ywl+H941JpaPqGLuEqgsXJVka+90ku/1hm0I+csVsAvvz08XAGLI
XbccsqXZQGciiAUoD223tzqs3ldmyT6ODW3Glupcjq15g3C8OOQQtY7uCOFB
p9pY2ige5/haIf08+Llo5HBe/pCE6G6lWoZc2efVIli6khioKHzEuRNURXuX
cCc3gID8HYDWw9t97lg7lN41OMs7eOGwW2NW6khUMOqUlmN5Iw5eNa9iBYy/
WDY+HsAy/NOGXcKIVp9LQpjb4k1+VaAxIXzICr5v+/XtkbB+mojB7OZp8lMo
xE3DCBCcqHenBr4zmcANzRxPcKzR24xrPO7FedBeL50IhvzFPtszKNdVogW5
SA2VudgiWQhRAAr/l3kEY6xOOyjQjqOLaA8H/30yN4HkB3Lmwgc/9I70xWWC
5HjYPu9LIp4Sb7XLt2pwgSO61btT42jO8yyzAJQvCBO6jgl9nYCJAJHpkRkM
qF3q6CtfYhtLbamjJvQ6iMZ2gYeB8T7nD5bRCCoPY4xwRtsZyvbGDXvjT9gP
5ooyfGBEkVAvBY7IAOHk7Abqv4iU8wpLbHfK7jsNRXmGjj0tHj8zM0hluUva
E0HBwn+NZc0UdAtShjpkGQJgx8i9kHtcurGth3rZe3/mOsn9IwunCFVSA7qa
amd/WVyj7rk10i3UT/reSXyzZJWqwNUYvsiO4a4iLRN7qGaAm1LlAmc8NNt3
iL24d9Qj9+7AFfH/CVKXNP6saDBISelurBOw+hFSEmoGoOBqAp3UmFtk3vHO
xQqhJzP0giD25udsnCK+4rRx1qbaEtzoPjYZ3ERASxWQcWCFoIDj9kjumkwO
gDKcKE8+E3txfSjRMzUQtcZiHfH48hpoLf2z/KuopGPvy4r/KxIKcRyyABKZ
UPxNWbFFsiMcqJanBG3v3TmAEBMT5awM4TSeVY2czkXPAkjeA4RnW5E0PGeT
HmDSHOyQWUkXaEnEUrOzAB5xEoz3F0YYdZvUkjWyTHL1WyQ/keFCco+kMWsZ
hFp/PZUrYk54yMbegg18KPOrvfg2eRncegJxVQ1FVaged6XPx01ASwH3Pxcf
nnpqFsHUlOQrFBjlgfPbwlX9AesmSc/GkC6HDoLadFPTEmF3sDiC7EGhjq3G
DCNYSHiTrikeTvMCMkboMVK2tCQNnzo4WcvUe/66onwYE2sc2GDnP2UpmcRw
UUWvtIAXkTnXJxaucCXNhI9zu0zZfQe0AwlyoH+cPqK9Tt3KBrEdY+C3FXyw
IUp4JJQA3X60bLqnjriyQkcDRGEmnOck5fJOVSphkylEDrWHIZve7VOifXHJ
H+kQw45p/iynzW1qHx4E8sEj2rExKQX3dniKn1aU1fp5FvyjPQiqliAXFlOh
STc3R+Me8kkiBdw8vYPQQeQbwnPakowNw73cbdgH8vQlGJHFebvua9cjKQew
9iXe3LpZeekUZeW8xCl9awHMHxFNDgfjnGb5oQhXW4WQZ6qjVBRXhz5IAfEN
TQy/mVT24k4M7zQ1TeiJ90l0IVllnuS0CGjv3lQ80uFSnHrPDUqdl+8cF+Zl
W/geyMw7lULRK9nwDwhn6+4FbIsPsdxHatq4z1TYz3ghSRsf81ZPslXPFxhq
QOMtOguWeLpJjKHpYZuaXQQgkOcm8DkB2kWno5yjceBLRDEP3hJuqX+LLwVJ
Fb95GF46S1gfgAzJwPbK8zZ86fCGl7AWsIMs6KZUYLO8Zu5MzbnWe2wCkp2d
vkLdFwli76A3fEiid7zHc8LKOfJ0F8ifgihdFx3QI5JaXCzATGa8fJyuHJ6X
TLSEys2XwA6Qo1Tv2KBtwTKa3xOFTy5tVjhan1uLNySE6IwNSHELL/WuNZ/K
AGhjmgICCZ7lnUqyDTilIqHJkj0UsAwBL546MLWtXVs7BJq/SBpF28XoeZO1
kFGQ6eDbKNQ7QF/AdEu4otLG+LcJM+1hpi/2oTi+MCXeloAi+asYJ6FY2sIK
fqFClh4NH/w2lD0p7YA3I7RtbHcdD+NfWCbxjsFQqp6IVSMr6xsORHgKevQY
8kr42vGj6237cqKKwE/Q0i/NlwGh979MoLmnKR52Hm1acPEdp3gFswE/ZW03
WXjOxubJYKcMiCQB6Evb8aXUst2QQYaLKfDTYzjtAzaG84kD228iTLGkXt0g
EJw81x79ci5HcINU1K3m7fBb6BUA5sa9VJWlRng+cgDEZcgbCPHpL5fpeLt+
qLJghbHUr6sTygJ2fb/751PZ65kxH0vDbNze9MxgNIWflAnkZlZxaOp9yFCx
KCSVyJGcAIqRwdKuySshFxkPR4scDBhQ60TSFWxvrgEC/AEpj+dr3Lr/E3Gv
mwBamj+QW067f8YU4FqvpwnK3k9KX4H8+KAQWn0U0qGNdEZ/p4OMZJQ+DCno
LbEvP/+wQZppgNmG63Kbltja/BmHgEXT6T7gV609NzhPztfq5CjipByZRsB1
O9I+9jK0zQJkJKb8dmxB31Rf3wQan58NZjQrrLKU/66sL+A/YqOTLfzvskmc
buGSsVvYmDH7lRvcH2ID6ylMHbV/NYN8xfG8IA4Dg/fJM7ND/2Ti4dzGNg0v
Iqwb9EZUxBVsOxgDWIdmuv0VF8e0ipFOsnGfRzUydlx7YouCb47JY98xWEe2
AqngV46/FPCa+QuDsYGdS9dkvlkPOsdKRC1LAcBEzG5w91kvxk8oCEp88txi
uV+jwq1DNpMTNIH8rZJeymfQ/Rvx2VQqWCc1Ol93nEpU9wxnMjB9WzBOGe4I
GeTJHpwLUXZIXyN1Ri6iNPJ6nd+Kcb7dZv1gToR5JdMFfV/s50bsuSHjeeNd
aGYdirmaFLV/cTp/KVwer2vEQG28DWTWpi1guKWW22XuRtXaKW4RnigWh3dU
OQH5qyp9UtPomzHot6r06dGFPywh7lSs5/zG/xH8O6MGN2EvwoI/zDm1bO8O
Zomq1qGJ6ssEbB+VbMdKqSYL+MkkDguD21Mu0nh+f68b1JGJwjipjVVUclAr
0UaG679w0gZFu+GrpLUnPeIX/2iN04L1GCxo75tj5KXsiOD/EW/SPfCGDur8
tS/IEn/vB6M1judf4EPYb6A2H/21ng8/exsZbaLar9X+QbISqYsTFV+1kSVy
GMshrUDO1dZPGR3zdYIhPKbuR+QIA/BgYLOsENOQnh4qRMlrrFrNirwuKlIr
bMdc0Ypy3Vz4U217igstsdOcTCFL8kt97Sua6wu9lK0yRcOc+sn1x+U3WzCp
qFxMTwwi5+sdWAY0vdiYCxfkeXhXMOzgfDeSBok4oSYSYexzRJ8YtncZ3AS7
+0ry3NX/bGd7P1PeUAGRqH96NyidpLaI9qW0s+xJRUJ0LKsVsxZiZ0bC2J5U
7MdihakezzuFmV4zc+fXzlPvbLue0M1e8Z3gHgLNx/dyon46zu7Ai8qiFlfX
+hT48vy8y/291L0iDWhVfbo33LlQYa3zsAfqm1js6UZnrgw8C/hMg93FJahh
QL7bVvyqdA2NaGo8NpG24JLuiNh8KxtX7btC99xbzyZnPMHBa8M4uaSL+kjo
smEqqHrsA88EQwd4lITBhdEITod3TNeq+BH5Av49E0YftYtVMaV5GVxbW567
Qc0xwfEDO3OlC1SYGfEq2N2bVK140YT2im6VVoZvcsl166iDM0AEmUoKmFWy
4dGEomo0D/H+mEDp4NxlWkevv4gmK8917ooJStVEhtu76diZEP+w17fE93d/
NfhpPWj0rR2dvV4BgXZzrtQX/lmV6Nicr0ST6ydDlo8aCklfmuyZhnUANp6b
UKlkQL539qaNtEcZHD6H5tRpCu0MLeVoqy/N61cqDU0JisJHfO3dp38k1UvN
i9thLp9jwArCH00462lvb0D9Iz9LQgQ/ziQpqrpNLJ5hTd3wPhney4kh5O9j
SND5hyGTOsBdOSsEo7vL+msD5es2/R6k+r2ouuLFK7LdK7RcNQo34wgTCSuw
Hi+o6xApXL8TwaGBdKQutXLFMWp7sVSJ4ZxZAtxOfZOPZdiT15HVOaTY1+/9
lQDaI7nGQZpOF29cKPwOsPjPMZIVO6ovfTKPXM/SyKM2gkEpXrG03Zy7QlEi
ovHRQFrE6P/z1/HYFe0lYRHBrUbBFxzo4vlPgM2BL6i4goTN91YoQiG1Cdai
bzvf2XZk6wYZgFG7lxVefpMtUepH/mY/wIc67NZZwxDlkM5xLhVSJJKnjApW
tBa7epYIuscf+T9tnqPw2pN2xPrII+cLP70H0RKGj24x62WNt7lEk8QuYIxK
nGKTJnJ8mKQ/pVR9yHsOMThq2vkRuin3ewskf13znIZ8xxgFYvxzMR+oDHyI
sPz4VugkAg34vvs0+jQ9gNmVri8Yi38qoDHKV3i5XavmQZphatEnHCLpjNQG
9aSVKoC7PLOFrtFSOiiBpjXn741+u80K9+wm9c+0Xg7rY9gVaahu8V9PpkzL
J1eRJ7L/spIeeVszEJj0WQroTDl4Z+0zwwZN1PxEUPHasxLm2iAUz51mkx12
w6WDwI9Bnsk3c24PlJP4ex4QDYu9hnz/p0pvuO05AYkYxuwSKhkbJbjCywMX
gIM5LNKUglaHf6BbIgifE0/+JY7HadUccTXC4erYzy5UJmNXsoCr2kgYl6Bl
3r0ffrA1eXC9SsDHMoDNh8FIZTvVc6fMuY7CRpTGAQA23WvhLBZPyhe0qxPM
oZM70CuycML7+iUraZnQVIOfb/cNxt+aZbPDYOQe1dw6t0EAKpmOz3HLPCdy
ig2hAnhR1o5kMHNviwZNxBWDgrp0DP8Y0cjpHiM9C/uXtaLtTP+bh/+Pdsgw
Mrsbnt9SbPE4/VVkZibwo+cecUDbTEom5tjM+3osvCsWTzVHEjG3QlSeGVQF
gt5UfyyXJv2Um6nn9qlda4sdDO1jkfxsNlSZB6bpWH0kjZ7iHzcm3wy6U2t/
A94IyL2sd7+vZ36YegxdQ2OZr6K/Q90GCSzLl52SeHWFyg1PRnolU0qGH4Lg
JZcb5Uftl7kM1YzDojYizBWprN9puiiXbQ+ceuoDqwn9+e6D+x4cf2XzzhpF
iEcM60D+Px3QXMeLQjFMMHNMuy8Pzcgrar+o/14/bsNdmMeZ9YmFdwkrg9Ji
uCBXK2uy95TPTgsM841wQh1dIHYgd8GdC7+YoiKw8AHbC9Ha5p0lmwF4y6nm
qGFFbwKCR9BBZZM1KIPPyDFR1vo2HHf79yZ4Ipq8Kn0C/wMkjJV9KvfNWW1X
LeaUd0xuoAQsFa/0nXD84SeyKQjHyQQ8QnTsjtjkTCNciHRoBtFJ6WEH/4Qw
l5BsvPThSc/jbonGVgI5c+KRHB/9Vf7/6nTvoXEv+sHryU9unfnpSmdoK0fH
qX264JIAn072P0tWsPs24RiNZ5CergltDR58t1YPmZA9PWBrDL6TSAC+jkw+
88bcSbh9ZvFVE8HXN7W2Wypw6FZQPm/3oVTAaD/S+FAvUvIXDPL3MZ27TSpR
ROXhrdvbetAEOHbk3HfO0lEVwDJB/HtSRo86ciq3jyyKiCqos7/M+QszyVV0
zJZ29lTMPfJO7the8hnB/89iBfBN8K6vkmLq+GTaa6VHzgiwcSRQh08xspvq
ACa6eWF3OItOQf7PFGQuNtVDNalyDoc2QLj/DgEi8QRqZXqukCK2D08k7/WN
XT2O50i5YjThqg/cNJKWMEjHX8xhfvTNfiw3lpTsqxOVOOZi9OVRj1BYQPbC
lHPtVqCRAn5fyblPF17y3g+ZbD0eZFnl5zlL1Mgjl4T87KwP1sPmzs2mCSDW
3mFse77653sxDGN0EO+lIlswhSrjoxkRIWuJOHeaLIuLtxIpoDlF8VIejRHJ
uYF/zNG1NrkDyipe/nHUfNviHA+yTMY9Y16evyrSOGETlVi/w3N9UTuxgFd6
OHreweEJEaZ+eCAVUy64gomxuf31wD8/R6c+gwz1xqePymn0+6l7Mi+smQRK
QWutGW7SGRqWvrQED9HJLYaurcTvUtEKW/xcsmZXnRiSNTH4JYcxLGiMqslC
XQIGV056y3+eBIhtQdkLuZUKR8gULvqVj+qrBWZfKjIiIngQGV5cSshTWZzd
TYrZZKGtxstKkT1eQIz6sxhmeY2/gErn/uVm2Pz8dV2JamNvQJ1w7rF+ZYeA
mAg494zFYvfX3WPMTX5xzGrebbfzDXmASqX9LKKSw2LWQpb2XC/8XMZ22FuD
DY/rb66+p9fLqQlwn5w0618YWe22qprCvIAaTQtlZzKjkDkHNZ4HHNco/NP8
YGnRnXV3voNDZDlYBAXQxeXRt7QGTRthEdQA7mhqnxm2yTCvBTrCQNxU9ckk
30oBTFC042UWmfnIJH08i83knPIKSVpgf4pRbyn0pBV5zh1mdbvaa5NeCFap
lAr5v+u9xSVT20tb1PqsMCLi/qxi1TuW4LuPlnqSjMm46NTpp39Qy/NcOxd7
DuG5kqattOiztweeDSUSGI6rN5hCvZ/JIlWAnHTf37Ids5PqJq5penqpInVK
JFqYvCi6IwcxgKc9xkV2z4/PbgntmdBAJjx0WBUv4NrAtb/iWlcBv50oIxoT
Ao7mYB5YQUomF7UeVH6DM35njIN45ciJr379nTx5ux6RWOQP5AXjpUM7Ka6W
qsNWuPc8pf36edom4xEWD5mgqwRZ7NBpl3dc7HzogHCZ5KWsheDCGG/oy1IX
mzv1ATdJy9+gUSQBzk27RgxUxTp6ZaR82OVhTgwASGePNW4V0WEIZbBK9c8U
Q4I8p8A02i6FHfXYQoLM5xvFsWyxj0nPLZCyKEt7B9Bms5n4bX9GR0STAyEE
6+AigNOWhwTDKYtTM8mFaSFcQwhn8RegAVSdbwQiMd/VQ1W3dsmA7wOtrxt3
q1Pi/S5lYzCOGXcYyHUpbkJgW1sJrFi7jJKAsQu5EP8DKfJj/o5A/aWEXbEZ
SbEGKvMkt3plCn3RRjZTqwJhW0nLlPrsz7sSm/BNpBvq4kOjlXVyj7MKkdRK
ZzOLSaLeQUEFUv5oOUd7tXerkMtU2rdUEX/CMWljMDBanB3iDCEy/nAgG2HO
a+A8xJFjtvSpMojF6pNmBQiiKSoUH6k4CVQDt+alsaGQCFIdSkOr3dOLHH52
FaFt3RBsWJoASTM+HkyI7DKBTGFpmioSf4w8wcUMRG3I1ETcMMK4kRIGv+sO
tlTjow4snUeVWEULUIJCm7cR2f2gF0EGr+hqfSQGmEy9HHQYIsfy+b46Qwv9
JGzL45khSDnMdN40djNXmBLqREWCl1+aic7lpoJ9ZE/u2HIwttc9UCC2KJt2
+h3kwvz+5DkrI4J+pzCaa/t/Ng7tL74alegiVN75qmwhXLs08G/WJUHzsoAo
YwmeYlTwAsQfY8ITv6AhKJoKe3GZwy+/f9jlOjZh2lnlUStZNxWLMB55q1DV
SV/bvhyXF1ZEecClMSS0ttC5Tm75j5CvR8WxEUURESsTnRK7tXILSxDrObXb
F2Rt1+NZrAtA4pp/OAtsH75AGqu+IOPj4u/MFGtdO2Qh65q+iF9TdSPcQgvI
vDAGQmdFXONp2yg+3QTHb6EANBX330BOE8n43KkbFXMONbETp7Zq3n8Wh9r7
GZXvyZej3e3g1Fc72uyquRPPmY6d1sejwxAotLB7KYIFiFq+iBv/m/FXIDvf
FBYyUFffWJvVQ0KQvAYpNSLmNYovj0iCQ/1+N17Ao+X6cyAVXtA2rCyR2gh4
PvVT5QZkcE7OfHRUgdz3pXDf8VoNXRgyHq86KyI4FY6CdHyL62lj6sgnxYtc
oull4M5+uqeZCFkq9/PC/NH97g7uvEy20+vH6mw7z/QVSCMCXN67AS0AYkWC
xSdP2KKaktCa42yT4NWkae2qH66Jhj3xIcN4Du4bw9uTJoaGAFQI7hOjBtWo
3mw/svQYsVFaCkvGsSe9jS0T8+Jup03sEghHfjrfC7/wb70t2fdHTt98t+vc
ufKx4TPhhGmZNDocryjbKeNX1Kaj9hY+9711waLJ8hSFdcZgtO8L5l8I2ILC
rBrx4T/Sac0MN/LBtrVdzwEbZQVg6EiDHsdaK29f4DTo95xD72Vdc5XCxmpE
VzxvGkN5p5/jUO56YWlQERmhoh/nlYqneOUu28RYx8qT/oFbyFIQ8uUo67Um
WVZXxEPl4nghPkJFcCEslXcu8DmDRBr6cyL2hYPKGhhoVULa4d7QBrBsx74/
5YcC4oLZVHpsS6SVWInaBfUQ8kbHKZ4os17NC9UhlWx+C2xZfoVlztfsvPUp
zrZvGEOS6h45s4OMJFWIW9jAWOY3xvgaonoKBNKUyAHu4VxwS3GK8aKdmvC2
ujekcWDYFj0ZInD2YQdKDU8+y66vpffwK7X1AHwQMpGTCP3odbOTy/MI1NLj
By3v6f0QY0VVUHv3LT++WgchIV0D8crSMGKZS8/6h5p7tjQc+sHk7DCGqHl+
ZXftmSr2ATHRefJ8x6xKtjrfxzWXaW194DO07CUyZXRAgTPMKz1Cm9Jr7tCr
GUfKCQL9aiWEqKQMUNHSgyVsg8oMdDpXxiJ26mzQjzjwNtgVHkXFajB1gu0q
Q68SWUaH4ccGqmxYc9KM0+GLp13/AzGPSOcQJIlOTF/E4JJosI7IwNyO78FI
Xy1HEIKX1bagMUlfbIDiR8xpAkC2e4KjmYUE0NxEMlOPZbxKo9eHg7MFcy++
ThR2gziphMwuQNx89JEldSchdv4Nn9IsZc1htGNuixPDFb9pYyDeI5jzl6Tw
294ETe/Kz8SQHqoNRiccSoz1SefGi++4eJlypQfoZbx6DOnVTDtITFJLGcOQ
Ev6yIqv9j0WssLwoCxdkP/44IVcF1oP4b/3X89PiOlnfTdPYeE9wyR4lYtGR
t/yb80kOzkAUFDyTHsH7jW2q2r2RA9CJjH9nuqU12cqjN8OjwvlOtmW8v6hj
HZLVstoTb5V6vOWm8nqD7EUSNIPUvDQNV382Bfk5Lx9SNC1at4cQ/z4LUvn4
+uw91sABMQInnYfbZ40FFQ1R65IJ77fO+sdwZXYri969AGzivjQ/415cxBIt
xqyNRIzDM9TzwPvGaVxF+++w/H8ERefGQyzHFowVuPZA2f0LE6h/HkO8V4CB
N3fDY9rdWXKIYhChEJCbis/hCVvSyf5BGlpfAVwga0CheWMvediJbpEzh6WB
1S+PbG2XLjlU0XMUd0vrLg+kjV0+6P45d+kPb1bRnR823rUhDzz7eN4rQ1VN
QnOtARL7fELvhM/2mxSuzCO6cYpdtsfauL1q5EWXFgoWdjcTO2yhrjg8+2sl
pP5uelUcl20n+baNwZQfM3iXboqJkXoBGDK81MGAastKHUOwk9mLf/OeoV9U
OwC5k3IPTGltPXuIWKXTrsstlpem80pz78e73EDuq/7/UNg6A7C0dd30wByJ
DDx1RcJEGs5/jRZNVNzTnKsW6SvmIr9DctPqqzLnMGNfPwTmXYBV3r3DeSbw
/6O5wThMF8H/IED5nPvyxpYRKXhwHMlHvx8c6DJreFRENrXjT7IgQfvitKrY
KuL+s/8lOHT9pzQjkj6BRlJ4Rn94vNKLaQKKhkl0q7UdGCE61stc+OmUQ3dU
/65DcK6dOqYvDgxj/MtuIcf1waLqpROYG8X2YxKkvdUpXr/QPER6pivycKvD
RRWUDwTeTZ4BJe4zuHf8bR1m7cQVJFz4LF3AYEM7qwtYlimANvKgHMf2pJw8
rKD53MWI1M98li0kBw2gD7Yw9lCd/F3v6l0I5MzVEkzSVJxzlWtxqQaa3XCf
FNXSPszUsQ6T1yIqm2uDf5FJ0/a/2IzCY/2ZDKEs9eyTMXHQauNnPnlYO68E
ahLUL81GgfA+aQp1ySbwbGUn0rSMKaLtI5ckp4moE96z2RUKJmsI6/qdGyUD
pjUPQLQElBwJrjBvpRjvTbe+slecp+exXgqPNx2lznJ+FkQ64FDXVBx7xFQJ
NElS16hFNd9Sawpr69Zlg2ML6bxrcNM7bLtMizcJ995WnlVMjKlJL7mC/spd
/oQVTx/6nOfAn3aEAEkX0StVpGdOwnbQ+J10H/tA/NsIcds5lmqLnyqOUUeh
zXpgF4ZDGh7KxyY2576hZIGOSatHmuIYbbzclmdSNp5NiRqjpqKgNgyEh1pR
j7ToK6Kpa0n4HXAWcRi9mUrISc2yWOCN70zneCAtjUa9yFpYk1JSoO6Ahank
lvem3fPixzel6JGswNuaM7Pk1xPFE2ouArO2cKoz7T9dH4OMyYN2zF+3nDPn
2jR4Nnxs05fhkN6YDcgmaJ4Ormi/fIC1FjDz7ufMaOCYKuDE1L0x6CH9XE1e
QthO4co6feIbd7zsOt81ewXIuJeDo+1en/JQzuQTmEdCXAtU9MC3GmSA+s70
+PnrW0u+DLm0ITZzym5arSRiLDJ4IIDyWBfBp9ETCSu3LzcV4BJQcTV2n3Ro
a1qkZOwUIV+RIDYMYMAxSScuRIz5hQXraqkMG2npmffskf1qICQWTOat5yvC
0eGFWe26X/XqtjCoRsTuhDGRmMkEpDNFZaLwjCXa35YERSwrWqlRj80c37He
qSB3Lj+33XwfABCC3fqHhhsrYk7pHaEh8U78tsQRGrFkab6sl3MQhx/WunLC
2RG2DIIzi30murdo74XeCp7Enbk2O4njyGeiEmCM/bzsBq5Fxmx7nJ4uFMaD
gcU69jXTDZFOVOoJDfmOekG1N8hqQEULRATZZOkQ6OEwv7JZ79xrsLPui5hH
fl7Wn06kn4Nwqs9WGyTMe9v7EbtdkvcYnPc2X4JEg9o4wq2X5GMiVTLfY3/v
BivMAtfXO9Hoe5dcVmktu7cmue43agAJqJLbSPfbbqHRQQk0iyQzFMWFYPzn
rjE2r57lCdeCsR9jBv8wgcF3Dw87O4f6wxfYnHAXALgFMQiCh+BebTxLAbQb
uZLLJ+lncp8+SZMaV+yfaHV0wWJYEVGmxe52AyVfcYDo4+stBlZpQQcWeG+5
iwPWmA/Ys2fFobUYF1kvG/OLTQgbbrV8Ew16C+ZshoFuJQ3gAXkqkjK3Hhyr
1QICBcw1LXOuYrkk1i5hARokEGX9q3q7jsmKCFnLITn2anXzZldAMs1qZsWK
NyqIa483FEdonLaqrOjjRXvXC7Y5cgubngKka3irn0xx1Ci0jZHFJwSuM3KF
BfU+I6OUFdookkmOJ4ic1QreRiwYVrb4syPN0CAzFktwf5PUKoxUIcXM/07P
JFlwvgO7HY4vzfuCr65ysoC0Rto80iN575UkZelJ0NPxOr8wRB+Yz4UYyTL8
er5Fn90xhlxxsTKb6ZLBRZK1tZKyufI3e8egXZ0b+6rFRhNXXgBvDIhnGErb
gGKlJIWOnD+s27e8s7w/PS+GRGfmwGVyoS25sloXhp86Xrxi4TYrjaHEEaiG
RpkL7hJh2V61BJYgRZ3h4UNYL3tLZGokWqgpxI1l2VoF4Z1gE+6wGUNIU//p
wYwQduYlo2L8msmmrAh01ESq0muIyT/3RcIx3keIq4wdy7KixsK+3R95eRqT
groYQSg0KxcQXNAvyov86NLMSiCHllQwPm33JczWtPc44In0RXvZQNMa5bbX
LqeJI2uSgDRYV2pvVQbQAedykM1sL3aBsshQ0/ljNg+r0fGg44EohF32MDCo
cCS+svuA78UN57yijpppJxxXR5YUtbD41v4Vz4BNKyAypQ0EglmIVhJjSf1u
7i6PodyYOqRh8sSFWPuUM0OusA5EcOvHqPEMuagzOQoHc1myn9dGnvN0Gp8Z
hQNjK4IlpF7ztD5dT8j7PpE9u0zSOTRdnYYywy9ZNnBfdHeGonOKcfp7nf7c
kgkLKFJQbV+Px8x5oT7ABRmvKEhKFkhDlnyRA/xbBoYSDumJ5xcdfT3wmkN2
22U2vPLvi/R7QLQVkrUpzuQvv0iUzDtkBKBdZIxnUm2OONKkFFhH0UPase5c
JEqk4qLqIhGUMUxh/JE73VT3UHT2m4yrmfgMIktZzZOCCfALkW6IjVqm7wuq
oC4CyRvTWWCluQ4rX5xnd3D+5RIpy6M4a+XbuCI3rk9xYNQashXIDU+qJ044
r3OrFtbrtgjn4wznK9KjIODIh/RuHFkSGQN1xY3Y8Pv8Qze2e+OxjwVT0vdh
NyOTPnXFOAXoHtP/0aiT0SX/d2rImRR6/6yXZvw5x7i+LzRQBYgNZ7Lvk5eP
Jg8slTxIuP5vz4bOMSxzs6Oaqh2mdS9ud0UQol92/QDGfe4VmxAOXbTxYgtN
p/bTIezwuajC6wW3JG3e4UnzwolSUTFW3qzO+KJ49cpYYK0PmrB61W5X6ZUo
EVjWRPc2Qkx6U7qyC+1W3/jzHCr3S3vnu9bKUrHk8eiRjA6Z2yua/nQn3Nej
qCUI9ZzjRDHismzW1Yt8qOSZlTyV3S/fwf9WP+lAGsx/d2n2Og1WiBelPoo6
p5MOIYxt0ENGAMitcGi3Oh8nw9L5J6WoOKby0so0nvelJu3iJXTqz/6KWi0Y
GSXyO9Ll5+jxx3yj56lFOdCpHFJ2n6pYVGdBITeve4sc1RXcl/6xLXco0Au4
PN9Vcchfn4wG49SVY0EMPMSvP5w3rMBohUWEm/waiOchfnLhdcpjCBnUQMsq
aUkuKZcYrEm5p1ZJ+5LlJnOV+2DMk4xfJIN+BDIqWyXKfLbcUq/ksaKNp1t1
tesOhUIEIOnDgl8Ok/ebh8mCmz7fRFHApuZScGPn64rSNG/uhLJI9+62ElkQ
wUrankH4Y16cU3WHAAcdQQG0dpmIIWwB0Nyw971SbDl0Yk9I+elu8esHX+x+
aXelBdKk/k/97GZB84lNf7mo6tCrmt7emhxy50S88hkZFxoGaoDuqrKM3Nfm
mVK8gBCbyOTia/3zrpZC0lGj2I0aPNPzHFm9a3CVZVUz1hxsFczkuyYqXjay
4joEANmqkDvYxHkyKQI6kW6zojsbxX9VC9iDlKwdkcF4p9GzGtg2AQWIQlM8
Ft8q7LrcuRBwCv/OXQINu1fePuzufLAtlGXC19UT1PfF8cIoLUuzOL9OlfOK
UoVmFNhpwd40gv3CJIlw1qefrhowaJYftCV3/tcA/Ifbf3OmjWSpsXHuhGiv
cZ5zoWiM7pUz78JrUlsdU3uMRyDVcBvkOeb6XmgDLeXOv2KW9a863wzoMkxf
/NL9zozMHjVaOvoqd488TYnDmZ9ERZJDptK6ZciONzqbhx3SBdQj/uK0oTP1
8P0nHKzTlUE4sz4TMWvNUl882QlTJY7pMZeW5ebx4ZurxPR+luRu8ptrQ7oG
F/HVtXYqS1/6DG7QQC/raXws8TDDRwEysvGwnEpc0V5TK2lwq7+W4tYr9x1d
ndy9YNhQ/pI4p2aip8hwBYgKJZ6ra8TQ8jtU5EVA4oP8KPyqn+2vRwc3gZ8U
9JbhZG2wvR0K0qnCsOvfBdlaW9cbKdRJLx0XbTKIrmK2OAYAfgUzdJ407gyh
xwaCezYSOe3WEtN/twk4yWZJN8sBbdU+pC1KM0H5gHbiRiuodZiR8mimping
3omCQlEwbQgZCGPxP38uTeT3sbIInLszVMfgzfDqPopxv0yavgUHJ+SKFF5F
mz75VwLLZuGWJ4Wli0TDudjY0OGUxkenuDtZYlcTqpAfldJBmX0l4qwOr/IR
aB+RIPj/REh1p2ZI2r8rhoseK8hJvSHuPwAqy2rcmP+bjx/4IZDf7rqIwH/3
Jqtz0oDCcQiCm1U07nnClemCOHZi/Mn0yZfyjiFrrOpbjiUSbsf5uA2RoQJO
RWAmvfe3HWgXCZqJ4IFxrl9zn2LvD+HNz7ykYb0uuD6efaNsEgMXSKnxll0l
kV957c7D+gRYyUgoKhzX0vO8rEmSFDG5IJCiLt7vI1FFQXheoRzp5SLCXVUf
iQ3ArX6kl9tmu1YXTiF4JCtpROcThzehixrH1UXLx2enqAjygrmhhQKZilOt
qCBmCjV2sTvtlJ57H2Fnvo+CtHGm6IbayZqCgL7LJtDm2aVUIcMM2BRfT7Y9
HLfb9d8+i0e76IPkan2LLtBzagnhx28K7r+rXb8eUM71gDxhd74Hkio0qqfX
7M/9X66mMb5NlLbiuCQINbiWKzBk+Gx5+CHfrpLUfEh8K7yMdaylxNUF9G4k
6nhronmSam/6RvhZq1uQD5yo2S7idZ5tkfhTigMj0iMHiAoYjPdi7Wj2X48A
RPkzLWChBPTYqNwK44wEQHrqaviTXniARbHSEmr5W3NG+6XfOg6LkCwn//+N
ZqAoQHSS2C9RtcCQ5RG7MvDoIiWgmf22A2v2zQeZK8xOFoj33MTXUxzgxfca
qu9aRsgEIkcABpQM5XZbF90KdnQjDpzWG7lr25/VSEIg5twBITguujoc8BdH
m+0O3OpsDPtbIF6XlYDU6pld9em+rpLDJ578gHgKkKqsNtak6xyd6uh1cGuI
dWKAjKTshKBx2i3AF5A0iENXAdwUEeaQKdZ2pszdoaRyrdAyIKf54O3V5koS
pAdlf50wLfVwtoeOujzi/pjV6xl7z2tcONmwBA5xZFSaukO1PX+SttZUEHxm
ui6zqFkF1NzCOR39mB08AKZiUDe5AwhKpluVvqK41aYNX4DpajD7wqOAdRjJ
PWixvnNLAAnGfcJ84yzMJSP6pVjeQaodnOLZbpYcwD6xuKk1ADqvnfUs922k
l/N1MCk6B0xPBlrjoDlxEze/BP0i91K7I5d1hmNQHZvTCVf6ZQKPMxtEj3mX
nvcIiaPiEO8y4kXNcsMibwPqeOYbNT3lFrlmH7lsz/RbvNjqie0sQjQRMpuO
ldifukUNvd0K0Sq48pB3T1Z3vAyvzND6KPduKdNJlLg2ZDOVTkqG9BLWi2if
DGhD7AynZKnebl6U6CSXTo7k+nxMmU8Q35RFjRstyFliOr26uUi++15kxv46
AeFVDYDvFE2XTug6On75TJd5rPQ+xG9s65Y73/dPmCJ9JmMwQ4JAVuj07YSi
ADq6QG9gQRmBTOpBSycsFQBW+fcDX2uJl7ZdULcSgsMGNGeULI3L5BAlc258
lFWAzJivtoMWZSrFgXa3CetUGIRAEYtSc7C6+EWRSpAnXo/fLRgWZ/euq/G0
DWDSqrR7PDBkTdUI3AVyACSwdetsqxTBBcBNEft0tVJ7ue0P52VRjwfSzeeX
8kDui9578P+se6jFyHZCBQHqt/o4Wsplbdf5ToFOjb3R6vQTsBcHvvZqxzA/
galGWfnFryC/ZfZAzJaw0fZFzGG461THjfnWo60Qn/jsVI7BhKJRPSiR6FOe
MWCDl4J5Wb4uKerzNlGe7EkfLSQFBIi0KdXy0edGfOy9UZRwlFqhLx9vfqQt
Sj+t+RvqW7KOzELw0LXcIszhUxvmqO7xiLlql8kEe/Bgl2CHPK7syY6jFNjy
xv2q4XLsXZCjyiJVktlN/6L5YvGEuMC4WAxoNLw4UutqDDqAE4SIB4SoZC2I
vi8RMRVgkM7qWsFRdh8dXRC1A8jyQaLfy+aOiZYPKq6rZmX0iTXvviL9BS55
t4rfCk81EDbS5ajjovw9UfyJwi4NUxT0mWDfV56fZTGbC424KTGoR6t9sVfH
MLftHbGSdfiqiPU5JimxnBeEVWRxDfriRGvQ+u1/8i8fEuhZVo/12jagjg63
IxPCMTbLgBE0KaCgpV1aLyGvEBzJrWQAB/NiAQQGey72l5DOU5xyfGwlUinB
dWtqipWqWrrYbGFQs3dVl7WFOnltR7anzm+KCZ0oJ5k99i120TuDSwDZ96zu
HFZIEbDN25NOd2Dhee2g0voZT+yOzl/gXuv1+zigvFmS3H5Waa91Y8BKmdHU
bBWdUgzJ5B+/wfMjTlbLF6JBWulnyRcL8XNENTvawpJUukys14SyOFswD6ig
6AwBN9SDD93FHlr5eWAK2XFb93NQe2s4UiFGKSaptWbG4erXV8rYfoao9jmk
eHWwQZrdobxGU4ba8dnChQpyNiG95oNJY+afv+qGqeZJGyOt4CX05+GmbN7H
Qx7UXbpRZs0h5fNzq4LJqJI6brQeBwY1bIC00AwBfmN6Kh+EyHfM9n6CAqt+
3p1Jj6P0qWf66w8leGitFV6KecWBalRRh+AgamcxttXPYUBuzGMl/mqAbgEh
J8wH/3FrhfUxseF0xXQvzW6uXjwG3Xn6VgSOfPdB0vnRr6NQpB4UF1WRtJt5
Hek2yOVq07wRAAcTymUp8TxQXNz5fDL3bCN5ZLDayA7ZnWoK2fB216mof2MI
DLHJGE0cjEjhKOXtQH+43fqkBq5VhIEKLiypDDJMLA1VDTw7CjSGQjAF/l6J
+/YQE7xhKzdTXNLYsBmQb4DsvpgGr47BGzgjjIBFqo7LvPyHPGecwJnSlk7I
xU8MPEpqF/lGeSYGgyPHYTD5oT/YU6Y1CFlJz5eq83ICAwItkLZDR9K7bdYQ
k5NgPQUGFBpiqmsMS43R3qW8gcjEYoARnlDP4JcmDt5yvbLg4kkZzpgycl7y
/IOloQon5KnFGliYf1KVYWrjCgJ9qG+sSPLy1kidQfnUZLEsl98DTjcGIj/I
Yf8mqcZKVZIRZCqGpSNdeJHiEjmfGvNMqdhnbqAWJDSGwmlhZldwb9SndrBR
KPkQogiRcnFVilwxhSQajpm/Tntfb/+rYLzSqxA8QidV/IPqB02doMPJAQkS
xsekINucs1tqQqxn5pqwAwZvhMZL5w8rz2E6klDQLFr/XTl7Wta1Zh97TpsQ
PyvBO/AXBZOCDiBAVswMsGL6N2McEjfcjWHmeTEsXW06yt1i0mqdICgLp7tC
4amN1o1XSNDSdv8ykFrbWxWe9crhmCQ92xve7bhg8ojdREBSPm0nMujd1nzd
nZgL9XHewyZdYgr8CTWk+s9Q+ViOzgIBXLFuR4713g22Nt1S9X9uBAlWgCVQ
kclcH5vHZopzFxYbZF4Ep5Cv2A09APw3FAJW/auBi38uUgjp73HgC9Yl1zg4
vKGTTzDyPUL+CI+tSkQ23lMi7Tpouy5uM3OldOMpMYkvYWVxNc0SLqCHEz0f
Dr1uowFJZ34xlBKsOdINRvcPaUjwcu1a4yrYXMmZPE56CtDRIBzHIe1jLbBG
ikr4F+NRVvzAWSTqHM45gE+9m5IcogqpYKJv9NP6r1eG89qK3a7AfxuVwcWg
Gj4cVeG6lVwAdbn6+NqcAaPCG8Mk6Iuy5a0TTjCgLRj48RQDm32Te5O0thNI
yNvfxDGUk2Q/0R0LtBLmGJ/xnTV8nnrQlDQO2NhpMStuAWfcB7fVMBie9rrm
luvVcJ5JGPn34owQgBEDg5eR4WqfMX//rsmzDR3VWZO4V2+oi6QBMdFhSOM5
cP9JOKeA7vdYLGFvsi+WnQcFuu9St7jNp5ieICMPhK3sbFWSeTRKQiiCQ+32
SjWmaK0Ko/7T/nWIj2FMGFWw4YLiiTDfJ0nrsc3x3jrLn++HOaYy4qn9v1eC
5SZhLwIkWe85Bhi6NGCKTBd+byk3j6qe39FDjtjKLOMwuHFp1wjGH2PrxNYs
HA17/kIvLCXDCOPpDmSwnOulLlBfKsRVxTEqgC6IJgJwsksEMVGvE547i/62
lg8gIGKM9mhFnNJ3Z9U3FObUkW+3T0QUlLcL1Q+DPL11ICIJYeb6Dy4NGKIS
Q7rAByHJeOp3y/GzZTRuit7QHAf6DEh8wVB+LwPtCgEEIub8aolx4TxmUR2n
mT9t0t0+h/ypPDuCMib8UNnCjeRE3j4HimDXS55L5uiTRGHog85gHjR56YKL
igsk7rBRo8NTCGU6Qdmo51d1YXJKGnVnmGMc7cYEgz5g8IpVSp3lBF0wlPus
XIckrietTCSeLsVvIhqFdRUqR3arC8CKUGe6C+e7DxsyDF56y1oYXosNIMKj
Ra1KPAu4vzu3/jh17Hy9u9sfaCO0hFBJcTritM6Fnnvcub+J5wXtxqlKaMws
kGq07GhiE6BblCxNqwNN4ucxXr59JwEYxQBSKMJZ7T3azrz4eJci6GFToR7f
Gb96kcX5lLBfuLy3F8cD+oeoSPe5BILntFp44o3llmv4SMKp4Y86MjDBmMms
ftyRyzPVuFS0AX2EBamcBkphK61raJdgaXNj4XxmoPF3xF0NQ45fBZeemc2S
lp3B7Hl8gaFHOhqATMLeiuteVFRTI2577lnz1rmFXgq4Yfl+CN2hKixpCSnl
Ie5beighfaCZyqfFhD+McSw7urm5fZA3BDV4U4iNhIQ0AK0M0L9Hbc0dazH0
nO4CgAryrZfLlFur1L0j7HyMR4MyUAih7glAo/1+mb/PHz3PSjb/XhQ9rSIo
eaHdUuAu6T1JBSrm/M53ua4ael8bOFu/io/rIxCqALzeFi0Bf5G7TrkZ9pDt
H3RsHVUeEk448dQ2++/1ohySJSrHvMvd4fa0sPMWjEVGUPXzVGZ3A/gX4ydP
4cN9Ot3y0ShURtjkwxoT2vhgulIL/SUbinBQPFEksr6tUB/AmI/rfSCD3EM6
qGOlp5epvCCGIVckMDbbvtP5TDOnlA1x8FZIJ9sJ82t97SdGPCdbY3sq4K1J
IQMKj7IaNmiOd1oWRfBHkJrNa5ysRBNtMGdWlvAgVcau1Rv4dzVEOG/Kh8Dk
NbocAr2PtSvRJrczTDJvTEJUTNnrR0hCT+wM15wIQtE4FWwtWY4wNHr6F66y
WrMvhi43bXOxxD5e4hsKpCdb4JvswieWxuOAI+A9jVXQEcfMGnM3+pxOlX1B
Wl9aUmbuh6xJ1J/ezoUhQLRRAKTVkYvN0rLaArylQiwQx2wq/kaGiS4DD/zl
kUEn4ojAiEG3BEzzYrgUY9WjJPLezNsYGwwzbnsGc4TcubO6POd4/ui1onGM
L7632ZtuJXdgo9Df8ooUVV1+vigWuHflNfr0XsHqa+LzaGKSP2/Et31wGVtP
8cjp4JYBv9NrXCYOMWJfCkArMj5pGBX8Crfui4N4+ci74mk2ipeycRjJgmAj
0JniN9GruO4xQN63ivF1QUXR9UrYd4z8pSUBwdhBwk+Ce0navuNZ6ZKsC1wv
xy20n9Pgj7h9Bn+jkx18RHB6gtKIBS0vsF1eKEBo66WZSXZbxBLEOoTLERIj
EMChB444Eb6/vB7NIfQK3R5JUufbt6JsgLBjp3Ro+PcEF0ajcEMT0wTichjY
KzZz0fb1FKwRNnu28chOBISkozCRJ39N2DT6XPkjBM0TMTq7y03PgXXpklyI
Hqcf1KrL9ejMivr9Wb3nQbzD1gD9DaE/Fz7G1B13bTFF+VCZvGiKG3bdla4x
jyMhMTVRhpXnlOBZXSucS7fZ/SHziSkxZhMAaAZPX1I/BaRpyep4JXwVIW06
JkH1hcgFLXkxVwBLDkfoun8YTXKtdP95rzuJjtXcjKDo6a///YR/CtkI0U6o
f4uFTenIwBbIIe0T8fAmAAT/UAjDMTUKU39yq88rpUzzMH77WkJoOhJsSsY0
2L8GHYhWtv/mSWHYlA51wSvlxEdek9s+iAp1ND+nAl8lNQ7gZYsrSAx+auQh
r9h2SPQ3F2Q/pdQpDFSmOtvdfhRYq0J32u77u8B50ZBE87Fb209WI/BmkJYp
0JhSNFLD07iYsVVVNSqY7MfnWQHVHaKRyWnSPhEYG3mPOyOEAcKwZOmSylZx
fFw43Gy/9DCBnfYOV/xIG9lBpo/ccmV50a0EvXYM2e4X5c0t4eEJHePCPPmN
oYJgLX/SAuQE8LmRoWpEI3IsPMxGP8HCQpj5KJ5HG67CQlGGsJ7vvUx3xSRm
SFxeBeKjVMYJHXgk91sBmwyo1nh/EO1EeX9ajvjL0zud/ukEXtqJt3gdyhdO
mqlRhJtdVMfjpIPEXsbykVmTc68bNqhO5nXrU4Bs1qLHUujawU4kHebOkhj2
DI22MnR/7+Uviy061u3QJO7+WZt0sMBsoADr35f+nz1FV8cBLA0W1vgZxuLT
VdLxRp19tmFMwD4zs0M/2ISoI9uRBvr45C6ZMrqGNRUZDCAtRc+A7/lBKcSa
1HzJtXpZX2fD7gVXQhqPUl9Js664b5rYZWIEM5msInwNUmwAt56fM5FEcFsP
JWjrUBLUDgAmPaCWqGcKaWniQaA67pvo+4Sp32HERJzlSOP/ZCVNKVgOtyeU
QmaPT5ThBvWtLhCZt2RqxNOMrY20taDloVq4/V4mRc6lCCPEAQoUWU/DdDWX
tlx3NqXiMETrcMU/yBLv6CpbK/EKsYIsTFXJamNVX15Q+GcL8IlKxr6kjHa0
wTfVCalXunPumgBMCxyjt/jrnEUmfLBSnDLO0ZtesWc708Dug8jtI9JdsLQo
yMnwNiq4P5v8k/iDYzG989nmtuHxI/Ae7e0KDcbAp7qnSZhYNYclkDZxEPFz
GOcwKWRMAX7TXRxNRIBSz5UtszgQFKUlFSduuWqmSNAJhK6gyO4j35Ta0BjC
6/i/e0SVDD/J/DFSKN6gGyOj3KXMyllM/2EVBl3XYKW57Zj1oef1MQ6Cu6SY
YS1R296S38YYd9A+EO+X7aZbW1wssYNNxQpOIRpKi7upapmIEJzt/xrktE5v
WtoekXgSXSmC/MHtX/oOteu10WytXjZOvZB89uL2G8A/f1QFuoTdJpOFS3nx
fs4Z2R2C2SfmQMwyctEGoK7yVx6zPNVSo9rgqEdxLkwXeffcslc+8e5dKE2f
6A3cQBtVt8K6/ppGtAW2eeVWDrOqpkEtNXhpkzyH/Ofb8MWgTLfOds2HeKFp
BPtpyBt/zxGpjQY13qepfnzKp+8Y4d5eWMf5DFU6NvXbtQNxVz1fPiJkwTDv
gBgz8zDLlBkPIOkYpv0fHHDDWezc8t1Dz+lEHBXy13D592kwKiJKF3HTpivF
x8rMWpxKZevFZv6clcaSquAd3JE882xOX9cVJcoC/avEs3sLQO6eyf6SThDd
rYl9Uyh7cOJUDdZS+sTRVUiqhMu75K3kRufZ1+Jiqd/ke+GfkrAP9Nf1sIFd
kNnH/edEra46hp+3ivpTSXLkVFBd3cCuXjx944uOo/1GhZPbPY3NpA6nuUwN
YHhlAoBNCaBFm39TA/eZsckzjTSz5y/UamAfLLDxQ8RhSikYluX4t3zPDY2W
YC8LPpTGFytjUwzPL5mtD2un5q8OBzgOxhRmGGfQOz8esFDeXKnbYUoYm/vO
iBVsWB0KSVfM+Y+2DxxXCz4+Rbuleh0h7GwJIxX2PuylMnqf70G0Hj/tM5NQ
k9eMviWjyI5skAfFN+A3VmyFulXmEKMed2AtpRNP4LU6gZm+yN1yNMgROX1K
AhhqNNt4mxBmVdRqahcb6JYnn/Ca25S2bw0W4AL34XufEhLKdV+g/zQw8c4J
9mU5OIXz2eBSN8D3SL0LDQ2PKxp2URJ6wPWldEr9y/2+zzNYtOtOgDTcq2jr
1vOO5jEMAMriI5n/zZJYSF8/HJURFHhCplS/fKXzSFUjwRKreak9iPRz6glS
RcPFEHGQSJ3bKi4Z7sNTFGe2xe8Rtl0dxhSls5T3Q+3uX4SvtincF6AgGWnZ
5XILkdBko2ANuZiT/inWleFs9iUSIp8u6XHWoDEvdwJyJvKNQhtZLMYj3uvh
ZaRNyQYp+p37/gbTmo+vQ/nkHMgCAjniY1PchkpVdl1WG8apWDdPzXSFvwmI
TzkO5HBknS6euqIzu8KCOos1WxdMPi1X1ixliT1CzKCBFGOSrqmNcP2s3QwT
mUajdO6AuJLQKmYsd7sXlX7rEEf3PtV223JpMkEnSaDNxiUCE5s2SzF+iByo
uJDDrUpTzyVCSdQGFcwoWlirZ/rI352aSRTTOLEPbIk3v7H8czSSuV92DdVD
3z20TFTgn/fX+VjTjCLf/qR6x4ULBX9npiFRWb3+gg1y8RsNmA5jc/juQTVB
QEvhn2NFTlizMz6Q4V/WQiSsJH4lNO6XalNsSY4E2kGFDsWhk2nhxPecJq71
GvwmyqHqaEuLPdErrygfunsItL4sIgE1VJ19V6ILpHhSsAL9fMB4Y1V6AWRy
DBqBhYL/E/2CRkVMaP8nGpuQoQjZGRt/6SM9c95BT2WoBZiNH8bsSwtN6ve5
6kA9TP7hwDWUmRXxAEXEmlWHCh4YHERCQPMSP2ByykW94WCU0l+cIbM33vwF
/z99FqV6Sda8rahACSSnAvHBlKwrLc7Nj0NYdgqLdlBDSZedWRxSjjtsGhek
ezfUQmvIldakzPKzvzaz0lupFNoizEhcryZgEdeg0YOM1x/Xsmz3O8S6S3Ij
Ag8BabN4K5g9kdM8ofYnTHHhFGmrYo8LrG3eOj7F7bp35NG+tsm6pc/mnRZG
vBbl75tR07HrYdb/2Df+cshjV5FwlBPFzlpnlVQz1Os2DwRKUloY5YoF5IeS
S7s6zU3UzgNz8txbEVwLJN6hXLJhD7b5yVJxl396hjR+UFsSn8O7aHEJ+QC/
fPNmjVSFSdeqd8eeZpObJf6hn7EMrg30dwRxVlNaT+LGgc2VyJwRWhMaZAO3
TysF1n0dgwn19hNr0ofjznj5xfWBH1o3pG6WWOBaZuHBSTaLO1UCqD+8VeC2
4COjROHb7XxbX7obv5aD13zEfcPBe7EwUYaygdoxt9mvkvX+61VAubEseCtb
o990JhdyFUguoIlBG72xIYjV8TzTCWmNPdI2oz9jsFKs8GC/6wkuWP1fPEK2
i5bCKha+51RWQNm4AxxqV7rfak1oGVWrWo5DmenKMjaxXWmN7THkoJfYm3WP
Nn1UoqfLJXmCm7mIMFuj9cvLrY8sBNxQ8xOXJVjdy4YIPMms5uasR3wkB7Tm
gMYZBDBusBTjw/4wecijskOIMs0MZWIZm1kTNmZDEYDn4qEgu8j5t41aDDt0
1apPgiBQEpeCZQfHnSHwZRANNb/nSiAlTCwy+eTFYgUXHrKdQbzhP1NvvgGa
lBBBc4KPNlOzPIIGCFgAA/9mNEJln43sJXb45eal2sNtjtQHIQlzXMYI80Bs
EjGh7Kokp4FrwjH27f15IpFfPW0CuitKpR/aMFIRe+wax7D5sUuy2qPz36/M
2lAl6PIHMg8ikZaXYJgCWLFrYO9LSQ9vmctg8QsQQzQnyY2Q0RNdAt3nj+HW
ZEZXQWMh8DNSSv6P4Mm8s9nTdWtG62b5Alvo9O3fG3Lr4PHDJntRhB0tLSrp
+dg6idMbBgJxKg+CT4HH/7zebRncuUEEDrERL1a5Fu6V9kYzLz3wVaTPpdSp
1yx9D0HXk1itSMNre2+tMx+o0v03otVWG9DKQH5+zDr5QnKev0KBjhUUlfPj
xpfMCR+OOrEjTbdH2CNSCuLBd1b4ADEvbtig4Dp7NBYqnHFPiNjlqMCBlLFe
l+JtLIcuuPs9z2eIaEYyYvZXxZiNw/SUNhVfIoBMTiJJVcvT72Qb+9ZIqVxI
cS1gw/rcxeYubVHLIcgPXQAf8thEdpJ65ROUCUMkSN2Q4Mk5DKGzrwFEY25n
Bz0O5p0h+NBEThp01BOoZYLmzE6FQ2mxc7q5fpGVV7uUsT4ZhNzbnZEsKGaA
sUIDchUnHM5qaaLqu/dOJ+sSlNmwpp1lOfaC6ApVtbA3ZoqZAaPvFfiH4cZu
u1Qn3eXYuh23VLfPOMll5+yu/CKYeV+sqilVkwrXLrYuIp19PIbCJwZL//xt
JBMRmlrX2NamFknaTjtLoaHveAU1M8xYioxgymCfpNJCs70gC16+7k1nZFP8
ZYiA0H/XwSeSR/Q+jX1ObgPLMpVg7xKliiGEzplo/Ey882SAwT3ZczZ1JHCp
Exag776h5p58jDmOPnYjmjULfbGhw7GjW9pkQ1mUnM3Y9JWKXF4/54k0UTC+
FmzW4ZcHJifTqg12btu9pEFSeIYiQR+CD4GJxppAV5WK9Kf07Exn/4nv1IfR
+jZApH1+Gop4YVDMRZtNawO1wEGKkGYROKbLxS7bRYt0keHkxLOZNSxIhqpE
LUBnP2QlY1NUkf2Mb/fuEphaqRrg00yUu0Uk8qFBVjTshWlsgwzg1sD8ml1p
614NmiJUVCwhSJOPTkF9srXPTUxgVZK+K2VgNSX5IXJwQ/rbewcSZJ72OoYa
AbEmsu8WVZtlR+FV1oFPxRabXxqVJSI0Jvmpo5iN99L7Mxk4v+13in5NLq1z
sWMJoOkZk2tORvRNf0KVHaS9nJeuO2VBpuIr6f0tW4t2dkYLdsBXFeOiQrxd
n8jTnaheG8kYs0DMBjK0C+9QrxlTyagM7G3MY7U1yGSHgnZkOegEGVPwmDzF
9NlV7g9rjYUKTC6d4sIOriXaG9NWp+ptpzFr6YOmbEJ22R+xoyImlYjJUXm2
OfkloKbe8fQE8NcuH3LySqDtMkXmNBl2WIlhokb0YMqxRqC7PMeEXXIw+adW
0jCfn1ekNalhxvudvmpsxP4QTTfdezPvw+YdiEbj0DdGkilC8sNOuG+tOMVa
JHb/CzSLvD74wEWegnYdVKc+m7GboDzx7r5AnQyKn+L18etGYs7JkEgZhG7D
VYAKHxo1P4ACcnATHF4aj1XhSCXE0gRdQnH07yz7jdNLpv9A5WnJ6D86tGA8
bzjcMHpiLrpgN9FEVZFdliVUuF33+REGWkT4rnydalm169522UddsQvnFyhW
qqU8QPci7J3eXxlFrVX2cRBPMmiK/mgthpTem8eGf++o81qr8cCKDETTLMMO
VoyLgYb0hFvm/p1Wmnfx2MCOiLvZrIzDJFuirQ5kxOKXKjFArRfa1Af4AWO6
sjFdk9ur2qbGoCcrS/OXE4hyVG7TLAbDfnLTMWpwRZu3uNqSrOiCRJa7FpBF
vCUExL7z4139MwAMo2dQd5OXDdH8nSAkogn1hVVtr+bmgVTO21YFaHc7rPoE
0UMQdh2oQGp1/Na0Zwmv8clMB7oxExMSfCYTtzIh5Ba8C/0ByJDXNMfiIxdN
Lqma6gPtbOIPnKO53VfD0nq7a5mkbSQsPDWLY8PaBL3ULaq6xrcFCR1/ifwq
XpBuyPU8Rw/7CI8z4HVtoixgALd1Tlu9/NvW6yDWF+tb7bwwiGE7GWflRF+/
tg4AvYVEtnX2AKImpG9dLR4hYLn0BkS82kNrY/greOE7vJNa3FacfysKqjiq
unUrYnjPWP7yaWzvYcjlkS9qbEp4gK0OyuOvdfWu5eKQDoaYkqql+xbVZk8m
qYogdaABdiqhVQgaKFuLIbuOKeCwHBNpNv3QgcUM3TH1YxeCyh3Xy+fZEDaq
HVDtddcxNPPVW5eVCm2aCCoXTNBgU6FAhtmXPUPQZ2oYAPoAGG2fZWQotuEL
aLM29vA7D0qVAvx7Q85mhRSZDMDmvTmotMFKAcIAv3LhtYxLArVmV00NTDWM
iBK6jqEW5xZDaky1CuotfASxuXRGgHXb3RFtGY4hDqFmNEy1y7AWXMAFRewb
XZLkMhcgB6Qddfan19kshS+YcwnH1QI9capIh6opoCJXaWTloI9jo5uc2Lo4
na8cCU5U8iy9tGOnF8F3w/gJj6Ru3+DSRECTtkkbGvsgNFGA6dJ3jDJrWmNI
NnAvOCUPCzkFclCZ/qs1CSUjWP0ETx77v6zwC6iJKFayHV6Ujm2rUenfJile
TBSMIwPMnhc6WFqZvxYs+KkRhQk0TeGO2eGgYXZdlxWfWwj0QnO3lP9Yi/im
00WXrPpql1EE7T2u9kI6Xr9Ns6SYnwlGmJXMv7MxjfFl4USjn6AtiYB/km2S
qh8/1jkhP085/2ZeW5ydZGcPY25OUmYYtq5oNE2Kj2sK3Mw7dfhyg4INym5d
+mhhCd5B5q41fLhIZMYj8stEqerq8rKHnl8e1xIAHM/4E7X6+Pxl9FR22L7q
pRLG4ysbruTrjzHph0/H2Dsa7HQLfigE/kq9nYIGPOoFOw070pZUpIrpaIX+
cGEp2B8gJfpP8S2Rb9QKrZ9vhvurtR41rPAnT4PKZpHfiF4FJwpGMJ9XAH01
tcEQCWDstBhGwHrdq3cW40lpk4jum6mg5ecDzV0grWK2k7Fu2Juqq9EczgY5
FLHPp4zGFUj4ggl6psS7vCpTnJ4oUSJELBafQvv1Jt7lFEcguGXp66vdVseU
zzSAPvxkZu1Li+ffc1Rtfsv1ZoKyLRuVdg2FgcvkI0rsZ7IlF69R42sLYVm4
Vk2xIDs35bQyvNSfshARDmD541Ft6fAZ7AE9hQatnHzWBVpkLkLMTmI5D1Lf
oTDgkdqPiG4uhv9W3iuwvColDZNAn05xUeLpdc5D3nJ569YIoFLO15V1F+hA
lerJwqLKlXCHlFDDAvoRGSaJnvS4e/JPADPE/VNCpzLGJ1b3XyV20s6d3aQI
SnqlWwnzcQVnUv1gO83AEANyhop8QJD7GU2yOjEtTCuwd2bUX8GJkKmAhA4v
5rvw+cr6CF5N7dsypsCghM/s36WYP/xKPWdgMwF/BTsNCOtMmdVeaNdsjMNU
TYHC++gca16//pqzujg2Xi8xh95E8Uk7xShfrh5D1K1g5d4eqM+tZFq49WLv
OfvbwPaMDgmZOBXjTZT8bnvb8qowNUU1lnpvw5xFPSrVvV3Z3hxIGBqqNfOO
+Q1I3M9TpsHKtxUdafv9/ONwcvAYSM/UBxtd0ezSlH/axjaqkoG1VxzJDuuT
Pk0uBsGMa7Tf28cPSpv8wriAffYNEJtQsCfhhy2ENaHYRCO2uEDp57o8LWGq
ZvnucKwWOiaMjZFwCqMbtVv63rlBRDKJRQ523+pnq49GAtvjvzoESzi2xuFC
tYMP8U5HxMRHTR96TiHTim3l28TVjBXhjgVlQHgehv6T1y69UHPEKUGN0SXg
ymOnugd8FLiLVJp6SVDZzbe+Uq7WhZQ2KkESt6AnTgHVb/5Uc3S7HdxviwQG
18EwVMcqAukyE3hnPEVO7uZ3TI95oxjD3BVvse/+GK5N12c1Vc8ZlT1kFNF2
h0lgGP5jkKjTVhSm+Ic0BD6QomX6DkDUnqt82XIkDbhY3vs3xK839rgTJfkz
Buru1gkcbdGIr8ffx2NyLvqQAXb4lMHyji+1BxKGHC1K8uXyxoECej+gEx9F
FG/G1Ua+E32aaz7v/6dM8vBKTCQTEOlftyddpYLttU/VFsjRoPXeXOfYjDyC
vbRzNf6Pn7KGJgsj3jJdFfX6Z4VjSVFB82AITXAcA00PyCdN2BaAWsgOAZPc
ZLHlFbnzJjtSgyJLj8h0kD45yfcR3JYjyCSkeUj9m8TMD/Abz8Itj3cJkRbZ
dLrYNvTMt8Zs36mmNpVFOu6YrYxlxp5HPliZx04NK6rRFimCF5YZSTcZ3gp4
BsHpZhIaGK11SwgkXuILernjRniuVlfzkbBei0Eo0ghqOivBxKkcLQAvHcP2
AZyvmpfrzJi47C5PBYW7yDKvQIQyz7Ya7Me/ushUZEVrB5X0oqSbwj3yFP3b
M8kCrdhBU8IadGwAC9JwrTXIijSvNu4BspBEECynDl0R52TCJZ5zS+Aw6nWN
tbhCwV8iXMShRAFidKXY/a+oNJ7UORLO7uXWIsfPrmmDPShl5XfBsmje4A/X
2U79x4E64yJxpn37nnGHGFKB0nVIbSNnN1OGAsJmxyFFXe7EJrS1W2WRNou2
FT65jnSxCMGHAFDLnrPl/1lVII1mGMGiJub4JCmOBiQ/W+C03crf1umg5WKV
GHOAOcR3iIUjG6NOk321sULH/UZkB9//ZnHYFLpz5zrkLps7N4mChW7FuAk+
f2p1bINxdhm0ibFIJm/I7a+xjilJPJ3jO3bHS8mmTVV+7wvDtbB6jXLTrMAi
8bB1ckt+6JdDuV5/rjokYoJRGslMG9Amqzkopbe3B66mGBaZk83bCb5wE3Mi
E+ifBXc3bEU1wqRJGXbWPQ47CQHfjthacQNH1lkEApvd/zLz84AEesB0qyRy
SUa+jIe45uxwl3KaE7V8fyWkDc6UyIxIIcuaTXr9JW+XjaqA7tl7usKW9aSC
kn1Yq+DyTXU1Wej1zwhNMBuFjCRlL21gJPW1JF0WWyiP/kJvTzQUL/2sG7fS
rt3RE1ZKogxrVj4YLRGkMnTqFdpYbeRePQksuxbBIIn+lHBVYi9plyTqmtIy
ygPld47HIGOVt9aOkFh0iZJouYkv68j4T8FI9D8cx3r9E7dvNH7crsZPvyqz
arFrMLRLugKK3VwX/xAsxNbwpTm0Z8xefBt3xztkngzDHVY7Peuf23jjZMlz
1070XrEXk4kE+/0adHMnkzsXMJqBT+9/NYSFyVgED+oXLfvg3WS09jiNnYWj
c57tC3A7ODYWuzFkkaZ0znjVTU6TkdaRk+riB6NE9QQX7Ebxqm86sZtnQBp3
0tQ/sqSITF/nWuln3TqepQjDLb68RFhB66yvVgNDkbEDct7LdeVI0Ccb1dAx
s/oqv5jZHygNnxvsbNod8wjV/krLzmGN58WJqQ6giFpMBFdqs45YC7Wt3VOC
oEEiCHavfJ/ySHmE361C4/8lvWD7WgLQ69ZERpbn7fayuM3snkO7GnxOd+GK
YTInpphfHKRxl201aWOSwV5feRVdwNtYfGWSOMYP28K+g71bPAQnUCRf1Va3
javhYiB8YowxHr7uvCa4yN0NMjiqp9ANRZ1D3eb2yXlR29ZyBBAKowtEeCAB
lzmzVRy2XQ1vzv/Xsfjw+wmTb8Xt+WNcqZ1mLrOs7CkaVCpNkCT3CU9PFZQy
2Vut5bJuYkBX/EIsUSAWo9D18+AUa7Vc08417SGou3r8LJQHdUlgmDbrOoIR
pax7i3Ufvkp4FNUYDFBGVGy8hJ4nVimVlw1/1XJxtWxwfzw4H+kkK7taeYRz
/bZRKnZuFeHSKssnbQd3qwu1fVcH4Q+snR2Ry1NpdXUAo3jQ1zfcJnOfrLST
yZtz1JkhEe2CONxUP6jyKLiMwyHySwGCdrQsvzSfRps3THMYAsLazoAjDhVK
QR1xVvj5GRR6dX8XEFxKkSRc8S3V6dxTMhCmyq62qf9LkfifdRoOMnZTvnsM
X7AOn3O70amEMzb/pcT0zEKRBJsNN4d28TS4jfefrNafEgFOFsGsjBbiSF+1
PKQr7isV+xA1oJEodcX8m1iUUhgcD22wVErUqU1Ik7Qo07+sfb48ajem65/t
Z3IvCS08HuDSV3phBlyXQj6eIujWr+eEFz/pn3Vjd8VV6l8+0SN1Jbmk8F/0
I8HR5tY2UDB2aS+5pgAUPLqx7HEEkgvkZtV5fwXfI/YPMboLTSOCY3/G0VPk
GD9234Lp771Ex5ayF28+j5penzoM0sNK3/88uelisAsHt5DG8Al0zBbvv059
QxK/TV/l6ahyE5qzj7pLCzPKbG7YXvs0v3qyR06nUW5rGetLS3iCbAc5/mYD
l65Gg3PQIIEmmSBYAcmce+vkO/srSYurKvJi8QANKkNO2ySJLx5bK0jECr/p
OdrvSHsLFDLS20xGmLOZf0ouwN//FVEO0Xs8pyvNz9cYWwMp4FfrpAWK85uY
Qi7wzU48laVfJB166FPged7Ppyg27FgviKWQlBqM9/1nGpKAza80iqoJZU9f
6RPitpExB6/IggUEPjKP0PJSIpJXdytaQThEMtN0DO7wln9W+wwZfQfsq22p
C5oQHBECyEZz5+EyBXtxuDzJz9ruILfUssIN6q6lVrRewH5VfdBrOdS3S7xX
QKtmnmcRrxItgq/8OcHZJVxCzQNL3YcHGBiatF7UGRmcEagBaU4MvKSQa3gf
7/wvfAr3sWB7vd3KSZ3+qTYw8LTFXdUOGKHdjk3wedxhQb+Dr35Vl/ht3KIt
ZntfsIS+YdRMutjh9GVEbl68F9CPufm9YCgql1OGCxh/8OWLUYQH2irE4Y22
39IE1uYkHWU5k0bck2GwHXWtqBnfXvkfvpN/tldjnOzes3+QVNZeT2cY8HkR
ZV6/u8Mtz6ZxUA6Jts79iiUgGdtqsCSiUL+4UtkhFiVgQ/pKPUXR1XpWt+UH
DdFjvDBOxwVkXRfvc+5n0Lr74Pj3ZqB+ruADZVPcpCb7jDK7nixu4zZT6kQA
pawc+x+Dqe55rBlSLEF2wHznjd/npoTeTu0tQmrlazGuIhmwHKOa6Ufvw4kE
Q+RiPOJqMqURVc09ivWqY2Og/4g77HoA9wUpS2xM8STkjCQ9cvxSV3amGQeD
sn34UzikFpBwWUUK4O7y0iHQ76O5BEyWdKL98Jnu5HWZvE41cNk05y7ZuDGb
WxSpmw0tWppj9UmM+nh/LglmqRlyffajUIU7E0e3bivc0qTndZe7ZOD8eZuk
9jGj0Zrit+a7uIKACE5atapm9jqL9/B+0oVm8q5nTkGLY3Jx68qj6Fh+5UXt
eZGG9bkhqg5JuFkCjn+aJUX/Q3tUri75fgSMttntAvcZi9ZrYgza0JpU4csy
h/Wbl+jYxGFaoBftzgcp2QPpCK+rd7+mhKknusOx4PxB2axQwuIMQ3eYvYgT
VGHcNoLla4lsAVMxRGoeatMnGIJTs3uIcE/8f+6sxAX+WDt3twxLdz3koF1t
3sqmTlxYs6L3jszBlGdxo9Ijv18O4i4cMKBdZS0e5CcjPeg55MsuumR6Ksu9
xqFIxbPFyiDOYBY8X2DVvTPKdZyCX9hLjV1m7GSqCdOoalYsnDDa68CGpryz
G3DSCO7PogLgT8TW3/zaji1Zc8GgW9UuItTwA5i8WlVJvUrGRRFxjml00Bqs
MUyXNOGHYcDNvq/ANL1xg+9ABpjTwyu4osAcR9pT2iZdq6IbIITWrw73CLbx
ySwSdwdPEgLnuTvMRu48JQR8awB44AxlqS8ewQEwZErMyrJ1qH+5f6WSfDzR
IqjrBxPsHt5ayTyXSs4VEOyh0qqpM/RpBM30LRJU/nQ5OsOFbSmMIVGz19Wg
MyMEsISYMJvlTXwEraSsBI14ibiHNzpy1IhIpu3JjIi+rRKY4U7NHjypw+6b
OAxpFNjJ9u9CTCRJ6I6U5s6mihrD14h3xmv1LQRvOGFFc8y+8u491tDwcMQd
UNfpKiU0QJPAF4wBv412Eo28Wl+TN+YevMUdblehpmNQZHEaWnz5LvyWp4GY
oTkpPInWuqI9AEz6/N8J16pW7RGGBQpl5KGy525xo/qdGnciaAmossvE127t
KrEaLx/zep1tFKR6+ASCG/TgyKWXYF4mCqfD4Zekua08BgKHxUSkZrZoXeRY
nzT1n6yQtqNwtKaAVT3q2jemplfNpSsCIKxh2AdHGRChIq+5nwJu/rV8UC9/
wwt9zCs3NAkRGVUiO2uxz7b+MVVW5hRr3YEEJOF8vbk/cxrMNRT4+b8k4HaZ
tyj8g3R5gEBFKiRe2MRbK75tE3CP0bju+lUY/lES6oLdhy8wvZKU3AvFlnmQ
QVm7Ix5ySyVrHQ+kX966lF/LQenOofZeRVAnEsg157bBiSQHN9ne+ogQwv3i
aw2YFGbrys2EV+Cw0NtXkgP/OHuGDiFmeFA7S9EkZrijKE0NkE9f8HxHeBew
6nBQ2ZuhOMtXl6VAPAGaEucazQM4K4R0IzYUdmqhSh4H99A2T0aHizVLkKnX
wRjE7iwUvAyd3JPCd1AWKdE8s9JQiBU3xI5S/gYb9H1dRe7kjj/HVd/yqRZX
L3hPByyglUMe2PwcUV+OrzPb85yaDMqlev+7HGEIXMyJlqGZIHNUgBjPaD5E
rU4fszH7TMo9MQkcNKVtu/ki4Zc58pn3zPQQXSHLFdQX5N6knQIT5iyLRtGm
dDPOHJruOT8661RFvllKVJ/KiqN47vl3x4YLhYRgdOIj9lFH2N3cNv0FiQUR
bJsvRrEhR4TkyTaBTzLpGtZo9mrI5nmdAV+zoAogHB3o20aeDWOSfqssPXu2
FUvs3PBaWI/yk8QWOiXUBDHk/J5rbLGQ59mCvcLRnfI71bq9oxCEyM2QE1hH
wk1qGyRwWpe1Q3II1yErFmp7bE0Ww9Vjz4qZBbrpWCbBZH+nk/7q7q/XSWb5
59AnfUxjwWv7PGq4aroJc2kOES9N9Egv3BP+vvVH8WwjZhawB+jyyU2DYoM7
Edcb8q4wo0jEePb1xdMWtMnF84Dg1byB9LaCsjmD5PKtEV+NXV2e9Jp1iWqf
ilY/L9hTp8hbaidXE6n7JMnJHOW9gd/OeHuup5oRfxgZ/DZDg1/Ze0aWaBH5
i1c5V2SygH0uYL7q5zTxHDZFk+RUs5Mm0/aX1ssTk4zqanFdmjJxJbbW4z1h
JrY7iSXks4sM/Y5cYzIKk8qZjgBn20fxUihCin2NAIGUfZxKStpOWJnNqX3S
nxxr3X3SGOrbYiZv0F0bJbtT1TumHxPJDIMOmREwUa4oY4P/iGFzGqjzOdnF
3BTcN4LjXiIBE2pFpd1DbCYurpPhbo2aCe0qfm9DPybldSbjDonjdudTLuWs
8FgKaLAm6y6K6YYV0NJLPfzKl60IJWI0wb8wnpz5MuZ+Ni0AIZ8jX1RCtm5l
+DTjqVwpOsec/+uxqe8/caeiYYBONflBWELnJqap1Ibwz4HKREf2r4eyMIds
sJdRx2DqLW8S/TDp1fkQYXSdATYtGdVt9a2rTUHue7bNEi8YCNXI7DZSMwhi
bCrhJVlcJ3NZkQPu6gEmRhz01P+HHvmvYPZvJp6z6zBxPTXgi81b0fYwax2b
u1kKUJovQlxmol03aUucEZ3r/3fnnHnUZwc0RkEAv2l6RYAkPcNBgUf0/vOC
It7hGbZScF4SPPa8+YLzQlRo7GB0suOWuQFEUawOgr3gSL7QIgxQBgoPQWHE
2CUFD76fWA2GQINNSZ1lUiGjwBeOje5ArISXulsWoG0Q/C9nrPB+GISSGocL
h/QMGME8WpFNbbk/A1K2Qvwig86nADrtHGQ9MLNoBaewlyl+mBzV90f0LTJN
/rveVveysWfmNcDYuctewP1vUkpdfwLYfQQzVE7qvSYQy89kxAL2AMxq3Jev
WmPAemcfxlpbd54vacNEdawA0L6isauR0JDs2gXe52hNtaL4wDfDehP0RsCW
fPZT/9A/J6TNVX8AzoV21D0PVYQKCrcUez+fB3NdY5NOvOe9551ACwq5boMt
3DdaRfCIoccH3oJgnOLKSuOHqjvIWhcmswwQ1KXFXhRxjkt5k2gtjgsaVYFr
H/oPuyrbbVz9Dfxun32YnZLTeIbM4nQ05a4eslFnR0MZ8jbcs7rOs02cMGLg
eyKMxK2DNDNcgKQ9fdN3iYWIyd4L2Uz0KQYxuWPBiQvWr4cr3UtmdQtS8/zp
XRbznhi4zitzrF46bZPd67pOzXeJ/e7Yxcl6faJE5relqkRYtoDBwUqfcE8N
UCuLJ23csA6ss2tZoZuSZE5li4HBrDCO+pHP4VF5VrsToqoCv9/zUY8jRXmX
xhu35kQGL+6JOhlfUCTJ5VTWE0n7V3Dqfnx8pmvSUL0CBFyjLCoyVq3NUdrK
nwbUIvHXGwd9hFBRkg6cAqbCVMOi4DaJUb5pCxhO4UQ0p4C3VAKcgaQvI4ol
nW/Yu+El2xXvQ8UH3KN2JuY1ZmIclYayMfAxufGwZszKtO9dlhh6Sp1gf4TN
si7fpBcVsLD4ZMZToFl5WFpPA1CJ1IF+zprxhRT3tqZ3EdHh/jRhxqzKAZFN
z4YGfhOvfvNVEmQCIEZ7VJmS4/9XaVjw+OWJ857WeGQQ0R6GZWXwkhtUimFu
BgGQeuZBNKmM2eE8LjItHraE7DPwzD5R3fKhRQ7I5aUWoGu02LHkl3cP7L8N
U3iPx0PDKE0uq8GCUAdyQCs0o0nYi3NJa4Yi7/M/ktzlATSpRx+rTbkapAB7
ASnRcSz8fzuQDLZK8UBVxPriTpa06tkyzCedeL1SvCTwFh/t277IQe9ov90n
1qoWXzabxT17YLvgzOlV6fu74sGyydCYhvEMCPsSAYN6+H4o3oWv7FkeRJWd
Eu1wTApri/9l/vW7v5wc5wZNEMwJOwZC20e8B6JoZjhV9F/u5CgNyLOu3W9Y
1DS14EWwZvOhhiSvbr55SPKwSHS28KwCVXMecOP30nYk7FFvaYyX9us95vPG
jqyZC3UDt6RESg9DrEUmusUNlwkvdcfDRwDqEdKYti08PkMDBGm6ZtTuVClI
jTzIEK/AjTlVux1NzUNNg9r4Tx//yfv9aSlxysb7mwt0mNLGZ+oA6pkv3vdr
epOZvXLsEUQi/T0w22hsNaWZy/42v4tgcQEMF+JW9CHOygZ8S0uUmbwKZd8u
anj7jpC8QF5bUrwE26N7kh5JBP0wBTkDFo+bEuqq1S+WmLi2DyFADVj94t/y
O0afqLiVsIOXmvfOoTQUINfYbXiGjwNDFKwX309EImuhRREEMlU9BRLW73Y8
UuwrmZ/fUIMNlHnS2/B7arJ+eJAyRauvie324S3EWUcmzWx27TQSXiALFLTx
okH7mA4q8KV9jvyNKqG8rUV/4hFwZ4OGx5hembdlDqfkd3Le/LuBpr5js38Z
HPyhoPP4BS8FOcC9Bibw0ZuCH+NAK2+bsCFKfuBfpIdow/Z+Gsk5JZMNxb+K
gEUcOBqIxohQhqwZFsavi59VdiyCJj9OXue2MT75Yt3P20IAlRxCtOx2ZVqK
hEcLB+h8vw9eFg53XAS+f1SwZzsO+YANBKjWn/3P+yS5QsMCHu3Kv/GNrfLA
GdMNakSP9rsZoJr/0F0EDy2FQHGsE84yHMmy45GsbfINV0uuHlMEuF85WYUV
4VAS62kpfEqabQA+HIAa9Dl9mcJpAZC6HOjtIBfMqTNckPLQRGG4LkD9gWGb
ELGalDz1oraqcu5IRuhn4z/LqxF0zUMw25hMniziImcLio1srMxvzKk/4cGe
J7JYg+DkT1k0Nyc0t8Evlfe67V7qLbdmAHf7TqPGHYxTSHiLJUT7UuYlY+LC
FKIMWrhrlmZAYxcUGhhrn1TtKJ6g3YX1LU+k09H3yvNL24ha9JYvO18UuxAU
YXlC0PoSR4LQA/noSkubKNiSEaG5Ak+SOt+8xaWeH+hlAZ6g/K5+2RPpDInS
1jVcP2gX+Bc2WWBqlGQAuBxxDV+Br193Lf3O+625y6a8piNjuWA97+GiM+Vt
XE3e5x2XfbwH1W1LgoeczGDc9O/5q4ZNxbFnPwEP5BoYhtLIVYB2keq6z074
fB6fxU0dFSx+XapbtRddoBg9fmc+Cblkk/RcEhkIfN7LgU6D1Yim0kTUjxj5
ii9kyfvo/LCHR2YbXchAInxhBXksVOXYUXKCp7Fd0XTcSWBnTxxgur+UvDyD
atitafwj0YSnkr+cTYOL+wegdDKGT3aclq9EMf10If8EQ5/+zYQYWmnkyFoA
hM0u6C10p3IwQiGWHR/+p6tVs9gLrze98oQDp0WvyYoeC00eoc0afwYyUhKy
+fv99OgU9zKizEzmGiLDw1R0WVREdjfaoD7/mdeAFs6Xi6xyc5feTsbArT18
ixynVjZvZ4NBBdG7IhmMXJmyJbiLn2g4CHV2v7TQOtks5KLLrpj5XdhxtMrk
qbYzKikgP/VjNLMxHgE6eKVNcvW11NcLjTO2FW6xRCeCOv7Cwh/zSEZPGAsi
x4m0fgb7Clo4Xtbcynm5CUrJLe7ol/8=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qR5W8/1q9d2gU3B8IKzK6DLErCzyMXeMJDxgSVTVW/9YjK3xKJ2nIBihxBVlmPGAn827Q9lCyUB8i9mN3zI6G99MGcIr0VqKfcoJSGL4C3gjs7XoRmQ36s99wE68Rl5iR1UonYkQHV/IG6dYmU8uLGl1oDfKIcOcsSDABiMvjtfLc6vNBirxIPa1yFuKdZPjuTK7BxDeYzhBUDKxXnz8TAhliq9lUbFt3W2ljj30erq4aPcHEj8fPrPANFncjwa7PUyUlZymciqA/bcfNzdeCJ1ujVM1XdvogYNJswxCGtyTghudY/jxXDx+siiat8SzDNfhpm9yg0WIf9w55omE3X0ccspP7BkKEnZ817KCgxtovy6IkBETHh4HuVmakDtqYTGEPnWf93pD8lXeYMNVN9S7VRIeprniS8vWQo37PLzUhNNlg8T+kJjcy95/oTmiPhPZ3fmzQE7p9LL7qTebBneOsGQt0R9QTuoMLLOhuTHZUT0AVUx9d4cMkR19Jvzai63A/50h+gw59MadWyjyOSIM9gHth+u5d5A3dTOzTZmGxE5U9ByKJJQu1bMZ7sBVenw/ePzfxhwhbVlMYRnAIKD4EK2TohigCYSbDVMEbdQWGDSZDmxTcR21eMm3hjxNX56b2z6NAozzBRvLeDcPVB9R3IRRs9cpmZZjGIXGtrnXDDh5cYpSnmDlPysg3aekJqyTpayXgk36f9BYCzNuecDxj+hOrqm12zzLvfHCP82qtd6XhDaGKEiNoBpaaoJJCkBRGDkxpLLpIRDpmIfOw20"
`endif