// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wE8KD3f5hPkVb0AlLK4emqp25PF0AGme/S96PBBXv6hZEniy1Aa2IljiVO36
WHGEOuUaeq2uZ/AQtY5+uSggZwLHMcK3cLd3oMqIWb91DP1UFdeIjVyarvtC
Hb9IBrH0b3insTcNaGua7lJAT1DBcSpEaJ6NZNiculRwle8QjZajNtIoTd/p
+EnSwUs4YR65qSvZkAHfnqAhcCxiJmgDyDk3/1oI9C5TS+J/B+LokfyNpIUU
7gEWJDBpmg+LLYU0BnzdJo0SX3rDm5vBWU3TTkjlHXVTNbrXGR0ranQSFUlB
weWv/kD1r3JH3FdetJJLLeFLxd0M9W7VTRraKxv+rQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Kf2uN6sDTGelzFe08DPM2CmqAqUX+dNMWTSOxSJRVGC9n7l9tONi26pzyVmA
HwIXni8OVP40ew1LSPsfbTot2Zvp/Z6NwBK8AUPPteurIDnvHbtckpVFgEnV
ihCOQuqIb+PlOcoUFRDa7wZ3eNGxJVUN+nYWk6TsQkv6AJlbIfbP5WPFcytj
3cQamVrc87RBXUSij1NkOnlKgMxw7/5YSEvwH37sFFl8aa6doVzH8x3MvONo
/oCcsQNCb0ldZDlsFn+6+C+nFxXSDtKuMK0lQDddfQ1yTRKvmtUKP88k98sd
xXABDak3C3FdhhCAb7ocu7w8f3qZQS1zUCPWypW9SQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p9crBakPb/gz7kRk0H9KyNRIxdWNj+VsO0iKOp9vpQMuZedwnbmikjnGMbg7
WzvZoKmwJ61AmnvbXqxT/4pakCMaciHCnXnPaeeoOm9Mbn/pbtci1aWTPSYW
AziUzxH5P7iGnRpb0I6O4NoRCiuuHHvnsqzZiN24z+xchFGGRbjABIAZMydR
ZfZmpZjyMKmIu6MfPE9ycghgtVe02Skk6XXEF+XURaX9aNWJDqI3Usfg7/V3
aPhZG6KBqbdnptzPMg5F+nMoI/RDvJcYon3Bug9CWt+oUKIVFC1U6n/2JS6i
9ersEru7hxKd8sxga6Pic+qBc93d52laqOvy9OowUA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KUtveZesvd0NKk9SA4gQI7BdUJIYabdBUM20QYCMbyBmEn9RQG0+jr/RePRg
IyZ+vXz2JxV08p/eL1kHAT7fN3pGIlnSdK7gPYDmer1Lh6QzFUsu4mdRVrUT
JQe7iKoIUjTT/CJvVuU3XfR7UdDDF/u1LTknsnJW8TDvj/j/WC2KaHZvTLSV
eB+o+gycdNpcBPEcNaQjLg+NlMbY9Aq+cBHWngCradrW5uzzIrvrtt187yTo
FA3dl7ONopl+6ftRuR1kTw/Nk3/BXe8XDuH68lnft39kL7UCpXDj/M6QzxGk
WL25esNbRVNgMhrhjSynqhci5+l2MoySj+1Yw845og==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rK2oZLyjhPKCH22z/ZR6ixjwzjin1/UntvHyQ4yLZU2F750f3Do72UILH8hP
Re5+IbM6Tytioxe7/wRw1RYIkL/gcagYtjHEs163Zln0ObYd/d344SIuoXRF
CvFyIenctkuDSVALawcxhDsYOca8d0rlk6yqQa1HCk4sEeaqLL4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cchbq7L5yHg3YOaA/843QDHeJUguWAo2/nrz7wi5ybhMUBWlDffFt8ZOdJZP
bsRk+0zRhr9mXd1Gl17J5IT83d03gV2fhogwdqrzrAKv1Y09bS3BBriqRDSy
BUTL6rKr2ajPMUTdramMfi9eKu0dxtVuG+gXHrId0mFZnhq35RmZGA2iYiQo
YP/ziTNEUfi1j4xL9ixMlt929BkcAxVewxeyq6aOqNbxnkHIIjWPY7BLrIHB
t52iWLNdNDSl+EkdMXJ/dGBgBvoGctRDRgZ05JJ5Dk+hXBn8DlHQ+TeYfcOn
wV40OsSZsXE/HGC9ymzRjUukV3xjj5xCIOSOaReQqoA+zxlrR4RTkTV7Imzt
V6jGWr/zwvh51b7FvIjiyPAra6ebmq2Lpvd/Lol2ZAT4kSQb4WWIJjaZFG45
VXdlONwuRUzskTtKnc29Is+mLuIUdesB9M1QKp7HJ6rsAYftNqw61JiKn2Zp
Ui7EspkfV1uoio0wpp5HDV54ZmGJP5vx


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hGl4FORQE8uGLkmCycrtvL3sbUq5i5+a9Ygm9DF1EBQQB+ikc52Cn7l5tZQc
ShNup1XBEB2zxgKxpGpMH6xr8RXe/Uu8DkRoKRI7/D8O4MzZpN7t2r9NJwny
YQUpTWQriLouekFv2kvGO2uZyt/1pR2TOjyd238u59vLgxSHLpc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AIYf2TfzHWmZWUwOaefJ4DdaD/7sbLbvkfPExpCyxaGB5ECAeso1viL09FdM
l3RLozuVDa4RDNKDa/o/G88U42L7LcMjQKGpkQv3fbVwWnqF/J08W82hakmJ
Ht7YitDeA0eOVYk0FmiVhR2c2XbRDGcJ2CiDo8dUGIOVMMmOz1s=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 29504)
`pragma protect data_block
XOpKddC88ZTVU9+wC4TV3f/B9NjS6xKvI7KjlHmtbLdicoi99kqMCZBKcXCE
M09Mjj7Q5VEAkGH67TWWizYNmnTEBvGhN7pkU7RbmPtYukwKjaWzM7laIJGb
KdCvhhWB9EeMkAOz3wptZFIpKpl8rIY66+l9Kjk3Fdx7vyJuwILDu1e5i8W7
gGikY2sG0UVe0i1ogwJ6vmSLJUCTwM4OS+ol89OCgk+XNauGXn//8Q/7jCDV
4CQCNmiSIkK3jbgqmqc7leB/pN4tmYIIn43BJ7AONO4TsZxYOdCDbTr+0ICY
nICTkz3VAgQui8QENPIZvjlY+tT5/1XlJCmRXpqUjbBA7qcbuT4iuXRcT8kj
JM5yRlWjMnZThqzIQE+L5EQWAadn6CBvFbM0AjrdZpdopVVReiWPTpvebGsp
wKJ5ANKp38HtP8gDQIzM0q/QtnGzEYX8dM2V6l/WpBD7ul3K6j4HjesVE4ub
j+95fixggJPZtgr9sSdlF0PoaOUj3Oyj9FyiYlunqc264CQ5irOcqQTiRz5T
kPBKAQg+LBZSsiQyYd6WHCqcepstqssKsDJWDqOxNdJ7gKvlfHvZ9MXKwu6D
PrPDxjZsteaV4fQhsVXBaqiv1peWFLS42rr48U+Qpi08VkSH2DhDqYuoC821
+HpH5UM0OWWPbIakdhey4ViBg1bctZsRsZ6ZjenYHCMSCEHw7fw45TRb8f5+
4RziRnRKdKpCs/4UdI0V2e9kfnoul5KaDEmjS1kret7JKqp1X6DyQgEUV/c5
5IteMpIQCqEwzJHnRDSHSdbrDMqZQACMlhQB9DNy4jWXIHki09yYAV2pwQtg
H0A1h/Hk0em1w3fR61+I0afTygz8rd6w18fNBz83zpT46JLTD6xW0JG9rdeY
Pcs2nM9dn5ew0Kno1EEVMTzlCFgXbJlMFJ/bKwid8wFh287I9t+5d3NDpR8I
VYvUcZYCRuKw0XAdBmnWQq2iilpFyQ9CUG6iaeeoiyTNG/HLGR7C0jnPynrg
6U725RiIDhpp70FzolH2Q5kJ8J9hndp7bQr4/bjgcDPRwFk19PKLNN+Xp8Fo
S8ELX3jtOZ/FAb1MHDHuqViTFrytNjef1ROFcLdxk12bpJ2f/s4C1X6BisUs
ievJ4SBFZDjtP4UDAC1KQf6PtBX2p6aKlYD5FzGc9oYVtUL/I94DrJMTTk6w
Jljy6edY6ktpSQDNOSVopjJMskxQUxtDQg1nkB5A8g6iXEfT9xzNAoThct9q
44a+8dBqk2ezmenUBQ/9h2ZGi5wd86MCJ86/Djn9Zto2BXZ/w+g5vyX9KrG1
McUpMmFKABzG7cyXt8Q0q1ro2UotQKG7q5ju6RnAJMTFM003pxBLlZTBpvHB
0pwhykPoXWaFcB1f/lJe1K6M6D9ia3XZDhKAzFF0frxcjTxGwKAwKJWzRPKw
16yn+aVfpH43UZ0ya7NgP4ekbtRIT6+xsc3uV8FdNp6SFVvCoBn5AztfaBa5
j70GP1kp2huuV25jaAUktI2wRvwwtahkmKs2AXxPKltsTSe57FnmgoCaDbkR
1cRCj7LDx7UYIxYsU1RPK7FliIMBWh3W88+ACV6Rx2eZKAeN41ZEpGYMMZij
sHsH39KVRVsszctw1kuD1lNME95Trr2fGB4/evn1AQ5IQpppBZ9naZADDwRr
BcCuh5TgN79cfca/+pr1UkyD2fKCqQIJjPQx2g8SwlmQEkpD3H9czlYWzfKB
gMqQNUcUS4P16ZcIXbLd1Tk0UQaJUDpBR5l0jJZ5hVfLgBVpwZi+2TJTRQUZ
ImoD9ivU2c3D6e0mF2q5OPs7WTjPhaUwDb1WswOW3ItV4uuEcDU1E7yjznxp
0vi8rsar+SZX51JpqoD2t4z6GznkbSQUFzZ4DCWyncTKPVAdi8Uaed+OIDOs
QD64Iok+/KP+QqOWxWlsnuTbG0RgoKppzr3bjnOr+BlxorlT+96wIaF5gG3L
u/mXS9aBn3gKAg0fPi7382X95zgmV3WysATS/lVlF9Q8ShkRDgp/sdjUBuCg
5gG+/rS44rgsIcmGFAVPfBmMmc1qMU33DCYjM8XPG34UtVls9d9r9+oxBK5W
4+9naOSqyW5helutHXgtsQQnkpR2EJPQaOY8iuMriaOi+qJSU3OqVJgYQUjM
kUKThnYidfiXxehFcdI+7vXPJ5v6gSV4MyjV5sZKEyr3QmXst1ujU0e+kdHp
SxFbOPUtQkD3CK6j2CzsgLFxI2llmcFbTZFR05pEirNty6dg8ZZiqaab/VK9
DBnAyXocTSa/VGCLvZxMsWjvvDbGK6foe4pHqlBRFzK1UT3VJ9E2oBd7Kzuj
re0B4hqvHdSyfST3D+AyJ7drfL2EF3OtjRv5YUmVRUne7C3MCYEUKbcGNzBS
6SmVitGFYTV4SplPXfZiukXBCcnv02tTBWnkW1h5LWqm+z6Z8DZdfHkkF6xj
0FH2AXx7RC/6p+KXwCUt6LBgakyx8c8cs+hcoI0r8zhlosvi8m1evwBZz4cK
Uk3fR9QnGadbKS7NqHdVI6N90U/8uWHQ5jRxeIQCCwYurfJHVqTPKWSJbDr1
6yVpkos042Nh/DUUf8U/WiKftdKKlxanooMyhPQU3L9msAELmNHIpnpN/6xD
oAh/cuklNOCvWESTnWLNGPue80fNLmhNsj/FCbETPskko2Le71J4eHgy+Fsx
dzBFtnHWF5qYFIF/g2C4y+Q4C3WdFefPjaL0MafzYoUSEs+AIhk/PIakFpSp
72kBXu+aUC0MiXQY3AaUlt2PjFqym68BwYKBQ4NBeKNZ6TwIR15iSuvwJNxo
gfVHjkmPHYOCYuamwBXyQ5vCKowkTXRj0fJdPrv+x5Aga5uBREAQbrDNtKQx
ZQSF6xZaQaph5c321revBOGkfgyi4pnw/KsG0Cdhb2cDfhbSJcmRd4ozVnVJ
tCpBY+/iQZsqicW1VZR7lpWCda3cxK6/jp9aj24NkTBvUbNPuSvcoG3Cv+B+
keHMFfP2J2mGsp59ycPyixS8mRzAH9EkwqAOVPDhLtZtebiO+MV4Jq2EhXWf
q3icYoWgZ/TT6wRZ0apmip6he0ZxBIgz6v+AjkDlr+VwZuh7PVE3apdnejRT
3U+2CUzZNYuDN9Bx/n39OcZS3xk9nRIN7pEg1r2TMmw+8GJI042G3HBN3YCp
NRybVZgvqn60e71mDpaoxp2H3JDjWrmy2axl8HDmHCzMdk3ubNURvNnChO12
y/HUI50+cyNXotgGhllqrNaiWtyVpdoko1uY7cL+LT/ZD4XDSe5MujhTmvXk
yu4jO2FfQzx2LhPz74IsEOX7pRi/maMQmmqFtZvvSB1h4O7J5Z0/e4BSG4kg
QNkRkZqU6B4CMdTF+abm+3H/l4O+rWYfuD5XxwfcQqzd5xY6uUGDmeeN8P6Y
i8PjtQjtOzQ+PZBHAH6+wH36tZbMWWx3LP1CgVE4Jm/4WIFLszt6jb+07LM8
OYVboZOZqTgSOJ5vGo0KP3P6/i7tXmdGluXuIxMskHmXO5cwh/s1wPMooo/b
ZUKuWb1REWVIFGBqSIzXiuCPQoP9DnYfRB+wHqdDD9H2fvp11cW0sr6RN6JR
S1W2/3EEEdyLQCMqZeSRIt7707cpMwMKU8y1k5mLNoGAySygeaJSHSAe8AWw
fhjeHpULMZpEyIYJ21rqGI9p/80zUWP+sb4T3Xxydbl27F2nC4s0NaIKdObn
r5FH6evfvaYGOqWPJiz8vmYSrHd/LOb/KFY1Dhmm+i34bRNK2eV99oxxilDO
ty7Q8GjgjkWpPfCDLI7mUOrjZxHFCRV8WSj5igT1ijDimBZgFsM//t9MfAE0
71Zzs9tM4TmH7lPfeAtbYks7ZLrtvqTIszsTVg2tshX3cLFC1ik2CG9RM/U2
aoH/En0JGmqc2X83oFsBzCJpZ34+NPrw88Nns6LcMP9u88gZMfm719B+VcaQ
R6ys5su+lmWE+vf6xhSBVtQFqTSotnxIax+ZBzIedMn7sJvPupzGGoUl7nfQ
v4zX4QIfhedxfQu4SDPVUsaieNbOXgTt3BGNZ1W/L3y/rr9+zELga5LDQurJ
1LqH2uNkiJR/ngBa24ZmI5gwmewHuqluwSBmyaMfXWJv9grBtZt+peCCNz+9
lke67t8lWQEfILN8kKswO1HSQNtGFVuXbmEJL8HPULBhfJcb9VwWri3EyBwj
6RtaJtEaxL+Uhozo0PX0xOgxFcmstsNEnP4IOzUJS8VcoH7L72kwyq9WbaDR
oiOGfYUTm26Q/6IScEdLGRBHruZ7+yZ1WCN3zGclV4w7Y+nKB+ZHs1o9uyAX
xNg4QOYtiyyvvYy+3zf/5j2H9SGa3kagHgqfzokAEL2CXFA4FKiUkGhVIRIM
gQOuDu652jKd07TH49nAPUyoDkEx9hgwSsl/oN/vbce4E3M2CrzCzhVEjMUN
qM1PDciN48mHwPFYGIE0zNBhSOFPweZDAm6cKeZ7SjmyiOkqJ5/olZyfzJhy
VMJ8sY3IGYfaiRbu4B9YDtp9UMn7YGNbU9W9KbQXDi1k9bwsuasIpADb8MUY
qbv++5FzNBocjJRFnFMzcxDqSx06VdUZkGAdAr9MIwJojpy1RUfj7yAJLCea
kVK4NIbJbCn0NPeWlJjMHpSe+nsyB38JTndc1XSWYxt8ki9DXnnOktNJ0DyN
2maUtvCuAlTfp25Bk040n+Qjg9AKT1IIv4FORCLvMoiGHJwaFPKA2fh5VnEt
5ILltJd/uuWQ8Eqe0Sed8KTzzjLztzZflHwustoZozxUg1HRZtFBFE5Nr7EX
vMpN1KsjKQm1PFkoLvTX2d4WeRKiJ3hUpD/pGUEMX0h//9q8KBr5lZxUTaLP
ZHJjbuZN95j36W++7lthVuvKcZwLhaZAvbs/+u2LMxzb8aS/ZYIMCCzh8a/L
Cqh6k/F2sgy2KaMkUY/cP9rp8bmuDy++Hn/YvUyZS2Mb1q048Hb24O0mzjBZ
jHhTt10Gxs4OgFoLb+TKYBrgLnlobvPWKG9YrD2lV2lhaDyJ78Oerytpjy2H
kTFZqfr5bkennBo1uRkJ/td/M8eRdnHGBhRfmOgVlXW04b1YxDpa2/KzVN1v
T7HLX/GrzpugQch6CEhLkuyIwwCves+nqQyQ8b8vH/mlfBhPkjkFv89jOuG9
YuQsA+IIQxuZRuFQmtImUbnFjP7bj3PE6YbGBNm0AgHxUU9ND969xjW5Od7z
+5uMkhkaHRk35dnsMr1cJicSFo85Lxs8FBkutYuH+2mBAj1gvFOG4cQyYaWQ
cLYDe+gvnKl4z4SgkPA15uT2zFcKXalDVjyDOQ/vlpp3VTH7SJzdDgzZQZjH
SOsSWcN+C6YZE2qlZMPEYjyfgcKnyc40plza4AWnK1SKqZJ7bENshjlR3A+v
lkyQs9b6pySYejrSF7uDcVHvAf0rSco3HUXLhMAdf2t076iawK/HscB7JVwf
O+1s6gAdITaBEbFQSGUKdpJPnvPn3+ZxaJF85SeB+np3zOKtuDxeZkjAd8T0
vdlVk/l4Ktqf/cM0ZuIhVHOX6LK5y4cgsCe0Ew4l3ezpMx7vo/pENwa4MdTn
GoMM7UtOnHy4XlpU+ih06HLHuFz/B6j2AvlrMkYdCKFAZk2XMPrQR3y/m7ga
82CdECxwbI6WTu/ELuQyYQS4m5NqlzQl38W3YV/Mosaes2Fir1H4OAZm2Pp/
m9tS01/iWfUomj+Ky/NlPQgpLXpV3thCMK3ee3Yt7wUD6oQ9UuOnOFrUcGRT
kzPknew7kkBnGGWbX800Qr1oGfQz4TUHwokkrCaeXsNwBtnaVaRHFjj8zpse
jXjgReSx0NP/v4ifwZ/LJcBC1etrZ0Tbr9TsFs9s04HaKIw14ljDSURcYPPd
9RTMqkf6QG/YvxvxfmLbCFhGriT3W7Cm86r0T29sjjtMijqShu8wZtvxyVki
s/MTDTE5Qom8Fn4rD/7ghNQP64vCNnK84hyu9fwYG4qKha3ccKVcbYP+YZSa
LW0+0uJdr/TBFNNiONiS3BFSC6kB9eN5rsyqicbp9UL79u/rvWP6nOMpYoAZ
+OqXlNDJBpBbkgsY9ByUriZoRa++K/5d9sM9NmvtwgpGS9kQi6zsMUF2Y3Bq
NHbhOlZ4p5Gs2/sia1dyXLtcXIeUYh3xOk/7s4ahFBojwQvnlK3iIW9e9Gfd
eP5oWrObqrkV6p0W8W+f/5/8UkaA+jppNqntEmD4WZyY/SsjSDkAAfzdgPmC
UbDXh0LonNRGXF5/cwHYOh/cb2JHjxxt56t1UZ0IJRVPZgFePSEm54sBiWBa
dEbjVoWtmXKVrh6SBQGOzttcPgSgGz/PEm8I4sTijZ57/m3A6XNuNjz15Jh2
dndq5WCa0tEFV8ZakaK167h4F5k21YFYpfJbWHYRt8OVBX5XuytICRD/zfk/
jiAtUaNCTMgXMGjX+V7oD9JZAAIgyhm2oz3Gm0cWkk0fx4XU67+mWNXXOC6v
phmaqPsmuqoQucu5XJarnx6EFzA5aOhxD1Aix6Y6wlus9RXoSkwOwtNcVLXp
Mt0JcbHUf3H8x/VqEcnWbf6SUF3eNcDv8XdR27FvRr4J38axeH7mxXx8qf8r
G3PF0yM+EYElyrtt3Da5VKdPtaQPt4PkONEyzNspQGEz+aQfhp3XtXg7u3ld
/rMtN8GYlhh99QXmDg/AvbwGfPSICfmS1qQEx+UaaDGuZaSHzpZMxjo6Htgc
x9kYVCejCL9XtK5XakYNBSvLQnXJlPrqYCWyJmv5spwKMpgTeJaT76eSOBJU
0f9tRwb6M6V6Vl1geZstF+14nqW4xJGkOFCa1xEEb2YxGNz2O7/sjWW9QtSb
SeGUPTGHyPzpnwlgpffQklHBC8mrTmc8s2cNZe5d+oWyYsgNNJ/PSY9YYqT5
vgfnza7oRaCo2j46Wtsd+vzy8ZFeX4C6OLeIAhv79HdDxGemeCdP++7ZdJx2
HST5XxquC/JenkC5o/8GvPUxS6NSkAlQIqgUZhRMhlkzgS+YhNvxx5wwhIw1
5EGYlnaqPR2/x/FjPQpGwRIRcN4gYKgF7Jd/e+XhAPLVyVRE+f7FzNpMojjY
aMwGJATaeARoyiQFZ8Jnyk5N4AS+oXXSYme+s0QwkeJzMu2iZeqVb6zd78mj
ufK6y324WwR0bizdSX+j2B4eFOFKkZWKoJFONmzuGKE9xdOCxDGXfXylq0hQ
JkiFVVnVGng4qpCITkxnNSgSd0HifVrY4E26ybFiKlRM9pvtMDooQDLHJ8rn
H1vjqo9IJOhxDv+zH9qF2ZDqXZLMFz8iCxjlYEGWqUWRHXFP2opA/33VfHfB
sj3q+YY/WHs/Pv1waQK5ZLOzYExZR7rcRtBWaOB8xAmmu3s/jRbny/LJnTVC
DkBfLoFtwGSUs46xRqY/KodW6KMo3JORxqtBSjroa4Pup1sd4Sl+yUo9XXnx
Iijtn8ChkuaZzW54Kc9PSJ6hrubejTYZG1qYEAXsqBomV0pExDDz2dOvUxFx
oVxW8yXaERGbe+dCH+GZDbtD5D8Z3Efg8M0h0kJ+bA42vEWlho3N7caDKgRW
R7gUXmJfqY4+rOMyNpLrH1QB+/KPva8UUuFo3AkBAV2GT0yDy/euZY0e3rlS
HCoFoiRDpSRHhlEMtHJymm/LUkZr+ojghXj7Q7TM3EDYiJApHFcgPndbaJoP
sUxC3LuwWywirbATGVGmjRQCCVCjuWDEugn/7ktUmaQ0oB9WjAJv90arv+K6
fDBuoS8xcGWwFnt3VgHKthucSMjZgVRwub7Bn+tzhP9wx5tO8B3UfKxlXbkC
HLYZiQHd6F20/RsdPtKLIN88lATHEHkm3Sp9ihYFTKax5cPZC55jwuvClaWq
mj6912TYpW/tFFyeI1/uyv7rUhkazHtM/INbVcxDi086219PWzeOCat6zdne
pafiy0fE8WHpabJ9u3IIhZbBe5IiuHobTS+S1zAtr5h+pPNPL6xOYis9aFiG
Ui7NjRa+80WuItkVYCroeMHRPcL2Fu+UWQYx6c9AuXdfVw9wsm8EFN0gIUZ3
p80IDyYJ6MvZFk2wcy4T00dd/AmgOe7rR/sYM0EEJVcShR7IXul0hfOb+80t
Lwl+Y0g5vIV4ONpDizcMbvDdcgfQRGOYNw6IlqZjfVwASutTjkWE+UwAn/v8
s66bDKNF4cqoliTnIykNbkMknaiHOrm7VF+1LlL+KPFsIEhG5rayKLSFRZ62
o3p2OSFda7uPAiLNucT9dRLaEam8fcQ4psEBskKXCiriQ/kjfLVNykSSJedB
KoHOc3ko/E1md/WkSOplsuBnfGYQLiZ6pPjD6ZBjUU7wx0DmJ74GYgNuo9i0
SxeUmEwrUbsJJaDxaTkgSaKPTfHE3INvcgCDbYuBk2ACLyR5KyJ6ZyILmX77
gONssSN5G64WNkyUU5xWvB2DeCURDVdScoBo7pbcOLzaX7mPoQp9vl9pabUb
TjEDkJd6DZK2tqcSfz2iK/0ejyhr5G+EnH71sFNLMNlk3gVU0UNjpsbQ0hfL
UXM9Oi9GueFekdPO0KkVpaowqDVzJ7OQXc0mRp1sLgfx63Jk69vCSVP0dRVE
8Fd5Rbz4ZZAzM7oS4jkuJSQ0uV4xVX/SQB/TsRB8P7AAKZnn6X0ceBtseCMY
9ut6ybqslMrjO6n/tA7tv8nKrUzsZ93EUKrjc0WaQX+a5Okq6rv/LZ3MEaP8
qq2hL6KQL0ZZGpJg9pB7uQWiZqyThbFsDn281xwe31cUpM1+eoAdJy5I8mXI
2eEYyTKq7pmv0RdNK/CliS9UjJZcsGIkayN+j3edC+WYPJJtGQoJxub2JfP1
PYC5Fom8hqcorc7K9hTpBsNZHH8qQp7HlVUPzMff82FZJBv3+VAtVvtFX7cO
Dy1MiYsmQb1PMn/ajlrdsjcR6Sp9CtrI62SFEdJt/3ML1RFhUM0ap97iZHEE
3cLR/i11PcvFfl5NmIrZyOavmXO/xanbo2Hp5SLExSIfQ8BP4DPrOrjGXUzn
h4vbYjEvThS/MgRoD6CGPY6kZhh9fTNxNdmIMqHskES1vRw9WyfprDcPsw3U
9U4XSlMv669xibw3OXvDptya1d+ghFck1pVxQ6W9USbUqZH4qvGU0W0YoyPn
LSD4sSnEz+0UwaDMTjAw2Wyf2Ff0aD0A0LMTP/EDShVUEAppHNy1hRQBrzSr
W2N5XMgNpzq4ond6/B3ZgnvboTd4rPae9HjsMBZ9Y9h7ABhlXQdhlVLAOI5F
zt/h/qUp4OTCt9SvCOqfZE6Y3EcyzB/BNK+DfmyCz7vxM+cmR1122FRSLhzh
Pi+q8nX+5vMhqOgkSDl6/ltPo5AWujNcoM+u82bQ+0tvvsQIELstx8SxoI+O
H4IHO7/1WswQm4TOPkMOOLz/srtYVd3rN+1Owv3p+TNcs1S1sX/OPLiL2lhp
9aRzojbwtN7y0HORazA62zgfC9PrO/Aa3YcMN3LTmCO4mXzuUKZ7BJ8nkPon
LS9DSH7myGOrInd50l8OptSa0dQU5HjvtvifGOrSiBjB0oteqdeLo+3WZ5lB
sWpK5mGpjusaDf/LPeO9fiIst6WxcSyRe7tCQXoCCtJWcLAH09187Bzv7QI9
gTMHu6WoojG9oWIeZGQB+vfH8/STaP+ILaXyEtC1GrTINPxGnCU2xB4lRoxi
wDbAuEfKllIbZZ6gvSSCMJmNA7ZaAVBz4n58Xk51coygs3W+eFJqzNrXL1Yb
KxyhUA/s2KK7RTkE8im7djB06xXCU8h1o3W5a3Bu76//WA3lNHLZU3vMc0UE
rbhMKdz/GX8/f+pUCMINNIg0hvvS+Jf+ZFrNQBFwStLembDqQijP41HWc6B+
50K6iwpkD3aq2EIKz+EZsvYBH7ctXFYte03zetveVLtrvB8Zh+j3OoG2nw5b
r1I7+bay0KgdKhg6Bonc1DfI4QEMqeEngQjupbRjDlUMrGCZglbQLJQb6Afo
byJee9oUW/gD4CKEs4reYJvNVkCtSl686X1+c/++39zkIy871RqBvxzUlQwz
EHz126WbZZbELHFPMRH01GH8R7ultvbT4n9MjUWYNR4ZZPmSEUzZZm7caujk
rZUChG/R/wdooHbENx13TS0iPFtKT4+8ylz7udnAbifXIboXGqDG49JaPFm0
XBFcgHqGbtrBmMsOVfI8swdhjHsp//7iZSxUamMx9ijBuB7D9bdOZOnxsSUr
L3M6vTXk9MGevEawUTrMN7H3WcZI873luIw5ZIGHdJMV1maIqp0ZBMSub1us
iikyQcbRpvt4HC1HJ6x0BPEwUHkjdPyVo1lwHxlbyWX6Gr1FCTeecYlC82Jp
BJZHIHZSj0vfRkkDss1I29Kt4sHaRhq8S8AcvZr4RTTRmh4sxluEla9xzJ1Y
lgRAlYlj8PnqauVskQfsveJI6gtD2AS+jMf8Uo1+pA3VVmZro6J50mxTK/JX
i3hR5TzlMUagRvA+YYJ6LkF/CW29m835oXUZV1jye/UiMKKLTw6K5D6EZp5N
Tw2OjbeR3fJ/iXSWjq2fIIOjhNj5Pg+uwU0XBS2pyumFy5AwkK87T+RviYqz
ZCmwEWT0658LsnxtuwDzFPd6J9JW+4crsTro+l8rc2Y0JBkN7tPb70/Xi4I7
muunySDTRAZ/XJIkAhtlwD3Zn9GnVxD1hXn83QFM6SEDqY9VvaZ5Hs/Y7m/H
96yFAGBBXlTlOq0Lm2bL09Yys/p14Gesy49GPtuRjg44pI9Xm4w7e7jW9/49
mYiEvqjyeuE61SnZTznJzuvv48WbVVbkFr19+m0FJCwMdP61rVfwno/CmZwl
aWCtnBOL1LQ3QAMVtdfCEi9qXb9ErAquBzFq/PMSp0gkRdVOk35vtMVNzolB
zNuWuK9X38lKbf2z5DnIMUFDRyTmzwc37UoFXH0rbM8SHJXH46pJrJAsg396
+73P0Nn92w3Sk91x83/HX29GaTBIMBCZfi9WbtSO/nbKzxpWJWuOeJp0jdsF
AhIRD/HGZcY7nNKPiDzwL0c+5HJylq3PfW1aLS1enoltaUOw+z/NlZsXcbu6
Y4QrrywOp/vZ24S7ZIgdkMdPMtcMyrmg6LDMiI7YHLtA7lXy627B0SOW8ST9
fSklZJcirPbufVseNPeDEfXnWgWa6WjsIx/JbTZsqQd8AdjP1Zt6Dwxo9DdU
eB+ENZeyM/O9CSIU3nlqlgoW96PHScWEIBAh4mS6b/Dr9U36C1wzogMYe4zM
vlkhvDJp+L1uIROr3y0GhaX/V7H+z9JijiK33fFnOcxlAYcQ+uRfGg9gLKnl
kJ6TjycnyjjZPQUlVLh9mwUy2xNhQ0qkT3ySY+mhFvWd2ap9xzasR8j8rwPc
GVjNdjKBFxPupoxZtIljiicodR5v/VxSAavxU0CZR7ICdvLJ4Q7eKcXcrlGj
1sx8MFCc7zy2wWz5iV2RKeZ777kpA8StzhaYnKlNzZolI07znGvGvn3LicTL
sZU/JFlFg9H/x6WhuxFxpvoestrhuK9qN3wFuEds/PxkjYvrs/yuQOdXBoZw
syXg2290THkCHnene5V4KALOsuOwMfhcKoN4LJhJQg8xGBDxowEVOsbfbbcP
4zgKQ2dohwnkdKq8BFzKHKEM1mAIXCu38jYziXKR/h+/XbpM0EApzBLmX7Di
j0Ak8z6n8Szsj89cruUH4evvUg8L72WNlefUh9aRqy7kyNtw3gKpFStEyfZN
KEiYDTwfMB58s0yNIbiIq/ZCkTWiVQ4dxOFhocHIaThGMRae+r2WE1nEUoxA
QnfGnzJbZU3GEcRdm8CqSjSGjqnoVgqwnXlvR1alErTs2YAr+TYSpEX4SRNK
mg9XC19NNTk3Wljn+g0ZroZVGvFbAtLK7qNnqxbjtcgfUnEqBmV38uYFZv3T
PaA0dDU0zCBVc2k39sTkTcc14F4WMJwfzMjMCa4H5muZr9ECiLpD1IrELPW2
nm7lR5CukzTgn+M5hXnm2NHs7JF7ZE1VI5fgX6GiAix3Ne3u9YipFPBaMW1D
/2Ln4+p6qDgGqXbkojbHm2G/yMmPjm2UPmAMeU/w+JVH3K85O2XjyAOZtVwH
6M4CFy5gxJsjxGTuMzk1vtuKYg8XqZxN3qnlXgvDbcV5ACrylR9eubuAPU68
SMQLZ+UPyyyU3lVOhlxGsagsxsmcqEOJJzE0m/vx6NoOhFcZRHutJG5wbUCV
NAttHG4dJUmd2cdiLKRizFzBk8gIO+5XQyjLXxqAYzlrwt29M+bfK1Ux9bqk
WZJXKvbxxb2XgWeAtWsPEQ/+UkAjIpr/V/3P1FggHBreNASIbp/J4F55CU8O
+xZ9fhKGNgAVhbCHKOXXNVhPIO1ogmaIWThgJRucDeMbOVJFjWbGjfoWShCH
6qoXGs1+fnUt4DyqaBeduYMI+yyUW4QTtSCWI/stxBVwk5oupQtJ0yLIEdVZ
mcJoptLwx/nyL7xiJf1/+osFPUNEdfwxQ3UBpakol4eyllzmgwW0Gipt4jtz
aCBKvyGB+w1YZYec6fHdVNwS5b80m8uEq4ZYKNcvjKMQzQ8M+qf7N9woEuf4
KXcZHvoUuu8hk+wLziZsXYk3PyMRqfGN4APyQuxrVlV0+B0PvOCPL+SrbBzK
AzArfbx+lRkDzCje65tvrM1aRR+DtjbBwVnkouCXsLS0DpKwEG0xeWjiNLuI
TGbEkLTdbzpdckGgrk2wN7klKzLvoHrZEo+uWEHlTOpjFQw+RY4kGtD/RCy4
QP8P3lx7kVNYMXmxMdHtDqy9ehIZjJIAqqz1SZEWCqysLBJJNZcnU27qgzzZ
EEd5abGddOGTZgqHDvV+Yc0Z08J03gjtQkB23Y2V5GvW/4o9ra0uOKs0LhYS
TVrodbEbjFAqK4HHfVe0xW7OOrmuqRVU4KOKZ8Rnn1BV9PzXc/OlVDlz6Dj2
C4AiWt5UzAWA9+N6NM6Nd7pYOL4oLO71oHS8EEbXp9FNXMk0nDf4hU3DdZ9p
De9Z3cbIFlYFxklrqQ1FqKHXq609/VfiCmwlbKoU174ykfzBp3JtyI2RTsrX
r2DmbLFMdWsXIOETESWbG3E5eToO01eb9KL7Ke0GaLM4ivap1TOwShQ4VRyH
3FedQmCKOgF9EJnEnpecHeJlMNwaM25+gfTx1JqI7eP+hVFV4vMOrGZrZW6v
EJ2I4Nm8K/BRieLtyTs5MxOglBBOjggz0SyAdf96oS1lQu4lryA/L6eusBce
gtNkwXI2kEeQs9sySag2jebEoqrbtcRTYqDMe391PvXuk15gHNVu0fGQUIGh
qhdpf5iH9i2xYbMOafZwTMKZB8F15z4isHx9N9XdTlMS1SldPRBKTbuDmepU
AV+UdFxuLjXBJKvIO4rozf68RhRY3uzbHAr2b6/VMn/nsbTVEmxP8my9Nprp
9EJtoml+LyhReqlBMZUdFGSlPtlZ5A0xwrDe/hQ2VeUE17OkMjVoHn5tsHhD
XhvwF5FO/sNtOe0c+EMRyYrCif+SrGiEg3R1l0hct1aN3ry/Zv1p0dYnLkiG
uDtAgkFOFNuiUez9LzQDnXKsClPeyXyQWtHwSNZRghnKnmY5cRu/gDf02oZg
v54fxdbywbN214c3PPzhtuR7mjKeb+PTMbOUZBAf7YDHZLxDbwqisMBRpTG2
U8h5WMpkXiGZdAmFs6phhXRARv4A0PQJcHkMTquSLsyd3PGgUCFfu8/bwNYy
CowJRZnGaFEwQwV5C4hlegsYwIKUKpdR9vzcY3MEox2mSnU9tfxDBygmV9iq
GF/PSLNvCPYikMieILCPM39dPBaT6kLWPYFgbCeKQ3Aag/gvsF4QBmSNaOYc
6IZED4UzmuWd4A2aOiDfejiYVhIZMUEeD8jE//5VDJ+h8KDnGJrKL76wOm2o
xkAFCF0MkwNQXMwlP/KG+UDaiI4NHeX7ON1b957kAPY4I5+6wTiNBdMnUf1C
oqLNCXLB9klnJH86Oi4xGWO+IBtbVXrX+lSeqC6sbLE6G0VVBydf5Ok9use2
qxGNVGSQn69DAlzBba4D81DnVAXIM0iBVaqsrKjWMcYACNFZ4UcOzroAvoem
tW8BMaaUMBAA6ANmdKkbMBXfPpVx6eW1g7Oc3WKlSA5PWGd8uILOKo2E1rXG
Ye2+kwVD67BtdLOCzdaFmQkambjJQWBDNtJYaz+xtvclTle6B+bOFtKET3FE
uY1jodLDkds0npDZMCuCBv+9KvMDu/c83Up4Vigk6nwKmxpRMwBvirc8EAJo
AYtjo2dAkv1qQkvQt4TbJK5OIgM1Ich6qEpI3aKszX2BS6B7h0lD+CPxiQnl
54YNjdRafKkYc7nqnhlRYFa0XUIk+HMoyulGflaysVZxmueO9dKQ3yMHU4zC
UWmeSyd8rjK6S8sQYTQUfwb0m8UrTxcB+dfS41tZaHiWIlTf6QlZK3LpTF8i
Q1bhy8OADfy+zr89ObBe8RJjBPcc6nWWoHcFeJDhq7DX7cejtcRUiCxRB2ff
IF8d/n+TP2Ia+QeVscuIbT5sFd8W59j0j03WYdPKl2dS1h7TBZtkwbIC8EGv
jyhfLabxSS8t4CobPMbl/ZDkWz12e+IrkSX+yXbDeQyBcnzfmf7MAyE6dg4t
rYdCIMtRL/LMkZMdryIqOHlcAhEEpoAF6UtCGDJ0y7vVSi6O4FS9R29XPIjl
fxpULzhRr9+vzqT8ryNil59n3Bc/4H9R7/UWaFSurWGWyHfZuPJCu/tgaTHl
peXBc3DGSLbSYc77csJld5a6Ud7MATM110Vc1ITcswV8VpUdsySkKWwqzVyA
Ql0dfINr/fwzzned8l7fCBU+mRE4w+jdeKz8XoAd54D01g42tOxxnaDi5yN2
VgduXtlczq8bWhfwp3veRf0+picFMmZqeRmUymM4Kgz7V6moqYLw1SRAQPIe
3/sE58kNpXdkytlfvW33+1czSlkFEIn7h/j6Ctun9Qkb65blNm6rc0ivfPBl
2gNshjLaSqwDPkKh8Wfbeq0mb99vDVH8aWVfNO8LsC9WNOT3JFe1b/+Sui9e
3quZFiyGCB8JV+vjCXs2AMAYtWr3oasRwpoHb5I8bDquPBjFMfXw2bgGBnQ/
D6fSUjfWJCb2B8OTbuhCZwp1BevXc+o9ogd5bWAZtiyKixkfYRAQzYy0Kf6W
qrVHIXxYm6vPnKalXG6EwH++hH4jlmC3PjjrolxrsNxzm0gz12VDx8wHBFmP
VC3KS+81EZjJuw1KBXzZGlakuiizGZweh4me/sqMuAuOV8W1wyd5t/NPeTLR
0wDYLn15TznOWCxpU5wm4vW8hDDTNs0O/PyHxJh3X6h8sjjzQnuTMsNFrtz1
gj2GtPmmQIJIdMSkE8MByCYn8QNRh49Lsa8FMh107ZkJszUchDmyxPz6dzx+
hnMNbbicbnmdxy92+yoR41/4wR2lWygqtTR3J7bZajgwzdEROsartUAcLiHG
5Wz4cG2XgFros9lHqxL7tacqzy2qCJP87EvTtT0w2u1jp1T27tWZE8JCSX7R
dDb9pq/yiCISQEMCsDorf3UzbKVBC/RdYMF90Xz5iE0CLpaysZF/8+2dReYf
S/+qR/Ho3jxbPiiJHMD13igO4MlwMMg9DzfOGUbana2bAOr21KiPBURaUQvE
11BnVnDWA9JQ1YP9mf713+3+3KIXfUDSMaChu4OE2fZ81kWe8DuM2cYjE0sL
lt/+asgdxcJel3jlCRlzTL8TcIKQETq0shz2veFVLZfsWP2PlfmOhJx9LxaE
bIYWaXpvZP2/qAsvLwpjjPz222lTio+Kg3PXmcUVP1u1Y4SxMgy2EHJBqOU8
UuhtcoLFbhg5TOy2LLL5CPEj615ChzOxdwq0qU3tw1CGFSVv5xqTCLZAQR8n
on+IWziaHq9U+OFQ6+6uYVrVKomU3eev/J8k3vlYuziSxgy6ySEmLKba7n3e
oxA9WZ83NcXBAmgJofYRtj8qgmnHRdIXJw8Gee7pbJ9zk1JgZjL+mruJ3JtU
ge2NDQfYaQz5I8fhM212KcgpDxIrAH/zQ4N5FCpVELBTuAzZpfFdz1+ADVw0
nHYCvNKJ4B/P5E4ncJrMiyBh2zUP+QpXozfqg+C5jpIBZeR1GitlJFAA3SbX
PucajjWVLJQHvxipcJuKG3cWihTOwup2S1CbRtotChW+PO9P3dNUy3W6JwRC
FA/VGt148Oz4QOfyLLem9pe255fH0jbf/SYUUSPgqlRZCv7IMArzG3rFX+J4
k9IO2Ya25U0aJu4w5neOlT+rTmWQGjePMGEHnxSUhkC7xHqbSKrI7onEygOE
6OzNjsoffLIg+7Y53SPaDGp5bn0yrniAbAe3yQyQwqAIGe870Y9uciDpUSlr
jFL6In4mdio6sphXJ2lC3S1T09cgRY3PFtchTMIEjNWFTQ9CFpzuUWDxOxuE
8WywhN5DiPFrbU32eyQ/vuQY+mIMsm0nJ1zYlzcOE8NfUAW3lsn6qLg9gaq6
FEOE66oQD2Nh/Uh35znCglAtnSOh4zrDLLWucP9ushbjos8OOKjO/qGHEXjx
wPRFi93svjuinMVCm5mFrlDM5dAFBPYW0/GZlAqT0KlhDUS9IQ1+ghzc0TKQ
zXJltayAaf2gQX+3l7k/C05igPUpNsIF5XuBwqLZO8gJ9rl6RZEsGYa729vD
/LJ1VNd1fA+R3ovTMIOMSV1Nh5cufJX8IW5gYzebbTEzUtMY71mXgM2dqLYo
w4OjL72pTcCvTrG9zoTqTmAAxJGW8ImTT6VUe9XEILNHGaj2uDm5HOaDy2Lo
pqPIOcWHS/fZiQASwNaS7mW99SN1lR6JHn0tmMsyYfbadOyN6P7oreYjUN2L
iN4AstSSlQoHZdJ1qXCcVUC1xW9OAr/ZfFLy1JrfNgguzRhx2c0ALh+O+358
9lx1H3wtxCBq3VlmT+Ovpjpf55z+u/ef4DTKKR//WO61IeOLce+UOeCsSo9Q
yR5Uk/1C+iUgZXdf4GIg/mfcP2vS15pirba5aoq3kqOTIOz9iCR8u3nEAEKM
4yPKSwYRVADlwD+NLoxxiDtuVZXLXRMk3gfGrLt77pzvDPwvYcSG+urQPwzI
q0XEGzMucMMty8cQHeScSkEK7oK2E781mgudEZMLw4IIMW5kknAAYVMxWV+n
Tkk/OHHwD4MY5ZItYzptwcCgb0R+GD6X4nidh1zcKgVqeM6JztHRGMVYvJ6/
wMaOw0Dt0+LJAA4subZD3bk5oH81TN3qJ0+AZLzlBG0OMXarP3wS+urvjLWh
MXy8Jg/ggWg5lUd7JtJJYwizQO9IRPNxRwzZ5yiNPN0855yk37qeQTyuUENn
1s7r8g8lDyGnS8uvzvT1EAomzmrTPqpikCrEOfm6fRBwQRhWAvCbbcEKWzs5
TZCsUyf7fAstE4ipiA++7z2MgnYru2VQDvqCpCjZE1+wDI67BQXeBafw9OQG
IKHlCbnTqVNYrPl2WhO+Batz0TDXhzzeg6VaGjbtHElpCWEkCbCKJMgjzctY
bNv+dtauf7RzBe/YTW9Us0K0qB6bNlYfprnBJfFOEaRz3sAFyRzUSFBoDW2V
JSMK4VBcN/ds/3C98h5mRIQm627VWBXlLxrbFg8xBRjn0KEVipIryRzb9xZS
rNBgpvFDx9/WWids5KYfnIFQN2yrX/XPSIvvD7lnMxQUZZvjk01D01TwQxu2
0tIGr+gMjXN0aR1EtN6AlVRZghxV08bVhX3R73S5MGz+4hM4DqHhJEyFpYHa
IhqdOi4ERZh0LGHcCgukhb1At6UqJK8XXSEeE6iK5djVsuxYxaz3WFrOgq5o
iBqKRaETuciAjbGSU1WPlLYewROvbrQ7LY/s4hV2WQbw0fJ+dD2H7GyfAdZT
zv1gS0Qs+D16jWc4DdQOGpm9c7gYM+ICwtp8VBLepoEgTHXR5NJRsv5Q6MGf
HjXjzBDQnbASYc2daKDlIN9tYhScpjGurlGMpnsRbDjanCkMHlEs4c5RkTch
407GfR6HNYzaziYGGGqsnj4UVb1+3nHyHusRq2sKg3jvFCCSzbmImQpOEfXA
2RbWj6L8/5ZYmwLGk4bMdDXTaxG7dvOW4DmAcwrgbmaDXhDYy0QaGwkdmnLF
rZF3GgXkM5Wv0puqqOFo2sevSG2fdatHnlrEfeOYqMnuG1FZi1RPxBcGnt6i
kKr+klfcKbs2GgcuBK98pjss1teCX+M3CMxbAY9N/V38jjlyR/RnPyBjtM4a
kBcdZjsf5l8c9tgJVg13sqJBRw9HzysCNGnwi6ueyOdWFk2sDwE7orGBo/hs
eYpXq8xDZGhgZkC4wxNzN5quGCUBTz7jcEY4h3vQrnWVL0Qh0nIgklQfbxrw
P3EnKlq66xd984lA3fLjWoC8Kz8X4J+ILcJ/A/jiEkPKdOl+8WYARbhv4YTM
Ocz2bw3TIGxeDvvDqO2OESy3lL+D3vgXkY95Cxw7pJx+eZvZjY9Mk76XXL68
wU4mtR9s88pI7ROnbDLqUj/sAx+tRzHqgyjeWUXvWBY+aMSixHFuWPrwLtDW
k2A5AVhPzvIgqiOzfLjkJFhSWF2uvt+aFJhogSyhOxHnCDPC2n4RWldbEGnv
u0T72EilsWIbpr1L7iVpXxLJTQ1QVmc0ezvTgQu/3+Zky74BcuUX5Pfx9ajL
7kzZbMC301eXUETOUoHBg/6PbYrGkEUUpv+zfEOiD0Ecfw0+QW7x8C0N2N/7
cmvVtRp/szUzlyITjrUO93DntFJuHgcYUNErZfkRy+L+UfXJdGEEP8u1+L27
69Wyl6/+I+pHi31KQu/rYCzgM3P4tJGB51XX/d4LjG1QOvsfSyjoSDPKSvrh
YmvAxJkFFVFGytyrNEc/xGoaQo/d3u2JFdJOp/wK3+DqfSJLmHntwdZgz95O
9/LqsVsZnqztyMats943b+FJZRDq3luvIo1vpcaKHabT6VCLLrWwXABkMR1/
2amKsEGiU6CKfakM5R0yOqKfGvDYqmb6mb483JCHd4jYl9eM8c35QZgCZVI8
YFqAZ/yrL8zRS50xKOcOvc7RrWljuuC4aVqAui94rF8t5RyjAochdzHEVxUz
u3Kkwi2NopqCtdFwKZu4yszx29VgREkEVtcwHwrkSOdvR1aGBWogGJut4pS4
bOsy4BcAzL1ggWki5+CedzaugQnhTpuRa/AZGC+AfL7lGsAnFbbPIzXCdPHx
r2F6Je1bDG19521aM8PoOmlFi8+vp19I3Uq1HmKOfSy2JkG4CpK1D+Ei5zwt
8BJ6lBdM39dXjYwuHSE83NCDBHKyb/isvQ1B8q32B+XJacQSSAaHK8d7evFk
Bf6uVfK0kds2snMA/ZYPdEWE25Ah7njcySi7w5GLBAYVVMGhmt05arg25jhz
e16HJW4Q8iuTMIjkfB4TpyabEmFityADokvMpHsXoO66Hz4pP8q5DEIesmjr
U2ZANI+WIj0PXmUIFayWfcE9am2D7k+1IU54wv7NJYQsI/SYb9nHxtgHXU8F
jbfhZdJtMJBTUatQEj12zJlAMo4eozet4R+DjQzWLpJuk3TwnXOiI5c2ov2V
cnT8nVdRsyL3Ulnu/Lca+B3+4L54qkPyl9Zs0BJMxkTiqHV3DfeQaDxRqjXD
J7pPwS1sMSf8VJaCoLLKSHKItUZRXkLwB/DToFnlF5rLfBGhXM4drn3rD4HM
Mb0M+l90vTo8t83kD+pOLYwSGCatblwhV5CC3kYl2eanHSNwBNh6Qwhspeq/
zm4BbKDo7A2EycfGzD5KtcOUZ6xLOdYBDcNS1TcpZnU/SvHz1mwDjZYUEaZZ
8JIghcOg7cPN4D/CNiAGMJE08DCgtiTDFXFkv+AIKzpFyg8NrwBxTlcTNnJ4
g6ZAmPn4o2iclpiBo2WVVFLWhLPw9rh1p9NodXa/kf/x6KHbXw9cslLdjlNZ
B0bz7l9AhpBVA7bPUtYGehIx8W/409KutEJnU60SMbrc2lw69ulNKgqddSYC
xa7Nohpp5Rffd5YA+b/4f2vsQhKYC+i/bcczg9+AMqvIdNlyIWPQ3aXBVFd7
u8dAzGzRoBVOMR5opf9zGGfRuoI79ZBthH6D/tN6MgP0PD3oIfqfJdWD5ZVQ
hH+Mr8xP49bjd9vOH2/0g/+A2iLmif7fHqKeMbxrZACKxwBLZJ4ANAe2AjVn
hFFV62g7rbkAUHWPTTmVGRlvLQ6DbMrI+OMbbkqsPP9Cue7p2/9t7qdiVriO
TybLiys1ETMt/UCGX9TiAkZUID0gq3w6pf6ux39JiDoEtwABFDc44hS8UlX8
kqD4dOOGFvYC9lccj+LH3G0GF104DFxu6T82rJWIP/nnCWtjeVYhFl+V5aDY
jn8yI2zsc6dkY12XrhxK6Fs+6RY02TYhiTpdPOPEz/oywANZa8vMX/YeqPWZ
CvWHq5xHtb9qCFKc2UFfztA9DFZdiCh/t20ip3SSeDXbupcaO+Azm/bTX0ls
AYhseJT/jaq0yX3ruaq5trbyronxXMvqJGehr1m5yLV2LevAi3UIn6blMQqm
9GD1zzS704QwYy7fSNO6ZkYVf0Ci7vPZk7LCltLuBt+YkZ3k5ctRqGX4V4d8
8VQi5qPpYBR8WLjJvJLjq8nW/ef2NTtFpPP9J4a9/HtORy1Wt656494crDLD
3nUy05R5lgEc09qiaxQefmsnbrQdk/297XQsAA267tqWUUloKbDUyL3guMFW
hwdfj4QU2lnRWZsfeN6RSFjaSb993bb3i5A0eTgtjdYXbPApHG6S6JI0/Uol
p+MHFXVnnfiBhGllPnk3QLXvu6hO46tB5lmIF0SBptto631V/WegLFVbWS4m
VWFOnvVqfTEtYTE4QXrMYOf5kDK2Q0Tsf4AmLKkz2q63jGkAhYPdFruLJffw
MvqZoQbQDeuNHql9S9WYx2VO8I+IlDqZyuW7lMab2QJ6/izQG5LGabCUwKw2
DN6OGobI5P5dpzI1AYx3lyon5/4VcVqiW4i4u2uvujS7E3vJXTy2AvTwmgJM
Cwn4lUZR7C5RaRidVuQ5lxbWhTPsrEDSZ7JVb6uHT6tL7Q5Nif5uRS0c9Ibm
WFbEkedFa37j4NUvl7Mg1Y400Xf19toKFRRzc7bajNMRgUPte5d9tvRvkPZt
jNJ7bP0P6osQK5vIPTYi3rVWBUl3QATQV+C5fyZ1CJ8ZnaNGxZ9jiT/BQkmz
L23S7tqKt0uNi6fULId+Tl4gRlAudNdSA480WQVrmRXK8Sg/6nfLmDXcqtkU
m2VodAEoO6f8dOJh94OkKOSvhOKiqrwHYoSNb+OuDKKfFvBM9mqTtDK8KwVA
5SoHfSaetxGJ9v8+24qa0ozjf9EAFhvSIjWm3EEc8UFIxZuP74zSuD7jVmep
R7oVZGS5Vffl2fvXaA22/GIf7qBPjk7vgJQ3F1FBODlYR1hCdbsCIvUUAEvH
fFEqQYNj0tR4BjfieRRwAd8CrHDPU+g9Ms1ckIXjk5SlJhf1NF+kllKG2f7J
kvRbcGQ0F3B0nnWEDbE4x0cAYlUh6kC3LFfTyvus0bruHQ/sNHndyGllhEOc
dGOZLaoOT3uIuIHD/BRDg+En6UJPCqn6z2b7RTbCe8NQLChTBe9mVi0103Ph
tS3FRYikTIuN2VamgcZn4C/FDVwl2+HXpAJTkwmBkdvrNtM49ZZ1at2Ye+/k
rNICaeFC/EZe9aLABNoQ5y/cylmAKHqfqNMQ/tEByYVmoGo+OQVj2vkUPPpV
qjsuuddkGyUkLIE/4cBtGDM+YBYYiZxSAPsaDf504LhzDYH57BitEMT0SaGV
uvaDVN3lTHxut5BoCuLkIDr2DGi9H2G+vuOoQA+wEMAfO3/AasFu8iODGP36
2q+HMAu9Ti4SPEsKr1SDfHVGMkP0qwyMJ0qifnJhcxPvpCySiCoOkqc/F6Ph
p+XHPVOu0j676yRNaWSEJKJmxLW/awkCQYRAgdHP4AMCyt9JGmW0/z1tu5b6
lZPWXx3pvZgHzgFO2dkIoW/81cEYQeVgOnHxX8kRi6tFWWyvgyKrWDHAYTos
tlq0Z+mNnY6T/7PML20hj1/Owfn6lqgdzDfyEg/SH03PA4pVVsdLjESgWvAn
gYpOYJj7zlxbmy6c7KwW0cSXCwItQ1qYc5iDZqPsAnvFmV2eHUfD29X2ANUI
ARVtDwEXRBEJjh3q5yErLVW5uRKbNNNDrYbzAszef9TzVpfjHl1ZruVQ/YGT
o847/cQ1kT6jYU/y+/gzEEap3J1614owUTwD1dqG1Iz/GesKnVaHMxmsDwbQ
IrtDQIgPwhYSYrPUod4mJlcaBIpmA2SgLdWCU4fR8oUl1lfOvjpNVA3GgxWs
j0N9CtCQrn7fIBwmKin625ClY8DnRx1tfN85Qd5MCTZ8TTER5LDrW+GgQiEY
cQ62o9YkUpGU9oIJ3woqJI7J7n2lCAhpg2shGQYFz7i+RZHOUCXFXLn76tHE
30Qa5tKOXe3c8854nPJeTAdGNm/+mT/9v17+GVx8FZstWPq3GQFnr3PUVNrs
X6XoBhip6k8LjPybA/1FqytFGcqC+6XXHRE5sYC8D0PfZfs7IP3QlFPb7kDo
K8xDzozoJNzQUDja1Y3DMlBANVVvCnm3M2vUxHGM3GVIT7TXuVZ6Jd9hhV8g
TzSpfyORP4G6924Y1QIvsE42fgDwUTdrAW3TAnqbcXudnSE9VO0aUSifZh1a
diCNzz9FvCcesp4Kk6CxfHl3Jk8vlSg8HLMxSTIJn/53UyUlsGseatlo/5LV
HxKAvHxwlMkxW7wvM5OUmeSVQOvjOaSum9g80kb5YqKKObu5zLIZAu7uPTaa
ROGHg2LiB8N3L1yvhmWUB1qJwcA/M02clav5fYIfFcshlYviUc8lo9wvPkxp
7j/c09Ngw2aGzupVAHqBOPW7dY0rRkoa+f4QnznET4zagb0O7Ch/Y592L9Xx
r+TCyYBDxm8G47nzvqpV0yZVWL0kxjSnDmmawVaKoVbxdRSNiKbTv2AjymBM
VyUyqeSo3QriHif+wkPwg///QP3n3DHf0vLZbP38Fr3tRvyNpArILyGFtKc3
kMLMELsASN1ZCUimmtr4psQZjUQ7LPsTfGiLLc/qBBwldj8q13oz9qWT2PEX
phyjC3ED9rtNJK6TmKOUAcoZtIMYlL0yl5MWVjkryrxCcKwtsO9m0hHkbmlk
kTq+cuU93aKUb0jpsA/tUXtKSbPOKyjMiWccEXYleRV5DpBpZ+SVJxRZW6+A
y0P5fTULZhjm5ifo8UAFD5AGpXEjAuhDYN2GtvXMJCdVuixV1H12gyB2zl1i
W3+/3wKkRQMKi8POq/gTANtkK5M8yJoyDlEA2gFfStM89e5mw6J2zU8X8o0M
PzIz7yYsJRCdTdvfzpz83iFXFI8F5YPeRNB365op6piuqzk0EAKZynMwDuqn
akbLbdWFs3e71mx8DuAcGkuHr34gN1tNPvSoRyEYx0t57Is179TUgK7Lx9DX
RqWvagA7UbJRzx47QqQdcdJ3BLtP9Ay8G6k51g3O6FHPk76bsXrq5N5AvPE4
/iC5Zyh9oTDnQYY6yE2hIJvpET9/ezBiIknCeZ2n6OLCiA4ZLRh1pEL37pIE
JOP4Q8ghS7narr81iE72yhtdKLqvWLPoNswr1ikgLNX4iwFeS99zydihLO1A
hv8kVH//U++F/BWI/B8w/VtT1eR36kRoIh+b6cp3QUvqqGUN5GmWdmJcmfXj
flBrYQc2dzRIEzqOqOs2xTqXanz/7/AvElyWKInsWh6Ya2valTK+SVrnDjVq
EsVTvNcA7MgqNInKodlw+5PTL49BbuYo7Iu34zfriEACHntSd6mMBA0IKD1W
qTMNuhOMXIah/LE2Nzn7+PNa5zCL1kA3CSKdfdAchdJfRq+RDzi2ObKQHi6d
EPYqfteH7dX2KcDCQ4Rahi+F2geWGT9MldCxr7zbhCfrO4pWwdbHQLoklvTP
dXHXq/8RTs5gJU70SdXPuNB5HnG4ktal++CdkWwe/Jv1cUMTKKJ++hDwLcxZ
IL85h/adBYe5eK8G8ABjwNMquYH25LnrB6/5OzofsxLbaWqHv6DFv8JHwSKI
gWx0pQv6Xb6X6VcgAn4rCVajnY9AtjeCcH0oAZNXXZ0fSxCI+kh+gL+TGnQl
6zb525Jx6AlcUIMsgMvr10WwQMm3IgzYj1HVx/JHPTcSumg6dK4LD8Lv6F67
dVQHIgq623xmHouxOYhMaMaFMdnH02XH3LkupHhrUcfGv1bVSHG4a1ei35m2
hgFKk3ocuL91Hwnj12MNoY3tCpPl/2n80gpRClayYP4s1skWSwiU+GyEBWDq
VaI8aH/FwWsJDCuYNtpH1OtyuiRvt7jFIQOP2XZZp+Son9Lf4yl2kciu8bpP
9l8JvfxXCy4xa0zTlUS09W1V1fqzX45LJByE3aY6jmkG5OWmaarCWQyLOn15
0U3HxLvk5lSvyGl1Y+RCS3xtgctMsVt9U8IMYsANKT6LfwFqP6taQ4zERkT7
fST7GJWt2gTJmWhwcT6erqHv6gXKdv6PbC9YyzK+d8x2bJArYGvD5rCUJkEV
rv68CezSu3BL80MgXTPhwLkpV/X9Jp8/779aKdM0YAGa55wdu7KkXM9+r4Sx
kIYCHMxlq9COEAUC/jH6dOA8CytA4Zrw9aIGDTlyOdYmVJXub15W7c+TkNCs
4R9HVjWjO728qwBQJE//x6evL5L2p3OYjjeucdyq+McJSpa2ZV96MzYA7Mgk
vIcmc2ihjM4eckm5P4uGryhUi7VHibdvn4eW8sgpOAXD0+ie2W8LlCGjkQ7A
wrhRTWpSHzj0JA071QO2dHLDqmJyrPTHLSscwbUCRj3PM10vsb0dAd1zTpaE
1jfSvc+Gazd2xBkdohO5dpiP+3s5vHT9CzsrHCmY+lp0YpFIXekCzY3H+1Rm
hviZlC6Fuq1p2Na8JDCMG6DdmFQjV/UVaix+wYQsj1P4CYTOTPMRRM6eFhtz
WW8NWCM85hxQWkuV1mn+sQR1ZAlUDDgQMsdJQAPiBD8fQqeStUDcoat9NlyF
spq7ttF765v9GBg/fXOB6+GJZgHl5XU1RlIZd73c5CBlkgyeZUfsKKdlCBB4
I1oyW6ez5EqsRpo0uNmBXb2sjN4e9NrZEkWfIsbxkJAYBkdyx9w/bgTP3DMZ
mnZiXp0AwkAzbECnhygh2UiCm8EOToB43+e6anTnmt2SzsGo+QEdVuzT1ClE
Xqagk7pgdTZUysEmeo33gvbuYqpPIyw28XqpP+t3bj/JTlGcnVlHj8zcZMZO
9e0FMN+X1vmjrPKrNaRWs8DDxtQiGTUzOdFEX12i8nWO9Tq3iXx0nT2TdyQR
X7T/ZFSB30sO/Sqb05VFZ7TtIo8TjiUVuXniCKbfl1jdnDuTvyrqyk3gjWYj
LEj1p8z5+lXDJzPJgfEbySxfI/wbggOpLHZC4OXuix2p2CZfIUyLMLGcPsqN
685RUtzaEK4ldIdx+cplUcpOamOqIWCMW1liSBi6nU/8ZGbknG7GL/hD6FqF
6y3rIojiq1Nqw0vXrNw8CMJH6hqQUlNoR2jgqbq72EonlxGCvoyIzszBLfhO
wLac19EE242FhKUj17WPqdURAmWM/Cb03HOjseJ12ih2c1lq+omnK2kRVPn7
r+fTvM83/cn3swME2lD2iGNZOZTzXCDyxYwt/iS1WKCBYvxBUxpj+0ru07eq
+h8N3LuISh6vC7+nhkM5YvIWBuwB/NzTJm9h3C2jORjlMtN25vjM/LmJNsAk
PnTpTap41sP1rErVaXXuWDITOSCkakxn72VyNSOiGKGvcmaDNlxpKhpZNRJm
T/G59+AkMoSrS9ep+hOi/yp+2fXDCA8o8kIbj/L13wfMeRCf3iEtKV7K1wd3
U+AUrSC4tUp13Sj84FAptPhs62qlfHawmTPQbFB/975dJuUHprJJaM11TBoj
EZdzFEC7Qrv/HULMp/ZvrhcCJ62M6vBEf1M5cyRMfAQS0dpGW3IkM2obTzj0
I/qlkWbVitsuC3HA6jlo41nN41eR7rCfJXYo6df2xeahP7q5UzZb+6Ie1AnO
BrD6fABiTAR7xd2KA9Q2kYxPKDXV9SyihLb1GMtw/6FaxTh7uRb1SDLWkFDh
ybnwfhUe1AQDlJOyvNrHHCX2taIWRSwxUImilxtn1DbpI/eUY/mzgMWYNov9
wK40WfUKRga2TyDN9dapKa2cRSpOlypNRHEF+CoZ98JlwCioiLKndw19TvqF
hJFiZ/aK114omrZk/QX3/yDb+xYQIOdji98FcyyZHkv10Jq2XxY4iowRwfn6
YVJsFkKKqwGhJ1Sg4jgnhrTv8GJhOAj4mZ/R1IY/6KrFkoDLVnl4myAtoj37
18TtelMV65M/Ta+aUMN1GhFmz/CO7qI1YvhWy/0SP3Fpt9KKVDApyTqk/pF9
OyHWpWb/NMVTb6k7yrhCz3khPu6HH3RmrtLbyeYELRgXUZrF/9mdMmtZa7yQ
+QcbWLqd1MwZ71gaq0B6WB10EGCF67eY2oOrMhbCdRveaiDfp84s3rEqzhNB
RIxXRRj2EOnhBpBTR9keVY9+0C5dZS740V7nyuRTthULmHCPQ5Feikrt9zBF
zH0lPl4n8lN/7sqedcKo7ahBESJA6ROyz0c6ASkqlp26F6wiBapE6nSUkvue
9Uk9HQzcpbkP/7heViqImSbgXbifR6ltzKiKR+w6JWCzMFI1PW5XqWhSBdY0
TXG5DNPMTDo5CR0vSt6PcG0HjESIxmp4TXi9IN9Pzv42SuClwblujokEWqW6
sF1YFGOfnXuTIuSxaFdc/uAR9XI3aYbnPYmordrBvyjHmHy2Asxsjsk3+4WH
p1pK4al/GXORMorSjxpKqM449F0p+GksAnYfQKeSi5hlN9f+cRtQ2xhaqtX0
2IpyyYGwNTwe3+FaNHpJgGZNpPC6o/VH912PZe/KNyFNJ3u01wXBbQPm3vNN
jl7zKiJZUGk5wc0JLoxMjnMiwDW3dqhP2beMbX6Dk0bOapjoFobbJwR0ZTpO
u/IpTMx3fKgucnoW5Wy+Wfp+CpqWUKy6GFXi6R3NbYuY9hmRp8Je5bQGNAPX
uIj76EDkAGaFjn9MvpfIL6gYqvG2cZJFy49ZWSiMO3hobR+CdFj4w1dDEAGn
pT9N+BXnY20c22LNvyhSW5SAjeOMqXlt0cvuCVD7xZA/D1x8kfGpwnBSQnMb
mUnVwjEPasiy99eYN4pbz7rSG6olY5ko2oTucRQIoIEG8OcWZSPB6s0LaYrZ
5ioqMCt9IA0TYcy45bMILyXHvg7j4GklL1u2M/oh9zlDAUf5tFG+/a5c1zHH
1S8w3paOeytPJzo3AsoC9hwR25ede+w4BjKOCbUtaYvhOWlagtZqro4NQD3Q
VS36NzvAlqnYfpfE6iW03/pf6/Veo8OUSzYc0wuPgZkxHTzpVglICXCZC6B8
0zABgB3DuMGGgaqpcc8ORuBEeeiFVsYhzy1RINyvJ+4r4p4qBuEKTmW14uBV
CmO9VUy7rh56p6EnmqZUg6/O6TiRCdHuTfgUqgC4QEYmc0i69FZodcK1vW+Q
YefaR6DhLlzdR4GqNgETMDxOdGqzEKGH1hImERaKk6wR4hxDN/OKuuNKYk4n
WudMm9M0K5fOhgHB7wiGDZGhThP1bvg0c/fhMichnTZKB5rTLrWTuW4ZAaZN
wj8mxw5DxAhwPoEfEMivxuGj9NpWftzbH36yO3126JHp/KD1GXWP9KCQjrjE
Q5TVC/+THarbo89oAbfQEnXeazMcdpLeRrLDEGSJO0TIZtnUsc8BlEBAdBQF
hH9osrOrQ68hekC+673YGoKZsfdyMPnVorSGZ8Ye1m0UfdV/d8nVWdKVxZHw
96VF3RlSXkkUFBrxiQezvBfH7FqPwTdmxfcfbQEXfAixQMU2BC3D4WFBrQNY
LbSLzxmCDuy5lG5NOnWHMoX51xxik26Kkb7wllTG2cQgaMglqqj7xveQvX4l
4ougILN+GSySJPSKld/AgHewdtLBfbw6QbRh9dYBnVX0lzsvbTSlPf+vHHkJ
wSsOmPhp5fDUAocduFRLFG9C84vmoSvtK90TdkqBGaStkZJSRln2gegvOGbR
2AiXBZkNWVvRnZagKlSAJUdWTlbmTaBwGaVplW3DqAg04Mdb/9v9AH8aIco/
uqbAlyN2zh2B964oUCZzgbX0gwySM8Wu7wJ/7OhnfnodT1pr6pMliq3T1+BH
ML6j+CUdJRpbY/scMuB0BvFzUsinDEg6Q4Xf+rBBN0AsTDWmfu7Ok8RnL1tz
Lvhzx0hEj7y7bo3eAoZ+4Aq5Ru722i7XZP14NZPmJPj42YmRtsBMfmDgfUAK
UaDGgiKYBCxDyne9jEauC0R1A6w5XcVCxw61SsJ1YRP3Z52LAC8y0RLssesV
QHKJRSdxr96pB/O5mbHXvJhwrFRFShurZirprGRGxtKsbZ2cucz2ghjk3n98
JpB7KnqXcGtghFMyEDweqHVKpwLVkSDOc/1ZhTcNvzSuatW9KvmIg7yYNPwE
bWqVIsSJH09Ig6oiVVNXUROq+2P8XX/+DswsEAiQGEaOyeP2btJz81ayqcrf
r/7SgvfzakhAkXzgR6JTVVV3Uio99FmjOr5d0otN2kEASwXI3WPqtHs3mvBZ
z2olh3QTcKocmhQtj3/TTKaut27dzWe2EMFBOJhL79I6GrhKvesoiQNaBeoG
y8FSsou1zmlN6BGDinNRUCeyJ8meBFOu8PKh5wN8LHn4hMusNWnrygyfjBWy
Lx/fbWNGJ3XZ8PnWTJsXCYdhK6qvnkh0aL9RI5YDEh+Fs4W3IJWTPCZ4/Lna
0bPC3RucQAZ2vrNFdTHjvxfEs9frdQ9a6bLTaxBYmQ+D3ZMSiLwCxD7vTd3+
cjxevsqd0jPZ0uzJFjLHBQ85c0S+spC0gj/CblemVeauQ13GaaRAmBX+MN2y
Bm6Ed3tqG++Eppgk9ZN4A63tPPg5tN1Hxnw9rvoiwho2Bwz2w5j1a2kVI5Te
xFMiN7YZqk95CVRHJNp8ee8SQU+cP2gI0jta7DOWWZFvKyx7iXJkM+0llxia
Sq6rYzQjJ2KxeaBNV/6fQuAElNt3imsft70LHyuazFsXLbNikzO9xWHmALR8
TsLi3zpOwzfYBN7QVyaxweyn8cIurDXw2YFPZpoU0mdrHs66sN5cH+gf9DwI
uJuSFB927pUDobT9YZ9jc2YVYfqdAQM4z3mThp2wrDW8gMU3M/tVub1rTRGO
0pDqyaSYsJ0Q2I8D3+T05GKoVBZoJirt15DNnVi8NIuE/JXr8aYJXBdTmkEd
oLH+Zp3BFkHPnY4+1+ofSr+TzPGveLoyjYBLuHrBF0MITr2akwwv2kTIwfOI
dHdxl9AZdaTKCWUi1nMUjsddsdJ/bMBLy0XCCKGcnEEoiGtD7RMvU5FI3RBa
jqsgCjE1/+cpmo6HPtWAD2MDz8hC7vCrvWUJYot6J+OcEAiMLDGRnLsqQiRg
WrFKlB0yMTjCHlcZ/zBebPtOgOiC4nB69fnE+0O9Rrr0vw/tdc84DCkTb48p
Bd2CdBwu2Uvsu4lDaBq8/uh1KfRB2GipPu06Eg35llJNTxgeWSeKSSetMTYf
4bLzN1rktzXBS11LfqQKOmd/tEQZ6chCIU0xvi3ZxLwEiF8h9APa6tS+ASNS
TjJ1XkRGN9+AZuqWC9bYzWbFHyiC9k5pj7xoBNEht1mKQFN/CXUSXc6Kt3S7
ocrHA0bmgA+PpSKkm92nPcrBbv5ovSLYszSeRP5E3ZiHXOfh1fwKluBtrA5O
U+59ZjnDVNdMAIrswknkWIdyHS/r62qZUcQx2cH9PVgHedR/7sJRnzxjdO3U
1QO3yKWMfPxMCBlRjV+7WUMRFAlZ51w7zgAdnPcOonAM5WODv6o2CmS01Fa6
BoPctPMY1wLxNLiyzfNwsfqPL6ugP/nxECknn3w439RTqhGYfvGY2OFaSg4i
uq4LcZTdW5pBN9NajmvFhwXmjUHsl+QepQOJFPRuA7XEQUVQVYwrAb6z6yro
Tunu12PKCWRcGoTpIQJJ7I1Jt9dgb3BD5TsMmwZ+90WGrpoggPakcoIRcEjO
720GEzH04fQrHZfaBqZiHswODo5A451ww0CKnZzgHA0sH3HykScI+h2MWJ2l
GHXFjXHlprfqJwxkyomgRRfhBaU+U+VIAo/EGlH0So5oyHDNiGEdDDFAfMbe
ZxzZJtbBBhA6SxNvsRUrXCcl0cowZkJkB2x28TjxYdbHTEDvqpd8nHDhMJQO
r6ru8dFTrviJuJSW9UbkJ1v611vjWo3AIa7IshHmFToi4U5DC3jTkcUeqzBC
r3B7l08kdTMqRthvHCGK9l422bBjoPM1icpy4fPUMDIQnI9fKWW8Ckgnbtzg
Iy3VnhZAilqtQHJ6NGLf72xUm9WfUynGq1gEOZTsaJ/7WUJt5KCWNUPdycUB
D9OTgavlSgrJwkFA/TcrH0Ad5+cSlmZdI0XVmlGMQv9/I2oJnQ3hN+KNWsAn
PMiy3Ltpzy1hR9TorXFIH8KuXdrEYoBDZ3DDA9HAGHj8qa6WKqB1/I8D+Xon
aNj+BfnJlBpEKgNDqnk4DR8snjReWlds32nIvLVe5uJ5KUa/RRpPUEnccju8
YX4mGczb57PTrXPtcPk8qfBPW6XH5kHR/NPDVICyQ+xf4Izb2kRNUjsEH9pb
GUoWwU2mfTSunG+mr0gYCQktos8LOSNVNnT7LRcU6K6bXzCWnxVzcW30Nw8N
twch7PV588JYwuFo403daN4RCUhOa4gyS5ZIEIZvJnyKUnYjOfB91pj9n/yn
pHDPRoCJ2cx3M2qDAQ3pByjDZ8YgFvRV2uA50YzIVW1nfkXeAgilH+Xt2WP/
4MUgojSIOo98+3hCELaaxaiwTgBpUtow+G/LMG7GXOvExGFHw1MPPYJoiqLm
xz81hX0hlUPdNRLbc6ceKa5n+m+N6+vQl7kNyoIK676XyvppV20Ut2Qx8sD1
4OWy0kJ/ROqUhHJ45EugzNd6E6GGeMK4M/zzuLCAI+WRSGxAI/jE4VBl5SmQ
yhMmt4nWudj4Xf0mWkesaXMN51JAncksowOGkaCk/29fdWRgGngyyXPTsq99
wdSRm0pI9T3AHODgEMYjIINIiiem+LTEnRp42qSOBdtqw7AGDp2s0KoLK/Vl
SyA8Bq48nG+TEuFx7iaLxpIzDsCS8VoenjSLgI2TJXbdieU7TBTGhEVAM1zo
qzEoTCc8Nfgvo5+qQUkT1pPFHESV75GMtrPKZcmEOf7vUCrW1783Jt9SbmSw
ZesK27BpIxTEl10nMUngI1p6K7TOXRoEIOR9SqhLLBGivhFCbKbt2GsuA3hH
4UP2+ef0oOgAqiITlWlI9XF1H6rYjO9d4FihnC7J7pUciQgtdwUo18d5sOyG
7esHtM6fERnyiq139Sfk8sWGv06OGjlUwKY2yHAiTUfzKOs7qDIRTI+yqyCd
2+QeXzr6bXJ3dsYYSfBleY1K4euJ5W8xBSCjIABvVBdMIyInc2SsFPl8c4yl
qkQFBVyutTEj9LvEJrZElH+XnLK7ltn8Zs5+cWuCI0Ui4aBmCeP3+UkLe4CW
RJJSIpyZJDEk2FybRcHHK2k6FL/pMQgowUyCe4NRht8GDpN9JP/o18IvvuK1
asa58VN+Se+JjLozBpqVRuveVRJsEomsLC4EY4ollMPcIVvzmTM/+etnQqWi
27YWtdcxPwAdVo9FeAq9C3nTXtxPKQTT5aUf2Cv6Lze/O9Ef3x1BujZlEI+J
QQVH6FUNrrc1DapMX9PcntncycQ08eKOFL4hGTAMlVzdX7GMCMWcWk+gD6g+
jWSHnRxzXo4ID1vEqU86oNaEnczc3ANi1VgBRbCvNwVyCLVXd1YSwWsunSmx
JFASd8YoSHPpxGsV1SuMboH7LQK/gzWdF20OKHuIaBfYWCJE08YxR/DpoCec
z3NLuBa1xKGxxq1xhvkKk6hd1ilAqNaWvmoEzw8CUXhZ8hTADTSoqHzxVl15
Kavqe49U0f1gHv/hmYc7BanaDeK8srtVyOpotbCo6q2Fv5Kw1QJ2DvttphgQ
Vyc20ZSjtVQR/SOGFYfb1DI9x/KycmRVHwCl2oVZh+ukG3xZPReLWcC1opUd
IBFEFIx25CNR6lSn+HN4ROKD2UCNvW5FzsBdzyRJDuMujMlFZSlX6TaKqV/c
w4plPwvIyMIvyI7lpet5jzQHNDrpVwPxm8NcUVWkTclyVVT3KJ9qxBPnPOdW
SPm3/+zeKD7Z4p4KECerga2ChzpRIRE1x/cuGoQ+7+c+Kk9k4EC3E9WYoTxD
eKywGSB39DDUJow0had0r+o24TkS1KdVccue/ZBSFhCSootp+NkurWF7nXsh
pq2Id15id7d7cfdmG4ZcY1tlCINCkpG4f8tGivtzrlwZpEMBZyBZOXvleY+1
4UVQIY4BNc7L53qleg2+mox95Fz6rg2QQ+MQ9tuHkj/KsG9tZJxDTN7kuhNU
30GTnTyUeLmY5aqS3TKrLsTrA0YcQrTkhlais/UFK2nsAdCNOes6hFT6y/aP
g7kPl37iD71HFcpCfohUlge/BAy3bbK8ALAA4VqkLNfgIA4OFKGk3jdLeCta
sn21uIrrjaQQKQWSTXk17XDhdqFK9/SFlHXrijD0b+HZjje9vNy1xRiRC/ll
L9oYGsKd2zeKo73qpWJEPttgxO2XuIC1OQQQOeDOD8kNrk6ENs/vA8dVzTuj
TfSeGpWZgQsGCCwq6WGvzGesMJnUKdtKl356zbb5QcJraqpXh1y2JljvtBg0
Ntd5veMkykqZj39eXsmM2qFz5s/bL21pm8igojQlFzKLwMl4w7c/Lgq5UI98
O8P+/HxqBTnaUNwrdOP5n0URqiwbue6FF8nwvus79jM9cDGjdzpVHsQCqK1W
NH4Iu/lFifbIVTPv7XxoQs3KB/QITjlOu0TvzxIAvJHBiW6HfaoppNQeOzBI
HLE6vYelfJI8CZgsYNDr7eRNi5BVOYW7TLXCnb1tEf3qB8vZB0wZcBXmXzih
/tJN6IRzG2BQ5IESSIJDBUUX/xIBIDBjYkQzRF2iant36BvSd7bhrFq6Cict
wZJFcKlrG2u9/0T4cv3v1w49QXK+0GCHvFdg7D0OK3ovWUrC0HIuFPuIzkTD
CcNqJdeb3q8lRcar1EwzgMUcKwi3mNlHQDT0K2+Ge5s7oGXimANroAevrogb
nR8jLe2KZdsrA5KP3V6NEZj/XcTAUtUOIUj5gAomATg8bUbCqv5fNpwzdQUd
r6+IVd7Q+PdiWSspoHVkwoOwLsKDnBqoLRIPkrPI/rLZCqA99kQm+37wA6Yc
J5L63qJRcziriO3Y89fCBoRtQ5RCfJEZ1yA+pOQR1/neE+d8NU9F9OsBBqlL
3h7B8yTmV7oU8k6PC7EY+txKfXt2lInkooS2wG6bxs2SS3rz3wijNtcIVKJ1
iCf6b++XRibBzm/y9BrflTqnTm3C9WX+ue2a86YERWCBar1BQ8mI+oJL0nFf
VtpdeGL3L6YegmBe96lxunNONwP4g1ZOi6os4s/5aS8hIj8gxiaRb4mpwU6P
EfkV+t8zNCEBw/6B+uG5M7TwyTF3Hw3bG8IOKHPfuYSXi+lNZIcxhj1iJ7+5
XMAi/j6tfi52MMBkz0I9+KdwvMw1yj3Oe8eLVOAp0APaLCFrcL0HmoOUn9Wy
Ij53dz9BFXuGYYssF0is8QaimwKi91/26/tTeObdain8vx/IvZ2RyCKrYWu6
ES0zHDgWK/5TH3VxX6zhsKrwJ6h0oUblqBA28/REnNMk04vjq/l45lb61rF7
uFQ9Ag9IGdr041C2mJyAqNmLLcCZbaYyAIzXxmpk+lbaMqWeNO7nBohGcnnh
N7FNh/MsGs3Im6o8cGOC/s4ecE8AlJAD6Cbx2o6ZlqB3gYaxHFmbd6O0c9LS
OSNRNs2CECceESVww0GicczWLU7t2lBJZ7mSi3ZTd9xOwacg0GZWU32XlH4s
aUHJM47WebFhulsMDBvyEhrAHAfHpj8ZRbH8NBPBJynfMVyEhbeNjNtW+tZp
dLyOnyKmX8eojmvyUG7Dd9gpvLRQryRaw6ItpvOE98dB/YgBwhS3P/VnlV9u
SsOPKTG+CSosJBTAi+s07Dm5HvAmRX+o3kABZlVS/UDgrDZYOEEFTO4jsmXn
q1SkwTREqEKDHNBZX4Rx2VOY776uz1ayRPUagjzBfHJiE6dQiXC1um+FboCB
NEuemnjudd0TWWAWqulwtPFbTzQMYgBkBkG6E0C5WBISE1cAPXqBRslZ0E6V
DmJ/aLdMfWEIPNulbgzBd2jN0ZQzaPMGrYNlNq52LSDuTnJDW/iprj+GBQyi
xCKjSPK2wI6zBWAhJ8uO8qsfLVG5Ibe84gVJdaI0o95OqSVmU2mbQEUXeEq/
UBy/UOpgtrFTWFsrSkCCigxsYo8KuDBvl5xFOveOo+Zjubk3dqlfGIe1CKNf
84R7/pVKwK+BKaK/lzSVPgdYKnc3yWX2Y1FRK8k3H5Am+QWswoPlBGREcSz7
0uqb3DuFBm0uIRvvrYoiGj36v2LrIq59Hnb2t/4KPayn8s+SCBiYPiSd2HfL
jRICUU750K1iWApcOuwRv5/xtJR80I5bJwe0hlTeujTkp66rIHUgrpcQQQHp
xCYOi4yQPninKOJQJfGFwEmwlMS5BbTmkyJA1Mzv5nBQbrz4Ql1fWv7PI0nK
s9/3yNh1TTrYr0U30kT+9DJUNxhRGtNS0UEnCOUka07vXjelAVGz6Uk/ptGc
YDTbKNVX6avlH6JKhDEoYfKbabaWD0JpTI3ZrOZGblPlVrhqZmVCu25eyOA9
xNvtaOhotiw4k/NbQb1pNWnPiP9sZThxgps+SD+jSNWl6WcMFFkFuF/mJIlu
1btgtW7EfwSG7W4lgv0j/oQjo0tmcI8XdO/Q+WIHq33dLXussSJk2N1OaF27
TykehHNEoczaa+2uFagW+jsbnN5r5SVvFc2h2zNihOOUofcSfDwj+CwOeKUU
3gKC0KJjsBOqv2Xj2Z0e08kGQyFpIQO6YslPcu3LVNGkD0rClvmd0vT50kbe
3cXTM8WkwlHGOc5Bqf0rjp4Z2bMtV0QiTNyP+B7qd0X5nhpOtrqnALeT2hYi
hO+wFD3OZC0vUdSaEX2ECVv2Xtl3DZWjrYjRaRVx/OFW6A42FO4jpVkiy8KB
mnK9ysrn1xK2FFA+otWr95/t05hc0YsmEE9Ws7uhO7Fi2TcOsAYsH8MSX2wX
ho5LmnsFzAeONcwcWgfES5VYtasmceeTHEzfY2a+Pta7aoejx1RvRNRJWQID
LdyfOPogsnOJer7vH6pUHZXNnQT0fo0+7SEp4QLWDyJ+Csi0macBdVjbBlCR
y+kvYDZY8ItWjOeE7SQdju820bR/+zJAD8vXrab/ok+LRntYA8GYpYBV9N+u
gu/XY7FRZcDuIq4CYoFaeiGodZr2uRmRVZdgLjvL6RFozfAwrFDNk13C8xB5
pPucNzL56W8PXbQcW93T7fsfehsFv98tkiwMV1CfsEvUiNBxFQuT3lSU80G8
BswcK0g1dijGtWboHwToNr+vFpsqiG5Mk9MK9JnKw7slGJ/1qjG6zyBMeobS
/7u8esQFtucz+hMVshV5w2zEvICY2eJYxeixj8gX6356GGO1/E3hiIRUwvy7
eDQPnTpDXlBYOnvJyFpyxnhU95+b3X1rMpW4gQyzf/J/H3O/OMAp3vTLt9GW
OjXPEhDhZJ35iLOwyipgncomdygJjzH4uojp9J63MY/o4KtNqnlYVHmChMnB
ZZJVvGXKGrmoiJm5E4lsnmuhhbFkHmV97r3PjfpFNkZyuCGzZ2YKJrkLbeLY
w1M7DA2sHkWqZq7WYV/oHatzYDchh2tNhwx61wQtzd1KqJ4W/jtKxvHrGdF1
hXH89rTheLN1MVwSCjLKCpEuFwRgecM9kzdperRB/OH48CLBTIUP6sNjcW1V
3nNLvB6cwpGePpQP7OIgYQFImjw0zBF6qjcDSQhr/3qFPrALBZfppJ4eoBzK
bcVX8X1X0OuhaUWjL+3EXVCHfM2KZPc9WI6vWOLBTzSscI0PvF0kWSXizB/G
OeSTXcfyOxKKBbxNgkmDI/vya9/nm3InAlE84yueE2wVrZEdzmFkpJi+l8+p
JYdfsM9MtUBKl0JOAnn4y6do15ZVomDCpQkn9ocMmHeVv6OLyiDKswH8lMlN
NCdpXUdfpmIxi7OfkO+zxNBqsdky1W8IzfSIg20qgk0Z+4/uXekCV4aBfEBE
qWl8afxIlqYelXlWIPQTraS6d1bSmS8BB3F6q6RBr9UEokhiwk9TxAnmIPIV
oHnkTQT4b9K5G5i+uSXXO8Qcz1YzZ8JLqqV9NQphtTRsqWvpsl5HoOTewSfJ
3+5zP21nRjMmYFbuZF1LWgs1hoCeG717n06NZwlQz3+r+DWYoAkY2+RAhMe4
w/5djpfttbGOmbBYr9DaxQvm729J5Do0GdkegoBMfBUGGunp48AkpIAcdjzu
hO0VtI41yruEgPAYjruH5XOAUU+5C99rd7XsutfC9VJjYgfimg8xwd6XzIWa
U3pcxjLufwQOhEKM2gBdp7ukz66nFmvSXwdpn4Fd6kf30H8urUKE54KRhnv7
fplAm4bPlZnET+3jeCnk4A5boxkXZy+Jp4czC+LkdWmLfksuMWYVAkUlricZ
XxPJDVOjUjfhlw00gzvEzGginQCHimWX7W71Wehi5Suspkucmk8OwIqmB8Wa
tpuGrgHdUjGEjtRg4HxBfkKsaZ/ioRPodT7t7xJDp+uA92cM+PtNzPP1Ufhh
uSe4eGCeTZdQIwH/x/GzRL4QTcT6sC4wc0nLIeUfRIxDmqdrzr+N5yhxekUl
GPNkXgjZmbJiVHNw0RZ99d1QKBbFNBV9lflsYyWxFHLBFd13cDQKaNuiJaIq
qjZiO6h9ROx5uYWXbXOND+lXNBVwnCmLmIDptXLs1bjKSW5ldC0UWMqRRWlW
Pq4w9lQ3WBZq5JccSW6db6vW5aNMU05AjLjP13hroxTtRu21SX3vyfDOOB5g
ASnKXgLiqx1Q21Zw5NYszJYC0aKR1OCK6lcnEIbSA3Pt5aZWlQIUMiSUhj3Y
VFS9CG+Q+dSMOgaXgaQmpE+SdsiNx8lzoqFwESVSamXSYe+KnUcnDaP2DpgD
WziaAcTCnTNdKQ8kk+vVdS663jTPPDZMgJBphX5sWwAuAj1D5OF2w5fRiACc
ST+VJxd+F9Je7KkEerv05KNxOy9Mzrd74Mx8D5HCdWEIY9BmFcszzlz9Jkth
FK06y6w6t9b83lBiNUbEqbdExE8yDqmdT9/rYyqKZH2oR7oFTxgbVxJtuLvz
5N04Wo7rrCPpBj0tGlhLsawoGn1GeFY41qCCasIw8SK8tCjfMI9qXb4KYkDD
3g/SUcuQKQ5tXqW+hkgEJX3qRg7owFvPGvvmqNL/lXbVXMIKGaqO5ZXB9RSU
RNcFhgKI31zrxACRW0D98mImuT/JLAWg+aqtfRM28XopHprK4OV0gCcWWcTt
xIQGtC0xrUhCkXSlapCOFYnVuDHksEWgUKrTsqKW+VcSI1JOTIHefCnR+1m8
+xeyS+8bjLfF8csXun0udlZv3yH9LJU9wRb9voriOme12hrbE7COJPz2kZwx
WtrbtvxJWCUN2q/VIxTJaKRlKPi+x3cVTG1IC/wiTGYxdBEu4ILSjVsvGH9i
TsvIe8K7E/67Cv5j4BINAN9dcSePqQ07c/EfXlnu4xcCMCtBNdvBSMW+fTTw
d60EwP5pgdhnJbpyZ0V0Pec/kWixVmzZ4mHdaOPKNrAwTLQi5yt9y0fxTarV
iicwNiPW70iHWEjmAgq8zV4JsLS2ftKJEI3ZugY6rkGWIo7mJxmPags0BdT/
FbGv8tTuRSYPHvKw7IZf/qpHPF4LkXUeaey2ao0Bm3l5egoRW84RJ2RHDeqQ
iR0KDlNrxCby1qSCmJScC9VGKiKo1+lxbVIsiZMA4HYUjhhoYjqt7a6hcelC
2ZYI2Em6QYBuQowx1wzy7xStEM3H5skdrIz/hQluFjjHwOl7LuQ9NNFBgfTM
7SuH9VB2ygYcI+Xn/18m3wuf/Kn/38vf3H0jvwPyJOsUhsRb04/RK6x/Eic2
15I+Pa7gTxwGZGJw9g6/3GJTfat9dEF6S1yTih1CLQYVKVnZCj33xPzo3iXy
JACbn5MydSAqb62Ns6oBMFE98rrdGwRPwwKyxXyKiIYr3jb4s14h/OxKk1pJ
XQ++CSD3pT8iTD8TJWJH3gFiM2uLigptPJEEQDOIBbO9bgmOArSfegBbQQKI
s5J5cN79JQMqC73f6k9rFw3ffixDbwarzUHajoAfpoXkF6nd5YtvP+Owa3jT
RBGThKASGjXVFugWjKyWkCwaJIRW+ogkD1/qKFOHN43WlCOMQ4069Mbyicbl
Em3wDQOTQ2fJUSY4n462V9PpWGc4cBfq8jw7N/e6xL/K/MVM3jNBDDh7lCA2
+q87ROf92rpFmgSBUxPUPGWeFLJIT4Fjx9DdB/mm9HSTL166S0jP7GGj/8Rw
cmzKfmk57XGJNWQ7t65kZlXxyCIjKthvUevAn1TLqT8i4sTvjD1N0RvF3l+G
WljskDmDLa5zS7rLx0KvcTYJEa4y1mfAfw/waxr9ZgEy4c9TAezGfuy+afAu
pJQrMa/95iseI2Bq4LAORy9FaM2q/bmb21oRm2JJJXfYygcneKtaAuuOZ8fm
pimFgRafaH/CdguHufRlXVebzbcQLJYVOSd6+Xe/OY5Qj6VUBASediQeqG2B
VdlOASxIdAb3Rx01FjoBseReEt6PrptVNSpl9TcOzbRXcg2keYveLSEDXntr
Vz0eB9Bo8p5n6scu8fo1i16qUYmHoDaqWN0ouLNjBJqn4CdFIWOtRxy3zw79
TKE9G6o/5RjqNe+ft4ZzNYFu0gW6yL5iklSd3QUghFK9JS1X6uKQorRjZNoi
niWTudaWcIkGf1viZzK0E+E+KAu/J2g8qrJhd6fhTfayH9GEhBczmSd8Hejg
IpplpfKIH8doaAFkT4bv5dBCr0XvrPY7KQihsmEVuu4nWqU+CpA10Q5wppFE
b9MJkSkQaNUQEzG6fVBn2CfhP5QioJxEemEnzLbAklkwAYOAIMhVO85a93CG
5BXUCM8d9hvysloicazkyFIZgXdZc7J+XtBsha3athIwvHxYpkDL+DY6GaxZ
kWG/pyswqsTFBvILG8puj31ZU6kRa1F/yvpuPfCJ//1BrVbiZprRZUa1pjc+
SYP5U9+BJrgla1hqXhNltqQ77l7WvN9jVZDCxStf7WYRXOOwu6N0vM2avDKu
qegWWSTma1CH7lsxqHewI0N2PCHQLk/0MF1qFwVWFFqn61fBgGDYo5zfBRGa
o5qYflYVAIA11VZlsAyHbFmeF/TXjuI9IODRpSA=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1J1VmecTA2s+b0jMy1p938K/bP6Lu647fLGyzlur3ZaWNPhf4RohE2DaNu+72a7kz+SwCLE8oSroA1/lKGL/dKuEiXLE24nm37ACrgNPRW7v4Xoh6nMA6I1JV+J59syMqq9D7RdG0CZZvhy87bFTY6Bs98t3Kfm/Q10d82MOqf4SRQbFXE9liATiziEvENIrs629NnMHirYqJqJ11UycZ5wd27NiyMYoayXl3fbIHcRFIXk0ThO3UBHfT0yrn7ECfZWm1bBS6XIWaWqu6uw2YVfMMvasUnLplQ9r97ykkTCcAonYHz5dpfryk2JNilkuDdbWxsaUaBWg1IIaANA7xMdhbiEElTDib2ELQW9ZW+RSDiczt7o3dBX/dq6OjnH/n9zv7aryZT2EfycGe0cU3WWMWbGP61frsgLJcFKj9aILkOnpzAzcqni/Y6g/BVRCMkSjWIogvSky2GYLgoBv1dDf6RA3kycV4msa1qtxOjViJO5oslk1/mESD3h8YInshUG0ALQY85zdhVq+0P3wEWieyeu5tYY43PR/RoLltPxCPpNfu7r9XMzuNt1AqT+0lBRjufbsEBJFHNwz9Kup+nKYnDxI/S8h+CYvaOmOs8x+qVbpYvLsrB5W4iCzY6ifPUnOPpEA4JWm1SMAOklBL0CGXrdfqVmvD1QG12lvMqlaVc0LTJJgDzdfsZ28/aeB6s6yaMnCczsxi50I4x26E4chEmFdcj2GfyxXdi1IXV7vIRomqD27/jsiCOtSY2ernrkHGpSv8fs/wO+q4eFBgGn"
`endif