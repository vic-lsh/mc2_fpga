// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rPXcltUWEm1MsoV7mt2RKPTFpstwYtcfBpHLjYhxgJA3eTOwUKCc/w5Sv1w+
6DFCE3vQFS3HQPRkaams1m6AfBoZz0GDpj9ceVluqzSoDfWfAoe0XsFJJxDu
6o5blAEbCAYexaT079h7V2aHPw5zX4fkj66W4KE0SNo2XSKBXsdpL3Eio8st
lDCpDCWNc/221/q4ay7sj7D47Khd9SyPhxxVt91xSYEn8HlyiiP/7Z6WOEt6
hKLtJzlLhhOuKyV+uIN4KGcOjCu3EAS/4s2xKT/jcQSWxJlsDxhcTsK6yoMo
GPXOUv7LjcGror2raNuTksRSWI8bRgwKyA8lfcq+VA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HBJSjosZ+R/vcRDwzkKL5pCQedrDUIfRVJ0HaXkrxZb9vL3YNcmFQ2jkQf6W
I+aPfnbUP23WkxL5BSuxsOVHukL5Wq/h6d+BvcpFq6OoDeCX+mFlMftluaIl
7d6uiwBz8le56leU9WlHBLNOGkNFUKjZSRLfJxzZz1iglElaWNLSI4p0fb7i
fzgb533VC+GD7mnh4Ovwf9xTR6B1Vs37WsR2CvOnZvdaMdUkuUECRJZ/0wue
c03YNXjWrfL5ICOGIV7GtyU31bNcI6mhDAA5NEVdt3Fk9QhSXFyGExULlKWv
E41DKO9PRyNd+LgESe9m3624CTsPhQ5luOzGOC+wbA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O9hdGmmNbVgknraapKxVhsAYq/3gGRjLxXDHCESN3ZjLF9PutrTUu4AX1GU3
IGiF/v/tF4sWzzhL5H9XXm/Kpb9f2/cdP+VillZSAdekQveXNElVPfkMXApY
MslKVKUOjomwktzHPJVGzvsx2hGfYC516GKOgFVmK55V1Bi3dEGJdQvadjOH
18BamOdvqOpMGzRW4R/AYDkh69QfCRYg/AkTSWiPCPwCDeN35exR4Dqi5imt
pGNDHZe13Wr9cI/s1EaNIp3ncjOnrKL/ur56jy/zzoN6/hTQrsKU6uWwrFgb
m6Csk2cbLx7aFY1MLkwbhAWgJzJSgEWZIBwSRVNY5w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Gdtx5EmRvxKy7AiTPXbdoheuhmd7uOi/AlpPAK3WOWkEYNhZFOyanzEPUu0k
5QfF2cBDXGu+asX0Wl5lD4CpO5v8IYaUg6xrRIBmQoSm+uDP43vhA9c+Te2n
Ks4bSDaP4Fx2ojyREe822iZhYiO4UbKvEcy/nFIx3weFqHjSvIYe6lbE4qnV
6pzFGUVfegDp+rJ7x6RgRxJ3M0puwbTbBrwKPo/z0vkeI8F08Kv/y4ItLRXA
cfNBQ2mPgP2EfcNVT9vAtaAl5hpWx/tqURIJwBw23zyY5qj9xDFAHKO2Ke4X
8FR8nnXIg5Hdi3c2CrXcL2n78AShLqJhe5Xi1qWXYg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HhJOuMt1iPV0IFjCddNAiFYgDFiw8KfY56IsS78iXxH/VidKSpHzWAy3HFR+
JezNUaT02VgxvKc/+sNePJ1lIuFybwXYbmrgoVdI6t2h//F4x0S93/JVhGnh
lsDvWlGgv201Uew+ApgAwhgQmIEYPh7B3Ymf/clIBWC7+FVaWdo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
T4go1ogeo4z6ap9qfhenoSgWkyDZi4ZPEqukcpZo1KDAApct9Neihy5yBU9Q
ezZdjubxxj7u15TCma3iePrS519qpznLOTNEbbIR0wRn87SbombzYxnnISak
TysBofOAAtSR7a4Q5FYoj1SnClCyIMBp8Me8zBVDpV0ow9OoeCTMqMmptmg2
KoXrFx0oAjeDCGCXnYIQkB0rEjMzYkA9m29n0q8PaHV0ECk2LePSYOuLMBHK
SVIfgEROhUsRQswB+raIO0eYriWOcJQciDBdaaIXY/SzoJyLOTGdjfZolXp+
uUyGUdaVemUiw+z3PfN5kbEHfp0g1abmYLIJsEgDCjsXg+HBetKWVt1lTUcv
rylrmI83hublRgq6xoavC4B3ZdpYYlStWW3waMEAVZn7/LRqqQMuPBLHEBgT
YGJCSzs+58vGuCH0KDTM1aazr8gzvErpvL/mBcNn12u/g1+WJhv325RoYdac
jVQSr0A26WnXbgOU7Dm8ZEovYsxcS8i/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tgcDmzd3Jf3S1HC3z+h+1bLl/aesFP1tu5X1gkELPHSC4m6Sed+2C1oh1KBT
UFVGCZlZS7qq7fTV2O02ymjjPlETU/Y+k0JASM3kzkAiZ/cWkgabPJjN/f6a
juH6tIh6pZiAKvxqbFCHMTi8emoXVvK/8OW8C5EyNmqylMSkQlU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
l/DvaGkS8q2ddl0GdAUhvDHSp4mSYTtZTLzNtodFFvzJ5O7haHvP45UEeSu/
6rVUMWdduPZA/rNn1AE+yntJo2E+VcJYgw1rwKe9EDBA12ki86NX0ZoJIsQe
dk0+h9mpqEM9bJJlpwblsxVBBWG9TdeUJ6CH64cpC1po+Lc5yDA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9584)
`pragma protect data_block
RnA1d4H6xAm5uuEEg+OX4FR8qbNR4tBKwNT+QVaIPKf/GepnM/j4skaHjgsL
IKatanC4BgeeFIOy1ANa9LTIPrIDYeC5FT9j7Y0u/fuD/sz2/rlQCQJju5mJ
xloWEMICAq0jORYRue1KlLOkNHFXd+epo47o0W1e0TVnRLxn17WLTT/cDZ8T
3huegBjw/ZwXoIXgLrIM8pCHDnjp1gSL9Fk7UAa+drFPwqeEpoa4PiZyq2cD
6XwHVRskZma7//I+yz/d44HOf/a2z8lIsPvz/kLUdy1zqXpoYzjre+sXTqTQ
UV2QcKQ6KR7DbP3ytLmSKoZJoqPSTn/IS9jGQZq0B+27hfFX2/7pAj/hnae9
myxhHsNryNBQaTStp2fRmfDQkNnC06x3KcAO6tWX1AZZxOSG1hS8L8MizdHC
n25YoD1Wi5OAPQXsJMprq2A+tdjE/dfE9R1/afZN8jMthX0kS3GX9FhH/Ijh
Yvh9qX8fF4h0BhRCC+MNTaeSVzgpYKHktIVpOVk3hDbHfKSggwhuJsFKP1KF
LyR/z8fFA9QgZt0B2O1y11frqNwwu4+hM3EXAWR9KKCRvwwBFvibSMCirqYd
llKReqr1svjeirlSEryKmyDQ2uSCJHuTlF7piPs95NyiC5yTncMClpDbr6F+
v51txwXir1xe+noY3m/x74bAKnOeatXLW/Hd3p5Qgyd3m3WhVM48OvElNIHh
TUvql7zzJI/QbizdH2fFezr2UPIDiun2e6meaNy0/3+M/62MFFEUv2jzfdY5
dTU4hTH9vvSXHOhqFMOBwJyMA6j1n0n7SpNEY4LaQWHyJvuliMyPKG5Sn3yA
OElHd18p+QKpZR2iJYvvo3A9/jEds+olDYTbMqmigR8hJ0HIPrvNXvdZ2ogM
BvCHZ/nG8p5OqK060xedpwF5lMTSgr57b74lJ2JnfxcPV0SHzIqKfMfIQCXD
9dX8HY822vXkRTAOQQQzF+gpskWD6fGQ8jCP6TWmxoU0YrCB6fUrBtPOmyOS
umuelQMPqSe/AeVr23vCdK4SMukT5dXLLtZIQBoD5Wxoxn5iOTpEevCqcyVH
JIPGiPNzg6BjFQPj2JD+fQtWDiBfXQ1BaFbkjztNXHcliR6lRANXc7eWZvJO
ejDeRc5Ql5/bjQil7bX+iA1kNyZjm3rCZC/Luta3xMsFKbu2m8EyDrs49sRp
dlDdDwDF2MB1U1OOoJyhP35+7tzueV48fCFR5Z4v6Sn0ijL3RX/LoeCuadHH
/x+/70uFJO69viemZfsaPG7MdP2u8jxzWwR64APPYGxnxP3fUj44WtvdnHyx
dX0MPHgHAMVDWnjAZxVG6SkwH1TVXD7fV9yThvoj+2IOlKFQYAwM9Uk+koZ3
zjuwbQpiOHg99fDNAD838dJBkcSEEaF2Lelv/WMlJjxDqDwZd2LYTI4KwyLU
4K2MHB/ik7xNS7ks5IP8++34niSEMj0w5fWZiRBcleX1hFT+GzuR0ukYIt74
8VAnGMZ2GCoT5OGZRaVMu8NhnMSwD/VP2C9NcAsqQYPvOyEB1/A5rvm06Y4t
mjBSXLlJBtcQ5/ZYWCJHsR4FNo7J1s9bjV3xUmNtNMKPON9hrykgzROMCIRY
eOqOWnedQziLcAhTXP2BQnnFHReGzJhhfkpeWm2tPBhEah5LoQ2oPxgXcxzR
cDlFGuo0rN+V72AkOQn1MjstzbLlj8W/pVeDFWbkFoMkYpGZK2CRuRQHDDRp
jifNn6dB2ya22UCSmeM1Iurbji+KAdDUPBRNMsYn5dXCKF/h0qhV9548mVyZ
oQPAWRdN4Y8UrqjxifXfPEQQmgFeTnj2pN9Dfx7rIXO4J9WaZSbwJCtENeE0
bFbZLM+tB1Z6X6Dc//fPzuM4PkD9NJRTGyVp3+JwwB1j78aR7kknhGhk16fc
Kc4WPgbWZ3sCHKUIKCa628sfhN+uqjBc7Hk0kgtl8TlbN5mkOaf7RioQi0aL
C3/GhG88FrqBp27dWpDUhlQME/Q/zxD6PB4rYShSCa88AwaGe+p8bg1+ATN3
WEuvWBYENHidE4FDN+SLPtYNyQv4wTtVADzkcOT3eaHAlAngvoM9sCoFmvD8
MCtbt6gAw71eDlnv5tyx4vK1hxNnWCvyIpYVJZVAIeqW5xdEL9xMaI6Trspp
OtrwdlkbfmM8IDsOxXsf3XTxryBoKjrWLKuXaGB/Y5oNGTqsoP1qNqIgvdGM
a2vmyi88ZX5bYxESDrw/k6IC9tuv3m7dikICFSgJcEkTxSZewCepUOdPgE7q
Tmo04HE92gHy+gmskFvuBgWtgsanFczSDvNr+Ch7I2kj51eGNIahcHMtA9vO
J7nbBFRGptrwSzwakBzPGusB58kdkaL5sUV+xo5KUmt+imOm11o2pvJ+/IgM
c6pAlABPgDz8I68SCGzp35GGes7kq984EWQSOiRpPv/YPDB4612O/Jd/IrsE
xW2aX15tMRY6Tf7bj5HyNsJKRotjjYuWt7wlviVdHMYJKov5/19dQ7wkG9dI
GIl/0NM8CCb2aXmK18ENT+eDtK+4zEkzHEllyWo7DII5McTD5FjiWEXWcsDy
ufT7SBJYWIVAogvPYbEA+993gNueriOShBN1le7VZLaA9F3+zTztUzFhDduC
gSUSh8usP6bYm80kKgVIaE3yHBzOr6J0KifDBCIwUNBd4gsK/GRqsEZc0Emc
mui3j04WgUpf6phR1IeGKvTT4UyB+Tk5iJdgialM6O0pZfPcaVy3dOkobx4J
JbJgnhbxbNffk0bEwxpl2lhbktooTkI7yy1A9gNgiA+wX/YLIdHPGVmZS5TD
j6NFdsdZ5Dm8lEBN4m2qSsNq7TjrhVv8MgsuEA3sK9aT5vY5N3VMftd2H4sk
I/tvwlKb8BqtTxc5mlPggWM15C5iTVwQz4qH7U97fyDer2+TU2+VfJOWzO5s
B3sVbi2xDnoTq6C4i5WhvEPARt6cEXy7uDHkMkX1mQ4UXcT1LkgzdPe0FESl
drunuWUD+UEAkkqPNg5AN4rzrKkGIbjMl99V6So2GtRvYmw8KrnfbCavchqH
Hw0kHt//9q0zBS1rIUSwpZbm/JKjH5jVVdRbIZ5tEBPrV4TvbTvoGLeaR/Dz
RxbYYvFf1nju9o5Yyfs4t8KnMImw1PWjndedMGGbgvk/l5ZFNu7LG0OlCKvw
v9lJWDQFM2Q8LHTZ13s6h8CEJnS0HBuAVW72grn3sl/mi/0w434AgY/Ame5Q
n5Ih8uWNsP6qHYSINDtUe5mh4KHfVzwJxiXwDeT4+KqhzZK/xYbcC1xtcEaC
DRKE+vIXo7LgeQoARYopu0p1prXGjiiF0V+NZHnvR1PRwCgfbJco3CXnNVKF
uSxnXuFH73dum7vygYFFx4jCGWiLwxpJnwnoZUbxY+SfclCIWbhMKiVKtivH
RBVb6iSPSApW9ZQQnbE1uiGfy9JuW4oWl0/6DaYAyeXKpBorjaMxHwu+EX0B
1jZUAVZRWlkZ9BPlTKOconv1fFnZ5I20QUyciphbqJ7vDnPGKoj7rBboNC9K
6N0S4LZtLcTS3Ffikn4f7eNz9D7pyi2jDS51fym8PXhbXkkGwB9/YM0/P6PD
ZWloWRIo5FTedt9OgUQ40IbgiQ//kJ+ArFcJCFKFulYbWapXEjK+SZyMkHEz
7xgkHiVK5mdLOY431ABV33DsBftD1oYrSxcP2GcOlaWp149N/M5x67AG/a0u
4dMIUW0agj72BRRwBny3+MLPlgbKzneos7EZrVHFwlMjJQlgpnwDUOTFWBqo
rfqdYAobLqx2+2JzaOB3A2mpUeTOn+2rVumQsF3rmmp+TU/aFn1LWLkNIhz/
m1tQJuWm+W7LBfA9JzeB4MPga21SPolpZON3vT+34MmbgTyGSEYvJ9pY8he7
zdXq6yDUm+bhnTJJwXBUcpCwNdJqnTbwiZupdryHSBVc5kbeTRa3NFt9b1i0
8AlPekCJn95dmYs9l15Xi66t8nTpmooQCyaDGfGZOkKMTtgv4jKIo5KIPwLt
jjLEHKFPEtI9O4SkIwNdXmoYwlTAMv4Yp3TPhORpOu/w+CruPwr9GsHTlb+0
KqdxQA5UUTNEfrbS9nmsA+AtMcYSu2Mt9Ljj0NY4Qq8Hynnd8H5WZF6+6enN
ATwUWPSI7Z6jB8hf9UuVl5g2OTkuC/wFOmpUNUryVmMtG0q0WO54eLMbVhoC
M90NW4YXxOuaB1LjJKLykxZvNHy3XAsRTrbNWzQmkiVIa1jo1ALfz9N7Ab8G
t8QoTHYLUyxOi0boJCGCJDZwQHcRABG7sCHwCccbvDOCWbefFVo/gg2h/6YN
xe4qKU3JEgk9ZRlPzFAkw41qRB+C73FtD5fsefldaJ16mKzIfwFyWPomlyDo
rFt3qumkCVGeiRrzsm4ckwEDybzGhDWg6A3sdQm8O4KdGSdyMmIgbGZzO0Ib
lmo4HK0DUQXtAkF51KoDJfgq2PEkeXD/6yyMAOeH3xWkouRD+67gjJdzm6rK
47x4SUEH6ZR3nFyhkNMUgwoWFNErViOsTSWkPOfF9sUpauAbsWnsySviT04I
Rn2TqKA4W0e9pk9K25rORtPMiRo6UcDnaDg8QY3JkqBxoibg0mtzoJfQTi5X
OnjnZhJm5BfI3X1hgC4DHEUKn5W9SFWxOSfJPFNc0Lea+mbYjGW/dGEEZRz5
6VSoXYlbxEOB9vvWS1Tmkra8JtJSjIi9q94nNXk5gQXNVYRPa6/z4rAKUYHd
wkIwvJToCDJjGGGwBRRVqEVy+lTZaUKHYo3TVLE8qqQrEgJz6wjt2J+rSAdM
uWcbKMpCqN1UbLRqvvXda3tkjxGX7aurddJPFHOWhJrGYtjKS4IQfUkKdfwN
e+WGNwpiJ66ouGFyLweKV5ueq/2cbsMMrsNkekMfHKlR2q51rKcB04UlhYS7
FqHjCTIj/rP8I3aSTH1k6ErE+tpJyyTvrOJnNmFenhDkK2Hfy0XDw9A7KGb8
9n8GSo4uKgTiQWBfRDjnyqleGlTiaFyBk7pU3eK8NA45GOQVPWrkOyoldHv3
Vou4IWf2UhaV1YBTkSsv6VixqBQWR06lr2myvVK4eZ3+ZhTkmalIG3rFelvr
P2LYoownMdR56ywZfSYaqFs0Y1DpYJCsRI5ySSukL2dPG3Lz9VfrtSIK2AYp
o7JKY4ZQ367SbcPpii1fg9tmnLdq6FChLnc/qFfcwkvbwDdsj/piJpvA7Yen
gAqDmpmezBTikGtTcHBRPAFKU4FVVwujRknLvRxzXRusL02tWpforNyTGeuE
Ev14s8pjWfRQySz4TjWekropNmssvEgps9Ab9ny/pHmP64DmVAUiWzIznJV2
PI7FD43Z+IQcVGJiig+tgTwqB5AQaxUUEhGYjfog2oymKTb4BNkwCOiqEeW4
3b7O4ShNdLF0qELIHlWxjiB2e9X2mAGSJ3VsvYeEUNM9GIutk0SDYttXi2AH
R9COA+7QmF9ujbP/QZm9k9hF9bfdUe9fXU5hPCEpKB1/N0l/Rx0dQNQUeE94
YIIwOUg24jP1DH0TDAK4ewa0l9A+Cz8t6okM+7CeJItrkxo4hbHoZZx7v9Kp
J0tbp/QB/GVTG0kNBkIxlPJi2tgOxy0/z4aPMehmlG744TMzKHbgryk+REcK
2cr8xKIIgEj+yBhRzU9pBMS5h1TW6c37XaRNqrhHTlp5ziI4fYDaZ2YdajWz
/B2V0suoPPweHfAMFoBx4XLGMKlfdroGfahK4CsKXITszKWwluqLu1sleKdM
muQSl+EEWEYyCAahWCjEUzNsH+0QPiapoomoa0CexdFLte8NSWyRVPf3XLpN
MVcb1F0bgKGA9n62gcrkjXIvf3SjlP+PGogx4odQ5A0bt1nJ6rC3PLh69scX
MmmPZHUaD90BQi3SNsZSa7nfctmB5al6hKiNTtTQmdq0L716BIDANq2SwCyp
WZmbLZVHa68Bb2oM742HMWD6fTn51Ydbsd8GmxbiKnwoDD93fGmtLaWatFc7
FaZN57zRGY2d6B/MO+//BbRl/XZ1Y+LgTbp8atykbLH5OTC8ryChChDG3+0J
8XJ29bjS3idAgWKpoKv0Wkkic8ByyGVt92STMATdxrj3qt6G/IVzzC5nfX7f
pCtBlqrsXGtu2qVMuO05uog9pFJHhryg8hCBPd72IyrN14bAtLdGAXC0UARW
kqOn1spwutY9EsdJtcssXRE38QQnTcB9C++SrLAmkMOTUSoxkW1t/J/xzmH0
0a0pSgqG7UGU4er6KU0t9jYAaRLpN3y5CgdxeNGgHJpCSCaHL1+Izk5r5K4e
tIM1ql7rfpPbB/FiEMJnERT0/Megzt+um0B91Ar6qcee2BY6MYtLSiwDqg/y
fds321slPWytjfcuBgPd9aI/XHLQFwuVOOaXZkt6c02fGHo4MbW7jzSOkGh9
/6CYBMSnxD+Dcobw8Poomo8cvSJfPoPXhizyJmJUw5dBFj0FHtEpNwrd8ALQ
dpfcdUAkoVF0wiyUAem40gM7uetOgx7EtEfyj8auCrdqjQATtev4eNC8ZL16
CXpq7tFGGydw8psTryppVYbDCCUReWTImgw54lkmcu5qMFfNcjK9Kx4vcoAr
RRHlvgJZ/7RuCX8zGHJdxAdi9HBMiN4Ex8bCZ9cL3KTtCjwtGqyFPXdN+0+4
kh78h5MnVazEZ9bcoEY+Dt9/uHmRw3nDxHGdMPZGWivqXQ703ZZgMCr8T8Z6
La1drjvATwOrKSIOKIGiYxiz2kC3iit+dLi8xkAPwtA05bsVIDkduAgzQBnL
F5tXlCwWRf0DsHdTdv+k9pahUuz7JoykHR2gXXyjm3bm3SuKxxx96F8sHetr
lS7d9XmeoxZIx7ENa+gY4UTD2v6MsrfPfr1hVf3Dvl8QJnZwfgPb0/Syp9Qe
sSohL/RONh4PdYv1CaLUwREHz/ah0wCq7/7Aat88K2vg3AN/KMMrDPFQ3YqX
iR4U+E58b7ecqxmk0Fj7Jm2rgcLXD9dSj73EwPb3U8NPXjNXY45Wa305C5E0
1uHp0SSQly5ogDBl09KkIDebbOIQlqVGWCXifAV/E2WllhSIjbcBe8Scs12X
/pG6mYnzZdWJPYyh0/f9hhvgGJS5+hbZlbNnw1Uz9LrdHwejBI3L7sCqCZDz
LV4Er0/ZTfOAgLlXl6QFSWeJtlSglZzNJnqw50fZLaYQ6UlcaLgtnCsB9CHU
ZfmYOMBP/j4CFDlU0V03eThi8A7qQfm+/20Q+zeXlXIS8WTutlJBpQH/c8Tg
I+UKpGK+wzBzq82Sb/L95mzDVofkbTccvOk0zhkjRPDvsPClVF7nAfDa3+G3
FVybp6mlQRk7zbnkyew6L6XISNVVkDgUPyzyrpbRWUWjIDgAcQs4gP0BlUmI
aw6hiKQxEh+EvZ54XkR6SZGIckKq2uXjU8Hs7aUR+p5qJP36nmbvyEsV23yR
CXa0AF9SD4ZZk1t7yb+akNQWU1OYipeY2QvRAAcWP2VuchuYPNFcS+CceIjk
+X7Vmw71XKNPELU0l0PF3tJ3sAjsjwJohyij2Nh4vEfrszn5EgSnu/+AOWSh
lKgvefb9iexrjjJAYezwbSNFfuLGY5LBINq4rwBkpFBgQMA/kMDRtM54zapx
oq4FdzaVIua6ZpaicPn+DaYl8Z+AE3TzO3Ux1PFzwkeo+2wnG+a1VkOZILHn
xu7wvcRaJ/gT9b//pihxF4Q9QO73uo5d37C0Sz31KHJeqkyNe6YC1/i4m79l
vxoi546/yaL7sqvxPEoQCfU9kbT/rIoolLc0qzHlNsTJ2elnrQQvjD8d+VhX
z6mfhrw+1aLKnzySQyZBeGP9gAFWff8YlMfftKCcVP3wcXWy3T9WjTheqbzP
GFgip5DkCqQF9cpNzegAohp7sPlwNv+Q5smNL2ucuI0tBM0JUgVX+Ce6uUYK
igXElZcN+RmBeyMVUoxHHqLj+xtgnO/jfz8B0yzJLoVbdpFYKiSDz9CjUcGQ
CzJb6CjljNn/Eg2glq/lvEwCciw+Y2e4rNSwbsQCmuamb4d4KxDlNBqi9K/2
/xkF7EST1+1/udRpqM9+40QNnHM1DqbmcDEaNtumbGZLpHZJNTTmkEW2MoCm
VDICtOJZndQ2TAf1/vk6ivU1uUZPc/WPD95VBMcEK7YomzU3vzbO21kF1O7v
mLgLC/Le58Hw2KEO/G7bznJ06UtyAVcHRGS21Kq7jRcdFaRe2tgMprStK2pI
IPLKqusne1ZkEZcDqTMmqhnqUhRntjb0y9ri7Y8E3Hh+v/tE5Z8eJX7+Qgs7
1YMhhM16WdVTVZGfabSOAfcGsiZR74myqFN5R77mQiPDcmn3oqPbH0PI+udU
3vke0t/MN3Y2DbY64574zfT8wF2j0lLws9wC4FGjBy/nvXqvYL+tN1YIao21
nQjBYFTuV1iL5P6aTcBdZ9R0tLIW9AnLBU6x1tV0k38SEr9Wf6a22rgFKdys
oeE7Ihy2EpgWdROvFXPprl75Y3ZAL1QaNOndN0vtPwP8EDO3K4p42o1w2+0+
0N/kaehYN5lKxiKfQ5KGQjdJFrWej/YiCm+Y4hZHQWp7saNhJjlHJEaa636l
+hM10CCn+c5eO97s027N1EgydVdxoMGDkh/cSW1eViCuS8OoCWCdnZbCpVQ5
XDeF8iuxcf6xZajrSfEU80j2GVIltx4heH1mngYRd+ip4uGZzcbJvz8ZLJFg
nxmh276UsDm0NKD1dV4c9mrjomD9wvOVl/BKK6fRUFBqbrtXEMKW90bhK4o4
O9Bg4NOj8MzzrYe8EX7BoAODHnlsd1djIt0ee7M9OWiNiWqpFHhqZSrT70Fd
1SjiZ6CHt9tfjKAqXkalT3lhlHtfEzEG5o+XMkDXscZMUcvF6rMONcb/Jtls
WwTol7jXOgl3WYCbTdgjLEImKkOj847xP3w6DFo6yVzO2zJRYwzFT27ZABu9
ykfkNA4US9kjCJ0I0NlrIFtm95+L1KOdiPvzna7QxfeoENvwaTMy4gj/JIrf
/jRzo7vrDem86vMB0cuQKTh81AwAS4yVk549eyti7QJg8SdfCyP4qMNYufHq
njZUgezsG6M5AEjfyaS9UMgl8H3Nwgpa3aCkFTVTspyj6b8Rfh4XLatLv3ol
kN0seE4yv8UUkf/vQV2+PDjl3DuzSCCswI9mRlxTACxgjPDTVxdcnuwa/Cmd
QkCsOZ9wZ+AknJzCk8cQpFdL3mwL+pL7u1D1csoT2AozwPlGLEYYqaaXln71
fiCouW3fMnBraCrEeJEM/G8Swkj6cik3WB2JPPtYlXRKJYM3VoMhlOZ+Kucb
bAdxZriUl1Ew+e44DX28R99P4Bg8nfQ1ay5xCW6M5xkFrRsh/GT2tRPfy7Q/
hcFe2hDw9of+FCYBqemd649hSij8YgECr9b7+XEQmH0suIWZLnep3i71as83
nQzmJKxvy49DQzIvMbxgq6k6bhNaY4dIfNyDMTEoMt8hMEfchruxCLQJTDxJ
PnAqjRor/Fu9xUgnPUTJ0WPASSZPpUbvawwTTBlXhfecb3O+AVFlMUySnXoe
u8QRhrkIIqIqPhNaX7u9tt6viLIUbTw4RN9ZKWBm8lvA1eMsz2R1pOWQC+nR
Ly0KIogPqQzANCuZOp8wswVZe5N6d76bGFlaIv2lDGp+/zVxKEbE9MUbiE2I
Vu2U3Jiieais/6KZkPcDq84R+5tyzH5EwJIEcg238YX7HvRHjcv6MoAyx1wW
HfdJYuSzuQ0yeWpYn3FeT27xQ0+tV1rtZ0By8xXcrL4t7BnjR1/W4Yjm9aJR
eIkoPWqtpzJbTRKbBZa9xUSrm0EOkIVWbr9zu82Q6PjugzofuowG9IKSQ5yM
6gZpOFWjGmKGghrGqntzAsOwUnTGqrudnwp358DKSofjT21KFN+QfWiQpt4j
knTvsy/L7lcERxtLAlY0VVaPvgEK2wFJwfhrn4f6Dr3q1ebE7WXmJ0fpyoN7
bIa0+F+p2ay2J33KjJtbN3dBq0CnumsqzcFh9PRcq76CrAviozn8cC2I9LTa
b+xe6lGhe+FNN5ho8I3CHszyXfufwiYY4Mxh6j5N83BDKCeXnKJmxNH0NfLf
RpsmKiRTPBBXTh2Fdcklz3RCzFHlpPeEypqpIsdMfjBmFdoiZbIfTtRKZjj7
8UlqEjlWSo+dCiqPZgJqh5D/2HgVy/yzA2PdaSDR2SQphKw3wAKy9Z/cqb9y
eGINPfEAvnDfor1qz9LE7q5a5WMWXoRancZVQbB5WYyR1nW8If/rdnDH3Zaj
64ETMR4cy4CC6XVdtb9d8lUQxx7in69+5F2Dm8NLfBg/Eu4rEGXYsrPaBLwX
pXjAkPt+KVCArOUIYjdPUEdF4pGQ6p2nUu+1OM3NK7LIwR8EulECj6S8J+/+
b5RRMb76QZOsYSDVqNlgoT72Sa6a4osYrYjEWHVXiIYsTB8U467h96LOn6WC
9iRR4s+SEjtfEUVT/7EcD9PkFWntql4wxDoOCGHSb19NmBQiiJf6RtLuWefc
vbt/2mYrBe25pWMQRNA+QnZy3X562+9jjM86Lg9i3w3buKZaug6Pz5b2taAj
0ENUOkYSTg8+BeiFhD+rcbykBA7eZPIUXaVGJ6WKdRZOgGnDPqWmYqAHFq1I
2jv11cnXKinjlpoit6sjE6QKdUf4qYc4ahKH4OEWvNhIc7ivFGQQiBlei+Vl
o3s3g1tizUwBWZKUJIodtHyLyVBZ937rX3X0dkcNTlitUrrfpw7Q/ZASg1oN
SpNH1HVuK4iDgYSyoyJy4G4lyP/JXov2T45hRtEEwr1M1JlylbIYtNJFFth3
HVzi2+EWTGqrGVTKXZu053+9C/Oagoi4QrIwKDKolbqQzqIjB0GyLs7WQ2eT
NPbpk5wWHa+ub+W26eFsg2aofn2tn1rWcCJXSSSDp68C7Kx/0V74LKLegcYg
yK74ukxup0FHmJa+Hd7vmP+NH5+fZWjqMg0KEn8aUMc3a/AbxOqkPj51yuWh
Fw8Z0DZNu0onmJ63DceOIVmb69wkgwzRkk+lZgYU0zdJxjeH4UFrwTcrvnGc
JK/98BN9+Nky9xRwYqvUK3PpGE/S6JygXNppyV5C0Ioqw7Q83Bfe7qGnU3cC
Rj7dgedFaITgNhEuJRInFPyDM2lWE2R6TeWYZ7EhoybFXLQmgu4AT/lOhcM5
+L/EJyRfhCKH+JJPdwj4KfggW/LzHM0hYv+v+CyGhdyeVfGZwLrlGu41Xr6G
G/pSFfRnyw4Rr2dK0ZInR8WM6dIfWISmG8QYIThpKt78q3R45nmvn/fbmXUp
luvruEzJQvuWG4puX4Q8iqhgKvYlNta3WanrWK3H6qoWB3iFU1mnk0b4fIbM
lOeXIFrE8EprhJ7NMZt4L7/fb2+isPbp/Rv2f/I+SsDk83gUPEpCWrlnMtvo
duDHV5Ut1cjTnBtJQhAeId1aci+p5ccZKlIlob4kL3BHTapHEdPxiITOuh0s
dYzIkVlTrM1pyH07J7kL6KcZURIBX5Wl23lvD/4CTV5lPUA+rivPijeLzHZL
qKL9jEnScMDVVg3AQhR50gJ5F880ScXGIkDt/xxv4DVCRa4QKDEDrO+JhLW4
oDLCqmCEUkJiMDEU23i4x2J3Ewq9k+UzIf7I2nK/DIK+h54I42N2dtzYKmn7
wiMvrwEymyFHG1YtBIjubx+BpsCrPCuapzN/w21UzdrS0ZmhCd1OonCwLOqr
3cx6vvsV2HDV7hMkgYhVb+GL6VRSzVDd1YQYugjvRqGIfH83NoovMutyRVl1
XbvFWXwdndQRbrSilqXClUNQfncbqP27ZZ5waDhzHDFEZWh+xCJeT3gtmCNb
wXLMTcH6wRzfFtTfGXIKsRbWZYPK7p/lo4B2+feINnt+4FKnF4SvMHZ1dRZ6
TrsAQJ5/44kIR+VPzUi+0s2A0+UyOpKmXCs0LgysFZb34NscZa3IFunbi+0J
rhc7wIIVpQSpv2KFHO+zACcU1PXBjavLj3IjRFzGkBAuRf0+4oEEUvmmFyBr
8reKCFK1pv5JdmJtHaK6nkKOVZYYqF+TQ+e/zRREg6s8ztHM+eV898VPS279
PIPWHLwFe39jP3ClMnSAIT8ZehMTEleiyCBISvh3nuNuvRs42AE0mUUeTvuQ
NrxyOq5SRw1Z2O9PKobl6bx1MeEq/eXxmrQyZSj9skLTapR7h+mdUEbt05BU
6tqif39GZXDhZ12Ptw1pl1xSjtSQB3wiBXeekw43I9bXJQz65ph7nsfow+w8
r1/EDa4aYj5iPkbBzvav9AhglaFjg5IzoxfZeCuNgg7crDPS5LdJ3aK4a0/G
kwoVf4wkbSujq7+XWHFOx4YyhDnBiGmE3LJPgYhafhMLkh2wESMJQegc4QG4
zSgxkkyV1+cmQWdAmxd0CLoe/wbW2Z1j8Kjeuut05wRqy0tg0Zf3sYV2YMY3
eNMMWMEvXeS/QZYl7X3tTDnypTAtr1mgzXN/WJuOlIBeChltEArx/tMhbp2l
AYehfR06xtLS1zMvrCf9v7nWYTS7VjWm5xVImf2wp8/H5mNe817eVdD4O4Vo
YAMX+X2K7bXUw6nzy+mzv9TeoBHwhkRyvKUV+bSLRsTs2Hsvfj5bb1B1kxCC
zJXJ3WnT+DR6eQbSFMhsImdZb5qhqcMkpwvhoRMOutgcK9wLJbcilr5L0e9t
xmtbQ/ugNfFEKKYNK4UZS5AJzzgo1DYEReZ7In9TgoqeMtfItSdfnQ2O4zPx
G7LLJuPDWLvurGLFSN0BimUkNDKKP/7fQ8O8yDh9CxTxIjQDGcWNyphkA1c=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1ITHxttW4a9NAjvn1ioEyuysX+oonelGQDdoTWCHA83iW7uhhSiDTrE1PVgUwVrXG/9OUCYuvrKaqMfuthhuNVYj9spCV5QxivKrdty7/2RAwv70t2X3J7JYmJMVVK4msP8fCjHMXVCyC5fonrUQUEuqgu1vpvPeP5S0aC4r+00JktsUZYPyjyuW2OJaRWuIROkjklf0R5cUAGM0sgXOFukpXBeIfOcPVidozoLAU8rpu0GY+wImXCmbKCEzUdl1tFxS63PhhVNS1MVHW++fEca1t17fHScZiAyRZjcmpTDQo0YR8hh5yfnVs6VmgJppvdXp1XypqalQFrCSnBRIAQWs2n/2JqGMTMRFh+TKZ6BZq+L41ix3TIMe0SHGsXuO+7DNh7b8jU/xTNZB3j49rOuPB/StyoMwp/r1eyUEUJkHtxb0uZ5nQFCEOtfi9Yfoj04Uaj/6U4OFXtcgjwjHS1IZ69udox1Gxpba6CanUQwAulsHQwpvCBFJJQ0sye05aWzyRnKDW0McxFsLE+17D7TCOYeOfulfsAr9nLdU3h547Ep4FVquOfNRTk4jg+tLlvq5CBwpqsxBNjEJDmkJuQayces4WRvkBl4k6mmAxmPqnoYJ9CQKP8pTnXL0d+M8sYXe4obm1BvIcsq/hSwK4JMJUHmDwsjV2jGteXuwnS75qriynDoDg6FuH9PZwXq/CMpXdI8TES+ktCA6ZCoggC4bSMFg//lGJihmCfJjXz8s88IQUkyjfwCdYYEvRCFNm95DFBmqFj9zFE3xaEJCA3p"
`endif