// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rAmWyThg58vmHT6umv5/Nn5Pq8D8hpFE9tqDr6gRmqW5BFDKM6kR6oMXEBrq
5WciTqgW9tEt1D1ebaPRMxW9Ry2lps06ZbnHIIamWhUxNawo1GDxpovRkdY4
tXpcSID1G+oAwyNy27YKDcv/OhJyc+HpLBtFOrYbzlcGhmtdhaKSScC+OplZ
DudoQFjQaAnrPlFXPmL42pqKnSDBfWnbeEfxMvrkTAiUsd1oOA0xSV+ZiPhU
f6FtV6Vp1xapK6b3zLvDIDMgnYxzAWcbNzv0wBiB9cFF1NbwHjwdT9Eye8OT
rMSVzntXnnD7EJVy60LOWidnN7usqzdQ9lHGwjQCBg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kWzLyXvzah+OeXxQToC4rn+oOSEa8xZxEHaLD/F8MoYupTuvjXv9gpgXqi/2
usJX2N30fZ8hC7uE7StGPRrja4yWRu9s/6AnLw2lG7SzIrPRyaCP9dkbcUkB
LX2hLZYmg2Uvuv0nmeNKNNrJSzxKlo7T3oMCEflRI5GRM0aIha+k+oT86Bw7
AB51kkhKlVf1S6UZC6yxaj5wcfqSBWWpJXIAFg0M1SBAPBPcm8QKsowdYVBA
XLxJOSZYHYxIjtPFYwHzMtHxvHlkqErn1WY0ue1QdR60dsPRzIA77f4JsVCs
8R1sFFaORPBsWiYYsHaPJuwP0dCqCr6humvzdmI5Lw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rauDdy4Tp2pP4hyqDY2DQvcBbEGB3goVdtPJxPM4RjD62GHQ4TG77ol0oUUa
kQfwe92QQCcMYIfFkv8GVkRIXISd3ylDDxIH+XlM/Q5+Yh7dzJ4WuCybai3p
NZCA9vJD8HGia4RV3V8jlt+F8wWm2JL3KhX7GoKXSM4bTBZAWW3hHEgsHsyq
jwfxHwXv9Le9DteJLuWPmfykidXvW/A7IQZ8KNR2z49gnNj6V9E7z5q3epst
PTauj/C5D0e/fM6GzzjHbbOdoAOjU2JBoUskaLCIKtGI6L3Mp99lA/GV0Vhi
ER5HBtn7sws5JW53D1m1egjGAJMeo6/WamvvQT7wfw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aqYkT/Lu+XUxA2DqREcdGWKkTY1FqtVgQ0jpiAKZc9z6A1gMqusDMrGhooBx
woVMfGBFcoJUqfrLhHAhCV/faO638EeBdB9B7VLWDPst8+RbFkmTw69hKPk2
v7gGi9+6nIOocutsvlYtdCbG64LWLGq23RUydMwz5PuswjwB76FVuxYmUjB1
t1M6nStK32X6yBDz+8nXjc7UCdcfA/kmsiBLZh+4VKNI4aS+2ehS80MIwx1y
VQz29XbtEODhxoiWieTcjeVTiY4t64TzoA/x+sWZnT8I+XLRgc6RL2A7scFc
AL38T9lydkfBeE8hj+EYBqNdrUouwcV/3FgIitwr1A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Maz7r1iKJfli21ib3RPtP4DHRRWXUEbgrHhvMCe4X7Zw+RGrcEsDkMpL1t9C
1Gi1Wmco/U/Z/xbMJBz2i5gtXB1FUWoCpwHuBirTarGacfCpxPs+2ZCJVlX6
1AqgvOfsQyGXxX8RTGxhtOcaTWNaRqx5Rw9LhP8i0MZXaq7+oow=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wbgcpO5VoFxUb4DKDurU68oDfjKCSOcrx65rpEQ/MHtXAQTSMNNuKrSta6CF
R9wvam4sh6NalvWPqNgEyJr8KCbXnbLnkrDJStka9oHG4QaoSKAB9Ms9wfmX
YqYKBSL60kI1WvTu02+ykNDj+EIZdGau75cX9pHe2SycNRUzUEv4C1RFL3AI
yUwc1Hr1xwc2/ffVMzOS0EG3NFeFGDsaQ233bQiW2xLKlsyqThImDgRntrhd
pQ/Ls0EEynu1Qbej87Iu+Z00jw7JdktC7gR1ocAbiRPtH6DJq6DlZmla/gN3
SRzlipnKZzLa04JPo9HPy7t5ydEglxPSCtTIMjbligxl4L9lHSaw5ZnnqvGZ
j/kI2Eo3FNi3tNlShWp4SndlOrZUugihDI04joZrVBiz0oaTnb03dlhgb1J2
FRQTJdfk0PR5gRCjpgxgbRUdkPjomS2AXXGbs5RlLzEJbDgaU2YUqZroRlzn
jbtWa059yYFTmHuXBXc7XLda7MhYSLKH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZQDLQncGljNuwWliTQ55Y5419HnEkSIhN/93pfbDYnrAMxG0XesSVHElcqj+
FiTx383NscFKSyY2QDGf/UwX0NqHz4ABN9tUC9mM2v5nM2ivMc3t5EGVbFS1
Gdql32uXsFnmM0aFht7tDlRRQgPY5RaznzU7XGMFO+/hHZgHwRs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
baRnoEM1Oh+VeyZwosAMqesIWU018Yv6LaXEyxrFOOYDTHbeWedSm4iiQjJm
j3jNmm6EvBfCvvRMoinyvPNHg4/Z4eLdiin8G+elX2iZ8EbBjk0eVjt9CRDn
myK+W4YiWmqd1vACmcvx/XAAZ4tdKyTDZe6Eg5e5af8Y0RDCsNg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46848)
`pragma protect data_block
xuHVygVf8yKxSbMELf4iZzr2vaLPbc/yrpk7nFglqS7LbCGEKjYOdAGO/Zb/
qIj8N2amyrvkZPmL9Var9SRvTy76JrYP7xGh2BHjDrCXzL68mM+C0uLRG+Vg
fEIgUwlHX8fNC+1B/KOSWvmm+06/PxpU4nACM6K927/1/Nn2/RvCL2GfWabP
SvaYd/M5s12V/40UpXfUTN/xdgGym8tgw5pKs/hl8VRr2IKGNguqfY2aGnyq
DvNGdLU1iDoTJzgsJSc8y4GXcfMHrAOk7R6umu0Kz0bVs2KRF6olsniZcDFo
Dh7hUxMDEqBtFeqV6joaCRS0PtPMmOvLAprloEQJ62LgW2v5cF8cW6oTLU5q
AsgEabRFero5+ABcIN5Fky+hOsKpSS7UM8TvvkaoQa+paf+8N9G4OIMyyG3Y
OneLvWLevQPkKR+Gp6298AiE2HRWP8u63sDxxlwXyP7+Z8Ws4HpQT4h/KHvD
WOPlY8R6SQS+8ySpyNgGhFTDTOWMAshPp18RT89sIJx9Xqrug30VoLOsYWOh
dOc5BShkAjAgyOYmNglHt1iYCKHWeHey2f1xTIk6oOwOxNOXqLTuglhqxYbT
RYnV+N+WRmEWsvNpHQBPYa6PXvIIui9qOp253t3ai4DwIoeyLeWyKDCuKYJj
8nXQ6tiGRqnVBiCNXLAxJPD5r08PSHPlPNq4OEUifcxxRCtb/+QwzhUCcFlH
fCF8E1x8nDecZyMSQ3bmzvVYRx4cVXnaZenYcz0cegMTMHiJCb0yau8Godes
osvq6361ALmzUxaCSc0Y/OPGhdMkYmfEuBjTkS9euxJGEn63B5zrlGINH0A8
r2X82EhcUNJsbRu9OxebCSMz/EoBeHrKp3tlzPLyvQPaD1EL5q8M6m6ul3sS
GGfGM71uXxyzhmJe4cvlWAWqCYIcSZ6MkIljw/uGE7hgcEKNT+t951O5hiKs
nSt9jljutCDOEU+cIIvABla7BtdUODhv1qCL0D8rz3St+CRCx9pnkm1w4e/y
VqB/A/eA60Iu7JXX6+CiSrhLMOsHgllTWtkN5ac2yJrC19zryyIp5n+hwnyy
lZ8cz4FwWys83yJFdESzW15+51CalvR9xf9sE4LleIflxkF2A+ANJXS8MIRt
zOnYeGACzNNuBPirflBNejDSY+/YYyl2gLLkEltqyn1WXV3+S2vt1/mKktiJ
ADtYf7m7pnuJ446SK1A7NMljCp9ODcLHNfYkKOLvfeKTA2AohcOOGqGTMiBx
SOHWHn8bnGkJ238J9I/cMkzE8UdKzmDBlrR6kmFEYtWdQlOxvDDRXJ6pTMh4
F0nn0b8Yuj7eCvcmJzt8aADMzf1qhvghd93UEzW5L6QiC2Jm+vz0BtZh0EeQ
6PfmGXcIru0+JYjiT2YuxzWSF/TdCqrezepKSqGmC06akhxXBYxO7qoxOwdG
gevwtVcu32zT5D1CvUnMzYTbnwSj82JAF/sAk33d18eetB1q3KbevmF7raUJ
0Ju9guBpvgAU27kPMtapxi2izHJKdz3Eml98yIzQU+LBXKRGu+yo4Dc2zP+z
inNaYS9SQ/BVUd9zvUsCuhcRVFR2pPhbff2VVjybIsHOFe8NIBHr3RQocTDe
Xyni3gufKQGG96NMb9+bTuQBRJag7lY4MSwRA+bVCEFcbpqdpkk8qnlCgqv4
C4w+Av4CK3j/Qr2Msm8AGRP2hlVV49MLB/gPaQjk/DcDCM8a16d5bTagGk/E
dl91BlMLMY41eOUAh8EezemNv1t2WHbGWC2VCovV5Yx97Ds5hwB/MrfX/QUC
oDOfySvxpzDhMtqoWuUXteq9KeBZTKwgh9+gPAoEIOkhLwI5k/I2Cyaos3bV
9RZIsRMpb0/kda+FYbC69qVegxZpebSPNu7PlqnVclFnzKCtJdUNW0fTY3cp
/jjUbgsXqgxMhZdhG5U+KZLUXDCa/Zo88STShDCmTHbjQajCem5Bjdo9gbJl
9x4/M5UNWf6QQ01lvtoS9eRbS/YlcxBXYyRVgo5oSklVNX2oEb2wuM6mb7qQ
lfxRVad/JlX/f33gb4rw6fVl6MmlaZkoSAHWLQwkDfTbplOFVOTOU38mZiEO
GhN56ohEThJASugqtgy+fHQwt69No9FbNA1SuqbaoKuxXRoVMhhsrMVWCjwf
/ubkvuvMcV0GJhoOOIUoXALLBaL80wnJk23wU6J1sHM3q5e3cexUvCYyzFEX
BNXgyYPiBciFXmFU3WMBJaHnWL5cmTZrEdJCUgr0LK7gCCukV/fywE3yq/UW
aWvHsM4zfpYc3pGECGcw0jIWAo7goJgPJX44FK/KgFV/Vjs8yVhSpw+8zzyj
RKZO+X6YPmZJilshbIjPV5+C4D/s982vEL0GzaeqIqkveH1ohXQCjKzaXGYQ
953iYxenaazpamq3e7JD0yx6/UlOgKSMJqlqi4BYYYjcDFr3w5XZfPOOpd2r
nphZuAeLL05E0RO7+PyHMzEQKcqNWdfDVbVJ4acH8IPOy3LCOxZPuLrgCIqH
/PgpjSGcH2CrpQ/Vwi1zy64pJl1CHvHQzSwLArCbGdbreK3hbcYCGACo8/R7
k8HSbmumJwn5/6JhVnXXUNlcqcy5YUt8gI17AQJqiNWnTMB63wNFZgCtLMda
O78CchA9GKL1crVF7iLRDIaMatfxccD7K0N0/fOU5m/9i+IN3wvzBdBAq7zD
B4tn+Hsxj17sxam1XHmhG48HNDa5x/GRWjYVjdY1jlUaxah2sORKMmtMOpnf
PN7BbQGDZuQhNq5Jw0CCwILUcfGA8SLVFIqJr7wr8WymtBOywB9z9KUAbESg
zVty0bj0y2rHvsA2wueE8ozB/mI0b6aaWjQ+vUq01ahAj9D33ayrrFqPw7nz
cT3wp9rT52xMJzA5Ba/RQJLK3rlC3ULDkFYTipkFT/t0e7i6K/3+UzQelKhX
CAFnCReTwVkvI4gbwXUyf+VPqEAFnt5izG1z5Kc8p+RWIlCTngbtgLfr787Q
DsRrgFR5c/t6sNWItVogWmCi+0TtQsR3AzJeBQ/NMqwJ4fKMc0zeRMw8dODX
Ec/7izkVKb5Q5MYFMH2umpC0iBxO0yma23AGDdDZnqx3rcbDcVV46VjOjBnS
pZbbHkityMcs+ytkwoTWqBliK+PH3wLHE2zyhAT8XCyL5lRnlYrVBAqwi3Pl
ThwxUL44rog6Q944Jry0gBSkqIro4sQ9ix6S+X36SXYYPiHXE3lfVV+OQew/
zE5Hmv7lBw+v5PjFJTNhE24vZ6XfVpLjhKsbx12HB+4xUIVzmAPO3CpRv1Vt
mfBYG8eXsEFT6Vd9lbmibUO4UPXzjI6Q9KZOR205dAfne0CnJgYYRbWpTLmX
6nwnfBU+AKpLDSOKLozU0wsFPSuebpptL+4MYf2hu0QfTcTBNHW+/QofSnuU
zzbdnujDAGbPEor5Gt2Kxp+RDGXsdHD3DVTFjRa0lBgakSP87fOrDQb5s459
TOK5V6mUfBmjK9tL1y+p81Ut9S1r3OrTpno/CI3TRCF3PE28dMfLF+EchZwd
r7HB+E/BZ8zSHg/au+C4DfkTDX1oziKVoTReDb9sbNHB5ghdU1pNPIXArvG2
u4Ac1E8AIv78N2jvau2kbJ1ndZOQEkOOQTdf0qj7ayqWjaoF59bf0QbDv5Uy
c/2/mx+8P6Go6m1TqLoxJQBcmCKGrhsxHCX3Hd39aBKOM4EkRSAyHrGoYf82
uP/FpuOuO0HaJpx/NXqX8LSemEHtMUP1h2kzJI2lJYDgVmzWDE2RGY4hhhSU
IhqqPV6im6sa9aUh27yAhLBmDyEClYeE08xOy9TNNUD+yzW3syeMQ1Mr3gQt
MsvydCzDO+UMp6c8Nr/1Jj25iCSKFyVQRlW2oYElJJcKouRrGYlhmzziF2Fr
8VtPRxgbKRLCvWbYYJBvzCAlE80UiOsoPkeIJOXEeRPrr8mLsPANQtjRsRMj
l6aHfHTNTEADolbYL4I6g6P39wivK6ejf2FbsJ9nKjxLPwQiNCkp8D1o//st
OSTYWmqKqvsQh6L6RwaqFHq3d62IADqioFcYem5H7/t8KjHRYJGrp2poDOVM
E+Y1nt9yFpWLCqZdmi4WM1ml9D26phzHEcvqlux7SslXLY6Qwrw/afMbnlXI
8RAuYx/HPw70b1PrdL6fCtaiG706zdhzGP1Ih9tiI3jyUy1jb9QNCIgLvnfI
gSMv65huUm5Gbj+PDgP6w1NbGOPUdaXhtiZeV+3E/PV1v8IXfyDHzmTz3QG1
F/d0nhsthO5Xqv1l0pg+SKtbc82b+d51ZWQpj06CZk61N6ZGJXc9u4z43QKZ
Zo86NQqTJYOkZNmPUNs1oJt/9ThrKjDhTTD21u23Tji5YW1FbehzFO+d0k/Q
1oJn7UM0u65hkOckopZ2FkHfcukSs0xqKYvFxFVIrf4nWmjNGxbI8O7KHykH
p1cf2g61K/B/A1WnUkAlaSx4IBcJ9w7jQHo8jc0R6IX+SlH22lhnS3TDKbVf
ZaG2grP5lZcIdZlSJo7iCE5M8AaCiZ6IMN5w4MDRAWFEEKSHt7Igkt5X4MR1
q88Jy583Xt+XcJT/h5cpezYxMzMcSQd5lccjbxKFxRnRlevKUd5onsSfFhi5
SHUG9NKXfEfCJ6A8O2FnhSqOgnz9TWbCewjEFU7TJaZ2TQMw9WO7AlrQY4aC
LQ0+VF7IkBcgmU5T4hVv/j+fOr9jX9jJ27mPhNmbXPjr3aML7F+AD6qMNsl8
4ssoJJZU2UebjhTPVuNj396+xOjtl58mG9yWX1Rim4ng6VpQaINoQVqGkWGn
oCz7FiQAYV+g+A4P01oSqMgC6/MBNSN9+yZpKh4rPIS8IOyrWWCYIGMXx/2w
lVq4Xflo7PBWn5MIUMHHhBG1CZNArUe1kneU96g9vHDvypgHwM73ozU4MTli
kRujJGzO0mFhDVDrIYe+9gS9loBByB58Kv5FCezzzIf3VpRW7BObwomwQm+7
4TMWwn4imasHhF7eF6k6lZcXCZAJwSQ/hR7JSlUDOuHFOWkWiHmSwtnS+xNe
zEh/46LfEU/WtE5HizIn7g94urWSW/RFjDxDv6sbn/L+PY+dcvBYRRNzX8N0
g0cu7V4EoZ0jMn0Gke5h5VCqMA27oqmLaLbKJXp3SxBn1rjK7MZAL7vlX2qE
qXbRW8E6uUptK/1LNQep+k1opLD4c4p1hg5wVTKiUH51Zxr6MH6AEKOGHOJC
rCxkn49qf5QBX+73IOwh/ZSrB6CWAOf3MswZgWjnfsvQ9L0O7o20a6XvDOry
c78GEi+3E/zgWTi1IiaBmNYuM8/08nTZGTuaGTV1KU0SWu1E4WfuB8sHxLGl
GKPCdz9CwanyQ8xCOXzgLHjnBJwLU750aJwD4VMuvrHy8wSu0S1nQc+u9l+n
9VorPyUbsiO95F9dsnvHjPTHvlc6BWekztagR3DPU7CN4nVvkw5zuJu6Pm1P
2b06Mi/iweBe9u2aCxxF5LePeOrO5dRNk3UYkSU4onAavTJOUgnicRXlwVj+
MN1AcaS8BTP/iqspSjGsX+zGVKHlWly+55zdqwJBnSPmxJd5eWBXjHCo84kx
ZGdqE5EkKtrGqjkR0L8dkFRpjcIW+EfWLuw7R2HGTvjqxOTmm92KROmEzOF9
Tq3Ig2DqLhG6G76zuhiRM6dy+YWKkTQeMriew22emeFGIFzvVyWyc5AyTmd+
rDGh3KeUqCXqES53tdLxJ4PogriLr4wq4Vwx9DE1h/mMGnsTz/JF52A0Cy77
Jpmaftv1suAYbaI5HIe3MSWQybS3Z0NHz1Z1tCizfj/Q/qu8GNutC+EGpz3y
Y69RMyJc4HeIn0DsGmO6J6zFjMM1ACeZa1i3yJRUVr0brv4rlPEwB4FXHdmy
9wrvKHdIVPenBGgJVJwdnWmHFwV+4QVTxTt1tzZUmTdW5MBx/AXgqaJbBLQM
U323/FDhcdSvHJo2uitTTHXoQJw3e0a8ro1yskJBVGJyoioDpx6sJOZICVve
DW0Oz/UnwSBO46BFAtTYvnjag+4rfI5pmLh21M4OUHu1zATVaLMoOrpL+5zd
wgMvHp/wJ3jAG0xdPZpwa2gxxMdatYt5iiMELuKfKkIJ/ybO7nYYHKdaOzEc
UnF77B5b5v+o/GUO/rvePY8lmUTled5LCX8B7J/rEg0/b0cokJu2hx4DL2TZ
domyStUD/Mu5LElVNeD23wqYjmLqdKyGU2Ta9DROYQu4CTckQN5r8bXA46Ve
v9qk56t/s1HTSUiHyfMNYE16LnfMRZ89qd66jYzHBRMqAXdQjUCwN7ZxPYwj
SO+jzTwitr/An9fqwXxltfDUq8YRAhUJHmnxc5zTKFGXvQKGmIV94ezO9Eio
jRGznGbtP9fU9BzWX2Apu8BxldYQzyb+EXHNQyVWUub3SzNtJDFKOOUqIfuH
5dPiMTjC8nqba4rq3z4OBz4B5XHUtXm0HHgdDyBSZlJztcnOewSD3cuMCSeg
3NADU0mPYWQbDACoagBS7ggOFY5Wigi+TPovKsNH6n2zUZ1+ZKyRq6s6ez8+
kI8E1SfpqHOIJcqWQlBTlJut/URciSLKVBfePGQ1jkbZLwyGsebxH49hFrEn
82jUvGTtsS1hTUnggE48Qqi86XbWwpRF2reyh/7xDX/j18jPQp5FHULpBg1J
BjhjyoIF1PldF4PJ5OTPAV2Mz38/hjqYINqHIv5zLUBRRGhA87I/z+LJe91R
LszuUMbD4sDwSKh2zcojMPbPDAR79e211TJ5xqCAJSq0N9pKTUIEK9z5E3eE
GalnufCb5UMWhqLdlr1hvGRTNZBPWolRLdclYkXQWFuM7fLW4NA5OHkseraL
wPA4nfnaOEFjGBJ7PpzJaUU2H6IfGBhJr9C9YRR+rwJIN6wGM90pktKg4nlZ
jbUSc8fOWFhsmljA25VHp/PBPBU0iWwkj/Ck+/3pkwCJhu/mTv9m7cadOq28
6mW0nmZb1cgpNWxaLlxCXMmvTxWbuiS619PHTFNwJAMVnxW6NiH7HeQ0IStF
KwmgzfB9DOGB4TfHlyx/v74YBGk1BjF6yznuLbB94A2NDcQPILAaSSpuZgNe
6cFx7YtR8dim5YTYUlCSUOn1oi1fBhzMOzJzU5adNBpf+cgxhbeNx0EZESfC
VpWWAWBHmYJoWQQvf27cjLgDM/WCDwskUeEjAqFjyoYN+ob7CUw58pHWeexw
sOi732JULJxduOoDVIOkkhbeJhJWBgW2fszH74K9QFFnF0Hc7V5/5p0qZz5p
9R/gbrpNn29o+tkboiJPoQpkWWxWUFj+5YSD/IJanI3vD4pBBeSyp7UT1RiF
SIu0gRuhj36yrCyE/bORy4MR8t0e7TrO8T3P7C+dzWi2wsiqOkUojKoEOPsZ
NOAQu92z/JGX65LW2ZICwEKsNQ+wNUXc7TiNclDPKTAzgaHbWz8MZe+A4wCa
pgjFKQWUpazsQITZdEkeJgsuafyuCWgeHh19GhHv+aDIa6aSW9NY9sD0s6fG
HkLrsBkj855RLGUcq3ozQAisOAneFMf7htPnCoAX22v1EgM13oMAR6ythlDh
vn3yQ7BMRwBHFl7Q5xmJyd9FZwABStEo7zDjTdb7lHEXE+IXSkALYa09pYpk
TfMxvxQG/EUP010jdIP2OPMuHhcGeutQIdmy9h4w8nILYMYnqU3yuRv8HAp0
SzszC0hYk7m1EpH73m28C7/b5GjqnIwaEMoTsOM/Jb0KXZ0FpHH1DbVb5iaA
GPxGpkHPd/ejPZDZNrtr6o/4IxXEcWutgKCpEfsq1og5C9YXl5sF+v1/ZcO7
9QKiLsZfu879ndsAadYO1QlCbh/wGe6nGEfaxyHFwM7OyBcruN5wSvSGoGCO
79J3iPM/N5ypeyaULg8tOFnbo71AvrIC9Q8UEW8QE0NNtxJ0YYtQIIZLfB52
UAzZfhQ5EHAjhii5O0XTF1eSVy4LxcKZWaW+105/4hcczF19ae3wytU7f4EQ
PkCsgn/ztmEmHYvzH/FpWngKC0ZJaM5+QSnU9jJcv5IGTA1clEwsZAzKKDZY
eOqfmJHqbmqpJkqjv8JlKwjIhJ20YnbvI74Zrw2XRa0q8bAUm/hD4PZ/XgBF
T1gvKVpS4eS+RqDLv4xU+pFsOex+hznxTmjTbHHk6ElVs6hzm6Ck9LGWvytA
16aSnt0ByrDhCnlbB55y5Zg1gGS08Eew6TRVnAXdYTRnCKvuPVpcgD8NvgWS
YS9hzRqaNSHKt/2jAmPT3jG4S2hp3ME/itMNcrQjdSEEi9Y1VHEgp5Uh3QFa
bgvDq8ebiBWxsVKrZiAnBQo+zbT0zTq05DdyFDd3ZcuHfIYyliHpjb1hBM9m
p+1G6Xa6CLS6MA6LkmbA98lQOCaxKePYLG5JLxNOJGHdOMkBFaQcWFelvuIB
ewU9DMNJTjDGG0YPGHzw54h24Y+96pcnpksDaI1cnN6+coQKtbgEkH78c9Eq
iLcH2e7e8OEdH0v0VX6JM6Bu9wfzreLy2NNtb37CJ2EkgcYjMkpujIngq9L5
pQDE+TKjeSQtdhEkqa/GEtiqNghWyQi5amoavMMWXghDnQbretv7SnWvqpzx
DyBFP+CJTd3v3F9VyYOUbGOL3Nb4f8y4XGW/Z92Gp7M05wJfYSuTLzqy0Wp6
Kod4a0jCtPm6oiQFeMrqf5sh6QxdHPL66RsAQlNOEsxgK/Qn6ynaiZg3/TYb
V8X/ATuyPmPmLGwKjqu33lHPlfJKHxfCkOEOnTglql6DhMRA1ToTEaYGPlH6
eajnfOWn55bmdHcDauhoDn47ULmTIYLPAka39eLcpV5dvqD1wssOeShHWCnz
oISNt04rX3eXRW++L/Jg+8pgODKF90v7nt3B3Caw6oN/X990nPuHG5PfxT0e
xQYUz/0ZHeMyP7wRjb05Zy1XXWLzvpLqK44jEFDXLjDES+LNW3BQpfqu6hNU
ucKDWorFsKAo6PuZ/xL7qtWb1t3c94dwGMN8h8T2aipKnzCr2Sy6ywYQ8CtX
JeLHYlEkIao0QsF6SQzC5ZOGgbY+IlrxitjNgZ9bxlne9t3p8rdj8qfCyoAr
sUEl8fyz88a9qRaAckIQwFPWTCVtBKHELd2B3bErWNj884lHl3NEVyKenfiY
YGNHmP8DNTSQ1n2WpmJUDR0oldXxhInA2n8IMdkx/lQ6lsxyyTg81uCFm2jq
HqyDneeamw8fmFQjNAHv5RNZr5bZBDB0mD+92Tx5Tt+uT7OLpQbf7Ml3jHqD
s5/x3Fq4sfbcyglHhZ9ym1jYpWi5XEATw+4TfPGVfWVg3vYG/sdnOeejMcVt
hKZyqKRkDN69I7QPLbs8HcFTgh/gKjlWKg5HK8TcN1vCQ1N43Y+QFwAs5c6S
W2sLbQWfEa0pUk/cR7pYAx3H72b4JXB5IZiEsNkwuWSxaR/etBrecpl9xWHX
vaSFlIgNS0xEvsZiXfEDJr1XWt9yWwNhPESPacBw/0ly/xAc0fW4Zdg/QG/K
us82g5Sy80EBfiRyK8bpk0G/oimQYODNISjxJw5tbjzs/BWYddXpxMvnGKzD
sn732CfEAzLX2qsyL3yS694MI4rq8eTfQA25CNXW4sVpoKOda7aK1Im+MM6Z
ZufGg+POlPyS+4Td7CEciitChVuZyePIxTozZu9sgZpvPHnJu+AUFcQQFNAT
94bi6wvdx8oh6iTcOtxDC0oQ2gZU5SXFaOCVI9PGV7mjt/CR3D/uMJo4ITP7
DMOz64DZSwsKKSqrvJ1RSLlO4GL1mFKIDvDVNCUYBjKyb/vtOQOayim2k79q
sFCt7UTQAdyukgvgqsYFpQtvEiCzIh4Yk+VaW1+CLqG4cBu/rObpQHVM3cAK
Ot+NcEFiYy0fmfGNZWIhRMWviOd20LPvYFsz0/hIUoB+cLCWE/lss79QGJdz
SrX+f3g6OD2aXZVmQUQf6Kn9LbBryb6sohjuw1FT9XoTZ/6Jd3OasakfH3lZ
BjzOebVI/MFgRW41pl9aOa9GwFJmFiFYD7vp+XT6CfQcDNmfHRZ+uFWU8mY7
64wFpUc1ZhSeybA7VCCy/UIXZ5F4+qcTCjp+doMr8TfoBw/9ZP1BdzTM4SXX
J+nHwWYrYsEGgtG2ia6AO23bM2ELRk8EByCKefQI87WhKRFKFcpXkSd9zoZp
0e/GR+Qn9Dys/RF3rYFSTHkVXPDIz5UrIE6Wl8OfiNraZEl9LHCHfOCMf3+c
ilyYi5oXCUT4fbEyavBT4f73Z80gqv6ZkUQhYsJDhB6RyG9zvo5aAIGD6PUL
UQTuT32zzHPF6HfXywwnygfur391YBPHuQiLyG2/nA693dlrn5421huTJZ4o
6JDTwNbnvucvZoXc0XUCRXSpt/Rc1P43Vn4xFoB5PZRlPBkuiiJaJJcfum+Y
647/AA7q9hu98PAv0t5labaofWr0T+RCti5HLGPB8bWGpROy6Uu0rwpwnAoO
Joc5J97f5MF0IL96MSJ7jtRxEHzxsiVuWBbQaKNSBkzARSX2BLCUJvXdH3E1
qFOUNwIe7zGjkix/MDSkvn4sgqVN20+ErNUVT1Ju0QxkwJF4XAYFG4oi467S
Q9K8I+WGuhQ4Rmsr4HMwwVCJUqgXDp7VHALLl0YtvIchm5BmNbgDnvyMu8IE
sX4sxKhFb4tThpEtvEhz+zrf4TrsKLf7bAeua1uI0tXoLoXoxBMVRIqxdULS
JqQ1FhIdgHgauT36b5GHLUsvBvX0dMbE+SM1bq82cUuMkFvO9/fQcvBQHkCx
7g55AuPdzumuYafm1135k0rts8FKWBoNMXzhfpw0IYrWSPDB6I69qY7cN3Rd
scuqkZI+d8rDQKGzmqNg9NvxRttITg5vBnjPUKHkDxNX9Lov5WJVjzyAMTyx
X6gmvyuhr8dELOzzUaORNpkyuZ9VK4hejKjajSBFxr17Ylvhw7r00RYex9RO
CpM8YI8SD3SGp59+ZWWWtVC3HxOPQGesVkZ5spp4qChC2BrdEITNG+GKEwl0
Yxx1NO1ycesX3eViYrMuoAg1ayFUP0ZSsyXAxNWDMGQVwrf3J6qlH5wrMD6B
M/oLCSua1zjhV3W3dJd51tkUpFvtDCn8G/E+Vidr2L60Rm0eeegGEIaRFOja
VookRETMovg8m59Dj3dkDsQ3oqsevmhJMMNzVR3+nMZjKamX680dXwOg27wn
fctBLephzDw1ncdqrtxjqFb1dtDhCIP37oJzIZaDUFh5rA5gUQQUI7+YKiPq
zJKdVYSHquDFJ+VcF2m2vOfathcWjrzet+rubN7mR9X3Ujfp6jgxk40llNSV
89XmGDbgJV3uX817iQVzxJgYCojBw/7VukbbuXJrEaxwP2U1wfhssJcXVGtp
iW7tUBFa+i8Mw2ui+jtub7KU6Tykji8on0A4wFRISMxfFb4Rnb4R+G580V/i
a5H1giwty1/VlOHKqXMTksfqsqx/imEpZXA+RGNggGyKeLmXEsVydCFiBar9
03elOf7Yt5m2dHljJBlAPboSwr8iCFaVxtYPTG/D3rJsvVEqEEH3K0REFvux
CXiXAfwOglWoco9avRwvEohl6zro8FWgwco8Lqohz9DJsKqyoEX9F4sXXilg
jMwTskkQcMaFMijewQWGcEIIecLRtaeHy7W4sT7gMRtoOOYR8d8yB+7efuwm
pFui6Y2cXPCrJOSX+r+XX2HkOzwzqWQtdIe9nngOdqGfxD4iqsX4nLue+N07
96g50L25Y2XPr+22KwS4iNZ9j0DB+N+Z2Z9gknt3s2NL0LHj+YDhUrULExtp
HbgRxNPJA8XzG/jDVjVNyNKXBVgo4hwjazCUZm86KVrhRfEEyh0yqYuh4OFj
2q6GV1Ye4iS9/HLMAQIbdrLJgQ32AUZ8C5dHV0yl/TObX9jn9TOruGj9sWtx
Zn8qBR8TjFrnhc9dGS0oKLpLFO0y+qQg0ygzj0DEKWV6kU1K0TO39hReSM0b
tHEGGqmjAayfcIJc+dQocyJt9WlUI6juUowqHJ/yICnoPjtaQtbRwyOzxWEL
45Z+Gsq/aoGJDmvD3DoPE7IFHiuI1MFf8AzhVDt09I0nSX7ZiYqbNszdcr2y
rFn8iL9/PikgZgLLrvLP+tiGddjdmYcYDXTmg7hTpPzstfJgYCVXayU6uAwH
R3z0inS1zmHZveWNqSq6OTAJ5wSqZPWTtb79Gy4yk4V8ChuaKkM7KpWZUCN2
ukSpu/hXvLEi85r7Ylu54qbqq4PyeeOmE5CQLb/z+IvCnsz+ukNVwDDimWWP
D2CTDfG3qsUU+jrvhZ0HPkhOSBzBj5O2SAihZOhuYvhcyWZxmyOr0tfSDTee
a8Ub3pxFwT/SLlh2P5ID0b14F+dPuoellWgCPJ5bUHgYteeErqaa1tHJOpxn
7fHEacqnU+oj3jQVrq9ySzJYaAX6qu5tZqtiK7VjxEt/6UsRusqX63Qfc7CQ
PrgrKhfye7FGmxO0fWisYnxp2WothXsTS2Xm147E8alqWccsuphEbUdV6MJR
rv8bMwGyMPaOWZDXk4heKm8TcQICeW+MdNJAtDN/NEevT2dd+CrbqB4zOR4n
xfszVq+kH6HWtBUr3q0lCZrMzKZLigefi8UNeLX718835j0Wn2C6l0iue+Wy
nKtx3MkQmj5YiEBN6LsLfq5UsOc8T1B9t8h4VPAWhbvDSQbKcuL4ZV3LTJ4N
XMEDD153XbbmzmuCSJzbNPeYUMW3anR91yYG4lpF54CiZwef/vJS3wZE1gah
l6Q9QNaVO/q4Sb8UuVCVdqvdMaTuNctYdTAKMTutusCarsTdOl1TZ73kJ1I3
d6XqL1Z9TOzKhOLVFPNZCRZJ3gf0EXc5Nyk/qChXEU5QxYCPC/rzs5UQ23u2
V+NLd/p84xCvaNcXEyZ08/Q2k+iLRS8WQEvuZEYsMlN9cTKLKKoCXv2dEKi5
/ukvIcK9f+M2GGjIdHqIFfOHKCKpqmgplgdECnnpjzwDr5FTL02uEdWkhi+p
7KH6a+mkfky8waD3lcILcPAPA8uhuDZh80G2twUC/93+c3Ix9HSNZjv1oUUb
K0FFykbBuWFFnxi2xPjD0S8u1vHtpf5RbSYa2jzDT0JoQLVO0U4ZOgZJgnkm
O9E/fM9GjHuc3u0AhDpE6v2+VrtlfTx7EJBv6ZJxT24mgWuGthiGXQrpt+Pn
APJUKvGupCETexk67lOoAZ++K3ssg1v/rcohan79nbjJ5bOT4JNXiC3h0zcF
l9UMeR2xpcWcapfwW1KPpOv+n9fpYX/yMD9WRLpbejm0U0BAXpMirisiYl5p
B6RAvOSC2KmnOBtDrSHkDxfALh1QOpG416ViepDk8gZuHG5k4nJdevLtjD9+
opRrtC6Ss8+np5PM5T5lHqCy10Bch3Qf43STK3fE0yvWSPRej/emqOjR8Vjy
tL9kUA+StC7WXYzmWqOYM9qazNvdbJYhUSoVxldpERjrp1bNR8RK9uGrwSow
n9xqK+zdbTLXFZ1rlD/jtTYpoFZ4UQetJiBmQb8Dpuh0L0M7DbQTyl9DadHn
JVkyTV3mIS9jEs1kY1YdmuCKYs9u099k/B8zglA/0QRxf8BQQc1gnxukC8Y+
E1yXGebSTsHfStrtavpIQHV04yDFMqnbL9kJ5+3eIrDiHeqmpbh+KpGa5cpY
Hi3As8qOVpEV7oeYgc3iJZl8YBfjoS3u6oR64BiCeSDmHreHVQ1h3KhwL2a4
N7j1YEK62AYFrj0J4kELBS5tca/1fpIywgVeTtwyr+8wObd+nRPE0U0sd3IQ
okBNbS9PcqP3BJPbXshIfucJMQjymSUwqR9mrdFDjEpfYbsGuezdFfImFBt2
Hh5srKUHx+592zgaDAjAgJ3jTW7VoFW7pIvgTM+hiEn6gAm7Eb5vEm+wM+RU
iTY7k4rSn2aEKfsND5gb1nxm3qqrOVceK/yYMc/fCNYZWo15KOBB6KrXWqb1
UFGYKrfFyuZsduD8sOXBSKgDHQr1laxjqw3+qF2a91zZVwsmkTaYCuHV/vmN
t/oj6v89OnDxnkvHYMB8vnDJe74+/tCND8tLkAmcxi84Bn+GBf6E2Vdd06rL
GYyROmS5uShdTxkzFAuMso1atjVZqhIr7y4h0qNX4vSiRGKrW09GlLD1JuA4
N8k4nnm+glaeAEN6BLUgi/kr+XxKRzLn2ow1OlV/RtpDS9NLBZq5+6fmlrEN
cfD3EM4cOS1KrAqY3zUy6GxIw7baIIyzyZoQX1nmw/Htv2aD4dKvW3GsOhpR
K2cW+Yt1SfX63sz1IBV27aQOvxD4UI28Qqx5OAGM4E90QDJTYKhl9r97dsFS
WnQPc9g3a/HlB1c6RObd490plY3i6esTi4VQCLr8wwrJNmoubiFTki4zPjJQ
/HITcFdwuabG0udqDJynqo5pTP5x1c0l9MZ6YwClc+QDm/AC0oxq5BeXt7ao
InfvaS5n6AhDp+wc2tdXVfkECo25M1ZnBs1Vp8Yr09ICrLT/0tl4X4kSwFLL
TiNngf0NcLI8r+h+Be5jhOab4EgyYHvTQ6BiqCHaIq7KWxAS1TfX0V8bNgrs
QRXMnvh7xkRwX0rn8gAFpP4rlCV855Kx0ifntGP+tIua3uc85nJjGLa2dSpH
eJqdsMzUHcyVfRQp/EjXlWNjgZCHL1vFTD0yLGb71uTXl0+Ixp8PL7pTBxI+
Yg61pI9I7lIkJ8qbRauvIkx8GoEgo65q3Y5WJfsO2GMae/OF0H1JxweOS7NN
EMaqDo+qgykSp2zXfr1kkM57l9I7JzJ7itUruDhWiovyxZ1F1XUYtClP1M+A
r6SDJf1ayPaL1DgZjAa5c3fpnyYSDXbkPLd0LOGDZQe5bicRffqM7HdNil7l
1OT83Q5seJSdM4GVx2V18BBB3y7JkJQfijuGQqdryL5gMqDNh7xEBrjpdMuj
22BbECJDlpeUKelr8AKNbtk0TqF3wi1gmLW4a83m7OJwCsXc6H5bhAep+cHJ
UgeT0ancapF8o+vvFKgZ4gwuqUC0yFFiqmm7S8tJ3uR118dxmpHjriAtNF0W
Ryuhj5Bcmte1lr9gbIFxh8zOP+PAWlA7GLcAebjqiHh9RrRU+ymgppJ7dvwp
JofvJGY1rFjUgwqAgAsrgxRh3WZGnQTuWVqURSYvpnqstBTSUcAvCa3zZ2fo
8sLv09r/U80shjDdb/bZvUQ1oGBIEB9dj8DujgSYNgIQLnaqWaTnsslxl9Da
u3xoe2y6QPSW3RqFHbRTYXvNPrYJePpM6WZe/GeaAiz7gUukX+FxGvoEM7RO
f5JF2DUoK5+3cy5DAm/MNXCf9jbSJuMIJdCWOwjuK1oiqalU9/GoKqVc7uen
AmFptgF95oo2A3bxXwotID6E91c1L8xgIOIyKXdUPMXI3nv7N5k6LJcockUI
wD6zhrr/MZUGPpHcMIi/HivsehO4z5xcscva2FdGll7AFjbYxdhArhXGjSwU
r6MQfE7J64RddMxMF2ohHM9RjCeNrcGW/+sfMwMz4pzrX6sC74rHAI5bdHCi
3axGyXlHwKauc0dYgOnSFKnla/p9OZgzD2o6OsOGkeO8W9iY8TW4ytGdBJC7
YBumoAq6yDIr/eyabZXRsYccW1UgIdgrvgWhPBsFu8t+dMz9zpRFneMLP0nN
7ag4l+saLi48RjV7QpD7U240svttwL0nWHKA/nLsmFrEi41Nnwq7iNCmdnzO
ir3vMGNDhULZe/t49jyY0zmjMWIGiGe+SUW9rseslxffkZj580V5ILcIdR3q
K6GzN4evsxEi7aSiBtIkbY9KWmpGd0Z+wE50pD3fQoS4czLoOw6bskDOvW0a
7y/1CdLjiAnKzdo9m3SWYSnzNjmvCVULcrV5OBRV1WwDrG4KbP6/IokfVHkq
0rdcuHw6B2qZzYxASj9h1KEVIYxI4KIY+PhcnDtmh73i8nBmPiJ6ili5Qett
NST/Lte0MIcBI/7afR3kWnGV3YFhYVoxGWvfU5LPA7GKv/d+LzaG5vMyUrNR
9Y8mbzyYzHDSzELp1OPn3aze/8pfUans5i3gifIQO4REM3sfwx9rkmK5Ag91
rgVTu52lynkjVYOzpxRUnRr0bhwtw6quGsvOzihoM8IyYjlXdgIpGO0eyfhX
NxV1flF9jKZvA8PdoaUptk0yvHHpt6FaT1E9uHqO62jL8ZMFryeG/GAu2WHI
7/VKVBpzOShngFJ+hsyyHYt4EO1PaorOrlixE8UmW6vLkwHrIpYdjVJ03li7
Den3bhl1uQpS6Syw2WhNR9yoEXrr2734K6EbfVmiVhGFpDvL5YvYuHVNt7T0
Cn10d93+Fs3dyRG5OLnIIsb0IJg0MDF8Q9V2zZdP9gjJBdpKP7oRyXEbEu+2
kHM4/+9ZF3P8Sm7XIuq53vKvLJAVeYSNemPQ+MfzhVhprjqAg1QAdj8QMrvp
UAHsRT2TO7LW8xvSHFDnrvxruMXmZqjxAZ+zLWEfJRH53d2UJs5SlhYh/hsQ
wJ3obl5FDWv95ioRccyJzpwyIhjTFj4H+h7DqYTbbWIIwT8CLD8u/UxO5YGz
JT0ncmGASD+iyv07EZfg2Y2VALR4tIlU2M1kXtrV6OasF1TPtxYwB4LLMQM5
lm8CfmUXK7Knpy3BBngbqPAZN7WTCGHKZvwHFuwzVwSLmHqkwUTMHdmx7+1O
fdNzp5SVuq5nQAiGBtkloZKI+aycXlJADzxhyfMslq2VmHMIdXJPORCgHCjf
z6EYb/K1MzE5w3R5xDwKCWNi7QI0Qa99Na8n1M/Chsqnw12Gz51+76N0RzQ1
ciFukAKnTaXHjHaQjp40dJEuABT6GynrZJcCciJ6wEnu/StuZLbzx0tkjpfR
VYx2lxnhmcu2GUEzcwbMX00Hu9fVe7ehyRp+ryLwT6GI3cKaDFcYkZdOYE5r
3weXACMT6sQwcM+85SVIgAo073MfwtKW8/3/wSScSLKbEJVBiR09fSEw+TDg
mnUj9/mgf1FkuX1j62bppp6mlvHGxnAzdlhHyc70gME4EJMAvR3Ek6y7Sc8m
0oVQkWkWm74P3fXk311rnBckIsDcgdV1/Cf5dHnxBWotkxjlIjcVhDl/QbT4
OR102J60r3/SFWm6CM/Dty3PAmBZ1hRIuxTthnHI+9HujoBNJheUJY/a33gt
r18xaWTChQhvBcjFzFwuMFwTf1ngCNkWyz0UGpNW18pHfMxziONbLOfF1z3k
5WyZyFNpEx9nKsvSD2amUlPlmoBk/RcaUQS9lvUZLqxHaQNIHmaCj07tBbs9
kGBqA3yJ9ssBrwF2Mzy1YseU7yu/dl36Qotkyij7PQeMGpfIobedCp34yvUk
KVErD4V9PF5j5DoXvJLEZu3Jhk4bdZGbVVFbPCyTLlTcEjHhiNXkxKvcOdeH
JlCqwOIsv6nzUhtoGcwgO4QDz8zZcbJvDCK7BLqxd3vx7qBLN9bWRBY1JAEw
oqaDJsNsxjX1VEDL37KbJoO7UJvzOU6CNo313LFB9BFQsS2q55rKeRnG0WGt
NeIlhK0C4HAcTZjK5gE3yOh/wwd3BzzWJA30wB19FrLl0hDliHpyrLXcEQ27
zyy92ewzsA2ST1CfVc7kC0Z9Tg6X8HvIQh9/1igj1BRhLlC1rLX5Taqejj4w
FTTywpXYdAd8Ef1tTmrMMgJUaDUa7IxgArXAJ2+gwqRRVMY6pPp1C7dnVKVm
7Tw96rs2pj/cbrMfXLdMskapl3av4as2DN1NOavOMVtgTPb0P/ancxhGygEY
efr68ZPPu6qLK94HdEx9js+O0LhAaAj9QGmXqo31sCn/pSqrSm1KgE8c03Xm
VV0oEsmB8mPaa1dex8nHlgBK1KsIXvGAG3cQWBPGH+DYKOP7rQyl4JT2Ld6M
Pyx+HxGSTGUC8toPUZRa3JWqB3Mu8cCWlHa4k4HJMdONc2vkSANFRZitZ4b3
SjCzuTnwxieCObPtiAHEBnhdRcHhU9KfZRNzKCzA4jY84SzVRpBcEU+9wULU
TNiBOosNyLjPNyXvsY9z/hT1IiGkhVhljfewM1auvmw7BAwaBob+HBajrP4l
e/6Zv3nanHahRihNMXTolxjPEs6i/N+9ZsKmpSsXDAqirB7yn6rkGn/Gd5aP
5axQHP+Kqfl9C1fxsHvl12tRNvxwp2RoO430TKa1z4a8jcAV/Yq0GIS50WHs
RaLhANmQdjsEvTLw5Hpgr1ceOYgM1dail6YMsQK/pHm2Csuf59HosaendsyJ
NjvAENGFQxEqBQ8u1Tp3zx+8yogdCEHBP/pY6zVnCEM40Rw+n4VK86D4WugK
d2Rv16TBSUJremjbKJPNvlOODr9WFPRvajvwx64FiSjTzOG9mOKw4R8uTPZi
P9lgywVSHBlVd8h9Pu4P3GDTAwhC/np0jfWXdYHlLVnk6Su22pbxTg/irXKN
oSLqVE3ADHJCJHJ0j69bSKSO7kN9qfoeuqPgqBvgRUGr6y4e+XxTu0tmOLkJ
4TvDKo7m5nCux0+2UE4e9sUKGaR26j5dQxYwxvsJYm1QyIMwVJRz+PtfIt7M
JM33ayLcxAZCxm9JhVTP6kVfHw4YdpEILvypFNM1mIeNOf5YQ29PsUWadMtN
qwQqXh1fYliAHdlCO6SeRv4BDRm8qOMGFY0o0yo3TyFkI5WdPOhNVgI52S5z
x/ZPsLfveXaG25pN5UHBuxF2C3Yi8SVU/lWhaYCR3HQ98SZSCYEct6gig9BA
Fvi4ujnoVAWsm5TfDoTirwf3R1F04AHRyqO/tzfvbISPc5HGBr9Ro+T0p7Iv
L9UQH0uxsTcjm6QR8X9CEJ+NCOIBQVn2wvrXBUIW2tvDb0WKGhZoiF36xlOV
BQx/ieEUO8w5v/o0RpUWZYZmgc7xxDW/UyWxnb7VAUcglrzPwqHtjKCwM7jX
F3lqedbVi/W+C0DG+vWiZyl9ddu7SJQaQO9DG5tkL2X8HQ0nrbqVv4t0pMg4
OKOIT8U3Id7RXdhpjsla1nDOYQdCiFJ7FFw/JDB+s0/iFALpPiwMnEFsBBdW
fPsqoly+WZaPWG5MzNj10SuYQQLJyi+J2bvO0k0fn4eObaGHYaYiSUaYTyPH
6fl5ni0sunQpPXAgndpboeQSTqy021cBnAFnZo4Q6cPFUkWLPZLeu0agJNLy
lmXpptA5J46IHpx+bcbsXThH2Krp4Bom21RQuS9QnWl369vZWq1aEJ0GJEbd
lln0CyfZcjLsULUKAWRGMHnXSIEG+24CahYv7hZ9+/BsVQnFnl2PI8mnDXIX
gU5giiLfGGzTgv07J9U5LRbPJHoo2tfKQi3rr9J3XZ0KLyRA55AE+iOAkUad
njfIVMvk3BPTDYipym5nyZkZu0ZzDE1S0zLj871DiUMLcdpsjFm+Imlu0EEj
bJdQlwinWMFPXGJHPYSKq7h0toBsQwRnb2gsoAcQsrhD4VAbciafbb6XNqdb
qFHY7HXqW+jI5NnN8ScpHiuC+vgPGG4gOOBOevIyzw52qgKQ0PC8cosIT8Km
yo6UOW5sdRrtFhYCwVaDZLIBYF6H4ztIPaHuTy55DNmFbxP3vDNhYzw7MV6N
PCuWs/G5MgqBsC++HuzP87sIeBg4lijxO06v50nF5FAPrYGxY8U3e7nhZHuT
lHiiHlHFaPbuuj6thj4viOfFHtR3eUHMnTdFpneXSuSirT3JdQWIAKYY8d//
Ch6PmiFOY1p00NtVAiboIxEr0bwBNzKgGCB5tcuihW1uvSPiFvwmD+2s8nQ3
oy03BHHZy7WFxPkTfZ51h9iPoa6lew7OURjcXhvFWF+ESGPXSD/H7sY5XS92
k07f8xbEmN/zZluXj3ooyAg2vAhsVQCLtBkQiamFvfgMprFXInYjLBU7/IKW
swwQtrKXzUvnRjhKpaEzBVVpw9qm/5kC4uQvQHxvz5Zzf5nrPGjG6nirTswQ
kYZAUtAPK7pFrT4el/TP+XrdBN0vY3sKSh4fH3r8koXeG4Un9RuJph4zAThu
cK75IEu5Lea5Aj6RAYpZ0F1KSaGpsHmXhBmsLWtdJ3jExyI5biK2QFb7EgX1
nX1EbFKnfmwb1UUSgql/N3cGiGYxldtiDuV3ff0PoU3TxTmyFUOnsdw+e0/f
Oy44h2wmSkWirzVwSGnBzafrJJdsDUMTZuZ18nD5EdabNrhgpthl2FRDOo6M
TH0W8Kloo05InT98RaIOJAp+3inx6LdNaLx2SOYYp2r8kKrRUpDwL4L/O+pt
q/RaTgCdmqh015Si61psPllDCfAib0WgL3WuFUluQI0/l6FEeKFlb2yFUGgN
Jo/mmhO1ANTzFYvTCDTpDJhw4qxA4yeF2zXHo/NHUo/SghlOBbt6YYcwMiMy
IUUeQrKeAGCr7MGjTKNIccBJkq4KtfFlgnOTQIUcv9RxtAEOx0INgT4YfNMU
iYws4H03JH396Ybng+rFpG6dy02oYPvBitPLpD+Ft1vr1M9sdjWrjWX5udGP
ieIlhbsuse43O4ytO8gycNm7/7eSz88nBrD1WP+rghZG3MnU9LAk1gSFYLer
jwx9+TqaPUOPMvpuEym+5sxV5B+sYvIBNCgnSnAc09QJxLYUTvlk1eliNXoR
VZZRIm5zsaKK+VFG2J993YNu8O0yCZE89JWDYrLmHCw/ZwdhmXXfQmgpj507
y36S3/wkMxBLJietUNj7kpnHMm/kKhim25KJLnqyQTOh9mwJ0re5G/Vw6gpi
lwLVmhNrxVZ/iA2i2eHOxifSzjIqWviHnVhJfFOAjpUffKhvlH9LwFc4tIAx
C/f0y2jggwu95ZuuxkcbJUrWi1F8kmUjlj+xoS07f3BXwb022m5uKFzKhpDJ
JzfigR85WwSMc7rU9o80aZXhbnXO2nxr2n1uwu+8VkSd0Apljy9p7+KlzeDS
Av9MT+g5x5BgdpsqIhkhCk6viY6gFJWj8wn8u2Gb6dQsLnxUtuvoMJWUaXA2
G82jY77ZlTwj00CehHYb1OANkn939BgMMhfk3IrH++kj3iMqkW+THs4UJmtd
axoPzeo890Pr2Me2zz8eJcxPEVOmCk0eX5kU3b5G4i16iUINr79uAUsXYGQk
37vhmAFj79aAC15KZVXHKC3EGcD3ybIsOnI2Kn7GqUbUD/YaJiVNfN7S7Wur
CYZ/a7lrHTab3vBgI1tQVX+HmKKqSqLZ654TvvwV05H4cfIhaf83ARqNK03x
IVWx06S3lbRp20y4L7xutoN0FgwETn0tsB8Qr9m2vGafom3qrY+wO9wFg/7c
DtjHJgz/W13HMcwWH+vgf6TIeAIaKB9r0NUKVzfiQ4EWVIMfioWqhba57lKw
4l9pb1H6VjmaAD8S7oopLrvsiUqlS7DVUvPu0EpGrhba5rafO4jEnD/vEWXp
yfev8YCPymlTfXFSHd0pNpwlM6JTm+7Sju5uAClEVMKEORDM0bLvkg7iMOM1
XE/2vfFODWevjYYY6k+JpruZQgj93tgJAge7JvOLVDfH8fmyvog9mrHWaJyv
1pnp1Lojzr1XLcbiJe0ua2tlhBAy2G6hdfFmRRt9RtegqAKRV0SZf8gTma1I
smcRXRqL7cquTltvYtEz+8shl2eQ+LElLYaZ1UJosad15r2zLQh3ks+OEDBS
phZhv/xlLYSbINbHdITMp4srVsTHD9WHwzAL1pNfRjLKCEeg4wNrzIL8Skti
usCz1nXVYvC5wsb54s8xmmbrHztPqrdK7N3IhWlAyXnDS3QzInlPh6Uj7MDk
IkYi2zdvBJSCB6E5E8TJEQ1ZZz5vV1baG6ewgXE2M9W4NP+4z7lG4RL4hY3O
LeTp5u7z/AsCfWwQ8OtNsmBtmilxr/wrmapNgpybP3BC+g42FktCJa3upfs9
6LUxIu4mFtjtjJTLA3zhNJIlKZUtRJ62P/47U8Ht9xCtE1caLBTKLBzFmUI2
1lUfCL/YrE/NBgR4fqdgykFoIViPsBiqAP+fyy37oWGoiAjkehkbmQtb/j8v
uHPZ8bphEqIHag+2lb5ERu1ooA4drWQMUyXSjdEHpKxaQmdqzPC5qw5gcPFC
+wodrFlctuJpnXss08IdGqFEn/TfXZj5pt83TsNlgNp5qPd1InW5mx7ZcMb7
NOatVjeWppMObcoYFRnJY5gqOmW50VjKeTkgRLk0D+qjg8+GBEXE3GNAmCDR
q1+kK16XdANVgBNB0c0y9fhSZnAX4honJnlL47Pcs2U7JjuiTyNGdHAI34VI
g1pUMC3S27kltTA4KXoJ7kLrg0qx83JRR9M89SUoPHSMreolEdldnx08ExOp
ovRp/XOqVqTkrCey4+RmMofoWu0WPBEb7/QJIdA3RRN+Ph7U2Qjpmt+0QY1Y
Gq8gAkpiLZqAQxPSZNieWaSWHcSPx6f7sXEiDHjt/Y2YuwnYcQzQnCWsxrVu
PrBdfrgbiF/8oind2BsD9l7ctACop96EBS/mLoK12aYGhOt7NMGoa4EThpx3
/PNzLBl40/JR50YsydHxiw8Ng9tbPbCdBsaZHE7e8qm9q8TQJIMVqkUm/i5I
rhbQUPKaLoq1h+AFh2dRr9d0ewp+H5Ey4YY4Gy069Wawoy6eyfJwup0k4qkZ
z5wqqxsGFDhp/nsZ2HH+K+wKzbKb/6uUwbDivjW0Gk1B9GHzZLcGo4++K0h0
EjvJC8SITRp06CnFEuKWoaKchYBYLjdNimHi4RnQPWvcDpUeWVpQ8K2KJd2I
01ziNzCMLN/pbXEPOzc3hc0FK7Gp2TKKcyuKgl+1MBdht9dH97/wcfreCz9H
niT+MVE0Am76bUfqfy9NmSy7me+VcYKDJujPXGTq+Uf4reAIECcpWnzvC0/c
cNKmWCkyG9ics+iLinLS89ejyCmO0pao5n0Ol4ULAVOQ5HboQbd/1bFud0uk
QEGrbElnqIbCT1FeQuOu9fmOJJLOBwLZbuWLMZ6L/HwVyLDVABtPUHxkOwWg
1UJCYGEeLEvmmQdB9S2rWfTGUwcSEDAE4nsmWXk0dud5HPkRm4cL9fteLe+0
trP4uMbhYxHJwUmPUiFFYYZdIWnX2PLI+6IStllhQI4xUMGq6t14pgiDCh+i
dl7Nqgn5Yjw5yq8JouInRKyCxh85z70dkqa4LTIQCbpWIdNX5EYy/MlIoQlK
7fsPTaakJqk+1/bAC+TrELcxCPbIpAyQcZcmdqs6oohrVjcVrOK0GrVIng7A
ChH+ijMeNSVM8jIgY5T5w3pDajY/if4Zvqc+xs1ciJPiKrWZzyaj1mwkpz5d
oUCNwaxF9kiketv54I5IK58OsGNAPfQT8j/0BWo51eSd9GUO3RLfTySyZ+ZT
F5ZzGB/YsIAEkPzjOwRebGLYC1w/GKu+dUTdM3F5pcPVglbkaT+eQv34FN2m
Sgg61x9upYWbK9CTgFsMnshgWCVoKHvaI/8N4vBK9a6MSuxFvCPdzMY37mdq
OyGwxwYEl0RQumrExgfSEXyXbtTlKBbmwCsjJI5MhkqHuX/THbcKB9Ef1885
ZraMIhe2h7dzGlmB8nhEixZTxnr4yBk2h9nyeHdwidgBdoC8yz7X9ILKe3kI
fG+o2TA6fxpWdES9n/HRsdXPLSA/FIEJO4/WJVYnL3S4eYxgqElloB2O/m6L
mvbhRTDviB8PQJrR5OWWSPnLL4okprbHFkJanejyb5uc1hdjG21M2puCq/ka
dDPdKyYFPR69h++AIpkeQ+h8UfOrj4hcwNzHfJZ/HjvbEW2SErZA30c7lSrw
xZdPPXlFtM3P7vheTktBLxj6TQsb4AHW/ry8vljprhpW2mXaIKhC2NaPQyFt
wfREzfgcFnsohMJXYt/ND11Kldw7DB+UwnnwAnjf5NUKJe/ywptUn3kYd8tA
hHHxRCmeZX14enjleyRYAyMgC2XO96iyIgKO2vKzkzEfMU5n5sLkd4caCUqp
iSm8x1G5mNYbVGB25EgEkzvHKwCLwB2oYBLwbmtJdc5hjCSTU27L0YqQwiaL
VSx8X0A22vqMt0kyq3kIFd0ROa6Gq1B69LyvhbpvUqXJSV7sQp+1E+5CMZ7X
sYYI/lwy5XmwD+m0qZCZh+jgAs6PEIQnioyw+7hpca5lIjiXnn5xbdEJRj8O
3ywMKW+se/NlrchTvFEoFF2FMfVHmKxf/VfyANbnIapcvn28nVIeBV6aHF+h
UKH7uuAHHnDrzTuXG+3Cu6esxOi+5ckm5cKFHvUICiB0vSHiwFWIcUOVdZ07
iMVlQc0+y+za8uihhZGofzgN7CymEpdjH0GxsT6sQBbBGicMxLALvHTXuWhA
ZtqSlOh9+NxyeORa2kxL3gY9DpbafEh1dDmMz/s5nOB8tRpccIBJBUPWezMi
sWKasjXqkxgiaZwjiLifwRohqUoJRSiVMEyITrhLlGa9QpI5DfKXEQGafj8O
xiCIvoRAnrFKWPCYeMthtuebyS+cS+5JXIYpuXLAY6bzilsC8WaZhKx2Tqta
3jcz/io+niixh381fsl9BIqFeiIV/2rChQEPyRYZx/Ip57CLtXiPDucnL4ez
9jGi/S+m+vQ7tGPkEyixi542ub3/47f1X6fVxUeETGJxzNZWgyPN0eIJDcIa
m16FhiEmH4gSR/ePBlBE6l1gl5Wf5skgpYEQ8ISZgFGE1BbM0Z7bFejRzwol
WAU4E57Q6SIXpyOreaKdlO4NzPdBhDsVrbArjkPEGLd3MV5nexJIvihqATCB
t0fUVd1cDWMEtLACthPYjVfjoPsIw+uu8vbrCGyK0eMiZZnBQOuvUAUZs/17
NND6yn4C+bEYyt3izQGOMgRU1c6exwEkNsTiOzXBHI9OsSI3RaPtPSPvmCUv
I1xa5ZYJNd1r5KW9QQRaq3vJnwSiu1/sdpULEBoFw/K/HEJxCaYK1JSw5KWz
JO7WDILQWrN9li2B3UKItE7WuwReiAOF+ygi6FZstPsdWWETTaLyJzvtonbZ
MjaB0vy1XR6FcAAR6c9l8xB2olwCIECboLPLJpqGMhaFotlk7Y/UtSqwvR08
4cHUf/PsSgULwWQRC5k1xJpQ92EwR1c7z9Mp34FWZy0+v/pct7gd/0yulDqO
XevGiK9mWP9eEODQWfoilHTVf2pj4QCDglprN64oCDtFgpC6JpKw4GDtDVSR
mYIxYt8t6/Gs5XMTS2r+71Q+2dvA9jh9AaIGgkdZWpbJ1U5uBgssmNJbH3aS
4zD5bgeXHuWULRKOMu/p88FM2iQWrfe9S/vDDoQuS/mYmDA3hTvv+rYPVBfe
LC1+aoflC9/7PtWpj/aR5AH8fQZ4ArLl92x1+bIQ53lpVR4/AzyBfQiDOzgx
Sq9Xdux1+8MCka344I6YA9NtMtr0j8L8OfDHlJ19BA8XpckJk4BlUlGntnto
MAVzGZIhkZyidknY3v0e2o4klu+yw9IA03zmlE/kfgOL84Kflp5lgfGfNVNw
oLxqe2h4bKH7QDvo06IWQAmwYWez1rXNozCPJqB4Rkp5Uh3+h69Y4Qq7ryyY
rdfSKEJcQyzWmNuDs1uoGZbRuxrzX9SG7sYSDC2r+6z2lDJu+jvE0quSbMbm
HaPr1ZpsyJiQDU92GWnXlr8kQHdttFZEL1VT1UJpZe1g4Af+7YJt/h+JvW9N
cEHqyBPeilUmdgUvrXQe+KrRu4xQVWiRUgdyEH3B8sBGPyhrZ1QQJMZ1PpWn
bpsuiVokJlQcJGBUWhaRjQSdnI6eSF9T/9r/dNgXiQ84O63tecOpBTytfeuV
oup26WZINvWQ/YlEaZ8lwiX7k+ge4aAXZTTrqY5aKy/9f+V3uQTvHdiv5og9
9EbyIwfgRTFCElwfhn1I8L0drAgUj42jnr1SaOCyjENzqzDr0E/gzMze70c1
K0mEYGMY0RO61DYT2M/u+zvXUfhMuX2SVbm+G90VcjzGDGXkqwH4MFwz4A/Z
PxG7UEwMjk33pNQm8cBdaxND6xg3dhYwfisMV7Rfk+oDtoCj7/Eb7eXh3Zlh
JL1f38y0H/IyzzJTWzTOv33GXEi2gTteAbCK6nVjTAmGB4PhrujXFALsg4Qv
4eHGBFyOnaQpTyTPBviRwMWTEByCJVCOY0ZGz5882c84CrCyGupgcnTRKiHV
dguuA1DyqcB0A5x386fPYncX8RBMBzmMAMUPFBC2bsoqbPuWnp+R34TmLFH6
A0qNhWSU9u6pdcgXjFrsf9Vs2PK5zq+ZjNKmhxY7wUzAit90UA5B+Xwj+Kod
ldgUVCd4kJTUEJjAmScanZ+AazgIMP9As99yfdlipA15Jjd7cYA8fPd4bccY
i5Xrlsf7464fi0/LR0JqSqJWZq5IeomaO1N7d7Lr7fpuSPTzVvlH8X6Pl5rc
QUXyVxbFxbG7p9ccRAmgBCD5BcHyG7mSfOWFMXhL9SLI+ylTSoaU18xD05n7
+sN+QbPWLGKfZndwvB7VnjsNPlyJV+iTou8CFuLCMUar981su3G2MOxeum5/
79egh07bPSPT/UwBIKx/jneCvGaz/P7tXo/pMItZLqNTE+tPn49Mv4DSu/sX
58YjGNw6/TtQGTAsflMtOc4dYqc1NIO6fKaF53shCS9RWvcpB76o0oKZO7Dn
n6pPrHnanqFk3dHljG7YFpozRLX9kfJBbQIsjSZ9E3EH1G9Ih3xRfyNho8Gs
4KvV/w3t8Vf3aFZla4ZET+4h86Lr5sso6FYdqGVzwab2PkOrNPrPV8ZGS+Gx
mXLjDaER3q9t1ldt0rPUgnrLWWdKhvVzbKTanAp/jPkS4gi0Yftf32L3YHRd
af7m7+9COTVNnVFr4Kb3c7k0+xgtAGdNKra7XiBamjUAtlc1mg0CkFQ5XftI
MJNut12Lb4bEa1poe5vj8WazSjcxeDY2o/eYgFnLygqca7f1JjF6mi00yKTE
iuT2WHjwGyhRlvlg0BOumzFyfGYcDd1FvHJaSlb7XYH66MJQ6cZwN0vcd9jT
w350i1saX3EcNfRLoUTBDAyzwil+46ugNPB0eJLmvZE7SyW9G4cyGCfzt/8W
mhmu7Wxns7m1PkcikbBwQVmubavLMcoaDWzBjCP2OJQzkKaDLdvS3Nm9lPFr
yWfB1J4VDiz/gw0DrCnlhyMtvNLUqRrYnQHqLH8NPMVNCeqwWNMzyK68+ZKQ
6Y9Rnw5jHlWUOnw/r/vQrgx+HvZut/wNgNMHLF5Uj6F7XD1CJQ7RrMCjtZ1V
uz3/W82r4SRsw7IzRpZpjFguEe8TNjoRTFoXQLX+IWYe73V+XbJfz3kCmjUm
+K9M1Hr+REMhpU2TSDHWql8g1tb/cJtAoD5Wbusm+mVHDuHlf61tEy7SXbq3
ehV47PfMvfuJrB/Htr7CW8VwvJKqa+b4job1mpbGR41LPlb4Up1FekF1vXjC
OIrAZFI+axdjis+8zpKr8eLEnIDazumip7mMqIvPQj/HmvI7/9X5oFyVOvoS
L29DLOcfXQBXHsaP7kppkuPUYdz240o9O9PeVTNAG2HNrNxcWxY/jyXuNzyT
wl8ArShQiIIZoxWc1K8p224hlr3kGrvOjOOs/iHLQf0s1CUdZg/UvCJUPf/S
3sG1nDlrJAGhXAGcd+UuiCDpd0x+0nBdYvfMNXpObqgpOIDF9aC+f8Mz/Wmv
zo1ygGaaJjSzDEQOUuawko/4wJ2HyE/FoQ/hfpZ+l5p1xkLwbPBAZFO1szzq
xbQRJKfBAFVAXQ1KX0g4dcTTcpGTQJZQWec0iO1Q/If4IjGXjOEKVt4bmNcx
VDNPVYB+nx/G6ZYgoR3t5I+m78zWZYjYt9I7ffEn17+bNb5/M+5TR0RE/OMN
xpQwHfeELaGeuMaDzKXEwcRCWibsOm0JryyRWPRDVTnALvpWRwwunG0KE4Bh
H4Kk1ZU5VlWO4Lkrks9po82LENfW9DRj65bZgqlYnWz1FhdT0gNOZSBm1odK
HYj6quBkTsTN2Ir+g6U6KsTR02/3RyzUnqhCd45U2DouYd80ydbgO4yei7P/
ZU8csaBLV6xhMJIZ9Xu4x+1thAU/FULIecjpAelp1RONc8AOPdsurLbfT3wm
4Jzss6qqE6c6btQzGzGKtcJunde+/zfGiCcyyxLSgiUazjikHU3pVppPDwKI
hI+gCi76j4aCxE7KDXwRdWuHxYLGxbQwM3sPQYO6E0e2NVzxhLOvvPoyKM7A
BTHZ/z5CpUj4IyZ1RMkOVdB4hP1a4FdO6TJaoQyqRhBFcf2rf1/p6S3sKMi/
1TlpOpOreyig9620nfk4PkMPz99Dfon0Cj6+SRw0ZmxQrwFO9y2PeXp1FOsY
tn+1h/uY7tuac0uK5mfJ5xcgB4axBPjgo5SzUOhIGmQXvxuA4ZxHm24lIrXH
GaKrpWNQP+nJFdqipm6GRJPjsPLYV4hRPqzoCj3ZMDCaXWs4sOUUH8S3zMql
cCzEjAPeJcwdgPWJjD70GO0+rjTWBHo55nOJJYKW0lzpnWVEEA63WJK0hrQo
7pgp1lzhmLmxsl/cT8Y3k0JY+f/IXFHE/qrCPPtcLXknNpXSc3QVXOZpqew2
DaNYG0q/qg+mEUhT4E+WyKzCi/eC11gtlkI8BPAuxNBZBxN1KB9WD4g8wxJS
l17x0MbkKm0woChubdW4iHURJ7vQC/Sf9/j8fUyA4pqH5wmSsxBBNiuym9V/
Q9Be6JTOqLql4RIsXp8MoiR9tl7is7u7+04x7MFvn1IN2A7mHOyDfU7S2mq5
Hnte20CXQdgLuXLhkZGNctrhSKTUpp1vq3iJ7YIn3yK1eu72Sqa9PKcMI/eC
IGL7jzgZhfxClTN2PS8MlETL2yxeDFBWdtrTW5hHNpESQVFdXxCP3OoE7XNV
3LOKEzd5c7kVUWKo66g3jxpI+2DM3uFKHJKUYjzI8YNM9YGkPavC601FGP5y
YcnUAhud3TPVVRArPz40OMwDyL5zhapzLjRzeoJB6yD+e6mg9347jGQ1PDZ3
ZiJnEKj0rUq7mf50usxWBk3GTaJc+RGCx8SgdgeyjwdRP7+HILeAzHeQ2uD/
fEhJfh9vTr6UF+k8DmpVoLCFOdoDCa9B7Ww7GRvsy0WWk4bk5Q95UxieqpaW
/olL1hYsc5P9geehWZg/PREDp/ksJ7lEVLNFJ7X1DTyc359ELxiMIbQ4y+RM
+GOTHlaNR8LylW3WK4yKpoNklEUF7K7MUpHeO7laJJCChkN+b1v/0rqAYvOZ
0BtvMWkFYw+ThJtY5KrEh9RTHII9KgMgEx+qxk2Z0GCfcfNnookTVEQj3Gh5
eexAMy+GpbCveG8lpkvt2MqTX4nfj90JdDj5HM38uoEezFbSJslY63AJerzz
aunVkqTSvzRc231y32mQdzIoLdIu4+iCOCFI+judJQfQQgkdYGLCPtPt4dyV
0feHZi46jU4xE7Pd969yJuHpfmdlzubW/4u1OFHE1/BZAuVfkVVgXfFlQ8dx
tOnfhpXZdXYxlURPtEtBRLdG1DaTJmPZRQ0ANyVUJjp/th+T/s+Fh0+/tJU2
aw2g/y02vM7avy4ztTlRXxlcSJ3X28VRLnDGxn2F0lAuBArzhLcbJhmmbFjW
hrgtpcxWSlezm26OTkQJERs7SJJ9cZefI05rUxfnRIqRHwOWNWRlhGYXAA6J
UYhtRu4iMZcOMKptE2xtijSAEkk/K03KHlSwI6JSBRt0qHFsJRxTdcZxfTPn
Z8v5PuPLpi4qAwelCb8H3cFty0twuC9CaujZzP/XESURsGdCkZKXh2Xl/VBE
gSOJz3q+U88Tlk126rlTPxVEvl7cuWo1yE5dD1FM9iI0yQReHomAqcqtI4WU
+TNndRQK9EiF3GB7fbdv6u23Nnex+zbcHVKVlsnhHM72MmVaQkuhGH0pwVgF
LlxmCINQqoE8usc4G2V6cFisHFokjx4kbwvdrM2jXIQYrKEI1juzVjQFt4z+
wqL8adgjhlccMSgKWPjn5cBFxPhVY+48fufLRY0cptuZ50AMAal+1WJkJtHF
I6UoU14QAqaT04J2Tlab9OFeF50rKRTjTBvDmMBKyMIek9V0q40IZKLivnEF
X2dFWLX1cUUG/RGkdLFxYMmL7KfOLhtCDex3ZAUfLSH7OJn4737uhok2n9oO
FJwG8/2orXE1LoD6yAp6g6rHTwX6lWrLxjMUPHbUYLGU1QKZtejvZOItuCY7
Qi0tYyTgUgVPS2Jz7CbO4mEObs5G4cy+B1NxOuwHpmQkNb056brBSggJj2Eq
vTctAIzN6G2cNFxaobb3/w84jqvf1Sb8wfGG6izK2a7tMrYQT/TKIll1M8R7
vQLflci+LC03L74PAFsK6R4PURkl01toEN6UpcTMRSiFqxMqyiYQjoxNrZvu
95iZrpY4cMtdNKmSfZZLsJiLhmPPj3Bg8SXggtj/bte38mmCeLfwt/w3swLG
vGefRHdQxfvevtLd0TPNMFgJYPw8xJ8zMWDDoBgcR3IsHcDDimen46/uUATQ
ayKzpSUgMBK+gPgyc1fYqmmDN4y61N7Hdv8PxeIvP8Krwdd6x9tcaO4+4teq
phLptPHe7WixSrqQjzt/ZL9TR9B/Lcog45Ud6x3Mv/5WprnLZ111Ft5YR9M7
n4QePhS/413VDrPRA9POoIWnfBl78OuFtudxY1IL196fOAIEFIJTUgO9uo0P
RiS3KvYPmBTBacK6JWNUUm5ivcSmadi4zuOefPD0Fdit1eSd7rrZqo5oi1le
Pk//sUjUHwDsNVQ6Z5PYp1Y3e+ODS/kop7NF8C+sK++F25eo+7zOf2+wtHfY
l1I5dNLqyYMYxH3vR1AZPlAafEpIFjnXzfZF5xW0EtjAiUKm85O6U8fsan+/
JN7s4zdg11l+s4vQD4w/gz+iq0i2m9jO+iWpjTuRiLtj/bEgMPtV1v5ijOLt
6kNSBCj2IBaIr0rV3c7Did3utPmt2kxhvBsy/KgSShCmjWqrzihPT9MmPTkU
g2XNCdn15IT6jN5PP8wKJzJi+7F/UWSy5pJSO5M6rIZsUxBtNqVevpp8zGej
wxdL8E7apl4418T4MQ9X+fLKT58/KcrUPSouceHf+BE/Yt1dKU1nnH3WmEr6
aceLVqYjDso85S8Dc6Fv2cJy0TtWx0tTjxA7h1Pp6w7dOLFHHpqNPucd/0pw
dJ8afiUjriUvzvVRi5sKr6YNIY51UfNaH22eZTJ3i/k9VnDEIeLaAuZ5s2X8
y9P/m4ba2K6aN5xC/E5HoKYkUeUy9fHiifS1OFeyib2281EtbZLDFSF37+eS
M11NHtLWXXB73kzy97aCImRqLjzUwA83mQgtrpOMLoAWz/NNT2ElVEvi0utN
V96QIZGPj9oAV4cqWklGLWjlM7hmQvoBjQni2KtnVhBxBL5VjgdcUcjiCKx6
ynJn47ND75HBwHZIMnQSFA9LpZ9qxxpixZr12lSX2Umc38g2+DOmZmhmh/3C
bcsLBW0bRfNhDmlIR7SqT1F9vLPQCsvOuJTKg+wt3GwOd+Km3yOF+iIxBJnx
mFSuIG3ndhRCh+lpz1eCdq8hbUDP+IsfxcJWPJP3M3YGUm6nojUNBRjmD5Hy
OtA/kOxdvaJTK1TibbWgByJ3zWCHCIX+eEbrs032cIcRdF2kXqfF70YPQx+Q
M413/gZHXBAMI7qyMOSn3vqlAv9OsS/GFWVi0uiJnPVp+5tazgwyCnJ1ckpA
oLUojwxFmCOmJIIvVDdkU33E+0NqmI2plmXrMQsrkXFPYhwNS5l92S556Ag1
bAINydGjiyAWALvKavO13Py9PxLwMcol3O9EInxHEdZSYTrb0Kmj34TL3S57
y1UH1H2Yokt22U29D1kL0HTdR67KByjFE3F3MMizdXoXuKC2AQ5cjN1PkSPN
CRYi404YGbYdO7t1/GxI8WTsstwkINa4fzl8HH77CzQRiy/Tm+YOdMyhl4tA
tOoXoNGY+IZ0aE7kiMM5HlHuEHNUWaPWjhy/TLUfWOas44waBaqGdrVgcm/n
DaqaOE25AGA8EwhIl3OOvx/EH9D5B80u1fXQ3OeW8M+LUZd2SszFLtULF84x
nHZCn0OWwm/8CwVxtU5L5aVABALs2YpWVJJrHwspcXNnUnUlyIJ6ITtF575I
uJrv7K1CNYjDZOoHqLGCGCcoS8En0dz9ZxLdmX5xG8xHxADU4YohdF6wQrry
WxDY9A6tiUNLzb5EOzL9siBElfFnp7m9Es9LTE5KBbvLFmLfR6257RMWcdM7
W5WSDL9bDAettqYaiakzQzdKjUFtVMg8QF5wKJQBRNE/yRQ7X+o2yCO/La1j
rmGBrmmZTawDkWCL8B9XEIiQQ5Jy+t6HbS4/j9cEJ4RiTrM1S6FW14UdqByO
UYY40+k9qwXMvOEuUY9aaU1SqeBKoULsXaN5/vYKHKGga6df9O4bo2O8LGyn
ARX3tcpoOtgrQkeAxWeBwEfgi5r7EffcMqrY0HILDIPlRUrMHhuPwXHy/e96
OhPoDEH9JR2CyrITbtQfXZc2xZTu6e16cN9RipspNemFs6PqWq2g3F2DXTnh
kfvVT3N+25tTfTnb6xpkbGxuGzKVTj6bw0Pun5FaIcDuA0B04LA9WNRmifqi
q2jwRH6K4/0kTgslBCVOgGnLfDRRQbT8UdDcldGB6E6pE/4F24x/SsmPWveX
lAwu2RRskStXXinWAsNXgc+R9mzrQUCZAENrPh33fx6GuaLefyses3h+1oJc
PUOfwFe+p/p3+7siDkNhkbNAX1RxMIH4GeLUMUygprpVBQ8WJORj91RF7R3J
hwQBdfOxwo9mvz6s0+X05W/GV4/thA3sjDcc77DvQw5MWHnfE419WQjXKPdo
80JkKjSMG5KHE8uUADKR4qjvrsI7YWlyPFISW7dg0RCYUd+ncHknpYr0W/T/
8mjeLi30SzLBuYpifCAT95+VIoFVD08AhTaRmJAwsXSB8H8Kb60qX6e00QAN
DcMqT6y3dWOCOj3xmPR0RtyRYghSSBdJgDqKiwGdvIuEC3fJkoz1/DuTH8da
NB3sCBHGaAVJblnoMbCXemvFdTNCdeKNxvy0SYbF18ZfPjx6Pdllhz1x3CMU
/PIG4qwgB3U0P75lHkCnjrjPaED5r/UM2g68XVh/mFdF2mHlo3XgjV9oFVb3
EoNKkzYF8zXsuYe+JVh1s7eFd8hYAOrXMABwq0S6YVPg1ZevH7JQ76T6Hcx7
13mDLJLhwqrKIdrgpTqX0cHIAjcm005oacL/0HFmVf+gW2wKgI0L3FuBD5BS
Alb/GrTMDZ97G5cxAb4mA4Zj0xK35RR0qdMVBqZFp06Ias4srmpqXBR5t85C
POSHkbIy3PnbeRLLIy+c2ANpGJdu7Tk2MSkfm26HcrxgJxORSxvteu0ps/rB
/OaLAtzGs98dftbV6naZdIB1VwSO/BGvvSlMI465ocuB/lcPEKLdJN5I6qmZ
AyRnUao06UIeVQcljroHf8ClUIzd26VeogxeBfRCKLifatFi/fomL+ZByDj+
/9PvHcZiUm4Ug1qPTKBzIVwzntY7zqbm0VrhuZq3h5CeAl+tSYyXVPT7+TSn
N0/bBzQBj+pq8UgIxGbV8riku0KyD8qD2mjcIIRGUtFOQL2EArIOaxc1mt5R
2YS44nLrB6OYt7gDPEaLBia3euLOhW11kPS4KdurURT5sIfV97ISbQWCXLCu
86TjF9RrFKogCjEItrrV42M+uXIKFg8z+cIS892vL1U1c9/hq9Zb7+m4+nNU
nxILnRqdlOznCXMKQ4iM4GQsH+fmQ5BNrD2tlXhITHYzQUPOJLyNGxuefsN/
0u7LlEPI5YoBMSp21si07XC7IswHf2NsXzh4QQieK97/vTtB55ERAEi5e1xl
8R4+ylrIY41s/KwNDH30JQOSb1dcDCOXtyldS/n2apF8OfjVBonI7zgXUK16
rbwZheL2D13XEgqXFBLjMydD3zl6iye3AfrxdywgZw+UkN3MfdhYLm03xEtJ
lEFO5Xv8QIn2ker2OjwvGfe5OIEZ/gPH66zuq60WUmITm++I/Pmr48gahRt0
U8lr8Afzyu69F40YUXoYSRDOJc1rhTdW7ME6UQBlYJmkrjuT6qmBEAuJ4+wa
09pGK6lhdkBLkdNRBg4Gi9wzj+VUrXckSQrzJ6d2mUWQ/RzrD/SmxBFSIqYb
Y16dK/1wG/Zs7NjMlYGtTsoi5eoxmsm81UgvAleMG6XNhH4wsbyPs7mhV0TO
o63fNdgafXWblb7smOn1qzQZ2KgAmDmqdhFjO0eNAvfqQ2+1Nw6oE+EhghHE
jyiTNE9jLVycoKCB8ghkPWBlHpucXZvVdC6/Caz9vV1qtMwj8d4xn3oUfBpY
FPtCdjTafdzOVuKhLGi2yCwVLhpM6mm5Q0xMHOWRFf7zOsZuEjj7wkgHPjY/
nLMN5IGIAcz3fnd+Rj/HXiKLZswxXo9OtC2uAmLViBPnwAlla8mBAWNW9pRp
4wi0y300vitrrTQQQwcRxc8fZ4sPbs3qlWhho4mb+IOlTbTItgckkW46M5kG
pvYKK0E5Y7QemqwLpl+0EF8PWPXSCU93cmfp8YUUF4Q9bQGYlwFvhfpJBD8i
1VdIujLv4xXvzovBQFQvpLZ7wkh2cEAEJuPVa+2JNiaSGTgUSkznpuJdhBrg
NeIVo+9m1yxY0yo3e04IFAcGfErRPFZu8YZJ7TyQV9gJ9gXsY9cr+RjJkRoD
IeHNeJUVhVWhNeNWFEKTy9BLNVSam7+mKzPNdlcwnWmw0a3iInSMnFtw0sPl
fVpzKrLxMV40Q8aP8YdCK7+WK/xbQkrK6plVaWbzrIsz5LKRTIKfm5kkSrXi
dRhuP1ebEiCKYsk6xjxSdX8dgV8ju1BYe+UJfrfZzxbMIhAAcedH/SGxYDl0
EN4tt9KZIKRk/hz8vtLVpJ63XM18ij4NwNXNX+yMkjtd3bZYRyffuQIklAgc
wEi5WI3uP+x6xNoQPHTGd6yHqEID9WZCiwtmWPvF1Wd8qL+aNWcg3pN8RlK5
02wcvr511rBm6vAototaq5RSYRXrzGT8AO7Jxx3FommxuKhsPXm8j9WrOt0x
NYKFZ5iML5e7mkbDaeqt5JJoRnrIcrGGXylnttg+Ew06OvyJTdjPVnehSs31
OIY1mr8JDjzUPXSiqtp+jOkaduBwdwFi+O5xqcEDf/M9h428PlX4H2UycFzY
dJF22wDszPw7wYtoLYPwxx6KNSyl5n/S17XSsn+HJdQCZn2YxktDewJANuWh
istJBMFbrA8tA1dzESQGreUsVSd8ur/XBGpxOO4oDKZU2lnC7EBomXjBr0VD
QR+ibSR4Q5Sb6fFqduAfcch7dr74fmKtUmFxEJPfN57W+mcpJK/vbpHlWTm9
2QbCYdkQY5KQRo8ao/1ix/Gae5P4qbyUXTxinSNKbDkvOwcm7MvGSa9EZQuR
Q06CC+ZiVmbyqGViP8+OM67JMwXPFHZuFwvrNPBNKN5mFj6OmtBqatBDpqIO
FQlzE6QMOq8+H/nkBCPGiETCWdgWkm5AN0A3e/xjts5tcfdo4/dUlEIU585s
eRqc9Wl4EU06r5/WRk4/pA1mCkw/a+FajOdBNinxrHoEYrwz+0cE2LJNauhZ
jTDdomXoHbPmw0AnwnaJwx1u/G1dmoka0todZkN/L2ocjNtI/BLGXgPDspqe
cFFLKYoAvyHqeKXhZ9pnCrxuYt/9U1je1PHeXIQ3O2tulj+FgYa4nfc6NxfL
9FEO/2UpgzsxJlr4PLgZ2ktg5jifdhEqXtkVK1TzYb4AbbNNV4icMO02aLqT
Lt3GJhuOSgFjDI46WeQ0uAaSDb2ZQnJYTqsdVh/gRYpazYjAqNFtK7cum0+1
9Cu8XEEuMm+Xryl1wOPcpx97H2vDo44bpScut7qwLzdhjfngX3z68v4bQK3J
tTvKrAEgOteuPKdjNfpn+iFKpGX53juezxNrpk2Pber6KjE2cogH+kNGDA6F
QWhCfbYkgONCWHWYFn6+MiqLDQqi8R9uhj8XJIif0eqG/6YxLPO0/3RoZaev
BD/TLeZcFnaQg7QmT1tHb6Kv8bywl4kIsH0lXweFoVOx6hSk494QkdnIilyP
xGSluOb3lzEsmJXrx4zMA9y9smuEydZ4qPI0LiZiNqFstvBjXllsNACj5wYp
WrIXeiWr3ciMGQhd310W6EeYKOQ/q+IqAHqyOBa+P7a/QhHFvEY/dKlWieMc
ABKawQpblNOhnz++ajIJdToLWgK+utu3l6o86ZX+15gvIOLTvbaI2MkBi/qH
GTULU3IhIe7j3YhRHmMbdEn/qlTHQod3gpoi0x8tMee6lBO3ifGeNJgrVOJI
dzbxg+meQauWeMOynVb83Ztyj6HWNd8w0QHH6v7g0V0vZajzrt14Y4xM8CK4
UQ+yjukZ5taCl3gyuDvlsuGX+6qtrCMSBHX6oDDiLpP/3lAkVZyYiXk8BUl8
kuvoJ507Q0xt76xZgQzMmhoFY+EBiJT4gykaIiYQfz3ECiNH6/lseiP//SZd
Kn07js4Fvs7wcb2xCaw6bUSyBJvS0/X1zews641wzkI8cqQjbbS0Jn5ZLZ5K
gU6nz8kU/pPs/psoo2LYs5U6RtHSc7gObzJELAg0pZXxJ41dADK+lU7tlRDN
55Twy2KaB5InniHOyWpuH2rqQHGl3dkyTSVTpYwncqe6gEeP21Jb6ieS3jl5
ya9nrfWDk3oIJDMGHJT+trT1BD1Oyf+l59X8BBKcvf5dzmi33lR2ez7qLUTS
k0SbOUvuPZIg3efm9Yg/h8lhd6ZV2su0BCVkOKcaoqDRBA0DCA2ISPTz5xJ/
JC5cf/qrLR4diW89LLQczZtR0PI6E2dq7u99rlDErU9oEUSN/u357RmprwQa
12lLyK7+o3tJO2TPebu/4Nl1jK2uDJ6Yjda2FrYaH6cpKf59uglPmj9Bza9n
ELApO19xIQvULUC6GUdnvuSRvjcen1J9QBGaf5E5AEB/cp6Y1XVd66afXTOB
6mGAt0wOL0kpMN1icw/pT5iwTu43xz5mT/VJxSc48ucAMdbLsJoOobZjHwJ/
sKWsF2NAhBV/I5RaYM/knxk+wF1zX0JL3F+WUlgejG+eg4E8BRRRS5PdGZU2
ZQHNlO0lKXQBA71f/hxhZxoeWHgcwQoGlOri2WIENrwKO0Qq48j0tyHJkO4o
IsFbAEQOVL1QCC6+xZy+9B4DShLPysfkZ1E7CzRrPxr2Yixrqu/dLn8bbioz
kYwe+vnhHBExsMVg69FyeSEBzN8gX/b5Kyij5MwjJSCS/GhL5xf7cXisMPJi
sZlwDvAGtQ8E99prcZeSO3jeN6HujSeh3JGvBAr5k++P1WZBgvSXILX1lyoG
j8JBT+gRctl9bi4FW/yx7Olo1biGdjUxFu7Y0QsxBodeH2Kqlnbm2VNFF1l7
JPpsL+bGuqqlRmUzlgzW5CVaqT0C4q0CEEJIhrS5cVbnXzdvmSLF9JwGunKu
sNjoZ67jQNAaffFDwcSZ7vkPa/TzEix43uJkZmYp84DKsfORoGP9bsliGgik
l44Ub0kYu0k+92X4MLLmOzybnMHMTdiXZj1Uq7pJSd1wnXgALqAVOK+nSHif
JliVwKLp8mggPybA9ZatjfM+aA4Sw4BtsFvfCGYq7bO73k+zuA+aKfLYtWIy
qxmpJu3dfa6DzXKNJy8Yu0mMQ5gLPCEEoRtPNyzDfsBgf4gDoW8k1BenOORL
XkzZ3HFM/aZuu4cMnII+wYvoLvPDOJwtLC7MNrXgMn4pgSHODCJai43jzibb
H5IDo/vwjK/nvvYFZc9T8ct1kzUnD39CH4PJ577NZT7ez4V5Il3ZWYrscxkd
SMDzbz4RNt9ieHK8KFEtfkBkBJN5dQ8b1ORX1bQ0mz3gpR2AvMzufO2xgrZt
AKx+guxhgq5f4V/xKt8rrneOBSfBNGi7CKFb//SDWIgHGBGikBrEdJKzPMbp
S3CQjYlzhkFPt2uq/me+CH5Wno6KJ0iNbXO2tX5+C6cU1BiEEXiTgaKI6E2W
gkzSc31WZKotHmEDEJTf8Eu6i47bg8AcAtcw2Q/uzeeT2fc7enzDBG2JGzCi
INRyrAP3gFn6PWQL4JniJz8jrlLsI7H95CHiUTZuW3/ivJvBjmNRGTLFYuhX
VNAGXigFckEHhu2YU+bBkbl4XOkuh1pAgUgO1Fp9M7ox6FMjl0KgppQxqeFb
tk9BkGaMdwrVE97M5VAnGCpWicLEr8+vbT93BqHZFClxQmXZR1P3xYILrQCM
Fx720SaPsDNS867So6+Uv3K6rUQprM4fZwYb4Y7F6kKIAZLUgGeo8pdnV8LW
rJnt18PsT30nUcnGaEjh3qo8sg8U8S4kh9PouT93MpBQl2F7do8IxtBS/i7d
bg+rhme05EYilI6HH5ShEFTF+CT4OrTIeh5BfkpPPyQXCnp3aR+uBjzsGWpC
Yr1uCp9Lp2QyBUFhxniZgU4NJ7l+WTLFf2N9AjtHLCLZBFSIpJMGXM4HDMeO
F3Uuxu30ngtQ6H1bEnXcw4v3UKmsnfUjbzQMO9HAuJQwm7jXMTHeslFLGcBW
Vv0swdt89NqJumeXq1eRVFBbpquu5W/VZg36gCMlwssBj5OGzJgHN5nHNuja
H4skhIZOnqDqKbmse67NrimpnM8P6soYwl0OvZK6Z3sGyB4rGw9ZL3ZmSyoI
blxp/CQRnC3qVxVwlNRw1TKYUXnXZM3BNo8jhsE2JL7YjAL1wsuGroiW1dPR
bSj4UnzMjKT5gcKWi81UgcsxB6Qj5NwOXUx6M3qflEaaequRTPTyx6FhDzBO
qJQaH7LjjofNKAo9cScpvrCOOBcOgNVaYeVJYSIGcf1+o1ZXnbAlgGslyHco
voHp8VsnJAUEQoif8rd6L8iLRj4pxUq9hESOgROziYNSKEXjdf6hX5rczoI/
aKih3bzT77HVceDg9yLx4ggff9AbZzmSyubh84FomHqt08n2HROathiz1R7D
CXNtskgjuIWgQuaHm1yLeop8uk3J+0YKLBadI2WnFq1DlbT40oM7hVWeF5pM
TAyV6yje4QynTLedIZXYwgQJyJbiPDNSYd26sCSdSCVaULDCTumkEs137Qvq
gJ+ru3NP5HeFiS1Bi0YHxk1ytyRlIdg/43JuC6RZM95R7FR1EKkLlgspDQB0
M3Ml7W4U/3LIaokXT5MXsW0m4fb5FIrkmzvcrZzPAnA6UreQ98Pup8ZMFaLL
mt5a9hLwjDq61pKkVO+hav+fjMDEAqEyZrPkTeyJOfRhhEv/ZOi8xAc6EvCX
XDX85UpXWVvBmdevkPvidPe6qigvY9mk2HLUrm3IOIj+buao9jaZt6qYOSLL
jeKAL+QE5GzXDisn9gzVkOSC2v720S5X24MO/x8V9ML6E3jdTh6rt3xZRHOy
48DWX1EGYUsjyYeTtYyRUhPSKodvQOuQZnmc7JiljxG1nd0OXT3DwSOuaTFN
gx2xDW/w8zEPOnn/KwPBB6uxpnZy6Uh7e73DkGfkoZmF0wI8uJDN4MtellXl
F2ZNhJ5W7Izn1/AsY97zPFr92AbdLLCUXWEfV152uoSLX98sCvp4000SIQog
Umns2Pzt3XIy2l5fto8PAjqqQALpXBiyN/vBCrJQw+8aTvR6nuJfWN7ogM2/
q6dgELxpZVCoB7KA/vguoJ1Pa12i/gUbHy77tHu+LB1p3JD27R4IznKFrrAT
PYdyjZP4e6/AZP8SfOwWOuAZX761Bissby1bCmaJZS2PJKgX6uHkh48Rppyq
aQzLAz2sBqIBLH+jNkMUcPEKDI0KPC7CJMxtX1NcladSSpn4jgFFlt2kKazc
yOFzA/etU66WG1K3hUwzREbwL8GhqbFNagT6P7G6iQkR6IhNLc58sRALFw7W
vJVte40Qj3oKDhB+/4oEnCVS+sq+3xiQHI7IghuVmYSzYkoqR6TAeBBvalpH
FAvoQBIVVw7NNK0PGVFckO68m9ZL4AyKW83bdNoyJqF4AMKvna1GWjtkMsXa
odVnCEoMP3KC0o+W41bvD6fDIlcR6wR7KWLTa3dFevGkDxvzjlSNPZlgjSIu
6MSTnQjmILjdTHZRc9RCzug0wLQ0L5ZjOKRJjfM67fj7g73GCaFB35SZG+gD
b5V5hj+Hbf2hOUB+wIxN87cZz1PNptU0vGl3z0NpgSSXgtHr7xaXryJMAlQ7
cheCtx/1a7MVsK80vHz1AR+P8V08rqXspx9IlY9ouAHyxIdwkpY5H4YFZRuj
fYwt+ZeDI++gBsaYWRdCrdI2GdW33Mmwd0YTgFnv2MTnbmxmycSZKNHiVKOd
YvwwNT1QC6XtZPIROoVgwpGOc6Cd0i6WQAU6Skg2croHawGRzy7Z2Mna2ceU
AieBW92r9MieW71WzD0jHm1pcBjvv/vXaocr0QdObXNcK8PyG1dHP9xEJkr6
ionvoLJIE7VAR8N9rNy4unW1N/SDPQzFH8BOOl180DqbVejPWaA165RvCk1F
W6Bi1xrZiD4VX2/jaS9Cdr03hfqS+mHybU4gGlnqDgAq+dDSxx3gN50CoQiV
K2JsKZfjwRw6za+D3yaD8WTCekko8NMat3nbvN4mO9uLc4fE2/ukqJvOr7Hg
r6kllEy6EJ58rd3O04NiURIAevKP4roNApV0BrHDJFwnLBiHAxi0focJFvCd
QQczRGv3CPJSgWP2AYjx2dMAU9d88gCfeNbo7YOap5zGqYFliyO+JdRsnqR1
xiR+6g9QVcjpO7soL2MxJxjC+EHy/8cNUAjmnT+roWD6j9vTkFiFCU01WxUx
P9kmuJ1eKSRe7EE0M9PnuFqu5mTPZCEWnJ5gyQKJ5csgmCR8484DxHrZXR92
ITBKSPJvypFbOTwIeCOvI1PPLTcw6Kx7TnTghITEtJWN4sqL6F2/IGUC7xEB
7ahnvhZXSWnUm6F5MBmlnTZ1im9alusFC9pIuhJn5jRhHOB99eZkqMKEkDsI
hPHKYy48weqKW9UDFkJCLqeXlFzRQptqP3Wo9AfXonV+/NYRkHJE7eIu7Vrq
H4DZSMv0dbgf3Vy+g6rzQjX5yRQY8L4U90RbnzrYoE1PWYxizApwN2W5bsas
thkH8g47qWsNniMGdiEW7HPjrJqqr2PCfzOuZO4LcBprx4/eGcyi8uG7o8oZ
qVdQC6SO0LXBJtTo4Zw5oxKjRJyGQXL7SBaWE8PZa74fCkQSnMZNlrPY+syS
LDDWk6TplfIm4nS0jNKaVGn2jcBq60hBuWObKTh2XZksiJA0ltsYDUIstAFY
LklCpX1XyQdTBH2AKox2cPyhcXuZpXna/IPt0i5uhvgGEARONF0QTiQRozLa
XTN8HcKoneqdt406f6RMLTxAGnA8USoH2nNCADFOvWAcJ5UDdV7QBzgIcxFX
9Flqj8/aQeUDll5fouVUShsAl8GCdaWckZNcnuh1uJmoKg6sOAlPM/WSO8tO
JnUbNjH0oDqNid39Ua5NPgVnNLcWKnEV680bJ9zqx0/5xwBFRwaGLHHVjSnm
P89hA+F4BhSFwDgrwgvh83ok31VzfoZcYDv2+3y/fbgAyBlY8gsv3GXfYVa3
mZNXHKjeFRCk0F+B/Xce4YqV4Io+PpzMI7DE7uzxVCiQADN6ej4NUvC0/5Fr
fLMtJmyS0vKwLU0VHBfpMOTveMl785QTwZTI61LxRea1lRmrlJ11rR/PLM49
jgDgtByPS4eECQfwdGPLZUagzdtZ0qPLMmpZ//oaEySK3k1xFye2+81gFLnO
8XIEnI8iJQAyfpK39xfTWvL1bHh1On0niRpsUqoky6/zw9UBruEDC0BwdrUJ
K3eJGUSzm6jKkNGUW1auRZ2dseI56Qg9yL07TDvFN/Hzd7/VvMa8yNgxg+IV
faA8XotQkZ7VK1AEuR/DxsXmeo6qZv5OBxIUMIL5hWsJVacipEIC8nDZXQZ3
T/iOa40k4tB5/zxm42sIlDkasos/4x2xmAc99dVPq6ckG/ZHHNH6Dx4/OKP2
I4L3EKJWKR2Il+RzGqkQaX5ahY+5sKcsEQbeuF6abXHLwtyL5EbQOvhi/7Hp
hL5Ba40ZZWCxm3pQj/TdXXb2PulZ4ZF3sUT+zlf0vRa9WDEpphqDoeFkKWF9
U+t1XpctXYHBQdrT2QTsKbyoPj64Br5/lDz2+iu5T7XjMuLxKolGObXNSrKf
xYtjp4BHqNC1imBJPB/vXc7mATHvmfVdKGA8KRdJNiP/+q96XKHQEQhevD3O
pphqqk2fDWZN65wKeeGgk/jSyCBjOt5gKzIb94GNS9ecog19hb5ZCQ78KetX
ollTwLu3xu3TI/Er8TNwXvkjpihc213aXfhQcqV473Wa5LXyisr7stN9AV4O
NrIpnSKdsrIMmqXKi5vD7Yx8FAzLNBmXV/IGfa0PDDRmOFv14GBOXmd4s7Af
uoCD4Ekppw3Vusx/IpDYQdkgwHLHq8F4FCA3ZVysqDN0PrtMC8B/G1dNBEo0
7egcPb4r/yk7DJF6hU8Hg6uM15eBu3w88K/qR6E67i8E81giXpeiPZJnm75P
2T1oQkCLS+64YBwQFrnelM3AUQK8Mm/l0648GQUHYQ+pO7/gScmWSW3LvIfC
wA+LEUVCRxXZ9L0eXyV4A0iiFxTcdPdm027FnyoOm3gJH2M17/9Ht8osdlu0
okfTQakKGm7jgP/OJqbIpJaDO7w8/HXy9ELYpJmkzkCmiA92/Ac4kEqzsICS
CeChFws5jd/zpq74XzwJIql8O/C2KgXIpTeSa+oRdMDEI5xZ1R+uBoiEr+Rq
5DEAdTyKv7OAmfC4ST1Vc1wtsFFISOs011p8Eo9prHy9MlvmQ9Ndph2SNosS
g89tkUXWAodl2AXvoBzSu/xHiXQ+7nQ8UmPjcWdg60s1oFyJvBlH7RplUz9Q
J9lMrzcjUfuco/Dih14bfQDrvSezIgxm3Ykbr3E5JlIVYXhk9k7mPucY41ci
guyfrC0SI2p7tJHGfmji8CcOh+ji7AlYdMIGz7nKOZNjuf4dOdXJtlncIs9S
A+NHQj5QXj0i1nfYbAhWtGU7/xRF719azmWZVv/33A0xl7xJ161tKuMxR5N3
gSjX57uM/tlX4JKasuPMfvlImcOf0EZCTgM6QUWPA/FF+v4X0dP85wn53VAa
kmugnjjKNJhoME2dC+yYz4f7rp5y82CYP+4sfz/kFfAQRUnfSLVnGu/NcIs/
QSDpFEqMVQEFj8F1QNMlE8gnZRvgN4fwUjqbYomfvsLGa/hQO+fO/9rKI6dd
03vuL3q5KkPfi6CFxvkxJmq0ID8isD/eGthKAgSpFPsH8A61obL4waOfa5WT
6kAiq35SIf5vvziysGD7so0/9RhAyWFtWy3ORDrt0Kil2oi1JBaeAp6B4atR
1cEIgZMlV9NzqSkEIdIjhFk6x00YE+8xR+A0uTNsoGvmz8VFfgIpvQEjwNsr
opUPmZLrFuFs+a3RLbeRazT24Mna3Yik0bErbu63XgQJP2xlATfNM4sHZEdH
a27UD4P/KLSBKDEMmpk3PujBTNdkB6BPCK0CAeLc48szPO7fZK7QLZPOv/5/
4iI+z2zls6lhMFB1g7KcYlEKNluIK+g3iyW3YFxKnlgSw/tGrjUUSDLeJqez
Ho7pyzJs3XpvOVMU1VgO97qaQRCm3kZc8Vv3B2eBHqz4yQ4509ecP1cTQxAV
7eb4/QIIiYGdNkwLWe4DvtZ3nmS4pjueLbi5DC8eO67qQP1JBsGdyvEs4rUR
XrqLnUQzl102+gLOvUWIpCz+qrLWzghRCep1uQ73WwhMwKnAdIP342KCvPsP
5z/Ar9F5B114i8abz7GyvZ3EcR4jVP1znwI0XYIGQiBJGDDmH7ueui1rShsT
fOM3IUx+rEmZAfdYGwS2RxFdNWYFJcaBfZhC8rK1Z2EciAvSFvs3DIQ2vmUT
O+/06gV79tFQOw7Vnje74/aURwUACHvSR+CW1MLBc3/oo3rwmqPvOcYB3mHH
cUFUNI6wWlwY/p2EboY1eADECVhetNbiwTMsUw+srHPODSyni/ipcDwEgNh0
M5D2YLXlEF75xq5P/fbtfzpsyPjTlvL90IINvMMKgPM6AWTLaIcbjPk5o61w
0Yla5SgLELdEWBGXeKJBd20u6EtgbpnKNyI2RgrCH9BlMCxe7RdRVblFt+hq
MwNi6robELHsyhTOzH9Ci665kbpNMVVXf25Ow/nZkEQ29uCFptzhQwMDhKEw
Gy7UefzXLXCm/Uz9IItiYK0Yvo1HT2bgjcAgLdGzkzIKWQO1xFa+PePslIC/
1iCqmTLVj+m2ts20s5vPBOIc4ySZQnUhjrykqg9iw7tw/XVst0Y1iujlNQd0
3F28TZErgP9N5KMKCEANvPHSXknBpu4hiImLti8tetv/5SgEstpNRJxz/eWC
zjo4KodchPfGiGRde99Z2tCD32wr8Z8f0gqFy8z54a2Ca+SY6o/mfV3BK4W7
Pzfs83eXpseArw6VPBnOX8C7LSHnQE+7LnBBYDwlhYrUerpb4fQAU0K7BEju
/MIwgUfXMzW9lQ6xoYbzL1Hk3rm16CEGeYFinCN1Noqb9VmmOC/hkczLn+kk
xHHJb5D3G0IgRCAvYEjqgWA0W2EI1jO1wXZpsn5T/gWhaOvLR65VJnvYL692
W1jk9zDLj79liO8jL/rodN7AYW4CFRMlpP9L3x4Kb8VRK2CFo8i4g5g7BPYa
mixY7BoVD/PKg1yW/KlEqlDm8Bbthkre3Z1+sq7T6RiWgB6imup7aGXh8Uac
QMb3h9Aou5Ns+HNG4FyhB3AwtE5Hr83Dj/R/EBaNfKVUODkf5UuhDDl7v+2W
vHml2mawCJM4egn6ia9o7Izm9FeHIzUIgRvhS95I51AVIIEz0vBE6MZpbw6M
WmZ0GUCej0NUcRQAomVMChEL9T2tg8nQYRNBfIgIT5KjWanKdEROqgAM3tU+
hG51ZPFsh9m5U3stOMK3dJ/QpnVmSpwFZWyK88C7GBVzkmpGwQaZ1nf3R16k
D7k7/gYdk6WoexY11xWuCMP660M1FZZQGcLQos5NXCAiLFKrZhkEFwVxGKRR
PFzjp1O45/3gOt6VebZvMt1CMg+ekyQULhbPA8loLvbziW2fPDX4Ri82cMDZ
AG+SBzEPXOfDMX5JjJUbgog7w/HnOYxKd/Vf+ssrzGfMhlAF9b0UOrHIZBRh
5iraowb42dTxYs5Lb8Y/RvNqcW7KUFjrAszY8n0+92k6AE+eC1hVwZN9lsAF
WFOgyxeYMLhYxB/5podpksRvSQrkf4a798TgpA6TSqqrAwrmwpXOs6TMONNn
05usYIYZu5in8K7IoCH1lZ+6SdhBc8ZhDrpF9eLZtaCyqzbzvqNFMvLVpqxN
JO3mHBAZ9fNTURlXMmuWG28BVdKXtk2wxMM5LH7gt8CfuuUrIpisamwoqQSx
lU9gP023umn+F/K32S/+ROrTz85/3UuiKHMaps+HZthg2XRzlF6vmpWwAkmD
8TmqClaQ/vFkR4LGGu2CG2lAN7WnaKi/G4jnZ57AORQh57ujoHlJkuNkq4HA
y0BZb2xtlhdXmM3RAK54VPj/G+22IAPcJc/4zO19ehe5FmLOr1y+xcQKpE1C
HnY7Yr6KRJQTqUSh33oJ0o/WNn5KYS75R0REHTtAHOPvq9uujDZJwjBf6Nfc
PRSIBzHOuJ/c20qXN62pbyhRTRdbUrHRjRHrBQApk4uqe3w6qqOE+QRoDzYC
0L3QwJ/2i7qQuAIbr3tLM6kCQISbQE11fnkX4+yBDNlQR/H+GPCZJWMGU2Ia
5U7lKs196crqJc7zEvw4zDFMP3TRjxB84X661N+P/vW0+ek12RlRIx4tlwjs
NEoskxJ9mSR5YoAtZ1eN3+59GarToy0cbKa5uI/v+7hMHg19bRxpTbw9YufN
c4TQK6+e5CUD6jeBn1na774fk/xfJskbTs7J75sAsogNeKol30JRJe4XpkP0
hfLPp90Mx1NzDH8jagbZapqoGwm97RTy0upKjUIQ8MWPabdD4lSICBBrMClb
MBMwCFu9pWgu0nVhNcYL5Ihkkgx9noHXWMOs3jvHQVa2FvHUjZTYkmYDj0u5
p9K0O95I79/X1ugZeDiff96P1XRLYIagV4weOohAZU0BsWh0fUkf7WRPG3D4
na//KgNQ944RIYDKlHbW8VOC8EU7GRVDKztfrljmJ6KGZc1+pB9sFeHO2iIE
xbve/UBc1tV1en7//ip8ZIw1fZLqlRp9yXu/xcOenvBF4YtcggQBr3u6WwVN
QW+kQO5b0+nGmfVaJAIpn8vuWNq8JDS1Gg2Meqpjl66wi0RW4OQ6INNAz3Uz
hHyC+GRD2O8U25PK5pEBSQWJLX4/fiY6yJKWzPWXmarJgc5Czl2w3vOYeJgC
IpCvUiV3lbVwfca+2gTaCR9y80eJielzvLxQXhfro3VHPKrW5JB8Jc6lyt81
gG8/KNe80GVy4O/wOMYe22KvtKiBc5QHQySqnmp1h2tDogpQcfvKHDPuAS0C
CWbZ/tx8Y3+N4cRJMc4hg0U5/n6jVuw1Q8S1xtgqLhWNTle+8/5b/szA58Dw
voKfGxvcg5LM1y+v7E1QnGkels6WMBLqsSH0cDHf8z3oItJaaedq+1m7Hf3u
C9zR1+cD03CdTiFvYYqC/T/M3SB+CL7crq7FSxkS5C3sD4pjY/wcznpK6qvF
bS4rA8sLrI0anna/J1UPNdv2MvmxwkxWOmtgeroSzmDbXfk6R0QJNRWyWtjr
VWt4IVERRmxQnRnQvXYFE+iF/19EukWpyWPBoGoM/L8YKi3djme8ST5SkPrA
joysIpX6vcLfxtOSuqjCnR4+hXaFE68SQygsOnxA1iO27XFmn0z/GDK6tJ7Q
LolbL3iWyrY3Wk6IBjYj6pSZ8YaJgIcxOCYKDGCvquQdaylHIhOlFBu2enwD
qwTF65Jg/3zgYQpDa6O69RmfHc4ql4mmG+9HErFGKpVz77mh0YhpB9/NiZKI
Evz0R55ufORj3vk0U6R5kQqDfJ5XTSLezmzm+I/jeWwNn0vq6u/1xB9d5Fef
EneCDCRZ7vsoFornNCA8ptbFaBNUhTgeX//JCa8T8JeKpzTYrNfyHB/3xNd9
qnI8t/JCWDrCygebZZk5+qgPIh5hkfnJUh8/82yxw+BDocQRGw+EImn2K6ew
8kQUbiotGF5Nro8BxGYyCwjZapa+uYWNTxNtTLyXXC+9jyxAu4/3TZQ3PM/x
YifFblq5AAU4OBKYF/+x7G1RfNaEQO5LsH/inN3Te6s4xK8MOl4zneqDdAxA
dJ3ekbyD9+8vS3+0B2GOWBwBSA8IGbmsjpnWKDbNUnPCmc+yT0YIlstAp6al
pqtIB5GnvSXK6J+Kz+moNdME498BqiIThf6miDruQCgC+NEglNeC27IUQb6U
qlM36r0mWwuWmtCYICWdN4EJJSGGM7NH//qrDYKQk+7bAxrylqXaQ+u3AEIY
eNpPfEpib+LJwfotTi/uTwTL3D7QIpJ5vd8AJJew7W8utcMqg2RFoEIOWyTt
VWXaTmlYL9iKWFwKnsSkm4Aa6wNhEHWBWqIeAhUXbh3wHYYirlyrjsdcgizd
PfFTmrpsK2xzMh7d1ZTdiM4lekQKHzszpYk8gxVoec4mW4qEPn8rOaBwbo+z
ETLzUBmnwL+RnqMpPJNxw9xHxWNtHreRbfMBpP0M4umrKz7fbrKyQbNkDiOe
Z9Z0Nxp4v8/AlLA3Rvmbn7mtN+SSBgXQ+5D7vCuPCU5MuA6l/hdejgH75oop
BEmwNITjG7d5zlGJvg2pW+ITEOc/We8GZSk5RwMfqpXK3uNvTSsxXngEBd09
tN6JvFh2r/wPS81WDlGjtenzRdYnTkbnSB+a1HegpKh7WGCeEFwynJWAkCYD
wYknbzpNsytyt8QqYrRYRl9JQ5GGRiogScgqaSWdwRJv9PVS8/DCgWPVq++L
wZSe81uaUc7hHD5wpJ2haJo/rtU5pCJcvkRcXkaUESUI7fx3EWQgNofizllS
jkD2aW4lNyVIyYVWtk394U9ESP1q55djJI4GOHBNNwO3MPVXdxGwIQHFydK3
mHarWuDdEg2fDRFWR81R1LoggszhMkgj2rPjUmOc75YosXtJFnHJkFnQxIqn
tb8WSrq+TC//UgycI3lxDpZ6ymQJFVLwqacLHx54hFND3p7YBAW14ubCYjRZ
Oh29w259iixWtax7Y/W0LIk9PflnxlMq5EIngNzxrTVFdWpMhWoaKu8s0tAw
EULCeED4/ZkGPKohd6vxMoDv17kABlqwFkCyLXtHsCrcAbGWoewoQ50qN4Ea
2ewlnRMEau2pqggr9YvuD2F6/LAl8zK/uHFEKF5jCY9FA1Er5GTx8BCiq2L7
aYAWPQnznCp9uN1eflfCwVkHWXdg3R6eiE7TeTgE6cTBvAKVmYRPPHwk+pPs
SVZyINcDX+tFn13+X/SWFfMVKDRu5DL8JRnZ/ZSm2DMK02aH6gQ79mlLD6vo
AnFCwuZT46IBsEVg1epQ4JJQr1s3w1UFhpNH+sa/QyyYKkin7Ddu13qXSQSC
tkPsKiboDv29OSQ55TaVlZcg0LMiSsB5qmk1p5ZQcXkys2Tw3aP7z4D83j59
w1K7mUrnSegu+zxxdbeci12XdWwcnOliUm6sGulbnf9SD+dk9A+lsgI0iQXb
T3e9hZ0agVweQ3CcaiM9GZ94YCCce1T59GvDBebnuiN9U00AIVYOvXLqMu7l
MgS4JBwtDrlTGX3wtMzHlK4sjL+vjuvtOVx+Ev4WCeg15JHLY59rQsKjH69w
XoWjkAwK20SvS14KjFXgzqHWFxGbmeDHrFwbsOSmtfsMNCJuARwlzMFhGNLq
27/z9ZyXkbwBShLHOmTubnQ1foQCelS2Zl0Dy1WaGDyF1cQkREpyAqu+A6hl
KsrvHe8OW22DEAyKdxKqOzKYDF1X9fJP6rME9QdKwJuiHjyCLZq79r+OmLEZ
18OuqEaghL4epwivsiEelqZjRqn57Lqf+kX01LiMkDC/i4iDbtUra/YGs6Hh
b2OgJ0pPZ2AV+8FqeSkzmVTQCrmXzipLs6+hshlGzRVZHGN2JASUgwRxtORE
JJD9zqsTrpJCwAspPIvAWjW2QhqvsNMrv9N22a58Q7sgXNqljXOy7j7g8E/F
BD9FLHzrJoRDVg1k5GoKCjVq6Gb9zplhaJKeJeaesqDiTxPbK80cGPWMMlAP
e1lgS+SeFFVAag9X0iXnTn2o8jG1wtHLpZ4WP9SsS9JAEmG+zvWixK2yjdjJ
d9E5Rb0U6lyZsw35WS5GafM33sl1RiHacbnealFJfPHCyu/GsxAFtag8XtKy
vzdb/LzksLigWSsUEheJ2tAcxSvM4J60YzfGAIhU4xydj8lBMzHPXbCZ7tFj
dGRsuE5flPBZB7TCeW1lC3fSiwNy+CnUqXHeDwlr75eLjC5wKoUo0NW85+c1
sm4BSNpXnkWrFI8LM/jAdqI+i6xbV9WjHrmXoL5mnA8eaJ0tPOrLcaaID5We
Gl5+HH5vAIZssys/DJHOSs4VJHLl2jj5quhYPR2Rv0tyCm7OShAMp1diCxlP
DIa86x9+a4WpZXkoY8KFBtwUidMvVq10noqRDXRIzfimlodobJHOkLae4LQh
p672wlN9Bf2at4AnM/Zk3fPY1ghvs5P4KpSjWR9o4BRMSB8RvobPO4XSe81n
Ls30XL5oDkotw/+QvBcP1rOOR4qiNPwF6vhXe4wgZx8Ac0QJBBwpEyljXSir
R1hRjpJTwYIjJlBWr5L6ILEWusqrEwAbqGWw2iv2J9IZlpm0THEq2KbeAie2
ZHy3Iq2bMHCOXvH3GR7i3Ju8nXPyzKfDb9ZHtdPtJ0rhixGDepXZ23v8tkAJ
T0CQpzSfmzyhGjH1CWSNdsllLtmFJ3SWodUuDxK0oKT8pYmLeKPusUaATnxF
K1KhbTaHNUZgxdJaGKJc+KEvwSgot6frXPAJRwIHwss8dW5G6oc7avBr9MCY
r3R9dXQfugVBz5KgUmvtPn9mY6em+gpcdgQgxyaRocGAnSbkKcCvyGPkHh97
n9SZMx7hC65SQ5W7RxmVtnuduGCjGI+mQ5mQlUcS+JH0cysys6R0AyHZoj+x
7/e96Yqym8i2MUAOkDhty0mbqbsOiIiqG3GVu8Kt65+v7TfHtbpxN7IDVjHD
rrs3Imqu6zxnwDUlMIM2kUwb/BySDtdOSQBcsD6F4AaKuTT9100gHuJXwrJJ
aZD8423HoAdVsDlc92u28xjfatUT2QArDRUPfX9yqtlyzivPUHMwD2E84QXd
uG8Zg8SaKxRhk9uLm1fpTW+NsWzSnhoUBUT5enyDyUJojFRgO2Eq1ilc4fr/
VhjfbXpFFYhOhcDQIBDo7SLNgkBI0PA3nBVXHg7f1XksGHYizfTYHOPm/ibS
kKZGd3SDYPzylN+o7IxxA17kRSFHdJLjYCpImLBmj7k9ZcgHCLVup/MtkXqP
nYKADSwIy0XAaE5WwvaIN2zER1zjobVlmVpBJnilXsXU1wbvphqe6CVL7D48
AebSpD2XtuQ98ZzRD578wHGD4ptVWMTyBlfUv8B9e+TkrB5JZot9aK39/j0j
X8zACoXHy6xLeXaU53QbXBca9kZhaUz/oXHBVsZUN8tBzHrs9TfFWxWvmpYC
9+LooJkZRhZeLzrHTOS6MT1Ep2WL9Cneiv8HS4AHDT2/9pelJNI6oIB17fVO
sOL5Z2E/M4AeeAaaqV/EGy71JIPF78dJ/oPHueu4XC8UlDxe8ZaQY7HeycBV
U19zIWb9ieMjKfSN6js9Z71mFDNBTow8Y1YsCIrQyRj6CpTAG+yb563HuH8b
ZfPKpG/VV2ZzlhxMEtA8FlUaPVPAtvAhDAaMOS77DMmvBhRGsi/aSkLESu9Z
ynCuH4k+ZC157qgpl7v5VTfrxMESKd3eywVD0qkzD4tKWQlN9IW3T3HjDtPx
YjG5UOL5hBfEkN8TSFB8zcdNG81Aa9XAUPmK4xU+yy8EyQ0Na5XXo9/ETr+4
jbBsVp6AppMhTfRGzyY+eVLxKrvgZFe93VkgoKj3tm7QodzPoCxoDFOiVpWZ
/F15ArO1KjSHkxeXF0G5HWRAkbgWwYPwteGTTtglcue+kEmQfWnkKA/s1wG7
COA8PDoJ0eD3+NbVE+ca6txDterY5lCk891KAAB4pQYVcdtYai9bmGtIbj1R
rNXoBIzqNDhr30aVb6sHFZ+neoRPbC8zMg2h7C9BaciiwywrZVaNBc8MgzDZ
BjUaQQOPa4NffMqI8iGI/pS/50tmlExv3Ekbw8j3kVg1G/71cKNBGPj5dA5L
cYuUuOAcfGA9sLaB03opVA+h3W4e4w+YTKw9SV1xXEiHHc2Zk+9rY13bKZ3u
OWRFKbvUCu5/r+X+iwFttDgidDWafkzmbmoNYgzJDymFtDPHrRxxO82UT16D
loH5uZW8gyjIw/OPREz7PGC1cltrYhxTMYHvaCwR9Z8jlrjQbcL1Ys5kKBPT
GIOQCbkaVlmzeIPZUkZmc3N9Uq/4CHBm7g+7eHCPZNjrzu/3eNfKzVdeAxL8
+2Jrel6qt6agrx8rNS1Bm9X2ps3Lbot5EL1ZdVg1Gdp1r5dVJ6mJ5AXzOP+g
VxAWVNvxUBnkJxECRoTco6mRkJ3QTbXKJdtFIXSUVaR96oQhT/27vDb1wLb6
hYdY68iuyGekzkLMkQuNzU55eAl8D9bOPzr621D+i0UtfrNSrMceCpzR5wDP
BaNxejcq+MGM3mGdWFYzBsp/m+hl/X+w4dyO54n75cWnMXQoio/fOOPQDrZi
EIzC7xdB9qRIz/v8RObUsPtrq+cP1j49LYzuICxZgRPoFda1ndjYBaRS0OnP
ePJ4OuT+lBztLTthKzFrI7boqS7mVM39oHy0JQnd4KsldT0da3q8veLloyVq
x/lvs5ILcv2kMdGcs0D7DrEHzn9TSCuGrNQ0O4cJKF/WD/SED7oOdSY6vaI9
47hV31Z/8VKKdjAp4oPp9mDwsB9b/x2XUp/8lLpsJN7RIRaa8nCDgEpVly/4
9XumWYU0UNMs0oUfRqcfxA3WFZpon2s6nR4vYm/QXAI6u5vYx293fo6WatGK
7SSTdUETiGEMqCnn2p5l1b+aUHqtUrox8MtJrNaAgzFn5GkNPUZQvn1Ead25
NrXEIbFoDXkutsmyeCRy58HrYAtm/ZB5MObEAljADPS9UGSBD+/kqf2EM/+J
bYLKn/WfBlqITAPLj9VV8S3nU8nrZcMu4I2P9kjnQNrcXrHimqUqkFfXon12
6ZTpzjG42BHacjeAuGErg+Ec9cCIk9plPlZdxOLgbgQ6j+xycCOBohMoypMm
E+6uXmnH8o4qn+zMsJYYNiGExCRSx4jTc4RqF5WFY5aeDhkJrLqyQHW8SEEv
p0GB2aBOF6Dlg6zUl5KVfwum4P0+powALAOWsstSlqaVlzm8dZnpngW1eW8I
nrvfUaj6Uv0GbPUCG/csEcR3f0ZNetZRi1tnB6t2a3s8cAu7u7vWgjUJHbYm
h23/YE5UsQiqYFbWlD8eBWiVfU++eUFmTHe8UVIVsyaiJPj7Xg5ooDnluagk
LKIPzao8z5w0FHkHG4cBb0Lp/asKjB/LrGoQB1ZB55uSHLBbJ1N4gLzRhzvc
AonbJgUIw5QuQ3Cs3uLYcGgaS5GCf0sd/h/y3L4oCVFlZl2j+ykMlWXztOmH
k5cYL6+eP1HmFz4dnu8zDAlTfC1RdBqifaAMwdmq1DpwAri8wdbtO660YGR2
VGXrZ1fh4uCZceImhOJKW9YeebXVB+b5tRBD6Xz/48n0WGLSk6zycpsPFGE2
efU9S8nr8JeByPR1O41F5Se20JgI/X6Wpc5StNtD6lUf57LocAMnA1wFkYTP
tYEcirPY5Cb2zV00CBzBFAnx2mTq64ITZo85eK82CZ3Gt0O87ujQwVdcMRwc
MlGLo1dOfWlWchwk45yF4CzLZXrtlwN+D+RdG43aQ4eVnxgcq9p2Aj1QyrVN
Ubf+97GhUAosYVwrduDT5ldUOcc9ez2ibVV40nsDDGRMHaL88DmavZTTMNHf
DbfZeMAMXgn8mYwd8+EpYhBy3iBTYDnCOekjr9IPZLXa0gkUs++knkncXn0t
RzOvjK0iFeH/va0fLux1uTTLnwP4OS7kdm2hAKcrPJw5DHzcstXZh1klW5rz
NGr74SNo74pHkD8xx+AWNQmNhQP7zkHcRwXISwhUeQRil2D1kz/g/uDnhNfC
KK9k2EfHQsrMu+/lGgD+PtRGWQIlrHfb8NB7WWl872rHqEmYqyY2dMRnkEn7
SIcEneu4+fMp8JB7+zNsf87hudBBy66PleNNC/TiHk2itGlFkyZ4TzIUq967
6YFv/EuL0F2R+KadzxwmWx27HuYyCOvT033M1M8y6pTPhlgosTDDkj93MUqA
KDXPnoedmn0N4FqMhuyV+xkWN2qyUx9RNYbeKfd8ZMaahyn2JmI9EVHM0Qpx
o682/drGGs1QL6I8nGR+LityJgAkXh8W3KDfMIP2HF7WAiPTNLZbNuFFKlRL
3N0vC6u7mQbj8TE1qHZFfwlP0rdn+4rFLVRT5VyRnglZ7eu4iNqBaWZJBUf7
q62P7nlCVMHPJqOlKeb/8A5cJy7Z/FC/h8tdnmCLJ0kKUDIcXKHFOwAXa19F
0CFMjqV9oqiT0Hm8b+v7pZod0v1eMFLPxsMVg8e4MFcwWZA6307dp4H/bUDO
lqSFwVFmkP2Z/wsvni7wGkfN92p5pyt+RTIuijphzD6T2/xIiE+l1kqLNHzz
QeCs4CLDyu+enBDNL6zytTqK9gcJkMQRsQ2ozqj8LPyIYvOnc7p9KY6J90Q1
Q/Zwul+89JVYT3qlw7U8MSgEKECkjn02lVdjsu8whwygDBFWg4Y24JNNP3eV
K/3LBOk/VGOT5+V20zvAhokCPPGJAlkfokdWizoxmxhwxJnKRaNZGLXUzqJ9
sbiDXdMrd2vdbS4HJ5QMOQpWaNSsRH/KmwdIGZgQi+K65DJTK/49ip3h6Sdn
c7Nbg8L66hYy3s3iM11ZbU5l5pALRGfT5MVa7isWN8WXgR4Wb0hTHjXJRdCX
LuVuWApJDg8pI+f/umsCGCmrXBQtC5rrVM1dRNRgmdwDSTXAvKPT9qjPcWRG
7iU8kiJA9XqNAr4/8IjpMnmq+5lHrDLFHoRMRLk3CBHFppZr4vXbZIjuEAid
DaD5K5ppFpX7tjE2ib2tH0uLzwsVIZvLKkTYBH/6dWRZ1cTeX+VnBBYW76jD
srIF8TMC2venfJwosdUCw/9tBj8lly7h9ieN/uSOrVgd6zNpUCRaHgjTDu2r
HYcFsGLAbttNT1H8DZ05IVZHmbFdjXKufmuv2kDMIyOeo6VSoKPqhsD0RT84
eex9SAz0GoVg6PijgOP+d1DK03EN51TsE1LgxwVlyCKYkrJFJ83TvbihaYYi
X5AapCH5ila4uFtV8JCfWuJQLxMgHEVsC6Nu5M4J3adKRCjBXWnGBiGhuLMk
aXaFlCGVjaebo9JD7xu1zEXxdE7I0hx71bLfMcUOzwj0Mwb4vQiSVslLjJgG
6eaANhs4B/yBWprvfUCQXo4vid+wuUMKsIQboSFpOXT+TOdCKo/Rr6p7T6Zf
861BzKcgpPV94dKO5KiUsy4lx1nqPwZE4M5sdMI5Wdn0TT3JO/aX9+iRRRPn
2FuqRPaIuFdOMzdX1gsE4lh6zMWBV+YlUSm/fg9FsPd2SOBklbysHphSmd/G
ia6pfHZJuZOcWChZL6mJJsmUz8gv2UY/G3nCSQ1nVzAhkJ+nODpPZCG2PoWP
R9HL7C8Vm86qVn7xtpO/dacQN/X3m3qVQobbVJadN1aEPD3BHM6zm/JkZT/c
3m30Re8iUoYnMmjOmTOTI5f1WZtztyFABebbboEWBxtumqTdJiOYhiunkELy
cg0HilKDn7eOKNHQL1T39wNl2gfhj9Dh4JTZJKEMIcCIKYsiDKVP/1AyROm0
hSFcADnZNj3wA1MWpJ39kHYFU6tE9W646Due9qGw6TvFRMtrjvtPjTLeb8Kp
JNCqB0peLKA8vwWmUiyebh0/j4ynDhUMIZy7rZNoROcEt2YkH4rDMJwI1459
BfEKkARyJGHRStk3FMhafmzDKNC+qcfVw5tjuVJ25DFQ5OWUeOuFCMY1O3ko
WAsLr+ilACbhmYpPqLpjFER9IrqrH2WqfzmcGmjSj2BoUGbqY4Be9wPz97Ri
yIQfIYawgPN71uU1n9jxb+YRvmTqEgY06/ME3maHVNTsy1GQCJxdmWKs6NG7
J4mxxPeXlzxUOBd49MjlzxhXVpbwKo34bwBm9q5UOHYCB4KiZq757cE0+/0P
bR3A1ammQCTqb4KbP9XNIrU8bMzZGzC2wtKxfZks0jFw+C1s/5JqSZ3dQmTF
wOwBPHjSZmUVmlsDcPIJQVKJt8uvgICNpDSwusIYqgxnPo+hCoTw5UCgjjgV
R4ROCjefQtWnb3ycl8YIUgskGZpPTqqiWcC/g7UF3kUDlzXCEDR/BWjJiDTg
unkEhIV2BnMi/nH/9+BDyw2ljsvMfjnWCM9rIYM8Zn0GBGsDrwumFlMWBbG/
4DxYsAg99M1S6rfT6Ia1EA/eNhPsDZX4e7ewJoRbczwhSX+L4c/4HbOZGfWh
b3im8+Su1duRwSn2rgIV9sIN22iaLh208XQ1eRvh7/Lna/M/Bssun0KyikND
x8GrYShl0vKUOUpSwpY7GZpfMKKkyyXDGrvJULzO96p+tg4w+DmqPKAt/WBb
Fcf26Sgu/Jnf8DIupSvRegi1DJJxMdX7k8BreIuP+glop/0SwZ+l25JDCskk
cEG8C/1UwKpzeCUycqMyZBdZ04VOIr50s/BsAwtqmIg6g6tpvOeV4N9kIgf4
uETFZJMB7SKDSI49uHDSId4o822I6F7VR/1z7rPvmr94fbqQc4zzea+JRqmJ
I56F+jyHHno/8Y7OGl26ipKQmoLKFNXvoC1eNmmiRBXMZ164BgbPlMmFCQLg
DLUAVNwKMO5dWxV6u2u17pnYNxRaozp9XV6DNo75ctwFxXDsUQQ2Rps5chfL
3lnIgCxX36bWUfNN/GUa7dpxU2CAMgfv2q37w1eZrojfCWRr4vOcxAyjnHgI
2ejP8kyqUE4WxllGDqk014DpQcpP0rbGwmbti9uoHWmvWslb4EUnS1H4xejd
xtKiUixrv+ZiFlj2Ngd1Nrm37TdMZ53CafPaUvEvLWExylVpTscYlZXf31+6
4c+t0aS/pZmgYl0fBxMZ4rXfRF9+J61q6rusQ7d2ED9r1flQQBpYS82M9cax
R1ipUnRDO/3OaTIgVf++EUDmJWiUwUkYYeYZGyeymCgoUcL6RZi8qsizHYqS
LA5Yb5B1fh2KRbndaSVq33e3P+B2sZJiYJ3grha+F/HMcVoJq58soUwRIV3R
CJ84tng8H/66ZCff7AHAo8LeCXid48Lv4DiDexPJgIY1Dh+M0ANZzVhTXagl
cuqln4dem3RhRABji39yGiC55cL1LemMB6K/f7GcIWtgMCok9ER7Q1tnUr1x
M5k6gbFeSwQTSFULhdW+cV6Ruxgopgle4DDbLH6TJrDGZps8rb/IVMMUQOk6
pTTNp2PpgUF//47VIFb4L0Qp8yHmmjb6AmqbaR1/SP6m/GH5bAjHRQQqIuK1
9ftnvkWgYLp0JhyljpsLCzcG3CLsEJIbGcUk9mnTZG5f2lp7EwUJttpOG/iy
gTWVlzCf/70szJUZ3trthjox4+FIBcTY+SmROI3mJnPClj4YHp6qXYvftXMc
8TxZw1T6aAyqesbJIeiM6MxmvHl8+X/+0p2ibj9PBniKUxkUK8xHzlXRIXkL
WyZJigvnOCaNV6ISDGCm2oT1izucmESE9nvEqFFaFP3x3mrn5c8uEQOFQbp+
s5UrH43QS8I4cmKl8ELY+bnGM9d+mH7eNNand6uo4cFzWRKRYaN2Hcr5NPP9
c/6QB7f/Gh0LXmNoi/oq8txbBmbrZx77Oa9CNVPESLHzjpkerYbEe7axUlWt
1f9sRZ7L7e2H2hcw/iAghHwDDZxhjefeG0Tr9dCHIuWrtCi/gaTnnGFuJG08
DFLxa/wXQGOMlQSPwFtjw39wHWvGgoA9+A6hvcH+usDhEsZ4Kvpignk4sl7X
89A3r8rbKIeuGEsvlV1npC3RTKjw3oDg7B6mwPBafKP4YxRqW6NwpbEQNdh9
0/G5kySdZoGia4Nit1eVB6A7vZ36nh3AHpccC8N+ayyMTS5Eis20kjY3KlUi
NBodFdmiwueVjF7z5g+Tygnbbk4MFY/VzJp7aIo2zibj7+w5Z0tt+iwGFWsJ
Ed9QBhgmq1Hpcbzal5J9dDBcFe/hQG9j07mrxZfBmI+iLXgfAby2XSP1Atar
QfZKWfV4kS6ayxoWqK14GcEzY8pM0ihuEQpRJOVQF8xfKPh8Z1zwmb4aop1O
evQDyR3Jw1+j0n8Rj93XIlPuvxDVBN47zEixA10bOLQG7O/GthmuQhD9G4bM
DiiVHxCyvnyZFPb2Plvsca9pF8XyIZn3TqiM1KjvruFqaoxLtkhV60rGBSjU
x/QC1mrdubqRsJgDGiGZyKObTg6qHo44kMcU+s7ZQVUSHLw71km7+SJdBBre
7GF4sm0FqXzNjFnddx9IaclEvrmKpZqJeb3HfKurMcNmgLwrOzql+Wv39ztr
fXTFUQPG3fO0+DeCswqPwZjdapejJJKAUUPjYFRyPilQWi943a1xjH1ZpVfF
fytLLz+vSNtg3ijph94pOGSIwrAm1xHyf14X+g3PkNFtITti1bAkx+QcTIAE
NQX2HdjhjILy7UeYXB8o0Uj4N93fHwXDv81qsughiC1me5PxTmNwZX1gtjvX
nkflQqKmHbeWyaRSpFfon2ZA6/cDFpvPPtcBtCs5SZ5NgI2qmz4eDtAe/pWd
qTo+Ksf6Pztd8jADX/UVfJdOwiEt55f8ZtrSz95sI2u0PesxybvwiZqGrMsD
X75Em68NVUgjP33qXyrNHud7EYTbD7XufsSHbgt7qcOVHJUz9sjydiWOA6dd
4nCVt97SZH1Vj+zHfKmBxk5FDqvx/Oe+zAnT4rZRwWrU6CwpyC8DCnb6zixt
t4Fj2BP4QzY4WmigQaMQYTSxVzF2rQMpcAAMhj8rjPg/HwHCnoYhjsB2yRMR
TBWQe5BFBG+jphFaxyF1boje62lttxFFlBc/QRlqA40lIxWnwn9AS+Xrw/+R
+x/MypaFw1NZuJft0T6lkJIGhEX/whpjbEmc+YxyuF/hqDqC/S2C+XQ30zq4
dqDJI1kLZ3XLfz7jQFEgCHvzbcTXalKarkYBwiAugpPMbmXyX4Oiu6YMkERm
Q5IVX6HuqVhBtJOY1qXNmAUJlV6nmuMivRKB5Yx88TkOmxrVR9sR6tVUJMqS
0jCCBJ3+AroO3oN3D+pcXUo300/j8qWO5JidBMOcvluQZGk2JhTvDj2bqnLo
Ee8VwTkhDSLTz45W4KK4ffELsVObYX7FW/4y9OZaVQsc+Wi1LtFljyGMNGlS
P2K+cjg8j59AEx701uv31SgGn5Bs86AKXKpmt3bbnJPJ2AdHL1il2g5jYrii
RujiPzOO83+K0gmIOL5wC5xvlkT8tHGLTRZXnxRW4gcpHNJxXT5yeXdfQN/2
9U9/EDDFB3CYwR415k9BfIR0piZaPPJkM4lHkjVj4xhL5V+JXqOwvXWOj6E0
nrDmlfXLNLzz50YX3zovfkQyRHIJR0wAHg8zuIDV9e6fOG7WPkxZhUUIAOkQ
jZNu8UC4ZhpkwFg6g4Ku99WksDZKjAkO2UOxCu6jmxnlS292g98Cnsolp5ju
q1N2lcXWDJcja29EChy3+vKYVcse0nwAIhWgApvhwf77jLHbXH3Q1yWXWmBM
ZgZYj16cesAjcG+KM8Cd6vQTos8/GC6Tg2ik03Vp/ZM1H4nPZ8aT0Hqfj8aj
mv6UpyhxqiHD8Lwf/0gMsyTyC27uBs7/fO4NbEASBv4p7liJC+0QnPNG7QZJ
utuRbZ5S10VkC9Mqad7EiJTe1zNd5v65j5HmPyU77X2QPhxcqFl9amYYOkq4
zJ2kxnNYawvhuwnZ2UIpkDiUe2axpphgl3UJazeDxy1qjkXtMVRqFVOorw4W
CH3xR2wSEl+zWjAspTNJRxrM7O4QDGzl6oaaZ5l3qzqG6y8+zhnAUebQnwJZ
bug3xdIwAz8AY5Xrvgb3lRPK5kf5WdJsdEiaQ2ty3molPX3EXP1mv+F8Mn17
xpBl9CdxCzdvlbeg6WICmNjwcfoM9u4PfLLtT/zts2T3t8vsYqWkn3McHS60
8oJGpVGJ9rDE5d8Dh9B4cAyN7Z3dKRBZTuiegfEWDeMNX6WfWK+t2Ueg+BRn
N44HKzwIVMtISSAaXxNxZvi/FneqfiCNAFOtT/37deLUoq3CecQuJ+4vzzAH
MfXevXwdHH62jqu09dCJ4/kkr7JWOE1tPNh59FSqeXWJNIkVJ1Fe5r166p2g
TWuugUofExIjxP3RuQEMaz0jdPd2hxxdSfuFicfhMDQ4nCV+6+ZoBHyCzXQH
XhOnQ6EA2PO1r3QL3Bqn2XaDf7RzSmGAzxEIHx+8vi02xZOUoW0XxIXgszbA
V8Dlm10lI37FoyH4sP9eHFa1XWNMfVaiQfw7aWuN4X5XzUF+0vCJ5Zy8s9m5
CJ7vCHCnHYTgbUobe1XwgiiIbvzQ8A7OC5TbiUixqyQzeFObYHOBcRmPr2P5
piSaFNryD7p4tBY5NUSC5GQe9+8j2PfJ7p+uU7cIBiGI0FIAa6YZ1Zu0Dudq
rFSFg+yQKIL3DPsJzTxnALtqGMd7sU+I1I1pobYxwlmPraeGfqhp8aY/nNU8
ukqploB1R7mLjMC04CD9SqS0RlrAlJbNNQTIrgPPUrJjPc1yeN0YEUfLojwl
nmXmf//PD7rMnQ63LVnOwIo55yLewXLox2NAG5gCHgL82citKKQD4fREFdOk
rJm2ON5igxiPJHRCYX2tt18s1RzQp8WZdWCLbf/FTIja07B/mSMQbbPhIc/e
ZS7Gutgly+ErdU14i+BGoTekfl6HYwVzt0ouzv6+OOY73Hh3ppohdtAxwGYh
heLInl3JMwchpCVL9wVMLDp2JpVafp9kpGF3LqqoUDaAuk6QurNnSEHjh5J2
Ct3ODZi20y9QqUGFxXP9VWbnNEziMal/QDp+QT0xxwnXQzkawBOfSGHaeo99
LDit5q8TeWhVnFSqS/10OEnKGhlb5dvkrIvt5Jf40Xjbwv3ZE7IbVaAlS8l9
CgAFDg8dAEAJQ64Pxg3b/W1R4WBx7GsaR/A7uILUG4EfTi9LUKxKah24cwXK
royL99soqcpt4oKWVXB+lbZ9hKJIBcX4uAY6fac4bL9yoEp9cAQaRJ8r5PrH
DmQmbX2SBX0Ys+HKVCpSR9DMrXIbCNLjZn8XdM76vPjTwoOjBIrCSDiEhA+f
lKC8FWSulpXVuXUupzU+G5lgtRGcawqpyjMPXXNl5PVdAktbo61k+ZeCXUwp
CWcb/916f9BCJitiXa8KCoqLGj2Fs1NmGnmyh8k9DIj5iy8KSs7JqRrXTkKn
dJCkVJgaFP1NueR3Jro8v0EXmW0MfmVzn9wbjBkrP+d1GODyrCNxj0zSktUp
BxQ5MJjtl12Jm+kWJJL5B/4T6HHrmaQZ2MzrOUOr1qupk4YjmLTEaKaIoSVQ
dKJbFnlS1WoafaXgQXdsqjcJshk2V+Di6sUVxlYA3d6xfyMGf3lAzX3Ofbpi
P3g3DOOm3Zq8E0NHvL+HofI+hyIhIpQlbSLsSLNymYLE0cNtyZvwLijRZWhN
qhvnJ37CiTHQXiMSlZJdV/YZMZq8wuJFNMTiKlxKnK2GEs1YHimBmUd/xGUN
cpTX24PmfUyv+WdUWgwE63Jo6UmmAT1z0VbqTOLS+SS+y/lZO+f57MIojZYT
Dz/QgXTqjBzMuj9q9XeAUFJhgMNpEGIRsQfhXBm7QFGoG49dAJ32f38YASTH
Daeq8IP2PnfSxy3hTGU+Mhpe2jbINePDHblYIVmMSyzbqFc5Psb4ZOfrUW3R
P0j/pmn8doxY2PbdrL0EYwu+wM7PRvduHbJ9cNQPkcPrky5GSJe21j81UeN1
wE/I/nxiriA3qK3ZhuGaZ51VxDoVjfglFvO4A/nmGwJB0uDHtXJu1inaJ7s0
YRP3XG+b1Jigid2P437phprPpvwaGXWQlY/18ivb/FQl6JIFNXFivqhR6gvl
bJwAgGbexfRBxJODCe8TWA/gEgVg9C+2reNfU6lepB7ExeUeN/CwSIc5+NgV
jqi8+kw8J9BrfoFMHJAPq8gMW9eoH2Oq8ehKzsR+PiQTSzp233Yoik33sMNu
v16Zq5XLyi+JyIdx4OkrEP4uSPxdTeNqgdVmp80IMCinOdsP9HL0Cqj2qQY/
5y7szMVJalJw4t4fSRT6L13qBB6C8Q+c8VTEp1NLhj4HFAvCuNZy8vlOMrqn
U/pMZzBuS3u0jOEfENgi3aE6xBmgWztD53JVsyRIHYguR0dSaewqI+8SwTEp
zsCebBCofo1QanFnUK32jyei2m4k+ZhHFB7yBRaOX/pY1iR5bz2zmqM/7dKk
5eLVDt4jHGgErbAnKYRxay5wmikAuIw6zUPv8A3qAlw4VQFve1tJoXYPfTgW
GIWurgjWhplGxwre6QA2DmXHJRUlxhNHtzA49aqBwdGKVfA1CHObhqEtiTE8
RI8SweH4mCzKaRLhN26/0mvEPqatGyL7StnQ4mQPmLI92ec1nmPe8ZtJ4btS
jrfFXqKuikqXcfBYBN7bgcSg3CpuOL9HPADO7a3ZQZz1BVtopIKYuvr/YYnh
AMO12ryigVVNRUR8nAtrRs+KfXGvtXarlh2pfDj3KQ3fOdaOsxEab1qVf8XQ
khcQNpEroWSpeNUC+uUDY8FrWobI/8wwYlc2tf+rp0Jr4s1ujd9eyBq9RxeR
4G4DfG+KfuL/C17zjZEjv3qn4LE8IXUOupwXXJHq5SMA5B0Bu8LYza1w1Z54
qo2h/qWi293/Cu8sBa1VqZQjaDLe3RhxQBtytiJi/WS3dhTFqAInG60+qq9T
xGbbrqO1gx2mVYnPcpvlj7Txv1BqFgZYCzPTYWpUHZn9kpqD+1nhtU5uFaea
L8kUlE2hphndnhDg7SwQn+YOT4lL4AVJE6YuOnlk0P0lcSrN3N1KrGBp2+5B
ahBInwZvKwGNxRim4WixXUTeTPpsMYjJYjFbEWiIRrLkA/7gpwXhnh8oydmt
i0O85RGPx6CYjqnfm5pmLQieQ4m97qvr+MIyqwp5Dqprbasoksl+WFZfWY6H
Qp0rpOxNocDe6bVUi7XudLz9sel159c9YCU15aVmXxsKothg6WsSNHyONsdk
9iixOBwWcikW4QZyRJI/FQVYOlriZ4q1x3efvPkpNdUnoQ48HyQXwQI21EUR
KxeUepFkFcMXNUlcobH/ATT4BzSPrIAEJjxLhvzBO/FGOGY1ErqrfcdhhgrA
4/lDH/PX8PiXv+AHSKrY5PSLTdhO6UoOa7dCuzNzr2zGqsdPv8MPA1vUd8tj
XGK+bVqgjlsvcGtc6PiLAFdtHRMSPkhyUT70Xqk7vwl8nMHpahbiWp8sLxKz
1Om2hJ0IJBXD/tHo8kVBfo/Rr587dgic5Dcy4Baxumi8E1J/X809NbNqfvk+
EcI9ccYuKeqff773GDCdBOWEBjFQ7RnKp7hIbIjXaix2MZ4SWDfumA0OlIT1
zyTq

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Kttctzi5aPKQ6vg9w+1g45z6Da0UaxXtt50QPmQzmLiVao+5Qg/yS2eSRK3c1uFoxS+G6ngDcAKHm0LGGibx4soakCOjaaRTqJmqblCXBo4qigRRJU5sOpNJWGKfxZC9LZLfFjqN04HCQ8ah5FN3P2yNU1iObRgi2dEkx758LbIsGmsSUmn36d6MTHQGWCnH/AC+2pgOY84Iul0q5eg7DNO6RSxNOih+2JmnF8szbMMeXCk2VKOWrsKBoK3CLL8vk+BAh0gIC3ED2B4aRACyIESnFAtizv6iOBJn9sTwiD6GaXHMQP8cbJZpIPEHxLZsKJmBypF4ki7rR3HxrFYOhS9pwuH56zVDNwPYc9XCVjCiM7FQHkzvdvmIPsmMIdex+YsPlvxNKyR+OH1+o70CakizyCnyItQm7JUOkFpZiBVZ+5MLJMV1gBZzVzzUlZ1nqoFP8WcSCiCdxnhf6lUJ25G3L4EiOKmU5Ztd0K2qjnr7ztHgiPq6UmWHSSINbgp0ATpgRqyLJQ2MkJhBwh8UEXAGiDHwmojanVvHh06wmwsgBw5jHYS9PO/YjUISi+ITecRWVrJAnJAgO8NYQ0OXHU/9i1aXFJ0OkdaOnTEPHE8HIOIuhAIQez5MDPUDmUKQNIg+QX2TCMcTfs0J2ouFziQQH5XriQNtxyWlJoWSeIOU58Ziw/nbZdBMaAcBU8BL+mX7hu6JMZoR6pf9anAJlsolP/awbYixY/Jm/EZIz3Mo0u9eaM/w3v/p54YFY244LmQjBMvSYkUqj3scwXezzs6R8NJuDk51m4oONwqUv+0epj2hYeSIpegWK2IFDk8oz8R3GZ8RP2rW9N5SOsZLBaDgPoo5rckfZiLIvuixQjDEFj8n+53T0kq1X0Dpqsi1KdZDX5vqge5fDm7DUuHNojiVJVzuyo2Odb7ieJly8z8h9a1vJ1dlvp3Ukt3vQw37LKEI4cLgtiofq2GvIbqKuw2M5afkfPxNVWPdtyX+ItnS+nKGjLLc2FVrO3EtOtZX"
`endif