// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HKvGXionms9JtPJQWxG57X9U7oXkz/4j0p+HlD1o9OyRQ64QKa8/DswkJUKs
MlTkJ2ToVe1WhVr7WawFrgs8rOWIY2SlY5E16A49N6cvQQOGFyD9cnz+1i6t
GruBQ9xq/qTKhzb49qIFA7kNhw62VpXhWe6vGJw9GBCWyBRvGrhC1cKvlUn+
8KVJ219QeWjhN3yBHVVx2eHqz/gqE6K0jvWikEzgYb0gmHvae4dNnBHwn+GH
rksPhjfqSMfYkQOufbHbZRjcuBPTsxR/l/RcF9RX44GzldZ+kGi4k7HFvcZz
YdLUQDe+PzWS1tdes+JrThIZk+ZO0cPfa6QRIBg9DA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YQP/D6a+jeESjS/4vDcso9LkrKGmlcwrmhaPldMGJzkF3kBGKntnO3iDDmes
H7b6ZKViNFs3+SuFZmiSqx71CWCaY5kozXOmuc7Njl4w+WTHV9p8Y8B9ygtk
lv5p98TOcRNil5eewdPT9mn+Cs3eO2LcXkz6Q638dbjZqll2qhauvQDQ0EQg
VXCUHnBcGQxQ9A6S15WvCQ2cC2csRxow1ZQRJMdY7MRoxvog0+iFR784fBqS
u0UM+IXrpKO+D/tMh6jgfC1fsS6ji7u97PXeidEkKiJr/BKoxh0FfZhmTYAE
5vcuAGCaFqngbzxzK6VcZGqP0eftUVzrwOhA7uuprQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
r/rFpz9Gfq4TvUmPvfmCqJhqyxfswv1razKQZlOSuhQR0nhaFPth2qAc8W65
c5m96PsN0PbQdRF2s1dquCSXstHwYqo9zE97/3lOZValeO9gCs29/bUh1P1j
xoO+iVU4OCjZWJrE8V7cRz+Ezat1AhLyrTfe3ALUUIoytNyu8qYFX5NN8Tju
vIoHiSynnjZ3+p1wOKxTbWGutn5s7JnUjFVKSWN7WY9mRA/+gKgHMX4rWRrb
pq0E7Df70AjirX1grsmfsWBfF4qjzI3KeJ+JeD/oEDwxYXdk12NR1ZyOO8iU
VoKHd3CDJnqQZ3IVwhVmEsFvv5oIMWMqgULhDjgfog==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WX8PYpPWZoPgCwqlw+6oain2OLC+U/1b8XyN1keNJU4ly9ciS5QBYa+Qgkpp
ssvxR4dbzgSGJCk4f7hO7x12NH+JP4vvSSh/eAtEZoQybqkmma27emoWmw5O
1L4OHXNeQkhRReY5kOEQkhn15HIs76ZQOvV+wGlF2wjQmxzdqmk8ipOEAqOD
P4g1Y45RFeTT5GAD0p3JNLECAlmJSZXTBG9Fw0AHT4IqMU9iGlH0IaoT4O0S
fI5POGVIlMR0ImHBh9iVX28fn91Q+ORR69kwDvhg9u506f420vINrOGTrXkP
jv1+xKuBTwQLRjm9NTm1x0TPOQhJe4jcBlTnJWixiw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MYVoJAxp6vh45JVIyTo70A+pOZe4Lk3OXHgU/jO2ge+XDjjRC197uJSjE2nf
dXSzkXHP77hJ3UPBFj15qMfd+0bEBpTLnU5QmL9UBzEh5E2Wzu97hufbmA7d
prkLeYPpG66zO86SbVh5wgJf9pKq8N/T43atlmWxnwpb4U0Ufkg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ouzUiE3vfZM1fCWhwLoRxKayrvk5+nwcsRESsrLLi/wjFc3Ca+31TJkw2zbc
ftceTa+WDbpRYqAi3hKjh33J7aESF9LwBOGXDOlYwQTlDlfc75MLxlIYsEMB
HxDbZKVugxVzToTM2EvsEenvCSBQ6SWLBG/qkFmFJuc+X/rBfPCmJNYHdUlk
xxIWFn7j2BLo82dojTkIVzrWQAqd3m2JZSzywSPrQZNcqR9zLu6j/aylmu1L
hoaHMJq8Ah2pneQZ6kPFdWBIFBYTRqhiJLHCH+rmIkoqEWoUu279NbCqaz4y
BhYiMGqL+6TbLJqUTBj8Zyl2FujWBBDW+DhxmdQ+fKGw5jhvf6TqNl2DJpMG
qv288+mj802eXelrWqOZigbP3KEJARKO9+snUDB874uJH0P0fvpO4D+BGfJ2
qQi/hKjvOgT7LFA73hylRmPEi0cde+P38L/rQTz2QEnUlZyYDB7zISRb8Q/N
iAG/kVJZ6kav2QKz76UU0uX646BYALyw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h7SlK2dkfqafNmI9aw7SppTR9Ir3zJZjEnttA1UTJb+CikV0FKsqRkUD/9WL
njFsBtr7RLCksWqr1QIVFPRkUpnyAU7YR/0J3j04MIONjU3MP74BrgrBRoyg
Sp7pPiwpIRq9u3fs9tIzX8Abwfrd+eQedySkXb4NN+O6d3SMJCI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A7J50SD+24yx8sPhNflvbg7AANHBfkmeoltrRW+EBFJpjElK14fnOyZYCkrK
qGG4XXVHsUQpvm9/eXHDjv7lc4LgzZzqFoHbLyq3Kz51zSL1nywTrC3gDjb3
Sn76Bpnqh988GgN3m9Rpft9VEKkJdhPBTWdwiugdnccWJ9Q72ZA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 99952)
`pragma protect data_block
ExZPRGi5gFTOR3GIgoNtizH4WKH+YagZwVSp7voxoNz0znFT1W6uBHIL2pp9
8BlxAJ/SM5EEUiA6yZeD6Ka0ut9l7U/5bhgvu/vqsvGXkSJK/3Aj1FB59lai
xuWcMRi/D/x0I4gvt2PgRldi687EKf4FRxoozjTYkosupQtqerOSupBddiM3
KdMk2IUmV27ft0CEJP08JN+shKX9rzQsSQmakx23fan13f7sM1nNIa+n9NQg
H9HC672W97yJwEdzjbOnk4PC0GGfZ2jUSgCPS57x/Nyqm/9OcTZliCmzVt4w
Rvs9jUbRWDl43HQzZUTSR8+ipQfMzZeX5lmqT1FRmqCFlR4YVxncjazQWo1t
OoYmMS+V7Z9GdsX12xgcO1XnenAVzf84QCWapPNHDQGGunbIrAPYGjtD20o6
6ij8JlQ5Mac4qqnDfvYrBO6aZtGQNOS6imtExTc7zE7MBrFcCGJcd02a+oB1
scyLV4u1eEispPdY0E1N/z2XFryZk3X2WWqVE5cXrl+ZfOyaNptxaxfJJUHH
OISWzHui8ciYHC3gki0oUFlr5GJ4rS6jCAIPgAq2MjnX6q1AuN+3msEs840X
bWsK6cWZ9aT3AjwdBis1ric5fzCE8xJmD1gSo8DM7j4chPPqPbrfVZGkzk0J
a/911VFOXx4SK9rLYH/jdkCDNyoHzzfEmZt+thzBYSzl6p5gqNw3TEMxtDEI
SxKjScAUSRtmVm8smeP5wnVnHaqccuYUmV8NniOE9O9bTgjS/dpbPP4W4mtu
hn+tTjCkk1XEIM1bGlO+RLDy8Rmbk1o8Y8eZvsxt9jH9Z6MR3RJrH18FwWAy
hxMLYnjAez4FUsR44hXztemhy4p9b1FH/77YgqCREpDt61MxRaNgQfKg9Fvv
HugXhS3iY+1RD2df5ZzyY1wdlhqcKE2eqi0RF2MT4mMvC2sXtYQ7C3UyoqGV
LPd/6O0qb0TWRuDP5/f6qFhy8lQZImPkIummPT+s2o+/4zGOiXNLxARFNbvl
y04A54K0EBahvaeEc7/IpDunGS9taMDXMSuEtXMDR4t1FiZBz/8FhYNTAfYc
CJNYzrGcrF0VbY1uNjXFqi6QILaJzZeJwbzyFfsIeUse3dqZcot2eIASEa+h
WPqYCkaMLR5LPUfjHTPCKKhsYwAIkwealCvs71x4rAeI1PZks+FU1wkqxX5/
xy7NzGbwhFa/y5Lt10eU96oEhi5WCRXa1N0Hnm8NMbi1W0t6tg4rWAqEsHOH
EqDMS3tVdhlYAntgptDo1bvvuBJJbOCtWfswywZfs/mT2sR+tMdOKs91dJ7T
pax29O6rP43p4BERbTBgXMw/Lh+sjLJoqNd2WaAJxDrxUN5xDnFuVxZYzdTz
00R5axz/yIeGvQ6LNlD917LabUtiazBAiY6oDx7ix4Iae9HUFBu2Xev7Dd0l
gK/0gRhkFcBw1oy/Nc7KNhpeJR2aOQT+oZ275JPWDfIKVCuGsJZHrWC8FoAd
PusQQb6gtZzyeEvDNE/Pn8RrdgsoQLEm/7PZZ7z+WKqUjh/+qrGIvqR2Y7Ru
mgEdMaXkRjRVFjEjbI8E0h/1mEjmhxbXGro4nn6HzRvofSuxQ3pNBr0aoYRD
3sqGrOiiHI5sP3jFWM0GlXCY9wv7jB759IWQ1t5SWjscx6qXMhdnDpPvkTkw
sg/aV2X7WGTIZjCli2+WqIJQi2cfbpFrnWhT2K/p32OyZ0C5oj+diBNuC3pG
ZWyMmY0e0t3Voa+bX+rWOl609lN7akuYx/jPh0OlQKqLhh4qy72jPG4m0FcN
KXUdxYak0a+02h9DtdPDVYQmxg3apntqyxzrCwAyXf7mjqAH81VqbZYjokqv
7V5DGCepGqKK8OXknafw1+NmMl3ByOF1PVDUvisb7Czc+0c/pfbLszTlTUqs
qZ7KUgqj4LD2w6kqlGyKgFmm8uOqCJNQhyBwOX694nVR2bR2ZpbruZ4DZ8Cj
72VaNDau5aWLKXeFJUFBrZir/zp1mD6vqsfG278z1CpxSk70NLG3Jhl+iJNf
2RO9HjyLUGhtHpDYlosrVVGdp5ZoTZ+Q37KZmcDqm4lmW/pv257jooaLQffZ
YppTBzHUqN7diKk3YR6TTkri/h10l9KxT4nTo7LdXR0V+n6LpWvy1LWEN1bm
4IKxqIbMhLnsUVMh+IdxqYHsbl8RfX+hvGup4QY/Ogj6/m/tN0Y4uleWnLNh
4jCgs/bQg8q37FSm4NICyN1hlDBlGMlOnsiN/w4ESSe7ED9lj4tkYsnnD20Z
RkTi1Q8pfgw45ubJM+hfbNW2uSHLpVcLDJIGiDbrQdycpLP5HejrWJmaTgFm
3flZgvqEW8uTlfybLlKQ+0ksLBCE4cPz1s6gAzujvI2t8QyATYeQxu/2+mqB
Y+ExpPNfd/EbaAzXuMBM0w8QJweoJw7tW11EnkgVr7YPTD3FSvJUx8FkXFEE
dPp4P1oXFAsmdZjItgiQ85v4H+iXgxJvOABWa1vvzILdu2HKrocLUlZ/9wtM
+lR+fq1McUeAA9KufQcoub9cftZzR6+kG4IoObmDY3KmtZJ+iC0A++yfdUAb
fZKVpMxbJhLU0Jc9A9n/t5Omvib380LA3/lF3La1gluZBJ34JtoNA+oHmk2B
cxWJJRIYE4ETmtIf6gJCvkQHoQL7k96CxKNZsvB0AMU1AxcqnvMLu90B/6qw
ISmB+6o5ygENV3iCqfDViQckgR8LF8Pb1J5ak/h+WkH1HTEkr7FffPJfgS1E
hFrxUakWd7lAEtMFrzxKJ1E84IbDeCXBEI2DP9HleHO0BT64jh+0CG2PCnwR
7JC7oohcB4ExKWTTDTMyjUA8L6t4OT6QvrQ9mkwdy/sTr8rtuoqUbUfkHXoM
BY/i5UjV5FviMeDpDAS9jqSkEaz79Z94oo7RzSIuPsoOIDRDBPBYdB8JbcBZ
OfbA/gb4qDP8Cl7EN6GMMH/G+0YUJ0vHKOLl29sxD3nl60fODhhVINPsPuXY
ZXGC6+Z9fszf2aVHW4AneOu6KaTyUA0tKbp37VTVXWI7mKtl4i/UD/kKXjRR
t4pplmJftukVkFnvWmW5Rnh7bRzR2wQAD2EmzorWASi3581D4xgYf8SZ9eXz
VpZvdoGOmrS0WqwVM3PB0I0E4PKDrjKv1fCMB9JaxLhIQohpWkRipeFyWV4u
P5+KRFNBRBTc4Vh/5IsoBPgUiVDpJaN0ZhKH2vui/MujTKIVNesTiAXvG9D9
gxt3cZQ8/+y6ZGVqne+nK9MVbt3jL/G2eNMZ4gC8FKAbdGEGjB2YmqV8KSgi
j1VKSa40ZSHEfnjhob7vB4q221HyU6xJ97TXIVB681h87k1g06yDMRwLWlPs
GDtW1gZFsHd1q5A2NywzzUCSp8OQhcjDNjqhs57234h302ywt8wTBpehIvY8
Q87nMsogNeII4r+kQZmdaFG1r+nL9htqj/cWM/gcWtXkrLf0twckLYsTU8qa
CFOumwO53jiscGdlJi+WPPVOIeZcQcMHPyvPuk3Ha3JlY7GTO5m2hP2TZykq
d2VcoIHJlN8e4La42tDop+KuRKy2CuAvDnpaLovtmCTR+TTI/6ild4LDbv5t
rwILIK0gwQMRgxAg5RiICZzXbY1hCgWWzbLTyHl0S0PW7dTDFPKYG48m1MSY
n2emCadQ27/lYAlCM39+XkJWzTA9y4ouhXJ67VZNTJgtlimAKQfexwQZWcjE
I/WFgCHevj0U31i0OngowNFzE95nI+/dhWmvBag8Z6A0yDRE0+/6kU01a/rY
yA+znup8ptlSiPRPnesw2W0HwBsZNuYcRHghPfj49QVXIgxW14bwAxIH65gf
XP9Df3MTViaqUGIBxnuCYruuzEtQjfC8vFx2F0BAXZlo7ZbEgs2tA2axvTpT
vDYItm19/8Qzk46y0e+RLzXaWWqlIV/1g/zydRPmXcIA2mjWeq2FvhrA+vV/
nTq6P8naLzN44VXjU6w1Mbw0wkAZZTLRuImQtP71di3b6FINeYxdLiHkXXaB
68y9JeuaY4y1PEjzgVzTsA8NULZ+LHHqwlMTUKr5Iu8291BD0kFSN98s20wR
XjN+lsWR4rvDeJH4ZgSP44NwUOaF3ptUUhOTfSfhLZvNCrdnssw3IAJVltP6
xxhOLg5eNPfCP25lus1BM5Z4WF6UBZz0nkiANSim4RIusXwC0K2n0VF9LS0W
E/vCn3axAG6PahsADVKxjHXAHUTOBkjcptKrjz0rModW/rO4hHqp869Iv7Cd
viP0Ix0nEVWgWEDy2pSayKMS8uyZDriqYKz8qjHlB0zYdKGCy6qmaC517n86
iEkl2F+edtt7YV7YgHd4pDb1Syr1M1laHyBI/D/PZPvuMK6+9R0eVewicJlV
CQskMSILRLRtpUnzhwLXgsYwOkrlxzqm7I2hJI2TM691Af+4usapBIiwwvH/
Yu0mg8Uy0qJ7SFHV6sHgdwyQSXFbDSnjfnLR/K4YPqLU4O5O/KSrlkegPGkh
agy4Zfd1IfFYaqe7u8IOGQvyYek8RDm8mblGsjojc6101h+XBeHe43RDhH96
GXwxPPQPPYrY5ckcT/h4TWzeArumoHqizF8TD6VHlA5grs6GH1h6U5DYgbn/
lVxu6z0zVO11sK/3UtfOeyKvyoZjzFBkA7XE72A/2q217F7TV8edQDaBP2H6
haVGjCm3Jr72nVc7I7ELWh4PYC6ZHz3vw2Kx7H3sw8cvQl8hExTit88/fIX8
PSZK51g7BQjS7HOIEuu2uEa0BP0wwwULFa8yV6yIwV7UwD2RHdHlVDJVCa0A
AC1IXJhKE+iywz8EOUq0uuFOpPxHrkZSwfuOU3WpdTQJPeRKpq9h2bD3y1RF
R1Opxk7rK61PY3MoxVltxIcBm5MOHBN6BBvaX5DREQeRItsB2HX8XHFqpJZi
Nv8Pkw+Qw4Q4KDgvatMLUQMGIvjuL0H2nR54WKNQ62cwlQoXouRAMeKoF+Ef
GdnGR0P7HlWpnBbBiruJA9yMOX5nRiJBDPiVVmw4kQxaMBjY745xxrLUKsna
2kNgTCuyJ4CErJRHDcJOEFEQPQVSCn8YotNk8ZQqumkHrp+Ru56p47SKNaIM
KGMvOgBXkWw8rZB1yuLwpO7F+j7rbvSLJdOJtYGVf5rtlnjAmXqGWgp+bACn
RALS3C3RfsT6iDT0ON8IWbCNZ/+qEA2bFNVpwicAhDkZWGLd8XFfgXari54x
WaLd1A/viZtKltwRcIVXgOCsFUhJHSXb1l5cYAjo09D8wWphi8wGbFcgYNaz
eHMki00z4k1duisJ9XdScuKyB66LeIfzwdLD92lXlA4cTkGTHWItaLgeO89f
wavdJ3m6lJ5O8GsdbcQ5tTjOHxdoA4K/d5NQUORaDhqgifQa5TuiRjLE6dg9
3U18LzxuBepc9KX2Be/EpH2FtOSkT+KKN/sndgpyNRIvoi1xWAJCcSuqJ3Wh
oLRG6Q8x2nQTdEHf+vq9hux2XK5K+UsUoRlyublqpj0jqqdYQgXq+VqSgxm4
uwojU3Mj25Sfyx7StnYkPDwsu9H53yQyiZBGBPBBghZMOZNiiAaDYkcfdjI4
V6ytICv1rU6LiUAs09B+ZThM4u14pHCgcd+yruHM5RwRz9JAUcpadSqDfAVX
v0WEbp1qXTZ6/KtPVDoH98N1ayVJjGzAHlzxZH7hnEjkLm610jaTIGXMiSPm
dkRWvvEr3mTtcfSSnqtj0RsB/TDE4AY891vU2j1hrF7RB+iz0j8EUObEt4cl
x5xMuG3TcBLzc+MhXQ/ihE1WdbSMGuqJOeccuTV/TEhUUMVuAJOe8aCVA1JF
aGXTqYXptMH0j/gze5QAKdgO1DFP/I5GhuJ8uTTRDPlwUfVwUwaYr4rBFM91
A6h1nf8557XHhNMbQM9WwjBADSRD7bPxJhVyMg6fmTQPFxkmouR5bVYtj7cg
c+DNGTMS3L35wnjABrwiNAsEEi73zvUYLTWaVj4ebJEcqTqaVkq+yzop6yCL
gtdeH/Kq9zdlmmn7j9gu+0FTWA+AzID2NX/zs4d6T0Og/um+239tbgMkAep/
dZIEghHcjpodngDzYj+dRSv//nqgjxmf+uKYKIRUM7wVmGb07wHOmmM7NdwG
h5wuUTl5dyauU92rIeuhlv7iqzeuudXb9SXXIZ6XxWHC0Z4exHnkTRmoEon/
B7lJedJm4axEL0cZaQ+o0scC3aLy+K8E4PXCcEXoGvcUK2YZ5zlYvQUVdYgr
2i0X5RW/jUGylTjtEypzXSr2J3JZWgcNobkGuFw+7nF7tilOJh/ShIpW0+Tb
0kH+xAxmyB4Z5auOvNPpwwxegrQllGhx2Ku62r0hrBCzakQFA7gBDFPCXh46
WDNOCkki8By3KLuLjaDdItP9KhsZFmNkuLXMpUJTh06ahFbS5hOwA37KVCeg
4oSGa9l5MODp7zzbzrZQ2hmTukybAaT3kKnGhZVm3H0QzpTbOOR1DxSMOvWP
xve4XKlxqKOWjEZjJb0LjsYAaQOTajdvo/k/ZeUgDbmUTh9R8O+nRsPV98n2
+dUNQXI0Luo/IjrCIwSlmupJR1S35lzZfNywES4oAsyUcrBMJW1gurRO157Q
WVxZCFfhqPiiC4g8Q1HKlirzkPHH8pSEEvJCygcAekdP9EFsFeLxO6Bnf7Tc
v9/YFDQurRdkUVHS+2H6zynJrG10fR3cPMNYCAHeiYnDzh4siIULue/XtKUK
nWmwU7DC6ddWUrYYN44hop2M0ND33vN8CS+tUMwIRcbnYLSlZuK8rZwIiFoa
MTAwFPHCUf4JpmnU1JYPJF+AfnZjY4yokvCQIKXNQ+hyqvGchD22N3A1Fmww
gDNcMOxgeoU+yGdE0kcXDVDoKbjYRLtR5h3B1OcBL7I7849p83KCX3ZKJ3Up
db4XtDtqzRaHbczrR2ehHrUZlOxFjSiSjXriAHWV5rY++BHRKuymyijjr19W
fUTwj82fJBvTvH8dBZD+YWqOwck586KoqhNwjAMUAyCPGFTCKfNwTou7CIg/
1FLKwiAW+fweLVGqP+CCP1SNr36LadYTw63BpBOoJ/1r2aVvxvgE3a3SXz1K
FsRU0waoC/blD3/jFPkdF84uMLLON7/BzOhDRzqa5nLt1pJplNvnT1UzYpwZ
hPPecJiI4BzNtif5umQKv23MpZf3jptQgchop96KwRL2n1tEtLcPbH7kVdo0
nxs1HTgm9LP4frnAw4u6RaRSi4QoII5GgeflaUcJV1u4dP0NhKWd2h0OI+oB
+xnFPq8on2+YJ/een8rqjaB4PUDwDgPpQy1fSUodBKDnrJNqAxMRpB1db/Sg
5JuUrJnojyQuamUtvYaUllX/IKu83KjvRpNwLBf6CGuSyceGbPOTGKQOKcVw
ycy4BP33TgASCb1N09by+R7pbIMrEPHeNA2pBEiJ2u79tfuwfrnAQ1QQnMUr
/d2Iuo5J9pgAhLLlMADN3dAuQTHbW1dA8QxRZUsDKv27nEubL3E0KP5fBgGe
9hob280ro5YQ3fW4kjt/R0hYCKx5xixGdqvpbzLkotBG12CRuKZQWyIGF1w7
DH16AGRw5YHBYtKVBJQ3qNr3js5DxFoaO1ygCU3CwRfgxEycjyPpMLckqqHp
e7IA4+MYzIgOMGe0gFj3x62RA4OAYkV7FokofEb+S8va/z+7j23evVFuJU4P
S7SBF2rCIU5GQBFdm4PpVT71Mp4B3CEtGB+DndwbqV6lmLKUvS0lwn5SjX8z
Z+YazbOMC9S3qH+V7nk4dJd5EVR+IoYojFOZr/vvS9x9cQ4fU9zR7a786qca
adwKWUsjosFtPhsz/Rb8nTTsY92W525Egc0EOnhjXEUeQ91bTfD8GJwrKVYc
978lb8UqwoYZcLicjgOQsBD8brponKmF5fyGWKFw5ZYh1gDfptZ3PIQ7vPuF
Xtc4b6yLcyppakIPWC+1JD2pMs9vLiREtwproTYYRP4a3FJkC+clowKtgcJc
YiyTsMxLCw+YcpqNwLVmHxQq8z+rzVlZLh74CvnWxLGNUAX3vkeyWhpd0Uyd
Ys9uNkV7MWxWpxrBOw9trwGOozxIKHPyEIDK74H0rnUM/PBZue/Tivrer2Ln
Mmq/EYBRM8qURflnK6YP8nCiDs4HUv+FISmYWsqhVlxhgTYzdm4JH9R9vdoX
cRTsO9chkONZO3CCoKVmaKe31VGj+C2yNXT2eTXPsfHPIriyLMrK7muEBRue
o/fGhSpX2t3z+wlJNqYxf4iSsF3lootbFOKQSFluPfJZQp4dxe07Us8zYeRk
PFMM272XJGNo39rJk3zS7C/z0NjuBAJJIQLfExHf1ZjaXzFPYbYZwH44F/x8
rdiVJPYy9AadamgfRF38WOrVpssd5us3Rp34btr44AA7Wgn0cMfo9ehUWJAY
vTLJRRsgoWjByLgkwykpf7FaRNSwfjuHlVnz9Dqk8JvGg+PU3PiCr70MoBpp
ndUK4KNJtin7e8ipVm9thlewRdI0sms1QogFQp0MiOFaz1ds1Q8kJDAJRvpd
MefkMW30SlBSZe//SMXuD8GxmpY0TA+kIujVYxIhFJgpg3GFEdpvFiOKxhMo
KOY1blKGmbVBAFDsTHhL/an0Vyf+GB1Tu8sA10UK+JWON0HNiroMwR4GURdF
bJVn4Tehphm6XfxlNd+sfO436UG1kft9E763HmgMppKo8DrTRWlTDlkCjTVk
Z1yOP49gHWBPmO9NwVDifHCGhuyEMb3doTcR2AH6S3D03DB8sSvNaoLghy1Z
C3r022gPnTZh49dLPQMxiWmFQQWhuYEnRlTmUjkHdQpduB1Y61PIaoSPwkw0
ID/DrDKakuftjLwXpNx9d7vvgJl3ff0TeOp2hMTKhz0QoAIGrhk/GimcR0le
brWXugur0eeDJv2HNB3LcB8CrAtLaL4AiwXficHxFNKZ/2ZgX4y+LDZVSuoA
zVqicVykQto3jgFlf6Vu5rC56XMsy6d9hj4OJ2RZf8fxLegR6o0p6BKTJ+Nf
FXpO4+osdf7nRXey52nROYRblTkh0nu8mqbSTKs9TGxZ3UfR3dLyy65WqBem
x0ZcEVhfs6BzpY3bGbaR518gV3nKb8Yc0HS2uUgvdOCP9DmgL4N9Gobsefg4
0hHtk0h7puO0CqZLUhGbclvfRtnF2w8eL4c1HBXJaLaPWckU4htDwjqd3Aen
M/oDn/bHdAf5KVOgzxRx2jw0M3tSysjla0OpuDwijNjecq0DdgIlq8KSW4Go
BvavoJs22nmOWcyipDMaWIYwY8garuCmgauYAJOqEQm8IUoNiKyuFVOVo9+s
vQTtLASA7Oj3xxm90+J7nG08QxhmjZVoit9nntl9+dU9tTeV6kThHbch+jnu
X3vTjeF6ZU0IWXv41T5FhBbkJXLF2MK2lkZZypZKyyP5mXCBJvIa4YkLYfyz
1Md9UAETmhVTzD//yHVNXSZp/y7n/1V3J2Z/brEYMdsEyuAzRE5ZsaSkAzid
D9xuJygBj9rD7YweaVOyJRu5ke/8a7WpdjK/7nIDsFUY6lKjXNN5sIRC6Jkr
9ryBNuTOCsMMLM2mexnEl8VjZN0aUi/HQufZhOG0sCQ+bxumaPdQptoSElis
A1VMeyeVG9KDi5pGC1wJKON0dNj8tWePiMbws39eMOMrEzYUZQkSGnVb2+My
XsBPmhbbLaNBiQhi+/hutsDdCh+dtMJZCLGTM8J3QIeNMeCeTAYrxJRAWqxU
9j1aid+e/XPs7+qNfBu4LdruM30+Gi+69vKNJPvqsh5lO5MEuKhIkcE4pHKh
Mq2O8gV9SKn7T1IkxNDc/0ZCG2TbzZzJnkeIFuSYGzNoBeVzJcXrJFZjlDo4
Go1dj+/XdjwOj/s5BBkMtUuMmbEXb4qMBT7VjrwN+2uHAnsq+9VA6+i963se
x5IxCqiG5P1Xngw3VfoUUmKbThApXsOtbSc3XBOYt2zYzHYjWkoyzdFRXuyp
Yqz2yvzaQmAIlt3sDN/GihMTaqkHEKp0XP0hAjqvxJN/iauLybjExAnfw9U1
QpwdemGttJGsifAKMuFy6C/tQ+8nmzHg+EAOiEnCSNg3pfEFA5aJoc191aAI
1FeD1BHvT6YYPO1WToS6cdk2DMSJbzeSJzU/Qgvzn/VhqOmPmXgiHTSSmdzt
li70wW/FT2tCQB3MLBglaPZO8WcLZNlbTPJeklHL2q5kH/Q8YefDXGS7qnAR
TStp8hNHXwg3uFRvuykU1iIwgjShA5DakyX+9Fd1QxD49HLtIYLaHfBO47Sb
QmOPpnNW/mw3+WLKT+Q5tSQduhJT57Pk+B9qvB5NtN73kJxV+UmHbXP9w/TJ
pwbQTQCPVGJqGFJG5OdEyjmQTEwrgPx9h+d40/z9IUjTsVWCKriU72tCC1WZ
UtKruWCpxWwfqHbQZC8MUy5V7cvWqIoaRXYatsq1gMUvaHIG7gHYi1Rh7EzY
2RsyjTFztECsS4eMPuS+os7Tv6krl6w/CvD1rFptAuGALK941/M1HjL8lnri
gFfy0b+PGnhM+AMAa8yorwvRYOEjCVA5BA6bgB8L1XdQo1ASw9X/ADd1+1Vy
dp0OkRADI4Y4FnihE0Wc63ZxFB8FnLllBYznOIXUjy/i6kkZ6A/FU6glS61b
BtWFpw4ZQlFmpxUT8pfd6EU84wBqj8dUmwbcqJOiHf2DCQlSG4W2DS0Y9lAb
JGrNPBot7V6nK1/7RrF0mWoLogWv+IQH9jVlP0c6+OPxL3a4Ro2NKpWPNglR
3iiKvqV3eB0m5PDGYxdVb5osOXcInjXwA1rJyTovjiBnnVbmWDtjJiGc9srA
/esC8PMcg2J5KJcOPTFZc8WAQbmkhF9bMveNydHi9IYNUQyOnSXXluPAFPqG
6FmUx2Az9C+lPgdpDHSQDbzO015tfU/FrNAQUx1z/hy3PfUmhL+nNR+2QXEL
7CvOvFT58lgvnMPGnZOUB98uTpss+XrSdmo9nB1YYoe/W+/Y8umSAeMe0zX2
z4q1hahi0xqEBGTOLbFwPIEZ7v+BUzIh6oIZNtC8LHcSGIJl3wq6Y5Zlysbp
I9hFYCMjVffmhUYsCvQbn+mV3Yoej/vUFKlOBIF9fcoRPAicgFoWOxQcJERW
Nq7Wb74XR+F8XQV0STQhh+jT7sEr/ogR1IbjwG0wHLf59eO2Ws8upl5GTSNp
RLR9MVgSK2Z7+kZUn1LxNhqdKMxKiVlGA10foZjGoXIJY/yM6Qb6mecF6MQQ
C85uNvEFCcZddEWDnvzThWKgdJgnKbxjfq9K2mcHHdPMbCc81YDa+CjW2azE
EH6tdNYSJXa82OaLLsQAAUrVR7GbVXBiHvv+mt6Nl/QDwIkuMEx98KhEBYml
nx/wWDCiyFMosgTQxEV+azzpbuh1aK7aPw3xXqgvcnhQ6pGhWiAqhOXcDP6N
UuaNNf/8BpQh0Q+HLrANN0Z8X8NieH/pIQhAcSlpmuyJgRuw2Eu5N1NSwf1Q
jnYy28ouhRg9+w8sGiYHKw98Mo1Q2KBYCSck+HGM8kW+ZqmW1RcqWq/vPfBs
KFiicGdpioaEhOEJsQ4jB22yy2DEstVz18U1LvnSWH82bVmr3ksWyugBpEXo
U6pmPQk5L9VPsudF/KhlMzMf/kw3uzWfg1zZGXWWKHuHg3EgzZFuZys5e5r5
WyWdLp4yW5R/iMPW7Gg5KgoKPjd5x/6z0gYbPRdamout7Ng2YyLmyXiTv2Pj
SvtvXAJAdpPnjRPEulvRiVeX+DcnF8eu0AYy0YVJnA2r/hNDXAysU7R6KzDY
VHgvEUKccYDuLCHegXuzb8tvnD0EwNZIq2wvecu9WQm7SF39+d6XPxv8ZQeb
IWdD5OvNp4gPYMSFbs5GxeYJDMFc1LIuH+w2SLbv3UB1wL8asfQsYLJMaQue
zewCvSS/rn6mSw25xwp8PTMf0icWUih0m7+TWy2OC2xglCICFNaM2PptFFTR
jQW5VTC6Fs9HM+DV6PBWjSOnTReVi2F+tzDgtwKS0wK8zr4qj4ob51l7YbQF
89HITPEYiE4oP8YUgyZhEIKEI38Iz4t1gEEBdqz3emafjzl+DTVZh716xr4k
mzlbrKs8GCLfgx7jw+hbG5M1ssZ1XSY4qM8cJankYKjP8OM3byR9y0Y6aX3g
tplsInFhoz/BIR7A7jLj3Ta63mscNAw/0TI7Euu7Qk3vKGj9jhG9zWYDBVg5
GgnnAmGYrqvnz8zR6bPirr2nGELHZ0mK9fTx/3xCj+y6/oAg+lJPH3oyFvu7
I3VpfGqqtRDmw6er79N7em1DJkjjyhMBZZItDZrIJ6ntJD+E6GdguEs4ECqX
NcRzpx/XoJ+lmYwTvbZvlxaPX1wK3KbnHuZUDQ2Vq1J5z0lAaO8QGNcCOPsQ
J+pXJDT8eN1xMhxL39BW/o3gSiRM/rewORiBYMe5lrRPyNicyVv7hqSb803g
QAJQt0xzLtij1TRuh7aFZusyrTKRfGRVDk1slJsbfnOzXWYfFGIeG5FvIeVo
8ISM15kwxCgBjrKC5alwDmq3U7R6P/Y7/glWBexQLE1frnaiX5gMARrmFL9V
CZeGUDE3nQPyrI9Q139ALhmzqjngikQ2AAEuJYPYQPGSX5U/0m/8YoWO5DkB
vrEugCnjXbAJbc/T0NPilpG4njEeP6vmYgF4lDrQGMCpuxoEE1ZUlMKMhGCP
CecUq+15r+sV0C/+lv/vKTTeQYuzcCkJfOJenrhMdWi0WDkZb+V9iHezRrOj
AQ1uF+TUF7cQ1WlMnkYjgqwwb5NyWNIa1v1lfIGNUnegHvr2MuQuexmUAFQv
VmZq2CxjTVdClG5ScK7eCchPPWvYfaUO5GAnVcboIpR9FByTa44SzJWws8v6
dY3H5f1u4Jk4srFAsNr00UZ5jog6AymQDY2TG2rM1dWBqkCHNztfqrTNFIEX
1W/jSFa9uxD8IvxQC2bPnBkfbIpsUxT/u9wJinNOIS9n8cpCCL75+0raV2g3
7hXFx7qez/r2iJwdjxM5SnjdqxSZCE77n1SrwRMaWA+o3b1o0emgceeJnakw
TBv2zddfCfoW4e5zBXiTdIuHbiUwcjsJxXAF1AQgDU5kAqkNTnNfo7Q7qJlV
JCWHMrxTTk40jGXohJnXM5oJpSiVXFLuFnD6YS5lLAAcY9UwnHa7LkqL6AgV
bCwtStKq9mNa4H/xrN5haGZvmYpEN6p25KLAUrnsENuMp8vdujotS6NqtJw+
09gk06FZg/ZNBBvO+GXr0eCG2AqiI6K5wQfUxBkOdv3z0TujlzZQWa6m0SAv
8oYyrVyTF5HTr5Tf/WOZGd0l0wUW5RSoRhFq8M01xrVU/P3DaNFyKWx4tC0a
u5TV21gzEWFOvICM0U/xCy0U/kjH5NcPI3Mw9S6Sh5WNR4MHSPNdwTEkJrVZ
srOJBjE+cQIZZTRn4+Nnj31mCsw6eqSlJ6SZjnYWwsfuPwx86p9IOVZ4UBcA
6s9etJtmR3cZ93yK7jYxOgmIGfsyBDKVId0/L9RZIk/cslWdaLYGGs5DR2eV
ykdyTeXUhCVH0wyApkalv/J8lVXkB36q0/5vsRDZVppv8VrPD3RccRT9S7eG
wmsSMALhEVOkiUTcQQe+G9Ue4h2X3aTj+GIyGghuKlao1FUMCOWyLplONDTu
Xt8S5oYJSzelsJGc/WzV0Xi8RsTVBO2A2ybS3KiDHIYWtOBf4UGZPZQm4XzC
Ag9rwKDoR7Fph8LJr8m3NZ2bM9KP1p80kJo0G5AnHvTK6TLL9+6klHiAXJii
kLzy8unWpf9smOw0SmpjvjqncDjmzdcBCc0VhBZawfcOOkePksx35kpbIu/z
D4C78xE0NuOEMIRfjfM6CsrbMtrkiHq7yLtcOnkH18c43uP2aMaUmThaHlx7
NoQHleDo50nX0rFrSVZcoBh4/ERoBBjvUYdZSd0TPCCMKHLqF6EbN7IxBriR
Vxr4kjnsKhkLcFi3CSjkNOLUWY94xB6DYQkJ8EqAJUXWpTKXesS6FIC6+R1/
Y5GUZ2gYjskXUPSUOC0crdxtiMcsvYY9rf58tQcaawtDyAIQBC5TeOwYJi4t
yv7WZ3+Bo6BBQ0WqVlVh1lAncj4NdcpsKBXjKc+2kdJwdYy+rz45D0hmc8bV
1CUaZeNswvtFZ6w2XW6CrGKEs+vH5HdZZAqMCm3z01OSi6udFKcF+OnMAFoo
NCzGpegNec00uF66cMfat6F4tSzrZIQdAUv3BnDzps7hkjUcGBMmWOmAzAn6
wTp9wyqMOZtJkW8qRaUGIcVlY6gtYw5DJR0OUUV8YfNJuCDSUggqZQ7KALJo
N2ABBInFhT/IG9uIs/sTmF9Da98WU8tJyyJqWAjyca0GUiA48i5mAFYv/jbM
rehoFCVmZ6K4LmWkRtdGEABU9y6hardUK7s4thPtIVpypqEtAiAu45dHkMh3
hxwvzq5jcqtpeGmMip7o1NNBFXmbg+esLeBnncTFur7eXJAPiCwgJwTT5Hwb
2kAPz6lXtK5OLqaQUoOkcQK8LbBr796f8ysLPzRpAsneebHAqPzSdrx0w5zD
T6ruJsR0p1Q7jr25CsjWJABn/THiwOvbYMjY9GkHW//qwkU50MQFr38pyok7
XZx0pqmC7GECS4ZcQNmCaOlGtXheKe8CpQMrIpXs91vKPuNS9Q9jtwg3rxLN
41vhW9iJH2GyVtVIPKeCE2IiGMRTkrq4Q5qprq5car8/lJ5e3IqpY9t9Fvxf
gjG6fKkOPdPH6N2KoDgFNiHQu6vdZLzYXCIXTIBqtN9GGSyYssqrBg0JGYrv
3yuJbHxScxuFhzdVEBuUKz21JZrR7oDDe8F4FdxR3Eq686OXdN0C+RCDZnDO
2BFBptElYBrjhIp+JerQJNl1SZsfYbL5kXJ9eUdd/5NT50kE9i3NOMbXsajq
THgZj9zQtM1RdwiDxJEHmTCzFQKOSFZqJBCVGctGpl1lgGJ7C0IQ8IshSCJ3
Vpr2Aw+/fLzlKmKVIKAPnbGb9XxrmQXU/x0UMsC2qRHewJeZ3qTRl1WC7+mw
LAmjciNCo2tywmrYXKqUeyN1LEsHasdnnClSQ+9UCgj8cScW2W3+LGk2Mvcj
l36NvKCchImsn+2tTb40bpnDB2V/NWVkmkNFl7b+hQbQWTeapI6MOTzztVSP
3/nmoAwnfMfIRNfEW8rICQInWNP5fgC27sKNk929AuqjB8A8NgEKbRDCP1sP
Xo8JL0GUa46JgqPoaAjNZXBZE28aw1P3WzNFe8F+bcUPZXjiZCrnXXAMhxcE
kLIkJkXK4X7GkO3QA/JpiWNPjSK1jPnDcibvfU4Ys/ugwNK/1dX1Jd2xUw2y
KWOF15thB1c38yv72XFJKi9TF+z+/t/vthXoeAqeM7oxC4PgwnQAxC52zZpW
WP33weC7jSoD32TGE8jWHL15LtygM45UspDmBWfDpJ/0iMz6jYdT58D6TzjZ
Z1kA5nSJVZ1FoUZb4sZvSJvbeLo0QqV39TNUjeySswwRytxABOY820zVxf1B
J3VhCftXPByrcIA9nxLBGhi61ZHvBUT3/2dlSB6IK6owruOu9FiubmdWFxtC
+o8kvFRyEcxErzMDC1Jxe9TKjTeVF/fzhe1rzHw39L0Yb/rn8VryQyqavFst
TOdBwHRlt0KIGUKbIJ9k4L1TFVe7OqTgU4p/1Mkw6/33L0yTVre2rs+Bov3y
Von02kX8JaKD71L/buK8B/DlE8X0ExvRaU6yIrZIQYjrhS/9QEPocwYslXyV
36Zt1rKcqs0Hu9HT76M/+HNcuKsVafH2HhPTT7s5QzCUQkOh6pBJNV7g7sd0
hRURy/tvKcTPA93tHAsPzadQNAZ/SuyHmVAv8WIB0O2hzjw9aunPaVRxv035
xu7BAXZaXHDKbt5+8mV5UdxS3xRvSBJVYAIne1JvucWwYA7Btxr0AHLgR22W
fdeovbvFlq7b1ZuyG8AhFbZ+1Ao2iBjrC6nhXTgpWpW9mOYfRqoUp1V4Crrn
H9x1r/vMtxPYIhtbbbbBMgwu2n0drgcnkkhlulq3k6egA8N2O7SRAqWT5Yrj
ybAnbNsNcJGzjLMv7jEqGim8ZqTuWjMemV0GqseAyareRM5mPykVjfTmK6UD
j1xDR8sGHwezdA5l9/GprtZcCExsdl8F3QLeCIdyIFgq4GygkBOH2hwRQRRZ
UOhzvyIgwkU+hpKhf7df3af2n1VKXkX/g5O3G6JCMO/hYZXzPWGKjNi6RHdG
S85+UwQfTkK0MJbSKijeEl1zwusoI9kzFFIjGW0QxfOiKn+FzhXAZVu74pYy
GotQ988lAuERRAuS5DL+xAT5yjqtGB7P39i3KES+M2XnMwbQjU6nJ3MJwXYx
MBrNx9cDVf2OOND2Qq6Dhg72r14YnExGuejHaeOcqRdRBvi8s1h7WtpjFQoZ
LcP5JU0E06HGylHE9pMd9G7SQpNV0FJolxHiX5gGVM6S3PjHVlJLP6SCGj8y
sajCsEuCfVd8PKHccHX0DYQaumOzjdn5DqzEUAtml7xrYcG8Pi9Aqki78QVw
7fVRvK/AGJEjGzq830H/ig37s7JrQhrDALsve08XylCnXF9KRqMRUZZzJFtk
O221hZeFoah0CNwh6EfILDAn26Olaw33GzXVBSVxNOO9ruGW2jmq7yqzvChR
Qjg2Mh3V8J3z4mi3BRCjN+fn2REAr7PrN49RKHmrhkPWOqDxmHGD1PD/7iUK
OKBalcXZ14szOgGrUY0rHox85cmz1M8Gqf1J3Um432cpKYCYDInMhH/ARelY
Tiqe2JcP0cFHkuLiYtDxfiT8m/jwf5IKs8LDbDrT+30Awy6YFveprOt5Ijsa
vgmKobOlATyA2U7aDHd0/zy5O3w/bMj9udeJyNSrBOkkfiKPwOODwxLC0/51
Lqm/4nRqfe36Aur+FsoWaWHceXu/bHCmb2q7VwtKlyE8xdfnZy9pLb16eaFb
LhPQc+ETof3jwjmMug22OB2uA616I0g6c/IWRjpBpbCRzfhpo/vBhvi+wIqi
Nkhb9mbz82mnqWU8q5PvEibAm5bn235ZdHv2igQu1IWgS708rKm5Vl4rLCs4
kldsad3twZhcU0x2p6WnowRlvM2mwPW9GF0kxNUnbCEygGwAGobI7WPdBInB
4MarCs6tpUPPPgSxAZJTxRiJIwiqdkwjBNc2eIwN/kQKd/yDZTPKkTIfluWn
NuknouWRqEMAmjHHx7DsRwtgoeh5jkKnivRED8g02VQyG8QWGUqN02Y6C5hB
5yuYC/MOc0UI1NFu+t/GhEcqIfO1j20gYXaNmTHyMKZUHO3Tt6WKb0pXldpU
qCPSrach58+Ljuhjuc/ksoYvh36/8BIek2+lxFp0B5MofJztc7euomvg8H45
SSiw25gtvt1TktPwxSebeBjulBUP/RvAT/TQrHpSfNo6dCW60DAXjmjLHBYa
oiZ4c7fTJz1ZAIxn9tfdBfHsSysodJvOBeZ63C30nWS8Pyqq+XXTRFtlWgUs
IvPDvGf6Mt/yPOhlI6ppRvWXCCjtT1EitSXotoUm7TipXuRli8Mpo0whIjbB
aDQ7v1KU6CgPVjTMOuKcn19fncGMH1Mpkn9tEmbF9dr18kbW2OgluTzPzwQ2
vMl9AreFENAiS3q3RK1RTWmo+cl7f39bfu6iXyh/2ZITThuUp2azGCvvbPUM
gyXMpPmQHqa7ESeJ3yYZIwxMrs1bHZQl/AKEYWrF7wTHq2uI/+zJoSXsA99p
zIgXAQWWlGRrK+MIDxp1QhtdnECnSnURemalVYQp2I7rDicRPsH3f/teHeBL
73cFtStxCrh8FedMejW0RZkXW/lqnMr5tHEZFVuxFrfGFGlCSlDDCOP56UmR
XTQCg5aCoYz+n5ahFDmjgksjrWETvTCJRUQTH9hmDUzIoXfoLtucVdpRkW0q
8jM3LEQbfbyqi7/3KlXKZ8dCSTVAmOmI5reavXXyYSvcdqzVMlwM7uloEw6W
va0iLYPJxZ6TRL/98MhfTUUgK4yeXS7F0BX+Wln4NYzeUa7NrMlndU+PJC0j
mLLfoz+0U7Yxe+B4j2m+L6H0+qPP6+CGfawexKgjKAo3KxxGgUDg+WouK745
n8KgqfG9jW0Z5WeoVzzth/6MXZi1M8lWjHPMmUnpLYEFdHijjeG0uCzm0CGt
CpAUAcBPTaOtCbcqeuQl4v47ud2ZnbMksTFPwhSVs4OG8f8Apd7VbBbIaFiu
rWfSIgAmij3kOaQhJGhepBeltqeoaXda5UPh5t3Cx33XtJY2H6Z+NrJgumvY
gq4Vg9vsV2zpw3qZBsTwWgM/jSnYa6CrVmH8apmyilt0yrqZCPHihh0RDWEZ
hOPMc7ceIfI5zjagNLbCQ9LIBEYSlU6oSv2F5Am7bAbW8Rx6PosG2rFAUaH7
4JUP1p6QrBBhDzCHELGYd+XnHUmrJqsLq0eLCFFx/REpmRtiYvA/4AjUgHZg
LAljwD2QY5IpiAMEAU6auTHN9NabdriFRlZVDsYrGFOECHmAe+qbBiSkdBdS
rR6K0Oso7D1hSve055wsHqcGPvAs068KObpRFnG3EHM2yydXDv7OtFCqxmpn
KUdd8jx9dRgwBz2yJ8JW4tFCxm6bpsHIUMezC2yxSNfdxwx77pfqlteNrmOM
LZW/TJhx0b64OgDtg2O+qoOI+9eWUT22n4Sl8icTxIi0bHVQuJw7la0DnnMS
Xew+CChbEgGiiuCugi8gp3mEEvLvTMca7WrWr+S5+9HVkBxiwDt30PklyaNw
qZDpRV1HZViaCtC5TIM1ic+4ciMqJYQk/S6IxqYL33w4ybeoJcw+uRdQ72vS
Icodda+seZJ5yz9C+mvcHmjDtlI/vVU21GBrrZKmgj00RIL4zmxYZ7CfKgtB
XVgzLBBDyayOZFjnkekkp0FFjybXKfZ22JHIJx/WEGrSYTxBvBLhRpGP3A01
qJcpsyo31MTOqEU0i1OoDZfXPPYF09P/DVS2j3kxw6qmYd7meucp9cwKB58D
oWihlNOun167ibPftkZNROuo9Yq7Cehw2wbaPW0K2EWwmxAUOqjk5IWGoD2S
NsAb60Ni7W0aFk8WA1pZHAD4fbxnhszse9/QB8mH7MsYg/h2Xf9BwHQUUrFu
CmppZAiNCmyxih9YPUEACzi9X5cQdO1v+V4DinUedNHxiN4rJ9fhXpav+oca
qvHZYQJkW/LVoNjvcdWEshaf4JPXylTKjK3yliJLRXzONL32k0S2VO3pxAxb
TBbTgeLE8zD4+nFac/2Q9XS0wx+61njxUTOvhZmgJvUDaN4jWNsvEA8Urbn+
YBcK+ImSj6kM4iBEB3recUvGc6XYlYSB2803dGKa/qJJukCpVCi5cJUfSFyC
tq6k6moY8Mz/eL44ijIufaSqbAfK61aciWX2BqxmVTScKpKwZBS6mkwaZBrR
l3g+XP/gXQdD0xsUqZAbw+gLJsVnwq1+j32MSXPHRtuseyhaKdpsTtVPbInU
bi81f9hA92llaW/UUtVO2x2lKQ2prNKK1PFAdX3IXZfGOqNL7IiyJXZXJ/k7
eshKJp2ZTEHZFaW1jkHKSeXSpxPT3Jafh7qLH1+MiLymamJsigyvoBbkDAZI
ZnoEy5Gt5FQeK3vitq9qlbluhe4bpizkRlgP3y6iZR6+6QrjRnGeVhsHk7Bj
ntMguBHlXxuf/ehCmm4mCdQqNRikMFFskAs/3TDbP3coUXEXp8y+bmY6E3OI
sK751D+UocDLE9Db4YeOkcHh/Sa1MkQ4HW2PK2F+cLzxYCiwrXWBLMTSJJFv
HpmtaQ8EqFHUi6hYSZM0coGpkNSN8tlXqmKdD+N45ps7ulA8NVjHDYt+AheF
6IzsdckawSnYhDDvAEpAZMVTmtvFwJMJW5o7/jjfLmTWPyPZ27mrw4y1+sgA
ftxDnjusc/1jKEPQ3Ve2rviJVte0mcMaRi3h0tICajNU71fTLb61vpufrBUg
7fRelLCFrTHkZXYrnZBYk1silMZ0jMUwNAOMo6b1VIUYOJJKhDHHeILYnqw7
/+Ys4WnYd6NzVgt/+E+dJaDPqSzLaJdWzv5XCvfp8KVWDZN5JAdRMVqlUi1S
nE8w7CZ0AgAu2ge2leZMzfwMxkOCtBwSSudo68tkTEGXY2BKs9vFJ2zJ3bbv
8vkuDgTL2+0lv/bmP/VucQTtYyztn/mc6l7/L1phwK7szZIP7BF7dhXcqPhW
08jXkhACVl/qleHInrWLw1Amg5bEtFZ18m8qOj+EYM+YdOlbQfdwol2VKpIa
FSA19gfSeukP8EVTrmTCbrMaqRxHjC87RwUWTgEPBGlpmE8P8QQlczHd2Mr7
NjtiQSbmoGvm8dQrzoRVgBW74Rb5RqI1psDBnJCyrh05jlqN1scfWGfVR7dz
di2yvW4hMx2ruAS/poJBCakuGfMIvZeS91n45KP2clj7dkqMfpZJ8B3hW/9a
A/KMo8xV+26sIsmFc7a0fRTJrdXXhsjyP9BMOU1HOPWV9lEIS+w0ynn2XUD7
Y+atsk65gtD1lG/niLsbYI/6GuxQ+ulCiF5+9W2kXWbfIt0ziRuQQjlfJmd0
TdN2Je9MgFZt4k6a4aBLWt2N+eyEt1vSeiMh5GwFOG4nO14DSe7iDOCcncf3
j+RxTvz8Uki0r8qInlb/lCcKLZl6Q1YVVHt1EFZAobPRqUoCLla1IEbdFXsS
e8o4TxwEaaDuSpl9ZeQIti74J1kcZUWfFQCnL1LJ5RUn0eTVUBAV/M7Vr/yM
lyvLEEkQhH0pq+laLl2kGTQSDknssKgqj3xnUnaU/1oxFkOOrZ68/nT0Lqwk
UkkE/fsgOcfeT1AEzbBQ94a6SJu1IqymJV9NsT6+5TrUXVJya5aH+VoakzvX
aFlA8m0neDK3We8nzQ92Qb1W9uJuVPTdmm8S8JN758CslTyPGDoDzf3ztHAL
sV5Ka+5fC28xtp8BPt1Ndb9o+vDDuS6bWcUKBv/EeH8byMkYS7bXOphK2xPV
bgiGDpzh2oCWR5mz0owDqVPZZ/cAy5l7dZvIX+pPKr4BC6kxoFTC1+CsmvHM
P7WcvOfgfTMkUdZwd9A8I1+cFsj6E+Nl9vCRI1dKTFO52o42yuJLhjODrlLv
FpEuSl/NndDYMrDYj4nPl3Eleyyg2hJROtvKM0TD3CQkwaw7imml9HYZiY0y
wcMJW8Al4JREspO2lnJWJWTMJ4IZXFiCRB/EJNT6CxTR1VefqCdrG6H5VRgq
rYZT3RT7jal11s/Z2ggvHBUxUq2d162ugkm9XEirIZOFOpCN1KcROr30FK4U
s0byPRaqVxPcpLF2sxorByIde++iUfqK9Ku0MYjqgClo/yJTmi1rjddrZjm1
lHUCKCrKZxHY9ML4PfzBcFbTtKAOHkLR2gFJP0YOVnjrygmfexghOP8BbcWF
LnvkHycq3K93h9bbKfE/RMR50NoTQV1rb6bp8fuuj2COBzIgrwjMOKhQWHMg
S8jlzFljWEvkCbsTrMipCObz92ipKvATN+GUk6j4zVkh91dBXJT52Y+HFwJT
HIFG+dJbk4GfCxfHN/fqce4L8tzDA+0uZUsvdbj+BlYVqhxe0UeSfi0MvwvD
ejgY6SXhXouKYa745olmJ9jkzBVvNU1tBBsk6dBEMen4oNu3CG6CRNAvcE84
nORJ6cgFu28upCKTHSDk7SNrcyWG4E2+rLFz/k/ILzOsE2ORquM6egUJZFYs
ko7xWAFubFQCJ9B9/kM3AFXtY30NCOJhdQFGt4I9cLCutIwdh+ndMjIevIrv
klAK1r2BQJzUg2jn4umnTOb+YYCeuAQUu7KXcGYpaUZHgsGUNfXZejDwAnki
dVOIDKU85zcKuPziA8xwbTqaA9xDzO7ehw6GvELphbTt/4wH3tlDHh3H8oRQ
+ujdKtF0s6aCf5k5P3wD2w/phHruylcS1XA6F/SwBPA+YFTPwUm56B+DhZ29
YuvWpha2vF7yHFPGB/XuPyNV+bjFidVdyGnBJfkqjxoQj+CBhJRtiCdcaWVy
VyTg/jIILbGAKsfKm1F+lwywT1zUbzKw4Ubv/JtzV5FCZ/kxDtShNtdbASRU
CBdZaAg2WwEKgyxHVuYjKDDwb91mA2zCq6SLbrb54kil9aaINBuINu8Wh04p
wY9/m6RTrTGW235BIuO32d61IxbWuD7P7xhKrSxlQUCANEv0h9iFy/3aK6kp
UQPXWGX/lnYwUPL54ZsfHDBCj5ViN6fFT0dCeZyDvyYSfuFebdFdX541lUeC
w9A4aSzVO9m2vlLwqcTH2hztIV2Pv8r9U6V767aSsyc4CVJqIYyQsH9mG5xF
i9oBBntVz/jfZZkNYe5Vxcz3GdQITqIUSx2Ftknpguyz0achZ3Ci11vrLy2g
9m0ZynvUs3w9UNIX9TVuk8mhYmXqT52yu7ThbfssNLTwN/rInSjIkGwDppm6
ZSurZOe9mCXxt7igrFLy4WqvUbiVfM/3DM72IuwmfgpeIlCnrtsW2gQ2BZ3Z
RdG4J1ASruWGBUho7/ZPHbfIwrTdozyq0rES7ECxGOQsBVN+VNzQbhpzKvT1
ZjoJySquu35rpbaojJL0XyBbtxIqjpU79Pubs5d1F4Kjp/ZweVwcYyAuTTJD
V144J+VMxK9yD5n63TgQUAkZtpTaoEGAaojpFCdrYV07U8vNvrCe8tBmDeGl
rMkw+/uikvosSuOOIWhR4Mn8ukIYrXK6Q1GV7Z/1eIgsKAnHjcltGzU3tFjD
ry/Wmt9j2oGY6ZFQyrdRhcJ2kyESrl4AxNno3yp8AIIuzHx9lDmRJX80wfKq
qBHgqMt1IJB5QOiLZtJDPBwK67lNYubfX46VBCWtg+TPSAtXhrcuhBAEIoM5
w9vzHD+Ly1hCc3i1wIV2orCmNKJlNUmeVdZR6GXaaOY9jwU5y80PmaAjj2AV
q/R3h7FCoNO4VHbTiMsEo/bnfGFjc4EDgdi89sb5yHwoj2/dpnWa3G7i7gMg
2M7nRT9tnVBS2LQJT6AiCU/FIWBbt3LTdtTvWx+SV5P5b3heE1+oHSo2yiFA
ydHs6VS7a2boZnPTYwSkhKb/PGOef7XIQAm+1NyoYSRpVJkqikkrjEQRczjv
lqGAW4sZ0P8OV9o3bVPbm9kgoNAE+DRCyI55pRnivlKFUOuOuHLIkyqboqbK
/GDhSqUAKjIPg7UdkWZfFyN4MfabaWyvpl+7OEQ6ybqQOxlue0CqinXrFvjI
a9ixbn7mEBRSoP0mSK7M2TolhK0XqxPPaqe+zEFIt7SO0AMH1YrdwyULLY+N
E5UvKnprtq5QVgMYTcoLNykpMYsDl3jmscZUABiVY7Hi1B3R1i4+BWHIJnSe
J43lO55I9nBrYEB1MFqwt7w54R0GuwkbK/G3aL42NseXjWtC7MclY9hiYszi
GPObVGr/JfXmSaguY+lK7Oh8b+A3iiz/3dU2lb28tJJqIjNILPXZ70b9mJBa
PbD/7pepWzCepDkAL3mrxToT4Di5oJZBtD8GAYneBYdkbKDfH0iyNGuFjusG
3T0V9s4iwjU1pGGTc4Ozi7xxNlaSL4jev67ttZF3c0S2C4XDgjX56gWz0jt+
IUrQMve9DNC5OQZz5vFP1AT4dbYj8G6sLV8DhoI17n32lWqxMPKO1H8uPsra
Yza5k7aKKtBaXlCNROKe0HsbvPmx2kDcThFlqrFEsI9l+e0k6i4AzzWaBF4A
Ma0q9j4eu3h9q5pXtfKxTLBbXHIErlRSj5HRAlPPNt9kUWyyI9HhHjScr6u4
4/+M9JCKg0jo9xZ5fnZ45rNNGaK/br3pvgELHCUq12yzMWd2pXPiSH7sAqiE
xDoJF3/jDZPG6gkZnJCAcBOto+o3Y/c/Q5hAZvKf1pTFkF2J00KlcDqwjzLc
aHQszinxywe7LMHdJJkARXqhNIexiyRGDuaOw4EPGrIWo8gEjcQfda/BNraB
69Yf3P4JHHnKjF6+TzWU/EzNSsex5/V9HEzWZXlR4+NXlUV5vsHj8SXTLWha
StSaRVNxMR+9LC4WLA2OmvRYXeyYjo+MlvLnmR9u4t+g98iph5ErfUWZnu3n
wUfPF1VFFqghCubMhmkYW4cLObdlqbeNg8o/EQiNNZrzJunpRIZUnuHLV4HJ
ftiQ7HEWk+be6qvl0T91I1MEk8nrj2rGjzckmOatWnaJ4A+oL/uZgm/IwvGk
97QRS/YkFjuXUgm/UdV4KNqWtApebptNyy69DyNDduLJUeCyYYDAEEs56Jg5
qlLLlUQD89Lub9DqNWZ0rShLSX0JdVYhVYZ21DSsY9tjMG7iBmq7LiaSjkMp
9/0wTOYO6roEQPjaA7rluZv7IQhR8MMUtEqDf75udyUPddgiORZzqi8W8DGn
PUQlPZDjV5KmkA5Arwkqypd5xaKhSSVidokOFWKsIsy9HpCutPIhtdSnX3tG
qQ80GZmJry5hOcEdlgXgmQQgTyd1mM0ETrC+4DmM2RGNQIXApU4TwiA1FTIZ
AdzLxHWSNp/aO+LacG6NyVXCsTpoqwVbXKojUSQdXH9yyIlFCNRKmuHn1EqR
V+2CVcJ1/UStwskU+eKpDYqlAM9syp7KiZOKrHfyQFfk+sGoqbPFiKfD399S
yW7w2KX2fC0RwyBEeYkWV0hWnD9ADwKQ7svjXbllh64kzGAredGYA4SWNpBB
vypQA1f0uoPY4rhsiD1mF8G9+pOz/SSvLccoBhWIVNggOfRPT1FqdI+LtSuF
9+/Foaj11vCSlCm0FQyWn23ElMnLdNDe7YxDMj8Okq2YG/rLhrYsR7nH3cLh
KUPkD8xj1C0NiW86r7vH1HSb6vrEJ/uDATPBRmc7RufFuRh6hzTPqtWiFnUp
UO5Z5A0iq1hJVe1HIurukxDRaar7iVn6eF6jV+iRG+XMvUaYrt+rKwALWar3
XvLzrQwvlR7Iw47HlKTCqodLsi0KDlBJn2IW78BPQxajEdp9WZ2n2fb7TWfk
sFscKqXtVKXuyKb5K6AxzOzvp6yAiKrlDXBfjaTWbyL21nNvRMwFay6Rkt20
NBIlRrf0ZU1nz3Gdt0/DTbmIwkeVwFPJTc8fGwF78QGppfp0o7OJQ7nY5ILY
eHYGiP0I1BM7Uj3mnNvgsnoE+B+8+xqrYjPn5L3+oLzzQKsj5n+M5ma50vrI
k3UO+KxqI7FF9SvWiX1aK/K40DWHM6fTVHXxqw2z+hfyBTw4zEKCJcK62LAo
kMCyNnhmYHSiSUYINY21YDfBOItaf9Y2/VPqZeZcKtDGs3iSNNNqnChYUFyn
3xdSwUwUm5ZEPH/piaAPwZtGbxStt3+M1wwV5WzYAIDWIgzmPGEBmNN41hVN
Ns7epiv7YC+32zwwdUdk9fhC1wT8jUb9GFTUhM+GpSPI8gaLUHgOfXjdGDDj
Oxnnd3gA2Pz3TcAM2Qd7qRqVV6Ij8LpIIyNsxUxaDfFIvqDD+qwihD7KMQkK
qR1SN2fZdxiyHDaRTWDrM+NHy1fB369H2Guk3dV0tRtkMGKwKLvIEA0c6Ez7
pnSBUuPRM/o7nIGHeJHTVs4UV9SUMYkxzjpmT82YivOHQaXacm+6tLOStJOT
baMPN7STu5lJrX/KokGyefficuerzz/PgXPRr9u07lisE9a1vQNL+Z6el2Iv
V+uDNUEpIoG7On+D2KENdnfBGMoUZAFmt1n2xF+TXvpcCriGv3Rc6DgOzt45
7TaNOEcWGbxTiONhPZINcdsPbHud3Qcky+l0ZjE011eude8ryhtKbKqbtOFn
L5h3Ukrnp2YNEsm6dbrXw9fujN44uM6dSErPp1NtGdOs0wWz4uzs/mlRwC8e
HgY8bprtgGsMOWr7SXDUWEUPOcT3398Hs2bFomjQ72rOgXLZqs/XwRe6N+62
0gvLqHXnGNuv+U9dOYb0pMCer0H4JU4GyZEdOhFo7yaWKQJrqQ+95Gaz/Lg0
6uWXlIxatroNS0zJUcVObOvBd+JTkToXMZLrTleaSe3ilA2hm8dU2fKKJDNP
VDtIwC95eliKkSh7nEi3STcKgk4dSRcogH1dhQJoNqE4al6olD5dd1NnGhLo
qkolryvUJpyUgYx/Z3dWBqok56kgOTmyYV8SxJXZWsbtD7KluJ/Ub28Dksn+
jK09kkL6ESJyo7YjPmgDzp8U1R9+G2pDiJZunj7RLyg51fN5Fgwsw89VWQXU
uCXJCG0OrPd9TFRAAgsFbwIdvANcUsJP/HURRLHVILe9MwDpeXCdz81I8IQg
hzuNT5scFP8SYAm7V68fjhtXU0sGEIwdD60LolXFmVvXtCMRNl+u8raHO9kR
rGJ6HAUuV5fH/iqfLplCbO3Sfihj71C2XfEkZNtzJchzb9ySYOmvGZqxr2dA
lAL4RGId13NGzkJmzY+77QZYDiZWr5XY9j1Zj34DG/gGZFbjLQUpu+D12m+m
uwm7fqx1Ht9HAL78IpZLSSsuxyMqkdB3uNxDdin1UgLdxtecMg42HFc/+DFh
h3bWrzWFyzDhYe2T1b3eUgPKGRIAwcav6TaCcl9nLxJQoY4L0scVPnDbuWS9
ujJ6D/Sxv6L4z2r/jPEqG+ujcKNp/nRH5NF773LGniqtYLZcrIGk1JrPM13s
KBx9oCyYt0mRnK8pQ7W30Q868whLcQ/mfnIAeSN1sieiUY+JPP7wkcxfPPxc
yWadftdpcDQkAvgQwSrX3UivA9lyAnwSY2tGRW1nlaIvhU06PGVWOZ/M0dNN
Sfj9H60HAI5ez9GEEc4INpgLRY00Sm5XFJDLktgc2da5DvQGjzvA3Dtp/+i6
ZDmnYjWc/VNiWa35uUAklTmdisRzB949yjtA4IsqY05QFTkzbNoXYHcnAiy7
lUM/GOh73xA+yvq6UeBEUM8u022zFHlPFqoxXd10jGGs0B3QSBuwtcifWXzn
U5gQayHG6NYqCmOiXwgZW+UadUJdawOOe+3zntzkDgcalO5q9NVS4wUVtjI/
TkBorNG/ix8gud33jZqInGdpoXFGehF+LN8Z6+FXMsSU4kFp45XrNHG0SmLH
84zzMch5Vmxzo1/2bjfZEscdeSuckegtK+SmS3cQajqWnokVgy/ectZ68Q27
ZUZSWYjUDm8XoCjERt7mjIre4fUQTQsr7snzusV+9FTD0U4qvyR6FqUMr3JO
GbHOupsccpFqypI5cTI80Wf2RvifhvD/rAu8FH9m0TKxKGvAiLymUpA3Bard
cRhoNPIKROZClV9RUlcyqOnFmf8+ebczbP0gctfi2z3D1j8e3bflUefZrR70
V2DFz7kZRy0PQo+YSOOvULTcN6wdSOkJuefIwp8pwyy+5QXPvHRmjkST4kOT
PbWG7vBinzMP8+7bfHAOxrQ8ta7G4FjTCG4nYQhikStT4kUHxMoMGMiWGTRB
rcn34S8A6j5XDca+KhPu3iZBNwgSeBd3ndarBBvHLCTTC4EhfNe9lDcrAtXU
uQy968sflHB/2au+jrIF7fROL1DiKeImiq3YNeBaBrvFKGq1cq5CSDHF1n16
Uehx7OnDMbv4BMJW4xnYfF3DgVWoIOZOl7Gp9WjIV9O/WAXe12p5dA7wmYph
8KMPFzMnnwsY/7Z+qh6w0YqbJ4IYK7xs6PWSIDAFy+pgZBlcRayGIq/pqFR9
gPd9Q8L6akJhxdvtC5CJUWwCg3VRJML+faMKvubyZU9woxcOz9T5GC6WSDMF
HSl3GVMNSPXz7gmFJ25fmgyZwB8ZYy1mnpjObrgRoHmPay/wwZuOMdX0Fet8
6UZo4uchD5+0QPNBoKSCXqBEHuvp0QtWGcLrxsgWcEihkq9D+XY/o10Pz+Ok
PRNLgP7exFmTDYZkW/IeYN9mbOTZVfkAQfuboAp0WbrQq7H4uHkYo4tFNRIv
fDYYz21iFlMBFgPuZoj5TcZqLSDvWjeZF3vA78EqogP9dGscYl0X8vptyp8N
fEOCzxu/GvsIbOFkG73tEbLYrMqT5NrC5hQlw+kr/QT2tEXg9XLYjgQtW3WI
T268iIswueQ8s/KgqtUd9Yy4KN5eAX5DVba1ItLm7PgtqYc8p5GieG8M6WX0
5KXcjslt1AOPhW+9YHdqi6Bt52U8SFa1gyXfQtF73qKfKyauuoJTKbG9OUPH
DS/Nop1LhYggHbLHk5s1maEH7iX/JuTP9kth+YoSd8e7cSx3cDjDpKQw0t0O
bwm7T83RoybeLY6zEHfpLAXz36PNA70rdUdBowgSE/b//Oqai3NdMRflNE5X
wWsCVaSJmWnRpykMSHd0Lcbt7zPTPPKJX2RQXqq9jK2KJRh5ASNFkSApJEAA
wE4wLSbHes7Ulu9V0vlZRzr1HMZozfG395LLj1xOoxXnewXwY4r4elRYtanV
GmIcIyzbqqrd0mNOLA7XVRHLM0DQmWmGdLEymbl/G/qw9kp7FpMsbv77jfNf
9PnPtlBr51OUyLg8qxEOKn9PSwpgE38PgNJut2fk/7Jn3J9PJ/YUJLFj7neq
aWK5T+EmpXJkS8T7No2iCOb6fJOWpsCPjyvA3B23tuGu58awyLMB0jZtQHuX
SVfrnm4/i4oWC2C29I7FANPJeEVW0VBsP6hSjY7HhQqk4IZdbS0kQp1ff+op
fOl5dklwIiuhN8sglTNBmb4gdnB01lkIl8s0VNpHi74+vKb0VluYGLhTVoA1
ickEP3jXTpZp9ndXxRltl8DN8IeDT0lYjNv/ycP0vdlYKIiqKgOuwjYlLagy
jYQ5QsNFzjXKdY/lRiPZVEbC4Mur8PgLreZc03MEhWQkfBoKP+I/ZhfYELFJ
Rkv74A0Wgh8qBsxjq4p2Yy295W/GP9RugiUbZErn4A/W4137nUaAQarJC5GT
B07NnKNyVpr0vQ3UuTBh5MFyOuNE+2cwRIMgIhxTX5I9RTn9j74SqdD6qm1t
axX/mr+cbydF9H7tnYhSZABtUH8gi/6gX2SSgaYVkvUM5RReTTZ31mownMLn
XAMY+nGGqnjNOWJiTL5KCeY45+jdVVidLfN9SHXOlo/fwdTv7xyA1WtsNAOw
NmLzPH7UZY9Zq7TUgGl3jReJNSDCOPm0aIhlBKdkmDnLBektr9mRhpZrKuE7
FRlRWusuC3LJ6gt2IZrubr5A3nQ5GF1qw6jJELl5Yf3pQwpESy7fsrz1zokJ
0FfovMenjkbExwOw60gx0woUHzrF3+TaKRQUdBfH14/G7+QTM/6u/M1IBw3G
kOrvn1x+d1U3BgUc5l+IFaA/3W0YsYGHilnH8VubHmnmOXmUT7oXhTH6zkx2
TICl4ARkpa/tneMYo9BPqtsUb8uVf6IBBJIsa5X+D2gIHSqbL37vzVKllT2l
vwt37idTZIsHfIUhwbIAdqQ6VkOXFXpXclO7mnzrPkx4EBEVnQOdeSldA+LF
ptARh0apLyHS7LdjLJGSC9dKByRh7QIA6GdoiSSwlrQMmYrSIK/UdvWwg4Q9
9ovL5bt+9QJ/57idbMaZHGomlO0gv+OASHMjeb5JZ80JLxUsMC0+dtj1iw51
We1oqbLuOumiKut0SONyjpe5vLeewYpO3KlEbNZ4no/4t8BgIj2rH5PyYhxf
We8r8ou7m215CUZ+nl7HQJiv8cx05ahy/wiCTzZHYiRQVmcYviWhlFsKlICv
aBhvaUQ0wUy9AdOBtm2CAg+crd8Yok087mjZB77m9zW8t25L/emDSgaENI+j
50DGgI/r504YxuiE2lLzOae5zonrl2a5E/Z/JZW4chZ6TqdreVVEg+E2FWIf
N+3dfe31KW5ZkO3YsHrmdXuPW/7Ljb7jfA1kacB3gVXZp1z5jWbbeAcXJSwx
1eRMBe99xpNGdWCpL8972AizlHqUDuTGaifvL6fuHONcVtPyDXxDWkD5nADC
AVOErfD1A7a9+4y6ckqNYkCzwiUI7H55dtNwk38aRnQqSGoSQodNzerXRr9H
b4U0XopijX6WZNet+HMxha/OC+3ijP04vZzVmZS4N7tMupH0MM386wW4c/8T
xYovpB0JxBYDioLfe/Y83VSuC3GroM/ZIxXxEvtfp8DoIo/7YvyAlOHpVMGe
qTf7OJu1yR3m7u7geLn0GL0j+NHV+ijiBWk96zbBR2rP9O0DRqK+pWit/1RM
5N92pQIF4GMztc4lmYZirRjtys7qDQU3wy5G7S25eIrOUpQoHecXEjIPhOGu
cm61exqZPBrz4FBpceenxqMyS2kVkCHwIBibEGHcFPWM6gXf4lAdMHB/pS4H
k+K1zT+UHvcAEykVn4SevXkh0/vG4+jioR02G177G7Foj4W9KbdSKbCerXgV
uGaaALWLe+TaR0FjybafX8GX0kLuLUdZwXdwdbuEohYuJwSrXMQuUvf9NkSL
hYc020VvO3xYYLFAPy+lvaE2GMKtWpJkIWoj9DsaqzJmwMUVihGaZY+3OpjO
rlFZbGs8q0XqiofnGu9bX6ZaY1N4SU+IHi9PpLDQRxNLmfQcIxImsCxqf9J5
kWuV8ctEAZdL8sw/dYDOddn8RvfeJynXylZQhQafyWOsLZ69hfvt7i05kN5s
6iMOvyCCOCjDB30j7WPYZTD7+GVdomskLCvPkxcQYdyi0rTAoCL1p9UqE5Zq
MAlvjbMJZ8UW6PyGrOgvhcf3KfAv/vOmqm4FvR9Ybc3lN5oGd0h5O11u0xeQ
PzjENS96Z+MHmxqxFWO2rtlFDbJ14n9pjfKGmpbxHTJLMI0uaK1hAtnDlmaY
zEEyOrwOHRRTYiocCB3B7ZpJci8jqKOE0jp8vF5iy9V6pyV/1DUNefBH3QyW
K9hSA3dpudTMYsUzFtwkQ3+KR1/3kCpLI57BL4BKBaVyl3tlKe+PxLLomcWj
Sq+RTDqRpTF07rAA22kqk3xjlWllNQ+paPAhIkOYZ4oJniLKRoYrC2D6YeIq
BXrxF9my3PwINJXsNyGAhpuNIV1z1Rp17sGNdb28psoF4mv1Q1RPW98U+RVQ
ab5YW1nuG+kAI7akLI5hOMI+RryPMAkwaQl1zCJkwIfPyrDmO3l+qYUTMMfe
hlI7zp774AmaX2IhlsC0TzDrtPWNxxWP5WCAUTv4KB+Ng/Qs1DUKwVwSOojK
DH0isN5/cN/szPASEsdD61gXA+mQuTs1n4+9M5lb/sZ1k1jzF85aw0FEWviE
6YKTxHSwc2v7IkGwyiKAyu676X++n4JGMFAOjTkpcAwC5sEl93aNJgQufHAk
V78V05kjRcGw4p80lwi2NdIWkd5Ajz03oOADzfeNtkPWso6Yo3Bd5Gwdkqtj
5jCI8NnqPfyPTFoA4sCt7S+8xZvq+hkqP4ty2ym0zxas27N0xt9406asqF6w
L/j6SV8ifC1gJSWEKFVXhC9womWlL+bie02oZEa3X/RJ0Nrv+Vr4fp7sp/mH
/wuwSG+6ubXLKS+5EWd1Q/u1XALKa/75idRv37cf4qHdLxZ3EZ6Gt7Zi7CLJ
oqqbuFeC3wic6cH924bqnEONYvxgDxT0VsiyZVGacX4iV1U5hlq7gLauEfam
qW8TmlJLXvWR9a9N+6eD+C5IZBk+VYX9C/2k3ORmNzKGUByRCDCS6iJe3VES
M8Z6mdj6n0E7If65j03XV4Q++EFZM82DWUKn0apkY66+QT8zeb/OxhoSll3V
E+h9ieCFkL1rp3hNx+BEH5jKbdNo+SsVmxA0sXCU1KsPcyE8HEl1iny8Y1dA
fBfAvJ5EbIXH43vJzQCAtTIE4iaCwIM/OtTv2nxZbFg+MevQxlWrPj4vskIx
czP2MrPPE6UICZa2/qRonLbSNhpBoFxAelg1xIHxb9GYScSSDrJ2zI1djcKn
gld5B1HYTAj+PqYedVe5Xgl5fnj6535G3qrQLDZ56iL54v0FVaPsANXpOpPe
qPZcZ0ubhfJLtDT1/UXnno0aibffzZyF3ZZnYhM0513JmH9ZwQM5JRakVGiv
Oiyuu6a8RcnmzLsgAKYntz0X4LH76gERGGYvzoDScNPuxa32F2GPSKEGxKYZ
QWUJlamdwXgUw/NsDoZmeSyhKualO6lL+2bUz9PaKmdcjOvYfvMesevU30Se
/EIfGYgQkP9DFu6KwsU9BS9kzc9Jn/56WdtOrC2ktaVLXLhwuO492cMiYVvt
dx5xbWxgGUNMnre2r72m/x2iI7gT1lP/p2/21GvcsFl1RTvC7gNaqdidbbVi
+z1snPRU2PI8UVm3oGVI8gEBkaQRDTp2D9KZCg4zEC3u1GjB283DLJgDI4nF
GX2aV9NIH+UuY/4tAIS0c98QZePk86NBfAfSWqzqfwllr2NGYybPIepMnlHf
e813wpEVj4HCBhL9+XF3g4aiABuCTBHKPpoS7bfeOTGKn3NcUNQDnELEWuab
NGYE+RgpWjIZrL9zM1isiXXXDgKHzpbtcDN/dQLDzlUv43HxlazHQomHrWZe
mXXy9Gw3OUM5SeHR/3uTKnMfHFB+4vk1UNQOdEATL+sYjbLi6Vsi35Ey0AM+
XE+mt9lAaJ3BmVo/ue41RzOi9vu27dnXlwbSf212/d0FMhKXlOT/M9qWZ+2v
9gPTA3CZ4swTqXgTRNTN9m6YlWAnO21r/cW4fA4S1RaqlpF9eUaM32zBeYLI
ONgapP3r8UVOm+dXCd/BD3PxjEKPvAh9oCyXTWSCbJWiewHKp+lQHTgNzkNz
KzRVdqNTfdPNqa82SF7pI3599tYlpUtpEUgzjVen0YmYPXTvWFOVyo5Bqr2e
ScaRGI2ulYrr0+VVxA57WmxvsBbRaf1n8w2XXSgubrVsOKwQjlstNggrYD7I
j75affT1rn8OhaehgOXI3FG1Ohb4EoGHHD0NGB615GlLa+8vhaD6eHvV2bZO
4TOi0sQ+CnRt+tRLS+Xzqlya+fvujvT/PnXk3tU49BJy6L5jR2E2nHQENHS0
j+O1tqBLbFYz8CGu7mk1VTzk0vshUImgs2E2DFUUSvEK/IrcjuXBUFj2duYS
4vOVdrf4LRQr4Ep8tbrLsYtmU7b3RxfXtOA3lUppKms2bzYGWFI9VRJgpXhN
n+rfiqkhhfoJ9w7CrWdrAxK/Rg2CTZWokUDV6YFiu7Htv7KgIzpggRcUQaPg
izEMgWLrnfaF8DNhZKHeq9i5OjEqGNfkPpDEl1PSTqsY7cVbxoONZN0+yahg
zrHVkfXbpRijifU4Qr3oDOP+FY3FOH4QFVQepZpMAtI6Iv9QNJSPAQUIVJ9W
NWFMP5oMTxQHSqi1ANjWH3Gf48t0bx1cA1iwEj4KSmWIEEG04BFfIq97QXXo
z5+bBml+KQkiBIwZyt5/yrzLUd/pXZ6T6pLg7FTi3azXLreq/3UDnhnjV7wX
vKEFmenJeQHElYi1IY1Ham8UDP26z4Qj6FLk6Wf4WT4g7GDH8hIaBJh11e2Y
gbOvQc45IJtMVtS7/Lnh4gWhSKbwO76nn27t7AloSuxYVLwD8QXBhzD1V3N1
WU8qBKTRk7z64DThKG0MDUMEquz4twD8nUaIZq5oKKGxn6AHmEnIp5L64bT2
f52uWVc9ybaQdEIAt71UPFwOnS3P4VAYI1YwJd+sUARIzIcUlF00fGhqNG7H
0F7/OBxEWUheqxdWC00rh0PD86EAp2d6BocDtuWBh2uomfKzaVi1laVl0v4n
6sR+aaHsPJ0xvK/ZeARLSoUl4LKlxEXe0KzvFLL7REk4ZTx8CaxkVBMzw3Pa
23Kgg5DO72lxa2d4Ptt5g4fadVSLLwA1YE3c00KBoG7EAcK+QYoESRt9xM5D
oPSB3iXAmyYv6g7FE7deniZb5qNpjfuRWNyaIFGWZy4zoh3FD6Iq2rIum3Wx
RwtU6RpSYL+BtoBJQI41HeIIuoWH+TLkJ3EPt9WfNSeQUR4KdrTbO9g8OtOc
u7HBLCbREFZJPPlyl7CknPRk/9P+bxT4ciWcwmiZHO2dsu9YKGtWXWnXM5RR
gOFGhbZf55CehAQCX+8e355ocaONQh7RvhO6x1TNWKIZr9KvXAKSr5FJ02SM
Ig6pS3lVOJQdkq57szEfSqBUcjhthbek+zxYG5LlFdkZ4EfwNppKQTupR5cM
A1sEt4cNo0NUv1CAOz5IIxtCJm5GdBqaPm2s8XkVrh2DxOkL4/gvXXT+H21f
BiFl4oG3epGg3mRNi69h0EoRQEXOXu6gNz2B81ujz9Ek151Pc3MYa+XTpmET
ivhPxOaIs7BJ66ROQDuWatX+ag3L1ypCUgiRaNrv2XtYLh9rujBph9U7k2BZ
jV4VwHr4IOytUI7DiC8Oh2OvXN8WuVk8vnS9MF8uw4MiHv3/xyfM+Bl03LEB
CzeC08ZTHbH7nHdMq5TZUv1ZLRThQCdPaSD4k4YiYwEqgnpsWy6Dq9p2hcc2
f0wTN8wx1ls3Zka4ddbj7cSqR8o9HbA5Wkfxj8xZDIEDK0AV6OEfjWlJJpMY
JurzApW3KV5mEuytitgzu8F1wADRMhi9cPwjXVvmcSnz0RIiJvHjYG9a3Zkx
jy9wl4YO1op3V8SMNem3FWrmI5zOmvRCD0qcQaEw5U7mYh5gGelcnBH0w8Ef
dIyl7pWJ1eHECYwnAeMiItHT0IC9XSEE4nHgiH4T/sBfsoM/PixD5c2HR35E
2gxp6Nxw2eGR0f0TPSP8GN6//zSnS9CyYsD1CwwHrUhpZdnV/mlnPGY7DbnV
E7olyXzCBDBjJTWn5vB/Ko9VSEbodFkY9g3AQJ9apxxT3kYwX0Z4MTVm6+eW
GtjEGIotVxPqn5p61fxkILqSonBiJHpUM2K6ZvYDzYd1YLtucsdeMKg75jqO
4+MaTV/N+Fy2cbKWddj39cPV1X6IVVofn8NxWg3L0sbww+5r4boyzKF4puX6
VgO3jrrlFvO2CJemFBeq4VKOcFUchBdwC45hYevqMRKrClFv4eMCkv7MkrG6
PKkxmCLnHdP35dXWerT/idEBx94DeL9qYKDkZ34S6qwACTaaR0JvI/u+Djj/
uMmrmh7SbV3O4Mlrisn75eS+64g8xK+yMh4qUiD36/kzckiaorq3AxvwEnsE
zJoqW3AaeyFoayzLtLYh5ZVHAoJVXVNGceLvo5juXoa3L/nLiEMWMk24evT0
34QCqXHp44pWJ3xnT74yoC4IboCiP2eOvW2y/c4pHFMfOQrCr37GU/gvanGT
GDU48Ih+FG9ksx2o3xEEyMPt+xk4sqp0goN8dUDLUJjy/LPZr2G3FvG8G9Km
GjUm/5p2qDKuolbMswqimJVr47Ms3nkwCufzhTLBHFOaQ6Bif0OsfdFJwp/5
Ybd96/NDH8Q6/lKioXKCykdarVY6llG9ZJ4ggwYGRxSH00IO/j23CRc83kjx
MT/IQp/hdK8KiCRUGh22e00B42QPBWnlIyEHQ5gCw6VIZ631hDRUvItFMjUr
DSB/Ym3ZdRNvHlhqj8yyba91MrNaTThVSzCl7oK0U0gnTtT7gptDdQ3ZY+H5
n6gtIPvN5qQDArjS0aECX+X/IUJuTjhOAY7vFZnh1bbQu0Wh16vYYWbSlAu4
9I4YVr3djht23da9BRBTxVhTp4hfIGGXqImbvzp0ESrE/bNJZCeJYF8iu6Cm
Dr19PM3/6bpbfiuvAJnsGf7ugYUvmv/wNZy8BS0N48w8tUQuMAeidel8YYQs
av/9dYACh3WMvMXmdHDV0ngwOTSUy/U+mI42MPMw6L/coLDPbI5BPQpS7b9T
RUjP90YiGtZx1o9I+cV7+9l3tMxKba+EBaThhMalmCer4X4HT9xnAECYO2vZ
AuCom13b6svfl6w/tYrIWI/eL3ksXMtswLCWMLY1hSgpUHxuHfMjt7kXC57m
qBuxVBtgu5U0nOFReqPGyIIIdUdCuffdvLZ2fG5EVszZWSWKQEUNrZYlX9zI
gB4rRZP0aLC4y+pwrG2dKQVFTtvk/qdXzjGLwG2q50EWIcKBj9I5+CjexMs9
paNhgatYpNWePVLyz3AUmfQBbr0BjGwTXh1uSxeDRKHyHp80ZUsmU7AHZzUF
pcbStnd42p2DNCZjpTGAZ9GYf6hoIoHfEh3N0TBpeM/VbG1JHsJsjm59XVYD
pnCFgKwNieWykLuocxZW0SoALbGT4wzZJ8soSyEntNu9SKbrrdaRVYm5t/Ka
8Vloym2IIXKoSWjTp4pmId3ZZY3qJVkdr/JBSMiz9QgbnV5SCcG+iI1dJMSZ
YkFEVlZ6jj8XEcTuIwZaQu9snz24wDrmgbuVRP1GIT9R/dIixY+odMO9/Zi9
HqUeY5EwrAoUlXwBfp9LJ7XHQnfj0qFxrXek7VJxcVipiFeqR9Lrj+0DprjB
qcVZHwutDK5aJvdwAa8+mE75ONka8LrsbHdr2EstiShxdVGXBEGFWFI6w+D0
TSVH0YBgQikcMGp1SUH0wC3MMQUyFEXlE36BKKws2dh+0fIrbDpArG1wY3Rl
7t7VxXIjJ47enttezR9d7OBQ32bAXzE8vZQzWSDNOFFsUXZxDK9HHQI27WnP
fVq5UMZH4CiiPQbB4NhI1Zax7mo7MvmZnJHo7tbJC49DWBCLTaVfYI5rD/sV
q7R0JBFibmNFc0XN6Xrz06XPhCF24lpIoQ4/SOHmz4hUfRkdVR41gA8lZ/qs
8Ra6fI9tCuzzfAgV9/QycDU4TVcUj7mu3lRXaWXUqbNyw1I26hwkYhFZS/j1
k/XLGCVvWTJws2GlTWfojptF/R4kUx82o5A80s9RfwH7RHMMwva4kl4sT23Q
8le8NvCQf8sOAOIg2xAHsQCY+q2ErTwIL4GvZBJIrltltTptKrWTG56Kq0Fk
sXnRPOq67/A54XwjhngnAx2t8ux7AU6JL2R0kOAQ5sfyM6R5AoaWtFUx8vza
b/y0bWxloOaeda2UPmVqCSUl8LUIoI95wTuOP9bU2EUZIUNGiyXenpW1wG+e
KC+Y5QfHQ/JfRwtAYLJbLh50g+qi7w4j2sgRPT2GdplANeOuXIlKrVonr7jj
a2CU+trtARgqff2h0dlDCUDASGFzIigfxSJuEpBxN8zTfhOyjXNJ5gTW4PjA
CmvvyzMr4yY1BTGdDrmN35ftcAbEjKCh0IIcVNNTYnchEBNiHiMlw5B20OsD
KRkj2ZJAJFxVovdVyb2jzHpfoEOyyzF8ypqtEpG2fSXWJp1aZbF9oPA8JS7u
4zwMoae2lEHL5qcrYMCEeEvZVrmUSe+6n8dZ4jnrVCZBlpgGHDQf6gOkoHBE
ZvHkEYSwmDf9kTmkp6PRTr3N+2X9BcTt1bwfHc30k/q7R9zy6oeR5kB795kj
TFB8HbwEptW/wTU1prFpX2ZNMlJfQBEiYMhMGbaCMrP6LuAIGxl5o59hVKGg
ZtsJ4eradAkjPwVgcgOEcvMTi7eDE/UyG1Lcm1X55bd9dRCdAT2nUWYUpxlU
/5Og2k49mpcE0xISRD8l9nUI6IQ0rMMrISGTL99nrogKEnZwvG+uCuHNkgVI
tESskV/rp90ahP8o9OuR6a3dfpe5j80ZiLKAdOHaY1O0nABienHVd99yMmL9
GiDBWcND2IJLfwmzn9l6OEO7yX7EdMLezKbeRKCLfOj2IOvk7OsN3wwfuNGS
3vpLZBkGCPExBG2fjS9phed3ffSUGFWKK34qU8FbifvYoZZTI/K55GOG5bb/
LHUBUzgKn0LEWLhO2v1EHjvtVjMS5FqsAIbaI9GcFG7ThOng8/cgCxG3rdfJ
vYS5X7WrYF6YYCN8W5JByIsq9t+9qqYmaVYwZg22MzuXVS281libFt9wyWJL
KSn63cCVU6d7ky1LeRagYv7k9gyabXzCUExPniQjg2iRCx/KrIh54MKAx84A
kvCrkRkuoGnfFmmbSQ5fG/CJZ8zLRy3FDG+FXDusOVEFWPh6lSLPJW6eIGQF
TE5giAvAe8k0oLXC/2WeelP3z5l65ldbD5ShEjjv9fxDpY8qOW9YmT/3jA1q
s0RoDPniqFYm9XE1vfF4Kr6HB91b1z9njJPW7NNpszOJ3/a9mz+3ZxDCgEmJ
86gAPfOgkj651LRydWlmMmIdHspec3TxSe+UhIN1Gor/UDpzCJm7G3XssMsy
Z2I/2QHVy6ynDCzPFFSDON6gxFLQFLL+z5o37Ecb1ap3RzYEHtk92RJMtfrV
iPMUA9JLtFowM6YBZqnUOSp3cc1ONhE/GixAQSqMKUc9Cwk5H2RZY71XWcSt
s8jUkE8/rtZyLGqKHspKdeYx4p1TKk14yy/IoNKtN2wMRRyuEw/kFDIqcV1y
zOsCgFJMwaa3EUuiZ6jUij8ckairK2qrWEC+qdbS4uIdUjwbS4h7vIlJubnV
Fecb9yQa8FgRPfNViDl9c5CUAmkYMPFnixNXOCzhcM503Gxh5MKwluEOGwO8
1t2m7iiuMFfvVigtjSOhmzOxbldSihqeASIqAMdXm+56L+Xy+Xu7K2bvl9SL
2Ypedmne19Ebg0xmsK/I2Xs2GgFxBiEi3rQQOtJ/etVXPJCZ0h2cTm2p/7qr
iytbwDk0DzUZ/0xYR+3DvWsG2QSMaax0ljv/Q5L0lpmkRh6zmB8rANbf0L4h
cXvpf2vVf1ThRjrKQWUjbCDEx8B2sYBmKEq3W7javWw99n7z1rh7EBtiJzl/
HX2HvX/HE6nAgBwDMr93SJVGCwJPrQBwI8r3ycFh08RRGfgJa2r8Fy6fXevm
FoPz4Yka51vkFwaPKO+u+bocsFtxdbCX1mt29H5ltTe+HkCX6o+MzYIteUss
GRdjY47hl8Y1lKjA7VVamHQe/J337/+Adt4xX7HQ6o4a53uDGJAhPkyfk+Uv
5gA6+U5Hkik7X455+237eVBYXD7SQNf8p96mRwkBeU/o4NDQhzpc59dY+yMj
wgGxWQYD0X9thnOzRThyZf6J7sYOqqBibXksY3FLhtbjAxWdxYN9BSoVmavc
ELTEU8yPcx393IMjSXlp6//t+5CTgazZro+mzsPgUdXqHBTMXubj6FVY4Pyk
/I7f/7e3Z+e5imYs8tzLh4eWg05lXJBn64iW9C0MCZ+/yGQDAnNYn1iElIMd
qDgeYI7eZybcUD8aZ86eNxVefdky0p2WJ48HMpv8MrPC48L56AhF3+9izbrO
5ZNJWe7lYTN0sOSep4s6n6OR8wSW4ykuw8YnV8ehklUqDcspjUmfgNx1sgEv
xNhpcATh1lKxXAIqvpHPzBzqxEfG2HVQItSGdCm26gmtniysdeoMtjZ8Au+a
fs9c5dCHUmQB4TWJIjsKoHFYRw+gqw/we6x+5RSoDNRA3wvKI2V8IOtPV2SB
FDdJOxhbJKW11xzLfLT9DuFCpl3LpAlLX62mTMVbyxWJEJ3zLoDAeLaLH2RJ
QE5PiuxArY7TmdU6tv7KFF+fzMgRvwTsTUUlv15UoInvriaeL1xbxKssWEMY
8H/TeJp1G4bkwQeCqjV9VXS7k3oB+dmidSyWOItIuBss1gtnCLTa7y1/V4lE
9QvFvVwxAALASfQq3Q51C9v870axL4yR8iy66vSJmLwQxpWFeQjN5g7sRjut
A0kB53anW+Ko4tyWp6+pq5Fa2hp13A27C9n++EKJ7AdITuHkzFk/TymjfbvN
cI3jaTds4N4tcZjw2otMe5M3CmfEbhSohpR0Toy6yaWohP9bC6r1PE2kwlX+
xs4DhJua2Cq8WgzoEyZozLL9fJQs7p1lNaHRZ9h2iYlRdlVuFidMjD3RxM5F
ly6jBIKNeghIuP6Je8YvEo9f3bp+pl3i5kQEWJdcbEmEefNCuo1kxvTdNkR9
NDUXqiqQDYtnrlWazZF5Yet2pfcAZgrXGX8IhA5dTpbqZdqzWIA8zpWmU0mi
w/38N80bOHCQKA5xy4nrfDY27J0z666qUhyfh3I+g0tRnnBvIuO+YCvg1uOG
9pMZr6S0xN7j+i1NOdQ9nt6YqUX8iNL/zsQUvTxrVoc7/FSIkanK6H3jE+An
vKDyUj2kmxBA3HBFuHUOxS3qMyJjYQCHSX+TSXnymtV4qYLVTPvXiGsiIa68
EgDzie6U+7//kXmDpNVoNVzxrkhOkg1h7jBWoEVNB6AAA2PCUzkDsi4wfCAv
01cJ0y++Bu2hdKLWG32+O86m/N8A1FtYBMYUcjnS1uSE4c8AlY6MsNOl0o87
jwEFkXd5xy0xBQLdP/F/BwzF7uWUMgiiiBWpiZvK9UZiO1wQTfNyaM2s9RCY
j2GoaKBL8+PdnA7cSFv1VhbN3AInMiXELlJ9dTIhD47RRbwAF/enoS1UjxDd
bAVgrC2Et/QrMCV1kOKeUsSf/bJvh5CO+TGt47pgMNbPfrYhOaK2UN51E5PQ
GW673I/XMVgqjHfSlVNDM+nh7gy0vOfg6BPi//DHiexGWLPwN6BPiUmlkMQr
ZeFTsFj6czBvW4jZ/rmi/wUs1pS9QRshBc5Ns1iMpHZNuOX3QTBwFjw+gK4q
ZSxan5IlKbcMppv+Ab9aFo14I32JG59l8yn3Q/eR2ZSqm8RpbGNO+GXlIhHk
sJV8XbI0KzuQn0izNHw84cHMdNf485N4kK0vD5+Eu5xFt6cDReMRLTGEhKVE
rxXJGptWYWeKuBB3Je51QW2H56DQWVQkHi6hqBhj9q6Lf5QbcqcjRCzL0kcl
uqdbLPcWxYU7iQWHGoITsdCuLaQRHXWsuc4l9ru/+KY2umaoTqRIDLfHSt8v
wqyVG9cBJtyv2wJ2ct3SyyZcDoNelmqvGtOG1656zyiBWeSSSBKmNUUa1lUo
NFky0oxaWlwXOtXErBcftfqHLgKU73qP/8830HXv2Guzd9Q32lRSHM33a/O4
FlVegXVrljEi2Ja3cedeFoOo0dyCDUwT1dr31YBF5d5GhoSkUdHN70NHPT4U
IWXzxoMsVdp5aCI29hrZnvyC/lfBFWRipnN57smvb6nck63ybD+dZJVwWv1d
dib9H4GkY2zMLmpGkTnLSiTEvbEyYFdEjxLzKtz9GQkPeW++PFRMTTGOxmNL
1m8BFbQwYLT/0lvvK6wkxWaWht/2+oEJf24WcKMdoOZoRvAe1PM/MtRsMw/G
CT0XUu0Vs7Gv/HD7dQ7uAdvbpm0g3EItga/FmSgI0hdVrBpvpBUDABoDyz7b
Raoswa/oNZyQ4axCW3fhnqAHwOB1wN+25C2MKX42fBoY8dXTCfuwB/7JHCuN
bD8dwrgs6X1yUGOJd0G+q81X0z3dpqF3S+hs0FXMV2Lvqpi8cgh7IbCyEESW
Y+iO/mi88EkRZOedAsKfK399tgjXW5A8t4HfQ8L+bbm87lrIfrlM6GLIbjb2
IuKrm9/yB3tvvqmHpyzun7WHSr1V+99Hj/IBtOrpR4cNt+tKxbzh3IlTmlt0
5ZV8wA0e7P5qR8AdMCZzIRCSE9s5x65cFV0ynSW5LmjlH8N/8EfW9ypoo1Td
A7BGUv0ZsCbpfOexs6LFpH7bDFux5jfpU26qW1WEHo4POyFZlMakpHrWx6aI
eWsZTO59j4nV4CgH9OzVEe3Ay79NfdP58Dzp7jjDiKMYXXc+Mxv2dZNFtn2X
0Iljhz3M5C62orZ/BjyLII81v8uazVstLmufPb8kuZuLUDUuqJaU8NA5NblQ
fQz1Ltrp9JkTmlt8EpmAnHl1+zYvdzwDPuapPShq9xE8yAovoAM0pY8wP2Uo
4D8pWwxxeOiHDYUyY2QTh+03TwwvSfN5IZS0JyAGVEkrakpS0gdJwvrXbCEW
GcsoeGrj9TJCeIhFSdDtqc6zerXXkMaJRT6KC3F1W1Y7F+Kf4KohKUpTrJkw
G4HLHYCbqhzei5182/eSKiyGfcGMoLl7NvzWhMbTebJ1PbOkfYGiqYHls4NR
HJSsedX/to9RGBLSmzMRacrvrSU7Pv8GxvNVT38CoPlGRO/ky9dC61G1+In+
Hoe9i5WXMry0OuVZyd767Sybq8GVOPURqy223pJZODM9mAAEoQLlDDymdHx7
Z4tjFtMtzcs8KrC7piJzIWhWGeq2wDz7XQNxDZLkShJyl3SSGBNHHJZGKaSR
zPEYFKTTgvkyF/ELtVnOmvUG1CfDr87eptDSyVEcSG1+Uk+z1usIaMCWFzyA
lHWUCnPCpAAOyQN7VMe0wTZ6QriGIyd3Vw4W8V56co4c4gwttWKcbByr1n7p
tBYILHzoreITpMKGM/qXiy13HKLSUu86GZ5HnKy9OhVXHnbEQbSBaKCmiKKf
KUYjFeCGY659jE1PGi5rdloPa3T+Qfodie2AcGfVWU5Ku5h+QvKY93NDkLdb
FPOLQD71ER1f8CMhep10oOoqNn2YYtt2sSxYfzHRKRKcjD8S5Q7E+Ih/wpUk
P4ZgJn5BbReVFIX+05NStGdkDvcDVBht3m+FpfZK0DXLuM5igLZBP6jUwN6/
UYbvFmNPDc1WjDd4dliMW7aKwq29jUtF3SxdK+tzl7K7NOXIYq7S4+7/4Onc
XkIYoKVyNpN0IK9iLztUgQX9a+AWlVvjDKKNiXxEEmv8iTt/VnKtdnpqHfW+
+YJZeJvM9Q4t4GpAyrtJHxqFFmZqO8VitcYZ6LVkGTYrprrEYU8cI/hIJl6Y
Ke+rg+sunFC3ALMnePCNiHw3JZofICox+sJcJf7xFqXbEd3KZbx6QsLc2vF3
xD3JKBUEXBx+RJdF97+8x93zloGg1Odx3RfbsNjuh3J+nA54oKgv5kQImkxR
BGlHx8toEcaKiYkrMOUOvxam737WtcQg4A/G0Unmt90actGvptyUWevew9Yc
oBJbNXarSc1ewelUN727Y7/ivFDM8YMQgkHnohUkLOCm9inQlashnkIUmEe9
RllNFdKPkPlDry/EK7CjAAqHskeif6q5zwWk796/U76+KZlKC/W537hyQVrL
HoBybKgqTNMd2ns0nBQrIdHDBXUe8oLifbLHaW6/bNZM2qfvDq+9wRTjJ4u7
5lzizzoO8+Yt+S1xzrMuwgOXOUQPBr5Z8aM3kLrZoR8Qzt0JPgyKWq+B7f+G
2+ULrGYGLOptHEmvviz878/wksmT3ebZUQKdUnqkP9NveSeHKrxi8R0pKgIP
nqR1RzpLJ7/0HRXhr0j+FmXFCau91UoSfcYGfsFUGk1MP8WTGP4BDXfhqguP
+KDKUhVDr9RN85Ovo3Muj8LkTBG4+HSn+EObFMOnBzAeTvLqIynDR27EWJv6
GsAkBsQ1GgWpqvKB6MWoj7FEa0oD7cyHOA/mKkOjpxQ2L0zV9mkglJx7MatY
LeJMdezmCtbLWsF4SAbNYQ8J1cZmfmV3nbR2LWY+ypSg5W1EwBfrbBTWC0Mw
c9rK0GgwGX8cpa3oh2alvpi9q0mWxygH9I/qtPf29hpfaN3oF/AbTN5hLfHh
7errt8gtSeiQLI6OWtu71sCUzgKnkZC6qj7+LOxKNePWHd1rG9dgr4fyINZW
ttJWD5tK8crWTVazpKt2BSAoXyK7uYpkHagTqE6zawZMKlRwfuzpvJRhgKLR
O/SJFJBpJToCxaWR1aRPRT7l3mh/EBIR2vqNhX4zwNnwxHEWq5HgGPL5DMEc
WXb+c9uTvnV4hO4ukFN8RoYKgPNATKdn028ARbGlryeDGTrjwR/dmmCHX+WJ
Fbj9NRy/7y+1IQcu99w1Yjd6ihMw5HVrt9GsFDkKtiRmW8Sc5pW3aTbhU22+
buTZCnCdhFYcQgigb9to3sFtxT8eXico3+AiE5bT4DBEW0MgbxU4FDRg9VW5
jMpHs/QLeDHGEgvbUDo37xe4dHB4rL/HsPZWeSUDSvqYhhKkNRDCecs5w+4D
GL+BdqqLCRTn/f/wCXk7fjRgEu8Ue8mqxsgB9T3M4GI5DVSjraRY8OqV3eKq
mE4vrb5/9qS2UuGXW9Tdx+XP+klNYwz/eR7b/leFK89a5+8D+3ZNtOzN7P//
VQu7b6XgGIEu0R9YBKp9OJGdAVYopf6D84E5fwKw9TI/eeVp2IxWrrVF3O80
03JCTWR71Mh3TwiqNQTPnpC78z0FdJWtXq3PljDNePqsYx3dHxUj1b6695v6
sGnlzgGdRzfc1xFbS0VsgRbbx/FcLIbGBsZaln6qNsrIRTDt+loYrhAOUra9
bEzYvo+UbFSNUJT3Crda7dzmor01fV4tsUebZYErlu1+XndUzjocg1mP1j/u
Rypahqae7CfkxjNDyKOpZjF/201NiO9H/KFwf/wJs3OvVHT2YuLCKxs5wBSf
XRiSZjP/xlk7/iZSheZa7fhTSNlUAd6kjis0yXygl0on1acYzLWpepk4+G1s
p3bRojwkZiA33g8bVaVnVdpPwYIoSajNEIX49K4ALOruf1LxlTd3+kEhiiH9
2D8ihXDK9s/mor9vRk62hh92o8N3FVyvKJCMhLQuWeTPzWQccWJ7lDOX5NDB
UBvfJcmtqwdv1rfpDT8zh+wQReM5DUxvuFxVKwDDlOV6VSYy/uNk7ycmEG/m
XrG3V1k+yvFklLQpsITceP8BfIljryj3pUcIYaR0V4ZgEtsLPmQ2QMjUfdUv
ioUI5FVO3dNXi7KkwHrJH72ZSw610K3e7R4UuB9xp0TbkgAf8E1MCtLWILW+
x8wLOwtbep08s4+LojmDL4jLRO4g+ujm5ICAjChPobYRP08EOi1hrB464eSJ
k5whbG4KB2SSINLK0pVuyklCDImiGgF6z6VOVtKpqz8dzZ4UTA7fKB/DTLmm
fRRn+yIeeu4x9DQx8gXcWFxwB487i1wdo81VrR+WdTlPukjU4S3j7WzQiu0S
zlgJos4DNPSrMUmJrnol9/bbr7ggPVaJZTHDNa28fAewKXDzzMxjD4t18ONj
ptGI+WwUS9GWs1XPBSrWyCW5WADEWlELSbqc/8RYArQmudxOjfB8i9oiGeur
6M/V1mf7jpQWDPWkjXqWw6rGvEt3CXLsDz9A5vUTNK60HpQrFrxWMs2a4vAn
vSE5ZZNyMwliV5jb7uSShJqnCLm+85xJQSzl0zD8eLz7wYBNQIhJTpOIxteo
DRUxqZFZmJ0p0x/jF5SQ4DfeWNtRTpmvLQtOPtIneeh8oJJAI1cParJm4LXh
MgZze6lsVrOmMyHgfRHkIpAOu/h32DzTdQWi6N3iXOMrNsFOI8HetS4Jg6ZD
jx1+icjRstF/tNesgMi0CQxJscJlzeS5wV6Cvq5l8WnrUi+EmewS0Jrc4/AZ
9zDShG7jAqTTjajN+0aS4cWfnMgt3Rg1E+8e391yos14kfrdw1pdkDrkLS7M
SMBSB+Xy8QjEEGBeamnqT+iysPneHOJ/oel3uaV/5I/0FIvqu2wpdyvcO8u/
XQI45i7b+3vTQ4umUMVzUR4zfRfPLvk69Zvt6RsH57apbP3OULgot+MEnCwO
mHHsV/O2OrwVVYlH7W//7dkVDzyKG3zdCNXWw3lO05EcO8lYjNffNKYEc8Hw
W/qLtFwZrjc6qzw7x1lJHG7Vswo/G2tZki+F8r+I4ZJ1In1wZkHoo/pOd6tS
fl4xVpp+5h44TASJkmQlNQDgFoJpepsWVCT7GA6xB7Wx2kCAlKVvACA76QKV
Winl+XtVuP8TITIlf78Ya3AZiga5r+gyY0qQ4WJwdR/qFndk2dMyTR3oB06b
/MOu8nUZeeEmJBST37bNFp0qvt/xPf5oON+5WIVLc8c8rJ0hIZNdGUzHqVhu
HVxa2QD+SowOtcDR7wBkQK/V9VFE8RRWxc2RqDpW1Dn8+qzbzSnbtYUzhSdx
7Ojh/7aRwn9Dkm3Vc6hX5K4TWP8GblFfGgsfI1cqabWxmsXdQl7y/kW4YxuP
6EQl9uxHhwvA8+/utpKLsWom/mQaTt4IqJAovo/vgH4H3ohPwi6WVz47gGeq
MPT9jADRTM0u7hn9U9mzoaH77qjwq+UbKiJ64MNDusY9c0J0cvfJWtVrogTh
d/HcQdXsfB/xMp7Tx9H7cnjKHQHxZbKhQrgysSX54PxJq8q3pV33HxdN+/OH
f/2dtHFFpdjB+dnpI9p5Bs9+JbvVetnNcL/lpNKenw6bbB46EL5gPYXVE5OB
5pD262N7jpGsmLoINpqbc2NgZ1HGAz87f6PsaBYeTWPffg1ZmQ/VCCwnTb39
dnkRdjeUOgUFlH6z0ijd85ItVGsaHOQUXDqlMMUj0GLG2BfT4oalGy//fqb2
q8jxhoV4IJMJv1BlEq0ntqtixQOaYHS9RmSyWP90oONODr4xjP+I6M6rFxZg
noEWw3rSqwyaLTEB9tSqMyZvWob2JgpjdNMHwEi7oVJqFlNX9PEYuPknsmOG
tKDVWzvyP2LffWW/tAXPavhDY27pQWW3QPde5MRK8Of3NcVPanyWzIjeCuKW
XvBI/ALTLwirxhIdGaILlZ6PjpQ+wNZR/biG+QBTMjAF7znuG7AFXKIC59NU
sNCjCxDflZr2T7boaChAkaoBA3fVHcgDa8YMLWJEXylIiM+sTCyTjTLxD1ba
SbsYA2pZBNpPvDa3Bp5b/OsRdMnpbyvVhoXfQ1+8MITXUAAooAT7llp8ELWT
xLKoYxCDKc3Gyyk8X/MPmXFptpx5e+/lNXcEUyJ/1PKn6n2OwoYmHuWbzeii
vSSaza6mKWmfgt9iIb8VQAnmURtBEplLtMQvDyIaa/jAodbxPid+Abhz6XOl
yZkndMwtuzV/+iOoaDg+ILHauJQiFVpPPlHjxI2NEFnWCQWkaWjfQKE4bLC4
FpPAQOnUrYQrSrl1BpeEifigPspfqmLnavtJBH2tt+kbVTHXTGhCfuMyI65T
fNS2yifCbTzDl6an3tsbAPwMlLCkx4E0SpJI3aSnKbOCz7jzEhl3q1g/BbJW
VSH+31YDwsEjHLtPlCFiRTOC5PWTuWm/JXYf++mtgFWrR0g4oxh6v6OkGkOX
S7l+kJy5VKczjrebrotCWpwj4a3QrrMU5zlkQiRe3CvcQKkFdgIvZAPqAU0e
542vA10q5Z1fjbZRJs/aA/iToDyzKhHBkz6sZDmw9zQcd20zBgGxiL+vp0bo
IZqd8ERzP6C7MFkIY45+NEXl/A7QweTeGHEc5EfZlBr461tX/zCyWVJVgfO5
qeUy9kngvlUyW9whMltyU7VWGryl9LiTPZ9fA93A+UYq+pA8DVLmPWnbMHyn
ORvi1EUzxK2aGfWey/Yxu+ppD70frsxIFooslXNw0LPEd4y9C2KGw+laiwBP
Z7V3sIb169zJpPYkh0CKwtdFeInqW/TUiX05E/Dr+2LlQMNlpTKqJNsg8dDd
ZcxH9U+9r1N1CCNFYe9oZnLiLY4hVo2mF+kCKTf26SeHYcF0ex9OBBGwYNnp
Av7H92cqCYUVutsI/4ld3uFxiofqX70noNf1jtimAyBnlWRSiO6BQTa4ijbs
m3BSFbkwP0s5M/M3LHaSCOu7WzuapWI16V/opQ77/P26TXyTz2JZfdTPalxI
zNj/vc3p3VTOuQfJ9iTVrHKIcsghyx97a2bCSUxHu3xqGe9k6NGu41UoisT+
lzScQL/MFVHxjht6E/skf/jBLNrdLsGvuZhh9LhNN/83qELEX2CiR5PzFtzy
Sb8cYQdni1mhsanJHAuKtkzbBstILzdPx4wcQXikxJieFG7sGxoeZ8hD/4JQ
dNy17qEsQMcE/p3kt7OI2prkmGVIEWDgAh7hp1iQ2tV0AlsBUa6qwNJSxVx+
EcEsw6PxCuNTiaLFXpl0ZfnFE6kyQoH4gKFcO7J1PCrrZF20J8MtaFIpx7zI
iLR9f7EkWA4NCDPqy1cOnyJkv6RDkkag4SkED/7lEQ+ab9iBrt8l2pobj/J0
KOA8cdBYGqDmucJJBgfpsDQgzHDxoN/zkH8fCb6QMWJN0KMpGEpAIICS1KWE
nC+Qt3R/G+OMv8J+4zWItJg67R0jYMD1wOMVlxQywvetSXt9L2liYrSiVm7d
boX0Yfdby53t1Yczns0vzycg+dsJZFZ83dW1PbKuH/Z1YHC3+szIl2oKYzMQ
Wlc3BjFXXmYlrh9+yvdANfBAcVlwgZYCl36X1i5c0B+/NDhR7RcSb/IuBwnK
0aTgg6FsOmdBrAT9VlRtwl0dFsQzGLtDa440gBYnc82iwK9tarf8nsghyFVf
rlIMMWIvEl7p8jUZBckbildwO8U1z/Uui9n83r9bjSjuSPWn+gEBWPPuLSt/
hTp+n9aHdbVnDttTQSnJDjEO9r0m5L4lC+tYLjxaYIcfiujLOF2C3BCMU2zy
pKvZ0CVxYjmzYGVQAVNxgnaKRmL1qdU/hTKf8ukChO2Qkzc/O5V7N1c0kB8/
FYH1AFOW8VOfye44ToZytRCIpF4jUuVP4usoSEEkywTsM+aGeUTHJcq3dnEf
zBniiISGKm8HwiafyezJvgLGVNNF06tjnURWOKJf1Xns5IRe2FGPCabx+V57
OdK6/10lPbvtvLn7P5A3T+zwPR/1zB1ifOoeM5kxyCjnkkbFHD9n+XSy8qZO
clMFBBEYiKq5Kf9R2lpWZYMc7/NnTF5Kz/no5+wFdMAkkZNxbAx5SVabQjhr
0vfYVD9wjvsJt6ZLgMm/PdbwU0BOXXqtTlxMCZJK8BbwmOyhSSSfSLKv+tTt
m8GBbmHz+8erA52OxgqtveZB4LPMD84MZFPJZuqAmb9FvgejXm9kSeL2omQr
cfJ8Bcy5b88laPYXv+n6IELkrglUDRZpqpTKg/EE9Rb89Q2zWBsohJMw3az0
U7S9nZyfh3LSOHS5JYB5PkcBTSwOPfULGXpIOB349u4LHaLdfCBbGqoedBZF
LswBPIR3JGzTEnu7W99/fAU813JRWe20sAdPwUpLzAV9AWXFzgq4LwtckbMS
rsRQkX8cBCRP9s4Xf5KabjP91TLOWlfHLxz7jwlWBDnYbPXLnZ6Lk3BywENw
SRIU4PMgtXzGgsOjeXkoNlzfMj6I4p5EkM2ZoQ6odnvqqXlr5QPU3E/NKxtB
W0Artu6S1J/OOgyVqiiVdAZ7gnHX8zgp5GNFjpAJKKUU0lwJylTa08oc4RsE
a0d6ZuZt3zO+smsW+HllfXUwrRsCtlea2k+oRGCRgfgH/aBwlrjTfWd1GJ7A
o8mnupCcUTUQ15EgXA6swRv/W9rwZAJo66yy+8jjRTNc27OBzneJtoIkO1HT
eqyWY6XNPiq0oegleRMll2zLb80tyIdT67r9Earw2FuudPTaTMVksb55lgC0
+cAT2XMsRm5HgFEqbKOBsEMA6luApkU3QLNJAsPS3SuA3O8Kj6IBv4ss86ux
ItuwHBjxIVLFHk2vEeogUs+StkszlCjBaSTqDCbuPQ0S7o9BxakfQWag95wf
A9RFeA13uRZB9ped208CgoWU8j4sYdWXiOphv7ZRpVcjFSxnL8waZogurBq+
/VSqlfShCpUipJ/aDYuu4B7DSK9R4hFCvcnO3yEKoor4Ul3BwnzTKcAvlpi0
aLMjw5q6GT9UXOsfyyeqCE6Fymd2n3Bov8m1jFOJzL9jzlP7EQ/Y7FSBmJ8s
a5M77PasUSdSjT3CsJ35UXRJAOx4dHZ2fncMYMsfkKPOV/R0l6qhrEsfUOlC
sdbI9tltHqLDclxXle+WfnrsAapEmYJtb5niYy08LNHOoAN8jEad5s2DmX5u
P0jf0FYjVrIeJqJ1EFQgyCWjuQyK8omvpCnrNTrkUMhoVpGgdw/dxMUXpUhj
+AhRf5WCRKxnnzeNa9Ii0smSvM7ujmnvv1pMyBjM66TNNLy+xMmjt4MPiHtt
SSkvM76zhGQX9JNz8YO6YMtu4bulLHZXsrETqrkkV0B4rHrNzGyaWTS5ezs+
DeQDWJ6yoCpZVeS6TxHV2hpFfELH1iII99pnIe96MCdLSfwRYQH5OLMWocal
Zs4JKKzBn8CS8Isn/bVVpXdGcuVXkTN5HqRJbsu0PutZL4cbG/eWdTwN978O
HE/VD8Lsv4DjTJ1h8iQnPi/d9MQqJCXn5JTh1DG2MjFp+WoPV42CiCYNGa9H
W+OEN61Gu6UslYL7Wgr4Adz03XfRf7oTYWUV+6y81p8Vhl0aeteqofVder/c
aAa6cZ6c2B4GdS1q+5HmLUu3A7v0r3P25FP3qnD16X6pWJvpbS69G6pGg6hY
rEdm7Mg/qXZ0p/A3NCK3x0LF687Tu7mOU7G4ncD1VOwq33tGJPrf0UgRIfvr
80NjxS7a4nfYfSOPOZXeHzOu84l0LWug9xRMQs2smUTaPYW4pixh4u0USeBX
WjtSyV3JFn7+/sT3/sn47KCvt0Uk2lqD6NmiGZNfvlHzqXtT4ijAnZDC+B+Q
FAtOXx1NEq/CIinTagR86L3yn+IF1X0XUgUNTHJ4Dg216U1totcyUXarUd7F
5+QYv13HICFi6GXD0sCCNnORQQJYFh+g22QCsbyb+lmgd41WPB25ejXfSc5z
ETFmwo4aexnVckJ4OE+PMzYaV9uuRjg9sVQuncPrRyePVCf75qxhu5IIRWmU
ieK721XxuDAKv4ol25rr/6dl1fi3ltAebYbK6t9aXifmw/k5rHGT8XVQYZ0l
TmiDp/VIGATZCVioeLgKTpCe5GVX9D4ry0wOF4g0jhMOSMueKx1oLdgtffgJ
YxN1pdgdYSvQIu/POlk96aliMtD6Q4kRNE+3WUzGmtQGdHPLOK9i1gE9iUyY
qdVP0kZKbMN8VoF5Et1iFMpZWsh8BXHQyf2ot5Om6RylXKmldf2cviprN2W/
IbT9LpaXXmJFhFtAVszSl9Hl2/Kc1bX/vQTMwGfPevvc+IQSafGY3/F5wNTL
gPe+rWvebCPhXszq7KSaigtpAw3zmTL+Go8q41QSccYwQI6RS2HXLY7zKFx5
RoCCnRYzFVX3DYDYTRZexVR0V2MEY4yZ2RtfhoxyscCzDdaTE912+MMlvRMy
oW0Md3O77ZoDKQOn7Bbj8zMGu1gAJZ1KgGxhA+nVVe09p3rKhRdvqGXakWC7
OlGLQv4+WCB9OPEJMNKIQupKOSE9ITyA35t30CPNWViEB4x43NbqNTlOjUQ0
riCsJdnhC79g8bAtGxxbNWDjwvSB0DMPiWXtypybvIADADMCyifb6WFcWYPo
SXwY8vNO1v7SPtit/eEgFrHl/6MHD7mrWlDKMusBBaE/QtWTsn9c7ahkZlaA
+q1QiDZOkm2wAxI8kQY1ef+4ps3pDjlSB1s25AJbuR/WfNOXgJJvoQUuZFE0
h/yrrP5JQDCQxmm3BNcP1VnM933a8JOPCiJRV7BLVVxRlQUBaLoLEOYDkLYF
PB/lYBGAM20YdOdOQJ7OUnZkNoThzOh9iULvIhtODf1NzlY8Jy9hmQ1X0Cyg
rRPIGAeF41pSDUPM1BMOj+n7QxSVyz8O2AYzlzSGxE0HaNEwCPHU9+l49c0Y
5anyJGaY0V9MamNscAq7Mm/GSt/us2DDK6g/5K5pcLUwp1bNi8WjDEC+SJFQ
iwL1n2KdTw8fqf0O95gRl465KyYqPM8fQ73oyojZYEFFz089e6papQG7iO/W
Nav3reVwQJSq32fLYBNMDTgS72nGsqZEqyJsXWtRRKQG8ZvnLhKlaNQ02DX3
eF+2yyf+fqwA+TWl44qq9B2ZrupX3qZ+a3PL5JXRvcRKl+aaGK3aLaqvx6B3
4c7uEWK1krGlDB5NgJEMkXQV98gQKVp/JECPs3gqrQtenA2sKtTNFQHPtKb+
vXiNvQh3XiJ7eVG1GqN7tqwr0/crujrGBZACLRQT3UoH/1oNhu9lyD3vcKrz
cx9dbC5RMyZ0kOKvGlCV9yyIDbC4aC6C0br9/+J9U9fuXzMzm89unl0kAOyc
oH3TQUXdwLzCErkjnYcLg9SwLAbIsXKg2E7CW0X3FCl/rGKMLAnJc9g+H/4Z
KrVQO9hJkslpGKrAlV8I7ckFVjTsXBEfzDjOyoHRJ4D5jStePyqVsvh96NoK
/czy7FaDArXKUh+GZetrEFYfm6/9ffk3KP6oWc5oTMiSRjRYU+5/CBoBEt21
bXJRMUtuklCxmlXqS135VlYGl3Ck/ydxyo47URVskCJrckyqvOEEYe+GEoEs
irju7iX6BLVYcZa1L2yh3kpuqunilMG/Ko13hLBLjp6SFRyWctInJm0DRYuk
glIPYGomkuvmPFD8VdmpbgzROHenw97nGOpGgvWuJ9bZqtE3fnhBApnTsE6w
fk72wDAZddUOSNf7iI0SoWzTUkXvFEAGfAl+gtksF4McsvGcNX4Ko64bmbRp
jdt+K+/JUIeHgAMReNRTgcRz9Av8iXOvxBdhu4QeuVgyP6Na1Hzxw2Qwh1Yg
QhdZ08oVOwLbG3O0OlUpdXcvPtzon/W6kltbZSTFMp5/JPTcUM191MRj+EkB
xWDS2cbajQRnZSJ1nnLUDmgu4+DbQ7se1sqU6Z0ZRquEBVeJkY+D6JPj6bil
DqzdraSlCkJSEGrdgZIShWCDTTRtm+rX0wrCK3hrUaB3MwlCk+to8MuzevxG
L63o+UYQV5URmh0uaTlXojNoc3Mw0v5gemnsfQBnn0BRZEj5FsjNPDTvd6ko
5AQAXnDawuQC9kNJcWSFw/42RdZ7b9RFNMbwSy1EoHAbFtsb1eFmmbCd8OrP
QWjaNLV6arCdNvoCNX7kBiaejfmTExVdbBTDTf/ukRrWbJe0rCAI30URhJCf
IiXvZGq+1JZAD4RJ7HR5F0P9IxNAiTOoz71uxvCPBMd66TbSsRCwB7SAK6JO
gzGgsbxKVVkanD6NndufCT8EgcdbkQiLiPfr7c/7nXRfskGpg+ylNUZLx5y/
72HVehXtlOVHjqB/aTW+iqDNODko1hoqw1J575nt0dG4tS8Q9QDQxg76xiAW
hbDLbdrwng7XWhJVcFUS5irzJRO5IKEz34uWeTzMtUnn3aZWXwoZrp+zzD1L
TiR+s/Z10mckGGAsF/lLBFnIjr0RYhDjC4VSe9gmjAvx5ir7SIr79+9mJG8X
dunmCvU5mF7SXzipkvXymAOos0eOfkJJY5ra0NOorRmCBq3/yZdQNIUau4Ci
8VE+BM0s8YxqNZcEBqFhao0rtgDn/VkGXMH2B+DXdvb/MxPurK9FUs1Qf7vr
XBQSzNgTliITy5mb5w9J+6zm0PWytmLIOFmExh4HFJwGpZGlRgEgDIBK0nis
mB9hyni1FR+fTNgHdaY78I4PrjL1EazqC9DT0yrxJjgT4fUbenIuhsdwViYM
4oCL3jyWlNb0VKMp0YvIiZg1GPqBx3v2eVlpb2Z4M7VN1hK24hKoQJr3b8J+
abtpxTt8OLiOJNQiEIvMRZu6WkMJlwiYPJYzGqkt9ZpE5gj6JecXONtD5WZt
hXre0brHoUOtw9laM3XbUkfAxB7nHtOZjwB0fUvnoeC2GWDC/qo95KSS7JTl
QRvI2EPspWSgoXuwNNk7CDNNGFGLV3gBGpx8c5RdqAwpuf1ceihIFhLaBot5
4jpLSp4w+8HLZjy/E59WwtqRYvR/EJygiBScHcPe8YZyQdZ9BFewSucfIz+i
/3hdLm/icjNnQVyp6PAFMy0rYkG0kmwAgQbVRnCc5uyyp+WW0P9gZXHbNFm9
w45p+Jf77ARo/jVLWcbX3TKs7g0SOl7cVtfnbZ8+ZYjkBrFFL+F2kZK8aXLc
+2fLhi/0hQC/fegP0zSIg7BjuzYsL4yY70kAV4mF7uZdM7R2halwKjw9qpZH
FBtHR6lsNSz9LozZuJ+oDF9wBoO/IVQNg3FQSov/jeq3AsP+qmFkGxptICoe
9wMZYICeN8ujKUDld6bDVjqyPl13k1SWl12g+n2x6wLD6yh+KD742HQKFdC5
XnJHwnTPJ9ZXv9nPBLm9i+kq0gf9LaC9eRXuB0ccfdYLnRP/6axNEc9dtdW8
tJGbrf51YtKrn/lPf6r9P7lB6eiOxZjJeOkz2+IjFRih1ydE5qrBgLaEDjcU
9cF7DrkR8si0g4ehigiGQhEVBkX1KLNlswCyeAk0OLFZtCIgkxOAvzoI64CV
InFh44EhFk5oVpNcdCw7cUPro3cXAkg4ipexsTMZmF/dvZTAndPFhQUO4gbs
RNa2rmYtHFlOl+xE67vAkYzD1LmSpIu8nJ9C2Q1C3LX73POG9GU6LkaQ4rvv
8NZ8SUHj/NubyHp0/ah7L5Gf7WC9Fq4KRLrMvWVkasNSF/hAhvpJ0NLs7NE1
WSwZ8fzvEEvNXKIG0YS1hEW9Sn/sge5xs8KTX/pAR5/dhccFhBpGtftm7c6M
mEa8Xqx+GvxYcfvq3o9nutf28xIrbsJ31nnljVw4EiAbk4XOiMxAGWvw7tq7
IQZagHVh5tz6Py0G9Xd5bi/imRxuiSBn5o81Ybvn43wqbXHf/O1RvkmB3H3o
fCvhlyouBgS+wr1ItVDWpqSqn6qjAJSHWxy19tHUjJ3BUxHjlyZqSLUmFcs/
sBE/34zUBxw0n2qkQBdvJ6BDHcw1d/rolX4B5fHLF8tIMTpS1LSq+VzQZ328
F1NhaWuuO35Vvj4+i4x8zbsC8fxI3Hjorgeydlz1yduQy2tRu+Aq6/rAx5qj
3kJADa5K2YxV1NftHDsclCqMZ9qirBr+0LiOG2xwh7NJUsAvBxPGwISS0UUF
ktRmWfubTLECo1My4WmLgCxCHIeOvPPDShb5cGH6OGQtRJBSizemkAQMROMM
wvApw90pbtim5n+5lzstWKTlnRjvt4/GoOXvJpjtfwQkcN0tBqi/+cO9G0RM
Pkmn/t9z9rSqVPCY/tZiNWMpMgseGon33Atl+L4D21X6FKk3mN4AYR3VMYt6
lGZT5SYy2IG/oJLYoTouWtHEIloBpUPoY/BKqgYtYF5LK5nUltLt1DWa6Z4z
DuCYZ0cw/VoeyHs7rwfEHvapfy2X6rVd7z1EQwxW3xMjR5HQgEFUhJB4cBoT
gsndsH11dPyIDq4kG7w2ATrk2VtbBRRXZI1izH521E3Ai52kd2bosLXJBsur
U2/Sp6YhaA4GcN1LQVRfHT+cFkdb5gohdqhxjcsH1YY7YseK7W/G6LR8FEFX
1NY2xVS7uhupmuJ9eU8P4BHZcELAg+P6r8nq2XvrQD7EFPDIjtrIeVCxWepo
hCKD3Cjh1j83b7vPZl4saMaeC7GMN78A/v0/4T17wP8ckxxgRowQ6wwksPg4
uvqS/TSN7Ar6TXAI4T8S6DwU15+bbCDBY5lFZzH8s+e1D9NTuc947kaJSD4I
s8uXuf4XHl89nJ3gv8Tj5LvylyoIUgwNO/qymLelsRXFMPZRquh8ZBZTjc2J
f4kOdj5ySvlwJG+/m/x7jk+p8KE/pXBUowGlAufWBIvAFPWX2iFg254D50gp
rpZRuPdQ8Urlq7dVu755odM88HUUqBvweA8qSLog2vTt8oOS4cparwj1kMSp
94KOp0e5LJh5Iss4E21guiMsoOxN9iSH2nHeuGRccabDsT9CbFRQA3tvpy/D
8zYEOhSgSfGgEBendTTt7RwwVoAkNC1wxfB/SNf2jvsyd8wAm+IXcdaF6uft
u7C7fctTBYQi9S7pChpHjfbs07L82wq8W/X8rC799TksnYH+aVYP4nPtkIEl
HaqCAjOMmN2CKzUS7R7F4KfshTuFLX981igNDRZj2T+NhBDSqoNdJBApsVfv
FPYakTHPhVEC+JoEdHqcsHiew0jnbzS/S6Bfo5vP7d3qx3r7hmsUlzSjTGML
IsYyRnC6+QtAX8K2Q/JGPPligKh2B5u8i/MGBlfvH/qipmlP2I/Jc0Ky/kOK
bWzkukuf5i9ub34s53mbkbV2onrmaQul6OZ1HU6KIvo0u1hk5OOVL47uE6wm
2/86fbBDdAdPijMa7wB/YPXekt7aWO67yarlJvJ/XQPUc/rZZeXsazNjSDEy
1N2ApQz58yoK5VOyIbCmAf4vgno0kBO64rXUCR9J5dJZhJywHJg5oP3/S2ZD
TbU1by/B5IBCtE3jjytu/nZwCq9W7TS0Ft34M8K9vEdgwBb7PEtuGdFrX2V9
MM9lrjNV7UicGtXQvpsdj5EY0QFXrbfwXbIX592L6aG0eLr8nsEOe+ruwJ4B
jlPJaLVacOSweuf6cDb0wQvbkkmVnZrEGpzSDWQE6ir397JUfbE7ux9C5O1s
iZqHpc6J3bIy5iQIlcVVTJmiJ/Is7tJbG8ldAdnGT6wy8onkbxMFbgypNC7S
/2ozWuGv0raC0bJQXcqCJxLoc0R86Pdf6/1mbCymZaVXU/k62gTYXBdIQKwL
gO6DXJQpCsemS6QDMTHz8FmJ9+wPUDjXb4Pafcfb6V3xDyMApjYATjsqojZr
us1fqmSl4oMre0mnNuRCeITvOmEAFJP4exNGcv2YttwUudUuceYAtktlsnJ5
ix/qldJBVMsxeROuU+GNZmUpOw2yzJoPjYfBZBfTLH4BrH+aaf/Hg8njd7ul
Ohkh2jKNu+JdEc634Q4l+Ze5qo5EcyGR5h3/HOyeuVzd8dvTCOw0o5cC2zFe
UUSOxJb3vwSL1c+nyw7LK/W64WnwH3LTn7PfXuT0HjDEZVfyJgE97WktgwaS
NJIQq1iz8jNIy/0J2pOYEH/MM0zhH08xvcq7he35jNxeZqtA/1raPMMhIIBL
GCB9Hhh43J49Z/3lLk4V7LXass5DD7a9JlCDjcJWH61L1G9ENJsc7oP9Gyvs
JofGUz4PBPPN0b6jtMvmgkT6OkZvv6YDpF1e5aypGH751ui1WC0LCyHfItLs
mzEbzWMBTUhXDssUM31+WBUTuhERuAYx7UP5Wf4wrbwLQ/ChjkgtDp+7dlW7
Dbb6jyCc//pteRCR3xtkrB7SLTR43+NcR8uG2FHIAC3s9Bf8LljulXctZVpo
spPcAwCzjcHrDKAO2lv/ydu34Fnkv8PG8AwemX0TvAMVk+pIcw0pMejfpsAR
+fg1PJ1/Ttng2xNbDB0I4zcVjmkMOnpSmtn4NMTMGICmmCfDovwQiuf9og5S
y6+tCU6dmt2OmHGggtGL4GC5UipA1pePnfBU3cgS/QTYPys3CXAIdem8jTLN
atdZVggKWQcqUCnWpzG91Z42m3HxHQMBftN5v4I56Ro0BvQFjBoiLztRpjE2
Xa7V9yFEBer5AYhl4dYYDHDES3+gi6hwbv6q9LAVnwFL0WiN/7FDPpFebvFC
TsG2h6t5F5phL0Dj22LsF2sZcAM/tg/0QaVFozLBRBKU5IWw0PYp2OVaa4oh
qKq0Q668I0saQUCcrrVyNrtbuM2PzD1Keg7clpjWFYSbxNXYqTE7EmxH+9bh
phvj0uMVRhxOS3FxhllGyHr2PiZiqZqWfpP4EHflhv/fRA5ZhzzGPNTfAX91
VSoT4umbPtPV0/osRIeHGGlBLQCjdxEJag/r5P9OGwE6h7HXxKcwmCakOvAW
gQkZyG+zmC/cFA1u92TAnju3qpDlmCMRo+6MBzvDHLd7QDDLeBki+FRXEvJF
JbCDPET+bZZKuNez1D0pPhS2Xj0HrW9tkUUds5xslJsrOzbGBO4yktJ4wo5N
XZoEmm7SN/MPJou9qAG2puVfBqpSdRtBOD7HHi3XkRJe9G7Z4ZsglU1NTBNv
K+zvQ4nMxcTa29EPgDkmxJeWCOH08L8/o+Hi/ZyTyd2Ypaczg2RRL6q5xPef
n6g9YXwnZ20qRQLYNkxQmWwDyfQPDlkJAhdSaAs+qmABzqKg0mG9Gde7ilrs
N+8rpXYW3p+fe+NZzSw/R0tQIj7mBkNohPbjngqr8vxps5pKWNoRuPZCzOvo
+5VX99sLfzifrkMtLJ0S5mK2UoKIoT8K/+qYnu/ltPjyTvMgO9Pb5oMDzQl0
+o30rTZIeUVQI7ynJkYtXkjfd2BU9rOHKOqg3qBf++NJy18XwFkIlIGzUvUp
yC58f3ovHWblG8kYWA7JSCrYXVppOonAjiEJIyeMu6ncYnEQ6+BaEYSDukCd
6OZ0HPArR62uk7d4oUVn1ee8u+fdiY5hemzEKFsgVIp01Po6kxiN3ZcXre+8
k5NwxH6GaJBJtNk5aPLuFYWJ9DVKIIze4wxhNjA75p5g6Yv6QNjzl2H7ogwd
JBacK2S0vGsCqfPZOqx0A35RRiaNRdMyvfbj8hYVo6lvSCeQ4ejuj0/w5fXW
6uq1lzog/ZyQu0Xhp0Y2Ymdx1eiCvM2ASmKnUUk70WeLpBlwDZcLXtcgT9TZ
Q/sbMjm/Yu3/CQdubKsk/VBntr/pD5OLsPKl4q+C67Hn/Rm4raYQgNgHqZX5
VIh40rAkdtDksMzBdcKNUmYFg1fS5XByPW3JqaYF68EgmSRw8bJ+aoVs22t0
StfxHNtYiMCdsjRt/uiSSWY43Jiju+2TH0EoeriB1m9Vt2D0BKKTrvEk6Aem
QkbCAbr3b1J5OtJC/kKvfnydrFXwNmzUL4qvlN/6tXy3lb9DNCrF8dn+BUvV
b+sOgS+E2Ps91rLnq70TpPKOc/xs6JUaSvkOYrj8yOXjd4uKE44/VGF5MZJS
sSMo5DysGLeLdbClthFB8j+FmkU8PYYzE8LhlHaCNYYiiZCY1vVQlNp2aX0h
Zw/zPTXjM6doY/73rUjbnVEU2NLdaDjZLy7J3jIRWPndPiYnSuOMpgfF5N5q
tCK27igP+F3If/n4OWllrDLNxZTZMCYsiRQh+CgViFcTifVBjI2QOzj7idJi
ab88LUxo/nD80JYiNbJOMMdpBv0PNQcTsnidso3ngWXDydzSydd13xYkqsYK
MK5sh41WMUGOrgt0HGTuZhLpJTIcPa9JG4QENcNUgR4fCQXRICgXa5DpVPb1
HoQ860ZWR6tXC1h4seWy6VQ1uVr3KucaC7vGvRpcG0P3TWREZDGsXq15HQ1e
q6xhIYGSA6YlaKD2hsU959Dmu/0IsOKTJQ2+ELHERMTcRDX+3c//JNM3q5IY
MyMvbj3neKzMwPppx74F+1fApb72kvAysPK09qTEmN+cOqzQZfxO/AFgOAtB
/+0lZ2dd2QaMkOAPFgekwX5K69tOSx5/blma17B+z4k8mW/LRtmaWngO3w3z
DjMcwXWE16JhBPrmffV8V0EdpNVyhKPz5oUBmOEOZpT7yWJoQqQ+FcrOq9g3
+l7WQWudw3UOuTiFMK9E8uTXo2FBak3u4IuI8guZ+ucdxE4yEbmZSlhG4Bzy
xEWD3TZQ9EsJMrMOmgsyK7Zhz3hxUgsxivBs0LDSRTUkyTpyVEEe90rtNqfb
UMeXZx4SI4XACOafvGfwTrscdiIOpJeID2KBgqiNfLQZ2IG27e7W40lQRvQR
sHYaeX61SiGm/cJrACB5NTiYKL0nYygaPsiHNMBWDU4h+j+UlY56rQtkMjfV
Q04BNTLzscSN0Sgt78OtPJ0hcEGSj2RoB1k7WFnIezc/4dM0gX8BtGixFqCF
l7POUo7q4avsYC5CLhJcXusCvIlEwdIB0aY4sAw+1gvL8jupJWIju/zbjtyU
jLZBHFITDOreZCVk/9g9HbV5kK1kimZTq90oUcVS2MAl+TXfv/ZJGFeEINSh
hiMaeB17wvxq2y4BxHTD5IwPudcxDQzEPyNwOsHpgiii9e1irUaCYLk94VLC
dRQOlX7SLgz3M2HHUSrQAvrfUFmL/X5r5lCrH57MqQ/JQtxGu7hZJJJ9+9hv
yQdHRhcBpYTUgktB50s789dXz8XOkyFBZ9sKxJNgSihCD5854gb8pLLUxTD8
+G87T+RxJr8glSPD1PIYejtG2P+GJZIS/Hs5Xna7w5IYdNr4JNYW06o8R4dm
Y5k8i0Ksy0ZX4KBc/eyWtHUqkOYoajWe8YFAUiWhIQRB3J3sosupCiG1hM1z
TKcKWrEFY12irR5YZ2qxy7B1yg6YHxyOiWuulGFk2qU+qUNgcPQDHbebDIzv
eSshyTabxiBiicle/sRexFctEw6j8M+E0H89H1GkaEbCvIcQKJb9eagtq+R1
8NfJ8aB9+AmAFsiA2hizSGuSG7yGvXx0RZJ6KeBNkX4fxk0o3o8ZrgX/0g0s
KSmExLRSK4f3Fjv9Y0GVcw52o8pKPcLrsAtycBdqW6RFa0Jqg9mZb9Kr0Ub6
iY7ntQ6iZUISoJSyDG7foyYZ7cT0+WrF+TQxAlqBfPS21wt2UXkxkwpFv2v/
hjGKbSRfCGkhr5UiVC3Sob/Op7mTBcJVJd83D4+DnAFTNDNgDf4zKnciXgxQ
6TPBlIRLWEFGge0dmJE5Tnx00blwDhA21N2buaDlvBmxp8jbVUL4hNvr4F+s
iXZm4fwgdO4kEo3+xVj6U+cFSU5Jfqp+LfaAC3ZePm8auKo+lEFaPmfjDlxR
9fjOdKExCP6lRXHrjOONExxb1eI77qZEsx1rXPjl8um9EBnEDxjIioFFdzYp
ugb7BoIigpiSn/AlaBzFLdh1BkDo6SEh81x8s96vJYNogIVgt4xrGr2fxacp
QuBTQ46/Brp8uD9C8UTcZ3hCjvV7y1AFoDKT32UXFQbsId0MCGCC8WMikcVf
jJd/j759+6aGsXd76t4e6EBlorK2MkiUw5CTzcbMZO4XCjRM9twivRIpFdgh
jpqa4YZ3XE0/bkiT9lFYsEZQ9QrV0LjpQLv66XTVppJUBiy6Lf3SH5+LeqtA
xVQ6mdcy8wfyB0KbsMAFv0N4VUWS3LJ8rub2mvSFzSVjGUOce3sEjFw1k88g
dNCHjR6Ug1F5yBjEDAlKa6ke/c95OPGEoLXskq2d5mer/orKw87raQVsnnge
iEDJGoeNcW/o360mvxrOHDJac0zxD7rjHbJy3FjWb2uLyqTP6MC0ddSxkAfp
99KERrdnpy4taAkNbm71sqUlVlOIRSWandBxHNRLBmBkDiMGKJu8DTfCsGo7
5SJkyquJ77tLnriUgAAaQejRgfHYkyVdXZU+vsJtsSQtR446JaZNvn3HmuBf
wgWFVHa82F216aNLzSDk/5s9j0wdQCdGenn941XWhUEXB1noUolwH1AMRvMA
7N5klNQsqzAI7/s4p+kc0j62NuwzFnwlQ0RJFrYmyMhI6o2LfSavnb/b0u6T
u+HqzFd9TjHlIpVMIqFRn04oV1D23xrg4E9ZdfHpDzrSqwHfIiWuqTqMqd6x
RYJOipQtTxORq+j5CLI9rerObV1lknyWwCamgsTgHm2G4fAKK9h6df/meTbA
Nu15YFmzKGWYuoHB4hUC1+xwSQ9iwbD9Qcv1aL6+v1/7FKWw5gA0OCt75lnC
Zx5BreB7w6wgSl7QNc5i4fFIBhY+fsnh5dzBdVXbAJw1iwNqhHkUrcHPZU3Z
Y78ehj17KK++xLWsVSwFJAUrvr7HST/ietkLCdo/2dD4DLC+ONrtASr0V8Sc
EGiVUg7nt3lm6kIrCt40pSpyDlyc77McihPOVC4oxkPuR2Jnkpbu0Su8CMl4
pjCWOXpjbqIo+KdEdjgwguYHlgjLawkg9sJN8E0eaVMGSVscq/5KMILWmLOj
z/x0fjezS026Bs+DHslhUzvnpnN3PTtagaOGN4KGp7h1FUpx2ecv39ucogyt
RN3vrA9nGEcJN7LHAZKgp//ZPky6ohpyV8O2EgJFoUXmJd34jjuPOhcHqpQ/
CJ/ISiedPDBFXiMBK9AuJJyrskx8jHbFDxtMycE8ssPvS2KR553SPdByOrFw
Cv1crhqusQb19u4FNzSi3nRl9dtPd7wRJXzTZE1oBuIh6hKLVkqvb1gLV9Pz
ouLp5ROvO7bjAx0xoIStpSzLis4e7uGbu+dqWKyUvtFB6HGdqsBV19iV5CpM
IStAn7FtKOxCC48NV4prnANe+u1awOR+G71QMYMT5ZcSkXyTRnZglcgWpcu9
isIcBgeoZ1Gl22W/h3u1EpveVAjrSC7RS1VGf45xdzl+qzCYHjMvXr4EufKr
GorUhPOcWAqXKo8HreGtpt/D0bILyykQkR8z8jpfSnOrye9uEoI4xmBSMX9t
HggUtYTp7fTctW3D8FD5aU+27LS79ASHA4eV1Q+D3USVSTS0DtlCuuqyhiGe
TRaMq4q7MXH+iXw7rp/GQpOQuFxxehFyIuhTgBpqxiPRqhn2UAaetmUn46bG
mtOONDTNULNCHCPtMmB/dXlhRyt4hYjLiOOcWGH9UXnCE2BrPjYFs2VfoyJj
rD8e1RaPC+7ZgNn70LYccE11F1SCulXErZJEuRonfD+hJ6eEVkhKLxCm+FkF
rc8gwQacrBzYqJCXzkFXNXy4y8vPjDu7kG2OnA84TLEHwYZFMP9YYD/u/I1O
+fsA9mxBrizZhhG4BmKGMuRloHqPyKTisTnqbcHy731Z9N/V5ScAbH6tfNj5
z3+qpZQWSFIXQW7GwuYrw227qU4QMYuPEioXdrueuW0tmkqHe0RRMKmi59lZ
yR4fFDvcxx4yGJhCPpME/c6QSHt+DYX9C6qdVdKPgNW+FPUd/1JwfwHkPDR6
z+XeCBp1b64uM8FAhAfNoJg7yBe3iH+t2YIndh51SVojOgvWIjxCaQ/9hCsb
cRWiRALcoDKBNRPv+v3GaUgn37v0K2+SqGp5a1/JW3bCGtV9wclMLuHpejrO
R4KmT9PNdSrIU5Pb1MjzXjrZmg7cotYCu8EioNzzdB3A9u2Ol0lHEh+zLC2c
aJgCrT8kyrtNuZfEipNB7SrnHU3q3TFvxgE5sBZTQraTwCxckGxSqiQU6Bhv
y0XXbk7cOUwFAlHQpIUpq7pWtTjxnyY/ORIjKRuNYRktLcywFbNsgdDvkCen
Otuh/YJhCfJ3EwGyohwGlOL/WMHurvKil6FFvliCAwX7vY8eAgrje224LdNI
NvJ5la+wQwE2RkEqDZsUvtge8VL8uOxcTCMlQTBUDu6Fk6OzX5eEKCfM7Zsb
cZ3iLCa8foNtVRhJOD9bqKsDShx0Gy0bQsxmBsZGlKSpBMmkOuLMRE89l96F
+CNga+Cm3n+ZR6aOnFdHHTG+9YP66AUt1k04UezLkV49L3Sg+lD5v9/d4UCR
2KCnDzaz2DIpAo1G7kCs2N0H4z/FHhN4L/FjIuVHjaZj5A88uAdnKWd+W5Co
Vjvr+D3SGpSRb74EQC3oVXgK58V8XuNtGdKBTN2vTmC6Tk4PyGYDOKROqX45
Indi1L409q+gq6w1mYm32ICMVlIOnLX5vq382V6yeWMejNh87Z4nI0eE1+Ch
gxHdeK0MlTBo9zOJMg9cB9i+h7Momc5ZlCCjw7GfL7k7CWYAm7weTzYp/Faj
fW+Q5VkdTjjzV6vC/6GHhfUnXv+v2hocSb58XTlveTk6Icye0naHxDJnih4V
kamABOV4vGJAOPkRABSCbmvjcet/4G165amwbQRaIyHFW3hsjC/CSp1IoSKx
sq/xKjYtxHzz637NJ91zZ2JZ7eNLaAwAlSMnTNlNvJLe6Duw83aXJi9mgvX7
eDWtuxqalimMFmXDJrbeT3wxWDUpHcme7s5luJXRT6KJs+z7u6HJeOMwbe1b
73YvgXTtS4Ri60B33Zxx3inv4kbkqJieHQMMSXRD1eL6VWcZT3ARL7/FbVk9
D9iUyXl4wUwIcK8q8qnBqxqrXerBlRtG9DTF6lwcMYDpzoeVa+RzusTnqRQV
R2RfRqHxYPnk6dQsnVZ+BiWi3RlyUMdnB2SBGyKpZs0WslryeF9eRRamyIK3
kffj3p0c9TPzPXwJEef/PkkGwzIP/DqtcuVz1XzkweNmipwYGFJPAW16dgy8
Zuj4JL///TgL8p99X0JzsnwH/DIkzoM8P3vj+vYZnsRG5Lsc0LcgjuVNC+YH
Pc75m3CjpnnKYdtsD6Q13piZsnaUPrPvmZAcXqIYZUAM7eTgWxHON3aue7lI
m2krRdeXVnJqntd+D8+dvIueJhJEhN7L1DNq7b4TChzqlIeleJFrfJFEzpJw
cn7pbmDaNufUfbGkBGwV0rzAZoohUylCbtcvh+OXwmGAfVLXKTgesMTuOJ0/
dyNmTv8PUN01PjDTjdAQb1DVYq3Uy39xh91MrH/3by1uOeeUISK5rgi2DyMB
ThyeLy9Om+xudejw/HPxLWnww1EFuziy6d/MVQkWed43q8DjsUXvHJwewVJ8
zaDEyvAf5FZecKKq/c9RqxAx1p/+0fiRF5SSsMxwmvEChd+gE4sDX3d01C2C
eiVwfkCAm35xO9CWuJyQXR6dPZ5gA6CarmuSvwDLitMjItvkqDpM1jF1nb7N
ph+rGiogHq8NAsEO8pROSqeK7ZFHXHClBnj19NGiqJjrwU73tNeshKZxVAwi
QZAYnQtUHssHuuKjmODc7NjM0a5RS9fHRJfIfYh+aiIptRW3u6Er9CFcD/i3
Hn8DA/QDaX4p5totudbqb2zPKL8wFPPOwfjh2WTeZAJXhuiwf9uuNZ8RmSzr
TaLyDDi2a0PvCE/LZwaWCA/oK7tnG9zHGcQW531gYCon1IudwH3VNeSHEHHy
7cGtW+48qMfj1mAG8/myw/79Ehi8ZeGAh5wwMteguK68Hz1W6L1rTs6BnIEM
urNA5qJd7nr6tW4D8H3ac6ppSAuL0Klg9RASAwkM+zkFRabd31B/VrwT07Wu
+QpjhlkYLhVV2aavdcYQEE7E6pUm6SbC9Qodzc3q3OaTpOEh9sDrw8TucIhm
4WCpRYCv6X0DcRKDCsAOXOL/Hu76jwWYq60SxRfuBHBGOROp0d66DV8nfF9+
5keZYlJq9e/eM3fic8sEUCxO+GSfs9dgXM3rN77rNRFvshRoIL9ue8dgqNZk
Qc7INabc945t+i0BcLn7IEr84FdwgUdIkGoCx1RotQ3csPWAwOQDxNr5p8jH
U03yTu4Y9lycBR4qqMMi3WVC00aFhh275GCJAKSMH1OTBzSGi4/hrwUZie4E
2rcMIx0LpHmFSmNhzaNGkwecgjgTkwnqI6UhK0M/jfxJ1cwVCTLKoKcuv9Z2
wsxpKPjAPzi27iILKs5gmK8w7BJHF60IGb/x8zPDHvRqKQwxEcF0hUVujQc0
aVuNWch/rddZDaYAaoBLnIg5ibc1DAw4UKvz8P92LVKysux/nig1/p+yoY8t
wocgxx486so+kzu5Sr2F9A+RjbokqV7K5PwMCgaq9TnPuolx9VXAr8K4HL90
lk31TnswFDb1Wjgok8xlfzgqEQdMEoNHqTIjzRlnMOh2Y3pLIog8dRdvtC68
JFk+W9tX3m0jZfBjoRyXTB1OJaSSaa7xzisaZCPeW2jNaK+pimWmIDCBCxfn
NiVsHIvhejCbDcnjuUBXJKTDE+RM+jKI8ZhRLWN2XXSLy7/quDl3XgehSP7W
84skf5sC0yUQ0Qau0FEeGuD4qFIeH/0dQf0njiqR5mXjjGC+QYdbbhcBhHmk
+4PH2H5+Sup1iu47RpOpfhPoHfy8kak29Qx9DV/avhtpgBSQS1FMl+FqOTIf
m0QPri+QDdwiOuCMEU5bxFKem2rgqDZjoJJTNbJV73YUAwSU+ezAcDm5CCJe
4qQD6YsDgAmZRvfSudMd3JyFnvckmgMIPNp1zkFFhhegdVDscv7PdpAR1K7W
M6e9UI6fC54MWEavmrnlKLiIghcMK8nVu4zcnV7fQsnv8Ow2HtbRKCUCI8gX
QzElEdDzI4YktVEj5BibZzDP+Rpiye8a67YUJnaylCoEobPvgKkllj3hDVPa
yn0CyCh8WDfwFwXlf3/yRWiNq16nraIo9nvEtUf7DOhdGHdSeWFIVlO6tsTg
wDUnnItbL9/nAk0MT8bfuig5Gfqre0uD8Syht7rx2bu0zIqtbpPTc7ui7vcw
zJZ522fLkg4WSfVNmTx79XAs3dZD+5hsg8Sf1kuoJzlbroJzWaNt4ACxd2Ll
+/jkhXxLErMe+H1i5ITz4D+3XmYWDErdAuVBs/+I42ChIyEKo/q6eK9oGlPr
xX3CymrD/Qquv2o6kUdzDB/o2yt6/5gG4/GsNs+EdGxZFC+f/8ZxiQJ5dc48
wMq7I0nljP9kpCb8FXTeV3Yovyc9wYBGphVd5YR35ChgY3DTi/IiRNJKUQvn
7Yk+L//JBh3rlRoa3+7jsxFHgkgK9Xr1qiimkMdVGIcI2Wvi6PFH7PZ8prvq
QjWEHyMyOX0rSuO4epfwmV7+Gr0jBYGYlF5Pqc9fAx6nBhmbLqwI3vWolA2n
NeFhMfjvSQgUwLdKvf9F7yoy6cHKudYe21MRRdHPtU5hN3ex/KH0RStVA4sG
SdQoIHo+YoZAwmOsZyUS9olH6xIDZX2IOXbqKGU+r5DTg1uq8pSOuun5F90d
CaGmmU04gGoSeYAL8nzgWY8xLvB+qfZX3ixtVSOgfFCHPWVPdCxI9eOHv+Lg
8U1EyOh/Tued8QhS3xNooxdp2ZPVbXbVYVyzlJRs4XY+LvgiPzBb5TuKPM/K
C82707xTGvQJHftCxbh/e0mzxrwrs/803J1dEd0pYUjm6ak1cHhkJwvClHjn
Hsm+8WbaHF9n33SAnUW3D1EqdER8trzd2YMEplyBcmcrFoe6RBRKcC+08Pf2
rTnJU1wav4ivqXqmA1jOGXXAcIX8sMdJZ0P7dD/zEyePebqgz+DiHC1EpD+0
e7VVuV+9oxzQugwd89BrBNNj0eSqkA4oMFWhQ/Uwcug8nK7DVhGSnnUoh9Xr
/l5UXj9ga5/DnB7/dOBZYW78NinK2MrNOneYlYkwB1oD9XdMBhc7nLPo91sU
ioEejFU2ym3JnzdDNGG7YVjU+hupE5XFf848YCyi6BvkBJJUqg6kzt9R1UWA
zHKl29Lum5tVHoibJDbZgnAFt+xk1Ch5KBQV6Y12FMv6fZ+zd72StdvXQ/Z+
4aeI5Y9qrC0UPq/oC+4YRyqyJkG20xgta6f+zUurwgB++3xIt4vzElH08AbK
c+3tzXTunERdnvXaaCOFsx2UCjEqilzxQ/Hi/guXsphpYvsGvWpSpS41+kPh
9zRWxLqANM0hpJZfiMNKujDULbha8l9GZE/e8F9T8L1T3tb4oydVb4vg/ZWn
1tpfJJnDHHNT1Z1QdfoLbfBCko/3Y9wBygevcILSB2aBpbv7OoaOw8uCOuLf
lsDGUrK0ZgPpkBRhpl/myVD+zbpljceuQbmHnrFf4+q6prdyl9/Zn3BAAsX/
h9acMIDJkCYmxWkErayOFnC3onY7oPSvJ+Iw/PpVGT/pSQpuxukLEugm45fp
VJCi6U3vaiSxYIq493ASnrdgxpuRR78hPPION941zgUWuwDFv5bAVkXQGwOi
lwPns0cpHXAXrE541LGO0YU6hqYTZEZXSE1wE/4u7nViiftmJKCOKRcqfe3x
/W3OxJaZNruSwt70sIbGs+iEnNY0YX2yUNor4IHamHmS8GRBgscxy2cYz+a2
5A5Sl5RTR7JWPgwakC4NcVu6wy0MmuLZ/JCAFOz4OU0MjntWef+32NmSS62G
HKCVFcA4UDNPWn05n7Vfpi22Fej0uCs3hXJRq5tMExBKrDj9FghUFRJ2+Wx5
YA4YgugtHF3PpTnGuiD5nhbPFHjM/nFWZG78KROZ91ZyYykmAKYARoEAlpPO
8OzKSACfVir0ByyQY+8lyCL3iXnItOkg1OIGU5PXbw3w4l7k6ni7j3VeaIOc
/HuC5pNRQvRvB8p5dLoChJetHr1Hr7QP36mfOw5mWtPsGHVM6YzwigECdmDq
B1T3NCu0V4oEHxfx7qnZghgWmWKJ6IXtqaL4zh2+ZFLdjwzX2Nh4V5J+AtJ1
L6G6RA0WCXw2ZYj8R6QSjJwfCh93YZvDeEGIVLTaosFp5ILBqMFE/BtwZreC
LhunZfy6lJTxhuu6TJ7gddiqHpL13KRkcK5/y0QYaUNRN7xKHZ7lY3vZR4b+
0DL31goj0/6K4Q3XTxcvSnqamkT+BANp/OYt0Z8TWoHOTGfeeVlybIa+/31R
LIPRya6JYGrrjDJu+3uDffkWb9xGfWEc/tGoa4a8BWHuP5/p7Be0G6EonHDX
x00CXsBj19t6n/1qk8+5GYZ+G1hTMXatt47pOk+aMDVvlpeuHyiPmtprbhLH
ZCct9dVSEGx/M9vL7CgqbqktGPSHpxV1g2VxuyWOt3lR4tOXK4mZEvYYlZGT
/GvfL2wqWjJebYg9tGFyEsLRIPyKhsOSO2lgIJeGS5dTMAmTe2Tk9r5JR4dw
Xan76/CSMk4kqo1MYrp+CQ6TFQ03gxq3t/qOSyi0hLpCorY253ItUs1/9bqs
j2reSeL/sEuUqAB06KwDogb4ovqt4EustS+8U35Disoyvsrq+KcGWKpZjEyH
L0TaIJ82VFX+83Jw5+0WA/uwvLeLrqBZ2TjgWaoKL+L2d1GA0bq+Yn/3S/HI
nreCUxVh04NGlns9GEqfAwLcES0TZ8OqqW8lvWBiFepxNRfZVSn+gJnn9TP8
YkRfZGpPtNoyeIDmxl18za82h/RgLIP1sOw1C7EOt0P1GRR9NizOZGFe2OX+
mGe4RQfbzI37JF+ix9BgvvG7uq1U0J6mBn1jVgAnFcZ9MGXZJtGi/jp4B/9d
qrDKZ4FNlGIIffXoXR4AaWCJaCfEXtjmD4AnLn/bcMKetnefcAFpsNeLnA9b
7oua8YfCO0ImtTbvCMsF+x/e7ml2WU5189RW2Ixz7224d61Ivv9joBFJ8fls
Regvg50pO18vV1yHE+OelK1Je0xd8QM1zpKKGOdJY72+8KH3AUWpv6WSLOmS
p0n8zbWdpHsd27ca/ybo9QmA0LP8FFG6+ytwKzoy8teGzPVhB14Mj8q9fIzt
JPD63MqUUVncxDDuwYAXSWjzUTNMGuAHNK0uaDZQhha9Z45XaGlQRtFiQIPB
9kJ0cwyzrA5vSfNdzm7+KKd4HxTMeyuGe3qiYE6YzipX2fOaiprfEQCZoL0O
OOc3Ls+WoIQQoo2viASC7lo5ewvbcg+4foXuRlLtabFo03DVW9LhTfSrqbvl
SV77pNd2/UVRxK+MbWx4FbZaOIQsh4J305QUeA9maYVp2E5B5QhgoDdRQcIg
L3G/E4b/PvuWdBWw5At7LoXEMKp4wCdFEIFtH0LWpRHM8msqu6ufASbnKY+F
Kbw6re0EzDiDS1gH53hYCa7ltFOn3aJPMq+LOl2fBdbT31f6l9uTW0paypn1
ux2m4xywmRWfT13CflY5jglaJjsGrg01r83XARJX1xdDDGbTWNNfHWzyR0kh
vGkm/jnuSyiyqFaSO4B00Ggq0Tw0cK9Eptji7obxPFu2XDVFRe80Y6Us6J6C
lODKRicqFg2j2M3qDMdWeCDlW3htMTgQ0j2h1bEp4NPjniTvX61kVEVG/JhK
NWmOCm4pxgQ5GprcKBIQ2BimE+lR3gYaXtNzwrc6Utqv9vsB4iHhcqSDBhBh
qLqoLDAaizb0Vrw1dcdqqtOAP6Jmqghk8BgDwCY/MDBqDWJ+xna0ta2YKkux
RtecJY4gQwWM2leHzhBtHbZ+Sg80r65F6ZrDvGYNRoS2rkBjBVrjdtnOcsRH
6f2bW2EXVeaQUcZd9OTMqmvW8w0xfSXvLWPV3lLMSD7WIcqMz238wWpYmjRr
y6ehmkcCRr2vEzGuU/GT0PNM8uK/KipwoBcFCIlG/X/aTxOJrBDgpZ4wAqjg
DFA3LFGYKQz6+FR1KlJl/8KGYt3mbAkOnKS6QGk0pXbSqf0FUbcfMwIE6WgY
HXeblZOlXe63dDFTcJaMEzq7U5MD4/XJNf8UR8VH9dvwmIFQOddActX8ZPzL
0J7DQ6MJSdOEi6XZypgwVkosUPcBp7ecHGzMFCG+GxBqODovBWl1W3dx98aH
E6TPBrcDKXypwjUGGosHKwXJJJ2VAt6GzFyCOtN2wgu2uYvyzDjtyy3nch+w
+ETw+VQjbh09+Aa4/dXurEJuhIoizRkCtugjaqNA3qV/ajhJ+JaObUtOAKRk
zHV6fZBgLHoLegYgfRalG7FIHFm38TF22LtGwsM1VAHorVe5RnMu4KLQLnnP
NvI7SyFOWNMxjnr+Ypx4AhSElh5vVVrQipXxto5GVRgdjVn5tyfzFXaGbb/E
0v6CCpn9oiezaqnZkEQF3xT8nK4tN2BhwiRZkz7UxOITinBEIemIECKr1lcn
ZQVjaTcD2MomsBqKAXu07VQH+Wdq22EhVMeAygWNTR3uasidW36fd4OrhFzJ
H0oK6XgTfxUbnvCa3hyhJLOMw5V6N8a9MNWNkUx/g0yc13CEMM4eKogsnlh9
HWIf1S7WcAG7J8LHvHWan5mc3A+N2DFZ7ekx54muFxgNqfAdV4X+S0uYGase
86GuPmebPOvuweGfL7tk/shieDcBHmTW4NjkSIBv9GHr41FfDF/lOag/qFof
BEPMHFdWR5CYvM4++zZfQbBwaYYDE0CXvX/nPpjrmtBQmcsAAPT9BsRW3JUK
Ofi0dBs19EqxQAN7nvPMENOuRR2Z0lOiBq93vnYoF+83SqA966JNg/cbdgUE
MrTAqW8JGUsMDJPdkUvLDUlv4erbgEt+Y9prwY73EICF5ydwVKYmXb4tdh0D
nxWAak/BqpaT2aDPdUKfGsMrWhDMLFdVwBmAKaRL6+52Sw+4zs+FbXgGMiYr
thNlnGkuAWqO3ZkKMq4MmqzbK9wCxImozy5WEipiv/X9XckrvQLBRnCUQFvI
DchZpVy2djgFMDN8j6KkmhPL5uXtXYMm4SmE/V8KAM826hDpRCV/KvVllQOC
E8mzLFVjIan6JtAtxO+EuXn3v8HtDrAhASDt1GOj/673UR5OfN1PrAjyElOY
s/MD87PQ+T5NFA5ingA0MxdDtY3KE1Z8jiE2cThM+kBLlf0Dm/PPajkZhMPQ
jjlY/5jtTSlYI7XBFskNiS2HhOzkLneAKS5VR6GRvpF86u4uiUatpjVJE1Pq
UUduoY3YAWZdlH2yKxj8bdOIV+fROX3TgBB70+DZNBy45HXnJNANIe9+Mz/k
xi7dMDBfz/CHIFZtB+FwXf+qQobuCf8lPg6tUP+c/rcrV1ue25M1cBY4v4Sg
YNYVLlbUiKrs0Xr7t9oR+tL3Ge976O89JJIUmCEGa6vNIGF6wPVMdMgnbo63
+zz/jxI4CKOaVy1zsnrtzSl56Zrmxcz/9EItwqHSKxKc5FizCGIXDtwlGMXT
CyuQEhhtAQt1GWoTywHS71jmN1eGZPB8hqLcv4b1bXs+bw5p3L/UQk9LUEZB
Zs6BNDydMa95ellCBAndjk4Noxj8cvxB0BXH3gSZhaGmWoKJLVLX6CcqqLUt
Om6CdOwP3/ZsqPbDSABR+w/MMT7F9G1B2PS35GyR9EKOqrMIlgVY4/Dc1u2M
h5+Q5PZL7IOPGaK+vdEJEcuBAcNVFJTHUYXNc/jPZ/c3ebVNdz/Qj3Vv8Yfv
j8xdo7TghkhKzzlBqQKbRjCRcj9/l+/CUF8F8+JKEmKX4inMk8goVfSD0NhF
H+5ab2JKe8VTsT7b/4kyVtJuugiqw16KPdk3+pIeizSBBy0WpQVcDsupMosw
eldavKtl20WumiQvtJYq1Ae4ZeUb/bPDteobZ7xKr6qGDiLOH1i6usY9+p/r
k0D0bgl6QmqIv0VlC1Eqtog5V9DhShx/0EjZIWwiLlpPQkSy+RcJdz5m7ZGk
LwiZOux5epDIKiHr5Gdw9VbSqeefxBo+122XP9ZGAkGJYnsutIxpPHIt0eqn
3+RtGwJPCD+NEzQZXNIB4fkUKlIbx8yGD2UFY+le82WEpeIOgp/U0Ct0FA23
ng3avOZeSVM66GAOVw80EA1Dathza7o2JoMAx0ieDGn3ZqrafLcZccz5Ig/B
W1Uhq8lHlQb65jZT93o52IFR9RKTDc3d84N0nALUYBA6k59ocKC4DbIzKaCc
CAHLsnjnmyrrmEEXMpVoDcq4Jz+dC8YMVo88b6ht8PmPYenTKSUfL+gSiYIO
8VWH+Ch+YzLRbfahBwkfq2FBKXoRi3Io9h6PeCOm7CTmUQoX4gD4FgCAnum+
5YmsIkpXwXvygg7w8knelrqbXUE9W7zlZxeckGIhHlb5SdMM6ww7T+7zGNWx
0/YrZSzX0YiTYjMZKOsrkslzanMR6YN5507ANRGC60+82ee62wKaDOoH331e
WmZyjBMNJJ6lbCrZ3+6wwQiDzjqS2St6FRCOfENp3My7PGC7UYoxaznJDVre
Dp6ZovNYVu49CRAgHBrNeucdnnLRbsQmJq6L7FJr2v2Q4h2zgW9fWh8aFrc6
989Wc4IMynVQTEjr0So9gppUOYg7novILeuVpNj1KlT34ubKnNteoKPS4t/s
ov9/4ynZU9AbJX+fd7Qw0sLwH8qzcgUquXellTlpJM7M65xau9sK4VGk+cJE
Cgay2SOwGMtNk551Xd8Ogs7xg1b9C3PboxyUq7BBZmpxyJ0E+9aSXwti6kJY
4N7bPvEWDxvkBng7oOxKdSjjHXwzdP6VfZwoB9BOBisQcEqyk94YtMepV8ed
FUUcArR6yRot3BquhlxusT8RDfpll629sk3HHVffoRzEr7Svzf+k1sYy9A7p
wIbA7kiI4fdjZ8lQg6VKivieQ9WMjrCTF2hYcVrGMtpDUrgXADabgM47VEmg
EPYgk+V9fB9q7eenEOyQ3ytUhIXm8MsRs/UzfBm4W5uoOxqQ9dXjSOVGZWBI
46lbns6D+p/gVafv+4f7oj7/1YESGE8B3GAWl+m0JjT+RzFB0O4D2dsurOU6
Fz92Q60nZoZSrNyIQPWRpXZZgWE4YkPa4gxDF66yuFtDwXihH6P5Q06OCmls
XXbzCsQ89BC6HTgnhrsor+xZozQZP1tZXynG6/8JZ+aDZ+Jki7xYq8jgezGX
dQ2owe0igySLV/z4R9CMZ7uhNQrlPpWoxa4PB1dPUueSxdPPOlKnFTkRzpWi
Z+LS1TVEbeXpB+DXFgT+oBDW0iOaUdr8nz7M+dPHsbXOsvPDkuOzv9MzhIWY
Myt+r/RaU8HQDEtuZOk8XjGPYasjoSOFxnDZr/Rb+27ho8S+RhX+rKRsCBRq
OwPHaZsai0gSIR2h0NHIevVM9H24v+AoCIbwhsfHJyQnv/styDnDA07ta823
1Ccec4N8dWZz6gPgsKe4A51POVUPcGtWB/LXlKAnCEeU3D5BbZWwi9s/YhU6
ltWl0s8N+7TLRo0Xdi++YheJAhOrmJfCGrX3AuYGKVVNSKbvKrxlhsAJPEhk
EyQDXraKrt1/KiB2nk/JC9gUkvPfGjE9vruliFMDR0eyasrX7+QZu9vplzNb
kXjH6GHFjeC1cMf32Cb4vdK+lbFJKfqVdThySFwuMRHgeT7tyfr9fOD6JQtQ
oo4I++2b2C0k3B3wHb5she6QKDqRcBclqWQGmSQCNAyBBiqPTaB3mrbXr/qW
6l/kW5OBLTJpT0Ski18vQmaZXWzwbKXiI02H9ARJRg0OPXRomieAWv/jjAyl
UDLqDyZUQHIa1OR84+CXXsC/FQPinCJOpz4Z78uLwJvNdlAfyFurtuCZ36Y6
gD7b7qgMkcR7u+P0sJf0mCofAp4jsne+T8v8Wn6xbUluEK7QX+NDWon4479k
VDwncdAy/9lI4u02YajTaWJjEC11NBMefRm0Vtrok06o7BD6T6ySon60sQ8U
24hH1lZR5RKQz/Kmvw6hHbolm+Bcjq47dVtD+0oopSOrPf2/wsTsBgYHvY4z
5vYwVvQeK0/13/RTUKENDnhRkpVWS/+saLygrSoN689pXhxAQ8TSXQJ+NVPL
Oxt1lMFQ5b3k+k5Z8/LHnN7dAMm2JMf8eZop+Wt+IiPHcYxAYrUSjGpqeHx2
ZDnKnBiYiBAwCR3XyhHoj/UwK20GE0vw3w0lUuKivuIS0+kiXUCULPTBUMZS
fpomL9G9ehfvM5odWWe922x/fxriOVfvlXOT7+smcHizUY4zGhfZ0Oh1ZBDV
ypY/AQXWJ48CMAM3je53Pt9x2vRRrzFcsl+6JgAFMF/yFnQPIqhw/Rpr0asQ
GKbqXXMCtPv3rjpEgwb1iSv/NAl2ScPiD6yFn+q9Axm7h7K7RxHHUfYtxW8u
HouHjFPC/wDAWTYYoxr4qF84xE0wKA0M/4RWSBYL14w/2LnKe55YvSkQB4JH
6kPwxqGh5ZzNQgT3sFGeMKsfS/hDsjznEeNJ8k8afPb05fnONsbgkjCMMjRd
thEcU3WkeN+YEYU3a+3JVn4i9ivfMk3k86sR245oICeKyOeETIZtEyPFq06x
Ko8sT/cwUbdpNkKHq9E81PFHp6+GxiyZ2Y1c/A6dkGJTxQcV+jaRl2cCwQC/
+hVUmirazIgoUYBPjv3ukQ2dkyUNfVSONBqzEKx6RkmgJtMtyLl5HRIQQVj0
FyzaJqJJFWht+PQK9LmFoRl9xrYAi/GqeAdn9Rhrd7y/JVeY9Maf+AOfqBV5
+6i1SpZRpLK88I+nl8NEN7OL7gdsUDdRZA5C04hqke+M6pGX0fsxOcm4seu3
UBkmXqXCPQUp0dK80vhbbuMktZbr0jt+sWwh9sNbkltuu2WBUh1DsC/JI3nn
H5I0j7t5pORBOgv3u3wzK2Y73nXCWyhbGFHoCSQVwq7S/4azLY6TIWKA7SF+
Bg56MDUA5Kz1bw/esYwOKEruk/4WKm2k2FT9jOmkfo24nU/rsk8nQAijc3hJ
hZ9Ac6gHi9IU0DLkxTAsF8TrNutrgNDsBk00kWF9LybTjvsrBSzIDDijze7y
Ecx5N9ycoTtgZCRdIxPRzkCVwWmV7cLfa3SNhyv3mk7kJsS5ADD6yW3f3dzj
0HiHWvZp+qK/tzpQvWOoJw8auYPCduakOl07ZHi+IdvVdgv8Db41PbsmH2L0
EetIkXDx2+o6hNFIISNsZhjHznqL2av+nsPhivrry7r2DUcsfEbgAhQVzNWT
FvNYvQsRTOR+GsnKsZlq7eFGxQ9qBSg1y+3cmKZDoT1V2FIxYZ/zq3sHPsRY
ssQxInatj3QLVueWWBEiiZ3uK1A+3khV8Ws7DXFbUo+Lcl2FZuGkmqwmJUUc
yLXUhUTIVboJaaumuCAwofB+CsUGXchIAiU+UchWlnq+rasIbIrj5KuekcHa
TukbCqbcSS87yiUuQyeVRM0yLa71Xd+fRyJq6Ir73F1cBssARPwRr9/rYHrE
s1M3W19gd8/L858UBaT991Hatt0PXu7880lpWuOnCduk+8y4V6Nz8BiJC0EZ
ZCkuKOZofBCORHI3NFJDFqpuqEPI1ERmjEEKnKe5sQLX1EoENcXaS4omOqg8
FQJleQ6m5k7YwyUMjy5BOnxtrTgXMkJwOfZQQLUZg+hWeY8uaJcyFD2Sq7gp
sYjqYfPiXWiSQiTBDMGDro7HXwD+Hv+g0a1yeu7m1pJ7R6+X33EV7myy8ttu
OBsMtfcvidWPPeF0gtqptAPtwBV1ngY4VTjE8oP0LaJEZDFNxljSMNGcih6z
nb10pARVvjamX4pVjiYVd6p0dJqcYcXPGwCzDGYlZC9gS41uVJqj2eUKIljv
JOoyUDtjWB52/Jw2Lzb9lFCdItI0FkazXwKssiroVYVbzkBHuLpij2j0ublG
8LJUp6ZDhlYiH0lDvEtfkj5M/iH/8iXCFKQ8gFWMe2sDN3o9uwqWqsPT1dsT
dThzq1ESfygeqrf8HJ4KQ8KfFBYc0x17Xrg8S9G23hY/B98tD+/d+2zsYMPY
blbRuKECk1eywguwIsoYQnWba7ByJgjAUIvcm4xUxBRTWVtQVXBFxgdRGHPl
GfjLt/jF4NFQ8PEj+Ix0HppeGknfy5LqYF/o808Ml20dyYGv74fK4T4D7dS8
Xfn90VIQamQSlZ6y+YJ9xnGFY2OYQYB+JXgsRNogxhF3HcPNnzOqSyAliOct
UMv6GJL4s5envl4/QyWIXGtg5kIe63CpXEAlIYMBehXUzMOfNYVn/UZOI8xY
1rb/7PMOLPPM6XCQQxW/C4vVeYzeNOHkEhGHw71YXTDPrQt1QtptLjMGkV9I
S6hten+899t1pySN8oi32gW/FBQnUSl8+HrisiyotrgY/DJHFG4+OlTQnPpW
NIgwVP4SqSQlFP3DuyUIKK0JqwkdDnc66JXKYxK1xqquP5sVsLVDuOJJeSm4
6948n7fsZ8H4E++I8902MaN1ckB7Rjm1IKRWBqt5PAqwVJkM1HOUf+tIhIQo
7hKrEKGgn5Mjov7E6uwcUPwH1LwhZgyg1Wc5iRJ7V++k03DNtoekrEo8sRA4
cLCJfqcC8arpgm0ttwJwNWPVe8oPvfiEOY/pmOaWMPrNO1xhIiWoA7mNZ59f
SbpNf1arEsHlcy0lEeHXj8Ird6Gvf+GD5DEPQb4F3EZ9mUutm1LcPHVes2Mo
ZzpZW+zh+6vCGkMBsREW5CuqH9GxIP9/qqcCbATdSp/HydPcGbWJmxvuX0kp
oUoKY9yKRU8EtQXqu0GcPNkepMpccMp7nP5GhTh63NJxndMGUEHZC1sFuqjE
HTlP6z3viyIIruU+w3ezAert9JlEQSlHXbW3vQdqLKp8HJfekLfETQMM2ILE
fyc6PRrOIWZv1oLA0lYMBJcLfKAWBLZkpobQN5S2CypSKCO1jseXMewcTUGF
hzJ4gstb75E5Aga8dEvC7M1qE9Qn8B1P8Lee9hINews/0C1Qe4B/G7rLlX8G
9e9T+9e5dJkCHXRFXgbp7LXofPAyY/kT9kVSe9MsnEHbFPM43FfPcMzSS8Tz
CZHeCFA1kkPcM7xGmPT5bg8LdPLOfW0aqG1/YlHSVtRejuBkUeuzB71g5Npx
a/+V/CWQmfWz9C/0sm7f6BVCv2PgF43jVgyzrT8gDo4yJ0q4XVurjYlDoNhd
Sv4z5hrPB2+C8tXR1JOiLD6AggrDtAx1CEIiFVZh/bUbdVH3M5GUPnVQ6vh2
BDisgx5kOFwYSAyhTT0TlOOMG2t3LeX3vJ6TGM68BFL1rhewOcmIorTojmWI
8kX3JXbLyXQ6teVMcw1HSWBy2JqVt/PaQv37RPt7RyVqJraNE4Thet6XoT8x
3h218txfRo4DaNfYfymzDcZWbE3159DgM02vxtQMhPKSHQlWZ2rLTHFg0kfb
kj7jq2qo6voDsCo0BziTCzLKFst4fZQ8AdqKyTp1MD4umnd0mcXwwVgLDMjp
JXtbGl+7e5HAS3+l+TSIS0iXev/+FWiQMSy0cXmdRJwsmXT4/1Yd62yBK6xp
CSttXcv0p0yuYoN4YaxsfxiRGpIEeD2uz0LHp3HlnkafhuZD9FJctj4UVcnV
xy+VtbLzepXQ0WoNMCRHVOHrK41m4DIUVexIKyMZuYFbf+L/B+8hKtIFj5si
lKODnjusu9k6Oa01R2dI3ZyrVaRqJrUZa/d8i1sMWKg6/k2TYdiASVloSDe3
qLPuhySc3T3mpKhPHsn7tGJ3oK9vkuCrteySEalw7sptvsiyZZ8FMTlQVaql
DB4UjK1MpSmCCmrVQWEjfP8A+kS+aOF8xup73gOdBm44g9PGeQHSxLcXwdqQ
EXOnRVsG+kXLi3Ih1OHUvS7QZXYGv38K9yr95wD9D0rkaoQemrES91T8qOin
GeEoXSWE14cqzc5J+5AxXbtfr31LOOxnHicysA7HwAAnv/2EQSGPoieYoJE5
uEBMQiEIn/5d9p1ssU8NwvBSmzVV6uPwtkYWTtsaFxkE2laTinQy0Foua9LZ
00nBijYWA93ttkTeBPcPd1BqP61aBgZy/L/hTOuspf+Pzpq5uDUVHpTUDk57
oxIgXF/uAUBAw/l08QESe76SWY9/rOEASgb2EKiqp15mvT99E2Rfsk/b6Wer
ORHISDjVDpbjfJmS9WwCf8LaNAQj2+zY+GQU9FNrqMADdFKLDMznCErNoEO0
p/oucaVfcil4npGKjZfNpVFuwc761varTpqvepTTItEeodI+Gzz8II9+L0la
yerVmCbX6RaI02PdoiJfotEPsy4/iH5SQcC+fCOP6I56iH3Y/TnCUMl5oqb+
BYw/fHmJQ3zLJ8uwBA8mXs3+s5kCl05FKgD91+zh/K+ceT/NL1kvvFWIzP+A
eItaIsK+gQpOftW+gN9B2eurS1eTu9+jO/hZIYDYdyFdZW7HWV5SK8SCbUWe
bVFt3O2Sd7hpRNMlWu/roZz/j6lgIghnzEXDgwmxNrpR0lydZWko9aaz3o6e
2SMgeJ0BZjHgNSsdNUKLaKNQgFAuP+no+5i4OHpuzWEVinaHjMCCpqRgf1uA
9GIsAHXFBQVxh+WAIca+M3uHvIcIsxw7xJ7RJEk4FpQgs2cwS9D4mGWquGad
AUW5QbNpDXTyYTm3krWFHijiRcw/RX8zhP9/er+10txqAlnabPS1RNmxndfX
BRdlns6xqU5I3xcZyhTVk/5hEv6Q+eEvJDrZ1d+mrtbVIpVuh9neJTdOZJGD
GMQrojIa9Z/17OJeOvA9psEOupq6UZ2cFEhwGAN94IA8D0wgbegqdZ8UN4co
fhNTxWfWMV1rIlECeastlXfz13bVS3b2VIR9E1bHOEeN0LpHPgeVDCs922JP
klUgdI3X45OUDeklvz++S8DTezRPXxNXTBnUEz2gDqXOo8pCuSE/dlDgtyjm
5794C0BwSENJ5uhHIt1Bh1d5JHVjBi6jgPEaPvdTKJUcTshSQ+ZxS4y3njOg
1TrE0lBy2bm4m/4g2NRL449/8s8KjeWKaCShqYsbIszeIUAGGPiKhZNzy5IM
dNUGmJ+YKAXCZBUz0rjzUjQ+NfcLoOhmuoHRr5g6Jz1WjAFsKJ9sb/pPM00V
AO4oyo9Ko9IhoalI8GQ7LD5Y4MgcHvGmSqFDKBmj5aX9YbhwmCcZ9uQNHDP8
6OCqjoFDrgd7YNpTWt1sh4e0B78lXInTUn0cQwcpKMrL+KZaebyDL+fH+BIT
/mcOHGPkV20JLNX/JHEHzFEd5AqlHgaaSmo85IledwlXKq1Rz/Me4EKR9Xcf
5XuPhpeTzQSZdpDRZWCF0tsiGPKrRkeNUBOTn+eC8kKng6yyIX3wqORLteGZ
+D6iy5lP4N1Cr5RpCjUjv4bISpNbi4QowY0YSVw/0580QtH3WkYmu9sfIG53
E/ell+5dakmOl/cJmVtFCSfxn3HFh6le15ojrfNCXn0jejVZNxmgmYn1uAkT
FW4AygMsNSu02VPJI09yVu/rC1ZqgbGzfRZBX9xhqEQSR+JzxlK7mq6aVmo5
tmYELxHySYzgpeVgB++358vWS1Y12KXUo6/PIhtKwroW+gia6jdAE4AdXRBQ
7IUJw0bA0zPAeSdQi06ccrvXdNg7po4kYmRRWgiqPbj1HSRrH7ef+oL70pC5
bUm32Rlvz62HVaqR/ohxPQKmgWg9axVWwmw9yi7hsNbwWibKdAha+xMXu/dV
X2vTl0+2yfWpHfsIU2U26pZJsiwJ6Dx7N0pU+cBcioNcbMaSk7UJVzZTsN0A
1v0SgZ1eFl1uRV4NFzbxKd5YfdLJ9NRGd8nkxAYxF0fT2jKlciVzwmWwtoiP
FvcEBPW8wtF2fT+XfHffZll4HGCW9P+dGIiDu870bPEFIkQGIiTnR6EaKAd0
GZ4UL5AsMqVhY4bIxmnLxTKj+vFDzyHFH9uDlorJKKViAvSvFX4mMrF7DlNT
CCYthE74y/fyjDnAntCCv20f+4UxsaZCQV4pgdScoGCL6ki93byBYyGeJK0z
KgyXErmdC1kck7cxHqmlG7JJlHTQM9i3qnPIDGUUEv7KUMWt5LsmNnzwFiV6
/zR+L5dELRR2R4YY/fVpGKezJk5nrc83MRa457uyNtdQHJoF7X0H8mMgbRyx
WPc88WAWf9xfnpjXzvM5gLrt0SiJFTBcyZ58vsTBZ/13UkC3nqjuAOafVn2d
XcmX2etfT9YHy9UQ8dTEuuo6luGJO+vsMMo4+O++NB4+LABWl7WvGyLP1xIT
kVHnE4KHZteF2sK8S2xRrGwjklfvdn1Wy7dXUdjYmEwH4FyLIpUVd2Qs2a1N
HRVowuvK5IJ9vjw7wqJU5hKBBfJL+YfOtsE5NDQdfPOOIqCJterQOnijwHaV
Q4Y2sqMFDp/AQqZTTJw7ndIejZRgMKgQ2zaKI5yNkHLowfPHwIbHyX2PmVyQ
BHfNe+jAlYrM6AAjIzyiMQtGDBZRr+CQEDzvTWQzAikgB6wdpHzQy8GVa7sD
iciOQ6Mj+Se2aMZVbOcrdkJ+5LdTExUYCMSwWCmOIdsUQEP1m5IFg4gInFoB
hEylMxDj/iYsHqee5EE/lTWU4ny3Dsn4T7c6Ph4QyaDLk17X6iyD9uMuQa70
SHkO7ZkfsAQR3sYHzv1n3Bs6Ly4owWK8Df3U4YoP+dylCJXtc6+bv8ML96jL
o9JkFm1KbZzDWxhEoPwPHEXmk3vEQ38YR5l2sVIMRtseKwKeJLsyKAIx5sE1
fZt6MEXtb5HtiewFYOx8XB+ROLFqIXQXi7JuLgMAb/zNqWbbacWY819/P8Nk
uP6FImr6S7wHawrMWCdcC9J8sLJCwNKARmLMZR/Hz7mA/3gTCgfhC6Yslpel
vb+vAk/yS4cjK5bTwBGDgukySrBKxt0Yq0AxPcwlv+rrgfLyVPY+iWKDvBux
fQgUkE9KRuivt6xTJIMmAzaidb9VYAmAMGOETFZYVm1xzJPX1KHCBi6WdeQr
Lzapi+Dk+NzGlJg+t2zQbR9ek9BuLoV9p+LeGHRU9ZumhAN+jo4LbDwrFDVp
WRJ3enqZw0mQro7bsYBAVnkwyFwSd+ZFe5/Fg19Ec8OXuLGsRpDJ42fHQOO0
19P8iqHipvdk3TfxhDfh3uHt8yQnKdKeNoKnpHJfxehrJBEFUQYCBqIRMXbC
5bG7ix7IN6MO+wf9nz+geJZZg8lynQ1ucWPJluGAFP/OyHlGzKM6Hc+eexGj
GBG8xtHUQFElO5xyPzDzjQvzphUnWIktgwWVHLMg6z4hiA20otCm6hlkpPV8
AyTLWy/YCRXCZ0+sj7JMhqGezbZXYSR+kTzJIMAmDcWGDdmmT52RSWR4prAb
qa/ZvQSjKYFzUiTTaf5b9uPp/YqF8p89xtG5U5fKwCMJOWZJX+QUijLndW6z
TpV9j1SCaRgR4hkxF5DmyYezN4V9K9LU271WlGatl5Ou0WNNZrSbpRfXoOld
fHoN16ibnQxgeOm8fnjY9EFXmEi670/ufzslZaNeL8a0rnVEuVU6R6bLs68E
U3ASjaXPdcAPJD+S+VygPg6DSN0NR/JfQOXPYjl4ZnEB0aiMKIZo/qKMoCvT
utYdDju8Mq5hEwX9dMlRmcjyPNc97+2PpscTF0mOoUFPOqDgLw4UOK4EbUGg
Hro1KNASrVekUxrE1Cr4AtqeSA6i7drrovk3vymwPcDhXhlfxOE+X3Zijk4l
q9RS3XsRtpyd8/ve4LBYoQ3kN6QzxGDMf2PQWAFKJH8FVOj+1g6NGLyiqQUR
/naCfo5F8x1FD746M3A4TYShmIB37ZZV4sMS1+K0+nGDXnVBoDm6hGmpBL6Q
IkBuUA/m615d9oV/4zGGIyE4lX6J1hTyz++H1r4u+Gsus7Iljk0Kc01v+ikO
swF+0R4HS+/VkMzJD08Q/dnTLgpPe8lvUgpJFAewB4q9QyRtGvuYsm904bZW
cB4gATcPcLdpAuLgxi9uu259ruoG3pMJ3bXLWBkLLq5LXYw4dKq5atHb4GUQ
4vGj9cw5lOaB8Um5YcC8btjhIL0GrG6kALL95+LnbQWZoz//Jd9I7ZkRd8yi
kW/gNzfoc+Gn6PH9YHnqHH5nMf0+BWglLCgIT6Nn4waxx8apx48FY95tHGtw
B+ELnyvc5YG7uDgdPwOs4DA0nNkb2CUp4aZ2PCqRf44Rj/8f01GWAUFQbaRG
DlvMyJfUsgSwu6t7euToAflorGJSOEsD/w8CHufvyuAsIWU/WtbUnteEsC7M
WqP8GdVkfmpUr1Q3DWnyqj7Ig2Mz0uavwECO8rH5j2+KNUbRY+Ez3ftt2RR+
U0vU0SW+Bfx0Uk4LutOFXXvgrsbvwzCjKvuBwt6urZjpme6y//62xjHRwtJP
k3K4xp4P9NPd0XFPybVLyFXebKJUMYWjPWQBBFTVS0gdeNYjv+t4LwCEHQ5G
0/DONnHGb74rkTEZjx4L9m8nrViwi541P0113800LImDLtfH0t5kGL5L+YoA
N1cMvz8ra3ROfXL692/4u0sJhjY5Ljqpc7YgdPbsjrLLRKHdpTwioAyuJ2Sc
SyXz7TJJ0UsN0VS6YmatJ2rTSfMBjzi5kQ+DLavxR6MkJl+YRshrCKOT/5mu
MFUW/L39p2KdutiUvPDlV5h2bLXg/iSBRSAaPuqJohnI8SKdYH7/dfKpZeHu
aDF65nPIotuhjzuee4KKgTltwR4+/D/TH5Aqp/0G3IlhreifqLke7mLCGsIH
t6gIcjaoj96iNuYTEX/Rm7S9NWK07AccEryNOSRRHAGu6ZNhx40/FMlDBdgM
H9b9L7ztDKWo4GfqU7uDCTE6uxnDtgINQSB7IIU7jNUXVzuv4aRmX+x+lsCQ
xR1Tn7vwl7sEKMNmbA3nF7xFm4yyho+jjA+7XfSBp6NkfHG2pg2zMUznhuWx
UTMPQYdV6jMLfBFA95q5TmoUiZl1wPCiBhtam/CPjNv0kE1mecEe0CXukL5U
UKVP/BLNbqNLgMSIsZtztJ1lxWIegZ9DOJDClpjibHRjaK3PJ+KND8Q25G/W
Y2Cth2bo72xO6yR1WkYXsZFZ+R7rITS/v9PCLj+Y1RoQR7RU39RlfM//t0dW
5L/a2n0gp0oKI2MVDv49N418mFCHsOeFhNNnpJMx/0AO3X90lRTU+Zq+B4Nc
JurTfis5RTDDLxAFAJBn2AADXo45CvOXDVqB399rqSN8ffST1zc/QlJN8WXk
vlX7G7nGaDunpjzmg/FM3brmQg5oRFdWeTYIeUS5WuT7Sr+gCzq2aa5RJXdj
tFiyN0FnNUi6k2xpA+5EPW3b/Vz32r2WsIhzvRNVFUpgUA7x47i37NPDohR6
Y0GiJkoIPmG+rWX+DxkuiTsMDGohigXJ6j1hcQcM1STwG5+oGDQfrLiMSYk4
LFk0wf3SjGDEWpgqCY6RvONTFWFquGEM+65jfFOqNp3mHojqP1EcOe0PNerL
GLk6boBpMuA7aGOba9dn7/40uIC/LnjocPhum3yNhwPUCmwQta7p1uFdjPEf
EZuXy2rWp7xrX3p5v+y28OZAvtWJaOx/j6BwI+7g+LKkSteGqD9lrNxurvTt
LjG/XsCHoda9rY58z79wGDLS+kbzxNf+f35g8ZjhQmKZDFGiz7UtpxoT65mW
cexGZmt+D8o+CvA5Lec9gGnfEOK4QpjD+FdILsoUiaHJrEIUUlbdQKqpWBun
6pP214t1EqrIeEcnk+RxLStbmxVZ4FGiUteTaKjiKBnJzPyxALpS21xwuu8b
YPPndWA568mtfas+FCOKwksc6heNw5IIFtquvgSIDd5piRF4RMNWzrFNja3N
ExSetkba9ieJZsb5mMtJtr0BT1CmRcvi63X3L4Shg6+arBLGZLTnJYzmWfhV
7Ceta/7s1lcItFrFMjy1pFdKGEmDvYVSdRdvz3mHzdf7qLmiz7oW6t16EZ8y
k35juuP8yjYWUsSFChp625+zdR3gyGy3m9WH8IklGDIRjDZJMLO97rjBhLw+
PmJyzP5de5xzLoLlbHMQTmsa8OilKsFWL22KTJdAY6MQWzzW1R/4TySz7EGR
F7XAI/VoyuF4GfpP+3DCyWEHRAwXBOLecosQFI72fMCc+svj/M6Sm4S9f6UX
p9GiHkKeWPWpeGNTDrAb2UWEgkY/9q5putbM6ifxdO7fFqgiI3ZDbeTeHwBt
rJH6dzf7d2F7nIOlGN6jXA28ySL/l5ycQ6bPFK7+3wpVcONXUryqQPkUe1+Y
CJfLhAGeE6JoB6z2RD74KVYwSLc+owZ4iwryRsMGh3Cb1eFFuUO97yKOJWnE
D4APVnIKirlnuy7iJtB9GpUwW7FwcttEv8Z9exacufLHKGW/zPDKTq8/KBH6
gFZYXGYOcHBDotKYTC3uoeQ6pBHLefb643h1AlFVBo7QECOBxZgLyruxom3a
xfkg/QZzXc34Tzw2nvnufqcUKsVKCNudq7zw/LekYHPW7i9VV1hFxZitmfjY
yZnjNXEhDwdXgXptKHc5jgfHOEXB8HfGwKPfCsMGJdyHfRqSVzoBx8PCEc8d
vJkGRWXFz/ya8SPBsNrI2vm4p5WVNm1qSynSYTQFfD0vrfMwsvrvPOV9chE/
Xec2aRDj6KsPrKPKPZVrdbqfk0FlSc71/fXCzzzBL/RtVf3Ajql94XTvEeP0
F4EnuTtjPY23wLeREzndUNww5LGl52qQzVmc8PL16Bcf1lDkjN5pcp9wURlz
Jk7q5agmtXx9aQ4QaM3IgGk27SlqwtLHP6MiyjOIZxWy7Ajm9m7mqrOaSlFe
Hv+bZrRBCAVy088zyNHC6lgOxqIxpwJllMlXMUdmUhOgerDdBYkeIynpkh7S
c0OVBOIzbwalfrqQ/B/l9RvCJct51htxjejutUyuLq9PzYLyCcotj9LQ6Ww/
3B9UfIaH7gxzJvkk8zqHru0x4nayIoNZnhPPJBbXk2IS0INBM+0Y513xMrD4
oC8PzjiX6ySl6cFMZ56yCaufOqxJ5uVF3ug4ecAjLb+2wmBvESS08TDdL0mA
8abW0rWR457jiGi6fgHgFej2tixFGWNKwoMgyGP7tC4XSABES4Md0F5jzyNU
+bSkFaS73WX0Nlwtq6RLYgpLIpPzhfUFcdBCnhvF5jJN8ZKs8/kziOy+z7rf
AVsbzoYp160xWDkZvcvPOGw0AnNdIv8wYGheY9Wt6fOsjBAtS3ZJt5d0uXre
qCMQ6ix4SKTz7Spf5rLksfTYaNwnObfJh86X2cOcnfcVF3FdikTC7690AmGS
jJ16wgcrN+SWif1CaZEPPr8BnyvErkJuJC6tnVzWzza5sRfTY9bD2F3Uy3Fc
pmYFvrM/6lvMGsUx5/4Vrm1iZJVyj9/gyKuN7zMfqTsjKzUJT+xJDsS82wjx
59Iw2fBAvPG49ZLcKvlBFxjQS/uGqgszn+An0fLo8odXP8J7mE8r9t2KqW/Z
AkuMDi0QwPyoJmcyriM4odpwQRa3RFhq7rcpSawQNEMTL7mjKxIDmFZF2gJ+
4suncWjiF+onIp7v8dyS7SPrxfD1JiTeQyxyFcQxsik3/sRDzpUlQGSwAr9U
o8ebD/M7F1GL3roIk3VYGIo7TOkkQChRzi6aG1ciRqr2/r7erLEfLBY/Rav9
Tz2CX0mXwXLaqQTlGG2JhUtICD82sl+IUw5ZWbtWj/oB2jWM13oWvfk05GKB
nKMkBBOtC0w7PYzuOFH365RiBB61YhVCaAf6dVUU6PNI7w5x/3oo8UttLvgp
+1lj//q3raU6ohg5WL19DyW6BoucgTWn8X4DJqhGdWHT8DUCktlkdvTmJqeD
eThc6LlCBYJjhUpUL3C1fYbTxt5a5Ws5PSOJ5Gx/mxoJLr/9zBpM2ElQ+ayx
rvvAKEOKH5k75T71ikDY/4/mY3Avbk/gztrqoVLIoKEJwt+g+16qQpHwk9Xz
Yc05/HvmFyfYFJk9tvSc9XPOko0k/E01yTYvSF11O4TG0sDf8mFaJzjBW4i+
fHCxG6MllbrDuJ3RXKMkOP+6j4G9UILY/SkEagfthvZZayo7ZAks9Uu7N8VV
/cTuTCxMYSHnbRrspGdCFLgZLWC4f8Kvf5FBBSlEMt8yGnAZ/r7GZ9T9oswa
UpjVMQTnBBekk+YTvEb3zluywhpltadqxxCTnIh70n6wHIKlfw4pT6Y2ObUC
CWXNnTYPvWQAHfpjcf5g4smbft/Z2Ebdj1PlGAfoylOfqlFgDuU+pCKI+hd4
m7xRpTilB+qbAXpOAq8z+Mm0o1QRAsnG8UKPwOtfCTuc+4RY9APuBajhQcLS
hX4geeKGRN8gA0FmT0ww2N6EpjrNzsrgCNrfPYbIJkwPQBLuNphdPyJsLdnn
MKKLUNO5UHKjvqwncL6xFBF8MoGcnjZgHqQcobikFe7tzUcuwOojF3rGGCYl
drCBg0MEV0U9HYiAY7SeRquInQhTX+iii83r4yM5Zu8a6sQ08uAIxkyYd+IJ
5Ef6ILtKABh1LDs3ZAC5RUZbSbztpFOafBQqIl12xF76YGyX78jbY3huoRvx
ieuIm13B2EV9Ij4VtQKUzIzmBZUCafOI9IFmrJJsRlFZ17psb0opNXcHOYTj
bbiR9PLZSLyNmauX1VmrDiUdGQY8C+31YWdJWpsV1b26ZxINFo55lANBb+jq
GF8A9U63qWwfdKei9nXF+T28XfaQZs7/fIYSd8rj8eFgkOOBjVuxuJumz+Bj
tpT1LF+UEqt0b3k4Ny7nEAlyCuqjJdbOAODz5kLx0Cqo4DfAPxL1ibPJacfO
5QtdLK7JzlkTzkTBCFR9AtYuWgetGzFQoi++ScrNIVK6B2U4DDX5zlR3A10l
SAoOLCqnx+pWLcp1XEDOzPOTg9D6nE3m3tUJNFkDKvbYtkWHkbQy5ka9TtZy
4kvmwKru1Fu61H6mEHOEqldHPp0VwIHhTBV8vFE6P2KD8lmc2595l6ZXjq2z
Y/F2aUzfs7ItJXE9JtErhQ4DjP+o8D3zzyqtiavDNADevqH8D6KfEbV/aotC
dtU3dtXJ6vYmeNuP3aoP1gyycQP9h3ETNlvzisVWVpqIcEQRM6IRWG7Kj5TC
jFi6VJ/mWC45zMKFB9qhqwq5QgwqSQ4Hr5n7G7Tpn2pW2FtnmgScGz+16NHm
yKrhwK1mSFl0kDvouT9Q0/bjEPWYXRIXGhVpM6Nfr/Vvy8cdjCKSm6efRwQA
OiI7EOXFiSdy3bZkJOjwIxirdeupR/ttmaRZ5Xeh/BbHhulG6vaoM+qooq9n
JZq99UPkCcCCkkoWs3jxXS61D+dZCsVU+sFZEmT0OmfCIqI8t9SOMBzIvjnq
b5Xi3417V1u0VtD4H1yKjLjZpRDmnw8A7e4YCXa7sRqAno9GT4e4cSEDrkD2
HMmQhc8ToLj/wgHoQii84YdwD4oT51tF5ZUklbCWeKPSRgrCKEEAAum0XsDm
q/sb81pG9/1cF/LeQrSZo4ZONro8rSFujTPqQ1FKTnbQ/bXxBMWprEVIzPw5
GT+awsXEfPBLXdzcfXvKae+fvjspnGuftOtI6YHbebtDgqMumW3c1Qed8j3s
0TeP9iW7kMhb1/7ZgPna/WWHlZ/tF8oqHw2SXoNzg0hyoRUfz3+EV1e8HDBE
zvwwMvUWuM0ytmpCYjMyqMA9jxOq9YTITGXyA9kiMzpue/5mbmnfDw1zKDZp
XCWhxsWK0md/M4a9IsrLoKuz2LfwzGjXe5pjDgfY0qRc3yptgPVxPAlrOgz0
8qmcOOZA399FPIlxvfJDEAFOtZjkuG3doCbbspaaDM0JE99KGuDDaxSFGy0E
kbMB6/fIHFPBxYezDGYvghqxguWxJuQfQht0EkHMhdF9ylOY370uN/ZEnk/H
X+gxVU4B+0birtRmcvgDjfJI02XlausJBODGATYD4bjAHOGnzridFVxH95aa
S3c1qoxp66PbcKianOvZ01GPvUVIbrBMngA7xQm6pTUfV3uGi7izv7BzEe8a
lqewUO+jVupqcqIzSRjgGP2BZW3stIdYxrxpR5BGCKyIxhDVnawXIdZvG4Vd
Y65TvxirRaZQSg+HWAR1OLcoI3a/7DlIqVYPiChfkRrkBPvbNuZzJfa6Sn+X
/AOq5aGmYi0S9+1q7/XzqEpglBD9T3XC96Kw9tusnQ5ElNehy4xcsaVXhSXh
C0OaT56hJ9FDS1nI8Ot9bbd/+s0esDvb4uhrkABc5p2A54A5n58lT1Qs/TNH
O0FwZweV/NaNn8L4zUseqsChS/L1Ic5anYq+B8tBl8pfsVpNaxUkevZw7a+0
Z+SNrZ7pOeFpxbokqOYlIXqghdFSeGaRyuqx4pCmGpdkpJ2mup8iDdRlR9Ao
BaBzRS0Z4tcNnB1Ub/ZnhoSFcsFXNej2knIJvF4c+4R0QCMTdl6zGdbSnzLY
AZxg573ACLKCPx3xKEDi378/el0FaWIv6VnxXeuxl9DhDtrDdcNPnLWuBsHt
6bkqnfmjEJiqqjGFoQXuuyltvKo4GdNSXsw6LQ7/wYbD/+dGASyF2J/Ox5SB
3N6f1yEjBohsZpUdY+GvRMlfnC+II92Ki1ot+QNunZIVv3r3HgVqkCLPzM7h
VUaaXvQkGQ+uykpwzD6vZLJJYYj3xEWiFPUdmKNuQ8YFE97na8XGccYsLDQR
g5StdMmULNCRM0I0iWynreLVrw3VWDztzjARQbFkBn5/PdagCF3PUkVVAhHB
WLvkkZdqqu1oiQPdH2iWdm3GycUUc972HQLDsqvewHQSw/B5cQgv39+bNbaY
r95+hdT02YhDHTQWm4tnX/EY6up9Z1kTLvlHWWOTYEjWtGrVQNL4UpPM2i+v
W/tqPym/efaYWmHd9+skM/JtGSy4U9WuEdvBlluBVnRu7t34d68xiV5RWyTz
waGrysXCwdR2vZP1yYWjGL1Tnfc9yy4a4ZXYEfjRLFIJyjnSwg1SuoRiwWuE
XFvtDpUPK0XbEVPbI5wFDC2FjL1Wcym+y5bWQvpfbq5r81nOLajMFOEuE8Wo
CsI0T7ZSU+zf5fbkOfFTcS8We8KA1+I11CiEgkZTliugG336lHdYGKWiTevl
HN3A3O0PfB0Ooo9yX4BxWdv7gr2BnWZtAR1XIOEuq12Wa1HbkIEhXKkF56j3
JuA3mBuIFvh+rO9vQSxItZEmD0g/geTMCPupTwWRXa4OTvaegnMqsL/F4kX2
JrMi4U1gkYEa17JmWpsGSQXU+oDNOg6gxS/2BDi1vIBqYxfKiruavD94F8RV
jmkIYLuC+XmxcR3dAD6xSoJn+6JrVw0u6ihMx1YjQHIxxPMN9UGcxkWUvR0w
iAs02tbesNwMYj62RROSgvEQhPkOWQNz7xawo4/exvLdygc9sbBcie2rK30l
QJSAQ+OsWdl3cRgmph4ntzplX5OR0RYVe549Yx1bPTtM0ZPnt+goo+GMz/jC
5nQulfzuMiZVltw0ighqvnr+2p//BG7R47B2IIsgw9sdTRhgkw5IYJcUIc2d
iZ/jEy3nr4LFEm3KGS/wsLz2GMeUXgBFfOBC3auqqdZfcD77bY08lXQ787P0
IXoQL/utTGrl1rk3kwowbEFUX7Ksz4Zu8uFj0gNXWjEzNUyUe4gFBX7Pib8x
N38G/NvXiewv5001saEm92nAA8Oc+9ufeKJ8Zl5Nr7adPhgadwkrD/CyKVi6
HPa8xLvyb3urVxZzHwTlNYvrjWv2WHVrdoovg+7a+QCqPvCRFXSy0Bk/a6NT
XYovfUX+6PYa/RTiwzPu365ohazuH/TQSy9W7fizxEbW8E04Uv82vPz+SoKB
J074zRjQInkhwbjZKUsxaiujLz/Grn4c8GeGqMN4/fwQkh/1pxf45rfDACFW
NovXvmmcm5iy0NNNkms//eJz5skiaDBPmti7wjDty7TW1U9LXSzMs1LUmojA
ChbHDtETyCvIISo+WNyJ8N6/peXT9Z0rb8ssTKZK3a+pSVp8UCV+cRpTAhbD
R5LnrPaoJ49GKU9+XNftOgP9PVWuRcCPKLR1EYs2ro68quh9ep3fZDSi5jMm
8TfvTKnmaLWXS7vzs0WWmx5v2HE/qvGmD+5GkOmp9Hj73HUfQ5Mt5L05kyvH
KM6tBMDI8psHmGWh81Iw7Gwi0i1B+a69hBdN7s4XlhnBGpA7s8WP4y2sKOTy
oMQ6+bl6EeEnopfx9uzwfcr4FZ5D+5pUFEiVn2+9vtvTlI/KVqL5VUiRgvX8
OCqOPkEO43/H7iXurZgC3QgygE+8MYjZB34zMTO9a/KaFrMsxTUG0XNl3A+R
1stzoyeS89X2J8C02oUO/MEXbA8z0ikVwGYJ3Hc+kHQaLM4OkbHDmwHmriZA
KtzIrtOWAIi9WK6N3DA/NSRPGqZPaAyDLxJIN37YxSfmBUSyR7mQUuBD6Yrg
ZYKb47y4LKjWMf2+O0GC4EVSFhpGFXqEAhDPlePNcjRWlmLR7ZU94X8PZ4cQ
T9f0VT4h2mRB4cSTzsqsVSa1JdputPnoNap8ON8LHQqA9UytMNj0YBbbD3kB
06EAgyVtui8GkI6fjh/5B0HloIra5OgpHdq8aMnuYkNBo7N/fIYtMigpwWJh
msYNm0BciPVrePlhqWvNxd91QohkOXaIaEm4n4LIJlsC0/M+cABi4apY5qQt
HMbRP3BQQsPHCLGUuirxmVST+lYHXJ0v9wn8P6WQ9CmhIFGZTVJfF4SM/q7g
WVx1DrX4zY05JLFWyUQoz+cSJVTumKlsM4UfVqsRt2cb2bEb8V8pQoLTQJf7
GqArp0GZx578JeAVLPw93IL6pIcdISti/0JChBj5l22S7EhFTuadGoYYQolA
oGTbwgQbU5p9hUT8uniSV7qRf6cFECCuvIBBMdESvK6iWSWcsl4ejYUzIlba
NvrF3odeUf5mO0GBWvP2HyE7IUVZUXogsoBL2mv8mWg4wuP2dJSXUd+ZxYTo
/ODLgxMR6xcazFvTr41B+uyv2Z+lbqRM9v+g/L4Emuh8+Yq4l47q8Gwwb4pg
PfgBG0iK+ymSjNSqWcYiMGzAyH5FhIYhOmZ5g5xLft61NEd48EdSA0U1F+8j
in8pyXbusH0dEdLkw4EmNOIDUn3HuWG5vVqo4zyeVI280+nHq3qUa927L77f
9bOGTxShkjg/0a/KoMglVPYFjJys06Y88t6qlgWqRoKwI2nzSA5/kFiJY6sz
UF1EP/x36gDD2W/C2WGubHLW3NtDBN0qeaCGKWrJ7HJgWnvHnb+PwKgetxzv
TdaJ98LLhsahsKayjYHDt/GqZe+D1gWxoAnALceCsRXqHUtN2097n85kyHMb
02B8+1gmTpw6/qBBzX4WlwicMXi4f/W4RW7X2ErZmHMbH54O4o71VAc++5Mq
FJERtzHjZrH7pfQkWsLGUdMyaZdi56T2XXyLNJXgnGHAQ3q1oPxygZdllaF4
+Dj8IK1H3Cu62eCBQYjmUzrryDpLO4aveyoRkOW2Q5KFUOS9jWaV6QYHU5Na
h1QvdcBCfoeXquyW6rVj2dLUSYynpjIg9J7XLb+WFvhQFvb3gdtmiktSsVEW
tXpAFqPbvbaL5uA7YccWckCnMJYkb6aaIbxv8cXvUdLzozd0/9NAORlFkLkw
Oq1XGbvmzuo34l6zomsdpXCSdK8kpBc63WGrYlF3RhZrOaEriYo89Z9uNLma
iL523qHEXZEn3RP3MLIKP72VQKU9BVaahxPbHLqU2Docou0Z7HnMDtM+d4mG
fRpdVYbexh66vkPXnZb+uChexFemIRa+MBD1MKi41Crurp4zcIKU1q7eHVV/
/0q6NR5AfccZEoUJwVqH5SLFNxGCSmaPrx9ThzQzkR7HpgwLNbwStnZL2v5O
/yO4Y52FSYAdhJgReliK7Qc6FncqigPGu9WxFRAqFVKRNSQ7QjGx2MtIjY0R
skbAlMBz7EMvCf6XerdstHfoL+qqj4SXHkIN2RIKrpkJ/L+Wq9kxiBacX4Hh
HrKBEnX5FduOuwa9b/oi2tFYz3EdoqFXVrOkgb9p+y2OC3YZwwezPZkQltrI
4WsG7lJw3PnGKdpeSXreH43FaG3GAcLJ2nvg1w0S3VCSN1vBpwL9UGTPLN0b
KsDRGOr6wFV8ug7QnIlU8aBY75Zp1kRqtZUcnkpzSix/wY6pPpeimYVIuTC+
Z9N0MGrGqH8uAhwasACbzks7GsGtyCY95kI1X7mu2F1lZxd1TZ/0Pqo55Sq1
PufqzpPytkC/lsL9i0bgcSvq5FnysSqFdKqy8a5+qbvmDH6eZXbyccbP7GCo
3sUBvvYL9+iB5RBcIQaQOEdRpbZlQM0NFHK5pGctKW1wO28YN9koxjG0iOYV
41hGX+0OBOwmbEAnxo8MhMXEQCLpv91L2q9i6mHJCxABEiWFUL6FOoMVwJcv
v0O6AMFQpyOyY38b4gpXnOb/yj5Xa7gQTcDnL7gGxEL3k7snPPIQvGBfQD+t
5XxGdhJsbqrzoQzFDlbWE2RmsaZNoH4Gi2xPHuDi5GK7g0Nfe0O3QMe/JTK0
trPMfL6Pz9rOoAT1aAyE7BRMCUKU8UbGKjY0cwv1yCKUxYQBQ8UzDK4eyBTH
bvbFImRf/G3odri+b3VjIJrFdnDFE2kW9ujAt54Lk1SpMfy25ToUfDuj6gZM
PM/JIM2zbIsoPJr18zT1s3dblhQ138nLwVDr1BvlV567/GRXML7i70yoskgw
mqdx1dJ1LONsqhFyz1V776HNpo3+7EEvWhn63mTpLqWoAFAt8hhyKPyIETpS
XqFdQeEvFmxQSuq2+YPPba0Y1gnqyF9uUeS6CKSYVBzSHxHLjqGnOh8OWFHX
86cVnVbdiPy3Ll24omKLrbDZbC45tkJVqNFRw3XZAxUEr4PRSlqphQEpckxj
xwFBNg79CB3WXG99ab69CMvcS8Hku2PDn7PjnY1bzhSO4noRFE4qX/k6fC4l
r81UT4ALcMfhQiueXlREXJF0fGX9mitlbVa2i1K5JVvm1zXxaiGaIcHTnQwl
6FASMTkwrhfnlj2DTQUyCDWXwY6z0PuG/n84FLFxbCqgK3nUH1BcdAzPxowe
A3x1lv/9cgF0BjsOgpiWO+uMwMIK36JmPJd3llpAXv3U9joqrsuxmFM6bit1
7Id+byzg+cmfoSwdOSeY0pDGCgwwmvn8Iw49Uxc2XERDk2KGhoByVVX3oTsY
OPAbrkVyXd8rLZ9yfFGx1MDHreaBKBBRz1YQKmnLqXdPRm3PAPHj6RIUSNpG
it0TPSQ+tIa4KzNlgjDQOWrsWgp/zDLeVVeB7DxiWVQkv4NhklMT69Z6+bHO
FBFy2KkUNN6q0VAEmueV3TrsIC1daxECnWEpmyOrkM3fFDAC3WXNlW4jUjAm
MQ21SzzcuPvNT9hNW09VLn9CpxiWwCGBVBc/aDkAIbAUcV7bAaCi4neunnZe
FJDPjfu0TlLdhF4p0HD2l3LjFde94Q8BOISh7j5PozjFrHHccWLbkKJokNwS
mCWe79QOQ0HxcN+CPUqCt6v3klg4XuIXX9sSeOteFr21eSbafM2mYwEPEnKF
TgY8ATOb+AvR1KJD0k1VoNtOFjHVvEL32VDL5AQE4TMwgPKOQeen7Z0Qwuoz
q1Jxwb8KszQNsOGJ8pGFK49e6XVorV1Ai6+BZbWBRffH5g7XLFhD1cPRvps8
pCgbeOQLtoLloWfWJYfG21nzyNWvVsCwa2w6y/3OJbBGSGVhuBFRZ/qQzbUs
vdRLwBe3/KGdqzP23/VlvH2EZvC8IE5LtOQ9eYu1xHO9qLrbLE4SiAP3vbCY
PQ8wuRuGvbQCLWX5e6TyXp7l/wd2NY0cBdM4gYBTKT0psil+ugMKdZTFCf7o
54KY5x8T/noOqm46rPRlKNvD/3D4wbZQPoKIvjjwfuM+sV24YnNreEq2r5ws
ppVfFEOjfP6EYJD30npBuNPONxpF/+5wEoQNUjHFq4qbE605MO2bZIWbf+rz
RqGXOsoNo4lAcRQUZv5TLK3ELg6VwdhiYATI4TLWDlyzQqajh7mwsDo/lT8L
MxrEdZYZRn1XlHE5HhFCc3VMHdsnh6nJwYB7cB0E5EJIIVpeDnSAndXXsLcB
Cj/fqS1aFOQlQOXi5/QmxjVOUQIZDoL5yYzY04uCzL2r4YYhdIpyoncYuQrV
ZZVSMPDLES+FazTNlF5TmK5paezr6cwC8rVOiRzyv8qgJ907rp47AlOp8FNx
FSwOqfZmRx5DF5j8vaaNS68Xeii8T+gT+idCYM1ipMipZjVuzoEQusVF3bzC
jb5M0bqgQK4bFDRO1Ohi8hY0k7PCyvAAp5kD3fDzRKCoTi/vVXZMjEwVc5CR
2H0bJISrIrnrF0olXRhyHGJBEcV1F5tqEKcgyElFyAyTF3jfkxJ3+YRcu7Pz
nzr8KZ5WlhHFl5zM3S3TlvZvLlHHzijMcM6z/6aLNzDybvisyXaKN+zRVoWn
Bom5Zqy5sOslPV0Vx00XaskReA35nL3/OLukVWUZUed56Vq0ljysXI4CRO67
PJNOtY2FpZ4mUaU4bua7vf31BFHdY2RPvZSGkHNXgpLVrn8SBj3hbL+MdZx0
3tQDUtGUvNJgp6NHtMrpYFtnRkk3J8XYhaQha46w8PQR6/xgjmnsCuiHzxPt
L3B1JsBzjerM0EBveFrhZOqFQH6uvdGV/CQpEYePwSXhB/jTMz4ZYc66GNUj
L40Mn9L7+0VV9vsOdhCONJV/zEiFolpne5QtUuJn4q1/yuJaqUBJ+wDFlCPA
rcKzct+bm7IoTv/opxKYG6SjHTeeA0obGcTwlj3S7qm+5GGF43sosBayTpHB
NIEMD5F36ZS1viZs9YN9hFJcQXJ35pZL17nZ7cFX8FkbpOFinnX0wBTN8rER
QYeJk/czGEwiOC9N58QXLqY2rtOts5JcwkJ0ayXCE/R1lFv1u16JL3hvERpI
hp7yxOrSo34pRLmrz/6YPvLYd0eYXolcEvswQY4f7H0PValWS+Wt3Nb5Jnd2
mnHZzz52LIDqkorq/ujDhicggJxEENbnae5IU3ZvaLAM39Omd+ECztJjMn8H
gWM9kHY462OUc2zdqndCMPNlROcEKivrSj9JeiIqTykkjiZKxsdoq2i/1GRr
ZEieLvWYLFNJznQmKbscTsRigegzogcJRsq/0elqgJYyom3D+2XeYHCGEVVc
etuWgELuRPhsvz1CJxCWuNaEiKZRJu62iwipri/t3EoGuwhu9idpTwsGfzbc
QULYiX1wR49Hx3qmcjivLNLcGtg/c7jbNIK/twEaKT2ez42P4Tw+pucwEOlV
6xaehpgIAJloBQex8SciePbXj5DCHGtdUIp70UzLxqscuncZOq2KbM0Urd7d
Na8rkx7NbvabWSTPQR4ZsdskU82ShEXjqad6WL8XDbyO2/ENfk5Y9fDRd3wx
OvA8kWiLkO6t0NSTofbYwJHP74QMLRRY/pIwtVjUO6nkZD0I1e+OqCk7nUE/
ey6t4qan3wgbk9Hpd7hfPhNBH1C89kGmfRupz5aIJrRIUeNCeS7QYK74yekH
koWXt3AxvceI3I6xhbYThgtC99s58fD3D54Mfx46m06HGJLoJbfWGNsfnuLF
wr1IvJvusos5JBzah2ofPGgMVRWoWYDH7zEjBdAgF/WuCVUwa+lpi7EMCYo7
TzG58zuG8BllIPYW6VJHFCmYM6ugWCQFWpNmTMDHUjb67nLw3z0d3O0Fgjrl
7Sbf+ku6MMcLXLiYwSuqPVxhmubzjxELYnloCwZS3miwaY5NImaA4JOO9BIF
A6P6r5mjwLo4Ff+O+1Y5B7OvPzF15J357cwkO+dCmxUtGBTOhPhbdf/mT31E
IZD7WHLqegJtDzSBNqHCZPKxSJk4b5V/PntUb+4OHK6atfbIbXxdY55WdjEv
jBQ6ylYra+6DLO2rlYS1+BBMIP6fIQfLhqeJ6fBwWgkNYf7QYgBExnyvWGqX
VImQrzSjKNIJce/xybnXe3zfEf+iMLnS0JQ6We6P3Et64Kl/af1f5gp69K9M
xpM2vCafAkpSihKwQTXT2WHk0sl6HLSUUOokweAmhcHh57DbQji14QlhAGV1
OYyjZJikrc1WjLxNN7b1aYB6MepLk4rF5+ZCWMYrk911dB7MwrZ56/3JUAeI
u3RlWXRnGYxJM49tKw7fH4Jc33Gh9O1An7/HKziB1YXxhS0tu1M2dFobwGF9
8n9kIrfOiOPlakpHOGXB+ohz+xloJJ1ZO9JB2jptdmgb8aSVW4JCcuHsOf2V
8s2b/5Vq5+m24jHCn9d8Lvh7LIEBGfCbO/lEbz6H6oWLqoeyzsd6I4C9LfNm
T5cy4upW/wYmlXsog0HDAxAKmy9RecFJl74xxCaKGE7hYThlp2HHclk09OdI
fHxlC8rueaRrtwqBGPbOJa/7WM7YooohYvuWaQ/DfRaozJm0AIDNXMflHJUg
sx5mawk1pbT3OpnI8OO7MsRuHtDkwei6ks+LlrDlQ3W5pDJ8ItT6oER62Mg0
Pb73ZhTc7wIr31HcIsCw/tqNE1Tjj1kxE6YALvnQXf6Vxt3I6Qu//UjPvZ7g
bgkz1ZzJDBli0Fi5lggXwahjIA4zXZ1NGmiIUiO8dRClmzbqxu+rtkSuuafF
xytjdoO7dMmrLEGnUnsNw9qWa4t2tWqwqHKXxgybXIb3Fa1oDrPdKCBeuSSu
5zSZdJ/F7jKx8gaoHJcgsrx3gzknuzNhtChRYRgZn9jPQ44XRolFukNgglnO
jjlZoS+EF/ILS7Z/bWNu7caGI9S5X/3PyF+rIU/Kyc7gFE1S4fVuGhXITa7v
+lXE36tALLN9BIR+KNlYeqmCiwqhk3F/ugGoC3gyGq5+AxWFbBAg/+r7qCKD
75dz/ocBslpOZDrRJ4+em/33Vwsmj+12dZaOnGxoEqeWgbocgkcZkOH0KtpZ
TbfaNlOs01KGB+f3Ud+Zjuul77WLJLJCWB6a++LZt78Y6Yk96qR/1hpOU+qZ
aFFijOBQlqqQ7ftGXO5x/Qwb9VDPCVEkvgQqWaDw3Rp26sX8LUTIfZ8rHHiv
LvuwsddmQmtQROfRPMnglNlhhjK+9fJhvR8O/J55tEYSrMlvxjfsIPgrQsCc
xkBFw0tpY4ojVAKvWvgTCZ032bn9MhnOPl3iknCaxRquhFBaq2EGYXpCMRmm
HIig7r+kkuAsOqY+lpjljoxYxEJw6F0UQOugtDtMFTdyDT6k1CZRxHdnLrG/
QBLr8PsVpQ6LpqezeURLXATtFhRDBttUAo4HRLVAshbaofXOAmK78vZ+AJ67
wcFZtpavmA6G/2O1xk/foP5jAb8PPtByBcxbuZfiLmFAsyu7wGKGh1I4CAuK
GvbjsxHNnnFbTCVIC4htlUQKUi1julX0oiU/zkTkueXMp+kKbhn8nPDe3vTc
RRylXhbB7zEHLgaDmmCMMwypOwQdx2TRZ9g74NHxiXS6PZC637QT5W9bzv7z
5zOFpwyNTEP9xXdZPXhMq0WJEHa0uHh8LBOq+avBCVX9HDjuTZK+jLc3vJ/y
3S9vQNUbIHCeCDdOPowFPZmpPnuTUoIytpMHOlrbC+8YhWsgYLD8SpiA2/2h
pW07HUhZ+bAnxOCLD0bZYd7NKC1emCXSq0rvJxRuDbH4S7BUXOwamUnmssqh
GUzHGhMFo+AlqGZYKMYAdF6KWstxQUQV/PLAy+I3edCEQhHaDslw3wNH2VSW
hfjELavZHVyk48wWt9IEvzYp3mE+SOdW0SeVieisykyNrTyTz7Lq9bjZeJGw
eFZtc6VD0duyGcLXitm4uArkt+aXNae43Lmg0abX6yMjIURKoY2Qm2L7XRxY
IW/PK/CIRDlUUVYQurQzDCJuRNX40zFV8NEJTK1u3fv7vauxuOBAXCn+Ec8Z
3m8fZLWAioIkzB7dIKgFjlzzZmdGn5FIlBvILztkmhs9Hzdn1Hj/jrrJncN9
HeeVK6botgrvlXpa07M73KF3bw2wvi+OefBADWeHqcB5MxE06H46bSdzfzfK
yLN+gK1NwRYkvcrMXxUZaVzxyy0Oa3f6sutYlD64X3ToNHJfymePlJTi5AoR
B0GniCxbSUIZyKWyiiUuF6k4ClKe4VUA75n2C8UAdHA07zSfOxF8AsNzY13u
fzQUasODnlN/VOiw8AAWyUy4sc/eDiBTf9hrzbxkWAxCnkpXlLuAZ9A0VR9I
azSfLcbETDNFp4tj+KzuigXm5sIzBfls48vbL6dX6Th3Qi5k1jZ4UDTYKghJ
UCw9ZA3aWvs0KbUf6XLqwyRaJRJGo+s+ttFEZAbOWVvyTjiybX3tjevAfNpi
gck+4a0KKwZW3PvnPlil7no3k45W/uPwm7FfLHaqAM+WDi8NcRIbikn81KYv
y3XBESgggYAyTnCHHSC56EUwhezvhm/6bBejYInoiUjXmPNapYPZbhT5Ypwz
Vb7hhiZ2zGAShxyxOk3i697S8N9VqJh6H/BvKsmvq2tIBz4zDM9Cim5FlmMK
Sp93Jo8+e9oK3X8n1faEhaWU1Y3zk8e9elT3BM3Z3krXlsfo04yxqkXayKFq
xBhux+2KDGSazNCIN9reFNv+bY09/5wZzDWhjtmOioeP8je5PHeirspss0w6
rZyEl+tfmUhUF0X/u5PdADIdRFeDID/QclYWIg7iAQVqOOYxz18v2DgQaHZ9
9Jm2+NgwOEMV9mt2wQhs8zQLpBFlRMBkZkxxCWkVrjYhGotd+agAs+jZgTSW
d+GLRcKMXwrPgXiidELiO1QE6c4ON0R6NeiZGDmIdqAusdAl0C/JBIWG7UtX
Gi3eFXjGd3STPaANphpyw9xVCinRrXy2ZxZjuBLKsBPiAdF9hfYnnQSBQO5N
vMwENCsTAKNuZzAc1habhD6OcTnU01woVl//yrJ/H4aB2TUgtyDckK6kLzZz
NYn6Wnh5gK1AX8jxhPPDTLWPVIUA+RpDJYfMTeUD/CGIMld+WxTUNNHN7q8A
AULtSm/+sLvhBa8PfPOy/C5AjD7otT6fCW54wZQlKtOlJsNX2y6NrcobWb0z
6olKRJ1wr3kSG0DrtHjI0WNU8LhTWLJ3xaUDwKivHwaKEy9VhOnCcdlufGso
BMAsgBXCSn6Tw5mC5/DfcCDWT+eD6dlEXxPyP2BehZuQ3nrGNZbOB0dzrWSc
9KQcUvaTA8m/SsYvUYOMRAjH0St+AhImaiayuQr0yMk3a6c6ypuYnLgilDfX
XRPaqgqWvK+F8+xWYNoovGThZdjFRHsX+dG54g3erbyQX8FGDNBAHCANh0AD
OYw34Hxt6RgYkuofZF6+BSrmCrJNakhoWoiBDmOf+g9SWZe63tMc0lzspYJN
Td6T5vTwqL+G+p8DTdMCEnnJnbK/1FOVjctZS2sOg4thUQ8Be9wP2cbpmg4B
/o3/HuKZoyL+hFgMa0jqbw+PTV/lx7wCjygrqRWc2GKa0DANI5oRepdoZ2gY
mvDbeBbMe2ZUJjdpC5xahr3JQDSRkBLwF3sQ09VQJ4g/O0GEqcUmfdFu4thI
1ZtnxMjyxxkim/9pNWA3wCa4K/2/Jd4DH8HemuZBdUkC5+ptxH9iclTUGr0B
dx8+TclbxSMY17ILI/Oa1/x6u4tIHUuCEIPIu2PE6IWZc9aoPr81K1vYhIwg
dFZzlhV2Y7uWjMPtLi5sObRlwzzWnRGJKjE3YIwlZwxt1fpn7rW71YtmoYqZ
KWSFg0B5ajPbTRuVuOBhVIcOjGn8btieISvf32QRa2X0Gz41JVnXme0WnaZP
lGIxpOqHfz9M+E6IMk23O50fk8D5uqdNFL7N9vFzNY5kQGcqutgBWneIBhp3
B0ImOd7qxeS3jT5PaEwncmcvrCns3RbtVhrWv2W7GVs2Q+sYibxQLnc1jHWC
y/o68Yo10ptmDB4aViw4mS8YDci08GnsyaaY0tosJDzVRxZT4d73dau7J+FU
Tzde6UmnNM+2nz+QBSVWQBegROQ9bTZk7NNfk0revUpCOoYFVBiEr4t0/wh9
bEhY1hLKfSl3xu0jcaI1k6FDCKoPPKPyZFv2kWT126iiSH3mGv9cACqejX/K
tjRzLVe3cFnWmGOT41Pd/nL6OlvG3FYt5tKMKmFG0xceKprwinbGIei5+vnT
r7KObq3OcgqmvC46HYzK07O3oAUiW75P4Ost5mUuwqekfcLNGfxiUyL9mJ/g
lIOpQv3Hn6E+tDwmW8DXH8jcd1tAh4oIQstseaGmfL884TfhkQMZdwiOsnZ1
HUVLqC3H7Ula3nH0Ck8p+oJEvCoR2NjoHLWPBljSObBzTmBlA54lOiBdEwCr
K2nRWZmDed15bMzJENo71+X65G1G0fazWO8+BVCe3oI7b0poa5a653Ol96PE
ygunZUzX+qJ9ckI+o37nAKtqjb64uQpQJw31TtaqPPWtfbykNDEeQcIZvaA0
AX6KD4DfBaUM2Mko8+LzTYy2Ge3++eUq6TD/b2+qt0HBdJ8I4GyCIZqB2HEC
AfD3MGr44mXgTskS+D25PGRUco+8ezhgh4gMSI89oTseKcRnwwTBf4IkUGGX
BaubcxaQYkEkefIEDalGvQCYymBHJDHVqcy25eGijdJVY2dRBYiZw8AYmLkt
pzJ76IqjMus8o1sipelDT4+9gSPQ74CA3l/VFxGeG3LAi1fNSoEtzAt3NqJh
s3uNOjAFu8uogjCjDWti60L4ShCTDbMBR3JYZbBjALtvKBDo7I+epsSKxjVi
faPZbpzSzTCoW0OT48rIm0lY6eLvIkeafMIjPTyey80d4GPsgWkw/C78Z++p
zSaa/qGJqgF77wTvcmB/bT0K2mWaBvPr8heFBlj+Q95I45LeHZkf8FLUOokl
OQ0TKk9Quw/X4XJMEp2VpvzkX31oK75SCzk+PXKcJubZMthgLng72uhfKujl
9Fo5pB5PGKt2nrikfcQyqYADFzlVfr0EdZKh7UZIyHbhYzUkLvYV5hgzB61C
8E1wj+2n98ZzlGSR9lxwdgEbEQAPq3S0hlneMyhsbPdge/2/MWAgyT3vainh
tYeP2G6706WpgtuF9xPKjET4/Xm92dtyMBzviit/GBFg2G5Coy+3joIWZ69x
//4r/0Py9XxnZpYAPmXoaW36Ik/2HCZbhELjrM3ILLzm5LliEFVKiFEijBvg
D9J7/Dg+kYtPwTOn6TA6yrFIVwI9X7CwREk+/pk6SwqGTSjb3BPFnzJZMx+D
XyoosZBgizKMVsbBlNjhLWiESSlRH4cnKizdQvcN6PkyE5owZhsrmMYkHSQt
TbA+dVEZQk6wHjN1xUu9EOayXEBTdakSAM8H6VJfUVr2Tzo9Myst0rknewWO
SjB3iRYhYyh8xNJmxjwhUJQ0OXSGWNAHV6oB5hbLlm0Ax0Y3j26GPytQMkI7
7VIoMPWWbZIgEgzTZbfpkOb0p283yqTcgwgAPlopsA88nW1WVtbS026LipAE
2pyqkxA3F3TBr3vxgVe+p1sEUqXMePo77CIu3otYufVpt60XILTVQIhF/UGn
GYaSD32DxagYwFkHNz3wWTEK6Fd7YbRyDl+4nxHbt2anh0XoCdgVjEhNFYfG
gVtIEXSS/7aS2wFGMYg5aRY7d1Osku8/oTPjLYf1DD0HqHj6BjYK0EOTEpkQ
iY2AgSb0QiLuLYYmnIQ28mOuGFTtxzeDIk4cY2/oVTOHApFQw2o35Fxmk96m
F1ZfgGkZJ+wj3wjdH5THeh4w9pW/SIwDi2/1VG0wS2XO9aM01avyuF3yrjDE
gK2uk06nf5Z/ZIZuJUECwLwfV2bKHQHRXgtjV3KUpJ6K6kFmwA2GtS+NbET+
ZG9E+kjmulRYJKPUWHo/KBmT//VlQHoc3U5i6lba5A0VXcSLgGBpGk2It4tx
taU/Be1Lc9V8l6wbLucyr2TQuK0310tTzHMfD7IriYithKpgqjuxzsy9QWLF
BCzXZZDoz5YlUOawFENNyRcVAItR6KGlNqDAJKNb0GAVZS2ZOBAUR7CE2SyQ
Lh2pHNxT+sRNBnE/eKy0K4cWSnmvlbC4I7h2dWogweo/M8yHjmeFQ5ostqnF
3aTjXMSe8QO8hWF+eo3b0YzwsK4aok6slUaDhfUduSRUD5KqMSfc28FXDhdu
UxXezAvLWDBNLfrheh+l1LmpsO9DPqIe5N/HABOgTCaoyDdiYsflsiSF8XTz
QqQrGloeJ1UXPGLZyaRB6coevCdMIxyMRbP7/2aH4xPL5UGHq0Szae5OZZzs
FNTgpmdwIjGmbkrzCK1oDko9F0dUNwLgXN/bnyrb/LJMNhKYZdfaWJpT4rNA
qh1Wm4tTFDb/Da3rwcCY+pWUy8E4Pb/OpmmAyZm/RuTTZCgCF1Ul01gALBTO
fj44BeH0c+vCv0ziUp7o0p7lxujFiVvR5Cwk+O8/xoEINLylZXtGsVwF92ST
vNXAGWszRPCwRsgj708jQ2TFrDJkuAGknamwCSQ4Lb07b56eWGTzu4lkJqk4
+CnvJQNrGz6xSjnBoRbpu0DKKik1oxhleRKHfL+dUn21OJv6qFenWSeGvWUM
O1XsfZq1Bh+pimimLPepglqNomBtQJorcbpydloApPz1NA46afiBqoEyQukd
yNgU3OqTYH+H7grxhg6A1u6mutDRNHos4wDIs4UJb79yWeAQkxqrDOKLB0KL
kXGWD/YIZmtfHynfV2PrxC/Q4DlqjfXK34+qQwIXMcmUYYFfxjni+D92qaXJ
bVloIRVxxBBvFXphlDqd0OCIIDVtQINOTOsDLGhkO2fcJGmME4TR5C5SyQQ/
T2YCk24otOhl82VCrkjIXYT+af5F/f8dtd4EFfwbtbKOme1DQCyUuTH480br
bNRXsAhs1Wb8p9r0t3ISdjS6gLTBUmnrjjFoYnuugqXwcPuBFfXH38U/AZ4f
f2yIS7DDwslE8eHVQtBl8x2g4cnmN1OVD3FBrnKhL2yS+CUmJgmGzGRFTjbf
qZvSYXLzUc8ZWpHV01jLOA3RR1fSwudrmxIoPrK3lW9JpvW4uZrDPRmCdpEU
8onaJK3E1oQbY/i2AcgT5EBet1+O3PLzQr0XyXrjDZf6mI/bRW8sXuvUNNCh
5omyzJUp9+HJD3kMtR6Kq3M4Tf2usJlI9futJ9mSD9vwYJ1EP2GGnRziQrWH
MeIIfUtc+XZF11cHLeLdptEs5O05kRDazzImKnNWZaajCKlKzqGhkMXZDZNC
Yh7PXbaBP7ycOrQOINZPHtH1zAS4t91iqum8+1s3dR8dqJm6VqLR6ncDJlBk
1DGqFYNlf/e1dhsmAohbOU72vTudW+SZwE8GOKXFDP4wGkVPCWP6Si4KLxwD
OetwVM7EESjsr7RCxYzNtCsEAQEwN+CcByxZP/UmCw86Qex6MgLP4d71R9yi
NmbzQhW60ulEFvzdSe4oElvbG5vBbUhP5QyL6rTY0nphVBF8qvcekTbZ8qVS
I8lyMWMmG1VM5VkyVVeMnuxnCHra+Zq5wc8sA7Fh9j0D2LZgxIAilCZgdqhT
koMwfA9qPCrISVm0gRAFdk6vmmS6SC6FONuKD5g/UTZaShcOdrJk4HowFeri
42GJ+26y0c6CbYNc2tM33T26aUBl/DFYxbbqln5EywlY0x+wIsdrViDajrao
/+nvBMtghPh3h00KZReScnE+k0K1FaHX92GAklwOjb64junGwuQrPp32HNx2
6D9S8P2dXmRBzx52J8EF8kRWuFvIaDHUq8b8viygi9VZ9xWZ8rf6XtCLhpEF
4EbwVhifMhTph60r9um1v53GY4ALgpxn0a/8uz+usSnjAxcsc5Z+EXrPy3yh
TUHk+31uQtA7Ab4gC40r0ZklIkcz4Kid5XpaYEsnEddor/+elssxVOD9S/3b
GXohDmavMbJN8watIH3xo5d19HnSInYx+7cJfv1sv276ESmmWg46dkJ9mt9E
dVN+rwYGHJLqm54LuZ0rdI8GbN8iwBb7Imi73Km0jVTKSEQdzjSvqoRu3GJQ
i5qFag1jDYNHqrhRXYMU444vT5YwK865TTS5Xn4eoqT/XSrcXlmPQEjYhAEY
zkBKYALZPLfUDMQJx6KmIFNVL2DsMU8M3voDkIwzGgL8dbOnRsm29TONhD3i
9CMNN0AAMW+qwSaRAPsCvkspC7mknEmqr65os2Ua8sqx2X5VUekAJzhfifc8
yJ7BKJHOah/JxtWdquQdQqCz8xUGnaZZK9DS6z8xywTW2jkj7DC0kHu+ooVh
vihAktpNkCygxkdThYaUz0FPuyh/ooPUdAANQnYpqA+OP1T8UR80BCDtHVg2
gOF9VUTPZvtNO4mdvlOp7ruX7kgVpqtNj6hpYYTW50kHb8hgJ5LA8if3ZMaF
X8bCoolCrhRBSWMQfpA77Hf1DQshaEq+k4eW4iev9chOphVQdsR2rE4XK1X+
TAXifLJkiaRHqzA1iDnTRPIYXsR95QJ2TQjfkdWTRjnAb1oH2PJ7okCciaiJ
1QI80DbiLae//YkBn8DwjlZgg8o19nbTUlJropZ3kwDWf2PZhk0k5TAjGhAV
BLEvt07IJ3qkzlxvGp1wB4kEr/4aOMKvPogvp7M7ROjEKXUmiSAO2svfamip
VeEivRbZscgniraH0nHtXwSlF0qUhcrH+EpuGINnc5ME9Sr8C+uAFUdBamto
AHGsiI3altYGw6GJYTfQzhsJq/0P80wwFc63irA2feGyrrVBdZ7YApVP+pt2
qvUtrPxYgSXDH9grLV8z5aE6yoIVJO9YqPMPJTOI8z0J+jgZErWFWHteJhh8
ft1JKMSjJMpY7MBdaJfYSRL9JSoe5vv5YbNn50slHUkUSD2PeD9lBEnKIGeI
UO8ZWQ6ZF49RepbyA3/QnRo2eb2OLJcfVvPuzc58w3DhiTq7lriFg9WNJ923
LafYhty4GbIHTjpPfVBYt3hLUGyLdDN36ECSXP3lTa0sxPWF1pSl4qc3DqrL
qOhWGwLphwWIv9cMgMdUWE8vQz3+/zudKBZtzc5kwWs5ULSwiwkNVsUyX5qP
lc2lT6yfpfzt+qvSSpRCOECEPr2FQliUtIv0WkiXiHOHGpMILC3xGltz4MSH
gJjASDe7DAInYE7dF/Z5Z0T0aI6DL20eTCzhtdG/0SocO92lrC7zQyWUSlkk
NA3kVsYxelIp2D5Orgw233+vU/kgy0qy6HuB5B/k7WOGbJ5BeEJYOXYOuh1i
kRssOdN6PvpVr8SXPg4GZSU+hQCb2ZTgNVvUANOtDKLdoUhofaZnJIiln9pg
7T5ua6h8rfOHnuAQ21sb+kdylRMkMrbPIwX3cU/frKBweaXT1z3cJiUl9mGP
pG+C2rGDnWV7VequzaEdvVHgfeAG2nXdow+GLaTMGIbK7MwqntxniwHgEi38
lwiZe5ShHQ+zabjrukhKicnb3j2biU16X6+ZRv9swlcZEesfujeIs0wKG3BT
V4rq/8eb2iIpNDSr7oaPOiYLRPzs/e94rVuIrVtX6Eu2PUmh/asfLH3JVkai
ZrUR2cBxmwElK2ltA+mPwblG8PyCaQD2gtELuWwP2HxuumsCzPM66s32+cVD
T+Bk5FQn1U2QYNBCAdoqJ/atWIBzodsHG+4yNeLKSj+gAWAjBNCKzWUaXof0
Fy9PzmJHhi9kE6eHqRWd24EMVr2csDEfz3u4Vmb2b6Frjn0aVMT4nnLcsu+K
r46zBlaMICKkxAYxx0Bmg3kP0rSbRKTB1Rxz8xRuVoPi5OeE+sMHotNFXdcJ
kakWO8DuNQK9eguGe4CUYlSmm2Ig8xYkJ4lGwLJW/mYHJFt5wA1K2ZprcfKO
TOS6w/PQjGG+C8daRHCbo9YEDrr55QtMM/DA1TOBtJ4WHdacKb7VHmE3Pd5w
XyXETKE7lLQJQwO+6M8PqXpKfbyyjaAYOdAKdb+yWXiJgEzD/UCVh9xZWZW3
5g2ME36fzm7Jj4Z5HT2sqk0duRg5ylc2z3W633Mz4TQLxbSIJE/8jha7y7Wo
dAvj3hKX5SNSXFiRyWPe9JCP3WamS+Q1qZJXCfI9Vg+dFb1ymlLsHfiAJ3rI
24WlThdmcxGZ2Tv5OV87lND5sfGsJK98NwjqnTT584LGj4q0UjSLDULeRMfg
J9FwjCd6M6+tMP2dvsd4vIdLddsPmIY5OvslbBJwTHezUZGCdNV/4lGaTr1y
rxhwYx+zQMMr6vv3rAjqLmBvVpHf+I96refh5JqfPKJsIcVTMwgTRGG3wCHl
61TZH54UiLrj8W3Cc72Nx4gC+t6JSnAxQzY2mWQXCqUlbt4IBH+AROD2QtyE
PskA3M9lDL3afWk6skHjIituWNKdfR+oC1QiX5F/yxXQD8nFD/ZQtqxhrmvS
JWlST8CU0wD8KyXOlXAFFvu/BpQoBVn1ersdZ6G4ulxqkENzBKyiOEVo2nIL
qXcQn+W62ZzDx1Cjb4KCMBFgl/wIDWxr4LnH4n4gTT1DD4fMpG+0RSfzatZJ
ZX4qdWH2vGLPnOLC0mBLZZHVKzs120bYO2FKOhbH68DXNpocWcGNoPlqCirC
zJZTU8NoC4hwOgW+ft907H5GLdym1CTEjkTE6GoBd1Nue5V2UZnHgFQJLifu
XWKxw4DhTk2/cZ4Xv8WdxSJc1ykC4NgQImSONImbKXx/leJo6n4etdNLefXj
B+28X9r97e6K0tEeTrFWKFKzFuBcbyzkxKpIjeTjWbPpmo6YXqLG71r0pU3Y
WYdnO70cJFHgod3CzLk8O5IAiAG1nt/EgC5/+FRy0/TDgON7vOpLCoAr/2AP
byeG3SsktGcUO9oRo6XMYdWnZLwrcX8Fl3iVq40znALKGgypf5dP3+tX/Hu0
vxXrx57vrJGEb9HF1yFSMQ1Q6RKTLNpG0aQ3au85huTtTu+EZYo8V/PdQTPF
hrfa14kna7izD18DJHAQsqQNpse90kZe5b+2LbpPdxlA6KhKzEERO2unN1K6
FBeo6CvIfacLAbg+UC/3c6LLXs5X5lN/FooYr+oFDMX4+jf8G795lWn32BYT
fLwEzk8YUJeTxz1RY8QBAqoawV64TStA3GFHBFkZko01pMj10zEOTtyzCFPl
e8G6PMQS79s1IHsT9JLQ99xYtOqerDHJYMDp7wPf2Pp3zk9XmpK45Juqe35J
TZRJkwVbvNpKPD5vKZja9n5MY0UVOXAbKYg8vjqAZvz56ReAVbzsfHrs0kZU
0bBtyoaLKx/Kw/z3LItwu+HD1Sk5w/N7p2LcxTohzgs5SHhyB04Tsh7RjvcA
0O72mz2hYbAWVKnNkFeaaG1AuBPo2O8JOKk9QGIAWGGo6xKZUQ6QNdepZoVa
ZX8T4M84ohhu+IuSycr4poSPiEPSMjJnMPGj5rDA3uSPC9HF0plPGfXozAUy
Me0xdbyHV16YS9tl2vVyAQhG8GHL1jf+BV+RIvDkF9sBEyrQrD9ezozZPiex
dFu+ab73Bn+SpEXZwWOlQ7zoo/s7OWRG522TwJIzQrXVLHmN8lbn/XMlKka3
kVqofS/dpLZMkFbaDZQskeB2dVkyVzgQtkP0Ixe/CyjhoDfI/CjHwWnVxIvh
cUDIOI8aD7ejxQ1KCC999UKUIyrJM2JttYLwOX20/XSMhCRPXZVpISTN/EqK
zs+eEmN4T9R7hC9qybsZ0smMuYhVuklRAvqeDkP7DYK6io/+TdiXyf0LJ5ny
SHMDBQpo915v7oA6/D5fAO9DKaCaEyBC5J/OTRtNLuM7x54Hi11/UNYnw7eX
4hOyf3EVid3NAcIdGrY8Er85+221A/VFzUhLXepUPvQyIRITJIYwpwlIqah1
kzDgj7DkicLs+PaW0QVKJts6E73rhoKTPSydrFo9t2nfm4F+t5+VmV/Q6bSJ
shi+MO0Xl7B+oCg9ES0+9Jd+6X1YGO3V3tg1LED2rgxo/2n5OUZ9r1cHHEWY
IHjo6IHdCJiICCr/rsB3uTVIyZ5a824ckJe3A7SNe+VFo2zMmxwKIBZ1uJGm
V+z3MxxuLkbX1nniti+Bf/kv3Ff1+GX0WLh3vGhdei6NHbKGC7UHFmqM/+T2
l4qVSOQkBLIWLbxyeBlkES+jWIyDe8HdZIeK6TSC3QAkhk1KnlMfvmIkY3zH
yGooS8tI9q/Uw0LT+wN+rbPN03Rdxj5iBvS9G+qQy6W61bCUtLC7vjJg06e1
KVe2loUSC6aC1B8hRRUboTCyi2vKENGDkVEHVbhGNTZY6Yc3BG/OAj7YNsuM
eXWmh8AmLESbeyA1VgyUvSL/kJ+JjdIMnHgjmSe3MIWfnmibe5et8WZiuXUX
RWteAi25tX2o+7YMCr5zjr3Q/AbIpRrRIqgK1THTOTtmeWVcvSOdHQxtZhQ5
JDrOyzeytbDiB31FIfa1glNpTM6LdzDktwt+8qW5wiCpwoEge9lUimY3LRc/
vbJTDDcUds1/eU7gHbLlGjW+ckJ42MYOs/U+dQbOqs3J/Noz8PUivANtkFjl
ZcoO0fmtN5oZYn+9LpGZtKPSCyo+2Ehzn3mB4WSdqCkJsi5PaRMxWKb39wis
PvTl4AgGS2tMDFIljILmEtR1OTjOix+yDimcq+OnVOqj+MAUNuubmiJ7Z+WM
xXRZSvn+4St15st0vgScDH+95AUp9TCQO+x4V670DjvmnOTkkodE77ApORP0
Vu4qp2Klh4TkZCmWQs4QEkFLI0thOOrMhxMcG1IEkwJ6DcozXMxiMAQsGN1r
sGh6rBnp6Pj3MSFJm/p03JfoT68DOwEkYd6n8ALZAEyfiLn7BlGixEAYaiRE
rgrNuicwpdgdZvaLuge8nPtuVw3bihM9Hy80tTnZZZgIY6SaFdcLqB5vu9QW
FFcO4biaYpfz1ntfeSkeRD6EKu3/2HNXnk9E9/0QWo+PUNAR7h/JUVojwoAn
GIaFz7ZTPBYzEqEKomEuIyDbowsyd2EjIRyKUXInPLIqndmd+bZCMevazD2h
G2nJdK91bdpk6GVHhqspKdKZbDNgroNVDPohksONpq6nNt2WnEWadppjImOv
7CZ/znQcxPPcYmVzBiGfbIvteMu8zby7Ima84UnKFd9TeniVAIIfB29YF26Z
xszuy+PDrP0A3OyiQ2Z76yqL8Odxl/ZG6y9Bf9buY3T8oZoIAL+OTWifBdc1
gF+mljSXVAeY3Qay4bxVlmvFVU3xP3aeoi7ikFOeNeArLu4ihZkz3XHYtW9F
FzXoHqsgNiT6nBDZmddi635cZdkfiI5hHqtfc4PkFWOoVwtLU/kgiladmNzC
vQ7wIE9L581GE+WxmZ21EtDTBtG/5j9N0LQ2wUaWLBJi2A8QACvM2EwOLymV
GiCsC96MVMVG7/kHhYhXEabe4+uINFzQ7XBPN/djL0IozIxwH+ZA5/Zo//Sa
atYrH/P0/4EE45eTuk9IQiIlxN8N6wW+gRLSCzu97sCM3EvE9R8lpxMGta7V
N04/kvqVXDXSk1C3z1TxuoWDY5Yfhu732ew1JfKzKoPJlH0FNGW8DOiB9Qqy
i7AN4NlrVFtHAeCBfHyxgzL78/v9ZlsuhRl8t/GPb8LlUwzOe5wxgBps0+rN
9O6ugMll31EVHgEI+h7xmpluEM3Q/CMpprYxTqnivCVDL/ooecWK9PyqmG1p
TTQQpT3eNe5oF+Rn2qQDg5QhH2v8LPojelJRblwRrG4Opx53a9ehlT+8feDL
tFfw6VDadLealGC+vDvEv0Em3GkrVd1uxPLZpYPHj7GISbv7ug0cF6F3R8aT
OjrAHsWPNXyJTX0VMgfHxYZmQ3+ZslMrREDZrxtVXkrtqJf3UBqq+lAiZ2xK
fK7hVvnoYSapiHTYrSH6+8t32vnogLDysllPMChSKdcP2qlmLi9lUV+aHcNy
n3fDySUhtwvFBBAr4CPfGExbA6KTOMX+lJ4efDNuYUSsMau9EByO6DJ/w0Cp
RO6juWZNziskWqqG3s48G4XHGXCYeeXTLiEweXr9WOGmHb3oWrj5K3zdY+AM
kHI5ppACnxm+Oc/r6/ehDy+RE1iP0VCvLcacY3w34pmBe5gW+4ew8/Dm2JHB
R/N/hEjmN1Lc1vSdpfAiq4hjXsCKMrhm69ul1uWN3fbC1cnVB3zaM9y2z1My
ipIGdTJvuNcftNT4/Ul7LYIIt8W8kxNwIf+y3cHIEfpma4FTLQL+SImJuV8L
8ljPUt624NvgriGPy7mdDB1oUrPkxqUVAGxtYI6v3Xr0yvs5CvRtIqZB1m1R
6Ppg0FwqMTGU93DPt18H26OSMdI4r3ITENWoHnpDeNDKxc26IEnVCB6RRtUp
Yujuiicj6bn4HJ9gKWspXPZyNtGBlzOTTJcQtgWQCToghAbl/O9KfdcN05js
Oq8p7Kh/2wFs3veNTgz7PYGc5mix5cvuAwJF/7xx7UmIBS2gf2r2jSxmgF8A
wAi/zOp4C0kLdpvRk+JyiCj4PfCCjnsZV1iGTEmpBaFkMdd7tqAdUgpPZdc6
jvWTO9hwSybuexASTEQDqiFUBvGdMPZ/WYmfoHdmuB7zUdXoCsu+BiBiiJQ5
iyp+kPE3E4cs1MaUoyK8g2XM6kKZLzpRZarYp4QQAe8a2lLt9pQ1YP0uJO2s
5WkK/WMf8olr99bTNgFI625g/hq8w/gdWWAJZgH0P51SgNwJex+fP/YTNhEa
+PtO70rusbiS0dNtVcHsOle94SSXel0RABeCY5WoxcM12U2DJCINB1TzfWxz
1OrmXr8btLAWpsZqDYeY8qbsAC//ojomhzdUsBwjkK8DIwSfcAMZaiK3+FRM
vfSHVkuT8tkPIibWNlsGz1UpGgYEB/uPROfDgJkdTp0aADlNBp44DcBsIFI3
kINRnRtU/1KYza9qRb5aQ9quDrYbL47/bjcPLEp5807GeIX6DwgnXLq3x7V+
nNtt0hLWfamzVF6kRlh2yN4J5Yy36RN7i5k6AJnuV/agOLfbGTOCEWUMZI1w
gvZY8RgujA4eQN7ujcVtkK4DHDWY8HCGx9XH0COXFDhTTBFA8jQVnD7dM3Si
X9Oiv5a/PiKvwwhQ4CHH/nCEsn9XOA+1Mwy4tKklNjXRt5O64wkU9nrjVFxa
J9m5tta/cg2GhhBGbvaRtyludq19Zq3OqXRDmTf9+g3vvvtiyx0U+poyPIAJ
DiZbK+D3JOHVpENWmjGV+FHoauY1nn2CfnZbJHPiCiWvujXvrlcCqMD6tnlt
mddjeWAg/Gr6aDqR/HHSRc0nm3l8NDSww2oodbfVfU0L0KfITZytkS6dQgva
k5avGHcPGhCVmD3qyrEVzTSbhjWLwpHvwzySbrmE1rBvv4WWTSEY6nYLkNM5
3LJ6LCUXmpQrqumBP8oG7CFLws/69+/YyhALR2OX0YpF/jJcFbYiaLI/mNU6
9tGHEXqNrYdzhNgwutJ6LnvOseUMEHAclsjX6/uGkCyduk9NHfZyi6bRlGXe
sv4cGrJ3myNCsIlvj4djinNqnyOJUwOcP4kcsHNk/Rnlw53tE20Sv+3bA4HE
DkthtR6cCg1gLPujz1oqoICQzU9AL6Y0TnipnKSDnV1Jilzy2Yqr7U1DB31Y
fJfbtR1uqWUT2Bz87s/dyCQXKOtlLOxhJU070NIOSSWTYM0frNJ2OzS0VzmW
XMdR0UcTwEOzkKY3BxYvOen4h0QcxxaMmmxhyOP6w9UbrBaVVkT3lQKy4uVp
S17y+dsR8vqYTgH/qXxTuhb0VKJ67nPxam28bNM+P3b2+BPMLqpYECaIs0UZ
INKTfoid2m5ZAYBfsDbGUXAPTg39tObNgMu5wOLT4NZzi0ri6GcnezQ6kX8t
0OxrSBfred0c//JtIXJapyCl/PNxenDOg46etfnvPwpXEoN2xYF6ZeLsNf+a
6bC1hcuk2BCqbGd58ylXgzhOCArXhCTK4wAYL7yN0+nCcwM4JjDZgRfQB0F4
U/cyI6cF1URnLLbalphqguS0RbrB8v2MeJxnsK618LhxEPkRe7/DHfsjJX2P
zcgAAX0Z4mMF9Kb5VvdSs3w/MBVkG0hI6RDxP4AsAqfEaxI1Z3vmm2zm/BeP
TRJA4cFNEUxLcTeKkGchnItMdNmwjjJ102giZnEmJBeIfrQcHDHX+JYv3L0H
KrpoJom4RGhiF2iEXqhF7jfmrRC9mMps2/5sbNez2JaxbDTooXaf5cyYBSUt
oQJoSa1VYZ61yPeHWh398mjeqZdL7KJTcl7p6AhtyfcuZb2Y52QcvXqi4J8N
duKC0F+7g/AV74QAMhAJROvnOsCBtYUjcV5rjxPfBCk/K69cflQPoon6TRRv
kRceXXA6TBQv1kkVd5nxQmhB28jtKChxrN3BkxuHVB2WEcefGxR6xj88Z2sJ
vmjradGf+QIbw4JM0aQTU7tmbtVcgHNTK90tfvHsXjsY/AqsorMHd7uM7kJH
wEWBhYdQoRuoTOILmdM7JPhW1vbOhMMsAKgf2JZTaFidifbD5PXJ/dByN82m
L6lYW8Hn7nfsP2uxLTXUFOUW5Yx/WXXLQHiBXAad0dU4jqGv5ooOmmk1JO6Z
GFC2DS43CkcCSPbwypcfgikkWjZnrYf87Nkxz8juKp7XUDBRzvPuh0VszJ9m
Ugb/twlAEjIxGo/0P1BPOfrvf65pMvsn5f6ukgiktnZGevA7l721qqrvmlfj
0IHmaqTdEd1WFVAMNKc2NEqwgRmrbDOReV4kMfwSRsiDioTxkx5NfJ0w3f3T
lK9ilTMUecbk3Y8ZIBSN6PIaohpSIFW8sKGa3r7jL51qNEDvKMr7pI8VJZIr
NAkwUkvUcWbVB+pIi6vqGKOmLuJoaT0SYhIp3FzyZrQ5IpZlycfGWF09hJd3
EezogQV1yJ5T4lWhnku4l1sGHKlHvJVy7vnzPRlhy/Jwy+YwMJfjSyN2wXYl
FT25izF4qjGflG28Et/3jnuWcxQUOU1/w3+1pn50zUIK90yJ90AQJdmXJyGV
pI6Z/hH/POg8wgbjlmu61c4xtmmfwlu4ojlh4cwAD0Rhq/kBUEhfR/IdaKHg
hPG1SNGZ0ovNFzmgY1IfZBhsvUbCLWePxtQuefkp826085mzDmO6HypPjwMr
g/G83xjvb86KSbaKVaeo2M8GNbFk0B8y9n6n8mDuoHwiZLVgThVjuN+ceGtO
tdTTkj8+dXWrId7zfxbk8xRU8/KPNQ95guIt4+41zr9q5uhswVTRl2zOgmo+
2xZ7Y1PjiIAX1+Yk9nk0x7wq7NNyHSnGt+ruea6HW0n8yJpBc6E4RpPEi5iv
B7I0Xgg//Wsg8j34zoFBVChGWJrymSfEQfBnrXuDZetwo+wENk1Qk+sWxAty
OaS3snAp1dnQG1I7nS6INg/IlVMjn0II8IB5CAVNxRh5oEGVilAYWXXznHf4
7YxY7kGf0dW/9BK7Ccod2PTLRRt0JhicaZA/YPWISmyxSz0L7Jv3SIe/oTz6
GwFprLcjU0lh8EKWOfxox85kTsmtq/0jx5hh6eL213InZtNJ6hFT1Ht6KXXF
xamdNfvBmT36IUnnZsGuxy8KhRhcTMP7RvBOKMXinnPzh/zhZLD33cfYHhGf
W/j64C4jMogMmxtJW+NBd9tMnYCjXPKrpCmpsD43Cejp36rugrTDEN/YJ3mv
rj1RZ31uyhNlX2z21Q3qn4WYkllt5Xbv/KziMseyGgvpyD0CKq4Fz+q0TlVt
yDMwmqGBGzZ4LAVl2tUp0wJk84MP3RcufeJZKP62t8cvlg2ULrTJzJy5Banz
krvmS8sIyDFfSUxqQ6FPEqZ4zDm5BIqplescF3rrqcCd+FU9uYrLjRbhlq5q
SCGeqsPjo3UzwiNoMRV1ThEV01sfP590O3/6qZrxm4r3v1MwShTJrodcP2df
tN8qr3287+uJTmt0F14bXzcj3LZj+2qaThakasW3ySJYdqETrMlHuGL+L5No
9rnQUzGmL2wB76IPtPGGuTAfN607h5Wz2iE2bn+e06kmHq/c9PLHV8cYnv11
6pB3FNB1TBZDnrx1CcsAhVd/pkOkR246CNJaF2mqGg7aFk8vb+tTb5fiTbMR
fXbroKn6/QUczhAX7ZnaqEVaPaCJbYfx645S7n89XPLRzem06NKpAXR9Oqds
AcAvWtPYw4YVphrCi/HyD7uUsbujKxhrK7MwZR37wY6HyZBtjWCyi+A455MR
MyZGJVvYi0JahsMidfRzbOY7RaYffz11lKGoZmqIlYwcHor/CTZjhoYbzJQN
JtSAAzJKYKLsopakPHIRBHeSmZlUo81fIa/QQEjIVeZraaoV6lzjg5C9l+Rd
6yW+au4WE87sP6BrZUucyGOxnTtHddcg+H3dZwnKVanGvZ2XDhTThSlMEbi+
M3DeEF4jPMaI1Nur8pvkIJGM9JA5UvSrjrSNPDY6mI2mbGx4VtS6HmuXJRrt
bbm7HTwPPw8PI297aYOJNFYKvcb7GgdQ3dpMg2ZibSyBJwZa4JpnxOir3MsD
6SZ8O++ojkCnNPouTPNy8cAy+qrfsImxKyzR6k0cLpVB8gVcYBftYOh1HgGQ
JfQZAme/q9+r7JNoJho2vtAHQzMCprgAI9GH4L0due0m/7RcYjEBR9ewzAXM
Ltf9laREpKr+2yjTFEmO27RleOH+/fBmiZsW7xFtgO+R6r4yhte7mJqw9h6Y
10jp9M1e/2apv7TxMD6gnt/ohkAmDv8AapxHf5dKbGt+WaTU5yNj3CC9U6Zp
E58krGZABtCTrf/8UbPPAVNOY6naJ10vOye6TJ5HwX/QXeTDQnBKHGV49J7b
5J3iQYvbZJP1+20psFNEsdGgBdpKQj7QaDRJhrBGATI9wcpolfP7I0GhE532
OjN6Eq/MsIXu6JNFWIMechA8QvPCjh2UL9oxD+CyUsfaLdGUdKwrKMkfTDLo
VxzexjWTgQJHYfhfQ3jLGdihmfyCzPZZO89bKi8tPVukGhtLy149oK0oRZcq
bd9a2aDBo+og/kobLB4fnhO8V420jc+Tcd6KGCqXnoZ6gLvYZviRIGnDaKFT
B4IMvcxS0AttEqXI01NUp1TNmjcOFNuulMChABWYePJJSRJt6f/uIbX7VFJD
lT3R5zXbVJiaxyPXVvs377NqNklwWZrAbmWXNOUCS/KA7MzvzsDKQXR/fEgc
Ed4yTPIlxDvIoXCb/RaizuSBYYY/qzJ6gI5pkKIaCq6H6VdYr1dWGkv0AvRx
v6qg6KLEiL6+oX8P8TYN1DP2S6N19L40QfWUVJZqGMnY/hyJRqGBMiiIVV/3
JktVzdE/Nrrv4qGeWCOOtCod0ZJ87Eh3SSlEWFh5qabfRbESJm2/A31eXPp5
eJUd9w/JJMnGbbAF2GL9tXO1SUbuBBJsgBeXbwUCp7riuDwQSkKBuvwzIxkG
Idbv6zWcC/tbGiJOG134xSTIidLywmOoCnmZ7qH6VOm73tXrovAA7Zu9WcwN
tnqX00zJzw1zDGlsl6cBOgpg0KB3qMOfHI/rQtEBpDG62kCiu7JZN/XdWTlW
Cpl4Cb8A5jZrSNHLqpt8bTg/0tXxPGlzmtI1sNSIix6HQt6fg1nMK4Ilmh5p
XNnvzurYdVtNwG3j9tezfrbDSSmFLMLXTRfgoTqZrMlJXN6ghKM6Y3aUw2e+
YGBrqF3892z6L4SWQAHV5t/1LThX40RLK/YYyVlxSP/35ToXmeuE1UCiaMPA
VUDQzxuoK3AtDFjCk2mo4Jjlz66YkDCAkzPSwpkPJMGRAGKdWAMgD5qqjoWa
OMmukdaMWLBvoEVPWdw2VRdgBZnrOtJmoo+qRrbBGE4/OIKxSmxx/WIF166Y
/zwZTITY6PprsWXCzyy5rcPMLOzi2wVLkhRm9g8/Jy62qBG8Z9+i/Z4z3A9N
PjnPW9KS1uGyjYOwl5DgY/VEEL8T4Jye+8qOX1ZX7sNvQ6MIfeLVbxe0/w2z
oPIRnMUKn0TYY4N7FrFv9C3zT6XlCfkGc80GOk2vvwPaCHbaWRJHfQFtAOdt
/Dxc78QXUhYNnUE/a2Aq+2L/Ld7zgCQ/9tnVXUUb2GryK8f9SP82DdPVGUsc
41Q3VL5Jmq3TqXhpSb3RhrAS0BRNrWPpU08i12F0qWBEY3yF1XC1JbY7Uj1J
sVuq/B+D8U4z5I5D2ZPFil1yKpisNox4sQdZ+IRV/apsqt+5VILdamNfCBLM
3U7oxI+cH3nTUtFPDMwXuFXtsxvnR/nd3KOkNcEp83FjBTifEGyjbutUigc+
GtLni45KGAhmOeh8rWkgPji46OnH/Ljf/sOJDC8R3kgaTGgP5OxiYnX4mLkJ
/ME7w7zXTj99oLHpCbjl2CBuwZeVSW/nTqsHC1I+wAcWJLl0ZCBeaTy0ub/W
uuAGpseRnWjGwImv88i/TUGv6budVyyZl+uWyh7Quec0A/Mk0ks3j1MH1UqL
ZISEgOmBpcGxSKEcyjz/7Hyc0IY87HFPhONRqz2CxyY1Q5yoB5MOtQ8QYkSx
nvsLvAR9mDS8iQFXykqWDCW18EGg8FfxcuFlNFbv5LQmp4kJMmiCbbui6eu3
iAKFoprXt2w4IdA4nfqRXogK+k0eL99FWA6dGhkprGkJ49oRLD8rDY9cgMFk
RKToeik8q8E180XrgQ4cDg27qLR+bjCrmc3rBZ+VMBVSvHiqPVtQ05RaCLZi
9V1l/Au4Q8H/w9oAU68w2HEiCx28JxQIMSvd/WjIY3Om7Fsi3Cr7vRZtj50Z
pzwP2ZFjbhurP7a+mM17voNmAtjyK/dK83o4Erne/I6ykRCL719xfGu1jiVc
PW/xPJHlB6sMemrvziU7JcydPWwjbS+3A04SC0dh0g5qLUK0vn9Gmfuf7Yqv
sj/BZAQ/oAaWLjZY4zT6d8qv5qNTKAnyfXRyxHO0UrpCbPrytV7ACQtO7L+y
yaOC8my67elUkdskT1oz7y4bUs4nTJBMN5Ju+2Tn8vDYmCW3QRVMfkCJqq3C
YgPslU3lUVs02dUi8rfS9sTWgWjhBghuVJiasMBJG4O+kyhBEL7WF8Va+nMb
dmOJrHRwBpBm2aWdy5jVci/5Y1bt/D3JNEE02dGXc7iZKRSXBd4GAXm/eGZW
gLoH9pIbvVwT2zImzElThPMXjv1QqmDr29EkxqRCiDA9Tc2nY0XKDeiOOojL
v6kkXdFmWPI3IiA8dHC8W8Cm2DUaCrM+sHMmwczl9wP3PpzICmVq8SblEdFv
E+7O0KVUtU6RW6Soi04ZyN+ZmSVWAkqqnxf6SCJ0AfnFvsRcd8B8I1fhGuk5
+FYVxYUdU/u9apkJbVd9nxpEcy7mXd0rhOV3G7DMn+Ojh8eTjB1wHu6vtMNn
TB0gAHnC3rmfvi/WNjJBfP2grsspZPuA2QGEslZmZnIHMlqrh+K1hauQZdN5
1T8+uB++S+To4tqqnLvthZ89bPKKOFDmOvSpG702QJJ0grMA+T4QWlveE2Wz
ZFk6bu+C7xbpJQknYHpHK9+dxVOdFHRF7TbKZ6shnmVBWHvX9CJS2475ofei
aOgKEcfBgxc//h7y22xhYfLPsFuPwU7sGmvqFhq/Sej4SiR5Fodd6lmHSIay
NwWoClkytD1TlY7xcQsrBKFFfx+jdhWiXcflpcFw1YwQqAl3m65Uw8sRQmWK
UUfGgYZTwT5C+uiJGHfnss66JBczLzANo7DvIsgHjKvUVQ5cnoj2vyQBeE7G
Q/DNItLOFxsVvRdgfw6r+8qOMdE12CxEjcmH/hXVNlTTUEmCvnT4S4Pu/Y5I
Yq5NPNzKrSbFgMMoINVbIaZ2UqqgDI4lSoUNHLmZKZ5cGA9Iszdrh9GJe5H1
qQYmWlbI/YrHLPNmSe3cFvakkmcVg35zq0c5eZeag3JN84I74j4VfaoNi1LD
tAD3AunrFowsygGSa4BnTe8spmiqdiDLYjkQ/PwgVVbuui3H+RNm+uBMQCEN
7c2/nl3hExR1KypOv7o8jfBLgkHkZ7Ip37N9AI0dgJSije6H0qaV2hFsYsvx
TmnT9QSF9Jd+sZmyrYEyH/Zt/CnO84CmB7o8aaw8gF0bLBz2n0fWJYfTJzWJ
Wl+4htaKOkErnV/1oqhR6xINMTE0RsZcMHz3PfzbE1X0sEyOjuiWVUXPu0MG
ZXQ4XobeY1sCU2r+4QMO1mFgT9bud39Mgv4VvHRzjCTldGkmBLAr51Ev79PF
MxwWOEGQcl9xzawBcj+tc6AvZwMWFhE/YAistn+ivDzGqjZIoNHzYksLAO8T
eXa9Ok/0IK9l+n8pJ7IgqIYzb8wKX6BLDTgzEahmD9t/O87aQznyAR25OxXA
BXv8w44NO6fdChgMiyKAsg5yu6RAoJmlePJu9vXR2uPUw9pMwzRAKaITWXBX
d3XI4OATkSceyMqkpoisBVhKr+aWBmyWhNQFi5zXlByU4okFhZxJahGOAdxR
AXen4Cgi54abJbfjCaRpl/jSnKYyfG8SdksuvULbyGG75gkCrReYWeoAf3H+
HbVXlxq/3l6VMB9L77oGiMssqWnwTxiIeH4WNR0OpxM2Uq58aS0Z6cctPulD
x7/OC4v8hdOAhhKDsGxkT5fk5FC2AHcMjWK2TdwpBeDVG28RIVjYuSuOmXfJ
UQ1TFW7yo/t4jKNsZBacaBKZQOrfcwUKpEbY2rLskoXHJHk2YG8PQuYlQoAr
R/FUwKcxo/RNJE0GESP/CeMq5VoQGwS8hFeLP07k+ZtbHibqpGM64GtAguoz
z9k7qzlg1gT6VPwX9aYn6CkyaEj2OfOT09ef3X/Yt3mUqz84msBtgkfDPJXn
nbm3bp/9Kmj5uaqkYIYgt+AOlFNMDnUyyi47wF/B3wRfzSNf9KGrR8hbihN1
baB+dwZRe7KqKgfcsyvu1cs7/IP2eVvePiewP/yxIHtD/oO1krI+Hs62efmy
dCfyGkQ9XmKrTQFpPo4emS83Y4oOvGVWZpFI490MGqKkDAzvTe8oeXxB0OqU
v8aws8K9072bnJLGxEAN4QqoKIyjz1eosbPydFMMGKz7DmMaekT+THV4+U02
fc6rnOQ4Y3oAnfP9DnrzFMVxdGRyZfi7d6yn0987ug1KYGq6IMCYB+MkMXfz
FE74mLVQOQKBRIis6PbwmpKABwryTI994y2LXqBc2PLDUf1YOtvM1bV9+Aas
iugKxU7tuxAn8StnYKjuU8jrq4QYFe3mT0IFYy4PDtCdiBRRStKOOy+n+FwN
MZF+Ff8qo3q0HNEyh/VEz2FkcOB8YvpByhdmHiLfC6/391qaqMu09QlwVF6e
KR1IIxTLE/M2Ch2b1srf2cAqY1nIzByNu8m96sh1X5KGRNsQkfGnwcqqWvB7
SyROkGiiMw5oGNH5UwqxNQcxEcPfQhcFVHpaadAq+gzqF3k6xO3PsMOF9Uk5
91cXQhpmDm6DsPobgrZ5NCxt7JneQZ8NkYflM4/dNH9mYHxDjlI/AnazIuNX
m6HHAKHsfs9/Nr8qLHsq29VEdpkVjPzwlQ+yDDUqUnVGlbAswStLVXKETty1
ETwmHYT1bwi6fWSEXtkb6QN8i2tijGmv6Gj4y+z/l8sfvwKfTw1GNqQx+S4r
EeAZH6s/YxP/mlwDy3GhPJeFKZob3hXdEbLZCYyXJjln90fXM5xjyrQp6Tuo
HXFn82QQt7U85ZlISHumoR7faM55eb80Uex54i5tWDvEypPzxCANSMOdqY2l
LsFUFKeLvJsnb4UD0ETsop0NHdBlo0jPbQbCNypCd+q3PRohyW7/LS9SOxD8
THqaAOxvkbK52G/g3C1VsxMApfRi3CtHHlX3eL2E8ddE6ggan2KcReCmmTq1
OcbTHYMJYBIJ8WoRk9qCuOF/SJlbSmN2jhzr+FqqLxJINxuf/3i2nvKx90Od
YPLOCoBNfdXKgWmbUXgx1IxtO7kM/IwN6L+M5kGcRCBzWlT9KtvW285LGtG4
L4awDypjnrL8VMrhrCmssnPg2YVz07w4HFBwSJyxdz7qezG+bRFOWRZiO2yh
yOiM+2k2VMsRLv6//LENvtdWxZG3xIkcSX/2QUH0nM5UBdlU7lGIFsi1k/mC
p60jg9CgK05WLvUWjd+gEdEKbu86Ko+ClEw6tZoAGFOUmzPvjEWYTR6qMn4w
sBNkKdmDar080enKttjNHTiy1j6Q+PTYLNAQwXEFiFjjTFpcIgTEmzNqk57j
B+rnpS1zvKKcq0P3RPi2i9Pcounwqu9DekjIpBi3acxJZd0INbLQSlzLpIbM
JD/eOB5SQHxQDTJyL1NoRrYLHTtR+5jUf5tPboWurazS0Vsx4H/1HIfIN8UG
88rlEwdTjQp0UCZrlwE1Qvb9wZqHxFKPGoVdx1i+wWpXjP/pCssMs+yuL9k2
OV9fonDmtZ7LG40cwFxAcZnmVl0p0y9C6Xpa552PM41xoSATrTIP9MiyxxkP
Cdn2eeEB0HW4Y3n6LtslzdhL+qpmUg+QDCajDiOKu6+1XthUPSwx2FfmUkrL
8FbxWKGXYVski/n6YCEGJTyMpJ5LE38R/woa4Wp+BZF5ILcm8lSmfcKWgoAX
GzVvjoH2UD0yvzFxck/kUR/p/ENQAP8uZzYw2BcFde+EI4epfHVLuF7cenZB
VWdiSNRl6KCzS/42kxB7KeqQzWtMbA4FynN668zrE+nso6uipczsW9EsEbdR
5y/cDRp9wteGmS3RitGMwLzrnVQWyzGOxyWMC7hvUO5k7J/jkDqDgU6rXear
QxS2u+00N31EK8Hm1rFpPEv6R5FzodOJ30S3ABGdM/0RhuOHtvpRHzzupCsf
2abUKdjChcf26rPLXfynXX+Cpgxx3QMYubwMcX7JjtV+BRjcMov1mpqVO5Tg
EGPxy21HPFNmxHokiBv2YbGdvSAay9nrPmL4IrF2j481Me12S5hzpiw0THWP
94AkOdsgGX9PBivi0wCcq/7aQZDQ3d2os4x1kAR6DxSFkL/ln5wnXeUPHH60
NkcyaF92+pqQ3GSCQ+77UpbJLmk9H0ai4JEvOII7W3wbRec/OJOj4hcGEYBx
24jTcuV+WIMJJLbBDqKav5CcRpdXjfx3sL+5OfRuYNvLqwifptbewHsSUIWI
CLgO+KQpLFjVbBpovYChG17UdTVnw3sL57hKu5ltzbeJ2M2NU+rhCaygX4Sh
8Sc/hZOQEav4Gcgvj0590B+0oNsUNy/dDU15yHcRzIzeLjFd9weIVmKv41ps
hVPBIqRCL6edhAC1uq2b57z8EBpST06A1eFe87OxyWwGt6DhS2wHMmKwXhsD
yWLwR4wIKlSee3UTOIk6ugoDBPVKVHHfZosvdOZPFoUPej3ER1RDu0pTG/pb
LfGAy59U3Q95LU+J49MdUEQqs64w9F4Qaqgb6HbQXLL71cQ9ANhTzP/Gyl6S
VIO0jxk60Z4Zxhzi+VHvRe0EqgUhcH2UV8pcnh+UGD8Hxkkfl+fi9fCKcaMh
XN1HIpGdcY3BD9dKnlWSBDTulxyhfrE+DUrmHZ8y7TZecSZ0xBasOu4ipTw9
RFzjv1cmXyFnL8cUgsbRD2zHUIXH2tYLOxXLET7jStZ1+somBrt9W58lucti
RBxY2F0xCuO5gabEWVeWhQXOGR5N51Swlo+fQxDDgM4i85yNq7p/OJYeQ8Rh
6jBvmToH2XzTqiBg5d+k+5dc8BAM2+WaLE5UqqZpHrQbXm0bgV61Nhtm4ghe
NS1iZlyQUlAe+QWIIraCKBkShUPlwp2GzU5krQlWijXxB1oUVAeKC0VQyuta
+AMKFLMkd/6l21WWtT36+BEuumAcNDB3WYiptRpkrLb+5ez8wnZflyudhf1I
3FnDsQiMDFHZXGieZBAfkNdQ+fYsgyO8HSSGZ0TPOT5sPgyOKmiHYCg89TAv
PfWgsR5rNUNswX2j17juOt+2j3TGVl2Zp7coZ22wu2Keg4sSIKnVkRkSp5L0
uOX/k/S9a0QKWIcBY42a8cftwP66QMf/BYPAFKcS862G7fQz0L3a1xTf63Ii
nUvLy5j3CuEJsKg73SW1oHD1IyCxL5XY7uAF30nmHYnzgReYXcc95QT/bHXl
jMUvp6rwHjeMtHah/XZPrRP1JcPcAJxssnDPBH3f3vEGA0c5nD8iLe20j4/q
xbjIqNDegVK6Ofy+t+hP6xteFlXY5bbYVZobFqzerPxRoxSmcDnAd7HXP79e
+S0V2K+q9uyR8lzjAFUxibvDjbF7/UBDiiyz+69fLOp7Vd0HB0FKveNy2VeR
sexCij4Iveqqzub3hsJzjP/wCs3UPDTiz6a2eLqxWsQ1UZtjss5TRvhOBNv2
EBjtxh4HzJwYnk3VR0/A7eHWg2IYjtINXDbJ708/TIh3zc9/EqHpA0WHjlI4
mtwquBbpAvnFbG6b58njFuHpa601LL+Q3gL7rS84Xc0osBT0cpX9LzUHUUN/
czSw4NJDZb2m/3hqsfTit7P1uIWjDTounl7vjknGkARbfDUYiPZ5jXx0YAsq
w11vHVoA3Losb5hK9fVR/QeC8H4GtaUM0qC8qLaBrhfvbgCjOOH7sozcqr+W
pXkXshCmRM4hVHp37Nso/ev9ksQctW3fLz8foBqcLxIeVi1s05w+RQm8FTom
dolTR6Wv6ssb7Yvh5MUkqm38q1QH4Lb97jC+SP4h3oy6iCcKmhoIMI48nMD0
O230FWrXhAmCa4vQmA1XrLQW5C7jif7MAQ4XXywMNTMZt0iv1YUy3RuNLtFP
wq6zO1tb2WTmMqLEIrBk5uf0eMuSYmaxpNtI3a3lB5tYABq2MkSZx7ACEMIu
osnjpIzX0yyRzBzybNsv62Afo/YK+BWGnsqZZCchYUD1cEIypXUKdq+LO6/b
YB0TbdpAHPafooMmHyfRFy2ctLRDepaZRSta62ifr0cAEcUWSDLLY864O9k4
SMC3pZp1pAXmYmrDTWaKM+T7p7ND7Geu+u9sPm4pn++DfS9aaaEVx6HRbX0+
olJMuCr8DxkIsfgAx5P2XUhkRq1cimmwiyF9PWDSYssv3fwcVdAMowpXqTtg
nSLRcF7joyWxaWWH90JAKkh+vf/ilWk/0TR0Ut2f2tilB8d1tTfz3XvyE31b
CmFq59+LxHiGVE9It7+YdwPW4sj2hQnMnvDEUyS0nXR3jFKk/TF+qevWG7ft
LP2zWfMhHvyVSY+G7rHmW2QGLvsUzjvLzc/Sek2ALnpjXtoIh649uYxBJqjQ
5SXRbXTMzGeSQ0FxaRkEIJklcCicDQBP/EjX3VayjiVQv3lbjLl2BntBzRzX
61c+6bS85KfcKSFUAyfXquDmBLRL8503kEqKYtfSgtIK7VxK1MNtjXne4Mw9
LQfubSvTvfAsK84TDjyHvPEDyV2QjfOg0H46DixNIDMbWva6TkisdUYQWZWK
Rc+gRTdV/7PNzTRir4V5erg+M9UNxgPfLvjNTNmYLjnYGvO51qZZE9HPbtwE
Ibwg2osOjiwlkGCGgH6HWzBE99FSK9jt58Jw/khE3dkolhQ7B+cKiWuZwvBR
YL0PHDX0c370GffeYSFRSRQa05YhRBTWHPCmbZ/fOzrSNHv639/7SAXzNeJQ
3L1yo2lid4h50o/EAlkVQguEL2zUoZL7AjnEYUcvSwwsYPnbx8gzVH3N5ogR
RyDRAMdXGQuph9YWSb5p59QY7QAZFzMHdQy4jeS/3ZSPp16C7cvRL7lNS7ey
wA1R1wLNzBJWTV7NeUSY7D1O/O0GL9u7/Pxo3R/R2R9TZiYOhSHMsopJN6IW
kpjCgasRVh2YCWeZokZlBBbtkiKwYfopB6R8ECtejmBcSeCVjgr5eRZGlZpL
YDkyCUdtnzkYWnZldaPoZ1HhagiiwSqJrD5TbznpUGd8DnWFyrhdZ4sEd0xw
HQkPwnW0AOb0cFiiyt9CMp4HuFYEFriH9byO2VBQtJG/riinTGFq3i/3Nv7U
9r0UL7xT+5gdtul/mlsH0zoi67N34Sfk9pwvlVN3W57DWx3/U55IXVVdiHa9
YMLCcSNJphoyrH0osY9rNIu4q5nml4PnjqQAVi2ENDtlWVI+Q/N1K09NQ0nu
wNUj3qZp4qPpL5CVWb2OARAepHLW6EnmCxSJfa46ANhhhYBnYi4uOnazK/xB
RNI4Gd75eIhH0Ps1WprPL8zp1TfeTSTWov4BBSjodb0X/wwhDzRg8kK6pXt1
24iKuwvqC081BaBZuArKt6z3LHmWYZTqbUtsaODm/751m85OLCyhu86dE4h4
q+5f3QRZ+mTjFwzQ+gwfqvcYwBqHqAwfwkXNZ02NbqFA0i1YrC8x4HypQqOP
CifaZUhy2k5XHQeWzAJdx39r798UW5QIyFeyPclODAmHd/FrLUWKGOh7R4HH
H3+jkyN6nOEVmEpeNwFPr8mmmSl0AThAoqIW2YB19z9nEXWUQ1z7ggSDN0VY
ptZdouAyIGqacYgD/BEEMRSGqxuEXC4wpKAq98OTH7yNzR5sl0bg04I6+CFm
L7oNIQenKfxEGCA142jqiWMHY9Z+ozlRAC+JwLNb3ynV60W9l6dmUlIfy6AO
KzQyi7jO6ehMN6WuMviuxQVtCkXUKN1iQN1b+U6jBWsgeIhk2yJC49uKswAj
jxn7TColoriJPqa0vqzUxHXuSO9Rd7qu3LWzU64YrUpu01KkIaPPDbDMbPIi
RJFMWkOrn0nNML/quheQTw+MkIBtHGmww9caQAe5wR3XiaixoKK4U/7lL8E/
qbQ+Izia9qGv/iJkrA03GHfa1I6uMq6p2P3kYor+5qi7IXAdJy1ZwjDL8ha9
06xVy5BcSBGhIOAI9O8eQ/IYtoXtVO/vyEeX2/c17d6H44JSw+3axeMAjuP4
MTQ1n/70tp453TKFKNvpibotyWjTZLtIg6QXmDTeFeE2ERdqMhUrRXjP3Bdm
8WwEXsx4pku/MqPvRMz6f2T1ucfMYDdxs1qImv9Dhaq9i2UrxvsasEFRwGhw
PqjCEfIqV9/xd/+/5NJ5eDus7eG12R3MuAe+r5PIbaIydEyJm9BZM7RNKn3G
1pmpimMG5ynifr0nrhUw+PuZAshjg4+Jxyu/3ElNEqOmMmUV9IAXkWh6YLrX
qzvVB7rZCihfOlh47cQvGnU1/2VDNHwnDs3qwvpOIBbMPyg9mCr/KYI9zxxH
njbAUvAfDZdVlZmnRmp73PGTO+ifpYq7aQeLjPIoFwlKChKASEDQsHok6lhm
IgEwAcqg4p0EBJx2yeR71G86iwONGjXJDFnbnkPaMJ+vCIqcCVWqfZlcbLrR
qrI6Ycw0FXjwHXjKc67Cyj/xfZrU5BjkEbZci+TphKUy39S7nAQVIe/I2RC0
tZYD895FYEXcT0nKGIJRPV1JAizmeMd+hIWjM03bDD7Dw1qv22Ksc+nu8llQ
GfgiaR6eCr5CG1geeG2kvhnTnH0NxNokiR6DoHofzY14D+odexscL8NsJEmT
48Fg32lxCo9HHB3O8O8COIMi5z+wRkPPRnx/wgauiE1TW3bSbyvEE1CeC7hW
C7y8hKv16Z8bGHWRzsUt/fPmCQQPxVqOylTnnaCV9nBZLQRJhOUnY2Uu+OFv
vKsFSRCSGGfCxVCzPa1p/Xdfeu0wo8DjsJdSaf4gtMraxhq12IPl9pn0Lqdc
OPYuuIPNBK77nZTDNvqUuNLJKYlv6zR7awgXQY1Chdq4bY1fY7ew1dxuLZEl
Z+cRGto90VItKSXm729yNv/kQdPblMxpVOJsEiDy8KMolic24/d/cD+AshPW
3mIhzsJHMlFwX+YlOCsJMxggeoSDs28kSdk4fF8Y9y+KRb6OZZggu6JqSoHX
HW7u2x1L2DPGnHEc6PU3bLI4mxEls5pbv/VtGZ3KMRW3hK4BWuVoW3B0sf4g
giyquWz3u6fQavTvPzlRKkgHgAkKZ5MqQFDr/LELVFWpp13tCfx39WQYxcH3
MUC8bPqeCwy0jLv/wOkTzxq0lMb3l1UNsZB4Viml6HWFfog/Ew18Zyg2kiEo
2jv6CQ5IdH3dZ2MywIXiFWJOdP6ZoYZ8Wde5i/nRpoOqg6hfScJlQwh35KDB
rl6YB61PZoAd89vIlnXLJ2Ghj/q/am0XrvdKbrSYU8jqFNON2nZG7L7LgV0F
ic/alWOjS162XCNNXp4j1exLYqouGwIv72IOJJ0eMMLCuq4KIq25Htv26F13
m/gncgCBZg7TkS9eOuW+PObsU5LlH0ej+1CtQ397PYcdZ3vMYRLcZdA6aUrs
1OKp54nVGjXrYwazPEbspGf9pxVKpIGrkHaldUlv7Ld9KF8+qZZuT0yiy5CG
3YsbJNDA1RLoGLPiqjbyG/GYn2y6B8a6slvl46UnP4EWaRvtbCaXTzOfdy0Z
aew8iI52FCKg/t0fq46NGcO3IbbVuWID7K4k9+uZFmcmCYqItTDBXo9BSINb
PaG96ze87iKYy0E6kktYBrxPG0i5eeyG9RenomC/evA+hdoezKwW6fyn21PH
aKW5PhyBjBS3fUOmLTVa4jg7sy9kcCiJwB3srVMM/KRwZWQOwj3Bu/N7r9lu
vVwrPuztn22Hd/kQhda7yg9bQqsD/W5PFZc5NL7vY2F0MCsPwjC/fbRQxlhg
jFDNCdw5nzKJsrU8nKbHbUChBqXdYrKzq02/hYB0siauSlXyiu4KNaDKYuq2
y2A8+GXB2gJBLdHVBLBnsWxrOBSwPMhdeh+IFTZ+I4pBy6fHF1rHhAEMzSy8
WXuKVdLt/tlCn+yQxCQtzkSbHtHvxJkSiWgxDcWwr4xj1obc0gWlvKa4gVkj
gUYPrGhzrjSjgTvLeYM+F+pDBZSCoK1KfH7e0EnEGLoEqpKnenj9vuGFFaR6
MNJgOdG+Jh55jHj4F4t0kXwP0GvFD9C4RLjAsaYOhmNXuzVWWi6rokdDejCY
dgcUxWYRob8Lw6y3WZHEqAI35UTNH6LvW50KnujL47MWLAq6RjhjrlGv0HBP
Rosl3EgxPrHUcGMt8gsqQWUTVsRypGB0hTvQbM9IOyFWK7+7X/eqCa8f3xHo
/YvjfCbywesvvUo2DOpuVBJT46BcrL/wh+rLahO+LLtAWR82C4ExN2JKm4t2
1QkyE0LystHjo4a5TV2Zz2CPQuNwDUtSBWXlVpyCyjz0vekGdHcNBk5oKfFu
DWUTL+BGnDOHAzUQs3P7pTWGHXXNyiDt8NW1DUgJL0TNAJ25Ycz02GwP/NHm
RsEFDl1xwDf3dpZwaD2vDh6ZJ9kCulSYqDKpLExxN9XpiJjbuQdovAYfo0m1
D9c530FA2K8xv6nxdDp/Phet1lB7HzUa80Tn4WH+rOKQf73Q8lI7BcwSXMjn
bun6lNbt7oM/UTCM/CfQUG0fytWNxdXgwFY6ohRwbywjgORHKLvVu2T2Z6yZ
tTyomHNZUSd9mnab8GMy6ZIElsCZXfmDG5H+M0LdnFUK6IqbnU4E6JKNaHJD
SVUSrV7knL0QxfleLsUvoR1bFa2MrX0WOxakD3xy21G7XWSi3xzckHCVcnst
9QVLX+b/ybMoKFDch0GWOuKmP3+EagJCBGBqM+Hgdo5I1dfmOX8DecNtbGBN
Wru7767OT/H+3GD57X4F0BDSb1ZkWB15/rAleUnELSpNnr5KNCwwl6/g0q6k
9veuHddy0m/XWsyUkZR6PzO3d8soIdanJFTuNr1vN+0e5VqoEUqSc/bHCqSY
+spe1ZNxVkPKU4iwsKeb23x0k5EoD7JYE8t7FN3Sm/BLVP/N5V3JniUX7B2v
5fEH3DG1eNmfUbw66C+gpAp7Pf2MKiEpLSYnYsNFNXPnCfyEhSXxBV0SxpZU
jZjzHCNZt7YXf5VHSjJ1ALHqC64q0SQjdT/XIeWYJHhRFlcGUk4JHa5PdfAY
x9ubmTJREJ/7o0X0tRO9ePvQKUrMGtqWiez9nNQiueoQ2WcgPbhNRpow+CQ0
sl12LYwgmu4PZXk2CzpvvV97UBfo5u5IR697uXLiEWd+8Mezefkw3CX4Unrb
TiJMmIU/3YJRGrVpb+U7vkm+nGiXMpDXxut99dk5oZf/3mi/xh/THEZXmUt0
Hd4a+KktMAUV8bqh8tLVBqdlXVhNj01Zv8bohukj9tay2Ukhy4ZFxmbonSAi
zTpbkls7KnU01VVPYlbKvVyPSnBqfDF8TMdzNn/LWH51YEndi8GUFCvY0iw4
+T8bSEO+iwkUA6zQ1MCSoFnkTiPND0Vd3zIS5tzt2pS1nGBR22LCTdlwS7E9
G7uO4JU1XuoVQGdthsRzogK/A6nhRfUS13fa5hcN+Nl8Y5FGhcjLX2ntq4dL
3qcgc4iD92EZehrhuwtetoDLkFjOyVm83QUd1n+KdFJow8FDnnvlVDWgSKnT
/4V4ulusx6EuM/bd2Oc2cibNktYX77xbEz+NSfJDVtu2wu8e+clnuwGCnVGi
uEGcpHMLkvj3ZpAlf0aQAFzNW0/tLUl2y+DuZ0mIHnpv2eIlnd77GmLvdXtP
4SpMtnsjaqTvUkXN1Sn5lqkpIdgV34q8noK3TKO2amOB8fmevckuCIflNX35
Kw89hDyT9MpBD43rGtwbqE15YPxw+LZo8RekiqKK0rzgXdw7I43XGfQWFKc/
xq+Y36mL1OTkVfcVupzDfkUZi24c9SwUryvB1f0rv8pstRnYbbam7kbIPf3y
5MSp5eg22huDL+rnMlfZanOWccAoX/lVGPpQiKq3aXnF4nb9yrgZfPhnE+Pd
1pmpYpso3U6xIFHCyeui4nlYdRb9YfIzWIjucdlUCrrWWFNxiTcpJCQ9jupa
nZgLsYorWRu0PBuVgl5uifavjD+PHSfKXFSMLRR7Na/7qAZAHgTHiWT1EPx+
RtZHDoPm27PJy2qtDmx4P08mgU4rb39y7/ujQSkI54dRr5VjVo1AASN5RAZt
Jg92wABq0f5svHHSOHFkMqq4iB+vMq8OBuY6IeL9SU2aeNPvlmmD0zDV1m5d
ZDmJTsiRxjoS2+cIGXDVbpTRqKcz3tfoOoXZJjSxWPNZX/hapYN6FNm4jdVg
EsalpxjbXuEx76ualaOKezMG5uVxfJDKq81nv7XuW95vspASdWKIbHeVNItX
GCcDehpcAKDbmqNcKJo7+luuI7i3FdjZd14cw9Dz+pTXvPNSpqYBvO/o9Cko
MgypgNOpFXCNIO1cAY30rPUl1LwPaZJO9NrJkGPE6RgcekW+4knLz7nDogTG
5q4OsfQLaQHpdwxsZcwhiFuOwkXFL25PzUJ92EGQ9YBgQvyW1lZp06MkInaG
P2Wb4vXFEyOY8CSm2kK3zWTt9n1J+V9hrZp6VRBtixCPjv1G6UE/Rw1i6JQJ
O4cs5t2E5p7J+9TX7apcELN5kh+9wgvPNg5dx0B9eT/bEWVxthfyf0DhMxUW
hIvWNVcm81b7fmwPvFv+4WZCmCzXgX2clzvdJRbGeurG7r7BWlwfZNnxLhuh
jM8Gnn2c3ooJEESQDfeee1kqqvnPo0Yw/YjIWGaFIygG1U2+59RXeq0M7nn/
mt0k1Msdi4nRjgc8C+IkidjUclJZHeF3+uhrnNrs+0aoKwlmA3Qeb8sKDGDT
eWddyhXgcxR59MHChz8d14pSkHon0VgLCiEqdMMTy45cZKF4vk//kAWFToO9
OBZ4HZPOoKwXZNH7SvXZIEZBq2YEGwWYTWPZTYzZ2/7vyxFdn+OIicHjs5db
rxUL1++cmRxFhijNwFTWMmnl+1NDjj/QbzKSPLV9yTSMBlhe2c6b9RP1gldF
f6xhLl8NB1XfnY4QS7gFfWXDUU1hLKzstfEfISjhEwfdRgWnCeVYCG5akAIK
+5gg8BfRzGJLS/5I8lvGVpS2wLeSPDf2EFH+jwepDrxHsNEf5KIpXx9sF0b8
RRAnuBaXGXXJ0wN5Ddih7CZ0hUyaPYI7oznLDvhEHdCUIvhAy2TApNrkPBYq
h8eensMC0t/eO/8vm/X6KS5hxciN0sWsgJaW8hqfB6CT0oDszNFuWXHFoQ/y
U/IqZOgwpM+yKUZsw2lGckE/59XkInOQg/3Bp942fAeBrxAnS3zxnmsN9RdV
CFG5O8QIr6WZAvYfO1cHILowS5ib6CmFUnDXvpFZxTSzeXctEj58Ok4MImVN
U8BbECtlCsEcr+/wGmfEud3WNm4tOa60reAlRVfT3C5tAduKTfLTXlmGbZ3i
nk0/YLAE3oNYb+ngbb3QErFpybDlnfMlcaSNuZhxKnJ+DExribRJgyOMmbhL
KlR3fyJ+HmEfTz18tYhVIq52pg/43X/sHDZTSwviyoEyf78UncptFIIX0Lna
RWtjbVKDOqjIdvFDU4tKFppITzhbkV0rrssoAT2WO9BcGHuIzpvMiE35Xs1z
tucUgDdTaP64wFXDm5jyRn19QAZxuBCCAjzmMlZGYdQmJqXldoi5Eyd5MjLX
EhzJTG0pHbPTtjeufXLzEXI6GjomtB7pAMY0zYyanMfoa1Togt18kP9D8nN6
WPRfWQn0mk1iqTst0os/x79SGGQ4qLP7ZEQOAFVdAKhdaJWavbTWn4Hk+KgO
jvIa7ghjqqgBtmBjt3B6Bw/m8prtjYiA+J1KusxWobBrL+7EYc9J/+MMoCBo
ndAPIKfZrflii6ZoIh5TIBFZwBsfkExG5S30veE3kQ+2JDDcgrCCf1aLb4o1
COMUsJ43Jwx9ws8QhHgl6Hq5USrGNuq/g52vNrRG9T3XhBvcGWliRtqqVq/q
3IlEPdwg0KpPj6Ci97YxQnYLyWdQr9ckCLTEsDO5DOJD+jlAtnt5JOVoTOPp
rKhgjMD72pFiuO3RQTT79hueDG7adHaJ+g4vl1oBITI8QnyxwwtW7cXFu24m
nCV9i2nIiKqxiLB8+jArNuI0zgF65c6ri7Rqtp1m2WDgU+eJh2FfpQleSI8C
HpGqBidMgOpxEn1rYCiWe8XEU0dBTFbhUbk7M1PEZQsUnaT8TvXTQOvIV0+6
cnIk8LemYB8HXc5JRPkkI2fQxZ9icDQLUuTXt/yOzFn5Fz1iKJYucxckAmmy
ORxTYNKr16fhIeMLYPU4U+IZmeEFiGo8+KJDMLGSyL5x1DsGT5x9MWxPQY55
Uz5DOb4C9sYvnO2UssiX3q8fayrYwrNtNLtVw2NxBF4KzEyG/ACaJSJqLQz9
4LUXpnAEgXC1QOaVvYIPsT1wNWLcLB92P608S7RtzBJRlM/1QugCCgdYVM3s
CjCYcmJXYmza26R8Ko5w3K8T/IIhpatGvcArwFi4rHmmfHX2QMfaFw6QhScz
w1r5Usk3M/T3igZzlGE/QWa8vHjl13576pPCfL6J8LCBuXpGlfpqn9SWIBlw
Z9NJEpiKqFPIG7jPGWajaLhuIwb5QzzCvQ4Wl9SYlEzsFuoPZqXtvyyEdk8i
WrTAEN+eM646s6sv7AuNNSBskr1MHbAyB4x4Kqi2XmHXX07P9aOLHpmq75ty
SkS10gAwuchabzM9R65VZ6KnxrkgUGSjpe9hv9hclMSFl1oskBHVpBNaV2L4
BHz9rI/C9Tnv2Q2tJ9/cDfa4HS10SY5uk37sIeb+S0PgOHw81o6YNSqvpUiD
Spn48l7bOE4ZFRhSctpnp/HPBNnuNPB2NPUBKFq5LQbLpCNEELF70+en9J00
Kn1T6UENtHr4fZG8H8WPHDt+s39izAhz8j7zjfa1WZcJECWgvB4RmtLYJeOe
n4kJ0BCFuzwbl/VX4y2Wd1b+S3ufFs9/5h8PyARkgt/H1k0mZJzJlUrIxoIv
D6f7Zbw9Z7SIQpf3kkLB90cEK5Js3Srlu5hnrhUPXjbbyf7A99JE+pK5k8A1
HG7SQCzyvuMTaeDEgYqt2LQvNOwVxv1B+UX7XuZmTxQ9Wdr/kZcVtrnn9LCY
Kvf3sWogDm61lYbtdUfzrxQj6iS5BIgSD30X95qQ4LOGpi2EuqDyt8ql9L+Z
EzGIEyKr5dsIyCek7PjBV1neQTE4PGCayhAhmv4YYxNFhegAwyi3JCHI3LUk
bUbui+h5y6BMC2wbSy0Psidqi2M6vDjZtg2Wfk2J5ahZXYVLrWtUE3N2GURL
LfHnfJnK6pAepPTDd701IUIxsCpL7Ci+QZEzkfwjvD97xVswj/FOViRD+5eo
+doHEu5PUILVH5lUZpHVZdGx/MnhbmPXWMJ4NOvB12YN4LuAK20e1kq8Kdvx
+LXeky9+ImDXs4e+/5WIn1SOfBAYQgfDrL2gUdlDGovqkUMrvxbKX240mJRu
tqLsQSPCwC+jjm3oogYXNV7yfYsTIW4ZMufyc5B9xlQdRHR9BWVxCAF8Al8u
H19nIhdvDiBcDANVfSQQNL6pyr1XwnYno+HLuMkBn+Tay3nahHjufTQaZ7dF
kuOpnJqhDn14Hs5debGw2yK5nzNpI60ONIBi1w8hqH8k+fUfp1UUXtH+KZJ8
wzZPuqwTjh7AFxNASVfyZbVXuu1uIg0Z4y9TMp1RrPr3NsKukx0uwRh916Z7
fnjz48b/G6mzoqurKEDJSNTVFNFUWBomTHAGnicFv4k+3hGfn/w27S9otvFU
ONKEojCgfTQxKqHbRvB52NF/o446XDUNoFbruwA37M1OPYmq+ru+4ZIu6zo+
Zh9oWKso2Yaw6NsmKqOqkYM+/CCc20G6Qvy8tV0Ln5euw65gOpfsypYjVbqC
1zaIqORMrZRigYmIrsVtVUoPzhk55/uY99y7oEboC/SJUC3zqEokqkHED4zT
2z+owwuMlDB8uPgGivviEXyFHlp/Vgu0vZl56tPBzruHzVZZ6KEgbTg9Z7oW
g1s1n6j7fXNDcOLxzM+skeoQ++/F3iGtkaMzNuxAwwXfEGbgnY3u1za5LPDD
AiLQ1s47a9vG7E35B+SV1onSR5eMLsM6SlvlocIYkszCfxw+idSP5GQkLLXl
EaW/c7Eg8qo394g2NGYMkYdZ550MLfN2d9+gu3aNa0KaWzSqWG6GhSlWgxuG
SWkdYHz5D7mMHTsk1kleYLFGi16SI82JamBvLiUByWyuItL+uaH2IjGzbBOW
5LGNNDfqov3QK/ILRbunHQvoecld2szNHgs2UnbyvFk2OWIbY9OMkHxehs32
AiX8mO3plLW0xYNWw3rn5XA6OWfCc+7pbTlZmJiluCWVcskk0NlhIopq/6LL
x5Js6myVtiJ/FwzU21g1f06txH2LlPbJ2GtH9Q/dG+ijOprB7n9Bi15jog3O
yb406DKIBfjfUW8ggsrK69WNct428IbFPWShdjzJFsjo6JG9oK6OR9ppxQTu
fsSqmSviH0stSmm7Pto+PcIuxTs33VHY1zekC7YB4adJyYUcXq58g4kIVB2z
y1o1TEvGIgtCIQHV4bGZRjWDAihfuW1OX9nlieGdJZo6O6vGdy1XqxmQgo/E
cUecKmd6no+WNPtwj2JAt9bsudA+XHdu1jrDFM5kdLnNnzq3OvnMZjLDvAh6
uqBC6b7tQo16w4wO3fGPdgadBz6nIIu1jXME125zOzMBx3vXxhsK9K4gOlPj
5re0T2T4/SsD1g7sHmTMyQecMfx3rWZMctBegsv9lEfXc5ofboA8HN1alyTl
xYLkJQRISCNfLvYGO34uKUiCOfbwgbkBSPGetU17WbvUNHTW7sKe/XH8ilyI
gDwiyriU4rNN4rSUidZupglMchPKBEjf0IsLIOe4IVQFvvD47wvlhUQ6TGnu
9tFgoKGfjaE5QOPOgobFB6cUNQ9VoDWYs90aXBOZYaNOYddGENvKznCqW2wS
3H41noRNvuPnVDfn41zPjFOVe2HwfC8j7RzcMvdSkaVd2WJj4B0eAOaGUeU9
an7bTRJebVb5d492Hwu8S0MnoN8B4nzhQwqWyZpZNmf27OpxpybdZpyyc6+n
AX5LP+llrC7tuV928lwuQIe1lhbDnHhEhiFwTKZlOkQevxKr3jXsIN7zZqvd
i2L8F9NeF12H4XmopkX0LVYSXYxJQ+35aYKupOca73oh6kVR5iVJaOZjjhml
RzQae30SQbAVtOnDOS3nETCmqmBAVMDW4/1eQL0b6TiTxKdo6uwtoGcHLPAn
z2lUnG4rHBULgLeq7qFnGwsgEKkC73Ny/pnDgjztEBTkk9Z4xPurpO38C8hT
g9fyfo6TO7HFLWG/Ih5i9UfXuECElpemaMQTj1SxwWZP9Tx6qOJBDMbaPCFM
iWio70IG1lkxuMyjfjaQr3YREMAMosWJNEFrL7WJouw2ITtEv7J18yfyhXVn
qWhE0YIlrnhAqRoZ3e/naHV1V7frDa1WWrqRhBzidylrrjsjI4ATaUli5l/w
IG2zCu3ntIxxL43XNJ0zTXEn8NqAil0iKzNpShc1R0zDiUtwZLKiGBNRQ9hP
CF5CjnIAy4xP70Ow8Om67WZo0C8FuHNKc9lPuGjaz5hUKTwW//VJEhkaVqBr
73FuxwXxOOfET95bJGOOZ/NBGZUJYXUZq7SIkmZjKsUANR0+zwqDjPbyuLy8
ePi3vpknBqjCT37l2KS6xvKPDqTJ+K8X210gvDKQqO1cKiZySaUvP8j+0jQk
pz+zEdv5FiN/FtBFlqqQt6tPEcmlRDMgy+A8YejWmUv/GW+g56wP7n4rD+OI
G7Br2LC/ZVw949tx4PkGVGASLxip9JCglNoG82LklDdL0+kIss8jvXnFpBMR
F6PiG/qROvyL8tJCj0FtXAZltSuwb7Pgy643axBi6AJx4hNhA71zEHAtLiZg
62R8m3mA4OhZ4CdY7OuYr24nieleZ4sDt14tNhcyJX5V3CYaTzj9YkypJDGj
Dqb9NHwmKg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzcw4hvQiT0kdyw1DICcrVjqaM/PnTizg+w/czi4sTEpwvmwJfXxK314CCBldyaFJtButMJ3w/rL/LqPQ6VoH6Lcq8pOYVsVitefy6jusgM3t3RfspoUNke+Ui+Y8h/sp+iQSD2wRIIHNPVuIb71lARMtwzKGX07/Dtmis94FOYVYzomouiP4+qliSVxaLuQEvtESz3Q9Eke82nmUVQKbgswRGFFrZMYFkGW4YchlfKDMOd0Vy7TxfOPSNfBwPxYPItbjgcJCIZu6zvC0MjmruKx0Y2Cnh76g3VWVMZVlP1xJWm4oUXG6T74YjkUlo101TPL0xLt2e38uEBfyCJVjaImB+1HIusCjEWVJyTweOK311OUtMcN3lsSSbkjoTz1o7s8ekXQ7C2mfQUSUlpYUsZ/ZeCIaMpSm/lGHAKvVEZ437aNsnsqoZ4uWY+jY7WFKuREHNdn14hOsGI5azxct0C8rt60dnGqD9fsfr59r0NUzjpZtxRWgcF3Y0ykp65gYRhukkjOa5J/5ygtEETZa+6VeNs4zkbkKV3RLwpDS0o/sPWxqYa3qGf5m559Ji/riyRiyyJrZ6YD5i6RROtwNq5xC/x0McCvIPfgbvcORGbupwbWzYuozC0DwjvgI3jJV/Q/3NM8Q6YRz6onsHxdI79sVYb7uLWKB3QAGHAOfKq9UrudsTZUCD7IlTfuo3NfPk3Kyk8qAs9JwGUeZ1ErvL9dzB32X3ITlAk3AyrY41cnQY+/+l5pHMNAo4fVrSY6NMMpRitT5wPqJJu0Ceo+j5d3"
`endif