// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
s0+OkWv2p6Yo7GjrfO9ramGHCb2KaRGbf+YiIw+kSIZBNS//KlI2ZcfYckFG
U/DCe7xpJw0/rDkPKYKX7UhSenzq99Xy+koMFglhWQJfxq8b5EIrW+QeegN5
gTwt6N6a8bRlkjQkafof8HHktfCbX8nCxwhiYgLagr6+iLDZhOke/pCwaNML
LD200/YyKpPk6o+DuxcSzoxUVDr3ZDc7gFpXNkkfFQGvwfX5zfY9a1sPxoxb
7pMABJKB8le39FxfecqS6JzInjZjShKGZuLth2r/WpKO5RAbvBZqtaAa3WuL
u0/CGnuno5IOtGOpOddRD4fP2/j//R3tDpSLWgfaaA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Xared3g5Fbz+HeoYZ8jio9eN6/31ifp1LAORcmESb9YvpFiEbwEe3t4J75hq
qHfl350v2fB8uEbH4N7hGsVpQzhzHUOBe2nhRN/5itKs1Nr+iVPaeYBqctLR
8CGmnV6G3JMGOXSjVFysTXWMCRe0rZXP1A/bgKlYXK7ZUsrmSgb1wz8NoA38
tQgBSJcM9a61dKodCI9ijuzhlDXCJVAXnnuoVNJk+9lfvATfJSqmSFloqYrE
JTnI/VnIqZcNXz8YrlMo1S6jZ5MobvzXr13wIVQPRC84w844SUu+eKtcdK2b
Mh7jM7GrP6xnpzw2m/e0FLwjtRauDg6pUU3fyHAaVA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DGleHn9waqXOCwyJghko0lC4JMJTgF8BQxw/amQEA0cYoJgxyz+zgWw0siEm
4kq57FFwsUL0PBjPTkijiRWtkPNq/YlfmffClTZxTlBeVj7EEaxTuD+LxEn7
uMa8/q+laT97g32//BISXfrDTfgahapfWbLQIsI6M+D2aX0yhnj+AqXH4U8q
Ij2PDV0dfvd3dsusYJxn6Pc6rT2nehOT8CpgFRGpvUuno+bntQYKRnRMqM24
/1RBO0pL+gB0iBWWmwRckDCu83Xn/NYYf9T1BQrnbksVDD00Pool8SfjEn/X
3pCelFWlRjVjeG8mq6Ti2ctmGPAJDjm5Ea4Y5L9aew==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TDDQPsSNNZef+fJi5fhzEKqELbpUnpuYunf0Q4p8ffv6/8R657hgZJtbd1Ng
LfK8tEM6+FxgdM+NieW89tgFxNWl6Ap59T+ZgJ/BJ6rYXb6j+BAdOcvDOQYV
uoL5DA4bF1DKmRb8EETbxCArnsuoe/DnXklP0kQ752Dd3xkqH7VDMYPS0MRu
9xe2fSepRdf0g1u+1U6JxpGeBomKL/KU8n3NnLhmt0BDKcpL2D0yJCdR770f
CjR63Y4OLT4ZkIQVWi0Y7KJbeA62svHr9cOc3AV8gwqQTxiP6peYBts32lf/
brcR7ik9G/Bq38Mfy6ZctfzKZRfWge1/L2lAHdM/Tw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DNfelrtRztwOrLkDAvpf0CSv7ua+kwv5mb9Zgpt9rm7HaNl94TdADuvLQMjy
iDvPKgv9cVNt2U8IXAGCE9jOAQZYOcGBoUtwSRjaOguaJ8AiDX9xJhbrkXkV
u5dTgEEFM2hCzoH1WRQFUUgdSyeX9vNm0ChWrWSGsw72DV4DRkE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HCxx0GO/j4a+/G22qFA75dQiLSw62NDCG4aW0yPTdks4Ef4spj94yhMZa5/w
nEROK2rdsGqW83rJJE7D5XQIvOPGR8rcK5cxdBEdEkbRa8WyThRomhGQTnEw
NBoStLBihSzRSeSo+I+DJS9yANY4yoxfS+U3zQzRMtFvK6mlslho0x1irPAi
pem3x6TZdzYOjdCBy28XxZL5GxPIGVwzNJUGPcEu9bDdr3hrkAj2b4z+vJfQ
6GFxSTYn1HHR/0qJc/C+CVwEQ98vx6/XtV7c2JIcbDfYo1IneprBXqM38Dll
mOHyJd5BNJTxq6t7Va9KLXM9nilEZRJX0Ju4uhnQbqMM/0TgLrE53gtb2sqb
69b6lO7M1CW8QGCJUjQIG5RDT8kexDo9+ZaTJZDJsQdbSTRGEAZbw6wpku0M
xwH7FpfrbvRZJUPP47odFXO8sG1O5IJoGPOhaJg3KRmS6EFAb1cEPFy7CI0Q
YksRsiiVtr+LbZj8jPkwmfiBrhhuCVXo


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rTsjacQhMSdvKju4T22EAjbczfbaXM86kz446YEUkVgHW9NKpIOa2Dx5oboV
FO8u83KAxyPUqxC6ZG1QN173HWzCjscK3UZJRU2ZjnBKJbS6c927w6/rx4K8
rC3+s0Xj3Fu11U7npOkSheoPRwk2wjiFQRJLMpQCdE8uIVGkoLU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SteTzJ69CO3/+t/Y5H2NAg78it8qGWNQvIbOrXM+nnwxMPXVkdvp40tTWNv+
OUlPoSskGudWLPt1AI+AwdyDTxJZsvZKw9M4063kyXJq2RAnl1yPPZGViPhk
TLTQeKZX9IGrBo9aWxi7rzhNw136a30A/52iUQcYSplt0Q9QiqA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11552)
`pragma protect data_block
YXdfgZsH/sFePQJDxD3ETWbBTav/ogLqIjkEtVLIQj3wS2B/yLrEV8xZDThv
8N+FOaBIExy4BDnvhXWDq/zJ73EH3t+lAhv2PywtdCJeBGhnn/oqKFTTGojF
aajuJk8KeFC+wuHcUtm9RBHSC7BNxq4a7AlFmNwsbDl/Er6Mb7Z92lCWBeBW
sE+4qxNX7gF7H9BiRbF8UIg3p3Dwen7cA89HwxZx36l/iqpzoY52oOwWRcox
vsJppb+njrk65KvDorMY457LevaqW+4JsG69bEu2A8YuuasiC/y2w7dWiS6e
XnW30WEg+0uJfUVekgQGwbgbS62mA6iPbfNYWW0HMB6ybPPHHUy/u81AZHId
nMfKy4Ynt9u8tqF98UJJq/NxvvECIgW81VeTMzzIVaJjVWCzKzs7cViUJu6z
g+NunvY5x0HgEtr0sg1tXxcwkLrK1wr96xqJw3q8K0pzxyKPQafzWkCwk4CE
lNgGu9ig+qLueVoPZZl1y21mwAnbEqbdoZGKOq7rg/vqZ3WkqjPFRH/Wa/3I
lez7AFY03T0nbYSuhe0zRWyFf72MTbWRTAMBgv/ZY3iSeZ02VtmOEgde9Hqf
Bq24BOp26STfmcxLqzyooIPWZtYkLDWct5Zn+Kj1XfSop8LiAaFznr9R66Zr
fcmoLXIfY5I2UH10kgLyl0/zDaMfPAddEHz/wt6L+WMuryxYAaSu9j5ZyoKB
BVWvpF7wwi+/tUv+p+bl/gHiUGntkfu/60/j6ZyhEolHHD+eFyqoS9XlPUZn
N9qcCVQRLrPcxR+IsTOyOrDeA94jHm83E54p3GVmXSrr7K6LvJq/Fyp2fNXw
/9avRzvJa5QF+3PtAfuKDxXlOOPpE/flqgbSpNJ0x76nKCt8DixCdPDF4BD0
kLsyQbZsh3OIKqpSWIRtPvWUMhq7zSCXzO+ZradDQ8wdySJ7JVLmmPcP56x8
ncmghagLqmIbXNKMwCwzWCBK1cDch0oDv5RD5CmhuBnHa6GN1mQHCVzsJu9n
+nOGAQDf7lb0L81bhnnTRt8IGNxY96sROG16oS6ujzTFDlLJFBYPOKcoZdV9
jV/MmyqafJuUvF4XC6tyXYBomVVkRNgQAUJSVT2iQfJAR7k3GIhJ09ZWsZRR
7SUehYAhS/DYTz7C7i04a9cKWkqVFaGhmbXS6VZ2zSP97eFockONsqnofNna
A2I7LU4NQJj+pz7wxbjUrRPBpc2OXLNgdQFzYwLHyiWSSivMFGBhb8YbvMDM
1O/VM4nMJJzONYm9DgH+G41SegSep9c+M6MTRX5kyE+EF5q3REKgg8/4IyR5
njMbbwWZse5jbEF7cx8L1NIyN9Kg9GDARKPvvsehRyRmxJ6FjN+amzW9yzuC
pgvp93p8Lld6jRIpz2ttsYWb7D6VV+VmKe0ydWkc4985A5RQy+wQHFionj4d
3SReU92uQfu5o6gMaDHrOn651goq9y642++3aWl5ALG1wywwHcVPKBLuP5ic
VCxfwGnnvFDyNzDDB5ccyczXzBtWkkSbpDPH5Ks+BtQtQ86/hEghdtD3O/6d
dMYzEi2WoGsmKFb95BloaDR5DsD98zhNQOzu4rBIxSjjr2UsyTPQr8SJH/0q
hBvCiEmT3cy9qJ85iCa98YuRdRovqDTyWuHXM8HidPRQSJDvrMMnG/VunaBZ
ftTu+Bt9H2VE2wRyUVJ+RVPMg1t3VuDffpmp3scyuyNhQYZxSu6pY4C0shm9
etfFQaVnnvDF/OxvLSZGCpbKEYrervCJGoSrZr7rTbyhnSJQXVIs3cPdc2XK
4hmAZ89ckt1ygyxYyaOl9XQ1w5uVvbU59GWUWw/mBDhs6y/lrxSHRK5AKEXH
7311xUkgHZnow+euD1gx/puzEoUiRxssg1SPYQ/B5YQE3ewaAIaj+ysDciM5
SnmF6cfYYDAxSa1LSzt2zV/lL/A/M/K5+ckZajd+tw2AKIAN0Y5kWFrqi+Ia
xnpG7NckOzt2qyFMw4vs7Noa5sCwYRNFW4IVtjhpY+tt6I6pVCenSXFh3QxX
QMuR6IWXr2LRW9iKNyxqRsfSu0rajGgOC7UMdR9/TF9tOfMNnoFCJMO4BPhm
0NogV27O7u4GFBI3yiPsWhNAah4/aYyjeJFNKL77fBCMpEFFQyeVA4TTVuyq
ANuChbgcbZyJYmNFq9p5XcI6xKJRaukD+EAs03vxEhvdrMs39DkQxCvepUCy
JvugVXed1FX6aHsecw4jLxThOhcBT92wJoPTzz4vVuqZZ/23ippAC1MVrP7o
2JhPrTnqoQCunGrE0ZdptZIGp4Tx9NOhbvTuBjDMuRQjBNd1q1xXdRiVsArf
qYxF6HjZwRMgrn8ZRC2uNAZ/m9X5nNu/vkx6ZP3TwSK1cs+McioTRJqEB1Qc
KQzlo/cTLrzyPK7K0cQNI0O90wb3s+UswkKDqPq4fMmZLXjeVqBDRcBBaJCg
xPRxtDQYmf0+OYCwO3lxO/xFuQFucAwFO4Q9T3QMbGcUE0ISL9ecM8kAx/mB
qawTxvYNTGGWOh9Od2iQDak+YPqW9IXdtX7wGB58LCsjD361Hv5gjAtWaan4
dNTCcclJQBZy+YyZ54vVDSTJZoRmaTjiIkv8iM/GRYM4ae95UxTh3kMLzKfI
2ASaIk79dRe5fKKrmWTcdgRI5mGbhFF2nqmTHjA0YggHsMxVOysKOeQZVIFM
6ljeT/ZcX1qBr62iXjixXRTZsD/N9zpO3dT1Pl7Htb8j9wUPMNLeIuc1N5zF
p9O/y0G5MenjJVHwX2UNAs0Ww5lNvpe40huTIbPXm8ASqNMhKbFVuGUVqnNe
+Vk1mWa75fM/jNU0c4okjaLV1XlAcXtUsb6Im0R/gBiBJB4ddTaW6D3QEe+B
BtzQ5Gf4DGCCQgPyPwzCPDb1y0MU8g7WXTPTOG+rbTl2SCxVi1n2oXahONxY
P2YsdJRW8qD5+18G/+gQXrwTSqkVnbQFsRC57SIHfxbG/9VeygFTkPpNZVaY
qG4R1NFqsXvLqyjphsNj8RgWNMtGFupcFwIOyw+UAPZ9gjLLq8wjyimcqUuI
uCD03LIakr6KxmVwY5tGjTFqPAdqOliCiBer9PtUv5KCzcltdACosgZBXKeo
t9fW5Dn/0spFDEA1NeigrZvOih8IF/ejkx5uFWQKxIwZ3KLoYmsnEfo+7gEJ
r+YLSGUBkPlj8PfIO04UsS2sQbcPEilPZunUgeJ0i8/wK+r3uIPWBg27NZ0n
+fC/As7ob6vpb3hur94X1aLAyVoK/js9L1O/eK0l5enMd9a0tXFi3udvagzt
FfWUeUHMb21JqzGq/Z80SBhNQM1K7MaY9axqFOQQA4UazdG85NIz9wAh1YZr
m+dcHn5Wz9Mapsf+pniq/PgZOSkuOsIxslCpQ/XFbhm2DhVXltRJxWCVO/aI
9UquqQD7blrMxmRtnnOb+3JD6Xhxk7F5Z6Qp+D+LMJz8ccQdE8CWjq7YdEM0
m4bnobbokEJBGtGhsbL1wV4oOFhlgzjnakIpuC4BIAfJlpZlCth1y9N61Sl4
ybmd/VRnff4zpDr+9peMOZM2/hQLIu85OM4suPgsRPos+uqfbV9KEtt8J1tf
EBID16jr6LVosjcsLHl0TtGih++9U+s+ElGuhpVuXc5jCV9TZdWesRaV1LMj
KpQotgaVEsFeNmTcaQ98NMt+VLBARrP9L3xc9c08c/uNAcBySDsVFjBhIxtb
k8mu+t5/240+APnt9Uk2O9BVXkyVsxDa371xbxDyEAudfaqwLBviQ6eevH40
b4qEP1xdsgp6H3SreKGnlc9dYDD8JhZAzl0BboXriRDBrZMSJx2rsk6wu5cJ
L0dc5ko9C0oyMF9VrLt84+cw1eVChXWSccCJptiRAoIpnFHpPKaKNtAvFCIE
f8kvFMPj6yeknx7e/4MxaVALMozfhhiLuvhmVt/3iVST1xSOjqX+PyyaEJVj
eNsRtVHQLIp7p5s0Nj9MhmZVHw9zvqHdK1NReFuRbM0nTUXmGDGD2aSbmYzM
ntpys9BKRGCZAe8YEErKvoRvWBqAsI4o5hEYhJxZPjkeZovhcZYwNiNqaLgm
I7giyfx5gvQY/5g6wt573DnDFBVslKyG/g8fjZA7fSQzJRfsoPV66tQm+dC3
7glZfsFt9IjQcCxVmz8LUKM+oOjDYTP6ZEQ2D/HN2Mmx4Kg42e+lI0OKaI9U
94eyyaB/s2WBrj9DKiEomdypHdBc1tMyw+WlIBHaUCo4wqzdEfvdLQKx5VR8
mMGJ9NT0iaRZMzBHbTiF+XTi/kovZyAeEhwD/tnxAMPWJJvLE3bmCspSxkM+
VmV6jgqm+7PYcw3LuSUKUkDIUioSgX8Uc6Vqb6qNjuQjuuyvsoTK4XPZHx//
2KDrVGbU3bgs+Jw2HVFflHUWZh0+Sm2AIdDFQkP8nsLXK2Kg+RAkvaq+Qcp5
GCd3Wu76quVSpKJ9nh8i5jAtXzAvkmeIMfZg7TbLeTI/7F4S1ZvidfAGOSff
jgTCxqfn1wkDYGR6PdMnFsJMAkT7RiZ91qMii+XH+ItrB7SoDMj5RjC8411/
MP9PNlAvpMCgrzz72Rn4UkUupeQgm59nbPeSdBerCZB6tLv7BjvOt36fpHVm
YTsyUfAemaw39jFPKdJsosOA2/Vf1eg17roYkW5DjedZw25/k5vYg06IZRAV
Rtsy/kHKmNT4Eoo68TGZVdG4ERFd+WwQtUQgtpOLSLYUv3KijBilKRwyUn/2
VRkuY3pXKlMwknTRLVzBzeoANXKNhJDtvTdVF/yRNgQuVirqiqqQIuaIhgvu
a4NtmIThQ7kH//ztoy+mmeQmbsz8GQkv8mesxIxMn29jk/aob9556FQMuU9u
NUzYgSKqecQpRm0IkdXcavj7wsZns9+gXgbUEShb4XDTSDkkvzSfuHxIhRY+
2qW6bYjoQFW470ZsxlSHrTqqvfK6hOLZ4XtOTDByQLTWidC/oUVNC9lHLb7D
VKZM8MhjxWlVHggR5pHAINm/sRxxppB+9g5drXSpJCkMVoJNJmpDV72MLCpz
ofUojq01Gxp9IxxIFe4OBOayIxVL3z2To75HsRaYD0y38YP/xMW9OUnc2Od7
YgtclK6LuCnfs8WvszaOp0fTtbio+r9YGHuFIEGSKhckx1HG8o2dzHPy9jV2
YMCPPO0VDRQ9XDuHRtf3jGj0qrxcP4rK6IKhivQSTp/19Bz8SmnmapznEhZF
uguKdNfJ5GyWyIuaUBKNXfXYPTS17tpBgNa5iyM2EJqK1z0S9zXbV4P3xfPM
JaldyfvJeQA7Ywc2nFuzAEKbr4D4zpDrZkLyjRgEF48D9mPmxnPuv1tXgdRQ
ppZnmQcrKAdIWOqSPAcE5KbKvnGcKyjoFHUQXhH84vqj0r0JDYJdA8yvV4bY
tuUkzjHyVgH5BmEM4N7tVE6r2nEwrpXjJAiPeBT5HwxELPfNOh5OPlMAF6nB
KQnKK0tejvTeZCofpMmUxglCgD0x4ugPjxdqgNDlQkxvDIKVdk1+L+DXfZiC
7SdVgj01vKPmtQ2JoORMTsI0+W/rHeLy4w2XT5hEoJ3wOrqU1QPp77ZDshXs
c9QD270KMFsNp7PAbs1j7Q6rwUQE5i2584+vqB3DaDf1G10x1y0uDj8MAS9b
Dl6y7B479J3whfaxVCQ7cDuqod3C6g9caSVjbhRfLHMmWf0Jvn2EdrSRTGs1
upV7JXlvm8xCC3vcH7LZ6Is+kWAUjhs8PEy66TgGSS6PqeHKKicFq06zeq52
ilPW4WQDXy5eUzZrNXmvfI2nEfPZaKoSSKMZyW6QV/kZI3y5N4kokGtJP8IF
LdnE1XvxACfCw9kCV/OomYPbVOuXWMDrD7UBoT6Y4QWWG/mFFBz3C+Ogi2Ad
swvcQOalEIxYoR9ngfRT8YgMDZuR4ILjzJRMAsmYI8+zzbPUIYecGvR7ekLi
o2wlYs58Br4JavB8q6RfMrYopL+Fjpi8FpqGfe82za2Kk9MpdZWUHCH2JZDe
4pkUQnl5YIwpJGrDJ12EEYnzIuO/EfCre2OLKI+V/DjZrZLhHZQK8EpdbHTn
0j2SlIOD/z7XbqupMQY/cU8mmqNLC+Df0EhCg5GI4bTOj4ol215C0JZ+uy4i
Y2q11sesAtUWBQkMH000VRbDEHXPdhSH2nSke3kI0hbf2V8V945Mhyyxi4L4
QXCekeypDRXpaYHl/3wNmpUtAnsGOHRK1Zg5nXlLhjEfi4sI7tjOmIUTu5oz
9LVz7fCM6Z/pdNjidkbVByLwBOVePTQlCeO72Qkjm5OOwRHzpDpPKt4QB8Dp
UMWDKYeIObrsl3PxsuiZZpvmhSvjaLABFMcQkxnPQ5EoG4aRLQhS+x9AF/DO
45y83RIYrPiZ7sPK7PZZDwNcyQ6apFw/qfFnTKaci9I4V6hrW5NjrkVvyQ3V
f/Tji1pJa72vZ0/CYMDdf9dy81HlPntXPsmHULa/Fho6Pq2qrJ7HKiYmMSuZ
+kTpwHJNCazqvo98Po+NvKuhsvnSfWEWbMQlr4JZPzfQFiGwjEZ99zYTMo7p
Ux8mJgrD3OakjBioJggc4xeiaBeMM9b2SEani3iqMdyBkBR8U/XpFFazY4VF
gLZpYevKkfZV/F0OO8NCVzP7Fkv9/Jh5qbSXgBkuv9JU8HYc5uYgO75A6KOU
DxcXani7XLddS9hQM67pbDSklnB0FFxAefe5Egz6y5WOy8EasX9AH/LLZhaU
LhK2xC+11ibETGBfs7Ook7jvSboTZe2au2yT+p6sh3evvraZQ/84x3nCcE8f
eBBezcmQ+FtpJpS57gLgSRLhT7Sv+DA7jSEb2qKG0MBiO/0j+svUuKmx+BkD
ZhgnpqLSF4ibeTXXh1CbnIkdu5hw9guncHl5ncdeEeE6KTi75St8jhwaZ8aG
Iil0WRxStPEULGl9lEsjU4l+EaX8iRjDZ5fdWwzGOnGE/xepjvX0a6dXJVeg
sziM4Xugr5DUq4UDYu/3cfj4XJEq2xsxKk+aYEhiezahrGpKXfcVMSh8X7wh
9hBXl1cPNCfI8yncfppaAuZedIoV/St2AM4nENN8K7SaU0xfKs6sRIFu5mdU
wIs7F0eaqHiXIctTKa+rgtn4yAd1te7+7BPAkPsqUk/r55lRAE/zqAeFNfhf
AUPIvJszVyMT6ZOo3PUthExKbNygvAbRI7FUHTnV/gXjFKjueVSia6tlvpOg
zLD8Ex/I3W43jLQrxQDpLEvf01jrG9WRAohX8SWGOrPDnFlL5uug/QTxlGTX
gyFrisRu3aDIEoLnsBs9RzKiBjzdKTBatPwiTaN13mFpRtEFeQGdsO+8bZaH
FnKusD+pMsTRfcbf4DkyuPuy+KTCm4XtQExCGFTcLhJGGdwQI8d3x4R2l809
pofIqMWQk+C+zYf/ETOLMxmftT7IA2npvy+oLeNHc0/YKxd88QwNicnu5/Ep
ZVDNAOdf7DttNwUO6z2dWSUjdZMy2o29xRiyAJfz8PgC/hBHtPgqfhkwLR7n
0e2pXP51kMjbpMLcw49RdarBijzf6IguCB1fCqQjgY8wZHagQv4+IxS9/dIn
V0WodxcVJHkjAc2aF3oiEj94gfTsD1IJ9IjRIS6pAaPIJwzkr5wzRkszayqf
BJOv0AQZW3LcXpULmyv9V/WFzoFf0ivXBOMwrCVMo7CeEGUYgw+6oef+sIH+
LqjsKfLRm+e921GBq/7p6VaXBhA5HFq7SJ2juemlI5TfZIRb1YV+hMqbRcrv
7YFGfHXZ7Dx6vc57ovhfPryOZ2xl51XX8bXSuYtXScLP6dTCLCwjzWT/eRFE
oP+JjEtdaHLTSmxRTdS3a49geie9jsaCZui6yq4sPrsqq+lzZRo6bmw463TQ
s3FJvP4G0F+FlULEKZJtcD1uA0B8tn000Do1I4bTr6h1xB/FPWCArKnLVluc
2CEBup3yUi6Hyo2RNCHe1FF3+E3Sw965Zqd+q405BDUHEs8p86yjjT/x4cc8
ih+c5UDDse7rSUG5/VS+4bX3cqQphKDGBdhR1ns05iDm1AQBgqc6qELiPYaS
B6n/LbOvnsPcN7afmxTq+znFuxkg0T3i2E1Smrec/6sBvD8hDfgyVMtxWwzB
SDj+kPKLewp0xd9HxcZrXHds7WqsSy5MTs9PJp+xIcjxJAlUZJ5PrUJ9eFXe
c34QIvRnfD40FcJ7+UhhjC5q6q5TKAPs04bIcO5/6+Y7N/zulZceSbkq/W+0
ZhiUcB4NnDP4ZiRMDAKPCfRmsx6O760ve0tr0hqoVmFPqgDeKo3Vs6zOXcmj
qKLCAbUa6gUJbgUPM82Svbyn+wNE8gu3Tvs90jWH2Gd+BvQ8trNzrHhrlxcA
/RKvT1RaYWrDvSjTTmOSeyaHDehQ6HF5E3oEjeEeRYzYzLUG7YitDpJ0WDo1
LZHe+I45UyiqaEetRa+BQb8QPmSKKJkbU3GoczH5f9e7uGo/Owg8QpXlYkw6
Xr+JTCEVQ3rEr7eedyx91Gst2MvTOo9BOHXUcZPMQ5FBa1r0m8MJ+KzMRAJe
0eTQMuspQbhPfi6ouKk4vvg0VYScwrRZY3AyuisMeUNsGQGyjv1y3dzWGHWt
YrLeIQS9xUOvOHY3YuxgCG5JJdyxkXNshk2QXMDaLEIRB9tNlLp1oTYvAtfI
Gr8kkF7iu8BqWNTU/lRiKFN2BPgXDUHEqYvQn/EaoNhjJvF9Igx5oD3ii9t5
dKMXrVzhArawSIrP1mJ5U5dQDIaWJyrgyLZQECw3wzjGhZB+F/4BR6w30KeN
rP9xKr9twLYu3kkFpACcyEgGNWddcHAZ1KhYRhmUzPR7pu7RcgJrAlcBM4UZ
sODOGzMkjPbkVOzLdb9Z8RF+wzche+4ERMaTSvKrYvriyN6+rd7pnROQq5lx
cvFJGKTQwPJBTV9pk0NThcst6xRZgZw87dCP1wib8YZVkVAZoJVVI9XnoQZt
xfRn7pcU/oh1OEwctLO1HnL5qn/rlOUXRnlvhQdq9/H48b3GXqOF3XKcvu3Q
qCK5WAHElXHt42PMRovZ/W2Pp5l8ZLKkqbAkU4dT5vJY6LEqe8yN/jwFotby
Vqdr0hXTPqWuPo/c7MmrN6r3X+SQtbwLM38w1M76VDE/jOZvHYKx7XvET0Ci
5J1oxAiQkrzW2AqsAx5w2Q832ZxIJTbdUnXjospV2me3CP4DuKdHs/iLHygz
Ej3VfRF1SziMGlRi65bHoqv7IVJ36Ee8lmeyZBGFvzEc7fFL7h6U7GlHMVON
O/IykBYJlk0EOl28Ae1LMrHul9zf7MNSwHKYe2gNccCKCpgC4WJtQaEpCyrQ
6dWBISSa4KesuCHeXUPPhRsF2LtDK8qDy/80QIwhYQteJ/JFQtB6x9qqOLQt
NH5ASb3U5TsVthaaawdo2w5Z+9whMxw0UHMvsOWfNuExA2me3w21yFwQu2I8
bS+mUhcqFlQydctgNzrHUboT731jMwuyFC99nEUc4+BK5MUx1eCymOWXcGA/
wvxUqV8ecSWjYZFrzuk1QFZ27fpF9M4JCWer+RKUIugPocw+yXjvEn0J9+Ps
Lb4ZqoPXvI88EXe5EGcq71DzW6+x+PBsUPzOJIXPII9B8hVsRy0qhIHstSix
4AT/3q6DeTRtfdKLYhQHd5iuIdiEucUMCnSCIbIOowXq9AvUPmXfRkrXsPJW
6BhPAiTOnm4F9zpYpVqY5vlajors7Dk+6HEqVEAqKehSFJp92pG2RoTj/6Fd
XscswnsvyT4uglg2abqbbB3jKhGemM24kIVJ+ymBa8iiD8B0T4H2Yg0W+2Na
ex7Mnq962qR5GZaqjr9wAkK4crTubhhFB3WrnO2XWl6Z3RgW/F/3blLw1lNC
03PwcklsfXOazgLcFueh29/BoUXR2w9o2HyvpkRCMKHdFGl5zqUAO98Dm0EH
TmXJLlvouqRQXNXDE9DXATcP9yrrPJ8DrWan2HMtoCEPlJS05H4mcb1yb4zZ
Tl/1qWNRlihAWHUJ9EKmyaol/rpIsadujUb8pBrdzfjV2fB/fIJMkFPaOJai
ngdl+EaEe9LSOMsboAGViaxXGh7ioTXXQdMS0GI8hRINEYHe0+C6qQ7HvxfD
xXXCct2EcQMT4mvb34Jfhh2PPKc+bg9CKA60ddtj7W9boGOiu84USanXfCIk
d/qTPib0APDrC2H06vjWKmSNG+Px+G43JK4sNk1wPTOSP9XF/ukZtf/r7E6S
x2cEFyhK5h2swG2MzMJIjnjwwLalGnclh8WWtMG/S1A5gbJkL7T+yfHD0VXZ
YsY+1sEIILbVqUDxJk86CHZo+af+bHSLjGHvaeII+uztF9Ih6GLsmg/1tkfU
j+BibBq611KSmkwEOVaYODpYMTKovn1rujF9hTdLZy5pC/WWZnnP/sC3Qbp4
szcPitIjSys0nV0wzpr0uwbjuB+q3xniFZbz1DVrUt4OB92CfsIMYJWGqIgO
Hedtg9atjTF5qsZJoMUTVIKrrWgPyB5W6ruzWWaxukDglr1tEthTTD3dg4fl
SO20qccHXTIyuie/yPXAJLtfjykK+nEBvwRZO3rgg2EpRth1QNzj5I78/76H
LmyQ1f+JmuuWa1L2DGWb13eRBXR2kco5emAqn5dBYvtoomtGjhu4oomSNgaS
fOrM94BugfuY0n+OBN+kPpjVluf5coWOWo9yd8aoZitmfOrAgA6tD5P1agLE
ajAmd0ea6bVOiyWm1cbTXrWFamDIPBODZPtdusPfI17nWMNKN1RU//DL0eCj
4QAL4vfCzKDhJRT0atqfqBKaav+kklb8FB2UdV7ECRO+7aEPHAkfW2X/uAQi
opAcDaHM91YEhFAxvMH7F6oWgkCNh8ujNjZnPzPB9rXw/nR3Qo7v9YE+SXOu
mGFImSuQNGK3ag/DGgIvE2WopcJ1hVPijl25ozLx9gGIUO42I2WPlzddHqTq
axdrEnCLRW8bwyVbMWZWKHS03tA9L6BHn+oUUNrDodE+8PbURjAJg91M/rmO
hbRqwPnELtZWBIjhAu7iMvYg2bk1aTK1UO6/Csb6GjJ2Y6k90iAFp8yhUQfh
zafj6elDRUbuJkl/7Kzv3tGCIFP6jJdrhY7HWNGtZIrp8Dyn3Oz/ZW/k/msq
vK1eJ8Cud+eY7i2mmaRsXvBp7rtNurl43ds95b4X+zWiHm14oCeMhswaSJFo
6Efit8y4pUwO9s/kg8Tl8oHyQzJffkU+/NxAn1mhdGQF5aHXLE0v4/ahKNTz
ilyF12g40iBPwQNQfJvnhvBNB4FXB125PaNxjFSZOse926DDYkkLermJlTmS
uflstOP4aVe66SxOQ3tu1z6Vzxp0pzk/oFc2xaCnyhe5M8+AkbwR7J5Hp5Z9
l7G7LO+F/o4EbThtJeb4MUSo4+CSDcuWuSEKIM3/VhKYspicgJXSjrZwm4t2
8KtyIyLbFfwdMGmHIKziZlSaxzLPi1HxFRNhBq5NCULVmzHntxb44+SwtHHz
7ionkd/PRn37Eu3DMDvyKXfO2NH5WzHmmcsVCEvbNAPExum/lrfc+NkJP77B
HahagCPqmfmP15XFHCn/TzNf2YRRPSxrECsWwOMlfQWxGx+KtBHv8LSYj8ZI
cs8z1gYur4Wl3dwdGRzNKx874e76DfWA8AKaDlhG+alq0qP7DwSRKRASc8Yc
HNgyLoktkNID/xDvXXWNlKVT34VC1vXC5zLXwSjpVcnUvp6aT3o0JMqzRagm
YCySaE1osbiIILbBmR7J7mt0qfqVMzTy7I2V0+/zXZw1S7wZHNIOkgoEbJ4D
JbFNzOMWar629QL4iptiKCXp/Qly7gyB7FDPKiMy+NwuqyDhkqU2UlnpVO9C
7ZxDOIDzF9YxRI1op65Vl/3nHcd252Qc15Rk208Xx1uIjMRwhJg0amAODkhs
E4WmWhsXGfjLei2RIMqsQZ4diwr5MxxrNVZN2BQc2dJ4+w3gKM0PHJ1qHHq3
6mew/+rScQjfMakzx63ve62EJg2BhuE5U5mYcx8GRfO91/E6YLlzX3Zqm+t0
PJBFT6ZoMZljQmQvG5uWHZPTyW507yzAY1aMfkLKX7jwJnzlu+lOIlmxfMG4
dK9fex506BLlnxo0QUZRnGO1Fb2l7tQkz8ClAFm+JfVcMUvKiAa0RavWjw7L
TJd147wy+y3gjrGiflqbyaMyWJSZ8HvupTTFoHHXbJUNdFBWRU9//FkXi6L/
53unqE/c46bKruuG6VcJ+pbC25Di+3EeCgzBYRNIy8yUNSMXksCduvoc4qD9
+HkZuubS6eFG7Oo6lA37WZsd1xz5SuUoIiERtOpKDzbmZ61mrUe5ik09V37k
GIkAsL65W5psu6zNq+CWKjoI2adg+zSqQqPfnYmp7owMb+NwgkOxDqMkWs8r
WiSiyc5A/zzuL4Wo3HUJMArp5pCmPdrc1ibX5eJfhVDD0idaaRy+3GXr5uuJ
TclWzf9/nCPUvtBSq7eW8a1Tajy6W4vJCbJWCYBwi052p6JbIkWajRXCr87K
E26cqxeh/aHhlcuB9pFvVEGQS0GqmHkXgtWQpp+sALwJAuDlmd42KDqET144
28fA8/+Ozh/bO+bzNQVh+ybYqMN9okH8JYyq/vB/JXkPXB/uQT4OEIP4TNzb
4pKo+Wd0StzCnvhH/MvquNlFTzI2FYY/MZmoXlJGQuE3T3pnJHG+ixKv2jEY
Q9vi29feS8p+D0NgbjbhPNj+3GiO1IAQK71jAxhDiu6QaJRIcg54/gzWw4Vk
SqlINhW8AnIe5uIMcRE8MWPfNnUjSWb+Fk3Ed5iTkgDthWoREvrq3Cqa9k+t
o7Sj1T+pTnxW7u83sY8ioHfWxktsObEoCfLaWbgQPqhIa0iypN+gAYC8xQ5Y
/EFvbpTr1ShaTQPznq+TGHXqT5P5uVY/PET1ebWiiXo7d8Zi1I5441Ohb3Fh
zH5tVm/msaHS+OgDRLxdYybtmowBEpkcrjpqCOjU/V4br/RVJp91mzenK979
UdkTQFxIm/j29icNYKVvJqNrIJYoaIj3SrA2WPWRxG6TBlBIaCIUFNV3vwya
Ya4mZwMYaUqTbOtEKpZqokYHYVo6sGJ/93WLtwJBpp1umoMROwZOyidqZTTN
lWQeL4waW5YPWbptMn3s6Q+dOqPcCkaKeDgsCMXUQTMYIMNdpt8tXMIDCchQ
C7qRsjkOKJyHpxMb6w7oce9giysNXngUwtzkJln80Tptoq9U5W8DWkMfifkq
Pp1pFuXu/4+GXSMXpVIze+xU/d3yHva1hY6NEL1VGioujJLG1vwTbUoU7LKL
xtnFFkXyFpl/Fj/19mJvoULdvweisPUxaLKH/WdVTeB5kBWHMBMkacVwLXec
2mDOrTNvgZqTWh1Y+u6TQ02xt5EeovWi3vvge9WkRUpYXEmdt7Zp9mQX4j7x
Tfpp0yoT9PSo//FvFCSJoEQ2gbXAPf6T56VcxaWI7JpvfXimHyginDZxPS9a
qhlQwVfZOH6BcoIg7iND3Vsrn3KWoD30xNco9ysdLECr8TOxi8eE5aYSW1qn
FchYy7Bq7An6+uPnCEFN4dJAGaAPCwkELnzoOPf7HCqZv3cSDgRj9pJtuyXd
puTO+TG/jNGoHxwvsXrveRA7nKmQUMH4Ddst0dyizDV0HwOld608lN7VhvUU
2Z6/eMNerXJ+JXd5bgl88w1V+EzAV0L7Eb63aK3UzWBABvCcfKBleIaVVyXk
t8d2XjScUKfrvH2hNnEvDl1fC5u9ymcDaBotKuJK8964Iqbb2JRQBOPTu//W
euh5F5JHp598qaBEWfX++i/dDFNcA0f+6c4qbuikof+lS08A5VdNNTNH6Eht
lJz8mmkxXX6fx5VFbZzycuw8OVIlMAXZ3jroLqW1kWaj2Gn55UVvOMgrnyY5
RL4o3iMfzJl2XONsjPlP3fE8O8LcG/amh1XS0DS09BkyrW8My7D2CQ7lMkkj
ZDhI8UyUtNnFQ1ZIK3Z7N95R/bTVp9YoTHNhD4stLjNp4cKbaLgtphBMkbBX
jXC1IhLKPhyA6wzwUFQSiVOxmXQ/NWCeemaXYEm9iyQCoIvrhTBW13Ud4l4j
9HGA1Jy6qoGpnHe+dp3+5dHkCSsw/MXr3aeJaZvsbjte2MZv45R8NGuqedKW
yKrMwCDslKVD/xjuzLiddBBO4qA+NRtfZJl5iDauEeNTYt5nc7uEtnHdDuEn
L7n7OoLYYsDklYzSUoUP8qMYw1N7EN5uWQ/sYfxs6XM/RCyhsqbvREQDk6oJ
il+AArVKg58I+eq8h+Sf0pTxqY3XfILdac6L2bW+OrKJ/bKnDYRgtdUqZsdA
UYPrM4QIZceJ+0WQyCdgGlUF/fry9xPqldr5hYBazwodB7DUtqshmr0PHmXJ
DtiLVB4r5ag2vYgbGw+C436TeIBH77XtXPhiZwTcAiWrxPTgrH4nK/aEtIuY
bhS+ZIdzZjoK9stmtGfjBM0O6ojn0342mCoJqFvkTYL6LStZZ7m8UCiOG6aa
aJqOdchFCdNZ5FFIFNyQFzitRwJyPiAhNOxFFABxxAn2Vcr7UfRYHICG8CqU
J1Ob1Wei+6PrL2VYVPS6BBK39ao5Ojd05AhiFFWaKw09+URyEy4bBlFuwTs0
TzJ5eHZQEZdkd0wOFz9tS3ZQqr5zpabMq7Ts8Ulzhk4d0dRgwYqRtLS/Lkpl
8ryfc+LOEyMpudk6IJ2TXQUjJpyDfoU9IY2qMGoLGymhJWcexR7Xf4cwI5DO
kFAbBuo64cIcZE5Xpv4Tw/3s2XekGULIVetyQE+Q9qnkSoYPZ2zFw1i5+7xK
yxBCNrrBk9p1g3A54riHOaQiyiL6BYN1VDJDL5GqXLJQkP4Q+r3SjsU43DXD
40APjvDdF2UP56WpEJZ6rYEs/eZyhqFgP9p7aeitsAMBJlLCckvumrghY3yf
6AYGeaIJLv0qusgUFztnNpnmHKvg0wPZPJrgwmTbQuaFVy3OHkxBwTHAeMGc
PDpU2i75CuElGQE4X98cOvk7AlFWRYZLVJlUzzyM0eFeJupnyB2oVcFW3fcv
WSHLRfiwQdOv6kZtHJYxEWLoCckf9x/qgJLuugcOjw1FgPomu6rtan22wdM6
UYlwIkR5DBc64/YdzJF0+GAaN2Yg7lmIhWFOe2hoBq3mwCrtjBX2CVTSmKlD
dyz7wd2Sf5yyPKLrEyNXCM+JZcbjbiRGT2w3PYQ4QEPXJVSm1lej2aYRVVVM
AOrYHMBwgoWcTmwv2RN6HWvehRxoAnvLOcuW2k9uZ7bmAaQBF/Fwd5gPvZsV
4ahlMB3oX0FyuERxLSVsl54ln/aa6P8zewwXit/5mkAzXLE8TyT7sGDxfrRo
enN3H7q8XwyPp7zUriUUTPurPlf2tVzoE9k5G0M41jlQrk7S7JONBrxW3lwt
mD1ikxxIpjWI0vjebSXkiZXaCQ5Ph1cYAc952/Sak+g=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1JX7aU/eKXwYecrUeevKQrleN+g94G8Zrh3nM5YpmxLdGHkB77YJmkJh3tQPoi0bab/439ubwcdNyh0pUpTu+J8JH1LHmHwnGNfGMKVRUQiA0CQNL0IR/BdWDxiYO22CiENifuDQBp2kpy3+OUE162uwmDwqVWqntDYziUXhYM2Ji5NYoV0e2EkgzPRZ7e3DoSvDQmPS0VEQIPtPk4SI/ZlPcLDvibBWZ0wjHwdc6gz2t+EIKqhQ5QQTkGjwX/p2ZEj2OwcVJFyTXMdwfUZ7gPjukgd2Wo3WtUn61SIKISgKezyvhi0kbiX7gbFTwhnx/FuRPEMeERu6KjAzdZJBr5F5wfN5JdjGLTqDdZ6cG4Y+HjP5COX2sOGAr+5AI4vf1BLrlwVNbxzCRq/EIh2X2hp+ORM71DnRGELutQsuxGi03JkPHSuHWvhlf00q7cD+DMBl83oLA7/XmPU2iSA7FymwCwPnPB7puVOVDebJbPFqH/dtoBANWwwfiUgArwom3wKaE5qaBgVKfsd+6QqtsPPpWSz+Aa8pqz1neyqz1bpiZsWyUvbUQF1pQBH5lUan3NTbYBYws1/DPBEQZiLrv97Lco/qggiCVpVg3y8wVKjhvQkXmhpU+/Bg1zgl7PL1LGgQp2lMAWw6X3vEa5vvn1UCCNnt9dxzymBVo2w9Yypxec3SIL+SpMDPijGQbao3SFPZ+RTLwTDIYG4F1DzJUoqItDPLzUt6KJ4fKYfaTz+ScNCuhZsKinNGmACIiKx3eAXL32M68COKnjtzSz8n0S4"
`endif