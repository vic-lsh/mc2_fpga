// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AX++WrAT/tTi0I2NoOYP4lCkT2bsp4yQhFytJkm05L9GkRl5I5DAKKPrxGir
pHcgpKuA9znaaLovabnoY/e/D6VuaOwx+NrSzmb6H/8unoldl0dFgEicsZpa
tvT9AEk2URC2XzV8mQS2Fb1T/o4VzbdV3fgoUkVsgsnU5evMLB4Md1kpkRMk
34DWbfwKBVChWb70Dm5Bb+BLTgoqx+jIiMR6hVtYf0rbvwc9qTvix+xGRk6U
WZyjCbOJwyGSut+wmsrfIWTnIp5CsM86Elz6cXfnPYxyk16FYPIVzkX238Ox
gLXvOXH+xAhu+STL5HkqEo8WFCBXHYsyxDd2TBSVvA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qHc+OdAu9unne/6xRer856pebhFejecMbrakv42MXEqElqVnHW7P4AyWMlYL
GnS6HO362oe7hx8zAP91IFAZ0bDXqi7Ek0rRcL24MYgzH5amQW5xI4CJ8yoB
Yqnevm/vDmlQxlJ9cXq6DIJwNDBus/ebI/o9ROcBzga06gfnASjFn4N7O5+U
8r5B5qisdzE4laXHyiY/5AVqc0ZykWMPUc2eNNwNgLeg41KWLFpHFBm0WC8T
1jLXQq0Wq201IKtgJn0iTgAIlqC0cL3GNW1ve+U+J5AmDyxohr5Bh9H3TIr7
Qn7FFWtxageR5m45mQf+kSft3GQTuDXAEL7AadVVhg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lPBUyf+QGuqsyIgnAmyk/AixA0lIGVt49siT79zsdkL+jLvA/CNFvj5puQeC
13FXvAtTMqZ6gDpoMMEG2z9TTa1zk/rvVAGyYNmv0E1iavtGJXB3Omjyx+3q
+7w77U/eWDkwRwzI93q4g+324OsAvdW2Q3qF0dF6RQgbpdOtHGtkmDB5KAaX
XBhLSIm2q4eHVXK4LvL10J2j+CMjMDNpmIrz0fHacOe6KVki3agyP4vrMMfi
NEKobf5PzaiXd5BVj80J3JtsCxMO/+mlEk8X8BWcq8qgfndigOhI0C8OqpvN
Ik7dcYpVBD390VdizndzsS+BhDhv5rzhRV+pe7tK9A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
G0LjMfUqkcYNdm8Np5Jvlc77WAurWtqwLFCyadDSAIxWUnVODy3BDZ/DYHTK
EuJMEd2N4mBEzinsuNTJBgbL66C9QBo528ZW50LTDWR3cUT9VQK0aQ1gYAHn
vb05Wp4GIFk7OfCAZLmWb4RjKGwcw7fUt4t3WF4+viYtxyfSPr85w8soSGIm
U13vgmr0Ur4eM4YDdeYl4DryoOSODhC6CK7Ptj7OJlAi44zKDJiWVTz41/BO
sLDyITTfe/hF5yPWRTABMLNTwOF/jABJC/6yNfAGInynNY3nazsPZb+DRyAw
Mtpp+Yjkj7kMN9SdxzhFKo33kpjCnfEw0aMTmkroQw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZKYDY82hmaMWT0KPtij8lyDB5rJMv33QUkB4Bky/T/NYZOgdOlMo5RJbwD4B
+xIdnA09W7smChrN33bOqWPlrsZxYWV6GDWXkuUuA0dOyNbbu/mkXAr/+8BY
zBuc4h3Dtv1KKNFIuMGEJdT6CkyBY7v045G3S9gg4qbLEfOHN4Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GYdOURwHOZPJJU+4tvkGk9iIfOvyaKK1I0fNy3uPEfAGwjCQ95zJX/OH8SM5
CmVZLB6stl2+x8IIK1tB532/+wl93ztMO1Cf/0kQSQHVNyK44wGBu7dutt4L
G27ukNNBfWyawe+Vop6TevIt2MjQEpuj0zEHOpWmPkbxQxcFJADDCxPihcAv
ShVdQZ8BwL0MAiXOmyx++zBCiRzpLoAqAdVgg+Jn8VKvAXjojhH3M4h7OjRS
3uOge4tKrUYcC9OSL21yjcjhHJFKHKfd2BW7StJcyWUZH/BGgdU/LahlNzg8
oPdS3WNU87rPdRFHGDCHWJ/xftpB4Nmoabxd3sBNo59ifi1wuyG+Ft969pGM
a5s8Z57j6EZ95JAgct78kCDk84H5EMU5oS1RyPR1esMnF6MAU+9CzG65loCr
U2XPvjRzhWy+B0pFLpPhcVtqKumbZTbvHUV4He+Bbp3I5KgfitF5ulQYhKGI
/MM/3cxMDKwTZPEaf7gq51dHm+S9CKdZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
u3ixzwdM2OQ3eQ1y4tl9w3hVI4PSrqU9PdbvVf2jWa+fv6K/oSccWrKO2kFO
/x8E7Uu5R/QRZHn0ExFRFEind4DmyuAMbZMjFwM76DSnqu/A682xuKVim4/G
kbuU2n2vcT3ShK8SlogPB3xXmaAHVGSbr1V6GJoEDkly90nEtIk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XnfbkqkF1URkwL/j54hHt9PQpE6T9VyqEVYwP7rc3+PI08WrQXbtlHw9pp7u
/p/4BVYjiX92cuWl26T/r/iVKDv1sfKUL8snSXFJc+6jxz/r/aJWC6n2qoAK
vyVk98RZSfb5Q+79YHowCQfzZ5iBc6IJKGBmOOLyFHykmZ6e1vU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 145776)
`pragma protect data_block
BWw0r1sIh5nWMlKkvWrd3FSTbCu9duGef9UVvQBiv9SzEgoHOJN2fIjwkPuG
4+5I2jUrP+uKvxkpEr66Q2a+Re4i1yCSpdZWWaA3HszzN14QkjEW+n/XpEYO
SCyif2v01i8Pvk28LxXGUOPEGWXS9WxYvgDRdv0FsLAmfoO7EcG42ZecERSw
E4EvXsWT8Myj3gFGxwYeKQMN1UBABCsSuQDdR0+FVwxfRDQUc/8paUryFc8/
fyurX9T4pb4kB0Fali96KSRrouo6ZKi/R5gz3se0UvwuVgIAa1ybVG86Vnkz
fTKFmay1S9nHT2KogHuk9x/I0XUGiV7fqyRksvbBwIUMxLnYyv9qnCeQwi4P
4glGYBW/1YnhOIi/hojp6bAHYYYdLtz1g0idYscR5INykZZBuoRU+xE/l7qZ
h/WulVfgBbpUOwNOxMtm6TJKMV0ua3kzvjS/lIvU/5gomK5iEfw9DnbY/YnY
yv6U/0UAFv/duDzAopDd1/N+31DqpXVbXfOt6mxW/c4u+j/XWd696yiPXN3u
AfipB1tsJJlHmNuu+fWRIdpo2aNNdfj7TPh8TpY0V7lbUMlcTnL59uDmScfE
LdtzEXR1dx05gt4qiEP8PlwlRJ7ea/8jeQ5dCLoqnMxmJCWMr7hSifeTatRJ
Dk6vfLy5drceSsGGlW2SwUMbE45YPdzM5H4604goS1yGlIiIR8HEQQrEZDdM
mlTTPWmKwK//cVcvPcM1RoEill5ofFU+8qM/WNZ9teW7kwOR6loCyERHaIuh
RMPHnT24MYMNHtre1WwOaldjiM1dsDMbAqZgUnlS/bCw0LVyAXuTMMEsA8MY
tg/J62zZvLYBbGFgaHGtOG69zxNGS32kkEW+ZN2nJ+LZHPrXeaxCc7XHn979
PJIL4EueW+lma+4+Z9uni1RDhNb0klFubqNjOu/qVFQTKSExr3m32ymlt/h0
Zdl+yFMXCvczr6SjpA4N3mm/EqJadR43pXn4oIY2Qqhzwo8mlpWoko6+INzf
N6FdXTM2p15Yrib4upVKYKkaOYXyHqVDTSWoKzBuBF1BiDkZFGLOfUlAY7Gh
7eossDfmqNBKeAEb2cUjhVTBNMjHV0vMIKayuOBHjfcSulF8b+buc2BG0F+0
2lct1jKFHjZF7Q9YdbcgISTgZaq065hyL3EqU6fxKWUluC9qE63dFJYabrfK
LUUpuHh0pxirXLdOJkoq6zl7BtUKqzkmUL54I2p39uKoSbypQLrxJZTf6V8i
vb0BQslt9tedrbwOEHyEN8s53q/JeV1+QwlAj9f+jNGTYsLfO03Ns0MccMqa
P6C2OavBLfkdpKV3safeMjst4WK+tvpQl3Z2BQK5fMLnYzYWGVXkubrzOmUp
slN/nt56/quMm7QD96YIWZpNUfy+jhQT3SNyxsAnK3xWSDa1EAevnyzFFyif
8EUCOh7X89ZwOFwNhcWQvONP8ErVZaZAAz0S+nkPl/Z6ODLU91pgNMzTrLRW
Gj9hHuT4Kc8vOn2bHib9D5LqN7aLaXbu8czSS9gzI1R0473JLIDYOiPH8v6Q
CG+f90OzvkJ16qQqax82OBM9UKRnAhSM14ont/7Plx5rQboreuuDEw3iM6lY
ge996vvggAQK99aJQsgBVi3LBGaONIgVeNl0/3P2jviLcSd8QJOMpaVjdSKB
exau9dpOOllKGf0q8D7p2tyvJFd3S1nbVVsICz13O5yJ7uYDj6Q03VD9q3LR
+uNiIgyOPGaxtt+ovjw3CXdCqItZEaFBNIeyy01VbwghsivThl7jm6KjFOn+
WNXkCGC4T1xbwu6/vDCByTftsdldhwQp9brsojlSIUolW6h06M/ty5A0DT1d
D0pNmX6qKciEsIe0e9osENFn20LUTnNHKwsW8fmejQCtlRcym1k+oPMl9aVf
U1c/HbWNvFupQReCO7vfmbM9tAKb/Qxkz/DMdIMAABFOk6WEcKk3hkOVizq9
C/CrSR7f9A+7oUz48/8jgjSAomQALahzTAXKXdjI/j4U3hYoq9XF+3Pu4GxM
adrBXmQSBtj6xKyOOqzyZxEPcqWP/jVQsxv7HswbGarOIbGkxbtB5v/vHtMy
D8UKVxeostH4ftEO1/ICEB5vvn0hZ7Mljka9bODSPKXzY+UD9ggqEnZ/Xd0t
dTlQcXwNdQdumvdz7uz/p9U54NDwDKyLLIxzqqvO4NkopUc7SVzxoWlE1+wE
0E2seEZiRzp2iWLzinkTdc80Pz5KjmaCi8Bfsjglfgl92L/ln6f7akEUZbLm
UyllF9cRcz/PssM8tZ/bTBKhhcwBrdET266STKIoeUoNAzJ8OXiVlAfkNPA9
Z3fxWbfWkpLNfmwpmH2pIKmOJGpipgItNIGLlB+USoFoDHk/jrWgn6ZQUZAR
wEeK1cDOSzMG4LnmJ/ttQk0QQqCv+vFoI1zIevKRJK96YL8l5w/6xeLeMG6V
J0/nNSIeqj6R9sVoHe4BYKO0akuRpdZywxUx8I1vWTltSuSdwZXeWtxeKl7W
gJHs/fjFCPow3+0YefaPbUeoh34ZDxd48pRNCxd/w+P6HVX6MyPyAn30sSZk
Ai4YiT2nfStOUQN+cOtT9DJQG8Ax4nibkVd4FzlaNR2oJUUuCN+F07Cdbeuc
ExHpnJ/gwDUXhChm1dl1scmm1dXXEdDFHFeVx720FH5aLlxU/tRYYGq6MP18
d/w0dkaKcQ2FEAD5VH8zoP6+HGA+FDHgaeBJwk0iRNOpoIqi9revrUPacZvK
jAaZtrVhxdsqSA5PpC+v3AXxt94trVWhEmyEj33Ji9DZLLx7HvagYOVghm5H
sJykD2eY4TZpvcgLKubh8GmIrUUDJ4rE95JFgyV8lIjXnyWzHfeHKuDgPXGa
XW3Pf/o+xYDa7soHTRFIUa73XJXi58VLHgPjEPpXkU1w8E+cPqoayF09q8aO
aYvCN2T4OGQCsAlZ5eq5B+BdLSU/2bWTKC/iPU81RxTWfs5R/DGOGXVCb0Pw
OcNV/KjhRglVNau1XTc+Qa1S9OWkG8+meiONzbT1IeLxpw3MW3IDz7H3DLo/
ElPP2/+C2FYWpkykT+IfXRhOVY/yBF3EEW+MJTDGFgn8aiPD3WNDQ1ENjE3U
JNH24D5E7I6a67udPjRVJ+OgTMfNYZLFsodtPMzed+piyE/HZKGjv4NZBbvr
cw3PXIB2Wdmfw423UtKu/06tV1G+yYlwBw5k7JzM/bzEw1EYtCcq4RfbghYp
edWdaSzEN8cwB2jjcFVN2srgmWV6O74nWpYrKlQvO6LkmyvXCl6SIHYKc/jL
RuYLOWVpHPG0NyRvLZeuM7evxpRF0PhG4wcKhj1hR+cudvQF+UwWah3WduHS
G49hKFJilHY6RSNVW4lwfrRGB90R6gq/H3E6UdIrOKUPs2LllL9HOdbObyZR
ZmKFWKy8qJ3Jc5DSbNlHb1wXUbTmoVLWE5Db8yAueppNBQqdfJUpz/opgwc5
fGyGNHvQ+UkwgbL7HuWWZ0DmLJYws53m52qWeYI0l6E54JKpEbPByd8KtgtW
/Xh9bUYHiKjFwvDPc99Qag0nWlUWKx8/slLm1ciIwBzb4KJHoKEzGXBcvb3w
slS6itxWFAuJn/8kLdEac5xMi9cCXHU0lhUrDybSbXq4IxoVkK38nidM7SHa
DLfWRamy1LMnxwkpPoX8djotpV54t9lHvgLFnPNGWG5xs5OaNi8dgIMAWsly
V1Y2b+OBuCi/DMfzfWfD8NCaIbY6VjoTcIKxat77WkzTvYUk1Lurw4/Kp0q0
dv4iBg1YZwpoo6GIEh9iO1aBS97fKqKlg4EJDTgucOFQH/RE1kpE2n9h7KWt
BhxeU2uutNoWQp9uw//ieu/jPVQhZ3UpHNipfPyB83gyhABawU1219xNCtRq
K6oosZJ1CUPDaB4JqKfJyGzBEghGQhotCazuYjiXxJueaSvxYxsGFps4FZrZ
YlBJ1cskXiJ+6iLGLdVH7ldQzQV1zgkQQJ89gdhAbjJJqkF0CDrrX/4DFVA/
8Tpd2syAE3HoaF9m0buJT5J2aV7aJB+Am+++VqltuME4lKwNKlzjAfsDHqEI
KozgV1sypfUnrx01Vx4zn5DTg/fWGFa35u6CVzTWfrSVpYvN4kBGmmGU3ULQ
nwB81p5pyzfXU7hApIoqSwUgJZqBsyIZR9g1Bjg8IOTEIfLGJKOFkFfaFwnk
cGMg75q2r1mB7xjFHo4F51MYOM7GLrlNtaJkIiOsrEArhVKqHbYE2bYlkvlQ
g3DdDI5G05ZRfmGCDfRySMAVge9bgB5+eqM3TUa17nHRWrFiOZfABHdiadGZ
bq5x3UPByZmRMDZYAWq0Gn/22YJsxq9szlFmw3gO651AeIUmQvz79JpWDtnZ
Js1Xq/lZWkaocu9R9q+2B7UDVdtvSjCHSgJWVhGybON7RQWXIcjB0bIf48Ib
8hsnTW8daaSCdOatCWO0O6cLbEa6ytOc0duuq6d1X7qKt9YxvPuLA68gCMX9
Dd76iZWFJT3KK7hvTdVhYFn0hRHESXJ8Jm2XobK1/iRzl5DEZlr56/7RNFzi
LUMVij6c7Q1zfZwWlO0Y2qHcB34vAeoyYuHEIXpdXaKUyGER6oFb5/7VQN3y
Jn9DhdRfv8o1I++HoQyqdMV9mxRQ1cz+Io3mbCiNVoGO6qr9QZfURGEtBngM
YbPCYWX3oI/R/jPXvWAa8YD/h3GmFKdvqdiwdWRxqOCC1mMc9dIs1aDE7uN/
wjnUZh4nhTY6QYpaB63ExY0YQHctZWxtKgZf+MkiNpgacdGx/Oo3OLG2dVU4
YvMbaBx75UQjJDo/ys4sDNAK81HyrjB30ySCCor9Rl1d8YYx8WT1d1+Fl+7T
wXs3jgXNbNA6Y79MrH+pJcJJmrBrlJngoTYc3ymWdOZ4Bll3EAPAfUMvE6iH
U88MG7mBDS4Rnc4EPq+f2CLEWcieK0GY05gBCw7jx5dQ8AHKIElveFr8CWOt
agQ60R0D9tqGCpYSUqtUqExEr4/rhLCRqmQE2VwxgBC7DIrPDmg7fdcFJq2J
fpAuD9dY560JDI/wdB10mWywSGMEfxOsYOc5ugTAYhD/S7ijjYOejvViOrKK
Ah8sTdfj5f1f8WrF5i3UmaRNGQWg86vZuISaR5BLyfHQAqOEVPe8LihUSxKb
4k5he4SwqlKN45iNTLfTiOC4vuYLYEbGyTKSWNS/il8qkfexBVy/9j8Ad2sb
SnyfqJl6bIHFeT7Zjgk4W1+UUFmRhk2Ad2EEb8o+le3fYqNLkkwCbwxNTORb
MUwyt+ewf7MESzOiUepAY7aUOkx3hjaJZ20kHDEWjj9b/HDfD/WrcIJKHo6T
SRWNXw1o7SLtvY3mFriCtr0XSP2vvpaQ/mfwiFNB68jL04r0Zigv1kM3KyfE
X813zA4SLUy1LbpPkDM3ulOUt1oXMuvZe4EhyOxScoz0cuP8yhD+Qp5s3kzy
3Pu8lbsnzP7wIKd8VdW9B6AfpxaptiNlR9euTPa+xw8F+SMHWr0kQi8I20U8
K2jBWqaYFz73cLAjuPD2nFfb4q9tZeZ6k4NGAxxyiMXp/qLk4fCP38HMJyOG
2z+NJWDnaa4Y5v/5iV4G21ACfCm0uAHZbbkzqkM6P2ppEKTGYlEhZz3cJjNi
LZb4GS/PNd/yda8zQ84cxi8asCM9NQ7y3INmBoiw3IsjxNk9fjZzMBIyvcJZ
zl0O0ICbS2qjJNyA3iwbb0QGYoNRWtTX5rtZONTvSK2E+AOdCYAwnkIykIlX
Mnrda+kam31v3D93Xet2vkqSuD1YzRPyCCfiys45p3Q3bMhwHPs0qtTWdEhZ
yuVVVC0AvJYSCYD3J9caaIwR6e4eCTWXYkMuCuc921LknWVjXZPBjJnl39/f
uRzUOmPOmsX02eKgXTiPLgTsrCnsYS2TM4lbaz5C0S43msLw9T+Z1PtlyiI+
NWVEPOFlM2zjHy78MndiKG2GRm3ftg60nVYwGaR3TdH4s/Fraq4t2H/byqzE
bSGDkVOqqe7Pi3kG5ACOdvxogiEf3SbYEwBsIWBvoENcN9nj/cijk7iIfYi2
7Ht53zQJtWwojyPhH4bv1AbR+M82U8qDVgxNaypxtahtZ+8tO56UXDRcHmXj
FGazVRYEtYUA+Un2/qXV70Cp9KJ/g3zS8R//EDQ6CotDuDSAbkd35YKldJL0
MLiM/ASuMUE7Er1EiI5qeO4qUs0fnqTA29jb3EccYuZ12SNhr0SrDJBnv35a
KenFWU+l2pchhIk5qkSSDw/PQ6gkWH1PYBYwJoYH1juhaPviF6irNMvqbPCh
yIpRhWOo5espbpuY1tfWcWPXzQGaUqwA9i6z+fW2HnYX7ppTzrRPucqy1MeB
VXZt21U4rrj4BPLYAKxduMQB+SquOEJ2+JMMalEBtAhrw8GmT6YCiO38I1W/
lR7anbOwfv3HB/O2GQviYKXW93SGSJT0v0H9EOqT0GIOcp8Gicw/Gou2oWAV
MXDpUouL/Poi9CyosIhUoacwAdwz7c+qlDeet5YqbrHnMdfdMPeKul6Q0Hoc
iJ11ZQGSyibyUjzZpmWeTZkTFGkjo47bU5n12Yzkvm3FLxFIyr8U430zxqns
gGC9iJj8a0Zn9XoV9juT+Uvrh9GAShVmSVknvStui0boPbLelbQp4AFlPums
ooQdeDZXbrGvM+8EYLXvFVQDyON5MCqlcbpE+eUStpz7Vb9Eeek2iaRSBdkc
saeIqahLdN6J4GD9zjbL/BmKpMqezJGTl8fxFHDwsZai/PevoawJmPXZMHIg
EJWzFzY0saYRFBuK0g96kxPUnlJVs+a5pailiT5vmLko6Q+3vSqBcuzt4t6h
c+MF5gi+xlLMfC65EQ9OFltAXw36OI0XaFmqfFbPL9WRjjPWltkHlGCvMbiY
P7GCnwPG++B2qvut1TJNy1S32ssskyCvaVS/9DDowt/EXOHDLXavIVHNZf9N
BLKGkf+kcPw33YGq2HWcBMsiIMREaOmBe+W8Wd0aEU0XlGhpuZCFy4/2kPGY
xuaHvtQXPs4oHSjB30clmvj0c6OKtS5UQfFOLwVslIIRPdxClsCYo4SG5ge9
N1Hb3ugDvKys3wj24W71eG0TBQTZo7QaShh6aYCmat1V0ZWQy8Z9ThhEmHXi
9n7rJxqpmdwxSOxKkA7b8bKEvet3TM2zYd2ZZwgMVB7kHhsboNtCUp/OQpbX
K15cpR38nI07v2Rz0Dahd7jxulIzmVs+0WzQP8dNP2u32bdI1pNpc9dr83At
35hFjedpaioTHSzbQ27YyA2VasSns+SwvE56VAG0A2qt2vQK62FpWdLP5+oE
pa2tEb++7Dn92aS40pJ6YhyM+y7/BDesiCyDS8NyzqJHq1Pz+66W0MGd4cyl
xw44MJqNyeQ+flDrRvvhv9/XAg7PmtW3Nx3evob4ugvTbVZu0Y/pBhgcRc92
05CPKZwl75SbtzFKW7BwY5lLjVzsBRn7O/nSo7O3gXNTkxvgvXrWKg9SNT3e
hXcavX+c4CkOKIzB5JeA56sXCwRdHfBif3YOwg6DupjvnpCu7sOllNV+CmSN
mN5brmu9kqZ/SuedMHKqLGa1g97e+3xgvJcWKCDrU3CILQd9jZIVqasFqIgU
twsV73huN20YoHOsMFG9U3/5au9m4rsrPD6CA3UWh5MT/Gq9q2oZu1VpZyI3
VQAsKyZkGFltWsmSAoqFpZoqu9IJkyQ+lQCH1icERkYaUmq6bkZUnIRbs7NR
QMOp5gbosKYPuagovzdTJR1+HlobHamG92gEkqKQTaC9Hw2gMJ41gKZbBu8h
1b7VDCzU1tMgk1UJdAegdcs5UQzs6tfCOGGsZKYleOvpaMOzB4PU2cUHIeix
+JoXE0EhtY7duEpA7aGPAp3qQOaTDk0gxiR0r7DHp7l95oDN1mQS4BoTs28J
zZbF779ZxQAQeGTO8whMiBR9+oUNZC8MvePl25/tOLhF+HAWFP2T8P30UlkO
PKH7IqMvku/c5+/lYPseXWiiQRi3gt/vVsrdVf3sL34ZuzwzGx0Lg7lo6M+g
dRr/4Bo/sGfuA5BnIBxn0USepx9GsEp74+8EWCO6DnKLpzo12/IoD5xKnRRw
qMUmSJTgXqwXSyE/cEy2oXx7SH17buSLOR9FrQiPBhp99asyV2OVNZQMdfjj
xY8de/9TBzTzEeX64U+lBceoNgyu19nDljXaFpsynLK/URaMmmLUcCsH1meW
xf0aE+MmXBPbponlQZHanRxR0WjGrU2XDCRkn2PWuyIhMYDBPP3JHbbcUxhj
Sd2MdMlXU3c/t/91NmX/cIoOTFYdYQzs74Fav6+204w0fh7yJcIbMJd20J8z
VTtC/KK9nn0udlO/+JUuWpRGgKAQdeQBY5IDfyU+sdQbzv7+aXuwdD4isaub
RQ6TLCcfikmfI+pgLjhWH2cKvZhC/wRk9fvyyoiLKc9/Tk3Wj/CQB7psS/Ea
csb0Zsjn+Eh46ilLLlaAJtRzl7a5nXLUxSDyeF8KM9LtKm/OvTy+UPtSMbxT
L12Oia9/mCWwDoMT3UQP7Z6T1Qh++72oAMcNNVzZX+q/6HJLOVoAMhySXPTI
EAQgyg572jWTFeoof0C0OvRFAl++JZrXQkv17eDFc0ukOk+KoharP3Px8Mrf
XW3WmCSxyPwfAeqf19Ijyhep6NkoL5L0R6mUCVxfpp85nzArCpqd3V8NF28i
kpVEEbg4dw7qFSUO/hZ341MZaQ38wTUgH5z4xSn/6QXXol8ybdU7aUdho3k8
bkO9hJBB+9eEYEXVK8pLZPCl3HF8PI/b5RriQJ+Yl2JCcqqX1VD11fIj0qf9
4pr6OoIRvkQ6y2uBRve2rhzZxA5K35Oc69otCFfoFyULM9BFGOG8rxvVB1rJ
Z/FRB/uYv7BxxCaFJh95ar1FIZJC54dcSnTtlVDSxA53ScbCrPD71AuvYfJI
2Z1wHYQ3dUPFu9asa03Wv8RS6p41QSZ8msrq3ieofIQXenye4xDpMzk0Shvb
ba7sPJwlIHtQtXYftHv3blFBGK6sN2GjI8wr6o+Cr6odUNAcjdlxrSmF33Fy
6CsllPHT9XLBb7icm9jf004mHyHF5wbpniHk/slXkeI/4a9q7ymL/iWE4Nh8
hN+B47EX8ysWQF3c2xBO/52y0Niqpu/ZQ05UyuaQTZCgyX1izFRu6m96KNXR
7cNNLBHXdmlNWWgheMfB4wC/whgbSeihe8oW9LuAy0pbMSGEm4azdGJWCSTd
j6NmogLS/+6y4W1C9QFPni76z47NZKyujTa/bsEumNE32/mwX8Pm5Szb70cX
toAHYvk2c36+K7NG5G/puZNc0m15w7Prkai5pftdHn2G1D0/bdUKqE+EIniw
h5G6J3ChpCcoISCuENWe1JWN2RdfAvsVhizRfK25jwWS9ywazkqZWbfM6qvU
WMzTL5sVJiTJLsxJy8VawlAb64GZsfpBF/1MeNsd56MbWHnumQML7+EozE+a
W0xEThLIhWoSK+FgsWMDwUXXuXKPYLqYCmLwcxYmnZ0OJgR7pyaRwcyoBj4I
nYLHtInVMnBUexGBeX8BsiM2KAD/KC9Ft09eMBTzqf/QhxZh40duwDzjSp2E
aAie3POIDWfSfHJzXby5szCzR+LU6CeQ8tYNntfNgB9r7W60oy9SF4wQG8lw
E8EHNMCljLgnWbwDiKUhfkjuUTI7xGUkT/nbvNhU7qL3EaFkkoEc/p3dxlL4
MwLBqAOCP+dqozVzwoWJ+4fEK7Vc59dy+viVP3Iqs0LljNglwkPuPLS5oF/X
Mc5OenDCUjpWwbMKZ/xiKtuFB+Pnm6taIyeDVKToCfOBRafXYsfzIzL+IfSy
I0te/iEuPZQ9Kv/MKajxUboZlGCINryeY4A//3IpIzF3GMrttJnptDYUt39O
MxzQG90Zb2O6nVEvWaZLW3DcdOqSLOv5kNlRU9E0AqqYVNAkX9n1bLcayQur
k9dUtJZ88EpTwh6FhfkdCT3fwfnlqnbhDcT7E6QaMtdy/vFpJ0h6rJVPv6Ja
UO43vbjVJW+kHykOVE6mgj+aVgHqrs4lQmcf2ldJO4pyp0ZmsxK1VD99AdDn
nhyVposk3agtcri0rX0HVA6IX3aF6yhkMOw8B32za2n3NWqx4kVRyEumqrc7
C57eGwOaIEYlWos32rO2dF9iJ1U03a2pQC4xkJtF353ZAHVFyuVI86QXuMhD
HB1sR15SGSbNwBFTb4rD4QUEVNHVKVl+9ihezxpUN6XQYmBoHsEBlj1grxvE
F+bo0kOkXDEWqGcsizCEw2P4Mzu4Sj0w5mkp6EWUa8ccbbR9lfeZN+b7TtKO
J35Il1c38wiV9fYoMAwe1xUDHZRJ4bSn/cZpKXqCRV6UDuIUGePze6Td+Tdj
qvB9TJDBRAlt55rmA18MLlz+AosxM3c5BkUKXhUXgpRTLH7U5zI+eHNBKbVi
1W3SyyPKpkhySUAQgOzTlsOG9u4v82JT2Od/X8Y++GbUmrpaY5jMUDIkVp4a
Hyac3qBsJjvCeWu1ZOtY3s4XfNss9FRiHnByFqrL0VeMHEqQ2nJthjh+0WER
fVoW9Z3DO2O+i/0jq6A9huqKMptGZNfX2J7YV1qWqI3ltK2IVDJOy7S0l7M/
Yqmf/7zbWNhaP3/QSIct8qXvpc2I+O4PXBq2Ywut5NbrkkJtj2nAgrytEz0P
e9bbr0TsWkk7Vl7med9dPHWxj5IGffMvMBpo1aQzNqPaJr200eTinfbUgp/E
F2nLfe8qcaGKxNoxDoL0Ad1wG/309BOgmYGarVYLzYRN8HRcBDdUupEHe2zQ
C2/LdppMjdu63vIp7+tyu7+wSyQ9CPvk7XmJNFh4/qOHkUFPOGlpmvFDh0SM
RQ0bfPFtWzBmiWaQXJdxkp4itX7UR1EyfEjnsKrAdesFwP79n82TRaTNdce+
r/APQMhWIS3cu6OX//nlELfbx4gKY9cAJSiM2YI75c96zNfH/XuGoNO/vaDa
qZtwiqDudKRbyLglTC8h+Utq5YICjJxAzXYMte97Aj8RFxB+czvrYesNht70
qyJ3ULfxN0IF8QTgvX2gEoFDZbTPF8boA6s8P6og6UDNiz2ZZkRe+YM8iW5N
xIZ6LPAhcadp/kb/TdW8Rw+GB/a/y/3dFCyAy5s2AJqxJfPKd+1bj0zF5evW
8t6uNrCBA2tfsWpT+LY/s0JX82ux92fNOa41phJQs4unTzTD75SmdAm73ODx
LRejWrtAryK0qSFi5mTShB78o3ombpAeJNAyG43mp0AYgTkN8JQ3hGHTL+49
j5XD/sDnF4LCJ2QFyJtdshECgdALkw8UgMPxVg2nP7IgU0KDyObnMRyG2Vo1
85IMOajWGBD9zEHLqBF/qDe8JQaXMWGIfHt0V3ALGeuGip8xY5cpr6oao0Da
s31e9k8GBc4NC3InRH6w2Cg6RAOhJpdbbmHo1SbDo79aSgeRe+zxxAHwse4+
TRPib2LDr+o7utZOvWLbjMw/qCzkDDUR65e1/7U1lT8PF2tNq6uWVMLS//Gk
Nvm2jU3lr4t2G7KoUqGfzg2ibMAUXaPvocq6JSaoZLpIZa3LtwoQhWRRhiY9
vVrFfylFHUTSVFWTyA4eaJpvWw7/sf5aUobFCKIfUVGRvXZVH/BYzMeDLBEj
0EzgUWDsTlXHFOCrJKx0Modh5zrmbjg8aa5fre+Kjwx6PCcVSmPBPVmKgDuB
rNFuR5JJs/bLYAL3FUl1CHITw0u+N8IaQ2jgA0d9ixzh27pxScleMgfqlbbP
+eCOR7RvpAVtPOvbA63WjAEB09DeiluAZQeAGywb5nR0Dptx3wntdqvzzUSe
AzJ59T1b4bboM5Z15EudK0n5vkxqNp9GGS4dTogJ/oeRk61a/5ZsDZq5lDMN
rleAQ75Ec0j4vAZtO4OrlXe1zkqceVCd4zyuXcKtmYNInAw501zIC9oYYsPQ
z1Tv5vm9xFc/2dAXhR205rf+Zq8jC3C7iSFp1qGFD/s5dPueRz89wHPX4PiJ
uVCEglok1fNajm+sysFbwxHVfEx4x43aG8SCDpIUyWSyivc05Yo/xDKTtev6
m5QMIFK0NpADcpugJEHsUTKzlMkepwreOGC6DPeOiJvUUVY6mUtwjF0VSzTh
rpAduHq3q/uS2r2oMTJi0ureuVZbQhLHumCsvcf2RpRrxY5emW2UXvDxTi+C
ZaCAkhE6B78wyK1Lwe0Pp1mY5mg6+tEvR2p2MROMxbWangERSeXDlnQIA1qi
ikVT/DSmwXukoldTcqyO6GLXe7qWrcyii8Kb5MCTc8wNYVPIb7UauH6D4xcR
X7M1MJq5OjwOrSC0ozZ9lQexlvQ3y5bbN+BridUgoX6H8Bvo9uyhR9cmo9pq
PunIQ8v/ZgfoXITUzsR4OK46Ir6X0ZOK/41+dnYmcRNSx2xGhUWZnOZURF07
tbnIYct1YyO6SQoYsn5zySVg9KgetDV8SFjDBv80QxQOsTTShAn3BHJlbIxS
tzD2P8vM816ZJxTChGmFE9oFbdaxaVk5VVDaI5mxatm7OPH3Qz0hN9Omwsa/
JLj7A7JlVdYZz2eVhcQt2vPjEfxmZnYYY7Vt+MK+srZar+Rqf43Q3x1RxbEh
or07VDIrB7CakRs7cS14B+yD21+1dmP2CCsY+RYLgCwliglMLz/hHwHmaHxm
xypNgMNWwh8xwoTmENywYJNNACWgQOPDHMnJJUW2l98qB3jbMYpoG718MQ8A
59CN5vtBN9KWqGqe9pBWQDI09AgRT1m1ODNtoFYDy/yMOWa+C7f5ZCVF4Ogo
zGp6uzJx+HuX/d4vdWLBXB7ktZMvGIOALjOYVnaDLO02rUZawAJT7u5Q9lSG
KyZOeFXyBe2Da6eJ2jnyKafI8NcG7+hLo/C70UggNQRmu4v2lChbaUsMril7
q08KlE9bSmeQZs7YwgRlJl5Px/VChDxefNjb5aBM5ot/yL6R9JknDYrKzVKo
5kTa+RgBgOAXmlPPAiHtcL5g8+tA1IAyYozGdEdb4Rr3KCuD816Sz385X3IM
BRaL0QYy/R9VBZVFLmw8SOU8ZiTS1eLS3UmXUjdx+OvPE8Dts71Dm8qXzTQx
+5PsN4LrrCxs+wEJERt4TSCZ0rgTC01pKUa1smjbp9vJ4Orz2YAFYMyoz9tt
VO05lKmP6xDEgGBZOU7M80rscpPoHuTaVE1s2GN+vmLWsxTbhQ5F2Qjon4Ye
029R+0vF5qGeHCF9sBx75KUwGqs/9ABY5oIe8q/nrCh7ESmINGRJLLyynwf3
bYPXVNDyyI/BAV/70eOvp3SD5bN4cHgXkgSRG/cKqTFs4K/ekIDGA8W1IWqq
gzlAlxI0SL8wHdLtOaAV4UdRSQbRZN9H7r9xGFTp0ntAVcMGyRAFFzurcH28
LX9FoWy4XIsAJ9hP6BEFJaT+LV6B4J5lbUkdX/k7Cqvxq4GDyHV2S+1IPKXq
wKtwh9QNb8bHGJFT5Yhif+/rr9hUyN55Cdy6BuG89uuiKk551BtAebjafeOG
oUWtnEZx/j/oJARB7/3tLitx6WJI8HNQwdNblx6gpivSg7dBnK23hfpSpGMu
4mtqvYhbsMpEQvyLPhbxPiwg1uRQPlXxIEQk5PkAc94fBgGY3WLT5KqM9SIo
kLQSthMXQryUjwAMEzMobNcy2aKaxN+o0D6hBF4sR4V1b/8x/pufNxPCDjji
Ui9D8Y0YA+b8FJsYDTT1+z13GSbFk3+nIVz3Agy6DHZ6YGVZ+ArYkAXPTUGD
T/qjU9xBJjKwlqjKIWUKAtrrp2MYq2b80T25x3dUatg8QuJL1f7Bed1M4tq4
tjQ9lyq+7/DQNWsE2AmyLtK3cmyaJ3i0x1sH8o7PlQHSx2ava1UOPfXuuXVM
6KEzUWsRqTdapTX9UNv9+7iV8dgb0eHRr3jY7tWXxvY4/8QUtIAhW6qYz23P
31iFTq/42/F5Sjo3a86zTM/RfZwWx1MrtaJ17TdB7z5r5nYzv+Oy6MHSEzaq
UWijjrOa+9uoytAGHVixIdd73Ce3+9Dl8IfwgQWe2lzWhJ7pGAWlmmFMN60E
X4iGV734jIAsbLA5w75j6RH6j5i28xFUL1DsBVGa3uFlxcR2Yas6szP748nI
Cr4uwCXO2F/TlfPst26a2t93NHFKPH5yuRUw2U65ZtMrrOjxQj/Q+rediTYH
8gN/fmGW5ZF3eFP7Pk13thsIqEi/NNEiqd/wTBfjgNr3LSXvELDIAWHr7Gta
wcHjsoZ2/pIw/C5f8W6QyIFky5kveN+XNyvzOkSOhONSVUoNipKcRZlUz0ss
1DAVpsJDZXbcZ9vAsqicqZ4WsFthBkAMyd8Bl5IG07V0ISIoFsUflVr63NUX
PaXNW+MkvFatO/uI6GmttnOq22zloiCN4gOHe5YWmXHmyro+az0djfdzoKqV
5j4QlNMN8HbXTF5x1/vQI6yJfRvBLDGi/93ft5wDKQ3qWSt+I9uXlowkvAfG
2Kk5oZJGxlYchZdSUgIpzUhrL3kX4cpZOeyPZeGjW3eGPIhrMNJq0tX0hRB3
yoK5i4DdDP47juaQRg9KVWErUh2/OiDtAVMtq942zx8Yt2PUnBELbleWj5kA
45KmLqfeA+hJvdZT6bFlTDQ7hwjzAX+cbYyjavl6ov+l/LqwUeuwzeBNlodl
fIiFp1mq15nRZEw0X5p5Lrun4Zi2vGAkchh7vEkmXfUpzhf+57D4DroeGhLa
vhZopJdfMvBFAQCb6Kz2++aFmCJD95MRhP4U2ZTWnOMLzmGHvwJ7SE9WDrBb
X7srDNfhfvoz0JiWe4A6thMpEOfdIbed6WrP0VV9O4onKkTOcrLMD5sb/bIc
xB43QAv8MNubanFNwjMswaoiHVxoCAHF37RDB6QaF12KgHW8b9JqJQUVNbEG
EBbbKTRo6dy6GxmuNNk4akT6mQinrMmsfbIK8GaGi4ACmoMOyzPiaF5IsBtn
aQxNzWs6Zz34urjCAUxfhL7ybXUNHPo7YZImvg+pIit+DPUJQSJtxRXCqtN/
+khBLPl8FFpyZiIbj6o3zq4PTkCCcuUgPDgR6caPvCKkOIRUz0T7oiccabpH
BOPQhUzin+OWwwQuJf8TsEZ+MPHtYlQsRkq28SewRmKAym0+Di8WKSpD+6my
XFS7bsn3wvaC75CdI3B4bSCBW1R4Et9RgUkMnhu0vhGvMYPkUHG/11ONRknI
PxdlL6bvmwVmlirVI79ro626/R1VgrdJWWqfrK3WIyo/VnvRiB+byV/+NQDl
FMXwSwDiN16Sj0sDTZDPKKiS1R+4SZHZt4FwwvG+4KlP5C8i1BiEjdirKjb/
t4hpkUMuqrgiM9VdVQpbFhttbolbn7zhlV883jZtMxZ1OmJFm6a46i6CkIWT
amum9HT6Jy0oVElun7YP++eNVOJrz2dlsoeHjQIJmxRLfiAe5CtdH+PMsK4d
8y+OPg0EJK0ldS9fgPRs8/YNQGi/9kKrNgfHA4CZCzFI2sD6O3myJwPC094+
se6HGdp23pne9wuxAQEH29TqI5Ask/nrVYLXypEnXhwSJxgufC5faOf6XaJY
aAQngqeeU2rv1bW+odVbOzKCd4lxtN/ppAtzLenDj70hebDLrKRoZDEYwG7K
KctSfcecvrHYr+jLngM04CWKlhYSkcOxDIVXeHwkK1RalMnNZ6hfLaqIZ50V
JHQvAapdkTurir/ohdQFUDOIIme87tShIFHoKT4zgjoiMbV1SaV+yYMt3tDg
MGsKhCB+h/nirYE8MtKaoN72MNyXMGcgUMRq7KeijMhU+cHl+MQpyk0OiuQT
e5resm0q/A1OHHFZpXgFr18e+8jpJI04+RbbzyEFPUwCSLGZIzzvW8PEdV/C
4L0BvDJboRkBOE/plgcAOKYGGo3oCxUKk8CRu5W8eI+Ws/bUy3F6vzkv5x1R
LnQzG3olpH08gUKxgsOcLH4GVOsSFPtrS1PPKlu4blNprPBJcpBH+bHwU6f+
oX/kDMbUPa7a/3eyjWdcPYRiZyyo2RP98FbKpSaN36cLVbAXTGTdn43qU/es
ObRWu5kxuwHL1kZOWnFD5r95rJGF1K8rV37MTNfhS73YGgOnT9n1yLrVprEV
VpZNfrNhb3kFH/6gkQ+rndtpvThX59TBkP/KZ7fGiezIM7pXdda8U0AOuNSE
NJqo9c4SxX2bxpszOVa6GCczCsRQ7Z4H4o0mWmFriz81v1998+FtZDGdQxr0
61xEv5cP9dXG0QROfGHkFMuNDF8a0sn0o2ieXjqbCp8FD3q9E+Km4Ae3VJQ0
IQCHGzlvNky0mboL2PiPhbCeivz8nN6mLz00PweAOyb8VxV0WJvOBV6DFEwy
n1DGMw6vX5loLtC+z4wiZEPma5PxeobX7D/cjDIoq2jI7J6vfjmr2KBJkrvm
uUx2TnFd5z8ZmKhoaYQDQGX/zqpKi+3cL1Li8glguDXi7/0paW1aiRDBzyAI
KN+LYXv+cIApDn9QNZ8j7+ZiPV89FqsbzFoOUxn/ThFSSRFrqa0empHhKybJ
Vs1lXuCgHy6Sqdezc2vjNYrhs0Pm0xiof7IkB2lCijciOhYlKP5K3C81Nm/k
PRKgryr6Q1YUBgdlKL20Mb+ySDl4E96Srtw1fI/5oWz9mxD3CXh7tQy0daZw
6ulYDFpHLr7ftXX4lvZQsUkTyPvX/352KeDHLZNZymQo7c35PKcjCcivpfxj
fJy+kB+TB866YyO+fDiaeRVZ2H1Ku/slsFTJP+VFtEhX+5UyLy6HKJCOTZKm
9TOYNtdJIupfifN/AIcbIR+uL6nEkNffBqNVyNWxkLUyBsWzxWfL9csNmCFZ
AboI2a51k58en9YphI1lijGpp1XVIDnTJjO3hZ2gVzDv/cEcPq6T2JFAmuiU
tekTsxujRJNVlpsQlL/JnX71i2YzLujaKXsnOYwgkzqWfsH5gNbL486XPR5Y
6LBo6K7w6SSDfPVxKzmBwHNgGUEJ2MHJ/Gtt2Ov1KcOZdRQ4EcosDHRXK1/G
vl6xYrQ4a8RcCSu9Zw/ZxZrbMhNw7Lvc27gFPzrur/f9pLDJECjqZFkmynUz
ZCN3dsOgigiTKSeY++hoJi1MhtKV58sCW8VhmmpggoCWp9vXcZzezztpV0lW
uo5E/p4CXq6XPC/X4ScxxEEvciDdotH4gF4qGSl6ujXnwXr1h2dNLwm9JcX1
zpoQbdhGe45K30HWcm4xJ9L3izD+s9vU4wJyi3DGFY9cw7KN1RtcdGi3edmN
C8VjIVgWbCpQPTAEqKFaImzglLjPUIL3dafxnsTSw0ANAdwQyXQRzudtatNt
8KQanzWaWFtuaU4mY+k5fqYoy+0CL73mn/12Vn4uzUC6mmNAac03+9nkJGmM
4Eqqs+4muoqAJclBE3N3SnPLXu3UZs0oUAzZszZ6poNdZ4Cw0Lzm9N9sl18H
YFYWVdGZTp0QGeGgW31H8+JTrpEzLV7Lb13ddAsdvY3Z3imrY0PWgJWjPkLs
7L6E8wKrOap72GYTF+O2z2KhhGl51a2PqffAHKgFlyVZvYPNTVWBvxIWq9bG
LxZ1cGDpuHHS/64omtbUQgnzn7k//0Zyga8gnd13XfwOukc3H8S9L0s76hGL
MaIV20IpBzO/RDDfmof+vKJ2mXmAJYpEO0iUQqG/XgqhKwZGAFEHTq00SBvd
ueBJs2OBCJ0cjjRYylZrlEc+asyS15FziXgKphTdjar+6w3a9YYG46GzAIq8
qcMLIFc9znuXbNPCzQw/eaas3+tq7b2MksYlb8HlZ6cEKoLdYL4BsYTXkcYE
VjApcMwn0PjBZW+3vlWnc6bh7JaMURPeyKrUZhb8b9kcfiZRKu9q/BF59tHn
DMMIoweW776/lbgL3YuTbqwj8By4RkvrA9KFNQ/I0yNfnBsp1Q4ZqIVrPbqL
iubvga+4G9O78hFDqBShhgyhApTMj0Dq17zaDX+2C6zVBOsfcjnQ4VeehLuA
+PbuS4GvewdyOZrcin0EUxoF45SBWvrF+OzK8b2/QjuxE0sHzUTJk4oR3WoC
Jml4KZlM8x/iHgJj+QRvM5Nhb+jIA9BK5pJM25MCJuStByGzju1WftnRzqK6
KxEnBN0cbBgsyncxm5QLHPtQh9VwE8u1dofz/3qGgXxU7eJq0V7lcHeKZ+Jt
sa2CcrLl+wcpbT2XnbjVbZepimTYqZIho8tCTetLl/3Kwhi7Y22bI4AYDGUZ
sLBiAuuWKB3ZFQK6yKQ9xd/pq9FbSW+l5iU46jgJeNTni/tx8/NDzW1QuyTB
EXHXuZHaWa4A2tU63EthY0oCcSDuFWPOa7c13W1VeTikBuRPX1Bmk6RFewrc
e1dd5FLeeZR2e6UbB7awcJovUKI9ubAzb+iYUimI3opLXZtb2hNl23gy0oWU
yg8yQQqu+jymCOgQXuhhlbsRSkD2+/OW+jqAaB3g21Uyow+gGdMlS7xlYiBb
NYQBRoQXCeeqwQjsboyMgIhQSUZCmhGkH6eMmAZTj74yw5QQ/4EVabGCJCyr
1Ru9zZ58CgMXaxojzL97txaWorgsvq1frAyKZabDduuFV5Z8TKKqfY40HCtj
/nZ1ttN+3IHBQbmKDLWyukjieZY6ikic3NRRj9pqTKGg2zUJcqLIl6bY4YRH
ro7KPfVOm6iwxFdLlZD09OqI7qcqUfjPxxMPCNORXEfmetNEC4XoE20tKYbo
wlLMg82WoBPZoyO/ARwNnTA9dJoInlhiiRKDpAyMLEIkUUZsjTjSiKRobnLj
WzsFaOmwJ/dNfuiuaTljgZAtLav86GwEk/2MWpxir77/MkTPTUZW8DT/lQaQ
23u+aRRjqUZoxY6HiE8az+Dv+o6k7Qn1yYGpVgM5TVFg5CuZicA+yqbOwtpX
psWvVk8DnbyH0tpBqS2a98vgSOs/RGxbrjskyqpTUQkNRZHoXigqT204FKVc
6aoUHFmn2/2y3ZZNkVl+seoT3ZAB0RGq/sJ1EYACUQj2wXfm9u82nlhx3M45
xNpv36bDqSfDOIdQuHaEs4KwonKtoAFGHK/YoXhHfo3lOkKlpT0z4wiUIUbr
eP3P/FEacGGD9rI+hzpZFRKDBD/j9HNwkbNjA6vU1OYxf2SdxgVQjlh9aI/q
+BP/OGxJoUcqBp46zavMSp3uFW649zpGUXTiJUckwQl+E7/aAoALdm9jFs8O
r1m8LZnnUKcE8y3t5wB57aGR88AX7l/E5jHjvGpDcfFewxxBVK8qFg+jN6xj
k45yWFId1MaFUy3NUldSBTK0gyP6Pk6q/pz6vonDiSL3IXbgnhqUbZW24bA/
DKXxo1j5R11JGOnFJEGYKv2/Otvy11F7nLPrtlfi+ue61SA+GrDSwUAWWXT6
Z5HjabG8HjJTROjUrnHYN4j6KUgYpXVFejysDfwFU7rye0xGyJR1m6Xrswex
UVYxHx5o5SS1ELNJZMKJmXOY92PfPiQPm3DicY5T+ET14h5ucsNrgCwWNTjW
HDHDjAnMm5xVAxPo6TrgCh7+AxjnJOkHyd+ziUQNUgkqUvtPd7fZYvQk08gw
ZR/pamGHSVtTe32gGwjaBApA1amgch+Vc40f+FHJKJQXK3r1zJfLA8tuq9Vk
FtTBaU3/iCJHZ7Bg+E3O0k7rxiIj9nPlD7FktCCvJhEGy9obkpODAjYU9MT3
zpOJ0yvZx5OA3ZUm/9U86NfkA8Huw0aBQw/prFtLG6/u4mS4/g/laajqka1m
kmqFLzDBJV0Mqr6xkc7PCLVgNwcFeaYhOkW1XoUHq7fPneV1zsmeFuSM+nyR
7RVUdttuq570G7ufrKAPzedhEerj9Jn4M92EIhubnD+yxXA3Iv60nuk568cD
tljvinrrgC9uoyl0Gq/6lqa9/HhnAqo7v8Z3kbhMW/KQ1zv+9g7t74xcZUTr
EzZA/9US79kbRizfe9pr/ssEcaifzWCIAuodBofsnuERTaGbD8U+/eb3dgFJ
SGhDhEY61a0uP2Kjkjta5QJRLMEhMrUtlDV1KWwXzVl4SaKhJ1/x6lkianio
uUy02L/Nmf18M5FV/jAdQzWLnAtoRFjKbPcTbSJNbtyTjkE23CdMnyBHbHJh
ajwDsRoxtzSRwupPO4fwhJtxDmd5bYHhwLfmYwrabOvboMWptuWqcHQLrq1/
WvY7AQi3UIWJ6MkZdkk3p/ReT3bTF9CThgZFyWtbSv42dFPor3W1Gf7pPGTL
GBko3S6s6ngETihhvMikgNApg9vOEc5rUz04lUN8BUqWfdxYs1Lej4HxpfA3
G29dtdvs4UBt+4dVg1pD7TkQZi61x9edjXiOYsqzG8xYvz41Kc/6M1r00NyD
Zzhu2wHtmm2w2QurS9ptgSg93YRd9cyCA+NkD62glqU4b9ukIogGfxNXCeeq
vsroJ5hU5TiMW26pBWW0Jyded94in2zMOMzYuU/7I5tyd6tJpF29exc2Izi6
wFUS/kTi1DkoTXVQHdHgNRFYu9w/8BmVYm2mRZg5141LqxuM4ARKFLsiUKTQ
YcvK8/WH+ylC21CngAWXkhd5Utl587KW7zBNeZcjczk9KuJO6iZv/Ug2hJA2
2HytUE+zWDvNxn3c/9WcUAHMPe815GhMKs0+Fyf+WoYyUXH3+zqI5EZytCGL
YOVwOtU2lJfmrStQ3DwoE5BrF66Ya4x/cAPE9PiJhXodIsrlFuHYBlwo61/s
Sts97Hn13B2Z2fnfQj0NPUm/wGpTQJav8uo6QtrF8BV0nPxYBExPFvY2DeyS
ONoo8mREG0q4O9wUdx975doEkM4CfzI54BKXydRRXAQ2O1KPmatZRnnTRQu0
e0f/m1dfugPy1yMZo28kF277p78I8cv4mV2ZhlbmXLxf9+dB3l24z2iitwIW
zhbC8tzKJGQL3gUHCSE1ph9zCZZq9Lb8nupT0VgRcjKPv9tln20+9f/xPP8/
uvwCFAXsqH8752P6/+3vJscVLsLdPpI+7ae5yVJCw4PkaGulA6XLIHWx9eii
Rxryuxr4Kb5dSOg9nwLoGnAxe2FrwMkqNDOk8r3fLdKPS89xODz6HF4oL01c
SpQ/kzawJkBzZsStcQd0lv2l+br4xwUzoLj7tzvA90W5edjWxAkG21ATlSLC
tcksrXUwqr+pZ6J2tyY7r/gYdM2IU3SOGeZJjAbYLOzRU3QSVzJ9f2yh1JX9
LgJBvSKHIlurTjc3QDc/WgRwqYn4RldoN/DpUnkku0L4llfvC/a7Shr4M3jB
zmwoHNfjuhHkD9/fSl6B2CxaASS+PvkygR8IqGSrZrTaH/KknJoPRJuXRTfc
G94pzbkirYVTdZt+8lTdQsMWYvtVROAcYCsB0kqME/zy8vfw22MV+OyNKyPB
fiw4FZ0wGzlcdAFCCS/aQ4yJlzPnhKDPViE34YJa40Mrhxbee7Mrqvr9bs15
N4uJFJMG4/LBfv4WXujKlV4BHtqIt92X0XgkTLbk8XVTFdzCKJgYk9Hz6Wco
cwYnAwYZMvNCArReRBj/hwi/GRgRyn/jhARKxCTWg5vggUNbWGVpU93tW4m4
BKIi+heXedt+XDhPxyDpEcjeaVQOE1p5voPdiZeLdRE3keFbTKk2+mnlUL6R
Er0ccTjg0i3ZwK5FUMTrMohMfqgktrT8KrpWLai5CbMUjO2vf7jkM/XhbK7S
6buSVaOpClvrobSefCVkxlX8YlhD78tlfy0bD4ecpSEi4g9K9b+HpIHS7BRw
xRVB7xrUrCFc16H/YrQI/wSJ1StHKumTYcGW3h1Qod57tehINXVQCgBmQ1r3
FVLCENSkIhxaqZlGM2cETCQZGHRN+u5bcFfiy8lcvotMBbnQeLrW40uwdKP5
c8yHUzYmPorhUKXpDr10b58k3ZUZqDC1BJPnH2R6wY3uNSYVqObD9Cs6zXAc
HrG/HS6Kf44iHExj0S91CTI9JjshMuBiWmSDxupV7Fpfa2vnkAyv0eMItPjP
CwmKW05O5au7zcMa7bLHT9mDuCetFBrNgn+FAoTGkGQnrsjDGJL6UAhuMzXh
qYd9ENWH5S5qZdOZexa1/tmwIpA5vQPNEWiaE4cMehDeiLDq1fJ109lk+ttR
wDqACy0llUY2SXRnjsMqCOynWZxwX2AvFuEdLXhpwhKevMPmKAI5vOnByUwV
hE46tIRL1ki1MK+KmvZDDiyBrRLAsYazh5NWMKIxAR0C3rWqYMZsaW1axanE
6pnLlOP/w24L8/eDbX1g22NGl2yDKQ1dIL7Mt6Edl5O3A1of9uchC/Au0Qb4
uarfuWMGOccl4JX+c4qkloYCtxX3Ig8qqVCGWF2ZU2I4x3Z1TlfJduNtGGon
xjmPEGTfOLO/6YHcQkI6hzXoyiQGbjEoxMEYnZDuFa/2IJfkjqLnuvYTI5Rd
BAO/WiHMLsEJPlyr9BmDVMd169RzTzigu8koVBOLtRSrKyE6AGd2+Ko8zXaW
/FjlUtK5uixVGfWjUQrcVY1yKIMajwqln6WxzpFp2q1fabsHtwOfl8GHcFCa
zknLvpESu4787k0ZWldCi9W/a7mXMOJ2m0lYRk6QyFHjiR5NXZ7VeWlLRaBf
EpwTVByevunKbf4mx+E5ZEakZrBs/U+/eokMaIPVXDAmIT5GuNUgTI5WOJMV
UxelYhEI6+EUjkIV52W0IHuLZJJ7RPuiuMgZJp+GwNz8uJBPmTzbwwXKVk1f
uelGb1sH0HmVg4xUFgU4wltEkokwWMIZ9WaRc1dW7/MIjcZZ/BBDd8gHrbha
5TRaOTkLhJ10/IfCmPb0dWdUbdzCLIFkT83BEhkfK1XHmlxiYhqFcN0zPOaG
GL+irP+6OTgUKI7us3P6UGXe20xL8x6QBNIqtluCmkMYYJ3u835BN0Xrl6OS
uWDe5+jTKNFiluzYybW+06jVebJPszOND66tIEnOlEZlHAsXvsgBXlr1FaGY
5VDqbv0DgqhhrMjvOvcUnpliRb8Vx520HfsP+OrSB6+WU35B/FDYmLGK1zz6
F+ZFNzArStnFk+3wGBmCjcgaSxguHbm1zqEGVF1pV2Xq/pbl6G0qkRg/mBLz
0JLOg6fSJq2tW3S80PD4KFKx8s/Sbu+Dea0/cjYtpQVvxjeeA42HGoDJepSD
ZR/CIvOPmmGMrKopmug3bzCskKz7gKth6oc3RyjNfEjc8kFAkpQaVcTgUaJO
QKdRGJh3J41jAvOQnlY6s/X1kiKsqT6Doy8udGi8akyprAyZ+2t3rbDWEEym
Zlr9YEPZ+mgJwvPwx0C1SRwwsYOxBxspY5jSbHXiYVeDZuP3sGYMciBrzEdB
CMEHxGO4mw9960zwjdJgZ7MxZ4dLgV3g7GXByc/e1d6On3Fg+t8qodNEZptm
MSK+1p94NFT7nzpVxALbIn5ddn5Pq3akYqNB92GEIwEStWmMT6QnWMZAC9ZO
XnH8Uzt/kpB9sgl4ii+g1ISq+sTd4oYJZVNtLAG7hNeY2Tf8g2u+vE/F2OSc
+QuYlRi9u44c7cOsFRyYx2clrIIAECQXfMYMUn1IUe3BKfj6Ja5HNKqaq9NI
jajwJ6m+PH7ec+ZxYuYFeb48jQuf0gudYM5FbkAz9qHIpPRHntZk2oHgnFJX
olhZr10m5aUgRDU/Ar2BTUokq0yMUtU1cSw2WAzu4iu6zC9mfBQY4gmxda1m
kh3oO5GkVqF/HF2uRn5RS0x3nEc6rRU+WR5R470MoOUlkgcf8RnLKG6lTsk8
QY+rAGwQhNUlfMu0Qz1+a+WHg0KBBkJEGvKWcVoRQnam4Z6A/VjGoGU+LtF4
iFadb0z0QszleLgRDIOymaI6x7wnurQvHrApmPG0/8VtdC/Bkm3zyq1CupdK
uUYxeikctvbklBcNHkJ7baXy9pAa7PUkYjPEcTHniqApsRzejhPar+MZYehq
v5lzbZSog2GQZUhL2iBFgdY1owVF3QTzWswyk0d6fcfYYh3vbvVZQl7DbPlX
BOBqYSvmBfuAFCRV6duqDFyJASU81dWvBE0mvNiXYA+RSQGILXK4Iyc1r18M
isRv9Q9DaNKRNXzu3rZgwo1sbcpKHFJZfLlxOPKBFdP0coVdNA64OHMtRAMi
ir9lbSblyZeGfL748sz/FUzzgWZxUl87bI7kZDoZyrHuN1YzNB5gEt+vnNUE
uEcxBbBkHuB0ltcyERdKWQ5N/XWkQH4M2NBFo5x1sQCY5UEWU1xWwA7FHZ+k
pGWBsZ2SOqtnzhvYDpCJeLSqV2rGqRKF9ux+UGluiRpc/NSTVrM9aLEv9q4i
h8u6SdpwxIVvR6/rjzAE+nmomCEOjWe8ADTys2u8lvanjnGs/YPovFhpYX3q
9GxPFXCnGZ8woz+SKL6aDOx2eB4kYxsN88v/2J5PZ+w5g6htj81k570N8di0
Cpk9OscZL/9xvtoqwcrZsT/xvWah6HZNMt/csbRk4i0J2+hGpHD0qnz8Yr9D
/z28qziKKomzf/n0rn5sZ7XplkqgTY4ApHXlrq5FKAZ3J5cuSTc3qEZ2or/Y
cjmBM0Is8qV697wL6JeGSYV1yAZkhe4lh7l6XwcSgw0h0nm9wboY8WbRnrtA
OX8ijGVEYcaFbw2M28H3BR7RkZStYy8WezJe9xVkz1xAOlMdluBbGVQ5DOSK
MO89ANRaOAp7rOW1RVWJiVod0+9eGdVbSDzGdvEC6n++T6oJjS4scws2l6UZ
e3VEwBuqXTJRfY+LC3lpzg/jOHvyuPNCq4xVTEJXmRImhSpbHhdi5ZOK1nxF
wJUaMoneVZYl0x1y9R58cvnX1BFLVDEYJR67SxdKx2m+JVCtcIYVGJN9sZKc
w+sIMn98sRwE3Fol+S1jZGUMCeEO/vinr1H4ZPpwT4DssQox7kBZogZTU4JW
rLf23JcdoobGROC3qmeboIzr8/9C+Mxcppd7O3wBLHGh+tU+4MzT/1KCyOES
U/vYVTbNj3JzBNjz+MYL7GC/LVSd/BEvu2lzdgMUxPMj17GVs32w6U5fOM4x
6LYNMquMKM6jWaioJi8On1dkyP/vESu5POrtM2hgm88RFxFxCpJ2yK6piQ+N
oaSJcYmCApqJnr0TaZHxdjanu0v65Gj/h4i8DQaYUT6Gz8xbWPMgzuItCxay
q0DBotOrEnUizOnLCabsbdawUB+FJVyawKqCm/5MVeQinM/FsjKR1h6Dcp/c
k3nCjT92TKCVLG6cmjFKvT4GVK8O/F14X5H5qfI2kMPVsCW7DscUtBQdQCqU
EDb87XFTt8im4ewpPZEPDsOmWgypTEgAkVsD4Im9w/+JU0Ola3rwIafCT8Ur
pM74MIZ2bp7D7KqIAPxy7vj9XoRdwhnrHBV5UTqqWJyGXBJ7sPKlN86joHWi
dyWRzZE/bI8whlL0pJzk5od+WHDG9w044hGJ+SfmOxLg7YMmrFE342rHjhwk
zuKAv8uJOi5bpEJJQXGJ1w4JXcFyVvsQWAfvhcamgUXnukfogdrdC16/AYUp
9kHc4J482VfaopUNZC3zH5sDFZFgEJq5BjJvPjhlxaMJtJyXH9HvINsrL5tv
5FoZPm8hiMqXU0h08tc1Ofa6/T3wFac/guYzgruGxjQ6BLx319GZssFS6wwI
zzlV2D4/+D46BL00lc4iZZ/SKAbpf8TVD4OOxEU8+9PQsGfIqbdE0ZD9p4Zf
VPHN9P0YW/WJK8m/KCc1ZCd+3Y4toqsYdO6jA17mqkL3LCQSBH1HMJJkXY7d
8uJ08EPzYRac3jkwlpCrfJx0q04UsAIbkH7CALdh+CCGxzvfRgaeC40ip82J
PSt2WwOFE8paegb9GM+4U8dP8W77M2OWmlwuLN9U+3CP5S6wfLOC+hsQB2JK
im8Yt8IZ7+OJuaRDkEEq+HH9A+eyklqKXjwbL1SfDhNqHOa18eZEKAGInWTe
GKuLDyq0qDIC01jb4eHPiAqKYtpmuLQ9GexUx1HwOQIwvbO2ZOFCBndAgdwg
tJ99rV7JMORTMKjw82brQQfImJu7asA9R8xGA1CBYAMZcxLx7lToeJrpKjzU
Sf3MmLVkAAPR4msNzoTWG/2nhd80mUKNAFwKaIjq1kVXiYn1ayHJ2t/Th1et
UY2hcCMfVSx+kUCiJ1/kyr1kbH7rb7ogv536JMcSn18LJ+4ZIS68k1nT2AqX
3kIC7+2sf0Xh3pexBid1qvbMCnnW/TuvE0GhIIXveeadg72XvUA8xKWgMHFI
aEDdO1crUxaQq6CHO6u3P9/WsafoFoHXLV/Ytwy+bwmCBtp92ieajjqCUo4c
JdJ3g4HCJvGKTTYIgdmPlHCSdO3cB/Zrw8YcrQ/zmu0xDMWpFnkO6hmvFgOD
9jZOkdebh2UP6OIVdQFwbHanVRhf7RSpX/smnMT0ER/dOL0aoegBsFUiUZEv
Mn54vWw94GsJ6kEMjtooV3KfQ8K6nI/8p+MZUm8M2OkXsvFe21bjjcAnb9Ce
GJdEr71wO9g6FbVYdgwJbM+OTX3k9BjfGmcBBAxQWGMyu3UjVBq6RVj7Nmoz
wjEVpVeBIIMrBwVqvaGGhiYVD3aAyk8wSFIr0zxdr4H7iqkNwte6aASytf5a
e06DRhSMqhO5GUZyGbDejEo0liIhfu/XMCOvFRahU3xbKr2cu8vwRF8ZYUcP
5ou4NYCxop0lRTHK4v1c6wrchlWS7SuqTWck97gTV81CJgWNJg/uUW/sM0Gc
Mfl5Uf2qii7Qvu/ysHsHB69Q4JFCLDtvMej4gDgGFIAFwqckBJezkFCU5yCS
CTAa4rGtP5jjlPicon0ya7VzuYN9cos5WLpzDDtYK/V3HrDY7SwzbjKs9oRe
J2epNiDCQpezvaJ07lqrle5z8FPUZlHl/mO15RUZ8c51fcHBmR60sYlly//i
+XdW0LXHD4/qAzheIE7X49tnfZNbCaTgvUHXKEc6m9M27wPnrRGHWrw2Qdc2
xV495g7lZGcc9dkItzukRKMeA84N86ONHtLltIe0L00ZGxqflSUSZ0HQN+HF
PdOEpW6R4DdJGI/aXuMTBSDG69dBemjjFL4eI5l4BlsOzUoW+quEZWaGAXgX
C4LMP6g7xX7+QMxJQc35d0lFdT4h+HmcmsDJu3KGUfSQRXKwnAHZ2H5vIffz
0dzeoYmC8CbD6XUcUfaPtn7kyKdBDvjarsgFG9MTlj7ankG/yqyvCramwnyy
Zy23Y+r4VYzwkYZf31UbaRseRDpgxh+saxBza8TcNvgEsiUG9B3LrovK3EXZ
w5alrlNb6JFkuTJg/ZM5aeBDPxR2I0e3quZp/3JEOwFkw5OLmo1Hg/yGVUgs
A3S/ANhc/V3Fdvl4LfkOkZwUyB6F2vnk/ZzivGfi9FBMj6tnyooS2H1ri+Ls
fQlyBZnAMEdf70WLRC225GhJsqBqszS7NV7gJ9jLMF1Svr9UaSyOumxxqM/R
8xPHFLS16ILdNhGo5xLowy6JUHVClhfj13KWiHGJ4wn/4UoUhS15v5KN9mGg
nj7Uicn6gqGYjFnXAgp3OjXfPNzHCcMFCk4wsH+fKX5lGWRdP2dNuD344YaU
AdlPLKHKC0Dz0bCZwp6Kxpx7txFR/73V5e1ljVup+w+pjoGAqINoRRKCULUc
D1XZA338e4lkf1trHSy8yhQczFYE6P824E/shHGB7KhMBvFWsdHrpK3fbGjs
v2heHfGLnXHghVp4WpeBs+xqImfwbjpSiKDURTQCkqWo5xoXxCMi8p3e5tM4
gfYcylXay+oLorWh72hpwXlQ1I0/znUkSx1vnCVC6LiaJ11Mggfa4kDwMggN
QEvKWwyEa/RDPUzQv7ZOS0bFCVtn7aemiorh0iL2ySJqmmdDG32gyZzA0NQ0
2xLA3a+VHBc5X5g+cRKEJ8NwA679OWaPlfcyxi3TRP+Yw4NG7/Syp0ycXYIg
+ZWoXugJFrvPzOYrL7sOtx5y9zPns4rXFGksypUOaWUq8/yeubI6iybhJGLz
nN2kwQuAKCe7QG9crLSHZM1/hDFw6jFpAb4ZuyNxrljjjK8XCduFvDfSwQiV
YdpHxyVs8q2sKGxhVh+X1KTSRa0qO/xIYeHNqGbv62bgOcOHsO173fNWplf6
Ln/efBYqRdbild7iSmOjTrv7bBTksEDMTsOrZzzPQG26R/VJqn5f7HSQKXIS
XkP3FqBhSloCg2ZCl+j48zus0Ks35ZFE4nHpFviZZGbA/AryUYllyDimNubz
b8cvoy3qnap37HRRFB419p23DbfngkY38wMK84tBiy3BTJwb64uX7aKzpVrQ
w8R8uXNMmbSuh0fEjXLE59qgIilYA7aEdYWCtVkkj1FcfB0YyTRSmGl7Gs9C
7hC5acoKXRQj8kkHLTqKn2l7rOjT5cK48E0nXa2i2p1cQOKv/zHsucfoc8H3
GUbVA8KAl0crwI2LVTiZfqczhEDv3bVwGJU40c6IPBNuu3kCmou7ww0iDjKG
2NljbiqxCK3ludIBDkDF/bDmVF5q1EGrggpMoCzfAgWecRv5/M7g56Sck9Tw
vLDD71mALSG9mjMeii/SCKLXDpPdc3Ymu1XotF3eyD7ktHFgZ8KFhw+GBd+U
CJqbkDWszO2JFq6T5qjeABKqZo8WnVMPsuVkcST3s2WOblIG1/1cn9XoPKtV
mcB60ZLi5xV81GWELrrbpQd62cuW2yn1D3qFAzOKsG/+waibY/iAwZ0Db3Ae
v/5HvUbt8U1UE12mVu/1sbd/TfHOTZjZBFgB5BZVK1fzRyqfA9e316crobmN
+ua3wtL2ZahNBpPPITY86a/slyE29ygxJuPf4DVDLJl/F3fOVuEEHQaS/mVP
8+WC5j0+CmTws79YWk382Dx6CrBtJrtVSLyOA9ZruRtssuTiwsuLVOUMBdrz
gsJmSXVD22t4iDdz/1JAb1Uf6li00XKu98z+aaVgZy32NjIspDEKaiNs37es
c+QZz4mN6dmpRiRiWbkJEkWXDK7MZ+6sVCxv8XUViGHdFWeuxWfmpvHgbxRu
1iJQSPzR3e5hekNm3AEt+UwqdyXb7je0P82JZww2UrhzRvFlZCY7zX61+ebG
5N6lx3pfKDUC1YRI6a00SyU/RiuSfLCn9bBurZoRqcXsGv/LMVUKU+WldYkI
5K42mlcuMqTPczw2AgNUaHHimZnD0125CHu5ueavuYFbCp53PQLnONij1g+U
qyUCQpogzzRYAz5c7TKz+3feBE3iSU5VmZFIV1uvu1TLFhSFotgOzg3Y2YnB
vIpV4hDT+/MTzdd/6rEv6FRLG2mgJrTvbXVJUewOOnULheH32Ad0V00l7ibO
B71xtZms4IaXfjRS/T39PWi9As/mV+/xcaWKauifiL9qH+ZiBUczbAtJrBmO
8T4gGmwyBr6f94ttd+eMQ6ybm9qU0E7D1KnsDCTwfs8drplHs6TrDo4JybpW
cOo5NmSRzYmzJEJkvBP6HeV3yccjkKI74NaPjl2dkdJlrI6Lk4vbkWL2mw9i
/E7tpgf28DoJms+89+Z4HqVNwQxlK6rjIMmTaV6ca8szU0db/wiHPtATA0Ji
pPyPZv/lHvkjFPQ0CxcriTTVCthXDOTCnriVKzgHdkoUkZoyrY1QzhANS2fv
gyf0WspmAjEarFqVaKURhVX4tqD75BLzIhZpDace982qcOzJvmwhvTuUeq9O
g8uH3I1SmLK+d1mQ4Le7vHPbCXm+sJv6CRTajBRHRCZb2Dg904IZljKAkc5s
Qz+/0PUXy01VDoGW44N0CZa2jh6tSt0ugDQHkPQ/1973LNG2VzgPg/cHu21X
QerR7EfBxHQHg77b0yW9+ts0LOh5SXWsxMISnUcSHAI4WC0Lq3nLkwjKO1Zd
RiHQbudKIIeU8iWpcEWb2QhMRim8g1rTuen9kwMn1SYx+z9V2FHm3FJzfbSR
/4VFCVfw9zA4dOlkqsnJVIwhfpkLwa3Zrt5AveMynjpeARGnBGKWVvS+rQJo
iWQeTEttV2hacjvdD0ksqymMFR9sLl03Wm7aih1OnlCzD/V6WCqiq+1sTADi
P28axWL6RxTc2zfUIay/WiGnAg0BbN2Z4k8TaAhMoO8+le4zMYFSL3LU8UvV
LUrwNz4e7AuRyuKJcZEfzOm8l52/5QfewZTKTBlOFGfKidtu2jMY/JFwJNjG
CwH8AM6g3Dj/RI5ahSIMfS3LukDJtCXIthR+1AHiCKvmELUcBc/kl/7niCa0
M2NCFdOSvKvJ6B3g7tCcPsoXdmkFHQNytle2TGRUAek2ai+QBPOcaBCY1ZRD
L6Opcz7UoTYJg7aZnEXh8NbBxxdHXabLpCCyTrHYSHb10qA1SjQ9OiZW7IGU
T7j1YMR+H44egtQXBlAelfmBJgkV+pSIMG0J8di6gVOMlYtuyJZ9iPlsvdBq
RIOgk7UnunO1QPKVHIwn2xHuDSoHx5CNmxfG9tgMNBuTI3y0E98bZ38/jlk+
K032MBsl/wlUugblUOiUEOo7JhG63Xq+B5Knq//NUIYjjvMWNRD61rSJ7GFF
+2LyLQyKJlRLXuEvFgaPum4Ltvhppi/qod9euKaCcAvIjb9dWpA5AdvAMP4E
EJl/63XjSi3jCrEXvIsIbJIVg645uUEg1KFyWfyb5HtMIDPyNhG7VaF3h2Gb
yxVzhs9M8NMx/FVpMRIemgpzqkCrwJoz1wQjgpEzocPFW+/KYrvQlmT8KUe3
XR4JG+fGgKyxQ/+xcmpFZPqykILUsfKChV7braiagiAHVIdgB2qmaPM45fvS
DRbaGFvd1JyocMoFepqHoaKKr+ImC6IIVtn+Flp/fwxNjrTaiEsVUNSQcMi8
b7ar4j8Fy0JWkOe/2s4Je2bb2zv0t4F4LvmGAw36e7lZWdwoDalzXnUZ7TW2
21/IKGi0MEK7z9m0Gk0AtzXT/vTvZ01WUT/T3U8x36AmK75WoGsG9+HuJ9DI
YkKDUXVrrky/NpoK86abzRD9CedaWt71AGLC2aDKM9a5krycksNDK19UoHDn
gVz+PdMXFak0lG6URnptwWckmwe9yRH3ZnpBYcZvaC9TZNv+RKWBHZvUbWM6
I5hiZWStgpK7IGhdGFLsadJ2BhTQPwaz94VrEceCGrwCJXjbSTVxDT9nYHyW
WnHNIg9FxPSmKuWPve2mPghp53yM+LnEafXIMoH7zolSGMY300Fba3McNrtX
u+KOtJuEBMySwHIUQKatqk/SXFU9oIvZTfvoIGxzIMVEUCjboTJIWSigXnq/
SAoTZUsVcuw7GLItE8aHFjUQC6p4V1sCkz66GsgD1SD2AnlZdyKeIaOwwXf7
fTVMRB/hQw6nNrAWtp60v0iB/rJ/ua4PfHMEaEAj4G2LivWZmevDg0QnBKu1
/ztSKVBMS4eC4s3tCPYaHQKXMvkQ87/9GUYnn2ytRe9SbP5NW6VIhbZe5PiM
1CbXEwBj6ttUCsc1T0tOLKuBw2F5NJf0W+Ek3o+7bcbedsxbbpiBG982oNy3
FjRtVMcvszH8KRvSptPN6sgSzW/IDOLHeqf163kgKhEri/ETWOy5imlSKLQa
HkW088mdJT0zlSOv9m/eC7eE0c1U8zXUIYk0lGCpVhgYLiIRWh+Ty8YapL4V
63BiSQ9SFANCCNasI97G9mh7CjnTYL1vRBA9SXpsdFtmK30h1VV2m8m3lHB0
zfci54v/QduNEFDaufBmSajM1WFvwaUdnUsJdOK/lUGllb3TXrww3Zdn7CU3
86m6c41mxRqYG6mhCN1r/jKimohKwn97AmQ7tbb7OT4BW5GIhmjvxAWE7ZEs
hvDF4CxaFqVpxkt56ZYSPG1aW+dCpIr49v9DNF3X67+Z/HecXTCnO/cAsuNH
f970Dk4tpzmejMp865sRLm86SoUzmJ3XECyRWu7IAHNe8Q77pxxBHxGdisgO
xK+tCrg3lbXXwr86kBi6SZHlVLRsMPaxeNK3svInFTGnkI5T0lzpuQKmSBrE
yrxH+4iEzXXeEUfVv7KMxW5DmEhvjzShKccWkh/U4gRBsoXa1LnhkHX48Cb9
9SFAkHMxtPbJEMbtbWWBhb6HC6/39fCD++VNrOXYec0xEl+5j8yGOg97gRnL
aS3vqqT8rN1sizoMKx9137TR8jX3EAiHJ0w5fe74Uw1rdNujebnakSFIFW2u
Q5Syp1PWYj3vjOh6XkkZMpQX6Ey5Stuc2WZ3kAlyywG9dNnhoHyjetAgGQxF
DQNS2nbCnsRv+9GfymqXO0oT0nEAPSkQCbwjkEUxhATiNrY78dH0PHfPAkip
PInAXkoMz3Eeq8xlt3XfMzPNGhP+9/IHJmw+IQ+AxU3xdRdyItyeWle/bNio
TbtFUys4tPDFGClIgLsg80z31wWTG+2I6KVrj23gT1kdW6mJU20riNZEhGdY
5/KqPQWonR49ob1Dou/zkQ3ReD77i5edrpW+1f7IPeFJDzMPyoWoWzIjpy+A
6HcsNx2yQ6QAjRpIhKO48WVMD1WaYlbweuU8wGu1y4u4wiRXTQTt4dxR5/oF
lnEMVDHHpgcKKNq6gAx76mx0V+Ql3ZNIP6ICcHxPA7zakn3JOvZKDH2X+gmv
p8tHdXr2MjjQ3z8nzj1c0+FMRwIc+02ITXZRLAskuHYHDu5aRMQu1tMq1wqx
w76dOsuJa9D9J9SB++FCHriYXRoYym4XEXi3Vrt7/PhYCSLm2scs5bmYZqTO
5dOldhrU16Xn+6xMHZtEs6fBTwH5Ke1LhUIfN1oCygmsZhtaGLGShQ4RPkaH
UaqFGLOxcKkJnX0j2PibJZd84bhieaQrWIPduUzmxr6gMXSVdUitIivXmr/X
dLjdq+xPu1PdDHcvU9SVsVSovUvYXYhBljn6y1yaNdpOlb7lQJBoA9WuepKR
y+fL6c3WOAZceeFbYh6TDPE7nFinD46kE9YtVAyVpBvsPH3mLYQUKvQqhCU0
wvzcwtEHMig/t+WdCH0ENmLGdx3NUm/osyC/c0e2kGOkE2YfbZRS4TwHOpUx
H4S5FSuhDqBjoU2Jr6OaXFXQz5RGhlOIS6d407me9hrd0ORkc6RxAtqfso7e
n2onJzsSK7US7vsbrXofgbd1FK/0fzQgkOqWLbL7dlFoRIwUeAxuAJ7vbMlR
OLNjw7HkSe4AWsee/Y4xupvxV+Qkxlc3bAuSg8wm5bKz1DEUQaoeI/iT59zh
fW2JlwNlR/haxldd23xz8kMMtxgRtYHLEX7Y6hl8ao4OR2ddXKN53hAkdFdA
mrqoFeeDn1aByF26yJFp3wvnXm0WA210TQM9bcuBX8ZAzdH7Di5z6Aa7MAI3
hXVfhwxuenEIl9GymENt365Ts0LJoHZNqVDtoVY+oiA6JHG+9jo8JbeuF4d9
U30KA4AhlOiCfBSub1/LvAKxCjXdwQbOba1/u0Pr452YNUzKNhCbs3R2fPnu
Rxl1iYgSKJwtVNHBznsumVNuwJIA7OuUGR2xZftb+X3DizkmMZwY+cJV0JWG
sgRxJs8rl7b1X3nNcOmvGWkK0Hxp/07qpf8mNtFq9XrkV/T7jxrv4/v3Ax/f
1fV605yo9AeYj5yogGXXXRYo9VNI1+3muvh3BeUCxqeannIRq0FaJR387dzl
czzk6pCgupEasNVC+DuVGuNDLGEjNnNDXFdFphEY8W3KhFgDbON2VFd03YRm
iiHyn8fmm2VAsKn+1rTybK8z0H6i4Wy0jr2U2LuX5mpXWMaLD2sT0vBtveQh
/xB4Z3D9p/oyu+Xa+a1Q5LDLbyQ3cSq/j3k93XUAX1ypi3M/LLxsepnxhoQc
ZGIyCYROj70eO6JDqJuVVJaFOPVx9OA1aq9WSwA7JClIo8DNjoYY+VHZ15Ky
7d2FObIJnxsdtRHzMbO69pKV8Gi9Xbt+hVsQV9omnZ0MyoLUvyGmOw/paxbB
LqKHf0B+XOqafuuZv11AJi+/7uxzhrA82pGIMaeZXlh8om45CJuTPk6Kv8SF
Ox4qWGFyKrAqrf4YG5dQ11Q5HBgKYvAOaa3glGRBtpevhE5qG1RRRJA2BMC1
7qRin17oZAslPjS/fCgtkysZbTk/8TiAFVoiclC2TqT7JqRc45ypCaXPdDch
MvepIZJesCBVURmhlCnReP+j3plB67vze0jpY7Qgp1mbkHk3x3jq6fBY2Kpj
sFIBAkAGYeZa1fwCSG2wDBXLj1V+cU+iFWRADgZ96h5NkYgstKGkwhPmvHXL
Bd16SkwvAklhJbv+cyaMzrK38c9OSOV1qPL9NsB9S5ksHPpzzxjqzsYLBGWV
wUCXcsVpGn1yYntAfhvZRFN0pSGRiY0D8iUBca6JW/nSJtquJ63VZktyMKoQ
4TFvx7KeH+zUcQQNs7KPiyHHSkXCxHZffNjxP4MvH6GWwr/w94z+nMPmUd0r
iO1fXvFhrMC5hmAASk+GOCNH/UwZ6iiYHLvFFwA23MMj5A16UNwuQpn28FoZ
En0ggc0jyG2Dr52sNxvCE+wO2+jNb++sUD5ZqmSz64iZQaoFThNI0oNJ2UqG
Yn4s1gEqd+XnvlqtcLnidosUhSsnksjTlQJdSHcfVgvFwNoYaCKQwCVseX5h
+yRpnz47B3RkEC/nOnmoYB9Fv2GTzDLhNTLdxr3+F5xTTX3yD7w5rVKRH5Vw
w2Z8kOkJD7ZAt4LxpXUri5oCubkUEYpAr8T/YpWVTsKtA08qgzCUaW4pdNsd
78hEP2n8Bao6nFmnrQjjB9nMHyP0X2+m/lYeL00IOhkHASAaZTQnpymfSFv3
tYL5IfXQaxfYpZXcNi868A5Yx3/SOCZfvk1lri6zqIUn96o/lzThKBocaeWS
YcLrdsnkZpiysddxf0fMovbOhSFuMC8f6WCPJf3jl3lD3PE+gOYu0Dd0701x
jCNay+3t3iXPg9DIoXwDkdlVUjTfI1Kyj2zHsPVAM3qfnVtGIydWpghbXBTb
2lmu+Z66M1GO7iKnLMc/OW+8Tf0wtRsisaVcTqIVPiRYYhUaY+TRGYBnV29Y
1aHaNRoDlm4cC24o913siFHfm0u2IPCutEdzxI1jge5MT+sQ58ZdwUyaSv2Y
MKPMriFRaOB54+9ku6pn7pTe9KlNk0y9RCTLFRler7UuCFXNyA6U1nmJ6n9U
AsN64IWY4FZJc5VRSytw408+7cTf85gTEtGxRZnTpgHMsHJITxKp/Wgf1qP/
x69vMM/FQlwSW/bNDiy49/37HE4ZC2Tf1+mpLA9XNLsHD9meFESLavcKqKyw
HIRNksXZlSCqPLwhKxpejKzDr4WdgwHtKLjp0oh1Ajd68cWc/hOrIiGtTAOW
PaycZaKpRQMmhvxrRh2HwZuMmH4sETB2uv22WA1WS2sdolwGzhVkTUQgg6Ee
qE2lp8dcCnQCnNbmvoOQYZzDgeps4H5pCVTuCskFLQhfy/0AqTcMeR6JQ+X4
kIcTir0D0fYThPiCNEhjPaKM7QgAfRsw9iAyIBOYyfH8mUQ6nqCyPdhnDrM7
43T/X6oYPdVw9RI+oms8DApJ7rTF1RAFq8an/jUaEnq5tBzzZeWEWMyx4ux+
0QE47HtVBNTPsA1dDGMQHr6yc2+/N/AzZmWOzwobWfogULCEBZmaBaryAtox
Yrutrb4yyUqukTTJJ3MLrBZltrgKjdHHGQcGwD9zk7SBbxD8EIJvMrb/5deX
3M9UMGj8H5FbFW1rwy2VtYmKr4anGyRefo8oVWCt2uJDGP5cVfpCqdwUbgTo
Vf89Zk+8DxOFyM+qZTG/T6KqVRmeEodJ+NL+b9tJ1AEHA/yJS0duWGt43bpV
805fBCjtK2XJeVO9azksjwE5dwUHB+tZCVsjyHI0wBt99ZmUH01HdWXb38Dv
dm2VDI5QV8fXd57WSehihi0Cq9EdvOOLg0RkSYNCBAkVg9QmD6xKq5JDtLGz
6kaB77dCzylmd9MdUwIgY0KdS4c/Yz4yw+hQ/w4R8BZYFGQtR7ziDTUbWZs+
CmNSs7ofy4pAvQCX6V1ON1MS9zhmbN8xSRY4URyeZKF21qbMi5rfHInYiZ4L
TQBUWRbBD5AHHQvw61ZVU274t1sduh8BceCNQzDci+SFLojkfHrvFRSt5GRc
X6TC7f0qBaOm92MO7hjfCbTZbL9AQFqWnUBOX340j0zLpV6/TkMr+/XvNcWb
Jkz9JG6dcsFuiMt5B89BiRW8SOKeqiu+zYpvLOcTYxwWglK3DwZrzTpiOMSx
k8nbjgVC5yMjgA3qkGCH0YAWvZmnkVLNMHlMnqNkL15wyJIWpeT8sHPbKZGD
XLfO4wR6l1qqj4SFQ4GNmHsnV9++Iw2w4o6hlFt8RUPBKT61xn02yKeuhQax
JTziBzqZgdwFtenKssuSfzMSEY1cCMzVpGAo7/eCkXcA32HT8pv/EF32QQMd
dx6Qj1GdAqSpB2sCXAuy3vkJos7j9eOcpm8FPFl4S/GwtUJYO3tcphWrUikc
IWJQq+HMK11EJ3KDvlxft9rzrSv6JtOons8q3anOGfet67juMvj2pkbJkZWi
bBNDMCdwEbAu6/3Mvic2fx9k6uyUKLHPnYuqN3smCGgPthfk251xdmXh1q78
4QBt4sJHR/na86Zg4rS4TCq+3z3iDYHym6p2fAr2NucvJfkmocCkfcUAIsv0
5tkJhrYYQNk0x9/N2hlZQTlo0kF4S2cBJpqn5v7zqduhPKIvcwInwG8Mq2He
n3L7QM4Lbnd9oC8inbeUecJMjf6tUxiBtVa0F281f1ZtvkWw4DsoZmUUXxa/
QOff5jMCEvufABFIiUZ1OOWLmpoudnw2WB6JEGnTcRivOLdwXB35OO9Qn46c
ck6OsaP+L2RZYoVZHPzvp7t3Y1PCd/RKd09n54PccAQKdTGlKVYlddv8wLdC
TdcgEP8GYK7vkQBv1ImKoQkRZEkeO6EfHHhcDyy+1CdJhMqob274PpSPZ9PW
NDvJQIfsPKxRPWox7SOS0julTh9KxfB2h7kQEpLGOnSThir2AZErTZyV+zGY
8xyE5K2T2jbM1ErnqzIb18wNsIJqKrMaynEHkKO2RXk4aZhnwx+fs5EG9QlI
sxvFEgTgJAGOmVUJ+0nK9qJr7aB9Rtz7NvCdk4WjMNYLuAwS7MLvkeNoWU5f
e6zXtToj6QNimAOyJHOsE4JceYIjsj9mg3cGCAYuTySEV0uHYVBxEGEk8IL9
7NgdT5lDVoCi9gQa0AqwltcpY5Gz09cCFHS2VFWZdrkzxNA+uTd+AR/gQBYC
OZo6HZ7eCzSwTkBHLrHYsMZRjfWlu6J6Zw9/yH6LDf6g0XoCPJyTWIW15W8r
Qq74/ZcP9wsgg8M3IYtk6JB3b7cnsGDKFID9DHlAhVZWP75gXRxwfrMFqiSG
kgmztZGV36+AePG1tkoAtRUiAx0N1qGRCSzU5QmXNwAe+qjW9ZrS9ayk25ff
GSyuv5GKQKk7mwfF7hpCPzwHO9S92jBXaeDvdcaibjjsLs8rpib7r0CJBSKz
bA1Crd4yI8CAzATVj+CmFPvB0+5JvXExizrBmek6U0st4NMWdxt14tVk8qHz
3K72WQm3FQKeqGMk+lOMMckhDKJfmQoiH6EUrQLAvHzzQFo+k5g67DOnn7Bx
aPSEgMh1MavlFgoE2kGfLtgzgTc0siDLhAJC3bX3lzEELajBaHbav0RvHfaP
uwb2d3Y5BdWYiGPUN3VFEp1ieI7l4UTCmAGz3BpaQZp0+n+bBy8sjHmxmr/q
BbkUkq/fOhMNlvK3OFMxU0u+0QREJMJdf1ZBvDj84HyUiPlQ7Tkk/WzicuTW
MEkwNK3GQw0ne+gBQYA7iUhmIb5dHUdKlueytULFovOAICBrt2sL4a9bXWS2
TY0RjknQH6cbKiSejfT9j4ZFqOo2iwpIh2jytfnCC2rroBSaAb6HrnKD7daU
s/OYwrYfP7cimFdRVH2PpU00fndW1wu5wg5iqTAB2Baaaf12RLi/NBakyDaN
l0fyA8QdewgU2CG3VoViTFpq42g8lT44IJK9NF0xNemIrEHhAKy4Ct1Fk8dM
zF40yixTm54pQxN1Q+1XvKE8Wz2XdBWTSVvnnBTsDvU0pWSxdX1NklF02sGK
Nhvo+867R+LM8VQ3sGToeiUteGiW2k1xC5YmtMzXGVrQQVrkvysQyyMFELUm
vCZQBuBDUkMHCr2YTxhYkmfoaW+zShEWvM1bCoq7PFl+iF0CWXFRn3yPjOwK
0MSS/xxC6XYUZpHSEfvZadA3rZzpYyY6N+CAXn2EodqVh4YSymyHcWKMDGRM
PuXqAAbMwRfaq+2I5uW5QSWbkNdU8IqjwtvZz5xhFPva84r04DAzAG0ewiJT
VW1UB+qFheSVVVSCYA7Mkk+5kRpSqPVSroMPMfafgn96EarhPEpblGYnu/Dt
/IavrFUvbU9PZkJxnVkoZVLSB2nEVYP9E2eW+UmBup+uuglTVyJ3+x/Q5TYW
/ksbJN7VfsPU/c2hZze8rw+ZDt8pzjmq1bomZ6y2xL7Ac2/j8SK42I50qncP
4x3Pw2RLNzQvh8/UdWFtwblTnroXRjPO5RyIStm6KOO1aF3t6LBpgnYD2MOd
f1Dijd9Lzs69v2Xk/Obil7PDWcAbHx2y5mmSrrxRxqwPnjJxHuJISF+TDI4Y
U3/30yMRg9TdtnjKwwYZcAmpBLhhmTfhyb5vGzZzyRblsOU1WFEdzE9G4FLy
IzCJvh8FyUtg2c8QYZaHQH254r/5lJs9Ia64MU5aRErS9ml4dzwY57vgc/az
Uir8b0lhRVYXgcPx0q+xo50vQZvpu4MMgddkSp4ZgvNYTDHPwetflwZhYolK
8cC/24qiFfY/Xa9h9FnOQBvnL35PW+miFmLxULXE6xelp1WEU+iJgyvDXh/W
Af77gYfDcZ0z5ec/MwwmVxK1qmhdm6+YSx00VjShD2TxwKRjTNqVCMd/Zm2C
RQ+SKBYelQY5H8BrECSDxDDKZEHdiwt0uabuUNK/CN6hASbHHfuNqpjUO1tW
+QudeVH3s7wzsiCPMMv6Bz5JUe12PYoLLKPwdphjuR3uOGetWxjFS6uDG8xW
YantnuQKK/gB072wEj7VboE4ZgS1+7OF741QoyjUZj0h8TEqyzjI2x7OQoC4
eLjlRZ44l5+I9NKdDFIPEKkZ/WaQ/0ue5qNxhIdJvf7U5+IiQF20W7UKtf6/
RW3+IBVD6+HuVLhMxYiG8kkikwtbQNG5vfCg/uOb0s1ybbUT07oiMHWikdGH
aleeXepRKxPIaqG3kiHUaXBsNBMcpJVdortgu36Ck+F2WNnFmisYiuQb072D
VaRA8mOGJyIBdfKdEsrP0DDORBIWUjVYtnxDHIwtqB1pkT7tgrlpd8zoYKYk
2+noIzBA7Ofoql4whQ/fv4vqxJ7RDOIL6cGCLI9HYlR9WPryUUCVaLGCKnSL
cj2WEfkOu2nIFpFoOBTyHmaTGJgXPBo4VYVkKGDad5QgIJLRPlHJ6NJQ3tdx
l/mQSQAv6CteopJ7wOcfdk0FrM4xDZz0wBVujSJ0s563x9Z1+nICzwbwYi+F
ExO5RjNwOhuGjtuJQzBV3MM29Fw84EMfLgH4/xi1PuV/tSq9NU4hraKSYSDp
vfYl/jYWsykN/g80QBRBo9ADwJwnM4Za/gSsmVyz5m1uWCMNckdr450MIokz
Olhtd5a/SF7EHiAInqgEieR12Iz1qWEqvjGNiwj5cWda0RcIVDknVgHzQTpw
idQPiNV1POjqvA3SLBpSrmsY3CHgUt+YaNg5gqTmq4W/BZ9GWYq/UDf7KMYp
kuSQOqMPwIJb2m7JfDdzmW2Agl6iKLo0Y5YAwp619jYq9CSr7yAgycPaRj7V
2slqucNaDX+CRJEcZo1FO0M4J5ozYGXEYhyVCh5pzlakWG2auNt2UVpZ4Aor
NJ+rM/ixdijg32TDBxsJVau9VCpncfKHCNj9LReAUcanGPQBN6P1RpOp6W/X
cZorEnpG4Re8f3jHY5j0R0r0qUjNyrdMSEfjsqpH5NiI3/fjm5QCNpr6vvkT
Lf9JzgiGlA1US1Ax7UkLkx01IXDYfPTyzl6Ff3KZjf1Fx4b6liL0L8xFoBSU
JKio0BBAGVZ3NZCIKSOM+DS0mC1JzVHSYo27dfBnsx4qPHQwkAsFCkFf2oGN
GPfECsAg5rWnM8nsBqQVEg4LKOe9ksMCnw2lEA9YNkmsKjlVt495JkFgg/rW
+Xh2lpD+hXmoeyjU429vu6otMnoYF8n8NlzXxzeUOX4W78SZmxTa8MJqIno4
/n2GLTca+J4L1qk99Ev6EbPUe86KyAr8UNu6JvpYLuFhfqXcudcGGwMIEbyP
GcUMki9VZHYxXbenQMGx3ez53T44jmgkTfUK3GQ0d1UtKhYegxTZ4NzZYfkT
TnJ5sPbHFV3jtfVybZXeinnM85yIMTaM5QZXwZhYtGz95TWhzj7x1raQtPC+
2x6N0P9AGK3KwTYp4MT2t+QIbAOk3i3KkVWR2pgrDGQnluouLuKjvbBuIOER
HhP4FY9xR1qVHWDzLd/XCzJ9+C2n+9hzgWg/WTQLpX10Fg1aR4UGlHC3XWfM
9lIAyujJ/y99+T4dnLu4N7RCnSZiWW2YQfpcT/hCcoOngbN/SldsXLLNR9M8
W6GCQuWFYZQ0Ecd10Z9MgMBL0XKxAdqF6ipE5tRr0ddNEcqjuhQrI9/El0SD
njg6gH+QUjYp0RS6HAwSBWTasW4yrSt5YVWvPd0diNsVGOFsBdnFUVIlWX9n
0Yiswq3HPn7qE48wauSnLygZYovbe7zm1f+VH3Se7b1IGvRVKUGfNf53zzrC
5hyTZVmfsQ6jHuhecizEJgzawxTHMI2lG88QGEm5Mhg8RLZHgxQa40DEGrIZ
XdyEDSpRb6KHE7pLyeXCZw2mNI7LvMBU7AtHWb1DTZ+QoEctu29WgBnMOtCx
VqerbimgfncnVUK4cE1GcoKlTTAbMherd6e0Ch8h9PoTx3kNHpWklcSoBlv+
xomobwrdJDkR9J5DD0C8b6LHPi8ODYpbqZZ/JyTVWQWCzIkBRVm6cl15XjAW
aFmtV5t61SkFpYpP79nsDLvEcVQAYhOyaQ8wWm4yatyxTFBxpAsvsO5xMeLC
x0goPI1RCNbXp4o9Iv8XAtoFjWJJmU+hOwEBzcOR0Xs942xqBFFHiPE7i0XS
qTA38ddz+H12ULoTncHo3qZyUhLOM2f/G1Blc+UnwJvZi/gEt6YTKMyKT4LY
lwacEJ47d2JBYvQRADqH7lcOBGuFwwnLHSt4WdRzHNdIYuUqy8ywa0K3qNks
+h/BsCfBOo+zmvf2iEQ8Ki2pChwK1E10xVf4SlT7ZMkscDtVrU6VNHBNcM13
wB9Qx9WB7aSP0zQzzatiFZic81jJqZ1I9QBFh+2CID62XYfSsSz1t3DtyqvC
OGZft4fPCdJ536AerQWOg39aKuAdEDMKs2wa4N0pC9hnUK5Sa1hMH/VIhNO0
To9BddvQHFROoCyQTO4hUEs0jxXdbXMjR+0wC7cWNauwlio5/CPMZ4c/XkiC
wy/y+o8i3CUomhw++X1+4vF5d0+AR/8QQ2+A4xeyVqXipGMrpKg3DqA6Kg0L
edc5K6xcVJtRJWb5HIGUpwyI6GRDgOPQVeP4wQAGxEIPMsypG9vIQHcY6jna
NozhGMvgi+6DvSxEVAnqIp3eqntV1Cpm9Prg/0mS1jLqPwZAOZTN+cex98se
MaQQuCOU6SRBa7I2ZUaP2slpLq50UH49hiMX2RW3IyzW8TPWonglfXJMqWC2
YDwVa36dHPVd8zVeAID2BxWh27GsypIUzHxjGpTXybRmlO2a5GBbmIWxDlZS
+F5tvcB+a0b4IFDhFgRHg4v6I19wNb+dXjQ0vF1Q44xyWCZ9YVhehB4IsKK6
rJ07tT1BE3Mm9Yq8ZSqzVawVslOheSg13y8ToT4tQBn8twCt9Y6DKr+MaZ29
XnEzQK7y4gLSLQ+/g0wr8Dbh6BYh9T008imJ8HTOWjx6zCQ5cwCo2op8kgUV
rDmQ7ztAy/Y1YZ9m1e0yHMfcEgdocLTdLeFsJLeLw4wXlyeb7iMGpm042Y6K
tq/4jFr8aNvuroU/y1UVU+ar8996FAnnwlp21HX7NO4r+oMw972OITFXFDh8
ahLW0TXjj+jFPstOHoupkaBQFwlYUA2Zf9G2pjYKMcSoACLZv/au4LyHRELX
H+g7QUhk3zKwt102d4mtp7XVg+dOy+Z1d6N3b57XuulgpkA8p3ou4VH8uL6F
UE8uwBkyJ1wz5I1yS56oO54cFJGd1PUEov/hUrrZiEDLj4DOw1mQEimuE5c+
85APkthWvOYccH5UPCzzf2IBQvVz0BYtdx7UGEupiqsjBzmCJelzvBcHqIAw
hnR1iD2OOdnqer/c6pz2UOPmZvMK77UnF4LSlan5gFoUxGttk1mU7vhVDOF0
wF5sYHZqyvrAPLME2siwOXsejvLwh0kxUd14XgMVK+YbJDOsEBlgKwkgA5rm
TTqaVGMYFffDktzD4xN9MfCPWwpWqOs8+aFhd5IlFvI0LGWHDeaPB8vVTURh
PhaTTwfUAkSRhjoD6+kMDIHessBQrL1jC7kpNGeVC4D5y61HYa9HA0Cjq1KB
TbHFzrS9a5DVsdFtUwRLDkvQ+hN+Yjnds98ypoRu/mIRU24ajJwEmZdPD/3u
GJLZJJw4taSagbvkZeYQFxrnwLCckIJKX/xuZ7ENY35FvjpVPaeGLLldQBFw
Q3RfvTzlSmBzqUNgcJ/bC4ZykIr0DuoJfSdtcvhvP8DCJILSedBcFZDjrEAE
KB7qJoQPuQOn6POF5tKAI4O2lC/cUCXkfAkOrlQwwilcWUksnh/X/G6lO06Q
OpaMPvYK5yYsQLHYefX5E5yZaKPKQlHQcQ3VmPXbNuXJjM6BdxWOu6q7McCp
kTVwHTNWfZq+jeR/EJIbt+Cb6F0CvtZ0zSH/LXqkAOTVCUR21Zkmq8+aDcQW
V05RyvkOIiWddW8Lo9CmFzMogcvJEo2s9kDy4ebmVPLeBLy8um/Ti9sJgXWa
xV0xYpJsatvsN52Hw8rA1pNARPIHI6klS/UnBXP+IOU857az7BVB9RsX48NC
pY/uVc48tDaDtAuivoG+FTx/HI0KDgOd3mYHKHSMeME/bUPq0ro5Ce4TxwEd
5AGql7l6hzdLhli6OhBIbPUkHsJKnNnEOKKLpmRH7/Kfnt92PkCnmZP4F5Yh
pCHPmjQhB3oZqs/q8vjvCmVWRUBZOHJyybTuayQze1ldCyyck3fj2rX76U9Y
+xPCWFf5yRudmLvmJ8xOVfCnaZlMGZsm6IvuKrq1IpqRbTmLoqwaAGsxZF6g
0BquD7m8G/9Sk1d4Wfp0o7EhWCYEnfW7Pn73McIBdIu3YttO2KJ/Jia0md31
Dyy1qPxM1XFe/nVtOun5+fbmhFELHOhtkK/l47mu1nPSMB3usiwMspF0Xm8y
FGOlzjv1+H+zI+QJ99/swGOnPoT0egiX3ZZpf3y2hoXCH4+xZ0gYW/F6R3zA
HF8QolY73tS+HY+HQKtI23A66uT7NuWZIt35630j5dpzJsoNg2OHO3GFIK+w
T9GtRoplYwnQTuJM2drfyQzj5YnTMHyo5sdHD55iKLLrYmnPWguUyNqxBaVG
KMTJHdNsUN/BAAtnDhAf+Dw34yJ5ukxGY/1AhctjwIMxyPNg0kw3FAD8FWg3
Cu12M3NslXsbbMrGVRwgzeiBJvtZl5jY/TxHpM+THsrh+hKMzF0OE7WEVNSb
g3n0zJM8IyqYyxiAsL1LDVfWThibDWbSXebbNCx43EgfT4IgAG4FwUnzsC9m
B2LI6NIHjZk/4UQ7WyX3G7ZjblV4iNXVj1Oaww2XXvQKcp9NCdJMoAyimbQ/
+OE45eD5kg3nnG4cFaSVDXb9O7g9X2KJvhZh1cYuqn/y3v4vtcTN6Ld9EMXr
Xfje31n1N586IpyFvqXbOMq9FWsuq22WfUTgrDtZ4W1tCNA3j8yCanoQOvre
IwGZ2Y4RmY4dLHdAqvBn4fgfu9ZF9eC471tg+mVvpunRMJhILY4nxV5gX1jf
mydFJ4uqwU1P4Qcp48/t0ecFWunKCJWJgCUfhkYwWbyk5ilnyf5apHOAXbiA
fWAmAsajkw2OnzBGp5MtnE+KIlP6ebPTvJmWSfow2BHrzyVtOqmwvxVLTsa+
Qk9bNL+9a4WJDkYvNv2QX0OEj6WRF9jdOn28oCG5QUAblx5RIifCiL356ZaY
X3wRfv1NHpaMNMAvhBVmWMsybXtybdGXsOACLCEub8maRMGZLq0MYkBaVKa/
nlJGyyRKsknk0Aid2UmzaroIMGJy2M6ifkZA9W4VywcXtygsKHZnPvvAW8yM
ByTAyJBb3m5KgRf0ktXEWyjyDP/XEDOK1lrxHJJwgbuNCs64Tkq2F7QDmYGp
vimBDq/fdd0JOLv7WZW4IGBa6t8K4cnQe5mlHe+Eohp78vpWBIx1GrGRmSXK
PGbpt9YjkGrgfjCJmCww38KSlYU54YeoiVC6XyFQM32iGVt4BmUTA2xhkhaA
U1DGZnFtPma5m0QL6gkPqfzHwvnt2maMCiQ/84vD0cX7f13bZX/FvRceNM+r
iit5ptzQbI65mpSSqsbjZcqQyPkQxCXu8pjuVtC63yvyW+1gP5ZGhLaGEO7L
zx23vM64VXyADb59qRqJcnfbXiWneYL5BzLoa8MQpHNaJI7vu/EfaJWXmRlK
++zUyLTmJjENhBZPLR0zQGKTDfLD8O+5pkW/hgeG6i6blVcuFxO3ptGR533b
PLXxwwUeNlglmCfW+0wn9+37qBv40CV6RMCXsHFENnZuFi7c+HjroPrLwkg1
OEiOZQn/ZlhvtYzJNjGnv9y/19SeDDnwSmAIAEm8m0uLS1cmejj4+Uuj+tfm
erz9BcpRTiuoVNE7kE1VnMtP22ZTLUuUdQa7IS4cPkkhOuZNyrM/PhUfBk5O
xj5kMrXgTMF5zS8XyyWFaWRWcYoVNLA3hRhuvPc0oRwa8pSKKseJ1cwc9v0R
8D/qvBQEM1FzP2tx4J393WCdAgcCw0Uuh9xji9h24sl7+gZk9FAHDDOFo5hk
MIMCm85rQOM0s2PgEbiZFWINQBbtzo7SKowoufeaL592PVHY9S5gk4R7w9gZ
klHT6QAuMhPU/GHcvrtdTXrlXpYeRR2qNqSApNeS1Fm7/BJN86re53kGn088
wK9yM5TQ7oGVreok3u11uaXqtWsnrCi8XQ3qAg/ilhLwuApqRKEHHK2c0wwB
6eekdW2rGfrk+kt/wsfrqBpb7zkonTrg/wkUddkZjK/DXnIcDGp7gtec1luL
A2gzHCNH2mPNaIOkaTrjCVpyV+aksYggn3kD692bj3RrsbuX4gM4JzStqvBO
yhsqN43rHOmdTOR/FHvyZZTshEboqdf/e6fmoxSubBHXT6sliuZOGDmiZapG
UDmHK7YL06wKIm5PMSkUMNhsIgwKWGTxvKDnuxGMZWpD+rx4waEQR8ICIBYM
yl8gC3bjjZ8W0xbR2XyolxpjnWtfOfia4ODZHUJyz1zxAhW4VsQOCDrlhkNN
peYfp+ZT1upp1VYb0FAA1pO6ihWkWQTQMf7rfz3SXUtYLYX+cabO9LRrXXkQ
OFuVEVU2rqsBkDNhw8QaNh2tHYuJ/rzLtvifm//FABQyYSQMdtvHLNPuJTAu
UBDN8yRqYsNMhz9UCO88FdBJjcFwxjhmwAQOWY1XJMhjqMLYnz9hXKa8tsry
2cW7pp236Jkbk5+TVDvuYD1IdhlcV+xbFj4wJ5TNL5KW/knrg/yWCldGeEcX
TrHTGjPn7SAlENEr6t1Y50iO/deaTYNDtoXQkphd0MKtvKiE5jz3XO9quDcK
OreQBBHqUm7HljrAiDTMhOF2ImUsOmEcbjlopeqK+84bcTw0Nw/3RSTmCx10
yLccybovJh41AicH4pnskpbarh2GVqSpivfQRt7RzmPwx4cMm29SRLN+yhOM
XYd55v4+eFyaU+deAMz/VV35SX0KHBlIs3ofF5C3yRoKPeWSYe8ToOh0+LvZ
TOSsffTZ/TzpXBEmZ74hbxjN/UqlG0PJkR3UjOoj42L8EFvBnngzA7hVPEvb
IZT0kMcGkQkOZVqXSayWASQJEEnPtSVtUxJw8WKsSJwAY3gyeiibSYu2+8f7
yew7DUCxWhlEuLv9Idi4EywOnfv5iQi8KFt3qXZwq+J85w5kksXHpIBAp/HX
/hWXy1KrVBGNCg+bFqk2BDUc9vOd7iQWPP18d0KjoViVCjEt0NiLiAzN63Kn
M0cRGMUoJxTM1AeXlkVMVW7/9hQyZtHxj0gTVOQsRFQBtA4BQdbxgZf3/9Bu
lMElXD08kSjVsZGsE9fXYDpjZZ6WvdaDz05z2rF5ydz/EmkFbl2NKFOFNqg3
YF2+rkDGay+nXGQ9r78604VB8S0RCHdJC8U/bKgAIHLQUWitWZmTb9Jl96yu
npmBhL7+MflQKtO4dHNJ3i3py57uv+Pnp8rW9hIXQ+oAqajgkeixiVkMu0U2
Ay/U5SZk/k7xnsaJEuX4w0FNYyTazYlnZO3NquGKfqcR+AwTEExUKQ21lma2
woaYExA6VLRGDoXGhpsKC+WqR5qi6o9RtOlMoC3RPGySkBh0S+XdbmdmfnUu
Kky9nADaY1tJDiJe1QlFjxTVlWW+lJuNePWwfywy9vdFF8wcnMXWt4rOA/XN
/DJgvUh9WMsIb4YtIrcbKBBmf8hOpRxUXX5m9XXjQE1DqyXoNTGbUUP8fcM6
wqEx72pckQmYFtWyEU7IkmF+FbQvUkCcD5mfLnb781tZemvbe0KyRVPkeDaw
8ehQ1rZAJxX7qyHSv4/c5UKA7nARykWRPLnB32xfmtSu7VryhbDaaLsFlAFn
AGxl57Gbe6SnIUWmIMT79mnE/E10syWNviW3Qq6JvPcS4EjlqhkmDXkVx+wJ
H6LNF3Ylbjxe4PmrPDtqhvGACYivWZzNMHoezGkcYVi9wycvLW11zLJHxTnl
XCtBS0XO1fVyzf9UfOZc7zxaz5zTXSpelyfGaLFKH5eMpmajrC2FLSaI9zve
4pcqA6HoltLLCCO5YQcmAlRuj6HO4H8SspweaJl/Ym7Lnvmv18GGXTRKMTA4
X75U2emo3s87vzZqVxUUMhvbN7+gQKeDKwu3hdcXt+zvgBToIUx7Ud4Zj5CL
/KwSBxrLxUZFM1m8wzogOTNKTQsqmJNJJoeVyH+gqynqLJWE8062KYD+C5jT
Atp88eMVA38HPL5u1SOW9ORMzTnZ7wG8W/X9omUysz5WzBLw6PA5+FVyHjIf
jnH6ch28e/f6gxQ+0EEhtUkE/724i3P5SUsEU3WvClb24cWKOWA5PQ9ryPMd
ackaw0662D1qkq3lCtV0MPKW/3xfkmP6kLfj2UtqpYkzZc7zTbEv6cms17Yt
o7oiwpraPMdnx+iGaq3nEWeReRWGDsnrwvmj5fUPz5hK2AWBIT1cWvER+mYu
cAHdoe3eN1KgXyxvNfGsTc1JuH1Ae/I6VM6cx1R3jvcY67xAAxZdcZ9lg7dV
0SF0sbagJywP/TglVPb6hHneNadQXUTcXYBAul/Z6qIzT56YCHpGkF5OiqXK
Fw1jeLkorxv+YyQjBOeZTxeShTH4n3JiV/vYZWBwvtMyKCc+CN/quOIoR0n5
E5/B7XnBnskgIdhAcjLKJQmimftEvc3oKdUFpoMAOPnYZzWhcthgeb/UE610
NBlo3EvqXQdwGQYn3NEiC2TFR/o91IQCtqUUGfdYsDGimKiAP2zBJClPczGf
MnTX9K4kkXACfnz41AVBaveJKORPARpjgOWbwt/CojQv2CyiIOt9qnO0sMjL
JTR9zJfpsOzsRRMiIqXcjcsFrnFMkBJh7o42ovgJP0bWPdwu7k3tiFqt/UF5
5Wm2K4IcQbgPcnEjj3aRGocoFmvBlcEjYp/Sea55GbBbFGO5GrVk9JNjBEKG
6eEI3cDO2s8N4+p2BhoaEy4aLhl1rINYcqQFSuo9Dt7Hn/aXL0OUGDwI0KwR
jB6CAZ1nmk0J/Y5X/jfSybZrE/X56am1W78Pxf+fSXAPjUzoJNca8yxolsJV
AHXL2YLMlSRrHOAQD+Qb1L/Lyo4NqXbWOKNOc1sBloXLQQ2Ityy5NZSiOiH1
BuDW0s0hHb2tA88vymGRspFYevqdZow63/mWdzJ8fiLKqnnHZX7BycYS8210
Mpk8sc9EQd4OY1O9Hf9cMcwKmg+H+ZLnQiykUzWwBBnqSbmdXPmyU0sj7G8S
Zwd04Jhzff/WjQB6EYsaDMWLb02MTLkcP1Y6aFoHCFwcd0gb1T1VJ4RNZsFZ
ukG/EVw124OgHzSMdWem/1K1o0m/EbUPXjcFb1i741i7PEO0Gm4vF8HV6zJz
Ln8Lb7YZgrMJKMcPsfYq5BGa8NdGd+AKrZAbHhn52oax0JDxGBVYydAq+Vnz
HLWn9zxtNDLLkVcuuR6UvNF5zPAATXBn5/ZGfrEtfK/fs5oDIL99eRK8ApDz
t+/y33atfNKxK/XvUuMuPepdk38CaU46yBQprxA8SRV0jRDieHLmxkszsDWr
RD2MVq9BKWwGazGi8AqYvy/A4DRts0KyVfZ54RLVl+wcWsFz3vvaiCKf+YgF
DaERUnJs57v52JKeEMitT5FiuXoGkqmCYB1QmHsjOVnFtghZRb/AJUkDqIVy
1e8Rhg1SXQE+o5wQGVgXs1hCjB54qpE8VV4F5uJxDQ9MQY4xMarN8z6biSF7
L6C5NYkrLDhoQpTgsbL5dxFuzzUsQzdt8aE6q/bhTvcMxJnn8RaYwP0WQSpw
qB5KtwBdUJG/F97TtevlCxGHjvQRBZMTwibYxc3+901OPYOLbjDQsvV8kPKh
CQWUh3/vzB99xCx3zZH+/C/cwx3lOz/brgBMIdPjFYALcZxxTcW/V8XfA3Df
ZS8XH9e+h4afwEqMgneMbOJloGB8KmCgL64COeo9fpyrkl0jEEL5i1MuHmMt
f7BKNf6E4Q5uZdjh+B/qxVCPlyvDjtkEX6NF+ouYInfwTOXoXpz8gUdpCiEi
2BHEiBD3FovRcI98XeqNpNLiUQ9Qr9J3Huy+S+hoNeQsZ1bdyJThRfVMAuCJ
GZYRvw5I72KKzqAi2W5SaGnGnuTRBk7gVjS98c1IurtWl6B5DVQAxD+nZKjN
B0s525LkRv611S1IALqDxHpP2Kmz3pg+Qnzvd5eD4GQ502Lkd+KyWi9WPYH7
NwzKkMNmEHi9VjL1cxjmheqgGnmJO+82zPEf5C4GXtjZeQ8eNutPxxsT2rly
PwtdWUaPf8RgQ1fo81Ic0Og5PltrLCvdJKAKwLODpER7EAWBikclFcxtqOJv
vjQMaCivyylaCDLKL1icGHB2foel95ggYZR+M9mcHlBxSI4kil1CvQ8j+XU+
cthqP7xy1JKlbop2ETJjo8x4E/j1gvkXJzjx52xlW8kbR4HujdIJPKHAgkZ3
UJS4StyWpv4VEYRwqQ53jGUgjcbcO1eFzZ5Kd6fA+15RO/rSGMzuYzYGiCwT
jWGpjGLosC6Ic85Seire9Gp3DCDT1CTB1vWDUtKgZVsv1qySyGlkHAv8M1pr
muZixjiJgPqzCD4R2KDmIPrjQE1H8wlAGOcWjYAjWz2DcSaBh+JDSUn+uLNO
EzqmZLsG/a3FqCDYpoKN9pAty1s91TQ4ylmHyeL6i2G4B+c0bkWb1RNeprIh
Ze0VLYOqHjXXXjaijCm9QVZo9K/Vs8tTnKv8445pZg9EgeA6/5eqGlykt2nV
bTpOgO+jX4Xvh9T4qF9+W4Vh/sZ9jQa9Q3XhcZOhJuVW7AKDMa+avQqStUv5
EEMx4x3ad/Hc+Sy6iNU9amx3d9/hLp/r0uD91l6lUCIC5wKGDBG4e5vZ3G6b
HPmr85vnyxyL2i6/cidbsdkhctHReOVwb/34FbYu4hjlhSNJaHam5RhpZ7H/
nGcOwXijGNwZG67ivRH1wkjB1HML4DIVmZEbx6iBcuJRtsBXIjSPvo9Hw6X+
nsl1qxiOm1p3Gk7doyDoeNnjet0JiqDR2AqZlawPgx25bt3yPWzE4M9IbtuM
ugTSDdkiHe1akAxXhUkoUwyot/0L03cIx5oXp+2wHsGijz4e9FdiFC8Useua
ajtE85XkZY8QLqPuhc9uHPDYu58zfmqNfOz5EEUKnv1Yl2XODy2h0cJF9WGp
dk9rkV78E5iHaBg8zKQp8kcXBxtxMkhalXgytwuxzrw4O/D7qKbLU62raF6P
d1I1b5j8sMhHbDrqzfobjGUd+gt77pfdXtNYQhh0p8lXwK8/J9UikVqlI7mO
02h1mNgpupbcdOR68Bgi0LnWrVmmA/ejlF5EnoDVUE+nUpsWLSNxMEbMPFtD
XxkYgXBqEsjkADGRcofdXL001uim/YskWQjUaD7RVsZl3OxinBxd8iPqsRMP
UV1NcNFr+UWOxK7AG6UYtGe4NGvOF7DuSr1i6ldBgcjFHlHmcprfMDI5TDAV
4lhyb7CrsdVJx0G1rG1pGu2EMzeDKKzEKC2HbjGTfYgsAx8+0Ro6hLZYly+h
5j7+wS2kVF+3T2JzQZboPcugaC+wu4SRWeqofl4Nlf9V5eZnRK0gKMShNhYU
lWC1zHANNNF2x+QnU0ldHnMtFDNi9idqSM7zObvCVQwhDRVf2gtFgROCmrrZ
b86B4tHOp7Vbp9YoYov1eaN3Dk7ud/erZppzXVSjQ69QIT0LQ+Re7QlcDhC4
kZ5gNnnocCxp15EN8pcS1Z078vxT/dhzaOZlivUp3aifV7mGUY4nXHtpCrdT
4g7ufNZ68zv0j6LaCOP7CBMty62KgoO0TjXNP1hvZWbPVCjtQcQUXUdD1E/u
Eg1DtJiTv8kDyOc3mnza+VkTTho2U4jbM9cy85Y+7Sb0EKrZG8Oc3rU+ZmJB
NUY/T4ZdFhnV5L14hoGx/ojFnvxGgyydPlvWUdZ0nM/4XEllE0Vk9LMSdQiH
ITu1SkI2V4GOvj82eBxCqEva0D7jA1qcZixpDgxK7+5wTXnshqkFcKvbuh3g
5Tjxry6ZN86Bd17x2FiWUSqMBylIhqsF3EE+utnCykZD1B0h/nWPNaJYMQD2
GPctFBTPZV1EJ5S0Rx8CwNehwJFyH9FjE4PxUQvMGroxY2wgABIUdfSf+LpH
/3ijIdVp2QLu0hbWx9WlwQgmkaECJhmKukYjcoCeRGeV7NF0ukbiaY4Dljxi
gdUhHtE41gTPhlhq/PLNVShvcD8e+On+izpdgxnJLWV9V7ZVRPKoKV6caq9H
4CwH2190hfVHh1Plo2vwZb4TqILFpK7E0ay0ok5Q9IVplynVl+p3VIFHWsAF
BTOUCM3o+BDAX6igpAdJ3Wrp1eJJ60GvNLU6HJiHPKi16TET81ZqrisPy5W9
AN6scb74LgbMW+ds3tTVKU6dhD3cMWUeuszNQ4BeivIfFUEKW4wTFfe7+eDa
XG26HuXJEJsrvaFT7cuqfNoUqECmQZHb5HYxIvV9A/px846CXd7XLhpKa/lE
k0ghNkIqC8st9d30Fj8s5M8b9GWyKDNSo06xmiOCEf5CKgHckpQn8gFBVtFg
bQ7fmDYG6Fd5VmplK49wlvXikNP5nhjQPmEtoZP6dObo7jbfTJPJxxUYdpFr
uDYu/3PcN77SWZ/IO7SEY3F54ItEN+timu6uxNanjYw3vlM24HT7eVFJ6a/O
KiGq04FbmwKbWpzoPCiPItI6OJ9XPQeJ00RB6hdN/91xJ38fWTKZesMCjHGe
jDdBV9XFXiitdiDDLDx7eEEJaDMigq7Nzxu5Fkm50rZAIp/5QMXylJ3PHjGW
eUfL3Kj7BuJwoIlzVjbR2rUppXuek8ftkwcUP57xzYMUa9VTDjhv3j5ggak0
YsWGiPCunYreVfI/jyChbCMFGFDBnQZgORDQZHzbHY187qYJcqcWCiPsn/pY
aydR5T8B1+FvxxHxMp77Z7bxCf6ETdCFeFbBjANxL6Q4iQX38x6iYZr1N9Lu
64Ept+bukpvFAu0YTFah0dV0skyqBKmXi9b00iICbuL7rKIdjvaEuSvY1758
GXrjvwQafd8yscY7M80bgx32MDBivFEZqU2CQUWDzK20VXOWrzqkdLyGu6/u
6cjarnmiqDiG4hzJ9AUggBQ74EeB5PQ0qIziRHcE4tkdfJT5RXb3O1BbNef2
OlwvdAsBiwVSx53ju5dt0zbFEdLXTiLr2KWdHN2PmY/9HVnMXWEWfPOt2BGT
sM0ExSLU+08MqN0LNM+lrTU+HTcnjLUDpzMH2A5AEsSEr2h5hjiLP05bYGk4
7V/7gtKRbs+yCC9XRX660HOHnTcaA335FdeJpjrvhDOGgsf9oiGz1OPWOUPz
kPdjJnLOthS9L4I8jQg0f3cS4EbL9Kp6IeFkVv35SCV0StI03GC0gzHhZpqA
NGjTKYXzAXti2LlCvT1FHBKWbQnEGXDLVAwaClMvD67rqen0WmwktLD0SFYE
bJlDWd0fGnQ/t7rmNV0aGWHVmPhFUwN3Byt/Xh+o6gnEOytZDX7WQbsPHFp0
f80jccsDHJPlKNAycPrUwDh4ZJ2w0sQoWtXkNqAFknn08YEHs2gMjMcOOkh5
2QH0pLUehrYM9QVdTcegUEXujYMJZ9Z/v1PV632yzqA4RGFfdAyMTe53iC4T
Zid7lIoQhp7megg02MmQgfaSZkluoWujnYxBvNLJaiQ4mYO7dZxlus/SzYmr
0YjGIw+rpew4CF+TofS+8Ghg9RPb0EnTlYKOIZQGtEAPTOBlirp6vRcO8hB2
z+HOEZeQenBH/w1GZ3Emx2t2fs6z23Xr8Pyxz/WIPQmw9OlADreBAnOL0MA+
4nIJ2BUqM4RtU+pkcPGO7bC27PGNooz9mK76WZYy/80SXswDK4NPuT1YJ28C
aLDVpt7dax92wEiS5/9gLyACTxnUBcGb8ro2ME2lbm/s8HuKxP+q9Ee6nKfO
c3sml1h7HlLsJkdvYgD8zFDV1YfYKozB8EXwZ39zfZB7XjqV08oTFtVXNdNf
hJGUQUg/NQV3Fx3ho2wyvGIQESRxZvPdpqh5T+qKaP+ivp0cUCbNVa/JpKZp
kSWOABG0LvJc22nyZjA/lOiOtw2i4zwZ+5iCNIJPmi89rMsUKBlz5EtjlV54
5aCkFRBccsYQ4oybSdJNh6m4Nt3GfzNR66tNW4ZK7Sekqe9OoLX73Tn+OZmS
1HWpTofyAw/q70beoImkQDRnC1ldLIr4N3JRbNvyQBt2AedTE4BL0SLzZDn7
pEO7ez65Z6+3ZixiN9Xz5S/tt0Z4jdu1egHNCaXuPbAS3cKW5pQEuo6BxESl
vx6JVGKSOFnFRlg1ERlqjzjNrg1TEx+6AiS0JkbgrEG7TsXrFDY+5/SBjzcW
L1nu5OrPnDi+YfqFWU6mE6osUpYhLr/XgSw+SzDHXRtpgjppK6J+OSyCsB3L
+sqWNZKrIuOL2ZHka60cbj1Ml7Bj3Ppq6h7eJrX3MJOusKSQsr6ZHWdMnWm6
/FdgQGTAn5p6BMcVH7jneQAafXek9m+5wHMDh0xrM/kf+QFuHa53gxgHNZOO
sgFIEJseHa18nmTGPi+fFWBzBu2siT1s7aU/AwdcnnZmh3st8UDFikudZB24
0SuHmTwm3156e82veAxOnvYHzV+jGUGNug8ELfYUNcUI72eppH/t5d3zx/c/
BH6Xo46Zzbnhd5nQgxrVSBmQ7C1f6ooY5pTMZMdhCuToULWLywXTMfA/sEwV
e0kHjXCDUxfqncY+Wbls38yUll4ugJNc2gt+6cUu0N7SloGxU0Onzs1+9jG2
ejyUhZf06rYYZSx3DRiL/SJ9++VUWSY/lBzjZ6jbo+42p7b3yvvoBctoDrXr
aC0IDxOngbNro/ZsnO2Dvhm9NHtW42fohvQP+aDv92GS9EaYNHKAj8EoTUEb
wWQP6Ayh5ZGpMMC1EdrNISVUvyn7sZdkg7pUgYDeh7vGN0bpsLNZuhqabupO
ADUFTdSwRFM11jjaKPPbveKZnwkkSkYVM825p7/eB3XyYRYg9qGcLelKnYef
CxvRGgbgkPpvWipDbgQ5AXd+TaAI1NXGsULoMlqelHvCi8Jz/MnQafMPq2Z9
ELkCJAI9ySKDBMpDV9DBoVuxiO34TJRbbF/zLcB2hz5q96fRJ8jrH8HlgsLa
8Zj1HnN6aPqHhIAyovc48HvEu9ctFAZG+R9S1y86MDXm12QbT1/hVixhbBpa
y3VWm9thOz0INiPpmYVw1gdQMKxnHoJQD3TjoqgOrciV9WkxNui3R2yb2PZz
EZc7yPp5eFL36iVvcEjevJc5Xme8N1+dyCTc0RW8u7oLgWf2rPtX/is/scZC
pOdbWJuzoaBFnc3adRH+74ByjljZ1Lg3Mk0vOfiKMUAethwjKcSm5aMMJrKh
jwnFji7q/SZM9yuqeZq+eUOKA/w+cIbkpr6r3pbVqhoWEcpLHy272Lk0aUgS
5PMc6u3qlmj40lD7aTx9z9FLL1nJks5BHPVbVFZyOj0EEW0ikVbJ/MGmTqj9
+SopOoI8aQ7sIZCcabN6pd2wKrUumRJmK31+1oVprk+bLX3bJKj3TFEcXo3u
EmUsx9uGK2+4FdYGCDERU4If6jKmQt6TiWOWNDfvnh67UwWPIAtuN96HFArP
m53EUVodY/SjXluOhwPKQsk0CQv9q1we/61B5QBNb1crGyq0Y4a4myRxwiKx
djV4Zj7dfc9fCoEKDNVJAYHk/dIEojAhQ2v0gKABeheZlofkvns+v/UGU54B
s8LLq1tkQ/PdtKeDHMAHGQfbbrKF4zRtuP7iwoXWphIUwfYBSiU6DvEORRc3
8F255Wcsasulvbml9uq7ve4IoPFszQdOBmRDmpJPWQgfV7FNgfIUc/BzyWfx
VXW5wEmJuCyxmjkOPaEF2viFMF+RVPKVU3AVg0N71XhO+tPG0tyrsQEQiSMs
hPra+BCOJrCxv2Nt+hDhDICoUkQWzrIjtYaYMfyMswva82XB6M9BX7mLIrkj
Uk7C3HpQfS3bdWuvX44iNKQLJVytV6QlM4cKnKyC1dIkWvnZwzCXflqU35V9
NdlOUxJHtjRXTXRLxBNHEG/0wWuSZ8/dkajNqJYkak3RXnB45bbd0gzQRWcK
RjrXodUaRrKSh4XpJ9hX+gIzB6+kOD77lXpIg8ZwsS3E4hTizlISAzGdVjyJ
vgbRODBfAzgAdRzZwodCEsSEnH8Lx1mY4TLUVducDDKwCamuTxfQr6DP7K1R
cQq6Mm90GoJbBSDawhrs+JXQxM5o10IG9ifNhLV+FOj4Iral3ovKGZIF9opp
EUulIyLTJhyCNKkejAZXtcGhQ6VrHCA4ldHU4c1UTdYfOg4TfZGJMjbNlqa2
j+TmOAw6O7RjgkaIrePPLUOTrJ9buBNuPab3/7tlLyuX4Cax0RUk5kU9i0Db
QJ5nhqWPjducS0AaaQ6oMrgW0zPlED5tUtKNG3QdX2le4CcEVYQdTEegx7zI
w7pdY7Ge75oQO50oMKqXPw3mMpX9wdjHbSvOoZCvERo5qJWiaz6eJ7ZHkY2w
uhPaeBqGcJDEvPJ09NfGD2qIT+gE8jEK2JHGM/cbDyGnmUCBC10DzoYPI02C
+T/mSCoqEH5j9R6ArkASKbdHqRjn9HBkMl8DEat4eSkti7JHoqWoSuqL/KU+
mlziFGDCP852X38D9kAoAuNi9UPUxlLqmtvyVPkayvnVspXPiQ8vW64WFUdz
kHpGpnfzVp74YQunepNJ39n0tHa17DZE77U97S28YqpFe+4Z0CHThvtu+/WA
gerOxK2Yx3e4GXV7usiNRqPUsuHf1F9jabppU0DDODn33DA+F4/U5WbCeugh
mI37wlNMf0qaCOonbjInOQ9wG3GxgVR60NkvsPZWDuH/WtOiP+S2SFq2slcm
YeH/t4nf8B3t6qh5Mnup+Qwnsh+c5JqE92JEu2X8ECEBT1Q7AFCpWf0KW0S4
eIDArxQ4/4v8EoZvsRZwCd7NXdBq5o6O+gJPuntTaeNmM4Q85wz5TipZxAtx
wiGjCIXuGoDRIFQZF/MkemFhi5bg7Z2eCyKaGIP9AkMaSSXyR8BcUl2djjSH
Y/lmjSSM6fxthxm+fWAUtpYuPzgPxXh9B7sCRJBuqwR9uPo0gD4JZ8Gls+hL
8mc5I0h3FPZp0WvwLvVsBo0MdktSkp1J1ZkxZofYQ7MiAC1+61dN1Lr0dL7W
DYV3N7NduHsBY4XyW0s8Ih9VfhY91MTvlYkFIHQqP5BfD7kyxg7svmulZhVj
mMc0gDJlJ+P2dDyZkf4bSFXOClzTdnrqDwXUo4Z5QleDucFW0QjIyUmWIxQt
RbGZskfoUi1suRPyOEtgcndGatgZibA9BmK//vANxXV2ch9O/VREWynVQPxU
i58VcHGefB5BgFMXUJwFgkO3Gcv+wsNEl1vJIpYTRgNvC4PAaceq2Kb+6PnW
WRy5TU5/UNqOZZsyrKk1wz0XnqB6h9EqIM0JoQMXOVzIRfoIpwyWQlRCiEBg
eIskStGzK9Ap7nzTnVCAI/9kP0cx6veAU0VWJXS19twloTLYJBkB8ClGl3jE
DVj4b9NuL16lOVPJLOVxQSlONsEBPOONxo/Q4VuCHBVVRLYB9wyvltu2i0NN
hIxQ0UaqDVcjC3yZVcii7flfpN9YXjJlCjNSBOgSs4aLuwko3rO3qFuM9S3q
5QRGUahs8kLqsDLx/NlL91sQmSf8w/pTtersTxcSuaZYqz1W7+L3vplmgm3/
y2zozpHoH50tKouSWaPQrXSi2CctRm6vCJpnaJB7u4eoG8qIzY5T4Axh0RFm
CE14833jKSFrki6bsu8/eNvconRg2n79/Ao1OFSoCi2jBjK6QI+zXhu0TxTO
Ij9w3cQKr5wF28trNffl81madovESAHzi/55cLWccRbdqHNlxzw/Qft8Z8o6
vm8EgFW09k14oCdr1VQI3/NMV3xH7c6AWWjOATglAvoBQsksEIhGsLBvwpVA
kylNkcoFlntBu/aJ6ieoyKCTnzP9CwSB2kxmGM/Mnge5deoD6/qpsuva/CmP
kzU7k3A5iHnV0CSu4JCQ5UmeQyzKzjOOMDTDA4cf7RulAjX4LRkE7/O6B9+1
CdkARiYz9mPKCuwZ9n/aGfMJGRUMXN6Om7eaiF46u1MCMI4yOsv24/MADY1O
eFj+idcUuiEuoIFCXYDZh4bGQp7JWXy+fYkM/LBXHIEqDrd3AfMXaICFz4FS
nfmREovaEVoeu/uretlliD0Tx/0YUqgjsE1Se7z1syqmQ10Cx5guBM8i0M6/
Ldn+exZtMrYlM4m+rS3FFMU7ssrl+CYiW55iT4/s6NdLqx0gSp1r4mEic2cc
7a0+Do56rrKhYrJzfSY8cXT07P6R+l56763IdjWupsqvrQ0hioH5TsTNm5Y1
2TKKbHaj0cbBMcyuIM4tgXtCONMBun/T73If48SmwienJwNBH6i7Yl3IJUEE
jNM19d7xhAfDLsZ0jernl5d6vfLdFOUHJE62CJ3YRX+sNV1wpwMeZstc/YlQ
pcCc2LRhM6yxIslpIowPiKgwxininvUJu+hBGYGhJ2ckw/FmJUfEo50IIToe
UBqo7fcaL03t/baLLPYRnd8bFfu1gWWLt7kazWA+QZiCU6cCn/fUaFtv5gHk
DKdtqStF7u0meyWh5biLlqxB9vgo9YJUTCgZBH9raLOnRKqbC4uBsvcYHLS3
Nc0o29AF7rxLK1G9bmDVBOb7Co+6JuDxsR4emrSrBpQ9Vq1OZ7AuLhMThN8J
OzG7SNJSQ4PzqKvCVWptg9YxhKewr9jLURCN7OYmIm7uXyN5YuEiu+fGYYfM
a0dOni5Xipil/ATaCSunQxKLbL3Rc+cgeT2yLBZJSLx8IPgeCSmZPfC83STj
cQpbwPstA3EhWBBxHT6IqVtX/JRBh/1qo8W2hco8V08ezJhdubdROMmfXLR9
i9HUYpOsXUF3cttwfCUJiBABuVBsuvfulUtA8QrBepP3yLjOkxs9D9rbCuMX
KEfqzMP2j8hy8uXrwSSIUsKeeSCaook0GrgIB9dQH5ZwhX0RnbvCmDyUpmCy
iWCEFS7olrF2bTZRceO9fB1lbFlKTbRG/Hqz3R5vKC1hr0nV5iZ6Ke/4nt2E
X0gtvlV5SgfF9NF6UNdOU68ePJ299Qy8SQV5xVed6rn4guvvtiPPrOzNfanO
HpLkoLRBE5CB/VwJegM0OOS0pS5vnDVdWy6++EyOghpSH3bT63lVzbdKet36
Xl5vFXc1fxUr8SyQSuF5MablaFDXbldkyTpBkKhHzJ5PbVIItEtuXYZWaTlf
n+uHpjwQIIbVyeFRroVbUQflHwH58FSaJ/HnX2nqCVFvLgLlteZ8a39RgaTp
xQqGvbSLQzKntY/WsqnoxmK/XwwUa8M3xtqUnYqxnK1cXsNgI49etlwx3ztO
kwHbd8egH34uxvm4RumgqIgRkw/mBP9e7bOknBcgt5rC3AMhTnRq0asRjrbo
1eGXw0Fttzo/piR/9PxWaEgYMD2QlOcvwnFDoXFw128osrhShxw+Jh8KcpPL
XmHzClFes6CfRiEY/XaBtclamR3mALdRgX3ia+dzytLB2MKlHdfjieEEkudB
yEfgh+cxrD83XVvwQsIqVHPGg7hqV5V4l12NyZ1Q/haVRtBOxj7whAcM/WBe
oPAcUdi2A458uQQQL66ZBH48OD4ZpWSIyxnq4N7BI+22qdyYSmnC+0jopBau
7ZeOCuqGGKFC1aQiivAdrtVgja7asUCSu2QLVVrWzUJeLYoe1sG1CxLGxGIr
jpcnLBvseqQZh0A+dpevoKsKpKMGrzETVBcTvFoLAAKiG4mB05JU+uJDJf2N
0qe7yzmpu0TDnSKN1eQTdHqJCCc1unLVWLoxgmUuuILvLp8oK9O3Y1w/Qrok
fdxmqKWpvIqcSi13lSyF0gNYvYIjzf1rL85eMyUvdW8Mgr90E9D0Q/LWziuM
/qlyYBh1sCv6sDPRo7e1G03wo3BULuDX+ZLsAvuaeYPea89t2Pm44ZA9LxSz
hJNzqyhD0A8ZKZJBVCwo99IZ6WqaKyygaQKxcCV4GoqW5PiRwoB6aKTuBrdE
84ewhJurfuRurZqUg5VuYx4dA8Pys5wtwsa4i/doo1gmXjvivSfasf+gGEEi
bqqAZFUwicJI5g8nyvKrr8BsdeV/UZ54FmQSpeC7mIHwuAPlqtdW7ce5OuuZ
D9sgWExevj7Bq2Ig1jJK3IRfVFhg6tLQuUuejoQ/xKDU8Eiut/gSGrc//NvB
q55m4WVYWlPAcEL4nzRiPW8O3XVbokIgnssSoCRBifOTv0wPO5sVE4/YuhxA
coHMenOj2Lac3Wimdy7Ov+rQON2Y9jK+9AMLHYKIL7T12Xn+lct+6+bqx+JN
iaQn6byxHLQ0LMARr8FNCibrEXyZDpv2MWRjN/JhpxwNHTJK0xVAtuyYrjTz
hQN5zbh4e9GGDvmV/jDzCtN3XAhmg2whebsKRppwWAoJNk4zddAAKZV1Wq8h
BZhMjdejHeVcd+fYCz8IT2+ffZzq9dXs8PP03XEEGPaREtodMLWI9pFMuVex
bZOUFYVVAYEaG55mN0b5Dq6XckM/gwaUItctUHb+R1G2zDLtY4fb2OYCb6Z+
MfmiyPGcbn7VPd+oOGHxCL1/jEUEBOx2/Reph60HkykjdkwSpo8HNJcvD+kl
cnhzyJBwLc+FJr0/4/SsK8ckwS1bddx/aad5OAeamSv5jiC3ERhJsEYp85Lk
tzJKPmIteVhdi+h9Ke0393tMBUAGiqc1wR+FKJAlAAJlhbzq38G0E5UonWCD
OQDMTIAShbH1u4aJYDDKstc+dQIcDz/R/n8leKeye6Oy8LT4+mmnck6Kn39D
Pr5Hw0ijgO6WKtLLXGg6mgv2/Ai929bLq5iumMT9bRDS+UoOKSq4oyZTpAjh
MKV8VgMAu24vJylprGzf8fM1Corr0aBTVochuNDjPS12BA9FajVIOhkjMn4M
UXwYG91lwVoGEVBd41s/MFAE00JpvClV7k3rJc6I2xEOLf4WZleo8YvOA/7l
KjyMtkx1isnHnMqC2MPioqSIAZKNJb6hwSzhpJF22OW6ulhq/WxlaIglFI8p
9k4Glsrui5Ss+r6cr5cOcby7kXXWKip9RlXul7LaE+vswk17JTaU1wKeHq0B
SealmKoplunxUSHnXzDIn1CZhMmcSGpbA+/4psH0nKGCSgdCS088M4s3Pq9v
jVggScJtB97UJwZgBYDjqBbT3mmwLM/c1EbVDHQYCmMNX2NMq1h6rLeWe+zd
TI7Ln9Kdi6Ruf8HMlTAUSeyoZUex57HrrmS52zyw5oaUQ9iAvEGxLL3TEZ0F
LcaATkg76dOcBbYL5cy0QXA+VLE2fzwQSchQO5P9oCvM5jsbyQhFOUupq7Uf
uKQRiAP+La+aEFJVpwfI8zG6OG7qywr7oTr0k4t5JhmqQW3yrpSQ+Dp5tajz
HfHvE14ulSKatkkeC9k0MLYmPQdM42JWT6G8NdG+ORm/yRVmuBbkyY5WNgYU
eWV6Zdi5HcI5sQgYVFNg5KVWMDmejf3qPsqC0cK5o1ttJndVFBtlolUYC8G1
sNO8fiFuYn2FGiL4j4E3AO82js1YAxjCVY3FyR/7hRe4cmiB6zdgEzLSJZWW
Dms7P0gPZ30TJsJBgIdX+oWhVy6UChfbqhnKVCm10SshsLUi38SUfhxxv1Is
bHQ0MLeqOVfu5TiRuNShhuDugiEmFE9VCeYtGtC6/iZVQds1vDoI+KgheQTa
1cIKa/MpTxUEmoid74fYZAkUKswjaF/sBT8kTSjNCwehVNb/WHCdiielPID+
fgp38lRHMEr+A3NrNZNsEQxk8ftQgUv40t/ykq2FNxLT2Dkpr/yoTOkYXlbf
qYRaf4LF9MGfbX0Xbw2clks25vrKS8qMmqNoyvkvUE2kZheN7Yp2MkPiPvOO
IykyTdvFQroi7mNQPW2xOLRJyuyecJ5nr1gv6+UC7Y0II9oosQ8skn79X/fp
mmadKYfGkECKu2A1immZlIFYScBLk8g1Bxhhh2tFfv7pqYOgu6FSldwECBUu
uRvxB0yYw6koFK+2C1jreUdW0Ycc83xWmQ7cwfwda3D/Wp6hR5FEv51in3LT
m8YLUc3UzOfjPBPBkcVV+oDPzdYnq5VbR68laSldRXSwr9gm9t6uOmFR6zzF
mrQ5TMxq6hJlLGjedzp0OF9934ZxnhxUI7qV1v22oW+58pi8ZatAR4biUcmf
5Xdj9wsE209QIEiRnQQqY4a15Sh2EVIHst+I6jL6C6z7r/PZqgXXly2K6j+L
8sgC9CDZVFyTjnH4N0sgkdwjDgXFcDZkFqSVRgZrRU+fIixXwzTic1hMCEkR
K/xPbhcDhtVzIoT8e75fqofIs+4/toTizhMDdsCANL1PhE/BRC3ed/1f/OEc
OaCqVFRXMqZwGCgGIm1NhpJ03KgQ4ANRYpQDN/LjryUpqnrJO4Ywjsc2QQM3
SS3b5MsutOASbWENfa8/zn11O2fzlCZE5wL0HcUmF7a3tV0DBBvGUIztRVJ+
M5rvau55vKUQx4tMuZ6QG1BPr2y3JbaFnZsIFBCWyik5NktUYjmVc/t73OL+
h09mfMzbMfO5AjOFd3gq4QOignOqM8eVkUiYoxJsGzCeXZrNMZrrBOBdA/Do
7xQQNuiym4D0RJBLlLKJ7U1kP2at6bAC3rVkJWA+4FxkR/jaK8cZSOLrkost
+Uy8/GrdiarHPiZuVx1dABCNKhLUTGanXOw+m6hclm9EtsAMEGsfufIb/N5q
suxBt7xW0H4BGQPEKishkwuhzpcz7/5FvMrU3KmB5mgiANsbuLOPNechM495
IBjTrq7b+4bDQxH3MvzaMQuJhMkNaT5nag3VYN7IdXuGOi/2P6Mrn0lDQEmw
h9wV4W1bett8xkM6viIMPvrLi0kFJBFnqp566O4cGkO4O8uzFFvggfm91uG3
jh+BVZQWPR0wsGfCh03Ywusb1R3LHSH2Dj4EiAuT5MMQ6etYa+Xs0Y199j43
3OY6Ym50EVQ4ZYVarx6yNXH/rnaa1jqPeI7ekM2Vo5OUS8U/CXfyQ8ZGpAEu
UeqTpJhmPGlFP3josiEtzI1PdV4edmOOaqFQVHLGwrTBA5vAm7oBtrVJnjPJ
RhT+DEBB9SvUPp0Zm51s0DTj2lMsbhbbAUq3KE4YLJbW8j76TxbUdbKM2s8K
0+w0rKBqkM+FZqiCrd2gi0TafihB1CFO06BSctDE0dxajzKknmaRi31SFAyw
w9jkmdy7p8Z3FDNOIncsxRu+0+UJlaccjdG4YQRuwaK5uKsxsPqNKUsPJsyq
R0CcZP6F1AWecG7SCpfJUmq4Wv5E21GmybE3GVYae3G9eoam5qPGAe4UMcxy
EXGuXoJmmpuqbCteFir8vLsMrn8VR1ymB/M+l846Ba0RKVWrl4ay98WblUul
5dwSbCu9ykMa5Pnr++MqJhgBwkrHcHWCznxckJcDY3hDVnIa7n0kuOpcKT73
RASAyDp2rz3GmUd4Vhq/aPHCRIF28sk7zffHuk0GBVv8Jf6p+9hfjOnsdPX+
2ublyNWPqw/jBWnDlxrwI6wn6rssuCtEKSChZpCSNfm76PPIteKvDmoc2Bwj
uZVI4ZCTWtOldZB93O5ZovX7B7DCceTqGzVATyMsthqLvqXeODVf7IMK9vnu
7a6H689z6IS5Ko8lLDDdLTJXrj6Ca0VD3af6nfEi0pdQLD8xKMwv4fVGwjzc
yvWq71CCS1cDUfnP8xqaOX+knneaIJPOkH9WpaaJTiojizPgZYlT11Gq9PUL
0QLHsmvWNNl6XghEmvGMs2No9OqRhtW4pZ2IoAsWijvR8fFH+hL+cuGF0CpG
AK4VpKYHgMZ4QTobCDCv1DekMcMo5e6ysVe2L09VWpBJMWqrW6orgSIyVp8d
S3Gdqa9xwJXae+fNrnMRpe/c/EPDpryagwZaOc/HQ8acm4/NwDTGjI98OhRw
yGUGqRKEziYBcAuZrLLIJIGhxIFfCS2iFStAYN1rCigGFHW8oRmVtqUuIx9G
l9xiQTbAfiyGD1oFAM7byONeL2xI+t3T/OgHEpGJdgnW7onUvMOOf6zoxMGC
oRwZHvEtC3vCS6nSwaWds/tyzAyNATCLuikXGzWdhKDYsuX0bSoOy5Bkw2/T
xgM7WaKNs9KM40tk1jBdKAOymWezwZz1CgNPrPiOiu5F4EsHL2Hleo4XXE+V
RiGenZMcuB61obpV5PU9PMSiy8LkrjuzP92cvVXQHr4KV7QIq+Vuz4cBglVb
6IHFobs7N/tidKTkYtDn9e9hjNZBaWNIz8J0r9J89yApVanQmSldzHLHQAVY
mG3WA1xNn7rLhZuWJrTLJMshDhXJi+V2mKWmbW1J+1qM3pahAC1G8oAXlvRE
T/81mmQOU+VkxLdOEe4xQcdjdY4jb7Gvmzu/G8x2nzaBJA7a8xy54CRvatnN
sy/YLc1ypa7N23u5FO8IjHMY5KYGEQrT2qXQZItGLcHc/x+lp0FB6yIG+jFL
F+XWabFfsFj/XAnV4fAB3b+pslmiV5zp9qzS4yUARNGQqT+IIx7N6i1Hf2kA
B9VB7p0tZ5ZUMJj2TvPSz7piT4Q/OG6EVMfyxbqsjJTAvFUlqEFcMr8R3oPv
p9fW3+7+/CsTjNGwO8EzK8TgDkoe1vrbz5USau0ZQ57ca+198ywDO5GKjy13
wW5+OlExEAx2GWjnuzRkYAEwz7AZxCwvVJS66fs2cI9KvR21XiwiVaLGnrEK
gq6nDDUbrQ9LjtG/u2Rqdde3GDanXliMx0Jte2UAL7SwlDTOoowd1ePthNeo
tCn40rYOeBHESqW/9R15x8A7prYbsGWo7r4ODITc2N0DnAkkOgeKdI/YPkIj
o4MgDMegqADQMelK/O6JAL0s/zL/K7K46I+NqmivDDyFR2QxNs1+tsqXYbGn
OQFxjFrFhCCh/pLqwh878+UxRLLjKj5WVKj7KziPT2QIF4O3XbhUrpg/Dvoy
Ins2pl3M1WSqQ/LwNSrbhzaxayEIFPB79pR1IibjM3Vqn20GXUbvSFQLDGyK
g+emEKMPTcbvAzsAuIayK0Sek2sPM9J+wspG+bqM7rAvJgBQqHFxLE2W8I8i
SsqSLDrO4qYTvct2ummNmk7xel+o4S37DJZpGH7TrtYLcWvwXQbYVQPNpGg0
UB1usxxAB8F5LEfWcd561hZVktsCCVNQ9azX9wlKt4o0PvB1iYW6rCQ2hVKq
BJiVe36cSmiQr+xK+s48dyEr54NOyLMZU86jJ4w63lajEmFEV5khOpAcLWAQ
filvRFJpvRBbSCBMhL6jngOy2U77bj8dQe1BhbmSMQwQHUDTLXAXxpI5RT2b
pPqTtmmm96nu34ZVgv+dueTiYRmA4rhnRLGvAW1x7z+99yzjs2FqJ766y8Y4
lkZaB6cCyrZm2dZXDy2/EsrcVJIFrOuGj3ZRt2RiPgGgBs/QJDxi/qYE5b2t
Wqb/pfHveoDgFxiwjwhHYfIxf1HURWn+mM76K/w/dcur+Q6qSpvWYQx718mB
6IX/0pt4Ig0FwOoC1Xf3GphgvNzKsEpChNboXjTgtVXv3ts4bHJOMimhMLR3
+O0BBQShex5IFn9OVDsRuq9kLaA2bZ8fyFcPAVLSJC1/p8KZnjxy2jrnOEe7
ZGmxCJnl0S1z91aFnCsWRFviLTWbzbkG83IbrTcy+hWSn2G7AC05pKDTeqjM
8Mt+W/OpX5tvgdWlfeplOpvOWeVRkw8SwQixBlpU9nWx6ZNbRNOsPPUaQ88o
xGRFdGvptwQ5wWH44EOa7Q6AqUsGkWM5LbEJ9HOzc3SuIf455oYeZgAP9I4o
OapElaCH6tf9VdFgPrZ2BqYm/RyYxyMuvY7jkrkVE3F1kvKGItU1lZYNQCyI
3rLRZkBLGnwqgNeX+tlp08Y6Y/hYpAghbr4iprG0uX0LrwNleo751hJUEj9s
XkVmGKuutFQjHsEcBREiISxkARxywzJZGV/O3xMwZsbzcR9sZO+KwovAgdAi
cCRsWbkvC9L8Oax7LnLcDlfy/ypSv6hpSvJG4PcRYAVVIcDaFR4/WfKRhEoK
vRxc2UCxUspA2ibV1Wbem9XvuwgXDOpzSEGpa5q09Hy0Yd61Nhewy/7cksAa
ZC1cE/V+azxxjxYecwZDl1zFt+P+35RniIfWN6iMkVDP/KnYcDg6YhGxb7Ov
Yugb9tbCwpGAAEDF2CY4drX/9d5FQHsUhT42NWXvosGBdsxnDVsCdjqGxqGE
S7iawfYkc1U19l9ZUgMOjvR711XiBjZIfenVY/m+atbRRdGnXr0yogvD7Yjo
Y+taMsJkdSXZZ9Ni43EXcU0EkHcpqMcjfmp2STazQJG/yMhZZEdfphyuOTAu
PkDRhvicxuIT22I0MGz4AfiYvorDh8OLm658Tf5hnuZdg+apQSJFteN0VGWa
oeGHxf8bgXS19bMcrTETHeLWB1GrjUizR1Q59CvOVuDqk6iOIN5vb9Pxumc5
BuThCxGGnC37c4Epc9oD2Q6lwsDrY5O9hzUJlGJBmpHAMcMB10DcGkXNaGUU
Mq81+UQYS4TXukKx+IGX9D/IB7u3OXFDYnZVxxHRsNrjgG1XCNUmhqLsfiFm
TEMdP0elaEo39mxCLK5w/HP+27yHgJaNTC4luf83Ms4CkxG6sVUi2bt41bFF
vMLf/zUoJkVZhP/AR+5dOQCcbFD9pQ1mKMzkNdTZZ00EZfuvABAaMCygTODb
+itUQqY/DHjHGAlj/ZbepamYtLEJTAABBquuq5lmGxRQdzXbZwu9+9Yj17ci
FzS8+l39aUXXpMU9qfpXfgdQB5Q6nbOWSa4dotqxwmrkQJT/jYBV6UET/+jA
msaecudel0R0CUwnyCLvhZf8qhkQV3sNhxL/VX2FU8Geo7jkclHBDT1YEKfI
D/GsJNlveXpbeFktXzFdqDHTZprsQu/6zC7y9WlSnNYbw5h1May212gkboPo
qHus4ZsWB3Cke/l1b0BNDoaALpUOSA8JcvM7hTT9P7y0FaS6IHrd0kxNHKfq
RTqPqOT2XdoKrS1te7rs8CzncIa3mRm/fRUsLeaRB2TQnErb97GRO3p4lanM
NdOVVeADzkJVIOU/iylahjdNBJwkAzg6A6/D/Bj4soIN1mjWzA+OZjh8aW9r
yNrvXmsg485F6C1B1gvWAAGksERD+hbmk0F+OFOvWZx4naexkB+W3/s9pKjv
uWE6DDAVYOFcCAzJrveR1sN8fJ7AXou+NoM8nyHFfUO2+ZvxJ3VAfb37D2XS
hxHjeJCPU6DX7lSNWY+aKYRiJmrqK4QqNEvCe8B7JYepXFcp7XyDsn1sTV74
iASoGHMojAII0BTyAUI7oNkUGPDvgsT7wNKOrvPVVzeDZz3MCRbTavNusb0E
90m+QCCGruY3RbYah7b3dQI7xszu8iB8UHk3fG5STwjJS0/+ThretTcIPG8D
n+M18KCi9UYXpnu7Bx06v3yhEWtI2ceRNEY+kjXxNzw9J0dHtEohzJC2o2aU
1CAc6yoQ/8P1OZXqX4xGjVnXR/F58lKLkvqWdVFNKhf9rcQ3xOOb2WrUmyf7
ZP648X2FSAYezWYwetu868qLVVubPMtYKqPmE1GkTMLGhxU673mmW1DhB1+K
vq+0mrrztBoJArCYzNv3qZmTJEFh9wyIBWG0es8mffTdi0khEusFMIrPUGrF
FKN+ETIoCg3UftwjG7VF09XG8vRfWXD0/yrCIWyPrVX6kMfbBejQN6lsx4VF
oGKfpE7hR393oROXOaD1k448f5jDOYH0s4EkN6bH6R8gcOjJe+D0ADZohTy/
PBRlwxsMewPOnAfLTXJIy91wBrgSKG2QX9WyPleLqOYN0g4nNANQCiHRXuY/
UDEqk74Z/eNM5aLlfyvjDDyUxMB2fJ8JfcpTR6S3pPnp2KhIzUEhSH+CAuvi
aVyT69E7h8cnrUGXBDF6mosIQ7Uyu/vOb+nqsY/GFKpi4gKIprJosbZibz5c
+4pgWY0Hc2i3rBoKfcmLdQCLNZEBQUPkRSkKLGgrFltUA4g+7e6hlViewkjF
jZL/D2vne5Zbo85MxoH4ImfDXI5jhleEJxSlbvTTLH+AfFBAfFgeHlcG3ePT
NCwWj4bAHt6uHc6BlWA5v2DX+vBs9+ooBoPF9rkVFutWvK1zIFenaJx/GIpS
HoI9YWLMMOewYBY6LrGppK+OLGLW/EDxgs8T0tczv6K6lcvo+1yVzn7FDU+0
nb7/rY2ha9ZGbB9i04cU1UiAoex7zl0ICg/5RSRdGBsDevKEEZRF7W+Qr6on
iJ5rcnmDrGcBPKzAVBaZr5jCUEL2xTfLlUFSrlgzl6T7R9mwOY0Ptjhku+mm
13RaM+d+hFp9N6QF481b64nmSNC7elD+3xfMt2QRY3jCTX4Faef2c4jwcnut
OkKV/S06dekSpPTT+bClcVccqu0o1ZOcJPkrniIfF3GSKJE7bjKeufc5U5WM
xAUYHEZOwuBToVmebl96Hv6WKxgnV/O6w9Qg/n+WzJyWGBqA/G4ZiUTNnbmx
Kz+lsVsti5eTrQMDZvNjRMX+ljaNjHlfgGsMnsHJaT9n7dLkd1I9fHbw6grm
PoLzfhMe9eODaRc25vDaR115VbfUtqGtO+sqz4Oi0OhI7j+SanM0k8jHvW7f
30YGYHj3/fPgTdYHKc/wK97j3yJ5wTT0O5RMp9QwT8Riae+1fMngEOJcuCX2
nSMw1U825o9HA6RhJinuLYhHR6qn+kDtXFH7KviQ1EY9zDxSdMYWLVGjw2sM
HXX/s9MjL1ksztwWNyUJcWuXTtwZJsX7lb3H5IROouiBRHdVPLEzgwAZJhSL
OkSauNGmZxj+uwJGiAE8foTBCRGLhXx0sDd4BP/QMKHM7Mm6yKaqMvVzba1y
dXpB1FWt2q7cc52tb/XaKLCvw93PuhUUVk1M5uPGCSRODU3wt3rlOYSEiRGv
KiUFwV+1RLi+Ic3so9ZIpvUMwGz3Q3MyAyKGS+I0rPdu8uBhqCFvAmsYmkLZ
bSeiWCARutOXkcCHBz5FxdlOVapWPAlmeKAPq/F5SmuOoEGMJx6igcI522WQ
0/9QM8Ah++dkRver426UDY45TNYovX4/0XBoWyQCjIT1L/dSjll6XHuv6eev
tijJf33UvhV/g5EkW4NgedAkrwqzxeV+HmpdYwVC8ZccX/hoCc2ReR251KNm
CxtFK8V3cO/0QknDKud5SHh8umFoYNn2HZHtYFcoPCal3Z03yiu1wAnDNBm6
ofAKmb1FLK87R4N4bh/jWZw+ZDeVaxwhkUvy5erE2eOmM03PX1eJBaUYIJk/
+IfNDQNAehHNqGEy7odmLSsvZenlIDNW/uTtdTaKOWX430DveMMrsDcLnmfd
0RvRnEjDEi5MxmwDqXK4UEq3JE2mwnFxstnnnkpHd4pAlCYTXeLcDdkUXX3L
ms2Mtn/Tk/k9lRgTwJ98kxC9pjRmC5Ofk88sOFoTLOa6OufAmur/Wll6IrrQ
06O3wHbEyusVgaHuIz/pT5NJycEMCCbGMz8czsbdAFT6MJNtuwmvkqR2Akwt
KMzD3L2+sjAYlk7QDJzClZkkVhVB8LzZZ8sEyukSXzn5o1/8RITnW1zFGZgX
FEHkT2pIjaLFA6WuQdCU0iXQArpM1k7IbI/0Anxwvc+UTzl/q2FUfe5d/j8r
RTkr3Y//Bn+ckjcUYQF2XpZRAjp9lWBkflVwkyDmndV26KW/zT+rmBvMOFUJ
7wCU5ImraYptI7bp3ct+8xzGlxinfF1tSyNFwjzbxNAD3Z8nsKXU/Ro3HILp
ESs5WOZh+0x8OO5FePAO2+P0gfrhQGNkD3FAKloLJCByx1apIfld2+OFH93r
0UqM1/UcoZ2+Sx2OxrlogOeNN/2qev7HgH3X9ujKaY8EuOdc1W4e4BAP+vU2
M8zquNFn1Z9ML3gqKA+JIZaBGZIE5Q2rgMWKxLk1rH6WNgG6fcR0e1+4SdmK
s6xzCJANZR/vZX1JZgegILOQ0Pxu9bLMVUH8AZXOWnWH2NVdAl6ZTHKtYaNL
9vq30IS9E9ZlltjvlnvOLUapW8Gj9V+OMa21FDOjBSzHqf84UV/8+DqfsGe+
Uc0YIHs3Km1EtrTb3FysPCcW6L0nCqOwBvCAwiw05QGihJcoRdmDXNuSLIf1
BnT2P3Pt/omHuOPJzZvlKj6W0gpWIEI4Do8b5VBo62xVe6fQU/VoiLc5ftTa
ujYUsljCj/KRGiDJd250mtADjuJqU/b5owGXnwCMbY4mUEy1WApwL2GR8c6q
GWPfPx0qKC6e21LU3IvZXQsRO0s6iDRneRRVF4ICHfslvz3iXwIFe6kHuboY
3LJDzaMeYCoslOvteLchE/gCkFp0cNNoF7TIhsQMCDmZxOB9+rcHy9usu3j+
XZVxHqf+uu7M0kPOGLyrV1q5VaKB4ha+OCVit+LeEuMmAugtHkACvRLQ+O52
+8vqec2hvQ4y3/FxGQ2ThVxmRjtpSzQbdqYxIvqnwAXI3F+7fRewoa27Mu7I
q2ZpS/BRvkzofA8A8fg02DI9k2qnIw3xdWSXFVKYqlQh8u6+zSibqpmLfSEf
UxjrlhEpoErXww2MqlsGQJvoyNOJbuYa834ESKgelSzWqzCUvv2cbQJ1XI0F
3JjeREcgq7AdgvjAf+W3ezFH9qnooR4hNgPiWwtbl5o+exfQNEkmWt84+PN/
1ro6c550W1788eAOnjD9BjhCgSU5vVA8jV8aNQBKfDOzVYyJ2RKEwOUkpWCO
tkIqPgj+82B0gpPHPC6/3Wgl4ay4raYX69YHgHxJ4DcciL7tcihliW6e//xn
+Pyzy8kmKTRoxAs3AJrczM6aNAVxB0Ag+BIPBnbUGhM6VxC4RAa0YxMs+Cxi
zo0Boabx2PMG4bZ62pCVvAQZcCgentb3k7V1XeaHzIXiQpCBSZCNHq7xi5k1
uo7X1HgDrqkAPt87XscXHt4VNgcP3ZqkD8s9APtrpP6/i5SJhurLtUWG7bsN
G1a9gOEH6zEqlG46TfWY/q+YmV8XBL+Rbx7JRiyCrGJtNmRSXMP3GD7+l6P6
xQ49mpzx/TcK781tJzZI7pgra8Sw9xfqgsiY/DyPsAZum3bPdfJtghTi3Ydl
MNT+0yrfzzpHTwQsTkosN1R7y8xNNyCCHXEEoNvtWNm7llVtb7rvQaeKejiA
YBAkByU7g8RBo1quwJ3++kPBwg0NpsyN+AQNWDxkJOltWuopJgUh9WzKY1Hh
i5OmRqKbmYtZ1gvj29BuvCZAH5oh1jd9IziTG8VrSpn4obP93NrUdksicqEz
2iTbiTG1fFd6gzot7QGYsMbd5cqQGlqpljjc/p6GTyCSw4DuX5AfDVQyOjt3
ZIn5yC1FWwYozOe0QlglSNE68tID1mAleCGjeTqPFqWxyaFFAC+1yelEbmKk
BIIw/deQBQNFp35ZVoDHZoranD+ZyQHL1c1YmPYCmWMbQQZP2hBpgI9FXUE8
u2RI11ma6qP99FwMGCsrOO1db6+ltYwtGYgIxw0iLH2Ge6YksX5wIu6HX25u
ckf7ViG56D3eBWYF99WLqto2sNMIJmXfOsdP75G/kiLoq5uDMjn9CsDkOv1+
8gLl/sYGBHZWwQ3dj3M1U1MZgu47xp4TUXxwMZzlYnM1LcIDQrdef8W4PVky
WcW6n1HzX3GovuiDKB1NrlWl8knPh2/hNgbVIJZdqmPiAIm8zd1fPQdq886A
NpoHoWDCjfVV2JVxjElIps51MyuiitVN87xoMU4Lo9Mb8+MZtw2yG58o1jmh
eYkEKJk9mjI1+MRHU5pluL8wP4Eka9hsMldSPTQco9myRQsEi40Wg26+pvuy
wVc5yEHdb0MY4w2arg2kmA1vhtT+HvKgZS2K5y36f3mmNlVGuWXbDXe/oi2J
RCNqJv/Mk3LKZzoVEBry83OiHB69LzbQpa9G+Ea3Z39tht4OYjUawkjqy1aX
FT4IY7Z9lVqmia611mHIDtavQB2glZMHl+KFHp42xBD4RlQ5fn3oD93eCqmy
VD90AhH6VplinuOVGnG+bJbTmoggUsJLpw8K1xKUSqehkeDcBwS2XMhVIsW+
ICmmPolnkXaTh8az0WEIhl+TOzS4isRTEjAIG4fMdFetdY2/SR1iO3lu9jBv
EpGphDW/qWKX8v+84Y97LN5maLX9ltNDR1Xv8mLWxQMze9B1e76rGBHBlYun
DBAlsBSz71zIIXOL5yspzFXz5Cqwzjzkl9BDtcMf4dW23KKJatkURR5GsGHF
dC8By1udDwODxSyHNLnAoBntU51Goa4EY3HoQ1zu+DmuGllBiMQUSFqdzson
+rmxvBYNX4Pij5RY8JpqmA5GQzB7O9LvfxLBJn/PYc/FM8+T4v3ZugVYG2vQ
tdGWjXvgsFwE4EdmEMCQFHWXTuk3QWsqamm0ULFcmzELd21dvLCOG6c/Aki4
/d6zBROeTUsHwqCirNI0XJpx4QlfR8F/bEm2Ivy1ODLif8A5RnxQgwOYCmw5
u8lJfgdlJ0mgZ9SItNtow6ymyxGS98BI7vU74NJ6kXMyt+54VNzAfU68TAUA
8/PeCU5DgnD2D4S3pISWS44GLNpf+mm+2NbS7zXKECOMKMSh7GHSWCBrvs5Z
JfP8GCrKbCND8EbYjDJ2HIjjn+H0Ztb72XJzuChGY6EuFdj92stUPkNrtDTr
42qPpQeVBfBBevPQ7eCSDTGRYu+LZolLYsZjw0XT6sfC3D6rpy78Ue9sKDnE
SkuufeDHNoDqlvDcDsEs/3wjoiOaPY18KPS7QoHnYkBlM5bypgYrV9/UkDhg
kThMBKrY+8J0H8FZpbQWH1cuSQHeuePeQOjqysM94u2eFgAsh7sEDVnuRifx
/tmoisUcgDunjaCGpYj+WrnEZaiMOZIX6VTyasn/QBYqAtX6dXJYnnyMgoGm
W9iw3adFyrpuUbwla/xJOOIVyUGHJOyCY3Ac0jT69twAG0mlvYsfZkaNDE/d
FcWoJgSM0lUvg6u1ct+NINdajBOKmLe/cpHTV271qud1MpOxI4wITAzNusYT
1ZeM4ylAlLAqLNcRY+JGgb8lc+3cygvdSxmXt+MQzFn1kGsSP4jPWElU5crT
nMBANAWyIQkxJ8Rp8vKwBthlP0p4B/4k2Ayv2JUVGr6IXRx3HZdlfOlyNhnP
aSXWfzi69DrKyfhy8D7/m/XI1jK+ouzYhHgwnjqkl537P67ERQ3q9tMz+pTC
7W7cAd956NlANB+9YvOto5o8xzwDRupyQKagpYFV+GBXWGa06z5MTkYQtVyI
gZGrPGLe6HSNixmyDYFix5J542u6TCrzJhJyVZCowh5JK+eJcQ3stz7nUUq9
1fh66gw0F9625sldiGTZ8lwSwUm5XanvrkB8qfV0lxigECOg0y7L032hYm6O
N+GKMRy6sp66HxYwBq9j8uhTcY488JsC9m9nj0sGar0McrxvopTk5kgYcbgV
wNWg8DewzSDt2ei8LwVO8aS3YYbyUWl4eWuGovtYOm1T13WzwB6fqd+mcE5E
lT9UsE1dTfxA5aIhJQHvk4te94jcOAAUhVLd4hPUEfK748VoIAStxQmRKB/j
pEpARU0sGkcV/iXEoTS/BSBYeRAFN2j26AAj2G/FKDDUSHLSHRfwRk2bw/Ey
vKVfZC3/HZRlPNQFJORzfEbWB2EItSEIQMKALUDbJHHkFtXqahECGC/AdqZl
1BYCnLwcdt19QyI8VQ6XIVkljpTTV2VdLZ/CRL84nEF9MVAkFOxSt+zP9XfZ
1/E7UNSTmTepbXDKB7Vvbb/ANq3OpMtsXvsICKt+cblDg1xl68iyrygh6hzu
5G1fYvCibbvS6cO2B6pi+KvelmybX+dLZxhQw9ccgSoqym9MYnmW0fPn9KU9
lewt3kslCv+JZfsGn3Ti/471SEJHyBGbr1C/g6lHxRsTDl/dUU3n7/L5JL7r
gSjUISneAmo5QGZIsWKL4/yX09k8Oh3C/VlcrvlxI8bsNb6uNaV++S33IpWH
8Pm2UyeaM4x8Sjil08ngEUoS/mC7NlK3K3blZ0f58pDhvq9hiU/SHdehnC9u
082Wydu2//zdf9l5MV0r/2XuZgHZeuRqKPhIPBcj4WiSZEmTaE7ZavDWApTm
CpGAxYJPfNg89h/S1eP97DM4DyONYXLGyzvWpNhxT7SJPR6qJIhw/cXe44QZ
vEU1xGQey77iDMpAV5akTLAl2vgTPZvFcL92s/cUwWnMtPUhd5aVMMOI6AaQ
rFm9oleqMAMgK1ebR7Bk/rzwVwJrKeHR2uwwYOGNHEaTtLvjh6xozclNZ4e1
radvIsT6rMkkElyXTSk5DtYU+G0/Sm7ktrmEYbIlGsmVwTDixZss/fto2yIH
U1yqYRZdIN4gIQD8b2WDd44k5BcH0xqK8SVRA0yWP9oooZE3NFcL4WdAryKP
IzgL4ccmGubSKsH4IgyvWkwXqGMS0YfeHLHeKv9ONdf5M7pl1E9IEuSr001Z
9hFpBllROLihq29SCXxTEyAqLEDmVItT+mb4FKMcshUftm403KpYaCm1C7v4
itz5epToxXbGrQNuMveAm4oxCe9SHwuaLefV7UPmWc3oYyq/VaODzxOWPYa9
WINOKaHRhUK6gddnRrb/msc8oElg0x0nPHbL9t+QdcVNU562qd5aeZWczj25
w73oTFffGrPvDLMnLcFtLxeeczShqbekfml0cApXLcxv0V0T0NGke0ARzW70
pM776k/7oG3XrWAiYJijJep2BABDV95q1p10s0nSe9HAYxFvYR3UE45ezxFs
Wzyi7y/mT/rJDs6LJcb9aeHkMyImAWjgxtFo7lZbcrf4MzgqfDxtGDzpE9FQ
FPBNPKqLCXN4R/n8GtFHO/uULzO9ugLg4WiK6Sa322G3obJCdALwHCPtmtQ2
26LneQULMUTgq4PYZ3ByTNbVSD3FYWZsTUp53sAsAV25qEYBUe8UHpkbSs+c
oagEYbyUP/X4Up/RtQkdkjLBvUQPYjJRcpsSj+MIhjn+TM16zXdfjhxkDMOF
3g9dcV4KJ/5zLyUiH6UesQpalxTLHm9t8jsANrnHVK3enRgFXsauLSqsJH7r
PMzPTy0Ke6RemtF25LPrVzk5d3z0y3dBbZAvlZssJ3TVUeDJOYFruyg/Qmcc
Z5LvRGaE5R+cnkz1P7KaO/9e57T1S70GNWE6qeEvIIl3qqLWH8NKlkRsrfVF
sw0JS52ugSgmGp+Jei5CGqlIS/vByNKnvIvYMJnqmsUzi51qNa+1KX+BZvQA
YbINNZFWhTlmHs5v+KBb2Oxr10aIx3ut6C5G1vXdIJFPC0/w58MIHik5SR6u
oW7oIxzHgNgvzAOBoAA/9Q/XZtoL++V5ULI0rnmrh8DynE3vdYOw3pwDDmI/
4kWewi8PCh084Itiq3ToNP4OBI1/B3cmNK1dDl2MXzL4mQpSKOKJhg+N+wR+
zTrTGULX8ccsqBlIPZ0WJTYHrv3VMM/bI6GoAGSxBCn/Gz8ksNWGcj3GDPyV
0K4V5wXHEKvVFZpi6nW0EgWhobpKBwBOg2wriV/cx2knrtS+U2D5K+UqEdF8
j5/MlAe8RFNxkVttTz1polHZHmt0ZUTF1Qmq7SCytM11AlLeDEPPcNJgcSUJ
KCUXHHQe1lKf2qkIwsh7XZPvryfU31dGiNDmlpAJ8o9UfwQYsWGDvWlfMk9T
HJyJ+GSf/TfYq6W2+m19myYDkt2FRU8DebG3fWk/7pr9lC4wlTwkZ2PuM0gn
MVTcj0Is2DKCA5ntko7UwhExHKpY0HUejlgleDOEN+yOMrx/EMHh05DOZ/RB
QLh2apc9hWPlzLizMjon+/jEgPy0bOvyWEryurZgS8S+lgC6eNHoHuvGfCTm
btpelpSxkijUQT95BG11csJDiHLo1oGHN13ir3zs3NEQiQXwc7grtq48b9mv
K971DB9afDa/SFmmFwttb2njlg7+sG1pVdeJy8pJpDFzm+lGlAJ6hKsbxxym
OaksRo6MXxzkWOfNlgIETOvZxcFI6drprrc+7vVx1kiscAhdnx5QGFD6XG0c
kUa9bMlKYY4vNFPqBQvaGlmtEjyVb348KAEZFtfPomaQ9NAyxOYRVHF0HOHA
/eV33gmRCFJ/EpcK0WrExBH9kQhcoW8cTryOI0GWTr6244cBYTd4IxMVkdbP
xtTiqwGYJOq5mtkia3urRYYW1jJLYqKZK5kRzR7x1fXHosygXJh4pust38Zf
jpKbx6bCMmcBWj6f5O9XlIypNOMX1XDEuyBL1+pQV3hwdaZdDvauvilclneD
OdwSjxHV2G064zhVthlIx807kzNp5pnGv9ZK6aJ35skKE2D5Dk/W9bvaU6dQ
1nsTTnyEHgXbAv6CaGORQQ/4D74AAx0vDx6XOJjc2LYRfK9GgNe6ODn/cLE7
u3h6AnJjRQOCPYCCQv7rcZmGiod6OVKqXbcxL8BfhhriWtuvD9JOXPaEaBU0
tIKm0eARFSypSZZHtSIAll5OZ57Eo6nIc/jjnWdxNOCDfYkJ0sOjbXgUpaGS
lFwJyUCUdmZQ0nItP9R4n4y3GF9HfN4hVm7934/kaItd2YjyCS9rIvG/39E8
MOYauzZtlZWlX2THDqRn+q58wGHvv4DpbURJrMUUVSAE+h2QqkcPkiisgTRf
dWy0P6dQ3/AyB/H5w9S4io8ZVee/peHWLOr3Ua5uDiH73GTyytFvcdlY9NEL
wtP97feP3BH6FMD8TJz5f/dNFi5/qpaCHgDKJZEPYCvt/ereApQoVprlG90P
sOlHFILdoktzRRC8pGz4fQySgDUohvEFq1JK5S8g1vacEMxMoD3G3Sc7IDpR
PY7HkXkxIJlyx1qRbMlu+ajSD0o7IAPlGTt0U5EXill8C6N874W6hGx8LhFi
lySSpMNvKeQ1S57Y/F88DX7GKEQ74eazYaKlIbsRsHYmU4azswTZpBGMTJVp
NMFC/J+tDPSEatb9hSx3soKTmKdjigvhh7iToWqneKQNoi6LqiNJ4gpHLN6y
7Dl9+9syqLa7+NcC2yiPeMIoEjop25DT2PD3bVzFvM6ujkzTQ8XG31nLKDWc
RysQ86foKgIxWyZx8bL5vqbRaxnw/FxhIW+mL6/3E7vNEbUR6swapesaI5/3
BCXPJ2v8/cYTEG0vW6K50ju0nvW8lDzV1j6o1qSHvrA0ZUvU/bVjFyv4k55c
xoAiPKoNskfbEwREWnIdjl1dr8sTDUL7qnkL9T2rQOgHAsEFelKJppnxMZCL
5ZF5qVLmwyaGqc5yXEGMN5pUV3TpIM6sdiFYHa/9Pbzr1WlWg85UvyZvFE5l
y0b2yAf62g5IGlBXaTN4428xOfd8OcD4ik54uXP6haTVFUpjSdOLtfzYRJA7
32H/ogCcfcF3AWM5lEZZsxGRF1DHhevQ/mIt9KvlqYNznEFHd29LbYFQJFv5
dTQwGjsw19ZZ829WX+eGGOPuynu0hlrPHuSpr8MOTx8Piz01dlllNOVtVQF9
jyhRKI30+h+M9UhM2Px4HK2j+XcWJiKovHbifSL37ZrK2eQRxyMsNhOn+vNw
a8o48Tb4HtlSu/WfwWTy5jr6cZk9BUrTaQZT6NSnJCVeLjupVolYQJOTsfFt
+d5XU79OZTvOgip1UKamasAJFPcHFKpCcsk/D2IG0Rwzi/6I6N7WYa5A9o6V
CTYUghep9nLpZdujtK6ud7fSwIaFgIuisEX5Nco6X5RyV+mNeuydSPD2Ahmp
ci7W7NnKtvlf8aRp/XW6MXuSsSb5Uo1Yc8G4rEbq9d8nE4ed3oeUpkA+Bv0s
nfWoQxWcFgT56/zaRUmPavJhh2D43oYwNxTyJXqpTW8xpC2UI4UKzxRQpnsx
sXtlx9ulejTVS3IY5iDA8KMfze+JOG/Ir4hOD2bsAV1BWTzCX9dbsfDI6Y+Q
l/kbArGg776wMyHjvzTnMLMllSu4PxHYUfqbOkCknUD+KNdLxBeTpPLnAfbr
vy3tQs0yd0/o2k2K46hIMENfEMtAVr3hDp6fQx/ljVpSk1ZtboxHzacJpiBQ
l5gIA2hbGUcclOX0NKVW0088mMqdgShYGZwteIGlZ71vw7N8qSXv93SRa4At
UPue/P9oqHEWsiTUIr5Vi1YhHfsjyzrNZIhaDpDWVE0xCPNk7sQ8V1xnhuaq
hGgNml06RaCWhgFt52M+EdhNQ03sOZvXYffF5/9rr3kkilqmflnRKEr4Ukez
8PXQgL0UhxzaZoyx+UlmOsQ/9DQtCnRGn4l2QBWVVH2Wh/tnC7p4KsAknbDF
9UeKFpk436kBlcJ34CFp4XU2pNJi+177h4vnKCeahqIH2OzSIIT1kkIi9bN7
VjF6o5+JtcczTbtpt6s5fbwQ0wmuezIITDR49B/I77QvrJlxlysz2SSCI16+
pKMWc2M5JXgJ0BI2Jb0jKnu2xoxuPIpncvjzWAwfJPpLmHGkCl339/mTSzn+
NjFOjsB0R9t85A7sE/5x0M7A/snkryt+mNz9AEOWxAzo4wezY51kG/C6f8kh
+uR+usMvCgOQgcMA8gTA1dNFFlVALLaX8FuCXd/d/wb8POUDbanMR8do6+ey
5X/4rERAJXMGy2bSHNNGRa5/cT1BAOIUvwS2izwsot17Sv/qegv4Uovt4+V3
/c6TIa59ZxS27BbQm+1I15EVcfDuOUzNp4h51LmmT2hosHYt6qKcqbcFOPhm
2UcICXTsiWBrIPAu1cvjYQhC9DqaX2abXODkVSaDFevZLM5CH1l+iVN5IpqQ
m5XvcoZ2qsBfspSeOyDkgNXOG6P4ms6RGoTM/KNTL9GiqqIaj9emDYrdMy3d
V+C3SshVTJ4XOCRduj0hy9IbqosbC3uw+DcnJ+Yaqnl04AUjIkOaHTJOmGsA
1xxnSVZJasgrvn9C+e9xqX+b4BYDy2ZNvTh6Ph6fhDvmOihCPGIrTqTSguWY
jpIBQvDfecwT1nNuAVbYpBft5P4ffiV5QWwlrKUaZY3T/nzIrI+3fh0+bP0Q
NnW13YuvjatGCmX658cLRYxvOChLNfq444XuxMe8OEYDC6yfAU9940vvVWvG
Dlkg54IV/KcS0htF3l4gvQl5+eN8ZXPXKTrWGyfy27thpbxVY1foNiHThkdb
vvD2GSzGLJtQA76or44mXjiuY1hZWt7ToqliRXQokDuQ1P69Yms/+0sO2ZRS
g5BIxEkoflEoNINyAefJA3m6RDqHFPriJ33TN5j/ophIwmYqCh15lu1BNoTo
YHFg0sERaJMQZDmy09tY9VwyAs+oVJkpp0OnWGzquKASRgXFOn2vRUusFZiN
B4/7shBUYF166cDCQSjMkZKTbKpltWwcxDdskwLYdmR4yTxeFRHUYLnorn46
Fv9rEpJtag32Nup5Esc+4uOCxikG6PTJhgRQkqFXE2OiehsobkZnszuZdABw
hVU6xFrwCp9IYcGPIBPl2E1sBxhtlKgCHP2emIC8uTuXcKx6BEUzKqi5p5Qj
5k+DDrpT8Z/3rb5IHzUos7xFaiowrEZj9K2xovhOIHUeVIJntHbYx6BunCOi
POl1wB8f7YrVQSWza55E3NJeGcXbURogskEdHKhGbZLcboGLrCkHhXYMO5bB
VyHBzGzRSYBe6hS9EoXKMORoJVaFtO9vTShyT1CM0/skIfgCl9X6swowCDKZ
6Xi2A9Y+wmyHNfhpCx/RC0w1jj6O36Qkzaz2i6UehiCK1dH9Qxyuen29XJgz
+3I3pFd+yM0UTG21fsynyb0AlGi5J1X8iPCW6Wu1slvUGpVOlhBJkzNlw/Fp
k3j5wE8wCDKJhRfrbHDg58LIW6fPQbLAJE6X8M6zVn7lmCaVu4wMRJBU1NXC
1OLZTY6VpC1LgK8ji7llLs4BQBYeZyCLGJdT0FoliS1Mi8efRsiznJcVWkCD
n6M1dF62OcTw3niSEa1qtXF2ZB0W6U5YRvryXD4w3k51ytvXLNIECGuQyv6m
ozTj6HbJn8kjURX74H3f2jJ8m+hlFZo2JmzTiQFV4Oie8WyNNhjUtwBKvFqB
xW2tgBP8dPsRLvVy2jOy67qywvlbrWLEoQ0Afz5/Hmw9UUP0IZKF2lfKh2/6
1ZeI2GOolXYlEjRDxzOsK1wjpUVe2wfaFUzqmL0/slrCKJqwErrMLs+YKlXl
MMqYh70+qaCyrsc0q/BOuBDXmqtkGAT6ca+6E7IibYtzn4mVl+MEeGZSu++A
JCiENLCpemYDENBt28x0qUCd+OWPnwoqt57a/+KdDUqfL9VlVOvnrixFXlCv
5MHJOhI/CxATlhNHA66B54+BVnEi5XprwOwMT/citMkRrtkLg4Ef9K3Vh4uW
X8hiYqsDSVPJW2tv3WWDgTutYAKJdw8rLgKdcp6CUsc0LBUqm7HjnjHbS69h
b9WUf72h84+i9RqChXBmF3kV7CK3JT9x+kEVsrJZZRCNmSSPB35TTK5yIhUp
DveS1lQaKovVnlEya90oYGQstVzMgP34rMku2ZIXX54KogszqPFy2BZUQ56g
Q3cj8J6dd7ybkJXnw8vzaSQ6KB5+2nFNYJXePgiL5O1eYsmAgwuz52JL5N4X
PugP0MIbFVindSMIeVvLDKJaM3GDzOdMfPkc4mLikrBtoOKp6dz8ZS2D3FHz
R6obGXRPsZF8PgXP/mbhsZ/XIiOBM9FI/FUJUKeDSKYkuRjvdeqhmSw5ttsE
Oz5rK5OQl2M17a+WEdc1irom8pnk34gKkY7ZpyiVDDF0vHdJfYZEcWso6UR5
pKajqkYCAqU9KgGJwf9WFmBNYCQWibdxeDU/xV1kOG+FaRNZ/xuuTx6OD0d3
HAL79DseutmLlbGbX/vK+tFo9+YUkuGm2lJUUMTVLAXla0xURRvX9iJidfW1
Apzt/0IbbpkH5Je/ZtS4XNOVgFJzYIuN///+rKdGZ9gYs569g1xwye1wsccM
HFKAIEby+/v1qmsFBSAcHxWD5RWFIvFCg42lBSGLxrt0UGFkKsY+EY815WWX
kBuFTOvi5WczCRVNjNuAupugnCX38aeAPXDTiqyGKZtz/6x0G8RY6kKDQYp9
irYVqIYxyA3BSdOxS0rXHofbdsrfMgw+rnD1UAQ80Nw2tzD6Rnkm7D2EgClt
Ju8on3t95By3jVXIKAaP0I8usUXSEqx6qZOH2kvdCRmMUGebM49oJ1wzNiWY
3DH/6Hdl8Z56Goj2PU+AzXfWWrkBj14uOHzD8rN7G9VOKBoEj6d5OWMl0jjY
Vf7A4A8hHRnmNWdTA5R8iXM1+o9A4AiG8bicPG4n6kfkh7JeX3uLoVBZYG5p
EN/pdq1jQBKVIoRVwk2FKUgtuxYD0rrwM09fmaz4z5HPnEIxVzPqJpToYyTF
mRH8/frtQke4dCG5YS80YYNRNzDSIYF1ksiKWPhIx1zzKUIyzB/Q9q8Ae9sv
ByDUKC+W7Vmgwky1uQwbovvze8RLf+luIDTTk2so220lovV2SBj74KBWTAtP
Z0BZMogd0y1A9Dj801LO6x98JKRabC/UPpY30dfBppdq17CogJZ5iyYtwIMS
hCq1mFyrKfqeyVXhiRCo/eshg5pUKBF46or/JAL5gD5ZfhGYhPUDN4Ma7QbY
pZRhWBCi3jhkVjPXuTb3ZqRZuYl/sJmYmxqfagQbdF7Qz1vRV/afCYkdUSG3
vkxAMCUnVeWSdQFOSahacgGKYpdW0MORwjGVxdvzZTVTT0hCv+NZU+cU9xQv
HN9+a5PldYyqvERym1mPZ34R1G5TDDRyP3YhQNtVZ/Dki7mvsfUJzFTWy9u6
A+lOjShzOqn+S4rkNcECYlgPxXBrZjYIkevHeaKJhhZZhPDyuVs/zzYSt6Yu
d/Z53AWULK4eov6+5yiDzkjHyKUUQoBbWDVgKZEmr4cHxym9zRESFhr84OQO
F6oSCQ/n2aHtAyq3eX3442Z8EpuVRuUnZ6Qp8PiAg1Td4kn6KG4Tbjth3g3w
HEScm+RMCosJix/rZlgpaMpjB1FrJLNyWdzp30kZF9QJtfCkHNOSPhV4ZPML
9snLFDwqrX3K+zp1TajHlV2N0RQnTp7RNMGZocq00vPnF/YEOYRWLXuorzYe
DXvyJAV9nEVyCpmsuxKUHAyv8S24pWgA8nDopA1kKtv0NEJttzd2fTnnD6HI
GTHlE+ylUJGMaNmLn3GiV0gbEpLEO3thE28uKVSGz42AZAUARrUGnCa4v32N
EwpDZTEswhy4vfwOxtgaxmWNUbchGyxi1e5OjR+SU5IGTNcBZX7ha3jynlqx
Dbn9YGRnu/JOmBh54QaSTrxycTWp2BB/3mlBB1kp7VkpW0aI7+8IPQt1MAzE
nuI+3ixD+0zHoLw3DDBMDB18MAuUFlbSTbATt0XxRaQahkiiJ9GS6NMAhIs8
qEVeGI6BmBhFXEZFxRzy0P1cjXz5YGpNOcBUMA/Ks4PYEGmIPMZnoWPNjG1s
1BCNLMX8SEU8lR6SkaWuYd1GZjzIKjBTBynVdJo9/xA+AQ1a/wioxbZRBVjL
8egiEQEb0GudVHYU6PkJalpYzhIDUo6IQCCnI9by3a4YxxIVj/WRpEDuQyN4
IlREaQ4+nE0HwTOwq2I2hBsmKBwFy68JVAWOqJM4oUgEwLXoZEE0DUMrfvGX
HlI14NUZsX9VX4P5ljARBxKwVxQjZdonTRyTldHnr38Yx+p/0DELlqQqkmGI
+SS0O+TX9bQhRQp+ktHvlVk1CrpO0+yxC0xMUBbMosBOcbPbND7VLJgOE5ty
pdetnH2ZSaNFlKQ3UkXAtSjC0Jd8a0KjGsqdaHYqxywmDEo6Hov1XdGtxqoA
7QTOLbA7tYo2ZvwVrw8d3c4CKeiz3fz38zGWUySzFXamud957EhuX2K1ZODa
eL16JriQBmSulXH48GEk3L5TNdWWUiN7mm4clpWZ/7oHcQsxNb/4aXvFtBOk
2972YLejsCEr6cY9/pOP1zlZYTCvvRu0Lq6uqgJrhphotzNrG3TBWzbmsmz2
psiRrGY7SqzxGPPyohEHkG2rag6jNOrxffwjo7ftfyELGdQEpZKkIsR1CPRJ
Ie9PEAI326oe0p+xODw7bxRwreYNyg2slc3gG5Oobur4q/cjZYOrAQSqLiKi
DTsH2Tk57vulXe9ncsVev8acPghkEfRF3QDJNJ+YsdzlDEJ3lUzTClW4gtkY
7HrL7q1PrjcmWFwazcOmAcjEZIj4cl/uAv+E4ck/dwNQ0suvgm37M/EN8Hoh
V7fFLf+XSuuve+q4i/joChlGUfj+7gxm12LQLRkpWsDlR3vV691eUnSA8MO1
txDSm7NhgMZlDxC6H/gJMqy671SNLBD3iuCBMLgdaFwknNNF+Glu8tLczKnO
6fkzizdiNR+4rz0dpWnRf8YYdsIK0zm0aBaysARYQ8EfXFXrunSqGPaWPqUI
kdFqIwLJypWxbpRmP5VcnUPylU/6WeRd2ZANpguoT1EYELcgBMt9pDrPSLjp
zdSWInkCmwFkmRRZCuQKwOMZjiNdXyuRizUI28VaGLznifXqfyNn196YOLkQ
HvtXJ35VkLy6m6jkkWLl8AfKal7Fd2q99lnIibOPbmnNPDwg3gNU/l0zcLq+
aMGHvWP+XhZHZYtssd4CecqGiShLJCTGRElOEZrozCttpf92k1x/XCRLxTDO
As5OGW4kJnO57Q9Jx0d8OI+wxmpkE1rmUMxMfChZyPabE2pb9rwgj1dcwpg9
+tnfxE9jCJAcera4bOTnYQvbVfNloFcYvfFb9yO9laCABx//WKOT000UjDJL
BtmxebQeRuqXc/7FpIpwd8B9VbBBj4WeTrh+afracDz2znDW/dIEcZozRf5F
zmYxN3cgvybxVHRVXE6UANhClsjEFrRk2VmXur8gIM9Gh/5kodMt1TjfPhEa
VbZlTzlz+alRbYAbz0ypBnH9i8btNFN3hL5pcw031TpbV+1JMQgRpk+7NkT4
Z9hMsv6IHFRUy07aEx5y5uGGRegqlpOjyBXcO6qjZq7GSIovXzPClr5K+B1P
X6lLtNJBcTa5+X0BBvMe6s5leStn0t18TtYhP/Dvrm/5ae6B4Lo2mWyPiMjq
hrPkoiOPJFl/4rT8D8TBWt2I2izyjm2r4nDa8kZlPlT2mBZI/6DDL4qA1PaG
m6aghLErQruZwzOeI23jag3t/ZDVZyewrOzq1Ll3VvWVI2orJ0+t3C+nZRKE
G1XUOdl6xAErZqfi0RdSI7KSEzT+p/3ik5bzz/6Lz1MgEX41vxtZOD+Iytp+
yZHwIqlKHG2DfIzV9hCn4zlnd8YyXgulw7l4nHEoIEk6bUxLvwCYSIFXJjHz
Tq+5rAX4peGKyacAa24jkqRQuH0Drk7DsI5UY8D70OSyJkVKw+SOCU4aT+xG
88Y+9ib1OU0PTwQvj9tXFYSlYIl6YrZjePzLV6gIYGf7dR3Rzyw7mi5snzPP
GP+C058MF2O55Dgz2+nl/fnG6J3H+fuU9xrHJFAbRR9A3rqv2FTBc7ZlLyJ+
MFCt2wLFiDs9CkzqBZ6V+fRGPUdufBvjGiPLf7yRI+OtQ+2HExD+N4jE3EiO
0b14rWRZ258uhxJeLAX3R/lQm40uCyMzfnztxzx9jG5fE5t/naKgp5GTfUYA
nd3nATGMsXkCnflgLzFAWrIK1eAn/x+wv1U+IPF+txewCaUoFz/4Uhr4AmXY
+1s02RGnfHXL5ea2trOUjAku9gDPqVxlLq/pG1mayLk/hghX4sXzRNFRQVpS
8hTTxAcfglnhkjIHXMWlXXRgmeDqq2piva2t2kCKm2bTYr+VRp78hhxDkgKt
5Kx76fxsxZsEGl2hAWeg2Jv+ErsQN2glOrg/GsiTFBp5U9AVyMSPTfl+HyHy
K6sNqMpGC06mgA4jhTgUZz5YLXvIM17uLMq9nYRX7qtBPbhA4rhMyOuOCWcr
4LtCR0Vpb87ecJs8Ozubru8vVPW5Cckz9tUA2VWhWciQjzCxMS3Avydzjn32
JuVTc53ulK5ah3q+NjA9vP5hXtCAeJ69Uegzqrnfeza/4MsVWZqkWJA8ILcS
r7A3N+fhXeNpUrz6c4FzG0LVEq80OGuLk6/Rl0YkWOXJ2l8lxooNzMif5z1M
9sdNFnVz1N8OYq852dTwTq5NYskq66070ZwJ+ZFwHxtLdYgQzZb4lcWTpOQd
VMj4Qby9L+S8tbpzODN9ovpUG3eta4f7ukA5a6Tn00OXxvBZObhOko3af0UO
jcjt/qjkwjCh9sfwRoPGjzIIiUhvapLNWGKsWNgq8BJ6QsIZFsgVmXRQt328
mpLKWVkcA3VdBj6LL5HjHyrjrWFZIW4VyxF+g4N6CTlLou2Sn/ZHCpcUpd/o
fCEUPrHOUqTuZrLysfk0RRns8hO9VqS44C80cXXzep/AImlLPpSmaDfGwmlh
OXcsCFnPM+V/E0e6kFkTBMJnH49yWumZN4B1rnjnezYO4q0YRBOao9cSubKE
k3efJ3Ah3Xr6nhjpuX0aeZ6+yFq9AVgNLUiQMjMQ/V27mnnCUpUJhwE90n8P
ed2xB0HxLkeloYyJo7qdukSpOLIpup3RC/KjFgV2BUUUEuvoPUOT8Gh9Zm3C
abHgpjNIm6XSAuygXquaK0/W9SdXjdWSzuBMHMJ+M8AUU+zJwp+YuAie6SGR
k6N7fYXKgHxB7syWzrnxhFSI+2BpO8Zn0EdXdJN3GSBP6Wvi2amw9SIgUsBq
PERAjieD+evuf8WK1iUR4CO2RTmjWaLiwNzIjKSSo4DhPr9Avvu1wiy7SVVA
36/uVE0/FIoidfRn4gXBUPdNuAYZJm7iUuPF1hFhKjb6EvtRqH505H/RNKbJ
ZWU09gcyFCKljw5ZcdFlH+vdjLBNQsrL2YK2I4ChdDfbhH1uvVhjnuxEPBfa
XygTDYZ31g9QjGC+C887+C3DArQJR5GR7mOg7nxnzHW7yktkJ5cUzyb3bjnR
IM2FwD0IBw0Soiod/gAS7dnThNrHt8rR/REPSRxXDec84xL/3hT1N+x2yN5F
3i3jOzAeBwbKZJMNHk6l1+mqQpDMv5qqQtkn521B0mqCMf1EjcWQdni0piDL
T26yzrDlge8tYyNtNdr3p6HXieSg731kttn57qvCUW/TxxSzUGJAK8XkXt+u
aioyenF1bYke7VFCpeOkyyxSUp2Avo9O7TpslBnnktskpBz5ppJCb/sltXur
nD6F+ZV6ldrTEkShuoTcCAlAoNHrCe4ML9kJlC2zY70BSSywTfGBbBZTXFfy
pUdfeGuZfEquZNOxmOAZALJcjLNYBi9FKpRMyhnkrGND3nqO5+804LJvGGoM
njEKtd0KUhWPIMIDUHF8vEIt20xKaRY1TvQiUwqJMI0Q/GTex4XDs6S4YfDo
OBnaocmp3R50aOnmwTRldJtrt0X1EUds1KyaPNwNPLh1JbarkOdTji1PW1u9
+0sYuQ7KztFjcUVJkSDdZ9Px1CuJ6l1lhSFxDa8g3zley3oAf0O8YopMZk6A
wLkWcYWNVT4LZO5jd/773IoH5Zzmk5vtS2orc9ANrt14McyL8jCRk2o3ZOG+
pGZCQj9rwoq+gHjfJ4P1rDiFRXlFzFisUNTaX8Q37NcuuJI9Tb+tu2smL3RA
Kr4mpg0V4FP1rAgIxFhCxNwBPHohx5glRwNWmkBYO1VmZ/i+V1ytV8YrtCGG
DYLRAPtMCb6TSTGBcQu9HX7nYcrzzIn4HYIGXnoXnxeY9d3tFdbGyfL7qZ9k
Qqi1M7M2vSOuoudsHyFvuUigmVHaBg8Otiv6fs3xtGD69/En0DP9s0N229bm
pABk7A2CQUtSR2Q/w4wjnSiH2WinkEvku8qHHPx8DltDk9q5miaET4JYsd3l
kgesAK3gVBhN8FVVOvkhNmjx0zPKr3F9FpBh/APxXjmIg90XEzB5iE1tL12R
KH6fJFd/FFQCC/qmxEuyyhmb3FB9aoaiPKXmCXsT564mh9ONMX42yKa8V6Ke
ovVLBYy7RpylVx0ir0mDIxJLIzvi+xD/mNujjQjc+TwQVW5ORKyH2NIxfFbE
q3C0CyqAS1qUOCLJBpzb7GZn6vLdoQQ21HWxKzlxNZbbPoTNabJrBVgupPwX
H1vE/VE+cMWY5ZdHpA99Wa/ogtb560avuadZclEz6cHyR7qUdNhp+Zdt9qUG
H3LFBbRdFDtK4JrQoZwL1d8DzXPORF9xxcI4usdQBvQISKJa/rpIW002E2m8
POo7u8IX9nzO7Lo1ehu+2sMelD/4W3yNjC43VbWp7ABfagH0l308fUiIX/Na
uyNbJvjrMGxWZ+LTplsSvUku0ycRUEaOrv0PVTgpwl32n3EmgidrTl9s+d3L
EzDTRUq+7yP3mmJ+mu5XENOwRed/XJ3TNmq5DdzBOSvoBRyWFwiYiSTFT3WI
jyDIUEfc3Fx/v2bFjmYjNUgbplqbTIwo0NWl97BJcKQtgOsO3m4WWyi9BmN8
WnCbCeGtSKas9PAY94UEHgYNdslF0yj5YFYdG8Kh80QLKNW1yv3641tb+2Ba
wdUi6MN8V95X1kYSP3W3RX2h2Q4Y8dEJnpzQ0zERmD9n6MQkc/tv3LqaCKe9
/liRsQUshVFURSoCQ4ZCTwxRNmGDNPjpfu0dc1x2L6TZMOTMK3tVQbhT9MaK
47WLcUbEAbUxjiVaqof2gpWvG4mF5t4/yzGwpgx3A0eSpJlaRbmiLvPCvmnP
PSyJR+fQ/6UJvW4MgNxaMWJNaiJFY3sDTs2mPmcbZ6tCZX3YXFbsEAETHT0N
7/54SjRqMq8a6wxc3aosCzA8WxqeZMHVlL8K8x3CSecDlZYgONcqNYyIq2YK
pXl46EifWeBlqxNgDQbV64+mAR6aAWUN7FvhCRzthvy7Fz3Nmjdm1Yhn36kk
j+J5w/tIGhRTHF5ZYbe0S+PF5Otrvwi1RwIMO70sO80U2O6HoOuAmVSi13e/
gi9h2YvIehkU86UqzdTFejl0wFJF4BgBYJQ0O90aBus1r3U+2Pu2VOlvaM8n
6UJV7fotFL/ImcVSw/vJHS99+zOaDS7NMXFxS2UFdQeIGaXEYiJ9zhTzW39w
0gVifwbhySaXwljpWrFVkh6peLm5FGKY5CX9m8L0c2azeF3DvMIYwIA6mEYP
2/gnrC5EM2rUJP7gb7XVRoMuy8mla9DI0YKlzFlGKTrsYdycIJxOa/CVM6VO
i9uR609CerE6LJZaK+vTuG2cbRFuIbhh0nu9uH/hhrJPqLdO0i4j4NR55M8E
qkZSp4OG9vo9ojdEcNMNj44Rbk1d2LLntiAPyHNbGJUOqZIDxzhvin1oFE6j
9pWPDy1kroJaO8MVskOBR13xRkh1lFcIcxCaGhxj3a3B2HbXBuEFef3Wngu+
eigCionsTA0snIR7KxZWw3mw7Wc0nTWrgYWHY3cL+B75FAeLPJY/ot1mfwfp
V0iY7gkX/xUmWCNsd3LK+nh92C9oByiCqdjvudlXTVzXCbgeQ3Zw0k2LzVo5
P3ZAdwHEsdzo7oKLbHKUDhgOqkJdvxBoYetL2OvX/0+PkS65qsWGV3c3wKd8
hMXy65vgos0Ulr29f5nnOJ52rYtKQRoYYtPxDczlTH2MnhLp+E0WISIzXDYr
AchCFMTQl2RfJklLZiYvABbxAOkuQhdUdQoteh4u3zS41TBzquMG3UlsgSgy
nnRUapNG+WvvyO0UH0UnRvTCvOi4xbwNnmvycEJm2AI/vsfY4qGSDg2pTTX4
YCRvWX0AQwuLvEfBT9jmwlw/7TLJkAs1M8PLApgNH+iVWTjdym2ot01yFC4Z
0aiS+ApTJfDvsXaVKZDwm81u9aT7MWGle1M3aFj6uOulP1qW66g/5YVd5G70
qA/d9OtCxao07lOKp+EyZxoBFj0vvgDbXkj8MSXWvA1R9ur0sW8cOjjM3BAd
+OZBzq1VVFkFREtDiK6yxktIdq7GzMMEbAx8ZuoLXV+uv5t4layD3WxgOTVF
Us5ZvS3IYaigZYtGtyVZWQtdkaVRPiN4wbFZCxamxHo8KT8zp0mB4vVvy98h
8LkqTrGvfqKSrQmYxKFmwkqV4l3dM+gxRlFSxel7+hFemsGRp0iHgXzb+JC5
LNtrxi6hAFxCKfzaYrpN1CMFc/Sf2LLsZ8PoqQrbnUAGfLJ9ZayUc39rZy0l
bxnrU8zRS/3vxrFFHTsZMsiPetUonJ49kUz1t5cWMeKnGex55do+8+XpI0jA
lOYxq5e0lr/83RoM22E2LYMyZBEOM/v5HyDmTGIUWo28F5e7ifj9TEBRZYOJ
hAcRGZDoem/VIAo85/8XnxXDmeGILJN3rr3ZeAQUmmh3RCSVScwZVJEyhCdP
I1oY6zDOw6RDmnjPKSxzCNfMb/PvBu8KQjwweatoqzOJKuJb+PV0LRGMRUyV
NcewdhxclxJ5TWb7CqRK0hbRopb+hW1EqzAPx/zyzUX0WJZlVN2Up76Anogn
J6IigYFJiYwfndDmoTvfHftRwopXjDb0jaAmz48uoWvuadZ+nnPCf8XenfzD
8A1XlwLIwlC6Re6ivGAafMZd4dFOKSGFgctPRhx/DSwQud07tLGLBXW8heu7
7mzo4GekD8UMlzYvMoxtPzYqQDqOTylb9IUuTDb4v+Mq6UODAWw+TfH7ISnf
dIrgRUuVQLlJI+me1yWI+Pm9M/ha1mCwrvuS5C86lklnYfRz/e4rTbv6HBt7
RhuwHljpa54aj4PWc/fXQE5u4VTySU43O1vWX8G7lhTb8Qsqox3A6lTJDnyO
KgXlr5d8+1ijzopdoZy6+9E5ciOkSDiSFDT9IehHi0M9tCmhqrHC/vlbhwcp
vqSXRvH8Wh06XHjLCk/S2pWPPh8UPT1I79EkZ7w67Iil9aBe/DYYSEvP8XrL
mxPwH3Ti/1knDBb2pv1R1oFMCNWlLJ7UVWTWSyxpOp+wChfQje/vCzSIgZcR
5Q5joE/+P2bjgEMJ2ug29GTo0MKsFFsJGsEiQp/X9/q1w/XILNjy4wgagzUm
cv5nZGIzlsD2fJNash0R26bGldEBk4v+t1mu6pyO2v7UdY+Nw226XRLp4OY5
55IsmQ4lJmyl7oJB02wgAftwEoRBbwJMaKM6yPIEtqvKC69dHXlsUQ2fEQLh
OJlX/HPzCcK1JpnR8R/9sjpGRQaIofVm7eP8oqVwGc7JubcfrYf7dh+DDHhU
+42wDg53TD25Gxljz1rJzhtWTMB7TT1X9epMpISnrJIzWnOArVZlVk0vWwN7
LaaMgfuuOZsBHBa9Q4ztvr4uNOWI5R43DzuAl68nRt3MUyoS+ndOz2oFucH9
VZzDHjTfoDnet5cwPZD9oAjQMzojTjpWyAphc/tCg1mP/nI9DC0aLnv446jT
1IfCq56+rJwG9SZOAo3yKp9JNbSnxfPiY7Je5lx7rJjyus6Av8vN9j3AY9eE
dEkT4hNi4dD9ynVW//qfuNqPkaQJpDeWIOhSmS0weaJpmq+FUGomgI9FQRVh
Nd85HKRhoJ4fcnbc96Bjg+xH453X/zJolIgdnbyKKXdeve4uwk2VwJqBdObu
vg3gW7XEYn9oq6xj9LVj1w0KpD3SEQrI70Ij4BsR9gmBoJjuBaPdtcXfAJcD
OP1XuxFRP37fFDoCCJF72KQ6NuTQhGK+rTKlJ/9pvIeMHsLpqR/ybEDdLYp6
FElo+//388R8weWHstPedWsaUa+Z263E3PaDLb8gjHetINTJ9NwuWoNga1ck
YbaNpmNUHWNory+VxAqGswz1eEhRLj/rdzJB7Q+xtmPKoewtt4VK3ta9sLeg
U1Ucm1ykHtDUJuOeTM4EpvYwxZKUyRkU93X52hJvN810jkGXo4blQtUsY5ej
ZOzX7OXvdCJ0CG3yGaQCbwt4XsUYXHx3Woz3ImA5nHuS2yKxA0xY19ku7vP4
vAompOiBnKkaOsjVKSzNk905PT8JEa0KsvymALODFfSS6VPNXugbFwzW+BJD
ILNgoU3vnlBIhYlssM9dSLUXnTmC4DceWDdtF/Op36s0pQG7mcLwsFwXAO4Y
wfv78kU3CcJURqkJTbGTWiG/ifCSm4vdpAiWVjpKM9XlK90IWlc6961j+Gnu
maMDFT+fKpKuCXoojbzYOAcZ38wPw47xJB6EuZZ2KQ5Yj9M0je+B+7jL2T/a
ZV+y0UVbHPJqZcCmdp9geSLCHI19tKVwm0dl/faGfUWMqC3DUMDugLisX9M2
aXEwFLJjGILMA9EvKsj4+cvSj/r2ZG5j9mdCASTt87jL1z50tx5eJcdaH4Gg
S2KkmLUL2PdqNvsp21xmRQPb+1cxYTShPpkwbgTBqKKvjDLIEjmSB20/CN1/
Yh+T1lRbfO9iPbre/sE2398sNPTDX980FYjTze9DgTVa7MWE5gPMkA6gS/C8
kx+TgBk7SowuG1voXGwlFh5ic9GuK1Wi8NggIi8bpIcTpDnNj9Y8/BTNyF54
vL4FG4lM4NOg0nvqSCWWymTjVJInJnBiMtqRnJdJVe9/C6EjctfJnuvVLThz
pE9KzHbjRMc+wE0Cf0hwYTFFu+fSbOI5E/9CvjozFE7HDGmVgcuTzzZ9XJK7
oq3XR8GF1dMaRGYbGHtdRoTpmyQ4Q9NKKyd9YsyCylG1fHX6W14vHwm9JqxK
9u4TQ4fYRdjZu1WSbTl5LWdm3VUclEcT0FMeXP/aqoRxtz4QkHYym8MzZjlm
nwLHqjr6AkTrAIPFYGLpjyDzz+wb/8GHcOSYUAFYeLEZCeZCgnXgroU5HPNQ
j6kAOp90BjxTVikOk9pDSbrHLUb3cyj49gPEaiPJf6QUw736PsFI3rTXWaS3
j5vYhtuloMOAJZ2hChtWvYK/CwWYVRv5ZtYX2d9GZJ5iVyG73IMoF7huCu9n
ti+BaihxMrgQQxdByBRupxrvKOt/xJ3TV8nSJsIRGjOZd9DNOoF4dKb6osR6
yag2uDuLHHTYG3t0MNswztBozTVYSoVBvT61kMs8O7Pg2t0Q0lJWzkt234j0
C2DKIcDnXQkz0zrJAx11Q+BaNWmOvwzHeuJim/QSVKbSy5MM5ahQASpzSvsm
b8YeHBAVEbQVYOMp2xXcUada7Rup2ZF1ZZqhvNb6p+sj+kfMJ3Ldov9yuHDm
qxi7tDcEFtjGV/2S87dV/WQledlZd/Geek598hcKCtduK51sdJnzVeGsCdsI
NMQ0PLgp8aySxvAL5kOkeb9p+42bf3eYl+UFsn+5aCfw2qYjqIgjvKTfQ/o5
70FxgcLFPmj2V9wEZ+Q68JaGmpam+vr9WHGFmCNftYBOxuQXJ+3NFcLYI0HP
cFVO3RV9H4cZQxq8wQw3gx3eve2L43z1ocZiGKCOLWJbaQ8me2xmxhAe56pG
FYXPEg6zKR+jMlTONkQvdcdFFpthr4tA0YSCN8XppzMOx30ARPB0waU7zcIa
E8d4otFBkkircjk9GRvfLRpnDo4EO2EwLZz2aOchJx5nF4RxzV3EP3CkY4tj
A9Bx7dqFUZmgUQElI+90FjLDpHhwNWPl+GAq/vdQFaKcVe5Qkt/2DqfG7xS/
Pm2+QFHQFwL6u3DzAp7mgNCM1dejZRJRON+Mi2UbHrNEaHRIb2zkA9xEctVB
dGyxD/pDO+CiG8oGVBFcTM0nuIjWPCu6z3/9oV3ToUwn3K1PGSonvs6J82nG
0tQAcUulbWJmQ5otuesgZPGC8pCxMht+YbgCitH3SSwZRKfdhA1n80wczfd/
giLsXkekOySwsONbfWArD7X8L6pPbu46CFRLsCHSWe6XZxxBjpacl3mkTkw1
BMoTAriYi6yZTbGLoAerbQIOri9MO1RTLLg4twNRUM++8bc6Z0a8dMHaJzQx
vJVHLF4OOBnh1R9cUjMMzRsZPT7ulFC6z24+kMNfpNt7f6UVzDgS5MCnompQ
8pfWz112nq4aDcArJz5n6tmX8RL6h9PwklNgKAGrvqIN4bBnBYqi2Eel/MQX
+gUAfgc2iNWwnD42YFXGxqiDKsmYtJjejngMtK+RSdUGP86zX1dv+f2RjurB
epCiwyqtcxp9syQ9GH9AW3IQ1/Q1hMsNO1J4KdmGosfoZ9Vf4TYkbQujburW
DpPQrHySKSKEbnv+m4NVnbVU7QYovD1/yBThSWAqtEEEbAQGn/P7SxAmPO12
cudLhVxD5aM885uX2kYnSPDVdkofDTBgN71XG3Rl3FoxGLnVj7pT76uTwDU4
oPCxrqcynswL0KY9xHDo4EzSaMqYGhSt8tc/8uP0Ehf0Cx2Bq2kCUFhNFbs9
aOF4ZQkuNrXEogao69bmxtOdGI/qjGSH0Rc/EP1ipZHVIvEl2eVjOrZPeCKL
Jh9GIe/CUFobNIJckupQzRbSijNRWIUjoal+Z0RpVnGjHmmlTVCvOqFU2t1H
yQD+jzSXQ9DWkavtvMSZJ//nKht5fbHCLxqRK15z3JdWq49U74EkH4XUSmLF
WNR487xVBVSFYb15Byo9qagRLxieuLD8FTcaFuURGeQFJUe3t+3Y79/+EzYi
e+ANCPXCRWD4+QPw7uBYpfRN3y8AuqJcOA+3xcBCgDF4KPgUQFqBr56Hlg0/
4p/FK7zUo+Lsmpn74y+0yrTYTT+GgElcT8ohtt3tuicWpAGcq1az2azO3Yqg
3E2GZIPro3cgB5bR/hSJZQeGIwlz1DKsQOuh+rBjdwHiuZNI/EAiTNGPtEUr
UmIeS2+neZgULirhZWbO0Pjc+xCJgRjoO6Q5R87DZMoO59wnB6RzK2tZTx3r
mXpvz6OOjMkwXiCZ9F+8frDEJRoCSq6hEC5kUuzk0NNh7HcBj1z7YuEytq3J
Shp0Ovv0S/IDG93gWftvFIHFovDw2lsAcjtF7AAZgOkWfcTRF5bHLVzRvdsG
wy2DwRtQC0lcSH1Nbv/nK+Nn9SbwHWBdEPeNEMlnL0jYiZXT47AHMNgJHCB4
blmATi15mJD1XDMmb990s1eY3keYmCvd27qTeclq4wYJnbU2YXgeqSvs9mCD
xkf5PXFcGaXyTuNGRFUEu0coX5GttLaywmrND2gep/mMg0dshMzS/mohb4wl
7MMGAQi1se79fy6rmDnEpzVN2xTl5mVYi6D2FTWDeBl2z6tod/kX7wlMsk8/
YATwOzCQ/DahqVeA+X4ftlbnLWne4mFqHnV49lEAk+le1pbl+3MsWMqNIAzZ
+WPhIDWTElsB/n3qJ098T/nVGXHMwJ5RgRiuXXlTMFRJn6TVpGuz/05CSdbr
zcMjIVH3lx/U9lZgGFUwNKGyUcqjJXRStKYBCjrABRSiqbkIB8oio36QhY6X
G/i0ZrcXwErjaGp9fF7sbBSpCyosmcpKs6iry/Q170MgcfRnYMCrMSw09u5f
iF2rgtdE16/mw6UkQYy0TsmxEWYGr6B8LW6wplMe4H4n03QD9IdDWBffL6ib
U+JlS0KL57+oa8yAM228nsELl2e0Wflq9YksGAKr5EIIIFg7DBnIow2OPCn1
Actf+fZqGnlLIIhBA4iUlGm/I5h0tqs+Q+65/MNJ5jolFu8Jb2zFd/+TDYll
CdNWxDrSzd/P1uWa/4esytU0NbKCRY+NzXYMn+5LMoR9pe34q+VJdeAZvR3P
ulnMeyQvhRnczmrjJGIZqeE6Ls8u0osUcqx12nflM3P2GxXS01Ff+evQxXQH
Vmbs3WfdG9olH+11D3Y4eQdZUz+3owCzMXXtH/Ws0Bguzo/JEki0NzEP0MmC
J0Mav4d2I9nEW/yp2ZWoLc94bENtjiAJw/3znJ489YO7doc54G1ZuBVUaT4Q
z4ArkNqPWb8cUDbTKa4+WP5BUaPFAzY7ZruQz3GKLoI7zDdKxZJaydcFax30
F2hc/9BgN/YC33bg+FEwqDy0r1LZjcdze1tmpq7aB+Oac+EaSj8YQNDlxx19
KX0psdoxsbDtSINGEBLGeUTELIBQz55vqHRSIc1dnhJP/rgily2CGOu5YVjX
9iAuKPO4wKvZr7WSrNzTQgZym/vxjlfgX6tedmaVV7sAxngBp00w6B0QLgQV
UQT8AgPW1aQsKyq8OhNesZq4hO+QUwYT4oCvdF0jJAn2WMYr5EAFMKQ4htsu
B+HkXLe7wVktJ22yGgFjoDy+zzeHEKiGa5Zpw3+4Ei1PxXRzUX49FTBc5qaO
vUlIMdmo9qpJqTTorBdeC8pM/JLWJmtja+TnRiCX+Syqenv+0GgKzG2OwtQn
eBknK3v32Xta5MVvMt3S7FCM6NGsoNXhzlnofiWhCpDscKoblcmVHUN9ayFw
MPfwR2wpmwPuXj1H+uB0guFSPst+lN0YpPtq9v1jF4otJA9ImjVqvk9mbpKF
khvXUJ6QU2rm9Tp5chYGpCmvayLquX8DwKPP9jaID8C+7+a/8vYEteK9QaNi
DjG21mJTppSO/8ELYNbSi1K/ACnE1D6Z7p3CYzg7iDHGVa/4kmvRYipJKLBs
Upmv1Fyd7bHbhxq7Alqmul0TYIGORW5MaLXzJui5j58tcxKLZBq+4EJ+sOs9
r5nnAghidwAJKNa80NejgmNcG1X8Qf3+zcYwh70dpmIc2Gpz1tuwSsynbcRr
MG47kBV/rH5fg7Ydmqpv6GTmRu+lZ79ymd7D0AlUwv4dDhuM/pyBA0ntBFSS
vHQYZGbYN3/GNDtwnfWGeUfG9R0vQwkI5vtikOZmcFpX3bMEOWMVIEcHraSL
BegFicH6X6F9ZUdX8kUQYTKonoxoJH15/6CenawGio7XfZ45jvOdDvrDrJWC
KkD4bZwv5+zk0YpH49Pu+SPM3DcPVZldM1JwFXr2XyJXhYyJCuNFDxs/0x1t
pq5CqTRupgS8NfjM0ojTKzLspUFR2PRflgusj5wl2skTCXYPdaLJX0en2ZuO
H/VubkRFcn0+BxGpG0YR6z+1v0HNiZPxsL3RkNfh1caPxyYGWrf5sqZCV0y/
uM4oa0rEdxiPZmPeYw9IJzhht8QowpWfzDeOXCuvkxV9ZE6yFPktrctEn1qf
Lks9YIveotFvaubeK3osG8OzZLvSquCySXLd20vjgEqVGzvTUGie6kEGZG5a
boKJik+OXiA9W4B/BADnzx3xuFr9xHbNZUzpNoz+NHHOUrZ1x0O1hOKK5h08
B6RGTzANL1DQ2H6hSUgLyUDIbgAcUhgzVoh7Rv/ujz0TdprBqPLwb1dAAurC
Cq0TXWhjDd85JrkLoFerg66JVQ7tK+Mz0M83fJ8+/9ymPvK5e5zziAWlBfR7
O50ykCONTDjejgDF4qMjVh0T/sCTwqJ3Wva6BO7YeheMriuLgLgTplOpxtBL
UIyzvfEkb4W+mjOsMYYgZj8ZhOB7/Iec4HRlZxKJdRCsgXux2RUYLqK6cl4h
23QYBN18czglUNXC/VacJ5UXWzceAMCsKLDNqdQmtxsTHXYuuSYypqXYKr7s
F2W66x1GqdPPNgbbLpUSx1h+lcF6vbn/SL5Mxo+40jxPb512zbsWXWIYWbeN
Rbrg/47l9rUIbZ9+O78vHRqJFJd21neSVec3NWPcx2itLBtmuOoRYUEqa4u3
yj2+8ZxKb/Pr3+wTKR3YfpeFzDUrNZq9qfSDtCJxR3ts7naMpAmt1BrNm577
p9YJVuf79b48ogiEyFz42c4WeMTUl+TiQWBKMmnVJgQScKwt4XSuSSa34ZIk
JRHYvdwI8hdvrLR56SsaLdGiTnj0LoJAw5dLtiCs0BE/KP267cuiFcShaqaj
5wO6NX9UlGeODhMteLjZSTof1/0MMrhW49kyAhBCot6jOWg17gnJKLDoG/IU
odklshV0zqMXOrKgO8OxkXNlfVqFGnLhXxh8T5a7Kl0/sE1X3JHyyWYeFVUl
ldL2+02FY4ZR/zCecwwrRR9HuJ+wdCh8V34Dhq4Kj6FIl09rdReI5/3tjbLt
FMxhIlynZeuJU/jMLml7DrUgIA68Vsa+ndcpqo6pntdBY+N/tmEYU4O+OGAM
Aj2WO6beSIBEYvcLVDy91yp11FrIMZTxURodBndAomEAqvTOYW1bPr4txPHy
g8LoXyoD/FCdcbi30PFCIyc4005ujQEeP6lGI1YRIRHjCyfU2hqduMF8hzHZ
GU3tnOOBTevBAsg2XsdYcSjwlEB4xc8k+L7waz9OJVIOwfGRLPxlQqO28YnU
F35hPZvlVQafCU99W0lolfjtdnTlv+kM63lClVPZuLkzgx9UUbtXhhvj4VCQ
pJCVZmpBsat95a+F0Q/Ubrp+FnNaJRr8NmMrpEdhHmIj2CnuMc2uvx/fXpGO
WOCa9JfjBHmsycXlI9zk+QrQGPFnhNflrUfAkCYi8tSAjYnqKV1iaw07N/xW
LWj+oeOhIi8YyzugnhER3y/Md0/b75cQoEGhdGGslBj9hhqMoRHPa7XCFYVF
Ogw9YiYDccawzrVoeW2tGjjzoaqYtKiQ031i4pT30tRmkJTmowRMZMxcWI50
LJFiORFajTkPk1/ymuKLfgq/I4BshHByrFW04j2eRSK+t2qzgS7KFYUGiKpl
4T29mwJbN3iUD07hIw5ce9EvC7YNVrcO2UX6vFJt/kS3gC1UQ+fsQE/V/4EN
vMEeLxZy7dScNKu8eyTrSUcj7SHpY3q42HZCCYCny+Ccq4DLjbvC0A02IeEa
x39982BZ4olXNqgoMRpsmdeEbF5QnIkZPgWhEENzWQUqCtWYctnEAKIQaea7
f6si629LPSOQO8a06iheHhEoosWZzq+mYVpTegNy8otoXmlatthkj+DkSIkA
rXrTIHuxwRFq6VIRSsHgVp6ACCls8RXjhhvkjAFdvQOZtedLuTVhOnrqTqOg
bfKFryoYH9T/iEcTk1KjCElQvEj2jb5YwjE0yXo8Nd5KVHVy0nslwu/kElWn
nZ0yD8/NSfv5C+M2o7hsgh5tEoHOoTxHGwdaqX4YtO018YmouwSrd9kSTuTL
plTXbvbJ+V+JeJkzhiXS0yozZlduiqIWBKIGMeS78HGza1lkkGneK2MnCqk4
ADL+Xw83gxxdr/SirV87KD/UQPfOrKzgTKjzpfRgvhSbDf9NQJxwbV4vyTG8
Ti29ORMPioUBbkBn1AmrOpvZrezFoYtCOKRRvGhZ9aEu8KzINCIKEWrr0ei0
/jotzViSmkNCXYrzapJ+pK8u86fvQEnlZUkAfWw98QA+HXKEocwSv/tKcW/j
4YBfJZEiwJ1YBXZt2FPZoXt8BAgyynjUfPyxZvT9zClUvoYIzaSHC+fCTunB
UbJ9fwqyi1SPhqE1mdsQx7QkxgN+xmF5R59y/qvLE4MtWiOVCWDzPuAa11av
BOebDkxBNd/WirfFye3wcmG7RLnpk9zCNoJVxFZuxefV77zwspVB15qK1gIA
JSBjGMHqh9UEQSVY+XsqP8J6QOmSRr9w/C814CGfbmTeO+EXH23EztVmO2Vu
ZxDijhAI5rA5mESW3fp1HGfNZDNf4ksrVU1n09J+FtqSmOL8Tl9uRwmzFPVD
+1X030BeHHX9TPgSrTz0dnUfdgkiavslVXsea5nNGSVjijIPrgklRN5lcAuH
13jl2iV64AfdDdbu8kIj5rjFMkvEVtwuQ47qdxdvj9rDTXUpqDfxvOxbNCDS
zuEXIiQrSIanXOsdG9aE9FUO06ov4A+cJ/jsOrEcZ4JVOeFYKVYWwcukpQxs
sL719UHxYNRId1TCJJA0kK8v3pog4eTQW7QcIvsw980hsN73q9/mpb/dULrC
l2OsOD1vqBM2UcJKOIfRZM8vRl7rRAsP2ml4i0rkY7Z3E27i1/UBXGEkZY9F
bbhwsK2P9X78noldv7Wj6g5FkezPAzvZCq+KKrwF0sPWzGG2Mhv0ofziwYUT
b64D89OJbcv+MAxZZ9uawTk4kM9uWmZR6PSYAmZXWXwU3vsA1+PmqOTgDWK5
uzIWaB7wzaQsH77nZnxJRfQD1UVhvSZT0yeNNovazjH02tiFrb0WbtR20tBt
9G3q9D0qSzJHCFzAG9pbU4XpjPtwmaPDWMYuXNQPjOffNxO3i+jjzLR891JX
O5wBirUkzqVPbbv/I65QTApY3kXBhQNWdM/Me/eMmIxeI5/EsU4+rx90+Ko6
2+X6TNOHR2tgWf36l1ahCGOCcKCF1/WYmBmEMHSpafzCVG6m5nu0OoHMSSgF
vt1H8GS76NJae72XmHRO3t/fYq2ZoiVbhnqGpB058cn3S1lbo1tCtDr+LfoD
NwDugK8yBUcvAXsymtXaA4ulVXClO+dUW6GQg3K6BX1CFXqOVMrtPF6wCTMs
CmAV/KXhgcS+ZtZHLw4CHkOG2HwaJUhM9iJIcHF1OqA1kWFyysNYhbGymgjB
TEEFq+5MLgv4LqAJvxGvYJFSY8hjdFVV96a90JKJtESESC2iPLnwdZwuNyTt
lvratRWYLU1I6iDLmuixWej566KNKcgALLNmy7dQ5jCvYnNv5AOIT+2ZcWmc
+FMVd6p+heSwj94mYt70FuZesQU6YlF61pn+ey48ahTloHpl042GbDVxg63T
RAyz/8+UkX6yEY7fLY/WTl9lFyUSe9VbBJiXnyHLuChc5Dtbp2X85plaFmbs
b4wxaL5nUe51Zh/zctj8x9KYnh/CqMVemRhY3WRqMC1iD/hIa3ogH09rGOJh
5tmd/ySUApxNpzEBp+DVISW0I5wT0HXenY9OJil7girHUiZIVBnZ+4NdTc4B
TInRdLOllJyCg4evxbxJWgTqEgfDGd6z21NA9OxAIpKaB9sOPN6mx5zpzKSE
oY+hkaKuZIT8MtCXmc9ZW+baT4yDtnr++G7QBsKppemtLJHj8cDjtIBjAnZH
b53dw+cAwJi+xK078zTi8m9bq8b8Mb+aS0Iv0ecHEED7wDEF9FcWzLjAGU+3
n9ghA1O9w27rOkzLJnvVzxgGp5jnFJXKaIgm4/0FijJQT76aGOYhqLnSERQK
/lGWd78ujOdOSHsscAVr/N2fPHU9RYkr+ALfLXSsTLM8SHU3CoBXrbGET1y7
Q44Xr0nvTGu8OBsm18kqlXnTpA720Ei94QG6lvUveR1ZYPln5PgGfyxtjhwj
A8ey1oWOgZgmXQ6vgRpZDKlggAGUsScXZ1sL7DD25oaEL//dzui9/UBfODbL
oISZNJyR51IH7MCk/jWc+pTicwK4nS/kQB7EPTGAVgd9ayyO0HMMx6Y0/Jlv
3rX4qU1KO3w7ocGlGPETC1gJ3qRLbD+QJaP7SOX6VtqyZulI1/xQKZ7+mw/8
AT5Kutr/4zktqGzwK99Ab0mKMaymLGej959iVeMpvcjzBZGKF4Ee5SJmBmsp
FKEAfLlVpayvEufqOzXP3m6DoiRcvAjFIt3Nn2/alIyXnzqGiElw5fDhSPXk
cQk1C2izfvAyO8fuwLL0ubgEQd5nSjkEf3enakJhL++kTM/FZkT+GQK+R99W
ZfADwPWE4lmRUQoXiZ3Q8YOxZgRjRca/V1DYrWykRHZeQJ/CuJqAvdDlE4m3
1EfmEwVycBlkRHhr2+2knGuGdDHjFfehe0F++so48QObSFx0gm4j2p6/GMHa
tBSjPArwDEOo/ImSOuGWGCq7jn+OaMyCd76mWyEVm0T0gCHIpwv4KB7F8FKM
v7cUoE5qDlNqberkQz6p4qJ69T2A0ZeNBuvydptPGDtOBxhI/O7E3spOeCJC
zqfbuj9UygIkdPHoQHQk+klONr5TIAcXDrMp4xI4DaKIGua/d4vtFsOleY5V
7pHo0PFHWmrAMufJy5ZlgPw9aBNE28F3o6XrQwVE7abYEwep3ejK4r3LKR5S
4zWeF35vkzzPi0mfnfYYRPwew1MawjcWfaEQ978b67N5QZRlbgRLn1phcXjj
8tW1jOrF2vPq3IPsCE0wPITfaQH7nlwIeoT6652ANNThBOmsILPDYtE2Lfja
cO3E0Eo4JEdE1gVFGXl6/UwEdTRnh0D9sNKg6UJNtKgKN2cwskDE9Yz0I4RU
ZzivVtfTftjRJBV2yEiliQrhdoQ8az4uZY3SgTkY9QxmQqMv0pHagpggmtNT
IylBfStsNT1wRbhFHqYN2+bpqGQYyu7+Kez83XgbVcX82xNqPHcT3ZyuCj2Z
xNm9U5y0YwajSxx4otjoeq0MszqihpFhAJFWHK77KWx/DV14IKhp7SP9QBLc
I72FwJ7pqEdzsPUYSMJRCYv+GpQ3SjA2lS5wV4JRyhpqRxmpfF2MR9wwpq09
0c9Rq5zkj1802L81gsqryyw3N8PcBSreFSx4SvxNzLsp2lC7NdALSn3tpaeC
NOrxOHqLpcKd6St94onTtA8Az143eVfbdF5DHL5UFO4VVPYt3f3lbfHS90uv
FR99IFdHyhr5YEM3+S0YQSGO2gwsKbNjN3ASFFs8zTcNv0KthrosD8BiEgmK
SP2vm2ggltuzGOCDxKNrb9/L2Xoi0+XpI5OaJjD1JeBraDIJkfmVuFcbR1fH
ddE/kjI729/Xpv6oGGT7j3xD92he/npcRclsV7Dul7ppsdU3t6YPvcOccUgc
R3FVt8tJrLRURVhwvoc+zCDbaDqtVXd9bQ5J0PBTuL0VVmzpgiXiqvOWeaKO
TRg5NX8qdaLfO8u4U8u93LTdH4IbubC7txqpYMQJx47VKsjVtm/M6LZjYpW8
mAYK4x+5bm+OoREITWPO2Pqj7QmRTGFat41aZgF127ChfjG1L51geH5p5eQ8
qHZu7KZVCEc45Vkh8/GFdXLFj2Qsj+pOgB7Btj3FeSApwkKkQ11e7CVsGQ85
5qz9KNuCn3basfbqDHU0ZpG0Lif+0CXtvo/cnSJYKoSfUd44Karjs9r+mdoi
yIrFGy0ywM/4DdyNDNeDNfTaPY8nhMs4gozvDWJKpM1oMNjpOX1kXffBl6+z
hB5O4GeXV0tHigT1ns0QqGXr1aNAeg0zJfROQXyNNxkMUlhIhOkaeYQdmNc5
CyOtUYKWuG3JTzZzrNT98TMJYQ9Pm3ZqQmQqJGOuNZYZDGr7UPXBZWV8WXsY
Ys7pZ3TLEr7bB9AdSw1VagmjNrSVp6e8ALJt3UYOGgYFcy2Yj6uV/hPjTUCj
sYJdlG0/dOENGDoWRY05EUZLPzL8S8f/bT9gs/KWaE3VaS/IUvThoekeklq6
rHTpF4YOzQIIqzlqNHSx/fD/pYDqJvjP3xdrbRS3WI6ttgj5q0dXBLuzFZFi
tv8jpjIa1IHZZW7z4LGrySql0K3aL+RQu3UzTCmwTleaO4VnfSE+pciVqshc
lKozAVechregUz70ut7fgZIsbMPcAB50Tr88dueyArg/UkAuX8KhXLrREXDD
MiNfLsO9b9jfgF/HtkCjKTDt0/gPxkk0BeCqJ5niPi+SFrv6uC49ilpRD0F2
LkQV8Qj5hMduimJO8i/8oGmFnohO5i0oj9FJdTLGgI0K0Nne5CfdLPCbXdvZ
8BkjJQRC7mdJY2tXJDXk41DGdoVF7Wppdgnul+TY5C195bX1K9/onFfG5Mst
0CScjuLdqkuR0jlAyvQwCEJxJSHJA4tW/XM9AiFegF6mgojGroZh+19brigY
PRBB1v9gg8u2vVMaw30yR/GcIIJumwy5mSau41kAZvyyQduUSjGqDRaMAPg/
DonLPayr0A/lXr8/E/5/qTEbO1eK1rUf5Ue11rHqZy5EKVuyWvoQR4v8j5+S
7/K3BajhBVum6SJT2Z5NyIx6DknMxJ17GU2Orwkr20cB7pld7u/pKc5WLdlm
GxuswrF6TpWgTDV7cnDs+hnB+DZpwvG8MYLmGjjXEyvaep30XVJ7QMOoB29R
UxmV1hLXGKZRL0Lc5CRajj5ucKVnE20G+CCeUaPrGbijKyrs+kFuX+8TqIWc
7h/t+O1S23Z81O8Bw+OF1bCxbtVrKZIa3WsWkIsMKG9komD7O3l3lKlKSuKF
UoSi5seswiV9Yk6BDg3/wGoTSgZ8fyJYsgElHLGPzr3SCVkjI0eVLthQw8Nm
SrNtScN3SXnr3Rs5H62SROpecGKRt4m+x98Pc8Pe3pNXUA3tNFe1g6dxRdsH
7OSz/ID7gaXndjp5njDXJ+V4IitQ6B4ZM22PVogwZOXTIPePxxyvGbNaTTo2
Begh9zQmm+tzfoLa6jfiVevVnfbMa1HKYbSeqjlEj3moRq52T0Ry73y7exZJ
Rlfnm8/I16KGRmkH1+Nb2x3fcyw3ABx0qyp6zIM4yeB0LEbyOK55RQNW5t4S
evNfIGF13nAgbI0RgzgAZC/QCVj2AUE4YACa1gTaXPIlwh2GIY4cnlHpPplg
2vIsSgSBSRq/f49a36vCqPEBYNOnuygqxGAHt0+wd+jxrwjuJ4f4fOMzInLu
124gqVnFCJD77+nzcQ7r8CABxyOXdwYIjTXYSVdsLE5hnFaDKETmIUhQazKN
q8L5owdg53XCLc8gKwa2bRHI3xtFjG5SWLhmI4iKLgTKAVcJ7KyUCxZE3ixJ
qcFR8Ov8V303dLhUJBEVAVUhIt0ybAsnbSGxxfsbyDpXvYbSEWSB3S+9RNZO
Asn0tNzrkHROaxcdo6PcKUErPzMG1hid66A5dacMuZgSjT/VCnBuIO2L71Zp
UPHa9KTmkEHHEV04ntQCr6jOWlzFXYA2oC3XuMX4lhE7SSLcXpiUecSt9sDo
PhZcCZ5hNSvBC7dn6+4Qtx14LQQmkkZH/lP4tORnSE9rMmfMcGfzi2dV4e+5
OobcvDnMiZMauQwq+rl3pYLapd0UOPqbmIokj3+EHXjCv5F8d09yWxqT7X+o
zX+0NKsuipEgG/1mQ3rEzp5shNuMjpuF/aM9SEUmMBxYA8f5sk0GFuoQ8OzY
OOsc1hVtcPycO3wP85KS9h1uReqA4vQ4RtG5yraruV/fRcGGOJ7hjXbESENO
XSEx3qaXJga5r8p4uCsbfkGXQ7IiWSOBFdbH35DdWf9LsNzA3uQRU7QUWfzf
7CYyZMjU8KM3kPwjDKYNKBGW0SwB51S77dGJeaYpAQdlx+cKPsX7VMjlvbWx
pNWeptq8XGr0gsEsj2oYqE+Fm2BtCXVL6laqEUZ3m5H98SrQxbunCqM1i/JH
7FN2hES0Sx9/CjC1JbxHWQ1E+S53kmfeBAxaJRqTbjTXd/MbzLZ24Awjj3pC
QeFF/sUVm5xUFDXrxojlSz8cT+pBW3GYkjVJoR4xT3lwJkBIiUYWWKwxK8AK
ZR0Nlv4yRWzdoXCaUCbPt7RpDORya8MST8MpR/b5G98gNjoeFq+qVYx/sQ3Q
6gBT+dICdeWK3kv5n6hbjr8XqiFOtTXjw7PgQEHrmhUgyzP5AUwHEhRwYCRO
AbbrvisvH4wCFXQ+UxWE6ZWXi6I7s8UK5qNPyvQ7ZRZC9sN6WQHRPhH3LZJQ
jQLJXpdc5qiHBEzClV7E/axghhzbnB5+dC5c5q3ANF7mvDxQ5Mj3Qxao13lJ
EJ+BgpzSKQcw43F9OD8W6bsKZ9PIRdz9YaAcCUogji4gSW2eFn+I6U0rjFVo
rFm5fK4mboHiCueq+eAJB50ZGVxnPcBUTa9OQk5NWvYfLnL3Cg/7Dw1IFeMV
pj7dhBc2yaBuolcYg0ScVwH3gIfOXIFs+faSebBRISK+6CMZlZF51Tq9HTQ6
16Uk6tsrlnfG/hdlkInTsjApkw6cRlDqdIck58VrMMPZtTG62x7N2LBiKgks
fd1Fvh8C0PK7Sce42ugSBHd0qytB4d5QdrMlxE0UsCOjoFDWh2h/v9vk1zQe
+erW6ZIOiJ7ZOm79Xnsx+oRQFhL4VDPCCAwQJSZgDfn+RZKR2xeZrC1JYlwk
tJJEGpH+MGLzHu5dhn96sSbZFyV3X/lvwrs8Qf7YotatvP7ZzbCzFcQRo0Tc
9g48FKHbB1ze2qmTH/ZH4SRsLZ8H1dOnKLSYB0VUbgoDV7sK+d5AAra4oOv6
mofDvYvjwdaKSOS4zMlwPBT3Dv+4NPKe7BZzZPZ/0UVTyosf+jqFUKn+VoX/
xDnCxW+uWybh0dG6xAH4AXMTlPPAdDrgsFhmAXx1ToUBf07DSTJsor3V3e4e
hX62n9AHOYkspppGYg+CCk0Onznup6IIdhtO+ikLuwWMBS66g2CJkMWTbvl+
M22yXp4XK00EDLDmC8wzq7Uc1uJmj0iRGNhDNm4chgoKyXjambezSn4BITTX
rozkUSXCJpSeZOVqFTjaz9fjIQeUmvIEW2G88V9MjzWl3nJ5PVjXeD3yb9AF
mRtfdnoPQPwilmCO1SvYNG/J5Nx1MV3ZL/gYZ0SZ0jOGpf5cxyXQJkH2/1KT
axFehlxClD3IhUV0fXHPKDj1yQsk3bdgmOm7kP4wXAKN5aU5L7RbD786V+ZX
7x3mHpyOtBx6P6zbsRZwLv89mgUrfGcZ+4bcSHvC8FY35GbKBrrfoJhMpJig
ED5SRDm6ruhdNHOdgN5YrNXehH8Vwa+DwXhxdCpAs5J7qa/SAIeo8AUmhdf9
V2upE4VTMaFZUYqV2taFZuKSTf9l2iGRzQo9y+GqCq45caVLtd0LHj0ISROE
TecJ1DKucveFx21vPzwTO3rCfNJinqcSHQSGvZkFHZy2E18soF6QZwfI0hfI
o8fQpu63CR46KdTnaxVO00s6CQYbEwVJDY8sQU4CMcSTwxfXHB3ssskw1GWS
Zhzc1GEjj1S47kCp/+IZiPSYq3givUMQKYMtiglBfp/Nm/gOIg4O7XSEmUV3
yNm2v/mhTKL2F2auDyNavQFAEN4g63a31qWpbyohIP9lz/MWg4iSki4H5lYE
yXU0ew8JTjzEFeJiQs5e2Ts3Yh82dhplr15lDPhI2LK+VsYsZfwHVY9RZnYI
4rauvbXwletEkpDpk2+CpJ+3b0tED4GaCQyZz9nzNwamNiZxLm/oHdfsdGEN
dYKkG8yA29XL16LNxKRiwNU2IWVwndemoeeFDtWEZ9Y7MKjvVqU5Mk7LFnj9
D5gM7kwOAJbx8U1uPEiyojT4xiRtTWhaqN+Pc4ZH70Y1k04ZgSdeMzQGYI0Q
uRrTMdZEBwt5YUyWFZvcAX/Vy9M+5RJhfIHdfWodtY4ijlrzfQSsjehR8iB5
nrtEupOqSFsMTcBY3ry9SCVkVMQidDoB4Ex1gPkRIamiV0owrYaScIxL56h1
KJPglpojk2Ua6K7ubSELtsVRTHaxn10RCklZFbJzajg4eaYnLkPUySRI6Non
76KHc30ewEMDQ+CR2ZpqyIeae9BSmP3T/Wyp46DTkLKM1WRCgdCXt4IP0/tz
Kmx3b9wNA9t1CzGeb2PSJ6n3CpHphtLPHopQ698W2DHO2CamNlIcgDzt0a4P
8mSJJlTHxadhU6lp4r6jjLnlgmQa422/jFZqdJJdDx0acUhVasmjXGWh3+ak
Zi/CTdVNfti70BpcUZblnCQ3FHmqqSsAFz2doST7ZOFjhNVubrdkWK7KJCAz
9Bt1k8OWeeKHxUin/p1S49rhnYw6wH9z7Dm/KGNTJMiWsBXKxEp17Xu3UgUG
7AzsLIfSrE0EoI5Jx6Wp/nvRTX9pTvFI7q+vqJD47b0ahQYsIMpcIxf9BMAq
amWNWDfLb87WrtRXHTK1LFUL6Vr2psV2jRHptXgcdqOpOz43AznzSIDu2TsL
2OQOpmZ1ibZCKj51HaOQ0dD5CgHj8i2HqZzeDP8HyD5puqpY888bDoLAnCT+
aj/UhjhAuUyLcYUDPqTDnYdBkUqBOfMNtrEQ3SAFJHczMJViO5z8sopFvPyl
yfP3dUINneevKu1cxEC1Mm5p3ZPRw1O4BfLPcqMBqX1U//EYe3if0PIkSErN
S07QHM6wiqjYzf4YydIe94vhx6/nIDKLoMzOhvwRwNv2sJcn6YtRlQftcJ0R
kQ0cuG7yXiBw7XaIsUQlY2oZB/DAntvKPQuuKKbkCtWViltPPFf0wljfMBtj
6VP39qc2648dBio8cdF8VAVIGBdniyguC3NZ2WExwL4QzzxMRIh3uQudapPQ
o5VYFoZSdP//SMwWhUonmYgVdtZ8zqxvmuB3jFRjMYGN0HH9gmZPNPczQ7FO
IloM0jGygKFF3uxDS2rMVjTY6VdEqfNhCkv75sL94JjP0CrgVNkWt9zFYQFz
WCHihMgSaOxJ0cWF/aKz1uQwHauKhRCBUhl0tkYEv0cnDWllcfJ9PyGzehu3
tGRZUZRLx2G0iQDLgiDgx2aAlhz5oOumSSHrZ0k8dR70kvgg7zrKvXdLXABQ
Agg4yvQ7ATQVikUipw7CGukh0tdfW1nXu4xg+HSKm7B3Ni8XAwoGPHBKMH0d
fO+i9r68UlN/PLSshwD41BlCcNV87LVjbx+RfJ1+zB2/thGofojGr2TPvwox
tuyU0T/sDk84QjmjZWqVcTMBthlMfNccA1AyxGLYFpXkjRvocY+CYrEeHLeZ
nfoBFI2VRQeJaxeQzkp8IM1CtWNSHlWLVagQpcwSZR8+E/3I0qXhCXJH6aAC
5pWpesTzQdsKiuEcDRVx5V+UuWkGNrNzVt/7DCSDmobL5NZ0z0Vgp3plX5BT
NEP9e53/NZRyIL1dKV3BKFW5WzKH4xh1/xHNqpvW/zPOEBkaavygmnZTyUC9
yWmLCgNX/3Izn7VkeYwnygi4JuQZmh82TzEPCgMx/fyVbUUvsVR7pOhNZGJf
ES33uQaH2Zcs87RVnAzEesm/HHHjWK5X93qzc9f2IwbtPbH4xLU/1g27beBY
o+IN9ip4NXdSzHr6EGVAeL7jQMj9TLla4rcodtiJIniNZZUhbQ3WHtvwlkc8
vrqTg1o+hYfJckh6hZqLWyQlNeogZfPB/pAXGkMBVdX1+jUonj/JMEmZ4FkF
kZdUwxzPvFqbYw4GyMs9p3yoNKC124FDoj44l5IYRxcYf42veZmMuOOUreAQ
77fObb4WaCQcxqLNrAPMmI2/gukd+aSkfizhjT9tg977ViybvxpiE6r5YIi1
M8zdML2ztgimRTOSw7J83HmVPzNIJUThwSXqFHQexje5uCO0yhm3jlbOEMyj
90raMXhaM9NvPVIezwvY172Ae147EQ5FCWq8s3QRcORsEQ8iHFPKljfIpBnt
lRt8uMUeZpDEo7TJ2BB2yIIDHa2/oJMYBKBxHHgfhkjMlxXCxI44wXfiM+vh
JjUiNKf8jE7pg8z+rnTb/GW3+IDZ1FwKDdqMyySOZUTJkXMUJyMtl2gemnRV
VvetxVzry2eqZkZt4GebfEuae3DXOe7NQvi7P7sea5fazG1DqZpiwNRGPMOe
6gtMNfXH638ucptEXo5U+9Mp82FcSoSpfooCeQs1KHScxZoWF+iFxqymvfdG
GEeb0++MXIx47N3FI6zQUcA40iwUHTIyN9i4nRjputdITdbsh5oDhTqkWCpG
xoXoFWowjuirJRybqBbFRN/WD4sp+rA7cklrMwZXwLCNQFPK+63q+Q4D22Y9
xBr1P4ifcHlFyanFLfPetC6dLjmYN95HACuClDHc8XezXAqTxm2yG3uDj3oa
GKn4fNuz55CFaGm2HqAoPCDYPJknisqEU6v3oaBnb59VsnqeqBlzE4J/dnWk
kdgO63X0ZGaZU4KAoHZ+9ond6LmliNwp/ct5LHoZnaj/eKfPfIWz/YsfEejl
Nw7Fpc2oQVeexRRuCjwXWuzXtEQgBHnCW25zaXH46vjBXV9qeAq9QcKZ6BVS
1idr2633tT2MOkkWTg7IEooJIp4qpen7y4bFw763MuvGD1V5ShpHBKo5P4Ye
htth+mUiYRX9qVsLOIasKDD5u5d+SU2wNDww3f+XPWLZzX6cNLOlIzswxXhr
5pQ9j3b4SydFZlFzXKKTe7uzz0e9ZnH49BTD4BVp8PfeiHTimaceCttoDhW0
y9Sg3bzQJ7Pk+rM/Ey0f2e+zVCiIJwYp4D+dQJuN5Cr+bP0gdfDf0S9feHOE
qDsPPRzCjzWIYMId1ec3fVa1K0S0qENEJoIrLvGm2Ab3O1w31xoRmefyyAuz
Cjm71GEIOt+p3iwUur7UDe1wuH0hIf1VNvMgyBEHGp6egw9SvSXU0godPxvh
dD7El6UV7MJo1Bxl9uEto5opyjYJNXegyC/9DX/quGKG+mNiNdjmdAqXqHR/
zdvaKURug6Are53eOkC1cGalBRdl0WbQbTFkoSz1AvAFO6otKTEeqE5F3PK3
3ahC/MeKHyMihh5e2TxWEcaMF55865E8lTa+ZAx8ghqm19mkTs2S7fygxZWY
hTmivi6Ma6J6k+jCK4rAOawMC4Dd1w0S9WeWffynpeoXrBHsDaAEChUv/JZV
e4IWyw3ePCmjdDqTedwbxHiYWrhOhMKBz6f3TmjiplkRKebIxdNlHqvVARY9
6/QFI4ZSS/z3p4fuTE1kDlHKFuyH4gQ42+0Z14iEvPbT0gtsIhxBt+VGCW3N
mJ0NTmqxcNZYga3cwjHDwGelrH8bxPwWKZglUALlHqHmekS7Gp3HD+W3Yr5M
AWTEFZT8KhKccMS8YjLYdsJ192vYpgTvErZHU/rs/c3O6mML8NJjtHHWYUiV
heWF0pOnsQzJlFj09A1pXGBNkrSxvbTE2n7qwHQUcgzamr7yBap5EAXzgNT+
9FNOyz8baFfd78v9heZtS1HhRRVsDsErmZGmQ2qOTNr4RGMaOwsePk9rA12P
nkz8owLVwL12100uVFrOOddOxLLu/ClXdn7ebHoqmMpHYBIstfKLAg7naDRl
DtFQoyICuaZeFEB2e24beFoJrHfQ8tPi46lGAAyhv5ccAzsgx0MlCfM4K3Tl
hqcBjCS7nRoYnMA8xNOvIdjAKC/ZJEwihp79OcRs7UfVR6K9jX2xt1UM+/yo
5Y+2gsoD6gdOKVikqTlDp0N9ENgQMbbodlNTh/zbQ4b0fH/zpwofp0Ui7Y8s
vZNwMvOheIh7MX1j+8PX0UGvy2dTnTCXDMESNA3l0K14qXZDfAeDSs1AwqJ7
W5wYE8Y4HBdCFxkBBhyzRJ03Ptu4kPmuY0Iu8Cf0hvENPSKhzOiAhzk7drnJ
p/m08oumzdsZFvd10UHw/ClUJgKZszMEXpoys4EocZQYTJpkuOsJbrWAX5wJ
qhcVVjvON3wuRucJz1CeYB/BizlgsbK7NkFWnEeaRkbkOOSCa12P5il5TkdA
AgfE3i3a52xRQcz0EJvPQFSGf5ydM+c+Fph9Rs07SK9LVrLS952ToCjGAkUn
FHl+EEq/919/6Kzmf1LPCXDcMxkkjoZcZO2llKANDo3OEfGFeskc8nDqn+se
/rEYzuOzDeTBD3qGHMxT3Dh6y3TRZXJwX0Ps/ev9AxmvNJ6T2OWKVJwaIr+2
mKCoizFsKVzZcOXOHnWO9ce5FwbnCJ7vNUgihWDGohmhYCedLDLLpHG50GXQ
DRlema9gb+67I5Y33P9a7Q5Jpm1jMa9kV4vTKBi+WqaTjv+f3LM02eUxmHKl
U+7Z+Oq0JcvYpHZRXj2BcvwTiXdJLRVgKkeRcNHrC4MES4P5qqC0SH9222a4
NPf1J/vw3kZxk0hftUtvXBNyIIkaHtSIfD7HMv4g+vbMFOA5S98x35J697u/
V5yLd9iLhTeqWtg80JEj7kWNubYvvNdHOxpOvNK2r2IMP10Omzohql0uNijZ
wImITiPizLWmg9fpSy4UpaebR3aqQf93MCOgjsQZpMkonwRai6tUnnTRY7s8
jbLaN4VZQVuqeR5ShtjU1p/hHeLr13HhsO/ISdL7GY9UYKNu3+BIX4jZraxd
9nx7GkUafv9+iSFo//ZXhr5zpNd1+4t0w0wp0NxkNlFE9DPqVt0iIj/baw2O
aiRd2S7JqAegJVP5lr8RDkHjERI4Q0bHEjjAF3P6/YcoY8GU8QTlVAnzTWMY
VfOssp4Ut5oJHAPllZhND4oQFEfaEZPwmZ9IrYTHhLhGJkbJ/rtUUK033uDo
EpIds7UE2eEjCjvVCvLlJuS7MDeJ5gFAIZ9ESCz2bK+aXNO65YAKtLDuOXaW
jzc3RnTCvu/pwOfmDBwvNV/xgyMttMLLfsBxhw8k6vQat6UgbefOF+YskzUr
Zt5gYAIyd82brO2eqEv6GQlUKnDWJOJ134yzD1XNzxuAqpdw/6egoJoXb4QY
Tfz6vHDz/xQLwVO1VNTJyQCq4iMdeERNYTCiB9q1CaFPQUUolh6cEhhKC4Do
szCV40mUqNa93VZoB96JF24Y0R+uaVdr/JJcaNPrAr5VZs5/eGs31SdSzMdm
tAjp0LGOgWgB+VP/6/StYV3nG3mUBkfUUgKTPBp95g/H5BEzGPSSqXzOQD6X
9QIaM13MxuPsNrO7lQWSswy/A78ZX9kBosNMJiJB0cMSagrEI7UUZk6XWOMB
Dgr00VTny9BRTQpVfRcoW6zmbRPY4qKOIvA9uQ4ugMYV/HrS/VsH3h6chhG5
hWsfDRqBS59/2jjVtWZSieHqd+GYib5h6KLOpOqkyhECepVvON7/Sqvyq5h8
tZVWzppGJz5SlNE9JS5hh9IH2zc3atFbl69zM/QN8qDw3pY8Kg2wAcMSw+e3
tIySaTqMW46HYaCbA43tGDc8KMIZBQ0iyU0UxAeJnZkNaWIbp0gnvJTc2sq6
egf7Rz5KhqogWyZEpA5YcBKNL81LFB7MtliWNh9Zgim4lgVpsm5Hdd4OK3Rg
i3xUdW4u1DeiSQuYWpax0OtNnHU7QU1DLPsjzHTP35zJ806vrxJiWW4IkBon
T9qSSAIcL575ouwxSA5qtS+XWXylVDxrsGQzaWZ0Xe0X+krdJTrzb+cSDj3a
MJqPL3RZqn+B353SNg1oNPn4jE6iWcdx4Pg5+RtyNTPNucNpG1/YdS6SdYeI
+Gg7QWBSOrheaOtaGXN39Qlpn1GA1uEdV7+ehLyzE8vxwR3/gF5cDuOfsaIT
zdUBwmnDyfjCp5hBLHlTOCl7o8EwG3D+dQjoy7LTAcPReQu9u9AKwpepjPvJ
zGDU3KZDDj/be7JT133xWLKg0M9Myf2F1u8NOdRXDDNmfFH855au1DHD8GyD
JGAhD1DWCgOYDzyVMTEy/S7qJSVCSh/w+kbS94KdHHM8r56xCBrxwXHYjARs
uiT+gUkMbceabyULeMO/7gcSUxTUXqLq5Z8E6M0ZVtlFeNgKIG6yrgnbrrSw
ALbqV9iv9uSdZULUsLnKIPwdX5tQZwA2FwBomJh32Esy6jd6+eaDVv5ZOOnd
LxdW042VuDDe81mN30dQurdpusEgC5lCEdEfyWn9MzHY02qAUiPE13C2WVAv
jduo+x3cjGqeIXrJ3EtiuRtaBnB1u8nhEk3d+Lu1xrDNqM9+Rcw0JIuCG1zG
Tc+6ftmBKGSFfFlsbrNp4X2bzKiGKw3YOepX1ZoqE6G8u5MQkdGl71U2EUUJ
W6pSLjDs42viRmSJqMFX09BuBmaMoeZ8Fd2xTOryVnnjNTN11KNL8jEBCPtQ
LBIv/G/VPawXzSg4e5CWu6lA02dZPWDSYWhw9y+ePUGWCaP0djnBEqRO24Ie
ZhIxcsVW9g9jAp3Pnp8mcOdAjvbhnYmoRubj4hHkAc9HQHo+2b9fuTyesKQG
+E/9GbSjsAevKxG6tn8QrF7Px0T7SEtsgIm7tw1ae3Zhm+8c1ReisIfRcwTZ
UrFgExlgtcUqKIXvMQeXywByKclpCFuOote4H6ndNB2J54gmwh/AVyZT5UpW
PbpcvlDicOoNdWAKUDpx3SLkeSkZmL/w3dthE9Euc1eXUrPq9g91eK4aVEPO
y8uoDPa327Z0KP/MIQd5JT08/eQotEmS3Nlgi/SF7qeZUe2RX3QDVJWKd+Ad
KhF/IHi4mXj4R25mHP2oOIjqB3WcCw3FO8Ntc4tUaoPWfd3q+mxy5sKmdIQo
iitIpeSXYq3kR9SJwF56CUi/9b3Q71t16vyQHmMNYdQg9rJZ5BfzcU+t/q7i
LhVgvRkJzYS5EaKPczVgKVa46VPiRzIOdzTxvBI+bNGfbnpGhK6QLFwCwYP4
LwKono9YMV8e+myIp33ox1RlpOYdMIN/yXIteNLflRYyAD/lZh51yWX3Vu5k
G4WF81J4YwKmp+NPrYGy+zUXVmqG8O/LYcbI1Luz8pffaBIGCjg61KU/T1HM
1J0sDOJOxed0ugYXvJhdIOIxwSW9jXLLx5lp/+t2hyC1pWMzH7gmxWtWPH10
9Y6AlePWHVLwjnQt1FFqZ801DgUZEOPhoXBZZD5lrIzA+K3TIPstu7D/u0IN
zAl24IXufkWh6s+6BWGgK1Og9lRh4qgrbBfb+EfZUH7DSkK7xP9NlSIHsUHD
eISR7FSdWSVxYUqZCaxsvm7XiAcrHUdbAQeVoM5GYRHB5YKFsznSduUatg0W
1czjCrmpUk4mrcJFULY0mxZC8iofxzBDMrUl+iqTCnTJVekiijlOMkHFMnkT
GJtSNbLDDxVLBFJMc/JgDF7BQOkfjGvNr7pR0GE9Rj8W1hqNseWD+33yr314
DQ6vWu0YTsQgv00pa98xSIin8vAvX11g+LCTsHG7BALyDrZGlkFk4+GjYSMa
PHB4ZarQtz2CmtR50an4P2ex715nN7ufhQDBxQY2ldBP76aUJ9MgTeag4IS8
PSm2mS9lkxYLSHqyyAGY9z85TQmjoMQzX75toEtqg2WOafujQn0KTiRUXqma
MPy21uVZia7ZegvV0J/B9BpJwyAAnGnRWb8uEcD+ybthnFTHtWZRaJa6e96W
Gm5/fN6k+OYFu7vyexD5zOc4nwPSjecJlDa3fEfqbxvQDRq5rB5QOlvozev8
7KIw20hLkyGZOrukuHEfOjw2jCInOakX21RuJ0Y/Vj/bQjlfDNhrg/dE/Oe2
+XJ5M5PZS08OU6TKw0oUgNsGI2N3JzleMgUJl8YJmfksyeKSQRX7jBnAXOKh
Ndn1oqPVzt5fpzRWt/+xLyA5NeTZ6QfXeHpbU7A+ivyJETkdGx4ery6TP4FN
UomZs2dIg0z7T2I1Y/l4Rizrgaas00XwAdoe5EhOyJyp7FRFN8yNZ21eyab0
RiPtCpLcrjeSy8P6PRQuTWSRY5zCWcrxZ9sQgFEcJICCR52sQxSwJgufJQvF
DCPB/L2ccaKqgcQHVsiduMkVOCtudQa3UAJCDXrF13+8QcX9k7HjdnJ+Q9bN
Z5x6Qld66coj29mgTNuEjz9wxkSR2ce0aVgUkFlCvgIFerA47eQPllBCSgP5
T1w3L73cm0jylTCZ5vQb3P+u1GbBXWFZXJq6LXwwkuEqYDIV8lCiieyVpF3Q
Jlxc5EMsg5dmDEmvyWMYa67rK4TlogOg0Ff4F+4eJ/psgwySOLtGjdEn1Mx0
rWH73pHAom8TJBA3g1Jm+mGx6Ureqjf/XHQ64ZIrgD7Qt/4+H04vVaDwy21M
Z2YOu0L1qnLdRcIdMJnrzEowPCiji+9GeKOcst3MAThS9t+wmcLrcDkXzuE+
t/JRDVkL4IIN+v57hSoiFqxesINeJ7r10qhqwZFPqoWX3VzmkPrGtFg1ZKms
7hfqtoq/pfXExMhwbtmBiqWZG+UK8GVmsPag/kGbVcnv9skGn+MXJJULjO2U
3ss+5tmD09wSBY82dKWoBQ1zOuIyG3jQpk/+CBcjzbuASRY6Zrfs5zD0fiNj
9Bjky05Y+SvBpVWFdBPUAIravHM1Ns0inY954vbSapHGmdpdfgcYAjpBY7KI
udYMm4aE4pGVAWiC7aHyMzF/Iq1OyeGbbdIwE4aCq6K6/WF6x0hDRhyhk6Hn
WMpyBFG5E9+dypAODjm9FNrEfkcExYHLYG2auVNL3ydN9d6d4jPOkOM+gg/D
LxufwxfkttCGWLrQydW/qbgC2RCDJ6YheKNY7xsAFtUWcL7nEnLkQPp4DX/I
m7qlfrlHSq/y7gdfhjOBrNMymka8i4Da5HU1ycFORaM4vHa/CsjavNQqbXIc
gXXaRdvoUWTycm+w6AkBhZJfuNB2xEMZd+iXEWEjpVUgmE0uQKqU45NOWrTo
zRBKHaAogXb/6IJoYnNofPUvY/4Awu3GR/X0lE220gdypsIXgVXkvVQCuieh
OShTUh5Q9WVWYrTPxNDSO484vzuNfRSVQtPw7algHUNj1w/ssH0oNaT58dHB
MGEVUnPx36KrS+HSnTn0v2sU5QkLKmHHSGeX56ZIkv0YeX4LGqJfBSzLTzwr
VNIZGvLxbiZ4MQL5TwPsHYDwa+D81Z1au7p84Fem57/6e8KgSNZRSyvsFqKj
B5PkNIDxQeC96QQq7J1Kb8ps7ACjpSuZnUkPD4ddiUkmRNmNaMJSFWYpq4aJ
EAWg9sWJx0MGQrjqPHDjWTOboNlQPQiNKizCTQoxfTdeScS0gDbLsqyfxnda
gmG+CeJA7DNYNdBXruuLSmu7H2g+Ox7Pl+WTI/E9rnx1uwiS2A+81reUeO5J
u4i0Y5R5CLz63wO9IMxGT2hBz9K1cIXH193QAvNHoyYYWzO8jE8YztFKnjPn
YVJDPlqwrH+1dQo2DVAKZ1AhCJ5qh3pNIU3akQ6otTq4N9WjUeHEBnFjX5pN
l6h46QMh6kFo4sNO6/FvqBy8VuxJlA6TuxU47O4Hz2XCydB16yIFy9/3PtgS
neClTIquwxf0X7PrXqgolddCzvLsAXP9ta5iVsB2EOoNm+faNLYGnYQBUC5H
+L/dMfg7609CT0o+jfnUea9pC4YN/HWBswVSZe8SczCUHCADJf5RVbVxcrNT
2QzTY2admoJ2LoT20x0kY7134sayxPEkQMJDYMiyJvdrNwesdIigrfnGM0Vh
cf3qPVxBLl9QKI7UqW5HUH7+raJETVxn/rSwBl1dxODSquqPSGjQDNo9GTU0
tihVvLT2+Lols7J6/Q+l6FrPxQKdcKxX9ErXmaZLjfwTqCBGJ8ZTGBolrEiW
YclaybOXBzb138ZR5tbavT87ql7Qj5kMOxwULldJNLxve3t9fNQgA6GqNobu
d4pfYUH/VjtsILg/xBtdRxhA0+knrv2BI0UpE92tAbXUXYtvQgOer3XW6DCt
8Gf6xtZMJSra4piSQ/45FrMFNKkomXwyRJyBO1Xr2sb/sb6afl7tEv5BnGXy
ffPD9EIJX5SICpd3O642xw/7rj6ZoOsMefp2Z5Cj1mIWfa2TVLUFplTOD8hV
LjHBPBDJunCJuhkN/H15Ty7hCcBsxv/MllknwQOHv7hspXSTPjx9j6oBwXy/
PzwkuvIK/KmzE/MUGAY4zURtj5T/N+AdrSsVp5NfULzsFoZ266tUg8tgzBQL
PYseuCc93N7zlOYiCSIGAScOhAp+70smSQ/+BahomDht2LtSNl9V1kurOb/V
qmTwGILBskREZ3OKiciJek05AFH+cr4/Ui44F5nHysl6VHxproFaz9B8mSQT
Il5u/5qJypKDrdCLOAHGC8XLLtr05jddPrWA7TL6vjjIETR6FCkfFjtcBJZ0
9drJ7O4q2sf8U0QxZ3Ad1tQcYpCT31hcF9uL1xwwzWsphQq9U1THNCbqPJ1p
xuTJWoFZ89PgydSkSIHdN+5Kq7s1KvUYMRJm6KgIbvcXhUe7buJzEm7d9pbP
aj9MqEAJnqUG387SNmvheNtS0a44L8nXXsxkshdgOdAmjj5Nzx8kUDTySkX8
Aat/iAbLCDziGIQscyizJ7F69BgG7SQW7EYg5Kj/MR0C96YWIPiZuT8MOQKK
cQPTgnh+lI/cKVQTUGc434OA9FGZNm/YZUXYV5JWT+zYgX+xLHcyG08v2X5m
r/VaXajT22+Q7iftzJMi9QaM4K1nQGkOoMToY9lA+Sr7ZutJEU3QcNSQLZCO
mT3+rZHZZsE5Z4jmCiSqpirH06EL6/kGskH4GM2FoCvT3Ink6INzlf/0ijID
pypzHmu4c/7tH2rRAUhqM2ms12557LlgmVy6MwKOhITLj76l2H7HmYeNCRXw
N7Ue3AoQXrFRLAESPCwsog3CCKDy3vW+Q2IhBzmIyoyeRFotj0PYBZJziR9I
QkDosUibzZOsHgxSodv5uZ5BkDx7C4tUTkbbkiKUUsb0Uvceiy7R8VD1BOqc
sYUCoIW6gJPSeGGQKL5TSNH962sWqNMoeR03/qs7e2jX7uIH083J00Ep1VIN
eKk3ySSPBxA7fEi8Mc8uZv9tBKU2cgYbdqi+Z+OSv1hSt437Q6FwHQPE5URS
une69dhbx89S5nudinBEwtiyELjptagvWf0YD3MzqpoZXtmpe90S/x+wKrD/
LtuK7HTtQ7Rt18PhchrZLy42D9EL/bfvH2SJtDF/q8dNZbJQM0TZGXWxjX23
iutbVDEM6mCGfqi8bCEm+eCX1NcS/VNSNUMwoqKkLP+/rBA3eD+0LOm7a678
b/JK/vt7OhlTkcIkADequJ+tn/B9Vp5YSP/u0ysr/BkSPbM0eNZ9Rorh0hYo
zVb+edzXH5o/lORmS9BhGve1uQL91ARIbH0uEvqYrgf47knQ7EvcVRYNWlpt
fGLfvV/xEZ7rb+YsHMn0jvlPX+GUp8UK+f4rhivnHQlrN+gGIGKJWu5Ytamp
ZZTDc1jH76UALSdXgyM9oCIR/srwbREGRMdmMt1wG/Uu527CKGRhtf4TzvpX
RQ82ZlJC6IAqbigVvvKEtMSqrzQtiw5DXtJ8yfcnd9wz00mEd3nAlDmnhCbx
yzHnHFHZ0y84HcEKbIKvuQe7hQQwVjYV/ur1GKOKcKmcVuaONdIOB6sNeuHl
F5ZuYtT53Ro8/4DL1e+EjMlDQlKI5hJbR9RL2DaiJYgiWSeDbCbWle7/RPpM
4FUJsxDSdgT1RKuX/jOdJe0bLKOLmsK4CpMs0Ytzf1Tdkb3ONiy3ov8Vo3/S
7SrWK6IoO0rNT8SQUaZ555RCLD8iX+UVGa+hT3tN1Gm4Hfep40bvtcP6JdGQ
gy5cV6J12IPrprX2VcKPXyLQLiYLTnrYvF67jQO7d8CS/IiFIWCFqYzEkHwF
S2zlcboG3VKt6w+rrheHVlh8s8vJpqcSYxt3zA/APJtxY8CGRBx2Hkzmp0lK
ekCku/Em5Wb7frs9cH3Iu34ASBQ6FNZX9reQtb3jZ7keLyZerId4Pa3VNrPh
D9F3rk8wuK03QIkocfa8MCQD9tKgzHhGuZJoKRJDbUdBT0a/TT26smmfDHut
iYRqWdUGSUjtox2SDSOFfixyMMo+bxe3AWSkRr9tPyFQFndCm72lZ/NJLqRO
kJCQ8RFGe0Ouqm1/I+yvpnKXyFKnBpIRDduRKTj+a4TnCKNm0lND4YYyvCTW
fComt4TDuRM0mZFxaSZucwS8yq//wAfkN2XaoWpcpKoUg2xyJUQvjf41oaRS
F4NE4w9j5vodeEYLjD23Gk043qcxuVup14SHA6mfnU4jlNtF+Xc0E5TKb3IH
IXA36nejvGrUW55n0us1oEDYxFjPKvynltHnINfP9OmtDXhmPyPaWQipoC+v
itQ4Ug60hdGrqW5xNwmR6U7lq8DjTOIRFrdFODjcXIt5D6M2MpRd92G+7h3I
2tbnA4yDAMspEstG7UZp6Vhl0MTc1GMMC2rVolhZE7ia/qmKPGXmXz8ZeEuP
gKa4xYc+OnqKCrnyJZPG2pxAIOirPVhbSmHPHUjXWWWt2+ZH4nwMA+nmMqON
hhquZ8jIt73CQdVxkovox3pnDB1po77r88GqemA49/ao6yGX5J9MofY+6Tb/
ZVA4TF5wAKpoZsr3S8I/anaLdL+S6JqKbuolDZRIgyf2NalbsEaJe8OJsggB
NhbPGr40W0juBHnm+tAiVauvOaExaOJuRQ+i1pGEUlURP8FqhjxLwODjq7dm
ugJ/l+0l9+Dzt59Oe4uUsTuq233R9VaolSk2knpikxkJsArt0BAVToJduyDR
KUFlxtI6QHtnzNka+S2Tla3WpKt/ocpRkSHuLOiUHB5EolDwWGsnUxVm/sFV
ewgFRaFTOmMmRzvL2Lq2+HuCgxRPkVI25iR5jLp59dR7X1cUGSj3ooyqAJ5t
lO9aSJcDN0N+iH53/Y84mco/vkSYHPrkjdCuFuQQ2OtApuXNsT6RoUfc/cIH
atbtZhMYUl+uFvVy0cC5052gQRp9ZcRJdh5BrQ3hxFrQU6n5Ej/TmM/jW3gm
XNtGmrEfsu3Vq+8C5fllLiVwcbQI+FvmyohW2zlmfhlF9wHlT/2bXXB/vTHM
92velEP+v/3k+WZR0z+QjEezOI8UXtVhTHCFyV+FqYwcguct14o8Dd92Rtnq
NnuzCHaWBGOKVYVgCsR3eYEFtB8I1FOu9wVGiTln6hvz4j/VqxYyMH1Dxjzt
IHKc80LWIrvHMWtGW1yum2nP2PYEyYBPsrJ1hcAJel1qrPWFBIARSulrH7Iq
HpibOmONIiUSm8uZAKuyuboZKRjBKog0d6obA7L9eM0NJjGTHCsT5Yf1JNj1
DDJr5FnKKbPujbvGjGVlUm/SGQ6jJN8eClrYl1Z09y4X18Brh5q9YyE4UDhe
c8oQojp+X1ThxnyingdNU52A91Sh+Z7Zo82bHT4bxJA2g/Fahb2aKW3Dj7BD
8siheZGKk6DdKIxK/7lCLZBDAcKK1KHI9djQncAUBQDwC5Z/SEEUpNzj0pLC
D0Dax766xnl4Co7fc9TimRQReSI6396pE4u8xHxB/LdPzhvaYRrIKR//w8a/
xwDNcW5enQk3kh4nv1gC9IdQ3sMc6+bI+Uqi1ioTKbtIpEtAFiFeVilAQUFE
KZU/Lyek8sEl+zbE66Mp+GCb5gKXc+r/oA/g/Kcy8iKtQDH9I7AHrTh2P7hT
fxaicIr6JyvaKHklw0mwVeSIK2lNCaYnnX/aJAksyenqNeRsB8JjvAoDuFqg
Rdm3TFnMkx9Vil/j8sC/qX6WYm4xzndhgT1QWbXTv9BmsrE7yM6BA6A42+J0
7XX8wfu+S/MoZbxWsBpKiQHU7uuxf0Fu9dJhIzcKuAO1v5oxJlr2JHyXG2PE
xum8ugtdzOY48ypprCQLt0TQx9r744AnC79NM0f774GreXiHe457geYKexBI
PBW1KbJCAkio6+pZQVW1ZPWvqKlELXEkCzmD1W4wtgI81BxEYAjYzrj5IcrU
j904tMBB7kg1d2RB/H5t2LzW6S4CYl53XMIjWoXz+nDEM12XMxhPMWY8Ockx
KZ9A/ofrONM1VIpaibeDiOMqyihIZo0aZHPZBLGk5xatDrco0aTkO8oUPWwC
mXBpZ+iwuhIoX2dLmxBDb8TNDv7lOUlsKYoYTJdRRvTKJ2Mw7j0PPCYw2JXo
chD1VnET7r+SjkYMufXkcdi1jo+M/cXuiYjR6G/zXOKC4jERoaut9GFORyIB
hp0YWwIqrcNDqgA+qzQ9leFABJKwx563DpAuWKYnGP9A9IG+7qj2Am5xGuZX
Fe7pPnglvl56kPoqt9/Hgw/5dxFNF9Cpn/VNTKdsm4gcrdMhh5YeN9nit2Yr
T4u6EpaTnWz2UcxCX6P2QBMzGz2Jq5i0EwuBCKsXzB7lhcR9QK3nV3iQ970b
qX11TTmmVNgV45BFtJegGCVX+81ZbdZwQLIBjsQcDys+FM3tDqUAaCewN/ta
H8TnVKCkaSYXe/wHxQ90NjsY3nLXcT1sEi7XUZW5/0LfQ49Ak64jhXIsKLwC
zGqlH5BSwKf3D6I1C8M9SHrRNhUQ9DryNq7bKg+5q3HCqj42zTRBK1HVWzWF
QGjdg9XuTctDOpBL9SUY/GMIAYOGGuR2KLETt6C6FQArNyyJViBN17/mBrnC
mkIsehKZo4v1HgfuJsNT2mWo9gn7Dy2IYMD0/eo8tHeFOPsDQvIpE0v4xged
lTl4zRu+p2Qd6NEdzZxwK+zM69JD5cigdG5w3KxWR2nQ6IQEfvcJup55vgf4
MI3p1U0fhbxTXNooLTxJanw8lLOTwfJ4aKToxjQxqK8quJTnbsRPlyaH43QQ
oAmCbCHy5fnK+gGQolCNWE+daZ9qmTEzDOIsRIY+t54Ib+r7cBj9HmFbDc3x
dt8KhSoJ+PMPEO8o8EBbE4WUT1UzZrF8CfBm4Ws3auDu5tnakTb4v/CSAEye
XQVwIXp0442aziVtX5vOcmUW/r4nNP69QPNPO09zJhlbVs2UBfcYnCpCpith
niAxygVy9dbgiEmShI9+onXIXbCu8dD6TkXP2jyIIcIzwui3foqCMosBUCuT
G22iI6osevo++ewBTNYR8+A4+oaSQCBmx5vJZzSKgf5y26Mih2iSL/+/enVC
Mbvw+JFxOpiN4TulWIMSppCqPlKt35XaPu5mN6IIlN3CHzTRbuiNI+FbF2lT
s2r3SzY8YU8x/HNTiUvS8Fw3XL3QFZBKXUlgzzOgZXN2cdEbbiccZ4g7NT0D
XyHBteIVduD/fUCOY0Y6PTsWDgmJGOhW0MnWYoJ7Q/zn4uy0rkA0t7drLgAP
RWYeZpjVzcmYxnKRpghiNjGtsnzUdejEBDRwQjHPyd7iCmamEafiP7XXlv0o
Pm0q+/mAoigO6KSNb2r0s37lew1HhcXe8Thm3oyW58J/hqrspCnqoevdI6PP
O3Nsd1CQJXjxJOO+jmNq/gVBlEfwVF06zIMr7rAGjYJA0Zr6GTAg0ZiC1cUz
dXIS7u4eBR7MNvQGg8JUecsxOojYe2aWRYpRLj/NVnNNclSIgM09sLmOQ+Uu
cDECsxwocVsBdPunLU/49mZlaTGniETdBh0YH3dsRQL9J2tUe4ooT9rOAbPA
alemq2wbibGV8XBI+eSR0KXsEyqE6k1KXnCq184meTxlHpZ8+MNI7wFZQ916
wgXHlp9xraKJbOPHvuXYk28gAE2c8S2T78llLYKzGS6mB7fJz7JwVNfaVM8v
mQ3ocINEseOgeR03I7sOhjZiENz9e8zj+vaomTFBSJLRD3AWixCdYAT8UAHl
wqeQo9lLoA0wKOO11ztVYzILeruhsMAbmj+4bggxKk9G/o/rkReXBlVr1qvQ
ZTm/Ne9D5Uy52KstE0tmlcFcBinzh4h5CxcPHG+xB/kUXawPPPqoXWxnn/c7
GViMVyW7Cv0D/jPuKmLzMiI4qS65IP8ANhs40lFr08F8+YT9inS8pcDFLkfo
/poy0p3SbgcFNu4/lBeeZH/dd9U6O3AWAREYLczruNAWGF1zAEEktzd9WPZy
HNRBNSGTsTPBfgR+J3LGatUNJqzCqmgUeZpeTSlQvQ+GCGETH1lVtXmE+zTr
TVwmu+C1G4HF/EDfzGWDYVJi5jwakc9nHOCff7s0OTzDhUi6lloXuaqBw7jM
yU82m4KqpvTnZUdjdGSr9fRpRbIv/ibkp9nAH99FFewfYcY7cK+57bnsvJyV
fPu55uozi0YTcUuEJLnXbIb90/pccYSdNhfX9fKvhsjgoSDVw7mYLoe4mVra
1ujKWfbDxIxwLlUnTsf/FQ1erSlasnSl+0OeWfHIgAhs/1N1NDWbTXlrSpEm
4qzguxyPC1zddnKjMTqsDZaBS9gd5Y2UGJVt3hgeL3L4sDgYRs6eyNQNSy2L
psjJ9x3Pjm+q4aF7EnNk+UdJXWfYgYgG/B4/MZqkL4wTm0SucfCfF0joaCIG
YSjs0yxoW0XhkpHHLt4AtQ3lBijIZ3O1VvWI44eItKG86o/e31k3DzjRfyw4
OaWnC+xulDg1M+gzSzcBPFxiXZDFiKc9WaEmnKPQkX86kB+nziUeMv5d8kzz
DEySZvY3uN3oG5exGLH6Bs6LRuheu7JDjLFu1fj8bpctDd7MJ8wHqspnP88u
8xI1hLBv4Bd35wwS670b8Q7ckXmyU1s0xLtkw1wJfR2HgVHpF816LpVKtfGj
l+nZswhjRQgJFSER21zkeY5WJiJS0blIemWaYJPAaKJwLAkH12JF8Dgxyiwg
5rP+/voapZ1joB8fmmftCJ5Vs00m6JjyzBbKYWfsotU8bPYKhSr6rntFmUut
VotwX6Nd/S06MxsJq96famDQk2SWL14/PukUoVc1Oc/WmUnhcfnMq5ye/NRn
RAGdUOQ2qZKA65p0r+JHUQ5sj+9fX3SfAS1K+UReRzC6dWq/z6Ax5ftJD3pS
ecEs6FVEd/MGkaKhMhDFm9gyDVJEu9abSGxIWaJJO0MR28hqy0I47/jxUnqF
ed5DvEa44mQkG8kZAvLeHmZt7Qp5apa2DP40pJQHgLiRk1aKKLqOK6S3Uweh
vz3Lak+6FAU3Otr/nG+CCOWHSI76mBUSkAP4bsfrFdB3Ar8FvlnGFB6HHJ1Q
94sgR1RWEgcAN9yP//dyMgmafp4BMyB1hSv1wl8b2MoQAHh0BK028S2TrrF1
AdCWz0SBVGALLWyzjVL4X8dlTR8EhY+N+L4fOspU/XY19XX/6byTVUmUe3Ld
JZG37fpmRBRTcFiq78UHBDgLZ4N/oiObAo+SFGjfljdD3CLDxIW9D4VPML59
TAq6dxkD3KZTGRbqF9a0IbTzkMLCekiibYZHL3ROPLqmLlkqFnxaxmvQ0PpR
rry7JLMAQYGFhNi6T5cvLDdyeGLrUQXqScMdPbMQNfqagiTsDqZOD6fpyUJ8
OTiSXSCjfC7cbFX+cUhuye01kniFER/D2rezd+Jfjtym0SJzZp3NC6DGQBCu
DkJh/xuSNTLoXB6kLDXGdO0jLpdPwyiGmldLDay2q63WurhhuvBgHNo3u2mS
QSI4qPvxd3Pi68iEm9AyCj4JuYpGfQ+kpqc+jEyVXBxBLahDvNH/N/9Shfwf
BYJ+rvRKkusXNF3Rzlop3aCpn6ROk2QERwmNv40GzP4Q8+y1VBkZdbLM2I8j
cn7T21Wek98m+lQUe42xIp85fSxNhgVBncBJo99x9B310ygM/3rgPLtPonUY
oq+FPB3gk7G7DKpMQx1gh5eyhDiXCfcqGJP2gJWi/a+yFXgJvoCYlws84ofK
SIrVdBNHWtmdCPPcmkpdqoQ+xMzVXRj/7ERFAsm+X+e8FItRcOZjxKsrP68h
Pn0HQatn+hyiIaYNTOmCm2lU7+YAjmZKnj6Yaw1dgdPH7hpu6RDWGMvcQ43O
98SYHgjiZpa3rIfyFAidOZBeHU3oYL8RGM8GDupxXFqii8QivJQQpkDCNq/5
uzu9kX/7KM2mPmzmnjvWNVgjm+OokHFXfBnALb8rCAtw9uyWEjWSx6GQjmnx
Z/+xTJI5+P5lErqD/S4+boDlz5h9OAxffPI7dQr93THLJwVSMIyRg8fVe88Z
EVIZ7pKXuKCH9ZTNIP6xn9eisR5/HwvRO+PUpWMgaUVt8tOGJOhcXH7KyItR
6ryCRaNd5zU6iCqRmWAXD+ALwIq0jW5d8q2ty0YjPutQy2obI822YnucL6YB
Reh9Mdu4i0+9DsV+9l9y7c1mbhOzv7dbwBqpL29atm5GCRh8mz5LYiD7iZLv
WFwmd9VtRvW+F99/CXrt+RrbeMKw9XPNnc6MocEXF3qN/tm2zWhD2109AEab
7OFJkdhNpH0o/tnOu2ynUFryJ0Odq0O7yluOAGb4WJkt7f7BwsDcqA+P58a6
1HZNJoudi7Rc/7HfQxaZZ9vyzKUdpIYbnlrZPjNoI3+sDkBIPVL0VbvWxJaK
hwsdl/+zNUzBSjEi5bG7A/2SHGywawFwW7ckrFAjzCmrzHns16KzxuUGcIAy
gzxsf+nwOqncul6Ucvnvw6YUxrhc2Ix1TzSZnTx6v7LPtC9zxQ7pL+BlGYi4
inlhPhT8T5lsLKG5Mc1hXdImsSDGPUnVN2vaBZsOfQ4fHKIin6MJCB/1ygC6
ReQGbXqx8jJE9P3CgeX7nu2jlosZ6oilg+Zsh9nonMYJ4bLYQ9uHnyYdHEps
Plvr0pa4bDKK2i6oHpUNVehWikBEThz3R5hStO0/raX2i1/C0X9BF0YtN0en
XrfFptJEDg7O1kvoyh5Gvr+sxXdcA37N3L4wnSspqg1DWesuhP/ofnpcUYEd
pkVfzjc0PeiTidI/vXHCMgWBUhEfz6GyqhfIOvQO1PCr6xI1vJS7pXbXrHE1
17zjm86V8a6trznb2M94H3Et/C90E31kiLjx+io+xJUE6++FQYLpX/YXkBe0
mZ0vhTfuixFP+6keOnbK8RMnDHtoor2qdDT2/Pkf+esxqWmNzoNeC5p7HAzV
+Ez3G8GSyKGZ1E4y3yG8aiC1D6cGTl1ImQ0LKY7cCNP8xVDPSG7c8B8pgYZT
IL4DC71r3tkXs80pke44RhZE6WzItfzc7fdk38vH5ci0+kiK+W6VgWprbLHt
/430wzStjFrgxt78rmo+IziEyaZl4dw0ZwleAJwlfib6w7Se7Nz6bTUOf1lt
Gmhw23ryPnwIVAF7z1N7jsD4YCp10YW8Pz+6SVjz3MpY+r0CI3rdTpFNG1qD
n2tpXS1BjNS+u5tMpLFZoFpODHV7ybcJW4FxbDcv/SEZDokuta85Y88ui0ah
XrO01nlbR4IWiFCJbjSJ1zx5VwbolQdRaCFxYOGJQyYUKqu9VHS/o4DWngR6
DSiFfFbXmB+A1JsOF6TgPCQBpMW1N+qC2Atb9nDjI99DU9t8UPWpFYytGCCx
SJxaEAAhi+ISTNjMUdu5go9K1LLN9mrWVtGHn3raAio+bZfeDLWRXrYEk4hl
9GVd9I9tYMwQDa6N/3HoyFQxgrG4sQm35zgClICAnpQxD521VpM0SW72vzT5
lg9vm0sMTsDFYAP/+TDDy0asCEOyduf6SZqXq/i/q1/mKqM6OYT98PY4bI7S
XZrKN+SNjqkqeXzLzQSp0bOiwYt5f7mt8E7SJf5oppwHfjOrWM5HC45vTl8P
zBwBSsoCXPiQYrrXc++4WqMPfxaLSXhLh+Msc8+B1XgJy2LXW7M3PXq8Dtbc
Je/sn9ZjHvVr5julWig6cELnHQx8zm+5ifACLc4LB5XiB0vaH2NHiVSMPC2i
ZaIYrR4AuGi9M9GLT34aftMYxWmXHBjyLsitHkki951FXVDpUIPMBS6d4cUz
pq/hsaxBUWX7daaqVjonWZQe2SityA67GnsbKJsY4yl+zXxzjxD5/5fQmO+U
ysA4G7/tNReNVStNt61eIRm9RAHbVS51AsyCI2RIs4yfPyzy4TU1Iu25eG8K
Cb7rVwZxbRiBJ9iWw877Z40mpUVrt9/OmtVoeClXuhV0kASQRI6R0GTvUjMW
DUQd2109zOPcL/aOnu6nvUtD8iEXNOFgxm7Xaiysb6i/gXmY8rNxYu8o+7b4
SQdyLBc5o58B69eTO6sdIe5wWhBjXoo8f5iRjeSVHcC8ovZR/Kq0/kcuWc5h
dBuKOS+m6mYVzLUyfAN/ab/A4z8nA5Uq8ZDQPjOaB83gNDOE5vDyRWpr8jwR
ji+nYnMsBIhsTEx6aJgVQXc/Psgqb/6NllO24v5c/++QGmJiPjJRYF6opZcJ
GL6YbR4uwEzVurw1VfxaIw24hq6z6UdLfD+yFXpeE7co+sTlLN6M4OaQZiNS
8WwloFIcbFZwui2egd+Bjs8ZMiVO5lImSzTH5ZOk3tWFob4Y2/T44AF4VlGx
SJLu5T7M5PLLWiI9Rk0AoVci35HHmCo3u1tWPTu2wXeE+6tMoxlS4gf9Z4AF
+j6bpWWQ//TBkAY0J7yMgBue7IBTqFhqEv1vzCS7ry+aSOahembRTPQpvdN5
ndaX0AmGEF7uW8sRsviMnZaWhbK2t4Zhu07Qk5di/Ek6omjOmf5XzpNfXg1V
NbnYklz4x5O3Qn+BmoJHiS/WtIPeUGTxa5vqRF3/jyTuUrAlmfpfqc+GzebI
aCQXo4jeu3o3cwRMBgHkAW4UWUAc8gY/F25J6x4DivL90F/CWmVwbAB4iwbr
28d76ww2cJ4OcBgHW7ULLf+rmKhirp/n+fHtSTqkGrLw1lmM/CeE1aPbshR7
kqxaVtERISzXfzw2WnZAC9s65W8lluNNFw+Xd9abXQA6v143mp+Ofg2Dsida
Vz2AExSrD6fz+SFROPC0bIusA/lmRS26yRzsoAJdAyu3bWGfzwDWdzLdlV73
SB28ry0bwxEwOb5D4ccBBxF5srnRhK2BNppRUNBnlHeNM2yegx0Fmodn4EDX
tDjhrU45t6XvHn9WEvRBRHIh7buOBQbGY0Q+4Rl4WiJ3Safk/7KxO9RLQBX4
v1QckWGjMFiJUIGVMPOwDxFVkfrzD1MYFZuiy96aibvte8hIA47y2fMMLkHw
eJU1NhtAAXdWivywXcHR8359Igw6uT2Ud1fgGZf0rq9PteMbCd18fUVM7xfW
BkxJlV+Uw+V8uwN0Js/30j4syPSos1CWyyYyz4LI/s5A9kzWDY2AWD58Kuzr
e+kxjDRMVB+AzzglEV+ZrpGOQW2bQ2hwO9AwJNKvvN4lQZ/j3eUxyBwzF+ng
Z9xI4g9cp3Yh0G7qizsHiOLF968ErffBIh85DsbaQ1jIz6qrxgDGLtOJeopl
8S62PuI2u+oVVTY0v1ju9asxuk+xn4QVWcMAR668MzT6VuL2VYrYTJOw5K+k
/EsAP3t/IzwqwoUYBiNfG2EKw9GVK/zw+Ny1VPvnTAeqvkzomvNJA2yj3MsV
hpoSksyPvwXDOb20PcgprVRDi4PpqzjB83Tf4az3HRF0YMGzl9pZJklGgipg
5Y/kn5zhpht9zaRI6ZW+0Npu0Bqz/ZIai0/Ds3SVDQLSE5qNmF+q7Sl6vgUZ
Jz3JUm8g5ZKWvSBgnglUKx48iyDB4dZhETyAwahxNGBkhGE+8ujY3xaaMamf
LQJQehbSWFabQWAzovkjggXJP6vQK+NyUzIjesSP4W1rHLOYX3AhaDfZ7SuB
nkqc9rLfWb66C4hKuNJdfA5gxb866pTtvdAcxJbI0VZ5skwiHhlFiGmWAuUL
+Dk5fuwjNWg4Vp00oVcpZAISJx2gVXbO3Xy/wZlIPxW6qLjFbF//HI41wiw2
Bn/Asjmd2FysKcf0NP/1Yi7EJwfVB7ziRlwAILN6Plw6sHvTofnFZ2F3FiR3
QnT67NRLcaJQ4JlPK3t7il9GvMyst5tDoGyo6amq1uijTY0uj1ueXeDbsgnl
ef0xoAlCaYXQfFOD16luzNKCjX52GWrMJSNmdjWXv8S6hQyIxIFp/lT8oBaE
ZwdllJMpUTbF2YgfNlbnNPV9+co6DizqaAJyGXnOhJuxc6srVElUBw1B36rn
QHROaJoVFhBhY+OLjDUIoURj14znnL0CzE1LwDnOOZxpizRXvaFJHTqkAHil
8jmAll5g+TO5cv97SU4a9RaTu0MzVOg/F9727wf/uvvT1IfxktoomzLrqqBN
FW5ik6Kg2+bADd2cm917UyA08Nq+H3uwFpAAVrUPrAQglUz5Ckgb0OJVW+Ob
cDT2+zWF45SpdVGJuaO7GsHWWM+XKnOcPizMuXytoIIWDzDU5ipIP/cuw718
rklZlXAlo8OWnAtXcTSmRMoIz28eie+uZXsSDEp1actp5CYWPrJ5x2qqqnK3
2wGPerjFks7JiK1nlO63zCIg39l3cKeTPqZjdUw/zGQXAv3A1qdw258fmgF7
CPlm8lZbyqJBQwWz43/BnArduU8T9nsd5sula8PQBKE7FKYAw594ewfV2s30
xGhmw1EZ/kSemGbH26BSwImrwo7dXE7L4O+vHPr2DcCrE7CMxvLZz6NLzc20
FKE4VMzEGkzV0awFmXfyI67TkNExGeq8+cBJW/1nmwtfeSDrCBnnX4zrfFZ8
s9e+Cjpw9zs+CfT21fur404GZzlpJuJD6pNb7u5noz58+OtWMSAPZOIyjfKD
1dAfpqEokFpolqrKvKw1EjPyS8m6sG2MeNwRALDV2LOdAOxN9LLhQztjy7fz
TO0KVbdHu1PuuF+xaWqcITlcEhcmypr6aQPqclKgfOXd2A0kx+/UZJBJErHu
H9Xuhh63NXDtzbyYJvLVswaVY6xu6YNYBVUVY9K4dc3RLYjS5AnfzJv0Fcqj
74b9kZuzJgw1fDPRirnoxCFR8nueOZe8grESJSitJ6KzuDE2TVn/EVFdxkH+
nIHG/9bCk/QXpmcAyfUmwmBrTG4MUqgEmcLX0bl3eUYRQmmbGvvonDKLycxg
2kGjg1BXBUfR6wjyZiP18tBOYB1vIjcKh5zn6PtWKmpfaU5SJQVAFMamXh5a
CUZKhLBJ0LR5hyKDIgg71RH3YckiShhEQO3UmCpwm8/Si58xtwRL+nDLT4pd
EtIT5uja4yWpuCeIcmABzeTjS4GyFJXJgGvSywg/L9nnPnG+hr+xY2P/jqSr
48J09zAyEJzwBGgMEhkjP6qJvp514YsRe0tL5s2682L+is5H8BrGFriiy9RR
1kIXGhInmBjtsiNY01fRPXk7kpjw9OGkPAJmdmSqxZvuLzosV59CsO3rwTzy
qoQQZE7z7/Ahyoc6mQTzw95jMSqfPbZeAfiPcEvzCmdXjvEff/dcBrhI9QQT
YmvsTjP/GyAIo39ZKOtR7lzzb2b19vPJL+uZjPaWbwpcSuMBJwSY2BcGqeMO
J3ApvQzDMcnkW3kxzRr5rtjzOnw6BhW/drNHXtgOvs9U/UIhf7vFaTKwth+o
mI00MIgiTuRgrh3oU0/XBsMVTohqp56t51qOyGzznao6LwQOdHuW0JM6k6Fi
/j73+GgImphWDwPMZtvvx8YUa6KpZ2XSGAd/7FOHVV/ezw8FzJqry/rOL0hA
1JZ+9xalsLI6eqUfZ65H3q4CqLt1T6sXnojceRKneCEL6zBJyyA2JMPcI2Bp
8Y+hSQgKvxkOchKYmeDhMo96YJ6qBnw8K+pvMmhmUek/Npuopzw4kUmOAuDt
KB7eHUkUI16swUAIBT+WhwE+m45EgJb5Md7QnqsjI0Y005uOpZtF8RPo2/2c
L3piaMvMg7Leqvuf6jLFHj9A3+oKkPu/k0XiTlD0k8pvuVBiy2Md+Z15f6ua
U7048jAXNBnsS98aPicWfYPIR2I1jOplFCdPs65acdBszLnaMMu2apDvvioe
WRdzk1IIolhMseTgUqI42hkE0KWdqboVEDiVBSjWCFa07ird+VTssIVl7Mlk
IiaFAWoocQO2yQPhO9/RjHhpQIpeKElsktcKnsDsUVCWfCsTFDZGurpfNKSb
W1vZfz9dHvSHBpVxGDBfxfUlmVETG69/P9Qjh7C3VM0QLib83Y+EvbfTZtGO
U1S1/XzKAiv3p8LfrWO0CiApoVHRlWkXwwGa3X9csHDa/U2if14P5MO1mx6W
ULSP60ZvO2/fM/bhWXrl8M/7PqfInRQsjUF5jxK+AAgAsIlj8JGpZ2b58UM6
VXaHD4PaoN3jughlEnwQDR2PfraDRJb/IwR318++7dp1QU4DOEK8EzDuFBJc
+g/bYUVMJ+hoLvNVPlIo236xDTr7Gn5Ueu+0DGrcYj2hd/8M/oBW7EpKPKhj
FfjrWqdI9K41ARRSO9I2/N+yg/hnYk1OKywCMRX1OVuq6aaPV1U5JZWrGT50
zRXYyTz2ELdvttYDqq2zPhYaeQe9Rsun1jwYzP/xkr0zcZFGjOaGOqbdMPhY
xz0+Yh/jXBk5VdyCwwude19WHXZv03nG104gQ87Jf2GmS0R+55oY6FEf98y1
sh5umWre7Vu14enR93cCfRbgK6fPnkaNFvgY2fdtCoh0cDs25lSwbQojA3NA
o0xDARTaTWaXiToQmQTw+DBeSv1c2J1EBY45dLvj/9peM6+rrycjjsYpEoy2
ePd6Sn7sdPrgpba6xNFLCl5tAThFwXkaV5fzkT67HzHrka7Yq1nkHcc470GO
5eaEIrYfSI0Q7xtEK8vWGrN9fmKLHdxB/bmU/nYmnYBZCgG5FipY5V2/CsKS
Gxri3D6V2pU3K/CMZnGQfG4okz/IF0SOkaz8Q7JtNwz0hMvmiwbIr//2YQB5
bIjuvF5yoGxlj2bdjjHORURabAdMSP3nwKrc3T+2Qlc9pf05exbJHyPjOu/7
NZD0KJPnBidAjFRXdCeIs9ojSLq8qh2CvSA42KhbAbzzU3yaqoUEBuRSyE8q
T5DrpsWc8mp+W8CFgEQGZBzMeCYIFlmnCdA9QHik8gb0KbNEi2daqq8qi2LJ
lMpVQ8wDN8b0EzwpLILQW/flWosFr5xXm/7l9W7OJhPAoK2hIev4Yr3B9y31
s1Dfldmfnl1fnSOHnxMksA8EYo31WAzO7zQqt8aFpKq1WwrQf+kZN8b1Klkm
qcbjazPvWW9x88ld1xIFm9zlm1cnCsLEHyjRiPLJCt6Ua+eW9TKrnZzhNEuV
pUa7cBDFrQ45DfJ6uRl1WdoYILOxzVmjm+M1HFbG0sWF7xPqIuKZ3k+VgvTH
wlbWZDrplh1/uopoITS32BYZTCJClZ5MUqhJZ94wo+0q1UDEKY3u7bquH0/o
I+66Tjgz9KPaGj0u1hdBlgYM7zhbrDUi4SWsFplzl6o0oNLhG8vxHU+ZndfK
VtlJAc/GLmdPOJUIW+ddzaxf5fI8qJ94OclSygi8BbZYkWInaCfxXn87yKtH
dlY2sJMnNf5dj1gI+5mfwQpL+eaqLb7WJygkby4pY7sVpAflQXvwTIT+kjgT
kn6HlkEjRxfPajptLQlCSLkin54goGa0tX2dntYmVt1IdRa8CYvMmJ1Qx+AY
4HU78Y43Bbi8bMhu5efgk+ELpGKCJHQw9xTTUeW8POryk/JuKV6WY4dl6XHx
afrFE4FOrlXP6+qS9cseREx2y3n3RVUX5jYI+lD7kfG18R5U9jCK1hRww5KA
mBktOowHxvVHxkZPfq7CAdtKPVg/IPZktTEMp4BvxqdBtxKr95d9n8QcRqIT
sGer0NqELIXe+m+aOR0tgQXyWBB7BGRjUH/UvPkp7m4Gpu85Af3kYP3JHVXg
3Eoj+iQQpJRgJquIUetKE3a8nwFwarO2/4MdS7DEgSKkOnC/XC7Pww4vkMzj
mKqPSne0HGDS37oSECq87pm33jzcIPj/YmZ0M2Se4+XE3kzY2u3W/K9YmhEK
/G8us6KKVcBgLU8yVBVSY6y58xLejtdXcocidgYijCzLgzceWTH4fmecPIbM
tqD2afMHZc681mqXuDNCL8IGTWGDcbhek1S4Qeqgo3/FfzSg5ag5lzkXeMbG
2NinD0s9bivpDSfQDSHlAcszSrtfkZsJRL/EeVmEf81I1OyJlvDD2vXMB9Gv
ih8+xVBc1FBNo3tOxD8+p+EwltdOXEaIXtU53DNxFuNQH0fawbHDMoYoVf8h
vZfIlMztBT6mo7hq83rD2JE8twyGLjjoOnIwvzAuPkk25sT73pCLjDAqfXW9
UKG03hg/po+TAlARBRwH0n1BtZoaK8rM3ROebbbUX+W898UNR1U7Cc8H6PVZ
j3L6sCddaR3ihd+9FIvhpY+5u+QZgPh6lE6nA4S72IBk7u5XZ/WnF6TpeQEA
T+Z/wXLsvrobD+NVwxNCTVOy930Q0oom9eBi3/MD4wvpdL3yreSz218qyaIK
SSg4zaLqz0dB+qXCXjBD31XPnwdb6UZR8/K/iDkG0fFCliWkdpu4m7TUq2M2
exZzfIZpZhfDFIHtOEiMtlghM3NN+DwXLXQzKwsZ1dYgDvG6guJ3G+Kyn6IC
k0pgDltk4/Yu/NyHTJ4Y1CNojOJtuGrNl2MEGAjcUw/1dRytpRqLJL9wxm1u
SSa4yWcrW0pXonnQpOLzKCwVOkSSZFuSEenXJGoyMiDKCnvpk+fEjwUU833X
wk35sIfmHTLhTqZ614h9CMH9MCQqFwxTXH5RBGZc96ug4ZaV1NAsDplxLEFY
FQXQKDboXajnRGjcs5CwaKvmg3d2VTkVmgGVGj7saMn3hsKO021zwSHIFPbY
dbOuspBAWiuLe3OLH+siHxyXCMvFJxvjbyrm7b/uPX6dMIFFc2bATvyKXqzY
uYnXvFkoziygGToUm0dHmz0+Bo4sKNMk7F/84eIzNFRdQ9VNHuG7EaeYHnLj
w7TQ9rp4zR6o9VMlcGqwVMGJR4nUqjbciVG3CP5OfFx1W26RYw557qbdLz+Q
nSC1bAThrT7rZEcdIQ7OEY4t0R5+WZowTz/rRw4lDsmh2iCGjzqPQtVcyFD4
/TbiapaaPKSURC9Vzey1cMZt1fPWd04ouwPyv6sdehk+iGM6X9zighCOVzC6
SQTXJXErQJmFibjaDQ51Bx8Pw8haMi/9R2+fDmRizaTYpycazB0YHdtovOZo
fpbfTFJt2BYU9MUz7OGBXxyGgYBQBCz88m6m+eeUMBHwZSIPtpu0O5rHgHl5
1kynNU/hsy6vuzP5lJUflLKX8lAef6YC1POye1PPp7j69xqszfHTnFhRGIRS
bgGMipX9Bz+Z3SO0/VJFTKQ4GSWnV7Iu8shWoF1qCU9M4G0kpt8KXm8zYsPX
nGs9yjEeiDPBX4PKogrvJZJ0fMX5G9rPY5cU6XQIc8OMwqDfEOoHHYYYnv26
IiWAq+Ckp+P99q1MXcs91ldX0XMzrli3l+OBJm4CmdC5ANDtFCbORxuD1IhE
spZMU2iNSuE+OsraP91wSrOHfX1k70tFvEaq1W3xarO0GvJVWSIyWecPfJKS
h5hXnNHTCuqz0sKg65gBG9Bq/hpxxsIgLVHWHXx8xAqyOdM2Qg3bZk8clZjY
k14OkVCf0P3RewdXzSUEp7MpNxv4UEb+3LmvQP0/F8edj5b7yNsvZDje8ge4
l3W5PjNTwOQS/hFb/dAI77G3CxgJB113TxdFgctm5GMXRUEGrAqCI0PP/PKx
ws+zh5W0fbskJiWrnU3tVwBa4sBtHWBN9ejTxMKf6lUCv4l2KolyDl4svKPT
xhm4QP65USiiNUrf2DHoyL28pM/uDKI0RH7TcOY1m1mcgZQPIp8f94xnNRMv
7ffh2AMiOC32vmjxzxrldJy0NE5klGcZjNWGdrlXn456tlVXlRWantVt0H9v
s64E3oypCDN2gxT2sVVLOjpyVNweRaBPLXnbBkMQVeI6ZKJoPEVQdWqXQVNU
hIwLUp15oE80dUrjKrTlewcbISOsCBTVjAmSbhk2DeZrFbOQIIO2uZKCPaLZ
io3FUOiLaCdvwX3oBHS3s+8OC8r9HmONjHoK5EJk+pPHNDtQwoLwbZ6o0kTR
YCEJRQRbja6A4sxw7CQBP5fg1cmv8yW5RKejeEEtkIscFehp/dfExulxdKMj
v+tSbno9XUvhBwxJve+nb4mVUhEObWAAStemaf5paEHsx5sijIc2XiPKr0Y+
V6Y5fg4zh4DSS9H0BfrhpV15cYKR/64q9lz4bDBQKP9sm7N7ZHDqyQS4K18D
TjUuXrx0Cys5xNIX1Lq1S/ndG+eDziVqETS3oXLDU/7VljuO9vwTqP4l4Nid
OdbxuvK5HTwiPqIiNNtOxLamjUX5Y7aalXR54rGvOW3Cv7u2eMNclDLRyo80
0+QENa3ddOs6fbRggNDUqoCj6xNhqIMbAFsjVeP46Rom245goQ19XKDj3Brs
S0iKWawiWwCtj0rK1CI0Uv32AidXjUfhEedmfKJqQBJ1Hptwa82FJ9G/Fy8Z
Lw2/97o56/nJ1xaE7BX20jNYOkkQ4nkyGZDSK8waZ3nV/9x8zOFU8n62A/OF
i01dp8IGBMAAYXxxiBCyFTDrvGaWmG87E5Nob66sWeZ+o/+94lsHV/UWtVOI
wEcvM2qtjn61+5ntaxwK0EZaGrR7ZBx62bSXOPEykAqXsSF2yGc1V45q2DPx
uXIbjZbArIPJYRIqPdP2SUw1B7CYnbfHIfPtpF7UFsXkGy4J80ZFylmyy6UQ
G8HKPFwDsbNhB8dFPSrnK6xOue2kVQ14mO+EHQlot7jH7cyXCXrX0ITzuj7B
g8a7K6ewLjtqDTvk6Vegb30tLPT4KIahrlwp6/uwe96mJeeQK4n9jn727q2G
2TThTzkLY7vlZCh27SUK0fA5kt5pfunb1aGjQ0pD/28pVoJ3gk1kecCqIkO1
gHaXMb8mi6o0h6/MWXmqyCla1950Ej3mYJVLULrugvGXD9Pp6++spnqCdaQ3
vS4ryV0lt7Jp4o4UuMUR3zSO87Y+nk1c1dJEK0pc3X1Ewh8BM8uSDuT6Sr05
4wGnKMAuf6Z24InneeKz4uFsAsONspOcpvdgPGtSZ+jCcFGVhka70iZpicLQ
oTQC5OXRDqF3K1qknaBwUi9vPQShChr88+fitvF/tJmJg8A0hIkLLklMnLvL
BeRWCT5bbv7u/y42iSMMYfBVVsE/dXjdDfdmo9q+BsbBlarD30MYPqBN+MJ6
dn6cKaTQlwSYYxgQpFLXL9UZmZId54yQXITGzZi+lqHLgFc8mYmfmCypDzW3
Z0j5HLL2TUc/2HobSm7dqqCnF+6Nsav6bZIkfFFjbrcfLpeGl2GMNR8xqwwg
p+RtohBAIBa0WbptshKNJQ42q3i3SV2LEN2Jded+0aQ0j/IUPOrXK1gWZOuU
4ULFt928erHgGfD94gqEOrX5mtoyp0TNb8nTEn34IxHl7RheO1q8x8Zfz74g
OIUuk+2RUApz0F5oFPaiJKvjmHhmc7joySs5+jgW1VUQC1jSEPJjzOwJ1H3A
HoT+QuRK2MzA5zC7yayAXHyH15F6G/joQSqVOEeYAdcnMW/zdBZXssTWyikP
S7D+9pSnqxAChGgDdFfvAIyXHLREM6NEjIa1klyjzTWT32x6Tr6nineakftO
4YnfL4cLqRIV72AcSNFGF4suJZBkJU/mczeJTDUUaQZsyxMfJ+d9kRnarZ2K
gtxipOERGMD2mRVVOTfg5KNLwjqDdnrQ6y+3/tv/2CBqzIsuCwmSePhyNDdI
klpdOF5RN4MjmLzMRjjEKNYsjrG2gSa5oX8pI4/nVIpp8HqKaI/dDL8J475g
rFvrGd9EkHcvY9Ysap3HbgnmM4ZlUrRbX2Q6azb6zw4bfLH0gXb117Ct64q7
HO50FDP84Rtw+fvLmSLUKlRNO7Yvgxrcs8C9nk3ozDvdH6apgJwwnNOsTzLE
U7iQ1dgRe4AmCVX5KaWneUJua2t/oq/ZZ976NDM43W9NYTuzWT3+B0ZEGA/p
P14lVhuTZW+19bF7KGq5Lk5xCsSiLH8ZFeZe9SX7IYB1iDDhwAs9u/pYlWRw
U6zxkp1+kogY8mpbpFT6bcKLnBJ8RVEeCvHYfJEGOOEbA2EqUEeMlSsTxoN+
hm55+Uv9+awEsXZwDOEpqRJMzkO+d56a0337yZYbUVj8dwonNZcZMpfv+h+e
2B2VsB6/74+qkZ6xRUv8I5tRt3PqbLcnvGbDCbE86sWSmkePXqmd2i1YzuTB
pFt53F2iRZz7xily6E/0JU46IqkoHULGcrwu2FpdUYQQ0PVpSCRv+Ry1/swU
PsNR1HTjZ3ws81QHpLhnR7Ij2Mp5A4cgTy0IaC1Kv6cO3wOa3Z10tKejCOw2
D0gft0PYvJyT6qb9V4EYXC3yLmXRJEZojQNWLQDpfpxXeOjBJkI84WsrNB+B
l96HqOboxUv+wF8t9IVPaoQuAUERxfvUcs6Qw+vPTVOqsSWe5NHOKj/jBSfd
VbBnDloowLbShbJIbmnJvPut7dQHTC44hR9Ybfbj60vqAbKNLdJJiFXUX0yg
VVc0v8umYR4r6FjNwTQBP3hpzUXd0W4mF5DVypuXVVR22PgP4u/PAO3+C60N
h3X4GDAo50hsJSRijoiN78F0elNa3Zih1DrwcI9BSLrW/NTo2FWaeVDZf5+Q
9osw87yWgiISs2R4j6F6Tef9kVjl7liPTooPJYrFzeDnAgt8e+gb9wrz0dCr
eowEhUSo6wx9ExSPqJaxx8EQvixMLgrKmkzjbrc599JJA0iPKkHqvzsuD1/U
Uc3jRKGlOEuRBcwUEPLlkM+4DGHhpCXGrISuOBu/c1+2xPTWiA0IiwCTbQ/a
fBmr8PSuTVoyhyLYBVfQMo7fiADCHUA7bJ+sG3TSuzOzyvgimLz9QuFVO/8+
NzfPUxyzxboaGx4baLu7hbsYfg/3r3L68RAdqJlapWNp09UZf+1/QmYlV9nb
pDnVJMapThoalVwv9OD55saHgPcUZ5Nn1HkxCE5Y1whalsVyrfbEXMzsZ8Uf
WM2wSKSQGVClnEfAOZP9yF+KZUA4SN7ZKKTUizIsznq91BcReHkA33QyOTqo
eVe2Dwlftrr17HaNtG6u+UNtQ10r1doBXJ4sBcGX70D5R+HoUf9vDfKMqBdj
a/2u/UG6q9M4hwhKdEtV9RLo5fyqPQCs7s/AH+drbAu/Sg6LjYiZtWUhv8II
22D8sxMqz5HW9981KvfA17hh2Vle4fVhQyD2Ax54147M+atrFYK8wEvZHiuW
jAWRDrW/UNFpXzvs8tn4exQqZ0jiF6Vzj0ECKx8dyzaoF4h0O1wckWOQtewW
7tXQMRKRz981Qme+Q1wbOhhC4ruvik8fPdArxh82RWbSKPWw9Ku1srmMJbIv
BMttMcMaECPcLEy/4EfOJH7xxkWtAunyCkYf5LxxxWuTaFa7rxl2LAyMJjw+
Kdm2+uhRSMpX0F7WOjonEzP830BeQUX+SkS/36N4p3WubHnqBhhl27Nwlenp
jKcbACwlyLw1Uy+n6qLAWfIX0ikWh01/Wv4kMaecEHnp+qCpRmyTybXH4x+Y
e6T4XG7eV1ATQyE+IHdqaKzNkzU+iBo3crouioE6nIbDSPr6UJhbm6+sdyqE
zsL/SoPyOVDZ4vfHvvmy9A7A/5JjGvP5SRPojc/2XA6ScieCxuc/fFMy9P2B
yNUrsbA8OGeM1hoqj97b6oYi1FSRFTkRSLVAAKPFjgkZXjBr+2wPH9bGCelq
oE6tmRFHQWGDdOyL6b/QjLbUmMATiIdxAZINKI4W7mtMbFR6bMxWZK6s0LpB
TWQcx21mf65rSBpQELXTKV04Hi4BNoQQrlfN9M0PhC5oyEcPTk5KIY1iJ8H4
DdpIfjjQpY2VfbgSi9zznb2zX/ThYQSSLAuxPMr+6Pz6Clj9Ssk6Dg8FkJw3
fDif6z3CeZPYCoexqfPdX9FJrcHbOmGkyn8H6emg48q4GKoBpUd+nTaLlS85
T5pUq7Gy+I2NhMePqW3fVMlmvEcBokXa7KsETXztrWEiZ1chNAHHz7tlpY0O
iAahZX/R4O2U9C7stTeFp67O2/N4E8tX+UEMZh0qHv1Gd9b4yGOLvediaVlv
ju4j/YOEeR3mTRtyIfM7YfbQYPWD6RQUgf97CdufB/yV8tayEnswBqVwcU2Q
nfUuXOyO/f5l8aEbJ8sMPtg0k1m8UhJ+Mlm31BN616Ndv5s8wNKQCxZMRDsC
kh+GrcHWOk5/Q8QVAxJ98cmn6skLYWGKcJvuPYLZxJGyBtKkFA/nY4uNyL6+
496SUT/kvPHf8gxe9AnK3nQdZitUb75idIB3+j7/VVFcphFeicScVSnfi+Lo
tAll9ldRD9DB50jmtkSJdMN5Kr1hSzDXWyo9BO6RmITaoVQPERD+XXQ0FAJ7
4IbFdgs8pudHDUVvAJ4RXt5Wq/9a2qKTYlwjEwOWm/1hqyg+x7j3bGZeV/kK
7vOZxb963AK4hTWDQ55eay8t4FSlgpN9dSum3bl/wG1zIk0vBUD9TCV4fa5O
7FYZNmWM4QCAtvk/HbYzOaBdwm6qgsk+Ubc/0w5haypIDDAaJtUF3WxaXZvX
fI9Vpv6rJfQELHo3gwG3cJY+DvA1YUCJ0xSnmf3qQ0lsxutcVwLvm0OVOTZ5
4XSNGsXbcH8UtJMWKoWIwEpeFlP35XacSPf38BJPSImtLOzFF5TrfbgpnLMz
orGdMTTaT2QkB1iyJJY9ZGh3tP8pZhNzE07mbLVQdtP0D4EZPTGuz0mwVajF
SnDBVmJEDE6DiveyIXU5PdJ7+9z39WaiYoLG+57jHnE04OM6FL4T0H0N4+Zi
CLSW3wuRYmBLQHcd5w1nQZVnto491Vcj233VHCI8HYloPqt+UEkRp81ixtHC
hQ8uTjyezzeF/gEjQx1ns1qTNt2QL0ZhaEOieuHH+SXc1PWipAXupgJZC77e
ysRpXLT7fh1DjoCxav6Khc8dGUGYrClxra1OM6iNmi05zr4OqLCqxe4hF8rH
qwKKx2fnKhFJiBcVZPAzKCkYkqLt55hmZrz59FdmA3C29diZGyupPnCdyqzI
fe7gauTD4qCd5E0nu5o08qrGH/zR3FwlEEJ2oU+sUsSMRu5u5I3AfGtfSBCb
Vkc/MOZC8nfY0BV4lDc5j75gEb4301Ziyn/EXgPOJ/ShQ8wLZq3sPNzW4dJN
Be+QF4Hq8s8wVc7vQ5zTB62KlctNscIeoBHXV4li1JuvIxx4N11CXu3oZjY9
tDe2vClbDywNW0gSllFQIGG+YAJhzQwGf+8VgiJ+xf0JbXY9c3ndPRlYnfNy
eeOSpKdttg3vWqMUx9NSJsviiu99MfQkUV36W/8fC7UmL1mn5FHaZoJ1FwMH
ewwV77IDD2A8vm6W/3t47O5c6ULDklt4Cn+bBYzpDO/+ty17QWrzSfD0sQ5A
060Lndl2WJurFAbO06l/xhubPxj9CvPfUiRnebqZvAT2Ldc73NYkxGndanaB
MafMZGbZQsKFy+ljGSACxPuv2BTMLtI/H6dZY+nnjNPr9u5SJel7aAR270Ot
/7ntwtatHq3ycwdH22K/Hs6b4x0yCwBWmJEPQOnZdJhom0DXsvOExa/ksWCM
CJuUrPJG+/pj0eW8HKOAq55w/lFUj2n9M5SG5kj40Vw2S+1Fo+DwgxBzl6f0
DW67nlJwvRBtKBHt/RI68kpqy/QzNRtbC78VN5Vdr+3XdXv0nJeglZB5ebaR
c0bUMLn4mOt1pn3x6y/afBSjLDioxMubPvt1zOB8WxSqNoXFNgdUfkBbEngH
cfD4vNHg2lI6C1GKFS++8fvhUAEs+nPbD1XvCZSnHsFaU5PSlL8b0sybtuJ0
zdHKJBbf2KLEjHoOyWRhes9pYT7aqz4gPNwmEJTxyNHUumHsGWtHkVpJL9Ob
/xUNz3lA0IPnEg/NYX+NJ0PbAj8LslFv59WpBROpSFr+sIFJfEPlSUO0sZoD
/52hnkt3NcRU/2VxwVOt15g9c8pYhcd+i9bwQzbjYtnybXDZWN0H8M1wJOAr
4Uo/aj8p67lmJWAncWRzpStxGdrqTZGmaGF0B90X7XlTLdIVrdOJpZjyIXsb
sXK7rzlbKlIuQcLVnhWPwYG3u8BRC+ayHU93BrzISjBh9c4cmCMHFjS/xERf
AhcKT+6YYNxlLy119shZ4NLw4EuPgW4sRHhxseAGcPErzqAMHNsN3NL0Xt1B
BHETKKkjNuKDzEJHoo42kzqpdRsi97PFCaUh5z/E6OCXcMG4i0WWnYgznTWn
lLimAJlBEjcdNEamEPVRjr+V3UupQ/JSgZXLM82WrIJvHqkOHur3OeFhGcmS
39Ra1jKV46axzEY/UHARsJOw3X/O68WQHPjVoqlPVeJn2J5KYVs4y0snSK1G
sKEO3NyYztQcD9hfyOaYvDMqTyAUMjCgO9aM+8yDUtuYotzY5AWlOjAkR8EJ
L4slLcKbxlxjbZVTAM3Lo2GuZ5Hh7r0JPLyxF7q9oKfHhzQXd/rpN2QWupP2
zUzsaigAs2XlYQoywR377u3AR5MMA8WVtleMrR5uqVQ8AGXBwhXJNRQoabX1
Dpzio+9QiAOYxS0xpxOhNQ+3mEc9LZSXGiExqqB+7asCfLSyihXpSCG6Zaxv
q7y65FXwxQ7AjxIz4GlPAigdTCF64g1OiImQ5FHkaMCvcp8M0ggXBxdSVRHT
rbkXcOBaR8NvTfNWXNoCBrF5iZBMY1ygofhaIvYInbSZ1uFtR+1hUzETYznh
VqQW7D8yp7lVWoXTzwNDymO0asBTVeDehVGYCG5B9EN+sIBzYZ5DtHogIehR
JLQ9yFQuXkb/Mt26etF5ctfMC4qDVfOJVhYyxR1jU/eHVU3Yi0nX6B/WDRH2
0/Z/cmvCqhrq2Mx3Y4/4M1gRUWNqH9yNCy592n2xsdCX3N+SwvRQScNy8FjV
OTBMrzBquEt5WWN7yGfdG/VyLNKlFUOUkopOo28EqtMHvO5lEtiMbM81E0DD
WlXkBCsIwxgIJwmOXc2snCOt7mFANEFJ6NpmEhPrGwJ1dhm+k7pzWxfdP9YU
cuASWFfLackOvzlwoqvvsJoRIJyN1i7tBDi340TX3DI1L8ZX6RfM8cZx1+Ue
BWJ3oHBAQQ7BwYP7/zt0nfzbOcN7oIJEz5tIhY4idJRsxiDDbDBUTZN9IwW8
2ZFDMpBPRr6WlpIY5YYYjerYvQxB7kI/kIEpDY+bMIztR41AKjCCauyitDku
vLM/IJ+OQtXCHlz5zMrP64W5r38lYFpEPo7zTNPue5iYacpCzdGXBmJ+oCHx
hjlafFVj08zAfbZ1OKfqptrDbyuK3QvMl5GAMc7apDa4ErvH88hRDXKGOrRa
onV+/bkwaVZglE6rJ05yUu9Y5sWRlt6HwdNqcOX+seC3D8an5Y+bNn8GpE0Z
b7DbHuWMqLHQd+h0CMTY9VNvNDVveawwlSZAhp2XDsfAAZxAv7LjybTg/iNf
TQQMl6XK7YjbBV4u6pxlgm2LNMf9MLQ/QvomDcBx6p5XcP7vgeuM8fLo+MqR
/LdjzLtJxH19ypx/Tu00zwcrb4AFwDlkIbIHKrQaV7sZTGCLrC8MeX0txTUs
3inqZPAg3F2trLA+OnOvt7UvgtvseQ0pSZZI4+RJKJcawTUm7me4dmkD+EtG
8ayBvz8ljjps441Qyd/u9x5AZEPX7N8DHMQbf6ycIVhSAPC/Kv/m2WEOq7C5
JAca4evBWw5ZOX1lqaPtuTSx4fec9UgZ2nAXsCUHHVmBjd3Bkaf6FSycSEF0
DWXtroWeZzvFAY4eathaP3JhmCeJ38DdyEHnvskmGoLM8VpxDGcq3RbbP54X
x6Ah3oZix8zeD6yZhTOHBRItHjhWKcU1bmMlYxmFujc/qVJeJZP0vGmMXhAl
tHmiH1m6HOPUsoMb7Zi9D6AAOubkwcExHRfRUZ5ctDJBuYeOUWXut6gmoBvR
kFRVbORByhXe1MmD0SpDQB7+GtrSRYGkCZ6gMeZdjNs+iYDuwdR0P1ZbKaq3
cmB4pMMUhY3mcOry+kZePVicHZnKaVgom8Wxd/YQ16jf1zB1PE3jgLTW9/u8
2H18C4irzhbHmqbsOEu/0u4sh2YC9d1Lk5J/6SXO6MZ7oz5Pw2mOuIE/01Du
g9Z2woMMmfbncpwVWfkvtiTS3kACG3O/UG1lSFLaWCeROn4vquiTVnpywWfX
dPeOfmHpEwenJSUF+6zC8IuuWsO6DQZ2YqMpdStnQjk0RhwZtJWohR5MrflB
lF5V4TXZAOQBGQiGFS99vYGmxdNmdKNTmZvyerxCx6nK+SiFP6y9/ej3xb3U
aSC4mJxkwtqvDaAfepT3iHraJglE+mon4cDX/o2XcjKN6/4cOmg3Zi+j9+3k
wAzEHe5PI6D31tFgW6G2F08wIwzeH390R7xf+FbLAx2AHx+JXP8IR5+RVObe
FhPVsBaKdIUZfzExMc6z74k8ZnRknUIE2p74VouaNfRdTgXoG1UYWBHDslRx
KEMcZAp6qz/3B00j+E4fQqyaPD0EGzuZwI50LD/2286qAS15LaAD1HV+eeak
yrmiLtiwwfB6B5DLFA3spKXlVfteerlKgnizowYXHuyCUlHTBB5w5WXKipWw
trCdcTHhVJ/bmul1kxutv1FR0nsijoNi0GTKe4xPWjgds0ab3Sg4YQiMEsQO
ugyVgCrX6VbO76fRbj1r2KCjlOUt/kmT76t9fpgA+AdlY4jjQbO/f3YiU6iH
1kLK1v/Ec6ELlsmIAY2RlcTEaUq47003+U8jcgFcw7E2CfyWeVdhO1OvBHL8
8iSNhpiSQOAzk54t75HUvoNIt6DAt7FRv2aEsdfC+57O69MSBZWggJW/4S//
+JnhpOwOWBlgBEp9mxEyeDnG9qzcfxp2HUVIutvNvTzm5ApuWvz/wzUM6roS
S5gP2+IplxbRR38w3Z4dsxXQyQqSRrkK7F0j4wgTs0JNL9lNIKZDDuXxsLBV
P8rgNFfOFZ7oax3L9rUoU5A0B/K8Ml+eNtS3Z/m7ECuBpRqeoBST2eHlooOw
seqpb89+T/kCx2LMbm9/aD8uEp0aCOp/9GRJEQg5IsBk945pOYvdu13zYsKV
Wu5XCDblrYhNF3UdQINKHBibU2t21f4/LT24mpoMnhVHcKpZfNfK/IavD5sy
tUBbjk6U0/qNRjjIuuyF65bAf0vlBkp/CR/87ws1R6aAKXd1aFFoFPEv7+pP
3bTD9+rQJng9rExzExNlcIfplslrODO4agLnUckPp8itmjEWC53ZZNBIXNhO
OVFsdEfQD2ymW1TefSTrtAo1aZxkqFdv9TW/iSBm7ycMW4bt89hGDcQId29w
/XBCqs6MARyZ5kl5D5KOlb1Vy/STB9ibKOLEU8+So7kVNnO9KvYcDcc4FSMv
diwefrjeGm7AyDN7vFRutXOjWDIviTzq0fgcxPsM0WKORQKC51kUvwWgeYnI
a/yfqgjz7Zs9bjkW0XTWH9nsQoTGJH6ox6B9DkDpTob9vGDDUzLW/hQ8o6O6
lOj8q2X7L+ElydpZlOz0IcwHXTUHPT3dRQ0F9AyldcoNk056ADAymZv011v/
aA6CZbSi91iEAjwig+04QTG6blexxd9ZtqTSD44DVJ22hhqaJJbFW0Ruynqa
DyMNxmd3kQKCpT2pscw+9+mwm6Z+RNL87O4MJmBDVrQfzZxBVLTbsH4J2+yH
mX4RJ16apTOdwMcGf/1XjMNXWL1TAZE9Vbz0PVQAniFAahGX9/+8yiZmf/1j
T2rL/aTo4IcPFquWuUtKcxBKXN2IujZ6Fn1bXZwleXNQ0sb49a/OOxBjLzy6
gQPPsUAizy5ZV6RiSeFw5r30EBRdJXx3y4QNsn/xCEcXJ6vELcPPUpbmo5Tj
s1RfYZs6lybS9/p8HvuU+g2janqhwIb/p7IW+oFsUoung3jIxxiYu9E91tJZ
1rQAb5xW2DUje1rsecjLru+f2aNA4I3FBVEOKzg6huOPebsSz758wq0wM2+F
SrUYe0SaKCvN2dI4XbULbuGxTJw4FP0srpCEbZDTVnLLL68r6huV5ecgsd/R
6xzIhBR7ZdSGR6DekbrdM1S9jQm8tW29+N4LH0gHUEmbbtxm361OYF9/TOQT
CNRr4aY88+2G4A5MdahoWtlvgJr7meAf/EgeNe12DThB0StdEt4T4MN4VFzR
jUUY8V4mFYY3SSFScW4ZLOc1871wupM5Q0Cc0frSkmdvC5ZRJIpAKU6AJT8y
Pn55+CWZ/4HlIkQCyaXE3rojEVpLgxNtqjCWd304L6zMHSpzafc7JkbIA3ah
e4RINvNlxSbxODZVGmsuWyTZCk3qn6Ryu+R7TabCKZsoUI4KPdRvNGjiObj6
b2F6dTHr017wLi8lpYZuDellQrUXpj0PHHpNdhgmfhCxHjXVeiBqKQ8CHZYc
m0V0B/DMtgOvR2EYBfnMYlPnltljMN1vYKyS/GSp4cPvakmqwyP6go+CqMH8
GROAydWR/J8sCBz44hT3t9SSHYHmW62cMoNX57QeLlIvS6Vj+5hBxzycm2Bw
OmNFM7NK91XboqhwxFtPbiFovogMh8Y06lit4FvQF4ari8IqzcXakmozMJuO
IY3IsfngEby1iNc7YkUpRmzSr9LM3HMwnfScdO2+9nZ6BMcDeCxGcX1qZbDD
CelJbZ7nDwMknh30R2zAZ85wJdQHH/xRHWrGo5U9b6zLytXpyutB1fR1+V8l
B6TJKZ691PqKYJPLeDWQ64geD9J5T92HDW+8uSkq6I7UnVWyzpf2jc0vOOax
gZtSDjo+gU6ovvoRyo/p/mPtTRN3ZSWd9Vvk97GzopaI1mS5IIFhgCi0oadB
raQifzPagYKsKgKK0tiHT5g8YF6eM4o+ZsByb4wSrj3NlR8IWRu+jSi4tQRU
WSC6x36smnO8ze1uTcJEaWnQY2rYjYiTGLc3Uce92ZyOFf+RIdua3BoJEtZz
3QI7gldxUPA1GJUaTzV+puuQducwYgkBRyHglDTrWFsYL2n9iYBoyq5i04/o
cXhkdOXlgAJJxEswXx5HdutUvYbIhl5sUKJ5E/+Nmdf7ZAKjHvrW9d5LX5w9
XbSMifkeTLTBY8TAJ1F6jilcssOorJ/wVnoRwiMWgq0FHdBmVz8j9YCVsbwV
NSgs5s4NJjxrjWQM7FwMF5cdDb2/0ve7iFsOYnR185RlAwcoDf11MV1ZYaa0
LrFCQs4GDX2aIDkiUlGmBZW6TraWFT8DWwgtLBOj8Z9kCfblDMc9MlEuZl5M
1ebijLTp8lQvV+yoVJqGxc3Cxvg2oIStDOYLZhEgiNFiXd1Bb8OuPTRtutfo
1XTNHX9ufMWjOqmStRm/vZIkNVrXlGDeNo1vcMR0N6Qsg67t4eB1R7CsRAba
Z4csYgq7tMaz3lhilOXshdwXkO9XqgGC7LmmGoqh+J/1GJVytG1yMntJcWiU
Hn1Y2n3i5r5d/atihC8lDHQdKbLUnRji44Lpv/Tv9mkIbj2sMu9ZWjlxPy8V
WPfsb0Kn6Emj5qSwlVFEXssSEKkH6IR//wE+FuW30ulBfkoo9wW5OVPFxhUM
0cTsEkPMmcQPjcCiUG45bNVkBvDIXjJIaXlao0/Rr6iZ4mfrffedSMndhT1D
COXKtp+wLQVNaYkLQpZ7WCTHjz31heb+9kDRTmp7JR7jffQ/schj+2s7uCvl
bA8ceWGUTEIv0s+UGqay1zB1XuS7dbS8MKkfrHvq6ORyhkEeq9mL6RwXjuad
jfKeP4ggNpZ6+vRKRgQpfUPi5Pzdfk2ce4L1xaWro6Sp/Ua2Q6CGeKRKusx9
N00Bo+hnvUawxz9lotrSHBbpHYVDBo4wvPs5hykbQPjC9EJG5NT08hMSV+DM
3SWHI+g+WNp5gv7D8RCHeugh3jJ/yHg0GUIlrxlY2MG+4W8jlud0HekVoNBw
LW0cvI9XfbWfeFXDJZbduF33eTxLnd1KfBDS0HJmHZlPsu7SLLGuSJErS/ut
WpdK94oHMzlSMrHrKaZ7XTPN8xVRsxD3NqNKrD3rJXQkSmVbJz33ksyf8iRo
Ryf7Eq+UIQlSgpH9rWjDqpR6PcabyLQfKohVCfmi+9wbdyyehWCErfIYExkm
ztc0KY+j8JqvdDiDB7O88npP92Upd35vBZmdyNDjCwsV5yY6OoZE9RrvuH9F
9y8lutmXXbO7nFJwvOCR7zpFD54ax0eYR6STOJToXeEaixvtXxNNt0xzmjh7
eCRrGVe9eYPN2UD3I0PAR6jBKFNqJIbTnVHTnElDI7GAcQfIuqQqOrtTPweq
KBv7dsWe3Ehdl6FOWjPNTn2i2XfCY22CLdZI4drLpStQo5cXEmH5MnfG29nh
XWCK4lsj9Pz2vdPgLkkjMNCodEosEIqEV8XrJklRQ7sNEeWmUitawnL7/LPb
XibXPCjDO4a20kNsnnZ+kx8vdYyIU8OLYFNrqdiZSUlDam1hwotkqbLNF2aJ
+BwgK2AtixEjCjFWeqH7cV/NGhnc2Gpd1tjMZUd0yzWDMVbdzgjY02VrJLeC
vMni9DMSMHyFOQw5JF/ASZISMCvyhEbbrqN4Cqh10DU3QbJYjB3Cx1NSRDR4
gQZB7uS+iCuhT47EUnDUd/h6kCjUM9D06zuIfRbQHsOQjw/Qej2UdpCwL8MI
SL3lG0fqG5RS93fPy+DXOKpCYWnWJvfSujI6mpyORRVxhuGfhKrQ47Asy7uS
WwCKtMOUCOVcUiCIKMwtj76DAd7hZefDOzyn06sBvqpLHtYJ+xN3cuTUxHKm
BVpaoCFtcSv1U0Fn6Qf0HGxMvkmMI5NqO8OxFhLr7Inl7eFKSV7z3kE4CIRw
jBqejwPTbt9jnZnZ49jrY9cegIMXKsCSxvkND8+AUw/VNDC+XGqdG2BoOg8P
TwlOMfbMK4SPkOZ82cjfa1CF1ryMM8Qje307Jb26c57eo3kb1hz+/cbmGyh5
c17m9wzXPc3DHQIdp8qIoc2J0MVderEfB25SFoD2Y+CEBwI4iuDLIYn/m/Fo
GEpEvPHCkR30bi2BSnuDLcoZKPswTXQWdT+7Wtfsy0XXlocFE48N0NS5RBJs
vsEWvNvywSy9Dg9KqpDKcZVsBpknAa2j/9Nd3EujtW5ciKfNXFFrGAD1WZfK
01q4ofaKzJBTz8CoJ+YOhkgVmw9eOEIzVykdRqYwRAJYrpBGRt3Xoqps7evS
G+1BIK7sSsn+efGo9YlksGvHIEEHFgLpXxh32UNfg1TKrB9ZcP7IIzS/CrB4
PeJj9Iy1vX0sG4ZcgdQ0bYPmHfWCTTti/k1w7WP016lIU505i5xoBCzN6cnR
GMBSTqxXBfzYvnRb67W92OkzFyatZvw+JjEPLXqtP5ihzQ61tyn/3xMBYVah
tyYbayxyzkQVeo0577E6cxGZgqxL3N/RBrCSuJJJUedhk9dRLZ0vLqUbFOj7
uQo8baabbkHGeJmcE6amWakmHwHI8656fpRFsLjiL0FI5L2qCzy6RMtnR/vc
gHEHb9Ag6zEDoOk0idBTpyAncJMEJGSSXgdeRS1uYG5EXRomJyxy0mJkY5TJ
Rc7yoxkfR6AbnhJwrBXlk34P6wHaB2Yys5e5eQyb7QNNQ6skV42Aeab5twEr
6sfuxzVx2m8fqn9Jok/2fs+/dEtBZKqZO5tBHLLNOylxTR3/sYcgRbvf+AxT
WdXqMN0xMwaEizGTZNkaYgc4YpCybJfVFjIl+8375L1AK2yYkXb8IOgWg+kh
eED4B6oJ0Hkag29lnoC5LR4uiN1gd8bUWYYeAwThg29jH+1AlrHpH2PepMW1
Gv5GHClRgskwTQfW4az/9yG9uK3zxg1WaG1jvzywJT3cBAi9imOgaF1SNMfi
Aiec/pBlUdPMXPkiRRhww/RJpSOV7g3eYrq7H9Ll1Dc+g/EdSbMUiv+jjfql
5yhvXQFYD0iaVtFjf7iQIEUEk4iUORbqomFBtECOxR9sndoxU+n7CLWaxAIi
965H+aZhhA094oXfM/Fzjx9+2YiZPPcczvA2ztq202Tm+9MJ5wLo56dknLIS
eM0MgEFcUlZ98rfOZDuAREApWhmf9Tc/ibWjxde1/uNOTG3G0pbMTl1ZBQIs
39yAFMkdd61vPCnJ0oqCgORw3ExgHU91oWnR5Lb2Xkp75gZQsE3ALMG4QUD3
dYxUvtWXGV7ogGqgsExr9o2BRXx0M8LYF10Zy4rPlNY4c9HeX5D+NJ4abhnh
JRL66tt1U9PgGRgPpU/uxgeQa8ZvSSw8fZchEaI+inIlD7Ys9Vr+UZB6+Riq
eDqUAyPWTdpgTyEAN8OVenE1bj4qsZSZuJXn6MjDk36E2DxAWA0w3nTB0wdw
vaJJLyXswctxHkpF+F33xLxhgSTlnHdriTBClB1q56KTMwC961amV3CSQ/q4
Kc/SEWuLr8Ip4L25UWbQEjPB92DUOWq/KtAIYp+gvEV3Qvu3GLRQm9BnfbzV
fZGpXRwgNimowkiQp70+mgymd+TBDNaEV1/yOzbqkWc0hUwWIQ7ezF6/GcrI
7sdvTD/v0cDW0B8aJYlPTJOIvf7QIpS4FsuCFjXjJrB342MuMxqQ39k0uKJ3
Dy18ocQMnTUdHNjQGkFFkxjGIJn9Fmh46aZmB9RWEdxmyT3TaSYoPi76wOj7
91SzH9PLvbhfRyUaXxMrOXxLTz5NzynG11AhWJ3bA2qITbVSI2dkUAz2TA3n
oqVJBkB4tyXrFBY3JGPXn/euTYyO3+kO9E2qd1/bmjzsupEsaHAGvLt+vYCD
nxsmDZDZbhuzvmbUOPsjGYzRYr/x+ajmcxc4hZnqNfgoQdVIYvdk6eoc4d0o
D8ELVDN+nnHJ/+zvCIXFJzbiig/me4iaX5X2uBB18MfSYVaDtHRrxrafD9AO
jR00bsU4I549JMTe/Rl6pSkedEOB5Zx91s0b/Wzjwv8Uyb3QDwfK5cslJZxz
vEmwmUP8oJRgATbabrXy3SuZDWwlnDOa37hsypNqITERnGd0J2hp9/V9TnVB
ADpwZiaNVqDshggsZZyXY7bLUHgzBBD4fcyq0c+s9zuDB2B9VsZMG8+mrYOs
xTLdYHruqROaHZVzQ4d5PPujKa/j+ck3XqS+4OHOrDWxCQ7A1fZ0ejjtoJQd
9QcVat6bjDmeyiqinHrZUx81YM4BB2Z/s3h+h9c52iBJVLEECTW8Yohh/fmS
HnWRtoYBLnullgo3IDz8sMBxePpfojSy4zjUPtwzM8C8PA2XrTZvegPk2HcN
RrHHiqwesCWvP5D5vw2VfKpqAMbdPgM+7Ri/py6/Frd/u1ldVFdygTEJt4an
TBdoRMWNvmduL920Xjv35vPUn7N9T1cYUw1GIfiMDAnMlND08QvWRjsYWZr1
o5Kr5mCHESTSnLoyNZKhpBYyF0nnwOz0ZwlN3ZSSOhGS7nOSpYLHnZyqq2cZ
Jz86uQo7EWlNBTw8o1U7jkZpV5PY2p8HScUkUeZqcc2r2QGc1fzKvQv0LMVN
365axJ8tgnc25o3EnGsTz9rypCNiCRchJEwHnlBbQhYdvPqR8SM1FyXoASpN
fstruF6ZDLrFCdzLJq12cmaHTHDMYp3XLKKDLRqObnK5pqyzMe10AiaN4sDg
/hQL+gAwkDa4yBQbiwroYAPUhZBKgViYyRrUfUauu1bHh5H+ADTC6j+VS5sm
Qs2nspjb+j48oocHcVXPIq+zgtssTt8Vq5CwhHx+4vbNiEOHlGfmmkLnEZ3J
L6R6UX7Qm7t2dvsMxs1WfHuzCDQqkbeQy6cHUI5EMAZt9E/QOt9nZ8ft5Pp/
T1u4mHq3Z9jjPlzRHE0gyGvpm1T+8DEthIv9bhUVAFsDtkld0IuhEBB5T/B5
t8MZFcso+ng1vnucnCwQAUMMrW4PWVLcJp7uOIarRnZaDkTfGCWD233DULWF
hfdzYZz/UYaa0dcwsus+hmEJlIGN3K1yK2tY7QRLtg2x8GUk1+hS5d0zH7Eh
9Ydqb4dS1WlthZEYsaaIXvZFom9xf41ByyOHXYYPmKKDKUAZTMTegS/G8amW
zbGsHT73OEYU/tkZXstVPWSI7o/iOKJ5gXdc1mWyRiKYxeS2gR6BpC1EqWkK
mmGNLUT5YL5ICE0PxstpGk+WovV0qou1f3cBMMSFQHSSY6mijRms0YkBYpW/
jrPcK+vg6LsCc2SgVUpa9R0XHhEGhmBYwTxqK+Zg8fapS56ARl2lWfVe/BhY
qwbpSnJkUUnCGoKTdU1biS+VpfoCX+f64xJlli3bOcR/68kDWV1Q+3idukvG
Y+0DynP2N/JjokADqI7cdW/nMMV0jtJJxqWMKWpvABCTjo34AXJw4wU7edv4
PlDXhEtqQH6foE/DaqEUFhEWmf/XG1dWMaXv4DYDcfxqkSmsFkPTyoVxGAdq
7m1cMdfzWhEwteNZO8ltqb5Ac/4KZkk1WiJYSjAeYCy6mCtptuOwMY+fNnZm
TheOCXumAGfim/8Q5tDBiBhmw2AnC2YJ7Tus1/PuyeL2uI1UmUtzE6geHzUl
i40oaoKuSATYiQYTvwnkcNt4A0Cv92v8ANrRnOfdd6MB0MOQ7+BrZ3JhFtvm
2sqKdv0l1u7pX9HGhziDyuhXHidhBMqV6PNAMUIeMCBBetGIsy0lv3kA8nnp
W0nWJ6dzysxV8WmMoPoewoq63j7ZyyI28SzLiT0j3V9eNxJrKWJQIDdUGH05
9gw62OpmGytQO1PRbuUErAAW8xvtmHhbLKVOpPTr3y2S/jt79TC3hZYU1veq
pg7Knn5lhx6FQFK2/j21KXbP8a+RMviEpOPZSlR94enLM6zWNHYrLEOoHx5v
oyC06ctHDef2trPvp90dH0f6jHrNj1Xl0M2o8BH2HuVcwYBZYZO7F4wGxB4x
rDNkWWF/Ay738P6oyoGW4+817G2lPbwCndVfpKJF4D8XM82NPWifnhUXxNzn
Ho3dJdXEM08BebUgudxhybeNPH/UNUCPGlRBxBtiW3dQmk4fmzCFhu6tNG7W
25DXNttWU+DctNhxtIQKvv58L2V9B0TAl2hDQ6FWf5a/AsQn1jmRB162fx49
V/vZ3Fncx5TEeOmqFdOytPcKUzPgEEzYKqYMSUElTIiUR8pnsHz6qS3GYWVi
6JPiJN8uBstpGn4fl/0L3ofWtSiM6T4hlZ+YVsIp5l+yK9FKW8qIJiAiB0JQ
ppnA3lAyz8zcni4CZT7BiKqFDzTTjVjP7UjCR+qTZnnWGe/kp3KZuoFOBNze
lq7rarhH4ih8nDH7vRSS3AXDA6iLo4YNkVJ0NWMUToZFsoDm0XpKAc6dEwXk
OhivML63qsNVhi9GrSS10NFsZ0MUdzf9q8sHGidv+C26nc1DG7bgf82CwLBp
l9Gh0JsL2/yZuHA2+zk0RQeyO5dXiLip2hMES0mYPl8YWGmVdKPi3S+NRE4Y
DjV+lotPgBhpkFvOC0nNDE96MG8kReljHykNz/YVIfq9f7EZEfKK78IUE3SX
wQTaSjXDtELeeApMxyENEgITtoinTQ8hSmFhoRmhAGksie7mOqYrE/lW8DnX
g3DWI56i4RRi+Pm/FWBxRj88Njzob6am3GLQ7zkG32OUGcOg/GTd2fBRUd4V
FySRvTibNDFtLQEZUX35rsfSM+4gVt+aSztBvO4XN4pjVfSSeNeaserB6Aea
UaRxl0vrabWnXJHgfijsEw+nXq6EuDi4C8K9vhpuM/+EWHvfuP7QnZt92n7s
gixr3HtUEW55CkbYMwkGsDux0tVDzKIZn4/AWKwHH5BytSp+htlmF0FGfd1S
l/7hLI2WuPSReVw/H8BKu+fYW1TLgdjbGoVGd0eg64CCNS8qwi11RSNjCcIa
Urb3PGzpm2zLpgWlqLqnQzYp06wN6zaMG6nogySPI9XOvFfyxO6Pu12WY1XS
DeZSnx60KAJB9oJUSoV7oAmcbGzwG2SO0WleMyZAZUNf3po0Pcmpw8pvil05
S0dWGs0NJEbZE8Cm1wTznwU9qSL7FJTx1+trY5ibRw80jb5ucmLMlotTJ3P6
ijKG7vskm5o89m3zWRUe5mg3S8Q3LHIYrr7/RKV6Q7r5oCLzD5Bj1ppJbQFZ
/pWTNH5I3b21G7NuJUibTtZQQ55XSBzkhFKu230amWZEHH+LRz4rHgU0Oati
njljxgeZETGc5fZCW03OttG87QmmF+KG8JmHSzy76FxUolrh6nOId4JcI0YZ
4dmi1k104V3N6UYngLv7mg7ZTbeXDrGUl2hqMT2/jicvSZ+Hl595VbngJI2C
WEr2vK2mlEaFwy5Ei1paSb353nvjDumcTS+ER0MsP8/kn/oPrnrS05Zz5NYe
pObmZLLfMcfNK3NuF75OzFLKKH9cOf+L0EaVPFN5sQO7xgOun8gf0mq0CTiG
FE5j+rJr/ndNZi5NyFuQOzXG7wJikxYyoHf8va+fmAND2WA05MAKQDiGYbsI
HQYaU9J/dhCT47eER1iU1TRoN6oVh5uLtazmL0eSoKoShHQtsxfruJ7odbaR
q9UnQz93jY9swKEEDpdN5dJODh6D1CTJOPyLLN7ym5+Rm8nFFzobbhQa+HPV
V4TvOIXGDPbDnc2Yj/cH69MehUDkq4kW79BccljU51WnuM672Sq8NgobPC8k
HvXCIVGm6G4X5lrX762I1e5UDAFp7E0kStTO/mj4mRaD1CM7Ei6JvkTlIK3A
KB3pJV7kaGaB/iEs7K6yuev1fNjDF19aoSxtshhq9N88tAglN1d5qhSa4fbN
dsk+g6ZRK69TZemPl8BDY/NGLGB7fza/Q2EWhtYBD0PVf9djSERkNCukx5TI
qU1kUDZNLZQ6BtmfQlfSqCqPcxO2ADTnhWl1LlgeXrvLJDoQj2ZFX5CeMTNV
1eYXqUvYs5x9JsoJyZqLrHFm1UXz7q3ScpIDeC77MQylLImvoA758JWof7bj
Ffig9+FWblVirmBPsbe1wnMZFA5H7mGBNfXi18n3vH953O8Mh9GOwCtqGQVk
ZKDLfB4baN3+SU4wgxTTvmsElIFaJaXq+OaDz6Qd4CA+IZ8RDBR1Ci8PchmQ
koizu8mt1VsfJIVaLHS/25PV4f8eD0jHD6jr7XnhCcIC/ZYB95iAN9VaDjtJ
1yuNwTwlHsoA3lOApwcFOFVgRHMGitUfKWdqlK3wjyhg1vTuDmjMrwV4T+6L
P5AGd/PAO20GDDKS2xKF4KMcukFAHo/tRV2e6kl1EPYz1dtrzPkFJ4mvGejX
PMk3Zth1L+OZ0UzcWLhKYYfvbq/+518bI+I8JwtAZzWEm3TmeH/2pVxtX2Xd
E51kJCssn/35TZ2wLXudgum49pJ7mvWNg/tcLXfaVWPgpjk+TcePUTpNL2ZD
QXecQiqs0jPyjBAncscxmreMJLhV+1kxD8uJWOiCD41yt7RCHeyhJP0fFbBw
aVCVQgMGO2aP94XTSPyrJW1o7kIFpxK/DARdcZ9FIwNt32NCw8NUGlzLWmvj
5O7wluY8K5Lk/jeJBgOpQkxcXXdJT9+yJp29KZNowSB8UE4r4DCq+5+dxXfV
EZePXW9tdvRcO1gOBOaN7zIuzbo7StKEuIo6jxq0GKuVYUew4NggHKlwVzQb
pD1K6IE5oh358Km9QfXrViuDdayxPNVLRHIZdcE9IRub56JY1L9mPpFaeDVU
Z5o+jNJZxms8H40vC97N+n6BxZP7zwiyR0tlGmakldM4azj430+rHe5Q5nha
yf7gmUYPb/6mL0TAf7kaTnhSMmFJDnIrnOoXkKKBQDTx/Daz5PCZEyGOVW6H
SmvxqSZClu0xDd8l7D6JJX+0E5nceyEE1fpf87ulUJjMILI2bMUZWmI8CbX2
c5cDASKMPdgjGiwIaB8dw89fA0EvwrhuBikr2k133uAb2+aE6KPtLoJZyACm
TXT7hkfrn/p2MtgdUY8+2JSgAaAsGmdpz36/VUA1reifyxos9jO2oPHO7Io7
fR4Ldxd7M9S4AkCBL9X24oXHvGpgd0AUzSNGisSgxk1PeLSu21kplYKibpAL
2lnstLu5uKqJ9f7udCIgWUNfl2IVSsIic3CsX8g5JbBf1bl6f46fApotzwnS
dFvvJ0KLRAoFhazC04P2go/aonzq8h4B1ng6Mc6Ad5gTn6ACCHX7tzOSWU5p
V9DZutg51sJvh2lfQ8/Mlr7oCCRXwz3v92M+lhOVKJXWS+bsm6Lw/MUr3RPC
2DV0QLraeUB2l2fgFTOcaEJYTBs6qh4Nisb70CwdMUkZ1zdrHjdSaXJSSwbJ
zra2m1QzRor+0KyiZzflfGbt2H6HJzF2jy9mxfRU77NNsVASrec9Na0JeNX6
MMxin20VcFq9lcrpL3NG/dvuIl1YYFQQvLdKXhzzVF+49JH8HVvhMIr2h+MV
x+PJAtqQhcNeTEby+der9BFejqjCen4j71sR1kgZDqIsNZmKegrsdRQ5AtNj
TJkco3SsQsVz7r64rf1+jOayFY7HCRSr2kF1pKHJGB97uQhojlCvaWmtswbN
LBk2y/t2gOQ2PKJREsj8fBozZfeS2DH3FeGNFOs8wLN2RU9uwCoN4+iKpkgX
SPuxKTm8ZZ91sUQ8Rs6LrEt2BxDdpiquk+w9Gb06idaYExvZMWWfmfJmgn6M
AkR7f9Io4JQGaBomHvqRVcQ73Qa84o3YwV/K4cKxtQpZn9KfOjMSdGwiW+b6
sDAPAdZcpz6ajNjfVGmlD3R30AzrCauqgFKlQbbIKrW6/RqKAvH2tfHO3fjZ
5975B+cwcERlmW2xXtS/4jkeE7AwDjGyuxhbaHDeue/l/Gv5dq+CFUw4xzpe
T1nUXt/L6xu7HUWTfi/JSyeQRDaBI+CkoenzYn6lmr328dgNcwGGIAMLlrV4
fgXRhajL/FfEU8g4J6IoXWjeoFojyTXCWlZEG6dYuCklSPAK7vV0xGPG19+5
BxfgOep8/xGCw9KoZi+6Pr92h6Yu6sx6FRGEUfVJ4RddYbq/7PM3z9WPC/Iw
mVyUAV6ze5lJFYjP0MSaScEk533d4repfdx7xa15k0q/ykgSdurcdwFXoYrU
q8T+MA8OoX7027dVDDDBM8ATg3t3qMO8b7yasfkwybvDoopJv43lwCBtzNlO
pq15Cd/GeSJsLG5GfNhtfZ3e6peT5Rc2vayadlhRRBvozFZbvYp9x0pRCv7a
/yL75BQh86c9yaCDjUbbcFLKkMZTLJPREM2KAuj5e0XRGpSnrXnAEhN6T/x+
IRPYTGetQ8Pv34XsciIQYmrN0O4Rz9WCq9/CDdsaDSJOCGMOrK2XF3DRzHz8
dNK9xix5ortf6smZOJD47nPCoplCPx0BKmcfJSq3q31Ec1m2sBTrAdNZHflt
iPM0BXn9g3UlMCsXa+W3Uj5VZ5/k+i/L4f6rhE6wv/NQcK43qAaBdyDudFgu
Uc200t1GWtXmVm8/aCSwgK6ih1XB/gKgEjf4QMPXnFIe8ISuellyIuT1Q1ul
X8KkvrjWJj2qmuoHC1MAQFiPAQYXKeKVQ3zeQxG4jRo8MjzHZsOS1GDe5hW0
55EaALe7bUsdmfUewwGhrEnxRD/z621qhbp4bZnE3XhiF//hymH2J9eS9nwu
D+Ango1IahIta79Y791qELQIrGos8LzJ3r1iK40FWdONX0Udhy84p+0BlsbN
AileqRAlP+gHLzX4CSUWeC+tG5A8T6SCcJPr8keHbe3vd6t8kgzgpRee06Cr
8giiX8RJbCpvVwNlEbsqeq5AQfqs3VIgIb4STmCknA5Z+WBABVg4I/LBQfk3
C9lqE9DjWNQmUdw9YJ+uSmCSpnPpkvJNE+ABKOXe89r5Uqh022zLcOnvAnrs
qZwHAQIjEK+7PlppJbhFvk0kx4af5dZ95l3KmVYlYRXKo676QVwf4o10Vc3O
y54fQdeiCkKGoPX6KlqIMOVM/WcBRhK9qvGKi2w2hRTLnvEHcQWXXX4/uTQ3
0mGqKx2AQEsS3iEBLLMW/u4jThwl2DGww4FoqwKJabUCakhP1UhtmXyZJOj/
Xotk4bcnNZJQtIvgAz832ny1RpKy9un0/TqZbr7QzVh2gvm5IJLihoDa/5OP
nmFxT8UVn8/lSdGjrzec/RPTg5/8ZMBrbU2jAspNO6WM7AvsDSIANzQoByRG
Ts80WDOBIzQxmrLNSsYmvxCZlGvjgaqVsSjskREDGq9x63BJVheVm8TzQfb/
racYbmXUpu9tJ0cvNKPv4Cv0jIbbY+6PtVZeBC0nE83MyLqDAh5FxhTdRiN/
KJEbdUoeZMZaKEt76P+Ee2G3CNR6p5N2QF5h+zcOuM/t+PZ3JFltNFqDC+7X
3jFGeJVcCb2I1MO/RCuL8gXMwdHXnfsq0znhaQZiAPFQLTAx4LwRqZvxXDSl
+YNGpSRP8xVZmmocGo96ip6094PfaEHz6gi0HqNefZDK8116yACkODPwUGPS
kxqaPWGntJahfQLfmHQ1BL66zscty6xCutgmjMnKXdB0F0W8N5dIrQlibF2E
NZGOgpt5lA1j591pF6RrMLbwAEvzqPj2at+uWd1jarRd9xMA2S2HKytH8wRM
xTVRgRQiE6cbE90gqk7Qc7SBoLMaiQIXTw+1LuPV2C0wLcWZ4b2Y/msVYsGK
RlBU+gI2uocfVHd6TW/rVQ9eOepMLJLZwdRSF9n45n1uiRC0N1ghn2pQJYAA
Z1AlWc6Msk+2sbwliBLXBNHwT6HnHiFkAJGpEEK6TAd6+oFq7CKGCGcAZcFE
qae+qFS+h8nK8cdyzNLTL75oFGuk59mQhCLxe8BtV1RokuI8Z1VoG9AfLvqE
cI2HPFJlXXqrs/EqI3W7zm/5tHlhecJImrFXfJrBnNO7zKhne72HyQKIz+Df
NGF7ECfBPowmeiSpigMZEtengFoFbduQhWbnkBPjGuoejQzenDdvNv0/e925
I6WO38xIhdL9vpeDAu3C18fTkDghFjE9/dvpn/vPMOZiK/QyBjtq3jqsfPDC
KRvYR76BEJlRSRmmoqY3PWURtUj3malsGqB7VSRPOTc5idHdt7UOilcsvTca
pFDqTePUuxP2j2RxGp3NsI+KkAcn8kRdkqCUYflJjw/1TXq3K8lWbqKaGx21
Wto3/+paqfy6tf/4gKUXTPSz7LZ66g4vilzpu9UEVPR4dwK80rVhBxA16gqM
FCXOjXYJfg2gkTuCDEsm0ogj2Wv0CmimNL4msXPJzgdqzmd9FzpDH3f/n2aK
ayZeQRLKpkH6pk2H5FnFX3d403GZwGa0J3n/UkptI25cTsQAVFRhUXgT03XF
ELY+zrn/uXuRs+4YVux5fC7C3hL1EqSbfclOJ74y1Y/Cvj6T2wHM6fHT4uLH
DQsVCCz3wFBSTVs8iliVs0UtNgtvd9TCBzsqAe6SSITnAm9f8VRCFjxGj9hW
7c2QGNs0Z/3yIy437vhYJOnXguPkB2Qtrv7mjyPhXBqEaobScPho09QI+1EM
qPok2EnRClz2O5WuaXhcjEvf57QBWqF+adtzZojm5+d3PVuR1GmqT13Xxg+Q
EMI/7cSc0jzNl1NdJSKFRUxMXRvNcXAykNU9DTKEJC15ugtvgQGWtp9GCBNE
OilOmx4R3rN/jrW6OVxkFr54kmlCZ2Fs+1glc341wuvYbutV9qW+Rij1UcM8
wtBYmKV+YnICvionpDJjy4GkqLpc47AOj/G3uqYfxlWVH+r+IEYRvJ/4hSoo
cwV0CA9C21kMyDO4yNJFpJu+zRWF4hRDGMDFCnFamj7Pcsy06VwHKxroyB2s
AYzgzm2jNLCxVJrNWH+2XGyr93tTV2Jn+fhqfQ+h1Aw8Cpqt0ZIlWjrTUVm6
+2HCARSQf+xNaKnoXaMbYsndUm6OWq3ksS+kOqCdwKLfjSoHgTekCgqUHsI3
cfIsH+ZXpubgV+nLhKenhnlKykB5+5ziOhIEzJmRohoQVCCTVTTo5aXe1f08
gqbJyblcv+1U4c1YtLnGRteY8n+s42y3LsSpKUMRHigu2jqzAmMPG/urKayP
FujaBJ9lg0jgAL2ySxi5Iskm9dpnhjuywNKcS1PjORg4JDEVSt53UhEUY1Am
uZNBJ9WePgi6pmCXJs4/D8ENvS5vmt0HueOq+98GyCmgCBhUuK1sGuWEhLkg
0OZMdVdH+fvuz4IYrm0wNMv9OdpczTGg3UaRSu0RJRRVkhJ1vBHXaFtInxNz
O5keJC4M6v8miXHhVbFdyr8lTvDNyrpr0q9asTPjgp+HsiPGTgt1F5DPxPof
qNfjlxvpiSRKGIL1kUDAv1mjyS+pR4eRcpGUKC47Rerm7q/drR1nOMB/nl2T
wghAxRc9AF6vnfgJLZnSQFgTjX7qfZ8iAd5JtC0xzxUh0C1x+zxXk5yL+Rbe
PTMUrGnsPvd3NFgIXrwMmtZ8wtwENOVVzmv60Zv++v1fqKv5GROQjr+7z0db
rYOPhkXTMpdvhmbTBQi9cmyLQ/lNGhaORsmtW34b7SaQgFKi/MdUXOowkN1z
COw4q4KHTKyfgPnWIT3moBMqRiPBcgEnWn8TeoPHL+LqQ31smf9NhCEK2P5O
atWUwCVIsGFUGrA5D6+2UPfjnZPVoU4lutnoZA3dVrZSQoRYcs3kcTfoSce3
O6e4l762dx0mGlxmzYIH0J5xnxl4EjoA+IXPTXzpLHm2j6HpALq/yp1kC0w0
30zpt6sYpMKL4vMH0oDfkROdOTuab6u1wWkyyFKwVq03UtffV1tEFMipaMtz
NYwzzTky0nyq8lkkHlc1W1/mPnhEVy8khz1Plt8SueJW0+ymPsvXeU+aeoiq
aI9kc2Fb728SADdHI4BZM2BmtRhfBXbZF+4EzmUyeSGbE4LndzVD5Kkr1VPH
dxzUxeo7ynZwdWRIybvIRGHcs/LiDHzX2shSpn0tZumAxAere5czjgPID1F/
jPSKwbT1L0k6b6u1o+wIKOP/nzTIWy/N6ERwo3UgX5tQGrwDDnvDdj5h/uq/
3t0LPKnpWJEZE7T9WVyUjQvWko0ihWmovzL0seSK9881DBD33uXs6h869ksn
Z3abShEkMu2Y1D4KLrIowjuC04XFZpqxpkgkx1RMhAQ7Ycbiw0XdJYvV82v4
cP3XtSUE4hoCkzBhBJsWME1puKRT1oE/W0i56fls5Lw2E1KMXmS/6/rhUyCS
n0BlJfXC0InbGBIW2aQZ5RcDF4wkTgXVDTJBbROwDCx2dC3rFGghlRfpa/X0
gQ/3kdfJ8ab9BT0U/NV7Y6AYBk0I4a82RGD8g4SptaWXLZx6EXy7BF9AcpxR
iWQaYc4qZbYJQuhH3nyeWwOCAa5+i2bVDUD2iIHOctjjtqZAepba51AlE2Kb
j0se1xnTx50/BJtSi3O/SUy9hLLF73vgtZGl/vdsKSDKbUP2kcW14HUMcBSE
PIKC+LeDOlXPw4LtmqvwCGzZKynQoWma9dvqxiL7pzLrGVdtGVfE92RVuBvu
5unV66NOQC3WOoxqhMD3cx7blYDCX9Qq3rWbvA9ozrz8dXtrsa4+nQXiMcSR
2zX7oWsvPztBEX9abRJ1RavlrLyZif7ORIko+PBpDhCE6lJi3SDWoXcewG6C
soK2m+sgBKJfYMwRTxEwUki9PXoPpPjA4xOZIZz/yxzxicTSm4eEz3gIDVxG
Xl9Sb7X782VkehjZ7HlUAueWPcJs5vRK6sL0dw/ofT0zcwmDKZf6cOfMk0x9
2kPzpw1AeAF+MiEhF74uOokTzN9698cHj+MHWi5iY/MLVO+Uw+csL7Ivj4W7
uNneSWPlqzUFUrgKnrC8576zvlnTGacci3E5gYSj7QL57FMWNzx2fFKpteFS
1prqcxpUC5x6jYmujQSjahBEEk+u3VQoETLymQ0jf5H3BmvDoer+OcgxMjuq
d75CF8/gVXskVx+9bvkCldxlIJPIRPhYQeprrFnJimxMvlJpr6eWr2l32cMB
ghqRBPYT5MnYgxr5Opf71edqSYPzrB43cmtxLCnvNBbSbL3tTLIJarZtyuoL
gpC8te5sQn3NwRpK+KwEsr0A/dIkIKRZMI6967spzKgmGZoLtP/mo8KvHXYj
Ngm43HIcETqKOEA1cIuRrkElsD4h/rVpJmULWBYeRUA64prIsoj655RGwGsM
bHO1uF5BuwYvZFnRFuD4SiQfUludeB1VMexJsjBrQhYa2qQ4KkwaW7FrEW1A
DPv3jcSp7vXkZTOCQE4/G+o7XZ8hcHF+zALFSxNgWc8C70/bSKOBQf5ssL5y
bP1H6lSMtaFz1kDn1PoC4CsZ+DVAvTRHx54+t4cZv17wKXOm93V5XSOQJoZh
2FIWiG5H0xy3oe24xmQZgQhSpIaQEVeYUaobqd/Lf4JOuhlqe7iRuztfu8KH
ceZBC+cRJs5MmcTpetjPM+sWUqtdhVYMCKNDu8gCIQL+CCeu1u/rJaLdODMo
MhCWce59T2uh3JuMks3RUZq58bbpAPz+W0dUPrH7YHUhCfRyaWq8W1Q9Q2FE
1B90zpM9AMexiC/yH47ot+jSqdFV9R8xKso/k8rAUNFU85jQu5emdgm+sTB+
3BCaWhC8g/+q9cM4d9Ar9T24yLBoOlcOsD7yJYlWavEZHEY2s8KS8GgWh0JD
SUtsr8ofq2zmnxr8T2M6hn8h8tsBHc7TMEifkjdqbRLqsohh1BanKjJ26nv8
i3cAkk6aFzLyEDPz0yC1HzVV+LGlouaS8XyFxmvEBaPUWSMcZkeESkH4Kwpp
OIK/ynrjNS8xZF+gV/NZ5AthcQBAibVkla1OU9bW+Pdb2/xmmm5BDlinzF4H
wFOmOgex4zMfy7Iw0arlxBTZbGg0otAAYVrcY6kUuo4srkECRNWgxzwhQ52x
WRv2qy7otLW0VhWEuWQsKlUGaVKwTvoAfuwEVuvDKoPCMl56thfVnIsGVWV3
z2RvYr7oCrt0RuL+YjQSmwOH2WAuQGsWGtZtKTOQtLJryZL3/ARNji6x9bmY
O5GsFebh86q6igH1jx5pOmhQN5jnVI/ojmP5PdoNc6zQCgqY9NeQi5WxnN28
qvEpBl1/SoP7uIgLEy87xIMANWpwOVMHOdR4KXWidFJrozNBOCVXAR6emgGE
mR2LDfDfN0adk6rNJBhCEw7N4YQ+T2JiNsSRla7bdZDkeNCLTLYNtPKIBWB9
yBkosCHI9ZEMMJULiDx2Y5kXtn7dmDY35XDez9sx/IDcyhXrRF3LjDI3U9dW
K5VrC4yH3hic2u7va4IawVJGBU2Yw2lG7HLUf6y9q8zFfutjX6HyOpuBtBle
hChzw8DKeR8m+18mzopkQXlFj+z5Clbel1upwI9bZ8TwzYMRZFsY8zsduj8y
aGRIdGKFKTRGCF17dcT4w/AL0YdekzC573TiCoI7Ur2Eq72ff3uJ6LvLpQRp
76hIurHl8nGDnkrFt4RE98FzHfH3kdzoVNRrSg7SqXU/9vXs7XPSfIMqN4UP
FNrT2PltNFb2zbiC5lNFIcmwi3/vxDxWISWV6ycideL3Eo9yUt6Fvfdq/gCA
LnJEEnQx6MeP43HWgxKbJpgyGuFeD4MnQeuX12ODhaeLQ4m9OlRVAiUIFzjH
2cLP8XIJmRAgEDpxsXlQ4TMw7l/yJyDlwd0flitSI0Cpo7doTQ0frZeL3XXF
Q9qo1VWjhmpAdqNMtQFgvIEOJQpXhEwxeYJo6I+yFPgeBqyrNqE3S7CGQJ16
Vt7vnvIEItmbr2dv67MDzaEZTRcPgrKxpx9XtPY/kCHgqk7ny2OSJIvcm6i+
HWYkTAfLznEefzXDAiDEv8DaGh2a6zn6rMrk9LUDjf6hp9sbUH5vczaVNr4A
AN5ZhAuqBmhnjNlAu/0APIuclR7xtdlLRJEBpJlE6NUMoD4I+3VK4bTfmooF
ZCqiDxs1RTR+KNxxc3t8RF89Vxx0y4S+38bUcsAcnKr2t7yfuAy2suqlKk1p
CPHk/ivQphrHKh5w1nkDeoFrRSs0cxJee+W1oYo7XSLQjG0MHs19rFYzn4Yz
cWwU3Ve0F+feeIwXHWDqMyG4PgoWx3h+xDShqz84qYDwhLquP561AfyGKYQ/
KPXXEfBkF6+qV8uOjNQqaQja8+fzcfD3p/gMxUdGm3UbPUaegoDfiUgVGfaP
So3ARptJ/mL92aAHu/mD6cwWSTCsaAGbyQsTAwm7BqWHe4VRemB9IfIqrUOE
oBgF8WA7//ntzBHjBRWGPE82cQfom42ZCN8yT4Zys03ZN/PmPFcgoqN99sx2
7LNFa3xiKUMxkhu83S0jYjYVbR/pNW96RnP68ctfHhWQZal0XPMVbCbHj1+7
pGALRJG3VjePTGUQgvBhjW/Il2aTG837yB4TxzkV4gfItgiAhbL2GRYbXFdi
OPh0ss0nUrAFvhAxwhn/uqKRo2wF8kQMmzT9sePX+tTITArG2L4uWo2PdMhN
xJq30mItVXYqXi9kWF/gKsY6+v7qi8t+7MjXJ1AJiJgpB8Q6Euha7GjJweRt
sBJnv2ZaniaRb8xUg7hIt9MRlt/RhKYHNTvnG7qxnaiS77ZUQcPyG5lOsuXU
KkToS1RZQyw+/G/riDxDXhmEcN+jyjjAebCPwaqgK1nrChy2hUHV77to/3E6
tcIroujd+924fqGtrVZwxAKF3RuEmG7TH8DJVSQe55fOQQnrU+/tD3t+JySJ
DXiu9xLyaxLFWw4TwuQ6nuJrKhMQlj/zbz7pXVQ6mC25aOZONQdccWZU2C8a
ooBZTEB1bn/8nwSeYn28282SK/XoFPhkMg95IZWNW065+7fYboTEkfytmdw+
1d6HlGEg120wDZaATfwXag5dqQK4oUM5wN3qsDK8lFDIIRX+Abow7bCo03he
u1rYlRu0Uwryq0yfjGnADq/YzcwSLhHBaHFTX2x8W9o/ZsOEKftenerv29ik
5EVjHxIdPLf9R219Xwk0RaDqnHNOG4ZjFEoRpMjfuA4crdJABVZ7/V+NqTw/
PolZagL88kMBLA6upXpzfXz4sQyUysFoZa1KbUqnq+gsg5iK6wNSQInKSNjZ
dXAWeSOv/0KU54O3BSd/TkwbKeAvWubK7bJseZ5xOOlFeHalSQtQCshryF0e
y/Ye5+tU2GbuhKyN278fVevUA4ufeiUfnKNuXa4Gb/5Z0BkF/5WRDePnNOTi
oXljfBXpZmUN3bysiXbjBYw2TIQG25/Uwe07omYQrJiVfBnSdbQ97EZLcSyU
hIKkrwy/AoobVl1a1zcoqtZ7FJEBpqcvGcC9ru9wyVGFWyJNZ+u3bmKo/dEU
riBdyNS5GvAVRc0uEf4O6QBRmP57VphiStaUcV+uh7FyCMUO75jll0/0Q3e7
AmN6GzW+wCqGJoXRjHJc3oR8vwvgfvvc0Taa7iqMolxq45JhD1M/fycFD926
ypBI9VyMaW3ya4ptzp1AvHec+3Cnivx+aePG0R1MK1iTxFzTsmnHkJquRtuw
qTvYhvtRlIcGu8KNW6jEfWtzGHyK+Qq/0PgmnFJpdqkO2YOifXEbr/cRVEH1
uWCn2ivohWLaTF7Wkvreakdk0O6t5reFfkYMVJTP+hG/ZuHu0a2epXYSbENH
YrFHnSGwoLSgLLQ48Lwn0lo98MBTfVjZQfQdxmztnh2T3uvZWv1vjTLUc/Fd
xEAkXg4RyEJubmUr1wu7jNU6FrNOkmFZiX71hUsOYJh1Pnu1lO2TCpfTRBKN
j0AgW4zxulFYN94W/uVtgbqp1sugWn8lYZs7064ojs2pQpaJlcyhqGnmbo6s
NNKCpe6CV0U/XtkhiO7kvBru86SrRX7CZGtNW17wf22aPnneE2ZK+qFrK1CX
CfvLitM7sguhnfCECeEACi4FaoHPdq2yFVFcevsRCS1Sexemb3QkDqmZ0k3s
JAdg1oaM5t86036PJPm66Y8soRg71y85uT64jwRPGjoEVSPPPUJZule7mh50
4S+OMsAV0O9MvhqWAIQBWDVdN+xAYf6d4kT+V5310JoWLqsx2tCR59zDSMb8
rtpv7Tre3czEKw1yNO9q8w4DpkXcc2kfeGyukOxsrgaLaW4nEpaYUt/OIGf1
/1LJIGkdpakqcDgXETpnacfAIULtr+jFX0irqUNd7X2GWyOyzgsSgvMCtk3F
BaLvcE3uujs7tFxE8ySiH+wpW4flzkOd3c1rep4f4jTdkg+gbRGtQQ2ASQ9y
BjUcnM6YD0sr8DJiOD5p/gIZ8rTABcyk/pr7BCviPXP9D4o5Yaygx8M+dXnu
uTayfm5vmN/znV1MedMxnB9AtBazvsSJiC5CWHe1lqUgne8KpIkLUbSERsyB
k2/a8KK6TO/YFuVIfV6o/JYys/TzefIU/D/shJj/XvNgOaQug9PQCr1/MMcG
wX0f6jwv8ovRIF/3QeKCTSvHhBSVDcpB1+lfiehaWVxF++rXsB5k3IVem/5K
smoNxxvduyciNdy/SlVd5l6yUIiTINI/jo1WqUI7632nYsgg6PmUhPU1DnPv
GEAmtrjb1Cqj3qa+0/HgJHwy0sorF3GkgjDizOQ6fnM8kQXA7k5wrHHvqvBW
cT7mGeV6cWON9oIVur2nYAwuJI1oIPUHrJvY0nCfrj7fMbDiZdh+I33cVfUD
VeuoKSiT4d9qIhvHbE21HUjOz/C5EIrzICjSB8EktxSWzmo1bSQ+b+0hoXBA
hjiqYKldvf6yRdJthCppb1hzqDjHfloDIusyQgRr4ztBqchVMBDsFyc6cPpI
Rzq0Zd+KZeOy/YKY7LSKGhlaFa5v8C6hpGiq0dPsV+LP5BpzQCBH881oUUgr
QLtperCTbc1Yjz7vEw+oVk0gqCXONueTYuiODCcAjTFB4V7U7swc+dBGCDTJ
ATXBQbZcnyzS+/Qb5j40iCHzqQmQn+HCmoaMk0wPELo6EXamUSEbqo4l3F7h
eU8xWxNUn2HsBYGMbGYXFAr6hxKVwpa2LM2WUfPbTjE5norqBvpT/4CtcliZ
ufNRWHvsmh9CJWLcliPlsAra6jpXxhExEWWHQ396X03ry9bdE6FjfSff0KI7
HTOnav/QeLn06FPo98fwWsEKZOA6fEZRvcnLE3ZbDKhkFHxVVyRVTsl8t9ZF
zOrPRpQcet81+habXHASshb8sLqzLFLsG2HNwk6agJ7jP8WGPvFjTr/n+oCn
u+b/4Uk1pupPVxMiZtKsNX6OIkNSixwRvDtgeghu0O95WV7hDcVUiCefT6Bk
iijmZwX4mLYGbWj6BqC3KB723uvQMC3CD2DrIr6KUAD10IAgGCTNeJV2xM85
LwvhaSMoxgNfLj1N3u6VqRF15vxIaceI+iTUixynynDGUSPPVOB3vHaIdJuI
/VxEgunjnh+L9TULtLTHenKKqQI9vb35EZiOadJmYEePI5oD3WH1OffxNToF
7jdI+OZ/x2nQ6tvHKHbCWlOeZNkZidahR2lErHEQoGr6dtPnUWn2T3JHjMOs
dddAOGT/WvgibgJ1FwYs2A0AwDb3wbz2qYh4zJAWPyvMOPm2DyAZhmAVwE9D
QUkWtUYp90sA0Ujb3QUXzj25MiblUINxTBlrow3VAtl1NiRENm/Sk9xsNOy8
K7CGm3MHuvunuufcUYTFkjx3s0rtqRdZRvo6bxQ6oToQqzuRNrTocPbfaDm7
WITCzuLd9KKOYFyf6tBI+ijek7i5Ii9L3WP6LJksd0knrHgxxEFB7+0mtWLF
WCVXfWRn72iBREoIl13D39vaqVWuuTR/KVdeKSnGjTX75QHBGfwTtHTq2fcV
oykSq/oirf9RxZOvTQudfX4zEuxay8R0d4mBAQxU7IIjV0XkHBpwQi7BR+X+
3OLw7U1GCpxCov/hxXCW2klQobIgN4k7nQWx21JJ8wGI+2pF0aLkPD/anLZJ
z+lKwNwF5G5QYnCUgPJqBE3zNLMUSD9hojAcr/LZafLh5burPa+x9T3g1NDf
qpywIJhmV70IMMw5MKXpdl9RueiqFgczFunMNhHeW+p/wMQzcc6F8OR9Weel
8Or5zteKMGM53AK0MPrEOOOwuGFImYID5uQWn7RaKW3+58UuhKKTZGNO3gm2
Tn8JyKzc8tz1o9rMDi3e2s9RumlnzEWuCoILS8r30Q4i3bdGvtE2jxReIslj
Oyp8yFu1HQRq6L96HLxzJ6Gmj5TQKxueULE5TqZ+hhnN6bRJiRUQ8j2OzlkI
xBwSINurIIzx0cs8yHGj667cz+GxWmkZOkSdrgdj+Z8fX0bdAVMirHSmeHvL
CnIvj4ZldI7N6m6v3Eznpjq6Nz1M3N8xjCWCQ5pa+yBvi3tdy7mJK1CPJeEl
G6YbMHUoZR4MUcWB0FVyL1MAj4A87lYQfG+DRCX62eYAdZHaeK/MTxUQETWN
s2Z7Vuk7QebBYUjiHxQLqkkWKMhgoOvYZE2cvp5vCQwD1uQKPYzJrFNzBWax
WGXJQhUIAY+Wg7pCzcgVp9HrjXPI9Hm3lQqVvDunhb5i8ZsNfG9higX7vJvn
3bnsckWrYD/PnKjanEcFEvAyophO/6A+jVAZWZ4L+RBCJOpdVFAnr7hDVqY9
qfbFuzO0a0AU9C9hxrteAiWA9XaealZkVRdayoWRs2ivmgy7tJHS8WDhR8Lx
2dzbzCDFI5odq4uQJhuPc1FXrcSc4j9e26wqGu9/5pBAJQZHfrfPfKNv9rLJ
33lcaIsecRzIut55ri7yo4FvxZdbxy5QIB7jccnLRuo1YWdTVJsPSPv/NoAP
kZphNTcNfpv4TLiqn6LO4HnD3LGlVM7UmKWxAa+jz3vBHaxGcErM7UUUCz/W
QB9T22soe0ndy3AE20//DydZXqqMwInyJFD42JFXnMAInMLP9Mem99UzNdXJ
XssKuhR/O9DARJgyAZylzFm2Vn78bTEMTxnwaO6ppUJ9nC0E6Iq3kT5aAr3V
92cixpBHfAk0PClJ49LRAh7fGT+Ib7+BsgdaGsZR94F+BG6eTaYFVxoTc/kT
BdydB53pwtBa7SwgWv+wAxnBlN3LKt3WnH8PRnbTiONKlUix7JOWHU4MacIR
7TENxtQMFCum5v2FXny33gYTHhmC9AuJKym6Pf6mdTwrk1y9E5YJhsXW6xIr
JHqOdU4q8gZOyJE48iXSazDj2gFe0kTobbk2Bpwo2CwesufC3beYowTE5eLX
LtmnqcXBwpwudfu5RuDIQ0Le8WTvtBhATwfMcMD5yhocZSePpMLbQ0FFvra9
ztQOMBIRCcPPDXYSTnmiJlBmxNNeCegMryLm/YuPquq8g403IFpZubFMfn6I
n2QXfsx3HUXmxcntHjkA3aOrpHT5Va1iD/2+am9rXtrIixcsP7lk5EVkoSte
kJvovTN5QKP724g7a1iQ0eq62vfi1C+jF4hevGoXnUSNwhB2Pv0DsbPhc7kh
IS0F3j1lL/uB0XE9ok34ZpllY6GzkURZSsA1xhmi0qOrwEeaLnRPjdypbxpH
JPcB1ZhWDLsI7f+TaTJ1ut8tqkoVBM0GorwLWwibPtHdeH4tg766uCGhnSpp
GCy+xeequGOGzIr1FjafcvS9OMcnYgpeYC2SMk/CPg8MW+flfa+ESU0MX+Ht
Yp0F+OmstUuLLxN8TTTi7smIF2hgM/a07sWlFlk523fSPwjQRDeAwkutSuce
R/E9eqZLHBM1LJYNz0tA9yi7min2ahf5KKXVTXzfyN2fLUpJT+YfKxxBpinq
7gXp89JjLph455ublDuKuXtDwFTBlXfYXKRxyx6b9nWwxxNHl1iA1qwSFsI9
/2s0nLXKzZSBHQ1skf9hTOLcSZV6XHKNl0Dfjfiq6vZXBQv5gdhd3aLUlyGt
RmJ9wv5EMsgz8HP2VcHQfzYitB94NzjAqQamPM42rltpmhUkAPC3ncEbuGGa
JyzzwomWTsbxX0sk94Z3huv4S8WIINrlheG5IqvRDPPbLP/zcOj7ctrRgqqF
YLuXv0vVge9395p1WrHJ7MbteL32QtdFPoUiZL4K1qOJVNMKh/0WfbyFKBqL
fFBXs7sqjHK+Sa0lFeMS3GhB4jx0NpRUtEkm3y2oV7XxLNQO1psdZAYi/RhR
51REuWLKuHpb4Z8TIT/NKG4i93VFY0u/p45qpqX9JWunhc1HPGkWhflkXW/c
/ejjq8RQsBL7moK3owr1Ro/SkBxRc/TNWmIQKT3DXtlnhEhvD/rmhFPfBhDT
PUhvrIDKOnSBr09HCpiipJ0Gxk9lWceDjJY8VVV/HGsuRBLhEUz3JBkh5/Cv
2Zs6YZQb1otUm9EY6GVRWlC/ch7KC7r1G/lQpcqVJ6u3nTk5Rjn2VmER8jRf
HDstDXc0ZVfg4KdNW0q0lJbSp9kRooGu9ggJ67r19+VRJgGrclD0rjohPnoV
nTWyfcMJdPWIBACW+LAQ/ET0uuNmqF0KBmBE1ILqTcYmhgnN5rXyPpb+dQtK
PJA34U9a/31lnsBzJrx6NRMiEnzwhQ9zBW6rVO4Uoi9DzGTrQDweq2SESB+l
RQwe9S7MZ6Ry+eA9QibmBcLIK0dQNMnKLC2+1mxE8v8tQI3QGYjPfRyVl96z
eUbfVd36N2MOtfpjuNS0z835waHelG0u/Os4dwitTnweESLzXM0mSgA0YxQk
tO6hV5ze713ZHhTEEcKbt3NicrVluxIYyVmeSkBLRIhihUcktKgbWT1X+Hif
7UZUfSS/IPon7e2GkXgW1hDGb9g6LzRSnIUHYE27ebcjBxEuHLc1ShJHWYXS
sA6otrIKzbHIcgmlFnB5RlFc+71ruWujQzJ0NLnhlnh9UkvysXnZGl14WHP3
BxRz85yJsY2dFCE/g65j1TBLU7/MrLwphdy5uuKDxOFYsHLwpFL5diRbHBAu
zy9N3ucAbhqFoUja10QAmHI9dimc+tVGb6EdbkPko18809Y/FuS3kMIr5TvV
551p16YzMWdPVAK9b+brDnEVjMt0kJqtMN9OP/tkl1+Zswhr6hg7n+QJ9arg
sv52iFjmvFywGp92hkO2cXeG9LsZ8vxXHpOdoQ5YCKatnTI2BHLoSQPcnqX8
Cjk1D5yKVgqLhU9ePw2u97REYLfBeFb+3iUanhGU6FMDBHaBEoHGdunSAW2G
KtIBGljyQP9Qkcb8dtHIBvkBWGuOlqtZcLS/2oOmlDr3p7LWSDuVVTTS+gWH
GN/sQVNStDzrIm3MQc421LAQGh5xQblFdi71ibcT3aUUiUBNulZ8VbGj/U08
OSd4xs1yPlKrsrBVOiVjJgvoD2yJJxTPpRs+2c7w1+5UBOtEr0dmSfBKXxAP
lRH5WXQRQuyPAWpdgQa+x5u7dDxeKwflFOE3LsiJCzHdVQbsxUPuyrJ1jm4w
Vje5CnNlo8AX8fmIUpMosnyGi7ZZug7R4Q1F62x7IREz05I0vtDG1vRlUI7G
SYJb5fDlNWkEAgGx6XFMKqTrFbj+KtGTMAn+glTUGLFXLf0nJQPaNWH38H6k
M3FgHIBo2UnUcDwChNjYGSBtS613Q0Zd4Qto/Mzq/ECrZfO3x8DDm4SED4Q3
6zPFTviXzljBQWlBEJTVRtuqodnbMPrtAue6rRg93RHQtTAjNNFxmNML/ic/
FX8IjnbJ2AxYbamTcvYfh0DD8gjEa28dhafebTTkU8Y2rmIePifE2VYSCxIW
GwImvWATe68rL5h5zIh11s/ezW891xbzZxkwCgTySpB3CjLjG9/v71dDEUhv
NerKBIoWx7AWwxEPe9tUutIgJo3nMs9OmZYHRXXD0mo98NraDSHihVynmnZ8
lLWraYJkCNBiIoMSnMy/xJkWahDqki2gRDR1PujlxwCy1Kv4ZuE5QtD9Yjbz
6qUEsaAg+PpoMBdBzPgBBA3Bxtrw2n1hCRP0in1ywpoL9hE3FU0843iZiJV9
UgxCnAlcqSYqtaGZ2QV8FBcDduFGogUqDjOEooJ5wEkGV69bnHsZsex7rw6l
LnTbufLrAzguWpuau20iJALFXnYjjG/n8LgizBXAzayGM6IyZheuz+2MbM/d
FiC7L+//VglrfmdpH4orKFpSe2SJeex3CoIo2V67T2ovGNI2MsQVmbtBf7b4
zI8Qa7Ly8TqnLY70O7zcwUzMwOmXFQESkJCDQOc3UgZeezHUus2R8dYCzDU2
MzrrnQkGR1lpQBZN+MSUt8NieMORWMI7UELEbKgTOVHIuWKLQBAyEI4tSIDX
8l5GMzzVY2gtZ7DBC9v2cZFl9Ofu0ywStdr1WUQXWahA8xjx45troyh2WQNJ
DdhfK1BYzXWdJPup51DH3q6hXYXi/rrM3Pqj9zuXRrpzYcqvBZ7j+MiyVbZi
zDJBwUz2f83eZS5ZMbqZwYPqt2C8zY6oXsCjthUyz4wa/ZeSEOrn4D0PCYEM
INFEK2W09AURHXgm3OTP4JQWbz5CEAgo+1FiiVYe0NxqxpbTM5VF44D1gAHb
owuplvdrKJe+cWs3yJEtXLV2pVqiqb2JormJNpI4YkC9zF+CjgM62gR7NeQV
IT341l0Q46mK+/+gUgyP9lUWC2NMV8teECg/bYxFh18/rAu/+IJltnFvbsr4
NvhHaZywtz816SJWPQwn7Jv1Ab8D2qhmvJQgioAgCqMKZ8daYBz03yuDmTII
8n3+RCm4oelpHr9c1dGdsEQ4KxxwZ0cyj50yLEpwdSeD547NzLE/pNqZyzA3
TVry9qwB85atnmzQRW9/opL7K3Q0H18MKbGnj8A5fFp12gBqld//ZiUWpwkV
yrPfbgBgZFtLJ7RNFTuFolTdlM1XxFUMymsHXFG5VQKxT42W1W5tqwJylMzH
BvDDuYQtKl/mRt9g0dN+/HXmbSRTrWCxNmxtxXgY2QW3oWCu37vcVN9VysQV
C3ma7HHKU+EkqmK65uvDEXOvH+8omfw2wQZL9XapjpGUB8KzxS9dZ41AzfQr
13eTSFclG84yQsenrOrW/+jFXWt4KgPdsNg24RPdAQGthg1wly5wEyN9DjvO
F88iQosN7Ikg4bBHnk6j43aq9h0M7bO7KiWB+kzvyfXOKneyBubG15IFKH+S
AORR4H43anLBxh4VBmujOoy/1Nab8+QbUjK1Mjf4Ma8rnWEZLGd5q2U1bizK
qRDzCc4yKZDVX6wSdQQKs1+diyNxs1lAin2Ng7fOpaPEuulBVupin6luBTGr
iWEMS91ii4wbVhfTiQUWbzLMPBHYJPVeqC0IAc4CvIqtn2SzhKZ+vkozh7ig
Nc9i6ERzXbZx9fL2XOuso4VBuDZrYD5b5vcxeg2/2HZigQGkSHrdFgwOMEnU
xlplpBcava1o2DtqsdUVk3lPS66JQhGth/+rR0eYiEBCwBI38DLMUAeq3oPR
wUtBhc39A6GzpmSeSltpSpi05PYI0hH4amNZUUCZxFzAbjuNZDfZAjbvrSvx
H49Jku5W6EtCRpPRgfp0lNCDd9q836eVh5BQ1+tRVSu8AUJlWHfdZugINmZZ
YrMeWGw1f3qHBjMJqKtTK585kjf53TfHYN6OHbuXUnaXRjn1ncDRKQbtBYS9
VTo/5J5B0T6aHjivvEYo8Rz7tghNskwgd1/GYFifqj+M/YXhCGAuVivU9DuV
DLBWRhpxmjyci3ShC4ADjmomMm4f2fZ7nVv6tSrYJuOg0on+4VxehNh61rTn
5VoM6TrNrRceHaIYNRy9tOeZiyXeNfGpzsAwpJ2dIJBR/KfijLSBfAqLmLWj
tRM3C4puqBdxfonkViJxUnJKAKTIJWNpFGPPFIl1rwVX9MMAit6Fa4VoQCmQ
5yILZNMPI3AHF7oHwuGWKE68hnwCV65CKFzai0R19LBCYIQVQgekPapY48rU
YnMjz4cGfV4gEeI7jfeeYUNv7ovt+fV9NrWRSr/r14XII8VYeCgKdYk5GHvb
k2DjKnARerUHiX4ePyR6Opwd7cevTkMnsT4CsQKJAuhgayJL42z/Ku7gF0Y6
b1hSncw/uHCi8R+1b+jLS2Q5dGLah5BeLS8b8fZeSsisXcyUhmKkDIuEw8tm
a8O5gq9Q/BmKjfkoZJAzT+XJBrLjHikd7B0agOx//kXtpHsBmoZ5J7/GLqU/
BAWcyv87px2vU7xvk7NTOuSpmaM36OQJdLIi1ivfqQpH+tcAdbHBABvnOpv1
M1sJX4IxMfQf0z1g14de+GHj5kKiO8Hjtn7ai0LS/38XXHc/hMZGsL/DbnkA
yS/bbSvpFiaAZfxAkDByoOBQsld3/8TxH3hzhWfMZmrrRqyyqd3tOkJOcBCv
q5xFLFgVh81agJszIAVap3PA9DFEZflMrKzSVBXzqi6s+lik+Y54xJHBGDH2
NyOuy8OleeFAIRPhfvKggWPn+zCWJvmiWHJkcTjlInnYm8ATeT1HPCrFo2mK
tDk3QSygjEmQJiC6tspScOQrCBHWSE7ene3Yii9zTNsHr4HiM+9dz975WZl+
kRCQVHhGWKW2vzNnhTVZOjq81u4RPpLlydhNiWIAcQlKp+WTqq48W49vG/rB
uSJ0GstalFPi1724f27uug5LphTLPr5dkdAGEcWW6w8YEl4+p8Zp9+6ztOYX
9DqAsajU0uNS6MxLCtUvKTpdfv6PYWIQkZTKA4sMxHWLLram5T1zzeBnqlUV
yGSlSc8ZiJeVr5WwOLXOhpzq18JCMpTXYilgo8IfvMNSGaJL/5f/lmCr/K3Q
lg9jpe+ZQcqfCTY1UVN7kp/2KFVqhIjNhSZVXNEUtJJYQpLr0jJZNtV6S1bi
VCdaQODfXljNruyBaFV4gXAVDcRy73Ipv2ls9XJXkZ7TC+CQ/FU8k24UGZ+u
Y0SQGqrIUXgJZh6u/g1yrmRjqSLVXMt//z01MXHqKL3gsaaL9IZFybCyRCYQ
nElRH2tcPNIJfSwrr2ry17G69NjMp74hzPiMXsFifobYIhc0E9iyIgFAIbfC
8J/WHQ7a6AEkHLtYCMgzCqwDm6zEvgU91QTv1nohC/cEv0wl32a4uEx2sUOZ
xcYC9GvE2abSbXJEwnWJZY48cc/RqMkNRdmS/zB9fFPDYLVjObILbjL+eJWl
BVCnhFxLA94raA+MY0Ku51bx3z/+nAN1FBasGNtrH20P6/5T4M9gM4HXzO2S
XvqeB549PvWmP6WlRf/ivVLlqlf4Mg0+e9wDU9JtvM0A1iffZIsAGPohaqgE
vSsAfga/cvQtJuqqSJwwJJUYaejOz4+CI+80YhSyA2z03SFSQEiOkFzx5kOM
VClQwTi2mO29CieMkavwTHE01jRI2iyotP0P+yuId9/qQdBbK1DnNFuBexw0
GIl/89TRYfgMME+vxaTfZxSq6zU4jDfu29ztkXp7UNiQ2ZM3nO/88w1fCiS2
EAoGsU1otUtxhmrohuJ9vBqRIAFfQ9MJcyWi5pjNc3qFgiP9cLA6PZWX3Kdq
fsTzrLwEq2S5A3WShkU//mYMOf3dMEKmk/5h0LOm3N2DhkAhijjXSBqq/QZE
5fFaNMxucSSxC7J2HqQuyxLOicBLSxiJwtfYE9+98lZZ9Hpf8xVwTEcTItlE
LSseSgHXN2Aju+/6CtFfErd/4zh5jmx+WbU3G+nN+5aub0dsuurEmnEZIY/u
ZO1nvbATLEX9/j8tIs1cr+KxMI8XxlLAmnYRMg5DPEeyWH+JQovwg9X0XHsk
O2TufJmy6QJvUFqNggpGbvQOlcsWJPlQEU2rIFypKTialBiWvjVT3YRBSYpf
WzOqVDAt0oyVSfU5sgAF5hdZIg+IlRoWwV7SSQmNhgkBy7SlKRu/YsW0rnSk
BmhWJI6twGk8KCYlE7rgRn0mD8sQ47ghqGxRsByuoaJWCrc8JxTqZchXyjH1
XJypgAXFtZFAMsjBtUTnlx0cZ7hfnDtAVpM0jVZrq56G274C9yYRNm5tuAJm
ClJTTgXTckqpm9uaLEt8+ht6h2uHkLUDT3dSlCuCisJHHWfjLc1kNbe/5d8i
4K06y/JaILN91v4MEbLS80Hy10XivH4KPw4kriUIe3acjSMy4qttGr+29SyZ
om5j+2p9eIdaqaWJU4d4BVI/falN7iWkTExYGapHdNliZqnvdpmDV7RXzmwh
x61CvdvZBGFfkoo7TtArKmEVH2iRp3B5twGGm9jKDcCmu2Ffo9+a4JvZW4vt
WqFxMrBcg0au0UI0uRY5aWIpvDYmf7pxvrDhk4noHypA2s/fQMqRjTkbaOgA
5ISEHJ7GNMEX5qMoWnLFueITZFPsDzdcS80wmFfpuYK7mljfwoaF8QBmIkTF
6t9UCxmiMc/3nV0Th4yxLJrXVd5JBXSP7t4BCFDPEbAFNFsrAEwtNJkOy5n+
xcJWIOsN+r1PbXTYSMwLLcZULoEsar+YUCfiX1YTwKCutRxsrYfePj52Y0E9
LOZNlWBcikQr+BWQuOCJTjcfKCjticVnxyYzFBf7p36d2cQLbRf9mmh+OhSd
Z0blKjHqE5KqzBl+xh8oyoRTgzo5rjqX5WbOVNig5B3t22omiSPTbSgiHce0
CrPT3+Aa7Fu55v4FVchQ2tNhVgYuReWWO70ZWPpZNQBtJ2Z4NMkIrj8pJ3d/
udD1PRWfJLnG54TYGBVTwuV1zitXs0p8oD55zN7dhE+/1tqijyEnARuzOTaM
QwBmyLj4yUDHZt5hafUJOdWEKoX9IcEgvVs/tn7XmqZINeSmag1M1QG/khU5
i/s5rDOgZ3ViR1+4of32duoKekSiC1dw/8MlWMxfPMOUGNX+stQCMbpmFABq
vNvWh+FD8gFBbSC3tKpED8s7t6GgI6JZEraDj0W1/PSZc/xlZTV79VILM2KL
YAseU/bgL0WqOXkwLxTCC6MMT8M1yat0nBUhmKIZuRyLXwlTr2nufzJQvJIo
OC+rFJRNV5hSER/2IWH03b7MmPuk8nti+4oHhAnmZXVMpvguxok5jjPHUQ6p
Nks7o15lWGbCtybaKWaol2Wu3vrVE9r0xD7bzXxoEX8dVTAI+hbM+lIQiTet
BmjdPpUW/dTQ/nirA0auUCAurYJJzrasF3/ZKqpTu/PABTS0FxpHb0sfgOzk
ABkP7B0zJrUptQRLODmP5o25QuxNktvHbCY3nAN1uxkRdXnVnTmRPC8hMRIj
c7FZMtMRzdZcxiWlyYFxfOWeMLyWQRlSc/vHlba6n4c9Q9cZo96oJ9iUZUcn
yV1iXGd10jmBY5QPr7q9uD3kSxGB2KwzwRqOvlK5IJXY1HvHmNjJfNYDhQWP
FR5UhUbj8FErl94wnC+zFcQPXXjj4GHxZybjwGo5OKTW7qJKz0zx9mLlH3QE
0FHylEw+fxAeQppo1Av4PXts22moEXY9FuOjdU5U/tqUEGxniFpOJVUZhZrp
W526n18AnvB9TbzfMk4mjjFAefKZcdJptU/rpYcdDCF/xXXeH8x23Lgcfu2T
VsY84m/w8+uifKQMN65Bmz+aEyFBR666R/9NLAcmPOFNHypPIE/BNIgUhXQw
Wy8fwDsFnQByNF37eKVHKi/RC8I4KLPkYrhQm6OA0hELv65ODkjZwTA+wGPW
qHqqRsR8LQhMTB3Pf/VvIT1B9VhsqBSdO1fj1ZMp/rnDpdmNNYVuZYF5C0ps
nZbR0Tw2ZDgprQblQTDU6rQGYgfY9AF07jv1EwpXpwKIW510o9sTXrH4LLH7
hnl6KZJVU7JB3R3o3yfdzkZywKA1XIl8f7+3Wden3Pn+fD0jZhaFf0gotoVT
hRBOLze3eV+c5PX1spUhiMbNkG+TQ3rJFBvICkAhiCrETliqn1YdWtsLFXek
ZhQE209Y0jTLxBLGw838ZjySmwFm7x697wnBLkd2lBsWu5222rMlJQVHRMMr
UbY7wMDmRiBK5TVfxUcmKMWSvxbCF+yCiB1oTzSXkuZCsKwRYnoAPdIXTPAj
2Mtppqa9/9l3mtiCfxv1XMLXZeNu1dRW++VsXFXH7XPmg9irSIHDiFpTAinu
gLJJpLgIhiI/s9zBlyEhfda3ayA6corgRmL8dk1ttk5CYBvC0Zx2qNdB6KFb
kQvbi6vajNl1cfTbZDZkKccjzaFIqAcYcvt74QPqWxPzPU/8Y92H4USjTP6p
yxlg/uecllVhWy/tl3EUr6X5iVLbPSZ5y4+RtoARMHOQIFgm0GQf4ZQLgwX2
nlrQ23GoLYEUmY5kFG2t5uksW+HhwY6/AmZuj+U5uAsFJGMuB89bzKi4+fdM
Db3QXJDvzjHmR5NMa9Y8GkhuVCU5NMf1jFXCZIc1f5YtEPF0iVSqZ/I5SUaY
5UhpVj+Y/p8QU46jnuloEs4/TTP/3fzxJhAKF0W8dX+RGx/g1EELgkNqgzX0
OYKeX+gqeDm7hFbovLqyx+sPRxxQnVzhES4kqGhu8aQ2ORGXDgzZftL7zRSo
rpi7wWw3b52pGMYEdwXm/NhhGf3m6aRHbL+zBE9FyyisrF+9SVSp6a3qnXQn
VmHKyeNqnLAviO3RCVs1z4OrRG17NQul8YN0f6rWJO4UFc8yeyzqO4t9gDxd
CG+FaAho/ul/XAtYuVRJQRuNuyRypxPa5hs7yl/+6XhU6svEBkB03mgWJuIM
CgRaL719nHa/r7ZCBaxsvPM0ijNeEr5PX/HWmSh2aVl+ZXOe7LA2VjTN4CHp
B6tfuKPza6lwBF+DTq/a0clYXKfOJ5X4Ni8fcoF+0PVZVSRy5AadZ14lCg4D
8CP17e6BXJzxzFd6KNdCI/IyNC91cn8xZvpMl2Qwx8VvyBeNw76LZvl8EetW
JlWfJiVmgPzafnF4ZKR3OHtX4jTv+xUY2eyDasHxqjzDxPqObOKbc1/KBi4J
fSwq0hxiEE0jC8icQ2LQDVqw9WCmLsTL1TOdPvVdLwa98dwN7ON92ETSAZxM
Vct3dcnUve/7vVcVYPZYjTi1R0o+Ox+T5DGq80LSiPEk8jAMCy2U95TmlhoM
eH57yFiVjQKG23qPoDXPRci5Q0CB2F5TNRP91H78eI+jG60FORRiqS1a2Eh3
5AwQbw/XiGKjq6ohHQv2GxPinJUOCiW4go8yILn/XqrJXGIaQvRppfl3SY1J
39LQ0aAiiS0w3C9Ju0SV645uGnm2v7f1YAqiXTNcZLo96hfkGRFCNL0mGZtz
23OfhbU3c/OCbt5oaS2YlE2XHRqYanGgzV52vxD40L/cJE8ih/RV94dx85Ym
RGbE6BhBGHT2N7Q9mVdnPfEPFpCkq+H6+s2W/ZO3i7YX1IH2JuQ1A9WpXTQ0
zRs5xZBmWcegtXOVkQmr+DYSXSIZlQzeCU3k5UD89CNG5dy1co3Xk4tR7bBQ
/6eSeg8wSfGEnEXUVd5yFvIWBxLluYTTKWm7YHXM+qS41K6ySEg+I/FpSrqp
17AI/FaBGQHq8SVStkyHcUKGwwipPwiiiHjMPLq05XB/lAIyn8BbuuMN62G3
kyTRf7s4KRl+ou5FtW6YfTd1LTvhOqjk/3s0eJssQfzh7de362BYRJqh2TQJ
9Fkd5TD5vvDPTBKRc2Doi5uZWAFuml2mk60zWMs9NNU8Kfh8k76b5ttvNjG4
tKT+M5FlLpCH9pXqN7/YJUZu0JnJ1NqtzmXx/KJ+JcjxlNQargSgDp/X7ow6
GBTaXSslrrhM2d+19hWtBAkkqPOWFwxg7XnDkj/zKOwSd8wKDtK6v/8z5ZWj
JFCRaFeGyV4nYv2gaX30QDNHEIEncJhiZDbS4lJ0w7CU3enSfxCQr20718OT
m5gTsM8epr/ztwCoZKBmdocI2EY35xy+BAeSl+FqpKBulSPQbaTJt/JtwdRy
/rvIOV6JTP00bFhtIahrEv8NvN36AF4DtloUSCNjfvmYzXaX2Of2T28qLCIk
JKKS5AaR0K3240fzV0LkzseNXLDzfkZ04YWyY0O8s/X8nZzEHYfU4oO3H7Ch
UtF7M+iJoQr88mf5IaZi6nIp7uBcAGCfbpmp6nhtC3BadiaeQlfCfUUUJqSV
RBBBPenke8ikDSfN9tGOvlxi/IBazZxeet990tRG3qfESZeetvPNwJ9s5115
3FVlblajGF+SW0jS52wrEz5lO4XYw+uVPsFdRFjfWNy1jCqAhSj6lQalkmQV
AR3gUICPJNQgdejgt9Xx6C3Wb3DOeplNgXetS5u2zU1aq19it97p6cKh2DFS
Qc97FWCSmCbN8wqVC4/PfJY3bVwBcAXDYq/t1FkrtrJ6GT/b61qifX3H2d00
kS3s97o3MDaJv0YZLfTMUdVEg10BPIxLoJO95mS3f3p+vq69GqA8UH0jSTr4
itKSERYoVHAkwFxioEeOFVn5C55dWAK0mOdI595tLhQiRyRGCviroUqmGwGA
C/y3uwmRVJiihxTVBUPhOZxjtlDC5zJEcfwLcx0I7HKJ5aJRiq1KEjhgVbq+
N6vdey0NoHhlgXZ7wsda1Cmv9C1Hao/A1VX6uO02EqoxsuxDIIWE9HIbRQ9n
9ZBgafF17uMwwo/wO9ofXPw1JxduVjH1LciBwcCbdEmH3aS4DV8XhmGAwL5h
0J+p6JN84yV8a3tX2P3ZYIOJm+LlqzSFnVUF5w6nwrHDe9Ssh/6/SV6O86/I
jtX26rqVgYYJaVP7I1dS8oYLW46CsHwpS3Kfx4fmLbDjoCvXemkV+6D56Hli
vNl1cuSoOQeq+cRH4i7B6OgK8Jy0mTq9dKMYkD7x9XUjz4Ig8ETzmtV31+KV
FWZiYttostr7iOMmggvuaFvCvzIn8U6uNo24i4TNiiMtg5mJsvQMJzwsyfwO
+eG5Vyjwo/REA52S4P9Gazh62Ulpp4VhNCfxTkdtoTfax8pBohlwd24ugZ2+
R6DhSLcMmTPCZfwX9RNdTsHaonb9bzi83lkO9jNem+LSkgJusTShjnywoYTd
TwXEmQAd1kk0GY+fb+B5bAsgG7TZa6nDgFz2OCkKfN/UvvZHPLr/y2AnYVx+
tODqEyxoYGcm9EmAefjlQQTnNoy9ARXY3CsG4vlN6rilBmvdjLHvB23ja9A/
bhPFKu7Fa6ETGS0hdKbTyXwDH5QVkKHRcQDLYARGwrcIriEuhN2y6nTOrwr/
XpDchMv8agU5t9tdpBghh9KicefJQayhHCRXU3rojEVTahLVi/q7y1fDJpED
Eeh4PPxzDtq7le9EbIXUy1NrhYFL5DQ7cpNz1P1QDNJucwgCnE091ZfZmnWe
iCK8qmWChElAt5Qr+IgUon/+d1gn8PjwEPThyrn2oTTN5UWrFG1HcplyyP0s
FEOtc9b6jrrVtFUPbD6dcoAJBivtY9cL3bUUUaWlF40L0+UIocIR844zQAaQ
fCVD4osekzrrFqF3zttcLryFGx1IgUDXtlnZ3sZKFBAspIb+qeMbvv+sk1Ud
lF3fMYyYr14sfdVfKTBlEh2ttQmQx3Zv3CGBAKifaZJbGemYDvvUKWeqc7Um
JzkfS9ur3lFGxlDXgrhbIWymeKjwOLUsysUK+la9O8CT2m2nzh0JqIUHRU3C
fRa5+YROFzuDVYthZFI9gm97CVAJpFjRqA8qehzenoFD28Ji5RAbkAM7ZI2S
QkhlioaOEKzMqZ7A1+SN0e/vy2t8xzlaPQoYnfPkNqUgI9LrrIm51G0Kq9a3
EeiXjv1vHIzJgh+54hlOik4TNVwUs9lUHCwzpaKeBTpzAXBdY9lVFZ9QeM7n
qbUZbeHsu67MiLT8doZpsBX3BX1UP8V16OdLtckEbSfMBbgFZHePOFFHhRbR
c9tRFFr7uAxopzxgrfuRUYkyp9JIkF/YVxnWXfO+l7jYXWvf7LWgOJTb8OKs
7mCGU8tdwUebyej/7lKhAuoLpbl2COKYI8ZhzM6jFRuEusdKd4RIykSHh8ow
QKAW/vjJfUbBN6t7p3NiUIMZP8RqiOVMyi6XqYzAWQmdpY+G/6Sr4cvJotaX
WiwRrVCu8LPgVR7HGBlPv465qbqJs6HfRII1CkK69NcUdP33Vp9nYb9uiDgN
jzt0WvdCGPyv7PIvQIwB2rWB7bvzlND9+3pcsprVgZXj/pUpOGnx5+HyK3zc
zHPJqKUL+fROOtIDLQulmD19ZDbEGDuLrILp3U1E9CpTbl8c3IW+7w2RhAoi
qndBtis1U2CivJpFO5yLuI5c4JAWtfRRc3pOxzzWZYQfY715NnONL/XZ4dFC
RepC2wO6q4Y/FQwzy6Ilp38SNCpaId5CUaHWaV0wKgugSydvMlusSO/R3/a6
f91N9cEpnAzTcGjwnTnL+1hdjYu7SXLWjihjFd3xCPBMjt+0QRdDhYECJZZE
R+DiDaGPlS7Fun9bXNE676WVflSYrcpXDz1WRgRDayPxCwq4pT7Vf9xznUEw
WQv6ylE0VYTfjkO5oLyeIxLSon4rITTdyuEuGmJFlEVSNy9283wtloXnEXnt
92WFugSxZaNYNxBy/60rZmzWOuA+RqIpX/ANDAklKp5mSR3K9zmeqSPQPpM3
aO4QIsou4URgvHVxEhdqYvhEs9p0hokSzfkii1rHmE3goOI0to+XRI5AzHGi
Ozc3Kp5TFbE9gBanZrnmX8YPe9CYEaLzJR/GPyhENXhUApsNHcnt98Diutzc
PSVhMIq0RYgHWJnTHEIYZJ4yvDQ4EFsjLJ88hRCt+gmkfnzjSubqLlSeP0+G
COCDrIpYInBoZ7cXg7c1bRBYvXQOTzshzeUYtqFG6wSlnJAXtH8exJUCBlov
e5WpxIT6Gn7FyOBqeX1gWMudSk/QehJ60klWAIXjl5AgszQ0RfdPmb6EI8Sp
sePj9rPer6cWoYzxgDMpnhGGv/mKLKh7eyYsgT6RlFjc9FsNmCIWJa9Lk7UB
nJWIdARAe5E3eP8JI256epTvVTl8UliVIvsl7DxzofUxOrn9YjbY+CZluYBP
bHJt/vzIt6DPYb0OGob1+jxxVuQH700M8uO09M+6tOeBqDLW3CcWHVoF1BrP
mRp1jvU1PupaRnlQX5RI589QPmAcfsp6YIdYHFRhOYXPGXPQVOPXfodQLPLp
oMADilQDOjOESgc1RhD9WjPA6G3/pebCj82JGjYmt0wVLr0kr7IJ9vD01lZP
xQfWFAmbXXCoYk7Q/M8ecjfS5aLNO0TqEmkc5DIPFcQ/08A+XhQ+CXkp4aXy
uJ/XGRaywW6YA4LfO5J8ZRyn+Z5z6xon4x8N8T21qWuU/dP0hqc/bZrhUqF4
u4iEwmUaYkwpIe/xJk/n4ddTCLM14LGnA0NTpWSvm+U/QPweb1lFjPTnPWUp
5GKrMzvNDCBDvxKguKq2c9rKB9pFeMcXMkd3LYoG+t6uLR4lb313K1izM36R
kW04WfOddqNDNOOEiGt4dfb07H5Rd5pQH34e838XFiWvXda/R2RsTYYbCneU
w9UWD7iRBZ2GYOw2hQj7Ddgx2URi5AWGuC7cyigsN+U/TVioA3OP7jIYtuDw
4hfUwnd7sh//Wjokc0mj/Nhk96bScBE1KrdA3BSIxUFaO2HaXzVr7qff7Iho
58QN0W5DZ7TKDj+Ie/HFeaNzRdOQLZPIMw5F/2M5kXNZctvCWGdQFx+7D0Nz
RVcuc+Hn9SLinu24MSJARyTHZA9sqs++bk1WfYP9jW7bL2NqlU64MHFOQxyB
0LNLF55TwJdmaB4OO3afguOLtpZ5X3giN2HJ6k+C1Cnc8+xJQ/9DBqLY34a+
SCdFwijQ2bBy/Mz8E6ZI09XTiheCkKMLcK5jMPlllxteKwv1uuss0TihwvAy
BL8Ca3NRxGNcVMkYVIWAVCm3khE9giUcxK8AGMtoYq7JCEgymSBzrTo0YnmB
iEY5Q3S7E1CGpINk270M53ENWqPVYQ+kX4FfXDdpX9vxdltdpi7Tw2wsECAR
BM6eykzhCgvIOh0YXZ+udEiYvx6nYbACSz0daS/ebiTCyZ9huVuR/HhnCNTU
BX3rgm4GZGnEAMk3JnVjkLEdqStQJ8mE2gImCSKaTv4wJmX7qbLfGVVwi8SO
NCujVahCti8iW1sZfxgyOqPmqpBz1S35CjBXf5MPxxLvKq02fNkpPHVVQDcI
ZGhhfk7h7+UPA900EP9Fk2Bc1wbXbSHkvdAL1bsfcH3MKiYLojL76B+eOuBY
bIpIJsdMHQAf/HgPxZyrTbnx9oONxG0OwOrf4p9sngyvpGg6SDplA3e5kzuX
utg1dC1fQkK5Dsc7oMwkz6ATm3nI/SyxFdG0IcXAvCbJgkK9t+qCowfW6ndh
qLYoEsCgxo5lqeFvmanP614ZYHEZiHMCFcjAwQiBH7eGoDVhRcdNfmdItBvs
hI0TJaZwmByZJdkVwAs2T5VRFat+YbVYUlcFUPyYY7G6XpZ6oiguQkjxSiI6
3UvXGtXEVYqLSddk3URTY4qoXNnfDY+ckk3RmtLz2+NGzpGydK4oBHqj2HmX
bR559JyRNWuTD7vpgPdU947czfHxq9FU+iHapL9bjBtlDSoydI2IPvKzv83c
Jwkzlw5gIzOxRF20r+tcnftJE4E7uh72cNfK1q6jQif6bFWRQvlD3vA2xiLq
bD5gPU5h7giuvytnCI0fio4LvT6hwd66UCzRfL0tJYwCRaIYlTGqJ92DZOF5
07UeSrLkGRJy6+bp6XN4UpYaRSi9HytbErznml6cqRJhR5u/sxgOAAgq+iau
2H6fJ5+khmuO8uC2hMCfL6f3xwRkPdcdycZlHZCB9+3eMwxwrnBuksYwcxnw
1IKsAB02MYZ2tNO+uqqGY8edYQdSkci/8WSbQxa7YMmDVLcQqEa+pY/ssOgr
kUFpitH3Qo6D7gsMK9BTk5zef9fmM/bW+uTQ8pH161psieGVeX3BJPkuohmY
O63vVcwFlLNBCHTIAYEcq/I/VZ08a7olZXs8xgs7d2urkbEkKlHmtVruTrCF
oz3DShb9/Z134qL8qOfGqE71emWVusQHp18ME2rWAy5LbNDYuJCIg5/Bq5fN
L00MT98XPcH6InR9RwzMPiAbWrrnPoV2pYIVoFjK3npmB2zdDiuOL4Nf67v6
mGgxixFcgxHyIx46X1EwFff+ad0JX003zdgWqUUjbxeB/AzQWx4Xsr2XUG/1
EccwTYImlWpjvdeZ2azgJcyowNsqlqPZ6IUoW2SZf7rluwXVj6jhXpncB82I
zzqWv+YrktZGkU13PH0dVyxGnn6ujSe8mP10vyqU8KqzIw9s6BJPJLgCUYFq
PvEaUoB5u5At4Ebx3nyc7Xb4Cy4dg/BCniC8/fIanJIxasa15axPnjgGpdRu
1lTJIs0tHtb8VEsFv88koD66GogN1v8HySbCrUVuaDP/ZSBEJDQT70X//tUX
eDtL8YjF/FLQzjDY3Hi2FWn8kwWGYflIvTBN5hwymSo/lJeoGr3uufA9ZNDI
LpzmkV5TWWAnWa3g2c5Hk1hreBISEcN6ygwB7EGCjMYqIIcCZisqt5p5S+Ac
iP6NatxGlRyjkrarN6phmYrr90kuTK4rncCXuvht53a3sL0FUUfgPtwJSKYx
6jLKFs5zcr5eJZ77UD04tvSVu9NCsAXbKJF9so1gSOQy9oy5sWXRikWD6ujx
I6pD4VSk44Ox5PnuU3E2SM0oa2klLegfiifmioSKlmL5LhStEQ+4FzrR6fTS
HK7UKguLkosVirLeZ+36ZRzM8zMyNa7/b+vcLEvKQVSBYldXzbcaWI5+kwEe
NA/Qjse81fPiT+sFlPNIIxUO4EHuMJxXlVbdQkPhpRthFlPVCpGrijxDNClP
Tz02FFSI+tA7KZd+RddKbOFx+x5MiSJsStcAl5CLOE653jSs+kSuSx9mvka5
d0CjGt8Bx3P3ZR/65RTugnr/d9l+qee9mxqRhSqSb+CCHkH6aLDpsqEcwusU
XPPLhGiVk4HNM09h9/+Tuvk2gSQnyUXwZ8j3PYoFGp3aPH5fbSh5fWKzKJwe
mkr4IWtweiI5sG8lUraWMPRnz2FyydvGTi2BzwZVwc2IL8MURfggrv9xP9Sc
/ma2HGgXkqwHRG4S2y8JRkk8ACJO9Sff3lOmCUfPJruPVSfQ3x0CbarXYqoi
rJEEHcf5wVd6Kj+FaEx8oX5hVxKhYCr922HbL74jQDr9pdcmIxjNhaHNX33Y
/NJ9fF3rUgEEGqVktvZqZG8vq5HTuN0EX0nExJyo+mlmg/r+dCXe9WYlC+bg
iwr38gD+jWR2qbClDaIGNwKNPzVxk2bhgtJrJgfyFrW3IK3+eHYHir5Oo+C0
b8aXx2Z+43EZE+tmaeE2BRkvj+P7KDtp18yzHodqC5D/cR3GSydnEyaPnMSE
NgBnAWTAfSsQ3l3KD6gWp5tt3yINLNNEGWn3FDhABH8pr/6JY13vQ107I/YU
VbJV+0sVL3vNdf59Wy0kF0hCza/+wMToWhHEdo9D+6tv2tJ8lr77TzVJx7f+
1X0QBd6u6kMbu2qPDO88S7GZf+CAfkbm1MEOIu/6prV06+tb0AKdo157PuF5
hVH5aELR1+x7j174do9mj3MRtT42e9dRTMv5XaKo7btf04gw4T4sLIdGBN5U
X2a3xRE02FhBo6hu2ChrQex+eoFE1IiBpYHT2R0MyFm6Q7cvye5jWYpN2ojG
Um2mr0NA7XDM6KOggsjxEWOZtDy9c/LMJG+A4N6VpvjWFJHiQp12FJO9yQS7
D4KQuJKN/AuoJ4WvGzi7dyCzQW90fxhP+hFt1VQQm4fGZ7ADhqVX2iLLE6Hm
qpnwB5C62+Y21d9m8B3hmjTAdHd+w59UQ9QV6MKeguzKj+3fiv/yzZrOT7g1
lC95PB785bCetyxVMxw39TXsEhJ8MQVYdkLwbPxcNCxCjH00Z963k6ny28O1
/hob9sSeOlV1uInmFG00qLn58IP7yMoGj/+vWihmWq66NfarYWgD4Lz5MCSe
CkN2UOzEbNfRv9eQqEAc2ZkiqzjT+4N32R9u/uMs5uO6+0AMhtw+dKGbZ5KV
tKUhYWGgy5ouSGpkwAWhyDW682/XxBT7KQP7u7cTow53+AQZjnunKlMgPdM1
Aca0Z14qv4+YeVAocIRw05MI10wCEoeKgNok0H/O8jH9FlEVNb0E413Q/xdP
yLXj30rVMTxgz6nRiQu0sIW3ckenRYNhBFFJAFb1cD6YPzk5cVQ0xubUcOoN
gJ3lCkOyXIeDTaRUCjN2CevLTx78IPBzKndRelcByvdq+3cUkHl43pwczGzB
YfhxQuHScagsX099X0DpGVLrMM3Ihb/QkEHYCS3Nysx74WigSzS1ppVcYYpe
p4KtqV6qvuiuyYoj7jetDRS1x7WvN1svbqeb0YJuv72CEoHLFprt6ofhMHOC
812Ct6CbXhmyl2P3BuhauRhD5SQo5DE4YLUXCperm/m45TqfA1vHRmqRwJFk
fQ2kVU3Lp6+6TDTFO1GTFKWoSqpnS6HQUaeQX9QuGI0a0xlcm0BGyhM8tLQc
HUX53RmsRA3ZO39Od936iypdTCdIbOncdj1qIfio0yrQjN/BQvHUrEq0+wr5
Seg6Bs1rF2CVQzIgVIk+iKcq/nJFYlMVXyF9+vbTmds0AJrRoqpuOmtmaUlM
PMiDQ8xb0OsMk711GtQhYcHar7x0Z5PBNVLxih7cdTQ622x6/OKcjIVp+0N1
hBSdqMSGb7DKA1xzvGEux2MWVx8gcTm+e/mnQJcw0xudjCg43B2tFbWpqj+w
ZxVDTer3jiCZ6cjY8pp4OR6St8pHwze88wJBkkU1L4CQwgRFl5eCqzLoRoaO
FLdKFPNjvMwCNQI2muyHIHtpr/ESZLlpYBuIToyn8hi4nLFBj3tEQH2gb19a
nUTVOLHqA76iAsMkzYKsa0NdPIPWfHOjMsBDXXujrN8qDAaLjL2sqTV5ddQQ
OUTYnpdrQ+Girmr5IOrLcLRUKUS1VmI3lbNP0gvDPxoZLeuJa+BLsd/3zi+4
X0nN/6MvhWVvI2dux3li8mIWh7fUCly2fxZxBPIfPjQdPZpKfou4tO50Ugfi
S4bFT5emvNvgSpf82ALqAV0VARtXUEpeUkxktco8J2E3fYmbOxclvKHuy4bZ
Z+i6GMb9MrWMkfsVB2/7B047jbJ3+P+FmgOvYxfarmLTflQ60S8AR27XEjlN
5tucAA5dY6NxdE2pn5iPGflIRPlxVZo4a/fDLEi74pqJLsw7CcOKVyh81CJH
MAKJ8pSyq0T1uVj7KzSNS57Yjsm0yZQKnnH8nV47KHy8cLt8jZ9v++OmAgm6
6UqlB1S78SD7TDWubwadpSnlArlurH+rhViM9ONAA0K1BmPSszJ3bOp3Lhdr
XL9AdBdUwuoVF5LfIISE3o36evBtnP68P6N6Al1LQtiSejX/Zey9yqE+E2Ax
cPGOC0gJ2cAGCMAiuMkHxIxwG018iaCeDYwLyrCCuPbt/9L4TAtm0so5sV/8
AIu5rLn0Ax8qq9KAzl25m7ec8e2LtP5LP8hrtxxryeyVQdDka7InoWpCkwIg
/siDM6NBBJx1MN3Ia7ltzz2jJIEhDOESN8tA+6eeQy2oQ3ooAzGBWfU0OpA4
t94c3wfGtboxfNumV/+ZU5FDK/C6xt8uC1CJU1t2sYDhqkIjrE1FVYBKgLPA
BZclZelqPketK5wo9t/JndEaVVgtRhts0oZNob95lmIA+QgGQZZJHZsW52sl
CSsF/8H6tczfdZdlyx8O7RN8ivpi++NoYEDO4K7gCpuPcuNh/ox5EBlxFWJd
4EXYceEjqwlmm0+FerDbsG1gP0FlgVWgT1nVOv+KyH+Cmmlr8B/Wgz9XeNkg
bEynXvCelOQ7L1Y+AQiMf2zRPI+FAZ7nMqlAvNBdgAUkWY0YZxcBr1Ipgwc2
OH1c7OkomS0ueXxfxX3EiW1tM/ofUS8vOBGr6nUUd+gnjUJAZsIQ1ZajEPD3
jP9CAafAa7fHvToVTkzx0kPXi7BdBCShlub/aq0c4UroFX+l+1La+9MT/Cmn
sP5ZHzrYH+KgO7h90t1bQg2C9NxjgBDtVwv2SNkQ22sS9D1ndZAjlapLYEyV
dxhtmxctEVS+lEvdvula2hvAHDAlymgcJZ2b2dIZySU5emFzjbZG1vpUhhr/
aOuY5m7Kn6nwwLhS4mybtRhF8fl1YqyhTbcgCP31KkxnzaZJYLuuao5NDr8X
fjNfyaFpUNM63mgCBPD/Rln3F+As8SOIVuNH+spQKtjb5Xmff33WUrqeM95P
zeu2cYpfq/aCisYXhN/J7YrqIstekATSmoOMTAVy+IN7fkJUdexVwF7pStdq
IiWaEDC1kUTrzaRcUBwMd6i1OHEleo8bDUn2d0fa121S62V1vOHkm3Z8nPfT
IEfUV8vJVq3ssMqo3V+7TxD+DLgZX/ZkheKHZarXrU3WGahb6mS0CWbauwGg
DwETuwJqDm7M/plp+EnFgYyTS/CBU7IaO003WheywyPw6AllGRr9rnXKydYS
OmDDKE8nGdwzv8BRwyieTdzcIrvTmccy8/fn+4X+dfLJNFeILj78SQDVxP2I
Zh/TL8xf6t8R+Gx/hQp9cyzppSSBo8izK0LJtxqTQOi2Kt5r3pFKsWM0TnSG
+ggJyAoc9148+QiLrOsmj9C+sIaAIWo9OYrH5vWutxT2TVyUsEq+fXSc12vh
4PEzRAcK289TVFqzwrZogEtjVqQUb97CckPO7WUYukBeEQI3MYOu5E9Wm2TG
2lqFgT2y2bby5snh/GB3JPydKRCInaYi0kIBj3fLQT9cRpCTzvCPbrssLuKJ
x7GpHxwKoooAzSqK8YG8pqcrYpHtypayAJRM8iE81xZdn5mPACRepfs/cv/8
scNxx4IqGih38dxNVeKpwBzS0HhWPbHdQSrDruj068JHfpTryW97Yq4pfrUe
MO3O5RR8mNPIOJ+vq9VCmbZcJAcR6ryWxtHz0hfi76VSR7LmA4JqpQ1KvTcE
zq1zpa5SqTkFtBMefLJ3GwAqNELQCCaziSz7oA4nhp5KsJLC9+wUdEPhvkvx
bEdDhNnSmqjb+Tqt2q1QOC8i38zpLJgu7um5ODJQzP12PHvdxsin6+oua61O
H/1rm7IE3klvuKWTW0fBGHsTZWUwYIG9mprJcd+DVA6xAhiqWC4JyIfwZxRy
LNKEKA3v2qHtXgCD23i5aFxooBhnsw0fYEcBr1vsdv5VBIC9Dqf28bgR/oKa
DxcMuJSOYQSt5iJ2RBDXWab+BncCIvxwGZE4L5vK6O9wgHkANMw8Mvm9nH6c
ro32PqJr0YcRCeKJ/SL5XN+XjuWptvmzMsdnFZFtD1sudaKnlxQgzYEcxPXo
IcUUMRG3bGRW6WU4n+Awm5IsENI9JxhgXKII5yrbftQfCVnxxiYDSdCZ0vHa
YNdXfF2T27SYbUcEvSy4rfvrZVuH+K5R+zEdZ26WTdQXAvSZtTXBcatwy6T1
s1eD0YjWB1py+LrcUDITsME3Jfm/vPXwBmewOZZhHWFMGM1PCYdZSCgrqXP6
FuClhEVfdli6jcxGKgEkCNlRUJkIXa0xNGOCQnLwsRtPdLJDixLesK4EAsV2
7rbWp9nVgudPXrIei29YgARQSW99pWlroFwEukDTd2y8JHIOw9ntcsHwhsKG
feLDpaNryX8Z9ZDcP6Y6ZZRSBAcmiFvElP5izwgrxnzay7rHf1OpXxbtAaDw
Lz32yjytRdX171jrIoI3+lEx7pioJraOafOH8vne7W9X1PIOEr2JdWKou3xA
oFMmjcvvVs8lIKShpiruIn6gSfbOlH5mYUKoezEixFB4/faz9AuedYa5LX/S
3IalFyxNokVih0/2bU5ygSzpiBXPbCkcdZ+6nztreXKomkzIeazEmC4uvGgi
vQOW6Yh0pDDZfdwGjLstSmt7Z+yN0gypNOdy+03laU2IXLqGeclNjLJeO0tO
8yWVkZGSLI2j7FKAm8HvI26KcIvYPdpdk/g1BsoW6qSSAfUais/xD143N79Z
ZLosTvCc/cGjFxQBvXQe6Nt6IZUte4iAZAL16sdQESok9ts5cotQsJ47oOVm
c/ROIi6aSLTyjk9VQY0gvA7788myHUBegulLUcyPu/DByGd9Nvb7s/66tp9P
es7Ek4vcpgrZGWNEan6buLiQ+Og29oYrZSw9HVSh0avsRFAmWlCK/8PAjeDG
lEFu0QaJfu14v1fO3j5OgDeT9zPxeFxgEXW2vn6SiOqcM01T3+qV2azaLjPT
SYP/rup2KAhiKPGT7JmbJ/0WCO88/6OqooFpWpom6PFM4mCpgieCW8UeSkwz
6F9QsRLZe5akdDErbhs/zgqdOWl49hBaLeOscH43bSEDLHg1g3H31BdqegM3
wfBpo4vYvBKxFvI6NLW2Q8RYbJZUiYz9in7E9w3PU+CQAp0OvsvvfUZ1GnvU
uBRV3sabKxKEcy/LQQsvZOQrzJVcJdszFWcNiKPoTVw01EqTbNrUfGTVZJpz
bLzInZIjnVwuk5n2FQNRws4jOV6N6NEY08KrvxpUix3xK3zXXJ4dtIJ5miEo
VJM08eD/gNtUzRuKP2XHQZpShAcoJmQEx1MXKyB/erv+4ram1NkwWafLDiuu
2lFMJRL2lMf7WvMuIsdPAnybI72JSsThGKh5i7p2O3lEUYRgbkH2ogv7je7J
M/mlPy6+qVqfwX2gmH6smrgN0wX78cep+mdNZ3xO62s8Ppw8oCU1wcZDthka
mEFSx4Mt18G18Ozkii76MPl8GoMIcksSKAvRp5VW6yUw5O6cENbF6y2kQuxm
3ok/gJnRPKeW0T+yu9ipTZNbe9S/YG24e5JcYMJNQaiwR+nC+iWfvslavEu+
BtPyjT9mkl/BVTrUY+/jU8EaqgJM0lV9NAHYAzoidR/A6ZPg/NtNayV5QQ2s
aijuQUvIk+cXBL64sb2RC793mkHCvyY+Q9IC9uUdxpMdcc9ysTwyssP6J1Y3
RjXnL4TOTjF4p0fu6JvIJGKvVjGHz5UjqtGazjYWq2NdTEuicrjZa0/bUn05
2pyB9YQorp+Vj5GC43BMVAfI+JpZ+uGfx5zQh2wIucdTMMCmktHtPPn1J68B
5Pi70h6UGXBrwmnK7RPRo4iGxCFTpHZR0SsD4dRzN9vV87u9HMa8aRtiv2Iv
Dg524ldXTrI93OhGcfUONZuUYdsVi6fRCpnU0juunp93+VoDX6pOX83btXeC
qKLsxF4SAU89faGyKMTn3oug0JuopeZFJs4Abw/+eXVLhXQsBhkiU2j2dnIY
E/gKkEtzW/sak7v1qldrcdhq0sCMSv5D0FGHrlFfG+nJtJ1Nb31uBfAmG5CX
TeMc+9GqXaTKk1oXsLYpsI/vzeLTn5r4vpvzDPIcD/gsP6CDmCdBOjveY9hi
7Qo16zeJqqndnEt3dtLbQUOwx+uWc68UeOhplTbV7NP9KEV8r1bzpDcIKR5c
J6X7PbACw39r3Wr4bExYpgIn5kvQgwpvt/pPGg2RmL/RXJ0/qvxf384QENYr
LwUxiY9mhuyo3zEqChPCqNMU7HuGmzwQ3aNfH96LTeKvSgFxqrSbagRfoAmA
jcvpb3I9/ZgomyMNX6zDeAT73TaHv6FbML8/3avflPs54MYBaRilcGBozU+4
yZqD7MRemrgHEVO5lt5qQ/xRpe9dpGuL7xiQMAIfOfsb1DaYvdbBltkUnNKG
2tsaisM1o4VUGY/tyqEUKnfwKgY/4A0qYuXpKMUxXSmSW9wYbwwJr/Bn1b6q
NZDWhkX4BeqbvHH7cftL16bf15Ev7tpE4RfGj2N0MNmbXXlIwNv3qjNSH5uf
ZYZGbRZJKsoU2nHJh3nCQDPowZM9Y69Hi6RPM6+EMQsjHh3M66iAFZY2NLqR
reQmpinhIYOSupAenIEh+JkgQqfR2iNU67iZT1AZ1rd67rYSBkL/rbRHKEOb
Qy8F+Hx/8LJ3LzH1ELzd8qJvPm6o51/VXNFZTmabf+kU5oZZt7lBXLh6UlaB
PT8zMaVSz6J04wDWDPpGCpKwOKFG+yvJ98KloaGATA7XodiL2SbzP1sSRsXx
IxKnxJBut0NvwqJU2DJ+TN3s/lK1JQyUaNTQmHKH7ZZT8+neBvMaE7hVtlo+
uFulYbG7uIG4G0kb1QRx8kwAX24jO5keFz6RemQlA4hd9JlYVt+UGlR+M9Bm
AXh8q3cS25SWuSVNMp2jtczczIPzTY9BUHefm8accLAiqSv52Blo+nrLEh6O
/SDwrYihJ6dQsae/ysiZWN03bNhtey9yeaZ+D1Goq/S+C3hgJ3Hd6i9g56X8
TJAih5+NCdGo/5Cl8cKiR2nyr9MKK0UV8Yz0UV06AeU2nn5zWGA/+Kc0o1NE
XTK4MXHiZNIqknranR+DnoPSa7AyEVko19PZ3IBrEmlZFE7VO7A3WH0Rrh7m
stmE/6m/70VP1v044o00sVzwUgTDNuOgAyDWOzXB/RP8G7uWIkpf00oxm0I5
DtUFjsDoXAcw/yugC4+iIbOmMGkj+5BuY4ofTAneibMk04twDchwQAPZXbXG
GNUQEqLD0KQ5CBRNWB3C++T8MpmyMRM7wy7CdzV3MInVxhBUqfiBu1cPAmER
pdH755FKTOuupC9bwJ6zrn0oKpo2XX3Jgmeo77LGj+uEsGBWc9cF61SrodS+
JltfvSulgEZ4/bVj1AtRNIbchhrQSx9a7Afz+hpiJe3q1kO/5PzcauthJ6Jg
YQ0qMpL7snmptv21z0wXi3IAq2K8bbRpVpowcOEf61fhdQ+asynLmvvT5g//
6/4Oi2WlKm30dFz/Shzs8YENDi7idMtSWb3IeFqyFfjrbw7iX0xGnhznsQKO
FJCYqeL4Zf9HXkLzz1thAH7V9AP/R/5vOmXAuIIzYy9BlS7XuLm63FbB7ejf
PlKHuklqQ7zUcu6Nljxs9lPSI1BsE1QQ+pCiC/bRiVOhW9S9GgkKPgAftr8v
mjFn/DGdIOrBDov8lDQnMjmqmS7hwxPaPDYz7Qe4uAoLo+vtX0D8NluMpSHy
5bo/bvS2tIlb2WBKcdKDO9dXTOP1hJcy8Aiydy1Cr+aJUf5QY7Tzc/B0/UUp
uBZq3UlUKyTMDhiKW0VW0jFMqgz9gZw8ebyBRVh+ipHtp/vGSpCF3kfS2A29
2RIuIZJVNI3d+ihXXtw9fqg1Uc8+ENOyVsSm8+SvFT2UmxTn/80Y86Mtp7do
3NpKiaNJ9rwy3/HBc5ZB8Rr2InNIYfXu9n/dDA+fp4PJLo6agCWytzrPTbhz
Cf92bogM8K0K1TM+skEnDDRg3pIK4LfSFb/EnI3+rbC0/b146KAaGj4hEwcE
Ucx79o3FFn8mafuuxR7d9j1A5kYah+ZPSxrdCuNFCDULJ4aaDv8YKLlpxXvU
N3QmLzcEfQ//SH5an8gYs57OO7GdDC7sroH7bwcfb8pKW7wu5DP2ff1pfEfv
9z685NywKaD5bnTD0crhfsIj/PuEJyymYEl7rycboMfARejSvFM3wcZxJhYE
CVozctS05BvhozHvHcUzKEa1YDgoT4RDEDTdsaG8leqJZ96nDL6rPRXDRO5S
EEl2GcbVDhHmmHGF3cY28jgAHBoPxfx5SBz20wqCNDUhJ6t4lTB1KYNh049M
yXMpmLuFL11UTvtWsdoGd86kJLv1/d1x9OFxH24zo3STkk7r5noJmlT76ccn
d8KrGtUkZX2kkBHssm3eYCuP19E098G11wLDkiMI3tXMkSOOIXzyh2QjEf8J
T0c3lW9JcyKZnaswFgx3bf1qbQFBntS2DlNYVImYpm2DFq/zJO0bAdHwI2IP
exXY/1mvISebQ7COKOw769Eh96Ny3qIAyc+lYTtQrBGMFsYcL9+qK4/cthKF
heQTKFl3XbYgcJ24dagUT8qe074hIJWqQzejTHeAeJzwu+8x3AZI0+YInfZ8
+1rFafgjuevy7mzLndYD+0TeuqL9zD9SqJZLvb7x1sYK/eCTMnd4vhQVZ+dr
y9BGzyJpWuKSAPIXJT9SjsivfA22bAFVQAyjR+cuRWODcgK73h3UZA6Otm+j
Kxbf3CLzJKFV57kKdme8UyyHWLlDPGy/KyScGZVzIi8+T47VqCLW+nK6S+RB
sJ+QlZ7OJxCrZMoV0E3vIow/NqbhxoHmutNZX0LhjqAT81RIlbW6fjkRc1iC
7GqDYXgLRSYM+cJXHSxuvdhaL+71+f8nsurzh3nRXV8XSG9/hEzDc0EjGUlH
7hTr3fwyS1OeOTfkNH5aID/h1Sg8ssIQXo+KSD8gPn9zSTNyTY/sY5vaO2jR
m+/ZDFgGpBgigxkP1Z2bwg3Q1XDw6rB8v5T443gqEnweCQzAFZTFf8oL33zV
1OVQtmoyY0AMfjzWk1Z/fqfpBVIjOwm2oOqid786hmLFFS2U9VpEdchwWMzr
1Us2b5yFjfaOMvVViFqTBEowaFBcEg9nKZ+x/i24cYAkOPinXIeVCaet2Pp7
4qpsG4NolXQjEyE75jdrIgn+uRfYvIyX8N5dlIda1RL2GA/3/rDp+47fVUZ1
B5SK2FTiJy83qzUZVTRykidy9fAlzLwyyTqD2U04dhKfJiZQO9FZkLDvpjDh
uFnsRr6gTiSNdc0BuF6fFV+3UFK1oeFSJx+30SaIdAqrev+wqA9gm/8zMuVo
czl71roqcAfupTxdLo3OibitFw6Nmyn61GQOIQBlqms13GlIvuvhYTEisb46
LxRZ3VqwmM2ix2qziWQuMjrCb4miYcz+sho95ueQMOEx07E9p6ryzLzxgLQu
ctjzhH1HVvtONifCcGU4YwOaMV1emjZO5FBTl2UVGV5RsTZ13NKC+LB2aI4r
MDBHwIXwr70mkSq9vjGR63J69VzY+bXVMseKq3cANwzlH/abkqRXUq16JJ3T
oKo4VcjqmiHVHMkRKXuZqSSvoOPUf/SMw2cmOlX2moZ+qgKrIu3IBHazUh9m
QG0lA2akgnhIkpsslEhwR6iRA4RrJuoXbifcpqFZq5IDYTwmTkDTflFhWEv2
VjKXjXvMEPaN2/uN9Vs27Kzsv3gQeHPcu8pRupncs+nilreI4rodffr9jsU7
pFPncxoZ6uoloDx4kRGatPJQdJNrQV27uKL1gvNlAGuHGTinPS5kXYlsaI3/
Qd0j+HNiCSB80r/BnffKwUTLA3lYXa4OJQ+yYvW41MX3qokZfCD476kZZ+PG
yPfbaYyk2Gf0wkrMZZ3aA7hq1uEapwZY9U6Tqy4nYDlev7CgUEPUntlby+6x
I4Jo8kLYbhlEMPS9TQEkYGoTToy7gFD2blRVglTi0AOqO9Ez2Q4ZpKnfWPlU
lKKFvGBRmkHnA9YE53y/pLdf9I1YuTm5x5dmzneFlJ5NlbYxsDw7a1I2uTDj
IwcQwgDRBMVO7UcDB1r4FfWn5HQDlIL6ge6qPW8INAahkMxwLUydVHgbFJGr
lbbNunCF0SgRT4wQrqrpkRC1O4/GqoemhVaehGzgno/FDZGP3/gSoymYYm68
o/An1lmKr5lJwhUWOWWX8Q9G6jHnyXAaCck+eOH4hKKNF0x/lL9aS/IQFjx9
vSCt1BMjY1YaJpilO8UW4bozabPDI7i1D+RnaJNKxGcSUoWo2rapDyZIjeXt
pBx7S1r5cP8h2DSZrIqomhMIL/c9YU3xcdDegq1ofi2MJjBKIaGlAkc0YxkY
xz1lTKYPBYqIn8VeHtN+aRqr+oXZIojHiwSuOIjt8jXng5euTvC/3Fxn8P0H
6aa5R76lnt6za45BtEraiF2DsLGuAII5JYAPXLLuGd1ZrBS16a/DHzG9kZeL
XzHehQGllAlDbGaFzs5nW6U2V8SSNustEA8PGrRxuxHex+AL2PvXtRsE678C
iHgdqTviz86jqZAEdpRIHZLafB5sG8FNBmuMnyor5un79THeIPjm81Tb4Q0i
0Zb0aQs6K4p7GzdCE8giYd7aCiFMUq2wZOU9FffecwZDna1ZJKyGBop5RZsN
Qn6jihL3heRxmJ5iiIbjWqR9oagShfFyRG1kpXvJNbq+igNUUYAmwHAbh0f0
d9FP2GiICBbqUBMT1ZESQsTaE1rzVlu0HeqFoWlOrxAHe6Kvr1ubH4iEtmZR
AU9PBWiBM2B9Qh0hWfY0fAd7hOsr/i9XI9WhDATk6xTOZ+51JOA63jJKOVDL
RBtemiJG7MyEvpJY7zJzAGuRtAbV07XDQWKiw9/1oo2xNeg2dLA1eRR4zVbK
PnHjjxMo7pNZj2C6hLPdjvyXnnNBiDItu1erUPoB+DB6GDB1JWcJJwtV7+lC
PWpX0WZqFLt4hI/Sqhy3ik7GkXEjwEaJiT+qFRJ7LEHjaM1bDWTWJiEr36Z6
O+aQZKklJn1VhgxsQuVnwe33kb6d9X+R+NRGfiZNtrV0vLYKTErLABd67ivv
AF5V7qCf4mzopPCoewVWYzIGq6az9ew8Bd3GSH+dLfHFC/G3rj/rMbRivDUZ
WTXtIPzLBUKUfUvm/h5dEszFV2yhC7TIizRbZb72HTGUj1irxkiET5dz4ZUl
OIEaXCfxgkIw2Rz/44H6ZuNONTj5DETkVWP9RekL2zz1QJpm+tYJIsFFADr5
izWw7lLCO+WDYf83VRl4mRGZa9FW2DS9Ph324PtUE+gVRURLwYRghigZGDst
ShD+DcD32rq2XI22ZGjloZlWiQ1FnJ/7VLTShXGXpMUoq81+wt9M+o2qwVty
9QwGbGBBvwmnBVfvhAGNWcyrxb8TzKjQQ7U1R41Pu5vtbaWsauZtlz+aFvHB
VaV5MlxwxEiFELWge8RkYklEpGU1vmSf/56Gpz7rKSjpuf4wLmUqOBPW0Mv4
CpIZ1NBn33dtzOs0QK0bDm84CRzpPAHg/YSaBfL7rwPIKHjkL/qE7kuu/mZc
iSNpHZ8blMBC6Ztjs1awMCUQB1IjKGLaQ3pn40K1lMYP8G8JeCzE0JmzV+Xk
hIaAMcgc6wJD0UwZHPgvMuOSIUOiwNSXlShf9h3INt5LnVx/fzgVDtdk8La4
9wdkf6e3CBRbK2bCoB9y8+DaYcCMW00V9IaUahf1Ywkek8GLosGTsJ1zQCQW
XvnnsrjhLedJWOjN6ospB5kv3/4I+ZV7bkxc+C0TvxumLDpSJMWCqBdm8DIQ
z5MNevP+SRIPchaPEXvr9qFL9Ct0oDlCRusBvb7orNIrMth0TgrE47PapHzB
FyCjOvO5oWMFtXBT2KlqdXmEGbxO3bJUKhN33lPpYGlP+H//wNrerCB+DEXf
6+lcMTut0sFsKwjVGcEI4wCCwa2Vp/r5TuXZVIZHaWsIBoxy0wBKTL4FWH3W
RESRfmRO4+D/J7+94odrEqgD8PALhiRcxejqX4Mtb9s5PJ2Iaw3v8nST5n4g
J9KCUYrLPo04MjKmniUMSUvh+2l02qD66zcqt1lL9dtY4+Pu60zUHn/1wsIe
XH+hAVPLXTBYuA7GvruPfgAQzNyP1qjVYTQNhUObHwOs0+JYnDVMzv4Wt5bh
u9yZXsTY3yCjbNeehTjZ6vMtHL1hfxb+Lg/NVzA7NT1/SGPGdlEFbtZD2/FN
iTQczpHsjFcCUxxD5rzu5JfuckmPI8v6BGoYyDG4sFExYb05Ld4yM5HraO9I
eyLEUme68+ImOtM4Q24vIotPWsm3utM3X54ct5oCjlYGk7vJHPpgw1aqksSQ
wEBNejxXkrrrBit+vnv2fIdmFSYaxFYNs8fSAYzLIeu9Fl6bJhiHcNU3rVOZ
o15+j1Z3gfMSt5yB4YaDBXV+Vmee

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeggB7g5X9N/aYeuO61bZVmh0qCncsbeY7qeL2ucN+vQ6YkKDTVsb7/JEKFT9TYojrxwox74eFjv1TUwgmzLicWu6yf91r50Ccs8PFQW4mf6P816m7PFSCyDg9j0mKD9dzyWXYRG8spFzjpsuNEGrLDCV6h5Yad6aSvkyV1+DGJtOnF7Tu8NGhvdU76crTt9er0sRX7c3LxCSfWKXnjoBaHrsuNczTcCPigAd2LYp1DPURbpO0zKe4/3PmLABUJkHS1BnruPvJgbaPx84aMzsFtAEaKXZGz6sjsOO9YFyFLdNQRqXbncxs2Zdk8z5fauhMpNZWmjh7OzozqK5Jc8sTxm1roV4op1vf0xhhUjCm7AnN7BsUq2IxNVuToUf/7WiEzmFz/F11S/mXi9Au5LWFEILtVOz4jtMKaYWjfdMXSUJXRJCjn/ANl7fLUCbDSzh5er4qiPu1cffdlAoXGfvgaRHpQ9/x3O6qRm4bFrgfwRZ/dpbzsW57K4CC7BpVI4YJCXhvmfcFhKJgevPezFsjDIxMwU9HgYjjtfyI4e16m78RuPqSelAZz0ikPhnv35Cyyp7LzsHcwwgnTxSq/5fF0ebMLYvjiDAj8hcz14vk1l9z67DCKEAu9zVQrIKS4/NJjSPTD43zwIXl5YHdhx7LWXdH3Hnhw5Lr9MwRM9l+FYtK7ldLOfigFVguiiNOAU3jK+Gc0hU9NYi5SUl18QJ57Gwp8LxBVscA0C50cKXVFCAZ+g4FprxNx8B0fxwaqsiCHcyYGgNhYpMJH7hWi2XrcM"
`endif