// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MH1e8cMQ96PyAONpartDqX43ShmWXEy1ifRYK5JbQeLrGljkM/CrEO5JiWll
BpKaYNfmEu3aMU4LZAtEGhS4JEaTXwMq5JNVwHqBopfolELtVPqP4Cltfs9f
e75HRJ5As3Y8KPLN5L+E9gwrEpoxDydUb4JUdAK4VBSaOWWTAwAu11eLeQ06
/OhEc0xEeWa18qvTOD0ux6aqrEDUadFvwChbFXL97huWuQRCRG/tLXhU1lMD
8d3xXiiWpjSwsjX5pTRKH8VPdzZfYfMzw05WqzQX6Kjc/CmQcoAJBT2owJZx
rKc+OaqxIdRB858JSNk7brx9zRZnZ0EE17WfXZX6QA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eqxIdhGqVJoovKU/j+6L+ZHDKbox+tUXGtA972YtK0YlrDheg8hym6QH5nBe
kMur93Avcg7nE2y7AHYt8CnMnCg4UBgobAAsxQ9QNUoIJCI0y2esfS7b7qA5
Ga/8I/VuLHuT30f0ouqjJDqLKAKvvbkgjk/un7rVse2o6n5MXqC0Xpw8g6FQ
Sw+R4W6rZvFCyUl+AQpSGX7szyR7Rlf6My0TvDSyaU2EXw9sXc0VE8yclqdr
eSnyIFwH6X+wl88YKWuq2HEVPJyL6V7Bq3EZqDAKjEwhI3lt06CAvCETT7Ql
RM5LYV8IewKYMNvw9s2L+Cm7pGLeRQ1Iw7j4ADDWbw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ueqIXUAr1YyU4L8ws00zoXmnSMgWT45jtxHYpaJc3dyxMg4x0PQj9VBQB2gD
3eFs/Cczd+4ino/fJQNFtEu8zwf/AvwSh666gu9/6Z4Ao6kyr9AUwqG3ZV7b
dVyaaR+YuEr/AJwXESLwWVeseFMnkbh0T7dBaAIdhVz+8Vgc+08EnrkIbiXR
E1C/Tf5NHwuxCAjRFXDp0jK8rkHFVf3ENko/pOdF/6yFwPuyW/JZfZPJ5bwK
REzevCZVAVPzQJoE/2w5FLPfeC1mDzM3b4+RHLWxcpMg+gSkc6Fr+2v9w8ma
7GzohTQHHYe9GpzUx9PVSN5SjoD6nHJbKlFKgbEP5A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XleYZjTHEbk7rBLKh148QFHTzH0zLl5CawTyXQ9WftDBjgH0RqnRyhWclo+n
tr0N3rZPYDpGorFXxko+iB/IQw1T1VUxi9E5JBm7e//r5oAjsRBD25Ja1pvm
cvTdzZEqBa1WPPTxGIM/RfrFfT1po3kpHIJkwp2p0xvHWvvbhzGKNYjc4TBM
kKMRSLhf+0a1iI1FJEx6mUcr+w2T4fU0g52DSlwn89hESa0vjDDV0tYUvwax
AAs044OBRc8Yst7oT4pG1MOysR1d9cA8lAvqslx9rZ/fnN38Xcz+3ahRHGSq
T0bQsA55IO+2fGZEJo5cj1CA/YAxmO3JXfnJdOomcw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dBSCyM+gZe/XKqmRfJVcIYMF2hoNUJATl75nPotSr/lejMwWTOjiGdH3vvdV
YZms41k1QuQU/mFKGp6pYgjLXCchic5NhXTJN5Yl3Izxyi7zg/Y1/npJQU9j
U/x4COER/DnhGFCj+TDUsJTMC9S06geFPY5hHHOibBJhj4fqoFw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ku66FlXVWxuiHU1gR0CkOHifo4aGzPtrQmPMcEa+9/e9uAr4f1hbp5eRVCoB
Hp2lHj9+PHa7hZFkNwT10EU+TRq1HE7PUwTt8SenDeWHqVIXa6XKVuP+g7p2
vtWlYpFIqMckNcYCdracK3ZuvYZBnssvfibTA48wSityo4SmNnYdvIyuR02B
2adCyxn53J7MTp/vfnFI5294LcyKZMW4nFPCj3MsTxY0a8bfqjN7cbcCljC6
RCU/+KF9l7iTPHvoNN7RxgC+cKl9RkS5AqdXOoPm1d22A68AEJAWGnU+7KPq
y6Ng3CgZd/NHPIJw2XlIZzdeR0CppzdbZsFyLDpoCKf/hcwXYs+JqtgQUHL3
offNeqtZm6WiXmsdqcqxKq35CoAbJphpYXnp+JmfA12X/Um3F66arY6+Df0e
cgY0DNass5m33V0a6hTStjkniL/LwtzFr9N2w4hQLy3mPUxlHrjiVVhTSPE1
E8HuZrXAhbf5b8bnhEfkIEpIrenXuAm6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Z1dxtGXkdJanqkN5WE7p64DX5Lq9EXfoSalvuBFS5nMhjIeeVhmhDzXkBVyR
GsyoEApoRD1VXnmiXHWNnAR3uee0wxCl2dr6fSm7TrnQJTeXBVtrW6JY1JID
CI46Y+7nzk1hhgxRqjMfDIzbZXU1lh2eKIvOUQawQgp/ix+JDHc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ril0BDXwkfKYDWKlSO2xELiZSdUSOGCJhaK0iGDImgV2JqzSdCTR0qFZzFXs
bbih+QU6gv4X6zFuaYyB7+el2deoPNWNEapbVCCUmQyKV0m5WWClLy5B152a
iAA6JSJw1uW/pm4sMZ1DQhIJ1wNzjKuAoZ3Zwoku9QlQtn4Mmzs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 926048)
`pragma protect data_block
nYCFL/QyqdF3mqm7wl3Ci3uxSyKJNKso75aqN5wii0stjZafkYFYYV0Iuc1a
AtibtQ89Id0B0FQVlA2KujPsugbbYkcTpUEAPf9ZzgUiZw59gQ74YP+D/avA
TluFzvqCLAUxb/C5ajGcHKu8cs2MEyoF5/ALv+gGrysdQbZ7LANYovOpRD3A
JJ5cnj4glqy1Kz/ntMvTcI3Kx4ny3I4wEnLSOCAFPD6zjt4uNxIHcB6RVnRd
DP9cP8CMGyVsHX3ALKnkw0QnQk+BFwr4RomhXcXna/rxU1njN3dKktBEf1Wb
5fuKBmP9YlvEN4Zdoeyvh8mYw1/bgF2I0FLggdElGtR2BYcqDB+TMDULFGaV
8cLPTLQJ0RrKumut8d/s6CbCkLu22m5DVHJk4rsDWpJi3/3EJp2Ew3XpCsdS
b8e2xFq0U/krm0OcCMhk6aKFpp37h68Lyu1h4QESaUcFv3XBWooMWdWIsPE5
Fp62dJCnXcRtpK5ashpXUDBDKCyTALLLijIUlR/pksbpNXfLd6KjJHrvMO/c
wveZUB3GWwov2F+zrBbzWrvUvF1ZGbKW+Ke64rYGb0u5RW2xH804D96KRRmR
F/v8Q0RWi80TMxfcWAyFd9rGsL1k27gquW2rimPIbqw+zBGwqhvuijFfgKkl
TdUGf1kTAFr/TL8ou8qPmVXTnPZ8eNQ3+KAHZaoRpVFgRgHpEM+GyyB2zwgG
xkQuoVVCwGYkR+8MlvWbtkDGAwN/Ah/bw7K1iqySiYojbLQI4nE+7gp3fLld
QZRMrMPGCeakedINIlH/Dg+yn1HqTJSvOOMAlkcWka8IRvIE8fOdjs7n86JI
I4/EOc+PFPg2WXqOm6EwI6Cusox8XBHh4PJ+6lWGPZDw4xhwEMDRHb684wSz
h+fdj0xmYw1ezEyU1I1jR3r4ZqPdASBD75rVXUqqn+pIX3+fhxKpGwgVXvOy
xPZcEGvk1Zej6x8SH5h/mSDmH0FaKir7Gcm71W+Bsgx+gU+oYNFdT/8ZbfKa
4vKYAYDF2l7jJEwg8VHuHqo0+uySNleDPzuXzgpnjw5K5dqUSRfxDNLfy7F0
0YFc08iw7ROrk1T+Ha5lCQlDzO5QaWBScG1S/2OOoY09DsY7Ybz2+DHf3Whs
6UxvfLqJCOo/Isz0QNdOmw6ztU+xukQISWlyXIVOE5CaRuCU+p0Ix+MMGKII
MglJDZF/Ry5brMQ5V/+yXlQvZp7hZ4XYfB2WSHOWN+sgsLz1g6pVcbMEMUoz
/7/GKQX+u5fs7VWf6dmmjf9OZovOWGAnwiGYU3/GTi5P+xFOVJWyhNRlgP49
4rD1MlYzf+tzaT18P3YYsbsqqaDkqiM8zJqMAZGUav4+5PcpnOVo7VtaYH3A
nyxikgvQ/T3vC8uBdNqnoc/fzCimeFZs08oUewzAZekr2xYKFFVujK+8m6D5
EwVNsa/XKlS/4S7tYClalgTJMfFgLAEVJHRSP0FsjBcI3QFMVOo16LGN/Q+Y
fiii8w6bw4eMiteRHPnX64pPCeM3qmsToC45gp1sHGIH6Hl98RmKkmfu3enX
XYXSqkhdFRwFsphtn/aInS0QiN3FLAgIC7lAMFCrRkjfzMlaiVqoSShutc3g
G9eEzJeWREbDVypJPKOasmiXoPpDLFV6VWveQ/29n2iWQjvPqJbVSL7Zb78l
gza5ECyTXM1C4uZPpd77onbA1cz4fvANKP0e3yLSLhsJZQL3xFMGXCYM5e34
ZhUOF/9bCCsT8ADVE6a/yNdKYD57xn1g7iQ4eJ0Dq8yBbMBqCVHVOcRZ2CdA
ucv+K9beWTRsoDJOToqRLeEiCgitCqTxKoQEr9g4twm1o3R7lK4liN7yFgQh
0wi0DyhscNJSIVlPwUXhz3ij4gpEotkumo81a+iizIU5VQ7PW78f9wsosCGi
pylJqPPkU/dFPNgf0VKMTfUajwnNbPHecWa+qHn7DcolY8PAliR93Dw8eMRJ
9wBnfb67zFkYi9bTUimmuzQJxEkNmKyuyM8L4Sw/IkkGnnUS2hslUu8xMQTT
4MidP1isv0RjgyjGYZNhf7MMqzzzXhMLuB0AhkiTiy59QlU4evVdh51vkgfy
uDV+lrBbBQ1+p5xP6KaWPblw8U9tGdSvabP9TQoJ8ux4ANP/rhhTcyUowwVJ
WXrpSi4iTRQsguowVK1PEEsyG3wWRKiPcff7OlBVdQFg7r9XrFMw0oVGozUX
eKuugHAJZeSI//37fCuArtBRJq/Ze8oy0gNBRxmJ/cbtLF+VvhzOwTsD9nWx
0CperzOGrSQ3rOdHxq3H35K+P05YGQcETz/DX1Opf85tKffe9wgjT+cgI9hr
N+5N3Z5Xh0kVzUdUqMSFCIP9A0VxIeNy0fZz4lGxYK2VNAztVM0VDScq1w9u
0dPyqRaCwoAVUtMEE+JrOFsn4DdPjYW+WD9M19cqCmkjVNo/H3gr0ngMnEej
kHWdYTgf3C6cyqQXMdBO72HiZHD/vpHYmRp/BVYRv2FSVkOjmfC/jezI4DXp
EIQot/ATubiYNk+40ezXl0ez1n89pF4TYHGFJY0R8d3uN9jsLn0TdUspYMQ+
hJb9XCtLN2rh6jwlvRUcdmOVD+w7MQOPognNWCODsnOzn98zEva1Re4ABVP7
WEBao1eMtup6Tgif3BRCDnIkq4GFBDxDt+yAda5Mn/rQPn6ymVMTx2z25Vlr
pXl3EPgK20yiuDv7Itoh8SLIhDdpuI/SvUi38LLOnroSLAPKQlshqkUVJRzM
4Qtbxx1FuOgI/3rjyFXceNTo4wZLsEDxKFjo9YHdlW4MZZwt9+x3oCCaRpmc
arHWYIF5GO69BMKqeBT9XeglFheGbvtavi0Uecx6wbbqPrc0ldd/WTbiU5jm
E0vIej5qbazI3iS/n9ETJ8yn1E9XVbnynpiDKRawsSf6E0/cZris63qGNNRW
YgR3nqm361UZo1LZJ+580fHjtrxIs/1nomMx5N+jLfQ/MTFoM04yH/fv24FT
lje9d0dUHh+5umWYw+4BMGRrKGo+TxFOn6iX2lt+1U2ttg46lCAPqzsIKjVO
VizFT7m0nce6NZRtLlwJnCk3wuiplfbT/JBeCP0xaGe0m8XjNnKZHNKQqoWK
abkN5WQwIv6Y6hdknzNlLcrLITIoEIDYOKhaFF42Wsq5qKqY5TXKmBwboxxA
M7SP3E5kfBuoUZXJcWwWLEFCZrGNnjJ94gcEabKY9sR2NKl03P+7uUz7fPJX
oyRy9TO5wDJ7X2tkCk4ebluAnxpx55B4RaPoEwcNR7ulyxf957ptV6eTDOcQ
q/+69o44U4Akq3oW6tiRDWXzbKY5Qm9KICXkCwWKuJcGIfNIuXht6jUIx6wv
VyxCU3uIn2+LbI1MDPNBN9dGEhTCvPN0RzYGSjM46H4MAE+MYiqnJOj/R93Y
SWUM/17EM+8VLOdPDP3Cf+hKBnBRTiHNDhgnt/cyW7N4tOO+lT4cJ4pqhA3g
ThzJ9faplgcQZNjSXkCfOEysNFe0LpTTZRyIuITD3L7+QluuG+DSjsxE2mW1
Ouh/4uKI1KRmwofeJmHG0luYiCwv4mRzCB/eMxkBzHVhvJ0LEsrNHr4QG12D
JD6/nfhSsj4HjXzJjYJEYLh96QCLBbpAZjByJ9g3OOTqckt3zbV9VL8LV3vU
ENcrDoKB04dDj1FpsMDOKotUQjDrx8NKbvzKKSYoiJHIhOfr7/G6cE+uryPC
S+b5tvJy3GQVjDfQundxOOxbkjfUuvQCtmiCr3JjjzYN5+TXsG2zS0mP5y+x
HpvpszXUr+/efxKIbdWSX92POdGYpEW3ydycRN0mg9wkZvClZ6jLuPfzeoj7
AQBmn5iyS0wozTkt1ZZDIGRzTEL7XinT83u/ARjArPi0Paj9UqIUMRzF3nmD
gXDfCv1E1FLsuGO/79vXkOhqcgAPLhEdwP1g/yl0UN0An4wat1MApQYPP2nW
Otk9UeXuBlkfg7qrk0Yez7a+SFGL3OHXrcw0dtdSw6viF1iKgfHQJMQKmGWt
qQXaFKZgUZ0DQNwNBeKgxLD1ESxy/B9R37Nf5fad0emeotkhvypokyrpKiDX
GJkv0HDs+yJ/OWIU5u5Q/ThHWfyNMKUr4U/RyCI6ohoT422q+Cu5SIl0htw8
PYaTBF/34Rq4es+jeYbCRF+chKlVBNH7udZTjYPxXG3uus1ec2+Y/n00DB6p
alv5iKWhtqGKnCLFt79ikDo7Lc8CW/PxqrPbDM7VJ2FwJnUWtV1BvOvYwOur
jHBj7r0spg4D6IamQ88GoyM6TYtpfDSlh3EOGBFvHQqJJ11oab2DvYLzN+Em
RDrHfAZ5QiU890fblqY585OZ4Yw3XMTIC9aNE1Q1VhSBw+Wrs4jtFjucj4dn
o6hTc94RYCEYxYyYjCJcIKVh4AJcdqQDLRAwjxuSfTn/l51VcR1cJJT1run4
/Bqz8EyWOKFB6lP470YN74N2a4se0Ktn+MkgE9wFUxe6GRpS+xj9fxODbkox
MqFwOcthMD53/8Kwq9y+89pU+8lCIMl5/XdI5EMtOvl6ASsA0csrgSzoeE2J
ikXiMIaGc88TcaNYQiTt8Nf3LOwx240uGsowt4RCJUyC/4WKU98+3RF9I1kj
iGYHvlqEQ4CHA+9bzsoGJYpoY6nQ5MBt5rmdM6ZS8eyWsYG1w0BKAAYk+wCx
N3DJj/UEnvwZomvM9xjn7f3MNY6U4NORaFQXVcHpiqzYr4RXmFMPYD5TyY31
mODEGufp9RDH3aJxi7qmK49jpnAj+p1Zd7ukIxTuWRxxKz55psnA9ZoQiszl
5xD9Jn+NMG64Ku9rdXiLJlcUsjScCn5WptPM6Gs+zhkQ8w1oCgVEgO//2FEE
mKjQfT1QGvoSLsM3o5cxMa/ee9inq2dP94N2RJ7CIazV2Npr9T8grRw5Q5jh
yJ1iGv3MIh00VgSwyzgR6Y3erkPaxtGAvXeOw7+Jphkso88e5s9NJlh6Lbe9
R1aWflMuMz3fTjDmmezpyb2Qr7YAC1mdvP8mRQjnMA89gzIE12isbP2kiWZw
EmS0LYUsC8kO51PaV8hfocBxmnUC4ewMKZ0GQPk9MklIR7Or42xVWc/iP5mb
jA6yWOLr+91BOukQkMuWVbpCTE/DUZpv9e9bP8TT+exDZTBFBAoPvxJ6FTS6
pI4WINLBvVwi/KKza3i23cutv7o+OlUqUIo+dHtYM0/2hGHn0mywGYBBT0vn
SFJbmPpSPlh4ERo/UHN36qGH/aTuuNFWmKpw/VzS7inylLF+37rsqGDa3lwE
7iKuYekBU9ee+saE0dLTA8PUNUXczbIYCqY3QTQqcuRdm3ZVPLv1AkXlTEr7
iE2zKy/T/Zqa7lvuMXd6CfeQlxaxnk/hNKClA8C8fnWamm5eQW9ZPmmJtz4i
2FgHK7w+V2sND3hRYvHpvv93Xm9aKexWwNOoGLat5hEAClgobZTkMyKMxzt4
NTgWrnYt84jSNQHaUZzZvzNV2ajX4jz5IrQCjMsu9S6Uahty4MfYMODKl77+
guEJ1hKHZ6C95Y6uMz1xdShj8rmcfHQUbQcxC3Q3akFGz+SbP/aT6Isx5ZB5
JjiEL9fIAdb2MjUJb+pk56/Y84T2l7p+K/SmcU0uhbb9FpMhpNPzqlhJtAxh
Qt0sf95ULxAF0qxHZbfEPuTwPE0VwXCd9thKRCnMY2ajeldTeSqrU4HiWOvO
pX2l6CTAaQHiDFdOHl3fyiFpZFbQ0o/TkvEUFHgFYWVL1dAGGi5DhaPH0qKS
WtWvU5AzjKiVoegFqzmTnRXMbj7GrcJ/qhKA9zRIFNDZM5sfD3uPhXVa2OYh
0vCJmEzYkCjkox/IBz8yI28sh470In9o6GjJjeGnt7E6pdRZbbwI98pT7Sjf
r9kQCQNmr9X0erCd+Fphwbp2UXcH0Jnd7SeUNdQNxBXwvPpOYmeHxYhH12l9
Hg9bOoQqbFOe9F3OytGhW/CkRmPHraeP48Vyt80211xaNqyNoqluEzORxwIg
uVVGRfGB7tK0E1gSkYyLtYEl1aWwSkoH+8OrP1WmW7VzNUWrhmnCXGw6sptx
WUpPohvLLS8fHzuSxttJydi1BJ66qLlacaoGUzRBeWTRTkB2woEEBZfj9+qP
cv8pf1niKkp54yQNkDGBv4ufldKBI5adMNNTfkkN4nmzJZhR4FPUzQaFOPv6
fQKx+4V7VUqhXGhz7ZdEzN/3+iX/wVBDqfCvk7Sjx/ynWroESRctTSYBi4ja
UMlFiZFySUDe3H/8vFsr5H2lpylcwvSB7wYjIwRFJWFwC4jGT931J6bN8FZX
RNLsTanJWcVa86pTNLu2E+wDyIj7d5KX4ivmp2zIj2RsSuJz2lpQQnWKoC1a
faAT5foXjDktrGpBmnBPSkOGWs+rn0PZkiCCclquYTR1xs6f+Cro/zLgkCrx
X+IwC9mGDzENcNOVEpTpbDHUOUYc+I58mDEDx81+AApCTFupPlAVo56msqqk
/ckqkENZhdf7MwXDtib8Sx3hhUnDUUabuSp6rfEG1bpQrlf/+ZBPQea6DlhZ
6rw9KNvnZeh3bO1sNfzTnJPuW2usMGy/QBchj+FxuMEbGyVtReG493A+Qduf
shZWRj7BYJYZLoiKHt5Ulccd1pvILcfSBVtw41rUMd2yQRaMSGz4cgahJari
BXXPvyoIHw5PnnMEe0cnzfHiMloBEqAEVFm9Dvf3tbYRn3ELc0bg7grLAcCx
MpGUZvM0OYkgIuuQAabWEQyNisJU+S5ZVOksR8qk2K7yhH74yjTnbxlAET3c
43XcgsY6A/xDrTHFDalAakic75WapxPVCjVSx6esBIkX+yh6GExuUJbp7aHz
0aeiQELxhszk6bwd0Q1fcA71STiDMuK/i3LJsMmnyIICyl9RnoPQ1ZhALTR2
Sov8UsIuavCpHljZThfW4rBuYUEdTuOxUzi/Gc8nUtdtGmWvaeOBMcsCQOC2
X0TOTeZckLCShbSyD19rkDEwVdTru8azE+m8KPVa1b5ZNDbAVjsAKxBVKrcA
cej7RFpUht0axqIXMleFNmf2Mh1FM/TliAsm+HIgZ+RzjrwogNCC4lsN8TGj
Cu0N5YzS/Xp/E+Wy3SxXW2T97xvLKqnOnJsp9MiG9nR/FEdsmjrWvC7mViTr
Tq5R/YNsIzMo63wM2m794Mcmdk2HuJzpqLbtLso0m73nCCcEl1wWCvTcURmo
iwiK/fqGD4jsaDJgkD7xbBbj1jeXlTSzfEmFcYWgR4vudUWrixjJzOdIhkKw
e4/k0PB1RQzHfBxG0RJGTm12L9wf0dG2JOEnAbPR3CDb9MyKDc7xcI6dJD5a
qC3jACmkL5F9cjjqzrt1gXyfvnViA/33OEwLHk5jq2HsPz9msBm2jKAPQvBL
2ihot0j7ibDj9DOYBQmkBrJaOreMsg2Y52mQ5WPZB/GUYBWyHSqcBfDx8hzO
7RPwGqKkvktnHWli6nEKIWRPET+cWe4al/O9QDOgHXu7J/jMjjofVZM2JRSj
10eYrNfZBZPjzgay8GazQT/ulcymt/xJ7LbwizrLjBnlR/jNw7yl0syEYchJ
S0QY9ksKsDB0YvceoiTmvvoEhie8M341Jh/1fS5ezyr3XngB03IiCf6UF7hI
QpgRoB+NAjLvgdepL/wrZl5hQJmWhK+0WFHb4NP0jfVdBhl6+A/sMZxqbJiO
eG+HDBSjo2noL5wu+CEiXbrY2Jf0wT0JJlGMIC2GpiXCWkotHIA7W7BPiT59
a1EFkyBygWnCOrMhJChJogYmJfs+gLTZXPdvYPsxOEta3X7ZES1cvaGe1y2o
04nXlnuXggoB8Xhx12Idx6W5PS0Zdd/wu0W1OUW2UGpPWRkdbYz1Old//Xun
EwuVDYO9GSKS9UAZbwPTM5yT11hYEppfW7VK7Pp7XRRfab9prRG97GG3H2Ma
sy/X7muV8LE6jbmJRJ9bYnHemzN/7HH+X5s/m5iPCbbJSIIv7UQz0xeoglnG
43v4LDHoY0vBXEG3SrC7AOhAy9vKAJ4M0oTno1WFVDOQKq87WF3jUGlX1UCO
PmJnVEzOFQeJywntiTuElNRevabwchfxsah1dAh37Dol3JRaGQPiqSz+0mcJ
wNGwJszYa52G41oPQVAi3q1GJvZjXi3vra2YEb5hRZZ2BbXWSLFdwyIHvjfR
8c5IfD2rF7TZQALBI2sKNav6NjMaEZzrISeM1VROOvvTYpyVbdrXgjvjjrTt
+vPuuuhoLeWPVzhHven05XjsgoL0NSLRQYkzy6BOcTmGZdGDAM5uMcabWhQE
CZ8PDulLqDIkNQ7NZsqOj574BLG5rZa/K75Dd+e8W4s+4ADM/yK1pqGoNcLf
K1vaUKoGiESx/c6cOAFaKoF4+sSJLSwlr+lnXVG+DWjQ9Bcj6rh04d8x44rS
fUMiEXX0zXN/O4JzEpA6SQiXoz52opKzfagtazqbqJ861wKmLWdlZ5sPaMIt
ciUdjagEKoi5Ho/EnkQOsxXk6POUF0uffgAyKvFGkoDbzOCnrrsBrIy/7UkO
4eVGidNSiK6QauDSL2qXA8v2MX5J6ncFPt4xh/wTWEA6YxqYIm0qry+KMVBC
Y04eZ5+beRCsuGulUscSBVT58J8PZIzHorRzwPOHo5O7kgrVgt8dSQw6D4CJ
ohmTmgMqe51W58SPnhGi6yGnVfcPhSqsCnVCRpPaMjH5Q/hVZb6fjIfjX4vx
+mebaV20QR76QrOLrY6uQuc3BLpSgnmspnC+wucVnXFb2jJAnT16JQCSWPjo
DTSmnXRKCJkOgBlbTnD6SaDp6UTVdbcVTXIp01Ed25ky7VQ3t4ajFM4SbbTF
7vQTzwWeuOhY1FHGEIxRfbkDw4/OgITa0MBrMq+GxSR4KQwXW7Id2Yg6cuyw
8rw1oSvvVe3FTWYSthPuLmlnr1QQDkZwThZPvEPrNTnzPDKSTAcg9YAfvfoS
IcKcoRd5JxWNUwyIvddf47HjZ0iYC5G+/BwYe/IIpE76ok7hJgvyYV9Dtgbg
tIJgIbBbujVgK344TI3sXxDGbFR44J0mEdOeT3e6r5yHxGzrh/gfh3BCPlzG
4j66oq/8hIEkXRjiZjR3xj/T0QKi2nqxRW3/ZoogPFkcZ2QvJwPLROmWkrcc
owWdnIBJYhUUZHyXSfS0nuM3l8uC/qLNaMPbpPzq2lJMqd7jaxKvhqd5G4iY
ZysG5JARjkOQ5jmUgG4kHg9D3O6cszQbU/TepVTmLqi/2T3irrZnaj3qpync
DjxOIr3s0Otmkk+w/qbbqHlMRjAmPIqAv31j1LrqfkqTc6vfh7EA0LT3VuIS
vMr/p/QnfWmPvmzxWTCdOO/f0JXfLB2Ohn+jzsTvsZFe+OOwz6nZJ4d6JAtb
gCVQ9E2dQZg2FF85kgyEtkHuH5PcBfqSnk4vNdMSShGNWGgclmGcR3MMHyqj
zwVC4RMsUicyw8N3m9o4rB5U2LW49zThdby91uI1mH8x/wceRTxix/qbw/wb
Lq8BkDR7lKFJzHofNin6cwFw2S/rDiBAJHA/K4G3k6Tu7+inbpGThS8cRJ+2
VFK5LOcC+Q8RHnq0QyvJCxhMGf25gPSHO+t+cXBANhaSJrG50bTb2taRCzjG
Xvpqh1kVdlrp2WmiNbMC8R0PzKWLV9Vltpr+ldsBZAIfjnf1pzW3inhbb0Ba
jfp8gdBprzOgv74NRi6DvMWiHx8UTw9HbbWXaNHOI/pzKCQsRZjQWZ0Ivg38
KjJTOKpTTqUDJ2TsYA60uRlsiJDgl0OTqOjl4HScRFabKYtDwgH+zlCrWiHC
gbvISqtPchVmx+apzBnb3cm0B/vlDJm58XvvKjNeaS9SZe07fAgsQONJs12D
J89/XmejZQM1Lc/TvBLs1GL7gSRutdhQcXmOluVk2lSbsY2IttkRJsPqpwjs
c5Bq14XPbnIw+ng/Yjmq7Qcz1nkDY5cphmPiLUVKqoo+GsEY/WHuIBaBvb5m
MYVYKy7wXxFxeYnygSeVf24B+h5odE8fpcrRDZiKS+kHvLjRmHMZ6vrGw7dh
i3efnE0OlyTEQFDSM8OaH+IBPLLiRO1elNIMrXazDU6MrcaRkPwXORshWTKC
5cdv1hg/I7vY5/e8uBoYueWqW14HYHAqkE0InK7HNiFW3VtkIKCCVmrZluQz
Gg5nvNnSc8miXMiSiwoMPXsKL9SVPRuacpqZopmQQ9AqvN/5FsM8kXMPMj1Z
XzOBK5e+3h9TERk1FVRjL0BGBj1bRX7F2gyawTgFOlV/CMYc7HPuDrGZ3SLO
ETMi1y7f851Gd/r+Ku6i4vgSG2xqZx6h0y/xOvNbnaCDlDEwA4Yue/Z4Hb6X
6rON/OTLEsDHsKcHpt4XSIFqn+3VRTsMY/lcHdZc984mauXZaG7e7aXeDG7k
w14lKilOVgH4ImoSgDcgAcBPHJLSOmPsgUoT2ySG7Fldjy4keZpKZFRHhjgx
9NqjdJPz5OWBHmBWtc3i7SzfZdRDPRMksYPKBMKUzWayQ/edHNrH0mjx5LlZ
h3mNToTnqRWDxN+X26PxP90nYxeEZLtbPLdFZ99xAvbZ88a2KLwVfRex9ZpM
DsXusJzr8uq9MB41XJtvPw8R06kwVu/PW5u6V5S+NSm7xsivanqcJwHnk6CG
uylUmGieiamohwjjpLBZ5fdkK/iaug5JeAE1E2glOI1w7nAWDnsloyoHTWTD
NCVe1NW0R6Qi8zpz79RusbgLf91aivcwSzpfIDfrxoJInE/DcbwZEWSvGGP2
SI17RMkLaH0VXep07+oW/QyWHNeeCyuZIrwtMzQVCX7GxeJ53uf60/dtjocb
rK4E6R+TLiGHg03wOBWFhmOjOIWBU9jAcFvAAVMXG3siFs09bWoUD1TtineW
1dIExG3Txg7NDcP0M7QypIQHNhYP3TyPHk9Dl4GzgfLW0k+eAwqyd5erxPFb
uXR13Zthx7sPpR3M3k7XLEmBtRJFqhV+dx/tfug6bBvcNCLZLlNFhK069vgm
/ca3Ny3Lba/bi97yympFdDPSTX+ki/yT6vCXVMnhwYSLOhtYoIf5iZT+2bBj
ClddTsmOCG4rk7n/a7evGmZ+85B/YRSU7TF1LAYsl7yas53o2clZLEqm2mdz
gSKPBd639T8PwFPY/RSOfObvEEqFigmpJuYMBhdjkEXAnNPfZH1/AwXwojn9
NylAVZBigDzz8KFtIIS/xxlwoZvqfq76XZ65WN1M76OtZFiH+5NmWC4bOAiu
RWa1+jyDQit9yDduCiQiaO4LkvUFCcN9UufHKlcnZ72x6ix2Wa+eRLuJLB4H
TOIc1XeWr2shLapk0hfBbwxB0rjmAcIdhcP39Mvf5BdsPrEKjobgY3N+0cTj
QLU0ZGbpyxnaJ7UtCDjwedD4UCX8ilNEGOZfqYhFMmqLQ4muE6ib2CqcuLTe
wHRHhkWaVla9QAF/kd+R2yxZ8PQOgm0+cENKWMnv3IoU/qMDnwZc32yS+bc7
0gFtJyp7FLc1uaBlwj9xn0bbG2DEoYGyAMuq/HYhb154yVJVu6icNqRpYIsU
zF0UCuYsHWkeESuXOjt3qS2q4XbhEbAoDnZJ/UKsbI9iZ4iwxC9wFCKhytcv
c1S3F1nyEmnL+oPFXRXN6c6c165TSqhce/BPCl18xr8bjQkxVa9CDUMIF5SP
gc5PLj1sA2pSB+HNnI2ormybuABiaRlk5PO28b3Y2Olf4mA76EcuvlAEtxQV
EgjgGdfUngP6E2ZXyM/q1BWHo07AMErsh/YXcHfkYx+Pugi2bhSovLmNNH+D
1v7j6YR1vDEAEoRCKBOVqGDEoEj+seXBYjgvukigjpPS2pIyZ6AxQVKfLEIf
ZFPi5adb7cpnN1oOlZ8ZJTAiXGGBKYeVN1IFGXkFpoQp/Cn1IrbJAP2T9qfs
r2gFGjhlQwTNglEjGSFu2vQRaMA27QizuptMTqJAIjr3juVwd8yXGQ9osEL1
0v4/qUPF5PZgr5fuhmU34k6FqtWHCslcOMuJ7aG44JTPTxYmmyZI0ZkXvRSE
gGhyFdtOhVAojaS32y31NRjT67DR9BprFIr0e0c2vdaTSbEqN2HfQXKbwPvL
q63YE1eqitJ/AOxWEu78okAf4zeRhsLCFclkj/7WXIpnqaqJI2d4ZqXfRFCi
qz59pGtoqdLsapYM1X0T7A1elGYDtv432+TH0FDVi/7ktcsDyyIxEB/1q7/z
0tzlNRxNFl4Os6U/6LF7Sj8rBFOSfm1XFNNvpJJnndGUljJ+BPQsG6v36vw2
Ppa2CZ9nPBbjwZ3wI+bmbYo+yyiuxLEZBf3wRpqLRs3Q3Z1CaNeV/AK7mRNo
vg8XCBeBw+gxVn1esA/WhvOeIb6vrQQN9uz7c6NIJ8c0hf6C6yIZoA190j7G
u8/GG2R/fRxN69/uX9zaGTsk+LprIQO2OmGR6oXI8/soewSQPfEvkBEziKBb
IedqFZpcQ2XOQd8wIBgSOJOjp+e0k6Uw3Ya3G5PdUj1PNaFmFgZhqd9Ni8HK
NBQnrxhh/t4HfuwjPhqDsGHwLGNlS+WzetsGwfbJjpFqy4y+flkndfdyDMf4
ZVgee9xzsY1VXs3N1yBDiZ+mfx5TluzT2Br99b6xDpi7JT6EMXUiDVuY61C2
F9lLGPOx0Hn5iARE0FOWpeLbvHaTNWRL8OnvrwEVXpv1AYWzVqz+e8hpYvjy
aPm2Ri2oqk100cVho2tOvL6OsSrJIA+T7X+l2g9gItPVRoCGY/I37PA/lAvB
34DHqoP5BvEZkKARCaIvPdXadWMZScNVkAC4R9hGNmd3XzTczet3SYLgNXJV
aVdjH2kynWiR5AFRNDrA6BxZGbBKF+XdX2qLGWxGbshMTtXL5KMJ+5keWFvB
pdwuEtevEGGDGvNXdMO9Zczt1l977o8BrSBdhAFR59mwx1PEYryrqfRasCDw
k9QJoTAG1VD1vpAbGy8h/Oq0MHovlsiVdmbLc9cs/tnHY+1PJ9VQJMp06AAr
HjxqjcydLcBlGnLrIK92I64UlwL1Z7K4AgRNAHWL+dBVIYsmIEmdeq/NRCFG
Xf8//4BIFKKPTl5VVgVfGLvJqt16A6eMZzv2L1WLOCFoh+67o5KDuYNRdeRa
mc6TEnFE95h1LvYoUKZiEfvCtN3c5RVM1WcSStA5qzUm++5nxk7j/tdWP7oO
7IynpAhTF9dJDeclsU+0aWiupFOe9J3pyze2H7blDg9mJbMUejcgEY3hEUs+
CKe6W7fkHKnLhDIdeUItXQCeXcO062SYgJv01EqfIOBAEBM4MFKg38FsnGva
sJMu74OksCtNkE0QeTSaCEldxnU4ufvYhhvtcUUj9N4KLhTsiHyoWQNKHhZB
3URQgkdNVPfDhquOkEAmH62fuuxR5ogYkhG40pk7Q7rvYLKW0/Eyukjkmkms
Jy3eWStwyyhxMTpU9at3/mJc3DoSBFoUkCGlctRxHDqw09ys3JTgWY0yWJYw
+AhdyTTbrHlEU1ZcAda70nNX+tWHBKGdCUafyZBwvO453avIRyPYSF45kMKD
HpXscjaVbr7PGhgvkjOAU7A8kxdU8uWqR4EAgF5/eEro4HC2SoRHxXg1RLi7
MIgpf3Byf9NqST56HLsefNJgAQnfVdm8Q17NpI1hh+az14t/W7/+Xsn9HUg/
qah4CmTsdTTqTtMGwTTZOGYBeY+IhQrYzgCxAvR9k2GzBe6JUCkwECfCFOmu
Vb2O9a3sMgj9tR1uhY7CUDzBrWiWvI3mfOmkHf74lPHc5nmkDujm3eWXkbbV
F8f+0Rsl5XGjaYrfDTiiRzvQwKSf20S9nEBrM1eowHRGwQYpSTj59jPuwFn0
FLGpeaCZ3LNtmOq0WU0QQlkQogCFuOsOkrxf3GoPxXJ0cPWeR7nF53xX1I8T
RbB3l1409amVYGK7hB3Gffd+5qlaF5hu0sAJ0bR5yITssJWsUkW71zRnO3e0
k3mAE7OBVoFNxy1P4SVDUotIFdUxr20AwZuf5SzdtDvHibeOd+U1bUcFZ2Y5
BRBe5At2xgdGLxWrQ29/mZheL+CPCy0YNuPikU+tux7Z4bDLt9hiijelqHBH
uqIOEG8wQAji3MOBp61AmHGLdMY3TfSGF7ZzrDCfdvtsAp25JPSaUWO1aQGe
K4hEAnLrNFSnIIsAPVkjvhsqRaExOR2vu1hGTozi8PQQMzSqQPNaNmMErb1m
Ea5Z9NTKauKby2ivbX89pACEgTQuaolq3RmLD9/x+k9m6uKfdbXMhCL5m4AE
hoybKSdWf0MpvlSbcPhS0sWUS6ZjNeuYMV5X46HejiCJqySDcgQh9AW+k6wc
fj6SsfsMMLsAFDUuYfOh4NJZGX7qvSXWN17eRvHuCzoDuWTjCbU5La+qTTfh
85nsZtZFG/9wf8zTYfcMxufk4h8HNS+FEDG8Qa/aKaIeyFza1yx8Z4m2kBb9
5btU9KVSw1VSznL815temijDYKV4CDxop61AY2EOksTBIpb2QODDiK9G82PG
otb/XdRxyybQv9SeLFYcsBvV64t6aNqHEjHr9/QNUdvKzxRKCRc0S/UnkY/V
Za+FaB8JKzgci9rFP36rvcgZxA8cBdAFWV3o7TFGT1pL6XdnRXFaEkdHHK6G
j6EJ2EH1jDHFImxqwM/fea793uwhovajxRVAuh+RybKLu5aKSxdCUabMc1tl
8LIdOud1CPi9chYDYkoW9jnhtiMjIU7D1o0vsnn5gM4+BqC7RIFV2RlHFp6t
NkdS+Uco2eUgOkadGf/yiaIVRDeaRTFCpetZshT8kpp12wl+FiVU4SvbYoaK
K4xQb0romtrqofajnEEGunmV7cm6lruM8FsC3OnzSqPpzDazvdPNYfThkIJp
IWY1+l/un8xpDR38OVYsvBgRvFpSFKwVQOK8Gy3IdershrVz96S0iB10QV7G
PzDqP9/JeCcruocmH94W/D5DLDpRwlJ48LFe4GfTdSSO5O8ojqwUPvKO04k6
C8fWRlxg1VrMa/QydYXbGYXUzumskqDVx7yQmf0agdOZrglvite1AoPOEELk
ZkShTO4VsLWyL6GAvxcfrhj25bcuBq51bCXvydfFizamxS+uIY8DrsnyE/DP
0niRNO8JuMYprceSHO8iGiXIQuQo3sr4tTS8YzoQOqJcZUZoixl+BmtZBm0U
Bg6LpepjOj+blDhlJkHiiN+n/pjoap++gibxaGxsdUr6Xdjwcu1GAeibqzKG
1Sb114j1A/6kHrbGz4O4anJRqW8N3IKcMFRvM6DmFMj6C/bDBtQvJvdRFJQJ
jHSBnfwY7mMIBJHX0hHOb/6APt0NHmv0OQxp0Pv0Bw1M9bdn33uT6BIsgTlO
he0IZqCHAnzjMveZpyUhF/z6VTEBWoZ9cIcYadX3InjQEGmjDECDRjfdPiP9
VAxxrn5d6zuMLW95rAyRSuL0zBCq6P1OIam8Vaq1btqSu9wEpTmc16GshyFz
pisN+rKgMrmfoq0EuVvA8oa35g8rg06lE0rWIG1tOQSE70/uHL0tfqO8swsM
DlxA1vGwHKrUbWRCMs8ArrUYa9I688lfBDdjdMnKq422f0wdoj2aUGVMelqa
iaZN6ynSzlVAkKxkYsQpou6t3ukWay8yuQT7juc6wt1y14nLUNMk9IU1UQFo
1wU+FgzhaMuizz7oNFHpOfqAXfB6QlSiVnmvsOFRiuaiipxZZSQrCyPyz1cn
whP1kPSdGIDdz19tP9fB3PViDs7y/lD5+JEYQYFKfQm2d/A7UPvs/anPnuhx
DTTVqOa3BR4d6BIK2MXdHenuwoTDVdtXSYjKV4G8J70YegsD4bV3dUDtN4gR
QB2hOtDoKKvBZPNYi7kxeg7a1YikHrFCbDbfbHJCu5I8LjW7xM/z5ZycLpIj
kQS0QHM0Hl1bvpzF7OOa3LpW4hXkEkceFETM/7jDVLCaMnwNYvHxsBoIwtc8
h/YqsDETwfWwuSDC88464ylPBpjgFDS0EkIskqon+6RQ2mWSn6YYTbzGgsLJ
jmybIlsi9ccEtvwB0yjZUAnMw9LEMM4Uu8XJkme2m6iFhDidlruTRAZSsdQX
boBlJ7E1SvY65EnlHhTJStnQzzRw/L5TY9qMTzMjQ+Si+ZItC8Ij/Ig+lsic
8FO36MuVwkUI52epKSD6BuVIWtxJ2/8A9tSJ8SSdL68GqublG+7qz+WCdfJW
So+YVevGchsZsSKoVYO6hDBK9JqtO/UqOw9W3jKsUIofMgQPRzs4hBYTdJcx
3CTNZTTV5jf4kt1MfPXiGSROHg6ZcSTqHC0ue6e2VXRV5O9ij9qxySumX/cM
578t4JTPQ8N0Ww7vCAVzpHgN/5iDvpN5dNN9hw/k5mhJ+3alpdDzUW20wvAo
DtSvzNGF0EMwpPi0+ufJiB5FrwB2T8DRIq3S/iTs3nwesNH48iPkx+tPXlxp
p9T51VYBB/7W8Vx9X5NR95jr4Zs245aJWFAkf1HOBFW6GrIH1+6tA1pXlM53
aGtN8JcoE1v9iCbmjKVlV/urDY9ufrGbH7UDw3IwxS7RxbGu9GaEK8tEIuVb
hWZCn1Ca+jvHLn4vDoHpmxJvDPf+br/4tkEXnKtAyKVa9+3RAbNit87UarSx
W/gfzdH7ejUUQ8t/cHFJw/PuCWRSg5uOA/54PUsfyyeRxM+S1qaNErO6+JMC
7L6bxY0aeQn3TZ8+LU2sK9/6heWldxJIibplMpWFD3yjzAWWeSQEAqQKcEl0
7VUVwU/pzJ27HfKRq49+WYdUDaUU0IJmoz3uZv9ky7nXcOtIEn4aJcdo3mLq
8F6b2wMKu5qiVQUPjn8jIaLUeye0HiimeZPZ3htZpZqikKdG5qwnafddwjAO
rbMV78iqWG/fe9+FiE0RQuPg76WCNmVb+kCcH5fNcRPfY1hi6uiuyy9FVC9G
36C9aRQFQr0AjsnmX+u9TDw+vHqJj0ms1mwuiWX2j1zOhwwZs4ZpE5a4iquS
XxBwYTSzsh+zSMUZNRuBDJ4xUm8LBTeP8/pOcHa+aWky3eQveQEf8fa9YXgb
jziL/BGOdgmNRKgxM5DgJoduu6G5622I2MbBzUVmtDycVtFmblWO3Brd0l/O
pxohvFbD2c29nC1hyBtD35VBnVzbd4cwRw2RrLeghgk+34qC6Hc5V6zMuXS+
Fbnv1Kaid6Y//gA53rozA9gh9hs+Rj85pJG2WKH/S46eMeUwTbUw1PTtZ70e
rhumIucLyFOI004IVGatW7jHlu5y6kcoig7ENf7X763BjjZaYUQXnYRRBRdX
mPfXQnxNjy7A5IMkMxyLUB7VcETrQtJtuhBXSV8ooTdI5zGs5GtCxsulX7lB
HFalOtBfW14CxSw+MaHb2OJ4qXQkQu7u2n7stuTqjhraiFwLMtglRztBcJGg
Hy8UIYNyfXh0Tw51sl7gfO2QvMBnJh6phr2r2Lj5ADX7RpBninyPsZvkyvrG
Xuau7BjOKwlXwC2Snwz1hlq+i/nZkH7s+/J3eNQnOPZ4I+Ay7TrkHsp8BiwB
QQlMuZQ7RcdFKymLlDMMdbGJQgB+jcncvKdQG6fv9XMIR6GVCt1L/irVlOjy
jc5+u3tWsy6Oecu2W8gDoPwYR5zeOhCbBN3lkzFZJ5WR1t+Ko3sd+ZN3Ol2L
yId/O9owXHuMPC5aMAjtTLKBvZu4qawsFXQWepsz+ORdwNYa9ajOc3BbtNet
8Tp69r9fIT5bF4SxuaxrbXwd9iH9eAsSsEMJGyRrOezlJfopkmcKap1cGMp7
nVAJl/HL0zoN5EnHA8ui/fEyT1n+SQRgaoZ6zJ/m5uAmmTWvC0klOu1OaDQr
tfPngu4URrbhVSdndZ5q33Qx6XmQwLgBnRM4PKXxVTQ5ARYf9mQ1XGRhmFDr
IhBUPinnwwibyRhRiL3c/o1PlM/Ib2rOUoIK3a81oIpQBQJko/u9fv4NpwFK
WkRbsqaz1vzfiUXp86Dx0Or1yQaC3TUF+G3/1esaZ2075b1Zw298fAGzAdfJ
eH7GAS8FqWkX5mlgZdv3HBF0DDxjLKqhuM7et9KDOaifVjxqofVi16J2hRWk
QXbZZ2OYuT1FgQLPY1e7wUSlF0BCIIgFBUpKtXyhqv7+OhYLjJJEZg+ndICq
v/UJXBqvZpwZxHACNIis8lCFNDcyTetjUR0zmGKq9HYO+5uEpvwEnjOgMkCy
BJWKHeWyosRYGWvU4rTTGMr1//Ef8pVu6HjE0CU/9xmsCKsD+Jgyj5dbxvNM
WCt2Qo1FxA44vU2mW7tzzTQsrI6ox9SEY+CeU6USn7ADm3cHh4xKEU9j55Re
EEWujb6iFNjOaXo7LLm+ZBc01HrfeNy3arJBfdEzKBXo6Gw01SBuaGCKUpWJ
lFKrokheGi9s+9Q+rr4CWP5BvfI4qZUsv1O8z3Bwknzlq3NHM8XzQnTpO6SI
i5JzVn77CLP2B0PyfNwLmSaNuWSgWcyPlip7kD+ppiP7WuXuXwXe8Ev0Fhag
t6AvOM+heP9TvZ5bhHlX5Qt/isTf0yKVilpeRr3Pf8okjuT6/pj1oe1yAgKD
BE3CB64vMPJ19yZgNQDNhAzwx4Z0xUe8diYhcKub7G/GsmJF+PP/HPtcjP+m
Z1niwD6N0J7ijV628/E2nVvCPcxAmFf5jej1qY2cgEEVvmAxyOJpA4TqvKfk
k0U+qmx0DTlGQl7trwcA0nlO78kjaGlUnANwh5hRubrvVxVm7lolFsKt3LLu
QcXHhTGV6SbPQOdnPiTjLyEGwG2dYUhUzBH+qje4kyUofbkGfCOFkyWHGh4X
OUOmlD4EfP6QJ8ppVZPONG2GsU3tXsR5ZAXVRAdNGcebLDOPefLd9MSIU1b2
fGepBXB3g6dq1NPkuB3Cl7YZFet8pP51HD4e8DTyK8PRd0nxtGjDvsukuSrs
f7obe68+QepFTZou5JErNmYyre/hDi7AvgrhgGAw06oSzwq2gLoO+XXPDSkj
5dPPssXaT+ZKMvXOAbwMXu6Pap11SyXkLO2+AALTG5S9lDpXxIuEciBxAshU
ERrSzIM2xHSxXTpZ97Dg1AXeeJOD6l2WXmeZsNrxHfdqyKigC3GyM2svDHs9
Nd/BN2LIT9QOjcDOWeOszZ3BvwOz3l9O7jmEoqPBzngaBMTgL9EqmJnVWj79
RLNnBZ5KqmAXdG1N8tkkYIYKrHVmIek6WU7ZkymDHswt3bYZ4JIpt8vWnXL1
JHVyx1vjZiSABHu5FLSmjlL4tWpRJb7tNQGMTzUQ1J084VbBYs5tp1rCDZkB
kzcSAI1KCCkqEF5qnlC84zD20G2BJHLDw1PM0Rw/uhs4W6E4IOhLH6CEYfR7
CWnmW7mMR4EcFzAbMxpccQYOp3my9y5VetbFOLMCm4zDt9N180KFOoomCEuF
HI+8Sm7cG5PlozxGW0iukbZbwmDfVBr/2ZCvDLUdt2bSHZyTGKOtoxm/UdRa
X33JFw7vVDF8St5T9Xy++RXIEFOktf9F4DY4kFSV6agr5+OZb1NzNdw2IBfB
cM5kuz60qiUTm/AhD6MaZMfB9HYIhTuzRvyvMMq1uWrhyHQeMfzLM925xomF
X4FMwbPpOPvRNzPxnAFlcE87t8uraGkAaavVknSfgDjLsYKObqq+kCqn/Y62
XtN4/qBFmsruai5pDffiowMNxa9cQIztP+h9DlYB5D9KA+arfIBGfaf6iK87
4+ds15BS7ZRAcQd5DBAE66lO50Y4NFvIcCwobtqxHGBwUyfI5yiKAy/P125+
ZnGW1FL3t/m/YexClEdkFGIVaaCXXvxyYH8cNhMcBNHX853UF/pyTjZMNan0
RxKmG5XOSbdTXzGNVSMXpBWxD4fUrEa/yPxq2ZwYW0WSj5l1oJsPJIZBPQk5
HDDdzn0bnamQP/hIf1X5KRwxSKyml5VvL115vgIlhgZQm/cJE/X54ADLyqQb
EfS5WhE+NuosdwXDic0yhkA0Oy7dvg5Pvg1mYiokklDWY639TCOQHGLkh4hX
CptVtOMtn5cGQeOMm9NtaeUdTfUYnrNVVJR9fA2TOMv30ZN2V6uXcCNYZ1ME
NqC4JHdLnxUgz4CkAFCT2Iyqs+/xGKRK/02GvWwhPbKIEBQDuuKnQtAarErP
KNGjEu0uan4nw9qd6OXRwIrb6ACuMk6jG6xclmJQJ/9DaZ/HLZ33i9H3jG0u
SL8pBZCWFTuB/tymsmYjkKnda62ic1PA0T/VLm3DpZGqZ+YNrv31Hct5tX1K
4Nc5Qfocus9lxwxa03Sdz96E0FcXRJw9bTbA9JfguBDOcJYcKgPgGWmc3CFK
0hz48z8dpstjtX6nZ9ndRWjmHQp9RcJCKKHAgLNFc/vhiUCq5lK+Is8n8Tbv
q+wpUs0kMvSjZl+XXXg0UpbLJqeZzUrSDwbVKyE/7QdXox56hJbPn+kMs/6X
LSiptKAeRJGZSL+d3q1FdAB8Bhbp1hXB+XQPOMvhDnYoYkX935Bt0zB5Sjf4
s3BnSeJvN/pOqXiZWfnUHzLpwmsrlsiRx7MPfQlvVRMQkPGrnwYeGZoLCXcn
m5WtytQkoVL99fnLv6pCKkKhCoGBSh2jTRHN/VWPOJx1dt8hLMAvmqvBDltd
AJp+e6n9IBUEQfhYuew37BQdzM9PWRXXSFtBRnyHTYSKSzSTizIxxijarq4N
5V1J7sOpZTKfhj8EO3weSS2oubmKYMqcbuvpgvvZo5X+p8CrxYPVDfFUu646
hMW8R7bd3Io+wbLHEErS0Q1SSYFfJdkQ1bRiEjpPdxdFTtegT4O9KXdDgikY
aid1i6Ve6ff8D0Q9SZH2f0FyceGC0Q2bkVSG7KsfL6sCJUXcCA8qPPl+q5CU
JldgX0naS3pmB0bOR6w8swJvVMK2vL/gASp76ahwwFjYR/QJuqmLDJmIK/x2
0gebaeBRRgG+jNfqSH5Nz1+YIO4mCDWTQC1fqHUN1H5yTYkqFhK0+YI/Qcfz
7lelmaj39V4EPhWkHx5VMzRHebwc0cpBHAHZ13+Kvy9acRZVSud1fTtTA65m
SfI1IpSgwOMYAzgY0Z4zWXhFyx0EvTMY2YujR0Se/W9VZZDuVAlGQdqfgIpf
ce02mP6XXhLnM5sR6O5bBPfGmzIJDzaxOm6AoT6Vm2eECWiiJVaMLuJP3VhX
HTSVnyRFh0cA8PSJvMM/jC0bff7H2uyaAH8iZTdADkXAjWaMRxQDhygNASZA
QKcyamqDsuxMQehrNGOEd7JsaJ25unTuwjl3A9qjG+HrGqrvBuIDsc1eZ6u9
U4/vulMlNDWeBz8QQnflffjDep5a8OXTcs30rq/rxHSgJiicqiC/EcZcQR7e
t+IkHf6rP9xpMFer8CbXnxGgDX84PziNfcH4g4bbpiUWuUK1qB12uVuqyWsE
t9OlVkrEpqKLLopbPxl0ctvqccYGIp2tp47ATzXnvnF8oEi0I+HWVmJ3diss
Vh5d/f7ea/Shhm2yznAOshZngvQdohu//ChszISL8dBYEGvvoOtjuawEcwIv
G7/d8f7uSAGLd1shMF3LrOt4UgWVsbUnT2/gmMeLqA2C7mSXgHskEPUaVOVI
cEBTY3U1HDyhEA1Fj5NAdZ+qnB1O8m2ratUQW0SDKV6X1DaXzzX3rLAQHWQ7
BBGfIAgkEW/z1C6igJPYfCEy1rHfE1tch/mauCMichv7rxm2XEsW3pT81Yu2
F2AavgBVwfQhXEbnGIYgvOXOCcLOLxZSPtS3+pfRfYV/L9L6o3St8HH2wlU1
8zwX8uI+Lz9d3I6pKly60ruYxHETfZF/wydz3Hzs2AnLYP8j1e2SJ89ThTWh
fpHx7PMDEJVNLH4XySeHzowYwVTy6Xp8sS/U3vvhUG1NuiT27Vn+W9t2JxEs
+pObKGabKX2ZVolrhxqoZchsBLjwaCNYoohcwiGhNmssEYzSgJQgL9Itqs3b
4N2J0OoZB0MTG8tbPWvVo3tYjJcQsB2IlZZLW8qEDI08JzmnLafVmawUmBa6
i/Zeb0Tjeh9ftHb+Vv9DJetGua4tcO1QadTJ+AAvTfhyOCCub+JDQV0SEAMV
O/EazFlEU2MNAepVFUqOmLHSlkdEA8hgajZAtIFs5cqU+v8OqkWDAH1Rc0p1
MT6WCm91qZYtvC4xiScJqANhIPASEqngDZgSN+3c1E15nnHEtLEjUJR4m3yt
0GsZ4DtnHj8lIMlIuYcImKndEETe1SSq1ixivHIvCbuXVcjU7RWjNk7M9DVy
JI7ItnvlYrjWK0AOb81531ML9hYy4MNvHjfzo8N8+rFegp7XeZiehhC9f5F7
IXrse5+rU3940/JTdlaIEnH6QfqYL7OLi+hTx5gcd5JYJPzCdvuXVr+X2AL+
XXqQCloAUPwL2/UeVzN5nvO387EUIzLuD3jgrwMhRrhdFm6yEpc9LICV88nm
5XX+kfIsPcG5CrcqKDR25If24R+MTWtYZEY7tcQo7IfZVDpRMZAJ9KG/sCoR
hTWXQ/Peeo0gkmusENeK/fwf9P9XFKud5S/9YUl6dNi9WvgTvkQHy3iuYNiN
dAd7DSPqqzXXwvZPq3UHhODqNlI4v+RJXMeXMmL7G2nX8zw4ch1aYV40s4nP
R4+WGACoGDBx73qt4lDGfb8rmnmIMsUBttoUlbG7PLme83oQu2UyPjKQwtKf
pcbAsXJfiedCRpegoYtHFCvdkXxI2ALOHpvZmV9Htsmi+vn729/HgNylPP1b
zvY3wcWFWIEUS/shlk0asaMtIfjKqqTgPfuOhUQtW4upUC63hINFm70We/Hf
7bc7Pg9xFQCyfdsgoefaihK3fnZVznhVrDAXREGsTXqMFy68gxZy9grjXL10
C2gHnABt7/ExsuMXWJudbbDH3SbNju3cVjuhOMivllVk7RggBOR/gno3kdaP
zvB1uBaSugAlzl7DutBApBV94mcZcXRGecdBuSzyrqM6rbnquNklfouIiu54
E7NifadEgueJldln1fhh2MfC2m42m6eHH4Nn8oOPzhPt6bVnB23SUpmEp0oG
JYxUE3okpofA7ExxFfGMX3wGQ0hINuUnbVLS16yi8Xz8/BeJNN5homW2FW3n
hqoBeCpZnHLEDjP6ZHuOSjtC/XS1w8jDck1MH6rrgUg9LofHMXnwpmUAyvKl
ZW29EMDDrDybRj1rZD4agmonUDvzUk/9ZhVuGSZIXVEKoSalqRuxZBF6WYMh
C9uOe4gGd0ATaRc4CUnbr1Sr3OS+VC9YZwiGSFw4g1E+3hSsbBpaBcBLtzwu
HWteMjv9EjqJG5kvZbLpDg9UjPWCph1zMoCp88p7QMc0U8A+3fNO0oSqEvYs
+ep9/wM0w+zJva6+Mlo1IxyxU7252Ak3/W0eB76nfmQDj1FH5Ky4hS0tP4a3
9oK1gYmyfnDc573lzFgCgyIJT9acXN2pJOxTOP1b41lu07ELqoT44pSb5kol
nbudZLcjgDItVQGTKE74lm/WDqdPPiGLuM1nNzUwPh29j/AY/XTd8CGS79Kc
d2t5JGOgcNvhNjXPT2lQJ+Le3gsQMlJVxdmSH05Jpw6eMtDhdPC7+SV5xJkQ
w7z1EN134uAve/dqK6nHY2I+4p+8SNnsGzWASutF89VdSuX4bZbDycF+Czr0
9G5e/lQLAjjUmq9VoiBflef1Qm1vUTaX/lSLxWK8Xg3Ot4SUg4FznU7K1RMy
uP7RXOMAvI+aa8N685TXqi5IGjQwQbwlIxhFQ3PiyQHPg7avtIkoQU3137l8
NJ2ZUEo40rp8UJ7Q1QV1GfxuN71K94E5KOzphj2viLfwsy3399J0nKP7GJer
vw0MUGsciYLVDKLx4XUy+HPUL6wzi80QDrJHPQBwOFqSYL1ZFIA/auzvNA1Q
4QFwSGvvIWD4g3KI9iAFgh49XJmX1PoyGmvHN+c2JyySYWBClT+Owwdrfmpq
rjvJmHn+q6oW0kN/LcmjdAoGdIf0izIH8SSUyANlTkdniiESx0/CzXGJz819
hdnseCD5UKQtyFzZwGrg5NJOPehmuwmo9VlbbBBeFCMQblSb2TrDGnF2zMe4
m15z7EbSulD1z3cIQjZiBvnWgQooPDERJZTIqCs3qbpc0IzohfxMY88Sayhl
B+GtRWgGlBKYcSEg3RwqKmSmFLMavnna7/vlH7d1vJXK5dnXz9jw5Zo2KFUH
N3s7egDn4u34shNnaMUATEr1CqiMVREJo0vYZzqbX57rx+26WQiZkE0sIFK5
Lf4OLguMTvHu9rihoAR3W92tP7jjCLY8vCqHg898pDMAHKS0op2YEwHLgzZt
Ctfvl0Pb+TD/TrAyu/3ClZaVLsfAyYK9QgVOJR/8vI4NXNwCATRFygrplf3L
JP1bxjrjTs1jiHiRbXCLOA3sBcoj9tNIlz9pAQZmTw9IkMk8Ay+2Ez+e2Zfq
z+izhTt3yG+KHlugNElyABPbze5g4j0R0NIo9mVATtDHvode2SgLYNDOnbms
GUK+BIlfVCaJCwrEziY7fmAh8GV7yLzHCe4i2xeM8wDLLU0tzuJmKOyJKon9
nUz8+M8LCBgJZcpzuINXBhQ/v9mSRS2zkLfcwpCtBwYvAZAW95RwFkQakyXG
5+s8D9UTUhbybG618lkEAYB7T2U9HV/JX28S9ja8ZPiu7lvEf/GF6TCRZ4na
AXSROUpyN6xBYmNQiyrtUdMAFXzKTC+OaZyBYh2BM7ORqwIh+ZLZmoSSHRP0
aSQGwUIk2yEvL5HxN0fVOV0I5/7gi4e8dqYC8Y59fW8jJOwEGLvpYbB9IvP1
k+AYQONNZ9zY4411vFqjdrNdaSM1pnwhAEeULNYb86vXOZgfVvK48a+8zEb8
u593IcXXXOIgUSUQp45HEUdaFZzEYioEfFUh0yw3eQDB3THKbagN1Evdspkp
PbG7Q6bmhiAxN/nXhcKJlJV5GQHCJXErCG3DA/bgSl9tw+qefX3JC+pSLc/S
9ABBDlinacva/T/O6vNqZYqRwCDDyj26VJROjEJWSzkw812mWsFmk7TSB2Z2
hO8s0pViLxrWszJ22WSMoylR0+bMIhIeQ2M3gQ/J2KzLeG+t5Dg17RT8LyuI
e5FeMntyoVu6/AazAzyBh84icF8jfqnBWp19ze20NQFLBHwegTnXQTpx4UA+
b7M4MpA/5mQtW7ulUQsjrNGzNIjdmOr3GkXD2NBsaUWWFmajnmwsL8YmAU17
AA+vWEk7MdM8uidEQgYI5qwNhEjcVeaApLeD+XR+V2e6hzszsDj2/R7dXVjL
CITzLnKX6ck1lQE2ZoMD+dNmkyZwyqNwwMelI1DiXmYFW0C5EbmpDujmFZYc
em6DIFFL8NACGat7D59ZShMD5y4wPtxavC/OBt94eXNqI9vMuwPqtbxbKCEK
8QetcRMe7HLLGq6s+XYI3W1JJwJY8/UOPbySQZv/XFhBppyZ5zo6QjtL8hyL
Hr5/EhAZWTlLgcJLg57gPwS0/8taVeVccZtZOu0vPiBqv9PH+2AHGtWI84Tr
uwp1FY01PSujibd0M+8pns0ZsjADmecW+AitTdSfKA3DjPKyx1+FtQM47ew0
PuJJiqIGGBtfeB4RTwB3nBDfAahn0RLKkKuGI6li/IRy6rrMkEM3EHHMCRqN
zrCUdmQQvhNuhEUZghWq8appuf7MbW4RjPlZPH4WL37X7EolSHe8PlEi5y3T
JagSIXiHLhi/v0znmMhU7rNT0Ub7lhKcIF2YlWlrq57C2RFZT1gwFvTiaDJ4
rxwzg/H4BK9txX2OER9w6cxk2HwWMKXgvGWfw5ETIcuGOvkKZOrfH50Bp71m
HsyC37r/qHJKlZ2mVg6oObDUY4G4Xw+DNBkbO0CpHh8wVEgbO3LSB2D+rbwa
VFlxpWxWhcMFO5Qwmm14KJyURfmOK0E4XILE9odHKH5Ntn6PwbhP4U3mMzDm
AgZ2GA8iexYKuZEEwrzwu1OsAMRAWxoQYfy1xm0DiaxTnEbwAINrCeBFHoJm
bzZ5U8GadsSOAcl9CzoJy3NLnX/yMtHzCGDmqcuTzNaTwhSk06/YNMpFwFDv
b7Qt2BCJ+bnGiddWHZGQiYnTCfBrpmWkZs4j7OCSTBiHLTGJzKc6aQ6Jeo2z
Zmq3ap89ILrknNG0xRCye8FfcuRC2qaZyyS7Q8+9z56oYnHoT4R3M146Wa8T
2aSKHRWJidtXmuMhriKOwC0y+OjNOdyAwmExDbrAkcT2E5qyi/BM3phQOS/y
LlqK+BFRTS2cVf3xG0DS1rZYM/LN6AQye7eqBllzSK7iL4QfevA4j9+Qz9HY
JGVeoK21LnGCT1panU5GpTFlgKtT4gn7UPZV44LY+fDnzRWJyrjnCoDmE335
UY40qpT6GvkVGN6Ymwfbab67nfC/LvtzlW9JknNpmqZBVazMEKW84Fj8bpBy
BUb9YsqNRpLVLM5e4VNb/yhkL6qtlAoLeTsKDzd6PqQi4NloQ1JzCBRosFEq
cBvFq12c4mo/H55o4NaHWliUdaJYDjRLhy/Kj4wi0mXfbNaJhHjl2QcbEnBG
b/N2z6ZiASx3VshUKM3tGJAPkQtQEpoPIInlejKRQKTBNpvcm0rGll0pA9LS
eilGwXl0f9Vi8l3UxwmCIooGEaLai7PB3yPVkG8OiB3xIdVJJwMeHWbLz7SQ
+KjZ4o75axSrdTdzkea1pean6Sn9GLeDgURIDV+jNpk3dz6v0AkWkFsbiU1C
oDdCaVMh23H3zcwEVxO/PLxh/hwjKF0C1oOSbG1NXZdmAHI4eTTjYFk2PRSG
NLgKHAfCGJgbl4e7wJPd96WFpdoFqOTeO1/jIJjaaz6KT3nd5vgAyeYYlLFC
NY4rwCJ03IMO94ulLCJDQ97Vv7tijQbOQg71DwaxNG3QWdF/tDyqZK//uXga
ITQ2wkaDDAmu6vrMvQ7J5vy+noMpyto3m0NwHjlszueNL5ZOMXHc6LqLXWlv
/N1a9zwzYYFiRzvU66sDLlSQpoTMHGg50lysKoueBuy8RTUTnH2Xz+4g8aOI
0EzscWKJ89SF2UIBC2yuy2TSdZd+/ut/OTasNDLtPYlYUVOuIMWKFwCCXALx
wfZ+Gu9C3g1l5EiF8Ci2sMF2nTEtRiGtTRvOretFWsq0+oF57H71YGLKjoDk
PHSemQ6E7XgTcN8qxuurJixL/g/43icYqqMR5CqdUTziopZz6uQbo0H82fJ7
ct3yyxYYUsw4KikEIUOaU5g0bfkjWfsdk27B5XtKMZ7S7j4CvE8CVBBYzmy0
rhmZHwAWdLwb8U11JHLnc/7d+jmQKRa8wahTeCaQJh7FvUx6GA9XeoYvnQgN
cwWdLbFQhvbM8UjKPjhZTpGno55naAsSqcy4E+1Ucdy0IEW/wUMBRKytTqOQ
WbDniVBsx0bdP1J3Y+aei8dhqnUXo5/LSLW97HcRxkLKOmtFQ0wdC2yE9bHG
abAf+ByZVGmhAN3EHT1QJkPfx0guhbapPn/pyRb/CB8fviW+qH7ZqLXQiYLP
d7f2pJXObnwTuiT9wd4hG4FFiYT7QVy+Qt8a1T8qE8t7jbZF5P93+uNo7Rf4
18wvSutr4/oUvAHMuEnFg1EWcsk9810etVLpQ4SFd8M+jHzB65YRmzUWY5P7
MqIjgCc8fgQLIhQygOrQUpVnFKj/jGKK3to4o296U6H1eO3pc4MyvGQayj2y
IB4BSTAB2EM3/XMgeityt/joPP1DfiRjC4hmNqezIKeX8LGCuhC3TfWZHe1s
zRhjwUiTBx+ii/3xfwhTmR85eyzZVUI8J/GrIWq5f3VpbIewaJ3Y0Bm1MZ+p
+rips36ODZ2IZTXw8p+4qgHA5dj5cB+A5r2sTILKzcJhnHGEosxg9gbHu9BJ
Q31cxdrX3w7ww1JQcJk3ZBanpIorHykyr1CCHNrv/OMYxe2kA5vssRJlfTON
LB+wSx778s8hIbTZE3PQQh01nXuUalh78MNxDKsNiyxXvI8xDYBWYUbzBd1l
mmXfQph39VdDM1+tyEve+ZSwjam2RrO5p1+N6KCNPx1maiqAXD4C+/3MV+s7
9nIqP1O4cLT7LaBuzyEmuY+5mlKTtKMb+YYVT5EqSVrW4crqt2ELjiETFK+4
2GO3//XdP5PxUvRSFzFYvF1cO4cPABwLzyDYxlt5D/Rbw8Y3R5h6p7FdRvUm
2+V7q96W2Q0CzWCdvaGJ/EaPDr0DXmpp3Q2oDDehyaatapgCoiXI3ttJA00i
amI5xmh4g0OftimiLzFtU3tM9/iY9NTDrhb2zXr+Sin5vtL4atC490fZ6eqZ
sIUUUf4/TQfD6EPv9IK2q6AZ/yjQkcpowIUp/dptmiHy716qswnrdnRK0O/X
co+Py5bBi0D5QX8b2cZJnUsAE28szlM9eDkjEvoj9rVZP8P1WsQVGrjyTcAb
j2G2PggmLqOqTcM7GmCAlVvtLWDEbF5fUb2K2JsCYC3nuXtropXYQBm/X2I3
9xzF2L3Ym/rd1zN8gDb+iKkRDqxVnJLjSJ/AMcSPvxM26DZB2MwPp4R6wUX/
hgmwj96J0o1ZuH2LW+51RVdAqU7UVf9yE6p9tsN5uIGbErLPg55OUQmcRAw4
krI1MRA28OaC0ThTDXwCG81bvUWyiw2El6ns7Nxr8JPEKalubBrFU5KM1G6W
CPBSq5/5BxMbp5sC1suLW/YeMxiiY2f/C0F6K1Wi8UJkoMpBPY/lBEOb2zWU
EXiKuQSxbrnD9Q3dzzkEf6LdvDJkdyYGNJU4H0uybbLYtBQyEgu9/rxhjTkQ
/cpD3C8aR/Yp3tT203WQ4Aege2kbTMcJwENTtW6DrHjTSlPnU2cMXQkzgUtR
c+hFaEHuhj0vWSm0UQV2dWM+CBAzrVnnR3MTLdKR0BKs8FBx39/mEjKRpqhP
o0loAflejoipDh1txAxNxhWklegdYRkqA7MtDLRXcLKp8wc9rzZi01FgKyqU
dlOWK2wxsLTCtAxiQkalHsJuZiyGZt3U8CRJp+cgysPpZIRUbI1nPdtVFLpk
l0rIRAJ23F4FSAVUS0AvT2jXhjud2omInkf5iuM2OXeZZNubq/4oCf+KtlzT
y0cwLiwFdvOr3D50nU4e+fFKx5kcHhCBcKQWPntsJ+VFsnnplEmMeQSDk9fJ
AZtai8AssanWcWj5OuedbsgWKgV1zUXMEYQ5BI+eFEdddccHXQV4jQMufTL7
lR+OZvcZHs5HgLgCXRDWQlrlFJhKo1bpJ2rAmBBHFWYzTDVFuMD2iXwSl+KX
yCgNs9Q4++hxwLE5eGjW++8zbIMnSkiPajGAu2dgx7s3e1fAgt11z3lWk9Bj
UkKRzcO4NgQYEyI10SoJiAz/tHZc1Y6maFPpKEkNbwV5IkFvCrZMEidJaQcO
0fOkU9gg4d07Ghon2aVdK0+uhe+UCAqGFkERsnfFoadmQ9S+L+VaayjXhn+m
UfQy1oO6YvVHRCt2+E25n5UYFWsr8ySI2lpR3bJ54eLbNMnbK6ovGMgb9lFN
YBZ+pcDrG1X4UB4htyixKNBHi0qpimIGkCdaWcH+StbS8ymhrd/aRswd/YCL
5euLXN47AEWNshYZiQ660sMR1xtKDTUc0JCpAcpaLCjR4T/t57fR0eT4DRvi
CMQXSwMPJuHq2b+bIJu+04ulYZas/AY3hJRF94MAxuy7s0zwLuDKk1/ZoUEP
Eae3RqDUALqlcWaIyZSba4DGPrs2c7rRSzCfdK7bbOi0EYOC5+HJNWPArVGd
40nhccVoGATReL+O4LF3F8FOW+O5IjIuyKcMRYiVa67TJcC8YS/XURglmQMQ
+goy+Zt0AKMDuvizNot7Wfdx7Db7afaXeamfGVv540FOqFe1DV1J0i5CBdk0
i03/FX9uDB00tjDNEG1PZG1f/L0JjeTaiW1UFG0srwJsmeFgdYnwXaufZAD9
vkiAkG15/1SymJeEj3txiRolHRQHHqYrqynoCtMaXRARiLN3P8u4BsBQpry7
ELP/5zjtapmtGeVl0uuo3KwIu56LP8V2Pp9pTDbyBmeNd4lzQ028Zj4cwex/
O3HJczZzzldoAc4gCfPueYngunULCt9o5900c3p5DoVaO5VOojnNzsrV4GZP
wDBjxy0CmRc4fyNJl5F5QvSKXNFiJXO3TVVf2qFMZGMoxm6VZudbkeoFIdKN
ioFa+hZImCGjX8y5OenHGaKWv/TIoOFTFoRPgCT1TEItyNUqW/F/l8zqH361
sgtnXLkrHV4uFGTb+dpuz6BUZqcR4or4Wo+UfPNyj/vM9ni/J/tR7Rwd+sjR
TmfbQgUoHu5aKa+0hdJUlLu+DKz4ghJEKFszegbzFPVKVv3KbzGgO/6pQcTI
H4pm3QOA9FnKoFJIBOb6jVc1sjem4xnay38SvLA4vvdpINySwT3vcHVQVVax
MSgRQiIllyUlVtEbrGMU0V7qfWvm0hoardAY04jw0fC4+v3vzzFQYzVU63lE
sxh0enycsE/hkNY/tQACOMDavnqDrojVx5+OofD6A/hr1DmhWpOlghQl24Ri
EQxHI1grcP3jwtD+D3G3jliK1VhLnAw+UCJpBNYY26TAbWCxBQ3cwHP0wiA5
L8SP5j0QELzI7pzZWi5GGRzlw1rRfH79j3j6PMsl1oOMmZ3ZHbqMTWVlksIA
9lEBPrMW80fcv6wsWU+ya/mMQR9xbyYbeH7FD2aOf5ouF3O9J+xrzPuIkeMy
hYX6dwQX7+Swk7oC5iUsVZKrPRnENvTTIM3GPTYdoasgVzDzR5/w75gKcGEK
9bo2aAoG+u9iB/rWLCE7wuldqbs+V8lUSd0PGEQhuR9nv3boqJ+OTbq5aFv9
9KqeWkNrkZoMBA/dApc6KFZ8E2zA2EGfx/2pAdIMnovoSex52R3yvTubCtsI
dMf8EiFLu2akAf/UUDrDXPQT7W1IHhvV6u3fHcOSNsOFleodL5vT3St4uiCa
LQ3QljxnoqzyFtztcSz8fCQ6mWE5z4Qgh1kVqzeus+X8gItPLo+AiOxarntg
pkwPgeLYvUuPamIk1SGCnDbK6zaEwGnqOG7w/auIKVt0XxyPIXiCXUlXO8Hn
77+A40DIBZaLtbdMkKqYT6s/n4pD3TAun9w2TGeQCHeaaYALI+7C6DdtUh3e
VhSLXgpMTmMgpHe7JCvHf3jYVDkGHjFysj2hFYOJia5wRm/ch9IsEtzjgnzk
wURTU2uM25KYgD9vJg5vRMB7buE5vJcC8QSKzgEe4TSRvWbyeP88tbXShgxv
8TsHD45e59R6pwzA7Dx+1aa9g9UIPFE+RffueUzSt9yw8anGiRYYowdJRlWa
aoCPx5KBi6dfb2iNy0qoy0fOKnMOMdTIRtrjJNihHWsmU9HOBZA8SJxKROct
NQcwO+IqjacOzz+Uum+zZvYJU2OrL/74r96J81Nz+iFQ71w6E4Bou2S6+ohC
T8AuEXQbO51DuRIrs4hfnpIPp0Bz9Stnct1TvKDma0kolLBjVdyGJB2DkQ7B
u3Ba8LUJ1FzsIeo/YTFdqw64ckqKIOEJoDSWZsrMlMl25/lXjkMSyKKbwe6y
cCW+WEn9fWmP71A17bLlO+UFR8ZntH8Gw4kVaJGD7L6NyDqoGA/9arRRc2/U
mqBHPmVSMJf2VqKRtyKzfEGSJNtWhjMYeJNzRnCvCbfA+DLVVDAIE3fjYdyU
t1vgBn7NKm5Ok1MuSp36mJmNFenPDPHiqjBP6yv3PnP+2Eyh+lZsISOTNle0
4hIZ0ileeizUJBXbtR6bqa1XvtE+IY9EO3fAksy4b/UpdXR+bhhH8ZagKACK
vCux+HzZdlCFNrR1reWuNqaU/D7VpMi3D2SA0nMATaxxPT//ehvuBSXOiGNE
3NnlG30HLaEck2EiLyzrjSl54ipm7GLyqgbA+Iky7ksKoaEUCebPORr7agpk
W/2VbumnxD0DlZ1PlXh09pBJjnzlKxCTRmDa+LZjPTvsPYDe3Cd6psWvMRGa
QFizdqFXcE6DGc2gC9W96OHlPrYdr4xWG8ozRzQDfSpZIVJgGFM3A/1c/M+a
PHUuapbyu/yKEoBN8RQ2A4nvkgGEgC7YtllkXdP1mfSf1KSmQF07wSGSEpkY
gpVdJOjqQ/I/JK4OI3o3M5xCdp1BPJsVUgN+UzeYZN59pkhy43hbKFbst1dE
bKkguq0VUofxPLie0zAsJ051du5cMlFfKLgHlWlje0QvufUORze+1OtXjDXq
FUXUVb1WmfDjzn+fgSUCiNRlN2p6ibvQQHG+WmT57/J/9FUVtOcteIWK8Atc
mETovz6TLDngI0UQNU7pNf4+AJJFbY+0zqWlRW4mGN+6hOdja38AmvOLLwPf
HLzfxZ0+dXrzuOsUj0czPoG3trmH/SeK+OzZBYZXLtkyxD6iXhgSQa4FelmX
PDocTP4ip05C00gk2L3AizC/HwSOoBiyuxULgIXNRvnDxjmmS2q8/99ltO+c
gs+tNRoYBw8OTfRt7JJgjqYr2CBMX75MeqtQeMbIkzfbyixIIK+zMNHHIA4s
3nNILeD49t1wbkHkVSlU4efgqfDYXR4QAES8E9kJMXhVyCQ+vm0SiVpqR9gh
ZRIR1OkH3uewopa0RcX3jp1aKVwasEgRmqFX/lCjWTwE/qPZ1tCuPmboIxeP
2LvKvnAIU/y/j138P56xPU8bH2BUGAOBV3JDggJxrAHleDMfD/Ju0PfLTvMN
eeY1yImgKRoJKBla0KtVeBWEUir5LqF9hQNnyp69e95n03YMKKWYCytjTr0Y
AUqTu09N9w5V87HzD/uBsdvzjmbJm3a70B3BWc0L1+Gop4GTIHIKEekw6W7O
HCqaDqdYDHSJtKlSnz/IvGIEVVQkArhn6tGAFWue3/UoWMw9/Zx+av+M0wR5
S11jEn2ZnpSZQ37+hlZbmfPrjFysKoPvRHwaOldCm3SjDfHJSZJBuz5YvEYC
S4v7CszhIK/3OawNgYYDyqela1PPwND0Uvly//WYo+dJ49MY3vLKMZgAMPO2
56EtTWpoN93aEB41rA/25m9sLBlUN5njzKLS3d6dIro3oQhhDLDEaqp3gV1H
aHB7U4CAj71ulr1Ao5Xu3CZDlUTP8hu7xvJrCTU7tlM5ZHmXINOVf/kpNoRu
SofPE31wI+1mpZaJzuuu7+oYKkr1/5oufA6MXZK5prcqXhNAdElDt4J3uJUg
Dw5pd1NWKGl+ejh2vS5xOT3MUrAlxPD13fr0lFVHKTU2BeG30pOMw2RkTMcH
OcJTmDmZqbFp28rX3a0rTwnSpMVb4dPAF7Ej7U2xk+J9ef7maM1HSdeqV2qC
N9CqrvmeuYD/f5ILmwgrjnJNF5i1Vzlu2BrneLzV/I5e2+GYhwK++sZYexCr
Zs7CL+snlOtlyqqrt5vkh3V0aiHnuLsS2iiRYEeXJOShk1gG+w/Yjq6pyYM5
nsbCCrDbgjjiFRtu6iOAOesWydM/Nm3m9yVLLggsytqad7f4iJIs4E/kTKFT
Ihnh726EuP4yJuiLqXSusORk0r6zHEuWBUBcMSg/AYDx0jmuxdEjjseJsf9w
Hyw1ulNfhGmjyqcKECi8cEk804GqsM1rSNkm52NGjJhb03bgsUYc3tEig93i
XihD1E3zeBjrS03uQeGXAm3NcIm4eKmd+yZsJA6668kflnHO8m9VF94iOAa7
bmUPSVtWVK2MO1aIclHL/g4Z4EOgk9kLl1/hfVnTvbnC+fXNLthUGiDKvrsP
E7vjEa6iYKrfcWkdRmh1tS7IQFtC1FKQTg640NPnM6vTE0TXlKMRzyDQlo+p
91I9gCnsK3mIpDXJX7UHdDd6KQo/YPEOWbV8PXAXTWppiiuZuFXDnS8+r/5O
KqSzCqjkgxZ9XUI3WxrqPAkx8RP4pgbnIP9agriTNZ/WiV7qXSZrF6Qyuqwp
9iJzYEPR0VtP9P16eosy5gLYmBoGU9g6WB6FTG4F+kB7eyUmEBbQVb6vdy5E
wmts4hQH1JecdiTBX8LdpL5ePFHoQmD1oVUbh9PEVloKxpRfKoX+bzSmXzi/
Pu8AauAYfZ/H9eTholdYA3OOV2s0WuBkOBCVVMcsawuCZc3iv9C1ezwIBcVZ
ztCf5Iwr+yN+O9kYYiZRvcCdb9XIktBA2BdYQrTedVX/EfskBNWg7LHJsTcv
MgMjIthPtitI57RtH/OAqsCoPkcGOrd61A2qpgVZpPHNGiHVJs12zn0gy4yq
aE/GKdv6yxvTZqC5ebf1tjDGCNE+Q1XmVq/93jJFMpA8wZwiG7bs22aTaY0I
CKJA/MkVhejxa1ly6BUNHtN3Rprx4u27rUnbQaYWRTDvXN2Hdy8eY98zKzr6
yFxouNNHfGQGWkAe6lsLfKsPpfLBlNIS3r0xP6Q/4hZOsmZIN2c1ZSsigTwj
TwkaA8tSCebLjZ2jA0WlOTHDAGqnA4X/OlBH7ezvuerVXNNTc+31bsDpvtL5
vFUGOSKLxqW9dsX9mfxqimA9YYenB/+gHQNCCbF8CsNwBCyqybVqazmuGGjY
kgO6kJBFnIY/3TmhaT/YnhNrafqz56WpoeDK0agUYUDPvCSSwBLPOHUig7O2
a8p8pIQPkGO8fSCBGvVIrqh6/9ySPEcMa0skniAaD02y8oTn/TIzUGHVtRAN
7tkyzTc+B37udoDpscbGgwgf3YL1NIt+mgqgzaANr5bz9HI9RZAFKUAlfYun
/bxKP5RAUhXdk6rhbY83G2o+krM4k9gtmv/s78L1z7HCH/iNG/SNz0wCRR44
KaBInwCef/MCILixMRC7w2jPA0HMsiCMvrxuNzqZ6ROUyeksA3vhX6dCE5/m
CtZ/sIp9Jt1vCDYD4zThqS+yoiXJDxQPQQTS9NUXefCDlojBnv4owYzIDP9N
82A44kVrfUCDwxfUFdPPy3onhx8qR9k7RSOSepgEky7mzRZyoC5Zse7s+1e6
Dwrl5lOD251HFAg74g6+NRizeaI6F9ZF5kqiYF4ztnjvyuhmyB4fGi827kyd
r0zEELif64mrzJXczCqAZ0uwRJ/UqlpXUyHjfIp3EnbN2tUMPPvaLT3rA9+1
jNoqQnVGeRt2a8cIwonzYlKQvGXtuCUCxW7MIy7yge51H4jhRsQYW5kn8iYn
FX6F1UQ/XMH6QIKtYgFPDu3GzRYgmvvg6imRsFepOhGs0A09caD9DvbW6XlM
hbK23yCDbrhKtyfZiwv9h4Jl34wIFCpTvupxuqA4owqshjjhz5VC3836mrjJ
fujuYWMty/X/yBjsYBVlVp/j1YWxURQgi1iRM+4ccF+6gDOBTZO6UHanGSfa
WuRzOGHjf98DEf/dsfZxgHEZUPUNLNcbnzXBDCuJJs5JX20jWdlku3pmqLoy
K7jLAAbh0JCXMvfJ1VqIvnIImTUZkYUI2zp919mBTJ443e+xfkPWzI8+x6F2
DnsBVeXQZvN+gANkehtuNadxm80dGxXGEJRNVs0p6kRr15nbdSmHSFkMsuym
HRq6n3A3erHzD4aZi8bkBKFUhYkKMSqwkdR+jETHiKvOSgPM52Rde9zaQkPk
En36z1VfEu3vnrAFHohczE39tZZ9UCUP0MRYTw0YM3o72BZ6qCrf8DBPBq/h
uuY34CtaFSvAB1i0FHHG/ZGhbUZ2Hz2+08HSvh9wkzjj6seeEH+Tyi3uBfIl
6i6t6FpwItwYWWmG+aWh1E+4c75NoVAg7PPUxPhyvCzK1JBClLzH7nW5XSm7
7ORbF948m58w70VzCZ1qgRPyuZ/xKVLqnbGvUEu1GyYxyus2F+VMrk43bVfx
ZJ3ZurvcbHNf7FXOcfFrA2aOnERgGPs903hx//GmzLPKRrA4s0+Xc7MElu2n
UeTYJwEeoHIhBJS0tSsjctseNFVEbbmd6OQ1XNY0AVQVJjjinHUD37ruZUi0
9nLz8UR+SZnIK0QV7p4kgfcHNcvW9ekbGYqMAMi/adtNpe+mYmYkqH4Zbh9f
TInuz4JA+nXEukOSzDVuPXjGJPzIkvrvCGQ7znkUk2qJIeLApnBp+sp/Y88T
kz4bZGunnxmPuDhyGuxWhAPcX5sb+ZZe6oz1pcziBS5Q8S0UB6QLXzdaJpX2
deP7t32AGD4m49dSKA2P4JPTmSHE1qSC9yZktbyPKMjr+T8nyKRlsbRecwfs
6H0tAweCJGAYHgFRzoO/IFNDuuxri+aF1Il2DwX/oDsSt9dUMQaigrCMC8YC
wbIJrHUTrGOTihKRd+iDYW54KcOZQ2bvXgzkRa2AzbNaK776DUrQtTzIr30I
tfryPBugb605UCbT4l9dsEFT2y9Hqn7vVvOKCSDANjxnYaNhU9OKibWfpdye
faqrKoHL6jEdh32EZouEBn5cchXrSnzNghNgaEWkWQxOwnbS5zOZwwNgv+do
Nth1pvB3C9APjjQWCyWgCm8Ix3hSp1BppnFuV2V/JFA7DJpeWOBBSAXuymL7
jwOUhvkxZyCaGA1TglMZNWgMt+Ow8EQlny71mmvF/ZonWZZNii2EPp9DU7bR
8LK6TjBJhuGg/jAfMbG3LquxyysGs3792oeZjhaZYLTZflwVV3nVQxNTXFdF
XJm8wDTZtn/KVu59ViShm+zEfz1wdSuGHwPchak/UjUmphfkficWSbkarfNo
KrhrXo7WvOVxktXoaLiVldT0oInf/hgf6MMtjSMOvniAmkICqjPp4nFTP03o
IXACwOGTBUlQezUlb+ckjmQISm0xSZT7doR9eDhcQChTXDwgyescHlILWQ9K
aQpSzUyb79QLQCxga6iNUDrNY4Q9nDO4+tTATbIPNlReGLPRBejyBEOn05Ov
hhdaK9Hv5ve6Da1G1J1tpkLwnfjtJKZQL1+I39EKKQn5Y9/phNc3xxnaQabR
WCrwEPF5cwXumO+a/YTr3tXScWJX+f2W/d/cNnTBp5XWBJ7hFbzjb0SxpQJZ
B5KYcHUjnNBUzNXUIYvReuYWR/d49FRaLkTjqWQZeQAba9Oxx02v/G+KjqGj
jGtrGZAfagwSvAAom54mbT/zLqzsQzLoD/kcCVy51Zkh4/U+RzAZq0wyK1nu
GMrTAz4Td+0qmEUZQHrI6/xnXsCuKugrY988J3EqrJ2Md9Xpajqem0swxQhb
IBniJvLN0cQCfjq32KIsL6JvY+IMctLgoJV2n3BUBUShiWWBOWi2InRC9q2S
gtNkypwSZSbDWPV7/04xTov8Q/jQAbPSF59EnLIsy2FTfKcIKzoyjWO2SSE2
BX1t6q6FKfhm+8bgWy2MQZOiPbCaTpt/t2/OXaiFSNs8STgWEbE3O8GSYSPW
9wyudguPCShZZupv8NvVvriLAjLZWG9uxXxAL3fFGJBh7Azr5LwLz9VNJbRL
3CJ0V5aQngdrF67AsNw3UzVdI+1+UCdWVtxUhIUTuEO/CDIxUGA61qHkyPV3
I4P2t3JFgF4el0UyDDp1XePJPoP7AOpkfFJ9WP3B6FGnwbWoWA0iyuydoT+M
8nbn0QYOwcfJ7keVN62gxrDZn/3N/plH47e/UyCDcF/xCgzQMWy3IV2vUa7C
5AwSsxWMOCyLleUb/LvGquVXewnVnUBlH++/DCxRzt4M+kYTopcBo3+my0je
qsBWpWs+Dpyuf4RlJEt+zhLKhIN2cMVzPM4gzePv4y0Tu4xklQE8HKnOlsfI
mb+811zt20S+r5JR9diEteHhVYjlgStFSgQYdjoLo3DlK8o24+C2+sEHWzy5
x/U3/ItLKiaFRDr7N3Jh9veJS+GH3UPEPyMIPb9V3KtDQ7AY315HWz2vjz2C
fhhO2A5tUVa+jk8MfQDiK1G1jwmBb2RylyBgQL2LIVNOiqoOX8j1jbPkoYir
fhWoLL0Pifn3d3fPoQrxEl3IulgpdCFv0R+yE+Cik1mNwMUZTK8Cq/tO+G07
oPwNv9O+smFpqykMApqMVFFeTeZnkVtRatdiDXAKmHK4kSgczJ8jrfgKKXbF
Go1H6+ujEKlhhrFAB/VWP787PkVp23FxNr4HWsnJa9PLnfPL+4XFMosl2dko
Wo3xgRMfLI2Ci/VKFde5Rb1VINXkeKV68RLqeF5384dPnLDTtg8cop6YipAs
pMb45//Y30PnRtVOXTFjT8jx6q8kvrCA2v0F1Gv5ac7PNx/v/u7Km2OoUWxZ
hWi9dBQGTcqGIheyu9p7Iw1wDeEkMnB04Uho/KDV2umoCR6wY2yGpeYAgVdF
Las6eKqRwsD3cF5kKY4C/N0e7LDUkQznIMXI9QcjlCJsZljwCUYuFBFx6MlI
ylSrBhJsf1Gp3Yaux2EPSC8eoBLpkVqSiy4g6JaWxEIXMzmMn+HiL6hUU+FN
05uBa5YzEAiyYJKHUZCGnioqzB/j9Q4oB3osc57Dfdtzx15Ig3PRi996pzlw
dZUaR9na2plRbCV4BL47rkIIoShyucrTWqh+u+nU2OLFuWfqqKbjGsC0Maob
k4lzBzmajnU9qmPvKbjDyz47gXgcenAvqIzJViZjg5W7AstNTYMvRI7wuoG+
KUCSeRCkYCzXfTtm8IOvfm+PcAMBigcM01x6+0jvBE4slvwzt/qSNXpNuFUe
m1dLJ9QkwOUu3D/YefMzS1CjnBreFWpAM6Rvup4rLjS6LejwJ7EpSEBA9CMx
QxmachTbH/iVNIkCgSWaEB3+ZzuTJrbc2tPscyU461OHqAyc0gmu264mGfUd
PkEtZITLF+2NOKbcAVkxrfL7uDOBfNy5CcvIZtzi8A1/5HFyJNzl+PO9l0bh
CJvrOd+yLz7S8TuRi+tdgQrKZ1WodO2fC9ljKeZlMRDLgEcOfODALaM8TMhz
nucrrSabwGnBUI5+/aCmTvCRsnZwv+06c9iJ2g1hDm0tv2BJqTJyHf2iwvXc
JpyKE3NaIa5TmmptjdmPWeBESv/DSfXaPT9CIyic22dPkAUj9RDaJleMggZP
1cuZZyC+TJX/cbsTnwe5u6e7hi8my49xp1b5mQ81cTH76fTQcAzYC6RbIF4G
THFY4OdtPv78PbbbwZlpWqBOATfLtEM04NiNHAop87G6XlDrUkUlRGhoIgbV
EZx7rbzibTDPYUwuLs6EftvyFMUjaIxZX7rg60BUfwQE8m1iaSFAYmVoy9pr
YV8F12maKGE27F/hJOJajHHBOSG2df/kpSN8owXczWPl0sZYdA1Rab/D/0NC
/Tq6V7Ns/DLlap0XMZDkMsLdspL/8qx6n9gwyTEGnvtMLUD+wsIWfS8RdxA4
k/V8BVwTYMU7Z7M1eGpptre+VVvoILYm+tnIXZnt3rmc8pjbLZ4cLHAKi39f
3pu50IhSC8S0fL6ldFkQcJl6SjcHSDPr638khu8kCZDE591iZtmL1ITA4kz+
zt4MvqvtPhpa4qFjFfCq2iU4h27eqIyBMHiJnCJB2Himx63cUNhN+U7ISar8
I+TGKAxNtxVpJO2r8qcf0grbTBagXFPbh9fcp0nT6Shelpe3ogrsQJnWTj7q
tlvIN+8SWpUUyPR4LvcDc2AQg8bXpcssj6/M+sNTuQRX+ycyjqPiR+Y8LY05
rQvEKOa+3z7n7a/eO2Eu9pt01I3J/QX2gM6a0zSlpc6s01klzgMfMd7XKLUW
y4UOqN+LCwUpB7fu7rIl2oTMI99Ikr6dsHIrZUwiLYNPP/3CXdYbDt9/jISV
vHhw9WG96wvcIKeI+YbNknKnUjGqHcmhJiAPG0nK8E5TzYMMWmHh3o6Td0xI
EjKaX4jRBlHWrALQKTz/GiK92HyE45ij3Irk84hC1p6ztTTDHYtJeen/jZsE
pJCw3XmFK1u+qL5kKJY3QK/OnJYIRvdL4zUvhISmSoCcS78OQUfH1O29TQWB
kSt+GpJFEiYSOhc8/BQDRWlOoPgKKpxGq6Cq7scCxaJ2Hc3OgymtUq75v2D7
ShyEtMOJnO5JP5JxS0irgL02w0A/qtdFj90KUtPYzq4LPYC2h12A/J8Er3Oy
8rySEVDtAy5OQgzOzS9gbaoU2xWP83vtf5EAB95GETA/vrSh8BtlGmI9C8qv
livrCmNToHDHvhbdL3GNzP+emRSqjsY+Xyslf1z8EgusiJZnOheRij4XEx5R
mWKJLvwgdkciQfUN4IyvEKe0ZrtmnNO4oE/dvQCttc/kgx1bJoFE8YDF8QbJ
w5E7N6IieuhcI6qRKvbqKsArEBtpMCEXkkhH4Fd5lKzPEDLaaCwqh+3WSAO1
yJ3TyuwQ6u1Y7Wn0d7Omi5zjhFBCSvXLbn/H+JKi5mgMLkFT9XYMr9WQodEQ
ZtTwWT4A1JnJLRjLinxqOIx4zu2g9EOm9vNl8Pbh+IGMnFDliypnxdypZmEG
xwJ8Erdh7cQr7US6Fl1ti0dlu6KljcldxrYbZHIavzHO14w7N6Lmbk31XpDe
x8FHcSBsiHPn3fV01libIgd5w3fj9WVMK+UmgF5v7MS9TDbOjKFXf5eXpd4o
BJHcO7i/54UbEPXmU8YDNp4jDIKzKcb1j0xVB6K8UAr1clNlNvGAkV9HO6Aa
FPpbAnOpG2HYJkBD6upid5R33X5f/jq2iC8q03PY7CSbOkOlkV3AtARnuCdw
A3KYEo+P9Fe4Z5IiopOJyT0UBHJxsTf3GdQgh3wf2LD+v7BJreetni5kh1GN
wwA/vbjtopJAfK8PpOD6krcT0zzj00nolwUMjwzbJi1h1l7vjKDsN6vM212G
AACta9unJVUhcPpZJtLi5+XuS+0tcPzMtBX0FYxMPM2cFcVTRc+s/0xtPy1w
ne+Y/y4O4Jg/UUJc2OzboWX6o/wSnM5v5T5j6irL+o9UZAK2Su6tWCuMpsRE
o1yF6nFVfFhK+yxoK4LbMqgey0xb1MPh8oWYK5DM8nm7pyFIG3nNBu723ebR
qv+HfSuGVwwaQNmEWAkMG8WplvyWw8ZW0RVLxscTvIrVcVWYbi+ffbHFAKPP
A+ppI3B6WXhIzwBb7qYeaGHdz9gwrUFT8ghS66Mhh9pLrSQ6EWN2+VeBwb4w
ThKHP23sYFjL39L3lZfKZjrfJyjeBJZApGwUn+wyDm9A6O3+jU1t/Uhna5u5
XbG0nNGQLn9W33YM/0yZdCQqeF9JB4QVT8cIhtlnmfg1UsXOSdhngBJwFHxg
DQhsmdcg1Q5lBXp08FPPyMgDYcm69XI1n1FlanhLUx2X0nYHPQnsiEon1HQ4
AYGq5as7/472112OT5fXy0f1y2NjoeVZuPdQ110OtXa0IrChcFgqpXxciXcU
WiNo1MaRd/mlmpB017TJAn/V5AR7KkuQ3nQ5GDHDbpcXZdjNc2mL7n0Gx82P
+yMXvEdQuBoJhPvyNHo9usaUyje+Dt+yRlWen/nGyNWw3I9q8LHBPlfSiV+G
+ggxLJmVZCKT/qT2PFi4U8NRtjfBFsBXGdK5fuNPeaoPAV21Rcx2fGtk6/uC
/aYjk9RyKLZXjRLEnWsFvLAabDA6OIaubaSnJbNnCu+21KJFw6g05QIz4prl
9BJYGSKTQfurW3kHMXXz+3z04Ux5SiIMKefkNxzxKpfFuStwZuLIxLPqnfp6
r4nHPf/3q+ypYcLV+rEtC9vLJ0BXFm20dcg645N271XgHjXcOWqTKiHhrs06
dUmQPScQlY5vLROj9+gCc6WPGNj5w8cx88U+5T+CXN7SCSx+NoPWY3TYm8uq
sVRWTbsanw/jjsltURAo5NM4uK9PLi3hCXCvsNb/uvshSin9LdWyT1BZXtax
xgSrBrNa/KRzJDgjgRD0yku2Q93YpJoYdAHVIVT1XYKG901vUv+QoXSD6358
7O/d7wwTjLer4P2TbeKSIzC/Q+xFF27ORrKmHShnouXIgrrrUB+s4DfgnT8a
9Q8JTw3uBItjmK9muRptwpO9+FSxTGFC1GRSyt5Nf5eYyxMrGXQmy+OacdHj
cbFS7GfHBt09GR1Cr4GAtk0Wv39mdiL89ypBRPBp6NUz7J451X+GUPKbUxZS
nbQ4Xdo7KbuoVYnsmkDlNwC7EVPiI5iDPS893lnstou3ja0DJQRSH+/QYFyf
ZvhHlAswsvKRnzBEgJstVxrDEujRPP1G4on5y2uZg/Vk4eGW6wNw+45/nZLZ
Hhxm8E7zBe6APYfAiokbLpbGlcfoAFhMnZduf4CTg1VugtFgsUgnoXjIg32Y
DXU8geSY11r/0ZC89PzYoia67J2wSjJJUcvvMfYQaRvBTOWC1E2d7HMZq3NX
U/HMyKz/i4uKHQj1o03j1bLb1SV5bXh0OsrLOl+zkeimSCOFWqpD739Z7th0
RNRsRV8u8JXyqvCB2p5hx0VruFTTpDF1tt8tZod0faMFDCC9kPu4215ZSXzL
osvZ130CKCVhq8Ktr5w3QSN0Bu7pt7wAmGgUJ2nGH6gZ1nP2T4sh1Feccusg
Um8pTNqk9AQq5NSwF4KIc7sMSF/AAx7LY4ZSasgKhFeQq46+ZdDRti2Xg7XG
8JT5mPWxXJXpBV9B8zi8CSZChxJqbut4yGl4/vpKU86H04tVyeSVWIA7xpZO
3BJ3tLBcGCJccmsPbmMtVms98lokVxaLwIwUMT+fenVofzrBBWxRrLavaUiu
32+0I4Y3tmf6lqFolCjzWjAvE2Anz7Zvw2WzkHKFO2TpSvzPInRU+uWRthXM
74sQ4W346rpD8qH8uxztAFU5AdslMnmxCA4TYgRDRq6H6gpQUdIBOAa/O0ao
z7S+luE2zzqPSUmO0Rh9KJMrbZ7yXno1wyJEe/mbEG6EYU6ykWi9YHc9DyCr
TiWkwFOwcJM44eZshQ3/51vBRu2agd/wQsI22DQ+GKwUKOvLthBwA33uBa/B
r6mZSYWn6rWRypneZCayCjsJ70CdhDofVtDQWKXTG7OZryHxnekTEemMOCeC
pHni8u+2M7DyROh4CNsIdoBrZ9FI28y4z6v+oQOz4ffr7BH+aKB122Z2eG3n
dRYp0RAd74A/OKD7uS114Vpz0wIkZkRFMUBXa74KDYfkpuT9QIz2qDbBlk9T
/jqOzcTRGts8IOAvahVj+3CefY+MVtDo8dGP+uXGeAttUy8uE4YK+nNg9x13
wyRPM7k8MQzXrq3/q5KfRyXMTiKdPGXy0NgokNaDFa3s6yng6D8gkMF1hHRQ
by3JZuKQag+HmoXsG6D0fcaxxkdiEsY01qKXkiGkyn4D6gRJr95yt5oZMUAE
l24Z7g7/3/MaUPp8AtD/NnXMrmgo07ybcR4oOMCoOvRboG29rsDGHLSQzHcQ
PF8PYRElxLaHDCgCbMuyjgGydS7d2pJm1tKihUALvtWOzTwfvnYujg9/v1aH
/pLY8oum5bYTyiayMRdhNY/WVkPJB4zFIvSW9B01Qf5GWtygNW7wwjKEsx+o
IjEU/BkDeh2Xpz+644FN24vKaYKY75CMvsZfZbeGo/LqgT7wW8qKorlq+C58
LERFnWOX8LrJr5EUIScg+tfY0BbTv/KsScFSPk+t/Hi0FAtzYOolcYQ//Gri
NX5b06Lv7bJ2ZfkIWBiPqtNckiALgSI/wnNhQuRRg3nKCeVA0S+cMHCrNydB
lWzC+ts+juBzLbC9ni0Zo4TY5LPDQI1SzhNERM9DPu8Cvtelj4MbqpRJe2Nk
LgMECargNo2Zdktr1vvtOSJeVMLqmMgNQMAiiy61U7xN5tdsoqWUXS3hPvyk
2qsvP94/+3PSPE70+JBMzG0jKfmWQSVKQieOS2uC/hurO/paYFfmu3zDSy10
yXaZmnq/CIy38bGJZwC2YWETn+fFBQQvhVoeqYFMShPiJN1RH7IIq1hoJ5Xy
Pd/O7vG/cwvjyjwCEa3tmN4iXYx0/UtVLZW2doEXqqAldrNy6BsxamPAG5Hi
PvRA8z7pfccdWuwqJb7JDCkBEHjkVoxzuUpABNL3+RE2VHLxtqQ70AD/FUkv
PPIBeUgf2JiKKRGVV21QEe7oTXrVVwGXr/11Rbp4+iI9SRFreXQn56iYpSwV
sQy/SRrkOPjfGXD8P2Wwkvi+OFGhx4IrtT+29qSqcrfv/m8o8sNIy7LWTZ0D
KpuQDbuy6AJay/4CHK/jrJQiejYLBv4ZxeTgb+XxZoI5OErhOEGtQVcAyW79
AJnC6C3JVFeFw1vIUR5QaQN+1JcGvP8g2bfhohAB84werzpJvD6K6AHLpT6P
co7j3jWJKx+0CQuV9/Y1VeGsuH4LgISnaY6+S9SnBYnJk3QZgxNpjGcCvDTx
KQq1LCgv5eTYjBAaefVE1sMTHK2qUYlze1+pr1M2nEQwbuzih7h2wIt6lJyg
pY4pbidBjbiHXQKxVGIgQhOC6tdMzvFifl1AcbIbQA45gnm78ziAQBHk0OWT
IDCRMHGw4I6gWg8KzaKlOnuDHvd90ocTdDQMRWzby3669/5/d4hHcl2T8VgY
pJ+NqJmccH2ifKox38ET4LAnHiuh6Qdo+7XvNqBG6t2wzOA09GWnlRJjvCc5
qMV2HEBxYHgltwxRbJrn75+UhSbmbPxVH0CAr/CVNWMOl5cF7JmcWmY53mRv
+29Hq1W0gsBwFntlnZWcqavrFOwRQjE2hCbWI/ExT0ouGNuCJ4rzK3sI5Rpj
BMTgmVph2bltFX8hPV9uHICs2aA8myuiFHQoDfZEJ4g87qgBPy0TRCeYXtWg
eDkmaz95dEh+yJyYdAYOmlutCLDlMk2tha0wzrUO13kFjm0nCpsmAShJoP7s
oCvXcZefKwlwZWVVRlFWa0SjWmTONLGRbNByRLYvArbx25IvTfs3OppzvNsS
Ujl9moeqfhiJ3iSUuedyw92Cq1r3ZfHyqZU+97MzKsCPZYplfuVf9WjhqrzQ
Oy8LPmdcPkzmRul8vqzNOwJa17VW+YuWcXn3S6icrPij/TiRHjKkNGKiJqHV
QURNsET39onStEmRjZrpiz4TXlWwGlqdNtsNwFU/zs056qXbp/Eg6IdGw2nt
l6vl4KJm9HtmPCPpXkja6A3s94+41VnXL8sJjER30GBZ3txTagUnUeHPNtR5
laCLkAlNNiVU3bKiwHyLHUFSNgVkq93gdkSoZpsBN1B/wydqIvVhip+aD0jj
pr/1qCQbTNVFGceqD/vgAYeaxCUOwtutDI5KGNEUWVQNJAoW5dh1oZZ2QvkC
I/glkYtEfEZDo3U2S89mw8Y1U8Bwwpk/nKBI16L9F5JmwidtbIWR50H1BvSG
sbp97Y9q5YVI2eznrFlhw+FzyiGRVrz9GLryldj0Fcvu8my4cXlA310Sm511
njDcsX72TLIs/G5Sc4GXztzGq1P0Iq8sgER5TJ1mIjEeya9pg8uFl4lRt/J6
SulfWt6NyG6/RsThsWzUOwZ+b1zgwXF0bwC3xFJEIP1qyygmsoorzLaAauoF
BR5zV3ARdIjTVaJ0gYZznYpy/4zaV8WjDEnvOD4bJhYk6DVxfFXyaZKwoKg8
3xXBsV4RbaOAany8rJccdOHK+UTYE5iZetyon6GW3nzrVw9neVgUuAkPsBIB
5aO3lN570rg1+gJwaUFUfJ+XShVx/7LKY/eulIVUgm27rCBT9zkSBcJQQJ6B
2Ic2BfKOTKTuUYiT6b6hus8WoPWv4JaZUlXMx7ywQdEOEUZFa31p1kx1uyFl
Qes3LGiXSLu3O7UHLitqWxff8uOAD91QnbVxJWd+7Yyi1n4ezcG9aoR9Npbn
ohdGIMZxiMjZvZ84pbbshBld3kXqhkUlnk85m/bt8h96by+0KsUxqfl+KxIe
FrWaQUZEsCle1dTM6Zs7//ruitN6fL9lNK1KHtX/Oa/aBwswRVlXZdMB1Wqu
V1IAQY6VEqpe/zKWBRLjK/ovtgCkjEFL1+TC+LKw5XpaHOFsnb8GdIxxtk9P
hrtR0C6g4P5PCeHhyYR2PmlDKTSty8abj47bZVypX222UQHMBcFbD6UBsL9e
lHVLMI/mtlS6kzgImf/vamlBHobeXV5+dyQA/4CIoo2ZI9Cb98Z1NQ8Dde4A
96wffj1ea4GDUtenXSZHA+GRxaAOzCnumpCZ9dSXHUWXCsSIg9fmT4MmT4dN
aVlm3zHZc3J+PqlYEoiAho2uy94t2CFjGBmiYpk8Zn8xQUvf2DnUsWceZUpd
6gRW/lpZfJFEh6o129toUJqIJSbo/5oVzy8abT1jKpO2sr8rlZvKXIRejE5z
4CNCrwK0Em80Sqrc1oLd6XVJ+VuKKgg+9O98KCtcuaYCEsPqYqgjX36NPxBR
kN6M7+n3zQdBj/j6dsSLUJ+kjiaI28zlUEZXWIMwI0gtbn/VF+zLfHPJIpZC
uk19NmI/55Iz0UQ61s0ZBB9dArDXnm+J4eiuhS3paq4Dx7lB03oBgwJigR3C
ZCGy2+x6IKA10Mtoz7Y5pVzo39lJwGlhvN+ju+oIJVpMvcdjms0S66Sou/kG
+F2lLars0EjjArgEBbolhMbyEJvBq3pcfrOnTuxi/C+SyIAWM2RYMVjpQxch
V7sw1MqmOAqP/L+t6E+xCutJzoqzu6Wv/1S8p47/wCLexPjja9o3IJNK6n4Z
iZWoJc6bVZrVhMYZ8IWymm5VrkZ3f4ViFH1rxj7WhbzYhB//a+GK9T5xFaRH
YC8rAvwZpKOeX9Av1AbVLri7tntwFyeZpy5qrCI9pWOHqz2K/W5sUWaFt+B5
xQE6keUNR4F5XsTunGHqa+z64Mq6b+jtPQarADp1vzWDuy4gggL9LlQedz4T
hkRkhB1zb1DNUrZjX5Q/LNxtAWco8ELloSsTB9rZ1ticxn2+jpUnH3o12e10
Q7G5GUdt61h1av6zfmtTcAZBaYgpp9kXvAiktv8JD4H6dIhmnTnMk8AUa4I6
TxlTTYD9vF9cPQHxFc3kRdCUGpJsIkuQeNAr7LzdcpCrhxFN8h+fVAqCBnEQ
7qMN1LmQNcOX47OJYgMI3Fzvi3W1Kmn/3j5tsJOQ9sV/GONPWkkfox5TP7w5
61zWSJH3eQOohL9zxDSpZbCm5mYfFxouwclqq8L6co+yF9zpYZNohIJayibY
DXU+E74qv7CLegtMO9JcySI9LWo+K+Egj57vZQWD9b2Qs5LkFdvHE+RIJBFl
sCKkYIz6+UBWyqcoMdhDRS43lF/m3p8hYcOvJyrFgVIiyji6E1TikkGA9ZvV
QVvwHY525UIdm56YjVe0rBuEQqSKyt/XBSz9wtL0Ie2kDssj+zI8xaBUEYnA
McSpAuNBPZC75ns2x+oqtZUtarNxh3gbX9xlxt/Zb1w8tSK4qsq7ULWQwzDo
HNS/esFyl7tqzJ/4iIUezkdGogHIB7YucJz9lHfBC59nuhjrIF9LoCBAvgvf
WXI8xb9DjRZi3XqfgdmVLE6z6FTCFyHJOIaeCiyPuV2UBaAYb6Mg4GWPawnC
/iaBddQtBb80x36GZBOSlSGWg6BD0k0VtJPnojbgdHZ5j3Q2GAenxjoEInGM
pgtszjLmys5Zi9qfZSIYJxQFYvakerS/yluCsJ3K+PC44JTLiRpNg8NBFozZ
g0KKPvAb4VEsvseyHS7PEcjD3SLwk74rfAkLBpFKSrytaYpEtWldWL9KJz/B
NUOPzO1snz/7xtehqSxwpdsdJOjHfWo94jGQSQV8B5qLjU+tCu2yhhPZofuG
VPf4TmOiJlIenqHR4N8oUFo2Y2Kmi2vMLWXlVHZ3D7j71uwtkxkn18fM0fy8
N2lrsyfqFthJnyxxN3NF7YpwuaZguQTMdzgVrxEqHfIHxwzbRg5156QAc9S1
/D4RYG5snQUV7vGIhqDIKZFGktpnf8LzLVo19Sh4W3Hk/+jMvZYkvdIYQ5+3
fLSTtEZ+4zL+n4k3GOjsmpsKpQtGxdcjzpQJ5lGqLD7h36xUcR/g3ByfuhM/
YMxKVz5VAldcvT6yxKB2sIHWpZCXkgyak+M78UwtsqW8c63mwgCZS/UR0fuX
hhGxS6Wd+BDBPsP+7B3OK0LnZAiUxNCiF6zqNlMO7O66mG5ZYH6Yq4c0RIOH
uaF0Q9ZoFkRZh6C5hEHP5olhEHNZVrlgPEGtWkC/XgESZ4LavZnc5raePbic
d5hyjW4K2M+3EXY/cW2cKwdmihErpGBkuShcr35ONliv4In4CD+FIPvXZlWK
+Lj6jnkJS1821m/F1hyMs2sG+2zzYRW295VhsE3RTaZtJqpz3kbg3+BbJsJ4
ic4y09R+sJBlwsXH/KXi/4ydDR0Y6AzZ0QV4fX8GxEzoiwDm1W5wgI1BD2MX
jwb6EDf8I8vXL4f04rK5mz1OCMOrbSgLG2tvWQMQnpKqWmMM02ZKbdhd1w0p
/KjiJ3Fxt5q5tP6ltZ17dNmbQc6oo+y6lmfKg/GI7Mn1+OvyB21aE9HNg9Xo
wrKW8ncIuaaip2wts1jcPEw59/c4kbC7/KKulHSExm0cxQ4mQOHEtuZZthG+
G3gxKt7yDkd7r2xe/+2EfzeyjQuARRb5EBpiuypAihX+fcrG/Vf4P9ExR86x
5JAc1Ci9l95Vo5xiJJ67SUHYffDBqAutYlrVC2HA8wOLVIKt103jaCZJ8TXg
QiF5bKp7sbo6uGLqMej4Dl75THlFaallphoHryozdBjGFJwhd5y9LBhpvzCQ
60PcWnFZGy04nKQ6QnODO74FiFF6OePEIXVenPE8EIYBJQiufWXygDj3GZQ/
lPCVXVVcuVvrV9Ofy5PRUKyMpdqnnu79Lu/UoO1VaT6RV75ja2yTVCMmGMwm
vNutLe0KHdcDkLCIz7CzHBiWNEt3WGdWPeY9NA/aTqffIrvTzBAuqv7+94Qy
WmxApGxZz+UWkZ9UxG9rETHe3EwI6yKaZ2zn7Wln61pgskk2J3oyqe5eBuCQ
daFnEzbKJuJz0eMMm2j12lCDdfYrHvcxyeXHaeJjuzrwSeYEtKFN11XkWuFX
3Qm9MOGk2ZTGgLuXP03N/DA8ZSoPCMrWwIJR5fp2W3V5sHzHxW7NPvm7xZhC
ZaYzpJfMpYD70LBgErD7Px079L/LsUD6SLIXB3YE1MkL01XsLwsKOlp3Floy
sD5fnxTeviU+4C/zfra3MdvRPjLty95YPpijmk1u31WK5VWZ+rXJMq6EZuvr
iLZUr/JokZT7vse6uGdpoNt2DlQQIcAmYwrWEIFkANH0WX+OiFhhNnBUnqmK
pEOhYm+J5VLrlLCd9ToYs3rkkX83BCmjwHwuo0nwz74elql6lZS8wK/+Rvyl
bkwp3qvEaGIDBT2sV2PKXfLds2+n0NLVfP5d/9oRIh7zH3Xbbn03PRcmGLl6
skKWcEtXUR8z1TgKk+T3vpUhLZ4OI6FkZE8IB+zl3gb64Jq2iEMdEtlAinBk
PWjkCWbp9HgEf4bTbejfCgIxfXhOryvEF8hibHnUOeR1jzHfos6FfzpPVQUQ
BoxGFfzTESntAv7eVijFYx3PClW1Iej57GtkTP8vcvHK83rZEI1RUQByiFFl
N2Afy/L/Hose/h8Aqpb5699Yr+DjrG49OKi570++W98HXLzzvcCyE9HsiZ9M
iyJZW96iJAalfFlJx2ZtIbKc7e0hPe5C2y5YTyzQhQTg2eQG/wR6Ym4/Qy35
AxY+H+jxChT6Bx1UF1Lr+zzWaqKT5d+0PCa4Q0Kr47npMHe3Z5fHE8hAD8I5
YJ3fKyhSk7xEnIO/WDc2LmpvMZPCU0B41OmX+y7do+8vU6NnMBog2fhGEl93
E150OkB+0gaDgfy1l6ZDMvt0qBVhMWX2FPIXuDUEo5eDUu9DPd61VkLZwrUN
W12v4psJ9ml4q7G0+Eg4TXXsUBKA8tAt/Wvokkk0/Sh1gf7ip6KOFBWMAg2p
GikPKxNoqlgAgNAun7o145Xiy79iboWmfITa2/2bd5lUVKdPy1WZo8oE0+NI
/8ujNEsUFbInUs0Iv3ZiWxbsKFBcuF945PCQBgbiwHokDPjARN2KjiLfDo9r
wqijPPQeHfvbHeUmqv0R7ZXChDP9U8aR4TdMnVe0g9iC2xoZL6L6xwVF5BQQ
/Vm7gXbJjb77DxkVqlpilfV7/x1y/Q0hcUFEf9wfUDGTOFkJ7IJmHcRVDjnJ
4sNUN+D0ZjqhAh23szHrQffcyaukz/2QJWehjmR+eW4zNjlGbwh5pFE1aqnA
KDK/dIEJtldPyXi1QWXcYyERmL2/K2Vn+dz94gRVt2Wpzt+uAllhzC2ocRWa
6dYZ9wsO6wTYX6JspsdK8y0j7edIOssIZVyaM8+zaD+z0Gdz7BG1d7f1vSaM
9Uimukh8wJkquK2niLycMs5rR9Kf919dgAO9TAZtjlMQK5V8NeDS6IC6Rgu+
2oFomm0d224d5zWmIFvnC4zrFH1hhfW2lZvxqOan9b9x7HFGdaFfQ19DdFHH
ENsHJ7nbw4FYGnr2u/ocVtwjI9GBcvD+dvCDyUDYFICMrftbi8MovuKJBrmS
ZZN6uOW01OQsYmyJ0lmSh++JbbuH2iYcjaMntbFz/lYm8XfD0sgUo563TS15
km7WeWClFNR23EagWx3/OsQivtBidqG3lESkPpHSn7qu/6IoEdmsYfVgOzyA
l2I0fIYzXTCTo/fr2ytjxDIc6ltql6/2LbXdZW/vBZrl1toM2h0cIP8AAxfV
oRMMsO5q0JsnTv3XYCc/LqSYxyLd48wdcJ0dwOBWZ6ErG3aNZHpfQOZ18SWh
2qIf4VP2Kctga25oCyuZehciGdT8VnSDXaD5alVMtvLz6R2X4poOoCNqeEMp
dFi8Er1w739O4IW99mGgI1/veKIpl3jnhCFlrkDnMeiqaz2SmuW80tN6yCmO
pFyyd7IzvmLob7SLuTubFVoB0eGULDdH2faVTMGSzgT1DOjUu9EQB+SXUXdd
6PKLDGwq/FxUV8M68+mZ/h3o8fouYYBaQPcUnxfMZrOZtPBpxVIez9Ne9Z9S
d5O4bVEWBisWZhXCHG6i8ObFZILkE7XYSGrIvqUHnkr7CPYl0UTItsg7kc5J
MMC6Ov8tBq602t/GZVOVhsefNmIhuOe8wc5U+Rs8L8Yu09eRH8bEqvPEYPSe
9m7fMQrw5US6WjmWyb6k0RfyraABw6KzzVEN/SEFuUlRJ0RP7WtSGzWX5wcO
Ew8dEHzf4EzPKv+2HT5uJ2Wvu0eLJroVqUZiSVnI1ju4i5q6kPPJTbfy5o+t
rk95fxhV7my9/Ca4DUha2zoyD5U5LGYfpvcCimYBLIouvHMqVZuYBCwBaeLx
tzP09E1LkUvHm93fBVKAlCH4y5Ffo4pbcB8//uNMvVcUCD+19EBGtK3bS5YO
85IVsfGh/9X0mOSlbGp1XUI2BLObh/NNE/aXfVZ03iJ3vAAEWr2JUvNnGiSp
Rl7baDcCw/xioQCeR9kCNQxRwCgEb7fMWPcEHzj1lcm8NUF7PoTs7Z7umoi/
Ze0KYYYp50fsrNxLk4mTu0kUgRr4JY8WdxBHndPrNpVwR47ztD+PLj4IMpnb
Dx92XzC87PBK5bDCuP+VHohWhD4cXcg6oCtcI/gQdVLgccUkn3T0mv/29IUq
sm1+3IPIF4dpQBh0C1GEGWu07Cbhd9mtlcgRv2HruJwf3NJipZ0mZ7t6kSiD
lq99X7fo3GeZhMKy18Z3dqX4V/vKQa/TxxXhqJ7o7W6aFBdwJmYlgKQFxmKH
7z+Kf8wBbE8xbaOqnZITqe0K4YawFJkRIdDZdXfbZZ8mmdGp/ZIgtwXaXTGj
mx8AHOXkcGfIVGgkDPcIyTvvBxlsRxtH0KXR1sAHDFJSvdmbsS5lqN3t35DW
QezeBH/Y6N2+nvR2H4AKcS8Z5HIkbw0y3H/i0kR97Xv/Ymj57JDACsNiuu8w
0K1ryhd36Wtu1ztTWT9nqlqLTwzDac+oTqrE3dX93aMzOnEbivwrjlSa92yq
1wsMzTwsVkq+ZlANUAAA6najeY+HWVsszyhB29tiRly8MLcjRkocm+CiwadX
ndXQJBY2YSCRnyQyJtSvUF+UiQwj1jn7K3mO+1dqHMjWR6rDHwsPFL1gqAv0
wKz0JJW6AbQ1BfU7GdF7gZ1y0jr2WvfNhsdakPsyxVdVj2jM5g/gsHVd59R5
h0cLWnXnwbIzHgnErVSLRPcrqprz6oWgi5o7dNHufoFNYNPavTfqxKJk45pl
ydjR1zRRY0Hml3e8CvYJfqRAv/WrKLxltGHpUlfWc14+pFuNgFpZjhKBpxIS
C184fQ0SNw8buzhle0/QBru1W8538AuU92B6rEkfx+tY+FD0Z7Snp0xj/3B1
/vrjTyWqa2C06crw8iw/9QJ1wl0pkgkKwsWSsvgLnRf9T7I9Oor3bMZEwHzi
T48erQHeqr4e4tZ3PyvipEmFckvbs1V7ewH80/H/1pOIpPH+Set9E4tEhNHf
zlPCWxv01ncisVgzw6bdgfdKv7Ndo60sNhQJfJN+Cu33+OoD89f8j4cXQ5A0
xS1y3TkMAzJtaE1qCJPfW8ngyXfGs8fmIFzQlOLhiya+35DZ+/RQhgbyE5tR
zuPTe+qSVHT/Jbkg1+2Hbxd1MwoOnVSGfMl4CqGHij02wxUOk/DvWZSD4N4u
sP3nVQs6M5f9VDN/SH1668gcp2q1mjxb6rx6q6Gi51uT+zeYnURBLwXNxARK
01S32LlIDkajXLhv/wnUu5JWj9hBSYEQdetNU4eYvEM+jDZQ8iEyRbbc/zns
Y7sOTa+6A44sGo+B9Z67ampuN1JcBqRWOgmy93przWh/MEMRYICFkb1sb2wr
lZsjlRyczoTS6NkF+n5zLsI8m/339CqYOO1fkglslprpV5fSrDPVgm3J/dyY
YGfScQmLQaNnVBQce6ychXywomq3U0gSvxEaKU0gaLOC+Q/b/zyKf/RrViQ6
yU5GEgul9Z3PYBx+HxrJKaJwCugOC7DdBsn9/z8D43aImurAftH2EahDx3dn
us5rxtI1Q2ionuq7gxwHSI09gH9oNPg+VLKcfNFbL1keakjDBzdiLn+LYmMK
23WDPQN56P1kVWSzrCOqFhEuSBTMHr4Cg4g5oT89mDH/aA91DdaUnePQtbAE
1jIZozhVs1sUk20Cv2lyO1WqGi7TVVoMAgD5NdIRZwzJ/G4bWqV2tiewapL6
y3zIkt5ALn9Bxu6iABmjxpOVaMyCpnu7rKqEk2+KQ0kcEq46gyIGb8W/q5LD
wG2Os0P7KKT15lHfxBIsflZwTnO1YXhigo+KQWNBb72ognmKV3XHPjpoGwVQ
fXVZeJTwzgXcNumFG3Mxh0BDgrbvGbqLHHKNygD1RkGLnYki+/PFcZcUGRaF
hLG1fKwmz1ojqfmm5BxRfW3jEpcbzP6wBfYbk567F0eVhG1wakSIZ1hd2BA7
JesI4CTA2h8SLPTHXSg0jnrabdiicHzYUrN2ALQmcWNNQ7Jd58TAocrlayxs
LehVHBnGoo1yxvKWhk8V7kXE7hZsEYVuiti+wo2lx0nlQ7GkCGnVKSVJ9Pgp
CMXy70JUS9VwSiT314ZC488AVzH5CTL2kq49MXuUHGehKpti3B37/0xpCOg4
DiQ+rCSYfXumrl43P67gj3BdkvxX4bCq/WOBXl89SkgpVjGwIdMMlwL/n+/C
Cl3DU+Ftk4oc5jd7qFR1FZ1oO0EjSa+swKRL9aUZdMix19jZJ8OfwZlOgEOl
EzlIbtavyJNcA91YlcARiuKlhhiquMlKQpZNitwG/jBOMhObfIIKHFunANIh
HnhmJu9cX8t6kGdKNiJISaSl+YADLzBVA6PAjF1ZJ+y1aNeNHTHzJsUvDKrp
lEhGK36cdWcROviIbjhnhOE0vaakfKwmDigzpc4r0se+2eqT7NBzRnecOEMF
xxQYeIeJFaBAXGODS+MIqotF1OzGcAkYJcESSz4twBGKQcU/wvt24yNlqS0u
kgn+G40R+IUY3J/YivVmPphNW3uBgr8cA+cQDugjcPG5mfBnp7TyhK9GIkAU
67lFwEeqra1YXXHpQQFOcukKo50Rt0dCKs/VUBtIrmrbD81S5N2HDmVwoK6i
nTOPCT84X7XSUlwpe6uxCLNxEN6YheyewuVellhWcA7FjgoCb1Y0RRstAhpu
EiB3BAv9SY0sq3e2aOlmu+UJ9SapmhZBzo9pva6t4eJOT1otIyNtVY3i7q2O
A+m7SzAuk9bGUAi3+m5JBqY7uholv1AfOQ0APHCc0K/QIyWQNYFGz02txX/g
n9ujrekdJhG9Uap+i8o5r/e077PhoM5GCmWoJFz2FLc7imslo4CWyOJcVyMS
H1iofYMHhH49NXIoBYvgL5dHPFMQ/J2/p/+QooGngzE1Tu/aXS3HcZlwIFgm
zcOG5vv3fpvtkw17NkYytySFWRSFwKzcPcBEfPqNJ5vTZ9wX7ildhWGdLNQE
ntd+3T2wGTwebkGxqVlioXvz6EMgvGrZafLdmX5QbUP119pD6DbU79TL4k15
DEUSkh/IuHnMMKCUgrdYZ91rYVlYgc+6mZ51CNf+RL2pLYlpVEx7klr3QeUc
83oXsA7leza4tpvClfokejNV4At2pi16Hk46VLVKDzx20n4nxTS5TVSHusmX
vEHT9QWYYgUs4kNBr0+qWFQ8WUc6l5stpUh596UydL+j4MYBxrYhPyQIC1n6
GCbvhUnFbHctAbTRN5lw9gHEkRaC1crbi2Sj+kxRDbmuU43nlTlfYO1K+ywG
4xuJGyGy/vFfksAwN20qDZgLchmhWQfTA7DDwUc7HykhVlrWDkJ8MR2H5SE1
G9MpI10L6j+mwDgPW3LLDDOnkm6pP6yvELPoRwp3EqXPr6kif3hlkyAdkHRD
8E9GWy35DJOnSyI7t6MvEBA02zp/UivNEXYSqxk/5DUwwMXOI/6QTy4IRaP/
Snxno474kjoDBs0Q0XUcrMHJSI+VprAXisRZ2Vuin+yshjXaml8T7+wKaaJd
VCiDcm6fup0yfwlePbgEncJpp3u9BDUIuKRD+mrf97VS3VMexMoT1/HunS36
/HW2ewd+88lux6t+h/MmMRxVFhctIghFJaqcnf6EUD8XgEXMuysjJPJdHveJ
/lvWORpmBsXwnhe2ONC7KsakIyeWnJ+EoqlaT2oxQZ/ms041q84w1mXTlRiF
MIF0BIQQL7SkKvw96BbsZHoyVqTePcZYxquk5MbqWX+xxn1oz0m8fCs2tLh7
wEHMS1bAgW3WY85P5N5np8ynetB0wjp2H6VCFbxriMeFpuGLqLjBngPqMYj7
E6q2Tou+1JLtOFdtMwHabGNYQ/N0ESi90nQOhBqaQJ59/QocW/obQy+5icDO
S0Ikwyz/lkRaWRJ8V034wW33QQmTDMJ7EpraScBnws9obMXmVZrRc0/EScyq
wASxjQKtfPRV68Ru+ac2vahZjHrYa2HLtgcOcDLPvQlukaeuQD1JfI/kbydW
puJBnNXAxeUuuHMxNhXAqT05RSYj1ckiZBnIOBVLXIkciPQR3W0sC4+WQhsc
8qyI7StAME0/4tAV5CQuUZhKW4HIjHhp4jfNgxaSPMeUHcyYC5BdGqeVDmBs
hy/xNnDsVo1F46pi0nWHJEmWclihUFuVZJsKYl8fqUC3EktjnebRfLBiwEdx
E1hC8D85f5WSk7IKmVI51KxeMpMWrctVUxASYpBBKfDwM34SU/wJokv7z/vy
hhFMN4DjTFx1Nucrr407A5DpQ0T4f/ATMmPsYqIjXHO+QJYXXWtiBrt6vEt2
78yIEKHykt3cyW/JJo3ohHW7i03bHo976La4eWNZcEJKIwZxBYEALCVr2UhG
djsIjan38xa3pqJYIE4c62zVfJAeXvs+IpxV57jw9zQ0FbCyNzrnLF/SmJvf
LFr44fkXLk55CRFPLbhWmXWxaXi0SOjeylYqp4U2jJhrUpF21yH2I8gsp2Ms
wrwHbrgNkLRYPX547fwdheMO91fkhaoVAUAozGPmVyjvMnim4J3rdjhTZHZ4
KtoN5QR7Si5gPfyRZeW7NJq8T3nB4FrALNEwa3BZVXUFyqNKyZ63ReVFwRdw
MGwyRplkhkBLXiFNLr1InS+7bNQ31iZyJOV9Um9MSe8eP2fdTlSMnR9IObTK
r5oMQveU3euqGayX0sX6QWiBNz0wyY21280mdZTr0ZjoBDPH88dQ1BWr4EP+
+DbdqHs+AGT6Pj5X2i7v7LNCx5pMNzLzapgCuvrXuJbwgMt5f8acSc9uoku5
3og+nq9TG9zfvUOzIx+md0UG8Z06QnhKAp0UTeFza3Yd6E43d1SkU7umCd/l
PpLXxItfLz8R4UHCONtBFm6gVgIR7DT2cGvyoYL/nGcecV+CjSo//83JVpSV
Fn5InfD0KD2iYnjSYAil3ZucXsXH0KE2sPFR7Qbi4/v8UF1JCZmERFnSOC12
KCAtN3gxziBS0s1eewwmNOmuTzCpnje9s8W6qZRpqKnntWT5BR+ptxBpcNiQ
vr1znim897Rdl6aQGx1zOBIUEBN1SLZYdK4XxQIggu9uKNShlYQ8KaImKI3E
/VeFGgvXk43kk619fnXdgLzo1ZETJ3KgMaotVFH+RLNw1H++HvrjzGF/oLyN
sMzBuVL7JuQ4bIkIq3TeH/oQJOGQ60XqdOcUsZURgix8LuhcUdo9BjN5vTAz
L/QOVkttKeitAWeghwIyF/fstziXge8NY3kN3fVcP9cC0lNNcZOhBDMbeljG
mx5D50b1dg1j4oyUqC1OY9LzfjzVA8yEXHunNjvLYULmZTpHgUCoUKpkRGNM
0DPz7buCCNsFSblmq8OHM5gkJad/FaVW2Zi7rCrts/kdVOocDygpAwK/NUgZ
xpYMc352nIpUJjeImHHeM/z1ie2Qra7VRiLx8Fzxsl9CfqyCdIRNywkLzxHq
GR+wIk55elgF8oz/HtLWuCc3+i8M+pPXQ257P9SPhj1Cqkyy4eJTSKQeonxx
4pOJ2Kr8zLW7mlmlES/5baCx3/Bs9i6l4E7TLmr3RJKaKv/94uKwWAXqzYuT
TlGAjtiXLhb1xs3ii+h0DSLX0c5oRxgs7sJsC2ImO8xgbFISZvq0aI7v+QF9
0ztvI4fIFadq9aRezg3zHwMABapJnHyTzyq8hA61XtasO/vd2VwFwNj5CL2Q
yxl32SVkXQMjOpjReoMhPg5lumB2OhPpfVIMZRfpAqNt1IoNhziUVnrONu9O
MA+HwBYjOQS/R7TBZsSJL3SV2zPGQAXALvl11aA9boRZWf4fqnLMzLQxNbfK
PCSVLd1Lsss5q8Ijq6mSoNaf2E8WhEFkxbv3T9vBYyY3jUA5iRmIShpTt4QC
sIjw9tTMx9Qv39Z7YOEfYHrwTE4B9MfnJfpTWvX+ZaA76q5DeRu+jN/2g8t/
qjAC9FQ3Jv9RjwQapTq9qy09/WuBTft67AaaR9xG66Z85xgJVvVG8AVJJMKO
luPWstT3YnaESaKV00acGHbZ4r1ASuUMrJcaocY7jF7O3aPKbL5LS2/SEgGh
4EI55rGV3G+OAogGFcqaaRuIawnyru3uFWgpZWfqbEgo1KHWvGdIAEAjViW2
7diT7+xTgoQcHxYtZAIfDXr2HwfMfRPnCoqwDrItRnJgBFu5b/xWM5/lK2nK
0Nb5hugdgSGPQ9CXGCoohg91KX0uUxStrmYLYsqg3C0Ma+Jj4BWh0AiAgCca
otmrFsAIhu0r4nxAY0QjPDyWy32a84Mu+QHu/zZ+hAAg9QTbTJu0PGdpa1Vm
JlRg2hKMe74emS9OHWpdCbbRp8s2O57zE9VqwIadWv8895tVJDk67BnJjZhh
MB/aoqeCeAmwnee9+1xD6lim2ZoYfo8zx0DjIxO53rDke6odQxfS8G+Uu5UR
clL8ycmF3AtWMJiQiCKX+k3OTJb302p3Af3jAMYVDfwnGrxwLw8rYQ6+blGE
mMXBhfJ4cz5eElFTXCsL+hOn+iHQkntZ27v0/HdyvO8mGq2JhmGJYT5vEYHh
uqBN25WS1j9vQqOu10VVAK1Kjg/sXNvMM0xUcomj4RJnc277ZqfGz3grj/4S
72jwnSm/j7VAqP3aet8PaorS0mkMsrmcRgKxQc9UiO/c09bNZfmZvt/iqwN1
rgDFwYNZqr0rnI/e2csMg1BAOGhmNVC/R38wVG62dJ4FbNdyUZHfuWfwZMnC
eDkGZYGVAirH95j39CwsTnpSjG4fpOHiPd8sj+d5vBgRa1B/HyWKE3KMGp8t
dFuaW/z/B9zBorT9qzLVrxOY0XQqQgBxxJz6FJNk2bwQRr7miBqCCmGMgyoi
YH9pJhaZDX+0gBpLz75JkI5jdFfxyvfFd1CBVAtgOOo63rjGNSGpbWt4jQYQ
XqjxE47jkh7cO6vjQoYlOHz499y7VmLIKX/QV7aIoJhQ4OCZzAIikh+8FtAP
cHu9zOvd3ew0UKj/xlD64ikh6YOgnT0eyXmQDdzmj9UfAAYcirkza934LvNd
aL4i08fjSko2Do6rvsfzdSQsFgaxpsBn/Sczdbzywxjn0xt/bRUszXvnySoh
X5HgDNLhS5MS/aqnv1uZVT3vc/wP/UG1/7TipZjgAkz9sOb/Q3/NNrcyc7WX
5RfkJmrESt+3VceiXhPh0v5/zIlrPI/K9sYM4A4spYkZn6BasGp9hZPAFogY
Tuneq4HjepugoM7Zspcom4XQII9szyN3SwpGuPnlIELRvbq3UAqw0nzyEB7X
4R4Whm304x+8F6gKqktfXn5xUgCJU3GdMZUQkjB4igz40aoFYhlEFNttK1SC
wxp7tLFTCH9aM8RansGuq3CiUJD1SQ9/T6OSMY0qTQpzMuL7MrJ216vhic80
8DiT031L8J0LRjdzi36wMKJsCgdZAV8qYBdJrcsxsmgr6erYaAGyON30GUfv
O7xXO9dFg8+/9HQHYjAQc0pYlZcVzRCm0HSlflnXS/3dckFeJ3EpYCVuqA2L
KWsYjk4OaOkplq1XUuXLKMB19eB0l06MZ9kIc1JaE8xP3b3kEuq+jBWGzVN9
H4dtCqulQOMlsGAcThspapTYJOjPKa0CGx/rcz7wTdtSO7F8r+aG3PxpHa1t
1HHs1cAgf3SZ5thFQLWEWnJFZyu7CGT5ARkqIwQp+TsCoGyCNk286KNO075v
fmG9EbBmU59Sup9FWXm0C/nj6TSS6Onks4k3WhV5aYItIy4fh2fXyh4phNTz
WMqHRYrixc5nd9sYNjN1w/JSumVHbZFYTZoRTLswIa2c+jmDhIPzjVyyOYMt
Vl/IDGytjl9W5Gi/ZxNRZo7rDO/eH5sNWsjk23mU7aqnAkKRb01mB709x6ij
tyRgFnixuCqKsNeCyOy9MznJ2J/+HmZOBe1uqMIcn8ZNkHdAlhsePsOIBuIH
pUK6lh6Cvz6b6nTiUA9k8jkZwq6bin8Vuhz05Zl0twmE14uyc615W1qytDdi
+WIMMfF2iZ8CkxuAv6IaS/c0R+9PXgO8C8VJpRGB2TvrLmz7wljyilhKAkig
fBTvgQ9tfg2TaRyCOQ467W1nm80YydX3+aS8Y9yPIBzRajHgcxKdiNuSMVJi
D3VXC2xwSPi1aOrYLDVh8VRasfaPJL7z2Gc6RB5AT3FA/0eBTVVEoVkFHo9J
VvRfZHF4a4FJGMHjOnkIb1Yi6aj4N28JI50xbvP/frKDjYaG5cfjEfR4cD1j
Y5NnQ16IcS2z0B2zCYATbbBEixRWpmLsp+n66lpcKi9aaPNzU55L1tMG95Jz
RHx2djCmDLyu+gy4VsUzAXbSHx+5RzMiVtRM2Xke3+kncMZB6maiJwAxy9lp
5LpLy1gBVjvMP3DUZOpVK+04cVtkVcuIbBeGMB3HgXZmsncE2mbyDzjF6abQ
vGEsJQsdJvhT2caQDtKI4FRkqF8VVJUpNiDJSmjpvZ43vKe7RPh1wvkLtQDa
u7tQUmYMveALdT3dfldbXqY6zj9I5qVX9KR09SxWTIqwizEMjcXdyaWdcs9z
TJQ2zvaiLtT1gZmC37BLsVGKA3H8ScKgiD+Q0tr5+4409LDyWf5lUhMOgtqX
fFYCM6InF87zc5xrN0jkoC/GUx7Jvmyk/UDHzInHy26ROqmYKXN8ubAm7+pU
zjueHG3KGOHQejeSKE6aa2+vWe5G5Fju/1Xfbt3LAx/H2WmVZy3RnWuy55SO
0ojEuwyIQps7a1qQKrXrWPZBDt2/WJMhPrUQNy5Yn4CNZw7gmj+r78VIVxEY
bDqtNZ8iCvXXiq3j6Vv24d7hzSegT9hD3gNwoCz9JMn65aK2Wo1fvMfUOqnb
uvznKwLzbDE35ITcRPuMwlkH/WflCtpb3tC9uwOeeCyBzguCWly2wolg77Dg
lxdRzxDWhwyTMdCJ7nD9eCc9rBMUmeNd7wNTJY1UMXqCImkKV+nXWfk3G+HP
7hC8YYbNw+JI266jT91MB8wLpkVGlsIYNvg0byn5hrfpGDvbCg0F6IdGST9o
Ag3MmS0lX1qQd7hBMlmNOWmtF0s+1krmvTinRX1dtIr9co8t/StB5+yhx2T2
4EojyHPMgS/tYNfaC3AS8CAB8g4hme/LSY1kLw//aeNkyhrhlErD2yXBlFtk
8ZPbxj1o7GyxJNf6t19vgiEL+2pDLu+GkyWfB5oODDrktqp05t9UDHbT4QfK
W98SRExHrhYhfAhu06z9qNDnugeShlS/WpZJGfIQX/bByet9AXN0fCDMrp/d
c+QNsx4/YkHIgUtMpFhwRh2CjLk/sfDOIl8orYP7ZOBkJbtjUmV4t2ZbMSWd
r5TJm8t8pkZKieZfhYcP/PMGIopVSunNOhLgoMXTVWsx18KXHEtVxYjDc+IG
400+nUPqThIsXuq1ej5FQrPdSND3AJT9y2dLhAzAx6g4Ubl593ZsXE+aR5HH
jZGuXt9XfVybelCXF4Tsts3a+k4URT/HFGUZuYU5C7jKz8Xh43RHZ0takRMR
NFBS5At4kufwtoysXrLIqtqNBUlBtmapF3O55uHDTN/Vulj+ZN+EfJtPwCiH
PbrpmWOU2BDFF3MJeCd3aLu6/jzeq2i6JAKDweEFEGRf3FLUxNcMLzFememH
JKo1P3TcWQKq5HZFLdYtRhAvd2WmHDgWqUdaWY2RzTyLtFPUmaORv+hDvOdG
PlHz0zrLg1BMGhaRtSWtRAe8pzZm5/fe8Bg5M1hZYqI/BCSA+euI6VHrMPs9
mXGjETg9Yg4cTD7loWTO31mrNLXS69iNXP7c9JWZBXT+xh2L/lmvAc+3D2WI
4wn7lvKTlZocrLXKUORlPhJCXOnCtaUA7i0g2v85UP5vWHe7zqACH8y0QdXg
SX96PzlYOtkq2dPIW/cZYHmZp81ssw6ZWHzLZhlBb/HurYzHL3e6CEt/YIPJ
LUKpiKOg7eLpSC+RlPe6xjoQ1T1cbxLutw6d967Hu7OcO3fYVWNJH9Yy1aWm
m6MjPYizPMgShiD5gZpiYB1tm9zZ1yjAPhiENcuthZ6tvlmkB5Paz5+3rcRW
fbBpbgt6yD9GyMY/igqbMxd1BymERrUpADnHZOCZnJatsW/YNYd0DWinzhzl
ADA/KnPHfImp3MjxcCKwkQBZHogMJLPBqZPtG6u3XigjnY3tFJmuf6bSb/jS
EVVCJ+YH0YYT6/XkrQ3cEkbDWzRUwkw7YQj2GhJzP2STMD5xdSIM57r/MX8d
j6RKpeiCsH1cbUu/M4DfRRhU1tlmKCjjMUnXeCdIx/DfViuxQU2zw/lxda8m
WokBRSjQ1tUgnUXehzIzIyA3sBjq77zLtpfyNVdyqQSvdSO5R1yvKywtwTAL
gOzHtDu026jTenFL9sK0ad9XFKpHs5a1gVB50czO0i9VW8ZV/EQ7KiJwldiK
Sq2M4SjXupPLMPebX5SCYe13FkKxqzQdgD6YDi2tJ/eWyW7rM8iJx0i0arXQ
pTcdaVgxZ5MTeqqBPUMtR4KLtxIOck+0lBNKdRzLJAd2VbAzgv70sOA9u/4W
3cK8JtTNPaXgAAl4Uwo6XOo0x0ApoEvcUvfZsWZ3Ms4y3bVJyw7UTyjCfCVd
THSgahqjwzmwgy2Nn49OP3fv1DjjPr744My2YViVh0fuIil6Et4tOG13an3F
sAN3zOsjIm59wBkmMVnzm+3zOvp1j+x+EbHR/8FDzv8FYHYM9TdtcYARAmIa
LkjVTGPUZEWuxidATYtzw9dOWLDZv6YX9pkYw4TwS5OP/YFeC+3WBUi5rXUI
XFzh/QjL8Uc4Cu3WtSug9JtslvmEsacLzqFt34evKxk221m3JEf+SmT4iZlv
6AIJ2q7HrNbw0NLd+jara1KYe1CXnyhOde6910u7Me23GlJi4u9CQd16qxDj
ssVuC5kx3lGbEFOeYTqcRRM+XtFbU9YWQLVr7XDIO55JSJFts2gXLsx1xomD
Oxl/x7WL9M7Ml0JAACiqhs+6mPH2T3jBGqxJWd7/jqGfECOk5tRS/0mp4aCS
VXLldetPCPIdhetjIzYZhk1jB0gGYsmTTK/I0Wl3iSJhDXEhTyCkEaPgx3NI
met7KGqtlDR8bRbFlsg9DZHD8aK3JQdW1KMgQMUX/q6o0Aai+cmYlUprWJxS
9Ko9VdM/MF+Q2CCVQpcX1vLMuPjlBNUDk3JryOFcnw2OtRylqMdTr/uvxH6r
ksN1AGOtGcBAWccyhcKR2Fr7CL1+km7QAGbZb0xvU7ecr4EeDPps/QwcZN6Y
M1uV2mn7FeCUV/XziZY1p+a5Z3Il4ZpDz9a8rFMAB4kydAW/mB8ML5gEabOz
Rj1LushZv2t3SFDXOFmXVqOy9hT+LEH4aija8G8XIwZ310S5BmzMPHjQmMQD
b07PQ/nGX5zN+4P/s258ARTqIY2DQM3lzH6h7rYk/IV+21iSHUv5w006KKbN
9WF+FxqJhlthJly20mbpu+qTJleAkYbWlpI5vkgoNF2RYVC+1dcMUMlM9okB
CZcJRjsVaZFFp8JeqH5GHUZ1sQEKlmFMJX8NBDSrmU8Kg5lNXsoeCjJMhXD3
VQWIbqTM8yl6F4zbKUQok4NhbwhMkY3AtScW/pfldAyROp3zX4LFSvN/EmoG
fUHOu+nmtNrvr9aNwllQIVOajO7HMazwQQDdH3CaGE6O//PH9mg2x84V/pH+
3I1j8ex5psmNuX/OQZEQ+KNBwB5uVAEcr3WSqW7uccHugP0GzLl10o0OdvbZ
XQ8DmdwryD6eInDJU+yl+ETP2A7M/cKaWiuXOEBPc6JgYTipTzasIjCTfObC
hgBb+H2WUKOdlyPa32gxJ1ZZ2tDfUhCDCNtz8LuC9aAPCpuXk1rdxZPQRfEs
PVvuqXdT/QeA0/AtMMyLiJvM0tG8rHaKhly72ZE/fZ7GIHvKnu2h7K8MI0dn
14Glp/iK3jhmEhTiGR0q2er28rEt3HC2zTlBlsXOfon/2To2Ds0XA9kR0Es4
hKYDx4OhisRfjoKkEDPGvsLL/14Tf13UjfUebf7rgwL+pPrIDmBbc1pfEL+3
3/c5h+siJRDlN7AZ6DAzqQSiCV38cKOFPJjVfAy3fZYI+pIs36kRa/UvmdIE
dcJjKnkLvstZJfFxaRP1/8/fBnZ1Doh7XwQ0E14oXNyRcPb+bYWmI2/ToMCB
5cqjjre6JE4bVetrenP/nj5oObk6qst5olHDS4164sbR2ZYd5DIASoPO7898
r50l6DcPCT6JeJi9AwlCV1YWjSav5JL5vr4gVK6+yPWOg6D0fhfjUsuOyEFQ
wQPSpQx26jhNXlEvlG6c8NJ5NPV/Xa+OWmPImOMyYj3G6lhXj45lrgLupa1h
S4Mxify57Neah7DCfyAzolBxSxK/6EwD1DimxzRspU24boH1UJvpEc0LWbV3
WrdjzfinssmlVK3Wdvc+358m6CG4VCKCWkN9yWo4FIuHg/rBRaVz6Zpx9B4O
p09281WVfZLbcViPGGP1SrN2bFKgEAGIbYdqh7a7xolpv+fK1NbrCP3IbkbG
vLrsjxBQVeSgVLnzR9UJwz/4Q/DE2EMXnajaGT98B+QH2ZW3IepvhEwW3PW7
704AmnHcG8g7ysHJ7ssowZ1WiW09uQ5K5B8s78FMRaZeev67gsbDk7yO2hDq
ty74P8fIb6ASx9QYYI1ZNXRHdwVDRmAv8bCMTWsqP4JoTRp+9UB2db0mypvB
XI9eIordehv2t26Nnwe/6BqL64DU0ty2YV4YAzGvIbEtvkLSrxy3evd8HDAz
R6PgGhRmdW/P2o9PSjGz1rxwl/QbH0FZK3ZStzieWKhgboOIyL0yvEUIvi4F
PwgkV+ppkCsl0TlbJFntTR8tL1Zvm0jNCveqxDXtoa6nANrOvkaeAFrCqWqK
SwRaEWcC20K+lAV6jEOEAFhJTeDw/bNfFhAh3FEzrUGnGbZNw5wdE8pjzDXa
YW+DcvOtEES8lu+TC62g/bfqoPmqp/y87K/00DgTZtviBHf6Ww3LPHTr/UgF
FWr6T2FNcEfpEOmWiAFtLtc4Df2UW2iqgSx2KfTOldun5a4nZI6Xq9oGWY1V
sl+cpNTeBkr5S/blcD1iDOhHnctUUcBO9U79KxA3DzEL5Tb/r4DfldhxSNEr
eEKO6/uRwDk908fJkxEigMNGsredttFApdVZM8iPha2mpOWN1h9X6qjPwTK+
q7t/uYv6U6ApEK1DJLk3yJ3mOMbiX/3UYz/gURprfkj4HbUfEGb4Mc3a5kR+
th++YHoPzgTG7DIbPWB5IA+SI015zpWRo+mFWsYJZmmZnSENfBLRbLhVJnGg
bl0KQ5OvMVjPcfjefwXUGdOptCxEhOBBuW8BouqurORG2p1fiFfNExytXHWQ
yL41KXiuvQ5+spMApWfBtcP5MtvD4xoYJ45lx4lTftoOYcpGu9BVa0q/gB+Y
FykvQYqlUU5Z63PRBvf4FNnHgi3dB3iUwgQ7XvroO4wi6qj/jOGksjvi0y8T
B7EHH/18ZIl5VAKAz7zptoZ6PdU8RWGi+DRNPEXg1nDjzquQ59cgSRV6ZDnU
6b6iUFxEAhOnqHEXz3nFAvXy+u02ujQZByik2ECRWC5x1r+LHV4mc8KimD1S
eSD5LVsEuEzhzAxjUvRfTitKH2WuE0SLZRcKbBa0ZA0n6lDxXMkJhqh1RhGp
Fk+e8cxCFDgokg9TKk/PFraWSsNkyGzcXxsoyRsMUjTyqXxkhVt1HOpfo82A
tHURRVpjPck+4gEwkNI14oJdsY2tjCINVzS1ZunO9J6mPjF9uCpOP79OUz8N
QvPAHmBN9qtsHri7PBy0iUnplFncJr7Ap88yr4PV1HsGPAleOUZP7s3Fjiul
or2Zs9KtrcWP8f1zBZneKW8D0kYJNrTZnaur7xvcrbui96KdOkQOfYFpPREc
Ln6ves8DyM15ZpZIJ4OQ2CpVv5uqU5NpgDi4sAMOApietqstC3bLlo0PJMbt
k/i922okkaZM0abNPpCAMuNyR+cGNXGbA0sbtXBn5HU2XcZ8olT7gBZj8iGv
o3sbQCdxGahaHTi/l5ToBvJyTD14N5x28XESdu1tzdGY8Pj8YM+IXVQsCfds
HEQn84BFMVFE3Ir1InF+1ym2ui3Y9ogAbg1yJ/nLPYlXPqAwroTjCa2R07Ga
83MxWjGich3CXcWaG3Jq6iJd+mfhnlvRTMn0/3Bj5etpIyclFc8KSo4EQlLN
hmSN5k2DNSflw0H860GGLrgmsgCTV1W5X2Go6PwOXTjbZhh0OUi49RwTndNY
PdxkERHDkD7eYVCeF+JbD8Q7jd0grw2ffLX8KhnpePDLIjBbBQPinhp9+AHh
wREkPoOwHw0dFg7kPk1Im+Ni8kB6gFEavNYxYvPkGDFgisWWJciSwNfcq/de
OOYSmwY9fPqHqRKIEiDT3339RKu3UQi9VO0wId9qqRKwU7eLXdyG6WG6jXYe
vSH72CytRb/lzFZMfokVryeFToJD+YZyLGRmSkAovkxJqhkUW2V5qSnHirHF
5Bzq3FUsSrrwFoLJm5dBzRbXficaKlKtm1CiwkRk4rtm1dW4vQRjJDfF6aqT
1EtInm5kXmkkzCTRXjgJogmme14ZopkIiwpSovxKRvQ4uVo+UZVnXsSPG++8
iX/JeBQTpGUWHgRsFWpF8j1uQLUSfZRFMe7hC2OQUAFiXnRI2XAEMM9Cvzzl
AYpI6IHmnxUB1eH+CvIMJ1wfql+0M2ZcOwshhmoOl2muNOgiH+B56enEN4gY
jCzgoW3hk0GQsDDx2RZggPp/rU9HQrsnoBKZKss0zN2VEWusat/wFeO6LtRf
yCTNz/HBpoq3Ay8CnFGqt5amR+wdTFmpLTp6ZhPneX4Cj9UDkSd7ZUYJx1LJ
s9UEw8waHn22Qqq8CXZdf5i51HokN6qMqnW5QY1O1R7kK6NcZpikkpPypGMB
6q7fPTw+pVje4UQ+fIrNJ077hj/368MGJuUrUVFz1LSgyEQbmraE3TJktMLR
PDRCHESTWFj/DCx20Nbjno6lbvcgfvMboqqKAtZfO3ZoncYPyeDkETkiks4m
kXA0EVh5QNvkCClt0y1PtWgijO89RIF5KS/dESfruI7YaSus0ws+ikOIimPt
CSo/i3T9mnvgQEG8nlywcoF8ZR562RzrxzIoqSKaNzmLHKyv1Nl45QizsMhD
tY31m7mzDDygegbYGFhOlwE1jDX26OdaRl2qz2y9DzXql5Ga/arGGbe0p64p
ON0nyTcoDSED0ONwE8sGNqGS92bCBE6Z9YTT2WQ0hg4c+ybXOlNS41OG9nPt
X3yaA9432Q5fd8JZuZWrcPuwMniQMxcKPd2KxFLnwqi2ZxMvvr9zf9rSt3V4
RsuA7/zbTVpoiL5z6nrosGw3LUi5Z8HYAtPBy8bfCMSZsYAQJPSDUSbiCAqj
+Mj2Y62w8p7iDmcWpCjrXOZQv7EVoV74+VmoSBPQ9y+Uai/i6g5YMgoxNbMf
lHUfdFr1kZyZvuBZW1u0eHszW4b+8pYoHqZLm7fJ1vk41inhZpPwFJGtQGg0
Jz/AkOGHQjHeLHlrXJhOQh2MJYatPNDafx0X7177/x546AxaAzCJ8gkD8tEp
+yAC8DJtrh0XWq0x1m5w62ILQ9G7GyPEnWUR4dkNbv3w755bSEe/YP2e+xTd
zuIDFfiQD7WXPiOuAgd7WRPqVSMjcvCt9umBGZ3pVa9b3qLLBUT5qTpsn7VF
chk+2fJcJ8oMCjBDCamMH7wuaCqaEj6pnz2edlioVGlIl4R0eRe7DOxmNNUV
trZtSlDeEHz5a5Zo9kQtGrK0mehHb9TIMZBZs2b8RM+k066aK1BnlinPxdj8
RuipBAHZLDUJ9MH2L8LKnCrUb3b9QFrgbYI3uLcKnfWtuqcTgFFjOOQGFkZM
dRQfm5mWSM/Q8LtmDzxD72kaPPaJtzTjYwFAIG0IJ3Ver+gmN8DqcM2LvXif
oAAdh+aO/MJDBT6ZvlV64HI0cjmr3OcKq2Y3hQi6gGuqZUF0yPKLlVWHn0hv
Y764ke17PrfnIo6yEE5ctNANkO4D/jaODkLpAv0hWCFcayCNze7WkcpxrEIs
EC7qWNrpKme/kFOptL3MV89NuAlahH/IxZ4MIwqUBfAci6PmGiZtpgHzKdKF
vvUU8vb9MZ+a2M1jTDm/ELXaSGfNwzndUAd/4EpqGCSvU3DEuAlEQhgteL9m
Crig1rAMOKN/9gbFO1X5sa1jCKj5th15ltc4nwbhMzKlM4OFx8DRawt56+Tf
R9KMh5Te5nF6V0HxMFwmuoDMAciTBPSR/KkVixcMbaqeCtPsBVlhAPGTR/PZ
QnpX2Tp9pqloHOWoTKE8HY09Ol6JuiF1hw1muK+eimw6yF63QSgdIfKNBqV0
Y9n4Wp7c0hH5BuQ9sybbSUyyhA/83qbNTDzNperYY/B5/KR1YycubaMLTj2A
2puqqNqHn/bFc7Z1gq2Z3p8NeXH25SVFbacome6sbzK3jV9OYAwSPM3F9lfD
V6eadn7ss+MesG1zmCx3WWUvsnRbFQOsYVplaFATafU/SY7YFfj/NbJH3mni
+tIk/INDnsLoLLDQpzXN0IZ6YQ+yEKdVY97U/sP5EmR3S1BwoFGK+cp/Bm3v
6pu4UiiHF6slZPIqMP6xPu8zV2hdejWW3PZxjiMCk85CJG2rpmU1d/zzLLIc
SKjL0q+dF9zXAzOKGcomGj9p1VDhZ8jE+wdER1noDNCbxxDQSZhuQf2p5pM6
1LPrGEn1mIgGwmI6+SC73ZRjm58RZFw4x0QcOAuYGTBT5S03rh2AdfRG1vas
IdVEeTn6WKbzaASjKJZT5tYXzMd2ufjsF1hTTPRHiA2SEOCWMNQQnwLkycoE
b33gSG4K5VQSVq5z0f0HFor51D1gvPG8p8I2WCCQYdRwRcVENSro+zW7tilW
BeotvPh1rQ0UIr6rFMHq6ctK0JBuFMND+TLiEUYnwDhI9cPXNzft6afi0Cqb
nyu8DysxBBm+JswSyx+xUJfOFF9ugaCjL48t6qmEal1QHVd15GGf8HRGOAKq
43XwjTAnfb5V92/i6/RW14AJu06Oh/kZRWTkLC2l1bMv8+h+5G5tdRe3EWau
d6L92GULDYkqhUuVhH2SUUKYPKuaVDcaux1kYmpDXQMZz7GRW+xvuOdTWpkq
AaYgif8Eqz49fUkoXgdKSkQQaC1i13c3a4g/rghj1uPO1eUt7QoqnOIOsrTg
p1+Y0yiFMTjzSDkDU0zT2z8pBXYdFYWmSS0tvuB1z10EZL9irBzCEkdWascE
NKBQP+T5URE7EDzRf00KmGkQz8+jEgfBleLSh9PZezjJxv5RWho3NSnlqI8l
pAK2IsldNkFTGRgU0RvvMRnLZh1mzrnDnP5ZK8gfAd/nemB4sL6V7H+6tsqd
A5Z42gHb1hpKBOgZDqjpv76CU4NhL98Xtfu2S8FxD739glIT+5yGQPALTVOu
ZIwX4T4QUmHrW6Pvok5DvfkCBlmLwpqvC03TxVHGLZNi/QTDhnAbu/RJRu4t
zKfbYXwx5xP4J/Jxf4GiXVA+p5t/G/23onKYuAG9XJsgoj7WBPZPo+Mw8eF/
xx/lm5PrmD+yjNnC29SPRe7XYqNmc2aAZ1shSSNkq2tNq9MWqsutjaWwz/cv
oJ6UYEW8QuKwWnQSciq+/bN+t9O/gZhNW27EpIh3hH6e8V5WK+6tTSe9RPkd
3g3dD7bptpnwg6xyHZQJReW54mwW+TIopGoaHqxvGqvbmvZDYzB71hBWaVF3
dHOehdI+H5DOYp5NJuhc0IFg6PQZJSYoNbuj47EpRhJmkYnvA6OpaEFGSL0T
g0gc1m4RYBhF4mr8Gh4m4ot3w2xx0ZsSMyEOuh3wVjuPoasvePah40b2BNc7
DwAWkD4c97mnYYEMxk9n4fRbnIWCYJz8sR26s5/4McnJwRQpPEX1fogUVrYN
9ALnEb/SjZSVk4OmN8A0/X8DbDGUafH7ToioxQrq+c+azwLDI7FDJDlC2Slo
ulcDJsNRcvq2lYrWl7zYuYDBvSLqRrGCnX8Pltoe5GSNTIZd6upxSnFeyDfP
L7DK+2ZoTKHlL5lF+ZthGhJ6epx8xu+CDZUwuj/5BPmmV/FLDSPwjg2/U3Qg
2Z8uAK8EajJZLGPoU+reyPwk4zUoPd8gE4mSFb+WQjqinG5zQYm27kZQkuHe
MlMe65smBlAC1tSeUdTvKFi6a6NiwkDknacQQia4EXURpyxsveoVNYiB+y8j
UMd+4gYtfnaYfGV7VQukGehwB1jRUZL0BH5ZYPBoDF9DEzNjYYW2q3vdblqZ
bgpvdgvjZdG5ngCyWmHy1Z8K7HkVfXDn4G7DJ+bSWVVNR2z0QV545Vwf5HfJ
0hAHYXJ27D2KXumoN2cykazsaBPORhq5r7m2lddUiugQ6XXrWyjL6pN0+xuB
Idg/KAqJeFj7hbe4hZH/dVPX/povYkX5BfqTlTYZFM0qxYz2qu0i5VFZtWK5
0ahjHiMbcEOixGO77ZPtxUfKvKW1YeFZvPyv6diLpF2xqWjp5fB0HUgZdUYS
CWJ9kh1xZWRNAnIM1PC5vkN24nM0wdOyNhCFWJud+HIFcNAADYdsFPA1m9kQ
+XJr8N58/u1EeI5hHXvYx3s2qYnif5KStKTqxsS/mGCHdDCMUZzE6SMsqAZH
GT/T2n8XYQlj0vGbXXvx2akasXlyb2ZDF615W8yiRlo323t/6jaQ3vBCeRzr
PFFsmM6p/4H7w879/pdLkIIQ2n1BhbDT4XssbuDeCtjyZ20yq8cePMucXbjp
AlHDjyzafFZhhbhhRezzfK7Voq/RPCAElTZVgQA70iQL9jBCzjQrcSblZic9
8+9NAUrmIa2uELAfeRDOZf1gZddyoe9vi3K2gAiVJLudEnNgdCZfQ7mErQ0E
eejeOnK+wnVBAc/k11qEM1zMspQSFKiqg45xZ7Mk1p98wjOcNERLTbAhV2Pg
7uZVwLscx0I34uf1AC8PVpobFQmLpvQdzq1TU5iBjpxnR9V3NQ4pdLu7Cot/
evHKDOsvt9+hBAguB2MZRskvUoLtE4sJFkYQpgm5lxfrJOJCmFqDtBhyk5tv
XMgXYFgJTa/dIaJIhDw7wRQF0Ol9A4LclZJ1FoozPsjXbOWT84UDs3XVMBwG
4DKBFvy0NVHvKW6EjKo6VokdMZZ35dG33W+oCGViNUtjLetSDsPrGihGezvX
aRpp3Ms7ut1o9o3k//1CuO04xrBnsqbHIVEsMLXcIVAfnOOY9uPuKmXLPjGe
NvDElvNAF26JisBJF598yCLACP1fina80juxr/dEkm7omCoCb5KrE0askDrQ
S7FiNorDr0qxYNUqd5jNEOfOg1/KTM/Bq/bL79m3KZVLQQgPgNAsq3vACrXI
UPfvPikEsPQgLyTsINAj5MmxbKIxsqtr1ZD1J0TjeR/34cT4X8w8Q7Bykskw
6VWHGJrXmt/E2CMy+w5rzk7juQkThLMszNhBHMsOBAgyf6mrTixc5X5i+lKB
2Nqde9hICOzL/lnrYQB6/fwunBwJJfs/EVpTL2cU+cy8WJSAohPK0jre8NqI
QLyA/EpuVJP/ae7EKi6n7qiZ0Lau0DeYqHM3DvpWf97zbyXmIpE7osgW+8Ke
AGa6IuZIuVD9rhgcnI0RWx6mqLyBqWWZfuPG53jWA8HqfiFUmLBwcy90GJuj
6JCvyrqA2bKai0Q0nJBzLGny5MjsZR3t1yRkd6A+CNcoTFLV48EK8yzM6U74
/4e5kyVD+SJSDeqANTLIt8nnAMKU8CJNFMcUwJE4FFn7+zziyZ77qnPWDVHi
HZNG0iTjMwExjJsV1K0/P96Ji2buXKsf05qfBOxaflILfFKBuIKmlQ5tOQzk
E9WqWLXNYX/9SQu3GYx4hIozhQuk6tYJ+RRdKttGJUpdpEuPp/EgGkDLpww4
+zWekaQqd2q6Qi71P7NQldPWwkMBic1glUk2MtijCtdTfXDAUoY/qzdLR+xm
3Xjzh73SIjm9WF6tp3kBQeAm0eJmZEJipfpXFQLUHZ+xAVkR0Wzm2uS4IY7t
rLNgdsobAjzLew0c6U9nPE0lhv9HLLfnkdlne5EbHrHHxMjHUqpjXc364YVY
2X19QrhpoisZy3JlYa/n9opD4A5gKxOAb4oKqXupCknwNdjESqek0W8LrVW4
5qKYWR7TkgeDRT65xOLLRaBMAwHlRFxbO2XrE+gSiNI5IMR6bDugcCdqN92P
ww5QDyLfZSCVckApM8FTgJDUh0udThYKCaPV3HkgAGdrlcIOs4fEmNOJ345c
xwq6MTED3mF5HWVdM6K8ayrmnS+DdJHJmHQT91BZOjPaHednAoZbjJo5g8IR
APyKF6SjDpxscZnSXhpKAY32UQkQwIf67lVUq1lFUL8ZxAuk4a7xlBtenaDf
UAB0yqXvho+gLvQZwfzXbUyvufBcU0S+m90iHMNyFeZ67e+mL0rBgll6PuOm
FzKJDRAahO7OwNa3GRmZltk2IMD5PO9lAArO4tTHYk9y8gNmFcKF7VvlN6qt
vBkR3THldkjRBBN2fWpkutECdaPLL9FbXxUk5yUjqEGtCawREbD4A91xOZIH
SG+CYg5AwcCwlnmhkyks6/3l+GYYT9EQXrH7EMxlVdN4I7GlOeTK43k5Z+eX
lYvwFiHk0lseuWYsdJAP/qqnPAaOwfyh8T4bCGDXnLokp5J3Jiyztjh19u/C
c7ew7GVy3okJremLWT2e8G5yTz7oEI8d2OfcSo5e6ILjb4iumHVA1Ohja0kV
fazk1VriW0Ua9BkYwuvjKjbAjKxkjPLo4utCcaKf0wqqED4Lf+gCuHdfqZ8S
k4Hzo6kyqK2Bb4DwpNyG2vK8BEKK3rLY1F4szo/4PAXHsEnC5bLnQkaNfnsZ
SxnICfCf+QnnCzcbpxhFZ1h8ZQsATt0vDoV3UoRdQRZ3AcNq0CTjC44r+q9J
DkMnYDZsmAAXUDY3PdhEp2s+Ec9mIXAD90UmMZCc5opIghfZTVGcOEczVd2n
kOJK4PE3s+xbVdr7D4RpgedV/UvY7OwrojPGC/G5mvVG1wSUVpaTm6fIYNum
fxKb+f++9X3N9K666ulvplG/7Y6AQdqKl1GBe282cFaC4DG5XcDZfex3mGdY
eFByuXQ93NHHKTF0Mn7ZkxyQr6f+xSju0FzkrlVuqtpgW3Bgjg7QWiTO+O0S
fNLORNkVJYMnQW6FhnLffF6/5ydUU3DHyfCtlj6B+sZzxi0CVPeske5xROtv
o1DSBKv/e32adOSoJMrMxKx15A4fxwSlWr2yLXGxzJCdp8lzD/jnirRz/EiO
P7E1B9hHuJc080amnfKSGWJdkD2tUzVmbYYvS80dtAusaLWaKg/0iHgQdPQx
NNNvNgSzWeDP8WZH2YZwe1O46HsmDEfLvZsOybrD8TQkMVJmdv/RV42EI5IN
7irB3KhK2uNx1cHGHJ7q4rU/+zlxZNhOxwdDDYp/sTT27iF37Egip0/jEfnI
gjqGTN8U+nl4c31FhX1XXvkmfraoHTuM/AbP7nHDm7r919JOYmSxHDb7VRck
SBTc5A+oYsqZnZkT4KNnjMA+jryZh3unhNmDtYKKKqgnLDAXh709ba3KNdyl
UBWBetx/anyuDTg2+nHYvvcEho7bQ3ppszhT/paDvfrpBNINfjhkYcsCcKeL
2n+myYXwizT+mbYBr7ktPHSLDuhcFz59J4lDrYBdGzY6FEjaVD5E5mwsxxo+
atlwfZzLYlN9G5eMYhoFJk296yovCUNLixCwqDjW2CXvmDeRP0eUM6ygKVXs
EZ3Fzs5Owzq1kPgTCogEj8GiCfoiGGCcOf0ypRrXoLSKAnUh6CsOkJVJMNo5
cxEmCqYPhgZ8K+kf3ytL8VrTovE0CreofI9hsKE1Q/8T+XbNXTKIGdpSdoQw
DH4w2bP487UdQ+XOnlzX0wC32NNmVSlERsuupp/hVn1KhKitugJRfC3QhbwD
44MwsaB3gBnufGKTfyDkVwz9zmNcOai/Lp5q012eU+IWCIEhfzx/buH8Kyni
S0drWEga9aJR2Bwz5W4UoGdRM3AccSvPKTUyrS4Z8+3PYiwLLagfDqhVmZri
3q5btxdY+pimApralm6wxi+LumOLSIXziYmeqHmJiChv72eVYs2FeewrzBy+
1vzBReP/8/caoGi9IOXNGZ/SFkiYqq3kmZIm82T3fC7mCxLpBFAWi8GUbTSx
x1yoirwczQWhl8f+t6RG3W90INI43GcwexxAJK/k7N9yuhpBdxiFxUeGT1jD
XCtELfhPIZSOYMqx1s9VXpJS8Nx7wGTysqmu44a0QeC9ojokRlP89Fl5SuSb
LFZ2PUkE+csUHmCInlxHa8dmf9KzBzakQkFQtrOGMNRcKCWKUfFU9trlGUZt
Z1TA4KpEsA+Fbhm4S67PvC9bc5QbJS+QgDP+xhl/YuHwTkb3ck6DdKd7oXqL
VCGIS9gyem26crALuPRGHq7ldn55Xst+HY8NBV7HpF1txvT7PQ2GopDMKmjU
8ZvY6do96DhtFeMR55FUybj5JYLt65GdbF2lD4MP9doA5jM9teHzdb7VEKW8
pACjWoumX85nbgK7HI//LCg77M5iFGKALtiW+UaqJ6TJXXy0hLLrP0Ggr0m7
4YhzTdAjX/HdwankZ7pIjzaXYlz2JhV55B+WO42dviZENpTYtWG07v+8wkDl
xoKvgNdnyifecRK04V7OQgZGHeJKqlbem+cP8NgikN68sVDpFeQV99cnEl2K
Xe6VvetP4IYcJ3dseFVfKq7wQWAAeNDECXV76m1aHNHwclGMqVYQBxFqFEfF
4lcmpXU38ngs0521Q8yoY8+Xewm0yJMNYiQmNo9sKiECMVl6CEmFdIhybAd3
pTXcHHDhPKiZC+y3ytuzRotLC4HguljNwsfn96zl2bua2YKi9mmcH1SKlxYS
mXkbe6ZkHrNhwpkvJ3E62yMtUAm9yB2qYxJfFGOHl4p9VFR0kGU+VT4AY3IX
6GANE9Sk+oUyOMQ2iFnDShdawH8aCdANqYMIBhXc9Dnv22zVKhYcWJicfrnO
6Mh44DEVjaqc0s4lGq/5uKCDXvDd91iiYW/PEjkKAOHbHht4jFNd3ZKINtn4
GGFv7aVBCnS15NV+LUuU+6yNEytK2LwPOmdxjiAWuUbQkESy5XLS21b322lw
pWXR/LZKnzefsIbtD7Yv5XOruDVW7NhQ6NnbiwQELZty+WSK5crdhWjsn3kz
0zzB+cPgd74gndeBX396x0q980RB3JCmqqhGYrNa3vJQZdMgjy6jyVDPHmaj
mO+Tvtt1Wnc81MSbyraCh6ULQj1xqjkavU7QfxcE+/ldemM4/9NcfWudI+Xx
AVMJ1rHn/gJjyLOkxasCEbWVt9SjglFXhNmVCNlf0RUKDlvhJ7Sdapms2gRI
xE6i0w0dp5HKRT+X/Y8CM8Z7rn10Vi5xZVLbUDSScAcpy1J6QvC+yeuWGapw
VNOTSpTHiG4stB+nf6NAzINsIlrif1iCFiCorNw06Rwq/4zbfuK4Ps8DPzj6
JbwB2jemeqIShWeGX7DlYYv3ax2A2vE5sHYj1eVD7QDAGAJqPXpqktkNu0Y8
3nLuG/PIQcOdxU3n9LQ/RaB5dcKTyxUflzN/DFqchsoqCvAg9qZwvVf9DBe+
2Ee90Zz6Nf1KOWr1Jcc+j+jFqnyxuNdKmdZtDJVrH7wdtALy7TEbo1sapbeY
x7Fb+feQE8j/6c4SjkUvL7926+BbAnub/7gX8qWzsk8zqMtXw6KIkUwALrqe
Zq8OWn4AtYY5dKIY6HhM8C6z6H9EI/HZQbbPF39ikEqXJpO0w+kkrSLTSONz
DPNmIMGTCTcZ3ginxVHYsI133T7jW0w+4RtJ/3AqvSY1VsWiLM2svGdoVUS8
VQ1098eyFwSRKFBNc9fabTQNw/Kd5xzKg7sRmZfvmR4v6NzXAHm8A/v8pUw7
cb8WFqlYzbegKGhXFDL1tAxIvlMTZkXnIw6HqrjOCaI1L6Ke40HBRyt15QiF
XmI/Bakc1NQAesyphvb2RuDaHiKqSsGhDD5ju/w944J70Wwqntkyi0ekwoou
IRlWvYsPZkzF83pl6qL+DDrqPZxcoFRfzcknOKgDZlizSgb2vAypN7W/RtqS
6o4dHB4ul510uTvoyTrXqDOsBUrJ1fL9MXVv5s+LvKKvEqtZZNSC8d8tMR9P
V6EN1QoR1++VHNGg5tZUApvjYCWd+CReIFn1E6mMFNJzZxhwc4EYVfrMwf34
oiBFF/7+ZjWEDMII2tDANmQndWlhJEtnpIMX1MeIXEuL9GVqF837PkBZsRBo
8LLgt++7l1An8B3Wl4d8Z/3SsAQf20ui/c/gE110ocGvKzbcR2SxMW3FoN78
RNZcppM2+gm+W3h9XjLCqDUyBYm3Wzy6BE6iepdnD/wBOu2ioTSYmHxUxvV0
XNh4zqI2VwWL6vGitiWsb3tG69qI/N8C+FW57MrsTWhsbqaDKAYvq6ipYT+D
n22wGBEb6iI1zD+MOLLx32ntXHgwz5MnXTkkqfAbAmuG0PZZ6PcmTU9GcAfR
DoE3Mg9toGHzjA5XNU0zIJxXrHJ8mcqdH3OkLk9vlnt/dGPxUsM2jknD86zW
AKsu+Rm/HzG234PmGB8HKWB31ZPMvrZEwlMbQFrvOgtkxMS5NX4WxwO4fbB0
wP32aWcONSm400uI3WvXeVCpf17Ay9Gi3RCOQgmbWnEnYuf/SHRSIUg5j4sm
W8k0WYF9PXDyedtdAC49gVkrY2fqPkI5FJXKTdSe8gHpKhG5eANILy6xJHNd
5+epVQU39UnfuVmPtw1J7FbK7b0+XeZZAejXXuF1AFLWiBXUg6sC9SGriUrq
yArWlqxtHkbG0YFzMWQNnQTYui/xVhpJef75dSuL5tItpdzM9MH383JIwmqO
7ZFaNCU+Mx6UDB3g0obGeI8jy7gMVJYO6HXmLp4+sEMnsJd6FO0h0Si5j8go
06LEf/9C4daBHTNA2awX2b83SWcedE+llABcP6JJaVfibV1NUMy7qrPhijIx
0yL4ZDE7PfeX4QhSgIBFsBD9OxczuxIz6QI8czjKYXSLoBPhQE1aRUryP6io
xuSl8rgo977WV0gsipyCUYbYur4FOd2Rbq3WxSFOllXa5QndKIuz0BYzCLPh
+xKa5PLamctRxLcLJOvAzhdDeIcoep83udRJidT0mqrUIlL32sM5dDrI3ya/
h/4PEnUu9TyE4fuKls6KZRL5cu1nUZsOjQd7y/1Qu6uGY7kmFScpUef5DoKr
Gn2mg2VEu7bopovKF37rJ61bDXn9QV4+CYIPpx+GqJuxBwR0XthvliVMi8hL
nEJIkmfDjuyUtpzwz8RViFqi8Zv6ul6OUNlIWXhETpXg2yAXVz47fp+Lmzjs
E8Pl3BiMt0lu7Aekm3Y7LqG8aiSCTH4whj3odFIRezRHSrqGt1fSLbuqetl2
BAntNP8s98D8vnujYGvmPMn1l5qRq/bLBSKe0/L8Z/3tst1Mh9fzMADjBpSh
DK8HW984sF4+5SOtb7KTUb/1JfTi0jMmfAUmBTP6UWBNy1LPvghCR9gAWlv2
d8d6WwMsbDYLsK7MAbxmlWyeFL9u/5F99i3d3CLTlu9L07j1VAt0c7TiXOO8
QOuf9ze2t3Yy1YdwLOK+qu3TR7XCQM7EA/nEHqv8lMy9TSdNv8JCpnd5plR0
0NG4jFW+hsphyWtCBKq9oMewdwj4ur2pCs6z3oeV27D/1JVMavqm3bZ0sOX0
wHC8+IjebhXCLaOuPKqHj28TqgAZvjd+gXnMIbz90p7X3SW7r2FQEo18g4kJ
2ifc1FtH46h43UprJaugo8lrr3Zgq3Tkf0jP7+or7StqNWin5GcC+cauQl0r
8Zm9BARwEjMa+si+QpSE5HLZKZ0jDNsF+D1FriudssVaUrcOFKECH+hIQHeB
WZf5zPOTSBemVW3YeuFUJXcPgil1e12+Ty8jvI0aVAsAa+anR+odpLjhIllS
dc0kTzjC6mSp2tcgNOP2GStd0PnihT+/IWhjR6sSE9WxbUHiEvJ0gEtLD1HS
I0jOOBQOBv9HWWRSeDt/xfwBEa0rfS4kEBhK9/vVIOuoNmNORmJW0WhMuw45
VXtF9/jyKVzQP4cOLAIBdvJPoikKy8bYXRlxWOfEJxWZDJ8U85DPmCI9XV0x
yi3fYwMR1zrKyHhomsIk2XyYjlhLzCvYC8ays1GwvfjZxttF3iyNIjFiGp+r
lLktpXSjEkpgPl3eQBy5xTMVTovUfVict3ZJyVzsp16SPYcS1PcyfW6a5H0u
vdTLp45fUhrpaymQQw2nqgwZyO3DF6oKTOEKN8wAb2TCXA7n420MwxYasY7w
Ur/Z+FzSVEKEmt2TcwDhZBAdvV+LekkBoximf0OcxQ7yrAQrUF8GZxA4FivD
NHQqJTWyoL6CgGfphypA2Dz/2eQhoyK2GDfzy3E6DnhDPkKzi5uWPyCGobDv
A0Ainb9j14Ub01ZgR+Jx/Qzxvm7gP/IAAwfvxrza2yyWAoPnkkm3/3WzLqCa
Ngqrfkx1iP0rYzeMNBHPlR5U5usBjLtRn2nMOWWUbrMDN6OjAmJCllS8eWVx
eZgBgou/z5U/zuNbq6YiJakhVwVB+EK6o74E0yA29fwIZ0PO8GWa3VUzQ2zs
dfbJcT/qIJtHyygItPHaJ882DoD9f5kZvxz/7lzlQE9qIb08B3wT27iVFRrB
xzoxqGZnGG1MvEbXatEvXW6hKlCf75aahp0gTMaahh1TR6rj9mH9PnFEAbCj
ZE6R/BfvzXYGEZgIinnRnUntgEZs09A5uEKBdFmkTFzbAOJ++7M1TdIMVhQp
THr20LcBezOG3l/tuM/bJGLHD3qkmftRIrubEOyy1UadrNP/iWQMVnG6TdNd
a48sLNPR5AuJmSGyiXNw/dZV7h+lufqaINnkqnueRtGk0quxeYCwh5rrc+tI
I16KDrhl9Rk6rcapNNoADSF8LkxLE+tEm0nMCnp2uGjC8/XBXBx6bohdQ5t8
FXqDdTbrMykfqO8hi9vQWD22AaNf1rrm6aUHy4oHYxk/H5fOKvBH8WLbrYKR
lsYlgNbQ2lB2HIOeG2E7SFYGrNuJqKecKuJg/UNR44ABQXgnYXS0h7H9KKtu
Bt9YPjjXrfFNpODWpB1Nvg7RUO2IvsZSHWvSQjoPqECakkLBfcyeGZP6Rs7U
8g+vdEWDzhdQMLoY6aQO5L4qnM44S7jf3N5vBsgF6d+K2+biq266ufibPBHe
xsOqtqmXiBm4oWwRLeALcMFpPXENNqJY0FRrpc0Q1FTuDIoSlbqztllvqUV+
FVPhYopYxik1GIawN6WuOVK+DESsakQn+4o6miP2NeDzJyCJUmXpUswucd3H
BopWc48T5iH5j1aKp5FVHw5q2eI1GZfoUYUp6qXjf2J22Tgp8bA6btu3YyXE
+WWjp7hREShmobrfPRP5EEMZYUGggsD+Y5t3j64X0zjEDXlFbLO8X48stKOw
YsA3ftSwQ2/Ry/C2eBgLDkOhrB82XLjdxX1aEcwlKV3qT4H9yhQBkxkuE0cj
fUo9cHbK/LI1qllnrTppT7JY9OErE3p+lsXCoYPj77fhTuRw/ajM5ZEC1Alz
teQmuyR0GnvDWi2c5cMiJHbDjAMdF4dLhoESAUN0ThS1zaDYrIzfGRhcgH7E
oc2YTecZpDwXovZ27cd5woQzYpuRZ+4ybHKpQePjA6OlcbIVaYurSsrdh8gx
AwUXirGeamYW+EYr1KsYxRLf1v9MwYaaB16+fq5XQNzQvhGVCDS7XFl0PlPw
XIXT2T5cNypdlAn/9HlZBPMu5tlSqwzDOAOqWAUYQ94U/4tHm3RNY5RNRLlw
T6oa7tXjn73JLzwBLcBnK3fSIHCNtL4Op84rWHb3jrwce0cguDmPwxjKi1DM
x8qN4E0YH3oC2CoGqbMzhi1fACOWpM6EDd/V5pEyw71jA0QQfqQ0X88GZbTk
iSJLNSIm4m+34M8o8MQ3KGHFjcI609NWMQ99jyhyv2aZfq/8HtkTeo4itYCg
fRwdUUTtiRHPWZ0E+MjD8ffnt5zbX0oLz9kYcE9cI2sy0btYyoIWD/eFNBxI
J7xfDA8AhH/cWPPTE+wufwv6G9T/Jbp8c7b9FdeCw6+AbPZAe1JshrN5H9A0
LL5MGgxTYyE2DxjIxeBUcKXQxrGOZrTC05VGCkUuR7ueN6UmoBODqKCOP7Pl
iLuaqEqqhmld3XRXqUxF2HQyZuCcKwkmxdlwQcN32AHmUuFGqrIOGzQDfPDy
ZJr7696hkKOoi6NrQPHeVK6n1GZirzruVmh+narH0zE7TMGtDSeri2FzP1vo
r3Y/QWzfkiGHrIh0wguqm5c8MzSE0p10oBvONOlwSmN1aVfXTfFe28jcL8pw
SAEbciF2k7gc9dw55NxZqhmW7+FvPZ+3plxVKHNVxnWUQCItBiRKi8hYEMFD
Xg4AsX/vkN+hFG6hrwPP8j6mYSO0pz8ygBzVUcL2YQbaXH/61zOU/nHSVm7i
rkr2p2VAyuW62DCDFaA3of3Z8sPrqHlWEkzs2mF9LgCevy9rFmSylOVj4WkH
R6vDzCpXnpfmlTWWuK8lgO53Obu4eYgho/i3DaLRAeIwPQfS1bV3LkX+XBce
5/0H1fdezb64bV3NZQEvomFwfAYlPp6nxzV7QWwCcrvpLUJCp8eg5P8BV/ot
YmPE7SushN1chHlwWzuZ2xQrjVA/uwGraHzZsw9gz0cQfy95aEdJzbhboiYQ
sysb0njoDWU1BfWSPl61ju62NPhKO+uUDF/O5+gnM3+DUcNoxybKW3OzRDZ9
1jhPy44RBpAi53YO0S1QKjYBVZJVX9+XWR8OtMcpIQXYILtKxltKnB4PB6oI
RsroI6fCJjxjHSplM64H0dop7Ul8CFO1qqHA8+TKlPlwkClAsGvMcSLxu3yX
DTd1pLkihzWqd7XdffCpAC8ib4YWA/SIysVuFD6muFjKTpctMfYO4nqX3k28
ktECpB5WjySZGQr+wvrHcLTaCGpVO2/uXTML9IADfWbLjjbktts+K1lRDVRf
zle3B1kPdwkVJEm1DDSaiJrTvuxhrSEXTxqRfb/f4leeaYs31w4hzeisduMd
SEUd0PzCZbuWHsGixSHeQbYVpDrt1FwweTpfq7qRCKm6fYrYehGZ9vbU89zW
TRVukDmnA8FcqUZglTF1psfeqHwRdJPcHd0ZpfpY85k4zgmlJ5Uv1eKUCDBM
2z9BM8Zi+EM/V3/AHkpwIxuqr2vg4meDqItZF6RvrdWIXCVIChG4zOBZV5Fv
jLCyos01Av5jdxPRY3MJT6H8efqR3XAfROgQvLtQSkPrsdvlEWjpfFICParb
HmPQBkA0VSwbk2eDer2duMHFNee1gBhh6noxfpLxrNbX+crX7IsCrvUMEIzN
UfPp562fDj5VdwPlUKcAOiy8c+afgvp1qqF4DJgXOB2tKjAuDGYgrM4K1Pd3
tqDNQwLAeXQfgOib9UNm1WUNNAuBEaC+wH0EFCLrzYkL5s+sOExSWjvyphBY
KmnJ62V72euhQ8v5DbinZiKt/GTe9iHyJDZ0rY5jZOBswXP2qfGQ6fkPGPt/
sKMV8Z2x/5CBmYotEVhhJt27goAx3jv+lPizoUDLSmJVlNSEmegOOWNi8WgV
IFAUNzr11PqDjLY/7zsGsvCcZYWd8J12uWSirY1vefrZTNV2knvRH6v0eBow
FH2f8xi++cX1xbOgFHNw9cA24o9+cGJOqTWBJKw2T6cYuifLqOGbwToXZ+G6
eh/D1GuVtbRdr54Xb1TtThDvHoEgdd00MQK32Tyvwq7xr+zujGt9ij6TlHzF
YWoXVDjgcQ6QVygBB5v1uWWnGjX4jHvOuUexB09HihYF9bYCGL5xejW7h8vU
rb29+Amn0sKYGMb1mMQ79vYlVevOQ35WMfQU9VyigN7MlF3l/HD2s2quPr0h
wBdlxNCUscS0Z6qSMrnKuq1t+R1vnGQv/q5hbXVgFPdQDRPf4edaMAVusgMo
DawMQDE+X6Oj4bP0aJE6fwPHoOXAlbLOnOek7iNQM7QiT70SFWoX7OAoC4eQ
eTcAwoplr9x09NJ/oMGdLgMvzUmzoQNw6MXxb+xxOtZ51DergDRk8Ipehe1c
TZzstEYYFOsRecv/9Dnunx68uvD9j8hPx1H7Tka2kj+CBcpRa6iIxeMOKpi+
eJ9EPlEdHinsT5oi8Cql43WU2YCqSTqsIvT9PjvbPuVvzwQvo6sp7u41pM2Z
SOUjyPCWTn5vs886q56YVBXF8+5l7E0St1XQQSZX0iE9Pzi1nZgKvMeRDuRy
qdJEV1bW9M1RHA9A0H9HEqrMRdwO4J8Dte7qStC+gfMxnEf3eFMaSIqO7O/6
YmTphsRxImkbRnrJsC9R7ojp7ZjgHqfSqwPCqKtWCkDe2SPYFZu4PTkRGwTu
5CwiNOqs1AcJukJWT3rW9QUNXNzOQgLCTrvJSeHjg9vp4nE5wB7kwFMEANpA
xJPJGtaj4m0DXPwt21rfhHDBjr8OCcAJKtMlw1dP24Wr7sU/EUdZv9rYyNuO
KHW+ipk/4e8Xj8RBN8psfbh8xAS9XYrODuxZQj7mZqpQGkSj7zJLmYhEFX3Z
JK8LwN+UBkF6OwtU1isXYJnycN67Xy6o22aeOL3uWG35jA5zpAPoAQyDSuPx
MXnWM4qXdx3Nt/UmfGDAFM8IG4WS2SLW4P9TGXi14AbAUxjND0PdF1Xad5pm
IeF/WcmwhS3kmAL3haFAqVixz4lJfESzw/wRZpFDu3c+QLScIdoMnwge3URj
laKfV8uOllHYZFOG4Kz+I7Pw21jt60ifQLt6C8wurZqWzA9n6vNHGvwH9VYg
1Lw1U+6P6B7AJswcmz9Iwhjmh/GoYBjam11/XogLFU+1DAKa4RiZxaZp5J0j
aKv8IO1hUivZDMbXdO2rDbNeGvRn/I98K+dDRYYG6bqu/RjXOpyLBE4vvbYy
eVoYANakCZVl0eDpYFNS1925L1SzzNWDaMQUBIMdDTKgnK6EtTgxp+GYJRHW
8Flvy+HVEoWoEBEhbhAowKzJTIEPK/0CtZPId2FE+OkADI7J548/8cK3AHO7
E7mymEDYekAXdYqgt1YENNZpobbqpH/kqryDTThEMgyRKrdNr1xeiEnWvxtU
qpw7YT8PMh6hyhj4S62LB2v4XvqhthRx+zs6o9yJdtxCTxxvZTFIYk/9EvwS
lu33v+1dIRrjpOBDDJ5WlnulGlCdNsFmCJRMWBnRoTfG8jQyo7IdxdSdvYqv
zMoPGsTREb0y1oHUPlqm8P+sWxy6KTdpOdYHXogsfxADbeIIX/jgnMxUNBih
lxB0uEh6k4ad63B7n1xovkA/GPQAC56kG74R2DpQlq10A/LOz+mffNQhLrXj
XvGW/vEpKNo7ipKkIOR8oadl68Ve1Y6AgE5gh6Ty6hUt0/e35cwGEx3hO6bI
4qawrlniFzCLIIY9L5rVzHsKeoRoj7muXMVdaJWw1OC6wEk9gYyLhAsvufhk
n0PEEgOvWhiuMliNllSWVYHpoB7cVzyqZDmIx9isFKzAHSqg89fNMty8Fb94
J/3O26t12nvVe7ehTKmtKeiC9YnQFJePAZkvLwMv7Hu/cHmxrq61T2+wQRKB
yZVmq0RxYunH65R98UHKFjD4Oj+4dQ4OELGGdyvwFdh93Km6mraT12x97Q4E
DA63NeVhLUHaZEabJcQRwp8u4UhF57JGryQo3KjSeQHtjaxcw7Jr5U9xR7Vb
IOWhdFF+xpVhQt2OPF7vrOL/0Y3z3yzJgt1m2HKv0ylg6S94FBMF4iedCAy+
do+U01hzXl5oWQ7FkLrYmvm9wECSICHLcCFddtEDl4KOIjUG/Dn9M1m9shdc
Y6WRlB7NxzFgtvFklPrR29kNcQYMA61CyBeEeaBCWIES7MhtWTm2+wcHN1MN
j5SvxvUQhKcEfbprKmLEkrU7cBCyUQPbbyL9x7r8NvdXPHClHR9SE9x9ar+9
6SXkrsIgkixDj7RKJjfxYHKuL64nBwTUY07WgoUIcLf9cPcTeoBadP3scIKw
j6iv5Kxxi0GQCaq5H0tW/HfWsBUp4DmpGF4CzPOWQjz2598mNPBhhq3AEcgr
EI0cija4nYTEmygt8RbUNtNsNWe85nmhcl5juj+zMlTlxlc/wRJqIXKXm8d8
AKbXYVRr3tTMvOlNpRj/rxk4pCTVWZrfcxmjFog03x7OUGBYq/9AxXgpgGn3
ezScILLmQGK92SHlo6tNyuMaamJQBGsy9apgL9U9jLiO51NFJqmT1WgsMM/x
L8BmZVDsDyQZXAiTyNMuGcjUzgFyss50KmajVpg1i2Y/USA60c4SKD3A32xv
VD3Y3WYW5awwrOkna/Dc2ZYI8+H3Hljcj6g+qF7GBV+rrV6fGh8No6Jbnl32
InYXFV1TWHkcZkrf4zaFzeJ3pYHJask3b+chlA1lxROd2arw1fwkzQaA6e4i
SBRaSzpnhcQNtZkRQ/CiG6ERf763uAtwi+hHqgdcot7Ss6/rhpHYswcbB324
Ll2TVSs3iOH90h5j7aK7OKGXQeBOfU+7ngqvo3yycmQG4yn4nuTjQmofB4vG
RFg9CRy95dSibjhVzlgkMZb8DPRamQp/bUOxmcizFap2lPdOZioBJsmaaRDZ
87bkzgd3leYpMoo15Nc1dqyoBBITDkUJDsCEhrWuR2Y1KameCWN0bmSHyx7s
QIeZsy87JajYx9YpDr8sLBriVmb/XKS/5O6qw29SSLNIHB4zeakRTTH+ys26
CrxOSRkMGy4wfcOQiiW6w0vFhnCg84z/xIhOKzJQV4jliAm6v8IM0687o+nD
YoDAfkEhhHcB4aIMBhlHW8Or5nMvWJSCrvW1VzxIOjILJw9ECSjdIIhzh8Fc
N8tzBTqfSXaJQWsjBfsZMzejlwlNftGSRZYCmF9cwEM1wkjVyVpW/Rg9kzzH
Xee1sPruEhEiB6TWGmK0ECeYLz6Gt+n1wR0E6rOi9S939uO+tCYMwr1uKKo1
99+UcKaNd1UTB6H2ZRSdww3VgytdLPN3CRp1uPnpU7x3RPMSJ/R82XTIWtrI
trCjFHDgG3MBrLnjr+gT5HTJWBcDlb7a8fA8kjfbH9i/CWtZx40M+9ay/W1x
Q1I1rNFa8O3nYmpsNuFGTYfyBeArEVZF+O8kvkIuDPN8Rh4BwjkILRsTh9PJ
BKuRWFKDKnCQ3SMNP7/YzoIKLQz1H5fHf2rO2+YTD03kR0G/7gWj5DJDORyF
v0YQEQ0sEIRtf8uU7lma7R/z/DM6ES+hsvzcghqqgg1FCUu+s3TbWGGRjQER
2+D1i/6/sY3IWH7qYqpDVQUAFhewKjC3xe73N4A1MqScOCaEiOBNzmR4S7f5
u06UM7BWyWAexduwduzvb4gFAzIbnuI3uLvYUVh2y1qTrRhxXFwmSv/YN+zP
VOn5GbAKI7hmsez1F8ej1aFkah4YwESMyNvQrQawsnmwpX5xUAWdnnvbcs3c
3fx628OPZZa8SKr6xJbah5Q9cfxTO4Xb/3S3lIvUfcGDfe/3WhtmamBUtntr
Um9+2r0dpogaD995mbxV4fmHEYhPX0/rJBP9nfQX13FFu1mFhL0osQQ5ZXxC
uSwjAclufntH58nD7cDVgvR/1XjyU/WP/sBGnBimVi3rTM4vJvfFLnROaYD0
Ls+ejB365UXAb5OO8rul4akQG7qgsOTQ1xB8zncqvPglIAZn72NNf8kDJB1H
d4hVBSg5vbe6EORaTWhCAekTWLixDN6WFw2XUntQ5ymmYBOHUg/ijmcDBZuQ
7kb0NCx9EwwOUPcb3cBQ59I3PesQ0ljpFKavitxEZwcWbYh4a60r3rBQjxVt
jXSegeBR/+wDxqTa0ijDvjhdBVcBXWH7Nd6g9SkPXlIBM8XmHtyFyvK7rRzu
EraL7CRyN3ZiOFKT12tqq6T+VkEI0O4ywF48U/MHKLFurZ83MkFR37FQHuFC
yNtjdRdVKsR2ZwByx20c8MYYjnvQTnkGzyj0brIFd5n0QfCN8ikConjZvBZC
bwfejehEy+hTZzlEU+tBTbBlx27C4LFeAkIWen5c59NRa9nxvC0ZfiSv/wXY
9LF1S0SQddx6whGa2Y47ZI+O9f+GDej1oNMoIA9lmrYo+Ot8E9i7wYOSsQcF
g66xqdGSzmzVm81Qh+j0+9JmCNBCw9NoqMh2Yz0ZakggeMWdYjNBi/J22+sJ
559NNVXnhBVP5BYNnNwDdcN7/Fbig/sQr5FZFiuxFLuGkY2R1sgSeJWkCppX
STiH/E0l/711ImzdGyIK3v7KshsaOKbH2UKsgaawzAmif0vvv8y3ZCQ1lZDZ
SnY3TV64XGquH+aLqqLW4jEjheIU7RA4Exxsrwn0fgEOM/NH+9WNBPl9WfyC
bnptr2D8n7n/jizsF63rcENcknEtRmJqPbrYWQcbM/7OyurVfrmF6YuR3nE+
QZksjXoTKzYaxI5Arjw66WYXoDM2dmEKDPJsSbccwbkYr6l8Aj39YGt0Bvlq
fTUwiO+h20P3VqCtgCZR/nfGMIAqaIYvIypK8o2u6GEc1Cls9eTZgqWLMvoH
4elJUFUCrx+L7A5F8U2zanaPudlSfqsOCzQS71gn+5nH7K/0+9fPw1/uHLdR
odLmCvy4HbGQ1iczVulr07STImiDFz5hnWnbYiX1CL5f/v+a5gV5+zb8Ojs8
TxOnqQDI82fPR6f5m8PjjJu7q0E6EqHhI8ZT2RYq+JHWaPqJBLB2OBK62hSv
qEfNjgXwiHI3yOiDRM4LQ5eCfHa6e7ki7YEUKZbJSv0J1THnLhrQSq1EV1l0
Z6WvkLGRAODEUGkxNEU7Iv+31gR8oiLkN1YxYRSX0f2vUzkXpSlEbzrbVqab
raLN+1SsVGT/NFzoe6m61c/ONLPTjKKQ5J/IP4p5GS6cxeTwEaQYqoItsBH5
b483JyOSDzw45nKq0Kl/RZGcVHqi8QjbEsgxzzyWvGfirtTGOkKYMiyDA+Ho
mPW5HejUBempeqkkfYHXYCw1gJGBkYWNBhrNUCf5H1kTQfHNalTi8MeAkrwr
ZJ7FyJ72aL2p7R2blCOeGDbbLcNCDZ/4XCoOpPgCfUwEILSYmX8zT5RT99e4
np6seiDRpHy4MSOh0pMjVBU1erTrbuHQn0gFp2okw45A4QvGkvPwG7l21yBp
nQqxNPnFXevFiwFrSYWiwhEvqUevNBqyZe4fG6734+Qt2UXLe1M9icWGqrm9
KXPYMUYGqeIDsNppMa3fZk4bnpPnotrSgl7RLGpog1a3XX52R9O8Ei9T5kaG
2WR2WOxcG/RvjvrpZFSH9ZfF6H9UzWEzxGTK4Mwf9B8pSBX8Itc7bs2nxXiE
uGH1WGQfr1ZptrgI3/9Xkddv/sPJUdYPeglxvDkZjkEq1XxT81FvibsCywvZ
pBr828cbl/YLM2nkZe97zfkeQhqHVlsvnmUT2joVqufoHg+VErPnFqf+OZ2A
x6OcwnnC8XaLtgOj2plV72YsOZpebJYpF/lXRNDjfP+JReRFeTjGR99RmYh0
1Q6ikGMurgke/ZwZgjjxJL0ImvogqVnzBv8RsBBUicygtkLm451hkYpKlyEj
yEpN7mhtV7aWlZqwJ6xlZfyVDxDb6nRjmbmRSx8qa1Rd9LgXz6QrZ3RT8jkW
duQcyWOJQMnGELsz3EZs4gwNWCe/8tjB8V7+EBaS0le8P3KBkJd7WyGSTnwY
ygPoDJKa/fqGyuqnspG+0UmwSqFKTGbTmHm2rPIxKtsGhOaqAK/gOjsmksKM
TTQz8F/qVVCmPwydtQQQpHkELu8W3BP7E7hRAFpyJc63L1Zs7xINgr8rRsn3
z7aXJDjuxhlOPqYVjno9usRW5DvNeeib4avwDZJSBgVYVLxUJqMFWdrOlQ9p
mXkyAPo7DfNS560gyKrBJ0f6/WtyjUcX3W+oYktlG1XbkcQJhdLW425TC0TC
jqM/Zfp/KRlMZatfTFaz9chg+yyN1MHw8qWSepl+02u4V6Y+b6nLKHFkVSgQ
42LyKYmOvXUDyKcuf+B9zwZRaOZSuzdRJjFOOFu5oa3RhGZHUgTw++hMmluF
x0dX0WPUch0vemN7PHcyjQ1ecjnmPfyHUC+i/YbCLgviHSqiGYsIwgtWnSoL
PKYBY8VLpNrh+TCW6LSa6awPmZiEQ2pXpMBOYKBqW78Ah9wDkQol63sWXvy3
LK5Mx2aMbrhGT+Ia5Oa+xbC2Mr8upMJwtPAgfMUYWHqn2CbtPmnqGclJnL+U
52IC7i7SLaQVF//flWNurXgSiYu6bu3eXh9ftpkI0yakuvuKrxcduC7tlxWo
gWBUM1bqGKbTlDoTyADjOapBla/IlmqT4g8LmJWgPvlFKWsRGAoWhDmS4t5O
oinbqTyFfWYgli4OaqIrFYXXGsacRe7Rw3B4DhqRFPoGkWs7MKzIKJotNW+S
lVS52NQEW0Iaxh3XGYuyzXERhq5mbk1znM1mIthc8zQE7gGVxXvLXKFodDmd
D8xIeR0qaU8UKBJiFc+gRmagZN8pNkvVtA0ibHMPGCxD31AGH+ASpO5k8mq6
IuTknzngiGv+fobvW0WqCMJh0vxt1E/kL45dwZ6s6oaNxdUXf8UfIMLi3rY5
o7+t+kM7Rfrk46xn+utdn4pd/U1+ayyVrYJtHMBKKrsBw6OuuXO9nvHP+H52
CW8vJt3Z/1X9on9m7lBTUITH7fLFWK/T1sYfrEQvaoG7UETaxshkb8sJOQit
4lZIAodGzJdA3sQZl0jax0oY2zY3LejwrT+2HEaEiER7WcbRVkAuAocCt7OK
VI8qjsRidItMzqzG0QabdevJ+ks/F3v+I8N3g06pRkBSzSzIPO6I5jB8AxC3
wQ0pUy6wJ0S/T3hOnBzSbJ06MvC1RILTwSVkMiaOTUZtFKsJ0f2p/VbiCqu0
203ccZ181Xo3HRAqiIcmUOoVsLmbQ5EF1t5dOiuAY4MrDQL0WprZfgfSopNj
T79MmhXEiCS8fLop+5bZYbCmmyUV1yzsBOxGbXOJ2IJK/l0iKoH68uP06ppd
Ai6xlWrWmpzwxVYznTUYzbBM8yM3wplSHXF/LZ8abY4AeNptrcZouveCQ1Kr
2wJGlc3hD98NVoWOgE6Pq7qxhw4ZDNY4hDMmr4cqOBZXsL7MzxZ4EMnv3hqS
XDi2wlEINZrZADlOtOHBFUoJ6aKav6apXfcW5TVPOWaknu95OC3aXhSSKMui
/P0AHpcwTTgpS3mJ2Z9TBLbyCDVNkIAbc6ryURTlBS1A7j3iF/0XNCYot6PZ
jyLWe/JpVfVryKdYVXyxzf4Rbohf4w9r12nfNZDvMqDiG9RedfHzhF8PQfbe
FzdqaUcaqYRUBWr4cFOayMWayNICmNqe2QF3CJXT0lSdsAYsgJTaijh5ACEq
Sq3xLxl7s3YW7c4YHWL0r67PfIRgnMSJrjfZBNPTRQO6CRN7E1MzFPL276g1
wFVe2SKFQwMzZX5tjznT+QvT2CsMBqnr5wQKNyiltxkhIgXM8K/CLYhbhrJW
1R77kiB4FB9JhI29HK+bTn40JbB9GhUPVYbRSE6xA/E9mE0kUM3gey9PWJ8S
dgHVRTVZ1q7bHnR8VgRLHCptGeldHoLrIkJagrOREEylmQb57OM/u5HpmIjn
4FPF0GLhWClFxv9xJrqBG8r8/PZvK+qU3IMYUA67ak5GAOAOqGUQgSp49oWR
WwfLeMYrofut326hMyBH6ruBG08mN0mkoubSA3+ZczRPkAS9U4m7vVk/0zvW
EabZR6BKObBkIL6wzdGm3H3jC0LR5W6MKX2gMZZ1YSWM0fcluT9JJ9PUWpwy
Da7L4jzA2+YMQBq3ItrIBsh/bqQ7pfTbtpvEKoA4/bDJjLjhRwDAv0krbDzP
YuaOvqFgW1w9Hzlbvd4BGQghmB+kb2NqMzCaXSFav6sSSCcFL2xhzKVXT51W
fPFBUAsMCP/sK7/BrOTbi4o7YVui1sI4cd+4ho1HQsmypwAcvnlW7pIWSC+q
DV+8cg3DCDED37HnDHvH9RrAW+0mjmGLPbpKRCC1Ulc7U81+7fEIY2hgvesT
SeTFDtlzNAU575ES4FC//mDjvqSY1KsI8sxVWQZvIAvT4xhokOUuTjw/0Hxm
tpiwuZJ9zgqUBfKElssScoRmdn6FkpDx07xGyB6I9n2rDPMxQT0DtvW95pms
gQ1+Nfbc9wtZ7Jd8bxLSm1AAqWvej5kla6z1zXfmHlv+79BBvSRA6j7VdJm6
mW+9ciCZG+x6YHMdCpew2CgSLIO76zbqO9iLrnpGfctrQEmPAw5iacw8p3Fu
Hpsl5VHDcyaFVJDIW96MdxsvchnbEcuBOGnUIF5ozNqqpKVq9GVkYTHsDCYQ
HLpyCeZbKA5tSDcqHant9adRO2bAdSNWZfb9nzeKja9fpR7ZTl8xbbjPyOe9
h8ur2YizzXoYX+xhKoWVCh6z8PS4gh5RsYg0G6rou7w34ABcfi24KlYtw4g5
CkvAVnJcjE2Q4ZVJc90GHOnjSqzB3GucJ3ITZCga1SKsOfmdvLL1GXJ6+vjz
cGSjsWXMnKvOgr5z49gNPgnCjU/lKi/0CxnGaqPBKdZJLOCxZpgLnpyj3b7N
wWuowM20synPr7FZUbR/upr7OqRGhdeQuBQ5j7nu9RyWoD+2q+GEWmWRoGEe
woEWHlFEUbhx0IUtDI/lp1dAuowDiXzj5lvH+vt79hZdz1peBrni5GxtjpkP
tMLznEvbQQPw+Rb8d+NprC9gxviS4Sce7M5rnnGmm2CjWMI03THqFHtkQHHE
W3LySgC/a24KE9Pd8ZcSwTl44YcDdyvrNFTInD/ChExPD2Bf/ZuWOH+B5Hdp
96YyR9amSOmFPW7JynBvzdIhLUhfVGOfVYitLCGqacs+0c7wnpK3d110l3Fw
Rc7HsSBfwfe1CjFcLf0eDqK7YJhkIkRk3xqYVHhOTKyKpi1y/jB+nDKApMgN
KlWbSQG9WIxziMZAJD+qGGtJ7Rt2KaqT9ZsdFYKibI6Tp0WC5SR4rJ5TakIQ
oUFTQ5Xt1R3HDrYuZR6zwadqS2bjVQibY7MuWi5yvGuOlm6DX9ikJvjifT6b
xKkWCMvwJ8ILYl3P3SygGUNjsZn+px36RZEoLr5LQsBlEOb5gjbqA7kopfwu
WC0HbaBU+CA5yCHO/PioAf8o1zCENa7rTcPOc5ENjYJwJ9UvoZn7MROJhYx4
SfXgF6pX1NSALmF8ZwBSCAXh0/y5Xojb7K8huKQtySN/xHAq2eGTHM2+2zBI
ytaqC5mRYzpwdX8GplC9Y3R0+G64TEFOsRQyueQkl5eQcZ1H1TYQWKiB1EzA
YFipxqn/24gdRb5VDfJqz7RVQxKe6Kiy+yMJjSid06/eb/Uku0N3pf4+GUV9
X5FzVvKSa4JSyPnffqzjWoD2TULWUh90SvVTWjWwHthqiYUVNC+rBypf4aVo
Wjh9Kgw6gS2LT+nI68ruNuOEmM+x9vc/DoIv+2CBFWgMTpnbSZgMF1F9vUa3
osij4JNpj7+Y95ql/cJS1D/aq2+SDpPjPe0rNuav3CYnGXov1iH5vAQEXHVD
fm2FJXnNU2k0WpczP8hP8Sg9JgDr+TCodiP5E8Lh2xvMM6UTkwZI4ZNcUc2I
3fGzOiGLjsOJAb82pEA5U7Wo+KFmcnLG9rB3pASjavC5ORPR8+ARLHM8FC5E
YyguJye+oZIhdf59xCI3+VANOgD4e4CHfBRxTwZQg4tHbHeEFu79lcR3tsMf
H1oTgV5RsIh7l2hqpiPRKjUhSjOSSJdRfsg5rcObzIjV36pUyqDxTi5tbZLF
6qS0RNWO6mlnjuTPqGwO1by8mUNNskr8iV/3rN8OFO0YzUCK+1qoG5LrpVeJ
l9mY1UE6oVOQgBysV8p9YttKEWXt4cJ71Vd/cZbVWk/qpxqWAimRRLC/L8qR
RXzq3YKyto9rEdK/vlwKR81O5x0+yLe3zJrP15fgDSLPt3PGkdQ5hRQRoujs
mumSk1qxs1PLyMr67qUFHfwUF65/piNXr7Z//hE69mmkk3pfYpz9205KAyQN
HgvcZNxnH3moFLiBIo9DRcQH7h+AGDKOwNgQTdHiKQ8k4UlKVMG6lmkDVc/p
NrHEZk/qj16F9QKl8Lci4fFBiZO3+cWjpWqdxgZtB2KzSY1ePT6rOUnXfOBj
xiT5IAesMeR9/BIs3vsJsdnZAs76IbSAGvbxGKMyBlhsyJy/d4GNtTECe2OX
aMOyrtl0XW/7rZkLnLB1lZchJnIWTwnETAx/sEd+Awgv+bPqMe1taPxcbT7k
oU4OBjnXiN8/ySc5I6LDHjkDz9Z3DhHKd4cnZm7/R9aRbeK9aWXuX6hy9LGX
QTXb304jHdXOIqm7PPj8uUJxQRxYyGMe1YGxJIWXHr51HDTHtAAbmdmhRgWA
ceT6fJHD1qWrpi5DsELz0JI9VwmvnhqNfLC9vsSSnRZuX9ID/kC+o9HwKr6D
s9f5k4ByCM6Hs6TL8KZ6GfiwJCSiXBjDte+RQ1FQRwTzzZLTfw1fZrH3bAKJ
zMV6uWgCu2r2HGgoz0xfbvd/SYTqIc6Ds4hmGC1YBczPqvi84ZVm3SVWSBQO
l+afC0B+MEYC5xLdCbp8K6CBGHA6yMTwdEhxZ7lHRAiqS+ayKhcQLuFSBqbg
mwErO6LexC2kN3TOQ2S5iLMVQlptk/Oam9lVFgCM1YAJ0Rwuf/tvduNJZDxH
ZasZyjXdYixKgOOdFJzeAjS66LBLwsPDMJf2OisikRX8j3P4fzp2RY/sj7+d
lb0IYuqGo7rFfbUn8GCF1lfu5SDE0ODKzA6k3A6+w43x1FG7a3V6HHFU9vA6
gAYgrcoYKV4A8DibxT6hTDDgIgNJEG1/WSfgmJF7jGvTEHO0ss+X9SMxjjux
eHhpv/v2RGLLRSwNz/jcUoIR5oxHgyvbfzHTZYzUWnp+Ezh0c0gwhUN2Ntit
P6GrCU4Ct3HB3IGUss0E2jJcim/O3xN9OK54lNSbzU2SWaOK/FuR4DjUszVc
H1gIl7CTtwBpy0dthJwM39UdLnOlbTx2Ai6/qr4sikkSi91iWmrxk1BJfk3q
FGdA7YPOc2jNqjutkeeck079eI2EtfMWgPd9fcAqwmW5l5t7hXHppmOvbaOl
s2Lt3lUoxHpnWU4JB6Nd9zribvQ/+gI8bg+Wq9mc9wzsjFTb4POBJfiABM2G
ajWIHbEsoInZ/+YMtk5AmK1hty5+F6nGAOpPsHH4HzE+3lg1gD6xv5/X/wOU
ygMnKbFt3b5k7BVomNG8EIIuN89PR/TqRWaFTxYC5F1DCfAJd4tc+F3uxZIw
2RsTJpOA8O1wz0DSsUarGm4FGp2uS/boVJRL+u0S2+V8E1s69h6FY4fAyg2G
YTfjz5qFHZ+GDTJnjEXRnkMXcmDAoKepha9oJQnWAL8vSn8qEDO8tOj3YKIu
9KSVyRnAoNWkamrJgxoubs0MDRPar2EYfN5S0WkUUWKhglVTIMpOdf8dIQ7E
wHeQsI2CUQSlpGoaIieSl+2UbyUHZKNpJ5Ez8yxX1mC5GwLij8gqsGo+ed2s
BEiTOvH4AKISXAaUu8nSQK/LFwjMDgGl+vz7/N/5qooEDT06sCuk8cTOJF7k
5GXJWNeGUZqIkAvfnq10lXhrPPQyst8JBvizLxdBLFXWhJe1TfGdF7d48xjN
YSL35/UZIhaUuk+grqDUBfjXuEfRp1ZFCxoQQoX6xk46lyRiERI7KxM2m7rj
s8wayNZtP3j1q3TXe5X3Wel7EtU1xb4nl6x5TdPVcjB6kVeLrtPxv/8DmNiw
f5VaDFSaAIQkwRS2l7MoxRgj6vmpMXHN1fgGKlMhcvlymOz3ns+dVvyKTsEA
uvy4y/gvbjMOln6EGXTl19tL+fZ8KD8UG1FiWGj23Drk0pfSQmKlbDprW+lB
U0ssHs57e4dsqtahcPBY/LtmUQal0Qsv9LQJv1wJV+7IE+HavXbYa8RN6Iyv
hsaDpQASeRnxxScqrQ83B+EBhomNlj+hAJ4GbdLI7lEpgzybRaqBw+uXjR78
9oykb5UFlLkHNy5YX6tm9CFD1KkjXRD3kFrY2W8I6yz8t3OsbNn7/UzdLNBF
AcqqFBBxQM0V0b7z8meLwsWeKKC5ZGpw/Mmogkz+zPj6e4SCLFqS5bSl/g7n
TdCXq91adQl6u0HKUsMDkToFlouAUUtQg17mm8hq2Lmt9Juf1mzAGNjcuPAD
iUiWUeoz/xnmaB1/PcS2bnJ34DfA8rP/D/FnYmzzJNovUd9uuEKbCqh2beRf
Q1Qt4G4zynoTfHyi9IBRV9PmikmyraJnD/Oi8UmgiiGOWCjcCPir9Lmm6+nZ
NfWMSY1A27TBelK70TM+TnSmRMSAogSEodDO4EyHuK2As++sXEsqWstY7a9e
CDic/bdOfN5Gm0gSr3e+YlzVkinhSXcyCExE61d+ggeVaWOjeW9pXn/iECJe
RYVyH0hj9r9eTprJYxG/DXvOEXs3gx6CQeiyNVejreD1ubBCe+OonCKR1ZES
9roZkuHT7C9pwxPwmeUmy00UP7ueL2aJVhi9OFJwAaP6k/7MYsCAwsN2dD4+
eMPhOhyPo2uStAoyubQnm2CiPMJ6faz1QrvgiBB5OcTPppLLzjGLyd/EYdpq
nQD0PI0RKlIEOWgulX07amHyXRcJ2G9WosIybdfka9o/2al+MEqlf7mfElds
vK0HJ/3pU7doMtk44vtGWSGiB7q9gq8pKbJkU01MjB03OaYals4o5JjoXvdi
DUTs7/TkTtUeCvcBN247ydtIhS2Ide97TeZTqe0mEo31Jhbo5kD7cf6BK5Xk
nfqhhOmTri7/0dqEIqAtMopYELtXCePP7OwdiYCkX9wP2nYeup2DXecHjGlF
3zCt+Q9dEaOvs+I7tiUO4bfQ67rTxGVYk0lOLZmnQx75zW++cz0RvQRXG1gV
nPDRhvMkrsaA9cj69R2uHsk/GQukhDqLD7QKBXIBapqP28YMSYOfCn3Z3ucA
6Tu03M17cI70BcDSyK9WVvkw2RXRs8dw/CYjr//IfVU7LsK9xhHaPsfWC5IF
7TzyNo1mSsD3EEL1965EPycGaG0ieRsNrY818n9AVdJSSZumBJznUxwrNhj2
eheK2T3nBO4maPcRq0yRFqC614/IRW1depm7ehvsVxvvKDErHOKO+gcLLfOe
tn0o5IK2FBl6F0lyfE6PCo1nL5q4JXEnOfbnHnIM7NbMdP+MrMSi79AaDiGd
Dkge/sy5VJdp5Q0lFXQjFjZAPdwAsQFxHmmkb0AtZSu7cvpsGcmxGKdGzFbF
Y8mhs64wR8eEtG4ve/fA5DqkN5EJKfFaAWiC9anFHt1TcxObfGGC/Z8L3jt0
hASSmypYY+7WpDD4hBUauQgRq8XBwg48HF/RC9DU5fZ9rovjTwooeHRYBl9C
kLXGctkGSiDMUwIvCqQIMAwNpb2KDNkv37oa2zn4dn2Y4Lgh8A/C8DPmPtF0
ttHh8hdKJugkZcIn3IY+rjzjRfrJGtFG0PTf8ohAJGlcDsbdE0VJKldLZkis
KQ6zJZnx7KCT5T/L5wjLczjnyPandH62xBLmEtDOqhS7GJ3KD1i0gBlibYlU
JHSK21LLRoPRWObrNU+ukoFoGcHdjYhDykMbqA9difJZQU3e1bYmSUkCYwk2
RMlB0f1DreYXl06GkpfdJVwYtGJwEV18L2KTNFzNmHEKj4R/aPT6tUmQSrnC
2NJ2TnquPLzI8EcO3Mf4Oko5ev6mDpb+Gw6vfJRghum9WrE/qJfQTYmKTszn
nQEvdZbNXU2dFdvubxTFF4HHrgZXseWOHOUtwcB5+mfaoCRE0cLswIKssIni
uQNI6+mquOdwD1iv2zO2DaQT4cbQH40ttIZAABKxP+kzeAI+3zFYVxXlOCmN
Ras1YI0PZhLFCDFdQfw5PwbVzVW9GUgdZAItJqEZjX4E7rlx0uEIt3/FwVZo
xYgKYrOyS+Wj4QNNkSDW4PHa21fduSVSQ8INjHLyb6+juGJ5nLZMAFtQCSYi
7BpO7+gUuUCmGA3auMG1Ky/OVvH9f7/4jToBA+Pvx6rmhSj/hZ/KwezljTTU
LWEWnJ+54goMNHTaldEcy39RNrRRiOwoQVWI/atazgglNXAK5tY9T5X8ov3n
nes58QQR2KwMxh39tkGH1eXLe7QXxEIlWHYvmcsVA6Srmtv+I+rZgGbmjiPf
IRkhBqlWiXoe44b9QiWuUUJQ/a9StOKyEc+kQdt9Jetf/BLRohHPqxNvg/tX
ocJ9t4fcUQiIJtCnH6tSjB5RzHFdRHVBE6YobnnzQab/a7b8EZdXPE2ivQlk
/1r3ZS+CYP3pZaAhVUJpaNReKCRjX195QkS8ptp9D8T0gfjncHaZig6UiQPj
mD6AGpx/mHsK68Lv4CY31TlJkedn9T6IJm1wHVxh5W1382PXCH12UfwZJHup
xickk3YcSJLfsSTuGJBAgKewXivlv7du7SVBh5cPjG3mG3LfQS8RjDWPynR0
QfuHv+gCg/6UXqab/HlGGYiwjj2T/zCditOW8bXycckyPfiKW1/n0+3yrr8+
AHWR1MhHUZN1PrBVl+WJUEKbNmexz+p5tmG9DaQ30jDx74XlxNEUIUiEA1HH
bPK+lltLfjD5equxseXFQTxc54PU2ASaPywPLGovW85wLlQFZP52KkqZNFxV
t4l4NZQ5qoQX/1fTarQkghp6jhALebFfYv/36axIuBd9HuG+/R7ESSwZCus4
z3mipmBskUmmts8Mh/E/uOQCPV5WV+jtxpyvc6TpIyBhSKs7NscQhwzOPzhG
7+AbprC9eN3o9m6DxeeDSis6TlppioQ4Csjel2p4Grzoo9j74C6p3D1GcT7e
SYhj04tKrQjyam19Qo145esGT/+JuNHTNHnYRLYLeAmet9RvYp6Eu2W/n45S
j3ZdYGi8QZ2hhM2e60Ddz8fUK+kgXQ6rE+1IWKYfJXAYWdlFvai9pm4+NcCB
WBLZUPHWCwKxOP9wb2UJaN/XS2TzymLAcwSGHrSoIzF46pdManE0Wwv2mp84
jpemRgM9ZXEoa9T0e4UTzq/Rh6s8FiYThpsaUh/FGTz6dYgYrX0Lp6pHXrcr
+fIDUfb8Vd39lPpUIn0+4uDIkvc6Nnw24CQrhyD9xADr8xGy6fP2QTvxXNhi
m7bagxiaFlqVPVBQ4DYyKgvr/Yw2rvqbC+4K2cQJzpm92idtP3888VpmXjq+
WoHmd7WUXwoZs4q5ZXFD11AmaAHVY1SL5HZtFDuVJvvOoqKf6cuIzPOKEO5W
t8pu+sFty6gN7h7fxQqbb3JYn6N+DVU6fKCENonswLONlztiu26ScSweIZ7C
x8zTMpTmBgDrgsJZI8usThYJ3WhzqrDUApWTY9vfvQGs8ESuIXa3eSfwvw9i
f+psO8CEevOyY/7QA/FSbeEoKXohLSdQkDBKEmuWWkAtnr/P0SoaqbVBy6Fl
uM+Y9JlD1hEgx4l5HDmrnsrCLwX5bGTELg0i/GSC9a2JoTTrHfGQyj6kjq4V
drPYke4IeF2j/gPwDwzMZHbWsF092xmoE/MVqglAq7b4KxuaowVgetEOCYUp
9SlUEt5X2HqdpOPuPHqOuENXDpZfgr62AApJxUJxphrfojO45best73zm6RH
r+CzfS40Xwfv1VKhMddlGYRyL+daV82AmB3z1D85sToofx23fqpI4SKtd6x0
3AkV5VRaKGYPjrpiH6MH1Mo9OHH5jJtzdcA7CnnuCOnn0sZFGXUhTik69v2L
VpQwRo9QfyF9LFS1spX88lyRYmI02sR7pBAS+CJI1Q2iuxpQ4wk6y5Yl4qoP
KapFbaHVsKT4TTZvtTOI4ziz9zd+DE5X9tTH8hN1E4Gzvg0dudCrPwnxYazp
YUnmiVWfyq4upaPq2pAVjSXssFLN+1j8zqCKfcWenbtbox7mOuzgkqFdmESI
oJupK6lSsnMLy3UcJu27QnZhKIT0L1As09F4HWEWHeZgkRTWL43lxUiJAJHV
BFsQksKuUspV3r8uatMDtWYAJyqJcbQ8fjUep96VnIUZCOUfX7KRSqAUVQFR
oummduhHpan8hFlvP6pu/FKc0H4Ijw79peltfEe33pEoFRHHI80bOjEbF//g
DClAi3rPzCehPzIcqJ/bU2NsYzt2TAuzB2QEd4B31nkSmQ6NqydhRm+wPsL/
+LaKAh/9GxQhZmN7yB1qtJhb64wYDtCSjHq4fAmLq551GX6NuV9Iv3Tn2tpc
oqNvSnqJtNxYk5LU5tXW8IjpTIFR+2I5I3RIhImsswp1C7fGPIL3J5tZoOT5
vK3D9xf2d7Oic05enHrYXwaYNT0r+h+HW0l2S1mbTGWaPnncY78m12Tgxop0
Rp9z0zhWLRvqG86bqSpHsNmlmKW2U0PipevcDDUd/pFuf+mvLL+8c2BdVqc6
E82mVBGMf3YH5paLAaYhOcHCO9d5WB8XemqAcUst4rTA4FKmOfidzDRYyGmY
VhbKevBKskwg7BGdX7ERGCmhncgmXFAV8E/C2174f7pMaqHJUTnlXaRcgHsj
UsDG1QNx3V/R3o+uHBBmJ9TNlDM0fXWvRBG5xRFEbCiSvoCeAiLDegP1tElz
tgzkJ8R/BVsIMWwJ7x4dU21B6naCCXvJnTlL9ToiQWLew6AHr7TNmlt2BW5i
gGuJiJ3H9ZifGTz+1+wJypK2XZ+vJ7l9HWzdlLgaUA+v1gVlXCyoj5pFu+WY
yb1GPVimTmL76QRSw0tpGykejgBdtWb6L+VAMQCF9PBlC+od66BEmt43P0HH
et5lmIFWnLfDNNDnVCSq7AQbjK8121eaRxlvZfg/RfC72K5ItkpAitlhwpe6
GY1w7d/9X8oTsuqXiF4+EPk6y1hhvqfmY3hco0OSU4p2+er8M+45zKFwPSJM
u5OvSkcf/8lMhbxPGycLAMQh00WWdJF3omhd1/KusZf3tUamMpx+QY/gmVPP
CZN35Q89Sz0JvjQq73mbMHHDHjdV38XQV1z7Io01ZZyRMeo0iGgyIKvR+o5V
vnD+v9JTi+O/zwFHuVXv6aiX7U4ijvH9+jcSgVzLWp8OZjKKbfO/7Y1z6ay5
WO81yZlcy8xk8OayTYT5T6nIQzqHdiFu4JKhIHcqKc2657vTUF6yLQm1ZAFD
+fJVcapjbfXGjVSrsgBbiRBeIuqlYrghaAuNZFJvHzRg7yOGWZsvNte/oYKk
8hnxuUY8O+c3qbWhMSKmG0DIzdLZG/2baJW/Nt0C4FpAbVbm91RP9eky2gA9
h/URa8bUcRI3T4DfnivMVMGJQFZYzByzq+3byVReNMYIWB6cbKc7m0uiT56x
PgCQIzqkoAgkAcqxojyTNEe5QOo4HVmEhqRIdMjqmJ3Qq/mUU3FPbj9F1tb3
Q/WbuBb3dm2zDlZHTvkMn24yibquDD5L/YAOjpAWxQr0YUuuHAqDMAEFqv7b
X6EqgmDg7KiS/OEDHFoXrSNA8UuIpu84qv1DJijStbsZIG0HBftw122armsY
ASHhQozBbUdT1QTEUKDKkMafilbPyDVDbuSjj0/yD8rJpP6xCBF3yc2sklgN
iQWIRIZmPfaCylAQX5GBCQZ3RD9W3LTI7OF3mL6DHRv43uuaf22/YdZjoVXA
Cq4/vixaCuWGUAeoKWUEiMdIIHb6ZXOggDdEvehy0BX2X2hufZ8v4qKnpPFS
8d6AcOtcuryFZmH9b0ZjYYFbTUoKOec4og7V15wkR0fsI8oiIpEIe6uT+pcc
BmJDvmCPElhIosjkeDrGN9y6pdXRn9l8e/1Fs9UvCTJ0MSHMLsqjeJ1rQrYy
mpMEjb1SV38DuCPwXQ8AQ/KBxf63M3Yc3fJ66ZZMrAJrXkShOuUhC99Lvw8k
K5RQJn/rQOhDuSrUfywm2DFBJDJuQ9apQBGZn6b4QcHysdkpyOdBbsdsf5r0
dfjXmES0YWoV5G0HvxTDGIKG6tNXwRouFEhCjK6R8EtM4QdKAZuIpDxO7LM5
JfTMX4gbxRWi6LvBCkuVEjNL7ssaaJVrpdpBdhBMRt2ZAPQ2aitEs+hK+y+Z
zALAGtDjdJ62mVCnXsXGlCd0ac/9kUYV/dY7EuMUiS0ZR3p5toZzBGhdH/qS
0agQ1P0fmi5p4Bdah7RQH/Ji+Nf6oTA7UORiAKD6cC6Psz/mQxg7a+18CHbn
KHDI8rrIHUyOo/i63EoUef56Hv53VqP1uO7ywVFaAB4lU/3bRMwCmWNh1bBr
OzGVxcfg2jIE23U/hyHRscTHsK63sDORter+83I1l6T1wmoagHn3r+nqCjO1
pYdwFAZ04rifCM5KYtD6H6ROPbAfmE+XO+SoPy6oaS671ySVGim1Keunq/fm
3NIJa79f3A5o0rxpCR22zr9n1pIAR18Hlf9MUkh51e9PtLSoDbZArz/E0kMe
/n6i0k6VNTCObco6elcuQFRSlckFWsCu4djyK+SCvyY7ztILDoBfyednZqDW
Dwks5k69uKwB+YJu/1bT+7i2d4JogCvSTTPnymSbTPxBhIvG1u91GGSmxwmq
2KPGtRPsKNLspnZCJC/2H+E5ouTZBwxEBuSYS/6DRg+DJcQwyA2LjpD6JwJP
eEvKLU9LDDmMckm8RvZ2RIsCd6zvMwPeJwUHiGG7UBaQm09ksxFhc3YMgNau
lH1PVnxOSetLvM4XmesCUvli37DJQ2PmYv77Zzk7+XXy8gv2rzxtikbUwfaH
5XTT5WYdqBCTFyd8avIOAkWpmW291KWtPnibGxWnazUYVMVauQab6tYsnOfc
OwG5RKzFYWDucPKOBNJ1FeddeBOpHu8uKR2F0+EtX/Mx0+J3pg/gzFJtnABb
PzHp6YDUdMI1ju1Gm8taix/J17LQ8hP7hQUg0mOrSXZATFXSXMWaiEHvzOen
l/e7Pp5ZBCdl7JXRmFI6jsglAZDpRx35z+8+ao+PVwa2VKgJOvUtCOmvAtxL
gP2ztzYYyWA/6L5HekFPCqNMHOtUTHtwL8F0eTdLzoF2IaMiPMTLjVciTXJy
AtCQWkAvJ6iE1ln/JxVpe3vSgcQDSXcCQEH8WVehvoPlCutSKN9yX5ZnhRWg
3uZwkVIHSLp2ZIKFxd5EFpT3sANOrPTl4z+sRYZJ2Y93ODMqTUjj9WB5277K
MrJ21M6YD/IjhwlFjU3v0IGXFNa1hCgG8uGT38ztfJetZG43Y3lGvtWPLcB5
p/lIfWNc09H1QCOazKCqBn2EZT1DEPoNzFDkY315nOEdWdsoFpV9QX7oAgSu
kgGQd6PfsQNL6skeEG/f4HXHBwyINJHCcZRGBUJ/3kG1pVro9e1i1vU/yrb1
F+asae77z1M5CkoMa8aRNWlQbMsxO8UdAN5ksLT77dPSEMANDJEtasRNNAPO
fx7GJfP9fu/2a+H7cmoHy3gOTlNeOeSahE8HsnQpulJ2Vd5q24VrJEd6EdXS
XZ84Qu0ASdqKGgDczrts3i0rB1kpSW811mmiaA/V5fLQsmbT42Cm6VcrtLOQ
cSE1U1gsRyj54u/1rt5DmwLn6si1AOvkFcyUaI7xL+sd3yG5FTZYWDAXewsY
1mm1HPCoMn+D99djm8N1GaktOdN+yfPy2pk9IHc0lM3aMM1m7oe+71UFS3OE
WYwsdz8QGLE1m8kLIMGQNexd5Zvvt3R37IFjg5BgFAnDUfrplcFtZMAEvSvP
CaeeGeJAz/96/K8JpRkDY2BNLf3EBKHXQTQGpwitQD/rpxX1KZiZbaAhkgj+
NQZnSBRhdHlH6Ig1q7jVqIyWjRzs8/6GrBUDFyabrQbpGHme6F97Sm/Z9b2u
7N0Yr9/4JXV6FBPf5cqrCilNNcxmvCbU51EPXNRQ7+61DiGTkOSZ7fImNaLa
IJFjBAHCR+sEkDz0XOKcRN0k7UzcRINTwq2Z6Df95soUEWZjBW5/fT3Tcp3L
g+iDVn/t2HFq5M6KcFI3FLeiyl5i5zB7/UYLz0Dvy0CbnBRiXe4LqyxcX5XU
B3kYwcKutSjksQCy9xEifeK377jDo+dpUoDpO16+qbP5qxDTgq/U5WaVMU45
56+EFzbTa/R0AdSUgvXJPog/hEKTUVy4Clmpzdj5p6k2JnwtPM1fyl3I9vfw
CIo2pi6mqVgwZafhu9BoEiU0IGj0lOHL1OJMBoOonY40ZGLO+3hzY2vP20O1
XoHxy0ZcI0XEMyoGRH42Z+rnwiSOH09sDaqreAmuHUZUv5edEwI1S5Y4/h/9
GW32xyX6q9Q4IlvL9oLX2YYacoHPKphcm8/DF5L8rANC0P9Yl/0QARDWXyOj
yCAXHAgSpVSRQgU8mvnoh9pRETx4nayaodwJG6PXiF4OiAyDtNXEzoenfue3
RNyuco+y3LZXLQmZrYK1Qci59z3VuiD4QtGDH8dz7Zs7GP2Nx5KUf1g2uAZ3
tyZuVJKrx/Llif7zwuN4twPrtKBPoU9Xss14car3vd6Acx6fePlePHI65KsS
LtVetMJeDyPQForGFZbP4dYCmtQxOtjw5NNK4//9LxRwSsGMcLbgD7Sg6zJn
ln+OXoaI7pQDb2ABDkeDvOa/04TA28Up1vhUkamXtdStbWnotMpvr2gMIc30
Y31gUH/FJAVSq0hwIKLi84G4GcvzPbfEzD4XVbGaY4G+f9wcMH+wMT4fypDP
M5j1yjBaX9mAGUHtfZZVDf7t1/tnw8ERqk7GkmEiK2uFEOR2MR4hkF0W5OPa
vumCfga7ulbdyNOh3cN2Iu6B4FzzMUsP6aFD+uwzaB6wwf8dn1fYWzu8K+Fm
gPgmVzdytjUUhxEO7u7tx/fgnb8cAvXAE6yLXGJOj4YVUgKCGl2GbzZzq+oz
X1wS0Asp4EQo7xCcXAgP77/CZBuCO+5jVNjLulNCLk8C5BqoiKxaCSj5ILgj
5SM6a8oaL8rWHkwdxi1eN7FsbQi8VViqVGczR6Zr8ZROBDvU4G3WzUNcZfmx
MjThYekjAtiZmP6SGI3igmrDRjY8naHqYxpOmviGQGI0ASt7Ug4vgyvtQuki
e0j8W24IN47f6loeUrPlfQ3jdJfoaJBwn8cr2VVQj1X6HuTTBgMuuSjSBpFU
iHVRzv+46zqFsBtPNL3Uf5zfGK6wOvND70Tsz70/QuFv3NZPQ7XbmQObFS6R
JYCm7UnKZuzP83NVd/qfAuZTjyekioebm1P6xVej7P67i1Oe9zUAeuFRXs3P
B191NqBRvssTbF5tn+r6uwZe80C8PEAV3kvGqzIdLFlEmKePzctfXVGUovvg
G1ZVZZXZLhDTwNbox4DElfsIIfUSNgBNMDRIAgIkkdcraBlLFfwBtjrT2a34
zu9V877kDXxhhXof1xUBS84UApr2nxO2UJ/K+CBWlYn1UMrmKBu/KlLv8jQH
xIQjgdctRiw/krh5QSh9KKNW5O+V6pg+IypM4Y4rYX/SEhODra1D1QWDttst
4y9mqBJHxpBBcYIfmPSMD6Tx24Fom7N27/TdtzIKG8aemcWuat1biKRACupb
gPkv97wdE75km33Tc2mZaeADU32rQYVt3xnmn1vENscR0rAwsHJ45wZe9qQV
A8ZCJb9891/bTgNTi7eX5f11DKPO4rmGznBtA3J2yEwicdr3rk3UC0tn1Zja
oHA0my3e0RrHOvr8Ya1vH7fvSq50k/5nwNWP0Za4UWEuRgR2ID+wfefjcEDe
FqReJ7T1AjbOh+/b1TldeEoDFE28wsF8VdWBDRz+NyMGtxwr4K7jfnCHB3pi
q7zejGyfl4Y4yjD5YgHU9fk6SiAYEg+MlFIiu7bLzWI2IowXNfX2FmvcLVBD
ES/YC9bkJmifmFyQA+UNukuWxlikQ8mu9BJ2N6qmTLJRSpmy2nJhRMczarD9
eFJguHbCufocdF3Zv95YZ5Mm6DfI62caYGmAocHyYql3JPVfJMU//+8K35ok
uv5SxiZoeR8M89GxgTmxStAno++Ce5pOgWaa6rkbInSEcnaybpVW3dEHJpfj
cVTMXTKQ1RsL0ewSutlGomkS4fVDfAwrelFzo3lq1E8TSO9up6pUgedjY7+U
o6C3ethiyymzxkYLSf4BZqZXa1NOegUA38wZA99c6SrEIp68WITjc8LfGCB3
DROQxRiozciYLPYdeJGqBEaRBk1eXEtIh2nDHc6mPj2b4NQ2FCqSogDruJl0
35AMm8dDmZva2mV9IW/alnD6iSRb35Y4yPpiFz8KMy8d3kSkhJhCKNrUkT7R
uREiOh0D2iiCNjkxULrQbK/UhBask1tHQqzVweNkfFHwCOcmYf8zGHSreLc+
4xVBdQ7knPTnRzVfayWFcNHH3Glwx232+y06bqcO5j4Ov4IXW6FX88kRUoR3
kbr/65CSGXv5Ybxkq1smXXo08mGpOP2Nk5qDN5GehorwTj21xStNUiMK76Fg
0he/U3IHKtELfjy3BDlj7c8Pp7guq59TxW8CIqCxfhJtBWFJRXwPGpBPftyd
Hd5JHAA/QiUrrXcT2jocy7HjM0xdaxUXyosV3HJJFaIDqQmYFm6GUKlh6CkG
3+jeWOmgRKWL/0ofh4r4kQXjDph59mqJsHMznxaMrEiO8J0E/AFtd2WQPmg7
J2SpUDqjfIAUx2a12PHLYouRxsr3CMSjP4h6QEpl7V/opvpjZZa4XkNFaw7X
D6HmOjma+Rz8WJF9uOsDtwW/i6/WU/xpvjduPG2VkK6+ugjgSzmNwQVaE/ev
aalUstkojxhA0HWRaNAMFTlZjI9Fmt847xGEeYNTOlXhQpRq9cFdckUgUsDB
rHUpvgdQvZ+js079djcPfTGN4T3jARRp+QG2TzPJ05A422VVVhKU++vzJhqm
kgVUBO8Aga7bDYoM7Az9TpTZL5pNR0rfXD8Sq4ZXaRuvfm0ZUXbukJiDhLlu
9wdbtbpYLPQPAv4UzX+8BHyfGMPj1IvfWo8xfBWyj3ikmCoSTk88KAazFFjU
7Wp8VGqylyi6hnCSg8Hv2rVOxjMBGFJAg5mOH491v41SLO6Ylr28b9KkACGz
XFgTQHmJKJq2fgLsmPlrw9AhqUwveVFcUD0TM8bpObJ5qyqxbD9hccnVwrGL
qWOSC19cnTTjQEphIIvS6SRbhUh7wnM1io5GoSPTyFitPAKksUJArjoP+2+2
4VUwYz77ZPaQRrf7pIgNCCZqpmW2bTE9DQChLBKSjRYaC5VezoMtYLug0/vC
Ajs4QkKJEesKKtL0l6LTh50+8pzX543fmjW+KCEuk1tUubekz7lY/1rXg0mT
7DXNL7YmqM5P1G73w/Jf8B30AzvpdifANMFbQEAYSBCk9T3FVZUCUaap3k7d
/md8WJ6QFFtCOOlLbzURCx9CEIjNN/WlHIt5c7huQSy07gUSeW/XTT8UQmOf
oElJHqQGwn4W2MQdHRXZ1q6qg1FVaZFtZUP/pqz662q32FzcxhOfmhrgRFj9
Z7gfXCQK+3GMlJHjBdp5CwLZ4XjARjpVFGMwOIxZgbM0BIVNSD9HDGBQ44FN
GR+wm5kgLADIvu6sVZgMaYWRtj3pLaGL/aBgUln7wTIPa/qALhVqueuLPLSq
Gt4be632qcJMWk4VQi8YxTVppM0lpejrriClutSdz4F9UnHEC0wYgpwQFHOP
KYDJOkWXZK+lBVtc77JO5dw/wRShTb4rba4kj9JR91/waTd8hqq5EztUcgf/
wv0Ca046Va+GyCAn5ELCoV5NWgJ1bghNyjCK9E8rttGM2TCAwWwi3M3VNcAT
Co5GSqOfK+yIXM4aWwQQuY9LqzybzZCHvC/2J7njgaKMwXdklOYtVBmz87c0
+2+ojWKMa5o3G1S6gDh8avz6r03MCVd0Tv4fnNnI5SC/Y5U2NG51jIZc3tZ9
Dcf+HLrNNCzmM0DqqJIpUNlZkP5C4ZqvIyW+9+IN/2gcmss5tw9B/lsVGstc
tKBsJG3E4P4Tc7ZyJ2ayyQvUIO226SDITY+1b6tEULEpppw9VyNIAorz9NUb
YE/DicB5mDGhlKHbB2ouuc7Tom24kvmmggRX4T3LxXtvD1Xq0zWmbnQcoIuo
eLU+5jhWm3zVsOXle4OeVZDp40Ab+LStknybnAPLjNTPj+E0GaP5ircc5kWj
wkXfbVpNRCveK57eIvEXQyclwgwLaJ9S5z+MTDsTcrjlwLP3jlyCNtKBfdsM
o9IOcMGNi4l0a0XlttBziO3wpuL5wNhQrr3yJrJ3J2TJ8bPQ1fgfH5T2yzjP
yfXKa8KtT3NfUkPqmFDxXRVBa1lj6iuTI0HFS8d2cRVPuwr1imAHxSRbl/n/
DVWjzPkGxRckTNDis4GHB0GshYU9NNCxBEyrH/IqalCY1jQmxPG+lGGAiov4
VuIAtlk4mf5qB8k2ia0udDTlhi3VS1tYoaQZFW0GuHG8KucNzr8hWPsg+4p1
uEqU44o/hiEc7OEWopXglsrQC5UEUbNzfDY99YBexf38XKh2OgxjVKiBU7ME
hN/ZBfB7UYHk8ke8nhloMUk26kKNJ45ytyN79dPUazx96n2AJgZdVF7pn9Po
FxVZqeTs8mN+c602NEqIx5aQWanYktViQgL5rRgEm3UB6PSO7NpbyGUmJTm7
UjVx0ITl7GpwzalHXIImGJ5nz8go2kc04NhLX8DTbWKNWdTwaE1Q7dUFNH3x
fz06vLK1djgYMv4++SVKyfNZ6Aij8UR3xmJBO5sNFdZjWSd3L6oeJBh1o1f/
l49qt96ApCtFBZ1JqNfcebghhWyNLbGejd0hqw2PBJETdB9PB7c5L08COZ3w
d0beP7HYUDlggPtFcU0TAdhawp6wY6tseTilwFzKPd5kzYdnzaBL4Kdib7bs
WuIqYJeTg6vBO8k3dksjBd7pxxDVv0Mw4L6DohdhIe/F/tVvKMPxqrfnyMjb
v4TXD3qLcZFilueOmtelKn6vJaERebS40RvqVL4dxGqDh8M+USX963uZRX3L
vKb5vlIXC96E9OMBTVSilQoqaoBQ8/17gG/gCmaFX4vmgCnJ0XFzi3cgL0VK
3dmwIS4kl2JX1Udgfs9hIiroAI+T8pI/VZnP0i70/aAoxzevGIyKUSDnd8Vw
zpxU+eyGN7UH3NTJqC7YBj5E74TY8AbXrP8uLWcwEGVG2mpFMBKEIAeotEGh
IovpBvNy8c95UeMotX6j+hDTANeiewACuCUqgVDxSnn7YcgKwf3o/bASdJ9x
UDJLiFxFCx85iR4IK0HhFt4vVAS2TgSNmNmWh8dA9HOHbMDXi4Sa4w46yzk1
/MVijv4+zg/84J3tlZghvDYy8g7VfUJInNLNv2NJgBRuZQ6YO23xjB/i7Zol
0PkmYjQXodjwlIwUZtKcd5mydKYwKiE1Taij1zi2ANgsi5mGdPrC+eHI5rI/
SGl1K+3vgA3yHZVlYxsi+mjr+2eRnoaB2ymRY7mkxsRa6ht07Gk64LwJoZrA
b1xRrvkZmgJdoRqaQhvM74mCqkUim3BWZrED+mPYA9cdXnF5qy1I3OlpvzOh
4tYkMIalLg6TDVM9H+W54yrfV9JotIeaoTO+HcPm78k2NhsAIBOF3As0Yciz
/amBXyypCtKeaxfofmy72X2i/PdqKESPPi6QoSn/K6guOIbvXY7YY+FnBWPq
LpIoVuCg3aRYkdq7k4AQK5pj19aH8H8A0t9PC+bZuopvLknkpOA2ZXK01iZk
PXlpklUde1GNZVxfHXFiievUb6/047VzyKcIvMtdoXhp2paigYZUs17Clgsp
tgO7lDrEz3lo6J/+fQbqO7zywv7XpQEsqZ5Dg3zsTedonSCAUYbT4uH+BCni
ZGN+36ur0Oge6nRsiVdk82Be0KSBwkIhLHPadmglUSJ10rZA/8iVbuLqZT7u
omtBGcEQUhtDBBYAcjt2KKlrrXWYxSubvWsuUM9ofzH2AfEqQ4IUnZH2Z2TQ
EzJL0ckaZRPxhmfYfvNy/mYxiYqHZOnzzdqqC1DfPzNObfMRj62QPJOaQH32
YT3rU6AW7HVycIzrPvG6IsIEVV8gCDcozPW6AUNAmi2VUsyPCsEz0UthfIZc
YOZUFMQ8e0giUd0AMRDWh5sCDDMHfNUVjglKmq7ahytmr0tw23+KjEN41YB0
jQ6UkQ/Hv28dOmL5qHBaHhMbfnR+BOBCXE/3e7FPd1l8LnysbgeJpUmg450H
JgjM75IkU4vxx8LdJlWvfEw7yroV3TfN86cem8c0eAcopKniQcH32j7ZUyfa
zyKBWHSgyKGUM/CaKiqaRFJS9HweSTY84NUnpP5xWgJeQ5axEVeYz37PgZVD
lBvvoKGlQ08prHEn6c4nhaZSClurRNNC/bmHtI7uEfAZXDdKRn+ZLD0HC+Mc
EXmuVU8e+pbvq5xncU+4e1sURXsafLjwVpQEFb8lFYtKPL1+GpbX5IDD4V+K
IhjYCwZL2JCqxRbzL7SX9bqB+xU/EqZLs6yXZ8XBzJea635lmhnWTNu4OJUU
4l+iZrm6AE+ReVYdsfYlmd0vyb7H9cFfgwtCXWS8junyC5Fuzs0pxjBMGU3A
zUc4o/jxvG3F6t7t0kw7hCYSKlPJCbWnd36qH3dMFnEKDJxjljBEAq/W2O4s
D1AbhLj8Cv87v3uvzUtIa/VaeveMDA8nkmywvkvwzIiXxKhYiyOdtng0y8mB
6wVPyG8J+9Sjbij/bHOpAgpWnGG5e2FIQPODL+PykGWeVJElOQmfZlLGwP42
GFD/qBJTEg45/S5fGr0KL2XoK+QVZHWDLapUjOubL4VLvH4ODmaHft59urDj
gDUAK7O79UeG+OvEjEoNtE8+NWgGM65ftJcW3CuXw+gCpdeIEnR/U73tw4kj
0FQxUVFo0P5MvvWKS6iSI+WA4hKmLg6UmTrJcsIwVo3xV89WcpoYoviJY9nY
j9R8foM/VY3jgwZMnK/DPuMRR8o03w9AQRIjUjlXvQZRIMVXeUpETRUxTlW4
vyFZD0JwdIMrAywC5Lsn5/TsJPjs1QRj4tfB78vyNV8lTKplL3wqLci9XnGB
IvM1Hsg3NZ7Hx7mfMx/N0dB0pJ4HQm7ootAop6ZYSh2+1ZUQzD8ufH25vUHd
ZqEMkzHhekkxoYQXso/QLu1RWWt5GgxAr5ZkewJ+8pOu7UMpfT3q4n+PQ7hC
r67xAJaR+b0Ym7A81+nWJw2WKBpyL2fUoYHRK5sxMYAU3DQz/rxK9pnQ2yM0
2b+FtwzIMAaha1rXjGPXQ+U8hGvT06uzqzz2xcG+O/gb4xMQVsYF14qUOCjP
wLeFh6c4m6uHF6t3Kq9cJLIK7TAv51JxmCKagurwXI1O1vX6lh6TngK/Tq4I
9pN3q8AaHiqxUr6ULrP7pyXo1kJxRsxh3ajNHCAcnmDzmCM7vMz4I5kcCgCa
1dq2AiLUGWw210+ZHNgm3eAILseOoN4/tGq6jVqrsRYoTH4Obe4L71BJW/pZ
rQ+TeL7BGASN9SphTv0VbU5DMQ3NEiTpSjqtCVEC8Z5rBJuR6jWK7+NFoyJC
5vpso1dPaIKI0DTNTcQ77B7YuusOisDF5H17t+GENc7rj5J1+zYZ5xYD0ydO
wC8xxTpDPeJEF8/1pGXcmdvP1BHfOmpJNAJRblZ/+DI5rGBDAa5RygLYV1Jw
DuzepcQ/UVZoFyW62kTY86kC0Q9tfR0iIYSH4xOgv9+mBLBVgfox079Hwq0w
exCzbtUnRMV0UXDK1v+wP6FOxBSXfL9qrKPmbA94+tptIFzhPGDGa9wYKTqg
Af2TiiHEFBNMEmn8gDZ0rc9FQYM7k9cLYpAcwudFofaE6QdFoT7NHWG745Rm
2l/UDX7fB4s/10B2k2b07vSUfRJEHblHtxvi+bGDRkoAtJ/SpzCNIENeLLT6
9uNV47kvQyhGX5XLUyoi59CTFyngJ/I1sfc4FV1Zg01eKLQ51abNW+vRrjzW
18dLpzU+yAU6/gmO9C887d58z0kDAypUDqPvt/c4vGl0aB4UEfgGDjzlNkgN
YE0/iZGp7WMoVySskPJA3bHwZ+kXgOmVjxRo1zn+pJtLlDELISCaI6Vc70Yk
liEF7CUg+ZcN96wrMPZF5TLOIc7biWnOsXVS5EeeK/aMoCEEf6WZOn8Tp+Wd
bK++gjoDOZPswq8APukuCXQP58aDT7sQzbprXnnzU+fI8hl7BFN9tQ3JuXqu
bMkx/0xc/NO11aNaeJyCpEtdn8uZ6Z/jldUkYGyu1JLBYgH7E1PIv1dX0cWI
WZ/yRYhCOwTYAyBZCdycwOwzHhl5ms7t/FGQvha7Wyb0kXtdaUsLFrHDUOAr
aj+XCkChKQ3Izn6IB8HUqkuCZKHqN6wJqjndeA2r/AgYmAyfUIJE78gwOzhA
37ZoNfVkWequvlY+BzjGQ7BXRTwDqJAuK3MJSmIu0yBeEN9+WFXBxhA5e636
2KRllJpKRDTPRSMkMarfwb94EvhW6jWgqpjPdjm/D/MV6LZ7hLnTKGAI6IbW
kB4PYiOXjtC9Pb46UXxib73MejcLtt73D3KT9bZZmUEfNmoN856qLwIzJGgx
65GjfvjEfFw11vWTc2R4nHWVYvNvQFyAU6keYw2spUEzeOx3rQoeTgdQWsSx
4Ec5UpBxteDQ4teDfYKtK+Z0aSquOjfjUfK/t02FqUauqrDD2vNX/h1BIF1X
Piaz1LjhEVbCeRpP76TdA483f/2L3PGQo5W6iVTvBuGnLmvMps9r4lCRM3l6
QkRz5NIOzTkmb/jbp/xDgdf5jcio49pBjTJ1TwRUgA2cgCf9s0gVZAa0AFpm
m1Mjj2Dqhi0M6CtdUNSHRdE0okvF1ljvKiagy+sKuEzUcFZG4zHta2aVPF0X
iw0PKFLjStc8F6cTHiyTZ4kNgTnYO2LVcP+a1PWpTaKhZxpNeuQefB7bnBHX
7h5uvaoHz/3XDk7fty/SjRzYRaKeHA7w67yCH8iPT54rEkTk533rGcZbDsNB
8KtcweQkR9F1rCX6DU+GkJ1eN2nOTV4yOe7Tu3wTc2qcmEduvX42YHiMTFHa
cQpq0wCP6OYrM7081B+rD0lnHvtWcSDw61PkSajuKxlz145MgjJSJyc3BG1c
CzLAUXW6UMUbdZPNk8D7JCqmhS/x26OeijnifNE6yRFoWObvm2reYATNg2pa
JL1GvKJiBA1eo56Sks8pVPNrqArd59nLCiP7uxwNuwaZw9UoC1Tz297Q48Ss
SjpZuMsOco1DenxPHv71B8nrVoR5lfWlyEPzRjPS4cwNrP2oPF0comQjSDP6
+CtuzyFktJ2FEeL3KqbKyM/0QOWtuubtyJOALfIUfnZY7KcmpBTKErLZr9HY
1c9SgXJbQT387XIfR+biSmV+TEc9mGLvEXqEUEhR9dAwGiOStCaTzBSOaRK1
ijZcMXrKu72Mnf6z0p24hhX6jW5rYuKTF/Owwn2sYOME27QPc6ogCLle5pME
b6QwxmrCg1G2eCzCGPDRkeL+jNh7d6DxV4wV/kE+HTwi1CJzfAUfTWmkKiS3
GEN85Zt47KrYWo2WinXd5ZtN7Fev/iCGhkgHKDyOfBsG3l9OyiZTceqcY+AP
3CK6vA9/ce1NDHz26ze9X/7v0Mh5UyLPwRqr0LsjVkzgsAYnlzpBhr+mW7uj
RY2dZT47kQqqUGReDf9RlWN5uYV4mSo1B9WywZoP5WMT8Unl73J9NCiVcvlj
hL8whE3iNOFY3TUMNCZ+UMJRH7iWZu1zPmAfJweKutLPD2KVkPFDdCTyd4QL
Pc8d0l9Nw8vlNLGvURBRKovXXuKT86SkMDhiXrzpSZBvMfF4Mlb+LyTVrXDX
CHdxmDnrtGgaivZSBr+g8/9YjtwYKqTN1GKdDbrMJtSyOVaMxpZLxUpycVUp
0dDU/gHZGRpnD0jIuM3ByZWEVoA/U/D9hkkNcF7YvFN/F+EXUDWNnV/XObKH
hjQF27VN4D2dmSYFzJkqGL9qZV1oQqZhUy6mwdXMUH9Rb1A4SAlOsGxpJpA/
7Ly/MjD4jrCpEECWyaD1XDv4vDsgPgaP44TOvqW1BV1gU1JCNMH+rv5NdWSL
Its5/awlPwjgIgZoHgjci7qb/OCDEk3z/NfygL/THI0pHtEVgfvAQI8DZr68
nHfuf9psMaEpqri7GPlFuSkfmM/TVLClIaRP/zKv3v+XXzvOoEgBYmHw16pI
mLOv0iY2gIWrYSeM5ufBLghcquEUeXjp3gFOIXFUA6nysgG7tO2zKi9MU3/s
QdLiqAjh8aIaGn+NJTwfktOam0EV6Y4/z2Gy86SWJGRmnnTHPpKqJxStGcUo
xVxwIX+eajLFLUagRlsxxD+gyRCfc3Bl9DPGNywq1uZzHEHKuvgymNFjMB6A
yEkiuc8qUFa3lxgLMVJuufugUvh6aCL7xT8elJT5VLeh9C9Cks7I08IPSDlP
LqlS3GEPQz3R2d7U3AZ16DTQUbQMliK6gu+JG7pv/PMqAK3iRO6hA9jk1sdo
kIQ3ddmfC7YlQL0g6saND69Xi+FusSVvuPeW6aj7HS2Hd0gPd+6763qgo1g3
GKn9y+2qmylPSLiZp5t/GSq2GtmKHcIJb1irY/AMFlqEbJS6kanjeNjWD7z6
aXEfTIvnaBmCt8NAfj9za6jdTtS/gF31BY07kj0WRAFCGhJBJzNNWq9I+CfG
q53KXRe9FRpXyVQrZY62x1PMRp/CVeQqu8ZRfGhlgI9H41AD30RGEmPsMhL9
3gOFFH4Ka25KKbrEvqwuVtrwFSBeaIJpnlSb5x5grJNCxT9ZZDIfzkmHyFtH
Eg/lNk3gUAvK59h7kjhtFNZaJLgB60mfrLZEtA+lelbXwdR755w2auogD88Y
UQsMhLV349lmmhSNn+3EcdjeasuS1Mp3Xrx3dH65e68yF9gId7Gym+l+JVfl
70F/eWwTqPC5QSAA4/WxFtwCTKDoVcuQv9P8xP+pFZH2sQiVVUNrsy8qjBbb
PKpYEJUkUprgwoJxkGEKfKazpOxmyLh8+VTfwWlBtlerIHvNiSRpu5wYTGcv
tkwaRSH/ArSl05LvwnICnXYBiB9vRL5rvLh9jnqqNwHoBmRydXJ6DRThDFEc
LITYlnI898pIroPsFmrRvDJDUNqMJiC3vaHNfalgpGhG8aeGfQZZTmYMPXRR
MTdCSPWFTtKW9x59lY4HgZImkJwEzqQVbbDQ/jo7uVPV+ozhidggjKxiZDAb
W7Ho+cPrrzsnFBmWbHYd6smf8y8FM1SFkFJvj5hJS0ifTWI6WQXBHG7gQScW
wZ7+0aCn+Il5oWTKOY8Nt+YJJiqT/sVXLYWNNZIynY31+wb42gxGHHP1dRIh
sRSH9OrQyVQX9B2Hk7IEcblizjYnwZlKGiOmzOFssp2LB7gJrMNF0U9P8+aG
5N+TqopJIv/OrC1LBhHla6ytHvH7S7hI6bU1SKHOUdG7iJZ96CtvrNbSCWfK
089rsTU2kKY4ieGHc8XGM7vrV3fvvGVFh63GWreYmxZP90olzzw44UgcDtP7
KRA4luAExHGrwlzleYUCCGzZLcGpk5Txtt+6vnfmaYkm8zCKfR8rr+cUTM6u
dwivxsAuuamPhk0TEwhl9e8jccjRlehxiqnD41PaKa1sEsOebK2BPLph+O1E
QvoQx/LUPmwau12l23jFCYCPuFnh4k/u0WJI3Yf3x3vC4LhPsihL0tr/ErH+
YSGfuOeU+AJ+KNe4EqtZCr1FjOY4/aJm1+y9PZ8q/2BlRo+xSJ9/3beS2nFP
btd/OTB4Rm7oIFJV/jyGyRPzEwdzN6zTZR1JfOBVZXI1gqgaAqV4l/zLiiB4
YjdG1r2SpPy2aXpQfekopj6gsq9lVdgC0Mj6TS1PXtvbK0515vvUAFhf1RuN
QAT+e5pQXKp0uotWuEnNuj2jYLZQugqg3qMUYtlheSeXod1TA9c+287l/STi
NY5/0VG0h4CfbcDX9JDUo2xb3cM6mSFPQbWAE7FqtysrFjaV6D3xOERVouHX
2152Owm/0GXPM+Le1Ok0iUSJEZ8RZvxhKDpFjjUt8/0znb5l1Zbc3KCF3kXp
maWLpFIk88FrWSDk8lDkm4PMbwxKtVFOCiDJoUuOaveT1ugXVUwLjIWVE2dq
uAlNIEyi55Tq9b8t6KRebx9U4qSmHIAO/+8TDAYP9BN5kEMOWVs6RQ4Ns0Qm
9X3KqBjFOSWFGiTBNqX/eLJOK+H1YyJzPErWA1xYmT3Z1YIPhL/AqzNgcAmB
BAWbmYnrt3U0cu8cBkMMlOObymIhH5E9RsRfx6FJPR1F+U+KHxp6hZxUgOwL
vopjL5OPkasrqTFT88YSsjlwYpHSc/tY1yUniLCGCi3ccP+aXMQ6MviKmlVQ
AUmadLc6MikKkk0jyWsSCJNRML42IeSBBLGT/wkR9KV8T0eHeq7sP3WD3Wmd
sUTWauq/sPJLbfRRgXZ/gEvhr8u+rsyfxFIhscFJ5/es0eV0J2jkuzW6Onug
n+aH7+O3qGiO1CHVat/JRh2jx+OwLKWRmK/P05ohdSmHoNnDIFnLpanB+g2s
WhaZKqzICkCdjwzBowvWf1yenvkXfzYoeOMv2qJTeTgtznuePYxag8q8wX9r
5MPD0ZelMRwCHPpwxIR6uyCQ9iTVtrihAjys68jsYy+OIxXYhuyr0YOKZpyt
OosKda53M6W8TsGV5MKeSq/tOklXCu0y/8XJne5gzMs1R1RgQiBVJYdKSiNz
zTe5eXZ4dVsNAZJnoBGGOg8qNC5zebrCwMnVlSXdmIM7QuHZ2zMOWd66ozfw
wCetpmRhFjzozQMvladV8iZ3FTj7cICB0O9W7pHcQLO8FVWppE6AMU+b+Vbz
vTYYPxCVZNMjXJyIU62G+UtL3hlOfXQQISZbHy5SN5cdez4VcjxhUfA/UvHe
R/SJJPMrhcuOKQuA9COmgvdP+omeOYTAygYnmwQGR56Orrv/HPFvANFwNCh9
gIG9arISaCoi+HpblDwxCeQlZW4axh0zSep2CCHyMuymBwSJm9dllProef5w
nnqzTginUfskbROQiCGGlKbcWprLtxzUdQqQJbzy9+OnzVUWVleAX1K7nPKL
dfib3CfAsHkiHenyNS1oeTB4odCn8NXYq43xXkWRj6qn9e8hZ/ADvrc9LSd7
xNkWcVGFMqplAXABkWw2/+wN2QDqHV8pglSDrnmPg/xO8b1HkrdeSiX7qQbR
siwOQgLtCIz7JtZ152frti9WINr8n54wnch+ZcX3rzDlf3XTEPKGxHPavoAd
cN6qOSkKlAVF7B+aEq4kiU8p0znzT32Ia+V3+YpYpDiRVnPrtt+/UeHFM5UQ
kXurxNcsd2NYKx+85QCMTHQ/nJwy8mScIjzo97V/Wie7ag8ITceTSXynXPk6
cRWOblLfm9l95puToZWaBV++p86NrzfoZ6+PqvzYf5cCPBfUNlOBnJh4yhzM
i4vz3rC5xE7lWhkl18GOGqA9Rj2/dTK7I0za4x9Km5KV/5txV9mK4TDpCx06
B9uG7bUdopQLqFJzs8ld0dY3VaWE81Zz71d7Sx8K0eXdGi3HnCyc1CwHQ2d/
bGLJlE+ktgOqMZ3uQSm3kpgb8ayFy6N/PEZosxeRu6J7QeBlYaTCKXNZV/up
xNu8qUNwW4bRlzfx8NKGh3Q9IY+JJ+R0RQWtKB4UWWfGk0SpQuKk6toWkyXQ
K1os5fLTb5z24HbcNP2m8/LDt2260nh6Oz4NXd7UFaL5DSaN9lBkXpLcUm0A
DdZH5meFRyOjMH2nWjKy+4ejxCk2JiNlqJb4iooL7jue3vVj5UsMOF5SPARn
vqTl3CmTKhKpVjUNOwlL9P2HQogu9ihpkBp7dZQ4KJ4nEWK1RyZJL76zgdVJ
wm15EL1QeMcgyICY2SP1e4Zp6GM9EZnjd+F70e+LJMOw3BUDjXYs7vmea6Pm
T2B8hGj5bO+kjiyUorQHR10MaGORVOBG3x8st9MGZ40N1zJCyqzhcHG2Cc86
nErZlBT1gwGMVHdJTXW8PXV0fkU5qt+P8WnvY1UK67Z4opM5kb7OTshRpxN8
w9zI0+xkPsKc8JWa02Oj45V92UDJC40aNljXDC0i+wvj4WzRzEx60mp0yLL5
V28cx4i75ZA/MaTbdy8mct6aOq/K2K8LKAdK4E0CwOfOr0nQHZ/rHsBUlaJe
0Vm8k/4X9429Eg8d0TTydI6W1YGTnOFrNjnl7i+5e+K/gwt4H+FEV5QkjJTg
U7bBm7+LYhj3lcW6tYjeg0n4MULu10zEzm8kjvtAeeBGXOY2kLVy8O75Yukz
dymqE405Cfoe026LBpJq30JO/EoQe/dKv4k8yE1j3Pn/vz4kTEG19tmafWXJ
ETXbCHjIAiorIk1IvBzAcaLXxides47C+iPJAUNE6kd+zdSnBM0CGaRwRjUL
c03ec6ITsNvh4z1HugXoGCA/xX41BZevBk1mDv4ATPbC9xXJsMDBGG+iZWTV
GHmGKuQqqBY8YSiuHEUTJWwy38wxFIdepSeVk2pCCworDDF4t5ssvihjJaV8
xlqk7sbeChDEzyZHqN3+CUEMdJi6PqQJRJB6vKPQUoTFUmbea95woK1hWvwl
Ds9hdkbB9CXJnvqGU6ChWeSKjgGxpBnbfnue0Y47PbqOAbxV/GKlY8OYvmeh
B8vG2gH/jkYaHlUpmwt8q3Cy9kObW8EdEZFykic3MTQQ9bsS4nSLOsJzHxha
pTEYw4MZzjd1fazFm4qTvXB3OG9DdLmp0oNS622krI4XTG35e9k8GRDJ29i5
YbePKE/MLKbR3t0AZUzVAuMU4sk+Z2FEMlIf5CfqHlRvjarLgG17V1JeH5g/
0fUt7jFtnsYwWyu/j+V9/aiYlWdk96T9RkcwrYNIPS3x766s/s/6078GNjWO
rFX2Q23YkYFdPKOuyTf156cNroZmv4Jkx4idTwqHD45z4h92sj+u50m84xLh
w7sDY4e2Io9jWpTn/Fj7+Iv/tQLQdUYW+pKYRzCtg7++A76VfAa5oMXdwg1l
2amvJiXJIWzKS4ELQJ6d1v6uYOqdu/LBlId55ECn7P0rE6T9IxXc6Ug/UzRk
ILny1kG60pw3aBRQTxFDefMoXB2LQ65gkpqojoVSSIcYDrSLRRaIrHsWdiPs
YGz1lYiR0Z2+fyKrHFhqKThs66ZIzbkPvDFU01Yos/MPYfwTjXVA1E5i+/TJ
6xSPr9/LzbV5Eq32X+Wkcb3Goc09gvtilhpjprWk7gbz2C1br6tuYG+la69K
zbmtvw4Yq0zujDJ951CRV8CfwBN3QqsEC7GC44/yTTXZ4cN5c67eqM33YTo4
A3M5YYvGtF/5n6OaWDbovSO/Z8DASB0a3Noe8eP1eYeWOIViDYhOrN3q9Q1n
ofvQ6+tQeEx22kHtEYM570dxPUMjEt3C5WABa1xqV6QxjCrKaU4G8ZX5+h32
35c1bY+rUSfboIiQbLR+zuoDDzL0hq2Je2Dwh2nET3oCEGdYMSw0OHew5Z6n
cr6wWSWkUpQAXxdM1YUuPRWe8XstZzmZ/pEicgmpfI3XX9ihHgUnkDg1njPk
FPNnUeib60SJVx428+0zI97IacC/upgW5demfgkSE+98XkJ4GKH1Ary1h0kG
Yxd2KYbpcO65zO4la6Rc5OnhBo/D+9cIkG7Hlyt+gc+P4E2wQ+rBrvEY+LN7
jAJRFOqVhD8liQ4vBLVNCDLV/rm4c5XcF5dBn/RCnlC5ysBvxfyZeKBBA1Yp
bCiVeIA/ylRshCUp21hpWkaGuwPHdr8rvfXwR2qM2cir+DHJ4Z0SJh9GYFdc
zmsteRrgqFoQPh3BEEbIDjX/1ze7KrfvdJL5jrJU0aPSGZ3GFqJ/vobhhGdt
CR9NZ93XCTJY0NbeZ7HSOcMl4NtBNLix/FVeSV46tBoEV0Dr3WTna4wULAPL
M4LP2P5B7/F5oMJKzccB43iZF0SQdVI6zNryGoyKz9yA8IL/AvExKJnH6fSf
AtpRiYiVVFVOnolVR96ybK0BctBDfcJ5ugnXMIU/WaDZTAx+FxNX23DbJhmx
d0NO+ALRRxEArJAVI4eRAnsivaqk3SfXiN0bq9gKdEFOZXHhWTnhOmVbgcz+
U1QW07S4SJOKL0dlpT8bU/KWwzYm85iTm+owLR8K8aKjKFRqZe+WBfECbMuu
oqryEs79RIjkPx7E4WJvt1faALnVISqORrGFd8iBXs74cxLIT6+oVNAx7kcb
H1f9111PpWnPt/FniX8xKWjuMMtwJaMA/ybXxmX/WxK/owD1F8qR7aVLN29t
Jlkm/uZfNsUsAjZs7GZqSm7QYKNKnJmgPG/fq3WAoHgU9uqgC+EQcg8M9uDn
/txgx667LLy6uWF8FSVoxFAs3Er8f3A9gFsUl0QZZZxs1P9XKCw1At3gZIyW
0xQcWvE3c5bB0wwopnpGtQz+pT9iC/RlOJACHXt0Yue/2UcVhP/ep4ON8E8G
Phoz/YBp8eEXkgW6dznn6umaS4iCLyYl0kjyCndBRZ5c9nuu+fhIUV6e3MyL
zWmvL3bPhKURqhxTG9k794ra4BmdKoCk/r3+4AI6smMS9uKJOtZJi8FE9JqA
7EN57FcxKvuOGVJvWRXep5ulVPsZHIQFdJfkPFNet2fUgvjgm7vf41lb7Ik5
wYEoka42ZUw3w208jmEctr6vU6JukFQ11OAzR6sVo76nf0+wGCbFrcO56Lgu
Zekqdwj0JOjXhC3upFs2FwYKNYxCxEXqIJBqDzC93HZDZIVYtENaFSVMBmBh
Wx0lLaXD1AkH+0tMKTZ4JRbOQumYkvHjsPVezzTHWFYej/GZE28V2lLoLZP0
qvmerEeSE/pPjGRXFWdlKM61zva9BqaldPmIY7T8fugmwtIrIs6xp1B/BMxr
bBeAYYKXUdF/oCfLONofWTcAfrA7xXEbA36nhWSHoTA8nRuD5craEROqvEw4
OrzNs64MFW4uPDucKhG0ItdvthB+OmdrQn1yhjcF91Ng1LtAmFKg71J/uV8N
Q/4GVEPllawbBLqRjKcnkRFI4AhRZeumHbE9BQL1LIV3kozr2lrlt7uvGfvM
yeTfvIoqszfJab718M2LSXerqy+hyfEgoLGQOWSV+6yY8A3TJvLh3XeNF9vO
xS3rLcqwC2oQQ9ylIUHPmibeKUgZdS6KwTXgau/uBPFPiNPAkTZ4C5T7/wwN
ei3iIfgorfUVCvWTO+WRBQ4WamL8f9mJmCQ6qd0khG+UMcGH2ciO67FcakmZ
2jqpCOdXTwX4lISAMUPIQir6IWP+KBPgvkr4+1D3dqvNpoxh2heUStC0HU2a
JUaaYPiSSDX/b/v1zp2yixgT6w5MR9hN4WR7Qm9Ld0deajvageNYbpglImwo
o8zqZQHInbiI9BAtyqbh3fPxQ5bDWIm0GX1QsfuStYOiRUh/id4Rgwwf/Ea8
4XvglWQigxxZqAdjcMns6yejneKLNCodX3s17wCIirLTfxOtrh+qgQq+k7MP
gCMVEa1Qjj5O9+cKZrT9a0Y+V+QhGRptZ8smmWudc82msPaYOCv6vBuYRoEq
idP+/v/TlZTpFR1MDid5JNwh88tazQ8WLPu3ZGb4Kk+d5q7q4p6umHDjJyzs
m50MK2Ypc0/5et1o6ERInIvHw2Utjd/eWh8vGfVln8OiW+sua/Dp5mxLPkFv
GTkZCpVuyLbR8bmvRVjB3bYDeJJlxBqfnB2AV0YC96opZcLtpbOX9g/umC/p
uDm4vRZWJR0+pTKGsU+I0GpRkHdqKExJh588fP7LwfYxp8MCkqhyCNXHoqO5
x4JNLppk9HnNHiVpGSjwMByJBcrN25eew/+Eb3b1hZbpwCtG+LOwkqVaNnSe
FTn2vwVfQ6glWj3nJPzMu2EZeB8mtxfGudBYvT2qQyp06bZ/bBSVrQ0IZ24H
6tGhNF+SwE62zvplbPvMndYVMY+jE7YH3+y6hJu+sC56vrF+B6qExODDfAQm
LcZXNU+haQ9FDA/CiFz0n8Yu5eo59AVho87Xk/PvgccEeKK7WaPmBWmOAhvT
OkaD6pGu4nPBhboGFyZZvaYlvp/pyHF3xGp/D4MAIQRVW8imWZdHX87glnVv
xHU5n3+Rfm8ngYf6eyOBXqDtLDB3Bu1c7ZYMBgNfsZ6IFBMZLJ5kbzcBilp4
7hxrFfJh54nF2JWPuEdaPaRU/o2UE6o51oq0lzQwEmhkgwKDxxa0jutia1FP
C6rjiEytOVIiEXwQJiqePYy2acWwB/Z/1keW3TZjEwkUMdd5IyyjRc00GPmu
AlorlnqG+k/LKcukfry5RIKemBLUEIK9DJNdb1NNMONZTqC4Sc+dDzFis1zG
misrXzT0JjkoVZtHZ4/dkN/SPNn2myu1+uDqNBNrJkmSaHh64J3wAQFdherV
jg53EOxhlCtTPy4GVznf5SBF3m3aot+HbHo/Ox0GHPnICOGrtQyQ/njrqLaD
wGGZ+BiaQPLXD7Ev43CrRCbfBZ56GF/Yt6dwNkJLG4vux7w16rX+XBUKfVvs
7X9/rT0Q3Lub2NxfpSar30266AAlw5MSlQgHGmMpyxKXQLzr7OlKvVqfKJL0
cRvEcc00AZz+1g+9w3O+Yp+52Q6YFliARfV/0gMHqTffNudbMZ6fm6hJY13p
5i07N0fByZ1RHGg3YUujm4DaC+MwQfEyq1orE4yZeh0yjOdtZQtFvRzYNHQK
msIgcC9BKZNqUARMWIoXIBqRoApWPkzYtSDOR6bm2n5pHiuFufz+Dd/xE6ks
xo7QEUujUv4JP5yjk7+efhz1sVG6M107cXNQ2buRx42JB/QewFW8o8wHNivK
6tytq0GZlje+e3s33d2AzzXxxXWqGmcKjGgV4roLCOaZGy9jv6Zoup5MsLd3
GT3xC+Rvxnm8lJ3XrAqQwSZ+rpC25vnIfoAcQGcQVxy5k7eGU0V9kQsJaUjq
RjBh71V2v8obHKAhxDozpbdX5gienerbPGq8xzVB8PvYFn//0QLYR77wtwix
SpC9UFccymVOby/YWGA6Aa0gSiceaTYRiEbUI79sp95psdPwQSjIFZdelBI0
aRpqU9LlcgFt8kDJtdEr5C0jZF8lW+14FMQF2Y45ek8tExuN/h5gr7FXxtD1
JfB+TGjqiXn+tG6JEMqsFnreVH1/8agYG4U1blwniSCAIh0M6iWHDscB4ZnT
+XvBEOeYZg9Aav6HODTdYZdSGNWCXeUles6cMi5XdpH9j+9CeQ+O6hP3N+21
s3/3VOuac0ZwpYM6ua9wkCoEqb4h4nDsQKy7bPU4jfCf+pV9ZnLYWjkD4t6k
a4k8WoVujIdkClaslA9y1j3ey9X4vrl8sS0xQ82tJyCLisWuJA33vQabz6rg
u8XXB169nsytjudVMvWbHOa4yoAYgkWBb1w0cMqT7iVRXX2YxOmTFL4ICePi
SbbIV5Ej13H5fCiEg1yM98irS3l3vAwFcp4mS5k7zOc1GUGX20bwlIEqRAW3
gw7+BVpm2PYBCUq/mtLR3d9AJpNdMT6CfojZ8AQpdz0lOkucCJPWxmxCQ86x
sq4EWCRcmgD2bkg+gUgA2hUnvvmT9RpY2yjRU0bs/wL6G5pkW1zFaKLutfxz
H1SetyPnEV4UA5/BvUNoRmpIZean/xTDmItvZouJczkLtd+5eyotRoR0sRjw
QQWbPrKezkrdYgIVvlXowS32iFqyIyZyBEWxD8l/XotN7/x9C6vaRLq5wMop
2RCWxR6HwKZvoYOWDPrJeqqwB0ZpX0RJMj+3kqV67iDuQzlo6TK2b73kA11Q
Q2kM85J+0HkueumrvzdnsAcoGIc8gOTcMbTOZYRVL7cMgM5S9eny93R71JtT
ppdmhojWvGajZkh2De73Dy8Xp6BwEU6FmytYDj6YfkOr5H2BsNJ+EVnNymJm
MkwPscWtAKUd7vnONmNvDodIhPjc4/qMljEHppz1kiDYI3qjwMFpR5IPvkyU
hVjlKigOuOkpLKdTAnlZrJTdjo0d4kBVRHhNCiFhGu4uQSvs1BX7KYagqzHN
O9mE8t25JTHu6MLkVzNBe7pp+n0ZsVL9ulfgNeKCiUUcUGwbGdrEPperXmZ8
xig37Nw8K5rcn6TpANbj8DlwjTqQHzQVieAE/EJuMUGWUDL2Va/c2Mc8TtXa
CkjgTORM+LqWFnjM0qZcoqVHaMXcjWMcP81WtCt6B2ZCwEGCo7zN54cy7wNt
LdRX/6VY+aYfDFgg9GpJYRIGQocSmAJMowfdSGYnPx+HIsDL5VLlBeUs+WzW
w2ddBuhb0TDJ/0kLzoNAwKWSX5pH1b9fxE1cU6LcmQ73a2TCXgwP777PUcrL
gtJy2o8t8QCo6FsNwrLVWTGOqi7fVa4Oy+p3sf5/0rx1TLRu2ave4baoZXO5
NFfkSN2Tt3EeuBE8DvQv7BHhR/aF0w07uUDrGLId2Ji3kvBpjP4CTeSyepT/
kw4cC5T/L9nSANHHjBwk2qgewpml2VGeXqeqeumHdpkCNia+5XzjTYe6FolQ
N+Qrv5L32d57SuC52AeWwYhc9oS2U1Npwt1BX9FqdyFWZOh58fLlE0zUUqoN
UPslQNJKeqJwSKTR8xyMuVcu6CuuBTYrQE1+fXZu54Bhr+0D/GMjDi0wb8yR
GlQC+puYxHmKM3qjAuGht3DRW/2DmZCzgMM1+t/VnrEmSutiICjFK9Y5vDCK
qv5MVBdWcA87j22AB7jucBdldwgaOJaFnfVLGPmkelw7N/fUwKJErDz4ewEn
b9sK4ix1O7PhNuU+L7384b5SPEkBeWFTEqjQBlq6JgSeFrdW/IXeQeE30831
5ks5AX3+RIv4OOrwXCoBA+UwPh/texGuEc/d6zhBjvN7qkT5+nTOwKsUnNbx
UQIzUN4G+gVpKf56rkbvrjpR3v/LUkLhkqeTHIUCKlwR8KSOY6cad36oJLv/
bVeqkzIZcfu40cg/38jf4+MVhN+7lZzgSzsg+8WTtwIjFH2uOP06hLEBhYYV
u5V4OxZ+CjSfw6cF7CMXP1/tsoV5W+JzyVWFmksOahALn5neic5MuOdNF/8S
DAo9I03fyevwdsjmxiYiWi57r1WC1rZunL2AcV0bkBC1qjYD46kMMDKuorOj
C6CHQif4R6Cj+etDrl20sYAuP2UU4y9SGrQ1WqiNsU6Yor3dV4d/BjJrrx8p
BeG46FgVOHzfrRb2IAaNZq8o6bKFbL5VNGuv779hDLY8VLlestYlYuude9Cc
4zjmwDc7ISdpmspqzwev39dZQ8GL4cVcSN9F7/aobOlaZWaJraZvQjRUn8Sz
47XOpOvarRAorqhFtx9Lq3mXDDR5Wxo2Pl7GTzzQTRE/8zUomfLDSwPTmFwE
yF2WRtTjJG6+D6W1VojY0arqS4zrMcZwHng4LZZA7V5IQqXDP/jTPhFlS3Cp
3tbB8VC+kRQRcAkCe/zBiTiWM3anqL1nVbkJaFYhzgd7mMWuGAtRc9kc7f3k
K+RW7ncYmJYzQkOTUX+C6QAvOywRB6kN541ss1inxobZzzFjNTWJBZA9UWX8
oETEVjGYqIEnxZfrLYz9/9sr1nIQnzPU1HdF1umPU8Jps0jXKqeMZw9e6iE5
xQRqgGs4GOVvTWDjnKI5Byc7Gq6/dGWdtEiOeZbw1SVC4SRzP5MGvIH61jmE
ib5o1/C6wXHMRGZ/PllBJNdN0tvkuc9qyRy0ZcO8BFV2b5HJMfKw2tajkrpB
XsOFJdZ23GFSEusOOnu307JQAH0f2cwdrR+inzG6xk6Dk1Vn2aCBE5l/Cc3H
KBSCBaSVmbbkO/SfczzTxiDz+3xVjm38QHbKwpiZN4QSyfNnpcQFO8AeXqZ5
m6AYvMo8DFTAjAvffbqrk9Tzm/SVqtdTRxDJrhAsUncfPzK9eQGj+aurxHg9
FK70ROTG1m53TeQlZriIBiJ7Ejgq5haqN2MsTCs36MFvN57PvBQk1NQFPvUp
pQ/CZx68eSDA4IMAgtrWmXHx3UdNHYeXrEMTFKdQvYKBssyGXtJwbOsjhl5o
y3ubXOzaGd1BgTOyk3PdEY7FHyTedptnFv5wWa9BDns8X+jJKgxHqbIawDtw
C5O0Pe0OljQKx5sfL4sObc2yC1uCerEmYk9TZTKIyb1yZ/CjRjtHnPOSBhhW
cGCvYJA3KgXY/NP95exR07k3LRcHAapyU/o8i5hcJw+y+gRmHeTQV/weu9uy
m1swr1si2lNo9cfgy2vX6st7B+aYPXwXaTwQi5rNRnFQdpvvuvPPPiddP9jK
MgvT9DZRsMS4fzkuen1OZeUbMm86uWsUzjoG1DHEcxLti0jhQ+wg1CUGRXrA
HpfWLHTu4BHW0QbgxOXVBYThZkpF6rSsXT/vlpyYkJLzY6gll06qfdbGcFwB
pBWZFRmY5ukb6e9dDc3nDBwTqx8tG8M1jdqvaEfPMV5rwvldh5ITQP135bMr
mRkm8iEgbGRG/jdWu82hsUgxjFgii7eSRrLc1j3JvV+4vsYG+YRLQ55sNVqq
PjuP6RLUPuzTE/NSMnurX/ICLeyHSAor3Z4GO6DCGrMfGsVh3lLe5Y8fcamQ
W5Y7vMCdWssSCuwfEqp1vBma33FDQwDppUy+5IGFTTtx0wot18f5tOSyQo0m
CrdnC+9FgOobchFF4e4q2+GknRKPej2YcMD6B19XE1qW7UYqgpi4HgNay4cy
OdqI8f0quotHvkWBaMdQoWhR9iScxvg1d1UARLinN4AbpYWfY4JoT4SsiN2+
OB/sq6X3Obz8wBW/HoL8xMLzBTQawSsOUGln92cU6bv7c3s1lNfPOwQyaMZO
vpaU8eobT7lWZj4I2uKVVWG90+eq4BIPrAJ2/voF//n011NtsgxTasTU49eU
uR6J5eNIu5t2o7FP6SCrvbebC0BITefwUMGr4Pd7aBLCKxoQeyqvfaXgIJJH
3N+UEK1JaZI4ikbaA/ZN0tktsaoGHJkwuFRRyIx5ZwvSxLnin1vxbj+jCxE/
GL0oY+oChDhsVi0qUTQgI/oWbuo9qy24TG9NhE1foVBpIcGbaWbA/+9BIxFL
G6QTRMOdZ5kUnHQOxCLoaPqBbvO8C0zcWq5URMBInxQNnfGCS6hI02iluHVo
3H6V2Rf9JRQHcjbeDJb4n/NRaKHrZLouBY1gK8/tC0+OCA/gWzn77Sqx02he
RGERA3QseSfWuAno2BB3CAB/ihd5mkc5V1p0PT3P+Tov6eu+pWuRy0kDeBmb
ubTRiilpbhxxI74laK2vy9bum9K5h2I2skUK1tlDwN3hHwiV3eKFz3tMcATf
9oCI4OROjKZq6gLhLnfur9eXuyOT5L77q/1CJvivfFdtVUGz3z2AQwLa8v1K
R+RHKb/XUqhu4S2l1qSrtj7Dj1AHH9287j9/P6sZTJmoGzlp65S1xcrr3eA3
pzKIVwPud31G9n9rCgX/d0/J0DA/mbypDeytT9sYZgCR2ACRF8cihL0M505j
kOUDISYoiV0IOgE3jHxoZGy3XQe0EGLKeOUfu8rPsaoY4mr6IF0mTECHfw9R
wQBi/kDKElSgHi9B5VGzOJGHj7n5IG/PV2WhlN7a+G2mlI9RAMi5te2YXPMD
XIpGItaTo4fbl0KHXrIhlB+pwq5vPRQvsFAKEub7QsSHxRf1KMYNOJH/3eaV
h6GTrKfprmnVzOyQGRsiLXsY5U39rJTSsWSuSZjqWunuqKU9CiWMifOUa7XH
YKp7WGsrPZcquozVsEiMaX7zwTabqqWksKypZhU8HOXwM1un2wbT3q2jkOve
GYUFzCGEtVAspcGYfLPX28oxw0c4Qe53HCWrxhNRVzBNdjQlYpWbRyKEffcw
jEpp9Nos1Yq8v46ryhsPnN5R+SevW5m7/B5PzQT1+VB9AkXHsdcTPMTSinDR
5sifjsZDWTl7sMdox4opk1lBvwjPdL09EkWefEsjcxCId4+zJ2A1R/xuoRod
itDn49PUGSopYvkEI9mmeWDp2q1kYpb2fxF+/IPozqI/iyE9O+OO7GkfqqX9
hYBRaKab7QAi8PCoHlq1Ty6iLt3MuegbiE6f6uDazkqWl9eGqkyLKR50tGJU
EcOlA2gakz9BjdjMx2D/px7044Ct5uSPSHxpT/kOWxieJrSKcaYvfmn9FFmg
U7nKrym2D5KVQHwPq+43aeyyn0h18KI3Wfa+NmfKbxi/E7ugS8XDX3AtbMjf
vMRBTauqwVe66LJ5+7lQ+EMsDH7bV5DiVYd/FVHjj0xVc2iRJPu6aXvVIXIO
4w/tMWxobC4Wg0NcOKR2UvwYzt5GZpZTPUJOZUx/PJkW4zLzQvSk6qbSkoW4
gTyLXQvij7V1EEpuRJYIU7vNIb8WArX1pHu5FrvfnTJI9BvaRLwl/rV4fUhf
irn1TDBKDrIX5WtRhSPZUOIovUyIAwx/yOaxVLgzvMiR/4dEZKeFrt6RUbC3
1A2t0EHinTj/dIi/s6UKAEM8q/AAVszLIN2bteGUvrt5T0NClO++frsg+ubj
yfgVnUDQaVeX0R7prUb8LIjX4tX7p4ytIJ6LvXX3/qQTgIeGdFQJblSkCKLp
/G9Uufv3s33wczgHFnooAw28AWlxKeEhR3Vxoj4zxKOfATmokUE/cAciBEvR
PAIF4N2iKQQBc4GTUlnDcBm+U4SUhphc6Zr7ncul6qtEtCJFbxYW8E3znEm6
e59dIQC/JeMAGD0FdytJNnlUAcR1OnkSi+2lJhr/Ug1SXpNgOxCGWmqVvw0v
zRYpAJOgRZQ1jXGy6pRnekWxTGuqdDrI2zWI8AMsipJNDJCvT6TUPyJoYdbl
y+sk0cegj4egQu0J19rzHdDg6xM2/fvJEofIWVh3L+x2k6/thDFH57/pJiyf
agbJ4bfHR9AdjKfF3oeycmzuDGp3qpeCd2s9l2pmCcMRBJrrrrbeRXSvaW//
3cL1Bjon3XH9nDkIhsoSiknYkVbSISZklii+ilpG7yO28wB1upJaeGkJr50n
xfuGG6CHgbr9Xx17TUtcC51d1UyR8jMQJom2cEcNNgrQAxmYqM/bqBZoGB/S
OTleuvWtHz5ecY5or9o9ntsdjboBx8xwXq/nCwAJpOGIHbjh5/V2R54Je+PP
oeO1CgfJ3VAzZKg5ZxrTywc7pI4wU1KLCdoIM67fkEHEhM9Ne9ns0VMNzA1p
Mq1TuJx5i4oEIW2BA4sgaHyMDUbVVixjFIb56MmQZC5/hl8kHYBI/Vfjjw5F
AszPHRHsKKDnbrPRufmZsxx+216Z450oOIbuHrPCFVFi67bZK3skqHd+h3Dh
c++2lfBnR1tHfnYFa22LXgbIwFAmmerg6ZVjFmLhaEpsVQjQLtloYHxYSVjP
2W7ffXntHmjSbyTxNwkDs4eKhMuSOlO/E6jaFZZV4HieNJ99B0KWF/bmoazM
3sX7awYVC2vCyyJ9YR+rNGo+rS3YUhfvQA4G+QbF1857MSnILMJ6y3LEpQgD
jNBWEuxvda/cSkfr6TDm1+fkLpHd9azzficEcyeakOvhYMccj9MAyDUqrkMA
tLfQbPlod+jYFHcQvyuH2I4U2nGUI9DlR/gcO0k8xPwqZBUTHOhIOlF55/3g
v8LU+RuxJiJlRY2m2zMoOL9GGFUdNBJcUKohlvHZoqSGGIbNwN7eKdPX9dDt
AaMs2aVJdIE3CU9VJ1Ca1Y6c3hFO2Jk659V6KYEVaz0fKYPuglDm8L3S6ex4
j9doDLRU2AauojqpEuCIG9UYRYmFhYiZcNiQ2BSv8fE0u3LlHSHjDpQgxeP4
4LSqBd0neEMFGPTYVacKSkbyvK+QaUxSN2tQORrKOoOJdsj+S3BG6tRmbT+G
j4Q6tlXrC+mkZQMkPWemMVxxkqSMun4Upi3Pe0AEIgOng+crgKup7kXeG0i4
1p9nvYw+eoz/aDlaNsSNEf0ptNLYPcOi+2SKVjfyJHjMl///7OgEgtmvi7ri
UMFJYZDdlPf7j5KnXrXd64DKpNz0RnTDrCdTKM4BLiEai6vJVLizVeVEjzT1
eo46oA3h+TGg6hIhUVmV6Ue3iyBecePD4tg+aF5TTxeqg10UY6B7RdNqeE2+
Islul68I1Rqm5kus+Su6fa1wtHmChH64m7unT0BM2sejLCSK0Wqg8qKCap6g
pRNjWuCjXWLstFWEdzYj2UIhiEJ+wAKiyI85VYB42L9wFZSg7N8EitZ0B4cF
OefZmjIi6nOWd5vbpzyDFl18gXrIaGqJSDnXwzrziDFhv+iaMLT+bqVafnsp
UYCNfypIwP1K+YQ6qwRLB3tkm8ViHzfsVtW1zDKB3rGzbF8zdyx+O7NID9Dp
cJL0nIpmE4l22UaBY3AyR4s8JnQR9RSxP00Zxu2WozBlyRCwwi+XghnAp4oq
KejP+YYGrcpyEpa0YICvJL+HolpUu+7ILaACzUpHX9J5gPE6uMLFP1nl/9EC
3VXu9h6kl/lUgRRbPPPcTSIUOGTWJV7Kvrj9kdWW279e+Z6Bn19w7P8M1xxd
uwRXsvC+68nU2Jnut1P0qkbo5oU7dvxcrTAMEWgCqxGdL7McqgySlQf6dfHB
nRGuCZbUxBpwdu53oRSk+gZ/9+Wa1wg6+E7zXcpKYOTunxpI1g5Wvfhhj9oo
86iWn7Ya0805Vce9KJHfVNaXR210SMLzHp1hcXGyvv5cOs2U7mLd5lCxWClg
UpFgwZSmZQzxCc6RhnE1YfSOg1yRCyX0iAnOb0Da542zhaz+/5itvJV5h7D0
lXnu+HINSi6WD1X03lXOwO7GtuhzopLjgYz8NRljIA/0pcqtn28mE9H8gF4O
rf5pnEwykoZRXP6W01f9jZtqOvBVxA5xYlCQe61lhCdH5tW29PvqBA0OcvPJ
2vInuJOfxIv0y8c150llzykO+7GYKy+rTRtFkHJfePYqD9Chyw3Zw3MDOwEw
m6Pi2JTS1d3jhPpUeXSNilwQlhGalMMXhNvoaxWsbOfGNjsdfZhC05DC5LKn
963WOgvXFiOzecfnW2dt+84X2V1IormH+psllGq4L3laHSkZD1XEIOWj7Pm4
Pui0iliJ27VNYBOdbiCF8qDlVxBalz/JrSFKYtPEa9AUmqJKPpQMCMqRHmj5
uBihNqptHZTR6n86rn+SwkLa8gItb+Z/e1GQMPrio2uaN0kpEpSCglvB26Gg
JBqfnfsa/NbUJR+TyFkRmikytrLLhpVEqtukMy9rFxD3Ms55f+LgSNnKcPuk
RcY4NpOUdMsUdQypsYrLWAENgzkx2ZL4KeJCvDd1rHnxYzBE1XXc8jm6bomf
YySR4jyRcdcke6gWPlx5RobUXZ7rcjGWRvpINX9p5KAbKDW8V++cGySRQiNQ
a1DsKERxtv5NKHyR984tF+SycTY2U2qor9OH25Wj782V6PTuoAWMCglbZMu8
h3/acwBhOLhl40H8Zi0RdQQCS6hfh6y1YXPKwGxBkRD+5MB2BzzX6ByWUaSE
79aIMedXXvWmnYr6VR87RH29WyRrrEqgcqm8Xh4D5TreHOt1NA3WtGsrisNs
tmSUDRTlrJveBvquc0bTCKyCPzNjYiFdvjuxakj4RSVqWKJ8jciVuddfghjx
6cxBCjNBwBvc/sI8hxWTx1MX/DoqWGbCTv+DUkgmAo/lMpLoTJU+SEUcsnkf
QQx87qIHUgHDVU6rzD7QgjYUPlytRSyQp4ib9H31a5E9b6DIocDCwCyU0kpp
XsUVQm61ckh3LSYL2mZZp45S9BxEB4mzY76iiD7t4jTmkhpVtpixk3wl9KmD
4R4L1c1N7g2mH5dAC6EdbilODDbPXi8gyCPaQVW8cWZaSX4PTNWnfyJEzF/U
sMHW40sw2vQ9yRLzZh2V17jyCBLyD8nP52kgIcaqkLOPo5U58Euw4m1mknPD
gOKSJhBDBdCvH3rY83LosrTmn570Lq3IV8kyVABrHUk60druoCpnWANXrQhz
kryb/c+hR+3aRos8WCtZ+u/VMNiI/ZQ3NHMNY5NkVcSRGJ1ZOka5N5QZRWt9
+f5is2z8/NP6nqdAgdBmnJdfurdONsCI+nB09o/ivsfqlG5nP/sVzz+s88mt
n31lNJuZoNLlKJ7EgGv38nXfbftfvTx7ZbhBaacZUGwae/X8iB3vEa5xg1Cs
A9RbLxfYAiwBrP7PLJdE9+6nKPQGLtFqm0VF0ARbCJCkQI3Rxm93MujV2a+w
i029sIHX14qQty/RzoXrV4O/SDzYd43eMqY3ZaSGstMVLEE7J9B55ylOMGsO
U1RT86MYodKcT1TbjEPGyCaqgxrDUuKcEkztHVK2NR25V3ju/PxvvSzUJYcY
ijK+ZZOYIndddXIVpZa2pxnRf1tQ975gJ4DWvG/Ljqo2v7kD3Y0DybUp2svX
nTY4OpjjA/AGj2IWpEX3MRyIW+cpbTmfWu89+HzX+0gekQx3p4HWicl3Sjcw
XcrgfvAuGnwt4SNxAnz6XwX1/yrvwaPX+MbnujVnIrox4RckQT1eY5SOyrrN
luPsOhw38WeQ4sLljpDIbtGDYefE1HQ+RMcIuZHkG4hyCLxyuxG6YqS79Gt1
OyU2i/7Kq1xgIJ02sMahg0+OO53JSLaCWlmroawRYcAVYtMf7u29NFTbfo8/
5cMc+gIVLEByUtf1Lf7Bc2iJzhsi2zg02Q1+ez5CelGwwfV8Z2KxRIEyBzZS
NFQXslSPApt0pD8fsQd9j3QSKobcc6hL28ypcEaJeOcAylig4qe9KSmBRvLU
9uf6DO9RC8Tpp0x3z8hR2c6JZT46PgfDgTSXXg70XhQ7UmhaNfPILVqhRgfO
AODZU+bdY188pBWYf13mLzmpkjr85HyHmEnIfDEsn6kOkRKxSH0Ti7n7VRs4
X/ylwtTsRtz1g1Wvk4h7GtqCY4MGm4fhXK9dwScnC8B57lM/91DQ8K9qftxQ
IDSx2xax8hAqHlVOdKuF9WASkqZN7JuzPzs0bXgF/LVdwTFLJMYKC40elHln
gaPojeDE3XwdGNEnrQGPs7P+1bLvPj+njNFLTCLxin75QE2DtpfvGntnDPF+
pKHYd7C5RdPCy3SWcEuySVdtYtc86Lp0gJCwZ3XibgsCrB5IgrNnmvtpXPLa
9O7woEA4tv2dnH5P/hyU9JqKg8xC1Hs7YxlDMYf2RlCRvAW8asqiu5GdHIOP
vqFgGFq1XMSMJq7mGdnW5YHV1c4ElArG6KxL2IByMVSgb5bDS4IRD3v9U49z
X4wwli6TW01Jh4FmsnBQ449SZziuOYvQM87SBG7kcXGJGSLlg6P78mgEvfYC
lF/O+JQfYYcoUpmVXRd7S/IiOPo7axI/fVOZGRzDB8jpJUXT3QuswtjKRtg3
Hl5R8fDsxX45FxLK05MqAVgz7UymSsDhsK/weCMasEO6OmfrD6GXyvbRB3kt
hKzaeGkaTfVMEArmOWv05p6JNYsHyMIanY6Z6kOeXqxdGGsrtoKGx6iYrMpe
zlhr/ApCXMNmhBZiEZ3bx0SuIIVWwysDzOn6SB222+CER+oh7mzCQKgQ4OIJ
01RZF5G++FjCrhGqCQG7Ffhes0QTMi9SLmrsxGM8GLZwdyB5yKKOcX/1saTc
qqbCopydKaDEViRJiojzNXJVR6Ib1Vu8WogyTf3SGZuQMk/fcrP65NjwIotG
pRNeRDdoZsCxAFnVHa3z8Ej2TJAXEOiU5t8K5BH8CeqDyxKiyW7T2FaMbye7
W20iqglGP3BLkg9mJvBkMdTaHgPfGChEXv87a3W4ZBIL7rbHqO8grq2FY7sR
Mrg1ulZDeLeeII0dMS4tkfcjkK578NfkPqIVuNZyK/XnYIV83c4nOotgAFN/
l0wM1Ac6cimemFfF6K8K27zafiRO4bwUIC8ZcYZJIzDikwFBiolicJYwyRDk
YPW3Cl+uoa6P8UjuJSY+I7ydamDSIQruQTzlZatEgdTb/ywLRIEKSLu/0XQm
tximxEAhNQP13rC9z1O1s0jvWMIgMRLGKxGcArLMYyVcHKSq1QL0EeeNCYE9
MqTI1UZ/QWQPIyvw70hmd77Vr7fX1b7RB7vaMkpzApI4s7JJaRqSd6hdgxJq
GWwTkngsiINLkAgXFiYJubnVZrNVo5Owmo2XQ5veCd41YphidxxVS/H9iCuT
Dg7N3lCCRKqklsNEHXU51WhotqTRaP55TievxSB0enT4i5SHAGUbFEK1cocf
nn0qQpkZJ/gtRU6ANUt1QilnoD+ZpwWOSn/1ygCBD5HWzV/ez2GRThOx5VU9
m8bpUfNTGhN72IwVwhpUbYn6dYg83W9120aoQEYq7CtfULPpYdLcRfSOtLpl
X4Ujw1Kpymjb4Nmj8oaMqkDmiQLX28apcAnHG6absLhvDQpf5bVDRXb9mFkL
h5LUX9AqqyYPyRBB1vrmWRlSGKvo6XpRXPzB8xBJTEjxlNQT01r/c0oF1HpV
Um/GOUvsuRKxjrEWeiLPhaCV5NDMcyLlanYvmp/5mAkL3I3Hph25/Rrg+fYo
+7Zev4AwLv6B+Ta1bFN3H9sPqp+1fmy1cclxwkE35OW/jRV4siTN1lxg1spO
pTPCXDYtjyBuSqXzRjvyedlublofu7HYqueRG52bsurarQ9UYiRMAcpqfY+H
vu9jz/Rv1epI3P4O2zKCJybjHLZFQmSTL3uyBigykd9H7mIO+lB1BsAahjDz
W05/JL9KawVsLCtOLHWCdOoU2mB6ZtHnmu4UreRyvLiNGMiRDRHYK+FfJJws
3FYfhQJRM+nwU/13n4vWZkLTQsP1Npw85N1Gk5LT2Evc89pnS16PtuM7m/y0
WJXeSRusNAISdfuLu1Gk5OhXRP/9OUZnuNLivsKf/o/nXDOF5BpIWo0TO5l1
gape/DF7+kKbYhwG8E18//+NwwSVjBOXX4+DkdsqMrcqJNhcWEt+Yix8e5NM
PlsaUpnLifTbpEqQeue9W9m2i3VUqUDGexZcUDsve109ociUN6BzzgFxoFhV
nu78+zNKc3i59LPMeutSxSRMLaD9DEsWm1vcMC5G4l1SLCI83CmcE6w6VD6i
ausrsV9GO9P/tXg33shUWnnZRtaqisPsGctE8uj4W9UgKJrwrYEDnBanxT/6
uo8KORlMNS7tyl7YdxdNZeUL1lixwpfGRZcQwzxiVNltpxvjF3VEy8Q38Y56
RHLZYEo0n1T8hjKnq7BC/h1d31QoDvWBeDZ6WQnmk2ou3IMiLitRqVVmdkCG
OEf614EpWjusoH/Tk6jnj/Zx5aXuXoToTDVDhJC6aMjNn1IYAlsWfhfxxrOw
bW3T58RFZo7oW4UDE5DlVqVZ63r4HllHGUU7eWMW4hTGuvd1/SVu31hu3yFN
xCbN9+7c5SsVI0mvngJQkzx5S0ZWR1fwyEdP0eXaZ/lpJYM4ZdkB4mMCHdmp
e+N/hE96iCVQ9GjZ1jiOjMi9jfkUmGpixMU5LPOrVTa2JhrIQz5WXE/dh8aO
xI2hML++Sd6eT0Y+ELIT++UadIoOPFwMTyWPQfVlYxO06C7mQeTROgMVCv8h
GYvsaj834ZnvarLpi3VZSdFW1Ud3NGLlhtkH9vo8w6PiZV/7/aGqm/n7CgLI
qNbu+zPTuB500uL8WKSp9wvqj9zyqHAgItaLTqnsDbzxD+flgU20qhp2rkIb
lln5vgKPoZIq2rlGc50YVZq2CL+Oyd3ruC5xF2GHft+HHu+Zt3uehZlT62pX
gFFrrcHmeKkbCIZPg6/GkUHhXRrIYmSztNB1zeYprl3dph5EGD/7VPtHQw/P
YnkpiE02njs4W8oEAZPVS8CQYVqvCe7Z3sLElfi4PzENVbp27EvPwNU0VTIp
VJd2cnu+wDH++X7pZgraBfI3NI1OnDnYDt2xTtd0N2HaLCHq9mPseYTuxzvh
XS84DPT3ChoOHevrKmPk7dXWTsCIi+4tT9gITrxxsINytsUcIWI8CK0QvAN5
29+tEiKYo9uAtKIWWwzLM586KMZNEyKiIPykX90RNAu+XiY4MypwI5YNWtE1
F006X+p0hfJCc1JYUFEyzJLy1kGCdk3FsQFUyL1te5wH+sT+zZEltwodMXzF
NC4+phPuomgIeFWNaCZUmq732V0JhDvzB3P9++tqh98L5b3czH4swnmIio+D
5sZG75AzTBYgNNtmRmvu8lTQbOrPp3CyDyFJTbyVFofs9CM4UzeJfIA/IGbE
1rJsltr0HfbqXwRkgQqpt9VSiF+8ufWoQK6S1ZWlyde7QhTMRYH5PjuOlEkP
aOYPKCid+xzeft6vAd78v8sS5zwyqjsxzhXXD0CmmUYCNd2MN7nuyxjtnt5B
kau4oM4pb2Fjn+lebnHsqYY2m2nXQvVq3K7SW/XQsiuqqLYl6MAoXz7HSvHh
ISIkM0TMRSkboe3Gs7tYq4wLsLKoVUBQm0U7DXLprZEUkgCj9fy/FUwdu77T
FQrkI+Eh/A5DeRPFgt5+QYhSTITYysKcIX+4UQPrEhAKnxY2TcHO4pKRs+aq
D/wodibtbPDNpeSRC2rgYykwzf+VW677hUpC0HSfBGK0oFf7r0MiPLjKJPl4
W6OProKUSZhMVlxmkGr4Z63haDD4vSsjbGLj4tm1P8TQm5WNOVul77pv/h2I
XJ+pB4FzWGGFogB1o+tFAkA3mNghYQSmOYJYVNCQorEeaOLSrRqR8P/z0QZ0
IEF/mCoTwt8reGP4vsNmjiftyq+yoG4vLoJ534gSNDDHBjrk1L/wd1f6IWFl
YIYRSHaT6/tcMdXc1ccwa6499r5Aa+Gy4EpCcm4cbw1eBTyG4JEuXOyUVNuY
q9HLgCRGiqVY+r5jT5c8AG06GR3PK+eHcC7M+Stpcb0NjmOBv6KGMuSInlpa
XJ8SvYrz2C8KpvAoEzxtloaLEEvkXZCPCpU3c0h40lBf4ARz5ITWN/6G3JBW
A0i67Yg7Il7KHHf4jY1mOFFE0yh0S/aRg8cTmjnY66hBpJOm6lnRgmnOc7L3
FPbI3g7JG5OUG2BlnQ/5nAew4JBv4+zHdhHH1vn20hPhDTZS8CeMmmUDojZb
UVxj6rGYeLRZ4jITzrpFhzRZS2FR3t6aHZxafzZJLHhriExbFYXWQ5Z87uhE
5CpdgXenE2C9XLd8uc3Jy70wxUhaI1ioG+E/40LVVXHvxGUcFTqk2U26KAAT
yd2r+sAzO157DsKk9G6DmjpEzrMQXbgrah8gZ2LVA2I1HSn3sxZ5UjjbGVFb
mvZwBWF5bc/FaU61fzreXCWrAF6YM2z3rxKUAtLJ/xjnhm7OwTIx41i3BZHK
x3PtP/92Qa2tTA2IC5fG4rln251EhSJIaolBZOkPYPz0vPaf4C8/Gfu4AAXP
QIHnNm1Kuwg9jgqBw1cvpuiRwU5OwEzq2FB3UPIXJvnzLn7N7NVBjLuPtRE1
pfJQtio/oV0n49DKXek/qHxMbKRp9V7ERt8EfmV68OIrIjQVO2p7O/cHgt5c
UT9m7oRUagUdOadJ4sucJiYomx9GK/l9XMr3t7zVNnCYuy/kDBn31YluJOob
H9YLmkW5LNWQrfpw9KeHw6PJsRzkLP00096kn2Unl/wR4csTQzCqb+cKJfOM
eb3y18cZcgC2Vy7rQvr2/Y5I1yDL4uzxjOa9Zdf/pnBQF2XfgFtDkAH3ojnG
F1M0xByvKXmSvz4psX6ufyDxLSkXy9vbqPGXCN/cqmhxqNMUWR66t7EOwquq
aXxViDaSFUDVmHIj87rgQqOMXdAINFTwIJEQ8JQ/faoj8B4SuAFle5vi+s3m
SK7g0nLVW+MIxikYpRQP6ZdzEWhYVg6m/UI2L6W76GQVganhW1p+bTL8nTzo
ws/4MwqH8u+BhRMB6ebeU1l+GCcSokLxBsZP+ORqCtlBlBnK7B69+7QRlLsh
jaRTghsABep0HGiREB9Yi7IPVXlw1Zc0CaE2ZGUIU3h6e1ZlIFJ1TmUiyrCq
Kh5F4Jgyf8pOuS+kH+wQ5s5WFbwydpQMoJvFiph0JKT9lD+8YGWvbTHyEjd9
de8b0ssVl9gXEwo20l5Maz1asMj5Hg7ob6RRVPIeoi88rG8FNnpuPqz2BCuu
fv8YPloFRYoAdsT5qXODgkk6XCzHuRi9QJPO3dDadB40rvXYJjni1YFoolZz
pudINkWUFIEpnmtNG/5BMSFVdMJ0nJMn8EXG9KcEdutjr8BXZ/zKZBbBbwf2
6oXKbwGDO5CPDwiy9wlPDsLgIzIgTH9z4LupCA74TyU3V25MRyYPzNfR2w7x
nvHSroT842PAkQ8TQ6bMXzLi/P5RIUWFqw89VyHPj5scO3fLLTcg2PUC1ANW
gGktGO9UDNkiVpfLvpfR8Dn+PZY7Jke+XVJ4QJrIQH3nJns3NsvDltrhvRkv
CXIRW70z4ImTJ1X2IQtPLWYVlUcdLwNqdhlI2LGTR2kWMjsMWXpjiv0Qgo1B
JTO/6OpTXvP+94xJzAStjz1+Zvt0+E6K23Wc3HIyP/9GT6iabnQHHX8l0xyI
y3QJpKUNmd2apHm/HUKIY2M+fDohQk0wgUyMeyvJsiOABoEeN8ucO+OxG++k
kzdvl5uOIaUbNvUjh2RmPsmn3sm6ek8/swrLeaEVvhmhf94jt6ewmXjUrHfy
JHSXM5WT/03whRupv19yRDQup1E6rrxr5P6kNXnahJELM5d6P/p5Ln3mk+hv
eV3ZpE+Owh8ZxRk0uOChU5Q4G1r6ZzbqPZJrNFU6axzNY2jIj5wMnZOI9lUr
OmX18akHFyKUda1LpfzM1fxt3Q5CjRXMGXoE6asyrvYajhLcCIFtMN78LmyD
qHdyJtt+5eNvXK3RppkrDsw+DYORP5U5o4vwnVfUby7r5NuXAlWp+olr+lcA
ws2oUSvTfHKr5n+0Mfek55jr/AGabm8ixK67k/gokQGK22hc/lbv8TPYpY3w
h2HbtEIwQoJZyVWtZvArpoGu297XX+D5DoVCiD6HiBOYn4Jd0hFGIWmlgN15
itW9fkwxhdFTp9mrM/PSBD9DR++W7TeseSn2Hxv7OMhzGBaFFKdB53HXqTDF
ZF3b52i4RHNuFlOn7Pm2RE7fjddMgAvImjryoyRxGDQkBla0oIhPcogMvn6H
fHJAjjzYhJ494j7flpS1GuMrvDKI5noUHko1XG4bsDAm3Ry4l6ZsaazYSnaN
PGxeINwHwNELr6GJzYQazJD0ZPASWKQXC2WbFMyFCcCpL0kK7zWH6P07Q9C8
Ew4LE2b3C4CEvUUOKUOQPfRud+vQkrr1wt6jNd+3Saamtcrmt+7GQ9ljAETV
JJyA0ogNJQB8Fg7ieLoetpcYIw4EoONDZsSn20nmVZXyTG/jqqfZQQCyKu8+
rc/ZlcgkXTFWQAjgioK0sZW0RSY3fOkpQQ5kTAyKfJUTxxyb2DD62Gu9FN1F
CxnusSnvtH5IQEMU8mxX8a0akN55GDaXW8ndDKelec3cwWd1kZjJNjByBuLG
S6qoA30gWQVeQ1Jl8NyQNjJAcM+le5lPCnbfB6SpsNZyOEY+uI5aclfS2Wjq
2YYRihEtC4sPGdQNrAhqiaqGpXwMkCZfnR0iA7MZOXulbfQIJ8wEQiMIQ22+
YJkwq2jMRdSLebgOxaP2z+Iqb0qpLDdJ42uRNy31JSFdmRD3zwpQuMY2TWgu
mkuv1r4ZZmmVE+mrZsdnZJxbPSXO7uJoTFKkfIk2nq7cTgCIGZWRYWXPYS01
s9FWto2+i/HjqNTbDyTMiMyyXRt6gutYqUGlvlmBZaGUphRbDUiByCQroQFI
RvEZDgvg4V7nw/k3CZ0TcA90uJm9CtlrEbOpO8EX00Fx60E6GRkqC4kc3Ho4
qH9CT3N1tIF4J3cPtJ2dmAZjX96XvmyrftTVoFr0EV4JxXdr2UDiujq27xAF
iTWdor3GOJ5/wvNfa9x0huKAZV3Wji0k89KqLK0KT0oaS7NcJpQ1o/34ZG52
jLnsBn8HQWfFwcGyPa72vbDHDcdAgxwdqtf3qJyobn/7IZ2vj5DAz4hQFoSq
Dk4U8ivfjUwvIM1V27MbsU1VE/8h9wHaC3mj7+vEqBXOGy/YIj+2h6hPmBEf
0IdW6YXFuevra1R7Xq+YToOmTGk4RGpGxs0o6GZ5JaHQmBwAHIeI+pyVJfbt
BCrEcSR4InzBwZgIfbVF4T/R0zGdBvbrMkGPnYYB/bZFoGBE0USZSqbqVSQy
4c4lZIsi9d/7/FmmhBj29oCPfJUJyHabSXG2ooyD7a0XaESvda7CuoOtc4ri
FVvP1oO2Tzymkyy04erKjYQGVvTJ6MQ+jNBxLzmjmSjjBH46yBz6yy0BdtAV
q0+F5y2CAxBWQzxlxTqds4QtNLpgjzHczg8soLjD4/AHClXOTa3OOGaIvG6/
nUEx/XJ1XVtPZQYNLoFbrbagwYoB56xhUCvwGxo/pJdk8Fbg8bVatMOONMzw
azmwIMDjn5VcWq0Y4UWJIXzm3BtKFEulJIwNnoUvrvJe/1CLdsKMCYX6nFlt
nv1W6MK0CXAyMY9aCP3WKT/wwD3/4B0C+Io+S5xf4nTg4IIv7BdsBoUwyYxO
1IW5D2kHNSBj5cvyjnHmBTbcIsv+EOYz+3piefCbqg1TT5mzJ/6dUC4mJfEk
3TDMC4DRrpwXDhF+eScLM59NGISxxSE4O1eOQgWoJvpcx3c8STk7+wDURTu8
UUMrsm8I8acLDVdYdmGaCRnAbqYz+0aXphULWBO6wYNYe7zPIH+JcIRwy/Qg
uHgx4G7JFMD5tONkVmnF7C/qKjdzyA9OYrqvcClp782hpeQMeGKrg2SpKO3d
GAV876gKnkofjBFCm1HKohwteO5HtYiosPBKfHmFUw8S8O2zMI6wI8b3lAYN
pl0dQ4Y5k6YTX0IYy+Eol8JmIWbPsRT0Febi0q0zDOQoTRht/mzuacOapiFj
krORERWEhYEYS0JzKAVknpm/LgMjaB00vzde30HI9IYHR5YkJrA6u7HuqE7a
xlu5OwD9ypSaQzLwNFpagMwTlVkVh/WZUzC5wuWFuU61vNSwPVYdt2OhikEE
eZ7wOgpYvH+PdtCGL4JS9+iFu5yoGBEMFplj2rIqZECNxzXpmfr+nB/VOZ+e
Zv4CWlFWARWSk1DnCigPGtpRLjEyRrztifH7pw64Pbho9MxXzmshF70M7i6K
9fIGXaI/n9mOqeeN+hLyhuAdpw5pjSXPbU3I2E8sh5Ir7FjsYN/Ja3Dh0rT+
t5iV4VBeHe/qwgw/hh9GHd6USn+WnvEXtOueBB2YKJRwVg8xd3EZXPet4nnp
D45OdbBrSo1gbqrF4rcpnVRL1vRCBLJ65kfkuYaq/y/K0K1mNKzpJYlfS7KF
3J4BvZyzfKWcBNxmu/5hd5sqf67+gIflXgKjYG+8XedZP80HqhIxwOtJrzD8
i04c/4MC/8229yTjibku1EhDmPkBY+op+rDsD9SeJFcroLyG0+w965GmT/YD
lF1mhAq+Xp8vaGNYuFZ4xaF9UJxqXGLpzHxQwh7YQ/o/0yZhXd+RQgT1wg2C
M3Vvr61KNPPZZUPdPmfnkTHEWr6xrL8RgwBaj67mLgry5R+HGP9kLc8vEhcy
GpqfAnPoAl5CM0Wf4y5MoSLY1JH3pprmgUd0k9nKdxlozA5/o8OQGJ9FekMf
NOfNm29F9RQrS7qs6wLmoZClC7til99aDmQ1S9cR2Rck/YNze+SnW+iFSvs/
iNqcs/etFxGM+XySUnGoBIK/IKzpbZwEfJ2yZ8SApk11yq1e4IAgLQTEXkOg
Vp6AGuBWy6uLZ5vHyNvk9EPB1unp6ARDUsFacGMQbQAA3uKKjhdT0OcIeu9W
3rgp9zfXwr3GisB3znGFOPfghFuKj71oxZ9uf8kJkrGPJWegTGD+xvac7Pxc
6HmPeCWoCZp7pMC5A7PbKfR1/xinpXKzwe9WkHPCpJdyjxgp5VwoyCxQPNVP
piEwLh0Avv8iL0GKtIcmQ76LPk7zqSSPkiLzPk2kqU6DnNsHS/AoZVMulysQ
YarEuI+/3Mz5z8ayQqSXYkE+UsExn2foElHosZEBKSEfKUSgrx3F0Ee6kI/H
bfADw8LuPPRi4srSOQSRyofPlM7lv14vWO/d4z3LU2cYrak5xmnT9oTuzGUV
CD7TWmcpsL36VwQ9u4/fI4W+7TkDQ/7q5vfimFi/ASmaV2/SjDYDDOT6ZEVS
IXsiIUMMQgEALsVqkpgwK9IR30uLQFjSMi3Gn1+kGsv8RBXEy5BxZxXPP5S7
kdUwTj2wAgwgP8qePe/+Q0moQB2mLMIGfTR+QeQuaVBCEpSBFRFCnfFZFOPE
6AW0XNge2Y/RpL/TFBIQ3bUH0U2EuKNfPhna/vlRMVhcz97qnj4lCNvgIDaP
4zAmmYETOos/KJobtrk9pYwftOiFp5Ky96s58W3MLWhQR+AmSA3u2JhaIt1S
3l7b6XZgwP7zg3OldoZaQ9aI2ihV6DHxircRZusnPbRtN2v4SZ+gHQtpZKRQ
g/k7SSzVNyLeERr1/hRfHScnJLh2a6r6HrG0w+0sG//aLIWsxErFlOhqrB0Q
JS/yEjuqc9W+CVibrb2A8YTiPq4kwI38hHItYRcXaJNcrWAR70/70olKACys
UESTDxkVbpnhBzsIhy0HsSZU5RKfqiTPb8euejQ9YYv0ZhdKcTsiWMCI2sqT
uIOhNvJtjcebzg0dTgPWCHIOhKMTyPY1bcP5kAFuRjbG9bhwOtB9AaTMbWoH
dBIHltOyxbSJGq58Q3lXPoOYJeA0lx4NwM1lH7Onyl2+/67Q3gXgTM9lSqEU
gcynVwkSwGzeSsVs8zhIHbhnwIm36VncRm0b09lPMvChAoxB16dPJF/km9t/
f64V+Jg+lHhl6kZ3kLiElaU58ygedwdPfvqKYYKlIZuyGRJb+uAfrJBMiAQl
mSPLFkBaDLm1A2L18n6qBL7OmUlLnDfzjdgscdwijTkrpeIZOARXNj7xKj9u
uJUP2Vu51DanDXaKTAO/K8Z4K1ePnt18nsFI4331x1GavkcmFveKiSDd0Fhk
gKINqdFyUx+fqjqJkJM5HXv2cdQz16tJ4QtyVWbfBPppLS2+t3FGP4GXo78K
2sBXpG5pbM/8Dqj6eJnb0vgW/Kqs3gdUU/IIMaD5F0wWhe2t3HOdmVXJdqjt
cyh7QSzvr0CHOcEtfXea5Q9garhsPe6ml0ilxlxs+iKiL8oXMstlruT0xpxm
iahmV9gOWkFbXHNcYPRqXK52MH7xI0j/739jcsxJVR0vBcMgCmWhPJ9AUkpp
Z0Ylxv/X6KN+F1UY23LycBDbl/KoX1D3fJ5I4Rq1i598QvVCcxTCoTu7T/rD
+pGN2MO4tWvXeiJalRkWOiUNpywDbY24pjOt3U55m3iGnKQaErkxIdU/leYV
hYEshq8Yyjf3WU2bQzA/mzdS0SHQ/pcAlZqXcq+F8YE4D4a3CpwS7DcCOynO
Kuj9VhRKLltSKyNYl8o7xJAzbtZBCpcOlF2Dn2MKYx3ia5P+eEDQrXivS572
05hj2ERj1/MKaRb0GH2TZtgPCXhyX+Nyi7xAxLswKg9YxMT119DrCNgDnoOm
O5NoE2t2jMA7c3WgMYF4+VIrVHclpdMK81SNwt6N3845dRkXYblrT+DimCHk
unuRJ0/NEFYfM0v23+Xf2SUXIp47ehxyJOcTJiAcWAW/bGn/xQ5JWQGKifIc
DspXRnQGBV0JO6c9o0ArHxGWfFSqioAtSUtsnPrgNJ4EzE0Zjyi8jYwOo7Lz
ErqYya1qiOpw+7cZiXWJEth3JJjwfLcfxzfkWZgXS37idHMSB+p6FDoDBZQF
EZTErky+sC/vK4U7EpvdVAYUxSQmYwjbBxF70vE3N0SvSnPIiXw/Vvj7udnq
8pl60xIsQcYvKEFwFlRYri9l1nWNgOza/37WTJk32TrPM5r5XkJT0OKK9Ekn
xX+uT6wsg4AnzoAPoebVZuGBpV7bKPcfyN3/xAU2ieZHjBSCj5IRlDMqtCUR
+CBFGkPQfcDWFxGdZHA68POfU8YG2oWWf63aV/HdE3nTaTWcH3xgnPh8JGy5
bM6V7wweV6AEEN3LvUoBgmtycfERy3O+24fkukJd8DR3Ht3JF3gia96AWRWN
bXvBd3r7lFRqNNnFt5woXLm/yZp5jLvsiK/eqRvE6R8JMbHSzou7sF9Rch1e
aeC7fJ6KtfKqeTMb9ZBBHtmNKKjGBT0Z3txTbQYeipLPd+NjYfzqlFhLXG6S
FQpj4+THS2CIBLTfcc5dEZQe6/yS7hIUQrQ76FYAV06NKnQ0wUF7qhp/mll+
ZNN4IlGRlnLqvrAzvk9+XLHAjh0OyLpGS6MB2fKrHq1G/NSVV7FXyNCsyx7I
qzkwpA9v0ZINXABvS9hMbrMbMZV6/Xldr7Qaztn4GMImXZldwqXdlmqZ5QSX
WVNr2XmyMJqS8VuUooKJkzCHuyaqaxkkJdhvQRYsK2N/xKxgCFWDKZxZPNeR
o9QXmp8MZq9v6K+rew24F7TbQn3F0vuHOzwZiL7wtUsenCz2XaQcaApf+MqR
HWSUSTqCIxQcYB8fT9ODPhOpXX/0BZdEvJQtNAaQZjV3QPF1KvIrXjNnoI2N
xS07yK7Go2eIlqIYbwylQgv8qIj5wRuPqe6kjHsYjDYISHiZe4nTEIad02Ij
yzGQbHRqaqonC2w9o25xg+KY4UinIWXoB8czYn4dSTVonUqX9vvaxJUx/Ltm
jv4vRJG0nQxvcYRtZes8PCLSJgcoBZOHGN5TygOg3H8vLu0EpWDaj7OdmCdG
+hSphG6CvQ7KcgcO2T3vhH9nf4SqfIxKN6PfNte8OWw5XZqRHEu/cLgp3wyI
7JQBOj142BT15SXSBE+aUKtFrk0sbBFdn9sSztZINMlVYutjIOiGBJthtw7J
ftg9I+/Pz9PgqIIzi/yrmvGUvdr5VkimZ36+GDDgDxdo+ApSV+531Ue2OGsy
EnPROD9Wjl5TY1BEm1fuyjHRlML/cAcVI22VU9yr2HpF2mMnFFacFqiqBj7Q
eDpAUVVjIrdsU2Bg7HiKSZz2XdE6++VsxlqmoyvbIVlA1csreMkS+2R04AfY
wdWiUwLe4tyI0zA6ItC1wqndQT1wPXB92qbDJarWrHSXX3x/lNHW85nrf3Ba
2vdfftEzGvqYRZzpHbRIqRLbhFDxXlICVX7fVPcBxcj7nHu0bexDhO5+Wj7F
uqxN5l6EIXgZMu3Vskggsm/ijwXy1s7iGppQIlAs0j6TK9c6h309YJcVucdY
/4l6VHu5V7H2mBNDJzuJl6yBvZJow6NGJcCxHRo7DF4FMAZFXDxDHK1kFQrL
WuDsAcwX1hf4nDLpBteCXJpOYwFLSgWZYhcLt1yURqiqN5SmfeYcgaiGV4F5
s/NNyAt98gIQe05pyr6K/Tra7Lxdr5xTw8GMJhcBCB0XfhomC5EzVEzMyeV3
3L118UGcbASeZqaTILQeD5f1jFRz8KSRMJ1vyx4C2/WK4GDZnJ6YcR+FRY+1
9Pa6FafEv6if/VVj03i0u/k/+uVafvU67wXTS9b0Wd05tihupgTUtR5FAbh3
GgHmYvgSF1DTKWe/bkVDjF41/r0gEfmnURis6rZnXQTpTqmuWdNIeTgj7Gq+
EVMaGRymWSDZJTply9EnwXD+HBSq4ILYXPVLi78TH1qD7k/ZZxcrDTXQVDeR
i29IEROElM7Ms8Tk+Ux7kQg4CPsBSRF7nonu7gokVb8T5TUjfsjPku5LhFn0
lasceHI7ccjMVd9ow7UUiSjOfrbtH8B62Ywl8GV9O7PJtKgc2aTFAfhGmdwD
d5qZsQ80rpdlizXdmFhDVFMGCpH9zu7Gcz3/Gl4pBiW3F2060ixoIuCEODXq
Y93o1WJeIuCBIlLcN35Pnk2dgSsXbaQ83gF+cU3WgNgbWRvSwghgpUEHALeQ
kl1QoUhp124PUX/dqBn+maVXJvRF2JGkJEOIauhOR2wip1sSOXdPyhpRGlEa
QxpAwc+xW/M8pgk1qOy+r5WMqIme7I/4COVAGnaYBIzcFsNXDYOTJZ/0kz3x
TcMVENot+oZaU8QQWNAqL0vZxx2/TOo3L4wqJRxx7+xe5O6Fhax9u9Z62HR/
1WBYKOyvVX1f2M4QluiJgsOhoVDc3YU79wlB2taJVYu4yv90B+YqoroMesId
LGhx6iYHnnB1ASF8aVP806mdE/bLiGWuxiIanGHpGoxFJaGGEOWB35DikHlw
fOwApeRdaDamnrPHvbDHLXhE9ITNWND1sezqEQx+e+ZbFYfEOZO1UmGTLRyT
Bi2wUOjZFE1U0YnpUym/HwCE8ebCtdYUK0FZiYDq+Vouzk84DT+YZ+ZNysST
lA4q+fE2bi8FjOyIZ1jhv5kqhGgtNO1kdY20c3tTG8brLIQegfIJ7ruwLsr1
SUQLp4VNzqIItHI2RJPia3PRMmv3A9VAl6NzAJr8Q7Cb2+2+g0g4u/2MVVR7
kZwSdmpsrWKndQPq0lGxT4fNLpLrHU30Y36jMuU5AnJ2HHYOBf+ENVUUGuLr
z1IcrAIyd1eP1aupMychTlYdrMG2RlY1Ml86I9NerZT73qZE9MC/6bD0Ub5K
14e7aX3MhDCsYpUihwSSZBPZ2NUjA5k9/eSOWZWu9aDAYTOd9+9sbW4c4G6w
nb4yI6cBVhGiI0nfhidfIa/m2elWTVL1Mf6ZFA68p5oVmsWhvjjyQVpdC3sx
HkoC52Gma/s/XQVMYwyS5+Sb2idOoLIZ+tG6uX2bcBU9r70ebgLXNR64lhEe
CHID0HUQ6rGXhHs7a74BjBhpAQVqLO5vN2VKmZvZq6JCNzRZkN2iA3pv3vmV
J7R1R4s+EzVQ5wVQkv/FsyJUZg+E7GvtKIrJrmmF8lWvmic3BeKCXr1xN0rC
9E7klYM0BzpWj9V8ALSmzLQ31tbKbhECZP5kmCTa0DwRq+1InS1SN8LN5CSQ
hrDWlHH2dW3FWivXisbTF2L9+l+ymDahtSNGN+DzALdHYmTjlV+kYXejzqnZ
rYSCdxY+gjrfO82GxZIM8roU+YVs/TnneGmfO65Wny7jOdL1so0uD0/pFzMq
YzeU5wig21z6Pkzuly+kXi2qx51bBXoZfjkSfBeQNT9JXOtegIkwBGQlVdQF
OCBd5m+/XGBNSUnVPPLY0LTSMohxZKjN15n7agff1ZJZFf9UV7Dk5Zvf3AdP
xnXGQhonUp1ESyL4WsM1xtRYhmiXQ4ExYnjJMrn1YuBe/G+BZEb0CIhpUh71
sV6BjfamRn0uAc/wKxgEgc8wkvLteojuS3HlDTfA244dhWVnoZHoR8DYy+3W
pHAEIZUusdUBBPQ5vaQjuRYHyj5arECBfYDUGtb4dEFCUEnO3XEhUZiAaf8X
P95NopndI+ncXQuWLI49YXsYwffHCU7YE47jn88b/XkEtmuTaEPjHvq8mIoC
V6OILtV8CVNqo630S47HSzIUi78mSXmWtSMBA6aVZ5NKQlGIZykglCsRybda
qIckxqQu79jnBFAPaI7RZ9mkiGeLsV00VuBlgJcAWJFXBoL48W73l6+bTkEe
9qQ/TPzH9VBI9wzUBq6JLgG3Miwoq8zJ/iV/tTT5sC1rp7nV7ZEg9RxN9zfe
SrHNIGWSzRkTCP9NAUKhcn5GXIyePDnCO7VoT79MJ6SuFNyCsbH1KWJ7fWTX
X8X266BFVn/DYX+qlpiXb/k6G0pnsHqljNYW9B+LQ29waob2hdTgeckhA8oh
s1B2IzY3u0cGzh78SEVi/blaMrqnnvz/siSrQLxZ63U0I5vXLlq/Pw2+RwHs
6LGSO3CXZ6bOqrbBsJigaXBtDdPTx7c+age518d7sJtFw84E7mULfm7QvUMN
pbcK08G7BBCPBh+sgYQLE6M4AoYy08SkKsotuHtK1Gtf/RdMDppFFBcFDwUY
R6qYLKaGs5VVJkGd1LJMUsYygrlK/ud8H8F2fErhJt6nvSZ9RukLmWjEFyY4
oESQQ5bMobYXXWRQKwO5nONUFFWLWrWuxiX5WDtTbhq08E4kLyD3lVko/dWy
3zBDL6NUB4SeQL9Qj8r8z1Ol4GhGwjOteYL8SPzE+0I2MpT17fZBZU9KZhkl
5hOw6HBFv2LJwL5xAUYf1S/YWLNyZ0GSXiYeiJSxA5+LfdvPYDZOwRGHASai
nHakfuTEGqXRgHGzqnOlGXwe4v0OTJUTstEkR9xPWvhAuda0zVGKTWoFVM4b
QC4m09ZoiEbJQEk1UdXZwPVzT5bkMwr4YVIgQECH8YRbeJgkOxAz53Ru0d1j
AZpFKzcu4KRoBQSRsV1rSAd/IsLw2szq6kb5AL4UYCnh6YVXPZkafk10ky5/
KwIf5f5A4Zfhufr+mUL2f5nZ1q+iEpMgI9JDLJWGMsagTmz7hPwuiNuiCAs3
IGEskuvr8BhCqGArK/c8hMfCWG4UL9l4Qdt7LYo2ZvhQP9M/zk3TKG6rtKmo
ClbdBD+Ep2raexqJZHRSPmmNeMvVKbcSNitg0IQvJTv4p5lfVAnGwhn3EfLk
YTFQMDy0Ou4BzGsQYJicWt+mT7BjHIUV4139WOGgYzADmYyjpb+BMJA8JCrf
C8DeEEbvkBw46Vwlliv4g2+OrtpFwWHzDHdijk3zeS/1DuIv1sT/UtBmpbF+
VZrp3TM/dyeVmMw3wRwgw02AN+geK+YflQQZ/0BLwV0tLVHZ6rz4nwbBYpDF
eDd/7HYkRgnbTTd3p7pZ8gI290L7eWUjuMovv9F4L1AkinI0zXk2HtlAxkjO
d0AuqHPdzoFqckgv4al6vJ7P0lYTIXG5T5cz1ULHGn/L4VedE9ZkGyIJmJ+T
XgXUJbZqta3Kq42YoJbkLeZS5h57bavanBNrzjf3/mcG8Kf0qSacDYujKd/x
7/I1RWp5BE0YNdFvEbBt6Vsxn87vebakkn7EXoGAPgnyCYxupAH+HqWjUCmD
gwROU9Cx/fSp5GALbq09YfaUypk996bscVE/yw6J/Os39jVyKGfCSewxyJqq
MrAxoie5/k0X0Ox1HFZKLRUecoFzPSVMVpOgoBdSbjhE7/OJDHbrDkyz0jeD
njIDnQV0qF/aYav9uxALuGXI9n5jpJFggvMKI06hZ8K0KzHNUkHnkg+CDHxU
uZd08nQov1wHheC2EhDaPYRGrOxPVPI/L0Rbnkok58chY0sES0PaOVK3FJsy
zRRuac6fVvDtfjvCy0R+Bix4K46uRQz8nxcv3cM/uJHDz555oHn1D7WTiD8S
L8i7kMRk4WpzQSqhA0xIJLF2Ks9RmKovWutnEudlV7+ZSQezcWASEiaczGpK
pbH/iMuctQl0mMaysMrMOBJlFXbNmgOMK7GQmbK4E7qNjWGa5Yqq67MS7hyC
CrnrSbV99HyFLPGfRqgHetOhq5wWPQ0qf/e7ueeU/D00Qh0luyGWXEYodpC3
fEOjkF++2XfP/MCVbkYqm3lpN96glP2XNESYwdiG0o4GvhqSnjiC0IqTzpFm
8YNL07j7DqiCU6iFCQexXBqMZhU/W7RVipz7knMpPeqmoFDQvZRyAV36Ake7
lZzh7p7aqfVCNoyrJk9EXDI3MRYJdhaW+BvSjxbgMNkdo2wwHOGtgHq9PUPV
KU1wwyxKxkG/mAe+RbVRxzIPtUIH4pD+I51oXpgCtuzLBbIbIujMSfi4H1LK
zLM2pA5C/ZucUHfgVSpB4M7DIc7TU+qXLn9/w5xVM921javd8xPQgSdSEgQo
Pr8aJ8Synu0b1/Z7MwEOwxhYBfD+ikQXZENDiE7+a0m+lbFGX1Kqv32jRNb/
vQfGp9WSB3Luogr6BYr4NdY1IQoPuulS6KQFOW8ZmeY3/VLNkRmfJABT02n5
/V5dqgYU4sL4hw2oGgUie4NkagebMvqbGqWEhCoD8+1Knza2m5KjUbQxd/Se
QJkLLzcCLFIgTit6W+gFTr54sHNw+xlA+rPztkbSvIH6BjGaWjdrhsU2xsuZ
35Do5YEi0qYmxm1ak9OigN2lefILiKKO1VSCWbfKJNlF0Z73FhEDZjsBQNOU
DzlyCl1/pdvpFG6SbuMChrhs8wQkgTFffYsXafy6AdffbySCz891AM0VKqGI
KsmxWqOC+mgPmM+Jw9zwPntvU+fH+p3XwQoYXH7WYsyqdKhg6jR/3sUVsaOb
MyQYbrrD8lnwLWRRpf1HNYPKLpYu/jbWNAda/23sCJM6NlGH6uHGx/oZsogK
yk64XnIm43fUxRQww/AoOdzMUY2T6HEzKDcFQ5DHvtBKt3lBuiPGYP9lLPTI
lUDicUGePOWiQ4EpGAJjPAqiidqcXFsYgD5fx1u3hK4qBVGSIYITUwBIk2dj
7LoH9BUzFofRyHXZ0Vany/SjuyXmWvDTPS3WdW3arm5EA7ttsH2ulDhXruHt
q7ftSJKtpJdJy4CuTtnCrR3NPK2sW+YGC/2sqWUm4tBqD2ipLg98KN2M4p/p
lMn6OnBKsq7fibJUOJ2UfxLOedXZv37dpMD03Rb2Rp8IOi6WUJagzQPVN7ON
F+dbdCcuWrFGAdmkqC0ZRivwmSUXunbUkgWK0/2PuS1Vkk6WJKk2hnHKapWj
me+b6HSRFt5UOeurrRmr+o4R8msDZGnyqHoX/tJ+J/Ryd73Xc0eXDsjJXF02
qfw7BepStTpyPbWoiqT7VvAaq3VyWHbOB3OhCU6yxye2sJqdfbIXm7+CzoPp
NAaHdc+6wWNJ96MN77POXNtegcmZQkSDhypUoYFwbFsyOa/h1+xRPPUtNVvf
S8Bjrhrarq4HIpXR72NKrOgupZhwG9Yt/feJf33MdkxOfIh9WHkoE9BV7IRY
QZ2nL060ygwPrp6d+vbUcslXWrBPGOxf29Tg39deKa8sQxL9UvX0fFS3Hzom
kBo2HONfNhhoG5tMe8SKjsRI2R3Agt/wtaecqgMrZwJiv4A25xqTpEZ+RrJy
wDu6l1cTCayjQ4PQbgqZ924IWrGTOfxRrIHE1inNdLVJeYXZdFnIEllhNxkC
1elZZP1L8u3xLber/A6QVufA7UySQlsr2pFjHMo1SISpUKZ1pIpiTAddfVv9
dg94GdUryRVU/6ZB6JUiewGoqhN8AeaKf2dfeHkF10lbFdeLNy9O+LuM/S76
HEqgyo9Eunc+ETxGLM5CXKBtJuiJ3UOEUJVWAmQbqlosVghdwJK2dP7O7wmK
bPX77vPROM/U/7OeOTh05Enh8/Xa10atAmZdr4zIPPE30B1CWTALzzR4+Tyc
hcJUN9QvLKjCrV0YrUGN3m3SpgigGmts35a6twNUCJOgKDquKnV9c+9XxT+j
EC7whreLCThkFAkR/Ewwv2B0Z7HQ/imYs2zmrq2mIKhXp8fHPA/IupTrd+4F
8cRd5rfV3ABOjIE6smgwFm46Kx5x9ibUtpMRNtR7dsTaeic73yg69CVccq7Q
NW0ucyBwRxZlt+NHxYb9n+QE3/Q4/1OYVu4ltLUIAGad18IF08/+enMXysAS
Cu8WvUk46PD7pRuEpEpxGJc5sDJTonlHHcLJ4Jjjt8pJlxAddfJt7zTSvory
g5v0tcjSgNJD62tJquUBUETfTITWVmu0y+GS9U42CFiHGGGKmAvfA3utCQj2
2f6P4szhcBaS470ioR4hQh473S3qkd2d011nhZdlMIo2mwjRxmtMTN+dFeBx
Gwc9qfcNKsOApQWBoECoPJYWBRmYlb+ZEIcubgRLvBRbjMwI5V8oPh7x+Nl0
dTaI4G7xe9uXb6OTacclhLkXJZAK1URZ9vI0osK+GXSKrE+Ul60A4vW1+9b/
pxQb+ZNwKqNrBqwQYNlpbnaEpkS3GnV9NXKMMuQExFgoCC+4klQjlKpNLYqT
x8ItG+K5Ay9liQPExsb6uC1iQMveAmErYCC9pVFT81Y6Xf90AfHqnMYv6rPU
T92oRlrrHj/1Z5363wUc6WiaWSFI2vmA9DiocWTlwqQqGEfegb1W+0Q3JfqX
LtllM9ihP5a7lygMIW3UuKzn8mTqRWlxIiuH2qK7DclXC5SslqC9IB1G9nf4
GULmyMDDRNr1xMGdqlX83PzUDj7iTzJotxeRmgWZRviORY6m/HTgiwklXEAi
4u2x/PldrUjTwzZyx/akU31qSOM4B7IWP5WyOn7LUkPTj/m64v88ustEB5p/
HDiF2qmkuZqO5+sJ5BZCXsZcTKGWBfMzAkBUk4f0obuQ0PCEU1h2vFcx5ViO
3CH5pPnAzykAfV+q4yODdVPNCBaHLM6gSIkiTQe1S05i/zanvTpOtMKKYbcR
lGYTcMOmBOOGXCiEyTBD4GGOV4nkEsWl8Ei6sYaNGa+gmO0fVtTqHKpAsoml
SAzSRAw1eqUWXMYqGlD610JXZgd5A/pDN0nAcOlnrwixczp/+Y27m50Vto0K
evOs5+PzUSe/pnXhYCJ0rnhA1pGphfDXPfzyBku8zjIQtrqui8o5Aqwj13Zg
MC9uFF4NJMpdlb/XYyQr1og/li+gzfwhR78djA3qDsELyPPaYo3Ls2kNptOL
s8Sb92yd0B1uavEDKDaJcjCM6guivY19pBWgllIqqNpzD0kLoTwntYzAouvi
fll8WBHBscofmwHN+c5XChYlJLv7uKWDvao3N1myzmAMkhT6p8WUhH9EIvg+
5hDrkhMeTGK+Xa+MrkOooqYSpPfOz3uGp20P6btsCdu9xXz/NNxEDwPVSACA
gBiT7bF34/sAYmvg5jXVnnr0BZzLZBeN7TxlL2WCXK1S9a9sBUhS5Xa8/GAJ
uCy7yscSrxJBx5zT5ZeJK+5uP+zvMyc7kqgBp3uS5Kjs7GnI9tlmqL136Yrp
xky23A0LaDGfwHDSjenusL/M9p1SPqZqvLUpJOtAFJTsUT0X5jvtAL3yEZGR
LevI6d4QzsxnfyF6G0nEkSF9vK+S8sKuGZ2UaaMgTllCmmgk2oDtP1d/XhtH
uID0rUlH3K7dBjGGrUwxFiMIj6MGJGDldd8NBG7qR5MLWI5dwpz6gjz3b7fG
RCFi6JWnLSg7cdspK6CGlq+dNKXbdQtqur827Y3k2QUHBN3wOYoPSU3SgVgu
B1/ro3l+rvRJaA3bGHLwC8ZlZLKHO2ON78U2PXO+YJdwme8JTJRw/Qw+rDO3
zNSL0TGTTuVhNLMU70E8M2Bbq1XQFpDwm0zOpCp5i/1IRgAbelWir4uppulx
B1FbY5Xx4imUsgI5iY+pLghfB2qWkCwd+4+C9dco4smDQTYm83oO/mnCLEde
hkA0JLEtSAyszPeJ0yMOzJoiEKCHoK+k/yuhNtGaNrRHjsJFdj27tCMD1qbC
MY0UEojLJBngoakH1bFfbiLetuJLLRsB2oNZ3QEZiLfgLgzTBNwwaj74stJa
C1r7EKNXNqIRMzn5j/qEOYCD7YHy9mjnM072rYGfKaUXR6qcBMSqdA8LRbTZ
MzC16yX7ASGOZda042x0LPAxWIUXGQumIYSIJsXwktSQqun41UfFf5YvRqbn
izoFcLQTCo0dLaRj2Vxs0XGBuf8V/Kt87t87f9n5ghpan7hIyxmUBSoPdx4x
O4SKlevXXYKHDsxsyrlqb+0IY6t0ithO6GuMDMKkDalu/2rRZTf2FEU41XZK
VzZIKysocfTNaKNzw/I3uHuYu43jycD1ll7u8E2Y6AQNgmmxLHmUaaSYIezu
85b8DIlhcvUU6XzXIpYLqhIfmaG9by0eLvBMyTaKW6pmBzI4xU73tfocd8FG
eI1gvok8udv/tNi+XOJmkD+J8ySDG6PBVWYD5QbTKvAx3q/DLoz+rDT4aZ6d
fTvGJc1WflwS+PKOjTwrbUud4jkMrMAtESeqpaEStoX/M0fPJf03h7V4c4JC
ciiUEaXaMEX97PvCEvEMWkl2nHrqfj6iz18zlbQ1V43BJYyU7oREtTq5tCa8
9zoYWg7Srvfg7JqSWxZI6LbGeDzp3UanQj192+kXnqCdX/Y0kgYxhvBMprir
xIuW1tbt9Umo3UZtDYsRp8ZaM0NZS4Eaa0KO3muQYgP7iLlU8v5Zm84D+bUy
i41Jx5NqoHZggUQYSsZpqYaaLotCsLFZos/vxteYo/IKptFxasVIUx6abr2k
rClT6vHRjv+qLvoU0K2WypRI4At3xyGAsPSxAYcZyd4uAu0Ty1ympSM7V9zt
0TSkHWn3OuqyGMThjIVMDsBA7hxh4hnXxnO/QG7YDXwmzh4DvwxgHwyRfteo
L9IloZjvGWzU1G8J4m79JxOaiDNHsuHadlbr1vJxZsiyolHPYRMkANyEsN9r
bKau6p6rK6Ei8Vuh8qdgTc/mTOdYRGMRw0gIPydRkUC++pA2koWpmGCimQUz
cTJLhAIv5WB9OywaYYjbzPHfwDyX4o2nKnOwXZ38EJFRoY9rJ8IJL3qNruoh
ClxW7EF7pxrv/rNNZEMjMPcJUNZSHkO++HZGeRIhM+ZQ0OHdVeEwlPKDpjDc
z4r2Uv+zQOM5PPsHJeFGhi2F8akEemF/KL9KPCT2AhKuZOJ2KzPAnKIucTuv
+fePbMtXz4Km4yykM2AzzgLWvwS1mqoWIxFh5lMEUZx6zrtvhtren5sXrAmY
BlrKry2qWZFlohaN5RIn7lqo9a8b1TgF6vUerpeKuXIAaStlUJUk1iwFshqq
/0rYlsuxsQPx/6tkLnlaW/eL96Ow8ub5UzFCtN8S3OZLSrnFQw6XFehrSFPN
H4G9SpTePOpMpaOFWfO0dVgzwP/5ucFfQtHktw0B9eqqQKydyT8I3blawpcG
PPYyYwbQO/1V1D+m8tIpTjX1cqvF8sQfcjEyRjoPx/V4McueiH1GZfga7h6M
FyaAyUcA+mVzM/FE5emngsJrcpbTqwJ0Qbz0g6eA8J350afYxRuCTWsmZx7z
C1D1NbY+xkX5MTvBHelVhKYddhr0sLpjyRGtiKDSfk3/JCi9CbJw2slqgmaO
Td9XyNQIfeTh4PS4CSdunvvlXc0oAsLgaxdoaFuFfo0K8Ix9YrQ13CgIriez
PMl7zfwtW+6c2lhhNC7us3tdfGejVbZu/FxyB3MZunandckpNRkgUz1rTx+S
VsLnJyDs0uwpvHw9StX356WxdVi1GTtJUlHSakD7FLAAr0S7CeMBj5BO3fCX
f/DxKoNdXiVmXxcS77y/cM1RUraDQuS1ZPWvtDyhogGAD5Sjx33pWggnZeid
c0eNGxs5bR1ZAEjthJzPyYY5GWLV+ERfIKc/yT2zVjvrAQoH0tcfWNQ0+LZ3
laf25yHBsN+aKBa+KIm12LHoq7ExNhK5jlHkxqlV0GVeEks0XrwAfIjzZdTN
Xn0hE9KJjZKUJhrSIuhL6K6V5rU/Lifodeuncm2JcQ0WDD7rF+p4mG5Ru6cG
T2HC+WoeifPE8WX91Nat08z2s22vH6ptwMC157doCkjgMaxfEMWw8nmnIFQb
hUoJ+bpNxwacT3liWckNDa3lT6u6aupNmE7nySf2ulxDBner3JGpTYRp3e+n
Pl6f0H+ZQ5Vh2VhbvJHKmgvkNJ4NDpRx7B1dcTvXBVV8Ezn44hmf6SWVpVAT
kKhN7QJZbuX7BGqqN9y+ehnrKg4q4e+29DrYMdgcJcCGkK1N2yoB0WNiAm6a
I2TnzWksVin61vJBwvCBSeLvE0tSiPUTwBBgl0jfBNk+kOy/TTSj5sdchWZ9
8EAtm9WZSte72TjVZZzrfWOsbc03HxciNq9GbroAWwUgFR4Fj2pC0oIiAGXU
jYLGYpcyMEHXAWxWAHYSZFPn3ppgRqImmj/dAabO9nL61r/gYpJpiuLJdhkr
Ehsvesr1GuY56YEYpibZwBiHjIxMEcB1hTnViJ6m/dULSZtR77O2EHkLB+Mi
z+4+ui/MkC8NtoPsMqqE+Qxjz9sY40OzWqBzyewcHjbm35D1gjaf1WgX22C1
7SZKHa1A5h94gdmOwvBkCoJ9mlD3kQv3du+/tfy6VlN1Y5YEokTMyyEC5GBM
r3UfcFsxvppgYgChFMCJQsaoUkBznc5fvSM2cTvgOjAU6wbVoxdNMKVAfddq
/0OxTGJks6o4eEoeCFEKZ94YkhEkcja04IjtQ//hG4LwpYpPA4ZAxXfmXGI7
SxdFUR8/edxLxjmRoIbY8WB4QM4D7Bu/stN28OVp6cL6E/0EghkrL+f0TGPB
H4v8jG6RYXyCay/IabX5AYX16BOEDLbSXr9a4EkTrUG+WPfDlpBpwynmOWkO
wmHnlWhkCC7k4pM5MCynIVHHs61YB2xZQkkMIqA0bsk7ANPH2U1q+xcxhA2R
f/BK4kTIAOs7WI2Y0hM6Q9aeFnOp7isjADDKyBXYXBKjDFsBu2+t+orNulRD
2XOTp6TO4K2h/oj+rB7gTiHXlLqF2vH2ggh3gTwqIVnhhbePor9HadnBEzO5
G/OoVI7Zd+rWxJK8jQ2h7VrSZ0I6VH2E/QWGWi9OhlUWlOX1mSlY3fN2Rpa2
O27DnYOnosiGjMRMnmYZnRado3p2PB0g0G4+ZrYLfbG+SLvjn86NxX+GBp1S
wDRft5oBzCjfOU9kgfAkFn363W+RIo5f5D5u7VYIqRkD7VhOYdig72TFWw8l
eJHgykeQ8QYlOnmMZdvty9wCA3OXN+xEG+prH4d6Va/k+YxGdXXfHQ88ekNC
x1nUiriXBS3zf1Lm+83Gpq/ZEzXcv5Lfnzts4T83p3qDmdkDqRnzpBRLjJRQ
oxdSaFdyKEGf7Ly70MoFm9Vkfp2Xb8116PRXoHhwjQ+GPEzXNsdSB7SDGI8U
DtdSaK9vyNlylBkY5nXaSqKzp0WMOXaVemD3Uj6odhKfJJyDotjGdkvABgEk
HUl5n9hVnj104o5z6dwcyHomIheu5JQTWylhmh4nLg4aQJ0U9CvVxgS/dqC6
f6xuIAwd7R/H4+yeI/l79LA66rr/3dULycZZCjM7cLxoSkuPtQ/uap7EuvOr
7akznYDcmYHtRNud8XujDnRvaDiFBtUe6oTCKAoJqCyy0UJng8ImNGPTVkHV
LgdQRmBvaECJt8DC/Q6oxEtN48JGEd/Aj9bgbVytrCm/xy+lbvjnbvuWwptq
9d5x68M9UCfywDVTfFx/Jrc0y4cTRe8+wPrdNIWL9aJiCjEa3CKLEMuNb4eh
sBlocy5rFgcuIUdkxGj8kSctSRdSZeE4Y4GbwJNtZmk2jJylslo0UlRhICEG
b2ASBr+J2ea12Dt2EiwsMpi5YijQLst94ACF2uOVWpGdz5rkwGWQqiYF0UiQ
Zwc1fWmKPoaB2InTtXTaDm/wuUe5nvMNqXmYQ/aC5/v1fy4CxV6Cy/2azSxf
IdiKVRtHOxM+F9ib42xhNNQPttu8xlZKK3+X1J+MkGdKZcOk0IqtY9BFTfYk
6Yj9JGzssZ8iW/VZ81ZVIOgLqg9gQ791v5x/Xs+o/9QH94HxpPYZhVPxPrOW
/x4SjZ7MhrdjszFOoOjhJ6ci3kghgRMNde9cqF588Am6IvbTgrel8GnrNXot
yZLLdjuPSKejGSRktlHPFEhEzHmrQIO/s9YDKJx9Cu2tdukvfzOskEnUx3Qk
zK4GirXMlSrugQ0nV2bdEka3JUiAcMY/65E+8djNWxAMnCZ1jMvVBD57ICkV
EBHp9d56FtZKnZLW3+vmm0z7a2ltt4C70C2S0rmX0XZZ/QPOhWZGK4SJ9210
Fk+YGPCx2fZldQIQA41jR3MKMpRhXNoQzwpdPE5TD1Dp1euBN5JfRWzlNU4B
Bm3uehnAoIW2Liemt2oRdGiDxviy0ecUerycFpBzY60Whb4WSpo/OxaV+rSe
VqDDDCXRTuCwIDvrbGvZcGpDipFnzzxLQHcHp73ax9W3jyjv0bH/S3HnTo73
EceOY6ZMveWcAEEYAMhjWZn++/wsrl+oeyaXOwaFUV9uLmqhmeMWIu8w6W9I
OeOaC/HqaMBzlkbrGFEmoULCOpBF/f/iyar1BsyG5SZNpulrrjEmp1vMU2fX
5Jcg7YUJbyc1HoiPZHS4K+q0+KJBCEydRVa+u0AR2jUPniNgDNw5CwFpZzrq
4grd/cUbdAwUiJZakQ4B6Ao028n5UByW1KrroSgLHeuJ4v3C3ClZHVZ7HwJr
ifT8PNH8ldlixsjPswQVac3TnL6PMYMnpWhhuvUI7xeXElOZzW61aiGjX9P0
lWGhzs1rK7asEK74E8Ixi0OzuCQlV8q8SeYh/CpXz8bhovlDVe133nsQ4aRR
orS0q9wubiFuoQyzSEUUM9nAncYXZM/5DulBFEo3SyU6N6M7CSSflFoFcYtZ
kJZS967Z8opyLX6TpR26n68EhJ1wbX3VH+iW4yP4KannbZkNIbZQtW5fPUrP
fr26kQQKGyRLpDx697vLR6BFUR0Jr/yMallTUYQsezth7m0eW9sy2/4lLFmp
yaSMyeXJFXOV0JJ4xoUcGB0lbZhErDoJ1t75nnqtjEvEjHsD7BsAhD/PFVn4
gBcrcjnarvTfHmdEVBEPurqrJSlenQFOHTRnJZKc2n79tJ3vMgaexLWpkI0A
NWGzz9OXJZNvLiOUcelTvjEWa+NNjTcqiD4iM8vLqFxoyDc8qGJLPdHsA4v3
4Z5CujBkKlcSmPR+tCG1DHUDAZVUfqglR7yLQZ7+Oh+kZvGSF/R8rboe+KGF
RzfERGSixK2EgAsJ+3254GMjC4dgXS4FnLBp6g4/ecq2Fa0AgLsdqjfjJEYk
wQFdAbcCHs1tQhLpqoNLFkf2uunq/v4mQ90OCmkHI3uUUeBvmuvNimnjnrFu
clFjO6ldOPkXrYXqQ2F2q4aB8milV5PbMKgO2XjkHIlPXV/72tF+8J2BKzUK
LTGZnZL+oFKDYcQFH3X2lyca8CvkTvQ5ukG8uwTPCC2/k0LD3EdAv8REqF/p
LbYoCHJtOWUFLPifNTk3GvvJyr1qvk/l1qRQd34uuurJERlgpzxHPILZjeNm
Mgm9ABBR2i8mYskUVEmNvalL/DmHx6EcglXqZ5fgzjITkW5+fq3XFcbJUyTD
pVxjsn9EtKK8ZXzZWI4ICU+iUB5tX2IBC/DQH1bfahoeithseawyVjJ/gv/D
yd331HqBhIipnjyuILgTVfmiFJn6jGGtkpNdf+qCNCOz6nGdyngzQKI6853F
fFgj1WjcOXFLGx3oyZIUA7VGxQ2EcKzaCr97IC7hvU96cCCulR7c/V4xk56N
17LP/gwFatR4yRAge8qg3gUAb6V1TmPwTCkWndz9HGkxOK1okQlvCaHUGcHe
pulpsc84qa9M/Az/IUUmiAniftPoZ1jjWFzdChMWGNMKCY2wB6B5jzwMfIaX
oUYl8QXGlyG+hB2Jdr9KC5oFtksVHJapdoVg1vJm5LYfBVPoJZY2BiAHw4cA
LO6a9WPBmuN5ooayIJuTxGfBnzGD5e+THGp2GPlV5dmNx29Y+FxERlG0yb5n
LY+D9GarvCOSnwcnnGW8FriHn/ffOI9Efk4bpMxwo8v1TldDMaI6cuwQTRuz
Q5QaHu1gN0nyRiYxHSfMzWF30DMEvDQMe3AkR5pD38Fsri+qxilDcS/+1c24
fqgvF6Q8XwY8U96I0BSD/8lf2DP5mRxDYUKwCmZS/jbSk5Ggim1PC9B4RbRF
hBVpKucEdC3JToejuVoQwFW3IhvUVezJP4+rY0yfBckfycbGI8y5mRWUQ8Cf
e0nmPkAyHaD2o6T9seMStX6qg2VL3EvrActxjbs+CWfHii2F0KYuffq0/OKJ
cwA9WFaamgh2x0yPic2pDDDu9FSQjclOPQQ26228aLKEcZuZPiTQtnaCfV7x
V97By2yriiL3zv4QL2DlVnnkM/5KJ0z2l9Y8OIgbvG7gx25/D5cZj5Ll0QCd
GtylkgjpoWHJDWYn+/KK5ult4zxP9fmTibUU7ikHOtpFJWTKswWmrrmi42et
BCfBFBs9fArXNwzVflKKhlEi+DTKjjepRFKjskHIUBDriMEx7IWQaSxGYHAK
HjiEgRvrKjvmPH3nWpjlJxUjoGA1fznjBN48B8tdCYTRpXSX+XymLuKwUz7X
qJryrHW4OXSZKvXOR7PN37My+LYkCIgYzJk4R08hd4LN07EuQKVdBlm/34pd
rLr3vLIMT+ua7eHR5FSbPHfbs9FB7NVx/8dPWVLOJYThbKj4kyRjyecQRfBv
M4lfaQ33jaB129EIJVOdeq0IuenHAkF2hjw/CIrATaNVtv+Go7EKPwz/wc7z
ZmZ3xZcj2cuJfik9ME+9MGtAs5fUojxx2fsrzCm9eaEqbznkd+pUCS8sVLQf
zbMUq+zqtmH3nmtQk+iUkGjYwRIIcSWKOrT2xpZGZ3u7MT/MBRSm5oZvk6JW
3TQEMxItGp62fAG8yS/Roi6SWK5n36CZBtyeulcPrkF8jrvfG8419NGju7SR
EpcFCCjPxUi2u5kMl2i+WL9EK2+X53dtXgXIxskefM4I/dDro/qCHe+hWpTu
u2LtZjt2O5WUJU4K0I1ZgkQfzvviM7/jn2+GyWKQGoNAN4PvCDS486ieAGzt
/tuNzYbHwEp2as3WafN3EiYhatCFI+KqvHLRc+YB2hHSLhJNWnVPB7jV6Weu
JOZzrQULFR4GSJ06KJQaVeuET13kCpvNZcmVnQN00Yn26+NXDxXy9G2fAhoK
N675UlUZ9NC7kX4CfSYj+0UPDH6nB+965+O7l2k3p6Xy0o7UCS9KCSFEotEV
a9rdcFiCRjm19bxhDvgrpjQV/5wIohnqOjPCWXdE9yzTHzpNN6fHonOWhOaX
FNWwtdgzhnPNUA9lVSDcAk0Fo24U9xZEYR6EixQ8Ms5p1uFnwn64JXuM9hS9
UxpcpvDLYwhsCv2+18YW3HDOe+3/G8wOKc9Mj9t9dQV83686cYUwz225ZsGd
go1MeY/DbmiFLGmkBZobytb2fETgzVxktez4xDFuGMXhd3Vmnx/ac++Kpj1g
VIVZBUHHOiNNY6kHHEPRrs8lVjpLMr01kDE5fO9FPMIwmlqXah0j6wP6mny0
38tnIn23I2u5CfPxMbGHwOLnXR0e2uoK6bYLelStP3Uh7lYtQEWNWZ4jRMkR
3BF9dlnkkUXyGYDK0M+8mYiXlFv7pyn66LftXdqq7QoyxnYOLlcg7RrzgVmx
tsr3rMuY3YiJikA9xUH4BckU6LBTecTXkEbMMqlWi/bSEBKCnMvsSz5tgXDl
1vJOoAq3jEqXsg1VjSwylG1ahz4mInnTimsDDzjySJrlnIZhf7LNNLnuQmP+
njVRl5cL8KvU549lTbETcUh9UACLZCQQA55jFflqjFQrdzGl5KILaXDW1tfv
glSfA2u1ik8w5CwHrvH+XD5VjKjlI6el0X9UCufVgJZL6MGv5LsF5KLY+mdJ
m2mXhJcsIfbDFzyrQ8hL6+zCDQz77CTKzkqa25bkh1UiUyMA53wQ2RI3x0vs
gOsvXFdJ21rJPcN6b7FMY1ASb3Ce5U+Y7dCle9nVEZNOl9Hg4O6K3c1WA0s3
EjXJrCLvnee1UFhTKc5/J1KkxE7UlvRQ3UZb0WXcJrD7xAwPGe6NNMS5i4/+
ReWCAUwa/dpzoVEX+cjUS56QymKJ1ihXBulitDiBOrljj7pe07dXvPjL2ZHU
ea7V6W/j7r4/W7iKELTwzla3Tmfkr53ZNObmb2TFtN25DstR70wABjUimWwt
3nBBGcdP4V5oBDTuPpOqLbvxpQtyLewKNgn0bNHmnWgaXrG11jOLaanUp6cm
5hSQyIC58JCnY0Xn3yVXGz+1odlkwOnRZanfQzGoML8QOrSkhE5ErrPLoNMG
6DdQAqImaiR45uOGmP+pG3fx5L/J5TjDMjBZEvLe6B+qmUKZFfY42i+WwVzG
WuWzAak0uhkyr7EVtbDMYrvBzbSWSXJpIExIj3fhvsTpDbgzqqqejKAyfK/N
Bjipxy/K/c8vuoxHyBqjxaLh5QbVDkbuno6sXOiLA3NqocJLdgrHBAuUsA4T
vJ7S9HApPBHo2AM595LB1YEUOubAN/1VxFRTEu5/ymewO/bmTAWS63tBf7+C
i0eDlNVKeoJkcl/y/RXZFmAUWNdibxaLW+2ZQW4L6x2CzE+4i0yzbwHB76zW
Hbf1kRQ5UijMSSO0ALIL9Jz/G6zA7cvxkaCpHKTQLDLovS4OSFps2IBDUdXR
EeQFs+n51IjPOU7cMfC4L8eNWv8sWZ/RywZz8UzT497rkPj2NCh6j42IPjjF
j9qxWIUrxZPb7ZajJ58fi+mj3mY0j36U/Gh3p43KzRrubZnVWxFhyTpeCcfX
q0Bz10lv2jdto1fRmUthZirfZVEjSaEL4rdJKXmPBXNAegKA+44SnvGqdKwn
MtusO7f4il6la4F2QvtWSF8yZJ+KKKOr3boTGSrSC887eCyLE7HqgBI42CC2
lVFBgH8ZGCSrlNYcmsUVfpxhQP3r9dhl1RFu42fLt5PzH5yw0Ykrhg9Mpx/k
Q0GyVS4Y6fvhRzwP4JVtVJWwhWnRVopv2LVfKE7zL3SDV6G2lz5jgYNzTctp
ZuwFhdkcyBeVWflg1pKrnoFH/qQmSYjCZYunyNIOWe4fXR/4beYTfAureTKA
0B3wcbeNg0Apv3fVw99ONmThLJGmw8ChE+YRFktXhOMs7s/ZI9PNhLYU+bZi
4tOezJFyi6Le+Sl/aqLaFrcrtfC3GmIn08SvdglN0dhjLoWtMz/g+aU/4Nm8
UslX1t4F9hK9rJysUEdrbiUHtZpd8uBeQm0B7iXbiB/zffSvY5AUx+K1pL8e
k4V3n/OdXsKwnKVel20KBUYQOxsT9c+rm/fDJmQX2lxr0VWldK9LZGVE3GmT
5xdaGvdzUbwTc5oOXbyYldgcMbe4hXIuWRO369myPO7KBAyC5s7uK/f4nLSG
7j95Kf2Notkfi+wc1bf3KA3Ya8hmh+0gvzXxLuZldw5SFY0lC0A0LpCGzRsf
Q3yGccPZ42cZV1589khHR3uGH1K3u9LxxDfG3imBAJz6RomweC0tuCjJZX5U
UFywpBUxThXMD9h87htR0c2YZdR9S2WbNYgtccuydEE29v3Jz8iYZs2tmNDw
A884Q2MG8VUmZXRDhUXZdsRP4mAPbmxVQei2GjhCoxa8xml39kGPpWOwu31z
N4fBbttcP6ZQ/SbdoSF8HI+N8Ib1TvEQtiQcmY62QuX9HWPCfFbgNYPuvC1w
5/yuA//Wd57mALoDYTmOlOY1k3+WeRbUXPKo999vvdBVsxHIY8U8no6TMA7S
Y/xU+kdCBgFAbzej0qNEdYqcKvbeoFWsPTdWktOrJ/4MK1f13qi8eGl1vwxo
S3JnGa0I8PyPG4N59/MW45iSPKsXAiRHQqfUa+cExhlyy5X8UKpSkLHdxHfu
c4QW1cw7kAqG8CcryUwcl0yyS1lSggMmNTerXaWJ6WJYjMyJQCQCVk17vIRB
MadRl0Xt+gu/rNuvgqEILAlVWmhcj4IVi+qHWAzAfmgDUHEA+8nv4M0hS1U0
QHDY/3+9k/kU3NOehnPURE/CNLee5MTIpNkDxUz2B6rsa41PolKNmKAxlJTC
Cftr1ZXShQlNm8yN0AnbPpojrDU9RNirq1RMjwN0UoRCHf58VpMyQDn6+f9Z
w+qBHd5vragvW5rCkgH6DnzeXU4KRWfybzZI14c3h4pXPqfDilT6565il6jn
nFi5WOK02TnQ1n1l0/C5bZEorbzwXpF+50ECTte0GnVoqMrYzxnob418xVHY
PyePEfAD0CbnixqUXdE2B3WrmRTdapcoFA9L/VAPUVsCdOk4TPHNafPkVSrG
wH8X6Ig80U+f4UlP8gZJEsE1oeYthDKnlroog1V6aqGO4DLuaIYlTngMWYFh
4GqYmONIkoGyZE7tHYYecKqHDarOpo80Q9dqgGYgFUXg4lCgeilv90gr5xB7
nqNgDGSMPR1nLGHJWDk87qg9vjj5hDg5/JeMjdOVdZ+BZFJ8OLhtwACEv88h
OxTunuaNhR31F+pNg2gaUgmNfQCaB80d7jmvEK76fNbaj7WgqSkh5viB8p2e
ZIbCVuwjMGPQDVOFfGJnoJWCa4cvxsiN3WaJQzVVPWmksaPmY9Iq9OEvctKU
PQfZE3iYmt9RlDb1QV8TmnOVOhdzO5ZtedyyWADOWN1KsvNaIMDszFdvUvjS
xzyvzGuNfuzOHyEuxcYHaDIIkCwQTdnbK3Bu6NIzrKlUUZo33flJ5H/YTCto
mOr1jdlToBFc1B6rW0CGW9al5VozR9Ngn7f+PG3ZqE6fdFtdW5Pyx+8d2z7M
BKmnEv+mgrSG6Wpz+6UiOD9c7U4J57UYnoRZBOilLab0ULsEDF4gDWWS7UWm
/DEpWP7yeUenrbTV4Q5uzPXFaWQjFGDxgpVFSElCyknrUItCyZ7tlY1gNg9n
1Ridz4RboMRH9vlBWMIKq5fTWs4bk3t/Ou+gPh60abNJoit5iXItdWi23feG
KeKRUsHVlAWxg7/XGljwUYxtiAJVxCSfMW1vpjjdKjd0jqaLX0ksKgdYakJx
5tunpILoBgZMTW1UVIeA0NdYo7X7dRdMud/IoBhLEHfK+f5j5Ehi1SE5scif
HhrJZZtM7Obiirancuw7RLQPevyWBSPW4VD9vbTCaa6Mp1Ssm8oLVfeular2
uAdpaeKbOZi6DZRQlKnoiHRZAADSBLI3wVXHJlaPOFpuhAWr6z5snMGZcjDQ
IIf9dxBLkwdMgFX9cF8hNjA8IwU+CbjgRLjbPM9rxs+NSjWePLzC8NDa1hBn
L2BUCSQPVlS1CC6oAjTvhhHNgeNKjd7pywXnm+d+5/gzb49p0lVoAjeehxkO
V2wMPjW77LQwsBofM/3bcx8fyA4P+9z9Ca6mmM+K2u8qjNQbGAvtiK6vQJ+V
0FT1uWgwIMG22oZFqVVuM59Spybxz1jCO5uaKR9Iz5LLeyvamyz4lrsvzuvB
YqDOACHzpuVgZSciGIyJ5GRnrWRRlTkJmBrrxNdumsh6CLhc7ETCMl4X9nSf
NEwZ9duMsZfFvb9qlbD2RPK4nhVh6fTtMOWOscYpeSrUeUm/YwORJoVXUEan
u2DHIxUgFIKgEvzUSKlR+5AMbLTYSQuKZxo/hxp6q4HIWPPjdD+7uz5lT8I5
IOcNjPQGbbxzsmUVT9na4ltEm6GR7Aj8q8N9YHzyFaQv1uYQtYe3aEEltq9/
S68BG22CanQTOEtiyfwM1vFobJtCg63udGgdNaUEOz+I1mLdCmx++qzPKtI+
YdSg+6ulNGbz2AyHtDozi+SnEotMbiCeuSde6zXJ7rY6fcPg7/fGRqUrZjj5
6CW7vJfL85MOGEvjXbG85TROkkWruwXb0Px5LlEPBPNFmza/Uy4xQlqZTg4n
bFrAkc4C0AyFYKb2CzEX7+Sdh3ZxyYE29L1RctOOvA12CpivLETcLsErpI/H
qipuZtfsVTGKJ/GWlIqiFRotFrGA5mP6ZSz6/hwNv4zL1XorAhYkL0RdLl3+
wx6SfV2XX79eY/uvjPTRZPEccxR5dVoZEjoRo42FAch041wFCSfROQKe1uPH
Zuijdk4bWMBUIF3CHYjlVYscqKDz+kpCCquyuW4w4x/hoQmx0BfeeBqVL0SW
bPJuWOXmQ7dwvZBs84TQnwo2K8u0dx46MYRDRBG4EfzfGnmzbd3lXo06Pn9X
nqeCrcdDRSfUlOOVZMupb3wd4LSsCwYy2pOF/wgcgvR0NPP4cOPEo76lXULu
AFPs5bw9xWG3Ehd+q+42Mv7uJ2WUBiP6K5rpdxxfX2GTynjaipm8Zvm8G2EW
Nu8WYLrpiJds28cTitSVXN+ExiQnIUCO2uXG9zZVu/6KhQ910lV8QgzfOfoF
7DZoew72b6bS3UOXJ+pWdsJkLSAUs52lIPRr20p6opdOoWeu3Irtvu5JX+I1
sjPAuXc2wBI+PsBUTTbcKWKlpQY5nGtSE3nLN2tcjXpj39zBXJ4wbxPCywCL
0Txd74iTXrPQk38tj5l5Kfcok280SK+KrIaoAyRYSr7ebKEc2R5PKDbiHWD4
4q7oPbm4+T5TpzvOmge7499MK7luiION8Uk/OZ1Rl8X1ax8EHlsTv/NOVIbz
1TSfCsy+2bhe1b/sm/EHIiAMtZVZesQXv27qZ2mNf0MMmmbWL9aqonCMFcqe
WyMFGaFxeKr/yFqDRs7IihPYXw1UUWjwbzcO8TkTpPrZs7a08ipbatPAB4ww
AXYncLbhIT7EG194Trh3Ck3tNylE4FPwhSgrehxJVoI+BSWxFrlQAi0xxEbc
3a5QwZ2njMMUc9nvCDuN1yMTIp/MznLOoD/wQubPVFMT5/Oscr4HFEIncEdm
F5pw/V85+TX9ABGGpUSxQZhBm6MEhvEOR76VNBBMSdzL4RV8EtPWi39tOuhb
tzO+IE8Q+CW+h53CefAWD/i9jOEGp1OmZu1BBdfM5oAFvII2Xo5S2/KO/XoT
QbvhP2jn6xsYPaxY+B+CY31jIeTkZp9xbZ8OIB79+95867M0ZPzCbpQJGaPB
vS/jyFf5qMnsu5Jm1LqesFPkLGnsM+wYVzgBmHTXCIAmT3W1vUqLrIx6Xvgr
oQlqQ9QGMwxakxVVmu9Gay3VRFQPJ0icdxk/v2h9kMfp4wK7sG+l2okjXedc
R0NJ1ItqT9wPWD6+qm/floH329CqeO2YXGtpXwqp/IrT8fDgivlljgvHlFsH
p/mXex0KKnd6QT3BYfaC7PQh+ARA3cqsf2uGduI54aiqBNpCdAY2dE48QIo9
A0CipWcmAccQfgqTTepIcn+E5FMuvVC73U0fmSd1OSpdinvfneutyuqYkOt9
JFtpE56ANdhg4wsa5eUeZRTBS/Nh7kmM2vkufUTsKuHK6E9dtUfgmHjnl1ZO
qR8y05wWcXS1+iiLDAn1vh0POettDnNtXi024fGfqSxRMnU4EN2niTYpZoQF
YoK+XB2zYA6KK9ET87AohPZrzwmCGRvw1p5VEi6kNWnZWYiZIeEJ2i9+Mv13
EVRg5chw6T8hm2kjDt6r+GtKabZx/XkSf/cq7V4JJjtcLkapua+mRecsh2r5
0QEfIFgMgcjJ9qcBT0jy6/7AAuJnLUXM/5lm1GIuVeSwJi7hvZDNFzArQoYt
4YmyYOFQ7cPAcnQZKZnGOjL+oVJQdbPsOgJcRwVlV+IHuD5MYrHv1eYIdoaz
oonrtUpNBLnf1U6j55145x3N1OXlGonnVU8OlexiLDjjIWQCephBB/7z7pEu
PVo004P42o15Jgggw5SlYtL3DvALqIiMjHfOvGsmy/kE0cTewlDimobqYVZn
cP21skLhdMepkepkvwsD2pdbSQAzAyGLkr6/+YFcjKzG90Z2wbpTZ+jqmgg/
lzPhuU2331ILf01EYxrcTnWkeG/TguZffXTQir4K6TkoVCB8rMT5IXc34hSt
wfeEiZaEldjjgX1r2IXCO0ny4aoJ7Und4DjTXsNedrPcfZWieJNFPzyrfrpc
jVWoGiVYOiUL2IVOseGH6S68Ebs+9shQqZ0pQk7BqVP00RFXTMQzfZNyU32I
eBcwNxFr1hQ0+KgDxwHTh2UFO29RE8zjRE0AOHJH42Xp38B62Rf0z8gMh+Qv
SSFcw35Z3wKXq7xewgs3g0drFDebG6t556oIT5jbQ4F0lDbSB8fPAow0pQSV
XT7hNO/FpHnzcAMhCTn/6uN0N9vRQpDFTzlBXFnsLKxIixC2qbY4l18kqS9B
/Th5SPhWdZBg3l0BR5paTA2kpUEoJOHTfFbRuYq6tfhVByGiPZ2V0L4csTXE
TEBx5jSwu0/bJ9JNFfDeS31LozVOxS1RqFmMhhF7eJVcvpk4jl+EiBeEsLHL
nOoLnCyFLXyD3T+4pT560u46oWga/VC8sySWws8CQ3NbItTLx1obkpjTJ2C/
Ez62AFcnnT3AJrYqveE6N2iuSJ49O2M3ngJsE7cjzrNQjmz3hHFNfYc4mpPF
cZPiblM5BctJCK2IuQBi658TaApZ7nwW0Qw29BW5gDR4acPASUxxbRsgyKBz
HtCuni4eFTBTb4kjUH0rHC0ky9fJ32krsgJ5b2RGVf56+cFcrp0lxIoTS9Ig
TQLpIhWA1yBca2hwf8AOdDNX5gI328sgjrkzwz+58SPRlH5bc3aS3fIvC88x
RjXW8M/6ajCNV40rQdX9YKvIEXBNaPucAy4/ocnD//4TGnZOjulZEty4K9i1
rbzHu0sPy70+WJjQo6HFz0YdtFypGeUPk1ZR6TgUgjFfZVfCb7aXwmsFClB7
/MHWecrJ1w2rFtV1GlefVznU7RYh8PMy86XtJaPW3AflCmnJVPcuvqALX0B5
bizr9hn0snXKpGdHY+Nu5+qWZwUytH/jIFbRLvE85SwCCR4chkla9rTSz7Xa
XCiBLkmjdkcpxas9mgmZ51DDKdjbvOjGkj9v3u1iRx/kRaXNzLnxK6Z2Lz0s
h1Wv3x1q5AtEB38M75iUMYE/yWTokG/HC6z8007YIueX01q2ZYlydhSuBazY
r66bIgR6HZj8hKjO0aAqVGJiT6s7MplcWxwzNf0MGUXLByayJcKT+om5TfyE
Qv3w7W+pTjWTfnncWev77AFJipuQ9OHMSH2xZRzPSn5tBQeDSEamkayyiNr0
FqczlID0RDzjqM7zCpgL51XlRD4Ush7ymyHEknH2Vh2Y6JJowE8p8Dbw7sUm
eO81ETKZT8PIZtC6O/2nGllgWLL2gVQyY43RVo+uiiJd+R2irdIuaNPV4Rpi
8iOBs0hhxxz2wSh4/58eee17mH6L4HNJrp4sOVjJWapSlvnDewiEIH9hbAXy
PAI9FJnnjTZuhpjmUHRtl1A8WMBy6APg1lUntk5XxBaGCSC7oIgmGkJ0Qgm4
XBKH8zTjVriUR2uHfGk/NCpG26DnKYX4hCTSDIR5aXBXFejxQTdJpUC5q85z
7OfvqIai5QvMlbUFDVSXExYN1MgJLlJuLE39hvyCHHlI8/WwOc+e3gZtFdHd
mNCBhTqAkTZMbiMdr/TVwQ9TqU8CT3w/Y7oXZ45ui7pEcSa8UUGZFi0I1oZW
dwBtZWSvcb9Kiz0Floava2Obq6+i4hTSVSuMAPaN6jT0TKiRtTayEKgIFhOO
w5bLNSaizv+qVpdTFhC4g3DDKEtVxaUy7hVh3IkJju24/fUbOviHL7Ag+UzT
pnx2JS0Zoid9WCToVLqD0BQQnkUyJl4Qjuej+SJYednjeAwOjhZd6+LNZCZo
DcMP50Lc/zeoKv9EhX2THTdKNVXLzDWSKnvjfVVGaxA20ab3q4a27tXvvqE5
Ne1541JviqbDb948c3F0k/ZaNT2Q1Z4Egn/3ZakuUeB7xcqdIrEgOIQAj7VQ
hy3cl/zxDB2jRmXpysWVkNcHXcbgGeVATxIUzE31hLgEFq0SLyx8iAvseUiX
fkNLylcfxLCrfbFoHlFzV34NlZVgjbYUQnl3Cpfm7ujKxFY9dkbMDkgX8Jju
p5sFHZfCGCdyal2VPOwBI5zCI2BTgOy1/YOLtpapLZFpvk+2of0yKArjAyId
lWjo9E3gaAl/YGw6DIcrcRigvUsdxo3oEflE5gFPuYh/J7vcXkTJhdlSqz03
gMBUa0eWbG0YF/xHjac5OjKwFtavUVpqBXzcLVSVGvmyodsCCPBlN4siQN6n
b0TUCuXxujkSCGyVVUTMdsRxan/8ExJOuBnLy/F+69Y6UTBCNekgSZTNqg1M
nDXkbjLPj1+EMmCu38R3UECD0yuno4Pxm1TRhnVjOgpnTlYmYjilPuCUd9NI
VqsoMJUKQ4CWWd1noA6ZHnVMUQ+zsixzR8p61rDNrwpSMq8hfoqd37QUCES3
nGDnTP9c1KiNYtM28gXK4FI3fbfWCjE/LcUqiMBCRxX440yYCXLbU4mifPcZ
MhjjbhcjnOdxdkxnEje2mxk2PtCbNoDWwpgoXwCuXV8+N20wr6i/UF8ujoYS
ho1G7CRBSaJptcLGMRZxGzWUlPMv2UKW5zC2ieeIWjv7YQtI4KBc48uW6Bx2
IXduFttk37G1jNVoJDNPiiPupNim0fIsp8Oq9YldP46R2rNxC6d0gBE6VQDN
zCZuvrSpyMSbyDQlJIroNobKJOzfYhZ8GmAkp5PIFyvtw0LBqmWuVkZlE4as
FDkgW2JartfbEr9FBK6AfxalOqCzQnLzJsrY2T1hUA7MWgQ7bT8acvO5QPyF
jYpWt2LS3+4ht4YcNWfCJn1Md3UzEyaN34Y7vqxd7HwHo7Y3mCPEyeiynNfk
+K2chS+YhiMrNcEUCjRtR/eokMBEgU9XRXGiZwWn7kxa37gXgBlynfp+IIad
KrbYEIv/sQAkAMYjMdlt0qY6vCyilu2HQFuHDkcAKnPf+viZ4lYwSSJV0RsY
K3bjsG7ZKacHbdTJqWpxN5Xj+dDvIzlpnTstJ14DBuYahbAXSrbjJ8KmgCms
9cz7VJRfBkxPEWuQ9spQevlvBmxZgE5qPRlLqf/a+VwRcVUkU3HTgwvPPPtq
4Bg0zB7Uy+qkpWR2VbzDk7yIryOrLOZHm35E83scu4j/zzciV7MdcK7PS60H
yLktqifaURmwychxN3qnP6YUo1wZg0tEaFyCDNLcOub4OC1PSKz5ylwHOe4A
Z2imqPIFRn4Nh45bPal8l7vnSETUKEAp0U3qCxLZEuudxy+80HwKxLhiJRrO
133P5FRfJg2OmRslL9vAv1B026jz5qhzEQD3Rtg9WqqQGW2jbbAiR8SRHASh
oBoNFBJp75fGPLrdFD//oRspRj2ZeYxFLfbqMqZdchqCrmSNnUuIH4EzOkKg
MHniJswdp/6RpUgpRP+UF2nDaasu2J0+Hgpp4GaBSMiToN9hhLpvp5zJhh9K
Zn7vGNQeNGUr2108RJGDYWOmN6VCDB1M7fuUW255eWzeYgaMmrdErZ96/I0v
auwFkSHMExdLBE+/hbnAb5NR9FztsbTSZooD2Q+/k6AM45w7bqFsiI/4u6sC
u/B0f64emFaaQjkH3sVLdWDG3FC+uqGzF9Sh5woCYtV3gbFZNoRlr4yRy9Cn
cA6ij3cMMr/W6paV3DmVww9GcBe/Kk3xIXjgw2ZriexaQDI0bxFkJM/aCFS6
XCI3AxbwFwJmtm8n52DK7IHO2I5DKPimrC+VclHAVhaAZKLdY97X8bM6DV55
BOJYROHaSvL9yVmqNkmtQt55G0whAsUfgNLmwQZ5gQ5gXF+KvLF9tkzW8Z2B
dWmrPF4vkip/O1llGQoIZygdgo61mh44261lwNrt13Tv5R9FpIphK36yv2+0
WqDPjsz+orLGRKtX5hGKd8ZvzYB0VBKt8ryLfCxl2l2Rj1Yb39L/oxxTqhCO
AVvUevYIr9e/iL5Lk0ywpvDaqmTsIFD6mtORx4r8MwoT6TZ+EKBKqGXY0r0e
Zzkp/fIs7w3c72LTWTaftd7ypYnv/gDOOnOce5axJ1ZTgqu4YvWGbGo/6FqC
ItoDoZ79v5AYP7NeM+vGJzWrw13pzUWDxUBeBsRy+7OlZB6qGxjruzx5Xqz1
ZUphFS04ZtxYGMsHJTiXquJQ7UrvvZ/+EYHZ/OF2jr34X0c/N1rkwDLHoB95
CVfiSKLTqGnBkC0itWODWF2XgR5syn1L3WxLRtocGu0boeJR9054YTUvGWTT
47r+JTtB8EjcOSWJ8Q90kFhxZq/yc0uEPb0UvdGG0DDys80/waMYo4rHNhhK
rNGi9HdEjgoru0phxYozOKOcTMqJO8hxmfdXI64L/rmJjUs5lIjZdc4YvXGD
WZjRbrjTeNt77pvQXe4Ukazka5cpwsgKGHQcIglTH6UN+CiVeyekSYy77lIc
g1ksWsHeR2rpdM8ATURXOkAVpaatboJJ4ZqPc9eryoDzkV2HBRRfH6T4Ij2t
9EFn9DxHse0fmcxOe4ngzAf/9fDpnDS+/43M2AYw0IfdsK0tCop8+ia3/Utg
LBMcvekKZ/3ONdaz8nFCht+QwjCiGiU3eNR9g3PIvenoJrTEsDo/nXFPFckw
LrtIqYwcVCkoHkBf+02qrkXQjiubzOloIdjkBug16m2Gl6mxnT3lowb5R9Lb
qi81tiUudq/T44mQghvFYrRx9xGel6sKUIW3BaUdVgcHummgHku9CiQgocdM
MZe0+9xABoATZ7jT9xNJhSIaBPRMfaA62SvKnxMj+l655/Me0WGvaICJPTvx
XEIrqNVChW3AsGvdyId2GyziJOn/6/2x9PeMNQ9whkD7GdY/IvRf7At59dlX
EbsEOllHyalHydIhVL1KL/uDvtxKG6dkB1uwsdxF+z8E1Tsz6VAw9H8q5i+W
9riigfPhOC622cy8kTm9DWYurmsxk65cKSh0bAIilvAC6TjeKjybTp2HYW7e
K60BvSzQyTSy5g1o48dwxHqUJgdxSjbT2J2x7ZGVhgzk1cyeLj9cKeZZv/lM
O7oCk1hRBflhKNzPOrW9W4y7GKqEf328lzz6JDfdNu+vIIkrqUTwfKkIzPIS
MUNF28r4mxBepMipdiOExCq5OJUzL80xSuVHvJRmctRcswvi+9GWAKbltW1K
UowC3MV87yCyuCxztpR2ulFCbWpvgmKeFl0xEKOFBKproGFqFeI8t2xK+2n2
DqpVji4vQ7gve8kLFl/LgtS4tsSIwKhp0Ips2GOvQVQM+KL7KhIoYbCbGS1g
gIOBf+cea8cmQFibqWv6+gNUuXhB4dIpXqpRJNRgUZCBonkdHyDksmeCLcEp
YrWjsYdzdlsoOXq5aECXsfCinVIuETV/zwpLLqJi351ZT6flDNBe8BEODOIc
C6DfAI30mTKGy7zMmqQi0WknwetnU4HS3GK4bXdgeTXCnuoB2kqK966SCT5I
fG7Sa2jy3LIrMTWvgjP2tDFWWVuR9wCw0Tq5CRPaPVEtEUXya5THWCdiVFZy
jBW2ynQm21C35hwNkUDyxOOhqSCJ/otoVHxf4q0eGKTYEPBbXtktsXn9X0wf
5ZBt73kPD5czo6bxusv4V2vCidaeLTjo/YEmGSsU9uNeKJVMJ4gJ90HWGAMU
Yyqp8o5U2bopmBF0LThFA8LwdI5uen5pgvSqMexuS7+ilT1+R1rITUcBcirE
8tJwh95rQvB+PkBbqWlaVlF3jSUkrV2AQdqc3NyzpVYPplTJ9w4wR3iwrYUX
iZKKVUj74MKU8eVXaElXQIiewbBul330CagQNb5fPJGzZ6AGafC2wV9Lr8tf
L47YDR6kCJdqktbzJ/zackReKNuAG1hx6YU8+OgQYKonrgPahC1Jby5VVLcC
q+LWr2kPN9xcdnZYjqY0PH0Kuey15LkXlOYUlUaS29dF4pWEB8kuK+We0LtU
YxrwnuWAixESU3QgUrRqAfH+pvJv+1XgVJKbPZd9vlzpmNhlV4U0W53it9BD
QIP6AeD7b2B/q4UZrMncYa9kWIpQ2AgqCs8WZQtpzPA5zjgRL+tvY9wEZdtj
s+DiiPK/2W1v5P0QzAFMDkJeUA1nksCwdJ5o/MR7cFaSGe27k/lLLrjxCfrJ
3WLnUm/dx67Ac9MkXB2rzTi/omHCQdEgcApwKfssMCXcD4rD6PJWUnj8vdvT
hS/KYZY2Ba6BdUXW6surq7xACSv2wc9TKsuF2XndJkNQcdJsH8TzMen3+n79
zjoL72iM4qUeV6mhlR2cRWSdkg5jkrjA0FVMwUNnUxl2kHKmemZ6tNYSvbUB
iWr3rtI4HobXbX3pjaAaZRvrCyo7uneymBHsQrGTrYmyXPQhwmXSH/EhhQVE
y28qrvAGH7pnHrBTr3OoIFVk4LZAy+bUdfD9eD3SDbwT5lljU5x/fmUmy0S3
SAn0s2MegVknxMvcDOf8922K2w2PXs6eiYop9JrQ1iJRVGtFcPrJi8HQcWel
iND5s06DZaZf3mL2zfnQhbXMkGdz6axmSONz31atcU7M9TZu5algVC8sfwQP
tsaH+dGH52mL6znduQAuTVihQf1aikVU2dEKsVgvT2rNwNBKLKwca9Du7c2Q
haS2zAezwo30Puj1GiVUTPg9yeLYuA6m24VNkAHE/3pZeX5zGTUJVPYIV1Hp
kGG7MHoLHPSjrXHgJ2Nuq6sBnLfxsVUsQo4nuPkW1R74P7fzyKFO+hdBPoPN
c1xH2M5A3u5goTzzSdp4AlbgeVk/hqqpqWcAAzXlW4nspWhYX5uOZ37cmLjE
jgiUUZa6hucB8z+SiFlXC4XZW3nCxE5gFbV+emzaJBdyD8Si2SAE+gsSoLis
F1qPto32xgdCMH+Ed/DVD6KOk+R7qc6Cwl35W4KfhejHvj2AdynHz6LDssUN
KaFLyWY5+39eI/Py27jietTRXAOEza2wnFwi+6vJUDzoBXbvTansZhz7/abg
ok36G8Ie8Nb6eL3yd7ge9BgfD2cOU3jMGeWqv/o2UYnNSunAhG/Trlj8Ope9
dBAcrJ0v0VVY67XzWZD7Q4Rv/Yr0DSbpaXLIL3/7uBXjjEBef3G9sMTBH6SS
Z2nTTP0K/f2APT6x2T1R3AAGa/cvN9lDh6fCuMz+t3fp6iVdA5Xr4F9ec30N
wBpJzOh0jTLkYJkVGHPR46Lbz3klR038gW3XaRnXSQ9oyTcTtNscyavAYeoy
bltsTq4MXfoAKlYddQDee/mYy5caiOgA+7rANjlv5bwkVhDjZSPA2HIMDSN/
DT+yY9LjPflDCQv0ulk+7wqSdgeW7Ij602Mh1L5q58yhllAm40cRyEm11SY2
KlMfLMSWCDf4npNU8AyZMSVAu453ZwT60qif08qbTPWDQ6KAl+Azy8jaHvOC
8hfjD+ElBvsC1rpYoAcVonq8E7IjvZ2uKJNys3BXnXcQycKjx3BMsEeenLJ3
YMrvZhGC+QM4wtt5BMo4o8m0MvLUg6R1obpdhmrkpgkcvGHIjtK0tc2f2cA8
yaNZ7G+JK6IkFM6eA7S7qijhUPD+HmawvEzw8NueNAg782IXhA9p8AvaHdSb
neFz4+F2rv6F698+0cRfH9Z9ijNn2HeVXhOhnaQiudnRrs5xBeGIvQbOXMt2
pawzClkts5P5ls4tQfGbiqepRNk+/nULkH+xqTSWN1GFvMSFuRkQPxGJt3Ip
pzev/FwVdGDke3JtOjv786/TDU7Ik8vCFkeeLrTCyZWUmh/r1nMHicWbf84p
Y2lG4VikXTAhW8tKKFPeTERWFJEu2TUBV7YNxr1wklOA5/ZITsezrzlmg92c
aqrbgPbVSFcCEa+y/CfBoajdQoFWEyweEwdjhBirtAKAtKP09doa3NwhSsV7
7cH7Th3kRGhfcI0EkNb2Kbr0oZFyOT/H1s1s9zGmWnHdj0WCKiiRwBOW1zMT
ljxKhTozDLd3t22q0udapVfW3sE5QiaIN98GHQhJM+o0TFC6nIfIQ56zT1eB
joHm1V5c5CybMJyLcxQ7IzUE06esViApxKRcxAj4xrZU5xV/3R/1Uch/tAY/
RLWPA8dP9pWMZRaOztu89JI1yc4Y/bfFV93qFYLea4m88Wt/rDXbZOPtloza
x5JQ0PQpjalSFEu91FSy4PT9ImUhMrxH4A/CrXesX/efLCXnyCeJyR0GJIQF
84hREvUCDIojCL+KGeNgyQ7Ff7Zi9Z+XKANb79lCu5EyLiOOQ3XRPN6IIPAR
tPkU50mU1gQ3DIMUP4scAWrUXyaLgF7sbXW5AX3b+PfPuMtUwL4/o9xDehvh
y/da8dez4RhTKy43FD5retQ2NF0RocyiOUj/aPi4ak58NF6bvz1EceLb6mWY
jFZZeaaKUokcsxSBxSqrbNLwB+i5+dvYj7cJrAAtZiVjnYMl18dwX/JVRKTc
w57+nsPIm2GFmmua63BMWsSdph/qY9oqXS7CqDcVRwb2hZ+6/xl0bvW1UVse
4u+vLa04L3bBJ1T1ba/g63+qinuPcf4qIxDl4FsN/rDvceYrwdP6Yz4A6Z9W
TXEkbnpFKqGAPhIsQu7p6MR/1awdTNccXBJmSF5hFuJXMc/Aixsq8t1WqkbY
T+yIyopWeXSBNBkAaXpNWN2Y0uZFJU3VUmGjFevEFdZ5EILanNXWr/QwuhPa
qYpkJeBJ7VQBGUeIU96CNLiDlyHVyF3NBsVC1Ij08fRRRnEJ5iTXiuRIlzcQ
uHQprq0p1lLgcTbh2gGLMR73S/iu8lcDHwKJDg6hM2mpy/oSFG0qCJdmQqTE
ImvoB0k+NInC9y5WU/y/H9wDTf8lZ0ZmjFmwen7PqEzsdQw2VVmg4ku+3WXA
6nrrqxrqOlRTIHArpwFsrB7LbajQWG82YYc+K+1iNwUzqZfFIpqLcJvRkw1B
DxqFf2UnGF9K93x+OfbCL2OmtAAv1LjWPU2M2t6sS/r2XYHBVIGi+z2OxsOB
GO1sntYX7PGEWG5/CN2ktGQGZNzZYTb184nNcZ+/OFOek0LKg+dCqOaMPDlC
XCZQT8BlpHQzAnikdZZZU/n4+mqoNPumbL4vP2Y9lRZ+0uOyF9XR5mngJr69
WvFxLx5h4mGrlDvmC1GfkS0wQS1wK2mtmyTqyASTZ0nSxc0uQ1UiJ3mTJud4
/JXnNTID4RmeMqiG47v8rdUjwFJ9WLQYkN3+2WOc8uSjo4b3hMBKBw0xOlcB
3n1gmfQ2XfwzbUkBgk4cmJOIY/LNwqp+3oIb3Dhqp1KaRLQZk+KzuKaoiyX+
9ZX3r4Y1pXPDe1p2VvALmSCOhjOEoGQuDvw0DQsU5cxnxB2yNkQ7vi4NENvK
vHJqyi5ejSXRpHcJCc5zWPwlZ3gbf1BnuguJ7tt0W8dna+HT2wR7a47m83B7
dhu8TOx0KRygk981GtFWJ/itb6hPw6t1FSil0DIclJwfjRafQlslKiUBQS1h
/Zd0MuaqQjfEkFZcaLcVRChi+7Oqk3E/ictwS3XA75fdfnx9L94JDANYvp06
1x+gV0hmyUpX6CtiadkVtPBqRRz2hi5CVFrxghZqLq31gradfSuH/aGiJsN4
tfHXQe0nN3HCN7DMfIJCH2jxmvyBjTexoLk/4G0D2P/eTkQYSxzvpR79MscF
kshk9H6Ny3Myf78wF8kesVJLCEtxo0Ni72D8Sq6aRuT6p4q7KOpbH8B018xC
gRcUhVscBzsLFvKeswEiXD4J1fffY9500NWPNk31EHRKGKWcFOQ9Sz9Bx2IX
GCySnltDiieee4HYV+L4J0AvFZ8Jwd0P9VlSLd7rZG1OoOm+EtDfa3enCGiQ
T2vRTFremH98JoEb1pm76fkPQrxzQ28l+8f7Vl1zrW3lr+OXENFh5D4brWxR
A5lQVqRRKDsR+8Wpwmb13bWx8TkyBi0hFrrz8/CoD9GzPbFJUeYiAPqDIucJ
URg0QQ3r8lCMMdzrrZkemoYKZ9+DCmI9Xy++Gh6/b5Aa1idMflt0Ofhl7gKO
QhbDFWgMA21X/ianXJtGkpF+CWlU4L9QPVsHwzVLJK0QlFYfRDJF7qVr7fIW
VXwbH6zGqaAVt6ayB4QNkg6O28gYYt67qt8IWmNnOm1BswWR6AbFF1Kr+1GX
bkqUCBuj6APLQfLazTo5VRrohpPO95dz/dA6UiPLUrNOYGq4wdG4J1AvYoDe
loNW3/i+QfjC4uktp4ZVk2/vMADNs1hcQ1qNno+UpkNsM0zOYPyj1TRr5otK
B58xfdk54WAwLcMEF+mtAqfMtxuVirOIBmu9sMtGVa0RCMiBZPDkTpEY/Ny5
Jbe5AmfAsIlzu9UzYA6Ci+63vhtd+VvI15/zer8QrY/LNUUSJkeJLtJXtvG5
JyzkTHus7jBAW7MyV7AUjyarJyQhRA0hrqL2L8MmVIxXO9LzyRGHrhp7Tj3o
uJx0OdF9rh+cl1/rd5MO3JDl6OARUR5bcSfWoBQ9jNe1TLysDLDdzc/CRTNO
SxV3b37WBKiZkEzpBNXQBYfB2lopdqVigh+95XM4ZBBIBz35XofsAFn8RoGu
0fKa6ZX31km8g7cw94WdwHEQLeZRv0pjRrt4LQFyn3+EmlHDErNyXN2x1uaY
yUUyIqyH0WSBdIXKS8bU/2vq8/L5SzW84jJcN2oF/XSfsWQvEjdRTJeQMOZv
cUHfmy90bGaGmfvUPKE54Sx5XS9Zm5cJYeKZ0TEP6ITplzJv3h0FlUbm3+/C
zrdTQDVNwWgqywEYecfki1Ig1hkx8ZI2isqxKdPnPFhu+dTBEIpX1X4XSNKy
kiLOenhOePGBwy75r3Q2oi9UHFaeRuAqhus3GSVWJom20NGuxP1xr/8cdzSR
0BW/cGYmMYk7+tAeJbLOCw3JovohS2vyWCWKtad0IoG05druZbSBVSCw8VDi
/OJAwZRT3ZW8G/XGC7I1CoNvubZL9m65YPuhTluAqtpTjuvIGZTzlMS1qOCS
sST29STnk5oavmNmNa2aPHhVwhhwl1b4q9UxzlfHvUmDmv1LqcBw/FVlHfEt
sPwv8ACFKEdkDA/f22QrQEATpX+8Sd4L4jFPaonnZG/uiuvX0HwMfT8GnoDs
B66NvAF7wNdaVWQbTcWsjCRJbkFWcdDaggeECdVmaPuGjVGqtCq9lNyfA5qA
Gs78+CtdJgvxkoDIwNeVehBplmN3i1Gc8+UujE2bTT+xamJnxSHAjdvZAdt8
l+JZLtDDHjkrG/GFiKWA132x8JnEBl3eeN0buDAIWBxRZBWXgROpHQYdO2wL
6P9xVjRZIoHy2+EkVYb8qpbXb52hG7UHCa/IjBK+wWMy7HaDijenI1UE+yhB
skYKPychf0HbSFFGAX6kLx78BL4SuyB4/eD9somMMvs/MH1xzOw/FZ/xt951
/aFTJUbRknhqRdlL3Rox1kTl1QiUXI2r2wPcG/so546R0JRDUksVoxiQ9P5o
tz8JRPbTsreUFV9fY0MEd5IAvKoI61Qxwpdu+No6GWjX1OpBK71ama/yNXOJ
2ZRDRKsX6acKBJQlxUwqOzi/CWwQuHzuQHAlOqU1zLFvTMgexQsIWHii/nhe
lKdeGUV7DtEZBGOub/DqlOGPpp14LEzrlBMQKo+k4oPwHCUbKkq7xhpG10ZT
Su42p/LJ2yMsMXoOHUoquM1WqfA/PlIJHnsl0vM5/QDUt9Wnb2adyAjlnDpt
gQFipUzymeyja/4R37e0m6ttVWgMN0MuSdVvlevBsOPBpF1Y46NVedpyuggP
M8+n513cQ7SCWcPdN00Mi+L/Xaz9v17oCOMUkYdACFDKiOzEaAeKd0IpPbrE
Xc9Dsw3zKbS8Uvu5tgrMZcSgZ8bL6Z5slfetVkcMV5t7e6WY6/m6FlhtGnEF
AodPPglcNIEWNpm25qpfYQce80L4yUFYzeWnCLQsg1qdl/XuXPc+3ChXlDGM
BqesMw2d3VlmdRAk2LeuwfXyHQYMwIZNvc8gkLsOSM4y+ETwnGZSdXG/Ta22
qmC6zfkmQ/H5u5k3s+LEPAqJKdN9HPgmULJ3o0TbiaJ92bwUlGhbqxxlx40f
nQRrh+cIPjcj99wcAIUqznTSE5MCB5kVRX5PiOX1XhMoXdrpSFX3U/ysu+BV
TRmvK4waEUlCryKjRffzMBbV/CeFRJzjk8r6O0tvZtI3wPiZ+UtQsX6tKFeV
kyeUJKQg3JicYMHxG7OkXG/cjZOIeMBZMFSCN73GIudRPLtsM7YIRCBinViq
bg5IDdw5BuxPK9SzAPtLsN7RBWCvg07c8ozt5dCz1dTNozEXkWmJIltxeyRT
tGPmbYu8Q4KDLmpQH2+CZwaqVbUUfb77e+Dp4zkiALIziqFC8iGnEd9yxr2O
iTAtcnfMnPqgbHLFAg2jD6WRayTz9ZD9Uk9N9dUrox+mxBBnk1RKy8kbmQrJ
CZRShMjDEJHkIKcoeQafSJ9zZ1jG3Y3nEW7ShFG4BEjZapaVHlQZij+jFflv
VyVZ6WOyIyHwrfYgrwj52TZ7vXuUD2yqRPi/N1JmCpsUR8eqQEBnl2KZv3Ny
F1IUmeVObU5kxO6VguvZWjBZ4xgHruIaBZRRh85MUy55UKgfWJHCD4OSsuHx
rdReN4Z+XcLnxe9JztbAHaCVRrU9khjvmWO8svRA1+HFYSITU+eCGKe3ipMZ
H2Uk60r4MLptukE2FVd5rClPaMih/NKVwEdZuWoh8eniKo4yJDeGs7w6cGau
EcHWTs6Dn3PsooH+Ghqw5usWGYNIKSEeVOt4wGq+m66RlUnRYjGAi8pT6bF0
Q/lRtjlQKk+cGNwglWJj2I322Gs7VSuEXRhMw1La3fRslswKd8zkCpdLSoC/
+U0OMCMrgE5LSBiNeU9RpX8gY9FARKqh6zn0JJETBu///k3BYr1Fvd2Kc72O
J6NAB7g89PQ+urm0tFYvwbycqZhP84NNtCM3iouHB9aBAa5jO4ha/ode1kK7
hBQyZsfQOPjDdyZQgOd/O9jkWg8uv1ohgUEPclcUpG35AGVQcsiwHVRvK/NY
JFj8fJ9PWsJnmegYposHveqF5yldvqWSAKJlBETn2W7+nCJ6LXpoYHLaZeWA
cVP5w9SOwyVmJxh5RNo085o7D7UJoGZ2uYon6PqQSyNeSQj5SY3myb36luQg
X0Ec0mwpFV0MFv6m3FNl1mjo7Bb0lbfDO4yKhEDPL9m6SwkSECAkuGluxwr4
aJGR04MlSDJsxCZ/5fQyuYubU+vo40ZVowY0PF/CCFvmFt4drqzSJUeRmkvs
aHDObCzX7+kXkM+GTml7cOsr8t5MhyR/l1HksZ+CQUVeKTjOP1LoDkBxo0s4
DiKjoit28Zr0Oam0JYBM28B8OVp5keiqf9TogISYqqePYhxVjoBxVseCG9MS
YgP1Rp6HE1MMupbkxxhoU5JMw4XLYu+o7yFQKIG2RnRWd6K8RFf8IJK6kJlo
b6yQv+JdCRjYMbfQ5n7R3JE8tsVFpZW3XPjRdquyXm64Er0ep4sQR+dfQNve
v6a7KdtCIieWgwLC/Gf/+znI5Sj4Jt6I//ptEzfQ/mOyQNgXSQ8yVHr3x+HC
1O1LQPXR1/NjBa2OpQeH6C35a1lOtXzhq9TAv5RmNpUCwa8meL6s5YapocQf
NF2CoCqgLYMDDRwH++qvp4qgp71chOwI04ZMv2UyEcaFkfCfYdkG1FcKUplL
gVOCR57/5Hzqnmy9PHI786YEaYHbsVu6ld66lqR+XObV5PupKdV4/BuO+lQx
cs9s8VehCcvYGM2idRENxpCwVx8yqHNwlgvmZuNikhYVwYnnsMFGCwqIedlm
LYtIsh82UFVdEpxnS6AT0GMa2GLAtw1H0+tiAsIbAPX0/qa1xzDLEPiPdppm
Q8BgtzRguqxk0uVmQidz3AEfD4MhVPaaCk07XOdn+eNKz+gwZjLsaVLcS5bp
3KnDbYU36AH6+YSYcKcCMRGphIbBohyZ2U4fRdXuj3qUpgDEctCbSU/xgkiz
NvNOEn2VuR4cqzv45c9k40tOnIV0fJPCJMcTsELTZ6b+M3BIcJ6Gb7u/6RGw
AmOa1qGtxkFYhDHRTrGQ7ChER16Vr4EbQMYW9IqcvwLuK1w3LkqWmKHPEpvJ
EpjH1lZ9TtIQwB5JTagCVyqjBuzn/niHFXdEUlRyYVBYhzXJC4uGSzBHmMgE
XZHWFvzB2YGCVFkwIzWMWdpP+jr2SHuIZN3yLMnaySaF0Gt71U3DSMsIFEoM
xtUlwEIzSpmv5xOb4zAR656zxhpzW3TIpqm3t6xnvp/wOgEeT+y03k9EBFbv
Flr9wnWjCAG2BTu3G8NFa/7TCLRYBu86L/jz2OWzPRDyfM3rS4/YkpstUW4z
Exh7fERLNeavfbCdZAqLTqY1MKGYz2vWk3FUDv39ITE3OYYqV4bNAZ6eC+6U
tChnArLrRh9QTduxdGLDGt7ZmCDEKhV2JvDvZQytQJ6gvqyM30V34h1oebET
PM4WVSuk6l3fm0KbmPVnhurjak0VFEWqYiILhkqAmQFUT2FSuic8t1/V3McT
NPbcCREOdpEvV+SCOJfd51kwq2I6tbh9wgLx295tIbRUtcO2gXeLVkFageV1
6CXDsCinvlB0I8kRYY7GwnFAFQClHvoMlv1NluXPgnPDD+doJhIxrrt4y6kY
eY6VjGZCKDeeQvuPSvkpi2K2uJcithTyFMZZcoWrthtaxUO2NJTykXn8PAqL
Uxi0JvSi4G9GaHVyvCwQvJXXCkLA4H1stRgkZvlBG40qREIflxF7aG4/y8O0
5UOrI2MSWVWeqrlHcPsulu9GDV0d83awUblUCugIANwCsrFgOXpD5yBeOZkQ
Qn5TjdfpAHp+uX9cVvBeL/BgJhjUqvMoq03sxLHo0sejephycjPopWjOfK1D
TzqyWNij5xntF2H8I9VVidsNAOgPnGfn5q7h1uY/JSPddcDjhOEF9K6lMANR
r6KaukhuOVNJxSGVKktYOBp8932NWnNoagC2paR6e33F6gfEOU/P5qoVt2Jg
64ReJm3MLWH993Dt0jFWcrXHoFxb60IbE/ZPjUOXwTtddLwAP9UnGAt7ByZ/
1OqCyIip9wBSE1dl9nGsSAI70Mu79ENOJQ7y+AAlkp4lngEsDJz1jw5s7w1N
ccg+OPfOs+cQ9wRfhv3ziukGyRIITx5GiT9UpBifoZE4fmf0oZsT0rd428kp
ocTkoRoQHOKQ5RaNQpglra1019ice64Xmm4EFRhicY39KUta/8Rjac2xHQoT
3/Wl7XHFSSV2Bh89kI8odasX5u1BlVTa0qplaMCLXwErSQviO2IB4SJiaetT
sHyQjHYDSUv8Ucozq8kl2+c9kIjeRFOAUV0L8ZG+FzpFFdj26SEzlaaC/XUS
X6tXWCLuoGf6nnTJXpBgRk1IMesA8WfhsDp6KSiSQb+kIkJ2WaTDFe/KKZZ0
Ak2VozdK/jepCHQ095U1lVAICm/2m1YXSbhzdZMRpRp0UCtXa5OqHCRlJYrw
4YDpgIN/AbTgL6uWbKWace/xAYhNLtpnRwfFQAN/VUTNGjgGVNOEoIph6rm0
nBwvQXE85Q9cORngQuvc43g14Uai/MxyzF/FHjZ6DACHGSNzqPNazFR+jnBf
16vp+in4EPuvJho0fJH6srZmVkkmPwFYjJiEzi67ui0D2prCJmc1FDmFFm/g
bOh5JodYghh8Ijotnde0qEZBUHPEoXT6QJmTXF5UotbgoioMzqTO3OlZCNZe
O0K2CLv+yY8EIwh0/Q2UuZvqZy6yhZIwKqnr7H7FEpxDlKgQMm5HzpV3iuUf
TzPknpJA3dgMMzxAjlWI+lJ4+2NrkH7m+Gt7yuOYXRtshTOGQkDohkkDroyq
M7N+RwsE5gA6IB8RjiwzqZz8Iv/SxmNwev6py6s3MxYT3KG4Kso1xIMRXdn7
+rPwiL3QrHhK5fTY3hD+CNFP1YTCJUDUFJrJ7QPDlAbXHUOqOg7ZphGaVp3F
fRlwjp+K7cWyAtZlKSjDR6uQJTCceN0cJM6uUFQJ/xObeoBhtL7uI57ovnyS
xWvhe9UP/LE1HUXTZ7+1jyqoeinpXRnBKFQ74DxpHYliN9lejUn93KMwY5Ah
i6UNXLsru2qwZny6kBwWAZ+DOr3eRL1nb6C1LIDxeQDzWBj8/JhHyU4rQZRH
1sZVutgZuSVnHDW9yzJlpBUzm6qbbGg4Sag229i33qRiBuAbL+LmRDVJ5bTt
4M4f7MiESxH/fN5pwMZ7DEEFImmbdyt/8Is/w152VbgTMs63f8aK6iEVekoK
2X/LPSKhL1pAP8Wu5Jk12bhVt2QbJlY3afSYI+F9eAb67Hu+p4DJE5//bN0x
/5ynxDDsg/hEI0zwJZi8+K3a0Up2B+QalQRywvlzoFqe2gJ3zR/2FOeWkymW
75tsck7Tp2jqNgCpdLm/YupvohmkWqvTaPR/TC1n+bCDe47vrXGRlnII8eM3
rlrPZhZMVosyhhsgGbSS/OxLS1k48OpkDtX9+9ct9gZqM1HYMoUvjXVb+/Uc
jKHNoCowXRzVp7JwAdZoCuOg7twc9pfPGmvTDBNAjV/3fsKlIwICAq32Jwbd
Ve7Z3q6qsxTDpEzGInNzVQ6UsiA98ll1gmf1jRDCZn9PD/63PnJXX4ttXisS
abw7BepBasKRvO2WYQuU8zZ8zkYVd63IMJRGG+4Qq3RPr7onGs/RnrVEumIn
s4LuK2HnwaTrxiLf6NrWaKjVrcUEpFxBso/1lVNSr6ARhyuhHCTekseYazT4
tNnEwNMVBw0pTes0Dd15t0F5+ntHEDz+HgtSS3XG09u7uPOjirO+gu5K3aNd
5lspk3ZDGQNpseFAnZ3iAm9dlngbzhJFHrKQ0kok4V0d5A0/0GmoYxbj0abV
VYgsZjTUpqpA5whRSmMZ1OLGn/Zdu1fAXwCrrZEcjlcNFsdG1bzfpF9yOkdH
Z97o/7evc5FvOhpXBdZ3GZyWxGRZ8kWVfIis+CAu/P9ZTlC4pyD/5bXVWWRn
ikTRtqSJEFHDhMK5GIzu8czcDHrpdehsv4tbNYOkyVChZmNEd8YBVSH/zimy
Lg99wt1JFoWnhC5TLsi1Wt/xUm+BrKN0EWa6YRrwVwFdSrWMb6avH51C7xHY
wpCcla86rMs361tC+M1XI5plBOdC/fM8xLA9oCwd3CaROda0eB6/ATYzx0wq
r2pnz+E5qI6t+vSc1Q8BDR5Ze210WveGeSW8ry68zlhJqEQwxUCSU5+T/OO+
RrwQ03SDyR9aOBABuWCq0vXz7dsy4vQXbwvPquaMgnestzvxS0ZhH2dke089
1q5VsgybOTSC5lWmiBR/gzxXvsEcfc9A98Y8xL5652TC7Os1Vyn3X1/GLoxi
dvEF8Z+d6WRSHNvk8w/n13/EAhlZB45lSqoQdP9TibC0lFP0RE46J9Cq77Fv
L+1uAw8V7E4+4sL6rEo2bvONd2g+9zOEbZ+1H+t8bxxwZzZKZfOYBvdKsu61
4zMEeyNwAFut3NRatJ9rSQrzJRSwxNOdUZku96u7rpDWJ/nYyrQCdqvFHG5k
u/buvQB9e74oIfWurjJpydj5CSFT0+LJb83ttjxOaVfqrSK+kMC691L0Wj9j
HC06mqz8jXWlavfgCj4DQjDEWttPRm5KH6SPaeNGMa61fDSs5B8AsWwZyknT
8nYOADlAEP2oSD5gG7THYNRXr0xqDhOYBXtGPNOBlla9HBBMnQPuCoDh+3AY
vdUbQXiXbzrDSunmOHr+owtaIt8MwEzXQd/+oqHUe7oAS3kVoagZg2zMqwrS
mB2JaX25Y0AbablS8D2dAM5pb/LNV5w5HL0rOPmKNuXuq0ImZn7Z2Tq5EP0I
z1h1OQpWGR9WWXVixog/6t0g8YUSp6Kza8sYLDWrVLN4UQTHoVoCS6sXHRfl
v+/HKsrVm6v33s7i55sRnOg80D8zKbnONENVNKrtg0iMew84Bn1wj22N4DJQ
LE/3qFQv6zRoTk5qsu5ZrcqwKe6CmUnSRk2ehDkY/Ri6bvzhGzvMrA4ds2OH
kFW0MjP6hiUa+PFUYtVDRHmUhx9FTbmHhgfpEZv1VXRXKE75dQLvjFkZ4nis
+kEj6nMLeToHXi38AxL+S0Bg+DBXXzdiQibrJD1+bCkDW7HVrAPmBhyBSL2a
NnLozot+xABv8M0eR3zSBLyeYv8+2L7m5lGTbPEjc5SfwT1XT2KM2MEG/hky
h340PKBOx4UL2jIKeUxXfguFKrQT6h2mX9W1xL6lgfnMLjRN3iF+TnwnHoFZ
TuPkBEPVNENO5Cf0Sa8eHBTQ3BVhtKbliohDp9ZCSpl1KU4aPCHnJeLGp3Pi
ZYHVVp6UaxLDIjbp1/ZBTis+vH1Q9+UsIEVxAYUiR2MM3aOoxAZWhWX1Y4x5
yu1pC7hTXAVuZVb0wVCdL6tMv53WyLLarXA83NG/VynpGtjqORr/ViHjoXcO
8g6Moi97lQ14zxZynVeNrD48FTAzBMiAquVOxZ/7mCcYhun/yUAt3iV1vqgf
W3itsJhCDZg4RSq8TE/bkxoYN0+qYylxZtQHWEoApJ889FvMYqTTPNRzyaKy
H5DEOvwTd/VOTAT1AudU5boYo7Zeplo+h5OcPpgcPt+t9g+8R0yrPgftlVRk
IsKfwnn39zplQ69HtntAHCZFHoHhLlGyV8lgnn0u/1JbpdQN1rhrulAfGn6O
YHCxzXHqO7ww65PNEjk6pPpiGd1IA2qgSfNG0YYfCpo2gQFM8BhtrURcWN1/
NuyisXzr/t9RtoRw+C+LpU/bcbZKOEWKzJsTEJ3GygQtsXoShFEd4w6Y+KFd
z9Xx6Hac9cF9NAhb5sX3E7G498fQLVK0QaoFRiakRxLznhFlgYJt7kRC22Ox
aUJXs+2HcpsD8/h+upydzclFQmfobVOLcVWJOOfX9cgBQfpvnBkFEB3p4/yE
bse5ImEDtsYRLPnplqa7v9vPLhtb2oncHoT8t4pc35IfsuZDQFI9k4g1tk4T
axtS4plcD0qNB5nx/sn0t93onaIjR5b858dN6l7TJ/hrftYGQBAWMMyKjy9W
fDaQBd96qj4yetfrY383Ji7zVJe+T6wD5pTFZwkhO1gs3Y5S9K7QD4+BF4Bg
zjN02teL8ecGK+YeEITssuacx7N1YyoMYBDseFUH7V6aLTrwg14H9YEGZc4F
E4CypVqR8wLI5hZZNZ2p172KyluxL8yPObDdLLUJaG4BAn7jlZKLP0b5qZ6K
yh+v3WFXLPoE4jEi7QnGaKh1XRRetbBs6HxFKWOOJwI3LS7Q/yALWzNsqaHL
lKx21sqaJZR0QbmuV5e7BI86cdhlaIDWpqPGQtPtujHVp3djybWr46BJP2Dh
N8+MSv/mnv47Z5JN7uL04vGDZHfz00jMZSngyG6Y7ARxJjBN5FVFVscchvF3
4gFs+Mx4enMDwFfYR5fcErhRjaVVFNMuETVUmqzGXNI4oFduUwv9/iXE2n4F
ygGdjkt9tcCd6WH2F1B2MPCTX54MSUqTYuGEm3a5x/H9cv2HkdXfO74X/qPC
pGMBRkTslIuDUBcpuGEjGsxkH739dLe3FvrzSGiP9iPo50l5PnfOI8A2Q5YT
oRPo3zjHcXiawV/31nqvdOnA+/MkenizOsBx8fx5WfN1BAybi1pTz0FMGTlY
cWz+wUhJHsWJyhqWodXNwH7qsv7h9j+JNjhyhZvdLEvF0yjz3SYxzopE6cBj
F2yjn2f8W6aP5x+aqVVmDaq1GdupKGHmD52OhVdA1P5d86QYF9V2UJ8rvYnh
U9ziXSzovAZzISPzoXebS1lIFAvVGQm86vIYPC5YsxV21szUsLAJAhw9RUzZ
njbFtxPAktyjOR+Yyi+v+6rf1DpmZnQDRWx4jwJtsenT1Xhhxiq9ry1EMt53
kqQewi5vmuLBSZu/SiO3YVcSmQJdciTaBr/ak72hXkumahf/Vd/EHt74LPx+
UwNbfOW4SwjajTe5KAekkzTynpKBopSXvly/GYEZIsBsM7dRB7oU3Ga1J5KK
3Ri0HmCsJRGbYTQHfvJS4x85JuwxurYTgeOIqcUZGjPCS1SOqunq27yQyCdl
WBKBy82EXLzMVdneCqGi/Gp6NSu3CzXXLjzKl8ZBdbiDtNXlxKB78iWGeKLK
3X+FzBLi5ysnJOMvr3H1tcbRbz2IRff/QBBirb9lGAykc2tZexBUD6Uapgk3
LYJnAswKSohBxXNNBs5EuokUF0ysjGY3XzHesTPV497QdWKMD12THgT6hW2c
KdxuGq10ZWq63CrlyvzxFkQB0ZSVaKyQ+tzp6GJ6drSGQgtPjP2E16rXUhE2
kUbp6pTkMT9DnPVbNl1RufDmaM8xPIonCFNhsqxiAew0qxjzPP65B+q9AkQZ
tv32fXxuhqvbiLL2xkSW/Zr58RCoqoG4tHYp+P0btrYqorOHMoUxB/WvFkl4
8z6shyZ4VBRG0BLYRCXkSz1JSPC6ZZNtNW/kCVfpZUaIeOJAndRNvJ24V80W
TmVr/Pxi9vAB0rmNYD+Vxmqw3zOTatATnJkvKrR2bcZptQAIKGlCq2BJCEb5
+R6bbNEwjJKhBb3skvb8kSG97QYRQiKELKTLx0h2+sDX8MnpgudpjkwgDkns
AMLoPDjlHS4v0naCO+yj21HwSjW2bCEJoqd8CK6XgVBs3sX3q0+e6oRl4pCC
vp9BlvX2pqlvmu0yM/Q4NqLWQtewnyg5ca43uoeoP32a2UK0KXOHskaNda4E
HJ0FjEJG5VRmV2sbNA2hMFM7c8ldxPCBunonwrAD40wJXLu0GL7K+FAZSZsS
PoTd65oHdLxsNWORUbMWvDpjwperPXZGnjlyP88y3iOEl8OCjJO2CyAZ4yBz
lv4TVssKIx2nvCGX5OFDghUe8PBNC+IJjmPr/1QG3SnfqdQHJagXs0YuCxoA
c7Ui2n+xGzLihqqoXprCsFjH/4btRcResc2C6HglFhijRcTEKO3QafJTiJzr
awZsRM39WNnDMvNXMKT4Ytdg1EBbljle9MLxsbtmK4IbblIrWOaYtNTIFq/s
eHPiCK8imMfEAk5y0jV91khrJzKi+fhse5bZ+YWlHC11aMEJ4jGm9PFfxRob
TmCrymdPthSLSrnJEa6/kdUMh2gRCR4u0zFRPr3n2/0/k0M4DuBbmYM7WsJT
oQA4GCL2wGQbdZqJwtAHSV5v8T/ZpweFSP+Jd0z/GBJyq6jEd3jQNtF1fSrf
GygBS6JVDXJNRAB/c3srbbCZBSGVhrghH2Z4K4jA8TzX6tpjgZuLod8dXdLi
nrYmbEujOa3oCWOAuTsh+9Y9yUEd4tSaKr6bC/5diAru7ZodS7JJ97CO7nqr
66UGRZ9KMMPofLoj+TBI7ZUvA6gOHhXVbjj/QViyVKifor+mpqIeeoq8x2ir
cxwInNQjuL2ZYYe+0APiyLQGELOQhUSAgBurS/vxeRR8bqWEJF7qyohzF2jA
1JZGHlUJYuMcXG4xNZZ4ylaMIW7Fg8w0eDS/IVT4FPxC9u07WjenXd4ikpNg
EezLzd0w5PN556tRQb9Mw79D3AOwbo9ZkjVfixETQxUkcT4LPQr9SW6PvvPQ
M5+jGxAESqamu8fHtGJuAM94goNy540y7gBOF5mVtEq0NCy4D28zCiY7iH1Q
OpiCKUC/XySGqAVy/3CrNLFyV46iO8hI37TGlSG2ZliY44FoNiSKhkuMqkWp
an28mv3lK+h/PqWjcKQ9udWMKamr6EYsXnWL//2avhEnQFWTbPwC+lxjJAIz
FmlrIPMGONoJvlsolqb7SGMngrseWgGM1xxY6qoBzbQlbfBDWHHpnT5oOu9Q
+KINnkeyjAZFDgNU6RMvB2PRyiRKudk/gvtHas2rkF0IEunmTEYRLYpiIH6M
9DISqEMMIymJpoOpF5a3qivFMI6wSq3OvDKSE7HnhJTLvKFn3CMZSzu2LA7V
pvz/aawTg08HL7o3Ae4M1q0xiBe22Lus1N7J84mLuQtfIUo6tJUB9lDybnld
pdGDfdORNFXP6A08NR5nwwKhR8AhZRZOVDtfk1GuZvjdAI1GLFC03Enrw7K8
Fep6KkeMcvQxx2yeLVPg+Lr29NlQmyvC25uKVmNZmx0iTygiNGQf02sb6d1M
7iHpKtgTfUECUKZ6Dvnor13BU/TNvgsk2f4I6UmbXUQFzVmP+BGRhp7FRhwB
aLtcXVqItEUH2MCWRGhBRtcaZiQKS8rxr178fOqh3obQkmry5oPx7i6MdGZj
ZmP05AVwsJR5TPFRjsm2igkuE09ZxXftJ4Zais1EXBT407quI+IsDjQem94A
Eqi31CQ6Qezljbhl7ogI/vuFUueYO48meg6sclj01JvEHBWM8xsBWogfCqQ3
0gR1UfB4ey8q9AfGX3dMCzgCl1gDomDdhKj96mrnlk4SwlSo2i1jR8t5KFk+
e9eTJIOKcb643TIUI9ofzmqJ18TZRtP3Eme/xVKrU2DB2+vUzC1cTkqnQUUk
lkapxYpPIX9SL85mLI4FnRv5Jald4XrqjVmty9zdJmhZTKK6VUSUBtzhUBmG
yWRDCRYTzIOnF9C+M8F0puCfI3LM5OyWE82mFYOWxxNsVs6CmQLeU3DU9pNg
FWrRz8GZ1jIKyZAM5xR7+wLxkTbuKQAeqxshJ5+6Ti2PFPPJIIk0ds32+YmS
H85xSZYd68EpjD9MSK3mHlxCmGI3dvnuPY7UCZRG8Hvtvw4vs5Ik9Jq7kNyW
jZUFMq1IqU7sT2WsfzkuCOF70s7mW3r1jflDY+HhbR59+fVVGaMTL2dUqj7E
ErVcQR0ZcSnZq/EIDt81Yp0XNyPldp2FfLEW9N8lWHXgjXACqpwxhdR6/+Hz
bIBJX+AYzP/6LKaKy4kWVspYilNL38zqsjAcLhXjejLrfMalN3Su3Oyp4vMK
75oRgZhmYBQUlFPLdQ9BbVSSo7BH3DA039geEWRkbgF7q8wnIUV4i7H1C1LV
ublwpxjvv1yq2cbZlET3wTkerbgM9hAbUFWzhGFFiFwF1juEZgfpyzfrOZKV
ixaEC0g6X+gLpXPJO8yWjeeEz1wPd2Trnz1TqwKUzvTPJKDBKQxCAuriTERB
nUW7jxQlMwY7r6C2fG2BFB2Hpd6Dhoy2YT8WgnILLOZAy26CBqX7jr4tvkRH
b2rWbMME3Cg7RLjPB/z+kHP2UOGd1yhDetbgyhxQ1LBjPU0CQGGJ90QgRfOa
542ut8YDtsMJDAUNwLJJ+WQF7yYYidTPwEDDyuUx0uz2bX/scJNBvWhoWhG/
7SeBOg2y7V/cytaZQjgIYpFMHWmuBx8iHxUoqU9Holc9m+H9vuxtoUcAk1es
+D4ufULzxDMp2R+HCaCE8Z0q6DMBzQ+CNRpp3fAkwCg58yzOWOy06iZa37yP
v/OJ10+Fuj7Rh3tZvPumhTfESQsssfaHJpxEiBMqOeZzAvNqb0fvjtE9gmko
NKHpFq5JrDHMEVHvUUeemWb8OTeo5QFnSfRDFMfMGFVQ+54/ejLcVjl5Fsu5
k9FeZZV3qyuFUHOwUCaIUom08Y4P4XEHBPyPJoMBCrmES+s1jrh+RDHWQwe9
oAYWvMXqwjgLaozYMtiv5oryl+Km/bPM31hIUCPA8hGnN65XtPeY5jU0FGgV
FBH4bNMtIrL8cYyRBWEDUwQO3ZskeQBqW8xwF6BsEJ32Nu16p6b+uoCtQt0p
K78NeheNT3m5NKl/LWWqNeOOHeS/c59SEprD6PV9AfRqlt20ismwQ5KjXydB
ku5i+JujR7MSVhEKeg4CS3DLj7FkWrcEp3rLG2xqxo0vYNkNmJwI4JujfnqP
L5qKr3Ce4IgwvIVi/6+0gbsZwOAcW3MYTNmvFnsBrBei8fACzpzYAhFAsTQH
rIJc/D+Co602ABA5aRKKeUR3yHkIaYbnYP/6OG1xDPSJOFhCMU4waSJc0beR
8FnVqW26LwFWgj8+pRFUOauxxmKfzxFwCymv4awCB3BIDRWenQUzNh/IfKH/
iRCWKgSjygQlQmxRrtSkmFbqWIAPIN+0r/5rz/TRB3ry3ZlesbcmHkRqFpk2
NnhIZo/Occy5fB2D9BzhEdVePAxSoELEGIal6yioLfUdCsNcDjCO1BRiyog6
Z7uDeiwrUwV4LXRwVqH1v1GtrbJlcoMnsKKvEG7XAMJTW8i5+wuJX8EvYgv1
IRb6ffgH+lAYl0hqYl2WXQI6npOp30j6pXuowHLlzNu6qku05i26GStQuVGa
guRoOsuug5jLl131CgmVNCu70fNEm6ZR8smMp5wkWzTSMElUBjiZRqp4gbNq
hLlu5ZbvIB78AZo7xp/Feu1fzBNNNfMsCn5hiqiZGsv/+a46viFpOMGByY6i
niz162eFHqLAPmClZRuUhFFPLz5TGgo+LPlS/KpQBPQVgdL0G1jAmJ2o8sUX
zlGjh+qRaxWp8yVgQTKS44qTnXJebox0U7UwTtfc+1HBiWgL5OMF0tza5Zob
ms0+xZGdppZroXMDcZ3SENjJIsWHH/QMwcHvRKLO8qkZxbINaxwvfSu1WgYe
G3Sbvbh6n6DfHK8Xeaa+LKTUrdxRXtt+0q9b5Iy5nhExs7lVT6Zkefb3pfr+
9z0jNKB9Tbyicm7WYUvkHkhUwQlJv6nYVrAus10R1IQHuKe2PRF47bGv2Kjk
46Z4pBuO2LmziXctf5eWdMH7VeqjVUsHq89TuNjU+mP2/7EWHlLKNOkpHUYW
jcV5NC93VrXdQIpWcYuh6xZmhXcnsfZO0mG6R65NgbITDQDLchG4hICs5ACl
//6QczE62BapXzh1nQ3fs5DWZ4RJHy1C+JHN/O3h56qHubHj/woTjbDKQ0Lg
d2QuYZivnR0+Wu2Y5+V5yPY0wLEoM5ZDRmmvSUKXJQLnckcjuIOb0jpHCvCZ
AwE8D++5OvoMdn1MjiQjej8QAs+sAh166nRUyteK4Jy2kLZKlH9khMpX9X5F
h4tlkPlB5NYZaQRIQg3avq/q0Zep9JBVAcIRaPF7JAzzfrEhmIMS0YCmjKZ+
5zCY5sLk2F4DpzDTCdAT+Q9wgCDM+VuQeTjEiXfvn85Mq3jfeZSLgig5lZM5
NnRWjUE8HM/AnL96fU1XPy2ePn9oT4qFWFu7IJJCv19Dw9qtbScmW4dtFA8C
hugW+rLfZIS3dCHIsFh8ZKYCW7s2nOFdYHVPVlhG/cLUsAXkmRAjm7iWF7k9
B05Y1aNTmo2ruKJbL+MjnY3bYxa/hcfFoTY+0q4PWTphdkQH6PhGIHQZ7sgO
mzPDAbF3nPLqRBgfRRjtUvVLggecgh9oUElRk1hIFFCwdjLcLGgqSG7akFvs
jt2gjwIWqK/6e48/dTJaDHNLIzyNg5//4yCFRQYDqfMwRkVX7TiR5zBDnQd1
JFpHXp68DeNIw9AdUXbEBnsy2sLfomQ/Q2TzDLVlyd+s/tOKdDH9upg+eDTb
JU6EqUwykIYkYnN9YyRa+yuvy6KEJfOT0/JydXEHk8ug426sAIrnKq1ewDFR
TSMrOmKw76dv2FkqJpW71mh+ZuIyW5l0KaC+OQCqHnPA2xGgwdU4+/cnbrjY
WxdPUHbzGKNvFgLJeYrxagrJRJZ/2yYcdVYvXnSwv5WiJv/xEcm4ireSOCyh
N4iWKVe9oa1KXO/4cTBt9YY/cC6fNt3tbI2wk8VpqM6VW8Ysjj0psfy01OG9
Qoksh9q7lp/rPqhvP9EQ/Au5tRtMzrFiqJLlxnK1bJrsiVfYElcM35dKKd92
4s4J+91B8yosLwaONhDljNOZ+PrTu7JhPf/mj0LGOaLIK/YHr9I/GW3NxHIK
AL4CSgmRhMGLocpkpheWoev5ft0ewQv4TIcPhNiKSE3NLtHMUv/MLJwuB2g0
w7ogXfKi3q6RZg63JeuHpbY/vt46KHlLPHRQdtKYt5KHu+2SmuhR4YwOAdqZ
KGuHLwel1hpBr41R+p4XbdlY31mRQEDAANEo/HoIp72iUffXs6ZOBp9cn2lc
yDRzja9cV3PeyjsihBn1FU7jWXpFu6WN1aEXa05yT+3v/pjQEpTntBdovKJk
DWgQuSzIzcpqo8zh/UM3YEBhg0CvsegkaL98jrxjB6Rc4D0IvRnFDxK1ax0I
woAsAYH599vaAhEQZFEfRUQfYVqIwDM3LW1AYEvpk98EVCKDp7z3yJ0hqP3s
Wh+7VIy9ZP7i7lDC4vCETNQijQe36len2zI+qRoEg96W+f19w+pyldKJN7Bh
5RwxwuUWfEtnZzv5wBR9dGla16ji2t7sOi/b+YFTG1taCeas/5hip7JBmc5y
qQ7K5BOg/PRyJAFXOmy/sGJoBOePQffPSw6fay0odgmq90LQviItdU7zSE5B
KHdysHgDSEHH93k1OY2IBtAcv02C+ccqH7Se5C65aEscQKhHX2uLxq6U1Tjc
ruzcREswUHKabRKZMMS2tnB6Rc3ANWi6FQlE9/nnf9ZlXdQ1TTaiW/0u2pJo
DaMNJ3nAUYdtzXiLLw7QUdNqVBtBLLTT2O8kPFV3e3DSUwwwtKmIJL2cdkb2
uuxjdwQV6emGAr75Cz8Ud2nN3gUvIrNhTmE/DII74m4uctyzjceuSUTGG6cj
/aWIWzb65VibjwoyIzxm/CdqV6PbftytNxs5YJMMTTs3++ybDrNjTEJz1duZ
BRBAeK7qXk3UJ/l9F2m/qE5um8b8EJyYLZycvJvjSP2T1Gyy91OuIKbYUOFU
ydm04Sw6rPpiqTWdzWVCFPFXOmnd0ddWVBuyULRDMyJ2CHv+9lHHmIJlMfs3
+G7igmLUH0wWikfUQOu4nR6XJwzNNeL2BO03cACTxgPK0XmnUSw4igO9Wh7Y
VBu2B5JmVcdDXnROgv5t1PFdD/R/ysg54vRIDbUrc6grRWuG12tG5i2eqRrb
ThqKlHovjHz2M5VA+M86UgVZsRWZRxK5tVz3Jj0FZ6qS2e2nxVFlp5EaoFE1
oTnqGBOv9elyaJbeTFunoGixurZ0Nk/TAGME2hHeb3YM3XLrQbGw6H2gsBey
O1+pPzutFf6pdHrIkTK0kHC2oJijdDqFa5yFG1oocuRDUMArDguUx0iV6p9t
oKgeW6WEUzWXMYh3YZIJmC1iZ/Jj+Wjbg/Qb0IrCpk24vS2SZp7nK5HmmOiN
01Mv/L4rhz2815bKP3wkNA/C+7oal7u3sYjlbXH+FMMfRObpMvXAR6FulHNw
yYEVfP93RDEspuhQC72FZzXG7TXcL1hfLUMLQP0XEeqMIh1T/Uv0JT07gN3o
Ew4CVJ7Rl810kbrugLOZj/eMti/S28v0MY3mYWtfvuBPYo2ITZO5URqzyCIk
Z0tuAkv0WiDfvApAhAhfmckLPOjIvhZoQREnbEiUYrwUp2GEJZfRk0KBoXV7
++00RRGmc8+slIqMelvT4LSNsGjCAiWpyfI7uu1i9xUy9W34G+g8gm5dbDiR
U2qfxu82Mv9+pKAmwfLZWW9WoLqdF9bXb85R+FIgBAggB4tdLxQg1ZaYW516
fUpbn/2JuR4z/UNltcc451GyDUb3QRkQAXSlI0USI4SxBmBMaqfcxi/TfbNT
4zyO+Y4VLINmEtxnGkLfYx0hiyFa5GPszEWERIMagZ8QYYlCr2ONAEgEsVDA
tCycCrt3pCNSwQxZcI6hLujImpmp8bOFux62Lq59s4+NtK2getSQbgbH6WGR
oVNT242O2M1T1ABjVioCQt7NoE3eJXjO/a/wYsLCd0FWMHLQ5GKd9Fuq+MP2
IfBobvV/eNpD+Z6GsAw4UAJ5olql9Q6pKGP43OgOcw7YNBIMMZ0sKqHzpnvn
Su0SwYjxsMEzCzTfqX0UVYv9mcR1wULeDdHSSEqP/94RrCWb5L9x+bd0kUH/
mV1jM53gXlyXPqj3p9nKK2EB1EWZE3yUFwaQTnKi12bIHCuSwPbWngQ4ulgd
l7VZiFbXKxVRP+RV1rue6Ns4KaSsMrQNI5p5VFWDfVxSV010ibx7eoPJ6kgu
DXt2OcDdcnsl2OMa2RTDYH7A/ZjF6e7vFFNPuYo2nGIsDPPvsC8K5fGyCssg
Q1WgUike57ZT4vhTpC8Y2tBY/LtKVB3WD1JUBq/DkbYkUfNegRZ/KLdWlEz8
IYOFLkrJsrZFgoa3VaOAEDAt0LIL5ytZScf2nW3DZBPe3RfeiRZWl/6/7raO
SKxmBS87Ju/Jh4eINszwT2vJPzJI5ws8DzCcQU+w2dj1WPpVWdQpSZHwPrsW
fAmpGk9skjdJSi4tDIRKClm3oUwXA/vpJ6V2gF3tn4KQYvw5srkjYFeWtW4M
uk0pofG8fUGvq6brefAF9gmy9dl5/RE8dAv4Ft051tkGboOcR9kG9K2onBcn
zLWhlpyXsF+Y+69uOWuwof/jGcGOig4eY6VXzRBEQY47EjLdJpMDEmHfM+JG
76MLIkNXpamOoyWeKz5iQ0Qa2nAlta2aeQaRvwDcYVC2AQnSaRBzfnqNWOwf
5c9w2zW9cIaM4xsJPQ8YMxMoDR2yRM66uwYc1nAbm/+nB66F3J7UX0rEKtha
JJa2Ujc7vxnP++3Yt4I/uX74k9cDlsksjKJgxkhjwBZMKkRpCuMz5gwUOElU
K2dox7gL2MiQTXNIf0SeQk6x+vr8caZyGpliRa7/bV3728uAjG+R0nRt7st4
hg0dXaifj8E5Q9cqeZo15WLCWoMrLtq3BCSfO7OLdANuYP+gyFarQMs1oKBp
GsvgJg5l7W57HKWd665Z7XTbUg7cUgdTwTFaSmUi+Vi542sF51va5ZVi0Gy5
w/BQta4YkFoBad67XWzMfMy7vq8REujnbkBDTkB+2UE6vhbKkWlPEyoYxw5l
r0lHbqJTc+xxvVvkK+E6dmg/RkfYIll5+onj3dIlbW2uQkpeJeQlzsdccxKk
O+ezTMmO0r4OI9G4hL6z8Cnwytn7RAKhQ8yEhgBYw4U7LbwbrM0qqqVmAqML
pVyV11ME8P984A+eWP2dzaMRoO+vslHV4F+onYYn13cDGPBjZfX6CLfVoY1d
2XExlfPBAje6AxNKhodIoq4flXdj2xIxkdjTxfL764zmBFFVX34rGsQBarGk
XsOyEYfOMIjy5b7K6ygRi/81u0m9bJ91vOLn6bDjeZjAN+r/mifnx/4B/bEC
3Ac+SbDoxYOYep2x7aNDjH4g6I5D7XD+TD9y3kXIbFhkCPChT8EhH6u5UJhD
AHdzlfK/GLWHmkAZp9CMOxe8s2B2O2L8HyuG4GRBe9Diik00LyKGN5vBzPLx
BWvTOidrjYmD6Qpgehd/GcxeBgWidgpYwqe5ocPYCDD4c7WVI0YrUcTlsm58
rFcwMQU3CFXS8SqeSiEVaRmHsqS8Z5EGw5Lu1w1M/Bk6mNKI8P3k5saJGwlK
dGLDQ+dmA7coy7wjZ1cnGU6hQ7ziwPEPZAbi0lskP7sg1F3jegbqbVXOyrVw
ZxonJxovLk41umyh62UusWCwbvDgWU0Jx9phNOum3hH1TxwtTVTP5KYKTpPJ
oe/1d+ST1kmogUdXCOkWN3gGktHBw1jytwZDvUOzdvU2TILAyUxT1s9lk//h
u1GQXUXiKHvLPc2c9TwmKxYe1BHitp8ycAa46QMahpaUNeGrHhxSOAd+EFBL
UEOXhJ9Ez/6NYtSlZa7RfypzRcGv36fWTr7fjXiUei14F3PTs7LYhi/wDzv3
2SRhDKA9IB5kb1oUJeLZzdd949DI8dkuKl6XwFqwpgNMlKDCKzmK7PcOMVIn
QV7jlQp2PFIhP7XEqaWEsZKaTGTR1HiH8PWscSpQDxyP9FdSjYvQEZZmoJji
YG9cjgYlzPh876UuReqy5yQiaucIY5RmQ3waQ4F5OePL8kVzuPlwIQ5U1lQ2
gz66cMkC/RK4C2XFXuPi0AhZ1wVkTklDxYTMBlIQeReceRyZNeP9TuX16udq
0qGdSa6F/+5qkzJS5d3cm4iuuVtC+w4VmuxSukIDbaZmSiGkxwSS4h9phOUo
fsiDpj17Dm3jLNnBtC9izki1a/szrWdc6csllcDdheFUI397vvGnXr+F7knf
FOyrvc3V4uFA8nJfrtD8+2peNhOamjjoEF8Nv3+eife85CXOVmg8wEZSeedX
UAhT/equjLUGJLF9eY9lat0GowAP7cJI3wxuTjFjezP1bKe0Ea7S4BuE6c5x
3CO3WOkf+XEv2RBs0VJ7H1cwQ6OlMa3ez3OA/MdyPrApvDw9yqdQF4vs1nvZ
l5Q6Omv4dCh1eV+pmot7o4i5tvUPn5Hx6bfStgNC6nhHpZYYrhnCzOzbN/JK
zdU+DdCsFADGR1LfTzBIFOhJOL9wIdEl/9k28ka3eyN3C6OzWQ9Rupfcgf9M
S3K8AXhJQRFuFNNYF5ClSuWY13bJB8d0kYVZjwotx3CaAUjxN5/43Cf0MjY5
5/NfW8t9Ihinb4NhMkpe8AJQ+gVSU/wVn4HHfdO4HDEeFpPBuzyhPsjX+1Q2
LZ2uPVwkB6nCJhGdOXv/85pGHufs2mLIDl/O1nrRD1kepeFn2lSdf5BEZ+U9
4Hu9HYIpOZ9hvx8ydGwZb4F/4Lw4uDAnudL4StvUSximiRI30IafN2+j32fX
E3PSEW1xCl1jUXj2a3Z790FB8PK6L0aG3Aapx0Ovp7N5kS0CSmvnQq1qsuwy
SNMnCWUc4NEhmRmfk1nsrC3Kckn+/KYnB26ggDCZTDwhKrz9XvPFbzJbqxn8
Tg6sHxNT9+mU09n82/lqELWON31Mlu6A55G8xXs5phsDRgaBgmI7wtv1DOBB
w7/BjdPtLww4pOsEm8uEyF7oVn8ChM70yTPsG2/1IKXtps1Ym5egeMT7u0zJ
92fZ5nvLp+aG9qDCZSfgfYUR+GQg+m7f1bzOFjj8VzTn2BgQb7tJL3eTW+oY
CP9t6IAXL8Gcam75d+J0gHEY+w37BSgJPnpSB4iJaRYVn199dOr/FKkSfg4z
Sr0XLSsJXxkUTdgoUn0NNrkVc5I4uqd+gml4355NLBiZJyaVwfkxfR1Z26sI
vNIuDzMFw5wbNElFTIKq/nAh0oPotalaN4vY3iBTnBHU0P66wSgQ63skZBHe
uP3yo5C+2Ar+qEWFeRfyVcWj6Ef8OOsFBsF6n2MVzSUFknK0T0RiU1U/Lyif
dkWg9I7MxBhv5KOWQfDSHH/BgHAHytCMPVVN2FJp/7/blgBmgPu+ZqQAjGgT
2O0ICSGvOEKlbz7gMFfMaw4xYJBv94EbuE7t/wofsnd5K/RBjjX6HGl4xYjL
ImBw0bnJtbwA+JRIgNe421KrozplVTOpqUD6FRSknNCaFjmaCmzTxRFdag48
sz4G+zInkguCALc3agZ1udPe8UN6nAAFBxgTqUZQ8cfn0FjfGckXTTSx+ElT
0ftqy2T8zUL1vovsJUjL1q6/7g/EK5NF83UJqRXBKAC0tQelKQwocMtFU3fV
QEAifNgazBTxC5ybHwPShdzGpNjACizuaRoTtH42WbRsYh/2ZOiHWa2Qhza0
uNLQvBHrNcjsQ3Vf9/y8iyeflE7eY+DXzfrnOflCOBeXDr8ayJlgg4SuD2Tc
72Y7lvb8o4oHNRpkMPTkd9DMANmUZ38qGuMI8OVJI+XlDg9QLaX+vJOxGUO+
kfOSeEsRaksDPy3VMWyMKN1puS3z7Gp58RQVh5PtPio3NYiU7Qdec40SXOeq
DKRzfdGA9Qcew04qsD/fsYHrximBM8S7y+RY2cW4/8Uq4Ana3xWtHcdDAW4V
GKEhWBwv7dxYjb9TPe/beZrnWQwMtkWl+k19iILfjrCgjpp0y1htSPnphsa9
I2pzXUK2iftumyxxPe4Os1ixjQFJNkt5HHtX+gv/BwX1BuJtTkbitT7Cs2/l
7Gp+Ibhui50y9l1Z7c3tkYrZw4I0PuKpvSCsMgPrJIXuXu3ugWv9WeRVBtnn
yXKC2RdltS0or4BERS1UEqaNLmcsKWraeUwad5tygV6HqUR3XGb2r1rQVsLw
rynG9/OyPol4KOedzjq+6njL4YVeVaSvUwrysPK11QAMg41Q1HymZOMpwsEH
VeHLjfqp+qhudrokUhECL5d97UcyAU/RG8ycNT5BgTB46xxgir3T7f2rZWo1
cVdx0PfXT/U3Nkh+8CSCmCi9iLV5VTu82NTf0n3pDAdcyBNZKoiMj8LcrvFx
gMIRxCUJ1+6Bp/bBgGNHtGEhOk/+I5Kws1B0P1fLjcQzn1SZb88mnddAWQAM
RIISmKpET60R1rVU873IoxWTt1ZMkuyVgn0m9W7XzrALAijiRvauJ1wg2hGy
3bT+Jvwyrty41lcBiZPIb0DKmqlWE0EUybszOd8wFOm/OL3FbFwl1ds+VXiC
7RNlqon3K0icKutElExIXjn4q1LCsCMSCS8kxyhCchoeALuzUT60w+5a9uiT
IYMl5NDAyxpXUExM8ZTVDTed9oQwxrexvZvot9fpVqKjrg0qFnDnjCTGsyF3
N/c4PqLbG3MUX6j5eLxaOH/0MM/Qe5I1xCVk/yB1w4TR0mMNShTynn2TKXV6
f9aG8+PUs9GEkT7I4/4R6uu4DkbFjq4gk8jMC9rTpauYnruWkrh6IhcskEcp
BhS3ceOlK4h1J2Ic44cDwDrzEkfWAXHD/CTAHlby3mom6PULksbjcatYnicV
JGncvQJKDHVCELb4idASGekyZn6iEHwIAjKPsNPwZzjZD0Axw10Mj+8d2qft
reHnd32WDvavBs62zlh7u23+lYI5qkYIYeJ2T46sYTf8rN7soQj3BSx6lSSN
NrpTaDGof/lxfgcr7Vrv19OSQjiFSVsLXE+pLbm6BAhNnkvMn9+fo7GyBRqX
hmeiNiMef32LfKqSHFPxgI6j/1GyehMXGm1Nr0sZpZsUZNDbvdccDFAH3ENb
P6HW2UOL0x9Zz/iPIbk5W0mRzg4xhtElxN+xQnJqNy4UiSV0IwF0x74Fvzql
tjlQpUH5o/ADjIwV+OcClBJgyqoN7r4McMjrDyDIefclRnq75N+m/00cnbP3
oKSoPUDpscsxL+K8mgjkn+NCJN0E6i+0vUCTIIe7ba2QK9hkImrPQhK9RhdY
z1FDLyLHNZarZOVQ0cqhthxJJC8CpCA51CavGbEXnnsokdbCdT4P0dIVy+uC
AsiE1lK5Tf+ggP1FeHZM8Mjna265iMs6HDWiRxsymYvHXbaD0tbwf7Vmyhnr
6fEAHcr+A7P640i5W8uDT9oCdMM+NrV2PXX1DKq7JEfumR8ElBtO+zZFh2jm
i7YyzcAN7wjNE5pguPx8ugU+HtD1wgkvCOecOzxRnZD0tI239mSLbOZK+9Zl
REKY4wRpgn/9IZFrfN0HsYdOFWTgRyRyf+3nQtJh00tZzBFCGW4bSO9hskEo
W0aJU3zF2YKhYnWh4QskCJh7kNLR3jiTnNRFnZAy1vxjsEQGdpfr4icLxMvV
XNmgIz4R/hoWPusoOz4AxH3hXH0GQAOC6YU7zBLTD6G1cOh0Q6R9MsJoW014
FBDpwQP/oA+3lXkK1sJfh0uyI6G3TrpRRfKQPL/HUITiFOoYT1nKgh6s1xnD
v9VkLoAbSqglthvYymA3n/xh6vWrNTjLgrMQ37kAfvGHTIShYiPSTKdjFrAk
8EOFOeQaQ9WEq/rO5p3fgyvG/YHZbBpLoI25cwLR2pMG903p79thhJrgql6p
W97Hmy6nXaa3/QwGGgjQcZqoiYvNVr9YgbIRnFQo/uuDHTRRqyV41kmv1GD+
pmG/H3KbxrbAvotkSNOA4qQtgQjSXLncmTbRoDuWSm0/tXkbNJtui4TrTul/
g6Jv/pA2gkC++sMLJiO8+ud9tBtCeNpcslI40SPdlKNUZdxxGBOUNQqDW8dB
uGh63afxvdp7exHkmonyTGO5g7zOlDgcDnjdspFEw4K2aLgjyZXG/s4TKFkY
nCE7lo2xGVH0rFHmX+5nHK//r9JSEaKSlZ0me4T1XstzCwnof3+SoMUdYY6W
Q0g9bI9TXWmIwDh8gwHc+nQBYMmk4IWUi7E7sh6nfxXMOJ5ptwWRrw9jIMqj
JdXC51m4BJGTyVFQ42p2rYC+ztXM7Lf+8XtXx+4hYWprKgrX53RXGUtVdBzI
zTyqUmyi3H9XDm4SN8AH58ud++meuNr6ow1WjXRopilMasiI8My+4b4KFOn7
DLxXtIt55LiQIZoDrrVdixa8nC3ivnh6BeIvijn1Rovv2YL0dFT3C1JLX73M
1Ce1ZzGJNgnv0m/+qrwjWGuoo6hDFiDTX+lvJoSrOCy9D+njmlM41U2HywUF
qHYFMVwCdUgopFmIrUkQH9saGMVcJQkMc6qyWGmdfeANElgdtq5OeRqnTw7E
ZF1DLx/35O1tMeL0cVsqOyXQiVi+iOi5Ck4W4mF1TVd0s71kzgLNNxpxd1Az
Blr5R9H72Ao+eAVwXD95gcOSmdTceLRPFqZWl/sb9GQJ5FzQ9B2X5F6nRaAU
yEEV0ItmENbXeDfgat1JjBBgc3YPK8nev/agnRaYRo2KL5RlwqoCTAb/znDp
K0ILdC7LQzZrsJMOLZDF3NhXwjuPoQLekBsjoL0WAfzkZZ462TVEFX8+76dO
FM/bJ3g54Z1xboAD4ULpDOe2PlVINaDGQlW5eC9Z5Z2h571OQrnZ/lD/7vwJ
cUrcRCUAYwnXNepZwxaZE8RiFfDGLHgpzzmpePhBj/q9sZAuoGhTjsnKb5cn
ZRYilR3OEhUMT9eQgRdkAOwK9pJzJe3B1OcSqSZnV1GdJDNDgBYgNFdGpWu3
/MTNJAPnC4qqBhHrQueXRll6OSqNn86tZhsMVm0nYTwP636ZPFTT9RSzICBp
ece6zLTv4E1jHmNlVI14Yug8lk/v5KVrrnV257jatfqMWE0hGI75nbl0GtUM
/B0YUxMbnWjnxTeiXz0HCbpmsJiYxk2dyH7psSaaPX1u0l8hqnCjOQZEMCUq
kQMBnApans+AiRbq/FbncETlcIOaeELeEU2aKKHTPxAsciwLKniRaUsbVDpQ
DXUzd4snlpk2Fukzun+AwqDAKVDpfh68OJ8Fdkv+r3LnTHX7kyhC0F2L7q6Z
CU0DM8u6U9etCJYlxeWgHpzV3Llz022pQGprIq3khzleNmcwvClELZGrGV8X
DsTt+eL+j718cQSnGtsFj5FwCJ8ahlRkQG/TPqC+qD+cUUyJuyuZZOQO8Fqc
jlfK35wVvupjticN43gIPLgb3THVbmhBVmxRbp4qwY9i4MlzaVdN9Xl8qnON
wnfTGJNRQZ/RwN35dCMCZnunPzWTa4ynil8wzaFIeHx3A44vNqVPecBVwu+d
6H6Ltrar60rem533oHYQhhBmSgTSBaNPTJc8HHELrfQ63h4BzOopm+t1YRdY
Ms4R+uuhTbGo3fnNsNeAKTdiyBzJ+mRPSAiPIHzQ5uTVpDHc2Ewd9KboNfTU
70x1S82c476pzMLftD6hh9RbPHNZS2pmfVQnJEbTjYhHtKc2/WISZ7rbLdE8
N4rwEEanQVbdSdfedIiY24KPEvjgiPgTchYKS19j2BYQO3kw6OGW+94MxEeA
Z2oYD+XmrmcqEuUct7n37a1bAGzF14apI8Dsn3d6zuCw/ebOqypKZsaeQfnl
KgdBRRi8sCBbh5uEkB5TAg4cUknNE3wvNWDNt9xdPOBBZkv1luOIUE9Kd0AL
uS1ARC4o1EoVZPKtL/uNmYWTU5mYbxk+Th0O21JAhnIQI5fEuMnUmRu80NkT
a8bSZAEN4fTXOorKnDRQZSCrxqBXr740QiKSi100tsIPEDY+hW8QhB2CxSGc
zzz2piiOZzKwqJQDsrSJLnvq+rz7SwwjxVI8DYVCrohAZoLPVwsKYiaWBKfv
s2Um9Jz2uTNcrJSytAJVrwWkuM8l75hbtlawF6u0fI1xwBs+8c6v7TaDSMoQ
IyDeFlX04gd4Z5rFkm6r4Aa2vMmj7GxiinwIlX7GZVfxwd/dFAFabgdtQfyQ
Bh4dLmwJrFpnXKpUUPCk6R4r314EAt9R+Si/aTTThM3wHpwUY1IN6fl/iBxE
1Mef3vuIHMxlBXClrPHVXd0aW9ki1ytY7BuvRjojiBHQYX9oR7kXkyJAV/I9
swgNgQHK4YDbc0iyizL4YoZgyihp3HcYDPcF1uYmjkVi4JEZWAphcoSuSwWC
gXcCjpTPo/eBukbXiob9P5UfnHopjsLa2DZ9CeeTz1i7eA3YDvv+reym+DD3
fZ/sow+8Yk9pzkpfbJMZPEWg28fqUfM4IbYqkGxRJKiygKEwF2rFDoSSrf0u
tOChucvd8XugwMak7wHbfq/paCbeZgmf7fs7ZzOAjaHow/14PzuKCUF9WtHC
Z95KMTwbhUX+DLeUMlorUprtFWDBc88dxx8/QLFjvRhjOhKrSZTX9PFzZAn3
jq3HTid3o2egpjLP/PlK8VAJ4pP4+ZtOnV4WvjT8plSOriRkc6n4X0HMtx6k
YD05MxSEujJWd2lZnhsgQk3uPaD2mn0pf7ydV4ciyFJrPbmsRcdyQy8pPHC8
UR/3PX6MaqW/g2DPilC+iVG6pM3I5ypw8eisj+EW0g+OiVtyUUIZ1qQbiWxu
NAU5FuyT6QOx90pT6J18qI2jAS0ij3oKq8TsOOfpmwYqfa4faQaFSZvja9l5
f4Xu+O2XDyh1QlF60iM2B64jcjcRUYNdOVyCcNckn8PAmY1ND7JSnpbInipE
QbeVO0KfzIFTcXaCOre2rshg+yaLUEzfY/BIghayBdu0gmh4SdvggxW9Bdww
Bq6BO1Ax/6tPrP5xKACEgY8kp1xnul8T6SsiX18IVfdHgl2Sr090YHxEK7gf
G/o8qfse6g3PTOZOw+//wCLuELvC7LCOdrzzBSShlz53+5wwtmuUY6dJ6nYW
aRCzimC0gp3l7xbtS2LP659/m3Tzr2OKyEwnNBLQlmTJ4iIzhPjgDkcJVAwi
T+vQY727NPqlGXB24TnFapMFGYMIlS0KjXHwr7zw8n9qWa5NP3EXh+x3svsB
k0XKxhbuUPWP7npkdrGJmCWpGWw+X6eE1PLMn/XRM6tKXJ04YFtNCh0Me8qv
tvktR3XDuUbS8Nwc699kdi/QNwYbtmb+vBC+eEi2PAIr2WNp6+7H50o2ZWKD
XZgSQUHZPPSHzDcwHrH+Vki46UkPe5O/incdWhc0Z71NGJdamO03WzEARxfp
Ng6Fh4pHYPrEMsicpYLWCiu99tAa9o1Ul4vHSI3rfKI+ysVmiHi5rGKO/au0
f0svKmLA3m/ZT88+O5Ihlgq1T92OxyGj/payr2DekGM7cY721HTXPGq6EC1C
FBT66RNqmGMxnf4H9BYJ0146vk7+UPGFCPt07wVf7rh92pJziHUyTgqggB16
n8CENFB7fdL+HmtVsF1TXSX2EvSPlKz+FaoVeucUUEhSgJFNXT875FaXq0uJ
0OS2qzZkmZMjoOdsMjusQ2JhbLT0vsZbd9gsUxZW6FkA1J7m9KkBocHooWgv
IJNQXZjtAqEV1hM2ZNDYliBmceaOpVPDJMdVQy8emLqdJkVq68mMRiC4v2Tc
YSl9WtknC4PFdLeYVkwvekSvzezEdFYYUfHl2gUuQ780G19wHUdoCeALV4nK
GSQ18kzH++d8oqqWSOWu4zxNMst95TnS4BSpsI39EI4C4/6cM9cc7pbJ2FCr
vgetBBh9W7aJUgSRO4xrmDSpVsxO11BtWZaRFEw9L/I/fpwQHYEr/LbOPNSw
6prV864SbNgHKhIM3//WM/xOro8W8J/dTCy6b7TFOA6BrbBEPm+n2DQYxfNE
7A4lCELs4wS0u44vU/S6YtByBLP1UmaiTdWN6t6iITw0KGlVvhHjd0khI71j
tfEU0NVZoV/EMR4iifvnWZUwWWYy/QywOXMs0qNfis6N2w8el0E+zT5AC89f
GUeX1zuL2cJG++PfaN0BcKjHR6o3eqL6jkrcl6liol3K+uFD6h159JcxjJeg
0vJ+AREbdq4jw/A/QrQntKpzw9XjXW3MvSJLke639rkHRz4FlxdNegmdYQ1i
r0X3CMdiAGyvZ9o3ssnvNYe0zSqYLYvwKZ18jQmfqEUs1v5bWs13WGaz8Htf
g3s/ajf3zbWdl4BtKSfc9Hu/GYxIcyxDiVbVmcUo2GDmfYvderQzQY2Go3gp
XbYp8Pj8ux8bGJicKfoacjc6DRoY1Y4MfFZi9gwGAAYgOWfw3vDzmc9cXfNA
pwOLZ2OvOiIghr3IYeI3xOBF7VY81odN5eC5RuNKx3imHc38oeTt3vGJbLKA
swkPM/xKpoMoKvZ2RpjG99MHmV4yn7aYC35YWBJAulN8AiLf4mP+debkWoNP
5QDIxuQN/pKIqMFfrCkotfM6NiZYLLeDpIb+Tb8CvBqatt/qtgEYPAUvqYXV
pMLSLf4BDvueGe616VPOEYiMi3it2FG5PVU/dqxSOWOXnFNXQXTto2mILA+u
ST1wcW4xuRWHmbluC7lhirt49Del9WyYjdubkky5wApMckVkFh3MctKZaYQk
4ySsfopoMYG0sb9ba9J7sHgTVqLV9MT/IE0rxjNxeNZTchDP4tLUmZsgPOOf
81OnRAlSg7TNMs0cuRBR+lDgK8o0vmgjkCeu2x4HH7hRY8eZ4hGqllylJ+Z2
5c4EkuY82oX0o+QBywMn9x+iY0n7/X+FLLuvKLg6xDz0s2u7to9QtnhIaDU/
eelKnekQvydrfFRPgwDku2l5WfaWheQAfnU3FQtuIW6BNVZ6sQzSlPWAe9Ac
UWyu9eX/3c5dm4UpQ89xp0pW5YxttyG6t+nvfka1qZFFZlxodopV0HTM/7xF
iUokEKWI8/fBeBehXtiUk79j3m2afC3mH0yxufDFKyHViAeNBeFFbsgLEMW5
khSo03+/EUJ22OSmVhD2Wf9shbasnOPDnmLffB7ucv8mPoAUAGs57xNabHnl
Fhn7I35In3t0kJn/OoAgTMhD0RdWvCH5zaSuRPP+ij6izgAtTQKVmT7QaEa8
+BBI9DWbbstGMi3FqTx/wfJXroiB12wePHzLbUriYZ7/ztGjWEykmDpOfvhk
FX8qMVXog3PzojbaUeD+NoamIOqvVgjUBU+tbdMMXy3Je6JL3/cwagvVnNHl
wTOGTv1PsCcySVp+a1bc6G4oeb4YYs9DYtvaDhU1ak1Ul0GmRFK+mTBmM1BV
eyzb+L8+oSGFewF9vt9ibaqNasr+iyv3asq01hBDVZ79/UTfp1okiM//AoHE
uJtHD3N1vPFfRzcoR4bSD2lrY7bu0+gTC+EYNPChtvWLTRzHYtpdtoo7oEbj
M4vkLlgLPbQMsdGds4gcpAZk0KI3HlkE9dEtMoSg6oi+R3dn0CvCuV+dkCJU
ZheUOkA12mDC8OUvSL1sYG4j+ZoqW0gRQXNENf5G/rAkkdSEQQLhzctnQC4y
YyQWDL8gZdA+hjcnKNh108MFmgwnnvwNgCVGP/q0uhB/0J2BnM+VW5WA2Q4j
rC/UV76pJBJ8bblpXLo4aNElG4PTP9G2CbzuCO0MlL/mR1+cfqTzu2Xh2Ukn
KRhkSSGhLo3jLgK5F4rr8hunRfw2T2iU6CHlNNTWE/RpPVw8MywVzZz21HqI
gdgTVF3fFEoOKa8nGDPVdDXVIpWxxQNlyIA5RXHvnaZpUi0z86mPq4OEqKH4
VE8l/OP/5PDrWv/5X4YgqE569vGW4LPkHA7RIbCNq8QAADDNQJklShrLzbzG
vDqyMCjT6POJG7vm5/I0GYFTuqD0n3mX6pKh1AgjzI6yNbIAn7Yxi/Yl2xU7
uelmCmSJFNumsyoK3pQLpxburdlaC4o2v2SJUvSQMOUhRF2QBRDB9yZVxKTX
kFyWqwFV6a7KRM1YKIsj/2VH4wyHgLeS14d229mzsBCCD6MFVL+3VLuIceYG
atoNV7wmccfrmzYAPRIYrF7iCElz7mLhpwI/VHUzpKlPI/uBvHB04cKgwL+i
Cto0zaAc1jhLlFc71IXFpr8VmkeO07nF0WRZAxVOOP8w5DYfJrEVqjg6ljRG
fLg+0wYIlP71StDqI2yeUsV6cpXi9lX2H9YKZqKhhyy0it0RbRh4w8ZGzY7u
QoZbMbPbkdDMMqRIBqJcdhk7AjDEgGtBhaebTXdrLI5FJCux2hkp+XHy26Pv
iDPK1jPaEIdCr99D/L2c31Fz+N6YCNMmC39KAwKsOsF+8qG1Rwqtd5Jf1Ey2
XnHyhNxj4Uo08hR/LWIQ1uAjGiWp8GdwoI4XeCPCK+N32smpDH96jnXqAw+7
OokV50QTYVifnlFB7V7jv/WMgQdRM4cQJ3fywaAzWxGwyKhBpwe6PuwTek+U
t7fTrdbHPzeatOcM36Jn+J5wHAob+BFHb8hwzfRE3s/fsHQ3P/2hyv2s/9Y+
SEyyLTxeXFNDjusJwmxVLZ9KvfXNSfDdpO7sp/fG0E8cm5meLRuANpC1Rkxu
KPRwiQk3SPGJXCU1d3osgDYlizJRdaC405YQ5dPMkXtMuRaJ25/bJZnPWRzP
VVT/Shft1X4q/tNi4m0GWi35Ew58WFhmxtO6qnexqkWRwQ3dPDBvaoYV0DUj
VEwrWxAhxChmHBpJnoeajAl6oayK4B5KjTdC9aLy4RZKOBbc+Bg179x9Vn/D
MpRpWjD1pe+xMJd8feoySYI3MsdM2JMYzbEpT2CzOsWpUQmPATCjvdz5z22A
BQwNydou4uLSbRTiKKtPLc7p5fZY7ohoeTAnBlch0LoOhcHJnAH22LzywMt1
ODaLkAk7C/QT3RSWvhyFBOolLZnHubTeJEZxurFxyrdmxQ9b9CTZKhmECqwD
9OCaPujPTtJdRqHVVea5HUxnlmxMpdDOcnedveypN1rk7TVX7/We7auEhf4B
m0l5evhu5CFLrP/Dy6mfvu+kIevAVvMOJ15aZ13RhiFM97Es7y819OqTCDAj
PEySGvKTe0guFfuQgf+aa6NyGy+nzX/FMgf/9flghMw7FD0baK9mCyitmqb7
otApGzaP2PbBFgXKwtBrMXuoAys15pALou5cmwifA/gtzlKB/qPZBhKUO0bQ
QMiy4+5GOVveys0qFkC5rh9GE9/5iO2WRyopnFWpb8wVzmdHo794UzCIraul
GZS5zTN/MyQ1arJqfm+9XvQY4GQa02EtaNz4vmxBq1c5a6Fm9mM2iqDVdC3s
ptJnwY21QT/PHTUywFX+94V0NTzpqj1CZD3gRJRnXD0cAByx9oV9BsDEYgTR
LWEgWEPEbV7FjXdPD0uXt0N2DCQWi2H6XBjlt6zDPyGl8Yg6xTxOubfBTEhx
NvCmN4DmO09R9XPBZjQKCJTIFGQ9UNf4HkZt3WUZlAJgK8cpjv3IAkSJQ9s8
+vEBB7GPhWaZujd+LrqiRSQvzCFGDXizyyxeZZF5eMimIj2EFYaTBbAYrIko
Z/DCVGpMtigjzqXeWXgfbLvbTgocGUt/4X0E/4ap6RSWU+MUp87YMW2ml4/B
Ppe8GDp1cUt9UoSum8wXsziQAaOEERsybRF+k8oJK1d641JtKVXUhRlgBZ5k
acCSkTiiP+t/dtk1k2QPY6mJnM2Jy8+4jsp48HpPWSHz/fVH1dCo7sP6ujqG
bePDgmVqfMZyuqMc0JlHUH5+Frb+GlNIkmEahA900s6gssdCFe8en5Caj1JY
aDP/+6Ner6/ympCEsktanU1FK9iyarEpxPA2V2le/rjgK49vKaQ1oF9y/mPd
UD79PHNweoamhKt8jcNKbDvvKSta0IujVcfhgPU+2x8kF34MGxFFYcU2FHj/
KSBqWOyZc6OCDpz2l4o3fWzodCJ22hfT/uTmTz3GveDrT8SBgYVnD0L9adtQ
ZubaAdazxgQre1dx8L0+mY5+TXgISKnyVvuq9mqhYtifj1WakA6+SYn1MQjc
lpvU+7aL0WXlZXuyhvTy91Vpka7cCRR+oIEHfr29lXQ+GQg8CJ1H+Bj5tDor
Ky62L+WE+faanwiakwAPOFBSXhAsrpvxfgxD0UDHf0jsMGBWVttrvGzBlGBP
rfQQBTet1W4SLay0YU2YfuxazVPHK1az+PKsC4dQyeiQAqplaU44k08xCg7+
E+VIkKwBu3GfWOnEEg/LQY7m+/ke/k/22WV3mCrxC9rPj8PI7+tmBD7o2J8V
fCCEFWAnRGItUiBz2kIb25rAXCOHr9WuVLq27NVZRfSBhzUAV4Fod8O0oCMh
FjzFrwHuItOX43F9/4ww7zj9JySBtf7vu3DSuEgk728DHfkRHHjRZAveKG+d
9ln9CS34+aKvJ1E/mZ/vHzrClNAkhDcjOllRNA2bXgNyj7E/povwmFVV+wEv
EkV/C2/VE8AT7igNd8TcbEiQdZXW0x+inV3zYUQynzOyRTEVWV6QDiGmKFmW
NKtuG8eU5ukXf4HssrwmC66ZKLHgeyJqfSkCJcyh1Z8ztmpGtkzM6imh9OVZ
u1QpqHjjQFlxWdZ/egVbz0XxcR80jB+Q8yb3yFWK0Th49Qgrs62iCwufsao+
sYq6b97JLWOy5/gOmeu15EWnkzxaNgAohnshhtGf+U6t15kJppbCL8Pp0tzG
3JeR5xSh+Lwc4rxJeFGWTmmfNIXE/qlcEGVOSeRnYFmCJIxjxKFG/yvsupmY
eXba7Xoize77S8zfiB/b5n5Y1b833aR+tRDxg04/sUrCKCPgPY194Seb5NGI
xkUhgiPRMtDFh6qKksWetu3yYf/nfjcIpVwivyKfaKKf9oCg4iV8xDRj06ml
cZ+KY+UoY5TQjZrfeyjxYljpqrsHmOpEYdSoC4RkgwgSuvXtuY9NKvw0bHA1
xmY7u2FDL8tlVGTin/JQPsYrBYSJdBJr5TVpEN/yKbvzLbdyafttSIj8Hyvr
iMKX2c5mGUOKpks9m1T4dch+XUxJfwUnTuGXg+3gl011vLZ7f7+xfHobdQp+
32o0z+iUoIBAys8vXEljhHqd9swE1hDDE1WJUMs6Xf7+ns6IyptPc5k9K+WR
OIA3uyJa4c+4QMbAlYlzepBHaaXGDHDEnxEgZCck5hyYhbtDy0SHrxnRZy4+
9doTXwfkatniw5h6J4JFA5pdXA6+IudeR98pYGK+DkkvisSPYLzzwSLoZJj7
rGNYqvgGbY3SX/dVf+3ek2agmbD+opwl4V6WgqFG8Q5WxQAwq78UdSjBQJxy
XZYqOppuyrfXILokiCW3OmTExxdolLNaSVO4Ll90SNoaVwLH6AKQP4cu2jPs
G+/0OzDxzA/bTs5kuNhGedwwNx7jLLVHpnCYjaDxRL3RP+fVvS0pXK4WApmt
JbQwX7XZZ/RjNdkjAcXXot78AxsSyuFRO0oAOi+xbEY0Cq/p2OlxFIPY3lyP
DIeVLt6ktlaUL2ErzDOkU7dyTLjbE1IlFXoeHg01KgCwqIiqdPZWir/pdtid
8cUvv88yYCZTp0MDh7PVeZOMjUG4Nt3QhKv2qXWQkK5q9VShz6yFNI0EMSBb
z3k9qgNHi/I7rvy1fa362VHC3r01LUzWtgr9mwdBTswaHiFLqHG2FnAofY6x
5wKGa8olANaT4TTX5ESd9kWQPSVbb3y4fHp9MXosnPiWBFAoNFZdAiic2uGA
CmJTSjM4nkbhQRVKV3RhLR/m4240+suwGexBkOd2WpOkmhxViDVeib6ihQGE
i5zmJRU4FDrlFKeO2FRhlOugrQMF3hWX9hQiepByMOqBD6kpq880GK1uHceK
WkNiVlKWse93kX7TfZjj15c0K82Zi1grk5tLGixTNWvYGcCDeuqzC9DPKWeV
LK7k/7gHZChQUsvCCNaheEEqbaJGn+9eXqgvz0zPnJ4By3dmUEjI8RFxqPKC
hE3YOrWPdKmKKpIdPBZGlHVuy7eVZhQwJ4efU8rqUXXRTo7IGzJPjRpzPcNM
V0zdB7Swocq7GOnaqZ2nYQvwVm+IJOtU8scpqZntJBRKR7A/azXtsXdtfSph
E9L5O7l1SqnwdXBVVrToHWKeoMEQAYxVmdMvo7JBcWhUskDYLthGJ8+68yYm
1RajKqsIOaSCwcb0YXWdFnBax7+48cruZNrf50FweTrDs41YFOuErjZ+Bnqr
SQjcKDhqThmUv3vBNzFWnLHmLBDDLRsKXl0J5kmXK0jIeYl8mVu3WeODb5wb
n5vdNB075NmlCSDnLjImiGKteqxNoA3hxnExEUgFznuaWLKt/HHt9ys1YGyl
l8cbOutJMJ7WS1BkE8mj7zfZlGGy/vQzB6xtAHpX+gwTCy5mM/Ie4k6D/7a7
4uOMqwypCzoVJ/RkWivTkTZfhC1XY4qgbj8KCvX2Nwr5JL2aaLwCgF0Ive7g
ClzjXpzNCeXo7ql10Hl/ZUfIl0wX6BI2DhO8B55Ub3omY2x3cAevuyYaoLaL
DEUVeoMK5yyvQKtydv0keW1xQVmKRPZyxC06/oFGkrN/fH/eXMTKSy/y05wh
QZPKBIeg2Ih8VVa+5J9XRYQGZ2ANaE5B3LUbHha2AqNwsgK7teaJe4p2jGU1
GMQdrRWQndUOjfPiK1Ojs0sLEr1hRmvXe6qJHp2N76u1i3vPp97L7hRdm8Co
Mrdph2lx52k0awU7JJSta5Al163glWRh6ZLe/GUz3OztS8nQF4I9+Ok6qso6
Ipq4tsiagHi2E7/e52Wqig78qNT5HUZL7BABBcQIL1rhFE5/ZN+/d6Wkk7cE
7xneJ4rFJPgyxNoMM0+/qDkzVXpKLxevCpX+m9Eg0Svauq/HIwWoJl3Tm9xE
sCDo/GZAtAXED4fbxNAIM0rMyuVur5RwsXlLX+1/iz+ksEG+UuJ+GsBila00
zyekH+jBQHiL/S0svt8kYLfzUIHmBG1gu/5/HyrjklMwZHpAh59r+QpUMfTw
9yxZQZYyOOAnkBV4RaxuMEuL8G0PsbnCzbqvnV6PLFG1JTXCJ0kwCxsT2muN
z/skDcchXyCQadXkQVHEzT40YNJSbg38yNexP6HWSXhZQXiXfTITikb35bCo
dWBqUlI8fqoNmhXvqZAxS1SJYMPsV8FLKMCGw7vXrO+UDOEeWELvW5evyvV/
1znCFKP6zaXi8lydTELfJNf6AGY31G5Ccre33kTQM/DH9QzlwIqRKwVEZ9BV
4KAvWznBNAzXIPup2+wrz1whcJpms+Ev5BXgzzmdi4p9h1HTYRNtDLMDGgbH
giTdiTevwfBDzXapsHPKaQtEdabdZxetjampDfXQu0O3MklDopDLu+gJBXxp
qyhcD3hLCA4FG73lJVmGLonvqlS8eHOpvC9wENK71hEio/0VRUPT3yAg0tQO
Mj0RuN9z748Fjmo5D8Ofi0rA7Td4n33UdS8C9jJQFTIgKVVl8P123JENpSnk
08JRE3mJwbJI8wm5u4PPoLsfBOn2XAkvgYnOZ+LBvhdB0na+c++PK/OyHh3h
iHr5ySl1uF9aE8g3LXOtnNwc8BeyYnpxDIKrSJhXAovDQn0bekO05aiqECWF
+g4jDJFAXJZZb4jIIXscBkk1MaSHrbUEcxDxC26+l0awSLY9t3NFiUS9IIOR
oAxqueHaDsNm0h5U5ez7urrPnd21yp9EvNKYYBlT2lRi20bNp1AYp3STVmHX
9ZpVO32uaQPTQRHFlnQ1Nqra88hG4VAtxOmaOjqilQ+4ylPFj5MHUpNRlouP
4iYEFxLMrsoNGKfkPutDXfhwJcQnJ/fNa32RBYJ6AfUlkx7dJMsgKzadPOca
kKTAB2IcNLhiNq5MLmPwb2llZfqrZOMV+rZl71oBBhVjAPwOguzKlhv1X68Z
63RTt6Z46V/xEmNbZTzvbaGrR0qI/aX6kzEowrdDOJ06IxTDNTZgf9WEoIIR
K93gcAwyKfi7T3Q605LUG8btOL2gEPZ1NgzQh9V30uC7o/bqeXHtuzGjWbCC
GK+uZ69mU7lmL8I8bAUguKO6RJuAk0f6rQb1GwCRkMPt1XNqgltAWYAuBOx8
atP7n56R1anx3+meYWAkK+mIx9ROnG+6Zo3pIGABR5kKPF4mUp6pMarrna1D
3cuEOxY7UO+aVBGpeN+Ryo6iiduRngR5XRbYYoKatTQy6W9kTtfojmmfUYGm
kCE0MeSeYQQJA5kWn0fLvltOn6Jw/rlc2tQO4i4mO/8rBodJvXSRiahRzvuY
RhonpvsmN1KNq92hRQZkR8PvybuCHv/s1R5pPMGO3Qr6y3hMV124kmPyt49U
kUXdd8/0r6+aK4xnhhzv/adxOfLJjjDWCvEEzxaCm+XLhxJ7jVfhHSxYMj7d
sa+BqL5cpbOuDWFFGA9Y3P9aI57/MJQ9Moy01SbGtRlQdpsYWI+cjvj+n4yo
/C4GGrF9iZZsc/6LmcLZ3AFKqbjbwYRgnetPxkCA70Lz7Po2blGvQFIz51WN
1FAENDqhvaDMJMxVG8KQ+PAqjYwJyFzzjYF5y7PmI9W2b4L06MZuGs7/9Vea
Pz/GteFtfRyZ+oOsul5O0MZ1iWENxDrzBF5OEYL8sL5VZajMnBoMr67yu5oY
KF2e2oWVA61OQhjd0K3NRKM/weVCXJ58UdULxwCzF6yAU6n5M9C0jjpRgIMJ
xAC2W11zsGReAA0A9T6OPfDmDWI/C5q020m/WSVTvKeKyvhN4sT7TDpiGMkG
LvRZgVwAcoX3oTR2fainpYBDjj/7FtTBRubSVt4WYghGQ9w70MqpW456sd3x
zbHsgieCASmzCwUW3Uk1kflR18h7ceQ1ip+OOSPtMbd59Bfuvvo57sMRrIAI
BbMz1otRkuG+C4zr8spB3vmb/mYR2Sk3W0FymNu3ZU1HjslO0pf1eJTZj82S
0ufhDdJ3TScH5rFCQ2lvIiDpFY8aY0iZsaNKVZjWmUmxwc5lZNbT7roGg3AK
ysEFkCF8ihHx+3hbs+wSvIiUQmuqwk8OBqaOUCHMyb/kG07pDWwuXRKcicdK
gOOPagAmfFq6aguHneyTIskZo49GffKGZ/vdJGaBO01IwVt3klO6TE7c515z
jcuF8x6QrXY5Yode2J9QgNylDcmVa+rauZR+FElxQRhlYbAHAL4xyDzHVD3c
tTBVfNzw0Si24/uctbh+MU/6A/Qc9QxszgQ9tlhP4i+9cqGIF5Xrtoho2e8Q
WYwk06MfRL19fUbAI2MD4cHA+nMU29AoZ0+N5G/k6FwYnsv7ImdOnX70nRX/
lItE2aPmTx9BBb2BJ4Z0cKlGhX6ZYPZpwpZRuID181NwXaBHUsOwTjQ/O/q1
ZnXwS+7/jZgzMbCopzFGhhaD1/H3OUiiR4rUvCTLiwPC+boggZznu56tvA1W
AIR0c497gAxW8+/XGkLm/D9QOrdm7oXzSdlZ7FnIc2ElxuK7P7V/hH8qH3j/
tUfOfu3SKiDMtlQNTMFRpNrM9aeK0wNJh7EPJjL5nuVxN9eg0daI+P+suLLr
EAz7SrAPyUoDYKYPwWk30Ud0wPk6PMnkjDtVXO0/qYpoWPpcnxp5es7j8b1j
eVirUS35Ujp45A+cUnIVl5f6/Nv5zTPHRVqkMqJJX5O0dw2uR9K39xEbNoVC
jm6fUxmljCte53kWz5AlVVplnBE3x+vt7yHM9Aeu18Q+wz/9XSwMPuv1j+Xt
CjxCcAmpiLEQdqJ0zA3srUR5zfTSZn4JT0lcRr1/AwcTKMG+iAD06CsnsOFj
GzuDMagYVzIiRcVqsHU+cK9wzV2QE2WywaqrXQ0YSRS3rd3rTopj4ih9MoB2
9P8bb1S1cUDdwQvQM1KVJhLfq+GoyoWn1Auh/n0RZZRfuDBSJ1ePqo7Uwtw6
WgMJ4G0fcc4FBHiTeJegWyTqmwdUyKijbv1B47j4vkVUQO5Z0sA+vmkTJwJl
rBGuAcJ4oFkVAdYwaTotbPYrnE4l+E28OjRpj+H3kn7Qj/Qo75gZQUTcoA+l
jygjrST/fTyB3vOdRsi/t7Q8I37UZxFyvLERo8wWkHy8ZTWErAsiTJ7MzF7y
m0Csba7y8WCEtZnAh6IuJKyrHBRN3Si5rsieYVf2CO9oFq1+z128gIu3GClX
qIWYZHvYNBAf0kjqg8xxl0EWaX7el1h3pP/aOPRZuqNpJ3EMAj0raFD4h7WI
j9zy4nPNkFA5domIWizp+2KfpsyMmWCSgWuoZj7x5CDCkShPW8gpXlx0vkKw
BjZnzApQbMMMAPbOj/DWhBkQCEoh5uxU9hqK3UbYkZgLsNjHBdwktvB/Tmft
GovhcVV+9NgQOZsnBpfYLPn1ziiZpryR7PzMO1AyApycwY55lugKb+niMQTm
exozID8Ol7RVb1GqiNxRDlJ9SxnofEVLxL3G3ExzOMjEUQSjnuLq1nLslrSQ
SQua40yD72rW1Jh/JBpjMYi/trOL4KUopsgDoj1hJm0pUBy6F/DT4uZ+P2qt
Cw4D9KTLqIfXF8jx7RM3dm+RZT9gRrEEtqw0az0SNshhgKp8ehqV9qSkXeqt
VGUOrStQ50iuJiT7uYyTBooT/0auz2GCRNpPeSkrIaONdgnEfRtIsYd3nvda
Tpe1bUMd6aP2x2GHyqxSTyR6x9p0FKWZjYEg2lL4jGdlp+eOsMYNXONzgQVY
BThPKMnpJFHB0y76zbB9pS7dSmubuey6qj3ZlwH1EocRiOXg3D5Up6M8/+9k
cd3qWG2jx2y5T08hOb8YJ8g7Sx1uWdihjpNbXKk8Z0/HCEJ8xQYns2VRoap9
uXlSMVyHaJg+YGq/HgZZm8Kg1S871o6PcSGaNhOyrZtJyDHvt1IjcilOcJ8Z
ccBhLNzMSmhIQnTVsq1xA/TuZqMh4VEWnEwE+sALmmmjy8M6TuIsPS483DxR
7DF7XvjbJKZoAWUCT3QZYB4J5jXWex2O4wgDBkIZgckUdTwgkdPslkZei9zP
RPO+c/SbJv+3+3ECYu2zibK4UruqVqQjz5rWGbml8+sR24H/DXHmRdNh2CUR
NR+V5VF/fOMk3QrRXW/F2wiAhrbfmi2ViWV+RGlWFC7sqAlhQianP0egaYuS
ziEmGriZgr+sd+RplbkoMDbljrEdS+y3YJq6JFZTOS3qOISfDuIif4tZPG/2
ALsJPuqvFy+JVHAhDQHeexj7B+NpFb/CM1LZbvqg2Jz6ICLha8f4XI2Drp8l
j/2luAAXxPropUuSLCW1C6EiuoJS83vDjHXGBe/+g82jv+5VY64SK4gBVlxp
jkNsQV1jBMuzctuMr1kGuf8DQ13fh6oyLfiwx5aTH7FhNUFYbxda3xHQ/Ddu
DUshqsh9LJm9vvzQTlLroo9Arxk7sE0TJW8UWVMmN7f0gp8qQEszsCXptaFc
QOXsCaVECouYBCPEu+Oy5C1u3gEEzULmbo9sjz+++R+YOye/3Zf6bk77z2ve
M+MMI67WKxvZcnCwQF9wikKMQva0y9nLBe0+x2wertmwjBnfobASuDIub5XG
IavolO5qbCZNYVywqFCOE+P/hRklTRkbiXUwQ/pT6zLiVsDpuaClA8yTxav8
QavuxdiK4ugqxKYXpaJyUTn/WGerl7P0xY87es2p+D76m9o8LgN1WbRqRWY8
uZEPwhiIsATv5DteDQbeDfRPqaRw7++NwGySRkzKQRYxxvItNX6MITdzBbGr
TT8AXi70v0VjqyNM1jNiMSV3b+oqjKIa9FGvNFEe/5t0ip7dRk7u4FlxwY0I
GvGCVEqvsfC8P8lm2/lM2CIGmrZHd+wpv3lzYVrR+pit9b2+/IfmQmkISwJp
X40U8mRJdNncSyIs+RqZ9rvKNC9qU3u+nscy1HX4vB73vbnp0pELjj2LtEXV
+cFRh5WzMDHOpNTy5X252VkcIdbQU+y4PxvRfOl2/4WiY1m7wgEcQazt8OrE
nS9jT3fkq0Qm64QlBRwcpWACKWKdBfDRKT1wvrHjd96JXAEAfo37qSiIjSxU
nN+yrKPxiL5of+uO3JVSx4kYOIdvH5qKXK4tVbNrXEtY/1S2JkaolkzepOig
/OcM6pmnH74TWt26pnrhs0rl4ARMS3qnmGniQiGw9xTxKxP2fwO0Wb4GYW9B
jbhVBr8jKQ9Bk2EAXE9HkFSoqUZX817FpiNseZITaB3fXXXOFSRMqN20Mjfw
7UruLc1umCMJpEoVKpVEaJsMqu5/WTMl3myfWz0sWdgdBq9KVVEw+1z0RL6M
jIOV0xu33wjg9KbIszF3stGQ7cleaSeZz00NixI9KgJO4jeYAIwGMD2F4Klt
aa0109N0XrzyYtVCXJebTI9Zpqd6ephDZGoP7yav4pY7S1fAXGWvaKNOevTj
geM30Dd+vw1xaPtWKy47Y0Z4l/JNYbDAuUlmoNcxYzhwhLXIVUQ7hZkPjUaa
VjfEqi+NWAsair7+gsMLV/qvmH+q+ycMbfd7bRy6UPpTQksTZJIlXRTyqReQ
8poyAA3Oec7gpaYy4HBCCSgRCZrDCBlPRkJSOuBmVvkVEN59329SsmGbiqlD
qptQSw1qNF1cSR6EnUD91H+z85D7P2ns9RDZS/b0zALPKynxj8H66wZmmXWA
7RXDtHGEfM0/X7cK3G9xiUkojU29vTTBavjhgRzM3NpBtyQs+Cy96ftDIuxB
3Jtbu1CgFAwev3SIjuc+sIT1sVGgunAB/zQZ2JFcjpKx1G1BzouFLRSyqTnH
Zw2q/N6ryddxc3NyHbJLAFv38+wldmQfcii0c+gWpjFGTzbouxC34S0hJ/DZ
ATohMb634SscODSyRFlj1YGhwEqQtLlZnzfkN8iFnJo2ASDO0VPg2CXbQRGi
YKN31uFCfJAeQWbSOKQK3yo0fcejska6JLS43dLHWN9TYjepeox1JPxQP2sa
6Zz+6soS02nggVmcepqg6gYb7yOOv1ekeMkbaxAO5D0qd/Wq0q/IkN6iOXqn
1O2DOg5I1a/MvzaWHHAyKRU3x2ZtjXA6+Bfs79cdeHVSwegb8s/IpEn6Un8u
eEe8vl320vLbo8IAm5KkGh6yJvHDZAcXc29PNRG0I3Xrr6V0VWANST7Hh3Bh
ZygD0W4TromLZBhs5Fh9WurMfWqM271+OIaO0LfbDA7LxSO21RBW7E5xvdZI
wE1SaygoDZwamAICYs9sxr13/oD4Crg1cSURt0QqJcgHVc4MEosptZSwVl89
FRGCSEAAwP5X/00VTuLPccTjZkmx0PGybzp9mKMyQq2aEHn8UShdYdA2bu67
SeMcop1YUd2dfGm7Ixg1nn3Q5pGiRUzz1U53Khhap4daaBl4Et9XIV5h54d0
RmfcT0YA7mUc1VsFXu/vxNuVnR6EE6K0e8JJu85LgN2R2Ktj8ZECToqhgP0w
TlCbDBFgULA/XqhmKd5iqFzI5L09bJSdGs7Adaf6LHI+oRIwG54xYFpgBnoq
YwbE7+fY+hzfATkJ2+3gLR+LcCfr17mj471BuvorG7yltz950P3pobSHa/1m
RkrZUNNAvXPyQN3rYwkZCfx8M61YJL/Bs2jE9EstVIQjUiBZn4J9U87wZNwr
qp9JsAa0xSCeI68ICUjghoVmhidzZOPY/+SZ1LsTnLfnPIgvv4RlcvfOg3Ty
hIVs+eI1f8RT59pyDZT78moNfiF5XXCWu1fWy8p5Mbl16r4b21xOt3yUmM+U
NqLsmsIjn498x0p1K7y7dD1wxQUs9MP8zTYfWYZdJyO1AHe5Li5ildu/QoYQ
NryeGPxhrDzPg+HM6I5cP9HxpghuoZiFnOuClCLNxHf9gZebMUZ43hJI6Z2/
I8daHk1tdflFMlQOIaB+/9fiXxyCppgSSq5AlR4xV3o1OQL7YTvLnStQGIhj
M8K0cbT7Z9fhHFulMv1+u8sY9mt5JNhQK5wkHVa9K69K3TlzdneUGREVqD5K
SdHnuwvaOBnjW2pO9rcW8C0wNNxPGkwGZxpOaBKTYT9eL99TYHQbzDrGExnP
xQxj6n++UgIBQXq9swnX1KTaGC3QX+juRxmnpgVs9N8UXdJnh/2hEZtmKTwN
eAMZP1Iw50io/8YCO3RoSXw85Ierh4c1zPHtzCTtM1BuOyIcuRKrsjDRPeJP
WMXqNKJqYoVAO1ugyBaC1XP3kkb0nZoaTxS7U/S1XuiqeeBFrCNO/SkdtLsm
45aZt9MgNrCrOnUbgJ7lERRaAzI7oS3eJvk6056GvHTuzHa5Gs6OxFYlVU4l
pgPkDEStpDB2qauACwlUovVAth0hGVZz9nYl1RDXIbxpWHXU51aDxF0S1yWp
m9d0VRW4C/ts1ZNNFSuzmnnBn3jBqfgTabzAFs6Y5gMfK/6wZ/Jat72Rhm2l
7IcZJD6Tp+ll78wrtDmXhMBRa1SkAUbM8N6YlNGhLYfl3Yf/2BWRaz4BO/Gy
d89vKObhP02ijvOPkbG9PR990kOsuefIEOXy6ajN6chYwjzamP9dsgQp3Zsv
3aYYxxpOSdsO2g/FchhYBa82hvznlXf1EksxiSA0E/8a/iUICTIQAkD2mNsy
2A8djYnb8ui/mApkZVJbXGDnOnpXEUwpqk+NVXKMw+s/Qx9FCc4c9YwbnKEb
YfJBDwKiHNB/SYUWFS7s0Fkz3JSUsF/F1u5OKYfuTYY0VUf+jKe4b1Pfet4d
4WaiuoSClHh55y6Ql2Z2jTKHUYWUEIvxcbfI5N4B+uAr8v24UtzZAjoiOYyz
3nohyNj2rbSM9k6bRfnZ+QVk2boeMNSe8fwjTK1mkfci+14qa90/URte5/r9
m8s0uUVWUPT9V0UG//krTlEjhnpeJx6VRfXoRJP1gSmCe7/H1V1i42vGo0b5
C7vkHxgd2LW1VdForsuh89GltY0o2LYPMDott7M5qZykcpcgjv/zVeFNDGYU
y8bTBvzmv3AjiLSyQlReI7m2+Q8mXzQjXXDnjgM5j05IE0UNcrSQXqX+u5hS
laesHlNz0o+/ySwFaE7HwoFGl+stLjKR29QdorAUfNRuGQWsLZnfWHZLekJS
7FVMc6CLuApdn835JUirAX668oiK3PB6i02DeYtVjwfXVa0sxNfRj+e1HFHE
rJYS2E2o2vfpraGt28rxl4V2BM2PsZPmZe6bUdVYlgvwJbaG0oDJrcL4e7IF
MsE/VnqQza6e0wCg6a2ezFhG4ZPGZduLKB14Qv9oeRhGKAxXtUvKstJSo/eX
2cfTmTsL2JmA8hGm9Gn7ek2iZ9s7dybc0J+N1PS70l6jv2DZGHWC7j74ZxHf
FCempUgmRPQKQuV6jTF/VLnDJF/ahUIzGD8542tlPhRmbToZYVkdl8x69pvQ
0ylhB8dmUgW8DIm79KZntmeTmWXMmaqzBOTqEu5aOAOw33kPWivoLHqpLxDQ
IkKHeqr04/btH2rfXKn0rtlbXP8X3bjvq1mlwY1uDvG7dWauwnDgaUAv8ppc
u2M4RiV4iBbBRgoHnYf2ceJyrZmad0OOuSgDs1pvjcDpayVT1bwlo0+0AneG
PJeGVyAOZ71h3cvlkKrxVyPtVrgJd/htLxMGNgUcbHpHc51SoS3urYV0Tpl+
RGddYRUWX2lG8EDbmyST9AdbwLJER4UHJzQ4HGZP7RcwPC/L3+voYh46kBmx
+DrhYvEBF8hmM+GUKuLU5aLy8basEcFU43JP4YBBt1C+pMPxPKnlsjYmmuH9
MS7OEn5/uk3q8TsR8d9TppWwaS0VK9sJcld4w5wVkFYvaT4s4ZztdC9347UE
YFJR40ToXWYlou06CcuTfrKd4bQrimZJs3RHYwFMa8/J4xTKztpKA7d0HGPC
JnIo04DaK3n8D5lYFeT4UscMoZnarJuFlD6KOBXZ8OkZWnmag7rFV9UCWP4q
hK8oKn7t1/YhPy77Zavoa8YZrGX+AV9iNuAxTz/6xQQ0Ur42/QAxGaS2ETYn
Am6Ayj7nt7SQ+NiUC2ipCURHKIHNYa+/ibhx3tylsa/zMlHDXd6msOTVAKMk
EVGdObKu19Ti/vjbyzqfJTIezXCDxuWi28O1Dtw8bQ+bore2YkkdmgutnPQB
qJ3EphO3L+ixVp8yKwB2bEH1sm4Ja9fk2dK9haAvEWGimp/MgxEimGIT3Rsn
H+AYsnLAFA5i6D8DP4yfkHlx7zxcKlnjEF8RRYUyWOBUfGcKzYBMLoAgQcg/
jhwBesFAF0OnG2DpD9DhSeVdxMxYMKh+9Ph6H54G1GHyR3z6k924hsbI7cDA
mhT/ewQfrt+pbUymSqwuezOgReBIfhpnq2fAyglihzKBOmgTqr3GL/GVO1er
qKm44/URTdcb2pvNTn/FPVVfqtYtOp8+uKi4syU2YgCRH/Gmdia7t9AX8E9n
PV+ft0Rds1WKn4UwMKqrbwsoWamRzFXWVzg4SzSnue2COM43d4Rgk7unQ7yK
U6zKHw4Lx3HwZlnc2NmMJCYbVGyrMEX44Lti4vT4OPlAmWXTI8tlo4WdS5+A
XxPLXj/HuX0B6OPi7IO2JNG8mP3qF0oUkX6Szb5pw4zIYXv0CjuWf4cO6afA
m4USMkfYNHyIbDVRKeZ+L/uZ/Gw1FJTtX+eU6Ez5jMqMyWoPk6ue3JD7oN8Q
2qpRPFtP2at73e6fO4BOdTe58CToVwoR+a7QjfREWePGCzjE2hIcqhn7YLIe
NBv26J8dZSBnM6M/P44zVXG6ijI6EdQm25kL2z3EuLmRR7LK0MaTb1aFmVqk
jHwIuyVLAcbmZaTsRCF4ZwLdov32b/5iYRuklbBqdWl0ob6HiSZu22jDNxOL
AYMwXl/sugN0+ogVxkKKQzGVq0R6F/LT47gs4jJx2ovS6h++3rqBjKRL8GDl
tySmZskqvbzD1dR1ZJs3NJtaXngOHAuywQ9WbIriW+FsRwY4EE224/GPARL6
ujkEosJiOnSfKE3MaBhUvVUBdkQXiUPSW3hj2usP3ifRcPqeHH16RDhe2gzm
QN31MLmdO1B4/e0vKG/4eltBkBMJTIWNRdA4P7AkWGe/2o7OV2Hg0KGhD28F
948OUur+WUg+vR8XpgksTVTuSS2IWCp5dhi73vnTfBFB0o/bTvKZu7OVRt4F
8MzmjO7RnXp8nYmX12Sq8jOTLaVTNVohI/Wdhu4zIHylZXKo5PuspgiDH8u2
YjkybXJPo1+RqpoP8m1dDUVs2kssZxMcXNaQKAJgCQBcHbPDsthhhT51S5lo
exjpw9rhhbHB0TyTC2zyTC3j+yvudjieY8eLaa5qf2l1k/3Ueu64P5PRsjHJ
bsrTMbhWzQdcNlT/5uMf0dAK0gzL0p3LcPLw0N7D6apz38Lt9BZZTkH6/bXW
CnTltYf6QUgmgTdG3O4X0VanxoAU7XzpYPoGCliElMpWHzcNthWcQ1Kvupc4
bhR7ZX49mDfLiQiM10DmKl8bSHNCEOjNT0vsrWT2mqhfwqkqMvvO/Aci64zL
UKCiUC2K7tMUHaQ4PO81vTOsIauOFGKastoPmFkgsW5dwAheUo5fR+uBEYDN
wYF0Uhm1yGBzYNR51wR845+WEngOLxGDScpGEmSwyckAwUP80iEENNfVO8VH
SnuATPdQ5+nGqomB05QULL76MiCrOQl1VX7VzS3IvpzOBeA1eH7xo0BM9wOQ
a718s3zfvdyNVBB6iHJQkvyrFAY3PEOxNnjVDiPWJzaGXJAxrPeJaazOzRq8
wr9/73xPKR9s9wpd+Czt66XoSYRdeJ006z4VDhgeqsFyt+r1b5NKL4DIVgOY
03kgN1GjefBdeKP7I+nA5oPP7xUMNWYXq17vI/QWSV+seuusg5U/VlhBcHSf
ye8Bs44O9QZ0wysVq/iHSNmLuyEAB6mu8SXBLXZWyhuZGo6FoAKV6nmZuXXK
dPW/h7uQC46g6BJxs78PYmR+d2VMNX6yWoC6hbGceVI9BUq93tPf8WzDkr0t
T4r0I8jx5YlSccWGrxSa/mE0g9BruvdxSTnRWUMkdnfbYTL647OJJqFu5N+g
a0NWEe9EXOkPNzHLXKEp9w0xW30j/cTRfi/3eehXwnZDLwhqTjCpOqHth6eJ
XtD6gx2BZ6a2Eu08RQX0V+ZdUwEQ5//N/wQl8f4jUdXAmmptRJqRCNMg8Lr+
L8NiSERdoX6VUMWiBaP1DFslThzf56CXJuTLKQgAICt7CAchWLE96bXolpsD
SXVVMkcA1Zmcgxpo2j0GoCo50VyKrG2zFwp/S/CCmomQuq5m3NOrO7eeva3d
qDM4eJZl0YeFc+W6Agk+/zg2TAUmhrBjpcMuBSpFPubUAMzfi5RhCk42Fy9/
YNaopbNsu6z2TtayIRxyM17MH89GXSkVVoY8Vm+m3639z2jhGC0DWJoRwNNT
sy+ChfT2P6amOimLgttQKSJ8ISehfBqtkpYouGIdO4Aj340DtYHwq4qQpMPC
tJfnih2LhwlyzKk+RBtZsRvLoodgZf4nANZRs9UlZfkqEh4hj6L1LnPL/mj+
WIUfOcecqgzTVzGm/dwEj6bcF1msIAGtkD4vpf0msGDPjpBaYipY2oCDP1Wx
uFz2V/mTdQZOMGw/10FUKFXSX4M6ZC+lCWHnsUttGW3igZHsNensBqewhcI5
qAjZVej+H8/+JBQuLH9D/A6O/1ajF2TfAqCscZf4sidIYmgHfmG7+KBSGPN9
C+Er3toQ4/77rT0c6sSICOE6IxgSDQJkAujOu4crUD9X0x1NAcZX8hZEd4Iy
Sk6pTI5i/3JxpZvwF9ONDqHNjbxISRWMWUiQXpYO9LJL5OMN2yEfvJd8o3Ir
/gX3wf7SV/bJzlblMl5ogvLKdmSqN+44zK4tzstFkSGb9W9skB1riyfFHBak
utkIGcHFWxkZviQox/MRi/8Rm1szxBG7UNtw2Ymo5aVIgOCSfEsXQvL05Lby
b3/EVN/niLrUzqb6P4fctHeg0Vplh1AOpSFoS40p+O+l1GhhpsPRf6RrOwD8
mCrdgCeiIPOeGm36l2nEbyI7yceGvZajo1HK/HE4gngfh+XSdbRU0DnbFzyL
SjWNuiHY93IqCIKQVAHHrlsi8GLsN026og/VDqeHjJOcpGLOkDnIIgFgLju+
fIsK5xcc0wAGVEk871Jg3j3QwvcyKM2jq2EFatXkvr6z7F7GFI9kIKLQ59WJ
0jl0IOXk+iLCm1tYq+WM0vrdjGNK429daW+Mbp58UQJ+Qd2UzgmoWscvjQRt
EwcmFOqirFaUCVrGg146krqV4d7zAp59fg05tmSjNL6PVPcdt6EP54JA0qFP
xNLic5mN3cNzIOQJaU/ue0LVwSWE2BFJsKXRId4DQ6bWkkcSstHqzfE+wLg1
KLGpl7B/JtWO9BnWByQEyBu2HRI5/3O6dFWbZP3o4Oyi9colSIa6ngH4Dg2H
uXFuTi15JYp4EGv9tMTcP/dMN61eZZxCr8AfQo9foXPvE+rVKV48nB54q9ji
PZqoxlwc/14Tz8xyeHwHLp8hgWhXRmBvpLsuOYihqFqEZVelw4ei1hgO9k7a
w8CZBUQ686iGMKP9NHY3C83cUyMpl+5IWxxtL5uIum3vkvHyYniee0s4CbjT
0+uEQztMgabLesAoLjmPeeMG+o8TFi19z6gf81xiGJdgfBtqvxUDX9RzZiBC
NYEW6n38nBH2aQvSg85b2v152eXIn0SRohrcS2AGV1CAwKpRYHOb8lSaNI29
jIfDWa0N9MuBswAMSM3f84TJCRmMOCIksBBTSz4bjekDx5A65LbTjwd7pG+P
iMpasp6GIoAzWViKO0DPsWuNZqGOysKllison80muofJZG09LbFMQzp0w3yJ
S/aq1apx3uQIV61yiVrrNXrbJwLctiJ/69s8IvOc+Z+4x/23Kihu43AOsO38
KFzztZTDXlv4vzwB2iQY0wwF0/VnB8jeeNyLniBmUBxHLpE9Jm2QaUzdlZaw
eBs2FDB1rLe42XxTkEGmPI9gJDkvfyOxKWI+chTEQmw1U/YCAH8gtysFfTky
4jJXwV3kisukccuTPYhSwJmWrMj+55KBLUn2EOKEk0aE4/7lMh0tD1RpX9gs
4wxUhU8wKOsq+4E2DOmpzvfbNAo0m7UwBIUQbgQEKpXe4AD6g4Y5PrHhz0xK
eC8RP4et01KwDJLnwK5tVRNjNoWOoTED9XdpQ72actPGd4g/+VJ+9rku05vo
uGZWTUcr1gOwSIXgN1gbzCyf/hLqnsKjsrYRzzBgEPNgUooCfgkKzhp4OCkK
qhfS5AMlU2HQgP+v1i3e+GXRZ5+7YRJfWWSexognGOLp6G++NQwcxbJWF5MN
pspq+aJAjbMyg2DB1qfgsbFQbCbBc3mxUc3nMvsUpR6dAcD9U1kVfsjgV/gJ
F5ipygXo2UP6oRjVcso+TQl3ubqDdk6BAv3zaNGj71LJ49oUusuVxRfbcs0x
2w+O3aG3zfnOqWFmVPKjYkdVgQNknOiGMnu4hvp2WnGtbgxJ+fxS61RemkvJ
K18jCJDUYyI+ijPdhDsMZz4dJOelYDYoSbz0miziNiPkdZqiwKPFstt+cbK/
WIjl0z2sGeqtf3MHrl9dwuWnolEMH5oXdeXlubTMgj88lVtQOxeIleMGeLrk
eNx/Bx/lzF97DKs4Is2DsMuhw/UBXl+mDwlkoKwELxgjZGt5kbJUE6wQNXix
PddOU5EeidhbMyOFfW+OmYebeBBTWqAVFod6IpCCBdduXsN6PxZNr2QBkT/n
MhpUkh+rup2sNlcUCSBRHq9SSXHy/xsn+jU3krl7QQ8L4T2oYMJeCJC8ERxP
lmZ8EOkuiLkpKw6+mFpEVTVGem566ug+6xri2HZ02pREixfC0EWPfT/g+Ya/
OvYbWC5aoXGVl/nhXTHnQjSkq4qe3rOjF/N24pLZ5ZvDdy92un/eGOgqZac9
8dz1XjtRDslxh/BwWvsLaD0WxfnPj4PrO2nVIs550sewr/VzaYv12srXfv64
42gt7tJqSfQMUYn1c/Py4kabvRKGFzh5ppIz/Zn/PROoj5uHrdrW+OSVeMfr
RIAL51wQ2sG6P5426fGzaZNGWaNioUqTieQcUqEgxH88f/SZcaUpD+CoKnyy
p0VtO3SUUh5/zZYAx29Tr/Z7VGJhOlznh9XopMSNDNeJ4Ye3ZS6RQdI6Rbvz
Ny3Ufw/I0QG3wBNiyGWgT5bBhB5RxfbmsaXCascIwZ/twta+3DP3NFRqVPZG
BBFGNuIqtrbfw6qg3bbeXSRguAO3Hj6+QmYPSx/ch9CTTR5uSrYyHNTGU4Wh
ZeGeHfNJlfzL13K/T4u3O5VNtarp4nh9soBLj7Ngb7tVGgQ1ddrjK9Ub7xi1
kJGYkVOQ27UWCLEw/F4VdZ6Nr3KEdlFq7xU33Hmw0VxalS8HKMj7EQXVjWYU
l2a/rFbAwHoNhYjkFSVtej1+xWry8w9Ey9NxiuHIfSKd6HnnGp+6BdBEtrLM
BDouyyZLlMUHwdXNf+CC/lDyqPBZ+5SkfznPTUR24TpS73oqMXRl1dl1qTYM
xOO6k6/jFu/VB4BdSukaL0IiNxdTRi+s4NFppQWKDoYv7RBUgoB8qT9K60dq
Z+3MWMSPAOIUc0zZ2j99JPY4741Mub+Fvx6Tf1ryb51ymmTP2VAz4k3hMOMC
SdKcHhijL5KIx+5ZiRziEuFWbh04j9jEyGiwie9+bd6qQHqew6hIKtHdDYzy
Z4rtMKsO8RrDnnCgR+PfiSFDdEepTrSdwv4HyDuhDVjn+vnkHF1xmy1wnP2H
QKjrQLxVlGDzcLnqLEatCrWYBKVM/zeXlUeRYAkLyk5DTmgid61YEicDXAwO
Z91JQF4OwU5WY3NA+XXsj/9IevlF4vTTun0M4a+JAc8kCtR7fCrJZqyboWFT
/49eQ54XieNGbqvRElgH2p/twbE19TNtbXEOdt64jY+NJIAKIk9S9YJdqeRi
D9OBIuR7hwMgkDPbR/IDPHQPI4p21bHEZfvaOVRBWQc60sQ66ys1eM1YUfig
t5q2xh4evP+vOyUZMMkyP45rNZ8HpTQmdTcdnh+IjZI0CNnb3LigF9c0BUQh
hx5QzEhiaBtO8GV+QDVrG9Cc1IE2hdPwmmRYbB9UYhEme2ihkmtMKiWokxMh
PaZoUKazAP9QYZixo3Ikj/x0Gw5ZIpx2V+ckqn+6YYoOkRRxG5AfZAIj0uDy
e4M+vjpQSvLBO+As+AawVVOwiEtafTorTKre94cjKqrFe4fCnsRP8nf1yZIe
zpKC3QJH3uyZg8xtdM6MJVDIAUoFg4arWYx/Vtza+jeKXmmol1+st4YwY+uu
HtkLm0vPmF8sxchCIwC0XYlSESwHVM4Jm6HmwfmvrGjxSVO/hKPadj26ymlL
XD7BK85IKWyfjM1EeRkDFdrDfQCN1bP0No2whdFBqe0wO6SbrvI0FFSVZijb
UZ/HibuiaBFZ3TlcgbR8dVo7VnQkPHqRaswQffrNnSWROdLmstJGrxgMJTZB
rF9vXllF8Ysm8UswAbR/icgiws6vXTxsyVbrz2poLN+DjjSOA3dCUNinbNKM
YqLR/qSruJuCMDWd9n60oyZd47fhS8jb7KsIgg4JY2h6acQ50hyJj3ZGubQI
8NlX3gFoWoKbni1wjaERy56cI+M5SUpEvjw+1pNHLr6NcDUUCv991LUCUMep
CkZSFVlsil0CKcNjp1A05h4cWCKlaUPsRHP1YUwryNu2ZUQrNNEzy/CQcoVC
w+iYI9KwjbzRM5u4L6wlI6ZDOf/WT4ujfhrOt9ZXQz6RTG458oYDAOyCuVjO
3jaAEL76Co4x0sxDkiykgN3ek6cbECOb/G8C38agBBW4x9tqMytHRdg/nedt
rq6sRWfzjlAroh/9zXjm7TWjjau4sM8xEB+txCFAvF5SmfjR90Ag8WzxcPnm
wLlJmnR2ru36Rn78vJN/cY54sEOLf0fP/UACHMILA1c0tzQRaRfwBJWcdInE
DwkmofKRZrD/nMUhA2eDDiYy6NpraA7F93pVM/70c/Fnbh33IuX8W2Lhrjzc
Bci/RzJuWEd1ay0v1CQlR2DmMS4+xsy2ax0I+mj29bCa6LAq/XQ7GS0O/5W7
fhckni1JGS2SygjgNqX4QASFKsLUnGGl1TlOz0FLjQIsWEJrTmHmm5T1iiia
eqJHsit+06pCbbuktPpvQYmlUdGsFmplqRoC3lB3yp4FZf4Qz5VKLSMEoqe0
3DQ53HmYFPUQeQILqsKjC5TwlKnp3EJHX8UsCTz0h3DTqP5Hhk0H2se+hAZE
7OQFUL802cpwBJ4kVl3mFgwE/y+VrLvH+ea1FX38MactH2qx1CPq7bIvNF1t
7elt150M1W2EPiIGI9wSgdAtfFYubBZ0yj1TugcMkhYfSjy0gitNP1DlizuX
XTsN++kmoTrIwzru7f7yUi1BEMiN1NByGfn4q/63SAcEWyJJomk+ZGANwLvp
o6OKollUyeXOkxAHo9J5WGgCrAtJJwh6E8o1CmbaNSxPr+DyGtUvS44epYGL
7D40Kgefpoqx+6ItRtAvuW1caZvhx0PYd4/SEDuVXZ2sma1payEDCO+fqIhv
ZGoMgeJiL2bfQqxdx6mpbtBVfhVNtnEJ0MMYIfAn3tyYY0GPu3a73U8EU+BL
HUSeooTR0A+IFn474k+g512RzJqNZWFgoUG8o+hQ0Lhgk8AC/M3j24TEgkDF
cH6E9muTMCKv62rXWFnxSQqB86V/BMLydekhUnsOdTs+lF2cjeoxk8evpXyM
RP5O+b4UoBHXFbGsSzkvc1m1Urk1NpCFiL06/pUqa99esCOGUMbyKOL3Mmlg
rqU3V96r3SyKvy2ypu3tiBxNClUvdiRFHpb9/pVj0nFftyOE7iARo/j5kbwF
YGR4iCA1MZNY8h8qQUqrlvMlISeMWzLzhmmeXlhFMQAA54fjOPPv8UCjiwf4
bzTm9u1c2BHi9n0/bnhVrfmy8Zez6v+xncqIl2yoa5P0RGPfuW9j0m6o69iR
YixOPwDtaJPdCdKTSZg1r3+Fs3Cx6XS1om/dVXnP/LZqlc3jn9k+a4KV/tXP
2rUqjK8JEU93Z171WD1r6osxbOpsV2CA03REjen+4sJG9kJq/5jAaqWRHA37
zKLxMPCR+WzD+CU/IuNH3WAlSUZ6ipY8RPeBq0v6pRK20LBYm3H04MCRR4Lq
cXtqMmY0UGESM8FifTxQZ9RJvrliZjLXg/od0bsBn9jgzM5d5VyU2eip2L6H
YyFtTwW2mAKCinaYFYxzvTk3yU0MCbvnJrxFQzqx4HccPtFFExluIZ5BQ5Hy
QLrExrsu4HTQ5O84nmzO9W2xC0KlQul6m9hGroWdWZSYAtwXsdMKtW2JYPG8
EMvUK2i5z1NmvZ7mHNYbK/WxeFM89cXrDLC8ZRmv0Vc+0QLoK/iM8xzJQfDl
gDj2cNkG/vOZBIr/5QoqaWPJMn44eVcE2t9vPScvdg8zAPvB6/jU1FixAQJA
yN+jmR0UwYCsvhVOhPJY9NwF8+nQ7f3ja1wDOKvvHc8mjUH5ureOdYX5JITR
BiWTzPU9KVKl5zgzWk9T61+2Tm98GbS0njb5sw2RTQ8e82b4lNNAkrsqI3+M
RxegCNVhPCOsMU36SFbTCVhL/Aj2bs+6IFzvJ/viTjKpm67F85hqjfu3chWJ
SrCy+p4a2FXccFYblU+BQwxruCzf+ETWEeAb48w/w9bcrJlcWzUv9/Mm3bP4
1lS73Rod0apzlKYpx0ni6+DofY3500GQX0jUqM2zpbFuX3/8YG+Vs7OcAwIS
p5vMLYgyi+zvn1NbzAdqcdbpWzZv29CcPyWMsTocnK8CBq3lxejnZTSM61C/
yDT+1NkHFlEZlWHpgbrFTtGHCWt5kGZMkeiDe3ZbcpfJFkGHPSzTGcUa/vfN
41O9JtCCZWBPtSHSmbsm9HFxCBbu/RnhUo9jeX7erLFzycw2XvIp+p43QW6D
7B+a7rDMZNPcADbXmYMEVysJ84PMjqdpIxYVP/RBTwXfMjrVJ+4MCup+AlG2
dJilYByr4f8RayZAhor4zoIesGR21SsEFSZAGkUi2DB63r30UwuDc8NyIKwB
sD51F9VwmMgCe8EYrM6u+vq0BYF5Fk9eatrf6Yl29tP1P7iyPWKweCjcMazy
L2Uef4kBBm7XZa/vCi1i6N2VPOcmGjxqVch6qxpOrJhEbikgO/LdC98j3mtS
SC/XQFNXJp4bOu+Vq8Gu6VQKHCjqAzkrfDWkCV1NjDExd6xUXcuZNFloEfqV
pXZKYYcKXXF8zNhtqhyT74DJFTzgERZ0uWkTIfi/o/BOzY8CBalr1r2ZFJ2K
DQ+uIOvVTtKOz4nLtxutqX2nm25UK1H/XqK94IUK4kU8Pn0wdZ6bXeBK/NeD
wThKzqVOdDGNXEGVdpS1P8N07e+G8bwhhupJavLutj63l9MTSW1BKAwTx6bi
zj7r75l8SdnIu6p64+ZINNVevacEMTPFWBdh8ajvSjjlib/tV1zZsKg8S0NE
ZA308oTQwSwEYH1T4MFCBU/sCdVH3q/j79CpSV0nlKlk17sgWDxZTkWhHbXB
SeX31//qIaH+TaT1ZkI3OHrxMbFmRG7xqX/HJVkWbRJKUDfzeKkZqFFn8SSt
21KzpDApBioeEV1MDRZRgSXgmihZSGCFyQrjVzh4SJ9uV5POnSNRYuTKHSi/
EjH/FCI9uFh+G4rD+At6TmYtC0dCnX62/+B+Ib8YxTQ0IDXp5vcn++P9vRIQ
KzF6NJpboFKw38URZlCUOL5T8Dtd5zFYp0SGUbexQZwkIO2k/f2lGqz4+dBn
IpKKvU8H1tf59lmmKcjhjaf+LcBWenv53ZS1jiVnfz+n7wOsOwg/XrMwxejs
5fSO25CDyE0juJwyC+2gqTE1pLh1FDmtlXvbzBlugZDpAqjVv8B+UTuudSqH
jy0WtNkvQBG6qzY/Z0DnBVFN5xlMRA87Xpe4jrFUPNOSbttvsoPNjufHNywi
UI8gosWtAgOV2jhiyxYOMEgVZg+9ZqYgblRU2UECywF+RVR5nF36v9lEOBk/
ipxHBt+IDPrGKzKPYXrF8QpwCLzmN/3Q2kJQsNb9fPhiDz/UmMw47/YbsNCS
TxelB0WCUTaMd37Yq0CXVUd7jQe6ea55TAipPcHTYOe8+fowpxKWNh+/V7ap
XxXgc+uw6aiEWEsTuZyctWFVMw1YCBBe8qcnGPM9f1x0Uo68x8+rO2fzZMj+
aACiPLAUnZ5HGb5OnJKbhqcxhQ4hgv+av/URs6aFkesAiImGhhdKwEOJa0ih
TBW1VtoJ8yHy3/U01IrrIVDAphlvE3pQqtgLDGwyNqwxYcMjf8FuVX0WNBo6
RmmzdO3x6vqd4O0FApoPUSH06hB+EivgP0+sOO4ts9DqszTGS4FNvsCrSNz4
Yr3OB1iUr0SjTr5JYdk+QVyHxkivv7TrzOEBeuvTBfdzxkW9J0HLhwJ8V1FF
bW6TePuN3MNoFyuBG1dVK/6x6dM+Oo1oRjynKi2pl0mxnngeQ1yL7L+svnRK
UmAJh+g8COUkMPV1UCFWHLhqvC52YR8jOmAO9IoL+sjPsNLrf2b6INU1t3qz
qoZjnNDe7+fUyZmxiCwcfvZxMdlU8csVDxp+MyCU1pu2H9vBzE6Z90YU2kr5
VxjIp62ExXKaAl4gex60HrB2lS0n9eZqVCe34OK8SRz9/kAfyolpsjxu6Ah/
a5zG8RZlCVU3Q654T57Vj3GFr19v74bmMZWttVBSLryRdCvchnIRqgPi+jWU
8CKiPwoSsRulA6jLrA8+DtFWBqIHLCcbRLRnot/rKSZQ/VEt86uOoOca7fw1
tx2ZoFMMs7P9DPx5/kV0qTZozMX+OhlsFccbAd/344YN0YJblAOHJ9OsGvsS
n9vFMAdIXaECRkApFP/QwEuyZoJ1j4MjMApobH/Ss7PHbJWwXl72N3m5cu6f
76NasNw1cHE/WTDjRY38veQzJPpi8JT6eOzn5pzCPs1CPMb+PqDGKJL20OS2
qd0Z1rK6KK3cZMPLBxjmfSJ9uHd8vxX5n8qH5MTaYM24WXx+NWSu1JgWQU2b
zuHYigBsBCdOkQzLZ3sQ8AMfsuB+ufGnIZeWEuVub4sNO3jY1p3Ll+827z3j
GcVfKLJkHPEp1PUO1r/EnpzqQf/9vJd8D93QIdPStNki/EA3b83i4xZ672bU
9xBTyS3GAJAAYHK72g53EuF5pVGIA+R8IEqSf6xorX/4w/C9MzMn6gbT9E0b
ys+95/pWSIoP0+rSURL+2vVixLDkecfarYFuu8E5avO5AKgjT0/NIP+xJBDl
0wpbwXsS61Vo/D6lAF7AnO/GTuWSip4mPnbwOFZwYUnPc24YNiA1DYcPLOzm
87Q62acZUuxOmyIE+ugpt7tc2giAl3gtoZV9TLtt45W7QtoawcI5Px45glP6
l6G91kuV7Hbl+3bR4kaIb3ftgkXFw4nmTdkgoHcT4FnxBUUfGJVd9cF4I3DM
SgKkab9Fy1PkAe0qHYPCaNwQTTx3ZCLBJCaZbgX87jUL08kchJ9RWsONEntS
BFOeEVIIHbpTaUVI18CFAbrKDrIFYubMHfb0PzHaJ4pBDCxsoEOfwJjm764G
AVTYhpEZy1l46N/CYK7AsvqZXf7SrHWvJwAD75kCcoQhP6XwgaHVYTa1YfJ8
/4zpXbxtRYNcm7x65BDZ3ve6+/rKhzYHtU86XqLOkf4g3pTv6VMwlRqz5rYc
OmXXyNjqZ+9GZguTqYQvu5iTFmIGBrY+WqcEkyWPhjRw9SmV/H8I2/cXVIUD
1HPKDchnfh622YejECJrWhQ+MBmTlkVhsn++EQZvmirvZIcubi0bFwU+3lzn
seLdlIRwMpXk3Lgm7Q9V7mA1VApEWGi+Nh6AjQrA5Dm6khaom0RSG47hJZPl
uJCM+WPna7+YDFGFD0rebQfjGXPrGQ+5eeHrcIiaczlDHwvTQ4NfAyK3G+hQ
Z1oZuBgJdY8ws1PKXYzummpj3k6v9YfRD71H86AM5J0eYSujzvW/rK+A6Xdo
LohtIFfAQyzVNDDVDfBWmtM4mmHa21TinZ1SdmL468yOb1QrX5ReHW3AYVrd
2h1mICuM2uz4rfsaruNAcgGxraS+vyu3KPZ4J5dA/6OLEKlqqK2xyJ36tPVA
TwPHBoQ6tH5vCLGq3dAkdSVU0dU5XZM14mUTQcUQje3QInGTHffpAnXzw3Ej
QGp1J/oJ2zc6XwgMGjaQHh1Pue7KOyzdDDSxxES+uzecJDoe2WInHZQh6wEB
+RPVg1C6yHmeKob9W+os/2rC+AdgHuwKGGu5tiFMwYSOuou7GiSvRl0AlFjN
j4GZi1Pt3lT50AQwBpcisTU+uHFLRz7iLQDBOvDNisexwZurlc/WRF34dcG5
Euv0jCSILLnIToNAWDZCro41TSj0+mHWd7dTEnJaCVXnlkNbIdSpgpMnINli
N/OPiFHWd7bghO9XPpfVCXhJsxt57/fPiA7hecKFRckiMN+RNTdUvuAvDf94
nLjRT06NE6fjjWGN/v7rxa0VVyiOo5mFhH76iYYUh8TK/Yg9PElHcvgjC0p9
NeM4GFdK++1PW2COG3lNPUTyyu1KSOGEEiK5F++wSPRFnGA+YvebTgIBApCa
ejlqiKTZAgFHnvtUnMuoE4TCMfCqymq8sQgaeKbXmp3SLQDV1SEufDljLP84
UWldeJlEAIGwuPSAvEEpK+Cg/fiY3wg+ADAwPPJ5O36f6oe8PT3Mu2oNnvCI
wzEyj7MbpMnXEk1SQfy0rCQHkX67QhnHYM+TkwDrhFz+/460L6wn+ZSukgBt
AUOHuvDXM/lNQWz1tjDcHVmUAelgltw05ST/6jYnt7pqedQuUha45VHzbfgH
4+KVPdQKwV2ZHs/05B76Nx3N8m7ngMoPX7YpQX5FjcmzbaSFS0t1WfZGwZMn
xM/Swe516XkSzl2rd4yglkjxwJi3we56RE/XBhxArEiieDRjyB6dr+SBy1vv
XHkyjl0h/V+13U7cUvmgydOSg+0N3yIipPI0rA57PgPfdSC/ULRO/NF/u+XO
e0/ruVuTJ69Gfkk6eUS06Ai586gLcbWhcQ48hj4NYFqr4ZuQE46d2W2MdGRr
AFiXEGdqY3bCD377CArfINsqJwYlfr2oT7fRwGOqPuY9POFrHuL1pZSyAMSz
hRNDSsFCdqGWZpatDG4qkLCv0RLZhCdOOLC5HTXxYPANBA9YVsqT5vRNVOmL
CdruBhxjoxxrexjCnkU9gsrQZYPQoPeMCRS5gS0M54/1TpCJMIhdp37qx1QO
Ss7bElFapG5cmtLEqhp1PSdTfRIEUdjw5odrMX6qepWTMxlpn2V6wS6U9Fyn
bg46cCMx7OteHxxTcTDB5OSiMBbXSco1uh2OTXf9Qk1mCGB9B6lfnp4rMrcP
RA9PxjZG1YtnEVaLNn2AlqdtX+LcvDR6Gl5nDVVXOFias5cRO4qIfN6OpR8/
Zwvhvqgf0xkGagK+PxEWrNJCQVjl/IxfYJda9sIbjB1h4jS8JFsIzJDVedC7
8cHRhixM27vuKM+VMO0FQrBqn8HyB00GM70gJr/iHsoSseDBGJ7xSweli2Ly
NfydMQXpAEW99DzHwx286MdiOggwSdR7JHKZmNiDPC1rd8jI641l6MIyuBa1
mkGkx9XeEJpiVmKgTgdDkfq1mtOrAKXmZijh2k56vxvGzClZDERXUPmNrq6z
ceXkOwNoyWftdb1hUMY4wa/ZtziM9fdfeQGOg2aBzUmsWKgWFDsBr3VElR8E
lzVKF7bOBxyvldhKWN7fwSOz9dIYQWTOD8Hce3kGunqKzaWQh6GqpeBIaMkl
xvl+1q76Ynt3rD5TGQoyM39Ku9qciO21jZXLpOn8EgRvOt4b6XBSn1duR200
oJf9ZjsDCzXQbWXz5M+kqbm5v5WOWoAmoLJjfmNTyp+DMAn7Ut/iqzE/svun
EPjaDRDAUdg/R/xNluis4erlMfid5mPiviHxQOtKZ20yocHyo5h0tZz86mdd
J1Q+TwlxSJvRHMEjA43eSc8FGgwDk336CqpsRsipqBQA1SL6BnTqKENDBxyC
3tRhSi0j61Dpn6UOK16R6wRFbCcltpZAdBNFEItK1JgBi10xsKtYRq103xE5
znKW6q1q0ExrLxcIAS3QZ0gDvWAFVWXoyiOQPA12Hb0zYndC2f5/0xZobIqG
BhxrcpbS4wfQ0ikuriLGgjAZBMjCHDVMoEz8dR26r6ECFzu6+J2XPj2WiVOy
HR2XVHR6KOjCCL7Mk3wgQ9cnhdOvct4UcP7sJIyK9BVgyHFZDAiHzV8Mo6Gd
wSGio5PgbN0PCoeO53cryLygZpoJfnhRBYB9hCzV6mZPDs+HvQ0QK9QRowZ9
01lXZiIp5Bkv+NSMenFIPrmxc2d0pn39aSv+EjqSABttAqmw4jTWIiQuZZox
ee2KwlNLjY2F7suVT8Zx8kdoa7utGuCTOGifx1epFZ+wGDmI1yXD04k6nbnu
Hqpa0Pt6IfHKojzwqOHOg+YGNIB1PtLzAkdSpYibccxD49x9SS0rnivhLvWb
z3dmiQFiYLgBUMr04M+x9iE+yAaR3NoaBy990kvvwiNLJTb3e5MFcFTIYtWH
JZV/FXRbP+0uhCKE8GaHgPbDapdB8f6gnfWno7bQkMHHrcd000gkTTWttC5R
aEJMXc4YBvRsJoedJMioPAvJf7tS6gcIMRa/mx17E6ZqyWx600ENk8bds4xs
apFwQMgqxZ6ycJeSUzKUn7isNMR4/iltq7XtITidkhdf1qi/kTBUa8xcSpfH
OpQUWrbGMGqdYKIQG9ISd/0fVzWT4shtlHr/8NMw/B0zJkRpQMBnEcNVOMO4
4csT3kVZLhyVtturVk9OzY118ixDmdUKshZe0qrISSWPsXokBtMB+V+Tzt/1
oGqcjC9QsnonkpMhje/4FAvSsqyHXt+2Fq7C07/oRQF1sK7EMCvh3gz1fbPh
I3pcW8ft4vgFx14VmCrs6sNynYbzxxu7mwiQDTqW1B46agemlvCjy1CEQOGG
txTmxbW7BHmXngt1t550JHUq4cD/StD7KmFnrfdYlW72uzem7+Wt78oUydGG
AdRPMpZJEMQdaTYT2JbhOWP0CRnrUVcIjDDXXI1n7Jr5hjMcVv9LGTzoXJVG
ohPQeDl5Lhea6qSO0VcSpZqDCrUMH4C0TiknnvPNddVrTnrggVybDPP4zdqf
4en39gxMRGf5HdPDhFyreZCQeeZG9ED4rn2xEZn8PDSoBXdKfxqh0FA9VVVH
EtARCaBLH5yDAY/QFS6MI7DxMul96u4g1ZoETaoGQyB6JTpje3TDbKLsPTGS
e7gj7Pl7eGm+TpocEcMrKisjtfjhiq7Fjx68E+uS7K89mMEQHhKKghz0zQ2D
dUSaysIYBQqI0DGTdmB2G8dZQVHcjwIoMQrShO6UEd2906y7eTZcteyFAZwy
gwMRnYahwBdleLCimeVqPovfoxxQOv22YCCZLDefuusM4BrT30ZxfnjOtd8N
dza0eX7VMLNokqtmJxwxxp6w8+ecFzTUQOjr2qRNuzot3VPigiyh39jzuX0J
M1pUcR6tb2WypbhGzFDSb5enD4K926NR9q0JS1/8MQYQdbzS1cfTVyh0hahu
CzN46ifVGjvFsL3XHBALfqvHQeD00DR+/4t5ZFpS/auGCPrknni/njHzgYuW
ak8xfFU1iNP3wxIgCNhyj7O8oGj3MTlgDfvg+QPAFYFBPYHL8XTfRbQArtyC
0yeVfKHmN6GL6cVH5zQ/oHB9O5Nb04n2jJ5CTWtzw7FZgUXZMkqqNGIA9hHG
icCICXgfH2pkqd3kaadlydONecbtvaPtuiUgn/Y7SSVfjQc64Hwb0YG6ztkP
bfN9HWL7ZVCrNBs6X23NCbPAfCAAbk1DPOmJAJXjqnDID4dxWIB1sZdoW67N
+lolhUEWfdpJNvWb4axOvx6o80NMvk0/1OpAHA6JZU8MrCE/undBWbF5j+fz
J1hJRTenIe/UDQZyddmwVLvQTasEGoTqRK2riKC9Tmv2EbR6eOk8/wCG0MN8
TffaQ3Z+JzBxItUDCSJQZRNL21c43s6Y2TNyRJrcy45fW7HJIPpjwdajWsD4
jDYB2r3WydXSlxpY8OQgAERISlWs/tzZ5UUPUWZjj8M1YBL6/m0GO0jSQ8En
XnmdHSTn/aFUUd/MghD8jpToFeQRkO4UffaA71+/He1WlS11ivsrA9Uaw9Gq
XYYtXetcgPg0JPZXySeli22QkndU/4ZkOimVAxLU6o2o7ShisVToNVvpDxNr
x+9w+aF4DFsVwoSSZ5YLnXmQpo+GJmG7BByh8zxNPgrehyciKoNe+ipi4BQ7
ccOX26cOQxEoYOGGEI7MKovkdnxIbgu1flGbhbvekIc/brwnu26vz3Wi6Z8G
Lxg15JvaOXEzzEg90JmyjGxm16t81mlUrEaiuox0qZBE0SdkwvxkZpYMS6Je
p0/4wikg9fFkQbiqF2Qin1UYBZep3dK/bUqIYO1LKsiLbI2V9GsJXu9KACe5
nLShD8gC6jLehWOSV2Nn+TBbEZ2WT36qLvxRUcEIy9+a55ft4pI4YRIb2czf
ATC+t4ozL2H/rJx+88SHk6LX/dXJZjSyme3oNotXSA/ZrBF1jHaD+4yCnDE4
DHD1BLtM1/RQBh0Wiuov0vhfbJnEHT2YFbnDnKCH+6R2zEKiJ0rU5mhxueXd
DcKHWPb0lvwTQmyc5hacGJFbo9HmXKkc9FvQUXwPiPb4zAsWmnhQaDSn2GDW
4jJV/FS3UqyX4/NBeY0kkjrHQPyoZbf8HeGeyTgUbFQ4K5B8ZAQrUWG//Qx2
rSx+PmeL+imISou0VjCr8yjCAC8zwZkkMEevc1KngXlgSoGpVK2ydWB0BYoc
22kF+8pnH3HWEo8qrRBc4Lkv9YrTnwtOozIQi6Jv59e6z7JRmT+SOFjHb7PA
gXfbWt2eXs4K9FP3Jg0aHyFSX/K8nIL2GqtEImnmSJBbZUs2UfvqCYTTfs0i
1n1TiS53xYJ9I2Ii3BllwM1u0R/KWtTX0LCrISNjvTLYR0lLGArKr0zlCH5X
21NAztoio9df6xFwWT0eDBCY/+hswUvIF+Kd6YL1Nl30Su5YPZDRiCIbxr0T
Aev9ruz3jxPWeltszjR1arf/rS7wGxIQAepjvpN9726ky2HndjjGmZwCNAad
mOLsk3grAlptUL4PEW49FUXbEBu4GHLLHnBb5FahJwpfYlGALTNMBgbvD/pQ
7pE2XbAumb7HOTP/fBloNZ4TgivYCGpRV5tfM8ednfhjDdsbvYYVZ5unOVk9
CqZ+yYSNNScMRIFihmZFagYcGS+mZYNlCXh5YGJwqLlg9sZFLxj9FiYHowEO
y3rWXWiCneOQxhwenGOxiHSdEayXEVoICeR3kPOtNLlsRkJD/W+TgSWpwVFP
JevicDEelzK5wpDndJ/2sPPmq77J7M9RFizKgj+ZAF96vuhynBMhtS/2oCQp
vD/e/7Spm6gVUThiu4q6hU9mnhJYKfw675Wjex2jMF/wLcg9HTzpYaBsZJE4
zfgv0urAqyDCf/Vc5nTqV34QcNYtq1VtK8d376pcLSM/vQabCwUJip/C1lgt
ADzsUS9RvUq9njr9epC3LZQNF6DhyjFb8w6YoeBOqVH5y6VMolIcylr58P0Q
gix1kqP3sPZnTuIAA1GDqU1Frnbzns28+KYVaJwI19efZ6auXLLeU4sCDKxU
Xc2M5RHXH7N8FeU4Nl0lJQqCTDeClZRXLk1BlQGc4BkUMxIno7Tz5XH78VDi
vnsfYwrfxPo774Kj8B+YdUIUgN6kMtQNkXX5SIo7zrr7WRACTvbczLd0Y85L
WskZhYHCUYQZDDg3OfJ+xBDlalOO/RE6lMBiqnKrzp2Q0aCw3AY7XMQEvKcA
HNsGQlYB0hzbA4+d9aXgWvmR61t4/jQCFsWuzuGNAeNAF87Lp7tdBtDaSzHe
c25vg5jfrnVw1yOW8QByoBA76MKRQqsepOMbY9VIjxfMfajT+oEXAvT0Fdfu
yhORK5aeUM4CRUP6vE0yk3nOTwz1DKy6QAG668NWOlO28YhAG4ui/5+jz2/1
B2LCJpibpz2XOPDTne1jNyVOHMDfuqjdGVeIq4GN6igkjZP09QsWgf8GKEs/
StWFYQENfz3+u5hyFE9MzMx9O8uBlKVrP3tuGijsN6yrwSeySdvy+SOgFmwE
g0HjKv0jC0Evyumfyx3UAgEWDpwDFKs42fhqJXFyJothBm6vJEphIuZCbOw+
gokpBSoiqc/oZ3dYH86GWVAmlO5Vn/wI0kKkP9/4gvHzravM1d15+ysDdZkN
Z64pvXgfNvZutsIx58NiwdicN1FDGHFwin9YoO31J+D7agzI+xd5pqc3UcVs
RM28rtcR5qV+V1Sp4iDQeyv8MIheEKRj6/GVHLuhGOkeFF7EariORtAR9u5B
iEdL5OTb63jpc9gm8EzZIW477P7HKTUKMPhiQK5VdC42GFzkbjcaPud0u5qL
ZKwz8iOAHKEqiRnMBSJjK0xRFyQnTCaGW5YmXA1JmTyI5FO3qaqx2QSWW717
IUDnuPLhO7G4I7/9F0uMUWuhlm2ArIVtezln/Q6ofuxbgp2X8jUDD8v6Q/en
fpu0IXqhawuFek2IxuquKvujviEwHvkweBxjz4XVF9cPvS06+J68rbOPOJ6/
kV8GP29tovs7KWJIfVt8lgamam4YvXE9EMRNgCAbt9tTF0c6IuY2Q3uTbZVl
0hg264tMvPpZXVzCD0EossLf2bV7IQA0Ia4aR7TJT3iDVJtjdDDKJW1AtCt3
x6KnhBveNOY9YAv5VBcFKL4O8jqYxQLlKn5YpsvLJJJgsa/Ki3HoTKUIOWNE
+G4fCBwWHfo78CzLrcVrL76cuOo2OKg0RGS17VEvrxf6B7eTzTiC59I2zjCE
1Por1b6u2GvMGR0kPMAzEOqetaVZ3gDNhFDBwQb+iqnsPJ2SkD7QzQcrPcKd
h6twX+1ANNarb64hZbHJ0GpvLTw41l1uyZpy3Vt0nTJzDBjjfHX2PDrhyHrh
7Gt/DyEOAMnJdjdCLYp1WViV9jWeFkN4GbvIx6pankAmxN9YzfqVCTKqlEsi
kaw/rj0PaQNMu/89d8RvnUHtjxkK6bMm+6Z7ArHiL3gnhkK6NjPEzllMKPOp
QfnGAgarRAFACD3rtWG+geVIIhaARM9S/5vfsD0cdX+D1pVOuvy+b9tZ/TiW
UvAveW7Vcmf7VXJPlfzUf17eeIlghGyL5MfqbonVgxB7HfM0TXqn0W3t2h3U
oaaBVbwvxMm986W6IexIxp+cWmy3YQ6MCXk4tGFrlHiLdN0zI5zRI4Ao7knO
I+Lnj4q2VXivqCcZ/yvUkbFMVhvYuz1S+bCgDn+6Xa0RvLZbSXkN9M+6bd2R
FlNd2Xd3plipPQhaiDD2FkiS0A0Me2vhAvbza5Bw3XaJhZT0NpjxEzksAgbL
ejv+1hl+3h331b4cfiSgIdkxUy8uG+rFuUbRz8uy5Td6nnA84gCKrzzW5s+U
BWrPzOmznw1IdfFdIRheFfwHETJPjyxcgKknfbv5V2ZUPfsu3kBSu/yoCB4d
ZBtxjtwcdLNrPCVBq211vbC+TbfYnEpw0BHCO4173gRHvurGSMN3V1aJIZTU
Mm5YEKhLJLeJWx2e7aapHNGxFtrwS7F0iaxogkjld4Uu/eraTJxjwECnzCEY
1pvFPfNVPMSQ2nBLqL0m/Rdpxii82wkBa/xZy8xJ0Y7OdyIY7Uk+9eYho6wf
xIAHDigRrpoRPQ0yQivKpthdUrb8LjbY3bC9Dd0dzEokQUGRHOmbyx3KjRWs
F/DmzQN0BJIcMdKqd6fmLLgheNmY66Ik9RWGoQWe8/u4m6nyUQC3hq3qf6OE
esdjTaGbTIPUDFm6QPulCxoan1nQfEL2wC2+F1XuoMjN/A4/IJgdwpwxksl0
+k2Okxa1o9Tniu2rqWFwk3hnmsqj84i1nrNdeIW0Hv+nU0i/wKh6FV519iad
cp3VFySjBqVT7ZA5onW1/vNWHBUeeXvd7+We7CtmiPLjEKGjEztPvlaZEsrX
/QNaRCK855FYmOrvncyRrRdQUb0JW2NG1GovK0zqG8Wu9jB8Xcu79HwqlOEw
eRl06htBfD9HDqxnlDIOhoiH+ntkhzHqafVTd6TW219KunVB4zHaXDnfBuuc
F61dFZL26iAytWCVhmuFg6hq6hyLlbqm/PfZQD/rQz+Buk9n1KCme5VCndfC
qGx4nvnfIlkkOC+srYy3+yWX0FKfxAP1QLU91x1RvDgwlEItBi7wNm8XBRvZ
wq0HmGU6irBl84aS20J83jXTpftSavA+bHp3liYg0bA7m87mZpT0zNfne9cs
VWs9cDIJ4tNzGSIXeMt2hwykdk4rOppFl1QHowO1MEunds3MUBm0KLji1W/f
rF7Ex6CwxFiha/+EIZy2gS6XiNcCXtbnf2ccWwtGsr4mTi+s6E3P5dsL6Yit
lLodROsNGfGHJABA05+cI4FkTms74YkpIgdTXk/kYmXIwu2tlYfMRKA7o9o8
UOb3zJHB9JvXvcWWEHBYW3sx2AU+f6W91UkxX8AgE4oY8+/QSmS4+VeMccmu
qpOtLIMueF4sfE+9Ys3FM0xQh9jtc59DIFidp3c9VVgy5gQ7hgFgnN5/2Kvu
OdLa7WLi1+cFn2T/OVR/Apd2f5uAFAM1RnseSI95AUbX4oRbsHtFrpReiyeb
WK1SBz2KnNvgvgtaS/StQBExw4kwnj8kmb9nN7LWvsw5DWlONsvPHpaubtHB
I3Zxna7mAUaw4nHh31PBmggsp6vcC8Xabzsbk1aAkLoROfXWvF0JrdXE+UbB
4dDRAkSBNEhToHl1+Vfv+Bd5F14h38rt9pFc/nLwejdb7gUupdSOEHBAPNII
q+6mQcTKVPjeNbFUriQLdG0h0QlqFQsfjdwVpiaZ7IYB9qD+l516ALkbzdxX
X5vxEqcfaGPoniydS7mj11uAsid8t3m+4rglUvnD9059F1BHo7QJ12ejMvOE
q8qqMsmuUemShuE7kg4YxJY1VvsPmCmgrEtZeB9IpCQ9oc2PWLrlUyEtuSX6
vAU65cAZu9ggQRty9CLyMmQvx02qVS21FsZwVyR7MNEFIFKchZRvn7XgDQrK
ELVqtFAi7REyCCzzMkPODUFh+YM3TCSsYnH/W03p8DAFdqzauMRhjE5H7g5z
usSbQAkuXfika1tyUh+fh3D0TSfpTHoLiurgQxE01QB7vmadVbPwhaffVA9Q
qkib03+XjuwDs4hGmGtpqnnqRuN9MHFc5RvOFyPtySRMBnrE/KTx7fC0MkEn
bU01UC/bdFUW3K5pAe/PjdFGY3t2GlQHck1JYGDMPh9Vio7K54d9B4MxFq1v
sk7Yg7gKhAhPbhUZx3un4KKyX/qTRvl8gtYzr6aCDqAMWiyfB0+UWJQPLlgC
wvXAh8X98Wb57m3DcLozzGoWcEsQQZjb5AhH0PFXGM/tKRLBfaSnMcSNeAoT
SgIhe+KTehJknLdbFcBixfuhOpU1pnxOnvMN9vaEVO8aNe6pZQRRdKuDCujK
d3dwqQ7eU/U4KwGC2gqQS31RirVkD0TKRERJsul3frZu9WOpb3iODvItWOXV
E7OQ8Q+FqUvDCU+KcI249GsYV7Ye7Lo25gmKgGrvgi9Ymf6N33RXJK+PkLRT
MRhhdNxjlBihLJ1HB6DAJwVbZ5/H7epZ5O3XQ23IYbZUhQaXCL8/Azdkq6PR
pRekg2Nh3Yrn0El9qw5bSKLpvyWMvjmj1suO1Hu4eTH0P1nAJecgjgbZR6QI
V2MUaYIPvfJ2SRFeybXbthLZL96yRUPH9oQyAPAbqUu6P6dBt8qvVDfYR6EB
j9J3VLP0CCWHg9oGAb2A2/WvHtdET10jElCV8N1pt/8Tnkj1Cyj6DlUdALxq
97nDG6If9ZWGP75Yjj4ymvob4Dqa6oBvg22z7PJ7wDLo7m3G/cY2sqT+H8ob
i2vRO72E5YBjvyPJMt6Tv0E0ymxiFB7O+EUvngk+cSmTWI2DPS9jq2sloB3M
T7uJNfsqhRxu7RD2pGednbukL8tUUVclrM6r/VsxJTVLWv4lS7qIUv5ei1JY
GDhY3/z8N1xXzbCuMPmdJbiXfmmcT2J7R2nJd9xwS4EF4/dDhA+iTKVNjK+x
Z2+CVw0fuf/dUh+qbDrS1Aul4fvpaEagHf/SOyYdNXl+bNR2Prz5Sg9jFLmB
Q49B2VMQUv/inL4D3+IrDxFOv+8gHEoRD8PdXOKD7AM1V5hxxEx0ELvwpvsL
71H79fWHr4WaCRAO4tU0PZ+OkmHKiFzGrpbxNpsEdUuNfMfKvqY+tqdtEB8h
xWvE/U9135mC9ufB8/pCJNL9UwAg7zCoLvBoM2fFMiSxbGv3bIT4Rb7Qav7O
hqxMzp5mTlfN4SW77m2XlkrBUMNsaPHsm0aAnLJwy0crhkN+UUehRpm68rIw
vhIUvvFxiOi04bIFnyF0eAJBUeCbQzSjZdHdPEvgaqKK/yzZ1DQT056pHriJ
pQwmg0jbSGwY+/XjQ6LstZtQ3RBqe92r3Higx5HRFpUsZHRa6KT9xoeamP0m
paY8Xo8GHo5idZ+ZO1yIefq1rEOP+XFBUnqcVENiW21s9jofG1hL944P/PMS
e3HN0gRpW6pZDQO6g6mbcNYlcaC8vmP+cGi805qExsOFXEhPpczQm+rA8/a6
/IPyeK3PN+9UMoRbk0CDM///vfGVqQlmscj+L0dt1EGo1fX/DXiGg5HbY27E
+jzsjQdrirgatMRGKTI34YZo1nhjecfJQsiGKoggB63IcfMT9tQLuSF4JQTM
lReHgaTEHkErsfHa7m4i0HhLLJrXn7cRJV4JYycqKX754IEKuXY8q0tnNbbt
+niYm5QfGE0uIEeueyGf4naS38CffL/Q+Gf7rWMFispp3mPZriJlry7pap95
otkHshQOyXt8Eb0SeHkoPXhKB0qKy8UoW9CoJitRJgwunLQzgjcgrLp2LLLX
gID9mXq01MIvYLqv+khLlMyI635eaHDarbOGBn0RlOMusZqpBs/1z5wvWFdX
HBiWhEk/ZoANoyzS+k6RJ6qmRpLWyzqT7/1dthemjukz/l+h1d50sqrfuXOh
wfKXY+fi4fgX5JFlBsTbxVJy2wsLUSEFNNKGHaTLHcJMYFzlBVrV1Ch8X6wo
4iMdY3T/kB6FEUBxjzg55L54sNYoCA8qq5vBg3XbJyJSW7pJq/JnX1Se52gc
3SqavYpYmVT5ChrdtAzWSwKhgBr2T3wxRWwqExoN+tiQjc8uLHY6dbqG3bBg
E0j8f+W+bqipxZB5Xuk9wwxcVaSBp19ihGlCLVav8pLYbzSRKtqNpv+ryZdh
zVCATkAnQIlAauIJyK3QKm/TVEHDLITi5mHM7HdhaHlephRN6QloCdLJIAb8
WLWhlWg3foB9jpx/a2GmoJrMptcxxFD8RJWAPbvbFwRHFwyeRPrnldZslzwJ
jSfwzQEU9afxb5lJERgp+YTUiRuOQXYJ2GvUgNFwA9o2PSi57zViuwWTn/w9
HmUv8r1ZVWL3kEz/cVeRUDRZI2xJfQfFfz0ogD3nTuvh14jw9zbEX/eOjWCx
klBnsGxv+/Lij6XviXNoqhMloOu049B/DAK8JAk0rhL5DYvXNIKgVdkOpYDO
IES106KpT6ecQxkoBRUIZqYbDDgU7QfjTjq5ebkx6LFJXoOPXsYeeBRQJu9L
oiyFQURTHpFBeNFFzioXpSsRSauuuYJLKUYvalJan5kElHy2IYVv+hG2B5Ky
qReAQPa1qP+5r9X/WXFpMdo4Zr1Q10uG20ognm5bPOscPOxL9k4m00b6emaF
Yl+JwBgQPKNkpqASEfZx+FECbgWazPY6YwNuFQZzSFb7n3oNm/53Fj9ANJWz
TNzIDXueWXgDzXlmTvqlomknbxXLBE0zG5LBT+dJHIH2bcX4mVD92dn2ausa
zlvRRu9kdWiocMl39MeEVJ4Cm7k7YqznrF8tdmRNfxn4o1xx+E3PZ6RkTFds
YIbd55m7H4JQDw03fsC1XouQgTFs8cMeSiXgq39TZpUfY/heOwbsKjwhjiht
qXuhg4OCXiH7+l61JPTMhYSdGsBtMuLERuzWFQ76o5ueg/wFPHqx14KViw7B
Ua+vRd0Dq0TE4kLyiPQ+hxDH5awazG6v0/pKTzcq7tFd1iPrekbhrTWLWhGX
/yXDGRr5RgJMV3jhjHP5gqwPjN5YqI+1ONB4ME4Lb777PatLuMoG+p5/vmbz
aPHslNBCGP2xImjifxxufxbe2Fq88UBpVou26ADesSdq0dEqCNyNM1pujFjP
oXvLMZR7DuWNvkJ5pYsr5phCsvwYf7xjwetGR2f84tmCUBWpKRTHMGiiMOgK
GSYK3O7Hfw7rKgFS+nNGthvvmMCKqQqIVhO8v7jBlzPVEnD+OYrsVQCf7ohW
HttJTicr90CpkbQsIbaodrpvMsQ+NRixj3bafBPjxZHj9EcQtX/SWMFRbjZq
MGLCYCU4nv2j7x9eFN3hAGBX3xl0Lv8h696oHDCXrv6uEffuzJ9Oq144fnro
v4Z9oqyqI/yIq8JJbtrOxqMUdnc0vN0Yoe8wqbC8SIMfG+kNIEDTPmgp1ANB
f6T5PazSJ1XwXMwsxv8pjO286QePdLgeEDJEHjMgcaM0zVNnLdR+r8jjorBZ
4J2BMW3zBFP8+q2qy37uMD7hCg+nnzIaNtLQfq9kr5c4w9st5I9y44AtRyBk
MOESFgJxUb4a8AuZx4/NfGE5O+9Mpkd0WmGBPAnQuCz5DnFsiyAu67IwgfzJ
ItXnNbTxh/ZGQ0Dfvd98sfVLp7jyff9IyegsS/3wcIKP6hn9ZnkDII10xbjL
P2X+h6iq73HC28g4yDCHNcYl3uQI7otiwF3gmHdnxFig5kwyfXCH14dF/ehx
C3ingZnedTiVZzL+72EZ6dABdI4pAz/C4Qs8j5gNkwLPYRBP5tdsqFahcw+P
WSo7ECdoaspXBbpwLRRWeOIyalqOljOVmRqImOiwN35oNr+tQ5Ait6r17YqA
zlIRA3TGa5Ts9DcX3afGNoW6owqGo3I2cghAzbCEe5IjZF73ic+T6BCKNNFH
EfF7EOBr48GrzWWYvsvJAo1I0q1t2JqM4Zpw3Tz5vBFa8qLWpuLSwg2ASdfT
/M+XTGsSeRSBVT/AUHTrcPeY6nhwCf+zSudc+YCAD4RapHcShJzG/TYHJoFi
yRcYIFpdLeVnD+MWQT2Ec+VgswF0BLJW3RG2F8IY2MpOZeQc+SfIRcOdqYqG
3Go7tS8NVpBXvCuYsATtzYAfxFo9h0HMtp5NiM55ZTfmsct86vGvEkQEaHXW
B0pj4L8DTfXYhGxaXccO0CSOB+qdcxJIJ9OLqCk3WjKYEfsOD0RTvwlSWrNd
a2LSLucNAef1m8ONaEFyT1TNciHckQ8BEhAwZfygCJOk/vTphFrJ004mkxfk
LOnEoS8WPTduCRrDnXyAAgapz7/4fJcoo0Jcx3283bDypASkYgzpDq2Eg6e4
y2RrM+5haG/3jvsP9XdEhCZyYGzKNq11j4AGxCTQWZ0L0NFAgbhXYc/5LaJS
AktVZY5AXki25L0OR+UtwTwkVdOYd3h9hl8RytpKUfcAxnrXyTMh6oG98FpM
ugxa85D1gQucBK4Rzg++Qx5lBf13nGG2OWzOGx/aLzCUpEF6vtH+9SdPaxmd
As6B0QoDC7lx1+LH3QkcIonpFPfroDbIn0yYVrTP2aEkw3afuJBe9M1cJQzg
JpQ8nIq84avrFbQLkezNke9h6vOClOJ17NmWoMg4xROfDmygwMVLUwiB9/yQ
xb0aE9p/lSmxCa4awzgC9HCwis/kV2G/dIaqQH/1relihwMHTg19y9QNflW/
r4UvbOe0SoODjHnD0n+GAfPuaK73tc5RygAoNG0LelpsywRs839473+dXhc3
OTAq5/Sr/qJgBO14JXNFwysoxr3i9SxgY3s8HgKI0w6qSIhr85hvFdDatJU/
mVVb8oqp/IHZxrLv2DDlMWH6qiAaVdVO2ZeqhhGteUIijQRIDsVj6JVcWE3C
D91rwi6PaP9IPc1uGIYS08Mc0TRBqCM3gaZPunkkDHINwxGU19Evc1v4ihBr
hQvGULBCOGIe8n3FmQEKswSLjBNPwImiNjshkX8oQQnQ7Qz+oXBA/DlQjCzC
IuWAZTz3FEgek7JBOFfqH3tv5UfNnleAtPC6ktrloyiZ/BS22ZvyBLfsLiIR
G+V700wOp0sm4tGg+jHSDb2l+btbhSppIUhOfTHtIOpOSVZIjSOIZGzhpQj0
pPArtb0tezf0T3wgLLeQOz1wZvodJzpu2sJj63dT8bwBPEf7RxHHyMFvFQYs
/ZXIvjT1h2SCfIQQoFjwkGh2bElfujZj4MX6/5OFgZvJwrPL50gZ0PBLIHiH
RYXN5hhZwdVy2YMTJcAXK0wFstkjJ0ak4vi4ZXrfAM+PUu4NReVhpRkwqytW
r+o6mo6VSUUKpMPR5tXr9IqBf3w0HGVVXViPvOwDWDNxjaAga1EDIwVn6dVV
vwmNfwF5bzndjF4b+doS8XjndDbeeL8o1aBUYHUt+XP0pLD/tx/LcaFGfUHW
wLCUbgXiAMuDuBdIQPl+liSAOM7sLRtFbt8LFaY1F3hHTgNKkrlAASjdI2O0
67MCykKDDdIbXZio1Y2mlWSs2S8PArP9IXhXxoECyeStv7qsWK8shWLSg6lH
QuU7MaVeFZQRdIpPw9iymtvEDeTcHtzS4Il44Kg/xMkj93Mtdiv9VHw6uJT7
EI4E26BZ36/er5PVbGB+DpMzJrpmmycJcRBTTuc8DogqB9HQxL/x1C6XduHU
b+P4+gDGgeoVHSkBqeMFttZyKhQCf4nBPhRYMAW3jTQWczLUeToc9yZtKiax
5zwrVnk1PgaIFUf4waeXGtfpHI4gU2SyoAdSCfqmFSc17JLJcevDtOP7Igtg
UJGtdpuwpLsOPqEVn4ANJsPXizO00Ywqo0IJS64wPK/FVggFB5Y02i8ukwDO
FCFpQc73Y1TUzSkePCLq0LGn57MHuvb7zajY9k8Ml9krw464dXQyC/X5AGt7
+b1AfC4dv1i1LNrwQfPHPiqaMRf+W2QZNLkoM8tXnWV9hPyLHxhmlzdQklUh
teZyV97du0EyUJx81eyQ+KwKAH5PMNAUDKL55iaq81l4XLfXEukIty/VXh21
sKV+JkFCTyqcwyjadQEAtN0PEpQ1/GRs2j8BfE2V4oCu41tdtkfyutlbvfyR
x5tw5nVCi90NS9ltKiGufJgCpFFmqwFGVDdSsmMzOXihGJMoKLEZV3dCiZAl
k4jJ/MAoxL490I0pCzpPn9Hso1ngKpBhXH18EDuj8OUIadjF3Gc86O61by23
evQIxRSRNkE2JLSusKYobQM3ameJqikMjFYEDg6futf7E8psqFqnqOxAQPje
crSjA0xXw9YDM4z9zuWiIPC7keSzG9OqfseWGIvGLZl72zEy4OejMzGCSa8h
4oEbclMrA8BiqUWtR1rMq2VrGa9HEojLxxxJY928wccXmGJz190zHCe0Ac3k
WT4kVbPPa+9NG6XtSags1lUPtnuk3OppxcfO5cTRrdtyouX7Snm+8GQsJepX
d4j/RlpevH3LiT/TIRPH4My1alrorAstL5hvDrSIResmo9dWR3c7ISmTwsTz
U+CHBr7yBe4blHf8EI0SZ/MNV8JFah/UjPmBZHlodT2rqiC0AzQqdGv7MIqt
Nl9W/d07SJT+nTDp/2xoX0nRK2AuxrJ0WkzwyO1bFxM8FBusgYmmmAiVNX2S
3o6PKmMbaFu4Vg5O8GjD/GiGBlXsVJOEptbASnwkU/0r3VVmwlGVVEdH3K0s
UGput73reA2eUeBBdjoYTDB1ffvfnHd1chepDCbLVP9n/zWZKw9apgpoAO3i
wh8VYTkqgTKsIN1+BSCu4STlQfHA+zdJIwn2IHtnLidY0JqnvAQJ5wc8CYy8
sjXYuw3EjMxByKXv2VHnheF51xRooeZnEsnbFQYSWr2zf/1MamJuHqcSy1Cn
rhY2ZNxgVg3D37MC9qrYxmPS03aWvgS1eTsaiVfh7lSAkPf48xj92nXpZGaX
EkYjZCsh8ZHKXb0zIiYiRR2yhh/3CYfvLzQs1969a9OLqY83pd/jnbP/dfdy
Y2z1G6ddthnUsJRBp7Qx6Cucrys0WX87k+VZjyAZvwRQcqAumx0VAqAmw/5Q
XzJ7ykPVvGTa6q8e9V6yjLsKuORLwkn1wpAycmEHpkcYNYtpZzIjPbX+NpqC
OgtT6jJRrHgxXZfX+AYzuldNc1Sbkoa4pTY8rfunLSsSog6QpH3AnT1JFjx7
NIJYihKsm2ryIMfBRYKYBoCyxec0lXMQdFEJmrzcv9mcbADpL/RzNT+Ci2Wa
+vrLQyjU1FdBmMcKc5TCzboB1lXl3xHyDKXYpfSmOKQSIhD3g8tYi3bVqYVO
0bv6ZWwTlwOUeEWV9vmMLC8nH1ie1M2Kyb6MqCXIUb/0tWAd8XeITzkxX9dV
vg9wxv/YGz+aqwpr4Np7SAbvQoX4zWHTfHTOiz5QHQp6I3R/FumEQg0VGMBJ
BMN+XvXT5cfMafrvbgwzDZn/ctwycJV9xC8rxX4C6hCbU7xdW+McaOvw/NRN
F0jKLY4KSw2KjVM0BSW1VYpY+vaZvlJgR1rDy4bzkTIVivBenYJnZJS2Xcw1
tIabENEnKiMwXK0JTjzIRquTSZjdQN9PDMHXm2wsCjS0WoQbb38fucObFzhe
RtbRbbWV6atJVTr0U4zGzhREh7Gx3SlgDa/1jpmr9VeaZzCOfDQLrOQezPRn
i6H+Qs2xsIQkLrcW6Q7McnFwDHO9zx5N9d1C0Y6H5tGMF1u0KHri85qk6Ben
NQFiR9btWwKYFn808bjOzixqNv6RmH+krfAbU7gfDswId61kVtDb7o4TW111
ttRiEVgI4VTJ+KhIg2+LX/1DW2af9lm+5dt/Y1fyviV9Sodju826hQ0S5h18
8NuZ3LqFcq+DpklnnupmdjT/ozN1LN6mfRA8N6zcGi5SQZYPVY5Puul4nQ71
C08lTEsjEiy9pE0+jGGlY45qtxI+eMTX170H1Og+rGWiGsuOOU3cPQTrUl+V
mMy6S8m9Era2ySMGSvAW81Wv0bjuG8qXvZyvOH/CICpF3L1+RlCHNgLXvbMm
JM3MyvO/AGDZw+oyYWma6ceTQmnc+cLvYw1cq/w/yVM3tql+S4rkEJUsAEt4
AyTRyfZ1qSIS9yn+om+BiBwdPJ83oqxY25DSI7ut/Jc5pw0FYRI1UhEopu89
w5H6DODbAzwtlxoRAdH070SApcVR8WvaxlWcFyo6zSXYEmpErRb22gzTp1KG
XTRjQfGniL+sdXYXjyP19aazRUYWGwbo1wmeAmX+uiwrj/S4h6JhJnuhTaZO
gv5X/eWeQKPsFqnyCvB6FZ/x5IE44BjuC+66rs3beN/X5qjzGhmi8eqaN+pX
y2S179xCtVssWuloSK6IKIHhNAc3iZyiSSSQGp2xcns7d4j4cLPiXZ3MLbJ3
492YjSLXYrtiSoog6bUJ2nsMlJO1UGyaP1yGBRU1sqncF1tT1T8oCChG9FXc
GFBMGDU3cxS2gnf1+aGOYQXzhZn3X/XgmLH5IRZ3Ges2kTEKhxMPmByaRWoe
q/QyUBVuMuY/OUa2tanuRgcNLbogjBvR3yVDKoix2ECEz63RQED0o5JhJ/D/
tgLK1S7fdv807dS7aWfNAdb5RId3ba+puHZZ/yUKfZyB3R5er5NzrPMh25Uf
SFztVEDJdhKjI/VZWovA63yu6GT5xX0Z9+SA3ZMqyCdB9RmZE7bldNUOFs73
yfOnumk385Xlkh8RMfxk/mT2Vfg3+ZtOvcMZ9gkIXt7xh7HCqVgHrlphi7cN
p+kfaGvyOxyfmopK6PHxtOPS1MwZaJGObsUZDwX556SvX6RN3yxoNf1aSYa7
UzcVIAmELxBQRSYqGU5HqALxjHs+ECyPxmysbvR85DlFBvxbIdATIAb2hOZm
72kKhfLmqnhiS/f55XuPgtdo9wr7+KBNth1OPTxKb44zK49DJg37WeHUgshx
2XyMFfsgKoK5SOkE1T4PspWgtVD0JLfw9zuoebk1Ef+pnjkpy2wsRKnGzeY+
RiIOmfDgxbO2azgKtkUCvKlvbbKyWgtVhKixClu5BwY/Dhdn5TJiw9HlgS22
bGAAs0hEzVk/cnD6GcMhrntDj+FD2iPI7d9r0xg+Gs+nawFz0TZXb//rsVfD
KbCWi+7t3FMsqM2rH22BBdTzKVtEDdipgLmk9t44PuagyezOof5O6KVTU3wR
63rXvKXjQrXU9wgotXascecVzxsdf+pXTaMSeEt9FvkR9+vzC1f+Qwmm/N8W
4MVM7bBSTERCisB7R2sQndWrQNQjsMhTTyj/XhPdjHpJU2A4va2lx71KqZ2T
ME5hIm5zSs1UOpkHxlYZxiStIE9qm2BSdvAu13qTsMShbqyobRN3FiWh6Vnp
GV9DBpDeCSDtI+k8peMnZ5jDO+c5KHu5eQVZ3P5ZT/Oe/Jh8wd5ogRTOxGgf
bP+jxQi8/oGwUdRMoqxYa9wurMLM0DjDUaNWKeycMmaTIgNAAFaQQqOx8z3w
x1uh/1vN2MxjXPy5jR4joTCutVs+Hm5e1DXYsqNzGEnPjtX1bFm/chksKBmP
S3QydoiK9qHuYsE6qMCYJrgV0ymg6MMWbOyu77k98ll4OZxeRNU4ZMnGuVKu
xLQfsjYMrh8K9SLihO3un73xt8MhHvwOho0IOgJSHUfVhC/40FXZDENA5cHz
jm7HVLNh1jm8TT6oK5JzLjWBGM/fE2jZ8zoAWgDT9/EuycMTg21YIlqHMfym
0fiWXLHwYzNokCxiwu7XcHx3rsvGkjYLAHTvxi1c5MkwnW5ZTn9qIAnzZKPT
2cVQKqS+ZGMWmlztGEsNe1bXFiJbgtio9gtIoYZKv3DuW55ZKGz3t6vjfu4a
hre6jB5C//U6KpjhBxIJOgUwvffNmVBaBYR/+Wt46Ddd8JPuJ2fBQOpbe9Jy
tpSHg9ejttPB5tt1CHOk8FXw1CAIXhYIhKfMXhxgLAvNcEyxkUt5AbiVDun0
vDWXDqpNHwOAbeWA8Nc4iJg38Ra1yq4z530HfV4DWXyYXvX/IwDTko/iWibc
dqeHfSrezQ9MQIDBfPqlY3LUClro+Rl2StnGB8Bp3XFP5uDLyj+hWQ4o4OUI
+KMjQkLibiCGV6GkCF7xeDlO9iIM6ms+wOhFkGtgHekvei46k9NhoIOzRNn7
pikS1BIKq8wVGUTTQattdLQLQ+DpgskSyXPSiF5QO8dngZNTAFoPpXx6Fm6n
VAgr+u6l+JPNc1V0n3A+ZDHB2Er+x49m0x+7a9VhpMgpggrem7+Wm+gkB3vO
5MLal1Tak24m/9hNLQsZbdVIf7FTgVUWKsePyT/hDQ8HT8vzvGm0qogeK3O5
ogxCsuUDNi+aUk0soj215SLiQh2j4PUBuT8yYn+/q8fgypHmwCEsiD4BWYSn
qfQbMEEZN2Tr2vtCROL7z4ST68G0tmYccpMpwgl6MkdE2JkjaX1OA9cnky60
wXEflSUHiSLMXqtANBzGkEaZ9Qe246o99PEPNDQ4z4WwZxZMyoBHrP3ZqYNG
3tV1q2wC4F4Aj8jG8UeU3iGBcPIPqKbs9HtbvDQjIZeGqkmxHNTV0+bvo+JR
kPwfrTq1agJdBvJAh4AHKAkmVxFqCFufTxWnXXxdYn9dP5IixcCdZ4Q2ubGP
2OOEprNQz/VLfV9/70teMMqx02l0whUMmGbi8lFi2Qf00NZWN1L2LTHcJchr
/2rzsp7cp45aEKYMSUx+5BA2uSjCusAwK5LdXA3bSouuyIwcS3ATnYIYSP7a
V1BbBedmoqKicAIXnV6BjA098bHHpsmG3UjQin97GbxNt9FupMzTTY9YxAaD
N/Xx3VsbcGBVtH5gbEZOr58xGHFlT1R+kQF9dtEGo5CZiOfjNFWpbY9XdSIN
qnffjfSy2uE38UkHNCZRqo5wV9/7xPQqdN3ChaqdeP4ic2xyCXvfYeBsq6oP
JWoJbDOj6dJijY7/877WoVCVOb9NPTXrUQu+7lctwiGIlY4zRO/ewG4f+DZ7
rtDQ2X+dhbX3NRct3TBIxlRLSvQCjfbtN5jzVK6LbBZXPnb5uIDKUsbNff95
7/Q888sU2Fnm2WZQtCvRfjEFdki4+6hhrcuBi6/obULAJKd6B6AehF//uxE9
SZ+KSf09Ultk4JZadtLrjuRaiimL19ZwTah8NoOF+i9m9y/ZqBR67n68DALi
NvfG5OTdnxqiOsnf47vma8kbm2Qs4VG7bHCEyGLSE68Zm6+D8DCZjcO0xlef
nPVn4yGcuvod6GL4vhSy4kPXKn1KebO7B4ulYjj8OnQgiv1Nc8atVsaqiET9
VyJPvy7183011Xtq/6u0Uj48IfFpZLtGldsTTN89lQphlAph1rBXJm4Llhu8
b+8jnbQNExohmpgYJnjEMRCSY0rqEsNJlOSOXpDSMKC84b69f3mFpRISLdWF
VV9ETpLQwIiHkc8nK03EHPMUsMlMV3YC9yTqpaEUOwg6JTzfe3Ri0HZe3QEZ
WNktMhWKX6hWKWq6ifJ9uep9CqVdu4DfN+hsJ/QECVJX3lLXGOGCC42h47+h
eXJjGrRyKO9qVOREQzcU3Hk+2RbplXBIbqau9BMUIawUWeccHPWx5xmRq0n6
x0JuVXokg67m4dtAOyRCeHUIZqCBXkD7IqQL6YFktarVi2FnKBBUusqcHw+Y
RHZyWq3GrWygTs+rB1BWP72QH76I7JzCR8sowqEjGhILqd8WPlwBYAHSUV3h
aRqZffJnRhPl342gwKaY9oEWV8MMKfWDXz/YUaqwu2hr43lWanfXkxHVMs78
ydIQgLxj5ifBdTIE8zfS6A8nL/YBZHKpgMwVBoaqo2Nq5Tjb7sN02mG/EVpV
tTTcaz6gHZOshiOHSPxu1e7U6pg74GC/HaoCSDBDmbBtNStHzv0ccEDmuSNB
JjSWxzTD34SA0m7fju/DYx3LstA1vvDX+ugY5wFsGqvwqZlYOL4/uIuJ+Ocs
5daWutFphpTu2FEq5wzQAsgulFB7z8sEUYjiSQGLq3gbo+0NHNZyVYqewsMP
9nk1kolctccqB9vtS68z5bFOK6a0fEUymLac/Nqrn3qZ5mM29MROQBaB5TW6
qNX7H6HAqm7nUcvkMIoCM757aPvBF9A+LIUOB55keQABlsXAagJBRr71XWxk
2+7tLdCfEzhE3EAjA2taNxTBIwUWx9d23ZoGe/XadMwVHRY21RWrSMG0SGXz
96W+VfDpOOQgxRyloFZMED+MlBqVanrJsZ/p1PUOPszPfKXzbp24Wn7H8SHG
3EyZOy+tiyacRzpVy9e+bzEXRwBmIehxcFBXM7rndKMQhCERrfbHehoJxIf2
PI1DK+Qbih+f4YrdHF1LUrcGXGh5WunZ4c0ca6yLjmqdzs2N8UX55AlxmEtW
4dbyVnsF6Rr4OxWF3l1lWpLVFdl6OkbWg/q4/Nfe+acjhGKUWVnz8a25Xud7
EACfSR/AMAXgCjEyEgYBQdP/unOeOWUkCZ4ve/RM4OvVfR6AtIaKNyrAy45m
6L2cJ1u/VEJhcZtVeQ5WzxNroA/806kv87fPasPmJcHcEOkgMhhXD+e1U2xC
LGEqof/Kk04AJtCbeTQi4rrGVdZkodG+s8DylA4z0qYi5k+Oc1+9vo6E55Dd
NTi5WhyE3CyM9jJMc3YXr5u0eSCJCzHeciyFhXv5+hoQk9gWMxtG/ArIPmAp
Md7r1huvyu35IW+UNY70v/U2RG9xFVB7xJxzaNNREDJpiUvlGIkYB2jF8vyu
i14zo8be8Qs9wCl3sLFNrebVypRTgHQdhy8S1WVYtYqI4+qRM1OF2hI4wpVU
Ftv4kfyhRqcu2K4IgMJHDTu3okTookHCHbdfcgdMyxJ+iTDZzQFk7sBAzlQX
j4YeiFjYV55dwEn6GhUZhMsBBbehIZPtbRTdeXbQMJrhtWYhu8Ud8LvOzBTq
MPGVqTykh4HHLytSoBeYUOsPTifFE2RQ3GcD4hHHrNGtUvvfRmbauTMSiEKF
+IllugurZl3oIV/ziFYFvXgcs9jdqPZRIJSl70qve9ANhuZRWj7bY87FFxcr
sUVcH+jUgXik6jIw2Gtobevly6SlaMeGY4VlDfFFtUBbjiYO+hgWNo21DvT0
e4Of6MJTAxTuho0oCm8TTf6YzjRxRbwZw/53Rii1i8hK303DT0qG9W7HAiCH
dUse3clTHq3xrON/V2J4bgmpNBbg+T/2781uursOMrCJSYy8dM4rdoOXxkMy
y9/dLpBSv1kOmue4lWkyBcSPQ7DApRjZpqzCVp85MZ1QziNcnRrGehJ0zHbd
kgPbRbCaYm2Z3/G6ApgQCJTS87lZJBW22Yf9cBlsDYU3UkxXEvaCekyA8mlB
tEVPFRz7k6bquU81fJp1N7Pf+AmeqBl303Iq2xj12LVT9wPryz6QYvDM2qOe
+0Kt6/MvGkdWj8OjwLvUMmbPvmpU/ofQzUDdJrdRfyXMPqKDCOMiPlnL7BEP
SvdL8tvpL50eICKTPKIHEuNtY9iBumGM2MG3iR/cB0J4sAKIxeblUSwVXPBm
CEsAzbwkV58VhiiR/71FSOlvSDNaVUenK5ylnp+CPnIKc9VPMKdU6lrK23S0
wkIhPVwOXj083MAnoLT96a7aAJk/Z2glj1YVpC+dMF5OBfUO0JlDIeDc2GME
99eexocUZJEqieAirOq7jYWo/h6HEQYX8GXAE9Y8NfJNA9fziQNtDDlQxEjA
9OIru6PDtKw+HFAdHEk4fHShoGZsA4fWTFlMW78pOyG+crbS8LDqyAKa7xTF
2lkK6JUNT+reOu82YV3uSpvD3RtnEUdXz5bt/MjcNGvv74+JlKOyO5pDSQJV
rtEHkh3wBqxGSOKiVDqZRjtxEjw6QN3ehlgBLCDhw4oLMY3IrABGm+YLCtFQ
K0DWrNwg0Jba5wV3el9du0FulA6HSOjYjV1pP5fYVooZYfyYMprjpuiQmSRF
+mOQriBrxjxa5lcIQYbBiGzUsBhxGVlaOvjxvzBqiLFfmzdBE1GXEJ4V2TXI
Fy2YSElI4IJdFy1BlAxRxEkbkAA8Z1MDA4TP/lgpE38kurRMWFHskL9DhIBy
XRvR8f4HDvMrThMGCGB9vBniHfndIdkUULaTQmznBQWKpe1O5wo0YZlADqkz
mFWmetPK7Gh4qY91JMUgFek4tM0SCSHycjMQgZ67qMU8kzpChJR0w3cOe3hS
uPIT+mChABVyv44H/rTcg1XLqO/k08MowrFfpwxQNIhayvSHx5p/ZJM5U07k
p0dy1KBNhF54Gv4c2kuZBi8kQFcJvx13GA6koTi75tfrTa+nyG/1L1HVI2tk
YY1r1rAW2m8qiaKH51XL7Sg3BtAjIYc7SmO3hTXqmiexkVf/uMh+J/jtOwG3
Js2U2x9Kt6/ymfhoV7rAG5+uhedgXjKc3X6REzOWYKYIHbHDtV/QQHhZLeyN
m6hZFdSEP8HtEC2tvNjwVAdal7wYfxhwrVvHmFi2ZQn9QvPC8PvbWyH7ChdW
0AIftrxmr/WBb9K2prtDMsGeNi6bvCSg0lcbuQ/T9k6tY/lwccNN2z1AfGPj
KDE1PqVYtgIdx8/2TklOAW5y7oKNZNbwiVHiXkKDO0bYfcJwFBp6KmQflaXQ
EvZwdt3d0zexuLtsFst20SQZUadggA6nFgJFw5mKRuC95Ao7J4TjSycbRsSF
O7uZRcynJYfula9Ip1io+FLXfvAIOxwgiUwDrPiM5oXuLHsdFU4RwylrvtIJ
d/ZJN2wREh0W+8ey+yzu/hv72EidD2VNeQr/X9aJ8W2/1bOTiRd0nLNtHPOK
HYioIsUd/dtADNHsE2ZIW+AUOx21JIgH4A9MAzHdhTrfTthvtYgTKwXAemRG
vm2fWfuBrBGMIZV9vhqg87A1+o62QvMGOWb6etd2HYQxVdZ1n9aUYROWkdaB
ivRwYilddRJwudXERtLK3q59MVVEDlZIy0siNss+bb1cLGs8+fAnO0ruxPiI
rpzWx/dsESVTh+lMChTXXFt0drNdPxPP1IGsS09ysNlnpmIO+F3IVvm76/4u
A7CWaxMslXQLp8xnhVsIo+e0ADvjNq9aZHixTzBzhUAxknvHS8UpoyJ1rcXG
yrgQA5p1VvBkh5wuzCr2IYRXG/bdB4f1wS1ym770JL5r4Iy1vCqkuWJ8O+VN
xftXlKybUSYJ3zGMaEiRmpMwuM8d33qG8vVP8evTrC08uuonfJbfe9i4YGV7
S0FjrW/dY+XlLSI1SXFtEUS3wziJq7Nnqzq4nJ564ThVi2mstFBfKymL7gDt
pPaN58REvmfetNWAvSEqgYh0C/J2eHol4bfUKR2e2FaBq3y/r1x+/zean+dr
FlyZ6DwO6Ywx4LXqAEQsgNZ6drmLFxCel5tu4yzQNbpsq2kzD8wQ4veEW223
2fq6+QB7Xz8O+C76XWg6VR32lbz4mVMTx7qB1sbqVHWw8bWXAtJNIdeEaCqL
UXmPVQ2UySG/zmyzZHosU2Nm13cRdJYbgOwwTnrRokUyLCfeG3xiEQ5nzami
GD5Yhmq0IrclWuEHsRAsxXwgSrnKbhSXUvHyoh+Mm7iM0jwfmREAdtBkQVxA
4MiMUrMBWlZ3jd95BcvOBijJVcMFYadsR2ZoENYcBoAqeG3rHPrw8e9oKIPb
oPc3mzgJHoZKKKPG71lej7bRfICySTaghKo+1RyKmNhAO8c6+/uiv7e0oAwB
gWjepq/D/Zyx7FRoJSa9ZlT5yu7Mz6TYn6O5QHbZRpGE/6tuLOFE2ZvwgUy4
rtOB+ta6ck4fIfixuCL5jjqTnASBby6oLkIiHmDd6nv81mo2J0TW6wXwo6/k
whV7SBAJWbxBG+zCb2IK6rEN7jMkKHIESq0VwaakW9rowLYW2k8cq1M2X3oM
eTtW8iyyL5zvahFYEauG34/cRoivvz+/zDa2XafV8W05KH7bHiiZ2Mmgj6iM
1cDX7hPyMCiEjFk8nBqkxO0F/C3D/Wl/WMLWHKdq/5iBqiPfwPE8KeSiuf4e
cd66NRcIHu+N37dkZ5hmwiVj2WRnuyRBad2Kjt84M8xlenkOyTZ42LCXeoTz
Vtoa4/XQppuTjQKWxLL9EHCxQve/6LV880oj5i+SqnZdtptNFcxCrNTHAbn/
2vortx9Jba9bQyS+kjeObkgM8LJWBoCZJzPqogxCsEcIYTZaA9yxrKaqoKR3
PnWR1ZvbgNfxfVJoeF4EFtM4UuZl2Ih1s61hyYd50X4wHq7VD1Q9NbVyYjM1
J1Tc1uRN/SC59hlhX6r/Q9PCX1ou01HFhMSwWoT6SjbmOqqFU63rdaW19s2h
tyuGN1DJbKkBJE65ERM8SXnSynQwd0l/qIelSJLp8Cnxo+AaJ0tIgVtvQaxr
QapxRDekYMkfiWO52YuKiMtCJFQMrdQcBvPCbsTOmquFnWjURfH8ac1k4gYf
Ns/PYb139kMW++NyT3Ou3/MnUc3yGDPxS/0aoZzwlOsoTG4upOG8di/xr0ig
lY7Ni/V5EHmbx9tkPH4ZiFVHEaHODcjvFvKPg4lF3n25Ulh6efXIQNclU7Wx
KUVE8k/f8sUX4YsO2CZCvXeVHdKw835Q6x4qNV3lxbGYrIxdKDmFHSIY8jKD
j4RpRhCO1ssWUxOrQDsCqTUs1gdYJ6UsiUeZyIkWPA5zFdcU7GW70XJSwUmc
EOr3SNOtYKxyg+X51lHvxdBmtLTpwErQPMjj/2iJfBhbCpCJXl+QhlKR4nOW
NrSSwV6ud6IynAC0hZ7ZLfx7Sll7bOBqeh/nCU4OGNf94RVIVpCcSfXkvCZB
xTSljjdjVE63kx8Vl5L0jIt5ohWjv78OyuQkxhcmpqme6bpsytU6XZozdlfi
21cunNIc2Reya3vkQVZF6TzkHmSwWwz33Kfgt58NtVQRTR5t0haWXdhrd7TO
19AiZkBN7/YODTFnaxrk7M9L7rVhQgNQxUcNXPB96pJ6xq77GnaM1P3tqFz8
I4WxG5Hfc91T3ps6+EorzNUsLiNIooOx2PtHbeEkVKh8OfWOuxNlXBeQkTrU
waFzfuXTMOo9HJ1j1bDnRzF233QhI3J9craWcTk84palsZ9AMwhsSWkqUUTs
4ooYP9xZ4qtnRVCBQqG17g3tFgh8vqviM/zC5za0CYcVl1x8XGUwW3wgyR2/
3RvFXP6vOBkxiBMtoGan81AdWdKxp4f6mOgp7nsWTZYT+T4ceuhrVUll1NLX
oyoAW5QHAE2ncckFexqZ8ioGmUXPFyAm42d8l2XukOSoTfvsQEQSjJBFkoTt
mPnxPsrx6gekDpIu460sLuYELsfms2/KtipMgAbCUSTBLn3zpk2SKFppYoTV
z8SAdN5E0VDdSPa6c+nURD1KMvBs5wE3204nqwGtRPsR50v4ykEvx2oFcNz9
ix3UYAMIJZyhtf6w5sABFzodkR7oqqia3z15Kvlj3VAK2+BDQ5Pfq+Gp0V+m
CfMED/PEpd/Z7BUlnp051RPHjbjWL3W2+hSvq/o2LyQ+E1zmIyjp3raoCPR0
USgGu9rrVKufzYs1u0hO0OzFpqgYypzvs5IK2AgvR/EJH8AuB09BXjaxhntN
gj7rVO/Y2K1dpSSxQwzf+JgprqoYPqlYHvtqjgDDcDvAQR6Oc9MCUui1fLD1
lHwODfgTzlbf0dUhl4cpMDQFMeZ2mTXfxGOFOrrahWUWi+u9iror8huOmWIC
jDjRXO0RlQYlspqqgEjATNkbv2zdiqj5LJnHnLAdcZfqFqR6W0ckcobGHJ82
9nHtvSVuME5TxZf2cH7wZZnjQ4yXnketXOJbHKyuxeYECE80y46llXoYXKB7
A+bxAE5MWXqiheM5wwbZk485K114gDPUmsZZ12Wcrsz7wUPPadieICARcmn7
i3mK11qklctEXUMyrH4QJtVbhw/IjAW9nxybbgwlgMFk4tOOQdcxUcD0lVfN
a9ujj4sa5bcROeWgNrWd5Sy7W/oI0j3lZGlRvjSUkqdReJchdtueHCtOIX9y
sHSE4cjrRWyVsPGhli0q1xd4t4WS44QZNF3DdPF2Xh/GeoNHQNrShmrENsiy
Z5zfO6qDQJYudreFHxd9QSMtH6lb9xODjibyhTI5RIzl5ro+YlWpmGI63r/E
EmAkXPEZ3boAhEzo9ykXkajp6mVJr/0WOUmGUhlKhOujuQBgn4366HygXXu6
7E7Pb/oL9ZJj1deX5b7cvYxyYLAghwd0P/y7Ve65ql1axU1vJekICPtF/xSD
CiD9mmmE5SkJx9kNTKOviuC5iy16/2+QiAsB1ANZDGA26DQIkQzWNEPJ2Ut/
V+5UCddsGxTlq89FWm+cgH13rDX1j7xwbdCQJpA4+c/+NL0MtchZJ8RYk02m
zTVMSq1CQOSqmaw/EgEWuyB4EPki3F2fC7dRPEy9PHmTflGnvdZTiS63XwBv
Ie8k/gsUjwME+3iohtmqH04sOCV+HyNh/ALfSLMXPOHYNvR2Q9Q5oE1rTsD2
woNv02zP4Ul/7EY7DjKw2i0ir96ikOCat94ouK/chX4BK+wnee4D90TwxkS+
/YwT6124aArGMufJ58Gx/MymD2aR/N+ytPaWdyOdkV/j/vsfYKlSJjiX3iwf
9K0mb7btrRpbqk/d4b4u113YB1mCuCWzbdHCpgcyFvRQmeBBfDeBMWgyuRSV
YncGCcxxokEuX0Fwa7+hMxdhy+xDH34RMWu9VaDModinm7TUKD4p6WPbI4Wf
c2VaU0QBDp9BQuEXPyBYnCuw2to4fI2b34B23LsubEnoxaXl7NH0zEGsRHYo
i8QoN/HBOGIBbgvv4KQQ9RTNydNMA0idXheggyzqfAUFxzY9qyGWfkpcAP38
RO7kjDUA8cp/p827EdOCzuz0misccOiLSxjzYX1Re3y+LlJzBVA6diaZQSHO
a1xXSEvFoLpjJy4PL8kXmaypGFrXv7qiQOvSTCrm0tdq3P84Qg3mrpnIA+zA
lBQRjg0MuiB8lKkNx1joD0ByRO1fPT/e6U4WmyTVA1h3JV0rSY4in8r6x8fx
OmwErKeXcEbpzO93g+NUWarKXyr/Wzjc7En5Qm7BitrKRABSUCEecxv0w72H
JVutEyej8FNOujEo24bdwsUUzLgQ0xEMEvk2uF1MR2atfyqHXtOPWOnoeqVT
Q/lWVRfOgs6+vzDLY3uLzCI+KJgTB9ksFrPePMGtdVqEJ8xG4IF5KWmg/1qy
J7WOitq04a/yACrrk7+Np4ii3NP5r9b26cZAz4YLsZ3jOOk8CJUbTzUGstFe
4plw/yqTVmzvcVLORVnvIJmWcvSABQC6sarWHeVxlNuIKwkf/OLyatEhIqJw
f09H81iKy2j8VcBp6W0uLGTb+Qb3JvKvRqkFyPZdTgeBeCAndHSjJiAYfZ9b
hQ8NywZyGU0fz/vtjRstzD+6kCsIG9ndQK85SCipyv4vjzIJy8JY7fSBZWFv
76+AtEZzPxWgWj7Ya8U0lBGHMBX9hJuUVou46ioL/7e4va1U9PwSiReAyXIV
GhuJiRqugKcAJtEtD+Whvwu1OynlIYrwMF8IncCc6akscNZvlgXyagbcQ0cD
6ZC02kJWXddsdBl/CocwlkEfmhuNIh6XECFSJMOvpzlUeB4JV/IDCsCgZmAR
n4+2sJf4/q4dZ4mQMoBhCdMHXMQwN9lMC6erMe97VmTK+eOjF7XQeN2C779G
g6+dHAHoHLxPUEBBTAkXgmWlrEoRD+pGiKexLuRTTOI1zBnlNK2/1xn36bWF
+yjjDxIuUCWx7yvyxY3kT0Inl8BHKiO7qFKANrZJ38oOaZXaXfLTMX6cUxnn
0dg03/+SzgYQoUy2zDv4keOZMEPBYiXqI1P5xDA6siZthzZrsQDutrsZATKd
m0frcfnvc7uMoOZZEHznUzIRqqnM85+hUSqBr3tKrfYR2V4358M/2p+sYPqV
T27WY8DRQbRhy5DqVWWEUdwvl7Kr4rzD7zDMBaqIoVRjnqgXXm7FqmBrNYHh
zLKnuNm7S1hi48yCWUz6qRiHWzp9DUk5lanfXgZw66pcUWJBzP/UD4YklMJN
Rvsoovze0T1JqiEpefa5W6ZgfoD5FvsLDzNefThh9hop0J9hfk26wwngCwpi
XbGA8Gd98kxrv9k9scSTTIlgXOhBGR2qDx2jo/2l0/KW8gSDLXUQ1z+qpzmO
lpYcPHIm6mMv6lJXSd2LokQsA7RnYEDsWx1XEljNeBF055HTyb3CEqLf/Hm7
fZiGqdu2xoLvZ6jyp9e1y5bHXS324o+OwpkOshh1k/CEDJFDDhprofr8VnNC
jXEvfbrj7p100qWUfGZSmLGMv12ajZ6q9i8p40u4sidR/zcm89XSrhdqXRPY
X/EjKEt5+EH1Fyhug+9Yx4xPTGKg+6AHy8OqtUYVCnnvqs+pQ6s7B8XkP+vS
poDUSjHm3XyRlZ+bhjxGsqYFxiItDjmh3V+3xwQa22lVNj405buFGdaOdwvY
Y+d/7g7HOK3ajv4vUBqjGyyuVWo0N7xUMeesDrCoQRFF7nHtk2/kZxGRtctq
NvKgSeRi74h2AW617q1ocn3hIuMrquj7unYYxA5v0A3O9/cMdcGlIVO34hAr
YzVCjdT/JANaJXJ9hmByoumPZH9mPFy7oQZxYAVgUbpVCFp/A2GF9Ukrxw1K
wBvntj4JuuVHO83dCjIuaQvas0cKSyf23cGTxA18Bq7H5S6wN0lEiDWxQIzv
vTDFp79ZKMsyjgga2bWBDlIRojqxiwDSQGo/T7FnhpmjJjHUjQ5NQGT3AwPd
ULow4D9Lfk2y2jPcNnlxHFrd0niASYcKP+WMPYS+I4wnjsA6faiC/fio/Ahz
XL75jcjgKptMW4XvvBed0Flw/+OvyNmj7Vt2c4Fraa7mievOszYrLy9q3ccU
ZxCTlu9wRMwCwVJ++Fuc7EQ5nIsFCyzzbG/qATKVj+rv1iOpPquV9s2fmtSO
EcUY/81smuWlfcz9Py69VhBhcss0WVAXuGWBQylUjMaWEp1cteVn6hldzYFa
R3x8KvrvzYGEMI4W+hfIvRCINNETioQQ5+v+J/FEcIIXfWOTRA3rvhiHzyGZ
EESYEC/HGHXVgZV/mkjMW41y9k8ttTyUNUHCQHc3kpm3vMYa7cR37RkaK5kt
T5R5RUi1QiUD7F6QO450kM4sE2AZOVTfHfulGqRy5VYQX/8dt5tzgGcYaLxs
wkWgGfAB6FLQ3B0WLzyQutUKQmurvCUxm6ocyOs3MUyHr+yg2M/4PjMubHqw
/cxLKXsJ0oVqLte3ZEK3e6ostx5a+tv+5AYlVl7/qHMfaH8tjsxRieWfBfPH
DgR3QBREMWCq8EMLlPKZiLAOHcpzsr+VX9fg2jv/Eo2wE0KLHh38cz4xbOOG
CURPgCsiYXwEQrMSLbsYwrvNzn9wjbo7aPCcwaj8SPYyG/328LT9zbQ7UIdl
ah8GDJPvoBobQkKyH9BJkbuSOh6m57bDBRvjBwOxUVtru/vXYOLUX3W97Xyd
OygTIau7pEOmgWhul6djKAgoPQ4IO1sIvPuckHkcMoI89IMWnBoYUQUhmW2p
IpsfKW6ZwxLRY5P1/LlGhu2j27ymyG1E9VeKPjQYntDJKhDcGDMzQx32oa4h
ApyBbkBVWEusgJDBch1Xnp/wuDi57f+FmjYZ4/68e19rQX6NY5YMSUq/e0Wh
OUxe2PvRzCI9nGnY+amoPiG/I3DEtb6/zuMVSJsaccqJUZ69ukr744TBfyWk
R4v32lIqDONYCa98CUDoVQjCMNcD0xka0q3pEAI1517+DLBbpoCcV+f2hRGw
GD2U7U+p39iAOH4i72OZF3FcZ1zodnRC87KSMMZEqs4/HlmlHgdwzYA4Qfxg
Nyt9/xF7Wa3F3wd/MwcJ3rnDksQhzGDrYp2KWSQpioC1D6OctrXrY92ENkfx
NFb078YYrcR8MFrBdW22d1DTcbt7YMOic6/GPo/KhOKSvxeH+KQEujkzrZrm
DeImVcxYlHtG59pzvCY5iujPQfYJlLUhaDeYRFxQWa8UJRUuTsj+YZebjlhR
EI7X4pk1+arIZqmqM3v/aAduCB4o+lLl1RUJqDv8czu3hFI4NkhgkmlFuiCy
wFdsLmbQcmTc+Voau4SZAwcCGTvXxjUoR6yfhVN8nIF9Ebe6/GDpAHYM/VVe
5rWvKso+njhHHwtUOo+gEArEP/ksTrT7aEAscnfBXERsQVNoML1aGMXwC6rB
tyk4d36SqHoOMiJsennongiaMwTsZHNpL0D1te8H4cShVoPcY8Th/qM+WQqS
rkIuapD3lfAoJcoj6vXe/MEb6o107VXUrJmDj50PLiEKYw5Qa2BdOvbsWc8B
iwWG2b1IGhWr9rm2VDuaD3mhC1vZZ3KibGLYxmvrENLYFUCwE+YKeJYfjMIQ
2trqKBNNZmqTe5RcP4pT6mfVWEe76jD31DR3iFKmnpIwhdsNYcMgh7Hv8fVq
yEndjmGpld84nZ61a73avAX/bhrVxhPyKhtgZmjS4l6ohBeAhtTi4yoaoZl4
J91IEBTA9peJ9LzRmLJj0q16B6AWv3h+9HUFqM5L02hxOi2g6dgg2B9wGXuL
XanKE0kOG0Lnd0wBVzbKPGGHzHVJ36DWaTriGWUpspiIHmnPqcAGN1hXW0Ak
bSxSo+FI0zxVfdHVn+2yqQPIQyQxQhGZczUOkPSOhnHaNWM5bmaoKtonVmIP
ddZ7IiyZbq7F0e9d1r/bkst86S/7pCwebSBwk/Kk/PiV7dLNHoqwojaOoZGf
xdKv2l7/09ku4ha2AXy+UQzKY7X8zniv7/HnZ8vrKgru+UEMnYNW4GlAUQav
v0wNKcWzNahPFDYRFFZVvb03nZ0vUY+QEJqRtkZQleT9g1HMBeGZVHPRiphs
+IsAXunmiYZHHsNATwlX/XQUMOKiTO01f+LzYgwVMtFXNMP9bc96WXYTv8VX
jVrDh9HKRAGCClxEk+o/V3EL9B9LG5Wq8fkt2MQmlVsItJomv/flTCj1jjbv
pVKiWrkMtywvir3Vv5+e/dX19DEytjHuypVfdB8EWdLk7svyJb3mR4GQ1qmR
nHvOtgMNNdG7V2Fvri4YI1f+GriWBCshWkOEaittymhF6P09369QFlbf+6B7
XiMxP+J62E2UaArmYnv8CaXDVP03XHd3yqZ+WLLkKXbqB2XM4l0c92ObgqNt
7C9NGKv5ScPzBNlI/OzFcNpLV7H+fSOWQh/EA3wfy9E4vXeAG2DRDypNKKFp
Z0IPve+RxRR5OXOOSV7fhH8l3IqYjYvZZbpkylULqoq74EUbqFUOIOFReF92
97E7nxFWDriKKsrUPDuL+2YcTbqZSF1Ov2mvKq0IExjkPBXu80XHR1RKFtJn
h8RFQB1+24Qkb8pGpoZBHcGobf9jb7+5u7yHmHadPvhODOBeoonxlmwzSiB1
0sFqzlefM7cazDtJW17w3s1K80bhgRAqUBYI9nH8L7sj6pkt9O9oWllsUyOV
IxRsa7igvTp5j+BrhXAsTs303SA8PkUtOznXBcqN8YcOPlNGzb1etlSnYNEy
OG6ziluSh3UnOk7MklHfACA8Z3YWbcUtL9lcRIA5sc6Rm0dFz7OyG3qdbjAz
w3Kurc9KSQjLx+JF+5a999qnpfyza9yZrjcec7tqmZNHzgvxHvl5E8JJcQDc
4A+nJj2Pco3lMIpOAaW42vM8b0DJnyYsfbpePmFznbm043Wth7dod/KCe5Ju
tt9MN9wHdkLOerfHcAffP6Fq+k5QKq5dpngGg/pSa4UTt/T+jWBn+VhZ0PIF
jVXu3sI2gufZo/vZzL5xUOHDQaoVoC58B9eBKtPh+M/AwMAfXD9hpBzLGjPI
Iw40EyHwYNLVsyInuW/Bwf/Lp1rMopj6SYjxcE6VBbEUCaQbGzIGobUOOm4X
/o+7JjFmk34aZHpMWg9Ch1S7ghZ+hjUPwZ6twAQMf7yWI08A/pdZPWN7gtQ7
2KVU8KM/o6XUXpXsB+aKB4kXszY9lXWCni+jXfPbuS9tkcvV6LxTpsjNOFNm
v0T9PoyTloUc9tuhJm+Dn08yekrkMPlejjTNQPxxC+yDshk2DUF9IJhkrfN3
vUeOmVQeVS4+kpY9EV9c9fz4szODY1CJF8o7NUt4GNB0oeSmcBpwUqnUH2gY
p55dOUidJVfmyIFdQqQnPtHl1iSnAEqQEkbLdbJS8hVRNGhoKGgK77CAHkWE
y7co+uDlaewjVuRES0l22o+HyqN4cZhaCy2QWoR7KxKIfeqM4HQueBRR5aLT
56qb7/CF65ItEw78j2lCv+lkE7qPTlwCJiRAwD7VC5yKUnPQPlU+/kPV1iDP
GDo49Xhfy7DmQ5qPGM8goxoIhSlXKKtLvp6BEQH0e1iwlhZBiyCF5weuSgtG
E04yuITHwogfhndQlJawo+4miYwuQVgKI/mHxr3ATVGCAthMJooh11I3SCgL
KnAVLJNZ8HQi/PZgUzQadJlkhrUbLxSX/wQHDj11jqqq8vZWRB775Pjs7Yqs
tQdlTm60u28mldX1J13EaAX3nNowD4+oRSGZ4tvZexiUQHh3mqw0IwMKTImi
fRHHYF8FsAdvKdWGrWIvazsDVLYrRtN6jg0MAoUZw098CMik+G9HguyBZBTL
bdHy95zfQVeAaXmnYj6L2977vtUnU70bYWnwfHdiSNGKnb9E49AkaZYiRbrX
HEa9ddj6YAb/O5xH/SSsVf50lKVYUXHgOZc5mEa4B67L4qPqFO4IkPhg7jzE
hBcRCC3yodwzRrDuB85aq/3Kdf57avVg+Obkr+ed5GiC9wuHVDA7yDpxTSR8
xE52NUHUzeXGQL+DDvUqWSIZwMHBrfAtHFA6FwHehyJL/t7ESGySvrsXa/oe
X4V7NbYcqW1MuaYhYoRFqZBq7c+WZ6HbYMxZXIADmn9qIewJTgZviAaJsnCQ
dmCgL9vYbF+4D1Xtb374zLFYMOITC0vGHIh+SFnsI/LYVjI8dNF2f7rCWG65
k3WQzgZDo8Z8RBZ78XsehMVwXdQbGVsxe1o5ghDw0caY1ompt8R91g7D62Nb
zFdpO2/r5qtmULDcDG+p0YRwxClXVcwy0jDCFxf/10BxdfUOwqWYJWI50Z3L
Z2NGCdnu/jvJOzjztAq9qybgWY6wsu7j5H46RBWlTNqZsHHRFi1duC4pQmg4
PquJffc2PYOf9W8D3N0v3nJcfUPWocPzbOSY+fy7Exm3eBD0tGQ8e5JOwgij
/qBaXhZ1vE13XCkLR47/2C6LwJlF0PabK4+WqWwHYjCJFUreHIGriuBxC0PP
D/nPERuQI+LMX6sx75MFvi4GulLXlZ6ucLJ7TmR1McMYnBSKe6i2xXBb8Jgn
vR2Ja1oPqGQ2Tmu3C0dgdMcXu7PFQGWXRChqzZfcQqFSyjTyua1iVZ0fhn7O
yDVYDL7ycQ7ct8SCImjTb94Hm+Gbjum0m6QPjBwMFYBPLG95/i6JU7qTR3KB
7T262gE9mly3uYI9u3fCNmSrPmgzANdT/XtIQuaKwAadtseJ48IfcOW18fCn
da1PnzcUn1L5sMd0itcM/q5ma8aXfRg5EETb+maKOLw+qnfre0Tmh//XmutI
zFT53Qhjc/KpIkW4MhOrkU0P7/lTL5SlT/myY6EqCFK4Di+NMVAMVcAr3KJd
iok0OR/ii7LGlou+7JYHGlZaZGO/wbopLgidL08dB0rl5Cc5wtjmycpkWXB6
AM3DdLSzq3CZACPo8b6hTAFtHJRB7TtF4qwlWd4fEgJmBFgbu+zs/IYKA3gE
FfcO3w7dJO6xF1w5o2L6U3ktOdf22TUHImpAo52/7wjAjxupDobv4XBZFq3m
DmAF1CA5211Wo1pXQCRdmjZSY2fTJ4Thskz222cER15FZ20NQzKGX7Kh+fsz
0i9qJa22Knuzc0MpSN5ZUNm0LXG/KTDvDE6Jg+fvR13vkxafXhBLa1m3+dxA
TJZU2X1ANMxyeqHmSGSuRwjG8hecJcmSNtkPBj4E7nviL5e1EzxBUz4dvtXP
6HG1O7hWAL76z361NG3u49vsbPgKFFcQDee0hc1dTV7eofMCV9DsrHlQVBed
dKWqxKSrtHiBVP9Av7X4Aan86iGL6PSioVLyF9dMlsxOmoHYkAZ3dG0F27mS
ZMcHLSlnuOY4esi3E0yd6jo8vgGz6cL5TLi8O1HqQOm646XgS6JNnP/71Ciz
LCDCYO8eLWXQOQOBlUmSwjGIMmj2ng340PKRztS0xD58l6FYy/qlIQOMW3Bt
7/MBYE1JhWb1EXBkjT3lydk8qHNaSXcjTiJPCBJf7IE2Oe+RSg3R4bEKBhgu
HHt28sGsasrbKnc/pU1xufjqG1WBe2QNODidt1i9mLc2sNcyEI2o2pe75sD5
CVOqvRDDw+vr2biCStcHj2NT+tBLkI6ifUtQ2dW4L2gj0MqJPSBrvjf2PS3L
wdLJ3/vNVlfxcWmpACsy3UzF2wcykulsJuDb4Ee2YtunLgbwDsZ1bng0hsfA
qttOq0vQR8W+0yX6qTUeOmx/NCeCQQhlVzxLthN+JfOmERyRJccNxXFGQhXT
WZ0n3pfwbslh4SMZ3OMCdnFn78kzOgDT0Mx0XeL0zZKwLT3FwGB4jqSlUYiz
BWAnuROazIHnlaqxfyRsqVgRzYrwwjIc0Rl3PUgb/6G0IefL6xRnwCZFT3x7
YFhjcQ+MgS/rrW0tcYSq9z3LzAdn3gA2Gh+V9sb79x1Qy3bO0WBbClfE3SPf
ABxZd/wsUPdk/pkxgvVidI9gczpIocYxMvqcz4YzAg0AFmD4Na3qN2LLWbTM
8wsiAYoXYwZINYZQgc7H7VQeoJKknz+ml5Ie7aiqh/zup2YohkWh6G0tD43m
zTHyvIXkaajVVG/HjatEmroIPaxcxwCLxRzrDVPOV+f1hUIV/1f/UW5W2J6M
fNdjU78DU032sD9oEa6AZINAsb9B7nt/jZ3o/m1ncoQNj7Zldj4qgl49e+tW
WkDsCIv1lRUbgd1Ium0UWRuzQBcmDA+Po7IFlgrUMDWH44HjM8toCEtr6Hs6
3BufsAL/JMOMIfIXEC9cxvnFOSoslvS+xAR6CbTMMBHjyhFU8S/CbGzlF8CH
3/riRDupbfEvSJrlmP0h+jsT3nHVigB8AQhASWahdp7LkwME6td3ZqHmkFjJ
rZaPVn6xxaK9N79jZRviJN+Fn42kKioQ2SCBwiR8cRK2qe4XiijiCBLcOFVp
FzA3auteXjHI4Zj0KWW8qz1YPTTvxSgTUj/4xfoP0RwG17Hni1qxIgmsm+O/
NYYyEJ8RC9lqfST87xcq5svX/DZZ0laU2LRoybp/Op8+1xGXXfVf76wVCCID
mdEAkGLKvLzzc2R/mMkKXJSeRhJsPvYElESuZ9nl7i+/zpnRz3m/qfq6Kady
jVv9ZepvhDVGZnZlKfk77Vq7QgHW3+JiRO1breVwNyj4tTquCnCawz9Ptqi1
rDSS8zdFml9/yk9+09da0sDynqlRFOzUFKrqMPnCaZ2WGjWRw4IZhwgNwgqb
1m0TnVz8Qpoh55m97cgfX4ckhK9FDGTYb50ibirAYZYz/6tr6ndelOddMq9S
MSWaxjh3wzwEJvSquxsMwdnrRJSyFteU/C4d5NegzYiT9DM4Uo+LGqe0FeZF
B7mOvizdKHKRnmeXmc6GXI1qWrAirh9/gHEkeQVFa02cu8nt2/mQLPxtZ/Ka
4ttTIxxoklDkLhNzImUcgsubX7BlsNaXjI5icNX1tIX2w8Y5oAdWQTAP5MoK
aRCLh0k/X3eaJ0cel6PHEPGGpfoJKlmRnK/jpHDbhaNQ9w4Reekb6rvHgmJk
MRcXyYY5Mcq5vVQbbcKCw/wzADuRzicSXWS+wNfMgk60yk5kls4WaCo1PVbr
GENhNJDo+fxX+Eiii6sZSEUoqOTK6as4U6a8CwryIyhgaVAMYCKP+iILHhew
rM4OasovCP71jyT7zzTLwrqbg/NZBZeUpasqTutfULL0f6vqah7JsFF2q9q9
OATW2jG9FsqyPY90aVuOZUAtSZk5Rq90Y9ftMmQpISVR2QyIhOu6PdCzBNa5
/Sw0v/ff5V3EGPdD+qBFtyf8yN/TYadjxifb3YeMjrRer75vTymPxFNa8aAV
gh7JS4oL1PIobRKJkx/eGLa8kirRHtl5wyEXjTVYEFQ5nHJs04fGg4JfNdSF
IfOMePjz+B538mfeJ36kDQa7LzVGNE6le1rGQS8UyZc7HonCqld+BZmU3QcI
UdtMEfpcnkZylyZlLw9LIUJwOIb0f6fWGEYE5+P52xq6VgN62w/pg7tT8jTa
38AHrff3tPgK/Lq6XW/yhXpQA86zAx3gKBY/j2+QMkee9voJLzdhrk4s73nB
dhO0ntALWHhZrMyCNB1A59N2Mgw7ywNdcw/kvJET53/uTtC3ePtKXkV6PjF6
iZ4cZpJRD64NprBttIx6Akp5a5jpNq1IeOpTjrNpWOPSGJrRgwQBDIcgxFyD
rjf25zYV5V8AlJLHOCsz4+TOFIrdQ6NvfVXeE7HWNfbPbwTHyJfl5aRlcaaK
AtctInykpUbUEH73mLURlrZF2fSh2s7aHAeq7filv8QzQDA/++P3p0VWLUNV
6rSt7q/SF28pjiDtAunuGaYuPuH6foD+61/Ya1OrYuqAdF2cO8EwH5aobOXl
iyUmObHlHG3RxMHC21PRU/TcuR+pPBoA5EmCt1awFFGlh+KkPJ/XsqinClLt
atioEOBFjczc95+CQt4u5pGeMqKWGBCl/h0lSqcmO1W8KWTKLu9ZYE7AJq4F
s+QGOvxyg2nbxplXIsrz/Ntct10JXvgmW593PxMIjqYhfQtBvqlATEXLGcC4
48W3jv03jlruNpAIlUtwMcE1CQwVUF0I6dqE4Ja+j42XvpXyIsFfgUYgBALE
arT1uLwcDwsUxw9DxUbHoQxYJZwLMs2rORO76dkyWYsLFb+y/Q4o02T+APSp
bAIIJqcoc9x6fIcssV9ZnnLBnYQuvcPco8hVZxm79D9ycHkWWHnjjT+fXGnG
wGeFqM6kUr8RwMEreyYmTWffpxG5c7g9YM5hCNY1W/nmdEh7Fm3okuTbh7c/
CTXegz+s4e/b636ZJ4QA1OVbNn2BiNz4+vYE+sni0lVyQYeVhgarjVhADnWn
iaEVeRFVBluPSw5It8rX0DRIeqnFSEF+VYP+BEDhL46pFv9nQQyCJpxmxNrd
WgA1tHIE3x/iv1RY6JofZsfhDFn2htIpsB0iIgvLZRahVSjLmPB4Cx4nC1HK
E97mMs35vWkVQYMo76IHVCdfIHO5Cyakx7R+U/0er/rfnwSk6jquGQXPRkLO
AAhkoFcGJLpFu3yiuYEKjzhTJny/Egch2AIZHH/nXpLQy0EYn5J3E2TxJVRX
gRoTGMGoV5r7dZyxkkG/+6KSgIAxJU/Vt0Wi8ZGTG0wJ2Gi4gn9ntfyjhQRA
m6rq6xjqDAjDdRTWEb4r2CEXQjyA/IO2UChFAHwDEjqqdcNKvcLjO5I25oG2
f2x2LWJssLDPIkp3hIRgNZEtfJ5ZqtHqVUyF2mWzrSN0yxqwxxrTXdyhqprB
Z2QjVRu5ZjJGvmVQ3RofkX1CxBV8p0FBdDa26/8ROWxglZcQigKTAFrqE1vf
PHuDh16pct2wpjdo+sk84X1HfHFVa28/r0zXiR+6qHZGdWHhjFJNQvCBrqww
/at1qQYagBa0PPe2ALBHDvOmwvcmCuvqq+YgHPGTeAc5fmaaZSioFLRsbqlj
IHRZ7oyXEwJEZYpRwXKv25lBz5H4HhcLfqnHSBZ49IWUX2GdoOARLAueZm+r
aQHmkq34UnuA/RiKDXy66/GeFluCmEzmSJQbbf0fLPwUl8A15Ou8JF8oSZFd
UIVkObHeTC6SB92fGQ5bTI8990V2Wd6y/oPCv9IoUKGUWYO4ZjQaVO0DuBBI
p6hm3YzZE++zbRzG+5uajELInPX2n4irLFVSV3xLOJvphD99u+z0RgtJTBoO
hiIQPmRztLDhQEuHjmnZql2yd+4SgoNc56G04CQk5Df+k1bKlj/qIWPxITf8
hnUbfWvCCAElIqEovjR6ZIzmcnunb/hVUE3ML5FQdmJ5K0fA7EyAchjBU43w
JQeMw4+52hBKXUyQIweTFmAUCAgcaubac12qqTHpzm3mo5ST21j92lsU4UHN
/YvXP9oNKR88P27ck+DdrIIZSxkfGGMvsazPd1meL0SbrcvTUVD6lI1njNtr
KgIu1wGrWsoQG4RY5+EYvfnCx38luWXppFthRbHikCOyFXMwGeAJbI3Yn80X
aypu3dAk0VcBzE5WeBT7CNiqvJjeb+e/BLVzG5r2AI47uoSUjleoLWYPJwbZ
Rb52AZHVSmUpOfx554IJ2I7/T+CkqW2Th4/PoQZ60JmX13jStomQucSvB93E
TJmJYT2w24Tzc5THwUwOo3AfR3z4prc7IOE3KsONzOJU+r5h1jgDFp2JI7T5
yVSLoL1tDLd9GBXDbyMyvKZQzaodTJBFpazjLVMsSYeZvBLB4sc/wRDT106K
vdQMik34wwBsz0hSioDR02NaNuWbTvbDGr1RYI1gjJ1ZyLpP/3T9hUsXypgy
lWkeVqiiRmvFDhFYD5tbDGdoiEz1yp03/Cc0K0W+VnCLKF9iwoXhAtJdqalo
xLdTPuQg5bQtPLE9B0cFtQq1l+vBMpOgKgS55QxnAPqzcbPXwBXTP73lo+MR
1V3x2ebn8YqqFMdO9Ev756/f2RCnJ1s1BreN5thL+SYOY7H9KDMfDpcGttDT
gIKPAtBupqiCPSjF8+LdXeAlqURi/xApsWIcpZGyaoe/tFR6bF2K1T4Kl4FU
bGWifz+wLXNllaeTwxWQS4s5/a4TnbgRypE9IQFAuP2mdYTq1sqPWIyi3g1h
k4cP3Q/C2nRdpfdQxR6PdV+WyFR8wQLNhHTOauZdvMipcUvWu7X2GD+2+gAr
v7SPDkoTo2TlN3HoVXuPR9WWfjHpjruKFnNTGVwb3FtXCOnwyA2r1vJzN5nh
F0sqer8+dnlc8mn41gMshtlCDaM7VbljellV/I/nEYHGq7+xmAA+OJIIBVVu
fi3JPmvoRxhUZLxEFkdy005JZQOu0IVy+GOQwJRGFoOqDES/KmN4juVJbAYU
zJbPkDNA5kuF1RmZqupO2vTIcT6mk4K7ojOcZVX7U6hQljNbOuMVbLksjhuw
aKZ/9r2L4C75Xl3rXStyZ4OsKVqhVfD/1gzcdgkAtcBSJsnLLXQc8RkCp0il
FEB1sux3zFYLlN5ivG6oI3ZCbZOhtiNGWEihP6/U93NP0l4LPbEw4vLwucul
D9ip/971vbESEI2NGJ5qyQFZ08fY9ePXHbeqpl9INZ5J9yKoZT80L62HWmcR
n7ByucwHy9pvUPiI1PFNJ2UeCTFaRt+CLsaQAVjALA2Xkp9gVtd08NSAhcr7
M9qBAaSppNGGssOveKOTxzpoMITyiTA9Pc336+EhLUcMGisiIOhbS7WO0hJt
IMHKAXn/OJs+qmlnUByfrknA3xB0qvhAwQnVrAz9S3Q4XlvVqOGoPvN22UE0
/szk8w8CLbTU61KwV3Jgv8v+FuBi7b59ImMvWRWD7QNQpsHLpk4WPGt+SbCm
BhagV88J0t8lYGmt8EIctbkMcsDqj6OmUINOmfIh8E0iWWABP1yO/IvOYH9g
fj617tTKRXvQcqKh870kBfq8Zn3GvZw4+7rEtzsAVvmhHY7l1GZxMZNC1hhI
BGlI4JBR+zkrIoGZgt5TkZW8etoHuf+BmpupO17Mi7umUNg9PMNYogVq1iHP
weEsW1KH/DbnkKAkIZSBPBEueFj0pwCuIJx6PtSdj848PrWWkpFRkI0gjORM
R1vUyorpK8i2R5MYliSlo7wwHgvD48172hye1fSGC0snkse7oBgs76zDzdDx
pfm86PyoplEZ0flCmHq9VaRWd5fkjBGAmnQZXj+6u1vADmJvX/nVkgaMy4+Z
Ixe8sW8L7XoudmJwVAuKMQLkKyn/PF2vmBkwJooMk7BsrBHpVz7UCNRzv231
7/T45bTpjsYkdYxuatw32Ox3xp0jh7kzTTS1MTME3rAB53dDKGxWKRwMpN3Y
RTGRbT8Fvc0FyMGuM7fnyOdNWj4zAdbLs0fW7B3H4Y+FnoMVYhtDf1kpnbaf
RAoRnvOEWliKnHOubzMorfPU8SzgNAZuGqsZhxbkpJKbPcBIKUWjm3uLajgX
LyyOh2EVQyom1umLWQsxL+cXjUrh9ova1yMmP3g0DjyDETlkOEZTLnHE3T3t
vJ/oL7WMKDqH8mKxs2zRwtx628bqSuGoiW/lIC7O+BCtcLBaFetBz/ZenG6g
ZpVkXIW2Pe9byUn8Tozqjqacn+uEo5wbl7IrIDXYtWpqtpAiEu5OT42YHvit
hx6axXT8FsIGt1eGhcm0zAdCNo4heclBbwoIiMc/hQ6aFWl/pFLCNEwYPTjO
blztUIcSUfaFoyers85sYqei2UeyrPaZpZ7f0SwGh8mnkCl9QBfmU75mAJbh
64aT4byRQLN9ox7jSqEm3xFeQKJOxgoICKZUeOx+kw7bkaqK4jMU5t2rFXMs
wOZ4WJQI6RthcsameKanRltCzN1ocG8yfZujUzjifh65Ma0C1+eKlj4K+Q6G
Avw++ScY9j96Xxng5WIJA5noV7bgTU0tWjDOhn2GNIoSFgkT7VWfhg1vr7Rr
ISEKnSh+eeWsY/B5j7xkU/tiKYPd/0WRqqFDQn5nygzs6eKEGqGkl2uQ0P2z
wrQ2PPTiz26xjnrdk7paGo9nivOHDsogw4IkMxPOBblBWf5hjaQDdtN3jC/c
baVVMRINtvtWvdHuVN15uNHF/MV1WC8e3xA3UyDy+pu40sE1BNykK8AyJD2S
VNUifC1jLrUtBskM7SicafVvSbdFhXXqkec4HS8yC1CUVQe4xaoAPxdxJLYU
AcroIY4MdfxjGNHrqL3Nk6hK9eOo/UIvqqGGUNyy9CTjHZ/OwvLSiTS+M8aT
LuKzis6KZT7rYRvwcCAt0gMtvbcnMOo0ughmlrmy0J2laIfNvQeI642u9HRV
7Rlg4h5i5Bk1/O52tPMfEFyNo6wRAkoWDVa786+8z/7EIwa29OrXcqivnoe1
/WKj8qd1vyUWtu+kLvPeLVySU/peDZEsw53vyTB6EXw0n1fuQqo54HfyrQ/7
JoQoIwlfEt+CZ7kh0Fi3nA3OwPAQTPLoEMh3KtsbQMOlE4/rpZTuGUm/G9CD
R/cfJvv6ifb7ocWAHULaeM4OBswOXSCTJQ8bCGbCmxshYE3Qj8CSNlLuNIuu
IG+l0KZxUHTcz6X4e7c6QOALoXbrIoulGrj5Uv1VoisPiO/RZydnaQLfEIfS
HdiYh3rvVWcOCq89see7BzHPaS5sAVdhpXd6Kg7OlD4jhFLFWlh/deAvUP6G
8YWodkXur+ncJoYg8qLgCjuEoAZUS3+k3CPd6L27VW79vu33eKWY23TRzpmq
021pelP9qs66rJjilnBb1Ru4qoVzHRvVY2Mdms+qGt/HwKxu8ZKVuEWnzC1V
dzthsaB42yXiJDT8PdGtzOrcBWPEUDzinEOm/IlMV45bxI3bV0sXFU9Ln9qx
mtlPmTKuqks552ypKWQQCx6rWS7yamuRdTOjGtbUkqIZ+Jo20fIg8A2Xb/Rt
TkJnqR3iKuiux/AIxeULAtHSktAqoAbpOC6DDXH1fFDIDu62590wHDY1OWws
nGCTba6Sp/Azn8a/2wQFZi2zxxeI0KcAH00uenSRYJWidIT5TJa218BFyncA
qxRzPRzMUEDe2hx+VfgLcwErY4Q+lsROAMj/gRf08/m62aoJ3Yi+7B0F+LTL
zfLKOB6u1m8F/hrwyBmZFs+1HZ9wUG0SoW/ombV6z/72qTOGws7fwWgQ9D8d
IVZvPRVIn7WuNfMccpFXhw7pbXJq9ARTdAn9xdxJYREWeg3MNLXVonQpNSya
yK25P8N5Pai4tedtyG/omR/YYWJprBY4kF2tSNLK/x5tqbiGrBXaZRU0UJ2f
IeQyKyn+fl6zGRbzg/RYwHRJwfl9hphCKVrcS6pwpexDceSKEJt/V6dyKs8S
z4Yot85NRoOn58MjB39b0rdL5rOP76Km2+pofFHAyh9N1KcvXUSNMJJd5yRK
j3e6AW3UoJ/tkt37SuAYq0HxVzPAy+vqZVo5j9WYM09ykQhR+S8TbOmSx05Y
2fwCEkxz8mHuFzcOPqTy9QSj6obvtT44nY0935YMcM/DiH8EG3XBW4nMzW9H
ObIfunykXQMdjlEObwcU1D2KcSIdIpcRT+udbYOEdO1IJ+32wG5DVgJ/t39P
MQMvtJXBFlJ3PuSKhpAcnN+EdjtC05oW9bPwlX4mg30/U5eZQpctjESshCuj
MFYPF4X0eLqOUN7T5UF/YKXnImRhex4sR8GDPRZAXo6OXmH21Zx8ftF3VeM/
XJoYN9dD1M283P/rP6M5BFjPpEoNzxWuVEiOEOLLAKDV7kp8LlTdPLsHBbmy
7EzgHIynNRxfdPXYhnSv0K5AnOlsTixku9P4RpkkoVATIsxz+aM3E54y5dor
uCaxe2uKnASlgkznu1wk03/DxJubnxomvxbBObDoSeaLAJELC0wuNQQ1fred
2/mMPRnq4TCs/i2FJcXEOy6HhXyOyUxhBeNAkEGnnS4NmNRCOC8YiZNUkW9a
eeWopM4PytY8E6JtpC6u9aVtR5VJ2cKiRA3iij1iehsD87/1TaWd5teym1Yj
fpCVGz50Z6+d56Hl3kL7YmMDBQkLNCVSz1fagtjAeL0MYZffVcig7FmFuNt1
uAci1WaF5RfJHu7zOkLnVyciQnEfb6B0G7IH8gRyZvV0NQkOYSUCQIYXnDYE
T9b73zufFIJ4UidLHdmwO4CMemC2ZQqRgRjaTRXxUiDXfrTqSaS+2TKBCnbL
6tF8cuW+LlAK3JPMZLvPPD3xKmD+8edX2mvJ1qi6eUgCT80hIhjfksj/m9nU
iVbgP2jazutA967VDlZh12mKf+WifKcwZBW9SP8P+snEFiAYtlzQfE+S6XMG
R1DlKQafD3e0+/KQpbXMKdx9KAyqmApBVqRUUuGhqsiSTR3eIwudNGUiqqYY
LMDwiG/+LmRvuP1dtuJP2OUDTapgfk9EbRkZ27kCs/NI3Cp+5FaKLDbrbj6t
xoSUNvR+ygirs65JTlOsktL3P5x+5hf4fxCSP4hGPmKjTiVnePqzQAY8c2U2
bjmdV71NFvGMtaF+8TxlkWvxrWy6Rkonm+CmJAApkTpzdyrsP/J9N58uwbBU
pF2vR0wRMeee5dUzqjJBBtWtVm9Xt8BsixIzf2agbxW74TU4dQIFBzzxW2yV
G/CJh2ZOKEVAkDuytJ1rXDf9yierDSe/ocKsxpSCJnzIlpr1uTMW6SrxKBNv
6m/fxFD13UXsLnMSFrpx2WVJieF7CTDVaKT8sFs4N477Xq5iqA0aC5Jp3BoT
YzlCDLtk8ZqBeMDUaAEqblJ1SsnudHs7MSbjor14aSN5RV/6guKZPfyxFcfe
K6Mq9uSdBVeCmHbvH+/BjEJIO2XviqKEf5n1OLOSkwiPu29sFaLT6wO7WI1I
zCvL+iIQT4BeuoEV+ItVm6cdSPR+qpu4KfalGmsMi3NXEexkqkbFRL4cPdUB
8WHg0dLy7X6ERJVo/lmDmg29nTKL2fHB1bL0763EntjEQYWOuLWGhA47ZNS1
HIXq6W3w2BmvRKbP8mWXBriwjcujnlIVxFHr4cT5uI3xcHt3QDf47RIfvad4
Z7R7TfgQN8cLO25r7IhD5byb/XXATpjPA9Ccdu1zjC+/teI8jUqlobXhpepZ
soeiETAyKNUQDlmh0e6lZQK1g7NTc+Z7/zapmQbR6ahhCy1ifQFZBWo0xTTy
3ITQsSpKJS84ykBbxCSZU7X8ES6pzyeSwYW8QlXM5EJIphKtOqeoMPwwIfm+
SNiwjcsCr15vfAOqzl1QioNbnvqYYXdIlhVym+iLlyP9PetOIYUKNkP6SWkM
m3u4B7S4EO+Ww54Hn3KihwI+jpFNPiFmSnWSkv5+REemQ0RrAZJyS6Z0rHaK
WNUgqu1xPvI1P4RNeDYrPpqKs5IK2Xz5sPROIlo/ecMGBRnXq+fWMujeznSf
+4wPq+GYmqsXGSEtm/rMoqvZGpYytacqitq+nptrwgSvySZsL3R2JY5UYMaH
2wyTu/b2vpvrUqZH3ze9PfohxrnhwK12jj2NIc1w9PdVHtIKwRb3BpzWDi+D
2Fd2u429KkdWk+XjSth26ZGHs/rLFhoKHegGvkUirc1gDUnUZPe8PAjpuKsJ
WfAie6GGiC/uYzmV1JRTGO20CMSexnj5ntr4e5Eq1pDksr+RnDfxMZZFP/Mc
qAYt2Rp1+5IVwOZH0xtZ2t/c2QeElC+hFuOMlgUWhA04wzHFwx1A+S95vwJL
4dTiUQ6Tdz2uSzGWrf/CZKwhtDXK9p7Gd1K8OewxejiFE9+6Wq3IRWlmu8yh
hFAbpmJAJmraO8h8cIRktmLjgle9/gryppIxEIVsf6kGEoAEhfmcwc2ubmg6
o2JHwzd7S4UrayFh2WT/nRRdZ5wRnXx5gOMsmkxKvIQYlYh/UYRznkXcU4Dl
bnxyUrvs6Ljlus1ZDf4UjJXQC4VC2v7NHq5P1P0FufBrJHAVFQuZ+V2c95F0
sl1L86O/iMgzmy/PI4txa+EZUF3MU17M+DjxTiedh4BQ6CBMe9a9WLnflwGO
UqKmVGTNuHqpjOTa5FwwqmSg5ZefhB7iGFhkD5ttf3nayTV/FIv6fca1wlUu
nBPUxvcv+OJ9Naf0Z/lXsPZMR7Ne2fpt4ei0f5d9BuQeaN+oYWjlUO6QERPj
YpzBrFuXwv1wA0YmF/US6wDgtD25wvjp5WCygySsY1uDKqWjMDG5GfdGXxsG
XTE/ls2/I2FUlMz1WVsaaJjsN94+i3dzZ8mDyh+c3C2NFCmmjgAZb7ScOtOG
ZQ39IQ6MG8ZiAHehEdTu47cRfyKqAtyyE+539NCIr1BxKNt5JnS+LoV36wRu
hvxdmeYWrTCHZSYK3Le99wPK3MQlDHZVt9k/xvU/ug1muitBz9y05spuKrz9
ZA7+h3bhHgaE6CcRtR5eL94Ab/WbVzMoO0K6dyyB2a9n+QmJ/aMbSiQlm3cF
+LjbZdrup45NbboeaMhAywXe6Y0rByrUUrNvlQhzAt0lfyZ8UkUyMpUno3oy
BXeXR7/CeqorB0hU6NjfBm1ytXDLQg8PpAdHGEvwGi0S3b77tk+/dLicvwMC
IEQBUjSB+fERETPOV+gr5XD1pzy62kh35bzrc0fSAi9/Q+mbuEhb43kmNHXT
35ibNllJsHb+dvDBgxMOj2Wc3BA35gvse15/s1aF0IbzACU5BAZZ9eVOuTMH
0XrElgIot/795eOABqQGWVFsyQYBdV+4JXbrHbpmVUp7jqUqXe9mrWJoTWYf
YBS37TrGZQ1PD61Jh6I2kQh4aPPyhsTca4W4ONrlr0KcuRV2PPO5PNEYQt6M
PyDPaU4IhIVX+mLw2v8C7XJlenFJbFBDQD18MyFbBypceQp+Z6cTQha6GCex
WJkqfHVODWpoYo0l3k7nRr9oUzwjIJW2DBsV6pGqryhxGbt/wobntJiO18g7
XwUVnB9W8u6QvslSvP/XPSSJ4cd2Neuzsv2AWJ4KO7fSMIFhZr4taPliMg0H
xT7Wos6JvL8voVPXxRV2ECa1H6TStH5G6idyjmtcrFDOOcFoKpESK6sFswp5
ybFR63/vz1bsWAqngROoEydXxkB8F5li+lUDwtAkf9VhfXd6dTpxoBFo5jDK
iXzJnlQwZm2gbWeEZ/ef9uH/nVNn69LU/KsczIn7PNYu8RV0CLh4Oa6vJ3Kg
Xr8GeLMgBlAETvyXXUkqsKMI3Av9tKQCS9AxPMXgCNiubQL8q8Ohc4znvLvz
Egv4InHduoRyNE1oeP34/IL7E0uNhC1IfU1ke3R2N3shZxqvKcHq22p9xY9g
uX8/4Lylhwdd2loF1Q+0d0raM46i37nesZ2yxbq2dlwx6rqzt0wdoCHOI/4r
2dvP1aURtCYzbdnQTQtyGLL0TMKmfVKCAkejMX2f15zKskpnzB34DKHxCZQ9
SynfM8mbgKfoLwMMSBMPNBb2L0GURTe5Vr7E5E0wGnZ1MDL4m5v0jOEV8lXf
KM4a14gpWTaeADZau3kU31TnyqFvC1mY37sn6hTnh/m57LJ95U96uiyq9yjr
ocrbsT9Q5lJAN/tyqj6fNND3USdlHj9+yuAQfur6JumKPejuSHWM0Xql0PVx
Fcz6ha6tkU6S6QgRxPVxMTBDTPL0rHvdya8H14n7o3JmHX0CbjrJeebfWPA+
YJIiu8kJ8eh/wRpEPMBQmunSyQGvluXVz3/unKuoF1nBtFYOO2lUVO3wH69l
tz+JMzUao8K8xnIwejAEnxUR0TXmwM5T2wyMoiJO2MNRpCCdQlgLVhP9v+9M
B9HzQxHhmX3jEAqHK0160o0XF0f04j6FSZDeIPn2La2EFcExkSB67YRZDpVf
XV84XeBNJXqfdXSu0mi1vIMADQ2/l631aZ0ILECePk9IbJNsSYC69LAGKSle
/Afqlah+ea2diUjTLII3GJhpo4D23HpaUSLfa3XNUpfbebPIndfpyhGFZKpx
+Quc12qKUNZW29C0hvhOn/l+FjojgfD2yKR0Ljoo6YdLA0bdSmpkZhR/wcIH
JoV+s5HmbfyhMS+/bmbkv7mwBtPUGfenJ2/ZHid1o/7bhpBTjLZY8vVjJKZw
f4fBfWJUCiKKgp+H0Gp6WFwwW7MeEdFUMxbaLZ73V7XcNvTC83tWb1xpo4Ep
wauOf0BZM5Y6LCvip+En3XZptSHBmX/62ST5aSU80UhXZdXbpJDnTFP/cyWM
Z9RrOFsatTZrnFHaFCi4CmC99U7Uq6ZyCBXZhx3la6vxAghfbD086Tnr8tse
+UAFEZD9Y/V3/Q4v7SBCalHmfYDkX8z+ZipSlXqZUSWf8o5LVOqWkwjdaUDg
bxHz80gh4qLcPcjP3QUE+MAfJHUnFtLgTghPR7t7Qb49PCcKZ/RvQJIdalNO
1v+wq5pMSAGFjPtz03C8wvygskK/t3qTvmWNTlIroAUsdSMgbLKknA/Lg/qa
WKw2bdspnF11QVFgFVagb/GxHT4NRFqUMIDIfD0vXsdAhIjLD4S8GD5sNpqk
DvW4BQfOWp/KurAojuT1ShzD3tU+aHj6jkRBANHEkZXG2VjWrPByAIjFPdo7
yrdigzuTgottq5jzlw8whN6zfYD4VzikXHiU+Az6WRFnnM9lAmjNGRj2rTqt
1UzYL39Jq/885K/cnsP0teSBuVS/X4NnaHYEME77EprYhcsJbHH0wVvz+hyV
oiMlbIi0ZccF32+sI+R7io1KB29KkC2g69ppCamp+ks7RXqHLj3OXieW+1T9
DrnBwf+xdUbmh9I1whxkS6kRh+MPatR6R9q22SNYb8xXN8FgJS+aTPBs9oOY
HvYvf9rfPk5LgXsCMCM7yRHjM6i6lczBDmbepFmNp+JB5wDZYgVzEdsHSY4C
+3gl1VMYZ/7ax7FiX4tRAhYkC46lDPMlQ6UmhpLbLU2QFzcCGygzlIlBUtw3
Ir+SH/eqDUt5DF0w39O33V8lIEZXhM8PxoLcTsahIQJPlesmGP8SdYvI9+mQ
rr99f58gLy0puLHsZIi0PREnJN0b7YuA4dXgIOdHTRf+26ZCJ2Cz94RDoQRo
jurQpbvpzUaC1osgdNN31XKrpV61sT6iJQPFpbC5MlGKKJmTEHXnx+ozw669
HKusNm1jAwp+WEn5OBTMizU0/XdN7X3S3qUIHdFdaXzgDiogXtO6s1yC8/4X
hp5acaZ5xB4GYZGUKBM3FvEz5ti9Gb3JTgnvSKh2krZIObLB+3E9a/+auFo0
GD0928lCHfJ2hiYEY1j1Q/a9EN4KT8xRzbYWkyXCtijeQM5ynsKM+o4ur42c
wlRIPULIAFZLSn6tITrXuTOParL7sXLyeZbxFcMZmv/3iwIsGQQ9DfFSrJpa
m+wY6PWQ5QN6/wa0inuIGb33pzdiizQTLqVKZMs3J0mLs76DTlf2dXzxt9eb
iG+1vgr2yfya/rPL6o1R+jzmPx7wWBaenb2HIEMYnk5PIw0chAl4zJG1THFt
Uum1AYw1hIkw93+ybe86mKDw3lbU94+PqfYKHezN40HLYfDcQelmyjrEn6z6
74zS/UG9EQidTSvCZIVvCCqEQ8e+7Sk1oo3ghzDrPjWFc4sFcNm6cyCmTwex
cGrwi+3ImHAXUSEWDCaikrZKS04YYFo+oXI2uKLkMIbaQkyIGROCC9eKTLnA
na6CS3Vvt1PLy5UCovxs5eMjBoBfWvi/llGyS9l1HoLJzg/3jDUxwQfNS9GK
Gmmz9Mp20Pjah2deX949j4EmqE+URxtoNGBwP9LnMKPueZtM9CgQZfXlVtE/
cvPG+Kx2LuRAZFT9Vr2sKp/CBMeRKaNlJbAimCI0naPzYfQxR0rxj5VFQ5hE
EItDbJEbSw4CjUUuJxrW89s7x1x8YnC3qPN7eQLCqxeLHDk3LSukxoSM/Gtk
QHN/uwwgmwLpqdmbYdltQKNtYWTiQ/+uEUFv2KXoaw+4RTD/F5yUXohI9aa5
GyeEk3+Yx8KwpORHiC5lerhn6RvzPf8ctZnXi2VX3EyeAtJ+i56aBxIyP17+
OMqaKD/7nZahkejeZtvwxgVgwHizLfYARe74NAzLWCQ/iCGGf8tg9ycSTbm8
/QDR968aTjTPe4pLI1b9fiarZkb0F0pckoHAnY3zZMHTiFNO35UjP8DMbg9V
dI/DTzJGlXvZk66kZd6w43a0yHTsZ+HP2A0ssn2Jr4nGR2hVDY97VUBScVyE
y6ksnTpBfDcrATQVR6N7p0d0UBxRBzDXJ3j5GVFmX7pQo0Mqx5O0Ay8oKyBG
fqtEQklBPc17dmiEcIg0KGTLTyVXm92DPSbxagqg1ixYd7/isiEaTUS5fx8e
MSnPWTsJiatXX4R8h+UNW299QdPLisNd97vJqUbIHIM4MUH+RPZOh2BnmeQh
IMCJ/hAsJrYWZ/deOWYS9Qk3nCRRpR5kmBnLMNhUKVLWdPkHzP5DlM59mcFq
KtlfCmvJJkzoyKJfv7WEnPK4YbRoAz7mfjl+ZDbricGm4dXbiOz3+8QIumx7
xJX5sZSHT1MSDM/kbU8B7cKkFIhjcLQP6e+/uqfYGl0eZ7qJRFllHL2YI6gB
UjM9e9vXGzn6Is2IY0fMevHhcGGYsJOWuVdNRzuwTg6c+LwBX2j5U0lM5dDp
k/Z6Rap+DrqQvBx6ffCvOeyDKV37Z3VYmITtswDVyWg3F08UPntTZn5ivIM6
icSYBJPD5FT/IcsI4+OIFJzaAp56363wadooR9GWau52ydQcSnYvSNvvo8qw
rBZMhCDDq6FtJF8yXgepi7D6DdDPTOItRThMwX1F42kEvnlR3dLIMGlT585S
sOTYsbwOPy24bUM5p722Yo6Uz+4qA0Ko/gpkhH9es1nS3QOQbgsbn+Lhw9RG
XaWo/Mg6VBr62LW+Z5J50rLhgjSxKvZ3DRy2ih17Zaioenm6EWcuG1Z+6H2c
QDR/i3VzZeytkPoI7P5ZyNVvMajcrhMVip9KgxqFD2Y+zm7pj/edLHFn8RtD
UTBRaY5tO2GUDZOtxH8rSuETDWhDIutac88cMHTDL59BhsxVDLqxEMhEkfr3
fEofwVcH0PyKUOAPGuAUPTw3jFJkOT3EkRHycp2W+I4I1pPdP/5hAjmvls52
TEBB96yl+Mf3Xa5JEfPckIjdJlAhrGeNu2lMkzRzm8ET2TsM2WE9ymYci54T
8F40n1BiVTzxYn1FE6MqBDlYqX6b5E+pprYcWTTIHFC0/6p67v7WQ5pC4TG5
Z2sbmupJenUmHlBpkPapAyIQDwy29ABrU6LnSPEK/hJRy+W9UKI7zwPIX7WE
gAJjbPGj/IEM+7HjVj8VabCbCO0SOcNoo0hxX6KJy5EaPKgSosN2YHwHKfGe
Nm6FASPbBNNw4n5hPHqqNcbABCnXTGUfCkqeTo+bC24ckD7vyF8tXr48IX8p
k1xCDZgf9mkP7a8E+Q0lvNCAcJXVcdDqIt+NqOTNaoxN4XEPFxrA8Y64FAVL
NkmUG6uJeWi756mEuYKsgir1BdKVJxnhw3nUrN/xt4sLKPhBCKjE6B+t9CPv
0ENaVLnsm3cv8E0G0IAJywItcKSShH/S6ZmK4dXlVeG/84dx3cFoJuJk7+yM
tUgWV6O7xiDz5FfBy4BxdwU8tTJmrPcYSOWrwWbAKCUdJ4Il4dwHdGMSSMoS
yWPXBWqk1LmPrySIq7ykdlh6gp9V4VYFVeXxknneQIBZCG36jAGbXDq1+fe/
dN7sl2lmV5lXlfJ3glJl/P7gNKSlt9MyqS07Jcif7Qf8mXunVgMInLeVN5q/
xXVSmk7qCw1rZU9xgBW365cD/Zw1xZQ5yamU7/pBesulqDww9qG+4ZbPWK1d
a8MdzfpGCL04FKGXkvfCmVRr/KGoSAjFDlJRqHgFhAiIvClG8NxbyFKR2f8E
gB6CnLG03JKkwDmcxU0gRuFM2jCl/5Yyfu/jKvEXTCjESMqd5kH/RitptuDn
odZK1mctLYqiOyyLw+Unkt7CxKJtPvboV4/eKOlRhTU4bq2UNssPnCzt/kwB
4Al+svPROqZ6ReOkSRe/j2yccnAG7+RPre4043FnBEhcxRwo0mOwx/R+aW1A
65YBKzCbVfKIAJEa9I2HPnaCGnXfdvoKq0bJuDj0fR6cqjB4qfCWae6aHcCD
MKThhUmb6aSvvdFVVpTsp0bAqNrYn5DFCNpNtH/51TAJmSAz+8ZVGI8sgogm
ChOi7fLJuMb3z/r3H6t5uvZUqjMHilKrkLnIJS98urZwFk4UDEWstihr5qIa
GCNxoE4mIC3I3CpMtSZRwfjfB95W+/m252XbU1yVvhPjgOipK9+G3yIscktj
p6GDtuhE4BXtGGf7tZj4DeHPTQ7yjv7UmKIqsoZ+2QJkq7TeXcIspEoZJLVn
OPqMWQJlDg/Y3N/dFAs5vZiC+7bhunp7cGFBpVngwLa5zboDR1QBSMKvFMHo
47lIShd15w919vPZ6xkEcEYdYuW+Qk5c6EuRX8jiK3+UL1I0BtH8EGYA6R1w
vVg4eIf3QMBhuEFIxDGcYb/fRT6GKgjdLpS5O9JgvvsmKmPuK9YJuG9PH0Zg
EV+PEsghdzXaOyaQ9vXBWv8OisMb50+S5272f1UWkPeODtudDMF7UeCSgaIo
8z6lLjfG3v32pxDtIUAEJWbURyPa3cCZhLG+5pP3cMtEEcBLzXyFSqma/fzg
Ol58HobQlwOGENh8PNbrwG044wtp+3bcMbkYtKoZcRchW+yF7Jn2nw8wF58q
fN0LbRW9lqdb2r7mRWB1LRS75O/qSLI0JLwqaf2Ubgv7Bl7uLx9HWwx/b6SN
a4quD+nCZ9g3vKU7o/MudTnJYqGe7UVXANYAvI1Fv2P8kEsb0RPcynPC0EWQ
1EyzsP1FOxh9j1rdwNYGEnA+yd6xz8eBmoZfoqpHCFST/9wxNO8OglocKHJJ
49KTsJcaRbpR52htXyWHdsDgAiKLltuiLK/Rewhk+xFzDYayXOrfiKm0lE2d
Gkn5fDeyWaJSuRXHUG4/B2r+gBqWmtbJBiytiW6gYpBhChV7QqK8bTBMmkzt
tT7Jzk4Av1quk6ymRHcXyTCbVQuVspN7vI1TR5Z8UYirlsjNyfvTdNhxtbJD
9udKlLD7wr9k5vYZW532HetAYqldQjBLR8hzpQL+6sR6HVtugVwswKck3tF/
2qKNPzhqfe4gUY8HoLtimEtexnOiDpyUbkEzLguY7NpLO0cjvW3ELV76Gb09
JOaSbDTelYUGEdhqRkUQTCA/mKNrZ4S0BcHjeSksUZIxaB9hE4jJCfjPyvny
/Zu1SOk6ksaoKt0OqV8ZNSThzXE12btkLg06RIp7lpDSKITtJ5sJ5wpzo+c6
m9lCkmSqQHYkw98u3/RFxrZ0yjfWGdvIUpL4GRlezGuzDizLimBH8i2rIlEn
J9ST1oyxr5TvN0LMQAFNIG9Cqk70+JV37eC7f5dKZPBlZogAw7Oi0lvyqgkg
ZJmaCEz8PpNnRYnQgjEXEl2TrDFc4V/85V6Q+wHNYIX6Q/AQmhDGhE9+wQSY
mj+uTbwZhBVjkV/UfFLG2sM3jfyPCaQPVkxPRgquh8aOLQqtTIfigVwfJSef
o7agtAF/WGFdLMOaTyY/1+9nvGPSU8k2HOfrftEJWA3YD/eukkdl+Nnoxdry
37GS+zl7nm0LI+8zi7Xbvsw2mao9RXvc8DpOCZOaIfUupUqAbZjWh4MxvX7D
RCnahyQzclpDyi3XJ3I523l8pDL/HRh0qrXd4kLhzq/zCv7KoZhv7p9f9ysF
2HVRTBWGBwtO7PIJ+kMLo5V8AzFnmiWVyImfLU3j0UV4FYh61dVeGA75wN2S
q15MV8VmRtOKCz2OarC7468Jqmk134RVjmyFZdhbqiTvtOz4BqEGdXy7/CBB
W+smt4G6ncC2GHJcopZe56HrmAE7PmRryMlG/aOBxl8W7kuwhBquVYtJ49SZ
jt75oNDv/ZtDd5Yo6zrq6LZ7F6AgdY/IzDL6+e/zeTWKC9spJtAvDwn/pDep
gRdLTTQmDSebZ2JwrFAqfQF9oqJUQG5Tq915MA1F+QhXOPaJ6H2RkT5TVyBb
jo5FJs9zh4QLnNEVfroXDP2w1Wgbq+PqNMzJl1ifLshC804WtMN8KFrlwaPG
ZihAW06pLAwaBZsQ9WXJvrzuXjOlZGeagNH4ohaNE2c3s+vzlLRoVBDgqtFK
KCeSeZhE8AgBNt+Wl9pzj136NYBPUcQ+N7zvDNBQnXbtXuU5In8jhtcQO6L0
I30VteypUfj8gxJrZmPTd4+yaAfj17rJOa6YR+QaNEvvighuvedf6gJoXu4m
TLJl18nm7LYCM7HE+f2jsJv2zA+nBdZwmBIlwu6rHFpDZELiA2vySO0W9QRY
Q1BB6P7EUrabyQVDTV1A7r2NNLefGtJP8A1dAZlrvht7za1WdSU3LgdEcX+A
cxG8sEAdYZNy4uUclzBEnkHDNyeTH0heh8erSJDK+4vQwk5CP692flVCXCIS
iYBZM38ZhGqWdUiZYwUJwlYy5roe2h0yO+nDYHs2DllpG3rjvE1lM8GfEBug
Nr++3Cm1TdSyL/KSC5liVj5HhZhmsZpPFR0aXjGBdJUftNsh5YmD4oXjJvXJ
tJ4G1eCKtKEapbR75eeVsNuNwpCCXKhHQEGFJw1Ojr/nocBZ3Us5ZiJFki0Q
YDEeU48hIGDZ/gh/uWddjjjmZFl9/f7meoypdUgFVo5560FfuWckNxe10Bop
jPyHGh149I90p6KM4Eu4Zv4f1UHf1F3miVeNjN4MaurAQwoK9yDX2I6rbFik
jGSUy1owK18okAJ1iZfWI94sH2u0PCKMhMOtjsePACOg4Thl/QzRZDsocmzs
Uwa3gD4FXo/q5y3mze2A66FcHpajEOfi6aFuXKU+t8AhrFELQbUkGTmgdBes
outjqHgmIGjulC49IbLPHfYdWespGoJVjWE3j8NE7a108+IajYZa0G81+1L6
T50sngV3+mtYVrXFbwSey9ko9J3GZW5/Y/Xbv3Po0fibUkAVPITwlcO86ce6
jwFZCxsSUcXNmnvPmX7PdSLp/x+wPwvF2jNntsLwNfEj5Kf4OunTiWGEJG0k
gHeZ6xUXJad4xKtDC1doy4L/6GXzYsjpvybfIuA9wQ/6Wu/Kwf3TD2y9C7AN
TwdkL5gEjwLnQE2E9/c5XjD23LA+carCONfwtOGWBKLcGq4WtkswRSjSm7Tq
LfZMPBu18t+5axNWMh3OywTRiSimMCnCHy93yk5nCMmT7eXoP+eJJetePLJT
VDCDMy48wIZIsr+k43Fkqm5N0mZ/e9El+IQAlzcqhtN1E8F9WYzabbKwxz01
0wCtE8rvJh3zapRXe5x1BhsuEeaIYg0CN59jFel5S/z0eoLIw8cQ/3MoA5Ok
+OpfEVbBMx0vZTaouw774gX4rzPY+OysEqfBj2iQFnApHlhNBj59ru7RfBpE
owr43vZ6uGyKeKgDUqnZooNp8eQjxBlasJHB+zYawP4RIu4iJvHZERabKTD7
gxBoIF5WDlr7l3RkayTkpuSvg+K+msrBwUA9YsI7R7Zdrq2TIuiVl+O+sGEc
obGG6Yhax9EqxNBv4ExLOP+McWjOgFGMuezsoy71JPGlz6Qdhtq3n1zmw/ZJ
y/w9AUbpTU1xDOmvgG/B6FgRQzU7hrsm4z3rgbZmQhojmKnHqD2kOOm8yAEW
xjIee8Vn0CUyDBZFxxeFTLZ5oQ9931GyLAJRMDqmIsDdayloAPPEAU8pdyq5
kJzWbxIcVOIir26Ju2UII9j313e0wKbnfBSVUwuJXRglCnAlHTtnFiVuyv/h
DRY6XeOeLBeK2YyM+SnyHs0fI/IIf1O0tHqDpvToXpJlMogPxohi8Jnhb94l
cmsVgjUWqlybrhcrTUWk6BnVODwfe6nxwGGO/4Z75EmHNS/fZvW0deC1vaO4
qQotJD75o3wHl8JSbu02hcqhMN+OiXGAUdI/EoZgpwH64Q218fBtUoRwtQyn
1MxRXWIKMSN6I52XOzxn7CIUyvECAApX5hgaY+qKNpbcCgih3QrqXCUsL+DA
LeA6zf+4z/7J9r8H0R6D8x7gmNpgDrv/aaDlaEOBuNdxkkBC9Rf03fM8ioYS
XLmpA84Q2f8WqjkcLDFkgzvfcUaewN7ou0xTbxpL2rgZH+Hdh28eedR/Brgs
ebMcJP1N9LjJfH/GHHWe5K4RwMV5Pe7kVGCPkmzceoR8ZB658tEy1GYTKdXU
/QPUfyREzGAa28s0ofcSWSP4PVeVFRSpeay09PZB+6VZBUjRXUI5fgklf1II
j5iW9+DirAFLqKRxB5ilhE6KLojJvtYe45uMigb3RKcKl+/8G/d7tCmKOHTC
gBXr8+sw9mhsWiBD1hTqbXWOQcGczxNTuyc+i8WL8OiD4ABpsngOIj/VMUi9
QkVFPztJhnnn4ldHFZRMfjABAP/RCJmsXyWKkPAuNScnXLoNTliOoFc2X3R4
sF34H3qGXlD+AFDBA0bL0RwlkmAZnDaV/8nkoLX/qhpDykiGcNchEo/X2yLd
cI3Fs36rtfZWYDAGv3lM9frL4iUTkNt5v1OVY9v3WMIj6bUZIGooIdyuutEA
R/2PNW25WDbC76kBvfkZqA+B4Tz142z+B6WE4KgUdv+cYgromHRzFGrZ7Km/
jXE4bhK0XBKcYBbkhj7FIKwhMzjO86S3F7cirBA40TnEodRCEXEUo6a0sGMf
RRpiTy5RHbQDexIfsLF/HrG5g6FfBzNFF4dLNy3BFpa8JdBQ7LkDz7ct+fvr
MUm09Rh7yNHqHr68X/FrwJ8EcArUUd010fVWAS6IZA8K+vNLwnabPcgsYpMJ
1M3w6hHBjs2jue1ClP38q33hfRtCIse2qwVKQYs9+CGpnbmipNVxXZGRVI+X
9kV94Ky+KpwYcPsDl60DXFvmITG9Pr8i5r2CrrHKd/ot4vGluBuPuq6Zpu7X
p62edW6L0smcecF+kCqoIehp3Ikl6PeLcERR3iZMxLcf3Fy0PnQFbMmIXFPZ
E12AyicWmwUSeUqjIXoK2HM1Bozba68zAr0mp5YJxBEKpgNsgLUaE9zPbs5V
2cHjcsxCVjI0N16y2gGPrcRMMCVApmLv0N1xMNzgxztOTUXURXfnZCSCrYYD
vapzhoXfXWDS8UCYSYcY4fp2Sx7SukdQqVr3GFCjx6kXBNbfe1ASd2rtlQHf
3/5pjAqjAeZoGtT07rYkwkZ2ur0Wo0GOIV6WtOF3LQx1rSUOaSgoiZMBxwEA
o0Kcz1hcFgb8nwQV/OELn/apjz8fWyLkF9rZRsGVuj5UPw+RsmZFyMOiNYUt
KVdzT0x3bGKYushQfrKtdjguMkpfzB2MXilKsAa2Hw1p6GohzmAU02i+2i80
kVnsGd8oqeT8yB9a4QEHUPUcInspbRFIgFXdss0BMMb/9NyJbgRcZhFWefMS
/bcTbZ9o77reD1cW3asVHJB6RfotroO9QbIomiKoylekKbqe4hKagc+Z2EK3
jsE49ZCK6lb2tdaojbYMK1mCPdJaFU23BUzhzllAdSnrvBUlz2Ur+gS0fAUl
Sw8QpHwPIXCSBdCRDvttqBHqfDXdEFwHR92GO3DrxMZVXfty5CQUcnAFG/Qz
BVGoTbfRH7G9tCjgkOf7i+ClZXhwfQ5eBfNqXnX0rurpKchkhXpOV14OgajO
TczB5K6hy757GD+en9yp0kzx1/pmSadtjBL5Edy6d8wt2Wx95tX8HwR1cF9r
yS2ialxaOxJzVxA9MsrxCIDlvhFkNTyl4OzT83ODuO0U9VHrwo2x2QyPpQyy
O1GlncaohuAsIKDj8AUL/4M/Eh1Onr+WcmK10JxbrzYTfKTQ2fcsXfVIN2Vz
tGkzhd16td6xmKiiyBtXWj85OAeI61s837ni4fVRW/IbehbyFT/EXs0iv2fD
BZnQsP+/qCdfiKjJkDxyndghN3TSbbmF2egKRo9CErFWu7fGvkEWFKhQof3b
nua2IvyvR5UUk/uv5fm/WXY5F5MybhVMhNPN9/csindWtAfzJWGz83Xp2E2z
oG0yYkqxPktLO6aVYI6HBG8dZNxHNxfFUSVAR+1WV3wYNrwOPDnSa8s0RCFT
UhEZZ4tQTGQW5h/r88IPwACrgPUYXETBvzbWZggHCiK/HaoM7ty6TmG1zxye
5cQu72T3Yhi2ACiPhLeWhY8aD1vq1PBBD8ZZa4EPiwM40Z8NST/d5Rppfp+O
n3v5sEMhUGVY8Vf68bWrdO3wgUiP1SbYJ9LjXf71cLAQHH03YR6S90s6Qzfv
qsIbIqXSaqQD7HJFNczHGeo8Z8bilY5/Tj3G7mkjzjd74ZNxjHxqoH3AZq39
mugR6p4N5MzrZcr2e4H339NDO9D97IGNUia5VjZzB8S8Qte+srMmCmk6OasV
Nctp+dJaHkuwG9pXv3+6o1eSF1avLyCz5BS9Deq3FYOTMHSPVarpmZf5ig2u
qXSkaKyE7dlhxIvNZ/Sstx/in3Le1xPagktxjXP9lLqxts/+cUutl0G3ZHd8
BqF9SLwqjKl4FuCRWM7mGwMLMeCPi0rRJNs62fq0j4xlKgHC6zROuDwDFaot
OJY7fVaj0NRbRs8GEcu8K2576ahKy4YHD3+ZS3BH6pcZmZGdtAB8O5KNv7vx
7GiMOAybyfrGoZ5wsUAL53AnmbGSA86e9Nm2mwWcEgXUIaBBStYm6yK3QKq7
KGugF4+AexJ0QzS/cG1l/gt9+Dzp5XxVghMcrIIp00naKRSJuVhxNoflrNKJ
Cp07hY5a+S6kuJrZ3k3YnpxJRAUqtmo8ahLLfi/YWL+JTd3tAgkKmzI2rh7Y
OidqIryPcTBjXgPvHohN50PfHdRdl+7JtOi7Ef2ioZIW+YA3b/RN3FDTQu1k
0wuPu0EGeSnPXRML93MKTe2fi4bBmsEOL4ZGg91NtqD/M+o9V6hhwT54pcQU
KKKQA/c+RxEcd8Gz2EkLOQzZLNN1WvvAxq8RKLfjYtkVKLo37ON2OLzhQ1rI
lzo/BTY4q8XrfvV5eQ008aznQByJF/2GKBW66W90bHxBXkGkJcBZsV25C06T
yY0nWdrWavyk1AaK8n8OBsA8wWEbg/bKYpeqq74xRBiq10pbWVnVpSLwtgqa
E/lMaF/KIPP8OME64obcgvB4+8NYilynWbGAHVvN6NMpqltd24Ihnt6VvHdW
sMHrMVU7zKzD6zRQwaDdInJo1JSyCDWTRVU8OqCcFV97+tGtBf08PHqHOkwP
4pJ8sg4r1jIc+ZjdhGuty20lybCnRRfEnZ5STuXmKXhQdIk41+MmlVazqFfD
88vU3MRmQFCluWRDzoGetLq0crBssMxWgZr3O6GeXFWCOPYlu41zH7DEPaUN
gPCtSiIl41/f4mPoLodRX0GXAL726kttTq3jIuQcqFEnNBiEivjq9/cLVz8M
qsrxeiMy0NL3+GWeqPfoAS+x4Wr8x228lHirj/epRaoXmAmcUe0qpuz0JK7v
XEvJkBTkN8SUql05pijmpupEMPRxEhoUPWZZnpjhPbW6NLFLwXtALdcdLZug
37cbW4icJ+mIohmIHzlyPuPU6MMDgLVOa7yEEdHdsI4DMt4zN6wQoMhmEEih
OIn0O81bovCtUnY1aE2rYpAK+c25QpNVdhCeGHEy+h8OUgb69WXfakRtsDrC
rKKKsH7K9ObZ+YjffWN+WqkB6YgtTOZ94/iZNx62wzDdB35+UuIB80izVbuV
v+As0ihsnCLxbyGt5XxSTlMcINA3+jQgAkY+qVoWSGnu2zZ3ZzcscMf6+jfB
9aDg3GfYCEyELRsjr+L44OO6ulGU+K9X0bp6j39gEu1nXywER15SmTa64roY
Ea20aEFJRmDI5h57uUCJW9Udwi5LJyce/j0c+D3jXDhB/puS+rEjsCzZW88G
QveVtXLkaAYK9C8abE7h6cTltyGXHKDcTre7/htaLKdc4rUTthcmkEMQc0/p
rGs7ikHEwTAvpwaBmlglpDt3hWPaGC6jq2T4RJn0jEvkjdgAYMueoDDcNtQK
IYoMYKEdzRoZPiE/b7QbILQ7e9L7JvJ7oSpno6unyaM05Y5cpvBKaW9NEy0o
AI2MAAry04/Tl7gxtqiojw7kw8o0mR25rTcVyEPWcwj25yEhHEvbs82UcAuh
e4nFHEBlkp2p6xjzRGML3KUd6nFTfwHw8Vfz/VpqrfK7g17JgLesIFxjy76D
F7v1SZhvirI3xlAOr9tubzIauLC25lwFr0+L+YBn7Nrv81ukidsghcZyKLBG
pQ3YDe/15cV+eaX/o/py6IABvcDEAoBu4X5WxrS05LefgSdDD6krmRAyBMod
ToXMmsAJHsFW6+slFihyXQk3O3mawP2O/TUV3V6EYOGslTxzQ46zyNajrXPq
k5Y97RZ+6DYm6ZKITsZ27mEm/TSygn/uD8lvYDyEUPxMfxqk5SE7yxiGec6f
Z+XtMnz9aq2DP03ua6iJGmfVAB6/MR/euH2V7dc5SBZQZBeq7zOGBKnkwZVB
EPIMWkwCZ139UpKUjcsdz9nx2ZkgoPYfr2vA62sioJOnLYbksQBg9RDdniJL
yfhz0p7JQCQI+RlVwU8zoEcDP5RSEi+T7kdoZX7svHJlanTCBGhdkmPJSZlF
uFIWLUbvPUs2tbCNVujQYBHaqVCz/3lWGARtQHl5l0ydhOQHpMyEeZD5uHbV
S4tl36of2ncxvsLpc6cGCr3TFtn2NTe7EkVnx2Aj/nKe9d/SDfXll3L0OQr5
yb8y6b6WXaA1Ywh039r5vLFq10zGZSYm7LTJ3zJ1oIKYIeuugPkAUv3F6j8c
mfgWgUWNSUTHkG0IvFFWJM9NbXj5L9LgyufVRV+BAIBKnWEmmLd2jDHMYd0e
kNxk69bqRf5JaDT4VXJxEtseGuSYDkD9KXT+uGT6hfYZn95DCqT9GO/760Up
ic9U53a0GPT1IYGUcVpZTKwMNxKbkUWDZ4VR83D7ysycvhL2PlKSTU5Jxixx
Q61TRiS7/5j/Nku0L5cX/dJ5hu1IUUFmN+tCqYzCpJZ7wJe/VRWD/705eZoB
CsAIjwcasu6tIYAnNQURFrvC33R8PM2ftAtAyjQoGZQPs92yvEaqrLIV3KkJ
+AWAY5a+fruUYrz+xK8SCAKb4wEgAB/MnqyqWKrtr7PJGUJJ+SzB+Pq6hGqz
n8fg68IpVOf/HxylmaUwMEicI0asn/3kiz+akxFrSmc31lJEXrjIY1AEuN0u
R7zAxRFSX8LMCXBbRIbLm/t0DzvzC5yi4y/7gLNdarSi7qDTcJb5vdMZj+zg
vDw3Hv29Fbu3aTrHoMQrjeiQeE8b6GD6nuZ+9QhR0AM9Rh9+bOmomxgCubRP
woczt+4h2JQOYcU35CuvVXI28Bj7AvN2fu31LOq/meRUPES1Hzc5QtTMvE4J
bmgyCkTYr41tGeeW8kBGg1sy+eDkBhhmvydauPUeS0f+2wVFet31QC4e9/IG
9We5IIAGYZ7V0WUHWjuM9fySXv53ZPdlt3UsZ4twk4Pd2IS6kRaG34t2PU5L
1q9aEc5cBMspyCrdL9aVQj1HSLyiqgrw+FPQyqJNJG+aqCMAr8elT3Omp92i
+LcfCSdoEO5U4jckjdsUIAmWV1zGRvT4vAjP6uLj8vy5tOZntCmtrR/aNTzG
V2b71E0u/Fa4oN8MdWa/iny78JAdLWIfPC2pSmzTGUJxv1TiOMgBUiFYvp/S
Z0RNdGz075+0CCsKhaSuy8vEjbkXmGWnRe0IZEk2wby0uyNsu0jGfXg5+sjs
GQBPXVbr/F1w9RSvdr1gcZyL0rY8hjkLYBP6PCV5mvjkEhnUZY9lpnvbmNNU
+h8KgCnEv3S097QvLm1P2Prrvc+13VGg5bZ/C88lQihWiuUcpZDquedcLbil
FK14Usf1stNOzWX3bbZVN4gDZnm46pl+yxi0un23XuAXqT5DStyqYI5sIK97
z5xem6MJxJGDz1M8ff6ViFrZd1skRBCFbBV8IBJmFZ0QvVtjLFPWGecp61j5
Imgj7sHGkRdNr24d5K5OQpMNu88gyXuc2QUC18gSAlyCYbPhbMes6arwuLRn
h5GURTeoU+2XLTmilwWD6z27Sm9qKxHCy0GKdsp715CZdU5qeM+drBuRPsLo
1eRrQjVslS/YAfqhiSLo8P8s3yeggFp4qsrbLcqNPKL15GktU/8hBYH/tX1D
PlYW4OQ4qkd3bk94qZknQnR0S3Hj7CagDQ+UP0JEHyYEDwDwF1ddDrCsYnjw
urSflvAe3h4LGulox1ENk/EqZhmSqlhUOfWIOpoVUms7PxZNtUZ6VaoTPXw0
5Lk/qNjVbJIqnmAxMKOFJLGgMHHDAMiWR1pUXQYsCS59Bp5E4RQY6f5kz6v7
nhmMbO2mTdntL+BMTuPor5+guflh5i/92lUOgC89tg9WFkMINzYJtLwImzbM
gNJrLa1Tx8bhjCVrkvx/XKJS5/rHSF1N/rdUzx7u+75vWQwoNZQTC2GJo3fT
9Rn/DJwapUm4VsRqgHKoHRlrXUSynbpWh9xmwm4OWAyb3NMQqXZLoA5PCz63
SIs5Je2IloxmdGpvGiDjTU6vQHwyg4hj9Wez9CRp0fDmPoZfNQ3/lOECi/r6
1junKdwg/8uMNO9hy4MpLELRBojpVpw9j/avPkWu4GH5x8fyQW7eLia4JsXo
GS82PeOTCswtLgfUFusyNWYStO/Lrgx8ghP4oLq+pP9uHqRfdPjf4jEs4k0k
NMz7KTUzEoiK9LcElGtkoAI5oQCh4OCtvyrvrgIuvKWMf+W6oMVxrPD5QIeh
JxVMHCcd6mmeun4nebsEIePjU6iqrtkxPPSdCPhAbbJD/fVO3/AmCkH6Orml
GqVPFNvbnpZVQaoB3MKqWXEtOQ/AG8az3g4Ta/bLD5tibzvoKfIFWbQf8jYd
ZK70ea+L4cATgbhQRt/lrLcLnxfk5zFEDxdYiL8gD9BqANVYvlWYLYqAC1s3
kfID9K78Zny3q1NZJ6+ZzBvL9WnUmRgBJiBwC7wZTIMWtJZRqOHJ5FoJyXQC
xVsEsIVkqBuByp9lq2FxNOj6ozlWMgk/5qQ6pcBoiG2lJpZEI9R0HaYaKe6Y
0Hbj0WnhyYJLZ6lL5uwHF2Wb40+euFW2+MwEJI2q8NsTnEJ4gTn5PsjO5frW
Td+xY1z0+WJs2xQq429lehHmTidZs3bqqc/c5DzK2nTFtONJ791St2ojgVbO
ekdYBS0DsKHMbiEBaSaxAytIu+kJZmm7iKzfV3acwUbP+x14hZqSo23KV+1w
9GO1h7bEFlRbxIZe8Yx1KKLAK1COVXpz7Z0dfGb8AEyI3wTmKXYsstr3yQwI
tjFhYj4Wm+CW1TJiFkydpicVwMxQzxkmc4upgntcGZYyrTlsoHS4YXYv6Ayj
wmk/bRwmuF2YuU+2/5TyuV+ZMV0tBXGBvkEbBE4oLcPD7lHnkZB0MXwPQv8Z
a3GTPncnc0UKm9LTJpkNQzpi9oASTJTpvbMj8KIIXwSt508zCz2+Sp2cE3RD
d9m+6+tmXdmmq0IKjqnKYElfHK54I3KJ6AYeB2cOuu16vSUVlQxsANrdaBxG
js53x0fPrPLwCQ+I6m3ej601y+ngfhH2E4ugD6Dhwpk8xljpSqxbda/bvnpO
t2SZL6foVlNUlYX9dw4R7BLTrPSnRpAIXt5wuZwBLCxWGJp7aorXgpB0UGTh
9w21ma97VjhVkpeXbEzsY9/TF3muDbEROEPSBGGiW59ikuUBKeTdPZPsavHC
ajrr0A500AdO4aBmfcOOf8GrvZEC4CFTQnYpAP5SQcluoJzAmIJgqx5noIMz
1V4bAZSdy77b5dzuej5TrVqosFY1DsszSi2ydLYY0yU9nDuBvkEczTEZ/Q2A
c0iHfXumUSUQbDSZMAH4Ajgpjk6SLKPO/N2krI8ZLNdffapScsCZwCqQcmx7
sr5zgPMZ6nbluiV82mfo/tQ0ENRuXywCq2qL0na5uARK5+IuI5/It4mRuSpO
xpRkJkcq06gq+dZvmZNxrp4G9EFtnIX8oMo1MJzXedyzqlIpJfISw9XBMTfb
JYbfva69jTFMbke5qY/f7m6u6I94RqMdmV0IujixYp0s8H8AAPioUVMRz+CC
Omv1FJTTEnA8j+27I4+pBLrOAbfFVMLnQliMPLiMwCjbQ+EOcMyhWINeIqXY
+tWVduKSS4ueVYXNhY/kuyvswjoKC4ejpXaQ9CtmZJ7cygFKuX2A+iy7NPTI
T3S1EU6opI8AEBD0AU4D0JrJA4oujq5+lAieCQi0NsKiley21/sz+Wedh25I
nhappt6tcB8NnS/VLlUoxQQNTyYV5SiPUjLbYPyvGeSXkaPnR2xLU3Um9KwS
7Gj2JTdbskv5+hg1UDYmV0m0Q0sX5VDf4GSRTXzS1a+gC9nNcpgauSrT9ucA
7UtmccbmwawyD7rHiSnire20EqvVThARQeaNoXkllM9rQMWXmPlRthrZyH1z
5c8jnk+PbnQ1Bh1RJOoniq4ouuMbemIEhuPNA+fT/TQLIydTyXkwvPTFRCVu
uGkbFWpdrApLQCHtZJokpsS5CqJ/moX6hDPJNeiZrmi0toga4hbxQDQgywjS
IpSrP8vJm+gOTyDvgIJfsI8T+vYrE2sRlzoRDynapr41lx3NH5kVqmE37uVj
OIO9nMFiYB8/qrnmA5bRDnH7IK9dCG3GZDo7SjVGjiRm4UCRDO7pSPfL5ZBm
PpTyG+nEnpMyNVXNjdSXyOfaHVolGzyVqox42x99FDF92GrGhvD6gBXBKEr3
OKX+0eeHDleUOcliOlb1y5dAq6Tvz8wFRuqBFVXqQ9cPLORzaAB9lX6kwOiU
5zhUOAAl0kJKcuataVKlo/xz/zT0CDtBEdBmVyuyb4u3QLFwa+xJN0zAbaFK
2ZUI2YTCxytdoI7ELUR4pnri8lVB+FnQAz41P6sKTv+Stscp53i1jHq2I5Wz
W3NJblemWKILfJpnE8QHILSGFw6lTwiGVcu2XCuB++2W7ueLC57HvXpecRTL
f+srovaJz1nMkqUAE+oBPLDiqX3L7yXpe+rKY1EGdNmQSTm4T3ovSHbHwycF
RFPS9xf0qT0KtRZo4MzL1BdQnNw3V0nz9B73ayUUULrn6vDfR3oE+yzqrVmp
FCoxSWho6bsfwV8e7lekUaNyf+chC6LA0JclCmO+E2H3g6veesShqlznJvJI
rpjCO6t9IUybYEGphKNumqXuHRINlSUBAsnqq3NA9Hox2wrZVJu2BfDCiHZn
/U7xkKeAmiW+8DS7jx5//8MEzn7gjzno6WgLmwgvWmXdrmqT5pTzdbeyFjHl
0n2J3Q5C8KvmkonNmalzt/fC5NDrKVxiwXlBfOE2QH7Jp7VnMBdqJ41wzLpT
NINe+erG1KwiDjM7G9bCSfVI2anndeMcwyBV4F8z6HCyRHa8Z19OOvq5Hbs3
20ysegsY2IprILRIpPPUZ3TwSJAjJpK5guhnBfSfqzY0fsft5icZXGzGbvAX
RCtJcPLWEOxwWCGi3t+Pun4Hc2m2Tx1WliTAdNFLVkhdts4Xo5ujkohAbDPs
jN2NPwLicC+L9xUS3RQq9Iotj+lt0paTmahVZ0UjYvdbIVZf/vND2vWioHsR
KjyRxfvsQbKQYIiyeOv1/hCKfBYbNuSnAf1M6dCunxLQUwYmKnykbtl3O5N/
3spxQr82mD+T+PMHbMunPjp+/AV3jTHlyMEQQ91znAYjdZMETM5XxCoNoLFg
JKDU7pwxoZkm0r9f1+2yV095j7iWjWjl3Zbg08C6Hhjz4iQ76C2wsNNL1iOG
E9hKP+a05MeoFrnZqI41GG5MCvjThHqhSKd6q2uveEefoaDPMYYKyyZL2W5U
yDzmvpPyOV7g8o0uqyIs11q+PHKBFz8Q4XDppGqbGKC3kX0i5ipF2jk6xTVS
bTJrUMmXs31ab0wck2g+pV0qoKeT9ZTvlG3HVCqXfMESahynI7U8WbUo19y9
6fWo5fN7WaEo7624Nj6Zi1B/EpDVNoNgK71wUkitJLRb6mw+MyhTmzsHhxEj
wvyY2SExBAVFLP6Zf+77+scT3iGegZwMfkXWUmsCMrlO+YxftEPch+UEcaxX
V0Ky+UwVHUlP7E9UA7REO9sXZi/KxRC/zV7cHfd2TLrsiURAbg8aNoNlSBoT
y9McQtT8ywArm9DdLV4J7jiJISwHrIjXnPIRTdTO5s7DH2G3SLxdkPxEERZ9
H70iYjCQbvX9p9uDJ/rLJb17RhyZmT80Rpz+g89oitOe5piSk2SrbMG1a1hm
j3M2LNYk9yBYxzWFbHvOsKo1kTrCF5EAaVK/A3gVP0Q1o1zVc7ygsWgawqap
kVYoh00CnaWZWe2VWe7ZO+q3iVDoqsrqoWTYOXK0BsmrhcIi7T/uxMfChIWi
Pv28oFV80LQAXogl2oTgzDvgW2igZvnAH1rYCBPgGCPgNt2ffdvtCaZrDQ7r
rlziFoTv/RyOiUoTx7DgFKV7CNLYrAerC86kku3kNPMcXfOSg87ZF9yLZg9O
hwi0i+NDnFOCgKW4fc8ciVqPLlFvUXjg16SoE4wHaMCsqOuaJrg6BlhQtwn7
1lzaxvFtSWB1iokTQEdhBAWmEleOlBcIHG+xwSzB6nxOFHTwKPDfCVr9K1Su
JYmDkHNkgIn+S9pGqiMSYPhJ7XeaTFKHzWNtoGKpWAbtLstf812tjzMYkjo7
TMOvnOT1ETiWTYGR3qv+0qPa0uI5RZCm9JM2fe4LAg0P73Jkz+QFH63e7KlB
h9K3uiiNKLI4A1mo9TBoY0M/1g6Ap7foNn6fGX0oSRUNa/uG17uPbn0ug+IM
GK61uq7cz+V0D8GhCQkSyn0xH/giAk5RA97Tt53wQOszE5OJhF8ndvZQ8J/S
G9TcAP22A6hBJ6qSL+XZ7iQjmr7bqaKflOPgwOYmRt58kfAO1ToOWh4EIwrM
s1tlzceDKyrsLTCEua/C1uBUAxkvYWiihReRfmUZYckn5hj0NE6GK8yOsyJe
+OL+h/7kZ4v77S5tLYccbNJXIGjYt4wbzHODPg3Lqpij2UW+KT9c0Z1T/Mu9
xEQ40M/nQuGP2+zp4aPV4UEgiNAMKm6ea4b18iAb6hS6NyAlhsQj6SjfNX30
iMEPP0guad+kSN0tdC0wYdmAPXfNP3PMMA8weYWs9pB8LZwMKFidKJWbNb5D
pePdIt4bTQGIicznSC3A5l+hKEeiFsEE9ebLSGi3liHVcn1v2vk04gIRW77B
zYYlpf+NooNf97zwqQItlz2GY51DTsH0QQFePsdy7EAij3BYvKIIC4o8Ux5b
izrvHn/XAO+UtJXYcVZuEAzSn08iOmM1VuVDWa1y5V84sRIZTqsTctNXVk/J
XM3baGiL1OEk5ubWfIDN6sZFl3x89SPaBtsSForYdOhFLqzYaOKuQlbXp+9+
dieHtt8YQlTG3WCuyV2rsbwC6A5l6YajXDozIIo5wc5flf3KmlCYLDCMnx95
WrpfFLHO153ne7EyXXd5teakRkiAVoeyc5Pq82DiJCo5jgqqa8TP42ulCWpB
LPEYhXfrL8nZ9qFHA3tMsX6FpD42YTlt7jfdcuEWchj8BRWba0aUd0h2dJUu
BPBubM8ZjUyhb/On9ggyVOg/egJuZTvzTquM9nRVkXOsnm7u0mataebyEgG/
TW2e0ez7WMP0wAucF8XWwjwvRhvCKQWpRg/W0ZMG94i4MPuDmubQmwcc3tMN
ZrghTV1hyh2lTMaP9v3gpExvgOEl2Nvjqh6GYlFm+mizDLhNLb+YYqPDffZw
XNCRYoJTVxK+RnjiSTw9e16wVfkpFFqSS4QAwQfm6DR8prUF6if6T8fE3b70
g0aXiABJKp+CTu2KAi2r5ZMwh7Ybk+nJOAXHOXIyuBvaMrtuD6pH0mRatN4r
Ac66SvH9DIraDCp9hr3oB8OOvBcAuzBCVXElearbo/zZ1FIeitYqVuUIWgVG
6aat0biB6havEiMvPKZGa6xwockWo3rA0oG1Tn/T1eGV935O5eV+//VdmicF
ucySQjXyeDerp+9oMARCYoKBmwR8J9Ubfjuli1uUcyEu9sYci55xOQXWu9p4
lkaTbpSiwV8GxDD57AZYa/TN5phDxukZDEBhpW5ajCkh7AWEkq16raEnskM/
dcXgx+4QtDTs/15uNLaXSjIePORGm6WBqqwESRfaLWyj21lk5rwIHqtDsS7u
4bP6RSmE82/hCm/y34+xzLCYm+3KSSl/5F9Z3ftle7NuGvQWJfNyu119hlgi
f5acOoVGMxRYrS4qm3FUqxDQa1Baf+FLFNwYTLoMGnq/RiR0Mrx6RVNB979H
Omrq+Zjh38XeZg4pmNxBwmOIQVrSPb7li534SvDoHXppHc3N7e65ZFUgpOlJ
11XvFk30/m5Imq0fLvAFBabjXkIG/48wI1IE3qNc1RvVTwcCJHrVqLJXcevL
C6HRAautpjIgHqminOMds/drH4erh6RZZ8/XD1pKQ4fSyAMNj13xgppLl4hg
CQSzNN1CYninMmgNPpbxnfz1IAIp+d9Ed2qdxhcK7z1s4RGS3QJYL0klDePU
5UPZKtiggL8ehjm2rOLCgETJwaHDBoaytsvnjavPNtLBZJNZKR5nuGEPSCCx
o92SrmbB8g0BlY9Q2iQ3fla7zsYboRcQSbKy3O6znQ3CRUR80WyYEZJBuurG
9en2rGx6OAT6gxcmZVl22kra+qpaVAyooE8FB9C3Xi5T5Tqs7MHZeLfj6MNq
xGJAhqy1HD+qW7qjQrQmJm4ynouBoQodE+DfuoBAKfxAD/KTb2fuVbpdlBEP
cTXfNFb1HcBJALLGboR3iwPjWx41PjT5pJSVQ/NcvydJZycDNVjdDIufL4TF
iz7pT46/a67uyWeoc2CzepIdGlihl48b9WW35jWXaLzCv0FSy1gsJFtcIkLi
eCKJojkLdAS44LJTsRlJGt1q8WPrqekKyyza0icLPHd6FQT8+pmznjvE+bH4
kcu8pbqanO7mK2hFPS0DiY916NTMOY0j5O7ddd8Y1FcbtJUpRFw0pa23A+WM
jYJdBIR3J/tMGGF3AI++lZXr6npySDFQ7/6wMvnbXwXBc0qSlcIr+eJ8hTer
FABK4ktLagtXAAA9i2iTrCzbBX5eaXO14P/rqdgjuRgsk6+q8Ll6BwYUiDOT
Rxe15+L1pPLLCfVYiTiBkQKBURHBM6n2Ql5uvPkOkT7JZzkShMQKQkLffeI7
Qudg955tP2HOCAFE3ucp1Dy/eb/evqXyw7ex1lCco8zsueIYrF6+Gngn2sL/
fqz4nf41zg9OQMhVdwrIkEoTkjtVsJdsCqzSEdn3N2zsDPYUVfd0Oo9QVn33
k3vZNueK06lE+XCsNoIGWdJETNrOPoTDLrOJatSLRfizR3LMOyzqNzV9joo/
ADnizHsSj4PJW50XAhOqwJ1tqXfUAZ6cLBWKCLLSyfzZ935ZkIo8PhsKQnLD
DgblRsfIT00v1GkD4j/EoEpWge+nQLsgeGq5rzDd/ySi1oFeZn220k4IXwAC
XE02hn1jCXMYS+FCZn+eKVIphV8NzhX8WEcFJVDcQd3yobSi7oHboldY4ZWp
EJusCJapoY543retDNSVwwVlB4EZemD84Ex5OcPDU3Ci4qb9FrKU90+KGy+A
M82M7B0qDjONcUjcDNpKdwrs55Y27+X23YpWUSNoMqBaJMTbuWGLvcUKmiry
gK1ZIRx4PBpnLSBTUSOLQnFg02h4G4jMa51llC8wJaWZh/NgRm3jKaKjHFA2
6hLOpwIfqod/aePk80jeHVvU+VdaqKWMgEYfxvp0UaYsw+yWkn/r6xnMyUtu
CGnRu1Eg7T2mK6uR8NiED1nj9Iwko2xoCYRhx5jqDtwdCXFB1/K6T9eRThY4
leehHz8d4xWgnlJaf40AVLnKaR3R9JmWmTmYX8lPM4FYJDuOKlFp0lo4zgqM
xdsgwr3pvengamuOG9Ah3pL5YKyMxUqMdvejd1QfpMhz3cJdDEGzSnEaPq9c
jRDcUgk6BOo+b4/r4UmXehxuH7mgFD7GGKh9WS4+e88vl6yR0XOcGkxFMg3W
HsUf1GxG1s3afD8sIagb0zYTbNGdI/O8LZJC8JW7r/4o3mkBvveHmj2L22Gn
bFUxRsBq5ch/8bhqA8zKWHXGSwMh0vVKPtlYxZLte2CA4nuK3Nm6oYabvdog
cl8uRZ1i20mgmpSSF5nVPcFYMWEZgD9CLSFLXhhX4pZJakCAQaLPe1Y6KBwj
1J+R0z1wLPVNrlAIhf5oE2Y8LPbM7BLyvKagF4+6Z0n1rt3d8SnGkukWgxDn
mPdOK7rIvVzO6szY7Eoqt+DVgUIuMkf5POEDcKtsDet/mZPCaI3yt2d4JzS3
PYj3C86Tw61STma9RX0crE30Z79SW+YWKyWOw3Az6GXCdxInh3BRdEWKkzRL
uaQvpAzcDmL7zKiiz5wt7BkUpuAlqVtrUMtAA1fI/GAGgqScmBXwT1FQiB2o
ExyGAr672qZH5wDVY1DiygW+ooH7D0E+knCovZh/oajCdvREKunB9UkbfOXW
sODM8ck1ERbGw9zQ8LokAtiVFOKf+/Odn/5IJXvAC0lHXPZbNs/LYL8etihW
ik42wQ981r2cfuCuDUZkaryIp0WqvuSITzjtwzxPcDujBjCzA4Mrfy3haDTK
w2Czcnyvh02w7QpRm7RHlBr37Xx+0z9QyZwDId7K7Veu41zEEBEH1jZMinm3
RCcc3umD2C9lbjJhDSs+3OIoMOcLTiKvczzj0RFqIAyBwzyb22c+gEUuXt3p
DcmSL83X6ehFmaOLWNfaZEzOFrGZybbKHjjD3saEImFKpphOjPdC5qVIildA
SJ/C2suN/UKg4xIXVui4Ukh6QhbMDvx7WJKJ22rjztRQQvDVGnsVW3ViDl/8
hBn2gr2YLcuWjzwxw2p5KCfDPU+W3KrWyjrupvcUCMRjJ5ZAMRGBFaTcDtjg
LLw/y02dRd6ObLd4AdVyTZKUTA0mniUbItpBi+Mvao4vsB2stWg35V3YH3eH
QOoYUFYbXlmsh4JqmAox2XqDChd1Bt/Y0g6owTSBlcxvNNpyuz+2nMubrBXa
SOX0/g97mrB46g0Ny49dlUcCH38RWha5rnXNF/5FZ6PlGV1eNoY5xoWvc1Rp
zie5Hrm/IQThMVeGWMZ0xAQvlwZ41MPhcpuffFAR/sE2FS3YgtN8EV8k06BS
nR/7nC7+jcxg1BmsMWwUDIWsqwBTz8w7DsfaWckVDcWB8WHsTLhsJdGLf+6U
pu3E04oT7PYklawAHK/Pmbr14OCtguHbFz8FzHYQmtIiwSUPu4pk0S4CQZoq
BYg5GWzP9+n8hPlTTT+q1KDfhLMOJ59psOXHnVq/EBbnat6nmXPlJ41dUEpM
ALMJwpyDwKipIEDY/XRiMcDgygbqZWES6tZam4gFn0B3AwP1+rK3e5fMrxhc
68K8fgWETIwEgOIReB6UdYe2xG6pX9DmfZeZg64ANZd3U4IjTNriwDaTJIej
hIKOz6z6BSMXA+/09t5kP4MbV131GtsI9KX92sgsvf3IMLJ2pf4B9OfXr4YA
C/XPi+MYdIRaq5e5jYUUSwMcbsXzb0UYI3PujLgwpJJ4+noym9ISf8UJE2bl
vFy+TMlY9D/a6lEaqoScDv8cxNyf3ve6+8YsX8IofLm8BOAKOtvMhvp/j/op
SdjSvYrJ7szrROumKoreFsMY7DDKl1jgI+KnaVe/uJZND8MxhY3V7aBzx86H
BtwI+4GwHA4pedV6ka/WrYyU37FCGoUPejN8lZ4l9e9ndA9l0QW9ZxfGdBkE
CGIdc3S5RKOlmUnFmU7u4QSG2dsyRZTWYE0lC1hg0rVKwSUVIS/M9FeuKWgy
kKXRQiVec7RJfFPVnEZNItkf7pde8D6H5jFhjJXGVcI0rw2oOtaG4d4fcJMA
ye4jJsLEhHWdHPBXJMEEeFZwcd3a5nFH0tfrXmxAeCpuZtiwB7edyKBiBmaE
nwU/hl6UyQ+87Z55OFPHoFBiNRUj67ZrqgTQ6+5lAvCdIv9mt0kJiO1kiWoH
Q/RxzOQcBGyXdfNVp9R9ypZ/wktSP2sMEup/YbzPlSmgu/s9ZwksBrtLrNQw
itR8MwpMJXur3OPWYeCj/8TzWj45WZaKhaIW7X15n4tWxuNCwz4aIM19GW/+
Axv+GT3lvVmCS2tbRAiMMTsY5aNQKT6VFZvZ69sQ1M8EKPbT5stSW1IgdYsm
loLaAS/5vfgLbeECn50mWaZMCV5cEsYMTwofGSUwmU32ErcDrWxexVkEaPIP
CsRaIMH14Y0W/9bqXwjt+ztmvxIQY1Qlc/M6PhkffBiFX/nWwWdjATYtRxIi
XXHcn7WlWATWBq6hp/GduLdNfZpU6gSEU/LlFaLwOdxAKUZIILWXLsFncuL0
bEnkMirqywbn0p6MnenyjbqEsQtO5K4rzZ5SV4tpzy19OyktT/1tbQyWjnA4
5+k3Y7tPYTK2bH7leGFTSPZ+IkJwTNEJPNqhECYxlHhg62NcyB23E1QBKL5F
gNXlFcU6fFTXd8qPeNQsVvDh5EwGvPgzASaSbDOvhGDGNxGut6y2ZDW1+91E
6Xj7j43Eba2HWZSegcvcbDQ9UAKMTMGH1iICadSWVU79g1dgXq+Q0KO6IiO9
amElGSb3eonMlf0/FNke6dUY1EZXiQQz0zE9gcBWJiOXSeCzMf83HVTgkme2
wL6gHuCw2y6ndauVLw4hqzfpyjJM215fQszLIW0/h4uHdkTyj57ph72GL4+4
fGGwNxpt+Ihw/i4MpSz6nW1aZtAz+1a/P7iF3viJ6uLoO2ADf1j1KS8QUhwe
79jZq91hG+NklWnr7o9DsDEUdAcKw3V6/ACSLhm/P/NTm2U+FqKbZSqwM6DR
JMD4DjwuA++9KpEsN7RF4pb02t1POtwHkd1hPUoIcGKrAUZqZCklSyTJwQ5V
uLPqdutq+lcb1zPri4cA6goJ4CgrGvgzZoggkkt+8VDQ+cdt9Ayh85a0DI7/
Xkd4M5nKAASreib7zV+LZN+zhhXSw5/ikYTmTrlAcjiQ4fR18kJGdCXrQFwp
bpBE6sDNrBTchBQy0Vhon6Pe4Uuax/QAYT4szf4cgdOmm6YwmAxf8J1WcVbm
fO6zTunPWW2xiZmFgG9/OXtOiGyg8nVeZUI/WX7i2gzwCHgYx0h+tJtCvIob
moWSWPPs8JSJYv4R6Rx16uslIivMCym8RnT+MXQKcrCii9jEDwkCU4mIcgOL
FhhYtL2opFGip3TjBj6zWGEw//ZuA2FEdlKrStxs7yXOhPMYljLQoDGvClpr
Hqup741FZVzfBF+0WeazmTVAOG1fMCU4q2xujtaX+Dp/ZB+cdTKArk65fei0
F8nTUQnZqVK0zBJ3rqRlrj7IDr+K1uddguvhlM2u/4INWQW6IzX9zyLPFP9z
LWQGx87VnplHCKUY8AiVr3OBbXRjSnr44KeyWSzpuwyT4Tq7lqx9nSz6mF6Y
IVUy+BMuc6+1P/NgjO70vCVClmweyCJEDLhlZsI0kDrivH4C6KS6yVg+zLRt
7kAbMJzmGh9PPpLPE8/NV3yakDOg/lBkr+CHVnFofXqNmkkVlSQyXdu84NAF
Ju+sJ7YgReUCHVQqkKpdNKxGSqOtHFi/cj8KAeiD6X39C6YJeI4cCmHWQ8EM
gC1cCMi0K0VSdwLYd6GaWOYtmh1MsZGC4iecaVZaxDdt+uyIrk+w+GAJY/d8
eV4rFbvDer36Sq0xqJ055RVUqrN+3EpTiVegayO74GxStP+DRoqIqr/8EsfY
HSjo/ubiHdLvoXxURNeA1bZq4jcLqX4hwJpz/7FZ2AN1nEd6WrytsC2dgvdx
B1GAZJ6lrvgDHh2YR5j0XUxy4VzC7C+mpbkfzVohJDWSkSEcabOPrmRhN4qo
NdrtUaxcrvfDyaa4OC7GyrBZewiBXPSOMr8YPC2nO6tmVdSBp2jULJKmN+Ja
ESess/XnODUNlnYXD1Uw3BKW1t3RRYsesKI0v3MQ7NRa4fmwhp+tgEmkHJvD
MzOOHzE3REtvYnPCxCuZ/J5mv+o+zfcyyru7ZX7kBLqQSrT+1a8pLR4hmVgO
6UAeuNeIwRxjNSYJtS7dxEwWkzks4MTw1iFjzF6UZxMiTbLDs+8fPvYbNfiF
2wyUywf8TeFzQFk7bMW9OsuJlRxYYV5sb6ggtkSpACcrGqU+7mvuyNqiLMzA
30glZYBY/JUhdpSVQQ7gS3Bk03ean4awo2iszFPrHNu3Q1zXmGiNxMTV2QGz
N7wzCfgePy+L+LRJI+m1vWWinwDRzGkPWfrd9+FN446n57KyD0OW68I9Il9K
ZEnGgvt7xHOQSHpX2n0V9YTEok4B3IBdssuR4UWK8Nv/lBQXYG1+qu5Tbk8j
NNYDnYhoVXIxDRQYJc2WCnymoor27sQnMwoh7+BQva1o3vhb72KXrMvUwi0b
LE3B6hz5VhIWlfJ73vGjBN/LrlLwbBLsSfkqkeSO/T0QT2nuCIrM1xHMjPFI
uVzFId7WZ4Trt4iGr7oyKOZvvKUKnIpk4KD7mNN35wW5MxeBKWpEpItKfCqA
PBlmflb3twnhF/++9jTfG2DFtICb+QtEZhlsIr6QNPUIxVpLaMHAL1bNIZrY
CrnZ9Fs76fk9ltOwcnR6nB07Om8L7UqSKEsswQeVYl14GJJRjwvhoAkhIVRk
cGZCbHMJdEL0nJa2MtaB+/Ueoi3VVE5t73InR+rJEZPuygMYP1/opI6qGxRj
09754+oxLRLqex+AeCYXCp5bkXhNfgKbJGsrxxHctfQ+3qlYRYRSO8exDfJ6
2hwP7V6ipaAMYM0cLuXdDO4m5bFklTKge6NPtVqY/kz/Ufg1+u5N/L5DBMrm
gKGEn+lHfoalZQfzrm792kMephMvBBV/RC2ypP71hogSWnMUoiY2A/07lwMG
763Nm1xOSGipHg6aZOY0P0C4F58deeOf+QppdOB6N7Nctr/rlybXpskQC0bh
9hJ9rEMjvtnZjbE7z109x6pOyvKEqcrTZ+v6ehg8/znqkYNrppg2Gza/c1P8
uP1+E4dcmhTnAl3pLVhmlfOBR574t62YSnxX5skS21CMuZZrBa/XyUIbLedD
yHwdu4YlVoDmgX5jgog02kZwvCcjrFclRdthLy5IX/i8M7UHI95niCBqLmiM
uVZUknGInuOVBTDLXysECedhChZFpV3rEw/kcATVxRyzjeq97fwffSNUH+BA
Hu/MQAtwMBvThAvJ2M9zDhltZMUN7CI56EO5/VcM86sVMzafbHOfCOroF4pQ
F2itjVqkpuL8bEJ7G4l3khZ3B6BcL3QDZ0s54EA8foxq2ywdLWTJwEMbF9UL
0xm4ooAoSgvs/yC4wDyOg+kuhFcdKFG8Y91GBfEBzxldqMvV00sc8EQfQYg9
WFKQvFn0QZ96GRHrxbff8LA8E9ffrOmtdMkEInmXNclEHX/VTCTWsEBCYeFU
pSP5g9Diqu481lufbgmSjcq4OND7uBErY7HDgLukTm2SYFnw3XZqwzvVV9oH
sFQa+lbBwnT0DTe3a3CMakKKJ5y11mwR7d5FD5wlMtsY5BS5IkSwDL0Iyzy3
0zVYvq+UB9DOAF7nzzvllS4KlPHBnuxvOFiRfBJuS9wJFTZS22k9uEfG5qli
kMvdMrHTHt628bTiKbSfbagmDIci5gy0OH1A7RjGjD3yRX9vhwlzruXbzXZm
wN291Xa3uCqs8kOWMpCWyG64kj7gaSe3/LMkkR3vx1W4QNTFvlfKTaljglRA
EkJT7yNMTRSTVPM4uRDAQ+xure8T2ek+2m2L8l3c0RcB+yaCMyUex/8t6qwj
ModlXnYgy6lBj1fhwEZDpfgu+3g0mNlPT9xDZk1aHm7YBqJrZPyTHDrR3gqX
B8z/W5lK9/AfT+XaCxPR5PhEfVGdP38l4MHg8HCjK3/1ADC9YPTJAES6jVZO
FF8RIF1tEHoPYIx2wAzaX3jM86X0B45L/3tWVGuNyhj1mYo+GvkHgtjtSbXG
3sWXOhlsrlYXQUsMwzFS5rHJm+IQ/JgymQ82i1/LKZBo6S27hBJTWeE+GQ10
uGSdMWRpILPp+koaJ50rU4LXQRv9+fvhpnNOll4obdmHLJkunG/k5ZTJGrgH
WYnEDsSA9k2gnTrQAgpsvZmeQmQvDnLgcCLvZA1VCCDxO/T+mRb4akyaNngr
s5vvFQBBFIoxNdw05uNjSOjn6YrEX7h3ISakdmQxcBgUtJcjtoE9L3je/MUC
dLBg9b93aCtZ3aoae+uaJnwdZ8zmAQngG1jhUcv7TpNrq37uxczeIx8RALrl
Icp/GrqWT88LXsWPH2I48IgbblGMp5XPAuffS5PlevCyuKkIwRf7wWnL/iDl
IwnjvAegNAnOEb3RjOeuHWtiMeoXc7QKalwbJaqjCgjKfBaYL6kgwChseLHK
1V0Fl0qAFVPIWPInTJywsbx9DQbEkM8e997RsaIKF326gTFObWf13tDTJYQP
X5EW4oMHGIJQoD/90Q6MyhNMxVNXZ+3vbjd9Tsz00ctjFQS00wYBL9vAFKN4
dHH92W8P+249DGnQfdyHo4VQZG9/q2rq4ut8Ll+Lhz4/oodJPZ1O2k8pgBb9
qrWgqm2dWoJXFX3VIhZGeNYShpCtw7NemTcDDnQrn++fynXTt2K4JcZSK/91
wxUzlmmmuaw20w4SXJ6uWP4wBzkKcPrRlnwonqLqiz6ocqg9/2o/IW8BoM0r
K+uEG2rIcd22a6kCPA1GxWknD9g1TAeh/JHBQrK2s52gD8hQ0+ToUpONYpz1
ENBM28ynqEvJ+j39zqupxk7WxavvUnOJZ06QeCEaPUJjelNuNzElxf82qhrH
fydSfisAH8QwBU5GByW2pMlGnISXYJ8cZLOT+GOqQvrVjtwWVDDZNuEJjzf5
fDpxwJCkoyG7H7hC98hXVCrD4NHPsvjlOg/1Ednd6t7hAQkQZMgfLxBO0Psz
fKOi3mzW9I2+PRREv1F/9+KHqf0Icw8UoP8SZsi2vRARxjME0VfSN+rfE1vd
V6lZnODenqo3KZRVWZExdxrzj6YY/K+x0UydEl53A8qFhGUURFg6FiKmlImx
kX2pKzbfQEiw6xU5XrqFmBwpap5dNgpT6dxT5RfYd0xUQWYijK1OIsPMBl6x
le0uh1Ua4nhqDExb9Sd9d447GitBA3VaqkAvDccRkxiw2vLOwp/HJiAQo9Pi
/USaN1ydKmbcoUr4CTMmbYeDZPUgqb25YY58LbC860DbLMUr8MgdQQxTpjM3
eEKa2w2dTpc0THwkZXmzvcCbekhdtC8hQ+/D/seAQUK29sdBEnGbS+/DND86
/2TjTSJQiJ3bIE6CVnrlpvAmJFUhsZLJ3+23p9VcfIHVR2O17WF5oPtTdae+
/+vSjmCQc2uU7iC81Avd6d4MMlzDxkE1g3c6hZ37iYhtXiXBxOPgaqWJTYF9
Cc5lj9MP9gu4H1yTfk9T7PSk013q+S3NM8MP3ZpDOgFGyHEl85yD3/LvXwqK
23XRvbiflcEv5PYmzbsk52wNvHCtHgYrFU7FpIiQO+PCHMf6xCf4dCxlX01/
o4GTViQDhHUgY9Nxz6E7XFZ14ITizJAJofypnoIKGC5FXE87dmuQYKjgS1uM
4ooMYV/0FVn6KUDJq8jMnv3o59DGysL6P+pO8KEO0LJmRRRniVBfVQjd75nZ
Xq3fs+rluqEq8OYrjferflrecUou1ETaKyF+A1lWBFQ/7qkUhch8V/WDcHg+
zFe+CjxFkrxg26yjFKDpI60HoVmY34gVG2h7oFQQgKLrvtqLwMHYYnqgWGlS
IiCtkWgtXK2OEeoqGFMeGhfFEMg44V+WQEfKrTlMlOpVHKck5NcIeawdzOAT
RY24KoKwQU3LPDnlWNncDjeQFg5Ai9u0bWdAYePFquu3WSA+qoHZHZ7BEMgV
s4s8cgCTCvmRwBO96eIqnD4ChVH9vFEYYwl+DjaZGL3pCTwJTM1ZYc/iUJqc
fBDT49G8pK5ntzmSC6lXGLWWC4ewon6A1ur42diYpWQ8SMoEQl1BzfU+kQhj
3k5uUG+WNuZ7e1ojbzeozok5+QcHNqm85aRwV2qzjwJjkTqjyYgpXXQxLaxq
YU9AYBpslsc0zf8lihTTr06NHKV+IaAXinCDA04JW5oIqp0ulrIo0rVDPoZF
mzg1dKwEtqHr+mU/V7FQ45ViK6MiieEIJnoNP8uhq6X5700ERlee1uCBOK6t
J0vRcPimuNmv6XJVlTMEzt7EBo0xMD0tTQMgq4yYGJmpzjZUDkya+PL20ktk
kgW8ALkZj7hKjuFBXpk4BFtUXDVc1ZqbsICF4q55ncu/cRmTdvKljNKtnxzf
HABaocD2Wzfn78q+4nDZx+ql12zZND2gaqITsoP4FGi/4m60lWvfBtyEX5mY
U4+t9+xUiy/sucGWXJVgbylR6/YKMkFslFn9FHrXvnCPTyz5DMXamtLAZmf0
Tsey8FKvAYpW84HsJHG7PbhjRuGoWqfTr5xFVZerU4WRus9elFvIlfnHkSy7
EGypwlImRa3oqqiXCqAtYGdUTG0Y2bm4pfRXZTa8/Fo/b9SEL13UYjhG8xvV
e3KSTyufcIPHQoainvzyxwfZsH7HtwNTgYGaWxefino683V+AQIB8IQLlGtd
Mh2LuNd4FppNKkj/SfVciV7JcBg7gd8Kyd2pdWfXcC9MMirdXrgg+7CvORA+
tj97zsO5AzCzU9b2HCDrG73b66/5Fuw66dGZI6SY35D/G+ThPdaD5MCiXANf
3URk9OUfMmnbeR9FioN8pq1UjXQyOLbEPIpUsktVN+k2o01WvED3GeEEjkA5
ZWtQaQgzxrMm/ekjlZqBU9hKWs47nAbUN9ohOYsLyVUw5j18McxqOEGGfffd
qwy+HDV4QvBUCgaf8JfUPU1CUHit/xOxpcNFJCYLU28PBZJBL8yAD7eqXRxS
ROAP0Nn0MkQP7okzDUP/oT4o7R0MMeflFlL99WVuXE/sHPChLbd5QOZDe4+R
7YbdwpY0dLBDfDrNBNAhkV5/tKrZFdvdkHFY54RIucNKL+z/efT3W6zwOYRB
WfG0GquXOV2wWXZGTZYmwMP33kVMcpfgldFIY+s5U2bajF4G2MF87uBvXNX9
Isc/U0t9wvKrscZfCtN8LUv4sVE6JFrOUNPE9yIst67IrynALGOU01OL2UQx
AKuzDybMx7SHSqpxyzOvoms/kl8cXw2phqwCD8mOZFOJYeU6bjnxUyDmtb/k
j5N47kuQRxyq4PWHZ+hYFHZlE6qevV+8vCSQepythdyPUyB9SzEZ826pD1a1
0plRxsdmG4PSktmOtz5jwnE2cvl/WrmsJtB6cWTwWRvahfrvWcOcqly7qD6d
VyyWAEWlZ9CcnwiMZBgLC4aEXjWzN+kMT9AILIuXPCJxpgjCCcFMz9mHL7CS
HD2R8YoskQPVg5ubVG2asRxi3ZhXMcZBd6tDuVXVZ6AAPHQmFZktuepuDlRM
nNmoESl0ahSdI1vXIpNU/io5DCEY2Ir2C2CYriczXWuzq30WjJK1Pnf2///F
zO1taLgOeGtHiJEGmeVIdZ3SaaWCkOexiJ0sTcHfxuSzJtcZLzF68Ag/Ca8I
9xuRtpSZoVMv32GXHR90UzckD6tlimqZjLIiW2ot2Sv0nkzlBT+RIU/6fXwy
EFAzsAZLGHqe6O7CWsgM/5WNMIvgBYpsdffRKcixd2aQRXuveNGcrSWNgoYw
WFwPZkQJTfMdfwAu8O6c+Op1rsH9UWB8DB0hw+TCJVIoOXapKhsCBn9usS0u
j41oOHhxIBsmBV9KrlV9+Y6DXir514wTHFxI/P7bLHj5Qk+nyZxaXdj/9MS5
n8HcNjLK35u5ceGq2PL7UKIUSTZYCcDOvEVR4nSXi+YNB8H8IC9SAAzbQdZf
u1Y+3q1pI2sIRXz8uA1ggqCc8re2yURR96NT33M4gcw/Rg3NPVQNfXGULb1P
hWwBjSIcU8Fp0nZYA/idtnji+1IS8u1djEojxjLzEQ5rbWEp5HdH6m1KmrV7
xX/9971vhsWuwzWoohdG1WB2rTCy7pycTt6ePNDRHZcWTa5NimPA8TK8LW+8
hfRR7pxeLAR5xHqymWUUlQCcxqk+BzJt6ts5WQXQaLUWxMfpgcs6BDChYV2G
2Zw1FPiZI7Zlh00eWiOUcIxuHE+2AV6TzzzebDpkI5njQpGcMIuQYRAeXD1P
JNKURpi0wZ4SUoI6k9TVF+Z4rBeeDSAnkYR6GV9Oi+L6x56AhTLn6Z6ERsdf
233ePnxPXZApUi5HZXTQtyors9vZOz28bsTw8+tFOD4OPsXhwQRxMZEcpUuK
Krsk6MFv1srcXrD8FcR6FlWG8LAqqezgm4yw4bhDlgtjcloQvjHll6wm1ppD
SMzzqyY2SvlfkO8o2ezEqN/TF+1WjnHqgu9NjPYazg87HRJXYDThCjQOPXId
Z2UcdnZc4e8Dwz8L4ZvB50lVSLQxDv5bvm0nNMKdCTSrbNpZ0k1KeLCXR2B3
VwxfSc26p+P5uFS0JU4eESIFtPapGIayn4SKP5JR6CeFMjtK5st9ea2vJqP0
WComM+2fjqm9UROETHD53ydPxKpiQxm/ovLKCNLmTJSHKIl4P/sF3L7sUwN4
gYcIZjpZbroHWXRKrGXIF5a5V13/mGoW8fMowsckuYXETdLmOVe3E9cn2CFz
hxQJzJUmGIVeBbr5t2ozb6e66TZrfkYim9fzn82fQMtI4Dqxc/s1LY7QRLPI
CuQUrDpjdJ/JlmZBY6dQerrHgf5JSRYrTWr4rZtrqu1IkS7jjye5sTBSuvEn
DWduFIxo/5w8l3CTr2aBmiOgKn0JUWyZ/TazyOYGowR6Mzko/nC0bU0jqse3
eQndgLePSe2+GaOPqQ8QZF3sCkUaOv+pePleWaI62jnOe8njE06LBvVq66Fn
/8ciyVKTpToqZhooTCyo169k3IrWXCBsh9wqwmlYu8p317wEg6eS5bIRX2Gb
vuUj/SSbsvAWyG+oCVutT1o+Q3dDVaRCt/vrA++AQlhEvuh6ZwfFhk84KINO
YsBWAm+IusTAVWeTlyqm8QQs/wa7aYEh4vya3661qGJzjmv8jOhM0mREbAvZ
R/iIVCFyk+9JW6Z7hSwiq2sckcP19U+d9pLifQ20KC4XDgEsDCUDNrZBQNj0
7rIensTmw6yACN7jy8R71aBexk77nmfF/UF34uJE96wuqfV1ywclLt7jIkPn
WYQREy6DT9WY6i7s7n+74gudsjD1BZ2w9EbKiPBa9UdhCRbPSsghj3Y4bJsa
GIhAwl35e/JpAde8QJS88rhSmpkxOBVu8RsxD4HzSa6xXIWgYGZyzgc5iiFl
fmifSZe7Rdzp71pWvmK7uvYB+fkMuS0VrRhCnuKPusL9ooZaOfBL7Fo2bPJI
QowWkKeO9IRtb0afwm5JIF1wJ8ObjtUkJGZzuzFtm4H+bS8h6jTrENdKNrll
4urFBAvTXvo33Nsw5GCZIoF+F+bKMF9bkrlvg26QqEJVTvcEbBw1cj70eSBf
1uq8SGioa7Y7YGaLwmxM6gwmXCXRHDO2U06nfcSd2ltYuPQhnaYI0e02x+x1
XhoZLUnNfTDqM8P46b8mCPuqLwQzaoawFWubc8XUJqk3AkR0GSDcpucXJUhJ
C6KqdXnqYVpPzdqlMl2ka/BGzjedlB7Ix43cGmHRfoNMrxJ0m8SwEydipM22
bkoca6LQoz3+xoHo+RtyaOzb+Xu+THzn8FIweW8cLAmt27yYzB/boIRC4lCO
oAottaaF9CI2RyaJnn9zaEX8utgPaz6gpoz8QPktYjTu2Hve4h0uK0uVuPP5
T7b8A1J2udsE+lIWs+XhGIS/D8L9b0Q9PxOyLbQ3Zq8xMb57Qnx0yYhJXv4n
kwHf7xK83t9ud7N4UmwxNlqn4JHLcod28Sf+R3f10vYXi1TpIFvECg68wdBW
luRvpNTQUQmT3GdCN2HbwXwAp/itLCNqkJNFZ3CiV3SxA2B2YSGcrljaWIPo
1cruRFHpeRzmr8uE9k3jdEVxiWndrBTz81QI7pvOMo5m8LDgYCbZgW8Wu6Ch
voSEFkXmZNVhXqUuXSHSfpGXexoOkuT2T9kSsz/mtX/Szi7FPoobjTqkHwWI
Iwmsz7uK3Gd1H1+12u+P047aUvA1ePC9MMDA3ehhdxVngZNp6NpbMVonP0Ci
tk5fnKj4+bHwpJUBfcohTFrc4ItQMOsg3RrF1YzeyuzKoi8xQoTqi9bxh5UU
oJyVMKsSDJL84wk0xV8+n6HtrVoi6MJ/SSS3u+1asTROGoYuOqiQLSyRlimU
GCUiF0Ti7zTkjhkWDaTWc0NtJPLYQlJedbZzKDcc0X6vp4c2me5xbf1fRj06
Zf3RVad3oBrPYrXlJt5yjBIxIfCPkbuRQ3o+UziAR88u+RsOjLSRT1bUe/Sp
rFf3hsoYhElCbQZmlaTkQE2Sk6zMbjjClAvYQjomvo1EIEqh6w8waexjmGHg
u80KOspcp4MU03t8MlBbfV/iJFXOD93cJytGItny7q8deZHPt56v7YOOBvWA
MX5E+2Wuyd0eJcFVQAAqjiBCy32+04Jw1YzxxgRzdYPE2ykOTN9Ck5W223lr
9AYn58DGK8Fpz8MgUt72pq1hakpo3B1ueY0dHrFfxuoVT+rnYTRenhpzCZFr
n5QNcSXxRj3jIknfLhnfbmjz79zbusIytcCfZSUURXyEqie4fKQsy6d/sVOX
DH4ohu1gDD/T4yFDcko64Uf/OwyqYpH3FuaJDoyxIsCnkyZIUVTcBxZGSDSS
Q8KPnIXJ0VTKC3pHaeooNrolWEB05bpvb22kghLpMMPCgkhJKzF+bXr6c3w4
1zUFi0oroud9ay8I+FMJ1evx010hd4CH8CaJtVgebtJ8XK8bjdTV3NWXGl1k
aXvuC+LlQ+X633pBP9qfd7hfDTzYSqtmXih3NDf+rFdlqfjOvoxPpbYMBYYb
GX0zosLtqpEwpdqeLdWEFuiI1X/p3cTlyQcTNcDU0fpN/vkWF5dp4cOevKHv
G/xT/kNCtJH7ybFjlPt1aVLymDWgjpYG88OF5dqHywu1U2FBBA+RNnIAevGk
neVhfLX3SjQVu0fpVEQ/gHm/dWgvpwcgTLu2cyv2kN7B6sy84En8cTfGdSIv
Z7MJciaKA3vwPBNwohdBv04th4tUYMC9Ivs+hFU1e/nyCSNeZSbxan+q5r94
56JuILTBbAguCNxHJhCVsOSlCa56pDOjpuTDejcs5ir05WgoTQ1aphtAw0OS
74GTDzga2JWXX74Iu9QwIxRMpVYZ998/s3kF69wT6yMvCrmG0L+HY49hXSiO
G+esn5vTjgeBUxVVgAu0NB41aY89qyo6Gc0/YN5UuUtbnwzInCI0MsBrSKF/
9eZSu3ibIs2w8h+iFJMBlJiGROwjRO/A1kpMlsZYvehv4GdlP9NjMfrrMY5L
T23G9C2Rh7ACFRnxlSEQZldAJ1MaKdTEvox2jfbty6jIPwY2aK44iK/Wiarq
lke5rIa35ffSy6R5tWFELdBNlHOIUIPWle4X7HDBUgeDnbodAg7IO2CGtXZB
VI0dCLCTf4hONcxLEthxKUn3vueWE1JVvDKjsfIR2bPTZiMKkEDhwvFuGwAq
iIZKUqLa6uTNRKPvbjbjIr1VOl2l7A5hC5WAa2JVAFk0zmCGpJHL2XMZVZc2
03e3Im0wjiVwTfOlcgx80JIZ//9nVubCOF65Ep9/VScGq/BFt0Sy0TRX1Bnq
T9sjStvYMcsCO/lRkQ2AcnA2JPrihl1WAspY0hxeCOA5XMbnA2Q/WKHvP6Bw
UCav9Q3f+b8b0CPos8r5unUGKvSatfOWnSMYC5fRrbUMpJQZnIM1Xcae1JLN
T3vNSSTuSAQYCc4BVFKeFb+JYk3N3acFFJg8R1Q6E47BPvMgSiaKMaJk5eht
W8CIWSJfG9shFdQjQ7B2oaCo39BM2bI200ALoozB1HJzE94qcKpTlq+iVfFg
WVGGDIlT77EHt+O1gAe7TYN2jqU/KYIpkZOcH9AHGBF732aNlsgKz3tBdg5s
IjyVHn40nLxkvm5HqlKJA0oMJa/62pBGDS/VUQuW0ig0JqkWKsH9krkIHDS/
QBd4WHmjYMPCorI95ZFBn/RI99u6kLIazkxvtlcDrhhYjwLx0Ug11IIv+Tsr
bfMz4spn7D65bzryuP/s8g+27MC1OIpgTPTR3rVjdZ8F+BoejhIQrSLlLr8e
5zwubuBk6VW9NpiByuPlX30vSl80h2sE29Koy1c2ClJ/QIoho9JSWhOyhVoa
BjuSJBOR9mmNQ0T71XV8fp0gBCAr7rNujw+VJgfCj6BlYGeqGD/5BwP989Qe
o0mjDvJtWqxvBa2gdO59vKmw8fc5akPusN+hywp5rIPkm6AxTgXfcPb22q3l
7BSsFIoDpzch1cn7gEOjqjiusA96mpmQhBmr5HDmTLFptXJv4B6F4468PsGM
N+jNP9OhERVL8oPLndIKZ3besG8HjxZghSvRK4h4UzGphMGf8V+7Gg4BKGei
OaIWE7kahJtbPrm2IjX0SQSXvZAHY9dm5rY4hKxy8HDZpWo8M6XBRWHc7G0m
fSk43ooc88Wc9LlJeSsY07VhMa3Ytbe/yamR14AwduPuxNgkmrQDlZ6GTQpR
U0i+HU0VOi/LjVlwHW2pAWbu2Jdy/N4YwLjqQKJc6B/aq9uE33zWggu2+ITe
K4Vxm2IEO2YAV+JjPy/pFqpl/rxH79+Zrwl5CzQF2MbohZm+pQWVS6zVILIV
L6YuitfuGZ8mVmwxBsRIK7QeKt29X0gx04iwoCpkKW5XpFEKKmDy9RfHSyot
7QQPWqZjkp8c2jfDoidM5yHSp6e8ms2maQ9J7vgirpj99wv9r+d5JxOJ3i0c
1bTtYPrGi4cISCNKwmundeT50YLJiqMC4/5QLZae8upxmcIT8iqUa/msxhdj
tp6yZsbBNIDpZyEM7wW5YKkJ/KFhh5caTf+EVA+KIirkMZFbUxJgyJDz1icW
BkMW0/2hZyw32po793t/5YuzgLMAKgMGcDSfwhjCcWh9YyfjSLmwwJSDu6Ds
0zZ1N3kmwpcv9w4budZ/jzB1DZJYnOqH7B/Y9z+a8Nw0UkhmR0YJPOTo7UDz
DnOluRqXgE2TMD51Kb41gAJ9NAAqdSQ7S40q7lGOpDdaQxvzAo6RJyWinrP8
bqw/v+IOls0ZJpprbVZg9HAGBxp+Z0G1Wpc3O3ft1HHh6P1psWzqFBNFWYDf
TMJCLaxR7cyoGTTRXeAIzTASihx9gKVKfINhWu8VpH35fjetfbZjRZFr64sK
1U4AlhvZ4y4yfaha6DBd9a7SQ0Y7UkHaYUxad4MYnd27wZPGIEns3M2pZ2Br
n4nV/w0HBn9FiJ4rn3YruO/AaRH11l301g/tT1VZ57UIE77wYWDmSUbQpTJB
CD5QIqabvA43iJdCiXV5KbW8GSKEnM8s7AFsfKzx2nBLguKiql3aItrQ91oQ
4r845tZ0hEKUAjdlFa1EQvaGC1AxcMQdD8RusobolthJdTz7le4rnXbWHfe0
nSwU36CNqFjq3lndeeGtRfW+sPUrvY9dfxEj+kia7dcX48lNccukuycJqL4A
gCqXxAVV6J60unqJem+yC1wtgDE/vBi8IG66MfiA3THYT/BR4MCtezvMQgsl
skBwxAZqgdzNUGDeCxMFB1yxiVUAZUNVD9Kz9Sav8ChyJB4jAPvkcNcJUWmm
li2UrE4fbuK0Z+p/wa/OW3ByrEkfcZTQYEw795IO/jOqX+BTJvIWu2KzQ9NC
/34t8t2V+Nz2k1Bc4Pr0bBgzVIapTcSwqaRi6fW5/ccB0soc1CD/dOd302JT
y5+u+aNdNFKOFncTFlYG8ElwnhmKJ7uKNDHiWFt0o6F6dzO735VNHqYbsYVi
AoPaCA2nEBMJO8sFAIqWLC6XQ7T9g8tAbavAiTVN1BMXxZ7ntl1alXo/boce
hmt58NVTmOEHDZJ0eJsIWMP7JQGxnDeJzs98kMulm6wwmfSiT6rCNiYvF/n2
93U+yVQ//jqvXXG1rdQ9/1cnWWVnSVPbe217/9gKLvzjVou47F6hvyy/NkiG
xy1iJhSLgveUfpcmKhC3Ho0VTDsFGkDluitCB5pomUpHZEr2dUVYzui4NlIp
21gPUbCCOqjAslZjVLHw1Kg3o2XF0rEPn3IuAMr1kbo4ulc836FbOxxiICIc
WMFI5NShLGEoBmsjY1P2go3xkrvZutTgxOVPuyg2/fda9Ga9nnOgyGsXOKx+
FeoHsJanETfuuv8S/Vlf1c9z1sujtDHMiCwyWB7MRASqxUmMFH1pq++C722v
nrJVBDc3hKs17F6R/Niix6/CBAJM7ETS8pnLOxgR/UzzhhRAFVUaRA+ZG9G8
UlMGoIAbAKgtOCN9E6NLDhUglDwmgfT/fSG0FO9HuFTMAJ5w8fJjGhnkgT6E
4nVy5LCP6RQSDIo7bkWhXaKg+q7vrAS6+QxNKlvxTXefVIBaXd6i373RyxQg
eo2lOu/oIjVGPdTjxqWpOGekFKC3mkermhEeXkeBQed2or15hPS+qXkWDSn4
Mz+gRrwBxr8nDCUUP+RskfTv/PiFsmp48dxcqQel8I6MhweLbzfg6qg8KPya
ahrulnBWLN30DftYES/QMm6DmYbp2ckm9aGkiu0p6eJi36R6BbEhns+Onndq
coFYahbGOAYRHjUM2HK0kFvGfqQCvPdkiqXqp3FeR5eCMTFfbCMsHLrmh8/r
3eiPGOKDWexun25loYHLjXU1hbGxJLbvQhitqN7g1ncgRCoELatCLKC2MLUX
tUPJVD35YwCNHfIDZ/awk4mrkF2rmfjdY+1x2wlaON9/5Il2PZL4jm3cPLA3
HemnnPUmUPtj34DJw1ysrM8Hpp69SALn60VnD1+rAUwZyhg36Oe5/i5IvXMB
CfJl34N5hqKBDIu0FFkNJ3hplv9L4qXtDu3QyaZ0c6MlnnRjmHFv9VobFCGo
TnfSZurC4UYbN5fYF+IbFVvKEcJqzEf6Qna3dZxy2krg8Bln2A3ftFVyq5sb
+I/9djNDY1AOGECMeLLZgh+sOcUZC/ihXeY8P6/EANxyjeiszYq2ufLQxNL4
YIj8nsIq6uufU2+q6pO8Ok2A5p/SPvJC01Nhmmzq1rl96FMmDt+IJzVwMnCy
KM30ooeT45UhCFoN4fXyPbSoD8aGthh0ioT6XqEAkHsjW+AqtHJ8Lsl1H7Pr
rAmBIjCobPPVKqca0sOEXG1SAIZ8sXZ+I8SjzVOn/N5/cYdGge6JRFOceXhg
oiSBy4IHCKDUY97NEKwnt0HqlFLT9N67T9SjKpsKtwXWZbtWJdh8c5Z/ART0
Rbb/EgLkYqC06npg3wy1OjprXCLIXnuXzElNMS5+73cUfTRu8m6IYvijxp1E
PJJipX1fJLN0rBxjgfdKfXOFc8gzU/UJ5YkaaV2oU9fXegb9oEr5/zVO29Ol
nuWR84WVAZ/gANh10wtXHnsqzGHZx/Ht4p0cBdMX24P8N/d3ttS4alB2amCS
PAERVmUNqexdwXqQ2lww0pDEUe8/Wppi00de3DDBiQmx81rqMY/DXRH/ciQ8
+7nk9i0grNDKenkiMk6SIX1knzXqZfbG2ezaT+CpNVfkF0yhXWLkBM1z4FhX
BdaJOTvbpbirRpHiiALZFt31F9El0POj/pI+qvApLnpDXVH8R+qSTQXOjKay
HIirbBEsjKV/USg9/PFDxGM4vEVVWCU2jnObbewUADPnCWVR3Sp3W8be3ugO
AHIsOAVeHVIwA7X3jo4NeAvBXVRYDbnl71/3McYy6NilQ1AZDjnQc5aF8pPj
K3X9oA4avN9XKt6qUBxTCJmClTq4wHtZodlcM/TRr3PolGv1RTMqdeJzLfPy
cE8UQ9rLIS1LVdpL4lYDXfNX8dn0emH0cb0AUYrwZJ9dt+38eO6VHAM2zhDl
kc+qfevvW13ViBDAHpTXt9tJz6OxtHy+zxw+iMDWqF2gXbjX5GOzaes5IRdL
KpqslIPXMmmComlRMBARWVcM7OtJVGO8Ae6GTne0mNvNSSQaoFINGDsFLNax
f6Kk+i8jCP5djl+ZgKQzEpMip37P51UU/uSmCBQXNEXkTXifsSRekMpohSvp
pu9jMLnAjyUn6/f4uHOTvihzDA0GDxFdVM7+uKJSLycrWdVA718JxG8Pl9fI
aBPh8Y4yO1wV3EATRalDxBFjie2TMTef/J5Vbn0uG5ukj8uj4PlAYUfdmIHJ
BEy26tasZOISnK0iioKN3wBhgd7QUhKEOGgkbswZNjzzWPBmjXSiMnVDQ+ZH
DLP3TMX+ns8jMmvLn8fHHSh1EGDwIoutLZtfN4J6eO/kSpkKOicGHTQi83HY
60tHjgulSQhVEY9/BM273cHRF+HO/QKZLC2oF6NeVqQGVgrtmIbop1wEifes
X4ub24ZPWsyPsWiGxWyvhHAxUp9MQJOWFngQ23QT6Eo3VIYDS9O3Z/C0F0Nv
3ucYeyAvwmgPTqo3zi614a4PlGn1aRDavuq5TZgCRB0jtxUi9QYwvtjkaT53
tQROu6H3iDhAgUK/ZJmz+aaLA8TKEeMqdNPkV8ux5xGSDIQpSPMryfyHutOV
XIcZfRn9Atr8YNJS1jTyJL1NJnmC5IHC0w4r4FxReUTp15qX1pzrfcAPdWjZ
XvN7oianfE7+liP0iWeM2bdUVHV9zoT3UHfF1dvhLJX1GRqVfPLcWXZqb+q6
BZ6+3+efZdaBkvXjudBcDTc1utGO56kY6aLK5lwDPiLdHtV8MD9fkM8jj7/4
ptYpFh+meIpGdX/yjlis3BsGmFH70LW9RQ37FqFteBfuoOWOMsx7EVgWcJvK
CokmhoPtaRfH3WX7dy0IxtqDFo9lJdVO9bpAJCb4y+uJhVwOqfNBngmdq0yl
k5TC0+FEy7aSLtjKarLPj15LOAxrkG3d9KFCCFEpayp50lD56ZliHAvcwfC/
kHe4a6fgCuICnNnH/gVY3mSNg4Q1Gne0H8c4OwuQTNtlRMo7GNtS8gNikKL+
gCeKbvG1HrA2e2kVldOF0jkhyyPiX+jyKybHWQuF7943yXMJQz68+t1/lZ5w
rKRXj3sd25V71NmGVQfnFZ8zWvLDMQQ0lGZelw26l/9kzWDkoC+N7MhT6YOw
scvsqM3Bif9unA+s+EZzhH1nEzscoJqRoTGZqJ8EL970ZPdxpMtnTr02Ys/Y
YxGa/+MwX4VJEcfJWkmZgpJFzvV5gddU+Q2vevM4WoQxsc5fjLxCNAbcDmbB
hjMWcuZqB006twWeK3bvS1xZsQ1ZpoTSmSBhw4PMOnzJSu3TXFz7+HeE2WPL
p4mfYbakCUxucEtBDo0FpKvHwTgIsBETdH2L+wzpeGWykB6dZuKJ8HWhcNUj
U396qkD2n54V87KGLXrGdrugodEFdjqlKwiFYnG9SdFrZP+5FJiZiKEPvh4y
5VpA94lqEkHVHK9BZHU15IvDxp5ZcDGrqRBjsjU54btBPtN6rkepuPqsScuj
fE+zRDbc6tEdRS4BYWkBaiX9sBMcVf5ji/MYf5jF7075lpqNyFUaoZEgHdzj
0Dhu53k2iFr4arHxHrpvFdJztJ1TjfVLmA3V3rZByow081ouJJ8H73cKzYQ+
ChWk2IRIfe9tid3FXhaQUY3DGVDbafiXVuuybkahADeYJO8ovwj2LtXaqKdS
+ClbvSf9JyrhQ74LGB856VngvL7M2s2TQUrzj7yf4iaIOfACz5cHisQwUXun
ma1CKzPtcEiJQCT6FVsy0ETOYErCU2HzmOGLUYw2JkXoCkbNlot2GKhH7D9X
Vcd0RIDUc81+evGBXJtFNsVVUw2sJnFeOwkyFBkE3hD9QOMgpyZ0QKs0GK3e
0wYeM07hGGUeVxL7zBMy3ywFwV4lZDhU0JnzfKkpHGlFuYukOuT2J7w7a1iZ
9LjFDzLIx2R0WOb3tG0KtXAsMiNjCdp/lUjEsQNVSWCtLh/SIaBmAVf/ntlG
PbGV1zORP9krgmD1gTi4XsZkX4bZGIy3Ni8IF2IqZEnMr1s2wXaq01lINjg6
xR/Av+NN2v8HrgXGT4yZGY6g8nnN9C4IJ2bKixUGxuAIskpgOsZTlBEut4o9
HouttozT/3T0AgxyMk3tXQLt7XnmSUIAqhflJh8M8S60pY7MUmau5aWcIpKI
SudZSFYJ2J5RBhVaCsjzAX7tKiFLIsO+nLJHmNdupDuMSiIWaERHOIuZcPEC
KOhVVxBvUa+wzxwjoczPm5KxnW5zOAZUjO+LMRvBC9fymevs/1JTNhuDRE75
k2GrwPbzBQxfWftIDqFg9csFoGbqLse4wcOs1dt0W7McmFQ6g3fZR7kot1wo
zce3iwHv1jy/fnbDlj+XL0CXlSQDG5o9v1KTanJx7p8qKPI/ScbKXK1/LTvW
jMWmwJsrgueu6plr77O21FZZxjtzEs/Av+PA3+E1X/yxocESHK2p8afIuou3
cniIS0p4viuClVyC0u/l1fdt4UzOsVSRi16kkaC1g/V4p+jrM516uHgmLeST
7AbjPgtkfhpIS8tmOLaAQnebj4fQyUhJqgAigHYKEgVCUXKBXsG1ywIMGMmv
jYoBJXA9MhdB+6LtlYyLljGCQHt/te+2l5y8PoVpj7dEyeNoczU98vSxs8cv
3ZzYRcrKbCaaTZQfBMkOBoFPM6PKJYVePtQHxBMRxuDf+J85zvX6OYfJ291Z
YzlJl13IJut607jJhmWmBl2kulVXTLZ9SL9WvxByumNC+xYD1yivcOOYdrQV
Dkok1j0waO4cul0SoXtRCYDlbUoJnd4nvEA4l4tPl6ntfkap9oNzztBFnN01
f/4z/Y3hSBp7jh4KWiqoJskQoA7ewXE/caDJ1x3EuK9xRmIXX5HFoMS07N4A
NeUkYxD8JP5xOIhspSycwZqYkZ1qnhTHVpkeoxtz+Z8KgbYNjmpncMmMBT4G
kvq6TkisU/FKkEZNiYjeEiT68TeORmBs4tJEjlwUr1cbvRMOAEJG8KiynR36
EZRRDjM4imMCNhLmDXl7zKirre2oDJjtTLKz1Bxnz4MXjQD2hep9cui3fxcT
SIOIzwKEz6o2hujKmEPY6K5G66ZVvWH2EJJh8XD0+nfGyfSCHJ4AxdxWdYlI
TQbTzKV1PcG6yLveiC9ago8DgspgsWBJmitVxHoWDp+5DUIl1kojbQFUJOfN
UReUNMzFlhUwF6IRUn20/iNDjXXmiLpn/C8+BponnAwC8YZc1vl+4G1yeP7h
QC7i1aR8Ltl5i2Kw+ZC7Ivxtex5PnEc9E9QQiek+Tr8jdBXDRRAbP7K+jZn6
itIUuTVCuxwdBKRw94P1F/AAoeGvWGjwcdKgE+krMHAEpduK4sIdsmpnJPdU
oLPZk1gwB2OiHLNBJyuojgSoP3MKwR5dDbKpfFY7e6NoRnoRPwTiry82L3tT
0YnLrp671SQMsnWug3WM1me4kG1lWA6QQUzhT9QYbFL/PAN9mQvhzXiUbVRo
XtpX7qeWvzpZ5N06Ww3BIdYE5CoqCmz2IhfxOHzIZxq8RoSQ8WKFxxssyc46
sz724+kVrS5UyNV18Qcu9xdIExDne9aNtyuIe/F6+COdfVrK04EWDH7WBfLB
RWktp1t3O5IRQmMMrGu7YRyMo97qt2IHdWFr64tmKJsSYXIFMbfy66flQjr2
W9hJ38D4yxq4vUWRJwR3iQKm/ZN12hgBBa2L48FOkRbtCSpzhqtU2dYNdQZ/
+zHPHB6r6H9wKQMug1SQfyvIl4cePupW9xSGZHuZGQH21OEQqVwVHa6iv/tv
hKgYv1+2er9P8HFxgSkRh9CxEfC1+7ialeDP0gBQRxi233Aj1HEXu5BVhJl+
zLA1o+6Knr9LKpkViGlSYFVismeSdf3xgWnpJdxzv52XSq3wajNFKLicMGIF
a9TabOk3SdSlGb+E+G3db8xmqmX6wOzk+OgG0RnVQybqCWYb98gQ8x8B48nL
iLsa+aGk5DEmRmrZ+nnusbgRwvHcEj987dA7T9ezWBtwhwT4L2vxpu6mXt6/
1OD6RO9mFMUkhx6oJnLiqFzVqrCwQEwTXAUyYh9YVTaQcHJXxTw0qPaZLl4V
o8bOSQH3VOi1eYH+kFOPMvvMpMfqRJWRxAKbN+kmhDchTgxN83TGcsIN2Xb9
ROBEKa4Z598tBdPQzzqJILfZGhrjwT//7QDHGTvHGEdJqtSm+8tk+gy9q7D5
xgAGmgp5WlkEKPMByjuHbV7oAVzSBkyTGxIWGrSyjBNmVL9n4KgyMiUUHATS
Onez7YP13lAtgrjoPPuoxbGFxu51OwmGoylg3k9qMSiMw1qnxaxDPWZPzT6T
FodoGti5qqbi+j52QLfIVZkhxGZ7KeIq1oX2KZmX4XQwOuxQvBX6aezmDoUX
GrP4Gxs47/iMkQlemewNLxPZ9lhaTII8y34KVmN0fF/0I3oVkhxtBI6DJGbT
plEVAUYvkUwy4iHp6dOc2ebt+Jd9F6yZ4kmTzfYt6XPX9qIU0a9q2lSE4H9/
iyJE6Jmk8irAaTMmBfQtdCKXcP4+PDwgbAwDdRzuKe6hIbv8PMVWhzoX8/+v
WAXbrP3hS/2SDids0s4SIZNm8biFYs9rqsNyrvy5afTXLSflzVuia1LWZkFn
fg2mZxrzOT6Kd+w5VodKgKbEZ+IzmaYvYxWfCsF3nc1gXhvvzDqqyHGk4D+V
MBKBPi3qqPUpciWl1yGIslo6LMPsiTuhoK/m1RTYCt5KZdeh6CSiHxutWoNb
Ks040IoUWoX0XLkLPswAhBv3haUFhUa8mQ++vnbAojlBAG+UJgMqmABtzaQ2
ZflFbIxKNtA/tYRhfFtoQHrJ/H6RK4gPSlyrrHsjOk+TWyrS8n1MyFdVYmIe
dzehS5+YViTv0sKSIgOqPnepZMJW8ObR/UDCf+nECwqxSEzvpqOHpRGr+KQG
CM7gq3Y4XFOEtbSZFdpZv92jm5UEqVKgFbJAu4xSZ5s4+25Ok5GZFS50rvsH
lbhPalbcGo/8zpz1biQ8ZW79mF2ht3XW/DEDzOHZtJ/y0hQeF3nJoyS43vSQ
UNsZ+7PaZPFBSabGC9+M6x2Tb8UfkFd5vfAol4gYVPUYM9MYw0m293gSVHDE
5ZCzk4w54Z2bx5s8SsAIWsCx6llGunu+volj9b0gLBmVQNMEWnmcCGIrJVSS
2+d5xk9vBVSnqN/2/Owb9gqKSPc0i50KW8T+KB2n68QJ8o5/sX8Z3A12vxAr
qNiei3puNhrqFGTK5p7id5HrrbXWI7hFnGuAv92W2iqwVoSV8+FsILSwNn7m
JG7KtGlFSS/oN0pFf2/6jgWY8gUPa8LFAGSJWgxZXp6fQdIWuljXi0EfsgPP
EaLClYISt4UCxfLbIjrLYSklL/doc8Rm3B7XyVwPWSQNMxNzWDO8iKoM649f
8KwcwVt8a8rMphjIrwaQQpBjtLtclrxzGIwa1ZXWyozBl7ZEi9zuzDI3MsO+
DGexqVJiJaZNzYSJIw7eeU9CIiv+zw8STDEKQUdPxuoXlq7gNoviO3HFeHnu
00dRMrAM+9NfEpLMkmTcYqSUGktcSXo9d5j69NUd9WRFYERpW84fMlUbBoDm
gxI2FtiqkOW+jGQ4qJDeHj6ALAlFsx4ytMm5O1Jz9TUhHA4KKX84Za/Xnz2f
OYk+lvwy40ctB3hAImHtQ1kqyNmpIOHc/l9crpO/77AvsgGKeh0GvVUImvpl
UUvSqp6pwApjphWWSMl8C93slpbx8XY2CIEikWnLtG8ow1omUA4T/6S8CSLe
Or4VvJ4s4NMZWBt2nY+jNDxXxy0/Hh9XuMpHecho6cKqhgJL7L0vbsaKzGk2
1LMEuYh7oXSsZUCSZQ0zuSK6gXdSxhtr59ztWn2WcOe9bZknx748kw6RQoUp
SlPjnOqHPuSmW96BJ3i/7JyUMrTPAbaEzYHv+GDmksQe9c8vpt375YjIW7BM
m2hHWXe2vROB5q/POysyI9oZ8TdOMTnCymrppAfrLtDG58Ug3xKOT6sYxZwK
tlOcubb5mCQLEKNIowRoa7R72rdaPvhUhjWcIHhM6zAeBcHLLqvtoNDYa1mB
v1s/GMmAaQYIJ3AWB9gZfQHtkrKAON1T+PUwsbITgEwin2qUS99ByoyTfbN/
V9wluBdpRJFsXbnBRz+1DWhTz5dSYvawp9nY72JoCL5CdJbt4mRjN19pxD+0
3TmYDl+Ll9IqOe6wFZKDdDYqD6Q4n/FOVJO+RdCENentaiQzTQ5Hoqe55jlt
XF/y9tinjNTKUx+NXfAMiiPKo4ebJq+TamcxMcUGJ8Avkb89iRrw/4esOO8U
zMvGwXoR4XtN0pi3y1bMBJkf31g6iFdCyX2IOE0xMgRKLKzIWrq+GCLYKOop
/OeI3gpKT9WXszEg8EgOcaW/Eg+teysn1iQNgZfOazuFFxMLgbifU0WqpXVS
twN4xG4AZJcc0byUpg1h97dRcgQspLZm1yAjbI30Pt8JcO1ZxF0FLac9n7N4
DhFE5jX8SXRaGtEK1m7R5/lXR2AEg4o/xKfqt+EwptkgCoh4c5DPcwLOkQLF
BrFS50T/vAM+iGoXoKNc6MoP/3ALvHjPndGiWKg0AXlw696zkAf7t+ysTLKE
EDQi0CZOwfer2nRtgAPeC5bzwWctLwqEUbdy7kjSldS+gnfFda34Yc+a8nYg
8kWs9w/1K/dpIphpytzKMH0KJvwSW/gTtTwA24uZHL+qhsQ4+h9Hen7+5qqe
kWrUhfLPW31UOOgt7nTNDDGmR3U3D3j7fJFyUZ4RrVOidFUUxjte0VGHRR1q
VhQERmzwVBEnXjOHBbHE7jY8r2vQR5yjXo5HyaX4pcgliyYA61r8OQ7hbbxV
FXuqJV8aM08vzPWGY2TAX84dTaK1S66D28eCjS7UMrel3N66Tr6UUEkT/zNr
JVz/8b7Wsgc63xRdDFFzF2Pf4h4qE4upn3Ks1HBzTAHE0Lvg8ljqWWPyYIja
puKL0poVPlkPnQNxeO71pDR0Cjx0Hqytysl1m6mZ2g0U4dzYpXns0gjEoA0+
q8sr+oiEZV1UdKtY8XaPPNe0+m+XN0ltz+U/AIM9G7mRTsQgYDBbvODQHmHA
2TUQSbD5MeTKrpGhHO04t5/lXgbWBW6w8HRV6ShP734T1xvO9hOyJEoUh5nB
04aA1NIbMyz/P9ArKoHGLhmlTW6yVlLEYhbFaHIxfjoAm9kGaPQhslZlnNO1
UxPWNdae5HiFMss4ZaXRWVZ7D9aWhLyh+iMgKHsBojiouOq8xp3dx+InHS6o
dPI1g1ejQvWMNh0SpepMmw64xnOhN9BDO+1rIAyQlihyFj0RWI05J9E8HDPV
Ox5VK9/P/IHuVDDvB1KjNnC+1GA3nZlf4DRIgZk6yq+LpKmPKKM1l5VrEH4l
OWxNCpLozVr0Xxey5oJhnEN9kn8wGPjnv9hZ40oAUOQz7zx0bBMUGulAI7AY
MqCPdn0LK2cOHIoiI6j5ll2DTGwm9P2DMlNRTPf9I9N2Wa+7Qz3wslDLwxXb
GDHAxiogLY5AcEmtKTEjaBDyqTa2ennbbaUgEno/RBpRCQ1YVPaEPX8J8bBU
JQHnC6JFYe86NMWv45kQh2nKN6xVJEghAZurq2ZdvuVnu+DOnOMsdMAGaede
YenDfkPi3OYvx4/N8EUjZ/ieRa2+iTMUVLH/bMSv/aacNCuh6MacIB0zyUXD
rPpwPzUoWNfI7b5D12yLHuOQF73XYEFqoOuT+OgRecmdO1T9qMF81WPJrPSo
skpL5lMKXSWDOZT4gtY7vIk008JmOO6jxpda7PgD/0d6/U80FtRDBP92kRHC
ggtANcoPaa2/959yAx16Gh+0rHxNBlhlVCw+S0QtrgYXQN5jV8FNZIYZdEuM
r6O/0kqmLH/v35cWNVUbHcywovtSaqOkANtEGpbOGJcbLsFrn8U5lrzrzz7r
skjYUslgDIFBSvmnUpISola7uJ3Sz1whUsoKhPCxlTJGxO8G8XiXXDL7ln9K
FF/cqfm3dhmB3ZmsbyjojZjEzzgW9MIiCbLtRrw6GkC/h7X835i5WroZJP8W
rtjpzkGXkiVze1pQ670hUdtEeUddJzYBPA3t13EI+526gm7qSPQt5sbrpttw
skiWdz3y0RV47VloUWS68s9r4oxLmtEIErXSWpAB227M+6prZkIcuRHQbkoo
vQe6bC+EvavpID/YgMOlUPU6CwlQEn1+5WfYpvT5j7BpHCboaNjD0KTEog0S
yULtrT9fHodCnTax67LgOZKvcA0CZnV5arRksA1AcCISEZBcwq5/bfqXHzEA
+rc0rvwPWIsh+w3oUgpoow6FsJwjnH7Ic6vE1EFzbJp03XtCp5sG6x1lOP0D
B3kssmhhAzoHLlDw45aWtk7iF9R8UvaLJfvb8xJVYSNbsNQ3TvnDajTrEh1l
UZTNAhiHDasbJsWDIisvtENrrlhVH8jjScSQEKL7zzUt0Y09EM1kXE+piBWX
LlKmr6D6PHdCAMhMgqdW5rktATbdZbmgtu6Op70F2i8pEuBy49fW6pRNu2kM
Sm8ZDMtmCPIgfuD+KzD5Ik8n37QegMptU/FA340C4NZaDvnZzBT+yMElZYIH
9iL85oPu9FODoqHYdwV+a2mRI7Lot934VfMO7T8nSNxG8+6DpoUASzcJuZY6
DCk+1HkW/71S943bkckHkGCPjJtJlimb/XbxxNWZA9F7iw2ZYQtV2hZkHoB+
JCp/dBiMiBNlggmWzPq6vwFUNCh7RYl+IYW75EqsiGG5kk/cjLix0lHz/5Zw
yKhZfHr1WvNR8DkLuJ1Hu5VfPMhJ3x4CQnclt0iAV4rvMIYPsnUKau09BD/X
OBSqDExA/qvVKIQpUo3ZOuxtSvdQhrAn7ydZ4a9msSNn84htIkOVQcPs/Ngt
PMTLR1j1cN76taE4GcezIbH5rzEMvbSo1BWqMHn/8o+b/sq/rK2CCu82v6nf
ddH/nTPaka3irMARvOm3AK6UMqdfuXI+zoy54juLlL5/1o1x/BeXAsqQjeYX
54x1iZQcxLdURp85f4liO8OKvPycsXcaUqNiXPM/TynWTY6ye/gUFYmew+9s
cF2XEk48ms4U6Rf/LRsQbvYI9iraX63evmEKAT5Iid1mqn5rBcXcQqEzuQMB
42ydGBp/i5k9S+pulB100enwz6EuHqRuZgFblUrVVSi/jcsBGyEp8b4jrjd7
FTpggp0ETHv6cxoV73BQU9iIGFV6HIXNKbushoPkNJE91TC0CNOk+7bx4Ahq
zRqVtqFZW24ObanxG/O4/jaJIUs/KZpET6fkYUvQLwr/dGzS0KMCPZBV8w+e
6WvMZ3UsCPFeHNTMFoqIEm6e8dqWUCMH8DPgzwH/oo/eGa6Fjv11yqcg+9uP
xm8X0xai8xLM7I15+b3v3dQoGsJXUFgnmPAhR8ArPrfHJz2RtWCNbLAtlT9y
kQ4rgQPaJIWR9QnzdhV1AU5TyO6u/vRMbFXv/M+NsFA/x9IUfPrbpnQhrK7i
2YiY6Gn/Lt8y/fozqnDVfaQdboss/qNf71L49WkP7NTGq09iiYbNbdJQ3OoN
nWF+mYz3ZcuT1tNCBn/jEmDWcySZaSjhtf2KSj2fVBTkvT0mprNegx417Br2
YRiLiF+iHeF+HuV3ieYmGVBDOtNTD/ooQQk6O98wjrG9c6lffOcaM+/hBMOF
WXDBgkGeTOF1oPuzIlOqlz7K8A8zrVtGwmywZILL86hBVi4jN3Ke/G6Zq3Gt
QEGSdaQ6FC/0d76+zszf7ybbGyfiedmnzMegojqY2aiueTrQiS72GNEC0MpF
ZR4EpMQVjk4y1MOYJOU918eUp/ug5G9w0DNFZM3mu+1YJtLAH6ET5MPcE8Tt
ZSbVzxuWiePnxyXSKkS7cBuJjGa09/G7FLMXRly/rOfzgYDlRjEFVmtgMKao
3EKplYeG8qeZ2WJT/iZvXaTgG5alq/QzPvaUVHUnp/kfu8CwNsKk+cz0adAg
VoG/3KS0NYhjRaFCu6JQlSRfuIMNHDvz9kloEpFO4SdE6UL0tHGrcUBO4Z/f
NwMRMqRs9RL+06XcMVnye3h7yEOty/sSVl/d38WrL8c9BIvY+ZN4xVvk0kNZ
UiMvbhZi25RfHY/QdyB9q4+u0HXHDjJ3HyOXz0B+MqZ3Qtc2+HBJ4JPVKWym
QKZQ1pf+u8/pwIbq6k0lJOPxElhcKAhW3QyD8UwMXQkvWTUxJG/XzfPuvSZA
V62ZWEh43vJWbMxg/lRaDmCojVWJfZC9as+YhHoPVkH1iInooNSrHKHldsI1
+QX74qntcg/6NYK6kJYK1dmiQZDH/yuL5lrkw6Vc79V+z3ECG69XXLxTJGzD
Lr5SAU+i5EvU+KY2mtHi0+md9g7kghAADi43ub81E23FDQ0hTqqI1ybt+bxA
W6Yn1XGtgmiqXIQG4qyGjPQ7cPC4ELKhHc7+XRoZrB+UAbFVMxG8TQSKHomf
qGGSjbngaK8ya2ZLSmsNydyzPWHi1LIu6E/viYHkZkA+dorFdxvFCsxbzWit
J3kZs0ojCpxRvXYcqGeNBAGG9uzYljwL3l8OzTx8zNI0nrEwXsNHWrtDWyEo
Hwd3c+hQJbgCBn+taRmhlR0sTcjchnqZCCgy35ZofJ0whxms94Ixx2jWqoF9
Bi4mRhAqwYlMlWztaEVkHjItcLG1dOW3KRnjPt/OEhGPI57Oo4sVljOO9imF
5qxAnL1GGWT66fzxe3BqGdp1f/nvcC6ZA7TFNr+znVO3PQNdtGMs69y3ib2+
OWzGole4HYxEgilHaYOTQGflJAP43jPY4Y84rFDdmXVeC6gz3iYczdVkBbDU
T4CTHtnajtURSY0cw+Bqr5VEunOn55WxhBXf/Tj63+LSjMVg5YshyMM7y8RL
5Ulc4ekreHy2GvoAhhat/6otHLkeInejqHM5I3kBMLxb6NMf2XIKSrxtbW67
N18vbe565wEodQyOp683qJou2C5Pz710vIXvf1Keu6/K5HUILg9gn0YoHK86
5Y1dJHI87dXT7KY9GBLed2lSEIzqRlpx3Cny0N0CXPgdaRRzfhJI4ksm5rH6
UD/dYjvS5mEzfnZhJVIgeTrp7XnIoRG08LVNOnli49r9+ml2hZEH6sHyMNMg
7NWqj9J5lG1GvBNE0nE9Xee33eh8gWnJmU3Y3MHo1jOgvK1fZMYXwMOOOpXp
1m7T6pNKPtS4dfeSTGDIaz3Ldn24yFiQscvtXJoKXcoLxTOddjxa7RdNRAE8
DmqxY3pDOBFlTkqccEJH9saJ4Y4sykCsu1J1n3XyAqGwibvygk4y4ISyT6hc
pFFoYlmJkEA7SqRxLcOi66kG27pduX+XKfYbCSWeI+Pzu8e1aVBYTaJzCFL6
It2WuruGWKYMKGWUEa3lM6jjumadWurhqGgrPA0jvCCySyWJIbwRj6pAiwWp
Qp4qzCigXe+ZRZtGBz/Q/DbGjfScazlXY+iAUsKpvzR7KanPxqAdTYvZeufC
qx2efYw7AX7Cg199ZHs4Aeo5AgCllIREHYi/a4BGU8Q4PsL4xYVr2RG6JyYE
74CUUKVaTyioM8/vRR940GHpBrllZP+J+OKygAUhg6WF6pI5HT2atvVpWHHt
U61EBDin4yk898tQG8a+b7Z2jl3hlrWZHLY7Jd6gWLnC9TeefiLJ1Ci3p8f9
avXknoNkRAfpqFBjr+nXJSulFTQz5dYTjbHWuClv4nBG0OMBm2GqHsNVQRb4
URmdNzSTGti/jmBX1XvuChQhEDES8x0FYQeelK9ruCMnnTuGgWg2zxTNMXrF
g2we9fBSYPoCi+4/yKVRwEkZz4YZrJd4WP3zT+rhGveDPWVORZjHjdc7PnIx
joR8tWxbixCIvi/1MKr6kNI5e1g/56MgFD8ahz2t9Fv+cdz4/gmufz5/y55r
BFhY/nai5QqD/xGZkt/fNqJfGrtgyJYsLroGhT+lG7+VhvomgnFk1tR4BS/P
33vZMFOsW2sdtTOeSxeOVoSkOGr/ve1IMMJwxKN/EFelWIUVw3DCadVDBv4s
NhjzT+yHLjUbcQOZ6MvIIJoSh2T7Z9RcklPzYYUQ/iMsxvwiIMLh6+wZ61oH
mFv4ClkzU5k7hgHZRwR5XzGfUHCJfQDHaY6t3LHN76A9XME/wOkmK4DZCLt/
eeQC2AsKTN4ChCYBQBclEoYILQOpMcOvPRPqczZrHmKYbFcNNPYvag2LtSC1
rLmKTj7PJaOrMhp5sOkrw0nUsh/6W5zHAe6eLmh3GDlsm+Hl292+xy4p8T4o
ONb1YXxh3dY0ri9crl3f3+PGgMLQ5i+I/MKK6gP921YZxgdrM279R6lD4sIC
ZMMRCEb1bEfsEab8rV3/elGCCj0s5kXMi6IN/+rPvh8vVNXuq1zpM/AX3ieK
YLhtoILLDHBjudRYb73mMgjMB/6P7rcB3og5o0loNds9J8oVF8sd0TbPjCi0
6DtpBUhdCr5NckOr9ip703kO4OTx6EY34TlizJJS+S8MTOBt4n8ztMcIumRT
mvsS9R3S//3RTbJIik2W0QfPMwfTnbTfMPf75Oe23U52lrA5hbOHj0R0SGxF
Aaga7O0zMFN8e427+ZYGWXIFf4bnvjd5DuTovHuYH/+TYNIY9CjP8VdjVqyQ
7ckfZzsWwwT28j8TuE+tIjzQgCbdKxyPUN9/qA4Vs4x/8URNNBVT1IFdXz5W
5hHVBhZD4jEoYb8BriGtZyoY1fjNbiG+LaJCpOvD7GBdT5JuI860jDqpD25L
qQhHJe18i1ZyZcjXu/NXVXhiGYinBvX40deB311BXhnJugDL/8FVh8RotCTL
3vP8uLhvwMCyhxl7sR7ATY9fgKCrcai6LCxHfhCQYiw0iqV8IHbtfQ0mGftP
aPd8crP+whb9HBBnD2P/PjVupMOmDdp3JTFJdEqTb1SnuYcX/CDYOLbeejmv
3h7af/CTU87wAOS646m1ODeB8P1xkcXMiuEr3szMpVnbyGg0ZKlYSbcBG7fB
BBFod7ivddmXdWB5Q+A7pblrdrNioLQoHcawG3U1noLgSvj6Ca+DdOb04Ume
WOUsZTg2WD35evLiFeQbhCVu/muKBSghs3pSXIqDK1nHgrlSYiQo/q0iVDiD
gYobkLixTAqNO27RKQq0pPZFmrWHb7rBTSr671wBZmMs+1VPjnSodE+yKMk2
jVS7BB/VuJ+E+4xORLvT67X1A2SW1nS2xE8/wokaRAK+TVeX3pHzwnMC6551
+xvw6yiywE+0Awla3zof37ThtqGKD7JIcl6Jnkfq0h38fr1lt19Zh/2LOmUv
+XQ0SyxEN1ToAXwxPIHCcGLI9YOchhPFXRpxvgG9gTEfJwUeHigwMaxle0UI
CzZSfRZG2S6Cd/bqi7IX8yzM6y1NhdIxVHcWllfRjU2L4uklu4GO7yh9/mYJ
UqGVrtMZYH9tH/D/F/s0b3UCc8rXVr0MjrMPai0f3JcvozGmRZzr/3f2UDdp
whoW3xONzDXRQJgsYeez+l1dD2nLaVC9jmWvtfIanzWgRALeTDKs43KJF6nd
M60EgkZyWoQNFhXeLzH0DbCDA8H1uJKwUTTELjs+dy5JOkpVmDLUai6C0+p8
jSCGXjW93NEzszNu7+udbkHzwPhkVZ5iUMQbZplQ+Lketw9S0Jms4iQDyHTU
DQ4VFnPgAYE3qi5DIBmFrWhRz5cmne5LYeu8IQbCsoyVZU1zZP+zuUQMd1j2
LOXAObRevJVEb1oecAd+sssjKVQf2gRerJ/TCdGxO0SEHTd4J2HWI/wrECL2
JJjY565C8BjjWEAckkroH7805UM4FMfebbpxevRmhlDJoqktwBcFpGnB4hcD
4BZ3wSYVdghL1Fhlx4WR7ni68F4kQyVZXkxBcMtWypSDTzz3iq8QaON+hAiN
yX0qkKNOHmkT2nRYbga8+GZN3Bc3DShNIOsgcb2u/yCDaUBzmE7y/yQcTwEz
/Ke5PaOjvtkXJhE3e5vEkotiLZQYr3GUjUHcBdk9rk54caCbbutQm+5I8cve
y3DWSfdtbYpQ6enL9lrXJsIXbePeT7PasCjNJZiXw98KqlQWAxnaEP/iIpQV
OY01VXRhWKxt+4qGpVlxQJaTl0SPA8wGnsvc+B+PU7f6XdDvOvNGsrZ9HkwI
FEXIF7VS+EGv/SL6xU7PtT+k9ajrcRMUT8Z6e/MUv1EfEUcGd+DkHmV6Nna7
1liJcQMP5auzk3ioa0m2uZUkehqcwhqr8Xr5vwM7VKHGaD5N4obD5b5niZ3b
/C/8wxul/5YCgFg6ZnXtMmtzm09QuCGbI1CTV+pcehSenwql9+N2ijqPbyQQ
1zkFsJ4VvqW/UseSiKkRrNtjB2dnsLxh10dGu7h3qj9arYQh04GsTOqkcSDf
DQpbeI03Z/oYt1M1ebXdb9NRxAjGtLSVNviu3zqSblz7nnbCtOVre/halkwh
A0IEGxyvq7SDFseJyIzyKKON7nZAimvfguYudZAmgqzoEL4XkaKbtcmJtTqL
Yml8Pgfgrt7+neJhVSMGEv4cgWjcrXVq1Yf0OI6Ly5xczkhtlRo8Wyyqr2FC
9bA6G8iWmGU0VmFcch1zNvbp3uLbK2fh/JiJipD8csZs8NUKatz5WHbL3r53
KHqx4wB274yXOG20BrcR0OpEFBTf1QDt1QrRzh+8bTKpH/NM5SpUElUXsXvG
ipQC/MdxpYenC/0sdKZhoMAS5J4kHixfiV7vJ7PsBgNylTzL6YeWbPWAOVaL
Dj6MDWpdgaLV4IBAAyPnoOmCLrzyguAfP3Y7zHmtuKDDHoisFnQINf4XUgM8
ABnbaJV7Bmj5soTM6eRwQYfZ2tgwyNpzKATiG885ue5XESBqhq9HOI5a4ix3
6GOpFm7YkXzP4gZkdJZI5yM5GmQTs/r4Y1dcN+94m6OkcD+CM9n4JK4T8gTF
yCYIBXfuZEw6LkqRGze7rI/4ZZT7bsksNwonfV7BOPWbjOAZR/ulPXZ0I1fV
X2tL0gTAVDUYBQqbEcabCkT3DRcgVvLYeuPuORQGJVq9AleOei6dgZBZz5Sm
V0d4qJiJW/bgt0TOjU7FMOdDQe1uE3ynovPUCjposgq9MNkFLiW36d9YvxLR
TWYUpVh1jzSueZmPxFTYQ36a+Q+pPmR1+i/PsKSY5FSL9PPQNZmG3CqzDkdJ
P9QB/8+8ARCSqWd2wfSeH3LrBbZrd9fhPdx5zTPgmE64cLrcCQyeYKOoFpK1
vCAXMQu7DvJ2FEUXMmmnjrGCv3QLxr0wBjYCL3alwVyW+WL6sf+eGi3Y45c2
Im1e71dmNupp9eVQXkXZj12eyAY1ALnrvyyjvJeq3DTmXUcezqkqsVVyReGD
jZEkU3Plww9S2aHOP/spRHz+QG2Lod3byiVIUvfcuMJHJNaUPF9/lKUoehOP
BHMISNHjEqLOAbSa2X3/Gr9ZsmyERvEXKUeZquA9VF3paVUXYF4AiGXi9Az6
XT/b2Snd+UqV0kmhm2WvDVHAmLZMHpnSQO/3e9hlsFvUNpqObWpFZGuWj4bK
sFIMkWjr9T6fMHWdT5c4MCnXS3GgG2aaeeqJhHVlt5rt/G001OE17jo51uNa
ddhATose0ebP2oroBZbhaKT4ydPInHhVVWcAs3MMo3dvjnN/Y+2RsyeuFRok
qOgBRv1ooPqDQMP265HU007VBDUIXZsiK742Y4iQ5y21ot0HG7LIhq+fpZsX
O5VcpZrfWXlizYHsPKw5H5Ojfqns5B1A/Sk+4lvJlAFSlCf5gekC8rryqA57
NHhAYxoknunszFIcFBA3BBPgs6m42ArikzeXK9yZcjHYNDs3ljQIUCj5r2c7
UdLjtpX6Fijf5bBZHHhi70v3kZNoIFLPDt5bL8xDig42fvWmgAaJiqG/ugE4
Wcvpkv6HJILBxfvoE8WuYVIHWqpwwsuOHXkKCwPwh1X8dqovHVyIsoAVCmpE
wWtWLT4nRntC5FzyTI3RVUY74YjFHgI4eUoMRL3VdpIvlvUU8Cyi8emZHFZe
UEMywad808CwKI/eOMRN1hydnZXH1PqpTHIioc10SgxZssM5aj7g8+2RZuos
MVjdkyhcaesC0rcW/20n4n34Lc+BQcZXpuFvRhor10ASL6RAIqlplTQ+zRP5
XtvfOwVA0N/1Xx9p0cVyHfck5X9kbkyNx2G5LDRGNWwlsn7zXPljzhSgQEHl
sPOgajkYJfH1uRkwA/Q6p2elWOUxsoQYTjljBhhx4hSltOLGhZ9na2Kj7EFv
acO69Jl09Ty5JWe43tLRYofqXf1OOPEX0Mi/S07z2bYQHECGMTIdkY6xd+ko
HdFdjbHlkU7HdoHPn/148cueRKwb+Cf7ZdKS07gcgHp2A1Tlj9atWfapkQwO
brOVS/l8KH0cJ+WBMhg3kuKS1BBKgqJI2g6+AOM1HfIk0FRqac331gMOcmdu
xil5oLLLXNuAKfpsSOZVnkCQlglDpXX3kly6Smyxvm8UvWV3HOeILmdn+K6D
glkZZZv/MVDRPhGDBh1BVOkHde2sn02lujDsn6w6BmLi8RSMlz/9WkMMdeag
meOTGutZWDk/ZviER1jdfIhrImNBafjiuhUfIXA2Qro/4UwgLmNjBZNYvpWE
/JIhLoD2o8zUQpWLURkhgUieS+4kpnv8OMlVhqC2+0lMo35f3L3r5JXh82mX
FUNLHgF9ybcH0l7RZUvspOAcHr5unFROAdWNLDkXD2c47bCD9bQfZSbFPHDV
H/f1+1wbz3wbtOQ9kY5yTrl0lhqIWfE5ry9xunxC+fElxIxOJF2a8KFgvATy
biWq5RWdcvUasQ6cxtnii4J/YYUT9uEMLXaGGoCD2SNWM0YiTbLxtRRNR1ns
5nkefuNPrS2HfeHJnW87tvYKhj0BnTy/rkuoKO8BtQiL8RKPzmfTSqBFY5N/
PIIjt9Xt5JD/C5APk+Wk06YLToX0pxZuJ2nRaiyozGpTMaHH6trkyRqF/M9I
Suhly9P32L2grNQBlFfUs/EoSOGhX2h1Yc0Oa8f9ydWf85ec85f/WdtUCeWp
CcIInf/C3btMRHrXItX7a5wovZVSFEh3TvmTbloVesx2YO54f/JQ7swwrdS0
QKpf3J88qrZUY2HSRc881ZWczGbknHqe5iaZ/z9ET97Q8hNeF7JT1Z/KqKvE
IjyePCzTJKIw/9Om5VS+Amq8SRCV/xWoqL5p38tdBIGVUL/+N//1dywSb0K/
s+HEoI7fiVemjkMiQOKq4A77h2qHm0WnXKf3arwIiQZgWVg8FshZZcqxLVh0
OFCCt+qYbsPIpZF71norxmzqXESZhEDy9tyaXMp3VbxmvjZhUM7JiUCQVjvM
KhPHu8In7vLgth6HG/T4nexcJlCQF+ffYQk8MxVKjZl3vuu09ezmBBe2THKX
t0snCGaXw+MMpCLGogky+NufJcnsVMIpcYyWmhbJjlta6olFe9SsZFZ1O6uE
l+QRl66upkqyJ939WZaFe/whWGx0tD3yuFkRYyVoYh/jjvSGCElb4CV9aZM0
3PQ7huPl6OLyuUrPmsuzkV/nXvAXig1wL/sTFP2Q3n3t4ACW2K0DmjtLLQ7I
by8oVLvMqz7auQ6M2oduGPU4JPFpH8BJO29WmsGXgLfoQlyRyulpiL8iPjmR
6RaIqY3JIaNykkZd7lJGIVm+zYkBi2Y3TPRyzFl/7LvGL1bvvZnUx93O+cQA
XLu7xMJpCMAtMoWS6vWr41H0LcEBHE3rKcCQ7w9GgCI/97pS3ZBhAunUtfge
N5AhP9uDxNnKCy3Jid5u5MuveY/ifUUdYEvwtd1hi+Zcv3yDafdfRsCnWM2b
tUU6QzFqIoYSKqTpjPZQLhLM6VsPpQpBbc03ItyANMYSxQa54pesPmX+PB0F
QN4W6EOmoGujgYS3DrdGpoXhWd7++p3hbtjbmQtanl8jlCpjwDtR/3stxPAP
P5/Z8xtrNXMe9aiuJcaVcGBLQGAeuqTRwJv2F54p7CCddXy4Cr951pm7Yz4k
EFOx+jLj25xV766w0NET/zv1Pf7IEXzaNOaBvhU/A3nYYDjyAerzwYRSEndo
L904n33By3KLAMK6wm1hzjkRVcW2nMl8Kn96TC/23fpe8cAovCMrcUSgzIzj
hnNP+yKBiDCRd6OONFNUOPGTeOhx7U63r+PxQVbGitOoNjEvLAGmTuuamfhe
Zgbm8GmrpWA5B2F3ICBzTKSNJ4A2JnIe5UB4OqdY8ExmMGV4R0gURvPAx3n3
g1zZML1r6uyCqm0bMlm+Am+ABpzYwJyGeTdGC9550QhF3jF4p1fmbz2GQ3nc
aXkdHfeg9KAts3QtYu1IR5t1wXaK5z4nHm3hOm53chLb8pQsfhdi3vyZ3VhF
ZfLmLDbSLLZvJnUT+wHZ1Zn/e5h8RxPAubfYNRKR5qpThj05uYUIsdltzbpg
g7HMc5KANlS/YkN+Z4vrTqMJjpW3GEJZznjzT9+UlG9+Vk5KULbvUEJXzaOh
V1o8oeNtvCrxz/C/ih0n/pWM44Dzrv55R7Gi0vDxKFIUCo9wn65kIVu3DXpe
z8g1dJWXSCrb2MQ1c24//MAFdGgoZnBwWtZ8s5CpL5yH/FAiQrq0tXq3SmQe
/zF2FCpeL2Abkw/ORry/L0BzJCVQuoC2ZXBHOVzV33iAU2x3S+pkt1++p+tV
zoSZvCWiWwvDlzVqEnnQ+D/RhA5zTkPgBs4oQN+nRzo/cBmEzSVlSEAx6wYU
I7KR5NFsZMuiq3hDsRkyzkBT82SNVmKa6MYLGQTKdRk7WITbUzXdUnlP/nVq
7ZBt3WpxnsWNb79a/w420F61mSFN1TK0ikZwO9nzZelcg+ux7OE/x4yvah6S
/uEVJvGJ5k4AJTKIMcV4jXMF2qg30ttQAT1iNpoCTKJkkUixnsEfQaG/FLxv
yU9dh7dl/gRH3xOSLu06Cj8o+MWME1MaIZDOPVE0ughPrOoY9NeDyKnVGY13
U1eRew+7HXhLogIFO+T6BTfTaor3LXKAF38pirpV1/W+eG+RhMyWqIDgjU3i
B7knQfTa2weCUnRVdpYXCtTibLhRd/AW+QoVp95Qm8Vfg8J2bhZW327DMRWm
v/ALSNRM4TCO27mlQRPGZ0YJb0E/XBGZ1Zjwr1L4nzY44cY2Qi9skF9RH0qL
02RxJSrKo2iamQ/zSGIzF16vtftTyY+a8eubk4YqAleD1CELNszdgU83N0Wn
vHQr9uHnk2QCCmgVOMFDUQYzb+j6Ju4Fs+PzcZeLDfGDqbXU0aJWZw1iO7qs
5KghDU6O6sLuHL6E8ROvOyzAMOxOCxFsn5o9VHsiS0cie34Mms79s6rBnC60
YpF2iv/WqmLX+GPQVqfSk9Okf3rdXoAa3YJvllmncBRwYn8ulH7NHSwCsA0G
0ReHO920S46VX1zzRmPrposwwZWNcEXlPTC50ieSsO00Rr9OQwIa3LjWgMBv
Yayi4AfwgaVGXb4zKnJLLTJoPhzXwphBeIJNgBhJbzj3G39fNxcpgxPRPD3o
1kuyiSq8wXDsF4ZnOjtX1x2JEyR6A3OU2cNGVBPDcdgNrY2v5aKEfhnZFMBU
lnQSIizmc32/qEhP8VloAdgmSUfSAMcnPZnvtAB37dmiiWhdsUJlN2GzAlDB
AVx2Et7UBe+XF511HiUu7M1UKM/cwI0fbyXHL6Opjag/ZjMCe8EzYf6pHvNs
T17VlJ+RtwChkHV5Q5VZdKo23z5lprNonqQ7MUMPZ9JQpIjou9ZpOLA3iNHJ
0vdbcPj2L/VrBkHWNrU7xqmnbG84ln8UkjMFeOQw4uUcnjSaR8SG4gfkOTtX
9on3/q1KCUgFxwZsK+7wQyd3F7YY4WZW4XxyTEi+g+A5MZhNrF9ohHsSKloZ
wjqAbCm/QWVALIxvCnevOgQCF0l2K+L9n4ywf5K7v3F4006ZX6op7fM3S2b7
DbpzCvNlDEVrrWzlFoUiySR0YcluHKAKpGeoVI/kAvmXXa6LLge5+upcYgox
AP7M7YshHuRbP1Ici+vdNt+GSfCOgutaxVNCSG91u2mU5gCaqXexZ25T/4tg
cyC0iObs0dIcaYsyfl29QpRPghNNmvzwpMXvNH9z7Y0nvxSI72P8qFN9960T
RYiMx+z2p0zR1j/dyMOK9M0vwjywG5ZN2xeX7JSpjbJ1Ls4s8yzx/FwnYzkO
GIDPHiwnX5KrFyTaBcf2u0JMFyEVcRAynxbFIJaUp2QOlR/u8BDfnfljQsO7
AHwIhpLc9XMj3ZjHuRh3BAqGDpGD9UR7SggPICgg+E3kzaAsGn3sNcKRlquP
3PZxZuBnhAhnpePEWy6V2ypEOkC1/zKv8RcrSJARAictTIDCUbK1mian3GpA
PZ3F5leD2xU4b6qadAa04NoFd/MU5j4b84XSxBKP7r9vvm7YrWW1XGCjLaBm
mBqoGCtuBdXNW7iUtDGx1saPKyP5CzO/lsz9pkYlPChn/la9jVieqel7ElaT
7Lj+j6eYyiF2HaBG0yamR1lk7hwQDzXoRkk9aDOl9PC/5OeaWz9cbTYvZyYS
ctFv8bw3DpzdzduhYAtvX7irlHnvtRPD3+0+mgHPl961u+JlHm8yfCXuCzRU
t1sVYpgsC9/XhuXqjZjxZUWmyW6daQ9TqM8S46ib48l3LeZY1R21L0mjMu5Y
aFpxGbCvlKHaABZHqoCs8nZLVy1kHZGPUqtMiSeAe+HPKNf8FCuj/Wnd8TYA
8+CFxTqAMV0vN200CTWMfWvuskCfbjODix5cV+RZzGyuS1xhmFAFjTT2x2gN
kS+hUv+73GBkWU/OUT4hlSurvYR4ECDCdnVecvN1FNs+ugBXgMEHCm4zgavd
WjRY/CRNkyPft7BeYBbwk3Me4nPMn3Z3IZ8wKT/yQMaCXVvMNimEyJImyMjX
tv3qEDPCY6FqG8kEi6wuuA+zMlQnH+n+afGzoBr6OYXVujQd/UbAbPXu0y7x
QuBNpEV4bDq2pxe+I284vC1xfp/kFmw944FO9yAk17TgV8yhT+Cw7wv9S3rJ
MHVet1j+ZoiZelTm35QWs13fS/duTdWjHg6KfozTBc8eKAGwBb3HyOtM+32O
tmCi+Bs7rwHlB9lZjOrV8Oc2Aqu5veXWh2qJzfV959mNj1CYrOinx3/44Rcm
QgLpe/0xZ3JgmFyGZrCO+VQcjOYY55Kn/tqGFvZPj3KDXiI6fisMvF9arI2J
cttIePdF+lqbu0zb60k+iD/BAPKqmqsgWy3LWRX0OizKZBQgiD9yS/aobCmb
GxfbbLz2LAegOaf6ohkX7LgrAwP6wjz78YYXDFpg61wesci5rEikw1b59qYa
5JzR9r4uSTRTVbYETLFXFg6/WHBH8eZPFJsuGw/l0iAjmr+TSwmsG7rxyeyG
y5kijC3o68uNfzfHPlukKZhnmpifM82zvVGwStXyZP7S1sPbznFi3GDJvDu2
tpEqTzQulJdT8+enHTYUXFTtZf/SZ0BK5yCT8mLB1F9mBovNDMS37Z6pgbRz
XPci1N+hSSp8ozGIC804uplD/VIzbWF4zzfClzUTpfVrmELSaThTOcja8Mt4
n6yLZaM6R9GvjLi0AeuQlWi7khdCi7M+cecZe6V8T68QrxvTFB0wuW/+Svc2
v0xWt963GJiwa35MwXa1q522kpH6E6fo3Ig5NCLkBHxTf8xEnVoxYJouGnfm
FDx51GleQx1REysKWmfS06GuDLa5BphG3kdXGI1uad5aS7tSa6oiZ0AnrOqC
SckIFge1+ILyPupdQsNdMt/Jc0PoeSNZc7EowEspP01Eh81/dUQBVtJy3Ooj
yP4bZNJuFx8Jxx1tdMTtBz8BoPSvh0pbXg9nq1K1FQXYCmvHM1bcMFV94yep
qFnauZIDgkMi/9L0GDNFeGmjed1Ei7Ptw6Hf4c01DY8Mc0K9K3no6DZhZi+I
U5OW98c7Y1RsW3O1zMDLshYYbdMVcviv+mbK4pO1tQYDzOVuPTRzrIgB10rI
9ooMBPTcqJy66Cd1+npkLPTDwWYROg7F8Cc8rWKq/ZkxgVKEJcgt2CY2rD0s
IhM84ARLsh0WMMHYMfwcJXkHv/zmZn84tTWyZhq6icqmI2ltYuJjAUJsaRxM
HXw3wra9ZjHjJ4lsYLgJtO6BmjnjJeDXB05mbJQnfKyKzQ2/yPqhqGR0Dez8
dI1xbcpflaelqZiKlOqXblxEVeASANlLMuEEo5sjRtrzHtZYY2/FAeIbxM50
g8XfVu0Mxcf0HUc9aIUZAixnzc5OPFPOen0j+rqO8WUm0zySzL/F77Eq2xNL
tHDnatGokUjt/L2Xm8wuonLJcWWTUQ18EzZ+VwMeIn4wGb0/NOjTkR0+xOad
0j9WVvChgXbjPK3myNa/HsyIjX0b/9QqZoyhR5wvIElrljHU4pTSxQgXG71K
wPptJre7U0so+IZ84vRmACvt5TRVb4USvUh/IA4aYlvQNxiD8mV58O6b7YkZ
5tnHfdxK0Sy+gT+/uaTeGWMwfOTF0YIBaM5gTBWkIDVBgMppf2BNuTFl9p5x
sBJjoM/o5MjrHuvEWq6vgoIJRKtgpxJnlIgVyfJ3mZ94AYHvmQklSz4nRk0m
vxl8mbHHz+/8t2ARCOw4i/Ua2k0i4vnBkesGjsXBMkwUdgH+Nc2fX9W2FSFt
wA1aamLP9vxrv3KWQ2z9VWeBotvlNaKIGH+lPomPgYE1nu2X1/O6XYBOQMmA
ZBW60TnyqMmHF9GukpI1HANjP+Laz+MKLadgbx+PeodUqK0ObgSlK/5YBfLZ
9Wv/URIMSjxAKL0VPfBWCHxowqpcHYYPcYo5yLh/ULGFGFj9CYgpK970nsru
iqd7U4+4b9HIhw3cV/OcYRbOsl3TjTEm6RaetfFUnurAhjADUlNUf6ZyYzGs
ntiuta+phURAQYm1kXPjHhkM9H2lk77/E1jJg+1Y48w0fldFcYlJs4Efepek
4HPQf4l1C9QdsfqAgCUlhiAYCIrv/K3Y48tiV7m1RQf3fI5NtElKXLmDbMfc
ZC3VKOFm6tw1RuJie+nY0DcwyAJIOHyX3fyd6700J6Kx0hPc4KqN6epudnbV
ftvmhNCli4JULQ/3IZnQIkoYg4crLlagWYs6hk4JA4LCUuYcr+SBtrV129wk
4e+NawTSsRuIczn2umGSvpqeU0uVzMSh+Swil2V82dY4gWTHAuTfWqmMHgfZ
Vwx89bi8WV2oCwocazmkrabGogooyUdf6NkUgT0clIJbtkYKsiKoea8N8O19
cOjuBRW3YeX2TqCgF4dXsXIoM7S1jwL8fsQcYG5ugxRZZcSHG5yorEbpd3kW
dFV+5Tv08lvkVPt9/yxeyczxMzd7JrzfBf8RaiBD9jCJWI7As4mPwEroNAKz
qGbvwIqxUes+KuS8FF1Z4F2yI6o97wC0grSpoHy8ptEVAdc3zNEKI4kSFRWW
xOHi0nJiuhjBqwaRySoSmruyoIsfgqWctzQo73dVJ5GHxADJRb/zrWCMh4Eg
hqPFIEbO4oCAV5yHI8QmWBmg0C6T2OrMTWDpexeHO1SPb+gm2HmVAkGhnfxi
4RZHczEQD6mf2RLvcGIcLHWCfdQwGSy2dX/s11tP+g55ZCFt7a3nQafyUKdI
6jMkcI8PXeIw93z9+rGWz8MpCZC7mb9lkWTq2QOM3hkmLERhLpilMPj5a0gp
EeYfXpZjE+4WL7Mv2Kn0Wq9ct6Uze/a2KKJNV0BM9h4frMLCw7RLHlYT8QHF
x0npeL7N7hPQAAaACn+MYLPO7kwFbwxEh6D2/Egor5iMfscAP+3E3k5KwYs6
paM4iLO3qMoePGa76IovB697ukcMKIAyhUhpYkja87vvQ/erXAPuGrSy2f00
ZnPoK3Q7ensP/RfuDyucb4mWpTE2Pl2M6Dct2hE4I/m40+XFcEyidKs7Idoe
VDbPY9qTxp1sI9e26w6vG8i6BAEJk4UEi2CNYVd6w4IHpfs6O//xOQ6lq//a
89wMH3jvKAQ3kCUk2S32jheq/2OX7Wvtl8uV/cJ/GwBLhR5KLRPpkrZziaF2
kpbqfEHLyCIi0fGYNkSjfmcX29oKH9uIlzVhadIHnDxbxEyOlpNLfpcR12n1
m5ytVI+BPtpOVtQOOx3L1r8v8eswDsxQrR+JDW9ECAtYOvfllZlJTHlv0EzK
HaupK8Wqruu2HHqC6tp6QVZ0c/MdhnG3jK9IdRur+od6PVYF8jMG3sbCB3/J
z0c+afRT5L/cl6CN6nVVFN+a7veS/sjpvSN0u2P1aM1TDG0qcUxn/ZnOtyL0
Xiyy1uVY6Rao2Yt/zYieu5GNww9UlBE0bcIjAql25oSmn6yQPsAxA/nO8jEY
Fg3C092G5oko+f6iuKv0FIKWEMhoJEnEf0M3g0RmYJS3oxg5J5emcyJ2Jwed
/qcuDzwSlJzXp7QbWwsrnwbECYjq7MGKHtzrNw4ylJJNpn4Ph8UnNuz9euSd
gXak5jTUYNsAHYNySU+Ls7XY0OtxusHKG32FCvDO5tfzRVFVprX+JkgJ9ALm
jtZx1XamWG183jRSe2yTs1EjIlP03uMwUQie/PvrqwSJ7v0GBD8ppBL/nX8P
yySlwRJKZy38KmcUlaYR49pSVkEfIbQfT5ikwRO+PF48RwJPi5nj26Hg08bU
FMgMv08uu0Oaraxd31/yOCAOrRv0hT8CS2OVf3ajNuNZlKpIhkrm5+OfnEql
0hmUUHXg7v187+3fRmMt9zK0F4KX9frbHi7tYg+7rSsWReyNu42eNJt7oew9
ZkNhNiJ1JFKkT1R2d0WYGGaVIpVrcEbrsfBHk+XVDylV5v3rQCH/JNs7dlDd
f0/hTR49sskZJl0Pz5Ib9P3yiROxFeSgcTjaSwMUR7tLd3qKR56dWaUPK6Eu
kyeL7543r6H2jJqYHmy5fWTC2OdrqT7XQ4ai79aa8jti1+M825GDniOGU04A
Fw4jMPz94dMDG7dz/PTIDs4UKUNn4xedTj67QiWm5ZB5Wor0hD5QJWIZjy8H
/GYMvfQtacfzWYXmYi/OKonl7rkkSxdHmUMym/sLRl7HwVZkkwyNH/Btn9VW
JafU4wAyTBHzABSGojFyUJ9mkNxBJ6mUq4N8eKpchyue6ZBHYyBw/+3XScuL
ZE4H1FbBofikQxnCFbQk/YmtWr60ye9IQa6g5P8YFQJovh1TLdHUk2pFpx6L
dNi1iA6qXbO8/UlVx7y4mFckIySB6cYZTlTHVFtvHrkz+9p9bkBSmgIZxwBX
tbquawHKFCbrFWpdtpz1X4Xag8qLGdJyI8wjoR5J/jGhKticotKfjFkRKZo2
sd4Bc5ESgIn9HOdlhzWGToe8Xb8GPH95MOh2Ts8RsG9yqv/6U0XNc91QoWsp
9+xXjoblfzafCzKBHsVwGrRkUgPw3xk5Hqx0V/Cnn0KnrzzAaW1s3smYLkSD
9qvcUUc3nSEPnA7kK6bKtUgkKQIbTYocVrFZMXjL6LZksYmxZCaqBbTUJsVP
J/1UiByl6dVHn7CMWSVdJn+DdCTwdzBNJxxEZAr+IvWb4kqDgyfzsFR4iwqj
uwF0gIRoDb4/J5idC5PPfMXsmjoYy4vqWwlAcHLhwoGq8/T4BlvQfliNXBs+
CBn3xsRFgHw0kRqLEBUwVx9miLDPqLjIt41JbtnCSzhTW+sBUdJLm4DIfWOC
Xy6MHEe8qLsaZB/5eQWB3fQFW4IZLhmCX0yjcStl1jbaOlsJu129fA1G+oAc
HHVC2gB+Wv0oKOwSy6q5Q1minN41wKhyUQA8r1wC02yLSsi3zyFxTLr//IZX
0Z2tvr4s7q2j0102PsxCgZ1JYZ9LUcQe66gWU0vr+96lJ8pMx3H+aQ9jhZ6t
8j196zzis+ClnJwf8pOZ3USynUlfrUcPIo6oLaEojcXxtxT9suH12oEs9EHB
dLFJPniIYcDFfiVOrtNfMiI5C6+l1qeU+SkskeAxXIXbLMPpAbywIlARJNOG
5grOgboRggaRaLENPC9drkX+oOj/dHzZX9LkP0h2eTR8Kj40cryqkb0N92yu
y5AWj1IV1XZeO0GufJMs+rDYB+kY4E0FkJn7wYIN3+3M4Qtu1uctTd0Xl6zi
UIJgT/+EQnwG+F0MY8oR+A4ULE+ckZ8NsZpxKwNvj81JawUtOhZqWCJFAP6b
NoVztn/6QLLXeMzDjCLQiNMNTeMk+O4yk7MNwYYP9BE5sklD6lNOSrThKRH2
lOTSpr1O1ItZXtglBN0ZDirfgXxMKZ/wWsJUK5Xh6IQ6VO/P2QZtyMrgs+P9
SDV+gp8/WtnhthyvGeS1tbu+AQ4HwqMNi6IenF7BBtXP+g3arMUjl17gUVOY
FwM/0mVxEer8O/ooKTXks5RzYHPgea6Ci9imTp4A8kKfpeS8Cf11R22x7+wb
Re/OgjeSDXb4NEOFYBaKDjoX2QfAExjp90RWjgmDxQ5mSG/D+u/wJCe6YJP7
e76Kbu/MXoR3FHEJc5Pti9mFCuiRFiSiuVCrV4CZHATc46EuTHTuCfeMivOP
j33hnW3tLoCCIdDQIz9z+ac0EMFb9aU0lA9QVQD5Nrd9Tjgj3x3soGsQV1+u
kWz80nPLn0qstLFWGFadiZ4PrHacHbTj1SynMHsnAOaOKGMkQb5tutAvTSQB
+DQMsfVFF0k7FgwrLM/t1Z8ST707TdQctCU4NOXQGC8m52sX5D5xm+vlkn5D
HkIWlj2r7vjDIsNCyAFGSi1h3xfMeo+Xa9rG4HEI0EIRQFt8o4SAvxbQIu8z
JSEUHPocseo58ybbMGCs2F82SkKI1vLB4RPAuJoDDXPMdW5kIEzIa9V9yidh
p0B9f6uQ6s+ilkcEq1/ZRgOgnrRm8uLm/wJuoyhY0Shdd7CYuh4Vob7PYqjS
tHmTdTFNLSIYXJ8cZafjyZK3Z0WtVDgdQPDJCkStx2uyG/bO4Zti/A8vyAw9
uVVQ5XhyM6OEcuEZxNv3nKJBTkGZGlYGB6/1Qg78GtWTSPTNAAxWKvI3jze5
5+Ztjyovccsz6Wu1NU4UVLBdmTyG5w/WsC2d9HgbjQj/LnxJRtkBU1UqsWlQ
jKmiBrBg5OuuirgS2UI4Zu+D92vrTSjI5jIDaU04VlUqTmYlDE/l4lmzM9Ef
57aLaM+9BgyNUXqYu9m9J/IhRKR2dJXAq7bObmyO5xNeKHbJMrV+1E9G0e0H
p7ol69vELsWmCPaWA1/ufxkj0W6mUV+Szr/7CBKu7mwPKDaGo9jomAp5o1z+
WYKo6CCm5+420ohz45xPfIjLyDQb5mDkv2vfgTXSBUeLNrrDeof5p0tDtyld
CZwTGVeWVb/tn0H/yCoPVX1dwN30rO5g8eqbpmHVip65okoyoFTJopcaNkWB
Z8gi51IhQGUvWEAGRRTuaygYqq7QnAEiMGXBeFRPu00BrDedXw9y43cQ0DxV
d6+AWFqvynG/L/PKz7cOY+fLj/wu/KyBsvY/N1KDmQ/MHAgkwB2H0Q/h3dt3
9k3eL39ymsmQ3hPokqBtlct6AKtmis9f2wve/zwxJtlxT0ccPxANl3Rc9k/b
+EN3Cmrmo5NR+tCNnjsRRkVR5sZ/nNilQN29JGOJ6LFDICCnwlMOLQF4Nnxl
u4uNChVJLcoYvYg2uwFB3PWRHL7elwx5OwFWYVmnyPCVaoLCvVqAj0s99AKD
ZbSoqpFrssDC59cbyfZaALnrO3VQV5gVXDSohfOBYdwldoslBeZegbVUBJT1
XLF7+zPTTKeO0Ljd4fp6QBJMVJ32zFktPqDLCvuOf0ivp1WBb3X+MZvYwzca
zqGuM8tp6E6AV9Fo2yo7MXZpxrjH07DZ8pBiiqEojF6vQj6uoNwmCJHO6QnM
vfeMaCzCDViII3hzimcN9PpGMtbc/YFmeFO5lHh65jUTrQWHG+Cecxu8UIPC
JvpG8cPh+8ltCG3trBz4F8s1ilVNs2fp5aDE9FOZjsmFY5wz27Lyr2uvIEyO
Hydtw+zxpH0jrdmugEKy8Pw465nhGMBjzekCpPSklewnGVSVUoE7iW4Lu63O
S5RukxJOI5mtQMBFMGPMPt0g6qVvvY5cAWyQNLDwjaJvtTpiUUhCQxQzmgWT
F40WjHbTSKpSYfBsATPiuI8bjjIXdBinl2tZbcVIjt4iN89vJeAi9mWt/8mK
qXpeY5IRMftDvzHFOYASGO+lSmGNPYD5TpA7L/AjbpCNu6+RQuJk4bhsWmtm
nsA2M8e2MtPPeKjTSYLQWiytoEDJ1yoRYS4wDGCluXe3i8ee6jmQGIdyL1r2
BFoDZ97x8WiDnxc91CYlbBoORS6MDD8IuVL9ZsWpEyXZVy2DMFXQesBmH5hF
SQnCU5sGAmt67l/DU8LaOW4pTacP6b1pFXKxRulZVuhSCun5BaImZwSI3nfm
XYfR4a/vbtf7wLsJbj5E2jk5hXrzD8KtGMEgoms9zRdYhq0vqA8VDDdXG4Jh
lv+5slp4/D9hHaw/+dTHxMfnUGU7X1hRj5bQEK3PPkDwOeP9mVRJCLgFligO
7Q5EvUut+0deJvqOC6hpAvDkbbCqpSxN47QxRei9VqGAImqPliqkseug3azn
0HPQ50ylUJU6VtKjW/HakzRwPLdTolU7bncMJlJHMqE06AXiXHmWVmAt+hX7
by6NV3mGc2KxXYV0v2+q6slFAMDrirv2i1hOjO9lTaivMOPSm65CLsJ0zUSA
gNUlRwML8jEBIv7rzdvArXCxHmpKJJHT1zHHQlL3WU0FasEFPTUd/g4uGIqN
slfT0dgi15leVHKumO31SkdpvoWrUnL9jfDq/+u9CN83G6fr0AXTet22OSca
E8ZvKxK2GjPZjtHuZtAPQfgg1PV09byEbCpyuLuYS4Z0BnGGQqaPFO/gZRzv
5eeZ/8MjX4bc7VlZV4GPurQns17nB3+/13j704QGTx29zx0DXXzpx8vGOQG2
w7kRpU0pZOtz3kIqYFk5gKRaNhWS8/w925VJxxWtA7QWRdX+meH61oq26dnK
Mv6rqf3lN+C757aqRQGnFGO5vaMkWeRz6aqG5wQ6CCp1Sw65ON9kee6Errlb
a5U8XcyK4bpgkVe3t9AmYqeF3IhHV7xyfjwJGQl4qkivgwEMq9TdX1c9PRvf
0Jv2yK5qk1VoQ7XWxL3pBZm9gMxGY41xaZjxhHRBW90BVFojGfDQMEYMs4S1
52QwFYkuzkjMVUS6DaqfuS+hEFSYIQxKvF8PxQW+2RQ09QsgjARVMBMYbOm6
NOu8Ro8WCT+EsTJ9l3rkcAwBvRNLbg3o5XzIEgeoecCpGBpl7Nw47Po4mPMJ
DoHh76RVv6se3dH8JiqKNVZaB6LBjMeE3FQVF8RwGOuxS2CgdQOg+Xyo3+ME
F2km5Fu1MQHm8sa1wsbFDOr4fwNzkyhFWfoJURMNzbySXBsyV+gUUr5P/Asa
igJ3e27ew54+6bBt+l48bXpBeSm1cJC/Mh8fJ0Xh9k+ZfGukbJbOOGyPsyjI
YWiGFhMEKqXN4NkxMrMBJDIrGIY1nqu1plDJaMMy4B/PvVar5Q+k4K2tQtag
EKNT1JBombsfr/l4Xuqr6pAqbJsgYA4bun7jqJ6IOwYF/aMGvMd3pMtsE2+O
MKMXRyYyKGicwfOQyN0OIoBFVExZtqWyZs/1Rp+TNNShePkNfBWjzhxyr2LP
y+qtc3YKTBPUhTfJ5ZzvSumeQh5hxiQ7EP9yGqG4phRBpkj9TogarMsFRxO9
ZklFcKmnviBr9QpZCy2b/rD5VPo0ZDRDMRQhSpDb90uHh0e5JQomtcpqMt4d
CgEPkAP/Rgw+sWN3MoI/LzHVLrr4+O3nygaIQxcN/IbXHgEapokLRsOQ3PC8
adnCMsPuw+0pFLc575baT2eUrroeW/dD0Fn2OEy9ccDVkBPm7PhXaFQlqFyE
NwRTASC0+X4wDoMRsbEgoevWFhK3IwjyoTBZhMy9bkfK9W/h+OJHEra59kkH
56RJDUo/HbWT7qjvcWU+LOz/znfVht1+67HPBz3eg8AAFee5hiysF5eCOM7/
u1iwkpoq8fnkpXZHjwgal9mkE+RMQW+y8X+APL+bQ6oQC+cDqa6KTk1+KrHU
Y8nJPhjm+COtff0zXfeX68HOOD6CKIvVa+qS2t1OpgPrWhYXdrzpwuZmUE53
VqCrI5Ye0S2H+hpTmdmRV2ZM6Wxv8ayXq8Qb26Np2XGdVySnPwSTXj8E2V8q
GKpkDOc1NBbQDYE/kLfWJb2594OyIy8bsFDGAdyWhe0AA8tsXj6DctH9QCFg
wF7OUQtkoaXXetSLbpcxIu5sZwFjqd11LkOXq5a/d2mOht/DzI2EM0gEb4dv
aDzzY2Xu0xoIIfsYxlULrU1U47TciTHokK2ZVrbHfK7sHvRsm9UvbI36T3uL
RBm8+V6s8VSoATjUTzMFBfwOWV+kPbHJYOXuct83y1/WZAn7t3m5skYDXxru
1wp+5TYoudh7kVTSsLd1rRcU5WeMZsLuxxRwOJmug5P2Ktq4H7LqYSUClh1J
RjEPPe4kdf2ECL0J/uwMovCoXeNV/ObKSToRJITILUo7kJHL4zVe7i9nOMBL
F3IihCBHTpuJvb4QjjdX4JcoGSRpi45TgP5nJk9a8RI2C3Beb12e56wu6JpE
ruoDShNUVMf7orKDZTVsfwexWyLqEuRZ5NXT2nLrRJUVQ4aWXO6fTBMAixoY
hwXmVeTY7LMaAtWBRSNkhek0o9lxL3ps7C63hCa+CXOo0LiRrrbu/cLczEwK
bi//fms1IS26ejKtPhd4mYGf4TGC/kF2ct5B8Y6enCKBEbcI/WC7HcGTVYZ8
yxP1YuFNLM/xxCV5oeOJZ6mJYOe+Vl2eUAIyAbfWHgZifS1PtYVwUcaqm/QG
fN8m8cVti8/CtcbtUebGxdSdqeIl03IpGAMTAv14dXAHx0aqEOl2bXxmwlms
urf8JW7uzgOWGzPu29vj3CdZeWRx7Ixldmo7OXFBEa0WvQfYp5GcNBE+jW7q
LquCDJtQKz/PZp4Y8lP+c083y3sFIcz1FrpEKWMd3ZYatfb6cpStTHqLjjH/
wn7bVlZqaQap44NkfQiYMQ8K0V8ZeYjCN17EKttqp9cLf+6qUWwD8CsIDTM2
Ig+4kGPFiJafr6WBGNLbuV2yMwCvdIwye/F0hWTRSdwW1aTkoEq+41LmJ0yw
gmM3lgazCKdC0zKJ6L4iDcoLBM9XCbTbj/dVgnanZJWuDwvF3xvrTWUbHpxg
DWd0BmqM0Log3MKuTqvOLN4sX+rT/8OLDeaxmM3OpTGr8TOe/FuXMANc8Gua
Nab2MhtQCxSjmiyL81aZXNAShFB8wOEtD7fqXy1ONkp5y3W826ozJCIFrPPA
I+jmu5HbnqylEpmfGm+g6zPNiUyOjLOMqLJyLl6hEXLjTjnzRLHkI7cIO69i
rBrASqVPELmRrX03HhApC4QUkZhnPGRml312cJnPm0+9GWKpOgBmh1vBlhX1
k4nlXxXHJ0Qv3sgJ5lxXEz6MXqdvInyEYU4n+Wr+M9Qpr48b5lv+kxJMlu2a
5h1KpPtT2XCaJsi5XaMcktr8jd9EiS8b/4TGu/ha/OphEfXIy1T08oCK5X1P
ZZYcVU0QJoQC1TnItiGc9IxLdvgnSYNiBqejJ3KuCGYDUof/1QbSpW+Ii5x9
WZxpVEMytTC36D83JlPlReJaoAiIxupbytdh5jaSHLG+gudyTblWnyGaToDZ
KJs509P+m/oUexVxabvwU+18Xdv+wVbA9d4SIX8y6bHNtBnjO+WkjITObyBS
JnSTrW7k4stZVZkTtAxDCwBqocjm578Gcr7iSZjkCBNa9FW2axxDCBcWp4LS
e5rST9ZoE0Jxk0Xdm3HhoY/BEfXIFD52H05rtpQR9TwMpbha8uiv6aDti7nu
DAZzgDBjYRPPZDmFU3kt3WUgDsHqJEGI3SH/5uzGMNHL6xzBMpNp2/SgZwe0
egpLpz3iofkm/v2nNPDteukRGmB80i4MPpP+ghbx5naILbJUGpbmBU3rcPXP
bon5CCCmPmKimTTIoYvRmWSA231z73pfNCHmSN6kqu6djV4V1Y2mLy3hqW46
JmwfjKwM/4i7Jgh0OHxrvko71NXFlqcO0H3xlQ6D8Q7RWnBJvOV3DMTx9eov
grZzMmAT6/VxZ7wagDwW+xzjfGqd/uQqZ8s+IJA67ojpMEhyRIjIBkEkBrlQ
b+3R9SU+TMpFAir9wamI6K8utlmhkuFr6d2RlvBrdQNgZrdG5ouJwIm+UAwg
3LzLnXQ7b+pvCDaTzlpz3r8OgiFNQ7iHgZ2j+oTFQOeD40+iUqbBiEdz0l9o
kAtBqe3rs80dPY1mAew5sOq77/A4Cw1OrF3uUSeh78Rlw4voz3RbqI2afLKP
7Wb0S5FRj5Kg8VDXUp84h0U4P94kg+dMXxPFCegcGhqB0yrMtYbe/SgA2TZO
pKI/fodQpesZxFSI/fjXsBYotPGIZ3dai6H3vuPQp/9RYRciDlXTSgHJIuaY
8G3Q51fTKfTRVPWrOM71rN+6djXI2BnqrQdbvUXsVpFtm1Wxei7bl7dw0MrB
qKhxDIPbrXpWqRJsteTR/hU1jQZr4MtZyQobieuYfHWNmSrcGinBjRAE5x2v
Pgo+exjOgMe/awjo+Jd62RdZWqM5ZnpEssWoSpv5mo5DBrwm3z4ok6B8L+/R
t9WdVycfkFPIBxTIQHZk8BybkgUuk2xAr252tutzJ1T54+ynLFNTT/7x+gyc
m3hT9YtOKl7TTIkenMHKmqMCuDKKenwKOzMDdRnDbx179RwjzqoVWh7Tha2d
qvbnx8RxNou0BJh62WCd+GmZLETs5+CRxqg/gaVuxoRUZNOCiEcaJ/tJjkGf
5/yPtYglyt35KlFREV1MwMnXtqiDyElpLynBcjQaf7oky3L/XuakxKqmTj6m
3RKFcFAmw9d5/pYxNPU04f1DefWPQHo06AYDcQHIAPK9gX7mgVygINr9Tgc1
+IYRWNW5dftMQNxNiOEddHNzkAUEcLQgiBUZu+1ubdhzA0YUhImeVSuyG8rr
X8eQFzMiid4GLlK/UDl/9ZmZdT+RYpxL1e8pmuJuiVq/o7F2ffQQ4Z84FIJd
j3QwUnYj91sEPm/RYTTMUbBYISYKf0tDWzHcjse/nJFH10Gm0ZkmBMTKVjLw
MhDaCXOqsWLgMbrpfuixyTtl38FfaZdex8wYZ1vw69KTSKbydPKLlVyX3qJI
aM3ISCKcsiJavtiFIg1hSFrf1mwu/M1N5ht00FiDL+0HGdOwFgUtoAUid6Wu
dEefdLRF9AFR4sNUgT+N9bgWwpjixafAMCIRj1NgFFUb9aUdqxwY3ZfSkuU6
znvvWGNmlWTxFglsWhm+qhM0lGlh+tqmWOvfe55kJeanVOl99S9Ol5qZX06R
F/jc4YeRpSGex32BpFaGL61FoJZpfYQrdIAhJ4fFRbm1LP+R8FgHuL4lwnVb
3yZH8/xYFVxt+GP951d4qDjg/hFmxpth0lV+mUAVolDmn+ql3TbOLGyn2NBd
srECpK0sVKEk1XixwS52YNPOaJIWIl/8FIuPC8BppL3Q4qP+Etr9SeWQKdts
YO7t8aJunLp3CJKYNW3MoAxiHJCceYShEAz+Nk1p4AIhQJerSNeKPGgVSupK
8UIouOtpuI8xiUQ28ziesQ2Ak8TmMzc6hfCu7+1CMN5D5HCqiOo+QREyfBc1
YVZpM0rIGyV2i7aeVoyPSLKS2Ij7QIViNAe5SC9Giz+Aw1Uu8ax1vrQbLbUo
tpvHkVoRH/G++GKA2tiNYZFvjpKAAKfJvyjXwUycBnswkP8jxbx6o5fo0hKl
VplKWAoWXidHddxJ0lxEuJXuvr/IVpp8cU1EktcX996dz0XRmqfA0OjVUPmO
o0kThFxNJcRQ0MqHPtjzPPrrWjZRkMMR348l0QxD4v0x1CGnZFw8Di4Re+mJ
ko/ZSj5JmiQhL125WHxPNjiDlyzPxc3G9Lnwa35tmAipaXXx9+rhrAW34Zig
4JI2GEswyG+n5uhoRZ+X18kxn0y/ux4mJRVc9XcfgZJnVQR9kIRp/voDfgwf
uR4gJ5t09Euu/bcH96FnEeToOu6cS7aWgz6bJuXSEdt3Zk58ZtjE4WZ3+uIY
+aYPs6l5sAIfl+sqRpvwhf/NzWA5YLx+qYNJT7nB6QN08V39dvWPTW/gi96o
jRWTtNOMtJ64vHDVr85Zm1CXCzGKUuF3pzNVTAd6R2vH1+fbhdtvM9EjCwNb
GQNV/lTwRl+TLnfBsgXix1KTA+aXeRCEIX1CbqrUbG83y++iXB12VPDdYo06
hhL3ijQWIHCiY6nYBDDT/xRTuGS7t0QP7BZh2/MdjMbLReL2Uom8g5ygXLRI
IMCG3ex1Tjupmute3i/YMO77dmQ5uCdlJZ86Ly3jWSV45HHeulkOIEjM52+T
krX4FfCYKVwkia5SDgjo1l++CU424v6OHwW0utyFuX0e1G2Sa6LPKBU85dqD
AUmyV5w9AMSlcbZgENFGhpVRteY7rdxnUD/JUolbQaeMpQK4IVXJMMPNnou/
dMf2PoZ5iJFE4ke3cRqbpg7XDqiRwV16IhlQOIa9VdgKlzqpa/CcLhcCxx2l
T2is8k3nqsAlUBA8z00jmdvxStVY38rNQKqPqq47sZRQUw0jLwSrMF2CayNJ
DbGg9kWWIxCmd8QkGaZ4as59IjGMtnn3Sh8kqOKt9GNe0UoR0q7T4Mg2B/xh
YW8viYC6qp+Il37X0o1/Ir1GMJxuz3Q12FAsRdSA5Sb9I1Wmc7/t5zkoRX+H
ZYvJapFFR5hPb3AgPOszapNxoGacxYN9UNbiD88TLY6Y8G7thTNfwOjn+ACL
IZ80fO6tyNmSgAoae+lWHNmz2NllSsTYzJOTyX0RqUncaHM6sqvj17f4YDwu
pRHxHEHV0QwK6//Wgwsm36uPecUVS0b5Cib83Kr7apmCNrP2uVWVOq10uPn6
ghccfnyfeKAWtRuk7T3N+ryZ3oocOhQ5DHWFvilyhAl90CuKfCjwuxkPGtP/
xhBS/RdGmNmpEbL0BW8kpXtK957kT4T8QMWRsA+FTMV0bVNGyi60hUmne+Tx
9+m14tU9iBuMcKx5qoT38BPSiE3wjHRhZkgFIzRvmgOnQP3RZ0zVLnYi2dST
gCMABVkMtxvG4kwH4YMQVn44MpnCKptskTPcPPwbgWS5nz53RXAxeWsXiQRR
ZT65C1cmqHG6noVoNcxAzL5s4E0ddsYJqdSvyCAXCemivtFwLJs2wlXnNpf8
v6YKBOCWxLTxyPR+hLPDLxJT/MMonPSTrFAmfTb5C+YMnm7N9dxpX99fQKzA
1JPIa+YN/gaVPnDi1TPfBXzCegU+F75HilaHg5GddB/LVCjJ8lbep7MJAJrJ
YQU4pJXw4qGr3o1UXmf6DP8qUfK2KCdPN5M0mBTcor6HpNOpuNmhGkZ2lvwQ
HdH8RifWjwtj88eIYy8roUrKyGB+8klNicq0BZxt66XxpTYlph123bqBSXdy
oClxMSgclh02yLlmT79inPt5Cb6EfeMOFYQ28fuX0zKdVMQp9trMcC4GvGiq
RLgHktpxliPWjbcml/qSt+HkhSCUltuklgDWK4GuKK1A7n9ECLHU6m4+SN98
lEfajgaPMlBwXUl5vhgrmWKcydAqtxt0b14Dm4QpMghALRUjwTZswAdSrlpR
bduBQyOJVgp6VRqygp1vz9mY8moAfb83S1TDERevPalqKU5Ido4lQp2Evb9W
ODYGAzb+4G8cMEA/yWQGVLjrPm7tzR6610Udw80xIb4Z5zN9uA9zU1Qv5fiD
CLg8YBvaQjaEXAdRVq5tBGSJruwnwhqf7iSgQlZSbYZoMv0EzJfii3Ryf2LW
iezhvVrsgwRCxms6Jh9nWxBZLosmGS4T8+Dl3ySCinYRV22BDLKv34Ny2O97
IZ9KZWHmziDKqrr6Mur9cSWFMdQplJbP6kcxpWjvR75D5lXGpNFZCdYqb2ao
S/lrzdAOoXxf7cFjTeg83cFKsa0NfiqNFKY6Br8oMQ0ru5wOVs3/BQeBArE/
ez9ARraAomRe5y/M6IUqU44dB6Zhg4uXs1dJ5Fuad6nScoH5DSHG7XH1nw/T
wuU3RbiVMVufk66VmeIImV2dXHOLne2VJJcVUgdr/9Veha/JpL75JEeaunD0
+QV6sQT6qSTq34NpRwhxl2wx+KxS6Jx/mkGHZMHzYMsUGN1JtWyKUT9/uKK1
bQBCQST8xLoNLCTicSNlSH5r4LkhAFC6okNKgLkWQNm65ttAKU6xlXwEEMNe
gb5ulA2myH3CDsVH2EVMGz/czO4w4M2D9BM1VmOa8ia1kcxQjaI9WayK2ljG
F0QaTWD8MdXUrctEadhAc8AtVFMGHUYMRA6VByaxjd6GlSyVKyiNRP8I1Bip
mn7E/tUV9EvVZ1R+dAXUKNJ78gLSiP1IoJcC+vi6Y87dP9hkxw9rWCTrXwA7
4inpKbMpWPCyeB8y/yKEMrU0qYK7QhUxKG4S3OkI6HBWMoRt3+j8tV2la4ZN
/nynkUtcu99rjoK9AvAjSg+2URB48/In3XcrM1idR+ysAxPKg54EcekFu2YF
f3w43OtsyGs598/fN5bWoEFAiT6vjkZ/GllUExNT+wr5ZX9BMLR3rLynz/Ni
FsTtLk1jXTLPuh5yEqT9FryBU4sjJ//rlMQSEBWslEJSJ6ANnUrEO1REUZ21
JQcDhN+IwJNeSBtwdRQ6l8dDZuVGBRjwFj0YfTGcHtHXxd9Pe102S3FCSjt/
hS7PiAr34LOtwQUpXS3c+S0PG3d/nj9Xpvu5mYQBovmnY5zOP7+sdmcvtAoD
yCJ3giGdBW0foVLxdxdryLSb6POJpBNwIUBeWTXbpH8TSFoYFIizsv8ZYcuE
50TMuHiFWEgPhheN+6Tkhup3GUol6k1nAP4SkFbnmhFWwlf1D+xAgrFY1T78
QfEDywTBQdy+vU0/AzwgDJYnn0D+D3Fr320Z/W7KRNU6HgpLOf+oaWl7jMjB
yEhcpBH7WcL9WEnVxtTCqyfyaxZa9FtC9JQR0tRDvXidQPrUoenBhJktA+Kz
39VQZPQb5V6e1SyN5p4MldPRmT8MN+nYRNl7r9Wdz1Pbgs7sxKoNFHp2GLgI
6cDlSUkEHchLiN9dLz57zZUfowbPJYkLo2fGkDBUhSispzeoAADo1hafct5v
Ig3/o/lwdUDVLhXT4hLV386ZvlBg9iSRJf7VVrDoYqFKSx0+/AdxHMKsTrPv
20QAMiNnl/pCk/Q8jmWb3s684iTj7tql112TiieLFFayl4/8CAzEmUlPWJxP
1/0dtnBn4brCQPeE3KCIRGsN/ZvU4SmsmlHF6AWneOI+wtxf+MsnrAb2qQ9M
VGKGBnCvuChbgUJC37L/JDukFGwhCngtrPhLvBeUa+pE9wDzeMwcXWHGbvAr
f9j+895LlbFw76ep47T/+vPm5NBIupq4S0xp4WAxcCoZn4ui1LOhxJFafaVb
Bmway32W0kLufe2il/Dtp0zuTXBUELXFCceGd/DiAXXTrz91rw8mzt/9jL/h
n++U92Fw7a+hgUHjwEJvhpj/dNJLQN4TipHC1WRDaVUDyXpF42cSCRWTy/pY
J5490RXd/NLFFXUwphXO2S0SkHvvxjEFvI91PPiXPDe2mwXdmPl5wr1rDTzN
tWqe3BGGpx1IA6FH0eFP/9Lsso4OFeWEAxk6TZ9Ll2zBmej9s7U14LG5RiZN
xUSefpZZv5YO338gZ1m4OzytQkF5PiDL29HN6Vzo9CfbvivekzAmdWcHG2I/
RiUxmzUyD/Y2qUdQqtB5dnE1UNETdYt5FXrSqI2VIvoC1ccB2JH28iKQ/srL
d0fWud09w9A4cFM674RJ5xJ9cjZSvzPDlcjGKc+Eq4raIvjnQr1SbYd7JN5g
u3zHMF1iBNeWfn9T5S/1Gp58vWjqvqrvkh2QSm6u53td+eoospPyFYUF/cfZ
a7yuHEQfCGvGEf3GgsldPmXgR/Cf4pRgesE2R+DjjB9FTRkIMVOaK4qJaERq
GGbkkJ7A1Ao/G82FW4fJX1pqfiw9klMxDJXo+HdFgHJ2nqdaYopbnurZhUIA
S0YKbeuBOq34KlPGW/00TlW/LuHea8gkCbgoovHP7fxH6xsbK3OaBr/EA3Xy
/voOOG0NmshijOivPzpDBVq7I34yeqDr6nUcQj2BQbphhtMDL5XQdjangPb2
B5PLLpm2/UkNCT4DabAUPKxd0jqvlqe8Fghr7J2rsx9l6gtHIBXrM082Nv8U
L2n/y91V17JtpNEj5x1xLq+KPpULV+XxC4q1o7ByDZnUlzWsJqE/0mA9tL/r
1rzdZKMmZsn/ZjPzHcypnfLaxkDbcar/kHYNri6Y9jXlXUtkR/goYLz6nS5f
A0IBGl6jsIym6l1gccxvEPLySTKh8uusOT4keFNMG1ODqyOr3yO6S7nA/Hf5
Q76iFz8YW8wnDo20FGhJPFQdvDiIDdwIn6JlcG2yy85yrMxhPszg0RixnxVa
pJclZZRlqy2SeGR5slxaHQ1KI3dCmoYE+Flx8QWabNUCVBlipMmOYUSGB3Nl
7YiXMIl5zQahGvxoqNkL0yiWP3bTyMtZ/+rZBGLLushdS0/B+1I2yMiVL1Fm
Zt/QmEeVxXFTjhGxsLDn4R8GPPDbnb7ZjDT4V6eKmwLkGSkoyxyPLOs2kajy
0pg0GWrpIyr5ViBqFJr0tww2IeIEpFAS/3rQqNiYqcdn1IORY9xAo5fruJxG
j77YCOMPQRzNRGR2LpHvwF5UXc9aXtl2U1ymQR0RsEUg9Oy3tCxC+Hc36GQX
oY/LPTKtaJOhAHi3mZtoI9Cgrwmp2s0QaDlXHZrHxO9FRU6efwnyTdMFtJvl
o2BgpnL35O9Hnnm2pb/lKq8bzXynoRo2wiHqqLEBTHwyEKOfJIBIKdmzbKhA
BkUguW6cWqi6oOLyAWrBdH082F+By3+u8rNVfLrdnXnmUiRue9kcagMWZ5de
jQkYNstpjJDTtzAfDQBs3E3zi9DyYewRvik4oRl/vGxsTufcTcxm2ZWtS/2Y
ANaThPUzgAie89IGV38X/bHi2NwHJIL2dpU74j8ScKPmb/HyhIWtU9wQ4XkJ
OxDoJaGFHvEsPlBID5CEHJTAecIpsgIRSpfg5i3RisyeTqe80Y8wzJl/RqAv
zgAfI+wDMLuLJiGp8BuVNg70XmBRn4HO2DB3cJAMiDzIWCWQLqgLDx+ow7cw
/4zfMvePvh0SoCAcoJ/ZxlwIjqq2ER+LdHZq4XAM9lWEhOkf0Qz3DCbgCSK8
23ezVRRCt6LZBtDQrIvRhRWOUftRhovW91tlPrL9WFMRnHOVLmtwleK5eYkE
AQxUq77TbDv50DcuVa8hpxMAeUtH2dZbpWNyYnATT7oeTc91MgsO8ZdIyGL4
bpqmev2L2naTa0S6S772tR+FGx9bA5O+ibc/Rv8XRuiDgW98Y1Tz2jY5ariJ
t/HYUNP9E1GGOL/DHhqEvC+E9YP8d0exqXgnLGRyFanNDordP7IQgn5e762E
DxZWnWMVKpfIIttt0qqvcoToKjDD0lhaRKxyIIf+YRMpkbpD9BlWLGtOAcmZ
gIvvpey2/b6xTdiTUB+VQ/h34P3Ok7FPdjJou5Fcp8vgZJpzOiDfKzB5YUFO
qiN5bwU3Owty3m/FQY33KO/ed1UHt3DsnlMkGbksU/ucSfaXr5R9XT8MtqJ3
yZCiX94qqPjpu/4D5bRMTZ+wSQTJqGHhyJ/sTmHHZZBPK6z0v+8W4cjrNO6w
qB7DuPLNOXQ3wU+xZdVF97ILe4FOMk/tSDGQfAisOfOpVLeW0rcdYg/bGXrR
kLE4JVylA3Ku6FTT366G9MUI/kpozeg8itt7/mX493e8AXO/9Uk7E3y9woaO
Kzm5XLnzVIkYMO/r65WhsJt0F1IOZWA+7TpmATNPb1Xm9vJA1wuY3BYQDhg9
fcKzKrGDwPYRZXDzdwwZsx4By6+dFovXdw7HsEoVYBBi/rcnnpPgZUgcnhDB
emqpMNhl1gMkPLDySvqGN3JQUKgoeesQT0FDkFqXnGnokdX3kNHXZktVlYm1
+6iZBjbGIWE/CuSEPz8/eXRCbkbH7ovPqQ0hN8ewqfXn6AKTO+oPq2NZIOtC
gjpuHg9HgefBtHAX+xHrMpJsfxCioAdsbABD4Q126M7KomJGINVlMTuQf7Sa
45hMW11bNd6V+U8+WacB/8rPTgKgCie7DvOChf8hLcPycpBKToaw10DaLrOa
y0H7u3cl+cz+eNkpMlp3X01HZvPIt1mnvNbQUVO1WvSUOxd25GZcdh/OcvGY
LiNliCR2K0tBhiwa/j5ej6C0IfkUsTUR10R9UWsEKmWe5ybY/1tJTRAaD1CK
4HwaWxNufew/94g+uVGbXBUXX46S4au/5uQfJB3aBpAs0YyClCQGn1n5NUcR
EYX0VsRZeHZmWVdxMa3qgFqE3/GImglJ2rgX9obIJfF4hHiByghwaySE5jOL
eCvAVoBmNaJQDqTjjChS0AGy7qj1sUM23DTNDAqVT5hNacDBhsDsNzM3uI3J
WoFdI7FnzTBZ74T4GGCeehNhmZRT+leUUanIbMBz/T2sF0pbrXqzDfYIY5XM
4vLtJyllDl7QvvwtPGiGhUZFYvJ1f4vbvsVGf5lT/qY2GrAa2vh9vr3sAzG+
eSBSpHMSOMtHtFWaiy5UA3wqHwtxSa7N7vXMFgBOUSiGRYI+LofHLhrmAXl/
v9phz3BK6l9PWTwQ3/HgdY1Dz6HTHTHhczBl/smRL9tWAeZqsap2VSblmx5o
bRgZefR9eeBAe80rRBEc3Rfo77F16hIu21HZ1MFp7sOr+18MocE/i6c2DnUn
k5oBIbhlw4L25GxlePs7mfeZ7Lc0fVTi1a358CvtbPDf/a2qeQbn34IjUsZ3
GpxHFlbtiRUKmopXBU9Z4i30IuCkoImoyh1UzEd3NZLGQAZ4GLp8wtuIKje+
f0zcRkWXvFiEF7xtRaz/Q40Tz9jq3zlcpSDWKFux4AG07+kuj3PSMpXFchb4
Ww6x0TKWo+fsI/+3pWGDrkc5Vrla9I8Bk9VlNRh2Uoak/Z92LZCuZLKi5U5Q
baKNEZm5yt86KazOtzCKemcuTSMwNgeY2kUAIVPTnVaE6WYBZtY0fmbe5p+6
ZciFsyXtMBWj7s7/lcpO4ewvDwHO8qR/4eeD0aLJAHgH/z9JFL9owBORGE1P
asRGi65lHRZ5s5eYbgkPRifnM79o/x1HroSXsy4XGzUZOIPSSsTlunQZ9gxE
thz7vv7baChqBfx1hdMCZq/izr/9PtZjDDmK8k5PNUfc88Msbs3F+J89agZe
svFHTktzbWkCaPK5K9uDHBNMH/Zo0oYvcSnMfPNeIYVafmhKyIwQMubm6w3L
Hk8fVvRhtlC4Ll7jb/7kr3xlH6FsPKq9jksl61a/ZqgoE9O0QEJGwBMY6YCd
fLSh6prt8dOK0FWCo4dTr7l2wOgPToun7vQyjXWp2L8D/2TP4f+3yBdUIYjU
fJzqZtIZmNJjlYrvDNOJomW+f+dzpaSbl93snops/DSl5XVTei3ercRfCPdz
RS19O/FpVoPYO3ZiUgM9n1GEcad4UUColV7R8+84Oz8+SRtrgZwUM8CQSaA+
F5y0S6Laz6ePqrpVLGdNmZQQcZNavXfBKWCgpOptv2JL2SQL2rKLLjf5VRH0
lUYMvo6GnH3HBqc69IkdWTbYPfffGsTnWmCy8MUV5Z9I7b2dx5CP4iLNuhuB
xQXcboY9FU+RFBs2LPiqMdvldt4LgxL626clisaqFnv2fm5eATIKB4YeXcxl
DxodP7qaJl7VZsBvXCl9R2L4yyRshw1Wp81cR2/Yo13G6OYHSCa0NBvsMqNj
G5n7mfgCoWwsjkm9N/SPVtm4jWOMKcvsUUTRkQKKnqs7RSXiM/tiSa1ZkYmJ
78qx+2mxaeyqsVrlHLYsmdqvSNvsauQu/BgX4Pr5QG72myWF8x3Gmz6bg5Eu
GEEsImJ2GFEtcZp24dF4+F7cYuZ79p86J97cAKJslDICav6OXpuX48EG1xdO
ZgmpYyjDGvs1U7lIvktz5B2DZ145LmzDnm5Lmcf0pMSWIk+nYWQ/Phvnza8N
Pc969LpCv7V+72GplYycVqAe0vYiBwLFLjhiSw/jV2GXblqaF9Hw3CSWadfM
3wCj9M1653N+arJDaDKZUTOZqmRAME8AAZzIBWwK9IgrS8tFbRyZ54ORSQYi
OB1B9nVFJ3+/cMAHwV7d5KaaaoZev+NKWtKP9ydmFL4zVHyVyoGKDrYpR5AC
W7i+s8ByV4+KMCZahwOk3F75Fes70wIUsf0G8RrM4Qga6XaXO/+MSWxtmk2w
MKv6AZgqEP9MwuWHbX8+/qsdqF/UfcquKToywRTpswWvsDLjpAv6+3iIZiCV
8pidexpVuW/fElDchdZJtjFZIksIPYMnruqGJrNN1q8lbD97kNLrA4Nactq3
Cs4fQUUWu4zt3orquVEta2676JY51H4US7VSUX5TVJkih3NkPrZoaDqNqEiG
yOlSXNYgKWn7ipM/xfnyzX3Mb8YhwoqANWDvltH3IUabz44LaE9PtghqTtR1
y07+XM5WHlf79kIVfQdVhwq5B0Z7+CorFFA1mMYjqLKGoSCh0OUrSQRtTGLZ
IVXtxrhET3IMQ12qGIKXlDoWmbTJwy14ugxPPCmcJ/XsIr+xwHlKV8O3aQ09
h81RGswvVuZJ1kgpvdgeJMn6b1DDHI27MaIrNlpMbNuusxuYWTcuR2bI2xCd
E7mfcqi87+a2Wg1h8iY+9EE3b3fyAHNKgfAXI/WOFsbMawph9W6l0sJQbBjb
YkzcZIA5tDz4ogJZkbDPnc/HBav+EHEeo6OQh0ownV/V5/XiJ38sinnZTBhK
DY0pSVjKkvpHbsM/vUT471ki2+fgKb/GLOzS4RS3501zKO0AOpnp0WDb+jxy
NvD0o1Rz6cB7EyWcBesCh8sBPa0VBqWNSMyihMI0Se4YWli5bg+SwyUmDK36
qkefNAvkbjc23u69JKVFcDY4SGpK9hOfmVcCHh1v/xFV5hE0qn16kTXdPg18
y8K1WCRVL5uEallW70UUEZ9yGMBvHg35OEjPc/SfrN8nmZqbvbcgziqmdRQX
AmFypqGdofhilELnw3STL4LsqcymEQAOOihhzx4vrWSiBuIDwXQovkU9k0Ve
0P2RX5qSnPRTclUIptSPX+ys52oWzxIvSeder0x2AKQKQ6JE1+ruSuCqF+Qc
E1h3cMCXHzx1Us74CuuP6TiIX3mdn3ctekkD+Y07lgr3OCN97bsoo106Lrx3
dJ1MXZ1RN6mjYjJKTcg762qOBKWH56dBMzwnWIKcQZdtACLLlEb+dus2u/D0
R9hOz/oZn7MNPcwO76PPz0gwDmOejZ7E0Lu43stSABoM9cYi8fKqZKVlM3+/
F0on/dxt09vjEZFn0hZwhi2Kq5pcsD+Ngc+D1n/zs+rzimHbrWb4+5NAOJ1u
2xjS/mhoa435MKAXxgzTBD370l3qsLQCWu0ZoAyxRw05FbGe1+5UeekkUl5n
VX9pPcFUZO4zewUZf1CqInsHzdzmas7nKxDEpK/SDk6m0FkBcR3Ofp+BoMZz
l74+afRRBkYxpwcv55gYPvK0NdqLYz9qFWQWHjcl6Wa64lWIjCDuHqUPfYCP
MB6GCcNkIKfP6e47wjofMkBrylwsb3mUDeA5/zV8W15pZEN2xPfI/VW0j6U3
37JHILt0UQbNko2H2SjdOVF3PJ3vFQDM9zyaQMq1FQSFxAfwmmyOVz49VJvS
BLaUkX+Wu/hccy2/TAB8AUIwZ4oOq4Igfbvp51YET+Avs1mCYkyjYbdt/xnU
FzY24WqjQfVCykX4nNOJ/amPBtc1nkvCfacgIFoQ+N3x0fnD6ZeUTI5o5461
XSaLFgKzMsYfbAwGzAOLygTpopLQE/iPeDq7eAIe6aDCcdosLjy/eYXf4vsl
C7vuj+iZBa+yg+Lf+o4tPTCk3bWWuULj/llPvMd4mquvmCUJp7v/dK6j8379
JyIKFO3hljf0Bx7Zg0k48W6gz6dY3R/PjqMFqJ+WclrrJ2yVuo7vq5lUMJ7X
VaoTRtcMwgUo+Y5tja3MO6W+40kJtCMwgZNBHBZZ0xD/BWMt3t43qw1QVxPm
kVgNV7WatK9QvryAxrGLbzoaGr7yhT+exJI6PX26RZIMU9Ow3KzzPX6dlB2U
gqrOJ8wWp0VYtpxu4Ku7B8mECC5BKcm729osJVn3tx+PuuzNH5d+cEiTa3j0
HYvLX9LTaO3mzWDnIbFkJaFQU5wE0ZGFxnSCIWUQUu1TCbimgv0kw1kCgZ/R
GNB/9Tf0TNzQtcsf9F4FMSDPifTMfnA+xia9x4AD3Hzd6hwpcegKGwkztCsz
zLma4Ln6Va+2EFZJy2MMnMIqMDSZs6OHz89Ss2gEFMfDEVkMSOKHrWNQr413
W5uXJE9L58oyUscVVtD18ZJ4+/H8lJnjj2nzhaHSoNqsjwxZ+tsBSIQo9JwK
P4s7Xd7KRLYUTsDYKXzJunHRRbjSqDM2RE9VA97PwPOl+7KJDXitR+1bU5fn
A1WRUgFGfv47bAXEgKmdIetcmcoVNVNsMqd7GR8wLzClPtY9is3GUZEW8gqC
Hf0HtJQYIJ0Ix/ewSquhNeLrDA+8okPrZCUnpxEk0alkZJzUXtLVALoPD036
LEMSpaz5R+/KZc/ULmNVQIjHyHyjUuyaIGfNoiiPz2hu9y0hgIa2AInFmOtH
iJeBAJn8aXycuM2X7GX2JLrlci2fhSnKKmTMABwRHroaTkg8T1kEfr2+oz5V
8JtLmfrDJklbt2dXGWQ2DoWSFTeaOqZTU8ckHoUPHwjKzOZyt/oUo3jn+e4e
RZk1WoBLMvz2sO8SW9n248UTYG+YqekKQLeUWAiHWFRdtpJmYhRVOI+AFLZ5
rYneWXlUAcamqC1H7sQ8/jOiXVJFhrXqZNBi/Sat7YfQ557/OGmGTLmupmB7
E4KaB2Qm12vRoE845JQh/QMHcIT05CjzlRpBwTQz9B5U7p4g755DDIQCi4Tj
UioLxqPXBbBS1udD5WqgHm6+/uZhjdB51ZZLzhdsTu9+RuftZc+hPgZayMUl
VDkTDDxjpUNIZUB8/RFsDXvkcEac/DmSsxWGhdsqxxQKO6JjfJr/EyW8Aish
2Sy67u7Ez0rF7pfBt8igLzRtVIwSDTqXBuylL32KJahybCLqGa95CcqB3UDN
ZfhKs3LDFLTsu7Ct+gAsF/w4q/qs9OwjFRhHfyB9o1x9H5t/WlvLvkxZlRyq
V7jNxKMQcWDFt913RfLIttExfVk/0ECjvVAXPbz8ZKC+zHiUkozESaKbVOW7
V4Q8XU3IC3afmjETl6zM2F7EgByLX4BZiSBfY3ukX6dETqnX0Fek+BcRd0LD
fJzqhXWJQRBmVPxrTAmD62E/G9j/xqpflXI33Xr5llJ21wzDwP3lZp7peks6
D/4pigx7x6la1qZ75YmUiW+OtaFKaH6Tk9ZfYw5+kx51JjAHtGNPirCGxPb8
z06X9PtbHsWXyS7uAxni2+sUpwjclWekbXawHe6pGa2WdqXXVnSFlZcE0ySY
pBfwGc1MmQEvZ306yH+/4bLSWUX4oaFW/djcjo80ch+ZAIXPCdc+lj2+XUon
P5T0e/ZNhaaV3klZukYL19yVPsATpozFEBSjKUjsq2z0oJj/5pPD79NETvaf
lW7nAiIiEW2B7y2jZ3Ezb9tycXUP7fC1I4slTYzmuOXxcAIuNVLp4bwMsTZ3
9zipJPFWZFalm55wVZgP7atrZK0faiM3AFSgRK0PMXH6Z2eMq7yg4q6Vsv1+
Fqlbf7DGCTyEQNeJ7MrW+rDJaq0TPq2HRsmDzPKH43IFNMb/C25of8m9B+ka
Pu+hgh2gyo+ZwEVHjlmAxSicl8bwOCfBJ91EUkroyKcU+QIBgtkz1Wtnevhk
jVIVtdjHIEXrRJ6gfRYmJx1QzFly6XKs/OpmXEwRHy4niM1BgNML1niU/1S6
X5pLgmfgkkcWhYf5ot/doGauO+6N/kr4oGMD9J7Yte/dD0VvE77PP5p9OTY+
/b6fhzrpWfDL0H+YH5It4xywzFAFloVe9TvqxlIxntUwUqan+L8DB5GHLQHy
pr87osW8PxEOOArGGJqqEGk0wE1zfvqOJLgJVy/PROvlXCgLAS8YvLg5oDoI
Hbw+Ow1umbkUGrF0vXlyFEnbMdOQqrebAcVeBiI2U8f1ZpzyLYsp8JrLquNB
2wrEru5/2lJ0Z3OK436ZFXE8TsgyTQ/8fpbbgOpya7fNaOElQyNfGGBLbfDH
YWaukNxS9ZcKYmvVFKkQ8pOdwr06hkqYb1pa7oyX0HoCWbsRgXO82s4Eug1/
FCL+yqkAdfSTkzVzY898XYwLjsrkXS+NjWqW+wIifFzfuwQG/rRVJbOtFsN8
HETJ0GZnv4tf0louArXc0ZinkqnkQ8VTE5ews3HuH5zVcVFIWamGzbFwmujE
31z/cB1MpFrLygVsZVmOx7Zs0KL/shcmiENdACeLTcFtwoL+Pprs7MhmT/8z
9rSSFuS2Yy2Eu14l8rqYYDYl1bYIdZU2mwJJvV38udhcI8E1GCfS+ewwB3dn
QBDDVHQA+uZ6ohJELUL7VMSAea5AQkrcn3RTdNXkIgXsVMQpSyj+q2kMeakr
TveXs9LXRnlKyujk2SZm6BPvggSbO4PcGbwcUBPmPuc2zDNZf6zQiLxfrJRJ
qMgf7job2ucDrnttASlyQqv1hPipLAB2C4+yQVoKYPCz36TlpFQlpt0Tmbbu
TxahG2FrSOF/Xr13mySKvHNGUNUAo5T7g/UEuldDxg3l6lHEWxNcQXHdY3Rh
X+37gqUgfIu/kiCyiYqkCqXMN2JmLKpDfRAxsnIsbgndvWpJmJy5XX6T9j1s
ZJqQXCn8N+DHSFx+xwWU5T7kwXMH1YXOMqDRBHVPf7q+6XkDJiH3yKI/1eLt
PhMWj0196iFDhzqkRJmp+4hSldpzaQkNKR26i8iTUrceKkdONe1dmxvN00Vc
82XLMuk97VdAnrmZ2ELSjYJVoScz72+pbBJpIkDUAHmQ60ZcBDQ58iK6eRa9
d/G+ykX1w78oZbKvdDsfsSAV5kA1ctDVMbaaYQ4wxxY4K3qBEfKev6SrqFd6
co67sC3b02e+aXRGVyezBJrj29hIHJyIBMITxFL44t42zT8fGFbZ1izkwGDt
qOtT5AWspcz9lG9GtRjJqNghc/TcwudZmEyBOnd5rjKT+BTj46TMit6pQtK5
Bbh5WF18ejj2ijVmr+O897HWdNSD0YAxkAL9oqiObTMAZBbrf/LW64BSLkoT
DrtY9anUdbFdVDRcx/hZmudO6quO0PNkMFuXtBax9K/iF9SJim0IRyl1CQn2
/by2TO8TB9n8N6/IMExRa7qFsi0z+uWNH10wtKbEXQoRwks09NZWOeKtc4ZJ
7vHqi++whTLSO9vVoCOKY42ElBNEdqxqzWlc8PgdhpZv3CnwVTo+pxE8/NK5
1CEq9txDXrYplqFzaPPEKU2qXKnPuSo011IoNU9CUJeS+BdBFv7yFtJC8HCn
DQY9oQh6dfvNlpbliiR5cCoo4jAHdWtWwNI93E3z1gb5wToUU/Wn2Lrt07rn
vdOK6TBa/vTrZMiFexoN0XhACjTFgm8lKCgzl/nOKQ/g2DzDDvOs78OmJgYJ
FD+EuidlTZxCTQZ8s2l4TqcT+VjPbtFB4JA/uzv+eaP/d5tGQQmyH0mBNle9
K7Zdw8eVIAtB3ocb9UzUkJuCrNpsSxNT6lWTxEEKjTMAHPTpxjxKS2PevTSL
rw/Jjc1fs+CPc5UOKFP/djg/bgPgr3pDiXMZYce2kIBcvwlwpgk2P/A26yvs
9EwK7XhBXthyaJUF5KQ8qfKfLN980epk1QgevyrZxPVkAT1eI34gYGaUBXDf
cfdk8RU9kXx2OdA41slYsdH+m8RoD9w4H0sWs/u12P6IZS/9uvYWtRRqCyRa
d2GZ8TT3Rc8jUcWSn/ycl1DwujQI7z+IdIF5rmd1LxXLYnSCOU7wl14IgQOB
i3x7f0jSp+sjMtWSFzROHf2huwowVeMX49vn3wUOlRIMBAGjOolwPjSZCiaw
21LK91IBdGn6z35UAHnZQpBRM31Vc87K4mRtS7F2RieDvr+88x4C3k2G5yhf
b6jI5usIsEwGeFYdQtyAxlHA/pq8wjIHmqk55iVY4sW6QbTQt3A3MY6HZQ4A
lrhKSiN0OLZkDbAyCx3IuFcjYaFsSh+y0vPIBRb/LYsSyqhhTV5LtsDRhtPF
NqMQ0HVM1xYmol4nOkNprE7OPigK4XOY+mChQODFORkfY5YcEMO3b+PijUc9
4oLzWkdtWUd9zTLPc/jofpLIC9nI5EKCeD61lDgh3g9CrDKomoWi7XFzZzHN
cYB2TJYsBORqPNBeY0NJDcX/sY5gApIk1lSrIF78B0XyuBlcxaUdPM5qaRRO
vZQoBNg+tUNs3p2LgGEKEsUjbtvkgMfFnqrjGK/kXL7HXqGJevTgmeFZM2Ls
XLszLhnBGa5YYx/9eGzZ2DA0GFrk7LE3Rfw1URQ1tiHzRYJcF6t36NYwgxtA
uGjYfm8vdDu/2r3tf2zuEvFFG8KI8NiS0uI9bB40PM0bw0vipAARmS5qj1r6
TJ31DBQxe0Td/HpKqyuGRhWe0/flCQ1UP3e/nCPChvnAGYoDrkYadFi+EJGO
VRGQ9BEi1ovVI4DBl5lxWJkppehlIGnUBnsk6L3BTVhl5u3eRtzGjvjnzLTd
5ZvqD6jDPPzVbFyd1F/XhiZrR4gVV2ulirJe1k3hYeESVyZPQcOb71SlXhpb
LOI4Zp92UTOuyz5kVhWbXYS747m3JEedzmnD/KvhEawrzd3ImV+8KgtRYVpb
2zHgyEnWAEstoEbmXPQuTpM99N24UaKOoZTEnY2Qc7VOTzTD+yla+GQPZ4FK
RrqX/GeFuQZaMDmeX9B5Aqx7+qDu/5LwXiw5CM5l75akSTudlgtSaDSejVln
wNpdhWCpiD0DtPG6Rn38LQupjofkko9wPrsfouFcn825GC9RJ4jie54xlG0T
8C5Gi1kt3oaMsLVkhlGEjurweYD689+erYcPYcmRlTfmvW1whY+iIhw/TwoL
Ed7bs+7vMql177kKO4Fg60HyUB+FT/DeU9zYGWwAia8mQTeqbcJO4LNIYNu1
hZAMdY1knrYC0ZBsa8/Bp3hesySXjZVzGS9nkg1vgx/RDVcK0QxbKCHMMU3i
TlNuQQG5zz3EekqDx0AFSYn/JdLmiVfCzeZO7b6vSCw0WepQU0h8v7fDz/G3
9acqcYbxZacXW8uEvOTr9jeZ0QDmaYKmyipiHibAoREoIPkqFYNcZBca9vTK
lAnt1z5LdjovAied2BuSsfDDyynruJHC5RdHV/VUpIvtniR8/4SWzs1iwuVa
gI/Wn/IxNR7/Z2WYUIO6WNTpQo6oEiZNTKak+DJFaWs9oPfd/bZGwnttqOOf
vb00xxId13gPhDiAODqkXgdYoECaZ/ad90MMffqjKhQ4i1B6PP5fCfGjwu7M
0N8k0h9wSeJR0cIIaHlz0uZaIWEPyPxr+WMJVIg77YlOR/2kM7STCYXdx5/x
45Dn/3SaAb7m8cqsNCa3KPghdhk/EzL/1EzFU0ZN2ekNBmpy6vtDATdLC76l
hhEIIlbofzusXbgpWoa/Az/KqBPNrb1j06Reg24T01OAP7Mdx/IK1Iq+1Joo
+rePW4rRFFjtN4JwomJLFse11r9dy5ArsX7WoDNH0Yj05BDPw3vH9bEqS30m
Gn2XO65OZgVZ7Yq3oK/ZAA9QSBkK12488S0nRrGjsyRCvdVc4SVpIeSPX+vA
fsTwCxyDl9ufae5LZ/maIeIaEo6AWshi0i9WoglVTKfqt0K8BZhPsii3GtMa
o0sx060zgdh/YOjayhXA7CLI2HsGIIkdNWI++Ip/UZODoz3yX1UwHdQhY2sc
8lszVmRA9VzBd2yhC676G8IB0ddLHFBJhVhjcpHILV0tZMu40bEAUztC9K95
s2plO1w3111kbP2cghKbeh1HM49KRVH4O3YigjLH+oDZiM+3YElSOlwxJgkg
usrdIlZ1Aa0LbV2GxZe5+uXhzCr2j6ccgTqp/4tg5K12GXKQfVF3H3k8YUhM
nQddr0pKXoakKeUEbL+/MHVnOVvg+CN5bLr0EfOsl2oc48sg6cdwZfs1MBKI
twtJYKInu0OdfJ0nuK4bhoo+/41vVil5Kpgk8xSjkaqQDSU1IH+Ij+tfJujQ
EBQWm4lw7fAYx6HP7rCqFsrD5UJCNfWo6gnbIA00JrxWlvwY/CQUbWHzYuCt
EPFKDaVvMsg2W3DLrVTT523UpceCIdAAdzrbkFn2kRIcQ7b5ZRwjuIzC67TN
u/xPNQispXyfXUSs/0J0ktKZNk9sVHTQYSz7kjNY0WRBuGJDV+p8JjeafGw9
xmFKR9R5kCJenA5hLsnJMDl6ilD6JIM1zAlVkgrnzWxS9qkYsQItHM4H3P7q
jghpZn1vqXZTxqbeoRa1Fqnah3mqMNuuSwcauuHkqIwpAoyVNKzjp4qCdxfM
hg4ntgDK04Qjdh6Zg5CGsIAQMsdOH1I1d6zp1ZOaemnCnRIpSvQqRli6d0ZZ
oeZfMyoOWtBR9lnZBkeWTrQ/OtgIIYQCxl+KDgm+UPvO/8EPjR8BH75Ah5Pp
Ty/yOqjgLyTVEX37yd1wV+/xBtFG/d4P2Z6bl/LEWWd9MRKgTbk6JJmd8Csd
QscT3j5G9EipNnQG5RQDBYLPf7cCyb1006Z6hCd6pa/0aiuiYHxMWi7/HAtM
bsaLL/Q0ME5JmWqnXXLb0HyBTRJPJn0KC9NRV8reAYEX7AsiMDHiyjcKmyRz
JV9tlDDTgo7c953HHzNvLyUUYDpNbQP4q/BvPHR6kZK4nAPpPtWXE/eCP8OH
odrMkUy5LXIR8Ywl6Wbp3Idz6U9nTKmbGEkP8D5ivcQViEOTI8LJqFlk8o3p
niQhUv4kyG+/buP0ToH5FD876OfyUNyN4SMTA0tKycYDClwOBlQ7Udu1+QDJ
T38lBtWO2L4QVFrE4NWwcp2LY2KglBALKBB8Z7+CaO7wuLuROS11l/HTZ/8Y
jMXLqB8mHzXaZUMond38Ti4Q+O78rAAR1DgoKQRZYv2RSQavB3T+XYgezEtl
YJhHk2X5iWkaO780QUjvR/RtGfsO24cmGD5N/YNJrss0osOjHU3SwrwZmHXv
auDD2YseycBpkMmbfvd9PP7Aw4gm8y2XAnpn3GSL+yML8mnkThvCXc6kELFA
Jcy1L+FkhcEoFXUIXbgYr6wJ+ZLTSodwdS5uUqqKJ2uKRaj4cntXzXT1oLrz
SwbyXI9jzo6P4q6nBHGbyNjTdYAOfWf65yu2+4eHxYfLW2lHo5GpIFsJWGda
Hx/Hq+MFQVLRkVdfefJ2Q0/RuxmRfrknLoZe4mVRKmzJw3j1rJN928DQDFrH
WFuEuBvp110VKAKDvf3CyWnW4MhwB9jCUGQ1hikDDQBcgSl5rLafsvLhSuwi
UpB0WvK/9DbGGlrz9mRGF02hKmXMJxZVXJnw7LLj+XlFmhktmV6W2oqO65RN
t4ah5e86n8hOxc9Ikg5ViFp59Aq/oQEmCX4bDepTDlJRuA7TnKNOcry9ut29
X6z6VsdH98uIGM1JSeQ6UMnoR4xleyrWlfCKkEZXy5J58iYMMLKAKtdWPcZN
RBT3MnmgtALPvVjNHdOoSyygg1e6r7bl6YeBEPPki5m0h2aQ2ILSFSleetQk
kh94F9xUq+hVArB1FTPrL+QIxZjrIujJFl8VSPthDcLUYhKpw2OrCPhXY4Wm
H6xmP8kCVHYkBV0OlAdH2RcRZwfCl+lXO8vSrLhHa26+8fowCIhXi8k3nSPl
tUhc0oo4ewTGp7zZO0M2lg/7hhtc9tFl369VEnvFMR/SY9te7855MXHX4B33
gz973Tu/EzZ165zcMRr+vfWh/h6pBLdGcCQz5gz0mJnMX5JcoTNhii+ueOlc
Az/06h6iXHtVfEL1IYCxVaqF4Hc6dXIeVUgseioQjrAN1K9wk8qESY6C31P/
NnfRI7w17C0sTZK7tQ9jJeEfsOmNmim6bOuh5rIFd5h28Gk2GcDsquQ3UxkT
PpRRV0f+PlCfQwTZA9Nf4Xr5BHKBYOxP3SXL8l+CzmkOxbPnOPQOCRPbgHic
hIH+cNBMhudv51rRTCGY0fjjfKXmFdBOjUgXbz/jQGeOhSIKmRdtLhB0en1Z
rF7yHIH+ktsz1F/gGK58FgU54Pf3g0YzyryF6xfK5IsV/pOoGAyBh3wTnVBM
I4gM4L8gRSCqb1WyEeer+/1N31Iqr+uY/qMZRX1RSht9gt8Xt8YHLERdsj6Q
QRed3a2zIUV7XzNQftltS9zAyTtHHMvR8/mYhkHZMbv/jdJ5D/AnbICD3NJB
4K5TrA/tnusqrswxApDAm9dhrRyMoEoKaelj57FWnYbB4/IFLwlwkL8HjxAE
c5Wfp/mN14C87rQrGhcwbkMKtwxmV7kM/p4PeeUjmPOveT108rrR5VSUFoxO
vGUsZS+5ZFzeA9gQWHVU6BZY9f8TelS0GkMGS6/OTGRAL++jamefWEsNYW5+
DBwx04bSFeUIT6/wi7YSknD8j0uqv94yW0xuds21nt70w/X7C67xphaxR5rN
b3I6DmrscKfptZ5pcr2h4i9PGiGHacwnJBm/u1a6iKv1E4Lm9eNqqzAyXFrF
7rUJHYd+34qpMr0/GaKj9a9liHb54aIPJHSmc35jqWijpSG8aSWqyPwk0HwH
sF+PCmzr5RYOfM8o9e1YEnB6PoJYNCnpJpn7EpAjVBrG7QxXctxf2MfluIH8
5Zo7w1Z9z0VkjBzHukLoqqDKw2QbnD9NVta/ShsJEDN2gSz70WqC4Ik8et8u
jkppkikrN1HXnc91PzdmRW9B31WMgLq+qpCxAuJG1tXe5AJ2ji0jEj4Lp+J5
RJ2jdXoj7bEE0hJC/y0f9eZsxFmTTgMY2sN1XhNrKbTfAGaa1rBewnMNLcNI
uKZu3qtPyv/J3fVP+bF9ogAn0gFNtgRYHCyNtdT2jrc4OMORAcNRTyOuCaUg
cqlQ/92lLntQMUEdVSDVuq6rAOHDy7zuzyiYRZLKAzcRJMl1YVqeF+SN1RN0
l3jW1kqN/4BgSQP6gDCYxr6Fe5wfGfv/uHRmpFA5amFk/SpAiAmNmdcM7Yhn
t2Ge+UnebQc0drgNv6T2yMpZlwyxDMUgNnPzuRbZncCtinZOSDcCHHezw8+Q
H4WwpHxlRDrX9WRzuADbySkkWNRfQLsVx2ivQW6TeKn+ISxkF+LSP0aOJEmc
puDBEBm9PRox2Xm7LBQpTIP6U5CqOFI4G46lyibn+FeF4nl1huYa/sXgzjVs
FgFKx1ujd3g11JoR2jCulGcsQCsjY1gJqS3FEBCrRVZchS/+4mk+bE89xTkQ
YhuCX+YOX01ynyMPnouvOyHlGtGU5aPIuyg8+9gH4dKKosEvHjDSut9z5pNO
0RS4JqpBDuMaBrOAxpwlupQ57/33DUniGa+hyt8S4FOkq5et19CwEPO8jMOG
xxb0vGD3/RsQxoqW5clMAwr6qxxmtrLbMQ0jlgZ8fkIhX9VJEZgI1jjLatYb
NoLiPfb1/IuWVZg68yvinUpw1SiESM7nX0ijmmCRxD9AAwEKrxq7W+ow8Red
qHeRMvr3kqUd1ILNrJEJ5zcOoLBymo2ExL1pbFat9RnAxRTsdWmWszb73a7c
u5MrUxHqxjdYtuT17RxNJ0kETa8zR6eVbpuSD8LZJ1t3wgzAwiZmY//cZ0fJ
1g/9d4c4/JhHMePXHUGDLZF3UshZTitwAJ/n0XaANEgNjcxfXOdqaNsDQSuh
ugcc3WvsFJPeMhAQTnrR+V5+HoeXPjV9hu5B5renTcZT2NWuHOa9M+RNLSAa
lehgZT5iWUazj6Uq0S+3IbL9Ldo+AAHVYZbJw4XpkDPHoZJrIF2KzH1pg6jc
/k1jt2AXswBBhMg45X/XrHflFsX2JM8W1bYwYNiLsq+RG5ahtR/QpU9P+0gu
5HWpneLepylVN511N2XPUcHsHAHcis+s8RT/SsnX0raCfQexoejhGpj8ANhp
QGJVH8cH6mKT2pAiGBIlMja0MM85V5oHFv/BQBZ5dW4COLo4RwGYJILSMtIr
GiBO/DsoSzmI85Yzrvn27CFvRGVfXkLdZiknZbTmx5bgupRZVTqp8NWuV0Pm
ewi0RNzdWIEfs3ma7VhNGcb5rrmLRx2vVVYBERll7QJtIJUxr0VmP9dIjnKd
1UYPJF5aTY4YWtejwuFd6wbICl160olKN+AKRsKd3W86om1oaKGZ3uatgCZ2
c3lXwXHDU8uLAUd/3sd/QeNf5moB6/11QSOgoKfhDXMNiXcECTIGC+Du4/w6
KlI8SMdJqq5+2QNDqa78Opv6VbEUkTgnMa0Ab4Y6GCc3hJTTqot9DpcPkpe6
hBf11mp+NaFBDSXFGPNo6rvzVMfNKJjUL3l2Lmi2zmEj8LTe9jl2WuPXN2Ef
9wTnunrK2hzqOYHBfQSMp52y+mN7G+xOYVOYKjTgGSv+FwzJxrREs+/Av/Eo
5nVaqI0SkFjH6+5tiSka42TXLkSJyhb6+iIXd9j+uC1iJpB90efFkqBTLvwI
LP0wmlN9YeryS3sdGJJeok9Dxjkb3kWOteMhr23BknBSygIghFhrRnZGdTOR
mTYN0Pypo2gKVOmriqqnThD8/QEJBqx51EFVlDP30hoWm/uIi0qYRX69kk5y
mXLNN8BucJwqUI0Lns6cI8r4yM0WvudWWyhEqI7h7J4xxb/f4ADvecHxFg4I
qfWwTee82M2PyuvQ4mRwfaxic+YzKA80Mav/SckVj1IjMGXmjF5pJbkR2qxp
qAX/QhtjlEPix06koHNqVMiTO15zuZ2ilPKWCgNgNPSdogkEad5oiJB9lzeT
IZ7jEHLahpvCb+TtabS13q8pEba+HM/1UCjEbh/8eKcmyDt6TnLBLbwDq/dv
5J1YoPnmuHzo2cYM8nNcjGyOEBb5q3UT5Ahss0f88UN26VNVTy0eUiGqXUyf
JXX6xTs1UVynG4z8ZAUCGx9XjDPxkgZrLovlkJj/w+i9yyXUyGeT2H0SwNVR
mHkM8AvcAt+AIs5Zj4FCCoMCTbp0du/eQSMbVFNhcglJpySFy9UvCGIOFsBW
8tImTqapz7VV3LRggU9l5pzRuuF7K8pVBzYwrw4z2FqbYRH2sMErYsXWTR/A
wUwzSn6tx4hjGrdUR4I4iZIp0ITsUo7nFJkSEGLENmhCgAuqez6wLTRxqfNb
QfPsBffd10Uw99wkVjBadai4Ogl0LIHCie2edfbTB7WXWB/WMjan6zfWMX11
DElV1HN/H6CCrNbVFFE8C7HhTtujfBiCKGTDW8+SHnbZB2/FjxIBnpG+cW9J
kGOOMQrlZoUVHQ5rBl04784we/QecThwfaAbXfypm8hgT7YdACDvbQqaOwP5
CC3F6EqvbgkMJOxLgwnDEV+pEKDpFqoeAKJtsh0PxJDRpjWIJF+wGWo/QZPC
5l7BaHgBz/F/pJeTnlcXydpHDGRQnL7yYVYcSIf8T2KoPFT71O6fhyXMvnq5
uRzksC/pq0OI8LX2XU8hSt8+YFNtMsHxvneTFjd/z/y+qb0TEbXjg+lFQixs
YPTOJ62kYY84Veub1Ta7lOSX0CQ4AjaCzTa2+ua7FKynNYN+E+k1Yuqt7J9i
sde/eHLkOHywPGdSpC17GovaNYFqzz1agm/jIkutE2ii2xTG/0pMln2M5eBo
46ihx7o72h3674QUDWV4ARx+xKmOAl4FRxsibUNtp6eHxVj+Q7vfkhUpDaZQ
zrRAm5gVAQtWn8/bMiSzZ40xpbK2BOJJ/HOUvTYk3EukUBAQqqi69lJxrDfk
nX35Wee6Quyc7RnVgEAP11i73gACkPmnqxOpymTgqPSFE3Ftq6xTsDDXcwQH
gAl8mDMCpTt3zk4sJg51mZUCz+nPhnPdSFFc4SoIMhUDrEzX9+uWpkgWCulO
PoXtj963MevjVDyicSFeL3Hj7j3zuXX2imAfDcqMyuMwfR0DyOlT8d0CHq2u
Xb/SSaLfhMMYXb6NFfBVOhrj8IUOA+4dACLdO2/3/HrwccL9WGKr4wWtaP8y
cqEO51Ywk7zD+Ma1DBwn0E3A1rh4RwXWmLU8nk4C+L/qBn3Dm7HxoF6Lf5SS
ZDTaErk/L9AxZMVUyhoAS4PZ6QQL3Yov/ZXT1k3Cu1QhP+s8H5G2pQWXaWqB
sN19q1+rOe+OQpoUFFxP1hGav04NF2yhZcqpfCAb235FduMZmPjMmm0js84s
2e46P9dO32WgFIP6Kz2HlWL12+Ri+VuqR6yf6dV1lVk+YTJEDzXeptQSIqEY
L/g0rES71Q5VtWsbIFsqpbzRYvrCvfUv2vZp5MPG4r6/GFOsTVzw16biKQ6S
GdRaO0O6R3AZUAnUbFI+BHjMEFh/KmzaHaQ3vAYE+BNaNd34N76YvMxuvT7q
m2/pDrx1oWUeVH+lhH4w1QbrZDvtIs9bjX8kYhIedwz2qb6KFnSFgfdT0Wy4
O8raHz7N1EO+jY579S9QLS3vFinbNSDCEENdI4IW52p2sPQkqL+o3Ne/Yk8K
DCOlY1wAaQFUtHF1XlBEu9XA8SFoeMimJnjP92W3vc7j1iHteVQNaAQ1qvjK
ldq7I+L9Y+p1p45HWrOQgifauvibAQFmKqJLZIPEyFAkLcXslrmnO4/s9QQK
5PbXGHIInm2PnelAKSTuZyk3g9uuelt1OWrK+Jc/FKU4jgp1Dc0lSrLOnBbZ
MnSokltEkLQ14fMUDm9aVKaLZFmbWmUrhjFJco+yalwnk+9Qx6OUu54+Wm4S
duRZU4+vXngzNE6XwHf+jWLDkhPorAbBQnx/AGtcli8vBd7vOh9b+t/oKG8M
ErGhLG1CnoGhToAH0BuD1pJ5FNKtR63Fr+BJvrFNkCCbw8R5eM0ogMFsp5eg
mugqTh/FNB9trBphW17eqEankORoFOGuyaXRkw4VwOui70HZ59fCTL/BnPzH
chiwF4yJwSjZnaWtWciNJqjD0nvMg1/ANGKaKxFlOs1eEyJ6LObu/fEFV4dr
ozGcEYLSXg6LJBelmYsKc2nDlRLDcvpLyGa/yPnrKKhvO9UP5jQe0KQiM3Hk
aezwnJwzTNfMxCvmlu/FFzgSzKEhN7IWoDFTZiPnNXECoFvDpmDHARhpfzEy
k8smAUHLulpfSiEOc2LeIuws34+sN7/1OobkwwrWP03GFvjX8CsCh6XMLWUe
3IuCZ38O6q2gcd++RjqrYz9zjN74adUBkX9mIiX7wxnPZMHeMIPUE60Nn6Qe
rsy/Ztc6BUKx2NLNXobsR2Q8InLzul5WfhZy1XGTpSpmlzmZLBpKnpYHU5ww
xixGN0+FPYHV2/oMgBxJRzfCBBY/hMZ1EcrOWInhWAHaxntRQV7mjmfGlbc9
VMjRIVkVQsjinQAwBBZSH5eo8EoaHMHL74RgFC8P3EfEY780DvVC22vbz417
6GqTiKnfczlxDq+H++tydKVlnKCJvo6Jvh2+lMI0Rn753CjJgHvmRQHJDVzE
xSFlN0v9eTiNYX/XpB/DaTq0Kmbh5NhslaZCwP+6itPQBfxDjlDkq1MQ4M9f
lH2r1Tsjn4qRHBT41fVkXh4451ONUWenIT4cx7+7Q2QYo5G+Xnv1B7ojoGrl
GW1Fz35fCHsGe6uQKKJ8433AxcSxwxmoc0yhqaJ2/QhImkRQIFDAyyfxrIKQ
2DOtgehPUFr2evsOu3+4PICPT1vXsbna930LeulGCIVPRb2Z6dzwmLYH1cOP
yj0Hf8iwg69sD5D9cs8IKaqWJOqINaiV0TRlj72Go5fC/0bGWGcX7xxJQuHp
P8MVoyLaj73CeXwfzXMoadaeDmymWySyRlEyvAIVX6al0822hs2nD1YsCr2Z
s2g4hRD0fnVBtkF0Qyxk4osTwhQNWrpN4qRgdFaRXmw1g1agQR5JB51otcbv
1d10tqfQmHQl4ip2pKvH4zex5FEUVlCKsxFXI3rTtCprR0lYSaAHS1XMt5dO
isii3+orKvdLri9hOSaqRu8dC7SpC63D8drktm9ximy6O66qYQvNhgZVBF8B
9NraXMQdcQ1mSvk1NWaY2vXM4/Z2CvN2LNLo+gHMuMRS3wsA3gMa84c1tG2B
CxVaPoyti9+TfC0ljypLuFHP7XnJoweoD0BOxIxAI/f+tqncCEpAo6rKZ7pG
4Ug7Tmig8l1JUp+V+wdnY/NrppkIeO+LxlGJzAHt8qLDqG+sbQ9CvDYHOzq5
j1K7M5EV/2XPmE2q81SUQ8t6scSp0crhik9clmojZzqjVNyUVOpsI9q3Zpuq
MMkfodGgTjwD6pWm8nhDX8NrpdncZg0TRWB+mIVLvXL68Flg/DQMrBEms3Sk
tcf9i2WTQ0DHtBydnR8jIX9s5lsFwEujPuwEMbA1665LvmFLX9PihKnFZn/K
iG9ch5Mwdrotp3YXoWiaKKmHs1Z5IRw6A7YcNQFB1JCUZi0gN8mF8ROlYo1n
jVyIS+lapp2KlxjHvGaAo+TiJmqRivh70I3siQtTafPYWoy7Ja0BoKAQAIW+
MZCZuLOwzPcVCKwhcszzV09EgQ4DdT3/6hXYHXyo5TZH+GJ47BvwglHRi2Na
ylDakFSvtHzuQUulALhVfrKGrbZdZrO2+HrL4+CNeuhLv9ZXxpHZ/BGFsU9V
4xueIzlD0Lc3g6vi4L5a6sFHgH3xy2hv7VGZ5wSwhG8YnhHZkEt7X+TAEmN1
V4BS1bpsd5WEbXFyVniiiSK6IdyRDbC+Za4ESkUuQg619WrfqaSwKU3WQgBB
6ONiJZxNc9skp+6tWXiYRQAZO3x5T4z62A0yilZkhegi9F+Og8IjOwqQw4Jf
g2HWCdL8VRdR2YTkOeuJobUGH/KL3vtnYuUKWH8X14t7BOO9lJAlEArTVFo7
ElqIf59kDhjilsNti69hT7q8ddmfjuG9yUssq1Bk6UNaJOy/t1yoEwZVK58V
WpArwe/ZoNUqxv9FGaihj/8nIrMGgzoJRIHz1FujxDdFLmg72pvFcieebKgk
cFsDIZuJTFWpTspXi+S9ldjc3NJ0QP4DIRrRE4KY8O/fo1+XdyiWaFcaYiwl
Pu7wVp7BTD0PfK2JFEmkhFEjOYJm4xXBxHVvEMbV0lrA6onlgn2Ag02U45Wh
Mr3zhlq1UJsFzxwJpTh/xCd6rAZ8vinTzZc9E+daGo0dypTju0uzu6Gt6itz
6c7F6hS/DCFNLJTyJk0sktbBWW9Yxgjj+0QHFtNebtligHsMOlgFp1l7XdHN
vGpSnMI0dU9E5a+s35QImqzxODxhKMHs530Sh5/EXCx7rgLox85ZzNaBUFX+
ix97YMtSbFlKNdCuWvgzcNMEIP8ljMhFmoyHF1mudBvA8xX35117E6ZuR2Im
vRVhupSJGol9BD2xulbMkK7xgmnfKVdVmKbvri0iSX6aqxJE3/34g22LAlZQ
F7LNPsmDlck0Y+FXmljByj+htGm8e34zfbeHwbk1Gs0h1ebUkHcoHvb1sB8c
ARMg2Rt7KJoW62iESXxVC1HlEY+F1vd+4XbEOdWeM+4BelMPkTJkUdQ7Je2n
UrxWaeucFFI+UNC1S4yODZ5ZFwl7Vn8vYXRUC6IdHMvzR81f0JW0yQZ5mK1O
DmoeXUHzGMM0QtVETBhD1wUYQsaUyiSMpEYT4zZ2+gRok/kHvS+daV7U/S0e
DzYZtd5D+dyXNzWuGOEhFjHJcTkSKAaTeXELrQlSlI1gXVOw7WJZQNqqDTxS
G98MZuP67larx95Pgf45PbU/wa5edTfWBJymuSifB4F96mfG/uYqcJdk2ksO
Eyzd6VbWRw3NEkWUIDUVgLLBdTVIaWij7Pr5CgUtReGVjx1alBXmsZ43kx2+
/iLGz9R6/59OvNtll0e7KI1mpupwq8NLpKwrJiSTbI3VTylZ8gwFGAhbwC9H
cbvoMryV4qXPDShQrdaRsmE96H3XFEXkvLC6WxsgzRPFa87h4EIRp4xdHenp
e533Z0QsbQ/hG4WvSWidMoFbpvxgc2Mj8FfY3piDluNE5hMTGmtAyO/WuwQh
zCk3mD7Bc9m/cH/XiLw+e8utcRhBqxe5g1DE3xxWIRvCGP5y9kbK95Azui1W
t0V5ovMcgPkXV4ynhKGIqLdo2Hnm3Oy8Cd7f4H50R7n3mWupJ4p1nvP+/una
kJvDmk3TzXPo/5fKkRNfgo83dfvHJwkYqs9stamWuw3vdimS3NnMZLCzdQZF
/8un/174tWlsZ2U9BFo4me6pFoawn84iRHMlxhr+qQNsq2g/8BgvB+EiO16T
LBUW1WM+ZuuhSCJv7cBKhRJqu7d8NsYjPLxCFHmWWCCEzt5VVDjs3lvOw2LN
CR4bNzfKSvudyXTUglnNo5iHWM1Hx9qm0Basi+FK6rkR5KfQBqpJOpjvv5ld
dCkgD87dH8r3vtNwHBLhlsMB/PyP4lXeHtu9sRjnqr2nOcUfgYp+TGd+buQN
hhFRk8zMTdnsMWQdcvcsvqnXhHYK/omuKaaneWff1ACaH7tt59PZV16sXAYp
mhD8dleeZq5B3xnOZnLxbMkcKQwUDywi37+Ey1koKtpr1c23S2Rp2VQI7LOH
Zr02sZBIp9xTo6f54Y4N4AOg4UiDouJHmbxYbWGH0nGOYXSyNUAWiJliweVZ
tB2/FS7hS2KxNDJpMqBa75YWvIikxXfp6UeoF8hMBKyTQCyz7SMdM1aqXFF9
yUqpInrpJoUHtdhvCSlCLHZrqFQZIldx+qgE4hqyssk2iXXIClwsWkrdIfBL
YDIDML1oi8pXjHr+k8GBZbDAL+uNXzJFQm/sFamHCwNsCpyI6RqNhEnUrfI/
Oo58IVsFfuhN/08NIDMIaLaFFK7Rh9zKrt5rx8wLnnaRbEI7b2hg6sFy1J7g
hr7r7WDjSXN79Q6grmq+mA8SHDS8oSwdQmW8uGDlAY/1CLpr+3yKNkrSiP4g
sLi1Loe2kskuRSlKnjczOhFAgVKAgBbAzahlvstZIKjVSJk+8acOlbQeHp6F
MHt3/sPHeTTbxe1E5i81wCFVDVntzH01zX3cQRRsBEDpMiDWq1WptQJQC8Gd
+F9QTTEYaLHmoszKpKXDAnb+IAvcaXcxKaiDX3omWsHHBt17iH6+cCw4YUaV
JWyM0alxTUw/lfIcL2uOl013gU39gLOeIbpiz1lahsuqjkq0OLh/LA9zfCuB
HPnOqcBpEw8J2fQBfsK/gbEVq4xQI1Ilx23PmNo7LuO6ljv9aBAzEoCXGntq
o/d20YmhCc++f8bF95b632YLVo8tzVnutJArAcPbiJkTdinyCdH0Et2xYHA6
8GVt/bVVDo0qYaz+KlTgwkIPMwOIH32ecU2XPisu6P1EzPCiSA34ngOzNk2r
thzWW3jrd665yWoEIrRdqHqLTRr4GLy7Gwy2O66q22gVjlCQFizd42ZCwxn+
BbAdfIQKMF2OHIPykETmsmMT0jcEomuXa3i6Ibo//nQQlpxSvar5wRRpJMNL
a2wdHhbjOrf91D0lfEyC8VdvoOfte5si16WTlCEkG6AoPQvSsmFDpOtf9HIr
yiDeUJzPssnIWZPQlyxtrJvLI3lKPbdb9r0X0zw0BQeH5mHGv987sIdvRaoB
E3MHUcnh2xHmp53XXRlUz2CcgM9qoZEVUD4jMGYdl73a3OLs2JAUuZyL9+q0
XvHlGZy4CDPGYtxF1XJlTVmu5UtP3atEtoFRXfiUcR7x+B7SIpJaMV2rJ6A1
i443nAiqe36PtWWJkGvPB5Tv/O4htXcoy7c/nTkg/DGjFqaD59HcokvM69dW
/v0NRYCaTWdhmL2964EhJvUdn0Q2D6ZbvUb6bKyUEkNx6h7WjZO8FvmknCBK
Fkh3fuL88ToabhFkWFEq5HEfNNZaPx2tqZ+Lazumf5VGLTh8nDkMIMV3LvPy
HlFA+pfxuqAmecU/zzUQAWu7M3Dcbm0Nj/57UPqKWecjZ4FT9DnJ7Q9Wx4nA
Bny2d7ix7113Glx7eB+jMqLaiwbdH4vk6fIcBlQVzP6K8zo8d6717W5iLC0V
lEK+jeOsCrY/V80jARXas/HCSNZoZnD9JvqmEkSGhBLC7qkfIOO1JntB0DN4
PB+ZiZCSEgRR5d7+N7S3IBQHbxWfUnrCI1IJxaSxP68WIqHBM+sfXXk00lCB
L5/aYeYfWib2JKNB4T17cRKveqWZfTUZppxk6oc5h8KYcRg8z7pna9/y2VXH
XnloPTWz4z+8lD7miay3diyhTZHcHN5xOv2+mJDoh8HDzXfKoOkWxqosUhq9
wFiVzQsK0lhApE1Pts1r7g+J2tPNC6Nfe5HInHvZbhBil3/okXXZHqK0YfGY
GzAado6SidhXx8Lr6L9b4YPqpA04160WzUTRjvnu/j8z2E/3Vv8+AWA9M34b
an9Os7cMk+h7h77uGMP1q54mAUO4Jrv+sIXO2Ef61Q9wNjbKCkKcm9+SzQJg
g3EagYQkH4QVGtaPoyuETzbCntod85GAE9zpMnBj9lqhGkMrIZBpOqUylk5B
wnA8JqwcCJAGAcTJCYNoXa/kMQkEXLOvfHfYMMLCkKZVGAXd9eseR9iT1VlG
51bZYGZipc4g0rSWkFym49Z6PwFLgpGR/7pplOPIR6keRv/GooneMlsE/H+P
o4VE9rh+0TNqhzuYWsoXHHgbfCeKvKY62Uv+up+a9k94QPgh9cKA6czufVQS
MvH87/hF0ZQcqGzYCU+7Rq6wJ0YKjV8LV5sqXSkW3dUd0hbo9KneoJcto93j
fgSbK/3wn+MWXjHqA/bDigAIQDeyo8Q74++US2g9jQu3sM77GaQ99zXOj7zR
wYNBRuqWZ9NaD5CIjWd60ZTv8ze+wu92GGwtLKcL5VFr53WhBmQKFo4Wr6s9
/kPl4WAGJ27u9X2zuWkUgGlaq9itGJDNl2YsZL6iyfDmjpeONx4ST0qMC7LA
TeJEuf74XMiwomBpH1cK0D/6QP2bT0YZq1sHI5ziV1dXFiBML3UXUzKURKcT
nhIXkR5BQJGCdU0KTHfvooirjcD5D85KlC0gaqYaiDUbIrNnKCnco8ePt995
D8zoQjSow2IF50LZvaE4kHMFO2rzpIwagxgBWT04wtvja1M78mocPkYQtVzB
L/BKa8JPfkgu1g67GpzwGt/Tw7WJLnKQy3YErFVSt04cX+f5b+JS9M6/SG1o
iPoAyoYYEq1guqdwePnaKhog4IFT1ETiG3Eyxfkwgc4fwkXJ+paNlNyq2YcH
dxSBvBRk8VmiEAHNM/GWgfYKt8cKjKHDTsd0GDcEuahaS+VPhBLXWqeaivFH
vuhqofNeUTy9VuHvPVELckUg8c8U3MNvoA/iS1O4PDGfC8IDpMLnjDeQUsws
2JxzNdrplri1XO6EUy/lhDIKZ8MqzHCIQmiljVIR4I5gJmW9d3s9+xpf7ZN/
SdMG+0SDzyPvKcDABGWIgf+692eKZgAUoljXMcYRLp4vHvahSWTqRHVfoSsP
ZrYv+ldsv71aOQr4AerEsx2S/fMdR1NQmD1nrH/SZqDyCDDd6MVLCItJWFwh
j0JYmSyP19i2A9TC9WPJaZ1cWlFCOlbc/D+ij3M5gDzp8Yw341hx6191IDtw
soZMeFiuAyO18tua6jJseJjHKnpu9MiJnwUt8qAmDjWfqnJvTz1f62VTKNus
Ld2BOC/fwvj0r20kMQVBIFPgZ2qBaNUNlbAq9cL2U8D5bOtaQuH0nH+ACse5
n5FowVgSAxzw8WaYOW3psjAHeuea1cf7l+stHJYFSx/2w8R+k3kVpQzt+z+5
vXP5gA36cc1NxzCnKg2qm+Un89jPINO4JIAYnn4NCpz/LdXfliXJaKBH/9lL
yuVs+3CysaFLuxn+kOqIBZpSwcUrXK9McozklUAygmuVDuwxgUsUhGuH+fJp
29fMBky991OkeU49Df+K3MV4JujcT6oEHF266bRU0ZUr4Kp1y/vNcWzlRar0
HUH0TuPkdYjEj7+ToyBlB8x4Z4KP34XIiaXx6tEVGowUMHU9RQnN9w8pD6oe
pDB+ZDfU4o5bxBf4vV9CvmM05xZBLQ8zjK7hOQmsnXbzPThWy/BpVlIpwyoO
3fG31fOOXlRem23BfqQXnZHsU3/S2UcAt1q4l4hjwtz4l4XllEnIKFmOAMtY
1yK5J+Q9heUPC8S9x9dlw+VvHRO3oFQoHV2jNY3eKA+rxWA4ncZj/HPSF1b2
6lAv9dKUNCHSRuqT6Mqp9cuz0afGVIjuxNKQpf132If2cIiKJRnCGAQuyLl/
drW3hjzlXviQBb9OMMoUCxCxsKdi+AGn3fJn1WhmrCF/VljS3FKkGzsa3jgu
lzhRjsLnxyUekYxNeq4Y0zHCm9exlPgGpHK6sqH1yLgNOKqhMGMVpo+OIJh1
VqlcP4EHp+hkglDmlcET8d4QmV82uNonZTagrLQqUKPawU/qqB3RNmrFj4mj
wQVtzwJYrjGHqwTmUb1TZTFrMpfcD8WO5tsLUtbeveGCvbXTY8nhF5Yf8jFr
mdaffdD+47jTy4KtVVvMj2WGmnJNwXKBFKI0S6bWBPstny3O2rMvaTWXtXvW
JpmeRrkvPE7MofsHWI6a7nLwyQ+U1+kVRVNF4Ofb7uoYMsWtofVhR8/3wI69
1zl8MM8nGSL4PDuYQ8xkIw6lPWPq7pizbUJdsSnGwKY9l4c6p1SScXXLtzV4
m20BckqCSpH2En6IYu3fIhzFouqAtQqzdIONsi1ZJY/flGg+/hL4I25O1aEu
+c9u90bqmoCjZLU4msT2W9OzfKb0s8Y6OIjo8ggJGtyZyZ1hrLHjqWVRG1c0
sZwK/pvo2UqUfXuoLzOjxgtGolWshSKMOFqZiPy/eGQvH5XbgHenfZwYI+zF
6jzxg+Ge7baI0pH1Css7dOHOjdYRYFEynzOyyC46W4V2hSqcZ9eD9cdLtM6Q
ga9NuycnRNotZCoL3p3qlop5hJzwrg374bzt9LtFgfqWgYC1z6d/eS9w/689
+5mXSxfpZaaJNbgk5kaY8WL/iSZBMFZ3/lv4MCsjVs6dr4KEd0x/JbbF/EYD
jTxLvqRZCTrRQYR1/MhOosgxsFCAIj9CokwdXUfddKzCmeq7QY2wURZsxmTS
aWkjfN0yTaVL5epDxia+Jh0bG4NBsdRYz06SJjWpLrGNE91MmfsO81KwA7ks
ahjap/qkztKtohkGLgK+79WELvf0u4ibYJ4KJMKLBjnHmdfhzyZBonLPsz35
wHwrZaesNWPrMUjf83doZu26nH8r5fu5DbnJM/uUnOKAhYhoM+dE4CgufiuH
N3WeNFKEd10rzEdpCb4IxndaSFavyan91Y+f6c2eSKkAxrN6th/X82zKF/O1
UJk2z8vocP9vhvH5TBcPo7gEUQrNPni46kvSKYOFd40PAPOxFbOqr8X1P5na
JXARXg0sOpPBBpnuY38yuHkyKjS4vNK8/21MReFKHKxdmRhzt374h+sxuLYT
BT3gk7PUcCocKZZUdzyWEu9OwKh7Enu1AFkMrac3zVEaWaCTKtwsVblFI/sx
Kz79c3srPIDfSKN4Ov+deuja5LJw+YC3XmhKz0wcmtJMF3gHilhxV/6/hf9y
w7AqLZKGmn5DUdlFvtQ2YUQFE8yJ2iwt58sCEhhvkkd7qyUH9aTyh2wbXbnj
XhvUJFTTh0NvoTOhkhS3aNh4fOfiXxM1OWi2N5Tcg/Yrm2LwbbwdSlWOOr30
n8+ZO5061ei6QF1a3nbMsAbQTqWD/hZeSsQc1PmNQvDTcEWyqnFOsRqiBef6
LMpuzRIy+FckM36wNE/GYnk32ohzxg40/Yw2sF1ro/R9s5ylwUytTUfW3iaR
Wfv+xsTyNpjSCUSd3qAd1mM+xaF2Qs4IRJF2ZMo0fHcK0cBVCzHHUx5r6Nls
GmskXyP1fz6QJiXbQG64oODrPIpPE8A9nqQnhzv0BzRZl7M3bV4SGjbD/57c
80OrPzNOSWtt6eWcJNWPCfdqV3j5DsVR9WiG8UG2Do1DGqfjOLyixcPcA13V
SOosGKOF4wprOn48emrZAitp+TPJDd4O9fTEsQd5ZgxksqrROfrWi1Xjl1s8
gxLAMv9YSTYDBIfBzC5jaHoK11orV1upS1rMYz4/apmu60zsZ+8rYi1Bnapl
rzJwHnTpTPDnwLkjAD6QjLpfXHCjY2h4f0XdBCNma69E8dcWEkpVzGhLtVNh
7ff1slx9xT1NB0Xyh2vAdXsoUZws5zZvowcFzw7ce9z4PjBxWiruMSTcubuQ
X8v/xnODhuSNbPcqqGoRzHDaHowosKrDQA5ZB4UKrbfEfcYGXf5iS9wBE2FB
A4gygMBTgQJlGoDuWB1W0WiKxqYwmquTT3RrXLF2LIG9PeealRH7JgMEhIh9
jepJC58kcaPHxCK1BaqPN4jXccNkEb3WxDo67s4E9gOoo8tYk0MaHbTviVeo
JVeZgw1JZWir3vp3RS+t519LNRoUm5Q+51MPf+judjUHLG2NnYhvX+s/8RxC
WjoF6WCHqfI7E7eEfpdcTmtCJuslmmEO5uIUg5GbtbF7MmrcEB+CK294M/O1
nMFPb87uoNsez80BER8KwipWZfllcwlP85Dapzueab00CWyxbMI7ux+F8nHM
xr7FdV4Rn8c1b33JmaTZI5ba8mGEb49McU83F0tWQdvjbMzfF32qLyHWkNCa
3xW6sg2SNKGGmiDumQ5SRKTUoxyQnxO0gi92lP6GQFrljikW6u+mhhcsDboF
3DPDAcLh5yoI7QUEtiaGuBxKGryaXQNHhxALNY2tXAo1ntfuHTTaBnWLGq7F
ag/d1M5ddI8FMX3L9JALbLLqYi52/ekhtwMaFo7SjnRTCTNL83BrewE4my9/
DGtKEz4rK9fqlIclQQnHjOeT/vpBOcFj/Dc0il1vwy42P4W5nWXtP7y86QS+
jYdf0ZeTrIpynLJUzk5CcyItUf8B1khmSVSWg/yefMkJg6KQWWo6iRxFuSky
rIb97UIt28m7k9hWUDme5FKXPnqgSVXoYCo0whqIVnD2KSNdhKF0WFoPf75y
KjP+JjMepxQIfdjQFm30yidN4pamuQxnNAiQfaQMcK/bNpjhlKZePH+hhIsy
KfzXujXkmBW4e3WndJ1jbpPtpRCj+pD5tWyyrjoSiRYE3YHz9x8w+RWIRV4s
9nx4Qch6oMmty9pU31DGVUmkp+7vR/cBKtsUEZ/kxKmXkWSghQwzrNHu2JcF
fxna5/Qwlfa7PeTsfK5PZ+Cp7/0A9gvpSfGa/kJZxk6x+HM8aXhVSc3jRcJf
ALjgVmGWKRnMcpFzPOhU0tpDag73NViN5TSNMgkIlobb4fuexvDHZfNE9B3y
y1YhiBSOoHZ9gfk/queiJudneNu3XwGiVaN9qQCd/hvaeYjuRgHjtKDIAu5Z
D71wm32bGtpxr2KMk43LKzFDtuLMXdLyByb+z8OXfwyrYBKdFduBpxtKIIuk
3tFk+Urh25u4TpBsCB7FzrX5Psr2FGfOra3BxVOGLiFgrXYiC+mRDuCA5hiT
V5vQCpmrI46XrmN3xI9fLzJvhxDb+QraGENB3mEevaaaxq/po4AroXzSJ0SG
+1LthdkoSu6goX3DgA77ku1qCycnu5OGanRav0PQUa8dmecLoZBSyQiNgMg0
U4vivYffHIbMw6bLV4FJzXHurl68fIjwELh1oiIF7+ppre470vnkQVb6BlXQ
mLddNf8gU0zYO3WJTfaclS+4FVJvNadkgqK1QtkgSCXt1pQGoG+z2ifrQEYu
t1GujL14kMtK8p1+dDhg6IlVnzGsmP+audc96EwEvTLP+h1UHlilv4emXI29
e3HKoDIFIRDzUBC7O/A/OeYwszISeNzZ+KMh6jCyJjWB2bBCBKr8XnVLiPlo
r1CNMbwYv7QuI7+1yPOj8XCU83nU71Abw/ObxdfyxjwH76iliAIPbctIMRNS
8nOG0zxphTxVhyX/oaMn9ncuBxPo26xfHodGWnPFra5bXXfHLp9xnESisW5A
JOsoKtdBfcF54HAUBrdqvMxzMWRN85d1ZIWFvaICPU2cottn8KF5e6I+IDzG
SecE5WMEk87Zn9SZ5M9DTWACiMIcKT1FoaCGXlrqE4UWOGUR/vaJCsWXz5O+
oZTqxwYByNIvIpnZTCRJfUaQR1CAzkBS2DlnkBAirtT9JQBBkaZeHy0ZNRu1
GuzocQBWe6Ol2rmJ56/MWcmMD3tSPNoldmx7ev5cZJ3xhU0dHbYo5zMFsdfb
euhH7rmQliQWG598gmVuCk0hrBhB7HSpFH2ar+sd/xVu97qteKudd/F2RHBf
K+bGpPv8dpb+GJdbEkMvgAtpuiqD09De6egLCyzN2zTsdWeNju+zw1vmVf0q
SfIc+Gd9US0CzZ+shFQP3kJJAdeT8Q8kMH6QUXIfvE5XreXMKsYA8wewgQZv
YyDmk2nWJkNqhBkEbg8pPzHE42yBCQqfyVQsBe5w9I9KmVbEnEOHcFqdm28v
Nyih5kiWtRlR8rWLjfMZGAt7FIpl2dpCuV9DFysp2XzMuo/XVAZ4//BT+Sdt
EvEgpzAo3/vdZAhtSsfZ3Ipm+OPalwgdyNsUlK/audpm1IHcy/KKv/NK5pzc
yBgIMv+jnnR+yBgXDVToeKj+iaxn4ZO+h7OHbWxzvWAdnUz59doCRhFZz8qP
YPO8dS4ml7yxELZRLa81gY6UmTaGdKRJ9geEd9KLlO7EYHPRNc5Gi9YJeVtN
k5Fa53EoG9UGblVPHu14HBwruQnowiknR/s3V8vB34b2ZD5zAJCv9bvJTFvS
KE1jOQvX/v6lWgDP68ZWPCJDLY8gSFkkdQ/h2Z8vwVmO40tu3s/Sh2LECTxV
Lkv8mUFKofmn/5eLMrWD19LnkK7qBsXUPBCrNxChGzPKYsiZ9I/f1i2voomO
NYcjsmj+W6OvdDzUOTHB/Uoog/cxwGHjh69R6QKjrYbH9BCtSfYJwprIDYDy
WlXOJPotTog8eg7VBsKdHGKZJYpJ+nvENmFxJraAmL9O+PM3EwoJVKyWpz9m
Wslgv9aTrxldGcHmDpTUA2JyvrTOB2cV+d8CIjAtBDI0K57N4g0Cw6Md1tP5
xgBBVkJtPDAPygqoVH+rJ4RFaliqFFFKCPstdMz2IT646lmdm2C6SBPgwpGs
NgrxABdsm2f3c46WY42ZXWW9ZYae97YZCvdZ+ohE4PdIgIagDeeq9lKP+omH
95FhQVpyR26rZOSKmKkoNOsUkGYbgi7GKZGghtXc5/Z4jupswuu1E1iwUrFM
81ueRKljjsyJYtOPNR7R9nQpaCUT/4YASnMO/GiHBKJOhZBQ//VTSXEuF9C6
DPgUobQKUIpMqMFshz6fGEtbC14qWKSACoRXuZ8mM7XZKIPo4bqu8r2PP52C
KjvHHm89fxvkZc6qFFzRlGDhlcwYe6sHUP1AoVhc8gK8tX/TSuOwLyTflG0B
LynJdDUXvtO1cVoXQlVAIA5Faj0axgm6uwNMgxM2hweuU6bVeb2Lt8/FYCq+
vjGODeaepFoHobKDnHqwD8Re0w/nRplMXt+Gr3Lg85PneRNUuckg7w4isstg
+PNYNYb0Vh4X4EAIFHYQq0/9zuVza5SPLeB6x5NERg41RL5QGAd0hgvR2hFe
37VST+obzfZhmzdCW1mw3l63Xjqog3QtzHQNu0TROtBa6nTEORaizoq3WSQX
AYghLmGaQ1ye1sPPYIWxmqxzrYoSryGyVQ5XbluT1BPTC/Lql9UZasW3EtY0
s8ukMBs2Jb2GhHTr05yC0M5YMZDMtsJnQIQdV6cvUlxcbJgQgcmjjdx7AUXB
YYsbBI9sfjZopWqU/McklrPicertU/qQgqCBwp8jfkY2H5aQT05PfWCs+8LM
/LAFhjHmNgkQbtm5X3IZhHHeDRMYNnxHfQsGMq6fmBCLN5tZxF1staaPB2kZ
Nw9DqCKqlr/Pa6ZJpqHmG8IeYQg1CEL/Z8cSL4MC0IuJR36PiNdZ0dh+WenT
+F522GrQm0Um2riwwlgd22WaJkLB8eJiDyBKVMNUAKEdxCOOIxodmEkkr3nv
6syIPnX+UvC23cpoQRmsIDw6tzRNOR5m94rRkArui9C3cCQLmDxmqWZptbaW
8aiTlesYaAEjLZRIGtM43MDPoC2i1B9kg6R///EMSDBjm3MFX8OQGq1HHMgi
CL/CD7Yidt2Jl/9xt9Vf0MPg+jCMAwAouv58tITx3tfux3nK5ePoWS9TRqE2
usweCJu/Tl74B4JLY9C5dEDX90m5q+QUO1O8jFRRRHMFUByPmK9X8yXGo9/r
+oLHp+9X4IlzT+3egsuWZ9bCr45YQqeJW72fM+K8O7pZSvGdmaCUMjw/TtSX
nz3NnA6gZjWGET78G7Okur1ry1URiVbI/BaBitfNYUo+Kwowu4YRt3eO0/Ak
2x1p0jpuqV1/ZgF62yfP/hcl3npK18WYFevzqf2rjxR2uxR0qI3yc3cXs4jb
IwHBMpC+/+pqo9twPu/x8INPgAeO7o+Nh9SK6esra66QSeTtulYSvOtIq2rr
KeyxEXNvScq63e2eCthqqNqY8JdRV2KZF4rva0vH/KkeXcgOOP8bFK68Pp4q
UMBnRo3Nud1afYVyba4DAfaWYRUknoV+S1/fvIT5MQfb5PEsgwOKGUaaqVPw
8dbdOPx3OEVASSrmmFeCwbKj1wzL+EYUw8Jenys7bjeZXHujX/0ZLpi76a0T
0IksyDO4deUhTrbwLLT9lYjRvKMTqQWhhcYA4aA/CVYg9/qerdU3skE6jUMg
if63AfW+TAbT8AWSiWqOECWe++SUogC44BJAbzfTfVaGs5TNDyrKS+bgBvGG
LLVvI/iwmsbFpGRgYmQ9dF9/V+jkGoxQE894vsoNTlchffE0DGscyeC5rwXP
936rlgNpmLj3Ekjm94+ckFe4WGHGapw1OfPm21hnGLw3GeJWiEBsPfnnO2KL
XlaKTGfNVs+JZ0sx+h+cMUdOiozf71qiEMiBB5CGFSsNqXpURTT+3z3wQeP5
zDhY4X/+ZQEEDE1qVKZZW9d9vj03eGMSQqkhH+0x9PgemRaw68mmPbrOB5b5
29GR/WkOiIQljHhMsBKpieDJkYliKzD5ta1j0DRbG0OQPzoeSgypQzCQ9A73
JEemzqZjTt1zh4Xz9yOn/ZSRHAj8BOAV0qvqtGUTfzzDNZQaJ0X+UOCKnZla
Kgfu85QAhNox6L6fv5UJzi5g0DQtuvlAk29zjXde9/zLv6LD9+uVyuyGkCfi
Xes/XVrTgd73B483kZb8+B/ByROLwals0EeVBcy6I26x6As9D+mZNNN3SHEm
IeNd0zxfZH+uqBuEdl0DJ6T/UFCaaiaTjsh0olUsaoMeNBZngbywPcmFRGUK
KShHTHGR5x4xnq90DnXIiv1/6fYxVrsh9sD2dZF5f7Wff5Ev6Nq1FpjFxNgI
nQzXBoVyitLqH+IUpnUJOksWT0aTVBAFmNRcVJZ9Ni2L7b6LZMBnnds+IpGk
sM0f3qkXEq7vlIUOEcbkjY0RS4CRrg8nl7jKBL9pVafpjFNQkEOx1BMqa+X3
37tD2eNh/xaN1HgMY5S92u9d4+fQIwvPwKjcPF+lQa4hdAZK0ywLW12rVIZB
Xeoy6tuefHUGtHPigkMqOvrQbC5d4my0qZHXguyrRJzVRB5bUpKG8uolfn+n
IrBKaIxG78tIqQQISm55hSuTqtvZfIb2fX6N3roEBmiRr/jo0wLjdszbKvGc
BXy16tQeWvtFohRNNEvFjMywgrwUORdGRB71IbSzzgzwL3UbDghpNDBOT2zw
Y6N87JXk6ZgEwnx8pijvzA7E3ztJ76TyBwvKED75Y0Y7EKfyqd11OpM4KuDy
54bF1SagjkE0uFQ9akCbd5R5lUh9ptady9SInBD5dhOiZFqUJmvYm4Gopsu5
F7TqeIrx3urzZqgLV/nOdEqfKR/vkYTDLR9o7TROiR/QWQPNwU7dYgIymw/i
ZOubmlA2/BC5Ik2NmN1GyjKF/z8Rx4BUexK+kDFR5mQW7t52z9VC0FDnhMhl
GM/oQyVWVsEpl/EHIVvnZYEqW986z15Gsaczx0ltQP53F+hK2Gat/b1nwuAs
cMBuxo/EdQi8Ktq3HHqubRq7AYqq6eQTp3p5Vgh0qHCdFRhh2of7sKrp2NbB
INoqh9VDP6oGth1F6uJV9bmGDkt1/cfqvrjEYX+aCPaXNGi8j7UdxEyGCDoT
njD95hoRi1cBBVPGV54tEzCVTO9QzFN/HA1lsXd5cBA3evPbQBFU3M07uAFw
SjPd2Ig6aLaLc6x+8uLrTv6m4ZoOjiP5OX1Sc39sb4/x8bYzRuMy2XQ6qLEc
rKukDv2+12mYFYegRVipLHFjhCA0IdMAZHz1WYkudMrPuqOdGEAxNqhNHV6x
loQ/sI8gFVrr2QvQre2q78Pkf2zhytYK4EjzWLH6CBxJKOz+CwmtVZxEHpC8
YlEbD6Vj8kYYTwVAUnKhmbKsSf1nwajLcwfr1F4iAlhY8h1xWcFQfOpX3gnq
bUB0cNGMcUaoBlk0Zj4aSHSpwZ5PMfR+t6Y2CDfPOc1mLJK/i7Ls4YKCHeP6
a8SpvA+/siNGPXVGDsesRdsYg1EvPHf4VUhVywXBiqxqiPBdExeXQMu0a4IY
D/vncBVAoXkN2VSPbj/nJ4MFvVDYLZ9KJhhYsEGIwQvZx2YhhFGrjsRjxw01
hv20dtN0ETD5Fy5HQSXUBIsVbLCXnIB3AFt9xrFdY4NaNv/SpQ01V8btW+mm
thY2bW7CNeBQHiJlAf2fCvRft93d6qcTxQFxFIHCEZVNbFIOGORc2Nmveehf
i74ZbZsjUfCsxopFKIOngwVXGhDX95BTmumaSKbuUi9Xf8M9rF26REo1GWFv
Oei+ClGdaWF0J3DlLn8NAmorUaxEMwRhc5EJxoPFByDdZ0v52tpPLVtMJwyl
jyr2IxBvC7AXUKzakDF2POA+0HujApdZC7cacib1vzt41lhtmVgRR0jV+mhO
ITYFnmVw5Az52nlFE/VgDUCfJ6h+NihSMhDJJ0hr4mqVy8V43viVpzlLLkAW
lQ8qf+xMFnu263AlmGIwnGrycX3MJ6BGv+fpNINvq/hsn9zlAvGiIFmxV3EW
ljd8w3Lfu985LjM1GTWZaivZA37qbomzOAG7Him6Fdw6suCKbxh+zLfDCYCA
UQt1zsauzSrhc/vga+NKssY2rn1NMS4ZNbjm57LBNrZ/LrW2PRUW2QGXIrEX
avXEXGxSbKjf3LShbZ18RpHwBHI2YO3qp0AfejSiKHtPV3erZh2oN0irtVY0
TLNsB2bAnEdv3MnpzxLZQI0XyH+LwsX7Aku51Xi0jL8jSCOC7rg5ggTbPXOv
ImuUAliFSn+GtRNEdXlKpi1cxY/wT19uEaPEpZ7bhIxgrl2pjzHJnWBLk36l
D4rKJrUzSgKWUaDL44RmpgunoeoQRlsSTbWuWArI4jKK/63hJoZFcigc8pe0
cl+od1iZYER7ZG79f7Qlxu5blNUtwPrcy6d7w4drQbwvz6RQWsKXEW909FKe
6N4O3IDMonT3Mfx5Bnb7oPIVF/q4hcDj9LI72754pKpIh/lJh6y07094d3Js
RVdr2aPfs/J5Ort1blT/IXHHhGzL/l7y5BUFcitehec+g1Q6JVQR8R3ExBop
nhoRlwqJbwL+fXnBU/RbkgTw91ui0ufdhFn1krzrrriw3Q3dU1s4KjqAfqtQ
glT8E6DtBJYdRaqHLT2RbaYbFId1oTjwUNmaO9SLnkqh0I+SXQzUHSf2ce61
MskLSeTH0Ck/CWaqs9oiFtBKh5g1N1tbBkV6Lq5g1mIxyMIi7I5HYYvRk2B+
Zl5yXZ3LdxqUsN0cnHfvdpiszJg9Zaxi37ccIB5yxXFwqlY8GkriRr6XKi7e
7os9xFLvlrF0BN9bA6a9A/TwX9vcqfcyFlbvqGE/eaGBZLuPh9DNvQ+tm1we
bJ6/esPL8nORzB4F4HnLwdERZFxVTLEoezKF3RQd1/mv8ERldWQtKHwaK8OC
MaFtIV8rilgltgvXNyh1C5ig6me41w2h7kCZFurtdLYqRRuqLgR5BlDbKEj4
CR82gdbjQ6kEK4P+EYSXI3LGC4gUl7EXVyB9FhR65+ozdyXXXUZtGSLS3lc0
ZaeptWVuJxegoElhW+wnPa6Pv3Bv26iL50Sr6/wf9gu6Syv36tHCwq0CfkP6
KWUTuTPRMQFHPrBHkt8APwA9L92WDXkg/ev62jdbSDYIT2WwBYkOAD0Iz2uP
iObVwi6dKs3M9OyCRzVD7vCsvPlRHOuk3/UbJY+/v/a2YLdHLnjFEaZnCGR7
QxBXzQAiYMUzyDeYY5Ygp7AJXu5b0OakP0oSo+FlxXcyPYnH/IpnccPCL9Wn
nNzq9ho4stAcznyWyrhr4Z6tIs4mjKdnjPG2a5+aLZd1fj/J+OlfraIvZpeh
7/tM202/hJ8x5DTsWY/rLuV8s37wTN2naogJU5gWqGDvwEP0KIK7CRog2SNJ
APYWKKB855kLxtXbetnGdfqbWne3/qY31XlCkXqRp2aFmmywyr5uHYO2+/Vp
ykYQ+/FTZq8qQfFoOBqTFSX/24mnucUiqj8mbhlWuiver0TJuh+svGJXZJHM
DZjXUwPhs5zRYkHxPIE6/Fg777777gkRtcQ6VBBTB5W2fA3hC/9cw2oE/8PF
AnGtSm5L3+5Gm0c048iz0SZMjEYl+o7/hLh0dMiWGjMi+XzHa19pIll9WG6i
+l54jBKJpi3ObGyAj/Lsf7Ldos3u/vc0FTR1N2Q+tqRmHIgfvvukJYdelmlJ
hNEP9Nelo5eyYUz8Vc/Ae/kDX72q28ZXxDE++QSrVTwMcddKN07Vik2gv6Yo
q15V2BQ+oVU+5CSywGqYbyXbS6kbKGGHRgLviF99Ubh3D1qCLOXZCKnEHnjP
PX7pxP/fA55/x7kHNYC/263AQg2oxtkuEOGhr/rp7iPtIpX3jJM6NnRb9O0I
nLH7IPiKCIcvzHswAuBHofRRbn0mu/+cATP2AGoPLyN5sJ7CYgMheRmK14KT
xx9Bw4ixGmUkwXReeBp0UNVcFjVQLoR5GbALa3lxKwixqUHXj6EG/UcX9XRO
ZkSnCXACrJXh6tfSshRJzM7lp87pjEvEhEIHC86d9YKnGZ2MFyYTnKVcqfal
OzO6k6pLqKbfnEq1Dx320jc9lJXc2wEgvrzS7kstQ4WbXXv1AsySmxPoh4Zu
74UWVblfl/T4eZoCmiNraabJ7cT+sPTGCKuftMOhjZP/NtG//veU2q0WMmCO
2E4Gm+44ZSZKD/cjPygPf4T7Sk4bTQs8dzfK3RC/cAtI7Mtulx4gcVQMLQdA
9HJZc4SDTzs3wPUct9YY3dfU/RRczUSGwPcYOhuvyy///DWlnp3+hEpGa3Gk
z3QWqUaow7JOl/38+rk7Q9lmLvsYWuBAF3M4Xkts3313qNCjpFnTwAOfg+wg
+VV+GLHB7wdgvEnvzJYZRG0fKarFbWj4N8VgDGtBq/k0xPE6U68IIon4hg2i
iLTsYQeW9EoM2m2T1Evhyn9UgilIkxROzalr6CZKTwwIgHPBkR+xyG+mEAfp
I6Xt0qiJpM7982s96FE3XIX3Q/s9+ONF84CUmO9T4YeW+dds7mN+8HjofrVJ
T+ATyT0JD2jKTibn5tbC3AYCDoKwuWSqUbERdLpP1hEbUl+wknE+1WutwQjU
azdA5HVyAuu2x+jVHTstWthg8dcHlOJ8MXdg2q9JY45/PNbWhEUqNwjYpd7B
HpJd5Xjsnz5/6rzVBngHcFFhoOD/IxWNmORKV5zrzBUMO7WHPUktx874Cjov
2EEZnq7Ylci80qMYwbAZCb3GUmIQywHHpFRHXmY8zkh4BBGjwcKnLOHmg1Q8
Wf/XbdJhmsUr90pHO8mSb2Yq+N4wmZmveFVeXmmgWYmCI8Ppv3Nlq7cToBiI
BwNupHq02thjgc2UZJSnfp+sZGR/JDT3zmlYiBvFzj1D2tIwJYTYpBVDOEyx
rBEH3SFmH4HBcfEb6MQ+w6fCRBuNpTX+ueb3g2j3ogzJaP6zekWs531h/URn
loiZud6nSI2bRhDTflVbSxuh9y1VHa16ldqel3DMeirRKn+uu5ewF11tF3Qb
MOeLTJzTedB7+xjTz0zK5HspNF13gy9koeh3PVnpah70yw0ZjyYsKIAX9dle
mjU72bbLCLOFeP5mhFEJ0EAK7bTK+mPB7s92DX7YPxLZj9qKgsWCK5l7ZScb
LQtuTj+7t1wKVKjwW5OWbQwQ0z6EWF63Iuz3PeE9/FM0RUOh0JyeTy6ztJ8K
t9yxdXaB5QzOQEZxmUVkKVkjBcqQGu/E9txW8QbC+5ZCp2xfS9fak63e9tUm
iwRlqxccrlDk2m0v81qNNAby9dkVOE859a6X2OcPqX9+UzQmw/KgGW9zPAn+
nCyPIXXaosoCPjoX+xy0etwXRcXXfTv6H9MmTChLiPeJNktKvwN3lHaoQSd1
M9Z7q0qce8Fw8CxQfkZA2Snw4M3EwUCA+IWXlbQiIwtNRdcMufLcBo/cHhkQ
2ZtMBcLdgeWDQM3wP4h4MaL9jy6JN9rHap6A6WWPr8Zk3HpHA/6SkGzXDfzT
0eUq6KdTNqS6G524o3P6vEYB3acb5grqZ9WAm9BExLUlyz7PM67a4lAw6ufZ
W/NFZT0b76Ig/LZTxTKNpC3Uhu+uHyy6LsAXwPd27vTiusAMtjV1fbQ/pY6p
+FN9T07qZ0At3enA94Q1oHA+rwVf+POuSiddF5DGsYchRm/J+JlUBqLMbjqZ
we0u461I8YCCwpikvD4CToL7T1hDywBrKRfY9mV2cTGCnnpxYCuF0yLDXuZy
sfXS2VHAmSqYTLXG0tvk2RfyEoromZ22sdSFhpcQolHGonwYNDQGyDKW5uoj
J9XT8bBtQyghhc9xGpaimqNAenvl931RghCpyatDT2+LSYNLL8L7sRdBPcCQ
dnRKMYuI4lBE3MapQQ2joB4P2hsbwsCPm2FMKf1/X+DSPM9x8dbYaVM9BKYW
lYfRcBWBLMhz1K3Ywo7i5/VYAnuusEcVRlpCp0IoII6RYTSYEOBdGJXag/i6
JDCvbe270tUvlzsrARyz4+dmc0p8CMv4XF8FazUh3VYWDNMa2/exoyO/+H2P
uI7HQy5wlTZOuBttb3CUAKqL4bhSuJcDLBGThc1h099+f3/gWT2KWkK3wtnj
0H9AELNNSMHqcl6b12s76FrVihvDsh6DUY0nEEjzKDnjIClFkrBL9gLuWzGH
lcvMT4ZmOMzTqIJUil0PHQQ0k0P8HGqeAFMC+CRjZ0CKPHewq//15hw79tkU
x9y1RlblaPDP2zIYzNSlLiji/oIzhD3suCy7Nw8EONO4mKLmGAKeISe2Pddw
FM0LNpCi3TMo75Z1OdNHr7Yo9/VzKb0TZ0FP//hbQWHZwjDvpPe/kifiYQ8r
f03LT8mlBTSypM5r+K419wzkSWAY3134B8UsTra3uiFs/+EL7mVi6eKp3dfk
SUUpUiL/RxEy2gO3FGWWwn/tWsNf6Hqvb9sgzcajD38BzgUV0jHGnjOWCp3W
YoZmzZqS9QdrI6etgezP28rjjyA9UrS/H5yvd8ZdvG73QgX3sJ3lAIthz8rz
WglE1x2mfLGnb1Jyw4W5Ozsb4pAQwuCB05xvYCM2USgs2eanmHf0y0H7K+1L
n7cPZ/RX8fE2u7pAFVuLw0G6+Mn3ZCseahDDp7NMKSPWxa766TE23s1vNlNE
DbxihaKDv+nM4EEIaKZ69wxwe7DS2ccjSkpkGH3pmZ21XqQR3wtaLXudHJXV
jvkX6XTufeEM1dULTWxcmoml6PgzKqhty/pIOe1gtQJrU+yRHcHQwjcrjE5L
/sSrPXlKlJTVu4jgaAH1X9XHb5EI1YgQxq5NDPU4QV0Y94jvqeTMX/JVaprV
eG0yuCBQIMgcX9qmkhjtKr9wZFXEOGpy2UcWsSbcVBd6Twnx1nd6QMtTWja0
+tsjWZNC8vmuZhRfO3Ceg2/FI04agiZy8BAE0KAdIwYJQtSgtRHupGBd33NR
BzPyeczSPF/DzQ0W5kzBVBesFx8fnaUkcxwwyrmXTnzj31TI/0MK27uataKQ
dx54YycvWjdhs53e0up8WVNu1L+UWLMLoJJnxCnoNUZrrKaolpHkXrNjZ3jp
KnVyd0K0AbvZ1lw84BaB6bfhfnrrwB5tKoMIrIiNXWhPV2gK27PjFYZjj+b/
AHbml9UP292uKiaAtpYxW0UQLw+Ht9w+1GUvAJSP1L3Zp+ijfDVaHZq7A5zb
z2CbAZqEopYmwUUPFm409KkAmQnZa9kz8jQBMtLpo6KGc8lel2Zei+tlHgjS
Cvb97C0NhQ9e6rcBW425AZi6QCdtphTzOQYlxNqbaO/+yQU7SBUCaeHOomEX
stttlpfPdmEUAQDjzRWz+BkVbxkFpLYxkB7DK4vgPbHqjU9x/ljOfjNNyGvt
QgdbyFOuo8cbdsJadg2dRbA6cBiaBrLvwaBTTstRe7fkNJH6kMMJKMiHF7A/
7/Z+q5xOtMksa7szZDbIvnQs0yXTz7CJavwFKGzmvNUOJNsMjWKndGTjPudz
6dbG/vO1ty63Bj9c7COsQTsiOAv+4kZeD+EMOKZIA87ad31YR0C+PnQuNy8q
2hHclaFXMg/BSg/CHTbpz3SdxmWzN3tQ7nCeW01Ri+0Gh1Sc/XBOVjEN6gkW
ZCQcploSLcKk0zfyYrNNTD/Fzl+pvc9/X+zXwpSPBfmWzK2Awajbcrot/yPe
nmazzBGrkhLmlAIMbDjIWawJFFW9JXltHQrzZ1w9rSFiNVA00vSIvmQ65sfn
GfQZjXNmwXzcmqx7TfVK/gG5Q7/T+iMbUG5+gO7lHpPfMmEg0HjtNzTmUK3i
mRpDHjEYrVDUaerydpKmNwEGkked3Kl5mYYqQ1Q2JAdlw+CV7nnPF/Q38yO7
irJ1HnFqMgk3DnV3VK7k9naTwNcGJyig4hxZqKwGUbZb1esd/F61nUzUtqsi
kT3VJ+frWyPXDKZUg5jQQwheGhanyABo+jW3NzIC76CvysYARO3Hou3AViGC
HDQRfaqYK6qBTijF5s7/2um2oAnmDGU29lm8U2JRf8VgiSSi1RcP1NnvJ8Pd
sjAodP6++M3v7YchcexLPftYx/L8rtPYC9JWK5yiRz5tHujwz+PFT3v2QAQa
ujQTACqlV8ZePRaR72pdETQvYpfXrIAmhQdfTbnXO67ZcP/9HyGeCY4hlcN4
yCxDgDU5xo9CiGP5F2wwwDDcv3ah0T0IToGq6xmlVU4PtA8LJxYsjMnTwC4k
mLrSJmyR3Gfk9hB7Obm9Ax0hSjYGXmpgJnMT0KCFYiORLfQvQ/Jxgy6pImmH
V51xCCcaLRiaXDYJPON1t3SJ69vMmWpjtIlp3GVlk8It8ofda3ZlFAXaFaNP
mCYvUCgprdXWDHWkVx78dmGWWeRJE+h/IYrA38v/451CgZmWVOj3pY/wIVJu
phVu5gIurROnZt6Is6IIgbWa1BIZK3azp8YNGLHQ3+RLt0xp/lfJAwYPqD7d
vejKkHvv5lIivJsnR6dBpTTNiCXtEkXiIAGWKTvSdkJONaiM09D+qla2lvXi
I6NUD6e6N5XutzrLI9tAVZyhY2tvyLievZj0pREqn3sODRFe/4jmuhGpYMv8
IhJZwv2GZJx1BF9JoFhuNm2EBb8L7xcAVpsvFri85bjVUzSvdwEZ6izIwWEA
4hCcY8zkspo7sVtb4tzKP6VM78U9kOtSr8XLv36eZL1VmXsegMmjeIOsGDJr
ax66MdAUJFaON4gsdQ3WU9tbQ+iQon1ku5iwnsHTHmE8AavgZQu91l33a7Lt
K69qkzPVOrv3YRmViau8dV0V8LWqUdfSMM8Ipzbx+2Dr2KqosHBOOQLf6p/M
HgOYQuHs20Ua8gB9hBzNkU2vuMn4JsX684slmhiAXNltyLr2jagauEJlzUHv
94QyuW1FR70o6JOEkcdcaTFrAVQWOiAHWYNqutViFneewNhZ/EKd0FWcOLaU
vjmYIO02M52+AYYUQNEB/BeDdwGi0jSXq56OEIXPcPsWVL3lGB2fmbAg2ZIp
e3uJeGKhjfF/8tcyGZBkXTsyscIdQuXM6srjSYX1eEoQDu/ZFn17mj0adqsx
sWjul61/VmSz0l4k0vp6efGPF/tgBaagzC8ZAHPDulx34TQd9/bheWUB0T2J
9Q0R7dsRRgzs3kDOcVkd9yiq4Pf9EChZf3+B92Yx5mdHk7fglB0+KnipcLDN
WG3vzNGBrQ6pACUgxgFmIZHvmyhKy2JWHTxZBJecZFpYMuRmIAnhzUSBNLAr
ZuZUelHOO/PaTGuDJyoi1cm6/PE1xKxt6DjnvskxOdO2Dmy5Zttcy/lHCwGr
PVW82REDE4Y+hgUIM6qtJlrs6PzrTR4Dp4vs9JEH2Fpy/wuvTN+l71HdRGDa
LNme0QoZwbDUQ23CJs/usxHSkBelsrFCbUeipvGr8NCBBfSZL1NWizpeuQGY
Xm2Pj3Xc220kggSGtXuUtWXFOSEywmuTg82v6gHoXUsynzR6ldK9nEvqwhtt
oIpmc6CZtKn29R7SMXqZr+rM0U3zTM5WzSiKM46CkWxjc2Ra5qhswRJqfLln
7GTWhfNGmZWVTg6hIYQiMjQFL56Zv/mo5V6ObK9G4ps1bgImguZ72JPJ9Chy
rGywDyDi8Z3XdHoHo/ITQ0YRHZ/XefSR8WsZBMTe7HO5nJXk8Tgl9T4x2fAT
zSbpLLSkCQKw6nK8o34LgbgW5meUsE6+go5MsReKZhvaIqvKvBX2HdfXcw2k
hLLGJg9JAejREi7pwiR/htNH5B+k9sdL8iOuS2PhshNkmNwmEOf7JgsYh6o/
hBkA3ANA8MnTD/6dIV67Zpk/67CWWvJ1FQHpN8a+4HGnEDikgI+yJz4N+5Z8
X3OAfZTL9MuSLYEV8MnrrTUnYZgf2T1yzW9J/a1s+fCj61RPJRrEyrInxjfW
xxGQHaUhFBPaLhUbaXVOwjD2Gw00IRjr0aoSqI+0Pyxb8W10RRdXOIgclyiP
VoXN62dWMnMdHx7Dr3YyRW+/5IflGlqKCYWnOscUlw2nPPJ0qCImvwRaD1s2
O7Tl29I29L/aabHc0TXpOiemevsf3oWmL5613pCwVxLdgBa/93ObbZmRsFw4
M7sHJCAt2CC8FnWJ36ElnyLJBsCfv/RsBi3065UQGx0r+yn7K4PTmS13blKj
3ddYbiosIceY5S12h3khawOJfy1PsJaN75+yZjCjYQQ0p7P67kttPpkbuWWB
MD6FQz62E4PxR32GxMRl1yE72SOXVs1UEDfge/1oICt/fjieSgggrHdUavHJ
YoOHbgM9rRLqNYhxJzukTcwDboCwaChydeXLJjT2d9cF4NxRPNNjX3zv+fMz
NdoftXABxX+tl6vfaLAICk5LsisPhxHlLROFbhiPXrGMT53Ek/QlSM0G2az1
sf66y4rXjYmsV7CHbnfDJv5wdT7V2U3QYprTRLToivUoCJB1E2D9jeX3am7x
e3yx1hiDvHdB0PVq2f5HqCWq7rAcjEKeeBnuFDiuX96ne8UsXGS45h+pj6io
AjXCfgeSnGowO/cCw6vpt5WsEKUY6wTHAhptF5FC7MRWyB0l9cjKLtDVn+DM
gu8yqVlEpvGzQnRVDkB1Rf8yKvjFhxcoZPjIQsMEKeo0JSR4nIguR+hUej/f
Ep40q4/vas95Q+7CmMhFl5DoDhjaDDjnzuHgnqo6JueKJOUFNRZPJ1jwkMU6
kA972m+5ltyiCth98pgnYkmWHzdLcSkpcGW861UXGyVgavksydQb7BXzWrQt
XvqrQHKTBjS6iCDwAZOTI/8FTQEzdzCtEEJ5NgeLWpzTeP7rFvY/uOLDSlY7
/rQtLy0VUCSjjpB1JxoD3p+fZa4P2A37/VvkN6lOHk9Ym+y3mreyra1qKc5J
DRLWQTX8Pbfy9oL1BPWJjeE0gv/H533WSZ9FgeM4yruHOST9SCiFd6Prt6/0
cJFvRDciGhrLo4r9wRc/6na49uZVW9BUgkL8ZztqWl6EnGf5WQ9iYfdvyay4
dLKsw1vT+L8jxAi/vY721rEWKdCjUj8cB1BIFlbwvyNGj0jfqPhtSYawAxcg
h5DDUsXsxfpaesyaJaas4aFEAh502CdrbOdpWLOsfbp+UIEQkAHsx6TNzGDG
3K127IbQc8YukNaWTugSa59vjcj2d6DNG8PqOvRwU6a52sBAMH8upePsF3FL
5B7jVuTlgxh6s2q7A+8V9Tp2hfsxP5NtHSZGN3eNlHLRypp4TF0t+OAa0u9O
aA9m14f0TPrj8uScZvL+RDP9/ELL1zkV2auSPki4s/J8hnhAKFtqPh0RBIcU
47CBDg2KJOLjiJcz8WITkWbSwMXjo9SK55egXmFOR9effmXHuL2LFXYWLLlw
Vt4CwfKlLVoGTmMIovNhOYLZS8jLcljbxfagBG8C0l+xi4GIcMQ0yoOk+KqA
zmtJiVLnHcO3poOevLq3g5SyF3W0ODk6pI+hhUVJQ/M2Xs8wrrAoJtNOhQLm
WGq+4p/CvhjrRshWEiw6HvGjD5HOBw/Ek33RSb2qBTgc4LEFHEibKyGhbYO9
uL++INSs5uMZoFgTqEzTB2Y5sJlgdy0RJ/gO1wkpaBu9rMbdm/YW8uNi4Rhp
B53CtJkKK7EBaXikrozG58w7vnrt3fMJp00cQtEqfWmo9/ulWRW21LyROkMO
d4VAsQf0RugfIKb+mrQsxpogd1pGa74aS4gJgUeIEqERPG+Ve/4amuXFjwRB
F7t1DVQSqTELxFs0SkUQDs9rmJIss15jsF3qzcYafJKg7YrTJh20wabqxqIY
ZI3wCdy5HVO3NCcPK1pvRZGhRx4j3IsWjIAOSaFRmzqaBAyelwREkpj/tEoQ
GdgbvEkF8twnkmxIiow+/SzrZyRhdIjjDwZEVq/b15MxmUQr93uSc2UyIitH
kpjLUR+Fzmu49dlRK8RC3r7K9sXNqricB1ZwTLHgcUpBlTU1CLzA0+5u/lqz
ap4yGJMt7hXVAA4dud0BNaGFaJFKLw/CSMLMlLSclg7bZCMNNbWE9OIGYRzl
0KRuEeqSnqDNp22cV434D3C1LGE35o6jdAJAm3QskslSOV7d9GgZZmTJlxG4
6B2EVKp3gz4vGvIWReO8BHdQQrLX71Ux7yprBHqlsbPgNluu/OnsHBLy1Tdq
tOa8YhWW/tEOs8s47F5k4yLN8hklfZfJQhR+65/4g86twC1ML3WIIwzCHzek
HbNO4IqBViTJmLI2fbrvLWqn25Bky91VhtyKSCMMLzv5bBu1y8Z+L7bIn8Ep
rdUSzjvSKnbs590bAjSP5v7iNteGHdVELL3g6peDEhhy9p8+3icKQvSQaqxI
+qvEsI5tngzX+SwjfWBD3sSEeJjczysiRtLioIeC8FrXcv/KAQTA60A5s7cx
0QsT64JvOaTgTU9UtZY2Z+rgR7k6ASIuDj8+qCvH9LmEEcJTZmStcvqOwDYy
1gGp2OBYvYlbXgcQYFyKjdzlSNK/b/UoGJkpbeiGsYXDj89Y69q5am7NgpGb
Txkhdi+xd/opSg8osjxv9JV5F1L0Jl2K2X/3Bxsb3Oel/d2yhge+J+e7Kbet
2L0dOcV8NAB0MhsFH8obriI/2SObpQq4okQQRTcf2T4NtDwDVxWi6uJZBwO0
vMlah4rOM30VFPmtJ1gthUqPlkNG/jUEDSl+1C4/qOvEeJwEZ0KCHEO5EwXG
uHZtPaniovRmSgPyXPBBvlihXhabItRB7mh4nmF+PcbIj+LBhE1EECNOowtM
Hmn7ct7xdSjm4rX3bZlRHbqf8Ziq4vJgMRkjG8+GP/IvFer1/cchcNii1TLd
jWU0dhWeenHs+FHGxfiezhB17nkDW5KzjC5TWBgAv4zhhot8WF38Ciwkygdi
LwTNcBJyGBvRoAeD/HXSyc4dL5AUOQw4v1ca+CWPZ3ivy1WRmzGTD2DZTJmU
o0orL+X15qpYOorNlkRVWf0cvyt8tj//xMSqsHCO4DJ/DM2yav7E+siODHQB
ySDhaXEl++2m+4u7dyZZCFIHp5sCGvdVp7qUhbNm9qdLOAvB3TqsPSRaafTn
T3D/j2Yt++l51W0IPRPkeO58bKwF73cehFc3MkNHfzKTR5LcbIFbEec3ACEl
C6s7WqYpxAKpL5Q3EVYWSVguHFYfrKGo7XolTTGVO7wAoAx74ulARwoQH+gP
UVjfRqzoy/ULDFJC0XcTCvGtf/VncIaNF3Yy/jJgQusbfZbNTKllMLaTO++e
C+xCvyGduusBGPPNtf7mZyF10JEYeKST5gnlhWISMkKw5ndnqmkFVxG+SmPn
1V+oMdRvK08R/VZ5Aay9rasBodU0eOYGLTGrOrsOOks2x7owE3dqPAkGl+0K
AEIJrGrC6xf+88FPN/UDZiR0X0KMD9atSz32qJVAeVK1nM8NJgV/75IvYzSC
sFtiVducZ0VnxCtCAiAQpJ/c2klWBKgEzQmJsHJ8etRJnSp7LYrxVnTWlY1V
+Qd0LNYYEZ6iMFHPpis9gXbk98dWoo8GYihjIDPgjkJEwLZvcgfqHsIkWMet
v1SiN0KHVGl/Z3iGxVhPqUK2D4jgl0tj2WcQ0p5Avr1JkPu6ThL7BR2RdJv4
ozlsjMQPgA7jIBTXhgDdJ1vW8xP6k5TlutDgDsNF2KJvcOlNIlNIs4F7SAip
xWaGRJ65XfUU4aImsBZyK/4I7EpQrlyW8pGJ1/x68Z0GEpEwyrK8iaPfN8E3
US5VU211gTMkU2miFtR6AkGa1SrLAdEy4GCgy46m7N2DnSCsyaTp1Be55IHP
bO/0KiZC9ONqLuGEwcjtEwhR0rq51gzPo2Aqr6cltpNViEtLC5fa4UyfnLn3
rqtAy6Q8JFv0wvcDs/7lQr0X34CswypAJzHG75E6fuU+RGbHj3SZ+6QVuuRS
MafYwv3dzuPAZInmAt0qwQWIDeRONVTnNPmFee3n7blJujXnGcD3UTeTv340
Z9DQvXfOdauXL3pQZsgzJATftsIL16yrCSAUATCY5YRHk6CQOO5Lng+S3Xdp
dUyQxVpPqa2B5dYTW7o3bIoS+Giq1NWDOBkDpdv9sq6z/LW9jdKhYXnYca3F
K608t2eOZ+m2e7hcX+SK3hl+UY4kGXmNVA3IfWNMLbGV7RvEk67zsVvEf9Mo
O/lkAndIldF6IkSScCuQsPdDQSBE+sx4nVNbE08L9b1DDorJi2R0huZW/Rdl
75A5ANt6j0Wp38HazdT5ZfhUDmQVKEyMTYYFQMYPPgq30ND0JyXQ8kIP1g5o
PrKIP0SfQvUl5zW2gn9z0ZjkretrY219dU2pgPJ9igvMFlW9+0vyDEj3QDJN
cSTkajQ8nqy342uhaCVjQ/K1+/8CIC6Im4m/LiVtzf4G64aI73j+NmAR+0Xh
q8A4GuOCvmhVQga8mB5hTCccHaVte8KBO8sUZv1BCUeEjzrGCqmu0cAk7z4M
w3+miqEqeeqKuM6N8A0Y+4xpeOQmUNlY/prdywEktuPS9c+5xf3TFFeHMT3t
6iGO0cWTvoYH20nO+Cl392Y5WiWitIkh0aaMMJ4tbNaUaXAcgeqFz4tdKZ/R
V97xbhO3iSl/R+YVF1zHzlwdp+JtSfs9VQcX9Jtq2LmIM2hbmdQRd//64t3I
jYpbPlHr4CMbigX8lt3MYBG9u4Ped0E31H/4BNVMaWqKPqQv2vF3+oaL3hoD
OpKW7gIL4CgecS7ZM0BMYmrcxXp0QR73A+J5ALzN7KvHCNd6p4PMzztfcTo5
E8gnMz8YFsGOlTuceJ9I46NtMRiFWMXFEqX5KNso2DaZ+ZLr6pjM6R8SxfzI
HoDtdDfohg5Ji9VpcBwLxV/XaIViHZyHB1Lh1VTDbJAwaq/YpkTe8gU7yKjy
3N1DUc5viQsQiiqVspuKVbOIRTyZgiMFzcYQnqUgD63F8dfy/qjer/qOwPmJ
lrvtGY1Up7b1lImNkX9QAeW1s1XUnQ1qzXwaTVKOcCak/dDPKQfTZxb2Jm/z
anSp+FcA9LpTOKM7OmE/e/1+J54H3RGj+A4tZr2qXHKAPTkQnsuoEn9x430b
0qKWg547DQvOQik8VEP0JtyOm2jiR3mjU8PB2R8fyeEP6vpaYHm3oNthBZQ+
gHFIhG320C+Ig55VPqF9KMhMbAKhEKPwNO2asCk6aWaqpI08RVcmM0vSOj8R
bIT+EqK72IyJ+e+Gx8bkw0K8aeWI/GhC5K3g/OZ0SGl47qz7xMU7nAnv2hXo
0QMU0zIe7hMZ382FEbpYyYlJBZ1NlhquqRJC3hzu6ZtimbeRTTnBqOTQpKFj
32FlE4eHKbSX696GyRunq9tr09hHUUmt+4ejTqLo3pekq3F0PpLjgUVk2fsD
AiHn1vm6zA+sngocC1NDMD9jsXmm0FQ3DQRk9oFkSwxcbQSGoRi3yksmFGfi
Y98dhB2PzAuAZgt420/kJS9KfLXRDCctoA776B5HNFmv5lTKLPiOOMPL5znn
t9v/8wePMocB4xTXuw8QnvcPDNdXhF4OFKyj5D989QI+uwiOSCisIe0cn2AN
sdNP7I1c8DwxWSzKzTVWzg2bc2uqs5M2GmsoI9kbGhr6gzF7L9tMD8TSeXd/
wYfdTUjl9seQG0JELa++9NM+P03N7yoLS99FTmMOU636Dj51p9FVBLrbub4q
ywrEEfCiaBqW5Hph/oUxICSuHVuALUr3kFggr4KeHghbUCj3DoZJzl6jXk3y
ceKjIt4p8wl6yxTwvb4kQTQwURPm+Mp180yuwRYu2W5BffOMFIfTh3IGomza
FgdAOAYh5mJDCAzvLdzi9rrVRv+a33XzKUn9ONz0j8MSwiPF2Fu+749zV3TI
5WOajeZePrcBo1rgK4DD/fbyKxEhRGQsdp+ndFuBe9InguWulayTVcwxFyA5
50LeG7BBmzdotR6PEXa3i5y5nPyvcG2JsTIQBRkJaS9DiQdSYoOZkFf6eJVG
f2ugNycAQ+mbgKx2GfBqT3elRiESjlmCzGSi+pkCC+M8dDGkgdKj91QvrvrI
Z3uFidjspd3rcGW8Et7FyYrpX5PXo8iWwibjXxUmthlrfJX+Wb6apTK22Gbi
tZ56hMvWaTuuzBdeJez2wKfSNBcDvHEGxotATPSoFOsoGZxajAuC790r4VIO
Wax7KSDI84hMqVH1W7SvfC/fwbEUp/lAMG+qNfpMv8aStpHxMLpd+Zct7wk8
ehtyWQ10FOvh+31hUgIKD2nxNr+gJBRbfp9kpnRJK7rZBQMyqauU53GPPNeY
i3+7sbBCP7PrLnEhK6hp/toil5Mltt1FyUEu8YOD8cboDZqvpuMr0XC/1tGm
kqjYcu+m7GmLC63U24gLQACoEu/tCVtAR5cgpUJwvc4/jqjMNrv6vvDphFdM
1x0RhyDNYzeRhZR9TZIrnnqglyzlx7nhlelxdeGMQBxmtITM2rUmGDcMQqp3
JLZ28JctgVchzZCFFLfXfoTMOOZt295W473m8G2MH4iT8TQPrxPA6NbE9whT
BK4re4WoqvfZYZhc3ERF8o7pZsGb7/plndklxo6g1hWbJELHncUtQDBYcL0T
qan+6dgW3EKcfXy1i12KIazezRtXbmo5aDvZNURYBdGg29lf9cCjOfWziB7e
dn7PFc2YBLT+LO/jh1UhJoyCPFf9unB/9k0n+Zqq38axZjipvLUSQgNv5sOg
RgPrj4DL3y588Jp7ASenzUJnjHNOEQO9TKECM2V+eMm1xLVBiqeyNmWjq5AH
ivpYj0xD4f9ja154uux+mF32JxjcQq6XNanNb1vv0ljy49Jgp4BuCpCKXicu
JXMXTlLuaPEf2z0JkQyQdumKEmcP1p3DTQIw+T+tFUqzAUWuR7gCD2WVVvQ6
n3TEp1Pc5vv0FFA9XqOsKrZFh0uSxrsysxxr+zVY0zZtib18u5q1tz539bbc
zrBio6+ZiAFNaD4j4VkQ05BWvoYSOtCw4r01dWAY8TbvfSPmHRJrai/3938a
RKjqkZv8CZzAAmfj/oJLmP8HFYHRLTC6IEAMIyPQzDJ65eLMd/MvyUsFwMp6
tQDWdBduJuj2x5yV7c5yhOMdlvJDVRGXHPmXwiX1yIw1OzJYFBh+V0KevowY
qO1MhqSRWBRivd95RMLN9m3L7fYU/8q8BTGvBtJwXeMsfv1XWXv0v4ipyij1
JtrFNh89kuCRvP7OYKCtnXcVUTmTI2uIGz7cQ7E+UKsdpdLloIvaIGjFi2gG
D8d2/LWVXeVw3ac1XGP+8rR9cWFEeP554JUgQSd5PSjgz7VeAdPkuTqPQmjQ
vf74v8Q4XUnRX+yfuGC0saYDJI6GyfUypAKAX2LhCUOsO2KffdglLkq2KcfI
okDYASxrOWGqFACu0sMAXJRA3hHQjF+sjvSzQ+Bn7irSVOKM05Z7VJRJJewe
Iv7zNykgmkX+jpZkrOdOnXzyXHtZVBwedC/HizlOBqfF+KfZQsU2Lj5Lap6I
O0QDN1LBkBYBHmDbbst15KguE80gnFgPIbKgarCxkfheHrZS7Lp/8QFw7VKX
w3/XCMCMD7yXveRpIkvQGcHsaYYYKokAcZr8YAuQ6eVv0mGiYYykdeU0lFvA
wxkguKIn7G9Q91911s5HqQ1fsUzKMFnhL06RdPlejQUZt0GB7NEEvbP44vj5
L9MPhkRdmoWDsgtvtjNZxakVtUZLdgI7EsYksxFsEDQi3lAXWwMb7tlanMGD
+sDSX1CkQ+qymmviFLj2RowlD7/Nh1CihMxTAB8D0x1SbCGFUse+dRLZWbZH
MV1FUvVGatNCQg3sY7r724c94fbO4RUHlMGjoXwTK5OUvw5gBo6e/TwM4NGH
+wYt57KHzo/JW+X9tAVCJUbANXoSx1+2BtjO8XuWG7jVCBmBOhm/t99maXPk
XAJoteW9leQ9S1Sr9kVFMIxsD6WM5pG80U7R6pEqeAPil1LuRnIAfPot3hLQ
0lJA6noadqPaBzy0/08GfoApmYyptMtPyPAiUhI0/9u9HVcdAiScf/oSUd8B
Fd0IS3vqQlzJ5j3De6eeSnbB0aMhh4HU34wXlV/qtEtTDeX63QQVOmpuIhAd
sMzA0IA171QIsC71exQhJIA9rlrbMiblns9iy1/w9usX5EucbjJ7PhO8uZOc
k38iwn2+XB/i9gZNas2fNfqr1UmBC6hrtFzkqW2a4Dq6h+WQxxkcU5rRuGN5
gJp4r55CegSNXwa4rRlAHuwLpSwaWHQ0wIb3C/YPkJ7wWmgAlTHYqcPeJwv5
JjLGiBnvCKJxAru995OCuhMXgK2rInL0/PErxq6S6irpuMi1CWNleA20ZU5V
vClqxh0bx9VZjwdeP6VIw7wWK0CN8OqWp3MumililxtoodSJ2BJjU8DLlIrA
0wbagLh8XAAVAmqbdAJV4/OS7St+wK/9ermELmgxY4odpidmJt+O9TxRvKQ8
UdP6LvTniRj86AU+IlaX48YyHlSDBxNaLewf3NZsLP38VM71ok9Fyk9sRiIK
ko/Jl4kgFwOTRUF39ilZAJ/qxiARoZfzxmiJgXHwxV05mPX7zFdAgWT7fHg/
nsYbSLmutlzZjndiNngu7DJPdBwLDrOrwKOYV9rY/1qXTVbfN1paxrQ9hLIM
pyhIA5Ii4s3rbhByDZxIBYDwCMpGTkBfttu4rUFDVmxCP1ri3g3OKFLgmgcG
dkXfjpDcdrhKycAGYhNQfrJ/gp8eOVvEGNuAP5nseE2zq5ERj7jrT9HoyMHJ
TNi0QCAQccUSDV+68l88fXymGKmCKafbYI2IBEY4xkVNdD4916OP2Fawpnuc
0IXBtY8A8WEvzifhEVApkxBznkHX8JoZDFQXftZWradDo3Zd51+h83QU1y6D
soKCpawncoQR38dyI786nTXYH5aR9AKulQTMQLh+0NXVowuytww4u0oLflBp
ZVmytx6AVB2eifR2HldNALOYaO95cQzubFaugHzAoaxC+AzqUd9zFsDz7gAU
DQbTwE+P9N8Z486fjowg8rthifGSb8HpUEB7hCxEH4rl9ODNAMSjiFWtGPel
iE1qP7lnU7r8xBJY+aPhaVgR3Z904jVKopx6SrwqmTt2QrmFMcSvX2cDLJ60
pC7MHm33P+JF+c9F9WHU3+WsI6hSQ7Vek8hhzJej18cSeNkmygZeKUMsFvgd
qZTwba43uzhsMV0/ZGyXJwktWgkM52cRDFtLOOGVuLckyUG4ffg+u+B2gvw9
v5TJulyofEcNKwPAFJJVj7oB2LLxuxrMUdx85GQ7LuOsP8v0Cjw944k+13fi
CjW4diF14wzvr4zB/HoESUetkK2M8pnr8YNnOjnAJ5wHKqFpee+KKXUY+qdj
PJPmjV4rqSU5ha7g717A/26qoV9E2Y8Rp59hDXfbENkc+cgEbQCiElqXFpYI
p4l0kl5xAlime4y4JQ7kCv+VGsRIme5gYcaL+BVc/e1Th2iA4m4SobkYP888
XKmscgS+SctBlwyEh2H9TbYjqqp5kIpbXjnPgBIUCI0ecwAT1YV/GRla0TL0
KgUr1YHjMt7gkQbVwzxyuWJc1nt4xiEt0O9CXysI+Si4lXe+DQ0cQrNleUqc
8CO2E6Ecc886bDlER2T/dw6/5Iyy3LUMP3utYqecK0JRVkO8JMaS1bYfRMdb
7RFwoJHnIXuMc3BD1yEMuV0HLZLdQr678x/MN+HlhxtCshj1X+bLjVwRgc41
3DCqIZyQ1lfVGmwgwRWZBb8ZTjHmVvTtsR12i4fJsaiFNQr0mxPCt8r2nDmu
JaO6DVjEPHIneyaC0xq0CFjERAiVK3HMvHMxLRKLce3/62BCfJbd2tBk6PRd
zj9fvcu047RDGaiZNNAnFwlxD8PnQWT2XYLifBSV2H3GCszyY1fq2wYTb5jp
2PKNgAIhjYvtzm/uEaJmGau4egeWQR+1jibl3olYLKsuhoqk4EQENY/HgA+c
gryMRKNa1pFSFuc1E7PY6EgKwjZJkXXXpLbVCVb/ob1QhRnJbFNdUDYBFOeE
K0GRVilnarE/xiQe0fbQAG5vUS9mEaNn6hNNuHi3IiuVKVwAi6WvQmuWIAD5
S/nbL5ixSLKYe5o9bmIPLRY9hRdn5KsdyFp6QH2FNn3nNzHQCefIFR33DIJN
jlYf7sQmZzmyT2fv1oXmSPDlv8xxnALyH11gbhxHgdbT37CGUzIatss5eKpe
P+bdHbx/TaSvzn6zDPV1LycQdRbih3TO69LsZDFwVra4XxoK8KQC8KfjVGSC
MQt1x9EdZhE6E7SQkCKgb3W+Zr+gSV8FsbIuvJOiU3V7RChyvGZPeRixcMjd
g18Ab4GBwkEz+jDreNEo0ypfmii5EwPplhbS+DxuVI5eqt6tAg34/Ka7BgA3
POeSQwRrD4JFCVveExjwebil2iEjfcIt+o/twsn/PUHvCCc8nR4bwuPsM+Uj
pTW+enl5VIoN9tC9vL9KVpTd+DLEXVR1ZGGKptfie/jCK9x+C5gsY4reNNhT
bqOl08AIwVlA4nzpL75MleJdqc8/TD4uKzxkUotmD7GURG0KIJ8ROPWRwH3+
l7RHpZnY+8AfLq39wzUJuaXVwxN5ufKTbhAXReK7dwT/RPBn7HpDDmcUEazY
cJN7iyvps4o0Cammsrvc+MBh1quLPcv/GFA+RZ5zGKtG06SuTbYmNhdeESAa
X/EjcQ3cT7Z6nmajT85EYkJOUXPpoasRr8xVXL8on6RMcW5nX9dXYPEz5odw
8mfoOfd97fgnAsXiqqtSCiwiicU7jN/zDfAhHdsARcOSAch8jrFwsbOju05x
Px+yu+DhnfEezp2I7hpsVuTaAIwcW9Ox2ap4c9lS+X02PVFcqy9cyJ1zpVto
2aBTGT7/odZFL0fNA0OHy0YSaDMK8JQ01XDgm3Qgpr2aKsOSaRaHRF8xN1Y3
YiYbJKYbV7/yuzdPkvmMMhg8ID1PFWmlnaE7tLu0P6X5vTD7AIjUVXQO9z2z
GEq6r+b95FPYScirzmpPyZhIgB0ImtS5kNbD6aASi+T9suRivfpH7oROxCL0
SsvPebP6WFHANESDavl9MlCY4xive7gy9Nx5E2l6jri0BTsqnKkeBodhwTr0
zcuQT8zSk4J3VmQJQu63VqoPDI58V6AIkoHpMjCdSActf/KB2Zfgl/DC9Hdo
IVCiiuoBr6o2RjhS0kF5Dtt7U8ouqJoix6m4SEqjFQw8XoXmINiLvChkLT3R
7Hbt+K+wYImAZkSzig7pt7z4WvTmys4i4eXT5UOwE1YPSa5fo22KvV3vwlIy
xTBftb7w7+XAXroalxtHid2xwD8G4xWxJwbaMxZGyEEqC0F9LTHKQ99A5OX4
7LQgEQb/Q+3oIiQzkmkW9MQj6KecsXTdyfbJxiLAbrOHCmK0xZMjMOiS0O+n
nK19krFs+4bOdZfxCDM0TqwpmArr9BiP8j0D7JCMvrc2zNKxvGyoWI36sG/j
KYx6mhtHztRijHF2pg2In7p/D5wlwROJB3dYWTHd8cnTLgtyScT+ylXfD8kz
dQIHu4+hnoqEQ6009cDw6zaeCGOivfdoMyNsdlSd5sqgap6PRBEJNzbXoLnv
etv/azIP50XqzhaaVoVeEaWSv2OnEysbren0QdIHDBzUdwwyeZk2o2d8Q2ts
Np1rhrXHVfpBee/PlErahBBENsGuGbbh1581CrQS/uzxwmreVew3zvy+Ti7e
vI3+8fT6/v7VtrtfBXtVJEcALltJ8DbCgxL6GKwhVF7dQ77OQWAQMBRiVnf6
WycH2XFDD6EsRDPVAZKxkcHOBUhUIf6WWEC+8+1w4Esaqony4SQDks7ViNAG
sRJTgJGqoes9DFKXrn4nyi2q3zzWlkWcjWL6cV2bWWj+WfqmeL22e+5ZwnzP
5ygKAz0BdW1i89v+tejpXer7Omra3HHbMjmlbT2Rr8cpmoYrSnT6EJFYprXC
9hD/sNxzgQmMtG/oUBQh+Vmh1hKJzDOnlEt9bnwHVePVmx/MUeJyr4Rc3fgq
w202U7KF13Cqkig1LxX25sLhFj1aKFdutVuI0mFCDY6CjKzPWqFLhjTznNOQ
BIzgK0RhnPFO0FyAmCBOY4nsCh8PNiq4i/QUDHN4Hff3o1SNSJV4UT2z2RBD
KFJTEMe1dBVe0DrBOeRwJIc4b7TDg21pXrAYrUw7+vFSulqHiucLpL6auDdc
gpaI80E79FB+hREghGQDgVtltFePJoRigUM4zmDDAs53TTg5UEufjSwnv/Jw
VklNK+NksWDb3BQeR0gvstzbKWgYdkQRxEwJxjFj82sD0oVHVOQ7fO1TB+Cb
8Qpih/ZUV2Mew8DzNPulIDmhYqiDPziwLZNAdh0dhbXkflfuezBEH53a7/xA
zlxxBenuObw3IthPJc5fr0isEwCDvCK+yfai9649CBg61qVfLRTGBnV+SkIC
1UABFqR1iN6wzF05ZPVP/gPez3IC4z/RGelUamUgI3gvw9ARrKBH4TQW7u6E
TVL958xScMCqEyybOyZKuVnQF9vZWXJk6ijIyr2OPLa8F1T/2bkvqlgJWTc7
lWOEVkJqfQEPPo/7/7+jjbpNnxZPz6hgR117p0AXceNv0i+oifh2TrBP2J21
KLoVlpmCWWJWyQeAEYLNBXYx/FwggsA+KTl9yAPWUDFRp4ZrBwyHufw0Nw/Q
Lu4Gm5mVoFIPy4OyYiJblf+lqfbzhtgbrLfx997eH/ne20apmxDNOXjWbNfF
vb8piQIM11xVpRABtFWgOkG38CZ1CuPRSQtkxozXp3P1Dac8IlbZ7fpZfNt7
engFX40gEUuXgznKZbkMlIKRVBPT7xIbZLHZ59o9XXCJh3mi5BvEoaGZ93XK
H6ZguUbMHbltz+QHp1hb2yRISrXgUvy1fY328+7YocKKI4uqy6in7dMOwXuO
S1SDHlOdC9S/FdOAoGil/IVAT3dfjMafZXFuGUaoIvXueWKdX1G8snIzwA1j
0kxBGy7mNIj9T2+nfcHspf3UPdB2I4Ups8v+4PIhHitl0cQ++dwJ4AazuHly
XzsCZaO8LldvIHG6PvhdVISvBXQPu0TFdPnVk7wFlDcWxTCoGBp1sNf3QcpG
j6ZfCf5EXLGTVmeakflcGsHfDX0L41pyjOgf6EnzyDFmraHhNxicyQ3cft9k
lJQBx645MO4S+esybX+q62NXl3FakllSDIpoM20jBMVXF08Kv4NHYPBGNN5K
V5rrD4uXk+Oe+ZVu7JLJGAw8/lOolg9oHtN6KbJkU/3EF4JqcTCJZvhS+W6s
WOBZtEy/21SG96Vi+Q4Hq0VjVIu0lSGwZMc0kUZGwmUOTA6yv1baCEoiaIo2
voPiTVwsJLPlMTtKvGydrfOA9eLcQkWVetQdOHqVN8l4W/CQzuM11yL/ixiv
GX19Zgh3eSc6H2JPvl/+kUkM9qQL54oR5V0ZYw08xxUx7cNmTXJmRqJEobYV
QPgnJ2LIcvAM5JjnIr56XJy/eXeoMDp5dIZQJbjVMFhi57kHr1HTavDP0XUG
5bO38QqqB5ZtF1HaKHQ7irkmrq79ho1mtXO4heh8CEqPVJM0+rKD5UrsOpux
orX7tReaDAfFMbY5f52C94riQ8UmwsgDeWYHSiVsicQwhOhoCVX19ObEfB4D
2PzPLYwDeE5emMtjfcsizLbgZlVCfsPOsKWhL/GKh3/Uj0LCjiXS5Ko4fOMg
1wkrmr4HC3UlymPabGCd0j+Yexuh8xK5NV/eRbwX6T56+SMiLKDWQTVJrZ/e
FAr3o8d3T55H5G5KR5pjaDhUjj11qUxZ75+6zba+LP82s2bxmdtiEgkZcJ52
lBi+u4w8v5geelnIpgdcFFIsJblj6AJIjTZh5X1wyNfC/4MAMIB92spYSPL2
5edt3cUP8ZtV8Fr/sKD3RE9sTbTSn7hR1l/SVzmXsqA+PgxB9SD7BUNwn4dJ
w7yXI64KNdqhX5B6zOU8qbOQtT3oQKHelohUqmsaBYVcORbp848HNzlLf0Hy
EK7jCdPYvzjSJg/hFWXfcRv5aXa7lNu5xjiwfSBkvizSMJfk4n/h9vEACIcL
5rGuHQt2kJePs6pUwPk0XZlHZxHGnUP3TkI9IsiyYWQnxhGNuravzpYJv5n2
03SsIgxwBfAHQep9AeapFcjeIne/lXR+HU/OMfvbmlKINgizYU9CTBBqXm7s
Hm0H0D8cyy8ICHMHn4l127snvTz+oy1eJe5aGDIa2rqO3UTiC5TslBiHB9UB
a2FoA9iU+Ko1JgpHZZEL7R/4LEqZFh8HJe0/RsEeHxXUO0xPRCPAB70LMhD+
3549KGCp3Gmo1HBB5nJezbpOmXWxXKyCcYC/SpvMgAcERxE+eqhRHbJJnvdu
Z+sQ098VFTCNpPR4cY0D9j2aUvvoCFy064N7eW5HSacEbwIN7Vj0juoqUxr/
z7LanxrK1evf3ZibJtrwyylBIhonmhP7vjiGg+S9X+/ZAaVULJbKPWE/6uUf
ps8hl+JN7GQjyNE/W5mf4WrEidjXyqsJPVMlAP+8Bm7kEm19bT2s6v4c7UfN
OcTgLE098/YFQKVw0633PFc/MJzFrk/vt6wEjrw+eH776h1TOfuK4UOONCYp
wbzGMYFN8jApcC1j7vW8iUemW1/gS9uyI6sYVwqhGJyy88bqq5AsNJ7bozBJ
J/3mWmy1FtEfZbggDqWR8yoMK4Mzy4Xv//9RkiGTfW4eVYtFb1sHtyKyJoXW
JqjkULzSJlb/yO+bgVjj5e4IE4uw5ymccEFUhXY+zop4YFMw8jiyqozswpqw
lSo7rVMhkhS84S4eXmfq/HkG99qwgYaB4aC2Ascv8x/2IyMiUKKi1MCieLsK
/T5O3n7Zz5rPUNB8a7+fWEHBGUYL/wOhFRTzPJA8RwaWXuJH5IB4xB6JoHSe
XNXMtEFQ3tTsOCdMuBR5RSZ+fZX+VeQ8mwycPNNqFk4vt2BuibD9ISEB6ZUf
93h7gR3Akr1QMeYyn6NH/uVSUmY6FB69AdmnTvWVAE9Q4FEamHy/IjAXdD2t
RY2eqhFXOXpFAJ+8fPv/ZdEeKFwoX1Z1YdzRVKgXb5l2apNg8xJairSZGLcj
EyYGqEJ87Plhu5B+IbrY/xDHMD7UH+lM05FR7ZBvVzCk4w/GOSHI2PNe66xt
+KRPJyzfrmzaQ9twA/b+cXCIl7WGlMS1mPisYsjMGqRtPgI4qlMO4GUHS2qA
45e0Q+Vk4yL3kc7R02WVZa1gOBsz98PGJNphosQ/oSkXp8X0WtqffPQjcjTH
CuIDqWCqeffk0RvkeUgouJfLfWL2Q76BhvTaIKenoFvgAOMSJ7sP4Cs/C0lI
iL6LG4yVDdr3IzhEYB92u/+UbT4pKFBmnH9nlgXTJZaVEsBYNrnF2l4WJ4Jw
duADm45aWAemi4WjP6jZfwd941Zn7UJiv8bRlvgEiOUbHWlWIdnxvHsV9GfY
vIyO0bPcZBk2laHp9nemEf78uvAUCSOKcHEDkEuSxxou9RutcB5e5fdJl6+/
jjH6guPoToFY4Zi+WwGLzScsXIW5lt5Fs5K3J06z5/svFOGsjptJFcjrklBg
Zh1IeU6G6qkeTLLe7/JuNhxjPapRCRImx24IajiYnBhX0Ql2NU+/SmywRFpb
d3eK7ZuJXkbCLf3WVFNtbqMqbFkIQcYbCKHSBT4CgKnqSuLtqgZBDfp9guU+
As0iBio8hiDyeM7yes3butus1C9bKe1Q4x2FLv5vuFIK6oF++zHNWz+gho+i
ZosjEaU3HhUDLyLqVnp0VAd8y01IatOfs8hzvViPlHgEpi0hrePW9GtLmIHZ
KT2UZG48vZTZZZ/eMigmmX0H4YRolj6t3fturDY3C13a5eJBFV75QWwe0bxw
v7Zk2Q9IAiFnH6Qo+LccWXEX0+Eay2A8RL2EIXTYStLjr8wl7p4mWQdFIGVT
o6wUs0p0lXnb+O0EM+2oqirB5ViDgrlagvu0BWC+OcTLXQ72UF3i4oz6G67x
TZcAn5lVHnf6LlIYTO0gFHv0QJgjtptJIDVEcUq1WZ7bc8MzqZnVhrUD/h4Z
kkNJk4p0HuypZA2gsnMhN9KFSk1bcMpUUqQoixJzpVkpSRjtw3V/7ldnx1f1
ZNAz7l+lZz81Tihy3pFZlLwOBVuz1OmJLDF/4pWCyRgBc0CTThtOHMoCm734
xhxSjgB2NvpG39Nk1gHkbFLqDd83UpHW/Gi21hh4xYtAIRkWafizsYnR6c76
d/4IDYWw4COKJwTbLB1al9hSMZWiHw/etEy2S6WDTA0kH+oxN8p0CXmtqLwZ
OFjHxALH5JGm6y1zFNABXPjOTHGi63bD0GuEPp1DdFPB76jLG2p3/0+RxcJ8
EeOBgpd9x4Mok3pu1mjkmczpBwaoJuyFtzy7XQJHzezDaEVlS4VTSWO8rtRr
1Nrq/VWoY8t1dz1RWh84ubXNZiuBa0ltUYiqt/emdHWFYK5O+z2nGMkQoRnd
GEonqZSCLP2ykQlkKEYZjZjqhccHSrBOevUI0fLu/6p8xJZwRZ4NYI99E/ec
5PB8NxV7DOXZ/KyLjjSJd0xQutAkb/SbYmxvbrfxS8htb3q/+Y+QP8806VKK
YfuhMYjdtZEb9azptR+VdT6ms3rp2Ph294kBDdUljIcTb7QnkdI3sZPJuux7
AZj1LrBVv9XheQ7cOoYICC6gOegvrzxvfEhH/cPklJ6IczMzqoJu9FcMdJW4
ZOx2vp1Gj5pGEIQebHz4EEy+ZKZ4Pb3pUbSHpAlm8oehgnEmfipFK+BFLo4/
v0U03EvzRR6Jc5ONewjFg3x6qiwUd9Tu7KNd7rdqNKkwU+E8hcccoqsp6zlf
hRjApdR3zWbazjOvRLLUc8Cb626+XSoVC7rfLLM5GYrRhmFOQL9ToOMeX6x8
OlTjA/DPIbLmjuI3zLVV0+nnhJMHEWDEfPfif/+Cjj8RwpCAs2iZCPLpXvTr
kj2/4xITjrckCiF79+ezWoZVK10owP9YBTp4dFv6/jQozwEFBR1Ou34ioLGc
0oGoke1Xz7yGUVle02SHTwUigL25qyUf9A4IPsQWEIX+s+XHvK8vjjmN1uA0
h8Vd/I3fubO7RtooXyCtlZFlGXDWZVJFwdcqKkrWtlZ+RMmAKRvwWjwccvM6
MzmegjWZ08tXS1jMsM2i4NwWzpcTlx8OHQd0b2oU4bDE18OZvMaw09bvAY6J
49lv+40xyL3OXkZR+ErKrcHFJUfWf1HkSJ0OHy2l1I5dTr8KP9jq8VUTl5/r
L+FAGQTN8o7+nqY+fzXc3JBZV29/MelFp0hu28ZSRfXHWhHtILgq5Ka2ILWZ
nvVohXJS4us+Q9iTMNj5KplpAnNU0jnHuH9lM1MHDnnoDg9hUt6Ye8oLSbz7
b1yLPXjmkAvrap9hZEjGG80PDowge89odbY9B1Z9My5OiCqrbhzR/AArug1D
oHr35vltGRNNuyV8buEWQ1DcTflOD2CH8McLFjJ6FaPmZnh9c+O7pvGC5CxU
wK+o/j93DfwE04VVwhWhKRAHNA4UEC1J2H4zx6V7IqxipNu5uoojrgTG1cEV
gholT0MuxQSFtyzIYlzrBoc1FwxXQOtI9HuGmXlNELnCh4aMumja0Wj8+I9t
mG8C5jOrtfca0uLbAsYTMGgiCZapaXkYEtwODIRuzahNxbHCILjywF6fhIsv
S+SoWflPPAfAzcbW63NT+QhG0Bklhwc3+ePm461TZKx4+X/ZvZxx5CwzAROB
IDeAGGxwyqjstBUA6rrw7FMW4+XJWLewGL7Oj1pGBytOqw5ettJQ6E6Amw9f
5BalyTH/kSId6HvaJ0Xxw9Om1li2pLQ/q+iV42kp8HYwSC9prmIrSMXgvF9r
hM68W9spYclm1Dqiwx33TDAyz03IlpG627n2fzTcYL/EBJz4QiehsBEXx46Q
QWJPEiCcIwAIPtOwP0QDudq0WPHN5R4RmCfaCULZYZuWRVD3Y/1Gd/6oX6Rq
XmoqThFDLmevCQTfNNt4im6TPlY+eLvMnMxaSERV5UlfS/Cr4Guw8pRfk8N8
IS2SZaexbtF9C173nIaCQr8zBLyZ/KKdFPYK7pjH6K5QSAAO4tf3fFAERZ36
pPS0/liAVyqwPcs9ilQPx5L2cNeHMYZ7oV7RzPlTAFqpxFBX9BAtTlPlmVyv
Nxaa8hWFbVS0otqo9Hb9TcYS1u0h+CQWdYupIujEq6gS5p6I0zMzLR4rYKn9
G/6CyD10YlvfqHRd3kIkjHirXHn4NrZLioetir29ZiDUY5OWFeBAstN4Tp3l
cWb275r6E4+4kZXjz/MCFypNofwc7brW+7nh9fqo0+dlVXUVgmhydCpmXSsx
sC7t/yLlSTSUgv8WsWRJmI27en7jNPSHZ4+ZEu8RLOjweulOzDQmtpq4Jl/u
zNnsocmHs6pv/Vd/EiswN+Og0/mTtLzelldfuKj1IFspVmxt8raWiT5EBZW8
EmiIwHgkBvsprTp8C7bmsMkkjtkRpudmaJ/3mhfIwzLE+ieQcun81kOt2Z1u
bQ7Ddg5yZNJf7Y0A36jE5OE04dEqqCrpTGpeSjCaG+GC9Cx5/Y5FC7Qh471y
3vbECx3tzLLCVxkYDaYB94zkA0Yxn3COoSB4hs1cAnI6jnsgyP6qh0jeluPU
uWJkBjIRxTY0T4O3voTTOX/CsvZJDImVPaTclbXDDv2kWc106n68tIQyitSt
yWJ8cFWL4/at1AvIc3J2n+Wtx3nn0TYl8KW20gDhZvLvQoAcVgnSBKhGWGDk
0dnNwsAvF2LFPAYIiqgD4kz8uFxpd7eVAqBxjxeUrQcPemKdvjcNDA6AdN7R
qiKwLYEXJnoB+kZlLniE9vxH3TzuoGcEL3wLm5UHjw9Z2dtdW/CMVrVwIM4R
773eDpeVFiFGIRZBCVuUsq9rBkfbu/dk8W9UTPT0//WsFRtOVSzkeMqgVps0
bpnZEwcNfPTRJ1wGkysWDtrRQPfWYV+BaX8RzWe/3T8+74pyaSHYFSW4eh/z
Dq6iA4xmXInBAnbjEysV8JGC39y7XDz3ODEEXsMqtJO9SXE0n5XSiH4ojtTh
ZfealGtreIuePLcCsTVtqY+4ppGu9bjpopLvcQKkjEZjc2MEYJoAU06BssfI
AbsIDc/VJGBYG8SshLmfm68joe3VDr1mRRz1XQKYCeG9u69RmocqqRiKkEXu
Z8XaYWOr71JGgmCfFl2SqepG8OYS/oEw59MdglFsawE+Om9xvB2AWlRwLD1h
bwysAgLjdXNfynHx19CWOdan1crTjn/W1475sf7vJUgwBbG0w9eljo1gUCue
y1UpceOCrrg5NyrhQVLE71dxAwN5curCu4hvAFxqsw+sbXkpxONlpPUUptkK
MrKmcGp/A5Z/J0H1wrmJwsmpknG8uWN9MqSoNhaTfBiGyB+cL0c5lajhttEr
mToEJlKhWgQG9x/Aok7UONfnJqZVRuPgpdHbvL1n23utS7wc68J9KtY81ZuK
+QJacjQurG2dAH9XfkKjZscWmCyT5Cre5mN3PMx7XKYHMY/lZAbjNDd1WpoN
HgeXWtowGPOFNO5gi8SynLNX5n6wWgGP9TXFi1/7j0lu+TIDW7yeaYqxW1XE
N1NAZxh/p9hMhf4C7bUW7VUim4Q31FBAZM8i0AGgxe4+7uE8/Yz/8/KjLcr8
UktzJifzmrDcJW4QTZWDoEY/UFcVRfXMGQBLVPm0lVMPwf1DEWbsTmOk6Q5e
2dJXC0lPn0ucfDQBMh/8c5e+Il3tOCjqBDMOqhu/O+iKAL5dAkGE9gKYckQH
2THB8NtwfGhSKD4HnJ6OXIs8kTMSZ0kWVkUV1dIFjt/Zo4kiEdomT1NM7nne
CbhfbbHUhtYiR3BIBpWrj9SzFsCExfGdIAVAsSqFgoZcnD9ZQSqjyKx6d09d
ehLxDLgPp0Y8SMaTcsrlDWNy4bLNBWuPPZHkQYmYCSvdEq5iK6byn3ccADda
3k/zJpBLi9jA3vsg8WUpXjAW//ZfTFUKyb+W0HOMaTI98lGFTibQw9uJO92N
dfCGs4bYNcID5LlHDKIRYq4uEwBw0br+EDOMnzgZ4pf4cWxNtfCENTeJnMAg
zcUNSifAwGRBCrx2VF1pRtyHRttMxNQ0WVoHAmPx8wDF0mCx0uW770E1OBQ9
9bKGSXg9weZooYFc6uL1UkF2ZittiyBWX0iwdMy2O724n6Tua2arqDYu5W23
KjwhbRFCDEvFJSAFSfaeiyyFzky19ImJXONVa8BXsEkcn8bFhonpimWPse16
RPEyTfj8ZOpwPEfQvceX+dYEA2viwsB7FpNusAfLRHbqB2S1B4Qs9xw2d7GR
vvJMv5l2wNA1X1pZvcvmyNS3ddK4+E4LMD24+sPkrKVnZmW0YOSVlcV8wC2j
xzI+78+gm0hXtMn4eyTDp4ZgBmTRvPtkE7cwj6htUa9O05lqV3bG4SRP0/fz
nr8+W9AcJLDYUyRDHLuCWm6O3FAyWMPg1r2s4iqqQxinAWaDAfIUNwLKxXMa
NRUsZ9ZgJzXeiw5jdZWOmHSlfkGV/c87lIDeDe00SCEoMGn3KANgny/KGDii
drXRF/ogLUMXUjuTAV4EO0/R8UH2YQBu59GVXFk3PRoFjfZ3KPZ//wcyF9E7
xTUxQHY+rUpmIH40wfiJK0FpvcR+qMsAglhFKeK0qnM2VqwrFDKZQDO/0369
AvQx6donvX3X9JZXh8FrxhlMDLP/ChCh8K7N8bVRNbVjswFOgjcMIchVri9R
+vueZCRTrGSmxD96JOjnYYZS+YPsYE/rCzaGkHSwmi8OljCiXFzLsgqZvG7B
i3G62hL+zdbwXph4aIYTeK8qjZCbYKO7O6hyXhDWwdaPLfSLmJJUH6qmttJ6
FI+X3SOZQtuDxG26XMrwZPfA3dhgrtcPAoIQHoclTI+wYwxzxpnfcN/xfA4z
5Jbl5l2l0zvkPr+d6ZZyZtZrYVFUaHI/sUIjsPe5a+94v8EElpBmkwFRIjoP
I++1OMDCNdII0WJ3tPurb7xgCNx9Aq/l0y5vdpGDyvRnVLYlQe3zzf9Jigd3
nJoQRgUZQGRLbj1bRFoFK4+SULj9PFA++skO5i2vD7y8n4pCPYWzpjEr24Pw
ZPKNx+yYolJoW54xNztepP81kuVUzy5e4FWL5Xmm9N2P/V3xC5vMgmE/jfRK
VWvbLTylKZPceBVe917D0fYqiLWPoe6KYQ4We2aDlipPsEAMC25CLwsQoE/5
rqbCVxWk84lvNNCo4+3EvoBZLY3+l/1PN/QTOvGjy7pl1uc8kjyF9QjqSIBk
r+bPEz+1nc5b2BsTbnhcQ+hbaXyVTrXQTJ/5A7qbVmEly1VM2WOssvavU9ON
7TghlAZQx8dbe2H5WCsa2Roch3zgAk6tS41CJAxaGEVZ0qX2WXvBKGFgEkn3
gvqHkqVpi7f7RgAe/0QMKwcGoDi0grpmC9BcL6+qv3V9hTRZbNbzhdAoHAfJ
zC4VHwH+YBPvjebH8hqo0x6Pamh5ZIrYqeXa05livgbB5mCIUnnJW8+QjpEm
6MLzkOwHQT76Q7DQDlHnXcvzshExtuK8covcmiKehbJQiAefX4dskLZBYuYf
deIAnPBW8A+tUAXombL41fyozfK1zPqtWmsUGElno8ifAi+Ac6guEnyql0pG
rdzIKnURfh3MvpJg3hjcxatlfWVrX53RScHKOx0VWgK/S9kZbSg6fHtxcIJz
DsHsEqGFHy5IHW6W607+2XZRZrlB2hQhg2TNiNu2RtYMsNyOHN0iFbWvXRTN
UAEwiFZ/ulddY4CX1MUc/CboZPqlSNfgqxxdqIOoZcVsUQiQeEgfg1V957y5
fcxz8dWUtsQMFeGxPEu9Nt1ifRPd4V9oZVf7gmd0kaHYHIIxImkHOcBnSjUY
1pqjINrXKM5SkCQCAkUfkeIEHPXBAGNcYoJNx/4XWxlBJlRj/2eW9z84Dn90
ZDjRiuFfRkVATuCFaROyWqgppM/9bruyVSEW0knq/Hs2n3hwqFO+vlzOPxDJ
u2LBjtJEu/NmdzwHSHAPVcsChDl8o3Z7n8OW0bnx+gO1epJlGwBmSCTkgrDr
xqXATwmCpqWCBStu9ygsG1+0WlzZeJifFfK9ea/6FHCLl3E2hNub3Q9t1jQG
dPwGR5k0ES+xH/jsAy7g7ollZpEYY1m3//2bi/gvGKCRWGg3uhuyNA3M2ci2
nOki1DRSDUO5psWdLb+yhjZPYb/fDElI8FxrB8uD3njGumDvlFiWAf0evswk
AfyFKd8wkctG7msK0+qJXofEx9dFChIEQWII88CWU3X40K22zrSFB7dPURlw
RI1n2RMP2t1Se2c2aUFwvT5ep1hRrYvM3rmc8b3W3vgtkbbbUqaC3T3HUvhM
RUg3ph/qScxuWIZ5ejPLAaSvp955aSVZtAexb33ScGCJoviYQpP3m2vSrpyd
HP8S4w0pyAyno8bxvNrdBuxLy37smdLfblofHfxFye+NsHlyxgt+cfz8Nm3u
B7e2EKhcES13cnZBd9xLT70jR9ykhPcGBfckQp6oh2LfyS4EdUJro9PsMEPn
d5f6Jv4mdku6QM7dZ2WvH2JcfC9ErclTmO99r/H378FYHXL54mjp4Hdm+XG/
RBzUr9O4Gj0f2yicC4mPFW22REFp/K3TGR3oOZe9Yq5dX3yHmM8lGcIyiT8a
AsXxunP/OJidl4jKbJAnnQzAqITzlZ+1TUp3OSKhamc/fm3am4zNVoJ6Gudy
iEzhf5LhbFYtBpQbOh68voGgMOpTHi2/HqYh8Lr2q4bNQoRdDtYYfwGnv1Ij
kAZYMAthUKDKOYToPHzHe/jyFW1g6m8y8dHe8/tZbDJbJR1jAC0iKl5LY4ek
peLOyd43o+oJagiMQxaOpFJRCi7U1TUMnbomwbg7AhXlyuwEaerRQD9IhD4B
gcdtlL8cokibQMpCIGQGN5xjPHcI67g5YYWbeeGIDXmmGGKzZvP7RyoJT8H7
/dvZFlO3/JWuIcPaiBReeA5Yg51NvnBT9h484aW7atdetXXEvOPCKmDG2GyT
NlBE2edbwt7MQ5Lc5pxqTeNw9pXzRvMWnKeRC1GC6HaylptF15d5b0aVpnkA
rcCyoXwT3Bec+Pd6noNfPR4TEqb+4NtXdg02wYwVAHS9/rD7NLklMNH4bZUW
EXmgVMpGQWNmY8N4TUq8cz4ngNWQAaMVCyPUpk7dBZBn0lKJwUq5qQ+8aBcJ
cbCyo4Oe8YCwckRqOAHzqeV0PRzBF6UcgnEiBA/l5+68YHX09Tiq1uls+gyl
vkoIzux3H9p1gSQ5axwA6er6KS38WGYF4WWSqyxnUrrFfZX6Gbcij3czpZqU
dkEEErVU9ZlZus2CjmLwNpYpvD7R5aUm9tLjByOcRHtxnXA7sCD3KoWr2+oL
1RAFJIaUTf2QrOvlte5iGqc5U+y5qrgW0ticfD29XumErqtPp81BevTNLsOL
dXSTTWKVLYY/1/X1neM7c1b2rbFa/UwB71UyqEgsuUvMcODkmmgpNupmmt+l
yqnUds8VVnbJa5So6qBayoZxoRH4JxhF4v/Ne8+ZGKi6g4wQED56rJIN6aNi
O36yxYnDCd7/oHEK/tek2ZrJISbbvBPZLDuKxpGb463PuEuCEZDwguTgklMf
4Fwv6ol2VGlxCoteFCAQ1CzlSG9u5m5jzY5qEpSy5PDvCo4NAWdMlpXyx2jt
bod+649AmEaDpmkw2H02tWwl7S0o1O9qG+rZsjI57YjytOKEGttf2lQuZTWY
NmUCaH52YZ+fe2eq5nNTnknvlDl/iu1VHDsKLO7MwHVZCnqt+9RDDY+uXpLK
PeQReQKh040UsLZ+WXKYwCJeZCT3Ob9zfFDeOP1tpH026vf8rVzo3RdEIuGV
RY/aFXxEojinV9/wBkHNB4oS5Pkp1WYOz5fLoeJF3DYjADhCrHrRpYC8Nx6w
HI5sXH4k4ArBusilHxqB8/gzLJRhAwQ+0VEX5HK4hcgjvO/IW9Hkp7bG0Q2h
+UgdWfZCYr6qHiyNEuuh4lAnQBigVjhn9xyZkkRWLOde24/X9+DbCwXdXrec
Un6hxTBQsDekvyp9N/b9l7h4CF2O5VhiMLvkOJDWyah4IzHvFORsDePR0qLO
x8hSEIeihapKACXszdXkmxrDB4m8WQZgh++b6OFf1y7FuTlDemc3DAWGxlkq
PIJEAwFL2zEwoPyJqbDqk/LleZO0iOAZik+nvvYqbeh7ZlMYYJzjHFn84W0Q
wmBnQCJCA4Dv8TK7C+VDCpmf7fmbvaZMlCMqe6woZYn+0lr7C/7XZZKwBBad
Xh46hanB7JahKBavnVzGpdXuCdIIKxXA0KpoUl6JesfxHlR5K2SG5Aenzx/N
Zmb6VqxnySXt/qL1hvOpQtWTZoWLqr7k7QrUYLAPPuhYwyJgaBhGGWtCgOSi
jrR+GaPN8gemsfY5P0ssYEurklLSPPQYIksjsUpEZk8VAcZontcdBe8nAgCR
2dnmF5bb2x82xxcKhe7uY23WGmYTlPfwS2BW9WiJd3QiAjbGgCmERWCTlk1X
3zM/BD3xftedq3+8izjzucElhDrUR0Gu1mFaOiY5lTOxHAnPR/FytulU4oMY
GMRwhyhzXvdC/HrQ+OOrXrA39ReSnIXzIB63s3BsxVQsExTIUwCEIhrvumgu
NtRIfMZIE3zTr0+btwCj62kHgwbtYo0MCxjpD9l9lD+etNBAu5/32HVl1pQB
mTeroAJEv7aKNj9sGfP7aRUBsttf7md9rXeMNL/ZTyabwQjZUHGPcNn+xL8+
5Ke+smoqgSzFgV9MAUR6eRFnA3bTNQHOzeg5Q0W6nimmjCHbh1TTwKTvvJ0S
pNzSYFsTXMFzVcE/rFOheery/aFvUOjETtbARbzAN56XlrmKD90jOHBX8uVD
yMk8U5ywUQ/LI5bHKb5HkNOi5CjAtNpcymTXJ3dIwvyzr8TuA6CPsPVMfOUH
FG/pjDfaiyBs4JULZ1I7cOR9gYbgngSjx5tnHTOkF4gxhXX9fhutrizGFbga
GzPag2MPqB7FyaKv2ewtDjlAqbjpGvcx8NeolKNOvWH4/cSasH+lrADjHVXF
J0X9WvkyqiWCG+6WDeYvWijc02xXVn4Mww8cpGZm+sMxL4ad8ryTSpijA0/D
VS+gmqlV5+ac1FbGpdxF5E5B6tUbi/Ye4WZPENSltWiDzdm5mRTY6GmP06Tn
0P8EdHIV3kYc2ITz83AbRANg48fKso4+u4gVG4EqxzioZKxS0OjXozwhQCm2
PchW3mLkwKzmWeCrH5Gus40AEjVzaEHyJD/Hc5FS6AzMRsMZKjJ5/3rjH8rE
n9ed8EplddxrYJgAnB/XcY7c4KU+sjoAeRmssvJ/5NlG31ccbYeKJFP5MOv/
vObQJL4955EiGBMqZ/6mYWeCOFTBLe8wWsXjxLorHlSTGElEviv1E79N0Vqh
7XT6vS0zkebCC3p8o1lzicWPq33LucB5hdE5X03Ssnkkpe318KuiCZjZC1Mg
6e+JP6aLJ+XeG90id0SC9emAU0kcl3sYVO6zwr0GV6vMxrkdQsQAHxsLs0Bn
oaD0U5IhMhC+3mO335VFaVZN4/qV5A/xTFbXEArZnF4kk3PFtBfm8T1vUFjK
tjohxlEbWO/molsqMb8Hu5+9S0J/7tZ/TBMMNrh7kGqohALqP3AkyYUfQXVC
CjEgUYmaZsyyPY4L0RxC6m8VwqhP8KTWwOvt/dIGDHNNzA2DqHNvl9JtgwG6
jZCLFSt1YG9Vkq6cv9Y3ttQ/BjFyWl8QZ2at15gaA27bP8/P5Txi5JxylNlV
KG5H2JasjCOYzK/cQfN3bstPQgh/AQ7rXChnBfWdQIV3em/otB6lAb3eQO45
QjaVemiIIbIK+Tn+/pyfByFEa5eh2LeTz0d+BP54yRKn7dTZhYOJtmhMg20o
GvktTfqZTEVK79MxWBLBuiiQbshAWgMBCwvBDUd9/CfO8Dvr/lLm7/oIwl+u
+P0PKPE1jXHDePK6JFYpCh0LD5Xzf6w+03uN383ncOMgkJMNv0g7lEk7EIhb
5hNwvwPJ6W/xRS342SzoJCQICr93aQjr7edt3bmKooGFSy4Jwbg+VrfRdy49
bhoRLGFKC7rUB/YGFEWwaOkGw65XzGtwtQexsZZL+fqgpqUiNOQkypxFvs9Z
hC/70iq9RXeKEsW9fh8PAPFl52YiqeeeDISbi363i9LLPEhVg4phmDr5alYG
3TQnG74YD6Mn7zObRQCRlYoZEB+E3wdesFvXd1SaipGyuMR/PCYL+ymeGTC6
9d4jkNLsEn3p9uwz6l9dpEVPvtdzYB9OU+OKl+KzGf8bEq52Gp5wg5AxptM4
4oqC77Ug4o+007CYi06Mz9B+dPPt5m3FWTjku5706uz20VIjFdM3Exqj4ADN
6oBK59nM6g4FgRXE9anvOmvwvdu3RiFoqlfddYs4POpSlYfioAjO0yqs1PFY
OEG0QlRXHvrhrcE9w33Tif00iEegiB3TTlCnAObupLlWBdxdVtKIamIBXCvu
WcT40mnOtua5HNA7qr+lHTPUzM7KBVoL35+RsghXcQ/xkHshInFES5/G+4Hr
RT+81aHWfrcI5T8olFnR7+9hpegrVYZNsNUXvjrwkL81x0Oz0DzOnwkZBZ8u
73gAQitdJhJjGOcNJ0kDT3ny0FVfTl/yCl0yWFg5SkGe/Q2qNRL0X4qqcukj
Vw739caXotC2IVnvgCWAFM/x5xoRtGOgldOedFIv80K0/m4xfMpjggHF1Vjc
ivjRxsi/hbTHRYJGO9OuwmRZJUqkq/peHvf/g079ZgsHxSGZ6/Wlk0l61rPh
VfgZHQUnLIBKpwgP5gW1yfWKI+7n70f10S3YCk+WVRoUvil41z+ScA1OqikA
fYJqz0ZaG9rC2VvojK2k+LdsEG08Slh6AgvTktJDl+OoSJEjHa5bBxddH0tO
vs9rWEg7LyhItGGBm1LbwrdPjxgVSK6gCBqiHVHLWsIh1hnoeGuBx+vOxLv1
l0yaA1XI4XUkcPkttAnNeb5RhmzpF7zapMOdpPFhvTtVaka24NRls1CB5ueO
hzPVVRz4iyhXuToIcpVo571Kr5QHO/dxlSJWOHb5ic4PK1dvo8sQp2BGnXZ7
r4z87/YV2YRlp02Nmrcur4oxq7aXtXQ3mcIuQ/pucTzKRbZLEsFSz8SgZIB2
aqEZPbSxlJMkJ+x7d2kTBO31ZnivvRMOhLlMICG3pTvf0P5WkAoFyzvITjag
A0awiUrqc2kPR/nnCsTXprvOUpWcF97y06KFIwysIq1sxYbAQa+fFQ3QV7w/
yOD/hslWPlGzQs+3umVzQjMeaf0TVGLVdtwj3ro+sSEbz9T7wqJ3baUA7R3g
XHPKgKbMQlCTb5y+qrpX4K/M+Rjuc3KJvKCOaawHzErk69WZdWWD58u8PO5r
yu5vjEEkcFeljO9Z4FCyc3BTCecXG1V1ESoBnHms580f7qPivXgt83Uoc9sy
z1lJA+NKZiclwDYOPzaZJ/b6lOe0M6E8Q/6hTutZ2CohPo4+ui5IamtEhKAS
9U6IPX+J4p9oQV1/oizQczQ9dC3PD4jKdQflWU8hRub8h5GhkqKosYJ5+fAA
1o/6E+/COTeAhRweYMdH6A/ogbG4BrVhLdvoMNA6xlNNOgmSVLqlzOV7zroR
6jmopF+gaH6GkcwTwvXSLbheC307Ra1pQXpzdOrgs533cAFHyrG6qZwuWqHm
iSbTyxCYevY2Nd22lA73cUW1MVcyxS5r/2Eby3XOWMm4I81TYePsBpcGz0PN
pHdGmJ8kA3e3RtuVMCkOBQmZ6qLkaxJ9FciJTrV5BY841RACyVLKDarru6XM
mN0aSgja1MB5mU0A6H+Jr+MEtKY1AsaSQP7RPQXT2wy5JYg7UxOi4T49QTLV
Ap9wCvjBLbYWG0PaAslx5zz6X2ZT2JXeyu2UKU2/U9KvP/jHoskGrR0kXqkN
l+LcY9qKAoOEYcjTUhOCwoDNggnw9GYODDbJndZm0CqLtwjcCEJLzAcqV0va
crcTm3SRWmhI5K3VfuH9GM6lYLjwYUxJFm5Q6cK7DmaiatLFO7PtoU/YKufk
bZDeOjJlJTQ8UkCZ59ygLPzvcKherJ/MpNlP0nwyJ+w+2qux6ZUeK4vQMJiU
rW1uzKm3A+Ae54SheqkBdQ9COfrZD+JoNqP6vVg2o10qU7cpf7MLO/Ip24ZS
X6nHJ/9eKAwhtf2FfEHRRknNBFBxcPTpcvS/R9vTTuxZUZuDUpJTqPpQRhY0
0o6Q/Rp/eUmqK8TNqx80okl7oVToIkDtU5UcwimUhqiIkslRDs9XtuDIvW/t
I+78hyCq+dxus5u82FctUJSQ9T82Ulezz7ODX3Xl/bMyQ68YUD/CKofpTb8E
E+3qcXG03JvRspWImOk7f2rq1G8nj+Opi4hqBYTlrRhSHQPYXXgqgtpn62WR
XkSqwNjdD388IDxZgBJiWXbhYOxv2Dnf+1jAcvdYKtWN95Fk4GAl15xXa0ZO
2me4hqTBdwDy9DiLFvM390lqswQJTOF5fQmxJ/D5f/05g2RovVzg39Gog/v7
5aGNTDhOjUyorzahw50RgYIl8FH5QO4Gfbc9IvoRg9l95zKuKX+9HgM3lPrJ
WbS2Qbe+qph6l6cFPsfWeCOTsfsiIR01xHevAC+75kOKQduTaeJefE5E0vtD
1jy81fPfll0XX/wq/jMyNnoa+vwuqE9yKTF01DPTacF1+0Lg6SU3wonvnXy6
d4oPhVaz8bkrDDPr38G5EapssCGmYlBDRaeigFwoWIBNsxqRS+8Hm/Pio3PV
cwTVJTmAwVxlEmXdlnX8W1ibAuQP79On1n0Ih2laEkev1s4VdsdZ+FT5ZYhr
p7fSHL2XIO6edeUApGjZ87IgOZUepVfTOQbwRom74cLcsl/svcXx48wEJsi9
zpzgPRA9+hwmrpNpFHmWknXJE2ZKt1zWEpLt6hdUdRefXPnPG55hRuWVza0e
0Ua6MtQvX1dqmfH6nL4qyD3V/Coz4YTmU4BT3ppjo1nL48HuUOjWtefZYpcd
dhNq8T6OkIlizjeLPiNE5JSNv1iDAOaElV08e8CVuFUSeASkMiwUSpXeYSZ1
SwO7NIGPhIhH6vOXTSBsJekDX0PmUQ4dhFwye/pYpNncd811BiSGLe24QxMY
pYvx7eMx3SrhfQw5HDGD2wsZoncanAGRU0S0bBAC2UifTcsrY2/zRncnvo1T
Sg1uPydRs/I98aTGKkQHeGcRQPD/Qv8qSdB7/mpBEe86BFlvkZQYlOtOf94v
EeS+SJ0HZwvDwPQ5Et2fS+HsTvUNOCY4Car9W9i/3xWwuXT3GUerHKW2SI0j
aNgIO1HWj/oqkZgW6Dct+Ka+9UvHPzgCjVEb1zl9ORVJh5dnK7P0DR/JDXqA
dpEPgxoaU1rg6/BMS9Uaap4TeYpZeFbVniMFtNwqHWHHoJwuOFF9cIkhbUhU
361756TDnRIUUokl3Nn25pEQVtqmVUZb1frogEB4PsXksAwJIrniPf6F27jW
gcQStp1iuI5lpIhxbVdSZOpZLXy0omFnT+YI2czRRMKFhXtuTcI3dcdthfZS
7dv/nKh6A46P8QVTaOWDC5bchKGYCPQt+fJH8RchLjJCalhWiDUe561kcC0m
pczjho1htPOC8xrwsNdTRXc8hYsnqqzGP1mFW/9vIlgemcIeRRhCGZ/N0uLr
/SA1Ag0lb88ECU1wzF6DuMXo6YSXYtcfLr6wIsMbQy0xjDDCp/OffNjCwj9m
DeNd43jP5rgG/W87nnmd/m5Ndtq7kixjoYw2R5JmrNCUt4Ap09dRxB043xQ4
EeLfYQo/bBfVz92Xozj+P59+bRCFy+6mZ98bLbTToTT+TljrpIsculsL61sx
BYfoiWd5vfYnH82tSSl66i5wsvliXYx1MXWuSADtkNzAi7TtrA7gnpHqcEsj
WL1by02dOnNTHOSd9O5fMYeor+4zZx57z1VtRg7S1dJ2xiE9dEIigsZpmk5m
pHs80HNykYJpJmaDJR2BJ26L8SP4AMDJ2wRfl7mTYsNli0fdHABuhHd7A+k1
CF2p0D/hGeFrkqq8UswYjQ8h46nR7kxAXKGL5YTv4GwEJdPLgVwZmR2nCLaY
aCLSzX/loqIqVpupQbN6KpiTINiFvHmffMIpHKy9cnUmF4cMWfLxMRxZy0Cd
HFhruQ48b6FhyjxLe7gjoflg/lltFWTQgb46zi7303HEjPS1+lZhgaJN2Y67
n7+7Y1zcBIB+bAh9YTNlWR8ICO/ImpvUPkb9WEygjbna7QUKm12vFsE22Rl3
EfDxFKjkTtn04XXx3Zd+wWR9ZW0hY/HIkTA4qz3QSHJ4Q0s5uCYVG7F8cXPU
qrf/1XsHJC9075/YAsCGlW+MkSYqIa0RIk7ZmUMXRzyguaiI9bfCSYV1OBep
xXDOtta7IgfiKvDsJdtNF+gQNnfbcJ43jFSbKwSS3XwnW2uGqD1chkj/rfok
9aILbBVA64AA5fWKmZ/HINTkForKtjFruaTjiZ7NlHJwuyCnQpxw9nX2r61D
/XYKpPOWkFSCvnsE43PxP5N6deKnovo1i523IAZh121SXF9hSnKtHVo3K7YL
nitTNvVuVkEuzw5ebbb37gsM8G4JkGuT93jjdZhrl4E21dGvFwKCYBbtgUay
ii8T7DHOW1knmVoWsARLNL1F7o6VtPRGKqk5fYtrjLWaqRLQd42eklkeJgAa
UnNtJY/yvP+dBtPTW3enewI6DVnyreZ7EX2kujDIk1BMDJRMwIbcJX2Xy8pf
W3yusd2UQni9ncbDTU2vI/I2jVimCVXu/HtTAoXRsNnFqN8Sfqf9feCfa3d2
wcMJdVdXgjC2JFyfDXb2rCuZeFZzAIuapr8A4hx4ybDBUY5ayyLDtUIN/cBC
/hgrxvxEfaOZFjfwB/jKLACQVrOiE6UVhJK8uIv60JdiM6Y6hrvxQkw8ct5w
O5FJ8R6VQjH8H/C70OYtytXBIyZDyXcHABK0tnNuIQ8Ccw0JsALY8nl/8+WW
hbeoYVRRb06bO8jOj21n86Xvu6wqPEAdEabEl3WAQsvMN+3GhbvHE0FASb7N
/4j6l08+KO7DjLg+I5oWocOkebmQlxP5qtZyNrchS8LWs9S+S/DMgiu+EFPg
wMKxUzTMS6ceQAGJ1POVJq6WlOCYVxRC/pF3JbtZsdHix3dYHRuPvrKlxl4k
aSdaYAHN7UCS/uFbyLZjMDkPQiSop7XiAY2eME6hv28x6Iz0KaBaXRqmwZy3
me2qL97QZtZHTGw+3ZiZKJkDlMpgCzQWSCHRzKmDO2X5OxUuBWXeYjW/fOMY
DRqMmjLTNOtwIHsrraCnpas4udHzL4pjFuotf5zUf/JDV2vDQGjmDPaRVMUY
xGjP1YAK6yfqjhADHj8QuGaM3uxfywY/Qz+USH6o5i7CzE+k7b+dqfMSTWyd
ghUk5Ts6qzrB/xUwH1Sa9eR48jejm/SNM4bd80F68Sgm8zGsD6rbyQyb+070
FaLvfhDuKoXy7ekqYtyq/GJA3nnWbzlifDKVzgFe270Y+88MaggvBkERCO8+
6F5jvrEctktp8BHxcmhtR+tx9C6gai+Qbu3pmu60+U8+WSmP+Qj32R18NYLO
RqUTbTeBNq8t9XDh9TUcxBDGwDX8UixX8juCGK5a1LAiVof+OIelA8SPmoMI
kQFE4P90O2YQFZDhMAkWtDQqdemY4DmnevXwSnQDWkeWMeuJUPWryeDC6LyF
8tvXOw4FzHsijmS7j8blTdY+D3gUf5kLqxQSVilFedlmbkCXxhk3gYqMtpyr
OQV1fXag6RCsN+Ht+V0fFOYurPFgYDnyXepV4XnLvCtZtUlngdthpU/YXKAl
9hmDGM5As+6NgPhyJE3AltQ0Pl50Kl077211kuLvQWCLo5ZH6wWB8FNn1Mio
lqFbwIrndAEQBvI8NjciHaiVokNUmr4nrHYt0DcwA/D6TUFhWxYvC3IvGyEF
QlE4s8hMY0kkZKxQiJX47a5lofurjivSk+AdSrVNOdR/bbQ7pX5s0cMqKDut
0SXOtSQR747M87p52wakoKSUwUx/701JMvD5fHxXUK2uK7/yTrmnlECygMYB
GuWyLnDoc2Hus+Zv85mG1gsjw4rjB5BPiQEbEVyxmFXdt9fIv9QyidiPCPc1
Jcf7iK7W8h+YDxvLkL/ErIWf6fd2DeQH9Wm7RgR8/renT42g5AHX1eTz8L8Q
bAkf/Ur8ZnlPDdMQoPjZNM+LTvV2seGJVFicmE0nKHWmC6pH6aIdMBpKrsDS
b23vRNxf7qgjz5Z1ffWctKDcxCyuu69XQtGKdSZnQ/UXQNwVye0Sxx2Aneyl
4p2uD0C7f4J5yo4gfJoCpZvtEldermNKjMMuWq/ceV/uToQ7AkRb9dtdDPBV
vdx33CyrIq0p0lXzvy4XBX9cbGZZhKkpAW7vn60Eo0pxuwBn4pb1bNh3rR6H
9Vhh1GSO9PlgYw2kvzAAFOJTWIF4qWfKG8tvX75fbSjZq95KfbXhj1Ybk1tV
8+QrvAd5TEJC2jYd9eRJeSRnRcuownw6hKsjsqRvdmt54mBMFtxT0DlxOE2u
BLqJPLol2MUNPHwMaqRmMPBYfrhMmBL+0OOpUSFFpgKwvvMyhF2mfcpBwpY/
QSum6lQMeM1oHdOUfXzvksXNVdjRthjz1WmcGR+pMlQO81VB6BTTf7NtoNRq
DxYd8Got04gz/drCbyJ/NGBZh7v7ukKfdPlzMcZ5DjtTdAiv8jZnqQqdQuhX
ULvQVgRvX9YUEetH8LG47rrrM/7TKY37qjP806DOi89Rt7Rf1tydHFFx7w5i
y87R/DL4nkkLN0YJ9Rkj94V0vFEFeVvTTnXYcCTK41S2E42Q60RFTakdvZjO
t4Vo5XU8PrjSPzHyFvjDDFrTOG4P21UODotyxO2ony5pn4wODhIE54NDBWhC
U2w5S1L5rCWh2LCa8WI5L2iu824PXNcxvno90FHnx6o/Uvx+i1fLQgvRSsHE
yBXtPCDZH3zBtJZcR7Zmp9KyTip8iyNDzbXBK05dpaGM5KFo+2T0uIes4o6B
nIdK9UlYLm9AGIA4AOkfIFiORfhW9YEhsn81tFmj6PQkcDdOGM36iizIFpJU
glbVsU2BOWrldguBxFASHexDTv5xpf/CpJHFJsngvckTsQr7hNHwaAvY23+2
w1U2sX6kV3RS1KFXmmk8iV24Xr+1bycjW1nRp8dbap0rKwqh6br0c42LRjPz
ku7KSOWj+vEbj97Rvy5QjR2EPG7ojHtcqi7Wz/miu2J4QLWFqYH9tP9ef86E
8mYaHN+P/V23xB59iBpB+kL2cRtfTbbX5QApecGAcFa/SE8Ub3km4eGWNlil
mQ7TMjiRaU8Hx8sXWP1s3PPIK/xPsOodffANGr6pTB4anWTn0sqHjcf5M7mx
xFeFenPTYWKeLGrsIcueZ20NzGmmlOg/RgSQL9xLhly92+K+67zImGritsEM
Bgj81EU+5sg5QN4VO24b3YyhxHZwCmtPJ/lzBrhVMfs155zsdjnfAKUbyg19
T0i3CBVTtYOxRl5yyRbnP6vHQTd4r12iZbdaBA21eU+DmpJtuAOxT4Iu52KO
hvrcCT4uetETnTseIi5qEHdrv5TNO/Vz47xxo66ccB0pF3h2w1PgoJZvIfnP
kOdCXEclunboDwB8CwZgbQ5moCdIeWfA4TdUQV5nrcDfJVXX3XycsS0JGKBK
INQL/+S7YAuMePCXChSVVESyQbaXa/e3nYR/jewNOjn2MCFJV0hvF9uwbMAC
6pFHCWVY3jgCKqU0Bk016dqDWnO8hODmAxxPnrxhdbNZQlZtUW6WFNe9C6VL
v8dJNY8Y3HMGoxRZabL2HqzqhRAY/ykn6/dpUXP8ogMCNUGkjK9zYsrUUwzC
Wu9NGr8JiJvPOJzXw1q4fJABKwjSqgdweHY8unD2IbExT3t25sJ3efMApVJB
P4AgEmpAHOqRFqytC2a4Z5OFXWYC8oD0X3G+lGXMIYCEcN9JESTNZwTxJkc7
f93YTQFQ63AnWnxWkwqoqqqBdfWRRczvQ8B8duka/NfSw5sGtcLvefNnR+NJ
DH6LekoYQ8I16eqIboIn8VneDnzmFH2JIUwSkMIIUumooaRD3MnsiCoV/dx3
rlknXJ7p+iQWgIAW8XJmAYGTSuLfgS7dPURGWVAxG0MqIJZlYENubiO3zxS+
Q6mGc79HVu8l8p0aLFrEX3cJnXB3vVGLAbLZ8iTyoy1uYYsUFm6QFN8sdqyO
JUyp+oz5Li1JzZPW1fs2TxJdK7FRE2lLlN1Wmg0w/5naNo8cC7ErQjTT/BeQ
t2yVwztKWbf0SVSmLA0hqAd4fTPa+H18YoqyTSpVv3GXL1WTpqOtj7QTcPpm
sfV7TZJ3nE2Tiq1A5fyzLVv99FbwvRXtQICPLK7mwGz0jLdnXPJRH5Efhudw
1MNsudiI1bcaZx4fLLtBCEM0bSqljOLCXB4TTlNdFHvTC35uDuMsZxXrFptJ
RRoiFNiN19DofEPcTG9HfpP9OIeGaQ53w/+dRpiBM9BKOMViZJzK4zdzNsFX
9N7hJ5Uej+cBaCoWFFjK1MDHMuM8BrdNVmfLqAVjnkLbYDm4iXAWIIaykK0A
uWUdN6z7xn2RknegmOfvo+93AEX2ox/WLw/HP0/TCbqPHacDSU7WhMQPUGht
qCMa8ILgCpkvXmxR6/OjqQ8Ri8d3STEJNZPjRHSGpb82+JxrN9DBxEFACu5w
+OT5Ds/Xi5uJdosweMqLoSTvpgAcroYvAO400lfik5Zcc5nROkvg4HqlynFZ
BuYCeii8hlFnoZJgVfWf+wFDugUTGp1u87DOht9SH7f/E5TxdT5EXMVCm4vd
/mqtSyJOFp/bdCERLBzDvFPq8mhtUbdAgr3q1PCXbhK5yHGvO/JsDakWPv7/
LSEPgyS9KmqM6D58tgKbwEKiFDWJ3HXpj+wCQVZDdpTetxX2so1CA3yYZvT9
D1xVk+0zJruSeRMCtloSjnAYzWD/vVU4FPwrdM7gtC0i3JYdkNtmEqyj+guB
am8OZ3OW2r7GkTqHygS3sp7wzaVoAD+9gwGis7/jQcmTp8SzVlbOmlzqXZD4
hSWkD2GLULl/kcEnIvwy+zhYCDzU46MiVDN9RiIEh4xbDiUR+aNkkTca3qWU
GL5aDpa25gCmsIH/YxKFB6jbkuzTK5IK7V0CtuqzFkDy+PwEiVPvFj/RRSxR
SiSaF5ShdQSJ1fLis4bki1gAGTvKvISlTSnDawSsp/PYxyfzMT4Mmywo/sXA
1DyCI0VFWqSBlzeH5q1jLQe+gZiLbm70vPLBAKLx7d4B6wGaiV2fVjvxU26W
96v8dobKIJM28EgPo6bt7AHXM7fLStUE9Y6FlJav2dorSeX+nTlvTMKX/n2Y
CA7jK/T8O+cP93ZyvR4WhmQo6zbATa26XSMSwx6Aqyh66yP4CL926K/OEZUB
LPpJ0kB3Y2F4W4D0mVBQXQwS9lhvojwnRiw3d7ujCgGGQTCbC0Za73ILAznc
LzICwJOKeJZG4S64yIx6TIvAwS2aZN0Xr+7eupgbA499kZpO5clIb/z3KFlv
Lj7Wxr5wj2BM8NgIeIUTYotU9xtjMF5JSfJ+3lOmqmHQfR0LIce3LDA6yC5O
nB6YxusMHU+3dZ6Pq5IshtcjqKh6hazwtOpVbaffKjIknHhEjd47v8JfXPrT
iNG5phuWFDMwe6W1gr4+UU730/LEkQbWaKboVRMjhi3J7DsEPZUo5Jf7BYRX
WzBMigjAfTRibtYeo7X8X2lmAKhAtUE3VlZBkIzjz9xB6vgrphHOdMtFTHXF
/Nanlby9FedgoxNu60unYLsFEvR5IoUpe3qIpevGZHk6nIUkGulk39ilVNPY
79XVLzU1KwVvU/SeV7SfX1Uei084V2cm0oBOewFIh9B+dbCArPbbeAsp9KF0
0tpNN5ZRbxfJ+y+z4e+dl6NUD4hjffJ9vteSpYbSsY+stRGta/OAdojDEEFa
XWTPrH+yzfhH6zC0mr+q7qK4e2mZrDUSFAjfqqtSUk9yzLPOdW+KheClSQF0
iwsj+IsuRM2L8ympg++vK3bWOlXqlT5ENJEt/8EKBT7Fp2hcf0UHZ6K8ocYS
mKFbaawy/26f/APCCKkYpWyK5r9f9xZZgOZuNHO2LUML1soMsAiEXGs0A87P
WeTQkNmbNzV0UOwaqKth4HUSNTLZqdMkHRZhhwA2kvVDs3qIMSo81RVctUVu
x5p0t/yR1EjeWNopsgOSwrpXiRiN1RNWtgphlBqC8TFn9uhOuivmgmhcb4mh
NIaciBmBfs9pH0HOl/gSinCDBeHc7+S0u0Uz0ngsG/iRyMMgqOT4bpse+KV3
vgp2u3q5GplKEW2y32cz4HXBwmHe4ipK8eGImi8ne2aaKJpM7Ew4pDYPQxYQ
GO+V74bsCUl0g4kllinAo+pG8GqxhrqbdPt8ra27gU8aFIMSC0ccGfjpOits
LTsHAKjVw7HMbGVTYL+42JV91kzLyZdPg/0FHx9Pb7ZasjSV0qWFSlPGtfen
/ibeut5yNB/DUUqAMGL1Yc2g5or18Tsbj40z7nwQ8mLF+/5nSODcatY1gJ0T
/WFewQ1ijdnRJvL2q78MHQcAtV2keQ04+PuZC3L8wlcPm6ddrHrUMo78o/+8
6XFANPvKFikLRjk+EqHzgiWFBnUMIWKZbYAoc7YsjlE/83Bj9YoMNxvst/ss
t0BQLoC8JtIgODH1zmA2h9iNKjUI9JyR5GAL/wKJtVPpdzIeaidByVvLpNRp
GXsu7ras6m36yQR9CkNDF2/afhfA1oudlYuK0kF3/y0CLOIHI1RDfH9I8ALS
W/pTCeFm8Bmhpjh3GfhlTD/k1raw5+dmGEBy0hENIGzjawdYSXTiDd48WC4U
/R1HzjC4WCFaZBqWx2lUzu75LJQNjiZn6Nj4SPb+9b8YHw/KQKmTfNCXCiWE
Rc/4CV0/NCI4xFowrWOriarpvNS7Gqcztl7QWKZtb7yMlno7xmdduOgleYPa
XewNuCQNcxrLYMvdjr2juZByu0d4rWBunBmT+maiSABh6RQMNePPV3MXpw95
5Eg03GtXf15TlPFG5aUW5oeqUUFFfxaJLAU5U70mlwcnP0QQcnyDmPBqMJcM
4VlRjdDvTDz6hpsGcF9+MwrrGTB6g+p/LNzLMUqgaxZfU8++aPtAImxVVUeS
J6Fcla1WrLtMIvZFYvsUz0IE8wkLw1RQxwAZuV26AlJmUpd2aR9osQO8VDy1
KwtxWFilYIjLNzUGCs+mXoJ0zrQPvH43zoALSMh7OfW6esUU6FRmL8gxPyT7
rFG9qQL0kDLVq5coTx311rF0V7dxTrvHc/Hrao4iYg/grPo0Pbq4UlW9J/5e
j66GA35+93A/GbS1IV5J4ehoWshb2srMNTptxRR6jmwOtpximLCSNzhS+7T7
OFw+Pl99OVZ5sBBTsZKQST0vmUPROUYmgm+wwT63zeVy0l6wJlp15H0IKRba
59kjF6UgUvw6n9LOQF3Ex5CqUFqzZiMizyhc6oDvoIVKdCnLSpgsmWr7OqUz
5tvdLs+3++MpQ5x/f3RvzT7h3jlrAMdvvTLcKuLYkWrS+SNMF3VLJD0FkKLA
1cgoPgufgOVUBjnIhPYya6+Tz6Lf4YJYzXzO0PlPQUAbXYmKTxhDxNedgY7V
aJTd8dpHXcc7a8KuGZ/q0L2X78A3qEHc+vUpdDIKEmx0ug0P/Z2fkGC2eREH
RVMkhZZm4+e3oEs5es8cZRHwSHMGpq100N42KqVpKzI1hULaqgi5je5+JNC/
AdM0YgQFRWxWm52p4HkVfMpRveEBF45B0gtR3kNJlHMfBDc3QXXsCK39mu4S
mmFnFxyF5ctXauMorIxu2pm8L8fIT7M9lok4HLzca+s5otNDBesMIVzqPlt6
SfwCgZ4YiQLvQmR/VnS4vQj3UBKfQC+A5a1zF/EnxPZqWp7fe0xSlMxmrJIK
tXsCgwvIc0PHFKZzHK9MKAMxmo570y1n2Ng5lyydpHlYfHSyb6ou+BAfOsh/
RB4sRvdVA+hq+Qw56SMb5MJcFYUcZL/ydN/AxWqMKZh5vHq+eD1jPz0wPoSf
fEd7prTEZBsdeN2fUxfh7t/HPKbWPzbl7r02aMM9HLQ0aHzXeSsUEZelVRw/
OzxwwNnGbHqipUXRCTq93+hpVEWb0ocLsQNQhqAuKXlSUgWXrgQh3/IPMvUT
NdBVvjZiT6FpasKdnQdnSuZeR853murR3iSQVGkt8LmUZvqKLVG2xMWTHUnY
gIH7PD4Ge1JmP2W2ushe7LGmeP+UDYi4a185h9Dh6jX0/qlvVz5FY77q9mOO
D1Fo7Ul8qWylI+PT1ptyjMwbI6nKpP8BboeLmjPwYQrKjfd5rntBc0NpUSkl
EKDntVpNsoOumBGJaR3XdIP6SkkKlybNt2El5RDbNuochi3zfiMGVREAvA7j
+3NjgzcrCsp2EWzaTEoP669UxfCw6UrYDttdQ3jpmxNYBnOh18YScmLGQ/1z
5pB0bIoLbujP9i4MNW1AsVTsj89I8ldqRGKVOOy8hAEmfX0TbedOiGQNoxe+
wYV+pAYiOLPliKung25mnKWsB0dwxN0w+DUhKU555be/4sbJqWRKWl0A78Nx
J47iiJdrTB68W7tRPLstPSrrc2mZrMwo1y3MjzZzDNfsbDNJIJIOngerz3o9
uGwT8C9mgMkqv1cirEi7UDqzPT7NKxP91MlkUCRY6nNpIDlxkTtIa+Ze8UUO
L9hvY7Uhulgx3C4lc/ncOxwgAev5+1Nh/tTISIL645LLInWrM9NEQV2sQsCG
zw1nCz7YUAQdgOFLlCr0F7Ry206we3GWeItUIpcm1EnfFmAZSvswPqk/wNAn
0AuDeyv7ZzIbLT4C2rNiIc0ffGaFYUIWPVmkShMc2Ej9/eFear13Rb4xfduD
QP27pR6o0gr2L82NeEl/UCIhXibITlrHACKTTvhYW+k1fHXcDkXb1LX2mdi4
EAGabSlcTzQ+I8icV8qdx8r35kdSo2mq/t7h0PfEVDq3r3DQTjnNOIuiwqA5
DsoWHnAME7+D7jTvJKGdKy7B59TmdX5EwFGIU8Z5Slw1p7EMW0EeoEWFueoP
fLgA7g0rGd/23ltE8Og/IMWxy3oAjM0A0bn7GQb8U089qqBaTFcVSYq2TDXp
1oAeXzcWXl8COnot11AxSv5ENpRJVoIRIoJm4pVDAPFDzPE66ppg97+Oon8j
mE9BJP2RWtsmUNuiKPBY3xNBjV6c1ggoUUNo12kORIZ1wRtUDADSWZxxLOrs
QGkewxNVGOwguzFJLj2P4kebsHFTv7LabBe8YnIoIzAoR40eOrMhZEvEdt/0
BkTCiWYeJYZCzMyiCyZfcHIzyKK7fPhAjhUphVpcegFj4A0h7K77YajKdlWZ
c7yDtFHVrm8gEExyRN0CDeMxN9IsrYs8l5SaRLRsL7dByMUE0ArYcznn221i
Ln5LHtiYHKbnDiUknSJUlu/JlXepB4B9Mj/niFot5HK8PR0H5MVzxKcfu5k+
ITZjnzpV6LNxK+CL4xNyPJcr2uOGm1zsbI34YuLILth5eNzbaON/hRbDdojK
xzJCBivh36V9u04Hk059JiiZ39mv8bt1KM6aDWZHvdrFDeO7fbLI1SOkpAMg
n4Tfut6xh6tWXR61Ihp+SnniJJtkLvmOGs0aXkUFa20LXZFppR1oGiBFf8LR
S02ihnMw5YW3NDIYeCzOI7klHIp/Qp53ocYbiSt7HZkYrJLz8ER1A69p9xMN
bjRjHLeT+mqfzxCVEg3zxU9qYcsFGDT750i0gN+Yv0oHGJ+DCYCfjUqrXn7M
tQE5lhQe7ZIKrp516HGhYcfrSa0acZFp7/tQdaYewfxmVc+e2SVuUGVRcPZD
AxXJv8WdJ6O5D46k1wwRlakYhvMSrjcFipQUEVJvtx9oJsCpDr/4HTu8Q6Zh
9RmORj+Y9DSfFsm+5/cEBRa5Ca+Jj+ChH1AJBNKLjS5GwQeIlT3G5AjZNJvx
d0q4AzjvPtqq4Ly5I6ozEUpowEvADpZLmbG8dUyeZpqD7Fgd1ORLW1z/0SW3
E6f6arc+SClCy9eXylNBTyuGRjUkDBhVTbOZ36FRGVWazey7R+XXqJsx+40Z
LsUM01Lg8QGi7E4hd27/4kN4JOirDiZJehstyflvcPzoCsplPaG76ae5yoAb
rK5lxDLn17CMpix8VA7pnXDww4RtloFDh5emxtAUvzLfWdpbrrxHzOhFzxS6
qZCkzEZ89Gx1Qgr4gykzb1BV8NwUywGdw/2LzQ8oQgVpKKz37T6bB9CLbsdU
aTVOePmu5s7J5yq4WKHlN491984Dt4bVE+vP0xW4vh5cT34GiOeyewZcXxt7
gd43TR8q+6dxHIm5U+9MJZShABKXQwX+1BrgqgV5UsQ7KZF4XElKiUv9uTAI
EQf2Ubl3Mt8hE1ef0NT/OmuH77Opf7CfCbtY2or7s5yWoAOYIo8nIyO8Hqgd
BLwvEKK+drCPP60Gq0wWqordaDOx/7XOjQahVf9kBxOhEa8pKR9PsumVqbu9
3NY5vocoIWNqgKGmiu7LCUzdl8MBvX1yZ3aeovjPFICG5iPK8om1nT6ToFea
LCrC3Jx0CeglSmwqanJz6iDd3JQqWHFFbi7Hht6Mgui+bhIad4Pf+VUBSxiZ
efOgUM/JCLSzQGW1aRihiYBvdjt1xPmNRVbAeOCTThNmNsil+WTTYiJrPup3
jlsMK4GR1c6nUSmH+VB/Y7QZIGjIV8giybBzqUnPY2lY99JoMoA3oIqu8sXW
NxepRjh2XR3XKKgfcrYKpRsGq9pOCOqxzICVk6sQdoigWeJgCQfD2hCWJZFw
mfEN6HwU+lSVhpKWM4yopJeWEvIdb/vuQqdQcPxGkGncqKast/sGuUQVeOsq
aZfZt0wu3jkdJuL6KRrHulKQfl038ijWqVJcWYfBNY7enyIT8kUfhC51SzYd
ach+GysVszAJi7YutlQ/vKPtgGbC7A/hCn4wWA7ksGUjQR6AKlIxoVftbWzX
9O+kGx6QpM6P8fUsdAeB8fIf7KcrYgdTsqOf1p1DNUfw99ogV/qFHidT/28E
e1D9dFh9x95XI9j9nQJrKDv0BrzlmxiZwa+ld4dEvO/DkuwnSGM82t5/omhR
mqWc3BAjYdlqslj3o/zkY7XA8aGFFh3gB8rGssEQSouuC+6N5m8bZ3gjy5hC
a6IoXj18OaI+VOa09HETXOLjGENC6EYgx5zbcQk0mLALxSREkWYpNBg8Dtb1
jVg5taE2Gh97Y8flpIhsY2vNk4BFBQWdvAhUnDNEXtnu6YVy7WF3qYoUvyDa
VPsegjssWCkGkJLvQqiMwLx6dmSPCSo3ts1/ed8CEJDBBL6UXwMYIGkq2obe
ahEz9X1jOx0ZIJis6lxeC/kAH1MaJBcX5qf5L8NMJZPpQdTCjpKip+DYJVvt
kY4P0lB4H7lGFdQyY6KEaB7Z4nOIh56ZNDhKwHYGPXjMdk1dB8ne0rf9i0yY
6sX9ndNq9nAGKe88KcEOv74Shhb8v72xNdyGEXnM4QYL/PDkZX6Ik+6CVDPr
muFsc77KqXnHpM85LqMacY0YLdxyaUNwpaI04MJTjEO4Uew8HoxEHF3LKU0m
hgf8aY4yjxcdbExdBCS315z4fQfjJWmuCRKPBWv/9qXOaEvFLymqfQz2QKfw
jp+1ryN4JnoVEtizYGnYB4/vicDanTNT7TC4Gc+aJT5v/vhQw26JaQpJZOcy
81YRcjxPegshEce6yR8bqQt/PebxFNO+9c+KBrkQkFQpJBvxtT5SimlKF5Nc
fca31IzkN63vkM+o12X+JT3pCXgKKybkmHtmcJDBlYNYqu0mZfYh2im/BURk
RIYEoo0Tb83rsFqCtNwMmpDTnMhUfVaub68GIdxMg3dVM1O1DQBSvej5vTfE
6ocl3NLeqHo2tgPFKI7qr0qMn64Yy0tJJHjo4MH+oeEa+rM8b1aRIDKef0h3
+XtXael5vEM6gM0OWJVItUI8rHzemY1WtkVC1SnVc50nzjnyZv2zKEYEV/Ln
WYd+ZjP0A3ePqn53DDKycfAucRhVTnUpYwOnJMkvtl0bJdsUJkf35VL0X7rl
YtNbtzYBnsyuLtXWKA6F64S789c613lvrCee/B9dB6XyarkSP3lo9UuLlvfl
nIaHgI1XabV6l/a3nDBC1d2isFLx12FwhmZYAdpcw06VeEANid0QiiPgC4ED
p14+3zUyFUPZIpIyg4V+UB72cj/KhSoW7coAEX0kHqtCrhhYaqCkwxOXTeC4
B5uQsqTTllF/LULofC0Lz1youtMvhkwEsQjH9GF4ZlXKzdWj4r9eusbG6J7W
0pUyY/SJbTdZj5dyS4AmxDDYMrcncD0z6V2HSJHRnVJAaccaGJmG3hDt+KwI
rsQ4fJCmyJoN7P3Bm2XCcN2kuw7VIUz9YHz7dReWVISsCR301CkrfsUrArzl
ktPIAY1o+Jlkt8ToKWdIFEU9iSkUDU4CE6PasCXjgQ5AEE15h7aYcPKI0OnO
+X4ROpVFvaJqFBeWwnWtKPV/MNxZW13WVgzdcNrudIS42Y7ZxdqcJ6F5kb7y
Jl1ljtpGG+2PCR0jBaXpaLfS0F8cW1XUn+wgezENeJ5UAqXEIKbJOs/ifubY
A2nN6iqfU6G4d+iJ6A9j6HQ+jR24E9qi8W9YVJfBOiLa0p/O7hxGll1BATFg
3iHbmRRNWFOMyw0fQrdW/z7vkAtM+QJBtc0hJeGRUfhalpohM/cEOfcVPftD
2/jRATQElkGDm1mgineIFWkJcwB0bJbrnqClnS67A/u0ZVFYcFTxDmFaZunG
QmeQn5jHCYFD0lpVHz9YA40X+xOvwL472dUAl7lVEyqs5DDbWeb40duKGldA
fAfpRpkiipOOhm/FjeN2sNQQkmBYGjGE1bkr24kjhMQ1Cpb89w9kaWS8UAeY
2pyR/QJ7JoGZqw/xuHDGv2vWR2pi9HRl0bldPgVB+r7Q+FKEOKdi99OIruSE
AZkSIgeAUFDIDHCyr3/qVSfR6Vj4vNogees981x9dobA+/zurwaDBr6OHzmy
0gr558b3PMwxpF+bbKNG/Fq/HxY2Ry6/LFT+c6awf23pYADxk4sR5UH7eaGN
1WHI3LJLEIeql9DucwtgFrJ3fIhI1zmO4A/27MrmhnStkZUvO8GDylnDzgdb
hsg5cDbMrC2JZSnIfX3CpvsxHnkTh3EvB67EagY8HQK7/q4dFDtirD6hdB9b
zwX1nIwAf/tnl4A0p/dAKf7S3y/GKvcLK3BFVdTpG/GBPCUB3Vfg4YOxLfsI
q53VpK0z4/F6iyo3lH2q6qz4zVudsVSoerRgH22ZeMv+hcI2rMHQoj/RV4zi
JmH+ng9Zzyq0fqTwVPDN37dCpwZ/yuSZRy/13q2rVYQdM3l9p813XR8y7OiI
Wk6wbC5QnP0Y65SK5kPbmCsPRacNJIokXqwTrm+B7SUsRBLGji/5hTiCiKCG
0CAal+72MHkknVf3S+1GawPZNTwTf94bvAMOOKeK0so4OejsfzbFpOhxh/jv
ThvzkgqJd7j/trSbZY4+VIYT4tkeKBCgXetx8ZD+Bjyto8QlLojX2n1GHPSz
ZBka7ERdi2GqME1gSCtuw/Pd173DH14o0Y7wusqzrWkkaYOxAJoz08iWz/LR
xoFMj4ExiRUhFadMF//BuhALqSW0tg2TgGKulDgC2qK6LYTfF+MoB+VBgJ5K
7DB0+bWcvb/RzrMZ5WezbnyBcw4hEuAhazLrVF31K+9o1F4ElnauFA94pmwA
pN9Iuoes8BLGqB38y8F3b7SlFAeKW7qb1hE4DfwPafuhtAj6tYd9cqpb/gEh
XI/M4WoIvqYpM2J4zse6N0KXJ8Zg+HCT33NHApBhVZvkqi6KyMOlF2vsfKVr
SHX61aZkNB92j+ajYHXesRkRNnhvO+arzZlsc/qjm2xPJtgPynB2cFkpPw/I
0BKy/yYjIMjkGRsICzbSmkqUYEcfC0kKXAmc+LS8vm1ilawafmm/m0cdN5R0
ReaiuPMjZ1OFE8eM8h4l0trShi9DldZoXBe8+p6OXfauF9KHHu5gYkWFl4KU
HYp6mVl6rPPEoj/lL0X9L5lR0dJ3sCEaY9VwQChqjlQ47gY2u3cWTMo9NAwg
s/rd7n8FhBPmUEBHV7egmdkIgUsEZo7huRO/ZiPcXy69LJurwWgxqOCDwYFZ
y7kqCPAZ8xUtfFuFNNgHceXFWQn81L22Sh0KAmEkmi/2WWPgQjhN9DXVBX4r
q5kOdz4yNPMlkbj81IaDqsDXD9Mqk1UMIa531QP3PSwI9cQOrVmATyIeFaf1
hU3vyOa5ifkYQWQpRnmHcCDwSduOmnztTXFELfxnYA340y20gJBHH/eh8KUp
K5gbauX6lgWgoMe+pZbbNj3/JoK3WtZU+pTW2X1aZ4AAxRgsdHu/w1jupH4E
Y6X9YeK9+U7Q4Ui6EjPp8Aifmzk5wrOVh0gJLRhJ27Tbt7cjHOf6g3KAj1c9
4ZfMC0JdCAel5yF280Ge4CY6P1j+WyoXgffABDULqkIN5XrUMDWP1DGd4nvA
Pn6bqWugyAmvnytpD29kf4Ig/oFI0jE1jGpDaRd040sylR3uaZ7zaCkPToZs
eZF/4hm5p35nLCDpGT5RpeO5ZvIDs4NSoP56jHUZTcnj1yUPfv6hKQfLspc5
5zJdXrMtvbbwhZ3JjGpbgqjvCrwx6m5TeH/aLlfydguk3b9L2DcxMRNl8OL3
nNuyW50IuuwhOn0CnQOOFsc2e0Mqv5wrQvxS3aqjsWSKCzRUT7vRPJPYLPLn
Jxqb2QplFbgl7QHn7QSnFGwqay8NYASYpc/uoHF7YW/4EqbKwNaNbNNXa/Y3
/ZmQXgOCdsz7WtkizRguQc7cHDV734ee6+SsLFiJ97dab4nQyOEokDQHzIKW
oK8wPISMunqns4MDR3sXIJnG5cO8nZwoN+YWsXXLgfYx/uj0aw2unv6eraZl
bBa7iOm9JgApY/Mu6ZSi6gFD7iyD2L+laH+YwsyR6E7XdUwSmbGgLJkHbZ98
1+6OXKRJH8NgxIwphQSAkEPi8wudzqDBUTzosZTJRpiLHQUfZ6MZMmZlMCoy
K6E2G0zLh2A6/m1NjmU4Rob6bRDAKv6f2dY/naDK1kvtjDrdy5ZT0+qRCRZw
fyFxnko5fmYrsNXj5xLMSKXGYYxDelkfoUGptdxckKnEPMVDk5ScWu1HGJJa
6NrEVMHcM0MFcs2ZCkqiQv2pKMblr0U9yhCofaEvi/YEa4YAaMwo1LHzpQyM
zZanvW0X0lUTITPgb3rBGzRzS/v8w22X5CIXYDIXuxTEcfpkCE7wDdEqEDwL
qiky2mXCBz0yKIC+Z3FMNMMUcsZCPYS1bX9zRxcoOPwNPp6Ppf7Uja5cXFq1
PI/zpfJiqNOmeHWEPf47nBq7nVZeZTrFAqAXVnZJCGsbvgwZdqDUWydB/e8A
IfASlEs4G4IZOaNbJRmv/+qXKx2v0I0M96s4wO95lqm6GPWQuEv+wsdubJq/
mapkmozbfjAFq5yeKgPysT96/hWfaegIyMP9H+tVygWv1MXNwFLSSXvQhKlQ
quASFG2GlraeB4EZPolkKmaFLVOJay69hnXcIp1IWGsOkmAm6Do7TGCMTEB4
fRxaN/V/TA3OtnxKATxgJKFu7hGAfMia9mVSR2zjSSlVgkkEcN0nHDccwqEH
EPEa+yAQYM4RDgfpGnIXTU3Tk6IbBV53BO2C9vlIO4QwVuteHUfrgfNyXpO4
lm2BeCbyVG4FxU9NKWXC/TwVBCrahsunfMqys1ZFphvksoPI0RwUNasnau5H
ybpOrLpI0z53d0I4dE7dx3ut70AWN1HonJ2CJXFmg9NL6kJ9rPozX6K54hTy
4cPTuVnJhVtu9gNSCBfQHjCumzb+vtEImOFn/27e1CR4aoc7Hr5ALVSFZcnT
pZVU1kuWfAsiTe9FmgkOwTFeKGzMxptk9+2AjfX8bbZHd6LqQ0pFXwF8tW86
JWGDNGk9Gwk/kyvdqFexonv2yViln8r3TjPuLTqYh1opV2gL32Sa0LDXluRJ
CjXF1LspudHFU9OHT/FczN59PlI84yJn8sQ/i66ioXBnCNOJctR0TmlifglR
jtE6AzN/eRNyArXP73bTH1Ngzl5WERLVLz57zmRf6i9wN/E4+Xk0b11i3296
GyBXkGxJMcP+V5IXWl573tzuELceduGo5D3DKGh4qrKp3lL84/GPSzCMf3K4
aW+CwEIAk91ElG4eHyuhuQT236/WtSKEqsYvbLgPAQjiJRJ5koNg7d9XVKv5
IWUuieIj2wpe2r/ekCXQNYODjc+E1VBrXKV9wvVFQMjKfzB3bHWgNDX82QN+
eWZq5hOn3Rreff8mQW0lDoXGoQ+KnOO8bxY+WFWTx0eNLG4k2s4E6Qg5jbxc
7c2d+miZ+XqZog+PXFBOyhZsPWey1YQJ26zkUKLOIoDCBzwsz21QV2lHVaj1
eVBniLOmPVhAC5UC7y5I09NpXtktbTHJCAXnTfNnU6SAKqWE1TH0ZJvebfs5
mJ5upyaJNvoBuvhbbB0OcAwBhYpNl0i1NJJ91idwUOJRCHrJOqhKsVbg9W8l
/oU5/CgomSrfwI1p2xHfLWYkzm6KJa7UlXuXHdnS/+fgNPL47aBGYRvlgW0J
XqvIKNAtNIJzRRx/Nph15Tk28M3R2s25W6CnWFGXginy48ZjGs/cfEeRiBmE
MaCzXLqDk0LUTfgdi1rVWN/U2v//lqwApsMF05uq0YQeQWGlOxtLnOsVpzkn
YAeCGkrhaEjVH4gn0kePjKANJ9BbLBKXY9UPDNUPAiyl5nk8DWpy/ih2STUa
CtlxvMwp/aD+6Y84PIiNsPTiYR29cX6Iig+uuEPi9vToDbaaPPwSCNII9swB
5NJ6A7mr5FPG5CrpCIvOPkfG3kuMQkBJdd40ppR495QABgh/zd8Q5WmY0rZn
sc/Out68sVCsf+NmPESfYCJ7RZ6g5/jYbJfJIq83j3nUo9mhMwJflZBFCHnF
aeCGR9cUCe24lSrEaDK7aPLUejxMxCYl0Ao4CzcolxihzKmx4pJ1+HkY0gkX
3PI8S6Ua4efG2IHDdEX0L2ZyglNCtJYxd9BaTGXB4iVLeI+xdhkuOnBusBKp
v5HrVKFMyYJDofE8GWXj3m8vzKM3LiPvDHiROBA9+IAY/alZu0dChbRX14cB
VcvAPNQNoGRVuuQCB5gFifNYQr4jdpUWE/jv8mGUTohb5T/eR/BacTStvKNZ
wHg8O7CRe8Z47084rcYGM5HNJDTD+QAZujbS/GIF4/MnDOBY76fajtEctQlV
yFzdxO2AmLqLB9tWRHqX4DP9WdMJfmba52H5QAUIlqMBXo+3aBZW/9CG1B5i
F62mRQsbeCO0mtG5asuNBYuYBghFJZvWoVskg3pB1PURZEdQd2ysxPBNiyV2
uGsrDhoK+wzScvu+HnAt8kxRfMXkkzGp5BN264Aq83XAKkcUV7tjWjKk1Vz/
tdKu7UkAWVwZTHV2iqm9uWyRI7R977NDDoIyp42/bvpmHR9fW7kaEFajoHdB
pXJBL4DTvyYgDFT9dpEt/VSSNzPs21qhGJjLHzpIQkNFeMtEoIIx9JMjQG1w
lidLMqtWSFPzv2lqQ2dLxyCGnjn5jAaj8fLqdKadjr2xndAg7nENKJvtbhF1
t0h2sUasqzAulzCn9jSYYMYV+i6iwXswuZK0hCM4ePyvUiEfyCsTq0wWWoKh
1M6PKFk4HAXrPF+JuUiyfbk/BFef3UdqM34vtQRQbg0ZfpJ9X7uOSL0ku+4V
wkndQXY3PQEpsXO/aM9VsGncQoHmxMhmFhzjOaSwEY4j4bhFhSoSzAxg52//
aVAHSnZZCCys5lMFfQuH85zMboSZ22I7Wr5L8RzJWjEqfhCzcsLhJAZJCDzU
IgwrY3ECnMnkJQFe58+WJcJGAhjXPoLbjmUg4Tp1o+P9DJO65jVgOpG3Za+0
l16FgJu5fCugNlYk98Bz+hIXOhRrw6Sag8HsZ83aXbFqXWeG8pymA6zXNdGi
i3PDjoobPnBoJrG/MoEmT/hHK/lryQrb79PV0Bycez54ZCQr45dWhVFB7UUF
SL0ZcRrL5vlTtcw0diLk0NdnNAU7nEkdgW+z6RknFFGp6D7UovVSzZZ9wcLx
xZg+HuJxXEpi6vLEtnmqEVaTFhm+/3mlq5DOZRl1tlcinYsBbAOYsOZ8KxFs
My/imJdd3bO0ok6/5E2kI2y28j35K0VOiur8mX+jKxsUxLEe20Xz3+g2iuig
TSYGu9rlBgw4s5Zm6FUazUmfpzOsooJ7ua329tEkVKpAo9VcriDsYGEpmVUu
QHSMvoex3ZizSRwcSVFvzPJlXbhTL3QfdXJ753qQ2bKSU8Ccv0O9SYNaNcst
3Kd/UlZJkmxbcTah8vHE3K8A1pIoJIPixoRUv53EeE1XiK5yg5NtYLMSYwm/
h6r3/HUFAA2Wd37VXGQoWbnxtk1IcsyUVYFNn3PrgbTmifSdzsLkQm0+TZLB
wJTnk13QGVIXMjUAk1042ejV9ecipshD1Joi0AWARMUgbC90rZxlM2zNRYYu
07tF2iUUkzujRPoHdlqjA6oHueFmwuEMnMvvZw4H2w0P1Nb08EAcb5OSgbap
fHa+nDc+8qrVobUNDly/M6tsyH9IZt9qyaCbOfK/UTpKX3QEAq/tuUJ0fNZ5
/4pQ0rB/T6w6WqFZBxUK9tAAnISNLoEF9TjTInfsExL4SXzH9PKhAey8pekt
+SfD2R3vUhlYf65uZDotKg7oOsIHpmtSM3GZc5kcykzQkYHkJxtLzfdUhPi1
BGURvxUaNWfZKtpEpIDR/Nieg7DP0uu9W7SU10s8/sj15O8HtBqyrgBCRaLB
3xmbTswqp5iQeRvgwUIjeu2O0u16j3m4R9BSjGpl0aC9uR5zB52Z9bASigMN
zqHTD1XgnvwoiXqiEWRHMojq0Vr+Px2OI92hAecJOPlk38NMu5DE0OZYPYIf
4wWHIALiskiOavWKTzEzBKCmuu30KTGtY4ijN1ONDPL+Z/CFenlWaUfCiO5f
PVOUt2IVHeui4uctHnOOzWA5JssArRVpUi+uYTG9KU27Udo8KjSCUEwneamT
kRt94Nu+3jq9b3Am3iJ1G9uuferLdZ9rU+uTyJ99mZifTB8KA5bPm5vlUNQD
Pudl5EJ4sNJW5jMilOOcaYUV49hZwxkeYmYp/j2M4fZm5dzeM7Qv3vMXXJs0
M3e45thxq/qKI1hnv4L39In3p8PES14Yx8sVwzlqpu+bwp2H7K0rKePByx9b
OfzaYY+dB0OGre+CHy0b4sWHdac+96pLC18qExkig9feZSPVJS+pcTRyWI4e
yX2yAxchrR/pYYaFcKb8AYnjp2hGuVbWrBK6XzPeY/sRCbV7/rsWz8Yj5eK1
Fkcdhb71z5d/elxoDyUTXrw3NG/0ZRrOmCDvz0dOgO+oIizxv/AzFoAlAERw
a5/yo1daIBZatsf6saGG9UxSUVj9+dPQ9m3+EhgJsfmt+J2gjNGK2p76LBij
MtaZGnExr5ZJX9QSpOCYDdBHMPDhzSu0DDYwIcSXs8qakfQ5SIzktWbYBD08
OO7nnSr15NXmzpjivG4d63iPT+tsy5NWgVlrhu0fE2Bh+dEevNud7g7YghGJ
QibckMBu0b2yihBLKK0sEcXaJvojHyVjb8AP3XAdbnPt0j9CpmqxNulxesVN
Q9ooln6/2GxSRUtWTWkNgp5gLQDTEZQZ8DXB3vJSyYW5lIJj3hsouCDpCYVN
bY22uGdhZKDMdy54qLxTpNTDkvYzsU8DjWnjzh4u04bEM6vuIfWfmZGPXEiL
OQAVvdp1aADzFnQ3301BQoPNIp+p+SWOSKg+VufoSYDJlWIpnD5r4egAH1nC
mSdPntKMF0ZOZKrHtIGQ9O7rzbyYBbJ9OpVTLp1T/D0b/W6eZuwLmFTzzo08
Xgz6S9Wg+3w4lFiPc0QpUW/1AI6dxM59DNIqACTD9o20IYNzubvzs1GzbVqI
uOW8RpLXnsmFHUHRu4OIdIpcOKqrp4t7lcc/zf+VVf0KngZy3rOm7zI4gBL7
2PtkgKHffQftk0B/s30eVH9ZTc75l4yvCo1MMa/2DqNcnxGmvdAY83zSUS+4
2laTuWtL0CzyMz8WrenCWmwTmwRGlnAsrx74osTCwD4QQh24/jot1apu2w5Q
xFXDlLzmk2H5tKh3Wvn15B7MfSP6rFY4fAUSMkxzNdVHU1ZFIRpOUf9NnGHq
kdZt0O8MxYsPuyUsy5JEAZ3RlsFqj9Y3NyuvVmSt37W8c6c+uNwn7OD9IOLo
IizlE+QBMwJj3KykCX+d2f3/82zfhx2CoZTW/75Tgiek+7EozYfAZYFBlxjn
1dYHu2RoAcM+slBquJM7xAd2ZvItMlE1if/rKdSlISik0nP4JWndteYQeSxD
zgqsddX8M5fai1x1yihpi0UgFDW+X6aYmMnUBdZm0rTeuuY2uIl1qopeZw3d
PvuMWeU//NRiLWGWDs6U5zP+MHEz/VtOddzvbypkr6821SScF359UmcPn7OD
yS4ny3+KxgiLpMba2/FlR+XHihuZOC1vMzoZuzAGpCmU1UbN6Z1IV/7/goig
v7XKAGAMW7PS9mzJf+nK/lmNy78Y8oD9bvLYxIrQaB+A+nHNbMRi0CK9hT1o
oO06zuDbIISwIl4xBzK2bTkkZer8RdO/Rkg4rOvia8KWkn9uSv2p89kqeX9j
i5L9f4cXc5+B3aggkbjjX1PDKIaumpeKh5iAI1+HtkHLKtJJlewIf5M2xu3M
Rs+imvSnjYtFuyjXJTm1Obna9NoG8A6K3A2SuyVLce455RbMMyZWwvZAwS6h
cTOVcjySHSB15bwCpFtYo3U8Xrh3yxPTGmbrFjaIEmT+b9BFTs8aahEvQeVp
WYq6WA1JPSJRS8KGuQI3Y+eTBipIjIawYDgXrXn3/k5buAsaVPAcfBGrYt4z
XGE1WYhGoG0HE1uSxkXqcc2mUVOQUBBt+/hH3h2yRSEj/pRuWCyQVHVoOTC/
qCtWR7ieHi4AU3b3Lntx/j8oJW/4U23j6jCHIz674ho73cjIvRnxzkndpCt1
skQNKsTG+JZjKZbeg2T7tv+fq/okq3qqjAV8+vrWWgMSTNoU82K8jGpxV+du
1G9jGfFZC5wOiz30nnoaqPsFoCFg+on+aRboF3oHkuDzA/l3Ee/Ax4RIEEt+
EFxSN56hBVRj8kM1/dkaWFqxxJ+mUIewuotfyceWqRNg0OjbnId2pAleUWxB
EFtw8mMZR80dkyKuqqiUWydke2vluDwJOw4oEVqHL7kzJ6pl8Rokw9uNbbiL
YuuG0p0xixmh/M7iJA/tUlJtlBkTffAmKnqd5MmPT/N+9n8+QRME0G6WaNCV
Tg+f4Ax74x5bg4lQQO1zhZD92ZPlf73HnmCFxoSDJNeN8NxfPtu61pEgtnrE
ppCxDT80wENrfV+yEyoLB1INeKtJnHS2XLyY7tJFIYdaU+MKx43iudJyHv03
s7YI/8BDdGXJfyCF+BlkReB4t1NbP8B+UlqQqiDqn0Puk3hQN8llyKzbfvNi
QodYwzS6dMpGAi3zuYhI0sPoiCx8yl6DIL7h1gw3bIjwef0eGHs8CpmBFoYN
r+jhgdLGfNQ9o6ihi1Zyvgfr9n0ynQPVaDfUHAPulMlUD782X9YSZTUJ09jc
dXr2dCDk0UdzFavMvPHhFszMu9YWBVJv40U8MCELSxAZHiUUgq+T9spsWeS8
and+rvqI0kgMwbHEPZcc6Q1/t+h/Mx4X/oSinUiEBfcGw/hVXSYAS5occCVI
6ipPtQ+5i9thKR9gIhdObwElM1BZsR371T7e3u79X2OWH+7TZM0FtVwwkgkL
ki7AVUjOOJQeY4QEoVKaa9wEIVr4FPjjp7CIsfJ90iZOMlvjhM5pGPssMaYv
jIAu+IcAOh9U5SvJ8y+rgXvngnDyi/YvW85bu5VwJ9fY7ngVEPBkLzpDuWco
AHKMosHsMiXi9BERVO0B/3pEADOL42DArUNKpDXmPBD2QX9q+2QAIYAL9e9l
2Tnm2d4kfLClapcEUaXd4Wk2JCl1uBekcX/H3v8oDKnbDYzj2Rob/BZw6a4j
RM4hN/kHF7tSTWd7tE0VB8SsJ17K1h3aNIp4u1AS9Pb0Qh41fBEuDtB+imdQ
oHf+G8iC1kZXO6zc4sjgbcGgkZRdfW/TuVWdoEkQsCF6Vd1bpsMForTEd80E
5CE7+cNXV2ht34qc2t6MVxVtoJNaivZnp0gjI+LK6oV9Bcqq7OWLgsZdXJym
94l5qZh81FEAWXPCsU2PsMFohOZzKKJW6o6cEc7KK8iauxtpYoQ/ahl2jDLm
oYgLb4v41vm4QFLO7c95k7JjdFSm4GEfVNCMewZStCrgwBn4OW4HCJkzao5O
k0P8iCuZc6in85cBCAXzWdiaLRhltaXCjCavg0mCp6bU8Cw04vVF8hFJZcD8
EJdRvSwWoo6eF6SV7BP+918XQ5nNzBe7KVDZlO39QiXJspks4zPcj+WtsNEZ
lULZbDxE3KK5biHZtKgbAbyioN+IXAEzn4xh+dzvU3v887Vt63a324xqM8q7
EfNLN/BZpXsg/OZIuSdMrYIj7bW62sldFQebJ2oREYZqOp2eKN9TsV6hNyL8
XieqexroMsTDUC7f/2GhTciJastbjzqpv1huaQovngJs3joJLjxHhXwTfBbS
g8eoPEU/h6WJ8ri2BL19K0CAeoZJzuIFPMQzOP4w2dgl9NJ5uH00P0HoHzB3
4bEPjKrvqkJaXw8i2LSHgc4IwXakZIdAiFHdmvBKdXEK6PhY3ViuMnGxQO2J
yYocY+PAk3fIAkZsG6RAoo6+pCZPxeYRiVoUR9vUdoV7m88QlE+minNYXzWz
rkZu75aBxb2HiKlYcKXYhMg+JTknLTg5N/yZm9pKkWKehdMvwqeTkOa7CvcS
G0s0VRd8M4SKlQCuqdl3O0qzuMwOecRvjgUyTha7KWz3HGikm4a/3QkKPlPz
wSviBI+oDdS1hxg7e929a01XXkplfQ7pUtsFVY3gm1jXEj9VYFHmTiBAtE84
8gBsVejuEUp9kTySmAw6D1eZPPoMn1SAMjdp0C9a48H3cZBW5Qg51Zwa0f2a
nTgIwBlretmdqxoIgGxkhh99sTZdDvraW2753tHZa11xCO3QalHt/AOZpiDS
s/+NWPVCgUbBzF+fK2/up3jVwiXWOt7SswISLDXHTWKNJdARn+bMh3bftOFb
tnlMaJJ+y9MU2iif8Tl13HFIXjVAwxXqeJKlXsUHPKdF2fHTNwsGcf0P1rrL
duEq7X5aE0PdC10qfFajHfZrU+ovlxN4zmjYuT1eRQqLAoOTj0BmzzZxHvG1
38kd5z1n674lMYZn4w/Hck4Ca+7cuwVTVPT2SWwCVcXavxbTPRH6ufKEC4s8
IMTsooSG0hX+NbkraAn0Bz20RvJISZkmdOCc9QgvlTxelr8C6DG/LLt84rEn
fZdA+z/3Sd3oY3jP85uvPHI1ysIWpMjFEu5HMnhmyhZ/DOsxozwXjfIgvVqM
i3p6PBM2GKlLLs2tiD/EEBKrlvcWlH1TK/0Wz/EzdkJI9X+2pV/9Xs7J9Y0a
+g7N2s/qIhsPTtcQutuOOowObQplZhrQSw/0iX58YI2F1KJMhinU4tdHDnNl
5OF2QugrNvYJh/t2FuDuWPf+lD56NYi3vXnC/QxMxq0Q7SONKvBwHogJ8Q9Z
gO0T1eSnj8B4IWY/yVwO3L9Iec2vOVDHi5ZZeHL3p1rK4k+Aqzz11p2RnDXc
3e/n1gh1G5Y74hT3t3Zc/3+F4hlppjNSxu4npu7UwoqsjWrnnRamc2WcNWFi
i5JqFNU3GYmyrS1YeKE6EwoUmky6ImHwpF0fNelAFGKXOdyUVq0VL+nDyAPw
ikPR985DbzM6lULflG8IB9rAXd2uGYX5hlYy85zzGAuXQFQ1GpBw5Jx5Cc94
b0tFcAC9ZlMlsiziIlhvJ8UghoHa0yZsy466Nv0h/tVdanIjra2ecFkJaojh
6JGHgauganDHzkRpEYbwZ5/r5iKN3l+5wyYkI0bvnwZHxulhKP1hqqTeMfrb
hnkmq9V6iji+zT/om7Qp5XpGXXFqKebjlOoZeHSE0av5YXxuFYU4MFB9OO8A
bXVE20+JEvPAGqSOZm+fy1frYSSTm5w9vSmGVAnvZKXcIqVe79MW2gWG76Sk
92BcGM5yrvBJoCp9ybUy6WqKdJsXrwmHbhkvaeOQyxG5lp/p2RXyD00ifOCC
+N+yI4KRyiV/7d21sTwmCqDiJlHhCsxv3IuNhjTzfWbUmOIWF11a6NM8U/NA
WMEZSWNQANGlyrVUmPP5qXs8ZI4FbrMoaycsaVxikKP7pjjbH66dbisuyd1y
qi5K+5DNAlI76dcAzjkzRPvlwQqtOjh1mkarTG5JvZVUR+5GD7e9z5yRCksR
EtWtCeJgtQzPHSM6yLtkQeUCh/u2XM6pks1k06eUo4IeHIx2uf76rJOzyxrf
ovqWvFv+FR5zBdctWFjnx3EtJ8pjOQfUDcKiywmIiROc+PO6qD3CaSvkH5Mn
nR1m85Q8m8E1qTyRaswiG1JNuYpFFKOG4/KBiHbSJHh4HTR8I5s9e4sJ3Yub
pL5WH94vKkJHQjCO+IAde9hb2TqM2IkDpWyE+eSsYaLPXC3pZr1xb/y0//ZN
jpXuqSoCrpXJc/vXSossgu++XPQxHbimZSo1y+tSb6q/rkM3/Gl8QxQrpPKd
rU/OlWMENBTCvdq8YXNgRDpupFvpILD5E/QS9sUipD6WOFOnscSniaDX+dk4
Gfq5CVSSLn2EDt625sc/igBqgxxUDXxQr6ZUOQS1wbwU5xUIoUDaOyW48lHx
VN0gTt3W4FGvKsBHVdluVu8uso10RP1FNNlXVAC5rBfbsQH7B684gPztJJ18
jFV/xe3qNzr4ciCuRJmUvXfPy6e5osatHuKTE2XIvFmcAkyXCoF0D1vqtEtl
U4dlvyrMIwrEaq+6Nq/QvKN8RTxM3AWMcBNWGSgCYgaDuJEFt8lB5ijnOF9k
0mbFbDewyGg4C1Hlx8rvqDD/31nAbkVOcS2K2EwYpyjisRd4OOHhKLryKYxw
OM8272F7DcQbQwDCy1HCsXeqSxu3V9bwic5M7/dISbZhpQe/rDPKT6m8EXfa
LMfvdTZX3YTK1c2VFj7YlOGjiNPTuy2rImzx+lf6Fa5MWIMVmip7F7VvWKlJ
IHCL334tUUbWzGMivVdwfycGzrmDybVvXqqG/tOQ+RxMD7TRpIROtnvj1ylR
BfebE0FRlnFxGop+aPnZjGZo6yo9oPPOb3BACQB8z4MPVKCCWzRa392ljFEa
Vh+bnuD8C9TnRdnA4fQoQ2M/O9mhmmN96gXyfarMuzNJeouyheBLgdHBkiKs
GebxxtXaw1RPDXjEvudbEvILFYvN1q3oTlJGqnAj6/aOTdQkzx43fOPnVKuf
THugl5KrCCJTY8ZTpk0OwDSxyfPIHxhPqmV9MpVYJxQaKSO2P68YdQvQyxA+
7fSixKaixrXnPXAjNiMyR1PNEyIz/YGWpKeWYlrj7RaJprCgnkR2hRu1ixWC
Zwvux51SeiZ5fxah5gvyz9YGUrnLhWxkrwYdXHtFY0KXa4GlXbwu/VELcIZq
h5Km4SbgS9AUrqwlekdrQZP/aZyQ1Tpd4ugQUwQMJXcB/2t3GeYFKGrn6nJk
+9nk8YLrrvOxTzvMv8yPMIwD5GesuUn5ybvfjKeSisr2k2F/GbdOmAkkhqWK
sL8KMFTYB/Oi26Tf8WwXT/ikRN7D8ichoUlJD/Dwq962UH61iMXLtpIF8zyQ
8UtZZLSU4ieoDNfaeqXRMRe85gwyW0uERmkNumqNCkOGA8kmiosWZk9FW6uV
xKhGODOi6mupRljb9dq28dXFV7Be/65THg+CFCaYf8HYpTuH4ueHbTXCmDF+
MCMIW87p07IQy84VpHim0x2rgEbkWiIxLgVM0PA6juaTqnss3Pk+4dmBzBl3
JceFU0DZhUZ2bLR6Q5NcBrWjO7mXXLxi1pno0ZxMAwoaSwjx2PO3D3AvE9Lf
7kKzXY058pghCNe1GZdzTjn1umMeoCB7EPRAHMEXhF1NImMDaAXUefNyRE0l
ImbRm11bLeVY5yPPmDKOTZKpRCGvxA4JIqXVHKVDxuf1SXUgrukQlNBfrC8h
VT78/jKkZSHAWkuVYNP9il2zgNOr6SOubbX1NQQXrDQdGdWLQeKCxkSWjqaW
Uj29ZtybZ+ioChSbn5cJFnUjo7cXOrOSPrxP/mMraPtxbi9LlZaebjnaQ9pN
b9ztggUR6dDTqX0xCjAQEjauCNw6YWXy4icJywiGzoJZQEfAwyejqVydWeaG
Xl5hWWWDxXoCJ7eMZO7TclrPRt9yDWp9SQ93CwfG4afLz9umL25nJSyHt6Ds
j8AF8As0mevvCS6xa0jqJlUmuruSxXb3w/GjFmXeye1eSa4kjhSvZg/Avw5I
fj6yT6YCfDYJMsQw9MT0eEVKU5JU9JHtVX32uo3o8FStcC4CK9uzueFWqznY
8bLzC994o8Ze3qX/gW4Ht2SOcwn7FfzlZOuSwjweQC4SD1MmMO8FwRnqjHNC
zxBWy+4jYTQY92Tu+Kq/4XB3w1FA9Jeg7RpAGrIQvqhUag1EZ0VVxhtPDDi6
ZckvFjqQ3jDXe/tuxUty5n4l5sOjNb6f/AAZhKY9VXBbPvlEDM0Dgx2K8ROn
gTI5lsOLELXwcDz7yWPMiobKduSlHlFPD/zcZSzn5P2IR+Xp8EmEE/66f2vj
n3axrCf73jI8Fyfzc3SgrMj+E3HNZM+T6K8BQOG6YBgzFCFXf40QG+X8C49d
zKhxc4T1yxIT144CVkTvcedl2nKaKkAyfMyDxNuq2OPlySQto6YR9byLR3kP
sXHlaRLa0J9kB5L3SQATI0Fa9dmGMQk4Vp0o6oMllIHRq3ig27NRVUibGmUg
uzwfA8YbOOqgHh6RIBPFaWed41Keiko2NlrxKTgq8BlGkuXl2BB87LH6ohjZ
r8ThYstXxm4XcBFxX9GrQ6gYLCKqvzgWLG5CbvRTSc4XZQU3G7CBuQbiZr52
TQEBJfv93YDwwPD/0YxjW4M//mcOdX9uGKuin20Afl5bsVS2m1xVt5KJdF1E
si34sQw5s3q/1cV/UeF93fT1fsCerB2tQe95WfdiN40GCs6SLHgciw+xB1Mm
x4pEK4DcNq1mOxrlBW9Ro6iO7EkLfNuHVnW+aRSK/AhVNEIrmN624RdNwFsS
Scjuj4yD75uAOJ+Y8RWncyZtS7fZeVZRmDr83XivOmoUc5K8GkoSTFMcocqu
rvOKL9xYfpJELIPiCoaHJwwVigRIkORpIxsfRW2jMwnSJ5BC1pRIyD9I0pUG
I61zR1TqZviOyIptiFGcbJbHSqhRjBIIR7UV2ngc3LT+NCcRLl1gn99qzb4i
MWGF5U84+mrBv16DgPFpTWSVYHaFYLiqOxm1xo8PCmYZRGqyy6HbIWMZnyqJ
tzP5ZZ0rr3XQvKnSiBz0c7K37X213xfX4mpOxuuV7JWebhr6tYowdx1Fl82z
msSMt+HLPY63Uzls45TmkyZoTk1YHoZU4LEkeVkyVsTBx2pnSSBRYPv8dmXO
8CTMJoEvhrcHXgYMXIpv+9c2A8ucyJTd6BBluZwngyuzCWaDbqtg2iF8ew/o
T2Cl+GEHS7swLHPxKHqt8hlzUUrixc8IzBRnL+jMI9T1qpXu67BjK+rCpAgz
XNwmsLfSyyeTiSHn1gJ6V/HmtwcjQtiTWHwNmvIE/C1jUKwZxnGU4C95kEZu
3S062D9WQLYnMpcRy7yI1AAfKO3tm6p8m3OYGfbIFGWx5KpFBj1BGvVdQ76A
qoWxuz5XsiCtd74wD/VQOMT0xcY645Y3of5yMOrX6doaXnolPukZCYpbTYBl
/wO6GhZV8j8FI9VKRcSHcJXKXmKlCkgdBUc5fmu5Fh8bgWUQ9E98Er+plsRy
JVfO3jGJMp70g/DsIMzwvSiaKhM6kcNYfsmIF/cF6UCeau00BG+aD0F2L5eE
UUFJlu7PrDTcdc32d9AbWJQpsW5Gv+Bwh/TyJc1xQRvkHLnOoJuWASmN4j46
OjchsxgIZR+HqJJBlg2FvdpsMN2exkqhxCXTTofPAwAWvDzjeWUh5ttR1H7A
kqs3uI6tmQg++Gd7IQLRvhDimQ2Ukzo9ZV5iAoHmsmUfQABSEzunAMRGSAWn
QiXorVO7ZvVB7o6VwZVp3VAQKFzMmYeMLqjz693i01nJj7RdZh2abTGwXsfF
QgWkTSsMYFhIndrWnlzIYkJk/oQugPloymrnrFHhhT6phO8H2pdvOKERMVB9
uZkZCC5gOpNeupAELG017PVG6pwYzMpuOYYU6m8o4ZmCuZ/FcH7FD09HA9Ea
SAMkp6B4wXQZi/rB54h1xIarO+ko7AbH4FmgMCOGbDYwdpM6LQmRINvYSQNs
RBC0/kBUjgawa0x6WoHNihhfoX+8n+YLbP1fVfKTwMOz3CPe8UYz0Vu2RPPO
TE/zA1m/m9rplt0Rf+5DLaA/ZnBTqytV1p9k2g3x/X3vSdEaDSqY9HDKNBA+
E3QYmFZ+2MfDtqrUFl0OT9H6iRAj57+OCgf0oF0v1w0qG+KFMqJy7P0nly8S
knzOBT7qFjBYUps0aWkm5kIOaVkU+znsOZbylOAVsqaC1TyP8ySGsV+aEvuR
UBMHJd/GZwXdzADSbjDhCia6b0OkS4UeHl03CXTgx55VbZopyBd/IDgsaj8G
zisYNMrwZ6bntWU32J3PaRWHXhtnpOw9kBiFCp3YBKI/zk2gNQ2Gg2bQr0fI
OLDRomEyyTBU25Cy/Zu+6rrhZaL7r6v3KbjXY1YEAWqvFyBaKps+XRbiW43x
2uQ6tThkn1R354UyMIX8RQDubNFkOHBTPXf1BvfuYJKGrw0oXySTd8SaegWc
GXHWpMps8tqvzA6ZNyXPZ2U9jJ0bpjzzzs4xdC+lNPq1cEmsMRQv5HSwuTMv
n5EGWRMU2nYZ3XIqUEGprvoWBBbHPOGbJ/EdVQUG/nBetnFJF8I49akl50S1
MJUAdzcmZrZHWNFWUgjYfaIcqSxcQ3GZUKdKNSMYXo/gSlya3ezRiMBkbCf0
TQ+gP+Wc8Yv8KIj2jK2cuGRz+qx4Tf2A4egjAVhj2wT+jIgFQYsM3Vxj9R/H
ceCbuxK6q7CvXKKFSN2KOQbVvED+pde50mA2qQb40tFcIpF41AjMIAy0Qvhg
iVxGiNaMQP4MaKIDe9PKgRMbUrTf9TEzC9kdu+nPoyrOSSsoF7C+NOObB4QY
Uhw2WHc061/KOBxO0LcNFNwHVlnda8u2hQrcStqPPO4Z1vAbXoSzRdeTICk7
Sy7wuaNb1y8XpWvC6zlSKDy44ejr20xUeax4MJG0yToZuzkN+e5CyBv95p66
GJq0UX+k6/47FjbyVd5Pz2waqNEqP3whPuMW2CfeMzIubzv5cmDrzM4LyzmN
MJX6kiIMOUzb7W9DlVg7kiRNagPerqDY/e1RVMxSaE5ERVoVQWD68LLH0IK/
1o1LloYvVIZgZclwrLUATnyZICOeQ7VQc8G3GY0J3PmuMa4WHxAL4zQyV8gz
csoqHjcq3NVxt4F2o7bcKPvjxphKKtFCkBqqSkx/hECGoequakYOUqj7ttO2
0MTJwwemiRo6Ge9JpIgEwB+h03CtngWxmjWuQRnefITwny3Xhjw978nkEy1G
X3GU6tpPtQesV4VXmDsId9EijspA8hV2cwsnHktmxyOSLJpRD+8PVWAyCj+V
0fqzGt08VwMP+sR9Jx9kSdgCxtKrCf+fXxdmZGFpv+juN7RNdHtN9DPeXIZ8
0G6rheLyYPkLeSVQF3IHF2K+mo4T82w0WImfXmgj+5NaexIHVKYSVrN7sksw
HfxoK91+VA8W+WsbgkdyCCailY6WI1A5pLBfCSP1OIj8BogxkDx3OA/ylkTY
5i0EcNZb0OmWP4Z+o1cuK7uEk9WrMwcyZkzYjXAsqx4GSMIctnKQL2xhv5OR
RBj01dufffOAUEv5sMIKT7FnfUpTkPGCxw8vI0rfMIyVEd+34ObT8cD/CeD1
rgVtAwM6aIoE9VZcsNXzb7h8JXO3KOsHC/7T3YkfICg/DmpmVdsDob6LLczW
QgRjP/1wpqjNPQ0d99o9FaJm+aSY9q6bsGS5SlggWj1Sxcv7vPr9Lms0e87t
SzVFl7jWN5PUm71sXAK38NIrbGkVGJ7WdpZChl7Ice8WZ5ahUWGFg4Yv9IiX
PNv/CwGVJ90RfHXdWSwmB4Zw0Dp85b9CNWg58X8XoLCbmJ7bABmg/Fo+4PpK
e64O3nWulfPF4znRjti/e59Dwt6UZ9HazK0MyPanA8qnifWjqia46U6baUCX
uwhnbr0P3aFZ4cBYf+8czhGa5EmF+1Ao89/v9B5QlK2G5i3+ern8zdYMGRuN
NBwHLn+HcqOtX0N1ndgmx9wH45wMhH3MfDovbGAfxiGaJ/nj+ND6cMwz8X9P
f1HamGql5UGcYm4uKu4EQ7EGQ6G6dkuV7SLJZ9iZC05jK5j4It/YWUGUUwVm
dVGiK3PVd80E6MiQyFbfeTpBPgK+yQVLG8pfqR8rE2HYfyyrsaSa22pDW4fz
sYO3llPTmeZOz+ePgCtEWIOZKNjnhYORlnfuwd+11fwiIgLLgWX12YasmPiI
viVcKYYwn92nijKjLWGdfdqxG2kpwbCSIQXAq+oGDDOx3ckDTWdxKakC1ZX/
ApUqegA/A2Xs8wwL0FHhkOCtLU7RCBg0QblNj4pK8t1WlTfPk+6VH71KRKXm
66lSDVp8x5i0FwJ8tDjtVoq1JDUZFcMZArbIjhvIgxEo9Ri4ygscsBr5KeO/
smxlo7qZBHAfkFZcel3hEWsgEhMxsq9CMzS7hSdx0b4vd0UN6c2z2T3Clo8u
Ps6oW0SwwIxNqZi2/jZUDyt+tdDNr86NBVlrm60GcoVzrBIoi1taWYh+umWU
M7knNHrOvUw30ydIJdIKcbNHUb9ZVWcSMgMGjFwPDsvCEqBykDSkA15OxPke
grsuyRHWjLOeD92SkMHVuPE2lsK0NXOLEklJu30JiT3iLh7HRi+dcuyEu0KC
kLNoU3X8ziHZqzKpHoA0fx4lX8AtoC65Pdpx1K1sIwPZHQpQqTWg6uNm4UwZ
ooefaN6NpqzUEI0qUA6ua8TBcPdcqBzhoEiClMO10V+Ca+8bUqUF/+AUk7g4
BjxVFRAS0KrMjYqUZ1Fpclvviqhs6a4GRT1Zfg1n3b1ezHPRrBxxE0T8bN8R
K9FE84bQ5S/ra7VtCH6wH5e+riE8iz/0hbIBANeTkQ8CquZrMfOjLjGdJMwX
+LpIZSDdUM8o5tyuaE/PCFkENij0gBTHiW5588njggppz3vtFrOD5kDViYru
UDioyrWIKWuZ3eIfQXImq/gsEghn8eLMkhdpev9wa3+YQ76AmCdQob95bsRb
bmxVTCTqn3pYaTgPAu7sX+Iv4rTE0gJxh9SGRNLmsX0b2Xd3Up3MaM7adPkm
1qfnXLwav16tVC4B2u5dXiA7D2ywhveLt0pSnfFMAscBw7fhe47kbEcawxqe
feG9Gn35y4qstR4daOvFraRo/qHB+Ph3EZMV65KAvBXYjdQxjp7YGAs9yZu+
lB/siN/tZYc5VGYKOOTKg2ocIwQWW/+eztZKmZfkv794XYrD9WahfBraCVbq
+rW1On/d2CgAtFff/KHaE2wVXIsgbJ9vDGtsnsScWIMo0wBTQncgBtzkdZC7
/kX4f90t2MWSNRdUHPt67oCeIwpuF9t77po2fKOC8Bg8mWJyiHs4XS8MeHgM
hlHBq+fT1W6dMoxjjL7XkD8ozVZ314DaS1ClzI8CY/5xaEgUnhEZm8jXlCHa
khF5BfENYT9y2cKam73OwsxVcSrDjwh+Lydzt4WiT2Aiog5ACGGGHaArSuzb
TeZF7kbcAkVZpLEwSlZN+K3hr95NdMOE2j845BtnpptOo2kNA+uWLuCHFgiy
FoqeZKe5xxYop2RWDlY/+SrQ1cN5VPPtfuZ+VooPXncCn7ePOmERDiROvi9O
N+yzfzqGPsIotzFy84MqC5ycaouRt30BTrKqCHHUUlqOpLu/zH6lH7JzQyYa
eQGWDGY7hgIcPkToqWMkxWTgUyGSEP7LCKJb9sPLQltYf7x4ijf7lEQR4Wxy
e8ghRqD1BrVhyvSz4y+fFSN/kNgzpYqwFB68YzoQGukMA1DKFQSPOSYCG5nj
xPgXxyPMAqemQ20WxkfWgF9EFQPZMLndI4lGME1gQ2+C8cFvHxbBw0HCgP2X
nBy5bFPIOXo13GsL+IVLWFoDIR5lkLVSq8IVS5WGlCcth3uRqWP5czLlPbNG
+9FF1meH+YbgFO72egXUYaZatVLHu2zokqPtcIRMC1PfbFKwFjVWyEl85g3n
lke6CNaUvIW/6Xu2NDsiwNbLfH2gIiLRrz1ej79mNMB21tVbt3gYBLgcX1dv
t/h1Srbp86jigqLpaCXcWguCe6s7RtZcDmofCtfDYPRbwvAJ3f0gQsQri6+z
XNmTITn1MN7zLsP0/rBtQ0udAVq2FqvS0O2N4P+0gX0IRP7As1yTzRj2mdUs
P8ETujAqQzVJt9OuMVkhl6dI993pzW2bVn9ptSxOOIqvRmrb2QdxXHPXQk7X
qPJwnYZ0d6IyIeYjMv2RPJdyDCF5WFRgxRGg1Aqk2nFKPkGNmk8YBKLKOeuk
d2W2UWUD26iCBF1HKcdNpaC818azQ46jWwg7caXvpH1uW/fBBWb7vatOpYEm
TBp4K/AWZc/yEwPM9HwGQTL2nUT1Hijt99PhMW0pMhLPTjJi9oc2AvmUNzcg
FWiXyKXPjtD3kT1pUkKGf6GhdfVDux5IDCFS16jnBcE3MgH72xQg6iHqKK4a
7gqDbB14NFlIuLl6f2iWpTuSNmhda1fJLOUNB8c+t2ATUsi/BxMnMjf1MY+4
TcpICPpFv12gzLD3buUzmlUwXsQjY5zVAkPK8ST/peISzENVVmMe3WYDI8Jx
SOU0UmHR7ycI6Mxq6fQcJZUJzwFx91x41ZsNiFdrfJymBqUbKfSeTqgiwFz3
QgmtAcIfBItyFMTXKYTFjAzTJDTeAcOogoo0udFshQDfXjM+3+G4Vt0uWdWS
2o91ysH4wCEJe+2Aj2G9lgfGFHwOxGRjuLsM/rTlhghN7J0+CUTZrlnEOBd0
1ivtklCWcVvM5R8Pb/9YeiIMgZe/pG+t8AaofuhfeoiK2tBIAyHCmPBIOxsM
sgmKJUHEx/xLSCVrGBjzlzrJklYrEwT3j1WnJddlZnzBNOMqWmUEgcHvTrn7
wjkyly2PPAOR4SDfl+bbwE9l/qJyg4869dfnoNeCbi/71D9t/bo15VYRdUhT
DuQ8UNoN9ZM4lmuPjWWgo0Qqn+HpSRmbjfV8cOROqouH1EvSq8aGnX1ehd8z
bU/DMwBtsMlPQtjTiLU+Nd/qehh09Scvd4ikf+Fzusx1f4hCJHrArrMTiViQ
dKQSKfWabxa0lKZvIrPK2wsuoROVtksWNewZ4gDeATerKNMVb6+qXUIWKhGV
4ZGb1djcq1htjQP5ZXiq8uad7pfXO60CYKk5czvuBAvhgSjIOPnBsJumpf1J
AZV7vDvWVsbkcWCqCpZsy9iB/6dfUmAwy90kJWtLXtvf/x7XdqNMHSu/iiH4
PNI6IsxgwgkwpL6NZ0Oz3NPeyvP/WBah24/JUCGX51xQWdoxjYJrbOTr+CNQ
4s0eYqsqC8CQ4861eqF48Rj2dXzcmJoTGr04GkBM1gcFQ7a8Wt4RjVGz8mkp
iwNHH3GcaG2wakUxDn9WgWEAOFLAlw80V/HXn6/syw5YgsenUQVQQDLmOGEQ
p67eEI6NzTxjy6+m+89PNR9U2j4jTqHBnXi7k/Adg3L4eHFEig85u41YgAg1
c3C98VidAcjVgxKYAlsTqkqK3AFptFZZy8sd0GY6V1i6hkT0lnxRvagVmROK
oEsEcUeltldc0KczKwjFkTxxKkCbwsn99XbCeodyl2YuvzB8k/2bBXipLyel
JMKjyHhbiGGC/MLv4zbNBu63bQzjgUIFSJMFPcmqhE8LFAKPajMFtA5WuYE2
8KyysW9idKt/JUSRkNH/IMTxuogsll90wRJdBZm3t31xqxIPrmJ412sM1kPr
PNZ/rB11a9ECTM4M3zrbpRG1FU4HNL9IMOgxvHNzGVtNbTMe1W3dM9/YEiuK
a/K2gqKzTiYTRzm8l8uMsmMgrsek3Tl2BletoSMKlrbd0FpFqSw8e01Td1KG
vs8IYw07zQxH+bZDJ12vqAjhAe5ngNirMOhGILWRqxIFNBjIICKmlhhdjQCS
TFgTNayL/CS1N0el3Cp/cUv2sNfA3l50TnaFClQnGGyDzpOMSK1GSm2n920N
44sNObNg4gaHBll4N0vFAj62DoAfFXMWJQEUFJui24GN3BHWlaOtGnkbBsHt
Sw6UGHepBuoO3kTQovqlvMuWHye6TiZewdbtqxquS3Xa915AFNgsXw3aJCBu
MKCEWUIUefddxhxvg1AFEJ9oZSxxc4ty0qUTnWQXIZ4ciFqCgpFCwNKwRnP/
72MWdU2XK1rRl8xOXv4wpIf5wtyOrpzNFWYOlLf9qo3rgDRlgykG/G3Cu+Hn
jl4DTRNVVjqqcCIraFH4fHWQmzyOPp+UJq/GrjTxNk+0D0d1yyitNFMO015t
HFqXOVZOw3Y6mW/exR1/sERmsK50bZ6Hr04EE4XaCUNCGH8+gijgJ9rV8bqU
DdtDSAuqjawV8rN9gFMVW2OAvgj7eWtI1gqmEt6jQTETd68A+Y6Xo6R5yl9n
bftpYC5VlH4B2LQHjvpBTEpVIlGDp8lUIwkm2epUuLSIhH5T4l0nCG9AqO7+
ZxnPJnbBQ9c0EpP4AbEwaNrieJmvU+kv91TKdH3cvLXCL3zfVZg7fFJEeB26
w7zEaj2i5Tikq6MHbkjnRsSxpmp9oaf5pP8MsuN9jJP4ErHBe5xC4k27PWZb
HhNvkuJH2IoEOf/aeoJlaxsOi4qnAQaaSjLsHaPovLGxQaPSqqWpeAQLZTYp
rDLIp0CsUMnUlUyLFx8EYp2a69AFtYUepUv2vMRHtIN85OJov294Bv6IJ8Vs
dYjS+GQi3XkGGOpDcjugeQZJV7oKQTg4kmP6awWQwVqCuGz487/68K1GMbzn
vvaQerfBr822oc5q6d9phmbgVQt+EHS5k9dNXxFXVKgFWEU0LhtKRhT1C+4W
E8TsN8Ez1YYk1PFk+IP0UlBq+vhhPcmPBZRFFHyQIYao23chPYl0D/U3aKCs
rC5K4gaQY4ecA9LUtnYrPEPQmisYGbesCyjvW3Mg52xTtQkeOG5iqlvLMalG
1AMYMWt+Qz1K4CLdXmiMvvoMFHKlJWxpAVVJ1l1zFb3xYtphMHSfq7EcMK76
YVMbraM1ffQODv6HVytlgLSE8oFo9EAYpG90VsOHbOJTFncZtStWFsb1K0kH
4vdGJk3TIDU+nnC3XuHxhXmeUi5CHofTv/pUR5YaXNUeD/mktIKjeWpAeu1X
sF8z1tGPQnjjXeYVjsiv25o6DuAWEhF9H+Ybv6lFGIzJSk4R5winOYHySYBT
GxKJpF+QebRpLwBW3EANcwHtUONNed9sn26Z+zUxOUIG629NQ2cL2yBiW+gD
/8sbu3MNWiR1V2cAH3nP8E/bVGlr5dgDw5lRNEox40xNtdXMJvCDLpFDgvQN
csRL/cpcOQ9jQQ3mPvH6G00ywoc1qOaFZ4hUjdisfJMZklOAUmJtHFnqI8YP
PZmhmGUBsKBhwcjpB41ZJb/dLce2f3FOHopybdLtQkQtwySzec6slv7n926X
kKacyL4l3iN6LN6haJ+u6v+QEFCxWMfUZOBewrQyZLoBku98yUr7e3T1k5bK
iRWR4qAmKkzuLDBFQU4lsLbgCjpmvIiScMSPzckE+iYMej1aEtBuYU7A3N+S
vJ65XfqyONuScPTuJ5xmskTRHH06K4j1+kudb9TZcLOQqNMEgDv/vhb5Q8cJ
y/EXDxkCLmNuMrVD7ZH98kZWILrn6oyxozMUmbdBQM+QA2aDy2oL1kGp/7ko
Q58fpMcRnC0jXjDradQtCOxQq+cVpOl/Td8vyVHIWctdU19iXNGtrRjk5hH5
8qnVEN70OJ61kDt4VNoX+mlX+TZDjCyJU07anmyv6NnN1qFR3zNaMzUrnBul
NcrUFikjW1hJUecSAd02WqYJxAHUOTiNSIzbeN/plE3OmVUhST2vwFHM0P9w
W3kTWZzdlcCq9hicC7HPM+AELB3p2LUcyM0Xya13nZVWFyBYkTKjLU33Fg/A
ERO3ddQrlHKl5GGaRbziM/AhU2LD1Gj0OSg4fm5w6MZ2hoL/h6iwNl56KkFD
XT0A2MiHR1/HuuF3jkzIgYtgn5eOiMd8lgXl9sAxcCM10sJh1DMEf6+4TscZ
5B89eZiWUv9CTYAyeMiqoVkS1H+S3KgiswZSBRi3MoiuPph7kbJt/+BtU56j
eOvRZbWUe6YWFESz75I12D2+yV3KUp3XSz8IrzeLvbpJlRrC7GQZiAxgCgxL
E40fjgyLpcUJ1bnBmHi+bbmTTcEAuUNFCsKTnoCDt/5bNRkm3LW/EzxeS8qK
LBxxGt2UvW7iwcJnHdSMAIIZtN80yWfe3nJQhcgozRK6wdjMV2/mZVamJrHm
LK4oO5OzfYgyHUbCxneU74uddCHxzXIE7aaESFsu7wPO0cQ8fswGTWtyZpjb
BTIRufj4WYJ0JG1HB86tby/89bNw3JxKwMAg+8w3Vh9EA/bCDR4mKhDLgoaO
cFfzXkQCnjk7Go0Sa8iACIhxe9HqH7HkZcSwfY67PB3iAzDbDgZUa/AolEcN
y7i6v48FPC1SWVMM/USCL6BGOMze35sj+KHFKrMxYpSXCBq9ADNSgqE3adhj
z6nJsajNqjrGx5rSZEUY7Kxzj0a1ZcYTxr64wA1IBwHXun0qHR70inB75N5A
5o7fKNPG6CD5L/+YR7Fjvxfc5Pi0nkdhNCt9b85JlfLloraOVQUp2CWnqS9n
1Wx58Bviupvw85nBHIisZz9cNdadU/xUtzkL1JdYWajqrwKjMMGwqbtKmCB4
CS8jNPTk8ipT+rV24CaglVdNCFD4OF2iA5O0rZkVD7y2iPvhuPkORaRATdP2
46TN+uVdEw2HLkHAQ4n6/WsC9Yl3U6B9PzYbtgNAW2TyTNzy7XAQWOCrw4+F
WJEpvMhaCB7LMSbvGi2/HxyCBTuCCKyMaNRuPgKKrbCjUhvNYdLb41pxUlfo
qBEihTmD9bzHODTsjejC/iCL0aOYZPWmm1tIa9hjPY0RvLnEAOIruhpDjSni
C4iIR2b0XUaUxIwv1ERVuKjO6U5h82WERPO6RtsZlMp3gzEyLyzDcL06+iUf
JudDE7LO2O6lfp5ZUYAcyp7AN58pWjYrlfbioG4zSxh8s8+ExnnjCmUaorFr
lWs4aePB4fdQCiaDA7CyVxXbJM5PluInHFBymC83FNsvw4RdUate+NuYEGJR
u3CMtFzyofUqe5/aY9eez4EtUxeD5DrUbA84nYRrOcEgkbY5+us+d9BymEy2
JlKjUO7WTzgZ7qzTJEpfWlXf//J22rpXeZ/xMe5ayOLeKiYyctUlLB525+HH
ux+kQ+lYHmFdGY5cFq96IcaSrjEyzlYOeske/6jXDWlG37nX8uk5dG0ZZRQj
sDAxeT71PPv/ry0GtTxiANxgYtpjksQ2X01XDIU0pVylNhzxTRRUKTOwLyRj
UJ5qpVBxVaLTuzr/d1PeIUDD8EKLq0ylsysu3KiOCaXv6Bk+laEevAJda1R7
eazyiCEBaM362yeEjNyBmHQ2t67RTiJyRyCswI+OA58BGzjMSpxS1GsN4kIw
lE99YEyFSQiHVoYfdq2pG04kQhclozh3M9Vb0w281Un4P1VCY8EtdcV3smvJ
msav8X+3ZjuA3GXqm/5Hd0ng97jVW+FDLDcrWzxgOaVI+kDf3fzHKlCM/4Zk
nUzlXMamRQaT5wiq5MA1UpG/ii5LkrEhnA7eR1ddRR4DJLTGfrF7w7I5Ddqq
YwMexerLAey2H/6n4mrq47NOEpnnkHNSFLepnWCbNkKDFsDWZZpjHyRk9nZO
XBvK1VV40eeVpTQHFHSyB1SjUhZ0JdFj540xwojoLRxC3cvs5wuMwZpHkv0v
nDruXoy43SFnmiw6t2OoiXaQVDwftavRtn8eUxMnRfm5kArjFFPsFtYL8Y3l
TW9siyvcgr+uWZcm/bUl9+7itjGzJwPtNOX9Ot07+xTFfOTncAuxlHWaA+tS
CegqTUKtN2GpJkpK3bnv5bWQ7LCiuD4lwx54VlWGKbP3D9z4NUn2Tc7fNyLm
0biE2K9WEH5GqEsekShBjrfPm4aSxrm1HEFxP87l+EgoV7NuG7S4m6wCkbxv
wOberc2We2AH2HZ/2TCxRv0oRWuSJcnbzIb83r27qU/S1wkloDSCXAZ+2C+y
jOHbMXGqFiMFvq6o0H2bTMtFQuuCBsd4aveptRvUQG4BfR9du+Zv2lxcrYPi
DYfmbs9s8cCuPpEiiQNOuB1WKnOH8senn5OgUNl6FEEOAU5yWXQkNGotURJz
4prvLxLXh9vW/zq9oQ5pfLD3+9SWlkBkMpKkpagaStj3+xIM+qi9c1rXaPEm
Ppyrp441rq6vvepkr4x79HVZxbVagk7JzMMS5W+7QcRnExB6tC2rpAzUqBZ+
gqp8BkdIBqptit9kv/h4MXwHmgIxM2LKG276iJr9m3cUtBSoZxNUDIP0eP4U
yrFS8lsxBArAXiXjZBActF26hO4hscD/CG9oq7vmnr2ylo6eJMmk7JXqbEfi
N0jEoORd45C/KkFUGbN4/7o9qdyu0SQScjCYG3j9qj2KsV3rgabs8i2sqPi8
mnF/JocOyJHJkzlEpyWeVxtQXISrldgu9YO4gwC7g+Qg8e+rK1cIeGIDRa0l
iLECrDU6TsDuzEft+wcEEqF5RXvnyfi29fC1SyJy2mb9atydvb2r5PN0dLLs
RmZ6s1FGYMFIDTjfAMKD6IxEx3IDNp7/D8PLFtunYZYbd3AeO1Fq171XRNt4
89mw+KMNKZ2JRA+YrRyeTN8RwtjNwNdSeK+fIPt8aMZpw6MwWRX8DOayd+Fh
yOScX3yhoFcnf8tCckBdpZo4BQFMRyXqnY5j6qKkSxCNhAtiFSVWl+3LJxeI
quWnF+fOLQtmOK/2vPLkpIwr6MRk4aRXT/tjpyCG/PHSuuF+haFOQepWp2bN
nojjXXLZDIFDDR+DdaMV6uIauHJZneooY0SIpFzBmY+PwZ8u5lSzSuURXP1M
tJtZ6RWpjtR3dfN1gFAI1enzPQNCe7DsP0aAhOx4+8AuRCDfrHVV66n+Y/Ja
QANG51Jqk3OeA160unDTFwVvnRllu0Pviq9uu9H4Vu+gTWShJcIlXE2mXJ0T
/dK/xtVGnkOE00PIzFON5XHAOHjZmB3JptLejLz9l09MNHZlnIEfE4oiHKUL
TGL3EHKIIA7UAYoxD9pgg3I9wOQsqezKghnDbX23Iexz2GM/Pao1sDq2IwPV
f0T7Om4x/ex1Y4cMZ2MlE6p1yVQLEOgOkYsUM+ZvGM6v/OtKddPdeW9sb0uP
xoH0bWMfKayrRvjcARVOExnRQ9PWecr+TIMlGkeyC2S3RuASIpkEQtnSZe8S
S3jVLRkT4KFBunvuy7qYi9P6om1He4F+YIkMx5VPJXONvaiURHO+z+LKu0fy
EZD5o/xFX+aLR3pLUnZcVyez56Tb0sKgMJw3njktSlH+bKa/ATcS8YUAY1np
dp4d46cW2RcYwJaLBUfoKZEIn0N6MAh87EQNnYZAam39IEl5wf2U4cTf3r8X
iP6BrivRZ4YqLPz75S/rBnC4SJdGhbdkVPYAlwRk8N6Ea0N83GxV/lkLbFYW
BSbi4k5iFegtBYn2bKu8pnQ5QvPrCLols6/0sHbC0rncX0usqk7JTuz6qrh4
qT3EvoeiFQ8OcRwLMpnMnGp+I6/VdzH0UNz3B7uYGojSj9gpcLykSYnzk+KW
craT/ypC9cd7Idecu7tp/dvFY/pAGwUxuE3TZR3yWCL1E09g74Hj8NeZr85R
DtV2X9xlso0Cd2agSLDUECkFKKBiTIS5tqTgecXIUCRokMwEfy0RA9T0TSkk
YbVLr+rtYsK8WChfbTeI4f5JeDKTPpnAQXJ750ndHDSGpbCe0aT4RMSWNaKA
yZsgtQyvVytvo4uX/yOrU7Vnb0+bf4vQCuOZByN939ans1plqH6/PS+0cU7V
WWIL3bEsPaURYaG9Iz/gL6/DO8pwvbpfyMOmmNTSiedB50sDXhfrdZpJEggi
Rk38lj81DRAbhVUxg3cYwNYKK1mLFYyYswDxBjTThGQDaT4grH85e/bpnZaQ
tcBElnr8vaGeryGwmYEQCgmhkT0BxQFq3FbuPDazbSVWuXKE6bMWhDxYDrDj
faY4YhFM/q/7MnLPeKb2UWsBJnVhB1opRQtd5e4lQMd+DXCIrafn3M8twkpO
7MALveSDwSROanNB4jlwxKzH3lsGIMCt33+6LAy5CkbCLc0v/P3J1jSqbI2+
Yu2rfPgBiKBxIArFfW0EhTVrt28Df2oY5qsbXbuJKryHHi7LgIdC5fNVt4Fz
+Mre6iFmhJqzwqxzRGBr2CEAPYUqZ4Hb/uvMG/RofY9S7Dr6bPmMP4hJUs7s
xUw0wqVKTOaJ/BJTNINFRJFizAI7cr6e29rLlB2d8rehByNRHeRekmPVU+NM
G0o2h0C1GPEzyeXOo7wuiCU4gK20hlICyNFJC1sVPHu7IFCNZ0UQ0hz/ByAi
ZojlOIqxQ+Q00Q4MZvO1davMvMNxvbnQ0hAzIb34r77Fh7hLHpeY8S7ffeIk
QzmJGLetRvvJ6BlCVr9mE7QM8OQCNf003Vnw0NY2fjrgm89EDp+OOL3KUTEn
d51u3ALvGv5Ez04JO7MU47ZH7rkdp5S9DaZgm4vEKj2ndUr5KgItbyCo+LsH
c6a7AtPI2cclYVVM46YPBTqF32/vtCHPWtMiTsjRTbveefQeX5MTKebbNnIA
QP0go02PGSSe1XuWkS+bhWFqZCJwuHaLTy0FmA8jv01cqFGNFFr6ja7wEfoM
ydP30hX8TM8koPZif6rAP63XK+cU+7OjoeMbYWqKulaHNpdBJ7Kl71DKn6kf
PrpXrydMFpvEEAdH5PQcz10FeXObhJ/gkUN8X2FT1Z9UgJCd+G+wQ4+oONRB
FBK2FaQUlqSUXRM6r5ZdZ8i/ZJ7a8EjUXc/+nj6sBR9RAmS3P3s7PYT+LKET
S7aUg8ankrdYoVVP6TRb4MKuixQb+OR8MxfXjcCpuHIr6qSYE2xtWgX4Li7b
7f+bdSoCXtX4vblHsq8oP4DPSnCnPDOKV8KFfuw4PjXRaABfFfxSmp3w4EGZ
++yJK6SMvMoCeKzSXnibf7hCNA2EJYOHICDb5Phxb4+WHqEHqAVFqU+TK6VA
t8xKWerPxlth6iLDdzfeJXduwUuVxLX/YEf7N7sUpvAePo3nyAUJosz9+GxP
KMwALGbefg5vtS09zTDaIzDd82aAGsKCpUfru3Oxr9af8XjvuVmE94qtW8hK
1kNVn+gqahuhNRvxpRpAWIHfuQpkhbYIct+vIek2TryQEIJy7jOfSDLWnEjY
qrJgUKZIuQKFzFS8JP8IRbkLq8H5JT1LsWlu7YHHaaUDS0p3KNWJTCJUy4iZ
IIRoTYdIOkx2ddQzg2kKnp8ElqO2QJcb91a645JW7ZyQjbqTQRLN3Q9+D4QR
qsVzrqxF751JtJ4U0sFU2o6ywb7lyOROS9x/yNRi/2yQqv1gOE/pVTIaFY8Z
6tSOYoD8A0d+ygQasURzCfRPkEBV3fTYUjaDnJOQSYq7CzsMGt2+Wngd/zcn
VMyuM4Axrjcg3YaGqaDowOLRbvj+xnQjjIJc7trWa74FHNOkLZC79DSyPoP+
AvJddXH/oNR2VVL4+GjPibHHpWb+2hYvU3tin6cCdhrfx0cyANvhDHoHzbuD
lHMY0I1SzdvKx4k6pDg/qE7LTA7k9x+3a1w2ANZrFVHE3pNHj2uzvaCk5ErV
2rr/SvL+X5o9iykYu45Ar1hgRbIqj3RsgrZGNDGOr42kmj8g9z6WIvRDnsNk
gqjHhAbGcMO3b4wVsrdZ+TnzBxHwPo0IChRPFO5Vkjgl1+nUK9i8GHDeRrMj
0W0k4k5rgCWCXuElolvl85h11c6i93QL6M1ToZtIDG1Zsb0rlceUgVYCME7T
vqqe2apIUnjPGhRtmHs0ylAv4QU7KbL/YRq9FF2lm7QLMEPgmLG8S7JK5ozb
MtrljVWrB/p7oYYS+NRSmd45Fhxx0zQuF56v9zJ4M3ni9TU8P3GzrUY7QHL2
nxQTJBDkkSnh05HYWvMJVI2S8pr+a6ASd9x96Dao3qMRVgfgb6SXfRA0+qe1
mC4C/5DHjkVsNcuCo48L0ty8gNbd2VVg5DC1Rj70tQgi2ZVyXZCBtg+hzqCM
UkpA7CmZ0BiSPmu55lfc8AmTTwyqqFI6F57XSjRlrUi7HAC2sKY2VAiMr5XD
2xUT1cv+WSZDcSIVGro07N74RRCYLAbqJ5xFa9tccINU1U/u7EgmV+d7/Z/P
knYdeQzz/fLSiUyZQ0ruMl71tbDQYxacb7+Ji7R6M2GINUMTr21176i0R6Gt
fXqQRVVMNY+r9nQ8jLZLcW4TTzgSFmCvFXycb9YwROGguDyM6DLJ69XNFJ8W
sb80vS3oASXpsQTCIJD5nq52X7KvZDrh4kUzCl0CCmiTo9lpZ/2Ro8llZHNk
jjfXHqABaUC+2rINy9lDmWlTjJL/Zs9dQ2Adr9L93Gr0XyxVGnLw+CudwDQk
PcomekRSUum+YN/6+ZoJ0OGSPsJ4C1OGqnRNLj1hJvI7ArGMLt0qtwNUDvtX
Wh2x6bNwDBACfuE8lhDJXX40OOSvPK8+9qvr/8EChrWWk+FuoZGGX9u2JcYM
N9a0VJca7rDjrxBTFizu1LFp6IjMmTVcIIdU7oW30eiPK2ROOSqydMn+aqmD
C5/Lt+jqBwRTh/1geJGzpyanGbH90og1aBlJwH6tG4uUfMRx3uh5OvdYNBwU
qIcZYD9Yg8P8oXxcxOgUljWdAwFAwdg87GXj2kU97hQduGSzoyXed5oyVNkP
oiZU9Su4sg9fBcxvH5POyGFo2S9Y915U7jCcjYhfDSpS/N61tP6vjoDhIe2Y
x/8SS/K5LZvS9ZGWUYNDuX82N9t+E7xlf4we9kVGFvgFkMM+Gj/yqbTInAjA
sN+/uvSPl9YA+hIihkfa6tO0f/y6AdWDjcYYt0+ooroCPdtxKTS4DQ8c8v+n
zgRss+EEg0Qc2Ez2fsZDB9p+julvwvSvWblnCfOgbTouzimca6r7VsQK7gYq
S1gRNSiunOOQwA8T3bMVGyBi6Efr8hOYfzfRlM4f9flisTxhj/XV0zbd19/R
6MXLZ/xRf85qOrRlkjPNFC9fD1BrjytLe6U0UkvsKxw5+QLMfZwliveAq/rB
5Ml1G2e+AkKgZz4fu2LMtGs4fOX4/iIIP4ikVJABJFA0aH1hSL2A+EHqEwuh
P/QY2uvrbCYJrjkaQFRGKy1FkEMHhBoZ2pOH+9ViQHQEYHCODKWAwmQUVxGf
eUE8kOdteowcEs039UdVgNseEc7qtgFxO8B34l44oWCYsBGnSXiIhu2/RvBu
l/FG168dkNcXMkLDJwVm0httAIHIgDer8T9dlM7vEJE1Yi3xmxuaIZjWwLx1
umFqc8B/WVqxa3hfvmDP1iuHOC0Wi7YEJrR3idTqrCAWKEQ3U1tgB9ivFbNk
vHqeTwur0zm5UtmdpshgaYPodwWOqk+mHz7tHWaEE/cfdviUTfknGAMLhalg
L6WWZz/0rniEXOsuPOewV3vicphbeaNY22w3L0bSapK3HV0ekpuq1WtVVUUP
zv6GFaRDWyyh4q7dmOGzKaHAKjLcoOAYyvmKoHo+IW9dZpKPiHe/R/pyIcKC
renJF3ocqVYe2KFy2IQqeTnM7HjijruSkyEJgOI7YSMlsIUlEysD3C6pH1Qw
GC0BaXMDFp2YFEYaPISY0xJk39LQqVFPTDSsl50/5gyPt8YxOsuIPkNnqMDF
sxjXAfOHIst8XyfqIScaqhyjJbkcq3H4jJBnPWVzGTEzfIPx4aeW7TnXefVf
eE0Vyp+InMsMV/wHf93EGsQ4mAEKBFTgBHqoI++n4fwg1AkqnBMuSLMPkV+O
MSJQGpUIubNdPrFiRtLXOaUrDO8p96IHHCYfqHrPqmdZpYjjxy6RoHh8Sdmd
0wrrecBEVta9ANn6Pc5z24oGSrix+Uv4LMjF29aJtTSJY4KRIyVQvSYaLC8x
AqrJ4us/VioYEGDxwqLqeP9emcV2z3NCrUBxTkWL5WV5zS7aZ+MYVgb4ag3X
OPSuIYQKPsu1j/HsauvCfsSOXHyd6zaXesQHxs7yixuAtwjK0eDJcEdWXoM/
/n0OkUX92Hn+sIK/3jf3J9xEeO8tD8ljn3CrqW36ZxP3nAMDFA3c1/5b+qkR
RyZYpMokcA4cp5xhLoMSibokY3+RPdG51yCjhpR9uBKHZ51aVMDJMUc45ev0
ZaSHtKV1s147Wrf2qHpOFM4xbA1WH0RkYQJfJ5Cn/g/PBm+0FFwIGKPJ/IwL
6ZQf6GXmBlmcnlygYrAs+QhcL0ZuRUtVVhe07cHFGyKPUMb/Lpba6TVYC9/I
slA/D/Z47wC4IXLLVJEd2X3YOb2SjXxn4Yl0Q4V5T4HOg1ojE4BeGk+5CU+u
W89JFSB10M6TmF+pU4yVizc+MxwVczwNrHBMd9OB6GSZkhOTLlC3jiuNPAU+
hxXHOaIq9XfkSLH0rJeSUS4djAAkC2R4kRYm55QrdaviI54QV0qJ3XoF8NF1
7c5PS83EZUluaCyOUtkLpr277DtCWOM32pXjA6gtMqrZtfKp3ltjl1mM1ZLn
72HHXChlnN9HishbYAeExmMsH5+UwtWkGD/i1/N7SYYBDlRtPi1AgaHSPYqE
yRNJDdVDww8WGaALxmdQsB2Xjje/3suZstG38tHDuyRUHrT7AgZ5FZLOZstS
yTdVfJjvre+/J22bFXytZPcU7S8Vyur5y3jKZhBhwGWQJhJD5+zApbgOIo+0
OFvXd9swaGMXnfAIYUnxRj4OinAJisnisda+750n5qX60rvXUW25Ry6kM6gI
D2z04SaYx8fJo8djicftOtHBaj9FleOa0U4lAXsZpa1eDRX9Q6FanQpt5rQC
UxQjncTDWbA+JIQ7ZGxolQwZGudjzJeIcSU8cpbXI7nM+HhsCwOFli11Zi14
iGXoRueRzsUBj7qUy7nV9xyHI2XpkpF568qC0zPJkCi7+8IAQW63vP+MkrX8
GM0mbM+VldmZYndfu2zQvVLZKq2CYlU6zxDlXiz5C3y5w4RmP/Y1e6jC8NoG
fBbwEkATg3bPbxI82o1B3AW+HbHJDTLSJY7RxiMTlLvDpED70pWgEudRvNfT
DGOczTOsTiO3d1Al6rc/gInHiOSJN9iqefhery2P4EP48xzywZ+FxcQIBVPv
PksT1yCmu7u5fTD1E+938XM+oA9yOqapFC0N6n/bQ1CFPofuMDq5xp+SN85d
OIQHayaerLxz+zus/GxS5XhtrVnLn1fOR0/dMtjX3yhq1pz60TU0zW3k5xub
aGTRDNLAZ7Fw8BLycNhb4H0RsOK0oKA7ViwLhLdWSeYwzfQfjelShUUaS2a0
jdHU3+BQEboJjsWc6yqbiOXfmnGkBVe2b3CEGCpyq0ZgNwyu9aXB3rmYyr7l
FzUx64OjtP0H0tyNC87zsdRFy1wmSKErwsw0v7TkiT9lMSfkLAP3egef8z7N
BszG+PtG99kPl7YtobB0Q7/KrX4W+uIQee86kUgPkAhB+eyBxUVJjn4YOrek
9aewc9VR8PxvkDA2drFt6rbFmY0+5I1aRPVsIumh2io71TM5t6eXkGJX1kxr
Uu1GWY1z3DOUUZbJbGdcfI0BcmPJfFmVUrOwggisloVVzWal6W+HnfuDoNzF
nSLP8nM4Mrs3Alktctgrx6lmp3fwkYysoKVFK2aSNSof3Tz/0p2FejUXbQjs
a99IWrSawMJo2ZM/+iGiAfebV5/G21qNxeHvlrAM1hRh6BaaB481jbWeazVM
d7W6o6/NQCGp4Jr4jpx8UIbFts5d3GMo4YJH9Dym9sBsHbAJ76EzemhMEGQA
y+9b2y/EIehlHZ2IBvt9hZpNHD2TUu79mROjkH2Ob/yML1u3MicafQaxbH7f
ppWm0T4I3l/cOkXVlwcqPGG8O42/W0VdTdZPmA7bJzczrSM/UsxpNrvOId68
Ok7CN5eN2b/tqMERVNw2gI6GWZKQvPcXH8uLSGmMw0K6rbTk02A9rRiRxaWe
y1kKB3QFX4aiR5jxOKTuohWuwVZhjzyV1waCxdVmGaFUG8y8UDbeE6qH2wF1
VC4agqttlPjS5Un5pNdf1AKh7v6PdgDcpUDTHgRLd70K5AoM1hv4ETQhylun
n5mj19DnEp+Bzetcd8whdmtppuzcy9e8TcyKVD7yMEARuAecnSilwAnS/PDF
honKpL4jwjqsie/cz9lsu6qax76dPKeyWoWdgdgfUvkc+Bdp3dsmJaepDtfp
+FZojr1AGdPgHSQDdgzzXwPXzUmu2WJh34XeOC2PIJgKM/natKrI1MZyeIyJ
IGHmKI67/KT4dxIoMROzeXe/6MKTVbiuLAFE0ya6OOHzmmbqSmwrNn9PMkpp
CqRCBXoK5s3D5dFRY8KL2sCnOW4D1Gy5CSvuzW/vX+Wepx7aVu0pDljwH/1U
6x/NMOeV0LXKX+mJEosGBnlJqqqfOO75RH+gYTROzGo3HuUFUQ8wDK90YENj
AeuyBAaqQZu/L3aj40iGdK74E1qSU8lsHuU3OaCmhs/x3H0v9KO/1AiOI5MK
VPr/JQxpiZt+s/U/t4ITCuhnFh7w+HN5snKgayYS0jaDv/XX30FsToz2Gwsw
mkVJy1LJG5SfzMD9Y5dgeD/do6tDbB4HciPylhUjxS/gESEZvAa/CGWyRwpm
gU8xJ+7gsOQa+qCz3eyklg471fGYa9c8Kq021ei3VNGyJfhs5+q4obA88xr9
6ibC4JWQXz90iOm9bnzMAnBtHK5NynltpUaFtHwdQArR4O5syJG9xabIeCy+
3+oF5L17b+crygT71/kuAK4sNBw0h46w1FPXvpDtqNJyHRbmKJv9ggOF2czP
mp20PCTdCV1n/TGgsXJBAmuHCJ64BZZ3M9uWht37Clhya/BbxRWhbzPt4HOF
mTry11ZAMh+tmJIbnWXwom/zn2Gy4mwAjE0uGl2MoXUm4B8JX4ZoyB+wpwJQ
JgQvXryBpJLVwPDObQIKPeCCozMlWcWrQa3R7gm1DNyjfOWRP9tXbtAwDJGx
hvrONSPayHXEcYKTziCt7x3RiGikJHqq4+NqG3kV6qaL3kyl+rmthOS+KbiK
nEiFkM4vpUTsDOm4cb3QSZ3vJDrgqCPiDqSox0kTCLMi8Z22W8pE5l3PsNxF
1a2/JWJbm9D9sW+zEsz7x8sLwrgJx705fZtbbrJSP3mKUXrWhK9L3ZIqV7kk
eR1fUxwzrvc5Lt0ybMuN3BvApbfgwEH7uCo/eNuIVZcgzIgkHS3fSYIY0Cgr
R4xgE2MPZhXv/co1e0eDAV5Zps7N/St/Xiis9aYuyl9fKsolJB7VJ4Md7o1F
LPA6h6+q9VI3+BSoVdm0MXall2rxuBcnjsQhgp9zPIGfN5qbLw8pGTrtfqDa
5qwGQjcF8oYewCAHf7rSfuaq1viAh3RcJdYiEOo2f8UIpm4qBlP/Q9cJhBA3
zsPq3vnr/VyU/n41fOECgwnmRQTRkQeU9AH2QZ2fXfPAG23z3GEz3hWcFX1L
9PwiIy6r7hcdwRJs6l2GawBquQNwW25DO11/QZQ6X6eEUm6ce79OUILP55/Q
Ov7tSJ3q/QPZRq63Xbdj9j/Weikg22UHpMLQAo4WbkTIzTRcuc9V9dS23Qdl
M05xjc9+bUT8+DYvY9fS3GKjCTYkntzzRp08eEnaJW2JwH2krkRKf8O4RUta
zbatJaAIAnlOoU+5Oyi7keciE5I7SGfoIRXVx1n+JC2WTdmvviiqcCMDk6Je
21r9L5kbMTfRzAg+uu2D2H+P9PorAMnumabKxibpWy3JZeHqGwYiKuR29a1v
ZYq79gptIbGIhhISedzXFNv8OVLS4sv8YT2JTBnUgVPOCn0itI5Oj2csDQwI
B7aASZlzbcMY4oye11LAwNzRapm6OHt2QGjMiep9/3ccHzRKjgmNYEUQ6uoY
MSA1dtRxi6KXnXXPswRi6jG6cIhWuQFHcpTQLKDKM+mow6zfu7YMqBpunNLV
c7oG6ghhVCnjFD/tajI3FPuGYB4U9aS2NSBCblB5xSjbLpIsCTPgt+aED/Lo
DsWU9tg/W5cQHC929kJuXcNFvNy3SGxo5AvqgNuvfqHReUJmTkP5sZ6aB5BY
jAKDhy7eyernyoIJrbb1Mruo6Po4JGZlf2YxbB89VANf7QWQVsEtTOOoSGDI
pn5UHN0IiYqu9v6kvavgnvcbWGZrdPbtr3XxvMT0JlzbVmR6jTm8vhlVnL+k
FLdVHZppBleVYfCnMRjrzZNKC6jVHmRfFuaesyrk36g/Vt2ywHmINcvf0CIK
KlrWEuOnfdOPUJsAmz1jZGEmIO+DVOI2mn7jZrQQX6CwV8HZNHkVO/Ros6YI
DJKd/IfEtF7Klv+HD1x8OSsoQyTSnl8QW8MS74dA7bEGZGVYA8JgQSYetwj0
XrcRkjPzVvBrJlhQbaTwLZ2q0a8vn1TTnOZniwsqzWKNxk9nIdTz83W090zd
QZ4agK0YmEnBNWngUsniJsUSgMMYjnb18M2WL2NvXxN7p2N8VDKuJyULBAJS
R2VXPtcFwt4m+xhH+ogWSpU7IRFc6frgy0eY0o68/vV5x4L+2bKzuLqYxy7g
viAvCKzy3rnm8K1RzRbwqVka8EMtz2mHEQFWj9Cyan+6kL+HThrob3NrKr5U
3e7o4/8KSJR89QU7Gled+cil/o4etpb09cfb8InfTwluO0SFnkH8SS20zQ2u
7XA2fUyyIBo8TeJ1YpCrAUn/poP8KWJGHLPchm0CYLGbTI/skN4E/tjYv8r8
EicNsU7SnucNwxlDsFUCXoSi6lTEWvo0jbk1WXrTKPddDfMdi2xskMgO00Qv
BiahCFPEZS8ipEVV4ffNZH0nUnfZurt/f7MztQ07NO6mcPKfvHijBimr5QNj
FGkWTLCZ+6s/X7gZtteyKyqDuR/U3FES4aNvKU1d6WfG6NIBx3kOmSD+jVUN
RJAzZHrDliIVThgw17PAv2GRaTInipqjL8rP8M8Ry7FmQfGfNfn2CyOMbn3l
ijFTZcyKW57+/t1ZvTxusrOCq6EXDwEakFSrc8SVaGJ22ICXzTPFrXwQsSpB
U5+9KAPDqIgjcLIMHB+fwAjXzl/mCdFJW2op5kCzpcQhMHFNFLHJwofPgc1G
zgf65sAE3cxx+nbiTb/bNMHGB37Sze3DTiOTr8U0SZCTeGrSSvdNng4aM6SC
ElZbJAnhALU1wk+Q2RgXcr3brdAFBvYA1XwrVpzxFFE90RIQ1bL6LuFUWZBa
pL1159tnoqPgTBWEwZhklOrMtttS78gutNBr20wMb77AbIOvS60NwcIGoGVo
cqHQjqGcjeoY4xvD/0suTGTiMgTyCgh0MNQw2MQkDO7wkkF9Wh0fiEvWe3LP
wwIURVaIt3uAOp+GLESmoQIIMoR/JrmmUCzhSX4BX7FhVF/u4DwvJh/lPNgv
nvD8ZKGRsALtIci5b6KYkdwVAxnQoWiz958HF0F25PwCQQgZlQZkdxB/fJf9
I6OSW9BwLc9whRwDzgd9PofCa0oSBdjajEILB41r/FkFCm0+jfH9EuCi8cB2
Ki0EJTRsd7tErEcz50IMtK7NHC5I/ojSKPQe4tHpQqFLYJLGabmMinrw4vdZ
r7nz7C+E4TGQ/Z1miUo8WjI3GKdBWjaFmJUyLxwh2LuNLCUKS0bqbuzRYKyh
ybnIVbQYJi8aOnDQOSNKEj4ldvMmQq5+l0ebTB0AkGMRy1kTKPbEGbNtYNRd
zzlHHJ+A3fDs9nXfjuMH7p8n//rZGBkPktzO6wjHXNqE6rC2oViYHcmUnbqG
RBw4bf61gAr5mbGlHWw2biQumAxydIWzxrCOpVFNe5xZQGguA6+N1lFzqxKH
OFaEDbZdXQqzu7il9ho+cLq7v+Dj30ldxdl0ZIFNIkBNPIArJ69Muvfh6bCK
wIygF+CEIMo0IZj2xn/xye//9/y7KPemhqZor+XYqYKoZeThgf34zu5NY/Ys
VNduVOlRKWPEUBaXpceNnp00dGmL9FlhLvc8RKzaj/kORBA8VT6L+xRX3fb8
utodZiSYcydbiPByD4qLSo3nrgv6WZEmNNDCmDPHiUYVNSSguRVvwZLK+JVA
cdIikKrhCJIOUjPTgYUlKvsFcglOt3Gd/CUdLbVjQnyPVHTRFoMFLR8M8GZ/
+E+jBBMvgkVtX/TqMkIsXlRZPCUleBbDJPGqnnx6QZTmYg55SlkjyoDcbUKh
LfAV1o69nQ8aTTdsXbADpC6BqUKbHQb7YDooY16slaQUqmKKEkEkqsyh/eEF
QfFVVa/FE2uRkjoy9IH7xIfwO+L5+vSpFo2MxavC3J3eYCXyFzWrnfQoOTG8
LvcGupAMqgiJIZwMJgCi6OrFQ/EExAO1eSE2AQXmm66PjfEbM5R+IZu6VVdV
HVpFlPgJ2XGqQofJh8OKBuQjH4REV1yGzbRaLMGuk441Ze1GcycaHVD4AkZi
5gKDEDPzsdjDx97XB+3QaLIyoC8YXIUb92Wu0qfN3Orv8ZiYXlccP8XVgj7d
7uwtrdY3YDU5nsKaVDoKNJo3ojApSuK68zwnSUdTo15A8uSgCsyPn/FjA9nN
8rvBu8HRFFtDDHH7Gyn1myT6ZAkHtamRzHBfVHPG5DN/lzCUSjey9z8Vllk0
BrjhiFjs+ZU8QXfYqvrR+9vP+4u9SXp+MiExsZfM1hWSEghcCaGSCnA8hoKe
x0D/mSxf85BDlTIFvESuAFi/KnBu5JzPi3zvlD35FzVeR/x709dzYHx/dH7q
/zU9SKDO4Y9pspbP7+9JG0NUVpk7O3DOiQcW+kDp/ucijow9flJulS2gLc7k
4y87jLhbqAG6GGtI9aE6QQPTMtOtDK32wzjfjiyb0nT2jJNVHRzMHBb0aINT
5UoqH25Mdg9gfV42SthJkPvj0JX3lQM2NXmIzhjJS3VCJUuDYl/v4v/UdXWw
+H3QA5x89RRpLc1KtITBSmAwsconD43e0CvsRB/s28NIvFRsypoLRYykpTqT
Pu518i9UrF3clImDguzvMg2OaddFWJ4TCwhnGfdjGvBBUKJw7FUM6Y5BPE4r
V1hqJGe5muNuPQtE/dazqWkN9a5PrKWwwHTjN9t3W9Kwm49R9I0wl/QeCYql
1Cv8zIoPkZVQUJBMkVSC1L7PRgXPz/duLwqh0g8oJW843OKsghy+sZw9Jqld
ecVjBvBXx6x3i7oK8Q3PbMPVlSbMNoiUAwWdxomySjnDYLKL7bJkYGH6TChg
M5VTcP86Fglp9WCXNlcEO5P1/DQcKmqMAAXmcX/XJtBmedcU2GLs0TEjh//+
UCQ85UJ929a7h1xnxFtOFubLP9u2n3gQIfJoEYPIDkSMrP/nUwS/gaIUCB+u
elqgFZX/J8xbduI3mqhw0Xwj3OOCV8YMItIgDoGlODIaTgejrXmIVJxv6YuK
lAkJmHr/c3DGdq1/Xsxse9O2i8xwth/j/9REfc8Rq7/F016T9jokMInnQ6E2
7NF/ORisgcjMZszNX9VIUg2QDXx4jaMUU6pzkOKR/7VWC38pnY/Rozb+Jo0j
voWruVyEMXRWG1HG5NMTbVmIKOGjCMD6uaxzLABKoJbzpfSmHuUUIhA735ht
sJcur7BAEixFbawy5aLdc91lAr/ZAfEVx2sL6zwGpwcHEhcShReKibLihzWF
YXlK9t13sefNoxyHfZQiKd2giOzKUU63TLCjwuVYMuRzslIRJo+OnjCXYNMF
a2s43a8OT9u+qzZLc2t8lZNEQbkww7O7CwHynt9uR2GuM2pXyJwpw/obkyVx
ZtthP52aT8bk9ZkPNILA5FChjqz4NTifwWgzX/dxRa+DJqjEPwE8ihDntKlC
SwUQaDzKIfdX9JdWDAquWcRnS6GffUCwTpJOlC4XZ3+ge/nq6chq00KmhEcK
KX1t+SXBzjHXj3sEa7vGoCQDy52I6Y4gtaSmD7NmPdiqYZtsBXj7/X+I3+eA
BU0uBM02+XmUsah8wPQG34zYqtaueXOnTJqGQQBCxuhc575E/ZlncxpQ1Qxm
R5yO1zKwplip63r87fw86+nxqIMHlDekZgXZ6ZBNbFuwsPGORebqnzlA+49e
Dx+WRwccqyZXe4H82IvqsYgC13GVmug8ThuEhdUEnuEr9qb5Od65AlOiVUIB
0TGR43eOuv3Po37B1yTpyiLxkTl2vr3GMBVnkhDjw5dzjiRPDDkUamaOjWhm
ui+jIwrKZG6btZ1w7zTyiTo+9o5Ty13WYdvY2s6P4kmzhchaDV21Mwv651Ah
LNewNwL9Vc/oLcYP/sVOrwhWoJ4FBns2YXppDguF64Qyi4xpEpNaw5FEtkxZ
j9EwWPipoOMV3EX7sRm4uJNBn/60EdtjVJMwOvWdEdQHuWXGblj20A+jy8UB
fR27oij4q0i9QOzf67gAF+zhZ07jns4EK/ij8xtalVjm1DeQ0C+eeqho7H6L
B6Xw3HQApgheG+DijwWUxyolwHTu+amueqER+3uMM1A0ALUK0M0vQUj1w48i
nV012gZyxW0oA+wO+LU/Fzo+AuNSYLKpVQcx1oYkbkPDNtpEdUlA1CqpcttM
5lpEUYGrc4bCAznYeVW5KYxqfEOIY+p9hMeHzamue2O+s8IAjGdH+C0S9Y6l
NOKV4k3FUrGwud1AdTAKcEiP+ObMQ5zaY+m7eadEUy9WnzP4/V2EwNcz4eqg
57LK1OvQm7vfyvMIfyjXiIq1GpWV8TcZ9vz1dY1rbt55Yj8/Yedci/qjPMr2
VNNsx7mdrb4G//1b3lVqWAv4d7EI4ZdDww1Titx/BjGNMRKd+NYNra/0k/80
HCHFAa0JFDDrIBvZZMil8KTC7RTkujjLpdiniX0bb94t/ldAG+B9qMRT+zAu
CtuJq+8nM4ggC5PhmyRL7BgoRUxr0U5GS7OI39T0TDfFl/NJcN7rr0PGnehr
vuUvn6J7BAkZloVextH9Hbp7DIaxygw+Xyh0GA9sI/qI/SNJb6DM/D9KR8KX
bGh0x6asHAWlU5FfSm0SSgUYQ/7lZDBqaq+9d/rqNXpqIjlC/0Vkw1TBonmN
NcWzNkj0bi1Bo9AWwAieXapRwJ8/V3FIcQ2RSytrbddHNR49gkVJFt3NRxHc
jBPDy1RLdgCfCG4iT3W4SY4Mtw+xJ54ucBzCZnHAHvNqrt4nEToH0dCjd/fR
jr0ltUtyxOFZxrScdWST1n/cy/xSo5l8gHSqj1l8ByfP8P3+rJB0n+nEaV91
JaZQFaMviyPMdVzn2vq7+Y9LWiryYft7MnBBR0pOhxQn7stCwJlS+CxgOcin
m+Cdybj0UQRa4odAGjuoSzeWdeQoPqfwV7qv/UiAPPY1CzyJlFUMIArFu5cu
gEy3z6SHhtJPZgI0TPUj70ndGugjVztQT/0S8IiJrLxRwFYqqlptm7EOY6Zs
sJgB9V92eau45bNa9ZWB+RdRvcZc1ODKuZCSlhM1YzyFa30DPqlB6TdZgSF3
6yiG+kzmqy7aLG6ANmesXjeQ4ME9rzlviNB7zeLn/nb1JCEIe+lmRVXxF4d5
KihCdvr/j2XabhSwxqr3N0Vz4x6rZ7zGn3ShBmLCi59Z3IMwv5Znq2Jq2Yvk
f5Mcvh1meElhh1ztm5EmQXGN1O1jwQ4fjI79PxmEGITmGn4zlqKP01V/hyIA
KcZ5fjiUl94/RTaLun9iLsFcZyd2dizZ6M526bvCD9ln9EifL4kvUjQi1YV5
XI9cmQ2zij00tNS9aRVQPnmrx5egsluI1XmqC1kA+ZvIh1HZbx4+dVUR6wX4
AMuma0L2C7GX5iJfAKFwfEuWDNvBW4/5Ral3DCBlkqC3yYGb/Jz+lWi45zqJ
xIx+Be8FXQPa8vOokObK/3C5bSIM68xZzA0EHmJiuspBa5kyrX+qMl0k6lqp
JcQrQoK++QAfQHKyuKUTjd81xu0OPdJePYAkplusFjb6BoUiTfTZbQcPMRZK
0V//4mE11QOSi2+B+gQSSyu8j4mlF15C/6QB6VlkywnbXc8U0cBH/YTmcQph
MgpTZgMa31BmNme4gZBDv7mbaLf39/gYglCBs+YkcnSW7s9Rlml+G+4Upd0C
xh+CnpXuVDntYWpSqHwufYiXrKYR9tFBF4zrvM2XZvdv2lhlx1Yi2roEsvay
Ps09AC0xfgtjucurxp7bWxT6CD0s6CMEP5ViQcrqaRKHJjhfiCwmOgD1y3mS
Hri3RBBF0p24/CXZOplmXCPxnI7kgqMLZ8zT1NNlByJFYX6TR2y1PZYI2S9T
9qbhxSggZs1mlch9MlIxxoz9Tmsa/AXOUyfiPeK1MuRhwN4D8kbSKFdgYlyx
o0ACOqp08Jb1UCITUuD2Yw9NMC8gVxE2NEfWAIvBecA29RHA4djbXbyErZ7s
2rCScS3JjqxFHg8aaKwg5nzADHOscR2fh5ImyYHkpSweSMhj5hy0O5DSTTKz
qv2KAo3xsyJ44jYWUIflAt/2prOi6awSCy5eQXKkIpsKMlYxxVKq/qKpOJlY
oyoNiY3BhsMhXSPQqYJIgZ3rxACCqh459LICnqG5nFvL1ys9+fIq1mf2mPyo
bH3m0zFQw+p9/X0pFwackJcSHNmSdxOW410lXIxobUVnkXhWXkXKKo69bf0z
QehijfNEehE5it3Up+akDOl+ILxQTJwnFhPiNPj6Sp5w9iZSmMlRJMoCV4ii
xlkdEsl79EWssHCO0U3MUWFms0v8Po+cQ0VxZsxx/9QAPhJIWMuaqxGn1RSf
+PuG0G+C2SQEz+mWDu+/XDYiun99kDzfDFlN6iyku7QPtARuIDoybnr+HvOl
TZ8dUX3A0AOEIpFzS4slgXAGM5nL74sLzBCmxg/iIp4MfNb34j2KPO8pUr7O
Y8Tc2aw+mUMrKhRAQ1NsYvWUc6Iec/s0QBRlTO0KpK5JeKuSZRckt5shic+X
aClfZIkRC+35tsZyvZqZH2Rc3x/iZse58zF12j4nYhSUN1WJ9+a8jGA+JQED
LbcxPocg7gMrsEXV1+epnBmvs7bEbqhFG+ILYu7gTNcRLFTNX747+LWxuAEY
+1MBN9jArhi1Pmk0O4BWf9quYCEEUHloutPb2PQTfYsJmqDrLWrr9xnAqLe/
dKVC9DCjWPF0btStWBjo0TmsPKU95FI3kCWMXN2qWjH9fxnMueNgdqrWOzQE
9wANPtrnlcXam+z+12hyi6qGXn0X5MsZJwH+dWzC4zuUf3i09psmz1iHby2m
4H3KQ4ArSXzVRVajlE2vqLGyOcC9ePuLfQ1LDSnXEUV+YpvQdEc8mQYu6eLG
Bmka8Q2FCPxwxbIAnq2uxFqijp4GMfmsJ0N1DMYAG5vOwID6D2Ppwe87J25F
rH7sWuN6b4EuVZFQEOoNQodQIKx/yBT7L252gdkN/em6TDd7bBu0weh/jI7q
EIqrVlSn47ss7smLR7FpiZoFYnOn8eQQHi4UluustR1QxW0zVA6FbqgQ7ObK
PB+j8eeniEtMRzhK3pt8Laod8NLM28h2gtU2gMmPyLbTQ4VlilCEbVe26ZHH
rfm4PpkssgQf/SvCnHncqiAtFkMy4ymjkGH11xRX2jGEgaYBm5GudSXEo4B8
euiSkamMYxYLjUfpXV3CrBUWKQyCf1M5s3AiF9hvgCa5M7ZgG9LDBONgRVVr
FFTBknBRT+Oy4Z1LRg1eeFRSOKLnvEb2MynLEWqEav3zOU8qhqwPpBtoup51
K6j1VlXfKWIoK8kgNnLIv69P87FtEdQTiI7F4qGFrUa/Y+TGZw4s9I814mkB
QfM58SdcqtFO0VUsyXqwzx5L6BKQJcR0gdyTCxwJkQaUxEwosW36jZ3uQRy6
tbDUPzYVlaEQsAXzE9gdFrr0Trbs3Zs/ufMfPHEOG18JINlqeQtIQAkRU0gh
Sp67OX9wpDZcsLOpP5B4X8otcAdxL1P3rp0OgnZOj1ZZObOq7+b1dYCZ4GwU
wBaWZNT70jBa5lSfk2GXyCxLA6RdCdU/7B7/5yCND95g89wd7hs1em3cYGcf
Nai6tkDOSxjIZxHV9KKbTVA1rannfF+sTXwMNWKSobJXWbYxpYGK7+5lcwwd
WEAIAkxiE4phaNRQi0Sbs8tLu8OgWdrfKt5KAaq+8whhwdkJGRtAcILW+Eig
9L9T0zUaLcX8g3YyiTgwF/rMV0V72O9j46dLkfI2GkMOMJr7dW6WRWY+Nicq
6N0NKn4VQEpi2slaPXxpRnZYZyUt/SgfxJpyw9aP9EOM89xnJ+GFkXViuq8u
SAx5ctMw6O4FHxEcfrZEEgiI/GKzN0tN5o6NJfehr0tdCaZDZK/8ZoX8grX7
76R7xFLVyxp7oef5pKSuwoyPVLGbJjdSniIFHx09pduber6/xHyHpzBriIRf
aESeaiBddTQ8HyuMl5uRMpo3NtZ8O+IFsQlfNRjX53VRD24FI/gNc5Z6NlRn
ZN+A8iqWQ2/cc+W99w0N/dEpHOB7HXoPLlH6rP9Vu4FYKTxSS6mf4eya0yMY
AuHWg9iimLWaSIdzcuBtr8qlM2MAOjsFuL4DDt30WJ/2z6B1PREnPihs3hBj
w0gmsQ3TYsPqWVSs4uDCRqJw1Ol5vdNCNNZIaFA14Sr8jX8x6mBv673Pugvd
xxT1dJgQUr6COEAB6YjKGcFlIc/n7I6IzZ6pKl3C/3sH7zcb/IiGJTpy9AkI
wqJvys7thPUzRvFq11ZTAdW3rutyVldzVtLHcSQMKhZcF9h5utV7l612Q6yj
IrNY4vRiyoVRiLs8t43gnYEjlmNr1w79Xuk1qgZdiHcdeeahf0Z/5Yi7+hMh
nXxJ5WbASaJYLKPtRTlc1seDEDRe01WgiRux4fu/iG6SKH2t95h9g2lyfHzL
MLYczGY0Jrz+2mzCzvc3ou96yoyZvC4xxq23nxM2k0YmpHhEj2hzgdqYb1v/
sIGfCsT7VYZG7M9OZtJeDLIlsEUuQK1Dm3MHLVEuFKTtZRtWfRQ/whZFjHO9
tV5ddapVCS6RRjj3nsNWF1WLPzKX8HxR7d1Mcj7qTfJssH5TkoMGln+lH7yi
v/ih62kaZ8fEHvc+FRRvyUfdXP5a/FrXgFA6ARbYMHKR89g1DtJU6QWDb+oW
/toLlxoPou1kv3hxRN/UFXenoy+AipBvWfdGj+xQrYkfJJbdnqDpi1CTIdwv
JCEE6agNDwZyka3NmIxRi90Hxfslg3Ws+gFa3ybVLq65w2cIMjF0X3GFxvfo
SKMYCQDKuaQnNuB0g8RzpVtEQ9MrX6JGoUw+cVBLwGU7GZDfEi1cmxirVglO
Z0zfHyc8Pf358RkK5ULvApSWn4yoc8vZQBF3yhCbVdDcQMPcg9KshxDHxVmO
JXw6pbUFdsOJ5lkPNuAruslEQ0AJQczUUj6rnPVW/Y+6LOR03Sqxhj200vfF
77YyySizabM5ojX2R9bPnEvXnLksQldZXl0NdI5tJaF+ApBZlVdofgznSCnO
0cngGlGsvrIH+hR5UPvfAP3u287dDHju716G9McRp3yl8OTwy2snH5OqjCpA
bStKeIHz1zJYRZ77XKu4JN6jSRWYZSvRmtLu3F4XGjXfBpe0rj4Ld18iNt58
wEx5DXycWKy8MKX6H4h6+5mBJobMK0cFLUdSbgEoXMiA+yIWcXUveTy412Ma
YKySjRjWwakXLEwIBEh+A8Z25tavAi1wtW28THLVuIntm+XU4JbSBIVM5J7y
uTri1ANqSoRoPjl/FiZz8zi2iFwY8HxnrYo3V1Id4INbN5JJuJvwzGYsi1I0
t+cBkPaYfSILK9iwucgBp9uCZtKl9H2U28bq8/LVhzj+ed0/f3i3VOv8oEs9
LxrY/587oIQ1B8BuGqS7xLZqibczX7POtBWup8o3405Pw39lGLKKlFAwGCPq
9On3/Jre1mIuEX1KlqCl6lDOxSWNyI2ur7xYTzcwdLgJwbNYSmH8OdDrq/Pg
Bp31VqXU9dD3boT0bn5Pz9uiPnN1YiKLxMkgEmgvEvkORykWqR6R9DF6Bxn/
0iBscrojF20OLE4falVhHX8ABl0yl2oqoSg51muU6yJjSu5JXy2ta3QDTlr9
CZM0pq2QPbv99opx/8cDfa/q8Y4NM9FUdS7WDxdgMg40uFpihZJyWF9nMmly
Ojg8tpBfaUSBaw9JQWumfb/85dFMo+tUkn8Uat/dQN6HGgNht4wZxiOxQhWX
Ecv9nuzzRnwsP3huMvY5B7NIlCNLPqoFzYbF/wi5+FJkZtKa0PMkhKsqTA/w
VkzTcqVE5KiaXc2OO5p/hwIC+jgfpiJWSb3Y3MdXsryq6jBMtsIHvXfXhGRH
x5whpliuNLpYrQ076gDDTsWBcBCuHBJ4L7yeWGSF6WlHs2c8fZw90u9YG9wm
eAkd0PARApK7oD7eUiOjcJzAC5d3agj1kT8BoDOl911qMLkVqKp3lGJhpncO
uX+kgnia+O7ML0+upYEAeTY25t4TMdWQzLcJNLDuXrJdYdOVCFw9d15P3v/3
yv3iIeRbxVBaNVHcdCiCEINwazmZLcXqd8IyAV85v9jijS1pQXDGafwaDPUL
4xK7hg3FctYTv8a6EEUi1+SZIQOpF0PBv26namf8kp0Xi7Hg/mv6hGLNUsil
BQLWXDafpw7CxMpMyH888P9wDrfjb2n7QB+OWBwaFeOLZeBBXv/ZzNb0s4cV
MK1WQOIa9vGBqUdZMEw1yDbCJkfDXjTGbfKEj77POYUMZ1KSKxNCLT+kHVz6
hq79cn8kokAYqEXz7hv+f9v2bp8dBUzLJMjp6IXDMLqetbOMrCAeO2GHWfCf
MdWFsMU99nmOjqXzZsQGG+DAQgFRJ4KloxeKTNxIH1n6jwbQx0ZZYoYc5s5a
PBtbiS/iryY7INMpDr+Im7HVva7nyVWB8Z636nq76U+jm6XBnLRER1wDXMta
sIJmXmxRRA88iEPMQoVmLzyaaQha+3JfI9X4PaMGCNWgaX+lbsvBhww+y4q/
H85MBmi3qP/XSGwOiTxFNdVDlGDn+Y4eo56cxf2+c2DdS16Dz79klgW6kqsM
rwOZg7kq49uEIfhme+mjgRNJU5DbTq3FOKaUWfK0/NYlsJmVCpTewcfDrkov
SBwQALo0HXXucNB3z4PCzBe8jmZU1HaaQ0Uj+q5pEWcP6rOGehCH8GnnXG0U
FcyT3E3nKt2Y1BOfu3DVCpKZCvX1E7WVG1qPeDD3g8hd7QMXAf+PVsiO+Inl
uzoV2LtuTkhh92+TQ8uiN+euXjXAUwMU44JwmHBpkUtpTqnVdetAfECfDbqw
Sbq7/ql3dzFaSd4a1kemjawn0u++RM88b4SLAtnH6PzLa2LfY8gqKCmn0DQu
d2kZyGVb5gHlDaypb1SqpHF3WBWm5MgWJLUQ20ekbjy0spDKCfRwtrsJ6QwH
w7/zp89Gfq9ja8POvc5TVYOjLb6HTtetIjNX/K6geQnQlFNjQAsDqRA7l+fl
vkZsI+R44D5wFB5HJWFt42l3QwJADKq7ENATnbQ58T5sjgsBQkJoAeXhRmR8
5njZH4CRDjR+9s/eIQyoxDqxOZ1Osamo2iJswMR7U8xGcWLCKqEJxyqeddCI
dmHzVelLpWUogDkVR3Gt48mlME1k84Ft1u7OuPGDtqvlM+gDUzBv1M7yp0hK
VDHZcpc1lebfOlr2hLIeUjXP/p34sucwK6rtDk+NSe5ecU3hCjFQ8AyMVKl4
3DBwdudnGELevVj76Lma+tjRXCinayDDotQ1j746EmVWHqjwjjjTIGcXmto5
I2CxcUa5gQVKhgnGZxGttXqR3ssMSoqYG32h6tX0/GueAPHvbPh/NekEUdSB
UG8SR1wdYNi7mkhAaWf8JE4Y204lQUloQP6KIjkCdVnV7EoJISOGsO7UIRgO
fIXfP9Tbf4IDzJBxs0GXUuPysdfzyFrpqXelA84ssrHoBprz4ICO1hDEGK04
4sDor32m8wxJstHX2Ejcl0HnUnztoPE1Q1w7jof4ShrKYqkFsFCSHQjW4tR1
Q7YsHAaPjHOToVkB3SuvfzEdotFx7oh1+4QMY6GU8AFSDkjXq8nPFHRnet5D
515NSgl7q2dTPkRZx2kS3c1A1h4+fp8GWkykfmCtPKeay6E4y75+kjYjs+g7
P4XS8DjEFjy0widZRlNFXoLpDjZWtjfhpFYcuZ4+GOjZQjgt3K24QHaDsvN1
VhQVuU9xgVNK/Marqdn4wWsXTTkYp+r9va9DPffNr5BpAidw9ftP3oU2UWAU
pwWFqG909XmaoxDu3d0lrm2Ch/XGp9iMyhBb6u2BmQ4pT9ry52h0J+Q5qW/b
G+lOfOEXZXNfn0AxfhxSyjVgoq4uKqX4VTZfcC7+uuV5B68G6YPr5X+PJMqG
jSUqVo2dQS7Q5GkYzIYn7B8n0qnKf/I+lFmZk5SPl4rEDCgf8NMJDilDQNgB
n/lp3bI4QP3daSlh/y5LkqGC4aJ/Fyo6H0AwyaEXWJu1wyDq+JA9teB1/7Kr
o1uTRN23q4DDKosbBg5t6DdOY33qIxpTeq46snrm1Cj/MJmVYWxSFvRCwQMg
FAFWPDnB6SyWQMGRKEFRyIqlj7PP5hr+CTSlJxBztdq7VQJLVO27icRv/KOH
a1UqYawKNc7HuQjYF49WMe3Fh/N7uvZQgNDlb0YblKBuhQMdXkqyQabPfAgk
kH4zED7PIEjoBkeccT9m2zbv1CaG5Nq28hgWxXEfoRyYoqP7Q1OL5TT0BHNl
iXPwJHgG8tybUD5aoqsifAgdezk21GZeCb0dD2XMbX/D+D5nu3K9CdMOx13c
DfV+iNTwgzRvgDjf0kTn8JKKDe4h/RnsMCB98H1zaAfyQEy00etKAGezVajs
MPFq2NrINokLw4SlahG0zCHeOrLCtKgWEmqBZthUWCvhtZ4QgZAzXJuh31B0
UmICMQGYbN7UsbfJzFKh7SDR5515P/k+qEd/3goKAcvLTw+A6yW1NBw4XT/t
ItUeWtN4pjslLFizlBBGHJ+9AZIMzuAP35n2U2zg+wbo8+UOPXCqUU0wJMQx
k1tNvfyg0nT2uqffgC0Pr+IDLKJ8mMbBiwZDr0ymwpQh8xik1DL0HgUwphxp
ISZ9gvOXi5ghvrQJkcxWMri/boFh3lqWMFvx8aabb6Nd2Nw+mu7617ktFDuB
Cc+Tjx7BPAvLwCX2MLTipeiQcDgU3K98lxGp0tyvKblqZlSkN2aMmRlnvJvf
0eFVuyF57OSNaWnHcbraCG57AFPeoZONB5SHUiR7pJvm3rj2a1YF8lLZxGVB
DB8jD/+wSr2XQxnEbeQvOep/FV+pDzUrGHaVlllSy/uKOwCZ3kZDdwB9NB8M
wbfX336e8QoDh9/oGWGJTcWrwAeIeLrkZdYYR/wFZnTolpQ5Cbkk3Dn9ArCC
Y2w4dgZWAV1B6SxLi0SFYfGUBRWNuzkxPsO4neV8xK0s0hkDQhXuQ/QrH2Ew
cUPr7XdTyGx/gEUcr3JBsyaYgYH7TWNL3N7/9KeQTwgdlTM4Yc/t/g6KkHF6
LPM4HKDx3vPuoz4hElrQb8nmMz0OFn2I8b1KBGy4/eLhXTXJQfCx2ampG5a/
diG/7XqO4NpK6Q2EClKiXXh/FJM5ne0SAoEIP9loxog66BX2NnmuAJcx0Yde
XM8IG0B95WH+U1306hj967N/CxOMDP32yyeTMQ2Oq/rPzNVzB7MBOhljJo2I
wH/tkrBOLoELS9mov0pNoG9pYPjHUs5rjdm1SFeI3Vl/pgVF6ZKCAfIWFl5d
56uYUCODzAAVWtILlOZJWp155phFJz+QaaPKsZQCB0yFuJ+ETeHMCwc7IMLL
oy0RSwXCNUwdUQfvMJvoQyQR6xd541Kcp8CHt1tRfPZ6BYX0CatMqer2p8Mm
FugR2GEpwSwRtv9wWogQrxyaUh67V3ERxzNSBs2TcU591bhhKAYxZcs96C2N
ukE7AViOH+TvEqJYiyNeY4D7vAcnnrOW9VsPltyU/q0NL3PsIHmeJpp6e0VO
gCnX8D1NXMCy+JhlxZxY/BdWrYOsxaZIGYs/DNq/yYoy/Omy17nvASqYYiQU
bp1cdO6amuMThv5no1SnpmrgqCLyYc9OTIj3j7BI4j5E43iy1YsTRBuHpBuP
Rs7iFT2tEgtcI1m4xV39xvjXLqNrixxSpC8JbZBjM9yx/kzSZT6t/KCbo2i7
xMCamFNH5AtyCi9VGnw7IP2HXPfwXBGSM9KrxbqYM7W27+qLWtGx2eKxp1Dx
wgYEyj5tzRhaZv51+doLf/HPU8fRYHEAqNwC2oSTtr20sGv95bkC5S4+xd8M
33vn0YbteIyzMkyGKUaINWTTh84kKYocDQxXHwUXHyrUA2Sz+sV/xfrF1/hn
qNLovMO/NWPkKNBbZ9m4FEI9PDRqPdP0YE1EqcT5U95DVzdovIVaEnrMGMEE
N5+OiEC+Nj7q2txQclmkWGQUG6TIg2eqIPF64tauOxExgvhsYvwjBVJ218Lb
74k/gMF3Up+3q3Nf15lp0LskdbP+Qn6VGwdj36p7spcEuZoAT15zKob6lD+h
xM7K+9WtgOB4mWb7NcblqQnJ9uGGnY3wli/esLWoh1YNbj5HZQnECBT46cog
VMbYdVZGpuhawaH1hF36dLDst+w+JOTsm8R9JbeniKL5LWXHt7mqwG5gKT3G
+1iy0jENk9t17a6zIZFuemJ9G/fzs1nTzbXBusFKaYb0ECjHPj1zoloP+EIa
+wzF1ev+VgaaHL7GQKwBN03LFHGAuywT/VWFzT9lyylIjdGiXMaY0Nw5TKoT
ub0Nfe8kBbITgA+5tRItHeOQx3EXrKJxDi43T88bfXgNbs8LyTth6F7Lz7+V
aSeWl8PBwz/+FuQT8DSfzKkcNKa4hTjw6DDBzvchUhVMtXJQIDZTESmko4pW
XBwtQZQZ6Z6Yai5KMKCsN7vH3qMBja5xKmF0xChSnG3aDoWy7BvX2FY5VR7d
es9NED9q5AnhUyWSFH5RBLJ+D12U34IpepwLFrflM4JuWGUq0Ci6VZapDASs
3HmyEJJrFdQvVPDuBeqcZUPneHZYNVp0LzMV8Kw2+vz43nUvKM3x+ZdxrJSp
3TA3di67CVfDFlgyiXfapF1xWL721/DWxwSZkcQqz1JpUznrl8mu9U+H3oPe
wFhwnS5jyXL9J6ckLxZjnno9jXtwynhFuxWbyJWXOz6qHrkysmOz2OYrFe4t
F13/svsjbb1IgvyWjbtev0jejAVoDFCmDXUc7cVd4KHzjOGNPbAZ5sfmkHj7
g3JfFh/Sb5r/rLi0P4jy2sJkusW/j7m0CijkW08mSCq3dUoPOcPYJgYXshrx
QHgp9nP9fIBUpzOJH2WOx/efhHvS5CLo7H8+ZFmxeBVb7rh5Ey01FkfBFNzb
tEHxxzrAiOqj8sPpgiZEHl/ygaPiEuy54gDOoh7u4FvL2BEi5MXB1y7iF3MD
0ctEDhtzg5pN8VOeqeHwKpHSklNCOMS4UDIF/bkAHa4QZg3azgJFAdiHIOMp
S8+6jeubW6Noz6TmnEvSrSmT138sI+F84okKt24ujs4oyHGwKULBpch4UTs/
cyD0uzAWoMvLpW+pSefm51REIvWgPSQfKyPLyQsDhSRqP0DnE+gcyLWtsYv0
KZYQGGrPSL3Zrao8towsDba39Kck0XrJKDYOQfTy8WEE4CNOMx/vwVnOynE1
pJbbJJRs3XHhbs7RwpYZyN9LCP4dh+CE89H6iTwHTB8fz8ASUTconTWSIZC0
WTGuzFn1dmvQ7vqTOr1YkrhIZtv3/bp3LPRQgBYLcgAzboZelTe6Kvrb8F97
jBKUTAZKSXxfl1qYaPm4z/tUUTj/f+vD1wZ/VgDd1n3U/hGt6ZC8h7mj3CEj
x1wb/M+5dboM1DA8Xlt89qMw//HFC6HvFKeRGOzf8Ns1ucetLYkFQ1SfpHQ9
vXz51IGEzjTq8zSfvfaMXhutmhm/i6AEZmWTxOVS2lwnZlMtoDoEqx+nA0E0
hV4k49BhSAUvdgAx/J2j7sjFCzT7pBZLv8hU33VkVrUiDExXmwTeCQmGUY8o
xomYDL4d12OQVrRPYVdkJ9gxGm+LynXS4zf0eNcTFoemz6kA1b70s9VhNsQD
CS1E4Vkoq340l/fb/IXa2xjrDq5r6hOF5O1Vo0ZE/0ylUefQcbl+fBKLoemi
5DLy3kTkM4JlxsnM3aNwPZjRJXeLu96QH7vWVHK4J4/LarmyU+EwyOHJYZeT
WoETek6Rcmpv7VBDdCVkxrjcbzdfo7/dPrSJgUjf14RMjr2SwM9xFqAba9R2
Q3x+5GB+HDHHapFpXHPJaQK794Wqino4xL7IVDYrdpXMgV4E/n87Lg2Pefco
BuI+WgfEQbPipMyAhle3n3mflj6nsxc8Z2gWUHH2xwCKPUwl0ovjaQscaVPS
yjELVfK/gjRH8gwJkJHG55649yYhRp4NLrXxuoZW1UyNJK4zs2/rF8SXTHT/
M0Uz3ETqg43O1z9rS9y+dd1CmzEPgsPEN25LD3GtKgx2x25CtHKAVDP1KjYY
8nD4GlKzYImIKTGpwvFXgszPyS8MBLkE3HZnFvm2vJN5efzBmtDOX4NWlWAq
pugcBbYzZara9T7Cm9Dguast7qH+d4v1lGrOcOZKIKqc+jXbBWFkPepUNbrm
jSYLuhVN6siGiNGy/9isXPJw9g6M78QHYHFLevdho8dX9PrbuFu1tw/PCeal
7It78jnG4Qp5KqdjBnOPQ4OJzUXDVsJbhwl7gJpFf2/08YuN/pbuqzrhi9+A
vPsRPKm0mnFdi1NTKidoZE9Sk+O/DVubYJwbh4D66+QKFkhaubdljG2ZyNC5
Y3udqqAmoBb58MgvjJP7kHLW8tdHLxObaasZ+uKweKBIDm1zLGB2X4VgxY1+
s/R8Y15Z7eaVcGWJ1zacFc5pBpKI8uCNShNZp/5C7ueFiRb+bOpochDA9aMd
gSPuO332uWKFdNihpxvpwQMmw2GHo4Ixl7aIhntMVef756QDlxSOLeq6OZdh
7+DskXCfBVSwIZQY1LX0BslXihTNJDp1QJc4Ns3z+eUoZ9zv1KdTZuhbzLnh
b2b8arKPMRUtypHKydnjxF6kWQRmBTID64NYrzXOspzkRCoBjLjewCqAqdEB
Y5M1C4dpzqlXy3dmDP49lh5rOMR2P6TSb1Bk/j7R8YtZLUq6eOczpSAHc4SO
8+gJmDdddlXcIFHfoQuTP9hcEX3+I5Z9VcnLr5d+KhjrduHvoTplGiUClnlt
q6QGjAvXcGsbP/uzL26/DOUJkB4bmrQ7AQw5/pZx1FQpOU4EksV9Yk8Nf95s
lugO9d20QivodjCwTF8ALBWRSherozwiVQgx7CbZoLnrKZ4w11x5iqQ9yvAX
nvqGssxvXWCH+ckp07DoQJBjzLX/YXDf9kkU9PnTkSOfJfq9Odf0vFleaytH
kJvPhZSyz+TAO3eM+9d1Je/Ll5WkdTGdFgj997PGZjXyLl7YR2QtdSxIoR7g
oRwAR5avIP7wQ+XI9mwxWx1dKwJa3A9kCet3fPKJQoEG/GCAwMlfxdWPUEos
hen9JdQZbv9iqq0KL52XpL5gCK9Zw4bmkz8nwSAXvnY9BSi1I0zSKMCg5RP9
Fydv74cMxgIyZ0PvxlR2Wz8DXWOqKM89NSkdWpEH8O41K6qiqPu4ngO0uyRL
7KICBK8tUg8CURd8PHBquj+09taBvknb5QJRe+NkVnd2tYNrfXWWWV3+zGpc
v7ZEMMZjmWe1EgdRy0Xd5251XiBpLzLdVThK7WcuWvTHuNrQuq3fWNEB0a22
4A3qFKKwnofPQezVzBL2qV1i7vtCxIhExZHEsN3pvd4teZ8bZbJZRlwHXU6E
EiPhI8+TsVZoNE/CPu64rpQ7YgNKXbNaihr9lYYzdoc+yjERstK4FIIX/EFT
q+45xpe5yAvY5SMIQxv9e9ylGspIAa+fWhjzQvt1uXvQ0tp9BYEBDvzDzkHR
hhZFHtuJlyps0JBxF+b8JvHmIhvaHiZ67RK1qzD+1+BMSHRqCJhf7YAMUiKx
bco847eO2HwJ2Vsi7NAmDsgYYLmcef90MAxSC43ucTStY7nz8PMx+u2gB+Wn
IIbZER5TfMRqvkadLX4Kat8DwGuH77zRMfmm9IR1tTv3PaaxteQYTDckNvQ9
WJByyGpgl7tpd4Iy2FBUWuTrsSD0LN/UCwfArFRcuZZAQ+yTddBuxwh4ZCH+
8NaXLbHTYSXASBXyBn+/Db3YNeVRCXKWedUPeBsJQL5vOPk22YqbZKO9PqzO
HMPB7UForNb/yQbHoEWYHvI9GQOv6NOIyFj1YW8ook1N6Of3vHHdRXObqQKj
iFcZ0+KygLfGcqPhO22nV6fXh+ds4pB8fslYmh+K9xAU4F/58Qv+T+dK9vpc
NVMvmDFYR5gJItdMz2gK8b2/NZ4CelANQNmsPfiJ1eZeEqV6qN4RvPJ1ctyg
x4dVPLuseaVp8rJ/MCud5njJBiV/Ogvw7hl0qEW9FZectTWWk4/ccB3geU3f
2EEqwt3tbKu9Cmwo1ZJ5LrZ5ldd86UhRBSvgTldTr/sKJOLR2iD4Zn1Gb2pk
Vk0ugGjumFWgGYjcCAZEbXH1zFP2LiyPTCDF9kBqkvOq6Qglxp4zr+iaW1oh
OwCncR3bDC133yOz4HJb5b1azL5dxQGXzA8gHig019p4JLiwKa7V9fW8F79S
I2QWYSE4rWA47QZ7XwIbJsyMBSoATb3kXyLF37zBkBEjfGS5jo9puetdSOOs
XI4YarLUUXNoBan+3eK+dUWCBTBtcsjtAWZA2ViTT1NHmu/W7cgrEQrpLC3G
NcL/wbrPTvoBScymQdsCVli4A5bTn4z/taofmWvgd9EuvQvFNNmqtNk0Bf8B
qzKAtU+lYG+g3+BLbn/3yCIlADkDK69m20LPB4rFya5gKjSJ1h+s6B7z6E1L
VJFGmKgKYcLekrjFyi8gACvCOAmBBvPJhhDk2en9hkP2VsANUxyOC2zafghd
t7M3wrP0uzxbImA90+7YLuh95fNraxhla0VNBcT2kxiENXHnNj0g7OY2XzDo
4Yp4U9xuLHBpalxXnkI/dXCGW1SAxaC9vpD7O5cdwODb7qC9DFpvUOiCPJcn
5K9o03JT3Z3dGMyHe5QycQVtMgp6GPgXA+XoM8ZOQ5MLc+OpX//CJhXHwjOj
JvOWOLqaf6+c/t6zXtgtaUZD0MdoHoljJgZ5gJas6UyYSRR6eRA9+V9icddd
paC71Mw5gL6jlwepgJrSySABLNeEjd/cz0DcwiG2VtywO1Am7fZA7a9omJOk
yOTnmlTC1WDGzV1qxsGdhkzezUF+vJdrN/r0PyWITnowJCrY11206LzA4SYN
LA6+Nf2tFTfMGtcSbUZtGrwU857TZMDleWAzLoick1IAhtag0vTgVYICq7CI
r8YMB33oge7PT79ptNvoIVslFmZdT1rhMDdJYo6VGo/U8HmYXooJV/yU0Xt5
JGQKnOXBj6ditgdSn9R7Ax9JdekGVpZ4c+FPvXuRv9j2EWXVhKhhv0Gjmwzz
gBEvbCO0aijCM1xzBldGlluPIBcbDbDga0ukXQPsyrkJxho02jNmx8x6NAge
xhC/ztX/riJ6eUo68pc8fEfFzsnQu4m5Qq4jdqfsmqChvVtXDkr+3eJiQ+5S
DcgSckhP3Yac7FOuuVPGGTSh8Lv3toHeVT/NS3EfU9FG0jBFp0c9axSY4Sij
OTOn0ZoYNJaqHBFyuSY9+vmvNDSIMAXyRqqsqMyLynRMKSf5jd8ATlbK0k0o
jSFRNqFJyIx6Wt5ORlstCsKhWRbqRIyuN7sw3K9sQ3NaJWfPFixonP5hWdIx
1T7x55jL666A0mgMBtbAOG4nkJAxOQ5vkBjM+ktUGdWCxOMZGhkO52fEv7Ye
s7SFS4YZeEskpwiDTw+PzPh0noSdWJi5fyxK2iwed8ooAgQ/7gJofcqP5LWu
ZClp6G7agNgUWyFYl/SlHSANK6e7LJ2C4aBbvqu3QXY76VS7ahj+JCy1TQ72
xIeqE1RaSHic/or1eCBqysd/lvSkJSI/2apXyr6r53spg2So96t923QFa3Mc
Pa7HkZpNm8Sh22lOG9jQPipO0fh9pJMv+VRs41472Rwq8ldF59/FDX3ibfj2
NSAPrDMubkB/Vqautdkhl4IwAIX5Zww2t+/DgOf5uxVmYMyBB3nALXhy2naD
E/Zgf8D8/EHb0Bj0ozkvfkbKelvg7VNJUlpsp6YIan7K+BX5K9F/rXDS0Zh6
QCElC3o2r+EZu74XLnUrmwVfNjdOqH77Lsf6Y1oDquujC8jdG+tbQmKE2hXr
wRdwxp8zgB8gwF+2dDO4jD79/obdI1l8b6qqI88l56YLD+H/QJLyvU1rU4US
O4E7CpjhbemWdlzBgPAz4NFLxiEtbLbsd0g1E6ImOhGWtEhV7gFgPoowqEOs
ycCN7s7Y+uz6xuwzsDxeDCdBJMQnFZZoYlJkK88FO9BugEYEJHeQwDeBJscE
lxv9ILQ8kdKZ9UJaGjLxTzhFSwfBydT8M93ztwLhmQuO3YVSaT2dV4UTl2mH
zCN7Ps43Nol6Tz2URBAzwUafO4NJNvAsWOj/P5FKJw/9wh6hOznaQFOSwXw7
sUmUdWRp0tsE7dL12+z6550CTHwD3t5JBeXqsumEs8c8U2cJ/6dDEFLTxznC
vb2Lt6SXub8nrxKWBX5MKE/AeaO7QuDlf4sriPhxenvAX+CcaAvYAkO70CYg
R9mLSmM1Aqxg09xrvr3FfaxnraWPk3CykV6GFyetK80HMl/MNZb95dVyCEYx
lcAs8mD3Nj/AveMEzzRrtbOEGLk47ofQNrA8CwPz/5BpIq78jYDfNznGpbcl
/0aat7Wp0wWvwg9kDZnsHRq3a/4WOT9yu1yB++uEL4RlR1sv18UL4kymexM9
wUBdC0wtZwSGWF0RCpzgeYYxuB3xmCQOPN1JqsKadU1ZmXyFRiSCrMYDJ4KK
b/+N1PlhF/qicio12dZX+JrS3T3yexwz5OMC1pOiuleaFPTYFUPnTn6L3gXi
Zk23uzWYQJyLb+zc+Ce+Omg8OBNhJb5X8lOWcjM5WIIik04apE8ynhNHm0RI
kpuESYj3aZPg09Lqmq5OHCR+YLqheM2/d1Y7OwhzBaN/0lAoiN4Wq7NMfJil
u3QKF+y/u8iVpBfb0aO0zN8XER+FM8fhGY2jIVK5V8ogiSj0kIrQQbFIq8cG
uHMpRhdCwNwXFvhix2L+fHS7/CJt87EBLbY5YrsBpr/6CcxHJ3PO/xG8XnhN
qahfJgRmiyzSligK732R3hUzeNXzuIC6HdUJcZaoHDUtKn95nDHwuJ/gBVFC
BeiEGwQBRCKNwr3f8fTtKStEarJ/Ck3BrWQbmnExbTraLQFY/hMgF2mR4kXr
lK8MHkWHFRy30cL9tpAL/CfsJKUU7ihCdHpevjrAcMFTzC/f/uV2ntQrTsBb
McH+7edgDFV4n3b/t41Vlv+Pxn9k1t3ifuKPXcShBCIHd7VSgJIqmj4o59ip
FIRcO9aU9qvpG1Hj6AmddqOhuSCBOsgDbozxs4qVImSFd2EmE1uERU4PFQ/+
lLa85obj38/ZJ6BvSaLimmQAngKtLij0Vi2dg4XXkgFeZq7nqS6NQGeD7eJ8
bxlGaXWv95TEHuEex2tbngJ3MTrOn4hftI0r0yoqbvK3wxCCdgRTk8yP9N/J
4GavJRUWgmtcdSfilHxhiOpcUbNaCo+REazDN39kXkpSdlLsD1aJts+hko11
X/Z/t2CIRSQrdRW74SokwaYyG8xEibABDI5OPXOkjz/mudShLmvFR0DF7P/0
mg7U2jiYGAzH8lW8yPPA6zv10lVlbe6f+GK2glscVB/0mxkTywsZnmCdxUkZ
Sk0zRCuGpTdxJ3HfdEm9quKZhIKtOJ6tQEObLnFAGmqV4uQhS8g5IlLeLzCE
vz3Hh4wz26/yqnY7h8wb+I/jRtSh71bLBWONIxZgl3AbbyJG3PQozeNlP/Fs
x6KJg+bW5ieNG8eGqNjcT1hbmOw52+8CH4eY1T5eZxqLB7INxjkAh1Letbw0
JchhC4dD9k3TH5Nsil8K3wqbRAj5L5Oru4UtIHM8mYiyRkphlTKiStQgkDcG
SoEHszEQly8OGU1oUieiMRVzJVjplkkmfwvrBBwcwIDDgvkhj58sZ+cAxlM1
Gy1utk+AaPNbD8G5aeHq3ARwVeZB+JT2g+/9ao8GPSHTDvFME49RjXhrP+M5
cfIuQYmyYftGeeUODXc1HxrxHYgbnlgPEl/lrcDXJjFaZywwxfhWdkGTY2wX
vquV8J7l+lIzZrfLN2tFSFaGEdjGea5SYorzFC4E/UHxrVJYOBgnVU7Lt5xz
w6D5fd3ngaGBaWiayDKUjaes431E/nOGpRem9lCOblEkZS/z8JRv7ZqRfPai
LmYKQEip+Ly47VKNEAdABVGFR/DmoA1YrOkFuWsk2Wk6F5A5ggP90+3P/VPK
pqgKbVJMU4Lw55n/vve3zogKhoU0vi0sBS88WE7RqVZhU9bdHKlMTB/OtCPo
9z112HWJVKKzBPAsI7z/a4lI2KjI43ujvIYv45HxMAllIrxPrnbVUxHIcELO
M9zhnADBMmDmyy132lKjplMaQ+vWBgPFzsb5FDW83lkcDVmZf4zYBeRxRTEc
0RKGLEv7aEunA4SmnQ2HZeGfw2uCjTiAJ0gjIfl0UXfjGiMb3uTkkgj+qBl6
DJ0Nng8G3cBI/FIbba60cF/+m4q2qJo7FobQbDOYL6Chkhq4laQmaqL48CEE
VrLLT+N4860wnlJVtbGkCm95CV24TuH7N11v9HBrqqtscExTRXtW/6zCOGgm
qofKgnpDcx3AO08xiCSGxh7n6kPp3BHUpCs6AeSqkugsW57f9z11kiYntXDd
30c3NzPIc5rhJqnhrn6qU7eLpHpvbeYOBkefpUGPSVt2rpBIRPG2ka+xpUKc
4LBHffg8v4caeyIV7S4ak7zt88qZBAoH98ZzcyBJ9NUaD/Lko0ZQ0rZoTvZb
+YXSYuIXL4tGPwGXL34gCeTaMYsS1GhN2vYynlcLU4NIDhv32xCo9P66bO/B
6zWQHxue+tvmdx3rtDXzAPb/aBJ5KR01OnY9a5RE3FZFOHIdPJzVf4Xwzvl5
k/OKZWXWRHScWDkAASMGl53yM2kORy+WiZcnKomm85VaI65qK4apy3RNNEeH
82mUHEhdVnkPXIB6lEutuAzJKT7k0FkaaYVyIKvZsy79F8NH1t+I/YsHb/HI
VtqBfT4FAGuc2Y3BgijUtpbCnWEfx+ecjwuLs/dh/8UHKehkBOVEl7fTQ2wR
RngrhldEfYXJkK7S1lJfB4x/pZBnRRZfM4SMRzePyWwzi8O9Vfj+qfkyIWCH
N63WMti2yipyL/b2fk2Rgm0AbjDF2xgfdQn3BIARQTf8dhkYyCwtvL0JYiJy
OlQhDSssedWzExmRzCsAG1r2kYwJFLYlxVW/ZeC7lHvaqdEBrQ4dMj7HOPnw
otG2gNkwIu6fgQ20rhd8cSKbZoKW0ygighq0PayvT5EGfxZduwLKFMIiiZUF
zchnPgI4jsQ6WFRlpnr1lnHbi28/x6yL2DcaWTVx9/M6LRv1ilcuYzonaZXc
xWpxISfELagGXOGHmeavMt3lORFwzYosx92oMHm1g6AEqErH2nWsWFN8X420
z/ANT/AYGXs2oP8hJVkf5VD/fk7UUe1V058di6llJEft/OxUKpRYxDRzYYIS
wcRu5v2El1DcfDB79oXpFHSU4wf0omTwlq3cGWhr3IWFdca0vthUcwom+H0R
wKFgr8aVj8S1C3r5Z73s9lFsCZtPlgezJVXG8A+qPJvrJWiyDrjTwJquHAXZ
JCeco+co2i62j0fZTd57tpeXZlUBoaDhMgTE0cAeXfNWisY3uk2xy6lqX/rC
OyCzuIfa8JYjR1GrnBjS2Y2cn4RVx8DQqBF8ecj8eFvPQicV/uHNizHRhRK6
f+5BesSzXjm/hdc9ifUWFZOGMGCKnCGZiV6v+0X9yd32hCOzviUzpOI2Nmgb
KClARXnC4eWZMFJUYYkpqh9LpkOm/UUPzM2+PT6yNN3cIJ/gRfb7MxjnrldM
tXAQlhKWvOXq/ooyhwCW2NhcvIzHtgFHl/OiarcK6ryuGwCf4uZLKUV8bGl8
rlMEqkhy3ErMsQsmchkU/4V0/8A9Fl0ECWcrZ47xdB3qdUiSfUkjIz8NBLZR
g7lrfpHt8Gwj6plTL3XRElulwgrg3oave2CgpSwQ3A5vjwn+KZrcG0HXP6Mq
0JmP7hZc8W9VbslYDGA/XYWsDufH+V85xErFUuz2WbhBxpNlknzGjMUaY+p2
+7MAzDmWUH9tADvXFmqZ3IdK23oQluQgbH0/BeJSWltF7iki3TPsdRT00jLF
82rGMkZy1qnQwdOcrQ7bal0EyYBA0yYGdm59dIec/+ceLMA8qxNUWi6mO1Bs
8kg//wdYxB0Q47l98zZ60zyL+Eb4COhoIWNeic4F/2W+/Xfi47xovUnUwCDL
OqpXRYoKCX/L1DWQD7SGg8a45uZaoDMVoq8c9B8dNC7QatpbjrtiKYLo8n/y
mwScR+w48IQ3gMxX7QUVbfgMc8977hu/ksGnHoxtaTE0c6AubGXhOcRFuF6o
qcmpInu4OST5m9bv/9jAxV4Vi5mBOXFEDGk+0bbyW6QS/CX1u/zoTXU+4gOn
pmbqfqrE+E0iyEdTlbBz6XYiXW6zKHFfqYAUkiJ0D5fYBQCTcYBQiQMxUzzp
eH0QoSryxZjGUSrtIcm6Cpiw3R+FUhLdoAyJpiJyP9+Ng29+YIX8YQMpeszd
15IdpveZvK7dfwX7B3P/e/83Udxhuqu7Ge0JY24HwtrJsdU4CocCYF43Ju9T
bHCZVRLXZ7I8aGO2d56KCc422wP8T79aPHChMufMaEd+icXD2S4emOtuZt1e
pOHArWu7VfNA/L40D7LMflEgN4Nt42C8GtlBK2691xtn3kKmPONVveixK36A
1kxIC/jeEI7P083uwU7KNZPcaOBktzrSE+ExGilE9OAcYXUduxv/07fq9EYk
cVl9bwr3Lh4CYy0Yn4sn7+K5aatomEw3Wrk+WYKL80m4fRRVnn2DXUu+Mm6R
rRCU+Q3rcExcQIzMel0+mSkxsI0w8MZTKs4dDn3/A6eU1wjmxdYmtI+GYuoR
HWIqrnbbUW88Sdaj1H1MFs5IQRtlsgDGf3gi3YwKtkQVV8luOcEXe027xw24
PJzb8mjPei17X/oEA1WbxqMOxVy7bi5xqQN9h32Q2qIN2RaQhc4w3cR0gVth
osORMml6bGx1w+xbNFVpk7B6KJEe7gYWtbKcpmRW83sy0Ts3WDAblAyla/rR
vb2OD51JNK6y6bzgfXUNG/mo1Feo7yzCQihFiQTjUJ8USgqQuruQX5mAPTuF
Gq4eZEVjqLJgn/Q5FipDWtaqmp4ENjl74Aii0p50Cj1a7jpEn/Hd79r9K/WY
yyixH1LWL1n/xQn5SdZSJtjL3xbrgJu/bRzTQHtmD6LJLvQ5v5yAp9Z0gn/P
A5cubvLAlewBP17IZ1v2m4/6hGezz6DVJiwlMgrK2QGv4ATIbJineo77dILR
Zz7L5xFqFQ2hjOs5fNsCU4He7I9p/JmSZnB8Y0r3IOvzECdZF8Nrv4ZX9p7S
BsUtKraxlShnCtndNsPzgkIN0bBSbJZ945CaXIsMVU/6s269V0n4HFDu6dNy
d74sKLc0CxghOAe/LgDbX93T2a+pOP1BFwyRi0iFQUKKwALNU5/bwRaHa+wO
GARmBhzrDATz0Wxs3WDw29QuTQP7H82hwziW/Gyw05svD5tuSH/JNFu3PqOq
HY5DHuwyASmqTgDDUTonhmuDmZBnhLiOufkWBvvEBIF846QpsYAJgNI22WNl
04vJwF395oyuOkcb8BzNNAHFJb9MsJ+GgVAqJScSKoWDZN8Sqf/SAcJCHTxE
GccOB5SAEgbAlu0s3o5Ruu+h29LkB70Jse64qGw+smXIdGtxPlcZPwb26wko
6Wv7W/DR7Jm9kGROOP/aQnK4SYTyIWewvBQJPYTcvGJne0xZ2TGeEr9C66y3
i4qoSwD2EOL599Ml/gF+6FlNtIZyRkUh30V9MN90nQBqf5s1HcFwPtNFfdh2
wk8tdXvqLQYC/r0YL0MPSYt7l76B8IkGW47vw60Eh1hEyXsjX6rmFLRO9iQL
LHbyeTgl8Y8J6cvSyx3n7IrH/GufVHYfnqCf0i2Gr2MGKdyhinLU6GzqhTg/
yvcyzQgNkx03B5xu3eiUpxSWrcLek0TD4zNolEFx3nCZuzpG9jeCmpRWsD0S
ZVLFwXFqJX56HyvOWyBLj/Uie1bzjD7cpXD/w3tA8b7w0eeV9TEcgoK0QiBF
RPjPRbhXGn67kFsUuupiDfznsaX/z2fCi12+LKDyRAhEQX949rLQKPqRZFRr
mNCe2zgwYkPCI9/07isvsFPVf802pKznqLJtvvLNxq45dGEcRGnVz4gfMKMw
oPITntlcp47NEGkdI8QBXNzlNP63jQjPNfIV2Xh7mbHPw50OhmhBGIi3iwGb
MIKSofpr+syWotLRi/9cwvc995veJgue8SSfiMYVmze4Er5M6dzPX9eK5/on
cPgC8UdmKg22RfOOr2EJoyElIKh6UulpdfeAtBFPKtDcnndqBvZAzJI+/oc4
RVBheKK1OWPiOQ/dMnkg6avqqkDHf8DyS6fRs69u4CgmZ6Bu1CBKjKqou9YJ
/kr8FKDVtdUJqS5cbVT8btF5osLgCUuhhs4DxuFQCrmXScvhEqFeHKdrX+Pz
Btk6d2DuWKiZfQCl4qBRDKskgjMpPYoQ0PhY+NZyIULXRsA0sXLJ+b7sIibL
bZKXbRZUReT3zB8Bz4TRLrtj5BSpLoQ7hNZjwcUkrI8i3VojbRVHeGMOgzJ2
4nGfzZkyB1/3bBCT4ue+nasM1YglB+3nG1RzotzxMLaMzQJpFRDEhPOBBjIs
MbziUtqYvnGV1G1/cFLNtjdyb27hcBtb0CbDhi7LHW27U2In4FiywF9M10SN
dgb3MiWRL7Gbu9GM5dKsHN21k4Lw5uLVNf8UIdolCyWAe2jjLXzLA5miDiH9
7k1cypuvYqj07l7ZWv+iQ6B8nW0fmnr69YXlmplfHvJqlGwaL8pfvxV2sx/f
+X6wBeYY6O2nFCYRP9Mniq0TnsX5lU5NxdDz9jIZmWn/RjOAPKwtMcwuxOQI
x5LV3ROjHCyWfDeVa7gF8Y4ItuJp7+0SwNff5pVwERFYgaP2oiLUqzB6T1DU
1nJqUpWwqfR+LzP7IhPUt4OTymkVIbTr+dmCcv5y/7qfubVZl9b6CZwSKib8
ygVkJbExvGFS3AkJlFVnD5ucUu35yB7c40LWmZvvvOhAtV9/4H7pCWie72uq
jCgtaW2rYXkVS1zXtKqQvK1+hbs39SXShfylrgkvHz5elaRvrU/racHARu7w
BFF1Uk3l5MHt1VoYpHMjYrXGquAJtesN0PpptMMdgBZtO0kqq4hUJ0EoGvc3
MHMXJZo0jCBNWZESzLqYxbGd/EY2+PK+TkS7Stf5hqAyk+rJFhZ2lmBaZcvr
CesC1CH4flhxhQZ4U2bEwBc7maLwiC9LARhrY4lmhkhF74m2C1gNtBC1p6Ss
/fKhrIXej/Rb+Qdi+5qh2tHUPyqCiSt5LWdfPgjthWeFmoK5+OAqIJsPn66P
gKAv1n1YnnYfCDIMeRMME+wWLM2tGD/39kLK9j3Edo+DsAWcmY9SKvU8+UCb
ksdrgLTLdlhTjg5lw3VraHH5n1u47vNnmiTeOyfRn77xwnr9E8U64TQvvMh+
UEqyfPOjcvrfMXSUwYuttp+D3CnL6wrkEl05VQLkJEoLO6P34ggIFVEjXqcL
hNqncXZo+SRt8gyEbsIdAdI8ouuOGgGgLsh2ILU9Oam6cB2gLTSJ8Z0jkGG+
YXdti3YUkWGGdIJdQY/ZnzlOwZscq8KEb9RURmBZJADrD0ahf8BxN/eCRFFL
DKdqXUX4SQJBR1mKXiKPdnJ4YandQJOEY0PqOh3RudW9C8H76suZFC6RpSBk
IwWnfGNDaT9SA4qHllB+Ya8k555d2ROPXX1MIlb13GEa+EhXjKk0LazCYLfk
BtXGTLCq0PdvH5mdeFDeFvTTUArRBbGZM6s03VI1hvjwz+sOnGDeBcFlN1cl
9bpyvtuTZ8qvXFd5m3fwQu301FXSg/sR4g3PkFcjDcqqlH/khbqd+vlG//zg
NhwwCdWi6LuvPwe6wBsYnjYmN3kp2X5pat3cCeb4VLWP2j/kvgIn3ubLWVkT
pbksME06NI2CWJhrECAj8k++94VWbn3SYKGbl92p14zDFcGUBVlurzR5iQmy
TMIN4sVDWqNKqoO7sxYYK/LjFZEXnVd407i6ExV3U+V8BaJ8e78PmPj0Kr9Y
PRUex1OmAHOAJFHwSf3eYO026SwdOIx0DjbKMFkPod83mQawCMh5sZhx81dA
yky9xTxfT6pKy0tN/Degr6GX8EFVoywMLV82yM4Alc6xp0/QA5MDTE+8p7Ta
/1Ru4qhR4AnSKTEWLhe2Ul/GQFcWHQX7rU4maX2r7onI+GI4aIAEcehHUMCY
YyGPahE+6Uvpx5wrx8/uvaIbOMQq5smOLwXnnQmAp9iWPU5a/itJZaf8R7ze
zZFQzBKdIDCwdcGNf79yN+rPg3SUogCRLA1qBjWiRoAvtqFbMfFr2/HacGUc
v8L2LIRH/YM4tpwCGWV1p9Tj6Cwg3Bsy6MwgveV4IpBkGVx2dyadqxSRUfD/
+dxQ00urGDcMqbvMi/oKrijLBt7yjUJSRZ5Ky/6Z5DJtHr/etpwtu5kf2HYq
YBrU2uX9vNAeX4BQsLjho2dwbISGfD5H6wniDBTcur7FN3YRTi6b81G4wLQk
5YC3a17S0gMcAt6MX7PKNMD9B1U/Q7YbCzF1tWhjWHcjmBIT7Q8Wcu0S3qvv
rNBEfuPvN4Ze/xR3ZfPuAGxUmP93deGLtXHp+j9jA1UkUqj8GWYH4GWeliBG
Q3DpDl2QlLZVCBtPqNef/Osgstm2BUM6H4ZpqbxqQHckC+zJpCBrMFLrZy/T
AufCjn6d0FqoS5XLeDLr+rbmuU2KMoFAVmmdlwQcnTfOfY7/eiHN9xc4C5o6
A54BVhi9Mq0NHSKSCWrvcmEnQ4eXZalrqXw/mOLkmjCwn9VeszL1WFBXO+wT
23LA+YWgnUk15x/7JxxS7BD5ulzkqv0YreMu/PlKz82tGAOq6UvAlBsg2s7i
Rb2O1BpgkK95Te3i1CbmUCFW58sIOm1s88JbH3hg5CO62DWpwkdWaD5bjWcO
xNAP+avC5Os6RXzhZnnhFsiKwH1g3+SoPAVJNHS6OTTx8WEHK5bbKhNIKuMu
0IQouFXzERrhDXhZVsy/OjcrOv1T4DRnfdQZaxblxowIOjMT2SUexrIgYZD0
wSHyh3BgHY0Ag2vMfVPzGg7SjnVsUqLoQSV4AOg+ukH7jJ42ANnMsuRqGo2e
5JdNjyX4IzHBR6XbD8JhbaFu8ov6yNf55c4LJ72ymwESj4mZ5rB7s4vkHR0R
9ZR7zX/T/qMWq1ZzQcEgdJ/+PQV7jRq4ysszi91ESN+BGafhC0ezAPycwaM+
onAl1FWcvVPEKwfIxpzw/7k8fWEFVhsUchuNmaQG/4uPhTA/yv/Tq3jMF/nE
3tLcMMirbaAJWMs3Kqf2K6xFJX1Q/D2t2P8vT/1oIV7X2MhKlt1Kl6WQzaSi
XJ1pbx39mT9o67EmyGc6KjwgznCfGHuXWf1DVN/ZXaEC/VtBrDV8GHC4v8BW
d3/Wcjy44vBQwT8ip09rG/yP0rm39foEK+StXzD9u9erRtDXmUQn/dV4YDPF
kXIlaz0VjadZZAEaC9xqf4P6dD1pIQMCkUxrbnAQduTeuUm0EzOBu0oM73b9
ewVQN6sbS4ufw4VefqFGQ3a8xh3Q1h+I+iVt7RV8JAd9WbO31BXqmWWitmnL
By+H2k9+nyvclqWC92dTicWQjCV+ptwTowCqgM14QzxxewSMCNE7FfRv2OjS
r5Y0YG3rI3OqMUFkvV3XhDAsorG8/G2WEK8LiQsqPPRdH4H+ULni411ghVJL
F6xw/DO6MD3G9T1uSl7Dtw3l+qdwsaRyI/3iXLeJJEKY41RoEGbXS05qKt1Y
65ThCzKnre6OkeoAkHII/JcZRPIpRO4KgGpThSRxK3tPmndcKtzzfGYt3R53
AQxACXk14f3/ctypDb72RpS4rPaykCgK7pfkZE2GxHhjPEWyNq1jtczxXwC1
zpf5w4oJEtKUki3R8/rFhIiWpi0J2AY348g0mqDtH8Bnke0EnxyBzwSj2tro
iTAohpfHXLnTgezl8mvPgATnzu48YD+zPc0eaJLfrkfpKQAwLX7m4te2aml7
WGKbf5Z4qRIQlejoyxMRcqdKLfsUTA3fRIfzqKhc1T4jz17Kr2pqE6GuQAIg
vHsyyBnzER6SeijVgV5J0PJMaNvpxGRliPlTzwzoKBhFRPl6VAxrwoFlkHBu
OrPCrw+LmdR/D6pJXQu5ZH1GJKyxs5IDGBLJyEdt7R3RMBOxf00I2dcsiMn9
JtKZsdgTlYRquoc06NEIsACNah+C+hvPoKdR2sjaGpoCViQL9BGdX2snXguw
Wp+ViMZ+Q3WJuNeF7e3AYWyec/mOdooLe4glUeQpvpQICgG2f+YxV+Dv/yF4
ei9V3vQdALyNUbAqNSLKSwzps4MlGbx+AOxb3g8WjdRKqFu1U6eRXVW9KCAC
MlhYa55hDX18KFGOHJzwNN3In5xPXdI3g4sSybsquXEjc4Z8XqRk5R3xgIJJ
2fFSQJorFho2dgY/TUb9DKrKvGui4Kj2Ytg3myK71KsiI5K8oEZH71OXx1GM
dL0didqDDCO6NfoZxBbtXqKPpGShfElBqZeIPgOLXJ0xb+qsG7JRwj6KguxK
ITok2CHisUPM5lCvG973UsXGfXlKxhfl3+uB6y7/FKGJZDx2xk0De9O+Egyi
DSoC7p6eXt6LvFXUQ0c1qIHgUY6flBF5rKQ4H3Gj4il2O/xSWGg+7VW0O9u+
OkuKiOSrHFToJ18I+Jm965yoy/PsPbC1E5XoygkkTmKuwZNXk9et4DaxuVNS
i1PaMpnwlpwr3U3i2MPTxcGyx0MO3eq88I6u1RZdqZ5JQPkiqndx2rBodetG
yHRuFyv5yhCiV5XeBFcDoG/o2ZvLqrefOD1cNQ+G84xtgyD5aMSqS10G3Uvq
6gq0kELYrEWFL8KYPBrR/v57gLlJiKVpGNJbagOqBQT8xOe8h/O1XOl/0+AZ
5sPLHPP7dviy5h9jzLtO1XY4+0KDxZcgVfE4fNajc3hCV/CArZ3zZF9Et/GF
usOOW5fafkf3MiJlvj5esH3dQYRz7nl3NGQ2SJXMeAhPIk2KgncdheRyax1c
agDSzlltrNaMe8hKqcM2tL5YEyDB6Cg3NJtmvcHa9rspi+C3gu4QovFymGMC
k0JHUJH64Wrt1Rgri+4G7RdBB9BaqJYybd3iz6wxWKEhbEOQe/yvzmLXbRhA
AQx8jGnXGnIa3X1pPCr24ieLwYOn7f0E1o8oh42pPx0pl86KfNwysaoLk0b5
w6ffPh7+S4cMfgjWmKqu0+xs97tlc03ABH+r9PO8HtHnM7HclLR+X8/STo44
Dg34wu0H1EuLuBvr76d4M4P1Do3X6Jt4Y3KpmK/CiECStxjrVw3LnBSbzx3A
snUEghJENHYAt0t0UZWX3yWVP8QwdiVOTqm+NCigX8HS2KQaqZ7ikMjjnHeX
jrfEdcGkpuGRpYnmrQxHXfZvG5yH4JMgB/KTFypFtGNJsc9nGg6ntcniYPVv
uNGFrlyvZeKxItkzVT3p1/DaP1bMUPQB5YeJ4Syu8O878pYYGe3C9VhngZxh
Rq3FeGTBYrVhcHf4PRIKhoqzFpXA029AHpxfOEPZFGW/31Az2TrRndQBpOmz
nzeUCV6pXZCMC/B6BZvLb6ojohvT921ogZVlYcD/pq04QmAco7r8CJ6a+PXn
kvfy+5Nof1fp4b8xwipSGVRp8GCBU3YsgUvWf1eQB76d6UG1OWaIZ2FzFAX8
SixxuXrlj/oKuZ9MtEQbm2YnzPdPeKOnAK/upsRqVAbiFOOSvs/M+S+udtxZ
P1HHkHsZKxq7h7yeqdXp1rSUihQJe/XMQ/U5caugkbfP+S01XMuyEnz8OU1i
c0GXHzNMCQ1lerFpJmhmf6cD/SpQizYA1SBzsQbIjvbYdd1pGNzj3HuetQfe
d2cDmfSpuAwf9P/DPjkxNjpWLg1AN1u0oZi6P5+JI24sFXMDLT6F5qOqE/CH
EnWAA+PyzxH+pTaVPARSJw214eEU+/0rZ5wUCtPvajr+9VglXhjXHFSNiGv7
V2Ft6RB5z0zZdGzVcCG8R2EFekXguJ8q88sANRKuux2KBmsKBS7YfdItFHqZ
AMZf3aCshYq8TmEHt67I8KAbMEcQUEZ/oXTapH2QEzbmdPlGoVwTtYbU5ifK
j3JCDqDg11dYcoU+9rneP6uJSyx4qThNK3IYWfUNaYkdbIXwUCynWufoIbTr
VwwUznLWrxLXxouuIVhQ3bQ4sSW+YPRxj5SH7j5tA2q1a4XYldz9ehChyNsB
K3XxyOGlRiSfkhxzSzAdRM0KH43i3mIIFYcFvCXJ53lphbyh3h2nhc5H6qxH
7+xw8lbP/DKbkr9mieIEkiAsnhcBtP5yYMetwmnj0w9aiIR2+3L5BMN/GmIZ
nWmXipdhBtZH+VAEMW8QuB7SZpWlWIrzrYq37dvpqD/Ajy3fuPa2taF8KkNu
lWbOT+3z8yBWfU9vYfhWUy4RLofirFT2FeKpNue2ocoSCtMgUFl8XrzPSgMy
aP8Yo0eGkYxDiRbUQC6E18ojaBm/kdkVePYvC/e3qwaVTQBlv3mZdVrd28Zi
hImxPHpnjspA+9Vdr1D9YWkgTl3f1kX7l6LOPmpO6lyuYoMa//JhXABXLgXJ
TytaB4dkVsOwqvPXSXTkcxWdilCNFcufGqBVhxfoWaaeBkaznSPFrx/W41ri
J2f3dMhpQDnXL4ItLh7Xo3pzqPAfVHiF0hv/XcPOubic+ciO1rT1en2xKknR
IizZVMFutfoz1wDYxTSCE7XKMrSaxe2qyLYtZ3mAKcjoGbmYAeEUvuj0hr0/
/hJkKABJUnCpXVLyIDIN9orH+ffGrVNuX09ltyTi7pjznUBheEWBsdqBrTws
KnYhKfyZNfKYuFCrjZnsS3K4fcXjnHQ9LKKVZeF+1ceBVMF/5WbII3Gq454Z
nBrIQc8cZokGSwify3dJ41tfECQDErhSc0vWjgpLJeS9E2/WIA/pfmBdqS0b
6tOjbEaBc5U5/zVo//kdVzbTVCmEyUrULQaTI1wpw8YkuDr8MHE41VqYjA73
YnfjWvVTZGWrgkituUYqwvJp4ArE9l6jGhIySUbhdYEDTQa4kfbCiCgRo+bR
Sj9+WhU/HMEPFXe6i8R5FjyxlMTrNLsKfxTuwxm6/MRC+AWMcoP3EcSjmfB8
jZSVah66zZ9lpjHOFh+G+HTYtQlg9vVEUxzDQeuPyeYchsjtpJo6OFC5sUo6
aPxEvmyKaArrREYZX6mjrSqsn8/nw6QFSoY6kvJlQdkAF+W/6fxfY6d2sMU4
i9QHdua7uJwNUh0kJD9v9L93b5b/7OiFV8eQLG3cVc9rUQ1cVEwDQeL3ukfB
V89LZ1KNOZixgpP7L6ZKBfqXZweUEEAF6dsCSm4M7aH7JonZ4DYt/ejt1WWb
IOTHpcml3NYehd0juAlOMdZzYDMqfAzVwElTDuj31T475WXqqXUJG4LnrDVE
YBp3cRnSyurcDKlBWg0t/IULsx1fX+LSGI+m1oajnTlDaaiecjo9uoXjNtsS
0ZcQ584A4+jMuBoXB6/sew0wSo48+iw4WkaWW3okuax1RolkANuJQ6DSLpUz
rgIFCSD68k1Jlglh9/ISGJ7uNpeLJJ6dfq10aoOXH/qcdKKdXQ6qq/z6YXGb
8CjtdImFqht88JjVBPTvwGurOwUdy4pihEpHr8YHx71B6lQRFYBL2ol+VWp2
inkt7g/uKckamF4/cIXbEANwErB44QWzp4m3Qa973F8p4LXV7zA6fZr/ZJV+
jxFV4j/mYAj18/XB3iKicgGvnalRCeYXPpPeQAlYs/n5f3rioSnSDpCYDCLm
bq2b3bkTGX31jClcFRxeEsldfV6kNephJCFm9dFCMjcXy/w4McQMM7Y6k2OP
OF845+W6Xfo24+WSIKglelBPy364MPd6ZNfIfedcIIGqnVnwRgbWdCaryqfQ
oUuzUjldv5wwrC8DGXl/GRBj0l6YrDsIKk1a2pqbSHBJmM63syRkEw9nAJWj
CXs8dIZyjWZKDGkRgVyVBZOuEPzhfOoSl1dGQTF7j+bBH0x8O43qksuCZLWL
T42r64xGjGvE/vNKU6bcYmvVPGMz5F+AUDIbyve5ckl9WIp2C6+nlVe1K9wJ
9Rh/i9wCYDg0+ihISPsfXNDyxR8ULFk9GmwWRqKlailkLD+2NsS9zyKPgvZk
iqYLuZf+k27QNsFJET8hx82dvANo86Bgf8fNs6t5IvcEKpI4MSwVgPuurE+U
GA9L9P4su3XPOOk8gZwA8fPyguMOFXAmx9+w1bwaEEw+o6UTHZTdaiqvFMAa
kKjNFR4yyNRYG0XuUoxbF1q3xgyUmPXnBCrdwcyMQCGbyDupZ1zhNRoL3B7I
J1+yRB2BWOzyzNPES8kB95nMxfZs4ukAF1pg36FEBkgJxltg0TUgi304DnX5
+M8fQ/OdvLBmcAKui6xHXra93iDTyQENJt12B6Wm9x3jUQRJXi/e4h4PLcQp
TSZls56QMQgiI40O5DZMZAsJqzQ7YXN7cz/ikAhvD2o3JgPgBc+fFwxc9jqd
57s8UEC962HqPYzQNFCbZVFjO/xFtKcSQCNoUcjEtT0npd3mEL5ojBpBsllO
AMwrzIJnhV3ek5OjpFWshdE7EhphMSWZR1jmVY0v54A7M1VU5DYfJ5yTCahq
xLEdo/1X1besO1wejpoRoFCW3cM/NAFe1kpNasFbegmudUxrdjnAbRtUJmvc
IATKjGlJ5QtRilu1Q4i0GxZ2Lk61/O6zuJiqkg1ke99Ppte6ylNd2p6f7x/n
o3ajbAuG/dWYx+E1gKTgi9k+oJ/XdhATy13sNFqqGXGh6E+Ilquy7hbkfYym
sQrrRgachcrVy192Q2O9uKOboimview93gKW9z9ZYPZhm0+h0aPjurqUCvHG
wcH+tklggxJyJtVH2e838Pged4bn8p+YCBLsuBfQlYOSI90ZSbzSosKCZS3V
jeC2x7lUKp39eqBE56KMp0H0V9z/eNxThDb5N6t80ldQ838QYMQZ1pLd1s0Z
vc1+domSLJmTn65NTrpG1+01/nFCdm64yGby2UosoA9xADW5kaJG/Q3fO8mS
OBKmIrJR49rtsnUdnuKbzlyjb293YZCNpk4GHQImXUlRLMPbxfytmeSW5Mid
b4SU+lJGzpRKEWujaCorvOeDvX9F7A/pR5owRyLQyGJaiVqD9fTfCzuOAmlL
r25U64wXX6NB02UcO+r9HqgwEXXdxFBoxIjYUrSDWjjGhsLAzA7476jtN/bG
eLmd1mp3H6QnTNJH4N8q2Vw8gkrwnI3aXyC36Gf4k3j3RD2W2mh9XBo8eWhx
1nBeiaZqi+IKahncAMPv/P3eVoYGGXDXzSYKpxOg2HPEP60/YS7FGxpiAd5n
RLu7r8Ke6lMRAmWuTT9vDNRGU1IOj0tHJFJN0d7NmHvSpPcBkK5w/Vwnsx5H
8PLn37z7+aQrs9aKtSIpXAydwvYL4jylPHt87NI7Ut/asGbgqfGX+1HAmIUN
PREVBb9FmQdYRmGY6RXcKFXhtpur+cuBh9J9tUuUpToFhJ7rq3pWuMtzPqgx
Tg56+uSuz1wGt9BglWq1OxdPs2Xs3wq2Vs6yaUiVXsYc9jEC0SZ5ZTo9Nv8Q
deXEYQSXRo0Pd6miFFeJR1VUBYIBwUdk01oRyVjbTM/hFNKdwmXKtptw6V6q
jlifN4Ucupxc0Z4EsD2ThOxPXiPtZulwTQt9YeMOsnIEKlRwDDySNABEQwqh
TY87O94rwQVY4HJPs94sd80fgA7Kk9GDGzli2tcgC4eGAMzsdnxOGPjOTtIi
mGTS13A0jmqCsE3j4895MhcM+aAhGMVFk7i3v+7qXPL80dzSRIf76mPzfekS
8/7uwOdTp6OnQbt/xm98cEgutbOYSX9lZGpDbjKVBOUJU4GAJVDJuwFUzfGp
qhIGone12kLeRqt+dNWcgn3EBgWN6HSSEDs7xA3VGoyxG9Cr1ZJoTWY/60hB
1kKkcy8yMRtvpe0CVZ4Fs5IudA/Q/Q52kgUnN5zwwzrnvqDPf3jA2ARTgX1Y
wL5GwOyqHdtc2kPl3n9yvaSTfys7UD5EwE92OsVjucdgcaxAvG/9ml9mUXQp
kHU23/F/3dRJRMuWT1+/i3ta5FZnEGAZa/K2nZPFlbB/f6SlqyT8zlMh0+33
KprRT6YBQvj6cjRhVJB7gEO0sTnurBxo7j65xf1xvokvS020ZbHHsN3zCeFc
I8MXz9IS8cm3BN0n5bt3YND6nkc8m7+QezHw6eF5DlG6vH1Et42EZia28NON
L910vNFNm0Ludyiefgq0tlrP/iHk6yypirUqaDoxxbUPVC7l1hl/iAf7G2xk
RliWcmw4yEs5fdaUveRPeCiupWZlPF58qrDjqOnRfQf/ejxdfwpPt4O/2z8n
FYp90H0pmkZBrmgAAAeMz4o3o+elntcnlHuUpoeqhpz2jUKCnlBXC2eF695t
jntaEVq6yNLnzmH20o0jr9zOCx9VOO2toS60WBRBZXJW/Jg8z/2l/tDOaaC9
RIq0FDXp4UCzGioNt3WoDirql25HDTgUHboKB6NqvyLVgZ4Cv9DQ7zJaSQhT
VD6NO/FkoKgBesQZXtMf755K4vRqYqb/4RYPD83qwaSBftvsRGKoo5Zwg6uI
5wtC4FFL/vA8kR90qh4yeydPA+UiABuo9+UgrdXygIUmTb5nsd9ELozPziId
0g8mrqegzAk+aZ5Wv3I/6+zxxZAZZpIl7SLvwaV2h66QyrwpD3EumGGLPhTp
b4uxsrCE7mDRUyVaWpJPiCpkC5Mo6/JZpZav5ySefdZfot6J8fDk9Hiponwf
P29evIKTGNg1DAHBhx5IxKP0u/cklNn0tI+ZIQylhLRNGVV0P5Oo/JWDxc1H
eI6XPjTjF74n63J8hSovcK6b7JLETtvmRgazBUOLf7gqOefrzWnW3ZSHHwmv
wpRmFLsnXwMY0Myb2N6UCElAV7ZMWH1wxAJoMDAW4mj8x2MmlPwDGYMlU84a
uQfkhH2IrWnZLV5vMnkBiN0yu1gfj4tSxsydJ0ZTUEh3jdUBDUQaesCoPtZA
pNsmlTNm41og39TqtfjXrGRLTNdZxCxQz4euAVyZIOxNycqOt2TZyExhfXp2
SaQjj1MeCbHfdMny/l7phLaBp6JgAPz3pkzfFJK/39Pi3/fmvITKxIRR4lgG
N2OA3bneaxuR1mESC3Ys2E+VsCmmClILvtoGrEugtLIy7zvwsOTAhpogHTY3
ZXWU5EFwPajEm+CnI2h/TGYha1+U0QmZxJagtgcAzBIssUg+P+w+bTEUB3tJ
ZRsggROzoOCorD+AVxCy6nGhqYhDL2C2Um4JNjJ+1vvO2mWqtcQMjVsDVJ1k
awI5Y51/N/n5dTh+Yd7ciY8AsxH/X1Swq8AAtw/M4vKoiX8TDNtIxt4lAtWs
R3o8txEUK+DqcTHJ2019mFZeuQ/UInc/TA1pVDR/FPBqr+xXbsNbWdSMtJgk
OaeIgL4Xn7lNo6yzdQJwqglxLN4VWYZ7daefUzo6IE+WR7PImPBamvEO3QxX
zykznZU3UfxCXJVllExFMBAv7aVkP4DE38CGk1H/QITSv6XydC9Q/6URLNi4
2PxUyPokWB/eWYNzzqUHX2e7zZwY8ooE2Z9AMiicAWbi4CB1UIKHTxcqYPXI
uGTnOHpuVqdirwqoU7ZfM/H8IdvYnnVucJsCPF0S0ujdCNfh194WRZnrzU2p
ooeHH1cDy5bqT8pTi/bXKH+xSX18GzSftID72JaEW5X3rX+BOM2ETjqNYVde
tDW4XKtOlGLSFjFijjxDHEG4iOkhHsascRTJtKvhXsmpTshomu9kEwksnhAV
r09gEFoijMKtTsrUyZhxX/X4n4a1vDq6LLvXrHJLgc+4OalGg0EKf2zynhqi
hG6UzKKbtq9zIm0nRVGIZhHR5bp9cEaLgm2JSYgYwg0LanPfQE5dOVfKqO4b
NXZ8MQFN6oZpuQ3CTsz9401RsvxRczHYfHEQ4rMvC0kd31xDU4/MvynioMDk
l04ww+8J6UCUdVSR5MHADMyO24lWMZpc5yrpKfjF4O8QYzv2owmVdcYNeebx
4qyjvaO+bvTsmOFvQzbDAwyS5UrSqjygADa2s23T+qDtiQiesVpgfdu860dv
xnag7kINPY945eFE5XkanfLXz2iRkVodc0UBAfbhS2ZVv9sdWEExGoXjgnlP
YbLq8UYMptP7FjpFQtVk52v/LCqDAnEucJKPoDaJcT9ypQ0zv60sFTmroKji
ePv6sY/viWGdM8RRVsb0cvw8TKc79K95ZmNlneQrjqbvxi4xmVBW/6L8U9Qx
a5O0UwZwRliNL6iu33JX6YWh4ncwxToQgeC5MpOTbQ3ludZBbQMKLNExu1zL
10ixxPL/F0SqMi2PuxG7hSiShBYBtC0Jg3JonS/xgbDFMkroC7wQYe5QfObZ
ZfmW6szsi4JFJSFweGI0kz1UgUzeKELzf+lFkOWKndMuMvIYpDq013MXZTNB
3gfwozYJGkryXD48I5azPylHfyxJBZ73MaIks7iQ8H1M02KN5ck6uinyCoB3
PnRlx8GjfPawmcfOibuSMC1rq3vxRmHKUp0fdQ8E3n77mPOgXOBVenB94y+8
M0lvyIVNNXD3nqMZ3RkinPVCMHZdJZCQbgp4VR87RgktSNYAp4GmKglLF5Mv
v5K/Xm5ZpWwWgI8DuG71+QgsdxeXVByWicoi5/Vrch46JfK44gbYI+PmCu6P
hy75iN65QyFCWFFn+5cFrJ6W01H17fUNWmcVD8uK4NjjtYiTqDUqF04FnKXn
KbyxCpl42y+OTNKZXg8B/HCLCC+DF91ft7FODtJMWw+YJxHURO1sHyvscVJj
L9Q3lx0AIm6GG3BvosQxOaEdoFb4zlFWwd6h4joLZD42UrPiUlJ3AQOfVt7b
hL/hkWrq4NPKKgiwZ6hEOkf6gokURJNoZWeFI9ty7RWNkw+h9gXAhc8Ulu+7
s7lsCWtPYGYD5yBR9F5GwgN27k/Ft9FTnu/e40S+o/x5pn9Y/eyPSsEE9aRB
R2wLMM+RzdVV97UQZOKjHUPrNQDr8EM+H7H1KgNrWkkOJlJ4PbavF7MQTe0I
N1RzLLKSafc7a/zJNPk+G9fiZ0h5Fo8Z8KBxECvlwYae5wy1qmiHpDd9Q/lz
Zx867A2OWDWlAzy7yxxg1bUGgLfWYcEreEbk5HXopOvo3yfjtgVEkbeBjxYn
ijyn7OAUUCJ4BdF9vGW+efIHRDUGSIJcTlr8m0KclsWXfuv6CjvTirUByJoW
hvcYgDjTlmIRegwI7CCL3/thOOuyXj/ws4IoY1igx+dRWe58gy4V0UM9m9if
nGmtUJSkksi0lecRdWoIywjLs6oGYxbh1Vs9/ihiDsY0o3aLFQN8JedN2V70
AMpGmyG8elDSO0qMNuNLkqX1ztpzQkeCYSFJ/GDs+w9fq07oZqM4q12/SsZ/
pHeC9w4GTXbr1T+McbJ52zueab6k3XgGlqbIL9ZRX2T6XBqLc6SRv526oDK8
HGC6fAnPGimKirJZH2HFRigIjE/L6LLPIQrN2kBBmFKOAVN74/GAC0M+oUJJ
EXJ1TmC4isOzlcPoBOS1o1P4qOHPoYkAOryIaEDcrHMEh0ch9yYWs7rab89Z
HqjiW7zJeL6x02OpXP7PltrmBgkrPL5/4siNOdWRMW9YQ4/Xz0cohuAOku9g
ugRzY9xKY/SVUdxYU2B0m1Vuwvy6ZOefCoS8RyPPUKiSOOcwjNnhZ+vghvIl
vyI5DfniUwrgy27a13pbsnh5iroTDjcQrgPKnskjS6E+JlLuem7UkLdvTTm1
0cmWYvUYx5HLzPP+VXzgETxU3bBknLOBxWnR9pxDN8d6p+AQWtydvj3u+d3x
219hCFRmQTGil9WNJU/YNaFSmmkrMYGZWToOBQpGRrH3one1s/G4fsvcbOzy
eLQDET3Jl+3u/tWRVfCaTTQIm4bDruTbS7qM2OdW/fYA4ng12ht8lByhsuWn
FJXykKE8+lPwcV3CWcOl0pTsr5lBAhx8GaZ+JKQXDbwqOuQyXQBfO20Q4Czb
nGnchMl2a6MrztCb7f6EOxNLWTVpgiWNFGzU7r+TlZkuJdPv4lOWjnZ5rnwe
cHiflOtvUSDSXUonpekGw05ZvbbxU8hb648WzoiuUwBBPp2ju+QT8FWf0aEW
xg9et2BwmCwHy7Ijsxooml5plR+ZP5OFSVjHkjBX3wAcav+hZSyYeAtrQHln
dLsTa42yz8/KWQN5JWbhKDGPrCFxC3tYYvxgb5N/IjxzPTlh3WscV6lD2tFf
K3fuIm5l1/5+tMIkd1Ae9mpp4QjatvtqFL7v952rILTaoZDC6Y2LsA5HcpQS
et8q9gkCVbcY3cieX09HqI6TWyBD2VkjL32QWEkv8psBBFimVHctcHEZMOV3
15PNR3+PzUEvL31GqX9FwwIcoIiFWTQWVlzssImuu+km8jSia7wFze9NZkAR
kv87JrA5NsUh6RSWdN/iMbkb7i8kyvQ0yWn7579izXtXhpFHBUFP5jLKrYI5
OZG0a3MNbKTs1t53kA6A+803ZHq5ecs0Jq3ulPP8Cz24Ti2GtnpVVyp6Von2
qfk/P6JS+lUVXaSdu4uJUa8oSP+g+i05dHigJG8rgZDY0fMCcTn2vShgKA3f
SaQj+t4bKODSnvR9TMfxoLqEnpFSyzcTGpHOZ5I7abGpZglwPFP+Ot6LbCQ/
RUB3ajyUhxMl4e8SZLnX403U9Gy+x6jYNRSID261gxy8kpI4p0VgLbwKoeiu
RklAReKLNJxiNRx+7lbXXYTYnbcpU/oHrdIiv61QMmtF+//1A/Rph17h3oO3
gy8pI7H02kv39Y9+LG6u8Wf2dyhTcd7aNa6OurTPBRRdo3c1JI/UkW468nPl
AO8E23W31Fc8TAkSUIpoPFXaDACJoywJoNQVWLlVNFD/fyTPJcEvD6O5+y+B
GkEP8UQ38Xmy+Y7geB6A3ljSEkOeoh+hZEYMAJYwLuyv9jWD/wro8uo5/9rg
rMwTGiJ4ottPZ7h09cgQgPLoz48CSw0ZTNNx1En5zZfn0wmby2smg1QORQ0k
jm5naKWQ8X0zgO1uhWn0d3YsO9fbXVvwpUMIeQcTWw/lxHAUDfKPudcNzBF3
iCaPxjvrj8JzwvQ46YSCmQmUtvllWVqpATtM53By/P7KKIKvqQALJE61pz3S
6Erxur1lYUtPn0j00finNFXwAL2bm65yy5ha4KS2ZqsgyOQ6Qtkk/4MJsncT
SVnqge6QSjrAATEWxwocZ6qexKOVmTFWZcTr3MV8Q/2/YO8oCvFAvH7RwloH
SQg5yHJfdULQEO8DqU/kwMv/+cLNOVZQyI5yCpWQriyK8OANJB0ZtmPmRi7j
tgdJmaLSFDb27pxyUyNZnpE3/7YPR/H5GeYeLNGCIarDb27Zw2ZARLA8EqSs
kortc9vlmYLFSBtnl4o5ju/E4fWK+h1KeVRtUk0oWYSB0gLdxweR23ki46PM
1auhKtXyI4EWVnmMiUcmpZZbfmcGZA5lG2XzNdGjOlzKztxzqnbMI97sZty+
A0H4Uh++F62q8RSQT162fWJGw5FEp4BQ716wbUWYn4FaFwn8el9VbbWDSCIy
9tyeF4KrDwESEOWkXVXt5Ec3qS33xybsJVHggjJ/rCMCx9udzkOq/AkqYqzC
SlbaNMZDhDzdKbQvIaobz8ZJzO7M5Zw1TzayGQze1+0hfCwoezT8yfzLYYFj
6sYxy1eHUgDUoI9rvqzAYRp54Sy9oCJpvimgVy+XIL6MrL/7aVNFs8Iy4tyA
MLxdbXavxtwsUzFq7XCkOnaY0mWPp0u6QPw5pRbzlggPTePGFV7oM7aOIMKp
Pz5q8zHuvEWf7evZaV6NI40Fh2WU9Xg+KqdfmPBvh98Zo/xikjD0sMJg9dxO
ZzUoKX/WOv8jcwOAh5XX/28LfYL1Xmb1GFJ0L8iVlIys1fGz/smZzsoTaNL8
8OXy9G1Z/jgCEhzdx7vsWxeLwESpQynUJ/Ln+0YgYp0T4JCebjRnTVD4askT
X2I0BxNrQ3sX33t2jsxlIlKtu6KM8vTRFOdSUF0is/Q2o69X3ff9TWjBNsEj
KoEwGN0nYuzW5hUGYZZmgPq6OsPvCb2tWoplufL8noRcwsrp1UviE2Kz9+4l
uf/LHcHy/+SgKZTazZr1pTnUVuywxuVv2Kt5kdWO6urjbk2TGeURosec5KKF
ly4j6w1xai6SsGXufsnZSE4h71WpJZF9lCRkPatU8HoPzWUDfbLSavpzr1T6
mxlLp2zfMDkm6LngWOggx2PXjkcSHmptKE+8/LbhitEGYlb4TMbU9ruP7m5P
VqsZ9h3mPz+JA/K/CRDeg6yl0QJnJmcKKsHKNgh6SmNrRJYW5TXBlfDqh00O
CT4lPHQ8HVS72XO133naOiNIWOMX5Q/seTsWyt+Ok5sM99ItlPPg5KqwGgLk
+dMAGjSs3w4NyAy4X0eJZS+n9nuSrCFCl/L1OQ+vmDHCDOMOPsnQT/tgoMq7
LEGDYvpN4BCv59ZBZMHnIQx1ek77Ze18WCrhqcokqFaDhJvDOEnKnSrAgvY4
wsL0hA3PISEnp4nPqaEO5E87+Yd/q84dJV+65KrRCl/G6zKpxbCMSuV5i6qc
VITwH3Zsflkwby384m6sizJiW9Y6QJeryLxVrynw3E7FdsVT2JEZIUUSJycY
5eLp6m+eNg79Cr1JznfeAYCNPJMblkI6IjLHHcU8qALhgTKDj9sApQgUTMvL
suDXHqAH1Jv+nmBFAWrmRx9skxDS3ZbyxynWC715LgFxgMHnNVW85/6uyDRx
IUu5M1QnmP3PrkxEWornBjarEDcDTOwGPEPl+WFG5366LZ+XskAyl5oE19sr
ri4NXVhhxDeF0dRlY/6HDT6qsCHODObEEGkbEjK6RqM365KDIBXE4nRKlpfQ
f7kidGF8O+6mjknRse9OLKIGesJH4ly+hH+9T9aLrZat2W9FbDa2CicZAKBq
w6D2qT4PT7Ra9dEPDoJwtvetVxDU+XXbZmDv306m2laeUVp4nbuga8HYu2Vd
/av21J1xHfYNhMbRM0dNiVjvgmAuwF6XPBupOVxwz7DpcFrCc52kWPz+3Fka
kvy88Pyce3NEozfDD+Aot6ij0kJRaUZFHNuYqCezw2T4nwF2leJxeEfEtLaf
Cr1aJoWBQdwvQtBsjLq6bxFh1pG/GL6rghw6Qg9R3qvpOIPDTFGsG57dYCQO
6/SxrxOSfVcEvRdntf/lQERdXMeK+XNoRWba4a1o/4dU7cCiH4Vr3KtwoJ2T
ANs1EvIffOrADcdr3w+c4HIWTcrpK7d0X4M/LPn8s9s0rx/0/mjlfuueqg+X
+xAnibSp/Xlco9GDwCTbVh/K9hPAJh6Jw8WW3xTdyy8/8MZU25OjZd5oOW1N
RTcIZxdXkbA21HEfQ85nHGQohQmp6PxgNPC9ZsPg0eX1mMmwMRfbBRASgUJi
EZFIqsx/53yYHk5pNALMUEpfqHRsXUTDK0RduFGm3xQ/VDl1f9e42gHD3i35
AInnloIRVfdzW8jsJViNDicQ73b5C9BxiYUk49cK/asG+UK0m2npkb6SCl38
l0IWRJKHvJUY0X4Sh+qHl4COiOcUDMdF8PUEOqtxBQX3MwrepQkyD53dzaV1
5zi+ThqoKdZaNUXyEWOr1Dmzb+qJHBfKL7oZfq0kKjG6YfFOYgwiUbcj44AO
ibwS9ruYRiwujFcIL+QqvDBpZFrJ7woVgaCBkiIt/Si+Hup8TfNZfT3HFQ9t
AX4Ji4lkZTK6RDI8tkQBnaCJPYpJiokdIxK2IuNU0kYYqN6diMhGxDcR5SDz
Nl//d2T0BOTUc92M6LCCcKhsA2JB1VzziHEG60OUJcbBfLm9OfumB9XQEP9B
rq9lvuBTnfM9+QDkE/091udcahULBFFR7vZmz6/Lf5cSuEvUhndvD0bXgy3G
771v9hIESrPRby5orTkfikh7HaP4bOgrx2a0CR0s/+LDei8aybtyl4D0IvWz
LsApIZmn04eEOfzWxeGrz7n/0p3HE5c5rmRQG+s8CXs2yvw091ag+xFNX2uE
dLuQs8r6eqTVhH8i9w3lxBRrScMkfz7Py0qUo7XRhWYUJjG4JmNFKxTDvmz1
PVDF4IpdbHx4R2sVpBXrfe5B5An/Gyliu8iAzMoKx4CZ3uSByJ+lwCvzECdQ
MVfh+vh6C9t4NAJh3FL2xc4V9W3A1pHTAKbfJViijGdcUVK92J08TUHbwOFR
gpg+eu+pEqJdBNclEvPoUQSi4/7Qq/uZ+5csHeDK6WvGMEgNfurk7hFrvQgw
Gg+VH7lBK6tQAuvgeGVGmXsWKTq2B2lDI+sNXJ8ZyQ7fCUi6AtZhwWzQb6Zu
380RGbQo14u6qqhCvhSWq7r9h+5HmPn2UbRZKZHtbkXqj4IDjlHpSbPvQW8z
yBkUfireDUNfniXR7SA2P2XXkzkQqK7ZWhwjQLYpkwn0tIboW/YoFgte4uI+
8q30sc8IsPGPd4qndnIR9cFGGT+QwVLT/BSwiIbryEZ9LpMRvPLgT8M9rgxb
TZByV4KG9ejTbPhyuB6LnuIg32zg5nVtqYL5RS4kRzk5GNp0fpRnLsMTWt1M
Oxpe6mqRTle0iy5ECG890OjovcjEUumZExN/UqO8yNS7p8x4VfqsfsM9V1F7
PSMit0PXsEx7WhiEMmnMnnvzVAtxwxZQV5GzwhJQgWIQEJl+muJ5EStDyYSa
vyw2KPYWj/Q+elT1v5BFgGIZaM38SJPKdPgz1u5IaUv11au/hC2d2ppRzvdW
rDWNDHup9TsVREj/B3toKz4bbb9JF1tEtrrC8zrlnvPE+LxyB90Dta0eBR6Y
AMZQZxVfP/bKXVWrVCSjEHMCvUZ0P6sMPTxNupW6n1ITGOiQI8/zp/9TU8o6
nslT7hPeaam6nvPMpsW6abdgsPLuwCQdkHPcHDAYVm35obo6LYQPqWBdmPuj
6mK7FTWh8TQAp28eZIc2LEjGI2xeKPwgneO4AEbZCJ3gbpArf69yEeJQ3Ey1
J/yBYeaSFGxrHxvv/oC1oddCXDdcCBsaxeBokd1rAw31caby2zssclTamNUE
PB/41zl9asy4zssTlYl/ocCck9UsVcZ/fhoVumyEXA4SbIFRbQRkaQQR99p+
cTr9fHcv5pPntT/tuppTkcd3z+jt7y3pjo/oGiQxxgV4fiWws5g1XLQ2Llet
Dt+VcY1LvVBtvDaZZfK8Ehbd12JvqWE2TufqaweasZC/Ej7o205gK70D1+tH
f25iPQUs/4qzUg47uMq1w2FBO1JOZQFHj9FGTBYUJ0hCL/jQGK40ks7BOLza
GX4UfW5QCEpBMPLYaMHuVezs3brFBUXG67mhtLQ8zDK7aP0DGxmUALZBUp3u
gQ8V/quGXQ3Rdxm0hJ1aec1d9Ku+GXjav+GdwGiac2Cs03GEpGG7o3ZyWilj
Qo9AVmk3tfvQozLyATgMgQ+Bt0xKnzdBhvmSdq0y/9iZr2PHSl96lii7eVFl
xhlA4lSmaLyktHqjmbwYz966hlyGoPL3OHren0NbpmKnu4tLzTAkxZjrITA0
nV9SN0LdsQetoJc7+6ZLUoOuLwLyaWZll6oT2FwABRrE6GiKKI95fRG/c3JZ
U++g7O1X4APJrQJDi4inJ63Fe6x2E1SKLlFeThJVcNMZYEVcbwTVD0K4l0G1
XU+5j5rlSoE5urdgzNREPZyhFh/814yfffmO7yZbhC8GE+WtY7OYHqYMlb2r
xkYjevZcpdd1WF1sDOKTc0trXdnW43TbqUlQLnTu/zunXN+YQQNVCO2m0HJC
ccIZb+4RDlyFQOWAveTFm+qQDlQRvG35dLBuE9/gYNchZQSF9/Kxsf9QAKdF
FzDsc/hk5ONnop0O4InpxxAu397sITbArCw3KKVFUFNSpcFhVuHrfGn1ojzE
FskUW4F8uGpm7u9M10hwDlhIYeCJdyg1rpMfxg/+kfFzy/NwfEDxbgpc0QZB
j6p5UcG0LbuKukKhqMzOGerY9LnbNvpNS7NCULgxjGf/d6nDy/9JKZP+AYkv
QooBqB84oaZzZnqxXnPqjP+cuI/dDbkVy0tc4zbzNr6XekA/Cikb8tJ9m+AS
r6uBnNM7kHIhPuaMFyeGIbbb6xzQsDfDnfl/W4eLWn5MsNIrT8WXiIzjBhDA
YYgR5+j+zOBsEa5TM1VpbjtyDCjsKYEvR7M6urJ/JKnwma3ijBrBm6rfAB8R
7IAkPWbqDORJo9M0+fmdV2/Lz6IMRDUqHJtVkblqB9AkoeP0Kc5wyqCMi3CN
X2QTSdjuRXbZrhfIGsfD1Ca2I78TPVj7TQZbtxIagVrHqv79s942uXr0FDmS
7l41Z1cWl67IYqAQfZKLTBdpPCCgJarIxtmw2+izF1CGL/yvgWnzuVoCelKX
sbQxY2awmTD/bMF1irnEx3RWfZzisvXVM8BdpgjmnG0Zbq/DdEm8F/Jmbdxe
HhXRQP09AYanqptf6D6r5Ke23+omcIE6wrKf7fEiPHLxSzHhSrN48cgL6kSb
sk3PHCO6HxkORYf/TF7WMUH9SrmKflTt5wrUpgJVoD8nhzpn9n/MSZJjFpZr
ma/EB9YUbYJrdu/6bB6/VBQBgu3WdcjC5ofjM64BDR7uT0gNSgUjmj1NfSZW
DqfeNh488dCV6t5IULR4gPlBQGbcZCgY4Gud5YjVudklLQmayeJjjqIvfPke
dR02jDtJNEf4B7qlWMq7f4R1s5Qcs3StNfa+REtrCRe7wEAGGvRImTWviZNH
rKy4U4lSNrR0TM8f6i4LPV84BC12bI0xeUJFoYqNlShZoGRgMOTWo7kiY3XW
4LwUdXttV2dU2lLdmKXesl3bnO+my7Hpwl1nDt8Y84aoJpMXG68IyiiCilPN
mb5sQcSscMkR0OMbdZVHGJvoZ8i2mrj3rafpBh1quIRQgtoZGp/8fpHDZUsn
i4muykmQ0jR4nClmN/N4QMVaz4TUCZW3JFhHO7EvIZoHh3c0wIKclp3KJrJP
zY8i5uahrKMR7itVOwDz43dNYT3jc3Yrcsw2SLhi9EEW74f/fEcARankaFrY
nxypE9i4CdqcWmCPL/trTA4cHfKYFVUbQl9UaSOByYvMZKwzv6Hi6RSObaj+
yywFz5+uiGt9b5npGWMurf4iHMmoZge9U8vhewbdIKKY9P9MCk1oB7KYWxnJ
DikwTRaXDeiRgF0hAzLq0JIa+Ple2HwPgRgz2oTamKAWwJdVk2tWSsP8CD0E
C2yyJNLlxYTp7j0kA626xX/wN9VgPQe0xqc9Gy0cWJGq1KKzp3Uju9lriwj6
p/K/XqvgiDPO9iYWa6pCWKNI8a1Ou98e0JY3YKu6kEs8FgNKMeAf5DA/BGLx
AukTNegTOKfiVStOYmQFU0CWzKz+x4TC+SOn1tRNqvlSeb/gx18SwLvZ3uaO
lgqLDb1+olNDyC6IWpY3UC0V83m8/JAakmkWsPo/McJbSsahTSX8Ks6xcwpP
xd5oY550iLxx5Ahvc3lXSat/JeV05CEIn9gTj00rg0Sdfluwsmk3mfB0/zrn
l8i32W7KZDkG2YBNCk9OQtfSgIJUXWd7NpFKir2R+rj/C3rCPQ3nq93dscRH
KvTq7b1+Dw6/A9R8P0XRQIXvL+jrhS5+DKRPq3H5v6HWRdbdVbVldL6Ozmib
E2HykxcFn81xNpyfESrdjuZ1ZL2XICpvFmC4wNFhs8j/q9fem1jD+SUhQ9dI
mGIomxHqWMH/DEdBxwOKsNZZSttV2nWnpw/C+n+wyNtAIjUoXZxy4t9a8C4R
OnUKk+Z9ZzkgRNejfVe4+JRmLyyo6vYSx0XwrdskQShidSBUYUVo5V+rFE1i
CWs/6adADfce5MbbUkVvnDoA8BsvQLCynhXA5O+eOAgkrA21aqH88sWSloTm
3mRr1KObZzwL5+eFWOn5ONoqC+tOhTtTFMxiK4NqvZjIgGcCNJrltBP12UP5
XM7Eo7ikK+/vXX1xfd3a1+wY0634o8kzctg9YTaFKTb5lWv9jxkMAOSDteLX
FzAk/bODlDzwenmtrvPcyYtdEwvw2E3JCVeolN7z2bWNNUdFua2UJaInzdIx
TWDNIRgE9T8XjSg8CubMgSD1USBKTEypnqX9cXqL+Wn6tHOYKr7NBX1YYEhr
H4qxn/q9sAw1OY3WgTQY6ylIqj62EkNiCNhOSuTaEBjq4kvBCLSdT8gqILYd
gkUnH2Qcg14f1gvm7ZuidkOZhfsaFcHTpPurf6+WSBqPj9sv3LFYYcH1aP1o
p7OZg8gC4efEJdeveiSTxMwFPDjLD/rjmBetcijNcVidjiRqA2dtOlUhP1Nb
JqG0L7S7O5dScuHw9tDql396ngdGbSF0rrzbFQ/d+lRuGN0fLD+xx7h12tg/
KFharXGkPk/oOLUM0A64UElbKjRiSqvAi2YsIUExCdAXjVKHWjVqKlq1/T9V
XGHJbed00d2PmgmsDO6ihoHT1xGR7aO+WY7rbS3FJ9JQ8Dv1whV5nRGhY1eV
PWA4Cz8QTgcojOlkrKTPEv5BVDRvfHQLAcQp+Qf9/W7Yr9wNbHw5vLo7LDXd
yVoAFPqUBn3z5vpeTVQzwnT8U5UbLeRSEIqw5k1ZemNUQlqiKpm1GL7WsM6E
Nr0NZlTN8S251Xfu3br5KjQOW/gbiG9eohIwdWx/zhaUjKijxMnm/3r0BkFq
xjZq1pXhrVvYguGwdXMevXAxbI9/AVfw1Caotvbp8lsroBcCUP1GjKHQQ8iq
gmRe7MhqH610hoEhHCB8hp2KyHGjHGoS2ATsa2BijUj0k8Yt5BN4JxHs324S
okbYRzeMmy7hls8Iy3LOb447NXZgmpe0+VM8+2ywXW86fe3+NF+zm5Hi9CSc
bNvO/X05lzGagX4eT2SeIFHfPmIQ1Tqd0ScKHLxzoXAPjOQ04UXstjQTkKvd
IVdSy+3ks+CnoSNMDFZ6KQe1WdXb6mJX/qZmaZTpONiihWIlbud16l267Idi
nGLYIKPrQHUxLefqV2XXcqxHyRwhkCs8mOLXqYEsimz9fFizLF/VBCCeq+b+
6dDcfgKe2GDGFwf8dUWxV0MmnNTSuMBE9DDiKvVy4uPTHR6qvtFofkphXtRk
gZ3mSJtv3HOPLG3Ywwg2kssXBUNdMpqZXhVlK+tb8sG1bkhWTJTMjmnFBkL0
mquyMzmIM8tIMz6M4RTbP/phnf1JVoNDPRfm9GQ6NQrZuyLiqMVg4/KyGEAf
lcx83BqMzUZy4WUkF7Shw6T/Z3pMpu1nQhwoypy/PZksupmmIL3Z77QecrES
6JrnqTj1YZVH00LyKTogwJJQ3mQtpM1UqzydVd/gVos8ztY/yNipiRff/rnK
TripV8LFfy1zntLWtCqqsKsu7QyCnwruNmMzINUr2xeju+2ziQlO9JpmCAWH
HaqJYLVQBxsN7mOB0u4FjRSUIqIcnYgJpilSyXGOSTY6mfK/pZaapcp/ShzI
logI9GL0LcYCA7byIU+fzJ74yvc1mgJbc4l+FVsVSZrsfqnORlpS298yDICG
lDjLeZkDsaQChdyTEROwHf26iYkWQ8RPEVJi4ZLbEyzTzJO5orQzd932J0q4
o7M2Xvn7nPwOD8OSiPCajGlWkcLFO/DzfJhl8g8bFrSJfe+kP3S9a9tLza4R
f4wf95/Yvzfy+N0yFE9p/mGt2L/vE9Xils21P0Ti692QWUw53GSF6wy5FXgN
FFjYYWZs49V4+OEcZmrNK4nDVEgaIWMnhd53HHXxFu3kgpvTuWE6bTGBifYG
L8I/TNGceG037Kw+s6H26uHD0dFfoHPhy+Zk+8Pm3OiizLujzOxyiwBxmPBE
QcZTGRewR9bWiTsUW13Ps1UVyA84wim2rH5P94Hpd07psW/jkmVEc/apNa4g
DpNyPIBb1g0GqU1j/bFKYPANsFWBsZJiJlh3yed9vsi4g4zvAdzeptiZp25Q
6Py5NmAG3dYQODVWPqsEJcS068qbirj2VHGvOjr3FnCcMdsCVY/PHNyYsCLV
i9UuSRPaUbiiHypZ9k4vB0POd6e1dFQKN7mmj0gMqRgeCXUmViYR+U1FDF2l
41ba/e5YX487rjbzAsgC/EGSpzRPctbah8x/qvuZiUi5P8Eq3MOxBaP5Q4tY
GQaEmiXr5330VbWtoceSADoOuz5Pi9S1txmnwCmfzbcnDK3l/YUuVoa6mR88
7q1Rr9C04SMDH6iFYdiLwS4qqoNXl6hBaH3SBVLU/fNpE70JmHTilYg5AjDH
LbLtwGGOkWseylc9zmwFnJEcpM+rmki6e4Du57Ex1ZbUSP2a7fgYDwlWTgwK
W+GAUEQtrKGJuC9g6p4Nz2bdqgJwMJKGxPNIWwNbmoww3v95jLHGRmvlOcQu
g5a/eFbrXEM0nEpg930ZfuITFFT5Up9ymQqsJ8NQihJ7v1E1W6+/AbKJ4fIJ
WVyM8vEA0IFZ4ZHJ68oCUMwZO1qD0zH7mgVm2bewKU/VYkDv8/QlgdNa2WG1
9BxIZveoVyi7m4MqPrQacaF3X+O0ovFJ57sw3XtUMUlkBlJZk2Wi2U9po8+Z
370LmmuC7gvLhv6vZ3y9tFm/JhJMkPy6ZvBFvIud5qzISHpf2pP1rXz09tdv
pU9wEWU5DyQzX7A2PZ0oBpjWk7yBeKMlE7My6epJJFg9xLYoP4rxA8BDkqzU
uxn/ZfuN0+xVh6iuDSVmIsDxe1Ewgq1/JTwfTyFYU7dK2rClNRhj9xTRrZ2O
jMZPUakWxlnr01UMfUQigAgPm1d3AJEdJjRnk3+ahyzMyOtLXaDD6L2fnWps
f8BlVJcxvC0BeeaShnzgEQ3dIupIUwKHnOfBhd1DZzmLO3Rfv8uaGWEr5TS5
WuoLXQdmHW4EQHYSQtu3R6UDGmF27Jt5BZiSlaCeqqslW2R+x/lzY4yrzaAr
7iAglIKL7HFPgBB+F7JLibFj9IDWumO7DoQNrL26fztcjupRuqgTDoXJmAQB
20V0OZd/6DSzXxJIKljELZHszEwIv9XfBK+D2CnHusVqB5JVZ+veQDdMOd+S
8umDVcaDSoWc6vqKPFFbEy4K6OVHbFXj4OmLPJ2C9WJixwHhHkmo7nlHkTGl
cFHSvegwIOQ/I/fcnr0++GJ2im5gTjfxhuoQx+WxVS/tv7JFmzs0or7Sl3V7
MT+fdiUu7+XhScjlg1rjLsUgDjgXcSBOQ7AtFrenQi9cF8B0c6F5eNKOzKdl
EFv9vJhbt8qHBd6uwE5/P7Uo+yzdfUxVmy+kiTX+27CHXvIUa537RDRVFLKE
wAlgxJnHw1Sv78+UiX8dl+XVMHFqUKoU2NWQCfOaG4tVflNimjzJtMxT15L2
HAPFkEVu394KFGeIua5nepP6UhNI5r+zrwZdzJshLYj8HB064m9q9kK5A+9X
TxgzxCYTCpHTlpZMvUYqBdKzojt8Ys7uLEWTy8/0pITazpIWRxDNIPODM5zj
H/VNI0f4p5ArPQieiUJGkm+mO//AcKWJK2LKsoAr9p+pqGsveNBFtPWeXj8U
ntW2QrdGJqy77V2Gt7DD2W/1t4COJWX/tQDK2Uram7/67E+1uNZG/VCoSj70
vFwCy6hG4D2t59d5ByV7ZO4iB5/FQJOrYNGM34kLouArDdeJVgQ5K+UPYD2z
MPEthI44UMDM551kDQUWDdmwh49Wh/xHk+0Hjfsj7rGjaHXlZEIl574QGNmr
MtzTMFwnbtFAF1q45RUmAgB/gK1tn78fdFe2tyqgJcX8oTM5/JEaB/zrBCGM
SWE/8CGxco33SP5IZB2gWBeWGgyseXoS25Il7qGuQagw6e9lLwxOspVE5mOo
ck3nBdKqMZcag31Oy14puLBpF+vJ5mOQRTeBN5CUympJJHZrbngpBUniUaRO
lUCykDN+qgM+0ylUGr7vhmJYTc9sHhprttgR1kZu3wLa9TT0pYu1+iEpCafO
w8UiYmKjJfNPowylOIcmv+HLsNyi1RIz1H3MLwVaaynZSmtVxNPuQ6zDOElM
HfcwukRBwZdqXC2cmpLiGppfcksYIGIAQNVoPSB9fzLFMBcynotUKEu5ij4p
K0hBTJKOsmtNNUj+Th3bwB2C1ORHOAaLJol3+PEc2QBScakDnzPlrVGDu01D
6eipGJWn/RDfEGOUH0RLIoohAYYIk0+hTVdBc7TWGpjy3uRFN6+BtuOoRaJk
CDJ+kMOBZ0223pF7W/nDiasQFrG5dsRhApV6pIK4ym3Fyv6cCvAe642wdHVe
xuxkSHQnZrgXqwKR3y8g1z3OuNyGPyWrSk5Rro4Mb93ouyP7ZliDz8/rY0j0
Zp5+deVfeY2POXcS6evYIsBs87BBht+A3Ww7Gdt7LxfQ95jHGyiSbXchGbbC
n/l2za4pOQPUUnUBJ5ZWT5su9Y559ErYGujUjpKn/1OQPv+KoVhLBbWL/Xaf
K4CNW3CzQa7y0/0Ys05++jGhip4k91gwMq4aSOYY+xuuX0cFr0shVCEPViUz
1DFqURBgY7KXgHvC4ru07p5xFpbPAcJBZPPzFC7KR/VLw0Ut4tI7XdubpVcZ
SRdOkSZvwwVttNM5UCkFdeRPCDCNsrKlDj1vIOfwT8eZ/Do6sHumsPK3+qVr
9aA5SAJ5Pf9U2D0SeIcEPOYiCdA0XQL3/f4HOlBWFc/LAnOxOPiy5DXnDVi1
TqWepZlrfpQ9LOmhdXarCeTFziFLHBYDB6tshANZ7LzBA1DPKaxjbDAPjpYo
mXs4vJdmxuROu4jLluk/ortW/uRdzof/yPs4+gkD3DrLTgNDHYeyY3Hrtuto
tQkzQoDrE529bCQtvgFMgzay4WTDplB3aERTgTNFj+WopIRIMeFQO7s88opL
1wiF3RRHiWV7m4UIhPvIh8G67/5jelVJRyNi5YnudsbUuIOJuV9opA3a7zmk
hbICmHj64QZlTyQ5uWX8hPoGIOTQGDO3zgD9Spo3c6mgIkaBxKcw8KFxciZS
BXbOplvf3a5WyKgrRICt2IjML8zRVbaST+2AvOdMN5d4eqgfLzH6L0VE8015
DhPeRKEEXJPjzieotgzpUtvcdbdmsKPIPkbJg5SFA+HiGSKKAo008sQD4wyf
Mhx+32SnsDzywIQ+x/k1E8tciqaY7MkFupZvhANBtnOZDZX1rJ/xFPZImMS1
/ZH5G/W3n3S4EIN4ejhfFkiSkZFSp/REoWpdT2hXlrUnts4fjaQnnYHmtSCA
xJSZnFp2V07X28QLcmA+xzhAL4YTjmgk6XZ7ZuXQ8woFDv859O/Qg7VBdCPv
4Q0JlYT1Ec2fFt1vxkSEwGj/STpPP+j6+1qpKg/EvmmeU0FI5OpcxgwELBv7
epBkLjTGnPh06d9m6oP9+ne1vVd653Fzy06BkXhkj9queNgHpVt8U1Voi5Xg
Ql+TdhZtF+xa/K9TMT42kB71btOX1D/TtKKEv39L7cmjg7sBN3HbTy7BpsYS
WzavdXZ40Wahh/CaFeT6C6Nn///hAmM65FUHdHJEHT6OLN8W9N88iKIZ+NyQ
ilOfNbXW6dGXl7kvkt7Jh/dCM3HGuLdfrMVg2wUNky7GGD7MC9whq0wDftFs
M6J2n55ZlGCfKKUyd5hUAMdLtIv8m8eqv9ihTs5Ss9yN2MIMWTx9g2OyVAXi
DIRVX315Q0PxfVxbnfxx0xxcdAaRih1HRMoDaioLqA8RPWWX8qqHGxkMvC9J
ji1go9dfVKsNZmpyZibfay1CEpZTojG+amUeJlDjOGGS3bSN5RNFni1uYye3
b86EWaLcePOF4Rh7T8UvZJQ4CVn/JtMNIMyl5gZmFGLkA3w9++uKLukFbPva
T8ZjQ5e9XP3nKIak6uPebi1RVnTKQgKOKVLRTCAI8uov+hpk6W96Qtsoxna9
38IKFycHGMLvRMqjXOG7PwiGwnxZLTuqHKUlLBHbw0etudHCBNmnn1WW9I1f
TgBIn/FbPL8xy//4TwP1i0YeJvyn+jfkx7gHp0Uq/RQ79SnVH/FSGgWe8vhv
1wBLb8jJQJFc+shetV13RpRAeEyBjku+tsJ036bK0ck8tClX1kkJWhpEgtxo
0QzBBOwHTFvdcWDHMdGi9Bp5l5GdE58Gsm4fxx++ZGBmNzG26CHPXY0D/K16
2yhLjV1l2dRg9RO+hEV8ZWTmDambZWOKlgKUgCrLsb6maWD65LiLEtvEpbBm
bbUO09kdJD4/Km2M5Bwwo+xd5L416JsoXhTR9K8LBj9xJduURg6H2DFQLSrB
0zDvRsDv5de1w+cEUX65kIG0Q4hJy5GomkpZGRg+fd+LIeroUMOC0g2LCT8l
3A31HwHiMSJBiDDCXq0dfGTOJ9nrhkDvx//xHxJYs2mP+V3fNV5aUymK1TEY
zWP3NfZXovG+0YGSvhYWd150yaEb+IU/3KhYVxyDByKpXUR7NP72uc0a2jbP
Wh6p4evGOYSEGRrHSRRNONTm+Dk/ozQd8Anmn2NJjLPW+Le6jD75BFLm78FI
hOh3ztRxO0CODNn1ePW/PfouPHjbWbU8BqzVk82HXXfKxe1D6v6kVZUSsK50
Y/OiPccMkQD3uC8vQZ4FL9i3zY4/WfUWshT3DKKrxFvLpX1s4/VOSOVE9p+w
lEw9WS5e1bX7WVqSwBVci4kUw/rAQFcW7kWhGYpNxLuQPBf4X3JivwX0IAIt
X2Sqg2tx5r8zrRMs82sJOCmvCuDhYDKDCPi24j+LJFrxie1VBoohhmXc9DyU
FurXNgltIj9QL1x8Itj+aLDUakVKZEcUirsAeJe1Rm/GbQGHOx4Fkc9jkjx3
Rh9cHkLzIsbz0Yn02yFOJGa5gNHAsqyb726GkoyYwP9kpl088+XbXS6dBE4+
+rZsENIsBx7lHAgSXaBeMTm/XfSK22sf8PcJLjQ+olA28xQ6kdmGqQrcqNXY
DFChbSdVt/+FA9fRRbRIMVS5lt36w5o5wiWWEyZ0eIQ/UD7nI/xfXl6I4B8b
yTC3Vsyyj5UNM/lPagjGS/xgy0no7UegA0a69pR/1KwP8jHuycgSB63sl6sD
N747TDteBQt9X5zgo0JRt9U8WJjjevdAXm5AFM7ceYrkQlvAFns8U3DwiHpr
TLOjDKHIqbtN0wJ3MCuCqGk947MzwRVZCFjYNu1oakPhpgMX+YBvtGWotOtV
weljTwQXVRuajiNU5koHlE1DUoJBrrRXz2c9pnEJM5JPqmcRvmgk1R2ggDXL
7C9EegS2u30jryLWF4SFE63EHGw85OJ+4vFXTdcF/EaBc7u6R+Rpj28VxN5X
q6EdfbIr6dPURSXoWq4Ig8qSMjjsX/ezamq1+3qRJRJGPoO6+NKBVRI6c441
gtYr2hdUiJm84Neg8WosKrFC2V5kyehI2fUK1SolK5EL7tLok1LBR9OD3IIW
TZIxw1bn6WOq0/vGmgTZmSlLwouz5/KAT1Ex6W8HYrCd/iAcdMLcngemSkVh
uYVWhc08R2RHL/kexAax5JpT6c7l1luNRnjAEwUS4V+U32fR9EMC6TJC3g3w
ldHUSb5ygR4v16YSjhVwpzzg0hQz9BWfanZ8AVx/ln3mO7Eh0HXGI7eyY63q
CRh6gSNJCxVto88Attp5eHWagnn+f3U1ItHDJqUibwE6tDNKREnQbCP5ZVVO
bs6knLhEmd99KrMog14efeEoNRyaJOuJlbUqBLzFjmVB5a0S216ZH3hKfGuv
cPsMCpaa39GFi5sBo5r/rv5KYf2g3VZsKV8Qz3KD++xy3xKvd19cIUcKeX1u
q0GrICQGaMq7OaF98f21qMTF9FfY/qLy8d1mXbj0xR+EdhaLYFfVgCJsmRvR
unoJYBI/77yTQuUQ248wgZogRvaJD80zwxv9bS6gAZdh7g6SHl1kNQ2qd4x1
GWeoVRxtEPUiqqBACRGc+DJpqLg8+6SxLVsmYE3uj2WTCGvkAup10gYOfU47
BQ/2ooSsydr/ytkPcoZIYhQ2gwTIR0IJWvm3WQHuoE1sWwCRxSRY76ECh8V1
yBRyTHbfwZk7uy8cIo0IPQMP8QbyDbulerZhOj6EPoL6yPG0/BsPfrgaFmLq
5vSpgla8RZDXxIgDjytStmxrp1LPMgvaT5DGtn17pnPZoMHFGw/gJeUpsFrt
EbN3opQ7mtyhQlpVsBe8SVNobMNx/fL4bgB2AhKiqGKiGGuUkNJVRlciBbCQ
K0pZtPt2nl5fBm+MXxWhuEGv07FPb1X3UoUetVj2DcyP3ElhH6/uUrl04c3b
+F1r7zRXtK8qPd7yQHBXYvtPTKFKlj2KZY0M0TVcDQgaGaOzqahzQGc4AnvJ
NJehw36KFz0Z8TB72GCAsGVuvnXtz/k3ZtZFfmcPIvC4JsUKKiQx4xl3hm9T
mWHZlsZ5GU/aPkmZIm3rtUL1l5pmu4Ph4mGS44AQ+dZGGRE/lod/Pv4VV9gp
GJXRTlVEJXIRh8VHYB5mRF3cQ1TEGnh95J0zPhOg9KRhGQdFf7XPJFFsGBis
3ulVVipACIZXGxxXPJOyqhBsfLUvsZhVX98tThNfRR/lkZkPgMCztU7ux53s
hVVhQajGKFWLh4uA4efFU2BjpHekSV0lciBfkFYxxm64Fy2+uO84ZfwP7sNU
WoBbJa2CyzSSNNdWSIYbpuGJJm4C5Mzc0x/p17JfdTZuJKSCNXQDk8uQDuZ5
8dDT7hDIiRAwBBQfemK6jOnXAw+jXT8Y66hmB50YQUhceR55U0Z2Jw/hcHGJ
f7Xu3YiG7Pj21B7FzF/Qr0JdpugwHbA8XEEWP42K5aheWCD+ENw0ONEE1WET
mbXk7IIf9TGTp/aVt4C/ejO2EXJIVM3mDOUp/YG+w9lZGs+VHxmq0KNlrkvI
JUB/N5IvnUj0ozXqa4YXUeH3kZOPb4cmLqLyD+OuanTn3Zr1hy4iVSkytsET
wPspbLF2A/0bmOg1qKHIfmBwm/EkaDGjkYUM/wJWDEE5P+mVF5yuEp/QR9QQ
FkKp8ZjoUmtt7wwizdvUe1CN2LQC7BxeeZcDXFNeZabwlWNFkMRgITm4wywA
Yp5GJvCzC61YUeQ6SBpRsgDkr6b5sM2OOGGbn++G3nNLVWdM085U57BKNFKx
nXvOSYSA325gebAMAVkRy5aK7Y92KByUyr1L+JM8i0DOVQwwKADk7qO2BPq6
lJp/9TYlPOvzXcTS6IaiHVB8q68715D0JazYQ/83LIDPMem2SZPNLsecmPtP
qyqnXZdm269PaRM5hTy1LDVDCQAo+geKyu1m7e8iDwYA1aQ7xB6P0ZpVjo6W
kdBskTrAWrkZKzMr3158Yd/iz2V5LxYr/ofI//zTV/MxGyCLTkRt41iPfxby
bi08htnwVKK5Wa55BOmpVA72CIFp2w+20YL0j9jhKqenaRUaOR6xTwUIH7ED
QcG5poDM8BQJYFfYJiYT02sHBKjmSxIdjL05kS5Y3LMqtdQa1Ix+xII/b/AG
sMVGegQ2jtxPRMVLb4wppb98sdDNTCdj241tNvcMJA5i22C0Bgs9gMlaARc9
NSt0R8hlVr2Fq1aXGjNYyaQkLDr7O2hk5LgFvmXpluGW+w3NmmjbcnIFuJO5
znjbBiLJ4x/9/wcyhZoDwebIj2NFi0owGj2tRgjmEb1eYDm9RWBbQj0dHi1r
bEFE/pUJ7/hRqqEfhSk3wCMbv0v7v50RjZa2uYOkoLylqI+vZbGgVbkLr8nP
/j11+FJKKlR21L6U4qUodhhRDC58GCjCSFfaxUMR4NbQaYFqdBIGwxPlFyZI
I0gLZ2slSpwZEWRX9L3jzjMqsb4M8DROTET70KrFexEN6BbYfJRU5b5jFcRv
Cb5lbOxg3gwJqcHB7zu1IF/OyTJHQtmN4sI5csupqVew81scN4JRTabpafaw
b3ZFOd3dh5kehJgD+tQYS6iJ5cWgH/9CzGXeSuGzNCJVJha6cAmZwB+05Uf/
16rd+4vLhKvRX8m/RlzO/0FGyEZOZ+FCuUOrKZlcn4yw3JYPQ7QIEfZ9ovU+
WN6pnBhqC6Ws1YfYM0aJHaN+tT0SOE3g3Gv4cBqdFqSn1mjXD3ic5WEgxkNU
NqhA4CpV0x+QxDu39ImS9HctnaWdZcimbr4EJN/XSmUaeYue1h8ts+yKyY9I
Ic8/l3lA6QC2YNoYbLcolcPdZsRioYLRTnzpNI6492WGjTQdDr/0OJ8IYJGt
pI8EIyanS6Zr2yQ9CDz08B2Q0vEtlmFQHOG3pHeElV36owYWfSYbeXGVvQ6Z
8rmZB6EvwxJUkk/duEduAFz7vjEH3v6IVCkDZ+c50rLJCH8NMN34i02Ea/VS
3iJ1M3KyCuKowWJ7KXflhgUPGtX9IoXK32JpovWWgoQ4c9ExZ+8gxNPWxeYf
8gLe5l35c5v4r5kb/dkac7nyhnmstPM7WrVEGr5nGH6b7iLHXAMm5k/j5E/7
CzMKb95ADTo8uefSrhV4kv+5BlFjDcvkuMWPtfe+TlcnW8wJybfg114ROBDd
NoqBHOo+qbvJwtG1jwCu/kL72BBZpi0ptkSJ4TToAWuMOKPtuMWRf+jCuv/M
U9wyIl9b9JPivj+KmIx/tY4y/E71OFLYMSV4fsfgPn1oqu/s1IuFZF0psu/y
gBMj+GKK61BWLBXxD0bejDFfPr9zQIyWyn3t+IPVgIbikYubd3Vat/t5yJkT
lwIyilfTByVqp+rWUb1RNekU1eEEI77Dj/8W2cpTQSoELaISMeJlalg6cJwT
iy4uF6ENgms6gLkDMDxu3st/bMYjJeoXF8Utu8WMxx/HI4qyadpSQEVKN2Gp
WFinrHwKybcETuOE00oPJbvICmojze+sROHK6Isv9ES9n3KtOpv1nSsRmErB
POL8davzG9JNozak8b3EJbFY0e/49HUySq8kUi69kciTHxOlKFTDljEuSmV1
8MdbcNsJ/hyBOVWH1Sbqib7PBGilInc9sXPNurHfjGr7BCPEf4QVc7YmlWrf
VRyKQup1WH2KJkPZZXkLninUr5zFjR3iwg6SlsKaSrTK7Zyo4LYFX36idoDP
AtCQ/KkRF5C3fS1WzTkAUjfdAzlVQ7q5AHaporwuROHRsSsEviglUAjcKr45
MFqjuRIJzmQzB8t4xWbfUmx+ezGrBkC5kW15gBtVEMxE/CjtxeD+H1K9UwyF
9ugsiKBB7Psk+Qx4d0ZQvSnC8eraXN/QTmx+VVHHSWAzYycNDwv2vzlE9qL8
mpIYk9EJ3CgvXlpHeLEEA2Sxo7rJIkBbdjIq6dbyJVAZAWOghrly8t0qIJrz
OAQg8CT1nWU5d6R+X9G5o2H0Qt7+BYQCwXCAF1ItcUiJ18fEbWhxSnFWsHz4
jWFoq5ZrLF3nOxjWn4MB8dJr4baZF10wdAUm2qeCZoX65HHLz7BCnrftCp8Z
081xeFLMMxkO14jOr+a1IlV7P+/l+Hi7l3UclJtH8kvl+k+6EDpmkpU0xr0B
sx/PuTz+9m6YhAdoMUZ/DHJ+hLQGFGSqrCMZEI9qnHux7aWy/da+w457I92E
qf44OKxoBaXbJTIRFC0KWx0ELEaLrehwxrxNUWIv9J11xLcwPxRGPywmQs6x
tl5ECG0tU5ko0anMeMmIj3KCJBD5K9JtTW/GMtuGG50xK1UbSRDY1Zdc1s5d
jrtKY5ghb9pdLs1V4XdfCcfucfjNq5R6NDIkrwH3myfA2MxhLfsNhTiFcbpm
4KZB95OeCo/0/ooyBXMJ6LQsQ1WkuomuN/S+m6StDKSTM1CjD0s3R0MerppY
OXQ1iSjDFWgsXH5wWiZYI5KjJzwd9ViI5696gxJYmUy3eecZcqUONDR/ZK/T
JgiuqE4uFzxWSLEXwPGXXTSHgwXZpjPeL6FZUR8/eTuMO/Vbo5YIw1eQnRHp
iGPg7gPXRHmNlj1SBWm9Zfcw6CiqllEonN1qOeW21BzLSzyHvT1NIobvPW7D
w+upkjJoVOlndsGi10f9pp4WHchOjQ+om8cmeEPplEiWDpC5c580jH16OYoa
WuyRavopAXOXWbj4S+ojm3gam0HFIbjFMsZVsf5aftrod6b3zlmYL3oEOqOx
Umi3jq7wPZhwl5Y2vm7XfTa2p/RPq5NtuhvkDsWBM19KFkR17iRZp/3ph6u6
y2zkKouiG0h/qKK5cqkislSNCIdhtfPM3Ql/0VaFdVqiD+LAfDIRVZ8Ny9vE
dxGzVX5dcBEDhr8FHRirRbbdKZSOCZZaI20Svv615+xKYQwGB3/En1BKERoh
s1S4AbXDKBBKpbp8cy45z0phqz1SJjMND00lTD7zziaqPRj8dhj1oLMeFHd3
RnnkY8deT2JeCOA8khqz8NcgqxuUico3MXrWeNSHZ+YqPKTfIEHSGFu5Z6we
EWeiUuoy/yJMkFTq32CuWGe7krA4pli5tsRI3NxljyUHZV8lw1O1ih3Ss48m
1XNFohjtVcdLiZ1DN5oC9kPg8ADDA4tU2LQ0dvnwrc9cK4M5umIVlMgMlSQV
0Y52nrpLedjHS4d/K62NaFtR4JfpgLGrMrr+wtSa/8oWkmdEIffOw2dCm9y4
mBfTK1F2TU9nBT0Ir85s2Et4gU7zj5AeCAPrsEAmLro2WklNG+1YlkdvBNNJ
XIkDHLmByd64WrOQVpOgV9S3EjLQtGozQWI/samnO2kd7Fgh/vW8lLOWnREF
/eLvLCUBZ2eC7sboEJWU8a0z/CR9QmMI1UIpxW97O669RFkkYIl5/QYFPwGS
Jgq++3FeL+6nIe17tdj8CKofZjZfMcW7Tz8+m20+SBkpmoQck0EdeirblAIv
HpVot0TaZEWYxoLW5eYjiPUrtzZRELvMIoOPFGtN74rpev4um+Lqgcez1m09
A4AQcj4ILOLSgl1LHuJvaEaLQKwm4OP6yzeCeszdOW7PqAkXsVBleNyhO+tv
onkF0rRfnNM0/mkqL+4+jNvhSeOIqYzo5w+sfbfwDKodY2fSCpHAvi03Jepv
W3DMmh2JR0Tx+WUdR4sz5Ajh66ZQl/3HItgrOuJ8GiWQZj7RQInQyFYjLoqv
Y4Iw84WhNUwuJyQTdoTPoD04IZSkT+OpcdFdeCaJ8TJs/0+a6DVgmVkdvPZv
wKb88ujVR8CvBlfpYJM/Fala0I0TMSqFZKioGbskfIhSNYfkcRdMRllO3LQY
cMkALSO2dpYj9V8QFAvIaGVYK8YRESZPKTPVD5ZylmM5bWcu+g2ZUev8AyRV
+skBmqmrwkMmqFqfaDfNZeVldpPQKCErDAjKt6O6Et5aUIQEHMmMjjr/i4po
SnnHtt0tr8jboiPW0sj9KMGz8cs8QHh1kugF3VxuIPVe+/bXaEijuHj9Jm4s
s9eO8CffA4eNr4HfOd/1/7N0HPyw3FwWY39liEg82SS1F7drc8xl3nPbVFPk
R13wNEZBBuNaeYPi6OfZk9aNrppLINH7DFx6/omi+XRqLVfBgkg2rHmuktx5
BP30c7HYupMmAmqBeCAvM0WIuLksgpwlOpXxS+7k3N0f+xR+nh1Rh282toOW
5U8o+bv3TjdVE9YFbAAzHSeRyhrlThB02MJOhVG2Po/u+uaAG6Ck7P8+14MY
lZ6F5YBtPtrvQdEoNnQsA1RkV/kMHTtWxbHSR87R603IFtquCDU9PJqJ/q60
O6yt38vCTNA0FwwePSwpLfF2mU+8WX2Oan10FzuNjhfX/X4WTmijc9JXk/jo
PQddfEpPZ8ZyujLVuHQ9WlMdkOD/SDomcgzE9qpLCyHH4doRAqNiDqQil+Vx
Bi4sgPu4sTChkHf1bofrWhAvdIZtBH5b4gALkOKM/FsDdrGXKHUF5Onm+n4N
jZX1DCNwqTx+A2r3VCm8APu9oQcBbhxhyicPAOQn7iqDZspdYy18VSam095B
0nzzyyvyV4lin0Cr2PTsehzhl/14fsWhEmcAN1GHHJwBY80w+P/O1hTBNm6t
GIpnITE0HeQL9+SWRaB4mkjUGuEkdA/IvVQMBZIWc/NgGnPe8Dir8ffZmJat
19+m4r1+cAyEdICIMQvb0Myse64DJkV1+oejYRbtLfW/Oxp23mIIWHxuNvhh
STAWQWa2o6ZcBfygGtr/FLRpINuWLMkigYekAHzBOJBWvJzm0lm/D9ch4XCM
VQ63zFvYNbAN/VUtl3o7dZ8PuzNGQgqOLxFZQF4UcQvEwstw3ajqKbPMulXt
yG8w6SKxqYDTi9vZc4I78Kvy+LDIUrXPdOy7Qi9sAFuJWNhbKkRhhYb3wdeE
hzezcDRYpFFu+/gwmnFsO917YQ8tADOzu9lJfBHWrhkgy2AeU8iQlz23jsXU
m5oSENf0LD6yoHGvtKKyKjHGoNMGyCTUy4FTrCOdw7BwoDAB6bx0mwr9YiUZ
x5lRibn9MOZdwwlngV8DWaEbnKAPx19maSnuU24Me/o0gaa4t8+Rgd6QBvwv
+5oN6Nx+WUoPb8DYJtCzoVdwZfO974VuNBUoUWb6fBREAgsA/P2GIch691eW
Y+I4LDjaDVNtayADFq8e2YOzLyVQ+56+4sPlz/04a/p/yal536llZzhp1Xu1
Li5mkiC4f1/ZR8pfUJ4GFaqWfFkXA7AVTwawY/0bIrfqTvgCuhyTiy/UgpUf
YWMCwU9yG0iOfCLNHUKnOeeEU4hU3cFITCWoVcoYPVyF75cwC0HWJzHWoeBl
rHRugC0W6q9zDbm4welub4Ad++yaw+iq/E5TKOAQ6x8oH8AdFUNImaL8+TWI
FbHUughOevnOXNpOS8S6upI6lSbuaxakQciymNUXylXacyefOZ3VrjVVoatN
BhBgLih3blFW28evhGUrZkLzGP9qCgE7MVPYh2Jx9ekqOzmdEsV4N3xL5ODR
DFlpG/VDzugWpKuUCSQfaY3O/nMnBpXjhYH5OdCCog5/BVhlaaMuan0bfwid
NFHFHnfmMC3K7WozRBgL1G2xztoDtUMV/n9aNOthHbOlbO3vrLzWnnde5nEt
nuJFrad+aDMJ5xlPizJDfJbOsLDNPI4lWA0lW9ItJv7/Gxjl+nsUzMClw6gd
EHx83W1ryiEdC2V/QJhmHcNE++Jjf1ONQxkq8DvtLSZnzyngqqMk9d5IA3Tb
JI7lDgCsiFMq99uRZ8u2clIpcvGkMCyi8hHdwz6FGzAsAk7rCNE20iTSbXSc
OeYifqoABd6XQE2yBcGkRvS2Th9humJk6zN/hT9+nTDO3RIfU4f4/BWYYmPW
5R+eh3nUoFMZLP3eKq0yFzZkZ3lb9IGfUUj0s4KSlp9TB0pt/PWX8BHPHuQr
YHSxdcpPxuN/3p+Rk//ddYqbuHeXWJmKnhU/wRMxcXvSqVij2NpH03U/8zFk
WkyVhPZWVrrQUknuukMC6tcwanBQHIFat9jdw6y+KiPUMyLcNWQVdAjKIx81
W01Q5uRio49mRFbrYay0dKPo61T7ban7yXrMs9OInhlo0Msf/jhuH3FVkZXY
EKmuTlhqwcXUQOwQ94/DCpVoiWqAXdhVn9VUWTl7+3md8v+IYdhYm9WlNHjX
30x2i1ZZgdZZ90nS+UJ3K1vUuwiAHsDq5KyGf1HQDe7X2/NtECwSLfggaEju
37MfNtCXebXIWixANIGIXE5HR6AChT5Mi68d6okz8VLbRP85zXTGjOUuctty
Oo5rkvVM0BWzhIfToAi9m8hpGGQtAvEjO32TUmHiTdacu8nFVUHvrW8afRI1
wul4aEFXXYkviDdz2TuB/VkkOxIH2NVSre1+R5IwH9cEwfp2FEGyCFD8Dd0g
XaTkwN3ivrHCu7txph9CWvgsT+5NWkyAi2LhkOAWQtUIPpjQnAE/U69t+wOr
X69+ln+6HHpGwQ5xnFdsqJODUtQVzZZrQnS5n+yAxdwH8lTfq178oLJHasZC
Pu+9NMQczM5KlIVrkSyHrkBaBNA+34AvKCMhXym/tfOwVJElYvApvdUytsqa
MXECrQzHhZzsF4DUWT727oKqBjoDibUTrwLtY6fBxu0lNRgVKBSGrEA3wFBM
fgxU4Pnu32yR8+HS0hOy76kvs7cQ+3EdhoJBvYzmqVrUXCJTWDo//IHaJoW6
JmCwasQun1Xwqnz6uPvq1UFWHdKojeFFxbW9zbUffUi02z/kUh3It78KtbtK
rnKyKgRlW38GmmdzUEwPWgVVuaTMfbkMHuEh1cHNw3PdLgliLs7cifiqlA5m
VaZjXmLET67rexome5otHY/GtkeJOAbzkMswVLMkSLHtiVY8ZLlWuByhm4Uf
3WSJwaViOB06oM+rjtKIQi8I+zy9r7gLa/VCXopsMZHufWg4gUIiwEZTAgNp
08FJ+SRBXeIALIoDbh5+XOhCHm+Ln2tyNpYFCHkP0t4EfZtpCn3OZbEPGs06
YUJ+YE5U9mZiWSyIOSV4U4legKftFKEh1JQjbgNoXv4MwfchueN6P+uq+phQ
lBedmjTKvlxeewzwyphDQeLd0G0RERYLo1eK7V58fQVJPv1rK1DMBnzp1Lm7
grJAul5TnHPzZ4397aCCRuVmcJY7r6l72nPr7vmWb+XOQgAP9X79ojpchTkg
M2sblQOxOYCZX3ioRZweFDaK9wBkgeyP5xW/Ui/Si4QPWLHlOMAlRXyIPD/a
cz6SQA26fT400R9+MgdrtaKlU15TsbcRDQrzt8+1OwYErfwM0Y4C7VJnR+Ix
heLdgLZn3nMtM/HP5gTrDgtRhMEDDPasZI4WN8H5haxZfVJH8+kPilC2b84b
y5a21nugtcEdK1pEfYqyvy8xQWXp7bFFD0RIBpaqQvBQ2DELj1IiqikY9MeB
bthJR6Lwf61S2XF4FTJ63/wk+W36IKbE4rHTRW+R7LYNdZdKxT0Fffx93rrS
HJBX+v1ezwpFpot21er+p5xItxAfxWvEsrbMqhOt3eiCjwJlAbqapwHnu5oX
1Q2Nb07Ib0iP1S3EzZNOlL/0UNhyEDBBHZ0ZPu3SBojXq+rE02QJtXHwjNFx
H3dZ/diUq0KWh5FlUHZlc++Kjp57c5agb/hHbUu9DYdjaqkxentp5erKzqNH
WiQo8T0b7sECG29thvdmgSWmrAX8Xf2hYLN4HwsziNed2xOci5kidGvFFj61
bIzkEE2PuvgBK6e75twU8S16ARaSkKvgs9ZBCDhzPOcBVGfLgMzuUj2yN+hu
hdLIkoBZM9GuWSF5K3mzawUSmySNuQ+A8/vu1LUSiWk6nMOr0H5MFQN8pK7w
wFVQW0btkx8E7pB3DyxjgiDK8qzGGfoj8MnBRqIC89GDFRTCeV7HEtqSot7X
b81s5y3ZgCdZCL4MNKFyYxb5rwb3K6Z0OT2aFgIWPOrPl4f4jwEvEngUmZ5V
JsfaC0JEx3Kb8ELr2nxphCkoy4/bSRNjZkiE7lI1TydMS+A7S4jdDk6gD09R
DfSsfX878+r2NDYec0VO+eLTPL7U61vECx2mWP4XPnARMHv7xd2MSRuDphBG
QoIlB5yWUYJyIRuNNlB/pl5YZ495NsZQ3tOo4HapfUh2gWPlm/KgPKFPcB7O
/3M0GiajVMWckMJTabwS1h1eD/Bc9d99PzgEvqeS6b2SWcjeH9Pvao7eKyYQ
3K8VUP1TX3vA8YbFhGC3u9nGQq59kVM46piRJjpllYnhQPodVeu14pmtc0Jw
CUUnXFdgj0dEl7DX//RnSFhvDyvOvfB/SH4OTPV8biQCyuIsJDYoWeoFe5Ld
gzChI1nIrnE1tbjX2XhvRleTWgwO/DIqWfBjZbOSBsmUuIVLskNqN4hAS4bv
V5xxPWwHjsEO1WTPR8ooewK+4tSsxwXAAgn/x3H1gP6fAtPUoYvd87XrF/Ho
7XHU9oR76kO5w7P01ZOz9Y1J9Wj4pyXV01xJDlOzEOgdpLBM36p6K8V9ZLWL
YCFDwBQqgQaHH6YVLIrWSacRBH/JUNqdbrbAjYl370Mww0ZxYEmLV69bU9dM
iAoBu6R72+Mlk8QEb62r96+hzViWKwkbx51naGSqbRMUYZgA03q9IUZpi0BD
EUrwjDSirVvn78mbcXq9n6jKDBVy9pUgg5suBCgouTr+FAHudreSQlHeqpPI
Rfn/PK3exKdi/B70Hxm6QOavV5Epkt8GLJgWRaEekoIga2TAiGHpdGv/uv1L
9xFnDctXw1Elge43EQhzg4RogBB7FlADeIZNDi60N8OCXVW956NjqK7yv3fF
MbKdpBiYmJb5JUivg8rFGHBzOQE1yJO52QAWPF7CjpYH0fk3qfn38PDhEM6N
1OSOtpg3foF3ZOwmpPeHW62qMYvNVddbDvxiwkC9D/a3FZy4s5aOuQ9FKyMO
7QOJiIouLCXD6eBrYktZXLZziCU56f5RbaJE3hrZSWJlgWTJmKwd25gXQEaU
Q0CIdM5+jFysmZTuQgBqesGhJM8UtGNGGbBxG7CAOKNHTOJPg004SV+OBOUI
fpbyOWwBojHIDAw0ZJ5+sWR93CDeedsFISO0tk+XmlH41G6q/7RxZicrV0UY
ohWJR5+dARg4KAOJvD7U3yIZrJ0oj7/nXSAAnu0O/36eupcXXtmTDYhtaj8Y
2pjMTcU5UtAJd8CrTHeyvB8EKkG87nm5je8DdsujakL6z4csHG0bW31SD25I
ecmgtdyQpgfZqPvdC6e4sX5TIYtjBXdfYCtyoy0n/Fuid2sb7qyejni9GTz4
f8yNlE0i7o2arlJWu9x8CFu3Dm2I1wh6H0bLgbz7V3jb1kEzmhV9YDQRxyYC
JV6SuRrxBXALKFP5hgGWEbtyuadvUp14NXOFmVuO6hlB8FojMKks6HzZvu2/
ir48dAuCM/DxaR5HliqISCJIRfDGbVgnZ+zS/y2mifG9Um4UHkh3Fz00U1Ew
fQqr8FoxZ9jeJB68Q7BQ3w9X/lXeFoyE5OGIkypkggxFySUA8GyxKVCCzh2S
STd39iUHwGZM7nqo7MiZYYkTVaBmhwNSfazKqfhETR23/frvRqCVEy7G7Pn3
uMEJNdq7THr3qemc5pkyoX4pfa/K0wVObZK7Cyo5vOrjcDL6WwhRQMLT4Utw
PQosi9FshWYMKVvzfRDVVnbZDtMyJOMw0ylR8M6jwJjTCRf+VswDiYr0wHxQ
f1ijr+stADPnMidi4CZRxz59hU1UnEsf19z51eznzAPZWze/DKF6ZB+5a6kW
OUNS326yLo4AkAsUJauuf2tLtjgmE3RfrDTiNQrnC4ucx7nclagkNgxYhYkl
14YKbbUv+nWi55shA62LITbtv9j605u+UcnN6x0nBBvvAa0KDuI2wLkq3hyn
iWWexNWDVzSpqdsOQW68aqbcv6KLbRLJKjC2tsYfS0icMyeUQ8lsZ158TkjC
wwm9XkvHXmcjrC7EdyB04o26QZbK6iu9DAFMWKBuqOSJFsd1FNyYlcLr3n6Z
nWYHl5bzuo8oa66Rn2TJNglP8lZrj6xXc9f+YgvQL2uEcXgLQj9MUltNKiJA
jtNMvSMqKaQyLQXitrk+9LWT4/NAO4cS6rvLUfrCJWKdsHPTMjErxB3XPVwO
BbCtWEoggQ5KTdGsRDAD4Duyy+0R0Y7psuWLvC3yxOOMTiQyG/J721wxJZIl
C1L+df6MruBymZDgsSfSnpQuQ5HCr34+bcqfIzgtcN6M87MOsxCTCq7VKaaJ
Ui8NSSJOmHK6L9LgMOWixtr5kRWtKKqmQAlZ5t4yCGPB7BzyYFEs/ozFY5Pu
xYRgf/qLrlsu3SzJdh9zRVTOwDIoVaZL2y6yuIWwBtvdQ4hp7COW5ReiN8Wi
VXyysA7/W4xzStoNe7mX5ho+nMdT7LqMLcNMBMXejMuGoW5YupUTIMq09Trw
BexYjjxMiCSloxYsNZxvruVbdXG2ToNG96YxpRU25N7vhayujpUh2svJe2ZY
rsm7fd3P7rAlG3Ws+s0J8JgW41VmLd0iHI2lUcvWBO74A0F1mza0tz7sxZdY
WvZpmpaRtLWCElhOxOJdQ+dOFO4t3FQPXzWP5twTBAcrc6HEonCN3pw0JE7s
BYPhx0m30YdFsansz+u3A92i2UC7OiOR+/PGkk4qYYetMh+wGysPM3pJE5ZE
Y64xAGrOJ2hoKW5tQ5iUxJWspf9tTS1EKIwUvkti3oZVva7j54k0o0twvJOA
O6QO1VOyWtoxrgdM5mxfuOdcrT45OKR9ZHVjP8IOCoWSy8QjJeOpTPS1BMeb
QNh+VnG6lj3+pRNHSRyYNi8Hdw+8jWfIDS650bt4f+f4Qzv0sPkaax1GPRhx
68sFviErnDCYRX6NORdKzPUZVAMQt6jrIXjGZ5rrJiw5iYMcCfXTy6RPzsMr
A4a24va1l4mzQvWEZs/eARKglG8CPV1Q10A/8LmtKMhPTvQUQFBitE6q/svd
pRoCxQhCsrP3ILY+ACVoFjzHLmlwXM88M7MgZifqX/75gSbfPsQLzFu3TZTO
YkohtEziiNVFUU6BLwm1lztqiTtVGCWuAmuUCs9Gj/1IaGnNm8G2tvyrPWCt
ej7zpurcATRaWIab1h2gE89PwCZMxkvqmtPgGnDmVAlYHwWAq15BVJrXirwI
YFh1YbElR69SYiFJIsrtStuoGggb2gvsLyJDz4EY+KeD3m/eZ3VCzxND+HNe
LSsIede1df81iCL6TqlECZG+BsvZdxJDkaXaDsw4CeJWfvqT5Bc3G4+bALlV
5QOhHO1tIuCMX1J3EDqYcss/Rksz0C6zmnNfg2R5l7Vu6C1ds49C0xllyVfr
w33fhfCrXrYSBjItGJLJRwyYOiMuFNCeh/pb7Tp1QEldUdCZRMK0J2X5Dl7s
8XZ/ixGl/MZ3h2OD+Fa/5GsFSfQvuJ2Y1+ZbHCy6hTs+KS7V4Ubc4cSSbnB9
ySHImFp27HkoGzrRgFgrkIBJAfzoCbpyteprywgU8dKKSaxOb4RkhYQ0lwUE
2lJ+isHk1jS41R5Asttcs/4BbPLKg8zELJ/efufVJ4VFcKHgECt23mk3AI4i
kQdHDyuEFTFuN+VT+ttQh7grphT28LBDm7kiwr/gSK5iUHgf+ocWjGly1imK
xL/8VZwxuzq331AyneXt0lnpId4yDNz09DAMkNdxNvZeRTcPZrhBNJRTv3aG
FV8LN5Cz5odCb1k4pOJARJNn5DoKvc0SRbWV5imvnIfhSURbQbEv2QvPnw6E
qVAxFeN35wVmPHFK5jsukMUjEmZqHoIqXL2Az5VLUzR507f1vlPPMgbHIjuC
s0MGH/a520fJnWUmv0WhuiVUfM1fUG0ADgTx1HlGEp6h2mAKsZOizXLXB8My
pojf5b0Ux2vs9iVDtQAPTLuLY4becQy+jULt0XD8Beb+OWjYutdmdckKVIWj
gorZS6FMEO2YSPFWVgo2WwOXxVfuH6VnvfWnTCZCoTBLkCOtzHzHlgRI1eCH
4Ye62nqzhTwR0mrJTync4uzrqUtLeYLFASVFiHMyMerunBJVxtc9mPtuak/c
6CoM+pehV9iepWzPo9EreYFV+GOHc2E59stGkDhanYeHeN65NQtaAA1aUr72
xW9+DPaLFu4bLq5wSR5chbCuHj5KU0F2eRwwhiAHJ7kqb2OLHjJ0/ejwSiAK
u9HeWFTzJZ7fv4P7i0QGFqNGnlERmktqll/nWhrsJSk9M+V0yX576Zc6tbFw
i49pVyQy9gV6vJeNfg/0Y20whcP6YyUN4HuyJG3ZPxZXlHOo5w+UDKLWN7Y1
gDgi7V+6iRTgcy83jjIINJJXM/FPnOy08WdJ7raaMH+uqiF9fpuCYRZi1zJ2
7jcu2uH8t10iLswHQS2FAf4AFMfBdCFeg19n4gvdNFYfmx0XDqOFpE0Ye3vN
GQOGIkBNtaecgnm499LOWGiguFTkVKrouvPeEez+ujf0RWYsmbnCk/j0DlCJ
5B/vKTFsw9rYIfMnCj5wrhKauqi3b3kgygyt6SdWKnsvCPy5M6QuT00EQk6j
qWlqxLkWcRwAoqs4HGqOijO7mJB7BYgcurpVyjznkiUdTKDWnrT+2qjoHBZa
lGv5ScRrwljSIKTz6ve9dE6aAxinOWWTUbbBEizm3tBPhl9eH/9gAj0Vy+vn
myfxfYPB10Li16pZNX+fn47IHNa1hTu8jAFGAdAUd0qWtYm1rR9GMTvBE61t
ABGQxuCWWQMEt20Q8PzBIOuXHh3sqvTbPfhpJOTpxLKTHEEsTu9zTYRZg5zh
uYfqPOxYhZgoKbTQAsIOXmUTpuhNgom1xmA7V5Ag8+X0ec9u6axpsjhvkC04
xYbB4gpSbOYU/cyS3eVkSbkr7EUt8uzvkJvahhWvxOcCpX6gTJ8KYOHTdGfl
wFyDORTSFtdD5V4uK27BINTz9TU8TpIPbF6ulF8zk3heL1fiMglQK/rD9cor
+wzVLf822w/vYX9Nul45hFq4qKOUEGF55BkvudTvFj5fQGcA5B+VpPKu/sOa
sOi6bIy9n0NAt47QaxHblIyZ/2S2sZt6W4JLON3N4xjcczUd7IylyAVBvR+K
qUwTq7S7MPlKGNj1q12jvKHD6BiWCgC3q3lMdALsOa9K7EC74dzQ8D1xliJN
+5dHY5jgGBsNoQ13p+AVI8OfQbpPweFJNz0WhK/FZPHdRjLfyrWpoWevBL4K
FRViPouNlLu9qLzkEWP8VhPvfhYktxD9m4uyyoGXP8aZ8+BoFiEWId66wznS
rKsZvnsY05f6qsel7edJUg+MrGAqandFpqrW0OHA8tdAxnX6gGf2r322LqAc
dgIorDNDa4BvO59+bsRVxN5kbXpFo31CHcrtUiZPHUa9bjZdEfrRanrBYAOa
x8OQmhnt2J9yp0GLzOyKINf7zT4ooUhJ5gBz1/P7lmh6taXN9VblFlTfhDG6
7ZfAbUftgzdXE0rfMoLzFlg8MTIx8xPPljikY4RIhoOnjlKg01I1n8/ZO2hz
VwHAGF1LRA4iVeJ0B/25gQL7aDxZJOlMQrtXkqHQWzd7m9iBBz2voKTxdYwz
XKk3ALQQ7C9bWyKYEJNw6vnNzx0vBkU2EZnIYc0baR5l/AOgVd+TZkkRIwVL
vFOdrVVJKEvrRl+Ff9OKEy3GfmycrojtifuoqKUnZQd4PPtcOHaENSnG+U2L
YjVrcMPeIRzHe6v8rZdE1VYL601EgXFETFYbskIdN1Hl0QcRu//AXAfqB2YD
k2lQ/u0kPCquXcMUlCzpgrft6Ms9tM16Je7URwev7aY97YOz8ATfQksfCxkX
vABJdBaIFinMKIuzXrwpPDb0BADt7jJNhdIjXAqKMgx4zB76DKWKHmvcPNWu
YaQ+Pdu4ilRh01S+LEHJrZ1wkLC4BVGzPPfiwr3OXYvhjbIPQ3yXvAE9ju4e
P7zF+fkyH2B2H3EbUXg8E8UPmuOHEqOUPBLbsnIAGS2XFNu3gI9oT6Bxzsif
/A95R+pz2B7BkXR+XQxwMaM4YyBCACQna7W4KSacckqhwHCr0I1Hi1zGl0Dh
3VtKejmqzRPDGCQHBbGShzFSWG60kOPXksXvq08x0DQ1bkNtgI+m2sJHesw+
fPuYuAwkXlYoBCGNjb6BYqPTJchitCMVpdOvgJtsbZglGHklM75oRlNbIUmF
D6Ov9x2D5U5hCeciVjhqRtDoHLEO4f+sXO4e5d4tmkoK+MYPXdlCwB+EpGkS
Ks5YLhv35tSqUJ6Cp61GMeJ6/GnxZMEouWCMoO+UIU2RpcyBYzxNoYQO3jrt
Qy0jbCFow12scZ0hiGARFVOeDEE0xkKGmz/PLRN1Aw/7WwDi+r6lCSXRHLHF
ABW16sWu+ZVhfvqYrsFORjsdoAIFGjg6EWpzNtiYGIEcCFLRueYen20oCj9e
14r/YNhDX/54A9Gk4oWeVrT6wtTmBT+n3FbpgjdXIgTdMMVW4akPrDpxFJmO
qmRKrcoJ84ErfwdVCZvpL5SCr+2FeOJWOOgZzqS7s1SrIlw/74KBOj8Vcsug
asnuQGZPqCq9maQfSEKMhP9ju0ztGkzJtAWI6ZFT0dbBqJUjwcHGNxRQ+WH3
7/wU+BwXrbAOXff4cUj+oZuqtydXF+N1k9K6OZRisdMGRedff+02V45v/o9W
J2n+IKso23KSgCnOoUJmbDtpnZSdZNb/vzv+TmCcxSKxmfH0UvmQAFwjZzjJ
Wvjkqy0WOjcAWvwzmcXC/pW0Qqx8rv8eyNQsGCzOVQzovCYciJfBxNQ/TsPV
htzGcKrBMxfeVd3qVxNrLavzBZfxBMoAy0kg1IpC6+m9F/mkeLhtmNUwphNr
csnvZ+gzr4Nu+RsHrHFzv/L1Za+KAAV3VYmvKF0VeLVeUFCJkttTdH5GTr3y
8pzmzgYtaeUrvJ1zMx3ANmtBf1FQZ37ftVXvAuTUdiTil1Ioh8AOploiGhzT
i/MzQcaXo9fbf5YxKBko1e31f3fJlD2okS/mtw4VqWRRhpqkGCYsv9ARDCOw
JNMlgK42cwZ/Pjpqhxs/HUa7f5ihMcWCFpowLtSyrZ0yq0QWRiRJx1xt6oJJ
wc9gqzicSKPPov9/jv9O2hhfnNRQfVuBb1Lu6v2IBbBVUWFblvddlBLPEsHJ
IrgCgJTuak8oNBxlm8H6SlY7sT/TfXbBbndtxl7vzRX/yRtWLY4V6b6+sWbc
vhNLXHeYXQksldh8Z7JHraXsqwT8/xDF9jTlEaxJGy0l3YXh7H86PE5ShE5F
gurBfDnbClwk15CMJlbWjVYHjDRdmchhYwwwHkKyT2rnpot6xUDaL7R59MWL
GJny9G6lRUQ4kLCzrKmMpxRIOQtY1tGoEvtYRtDfrp8Pn3ZPY8kJULoATnr6
LHNRhvhq0ddOKDpn3OUkrsC1Q/Nc+wJdPVV9lLgIv5XPMIBUNTcWidOWOWtU
bwSco2PKOzLMWb4Ig3P+Wfm2Ej76nYre70IiEV7wsCdUs+acyw6/AGgaXbt1
baeWOMysL365q5Sif1m82GVgN5hnXpgx1Ib4c73zGS1FG6UJ1LDqRr7vJAqz
gZBTtl7e3VwBvP8d/ifBEE9W5j8np0+F2Xzw6JlsSgsmEugnVhkw+PfRM+JT
nqzzG4lzGd0PY1DGTSa13AxDoyFOb65ISDVSqc5ds7ictJh9UJV1hZDTvcLT
8tbvJiXpRjkUDhWwi3uwO3CY8AvqK3sf6Xk1TG8AT3/MbPCP5oGY9lF2owAk
9RQpPEYDfKLeLRK3Yd1ZdohsVTYjC6vOOxtDv8WzplB+Vs8q1USC+Qd8nlkE
YlbMIn9gPbk7DEttmw0vnU5AM7LH+mOep28KVE3wFUFK6YXd4V7LGD0p/GdO
OjO5WZ7ILxKLYjUVcotf1xp54zRI7dgW/lR3jSp1PnfxMYTYkOaOSZWtJKW5
RXZgdp1g+HjCN4+HdlJG2cuKmQPp9c0bfUTr+AY9r57VbsyslVsoA6xk4qZq
LuRkdzPBboKbiwzaphAd57SqxaW2qya7lalH1BOCyNDf+raSvZy+NQbf+skJ
AEGpSDXTwY/O4fKY53ySoKm11F6VT5gyjtpyhLY11geVX73QkBaVit/XFvK0
f4TFj2LjsWLkDUNNTCJ/lENDbiEzElKz85tyjCHIVOHk1neXiC7iSZRiA3/7
mecvEAgS9P2MVYOZE80uaB8r0UlOuEmTl9JLuF1DuwW05aCfpYBqTeHfwizR
7PqXTIArvZ6KS4w/2tbfOFCCHGxBOv8fB0ceDhWk7zpCjk31PsPoqjwmpRq1
TPaoHsArKcuxM3zXv/Uo3iyap2vVF73DwOyN8TNcee4IRRBZGo0UhseI21ZF
aL4qtHc3gO+8wQq7qRsIYGVqIIXzCXFn9ZfqjPI7D8axQT+Kk3afa7ebPyHc
fAEsVM8XvHGHs/1fYuenu4OC3OlaaWZPf5EPbw8FY/N1otCLLLMdv3pe/14X
SLqVJUd2mDYpoRJMGvthpXNorkZpZ0+3Cs0uOvecsk1ZYUbCIxHIyNK7a+B0
9xiaFw7E/Awh07saM33PFGaDNdg8+ai1GWv3Rfh0JdB2gegeyreB50llzzvG
vI5BN8NIkjsTUixpHUW/5AjrqQePjHl1d0fU/ZeJDrr7/5yCyEUsCzZaRC7B
3b/fl99PrF+p5dxKjMcR4oGtJoNX0lhMnH6saSjjVQ8m5/k+JkxYqbCWUfSf
PcxsdoQSM0J87ylNxNzIK6Cu+d8yBJ+8DfbzLFge+pQ/inZTAXmNmR5vqgJO
XyxRFdZ9OZ8t8ocBeE9RGvZoELM7BUfd1JE3h0vdTtHJCpUy/vVJ36DcjboW
5rcTKwc6Rv+qK9hrf9dwKpjZwGlGjDOwUo8C2YunqJ/p/u+JmP7Np9gQKZPG
fgM+UhRbl97h59SLrIhA61xXYJflDBcBWT9lGWclZoqgtlgcOvPu+YnCMj1S
tKyD1R1CiCpyQmn1EpODAmeLACT3EsqyPJHodXSU2SetL/ADdTV3cfeB3YNn
45OtqR7Owp6aWhC2acMzrbcVxYKKTu8KaEfB58gqixamp+Zy4sZbCK29QalV
6dQCtiXaRvwvn2tVLCSgZGHKBjdWlQiqELGXzmqWisFqwGm+We+HxQpgv3ii
IAzPzpb40XJwRi0/x1SLzcjQaYS0SFAl7+QIgC2N0ardQNuVaBGTkSrxCYb9
N+guBa2eB0yiFUMcH1lWmDwcLytsdXBVjRY9Q8TsT3qFhRbwesD/u7HbOECF
kkiw4PWLbCFcjq+JcoTQjxaDAcyhvNg7Xl0o2XV8vCD42t4bqsISfPkbcrWt
TAA7KwwFLycPCsEuh5pqI0vyJXD5U2sJ844JjZkH1M/pqxdzOMfz5VKPGUG/
W0HuNTXlJkgB7m/gqj8PqXqDL6Fc/gpSlLYkH88e9Bg8gs1w+51yNfnAYiHg
zqpvIqM1MNx9Lmd/6LcKaJDxO78XmH7XzBdQKTJ6kevPl+MzpswYjIyCpOw0
PH5zJJpveHqBh2Bm8NIxgxq0lLRcYdUa1a8J+uu0mXfQtn2ckom1CTcHCm2W
7wA2C0W5uNoy87ng3SeoNUDuwVfzsSFOad5CxBKc50Y7hBlCGAB3V+p16H7M
9moQgllDWnF//OBLGrXgOIh088X1AcCXCzXXtRKGUYHp5uwdd/BcmfJ8zb6N
k8yLDLr7m6OSQohrdzbQclQg8ojSkRaXgoWjdnumMN6aJVamiVoH/ZYLLYv5
4ANEfc0+sIGbxarJn0PC5U5ImFBrvfwKXQoNKodWcEz2/xjIxSCfNhoM10fT
ugGVOvdR2Bc1Jz0ghFXQ95JybRrDj5Nf/0N5dMnAbV7JMdphg/9NmubsLvFi
4mJKznynPl4Ni+isJdGf6TK/JacmTgEdU7mKHjcBWxpB/TfUmXqLM5MclAF0
eEzCtxxFz452OT1HGvc6dBqTyoRuvVZB6t0e4SAZD1ST9+uBtzg5kfgAV4XM
e+zjPgja6yw6lPaUXOvpgjumKKHUsygnXXxei5YbJzWmTNzlRoyGb4QHb0Nf
j2a2V+hA37kvZ9/taD50eSkam9xr5qoyyoGjG9AQ8XR8NBrsyA26vB/uwLR2
8IJUItnZlxjw9UYKLaXWSfl1h6rf6GWv1ZXYPNQlXK1hx11/woID3XvurfT+
ex1qPZKbqeD+ONof7dolMbp5z1HDX7r/eGBXq6XFadVMzldZMpsrmobqlfF5
gA0q3LMC8WRaUwvdCup9X9E240cPstodVJaciYVEQ1ZUzXXCB4vkOEqEtf/a
yZrHHrfGDPL7htSB/NRbkSt960XkrQoJuUsFGZ9gnxiaxiXftaBYcikTZaY+
uGs9nqbctQ4MDxijhjFFClVXiiwsqrYiOhrORCFFbMVyR1UTp7GHOJoPUor0
GbAFoBmX9LU3KhfXNOgzCp4Ud8pvcstggklcPvougW0+feBZ4QoBIllAp53M
VWXZMTS5HMd6blNmRdx2sR9L9f07Ek0Id0RKLCpwFzYpsvuKHow/br0RVQsG
BMOUA3ALvDZJvjFnZHfJ57PmSc/Sut5mXqvenVQjqhnPPtvCes82fuu48AUP
lQkOxWGjrVZhZM6GVGa4DseTwVQZlYTvIz6bUBCzgfDesb7cvUHzeB1nBNe3
R8gTWlHy8ncrLNIalxD6TcCi+dbDsH0K3GynPWwzMOFG+fqT773iZ4DUcKLs
WrJJUtE7ZpfwNEymjpJ1GwJ0X8VnVRXbWoZtd/bzbIlnbT6RMeCj4+jM0g2G
QXfrtXI0Pnq/XRB22cAxGbfYz8iOf5Y5DFg/jfN0XtN3fQKzp1ke6ImcOLUE
4DXx7ZiIwaGvZIKpfGT7sE4YA8BgEJYAyVY+lWvHw0aspyFq76w2urkPQvBk
0Tnr7i/4EjvSW8Z21e1+YWkQc7QbK7a0Mus9nKeoLkIBx6btA8wY4Dkq4tzx
NU1923xoMYixAsU33xIyoM5jARPo5zeVqxNi5HusEFHGTYYjBOzFA23AUziN
mFPRlTAPRMbfAjDfDvwSyeUGdOAUH12mJjIUT+2r9yTMZjtBjiWI/62XSJQQ
4aeCSyuAH9d/1FtWYMzPTCdfIP8ONciFUt5VlAP0E8tH5GcephQblpP6IkRE
WHs5vXtoOSIlukzR3LKNQMKLr2rVp01bqxCpVcmkhHEUma7aOw/SUiY8Ur6O
YYR/TS3PFz99rYf7POYoHpCjZvSISGRnR2tEqPCkdH/ll7rZnZu4nBiUwAOr
ORAO2dnyJ9mfqDEyvsp3Okz00YvqEbBQDV+6T1B14vjORe53dawd6EWG/j2Z
Ni7bvHI7jL3ps0gIqu9yGONh2yeKJWBJv12bT9CrOWcRXbJTM/6MLao0NnIk
sj69FH3jywsZndjYKbh0FKVytplfQ/iNytflss7ncQgtIFvLKkl6P4daq2Ki
YayvZAg+JEx3A/vkh4/RLBO0UHZExUFhIwvX3KPXKb7vMeG7nmtuRGVV+64M
Svu24awcSKNfiSfS3XBgd8LDKaW3WUDW06XIO4SXCOeoJc80MGvXp40+2GOg
xMlwUj8dvgQnpTzbNSkr9x4ISwP6aSOdT+nM7WjxB9ILyAXT8Yohrjy8ZhlZ
GtMsjHsr96ddd+vWMgt6zTFbYEO5qmIx6ojvH0tl7/MPsa2Ua5betno1RpDq
zvGoy/w2A4a6hjkv3tiEoIfosi9xfAY+z/oewn6VDLJ3tfpTzv0tu1ZSa9G1
ElTcxSKeBzgjAdmo5+oOxA1CUEtWVeLyCNcWgh+EJ2Sf+S6NFVUaw49U/9j5
7wh4fpbc+zprhS0lfFKGXkbkYJinN9M0P8kqMjZlfgNyJ7cgznBqq0ALZqJc
Lq8oWSvePiY8+2QQjTsJ+7ZRRkLbwtOzAYdC34d9CA9tjxBm7jOaVSZXPGCX
ORmn3o8nXBEr4swPHFc2mw041/lkOAdLGVgg4WgBZWWtD1MQUedYRvY4xb2p
eperY6mVZnVuhYB21fUUmBy0vzMgvMsB+EeGAJLXO16I7meBRK1gj3mBxqBg
GjGFhKKOduH6am1xLRQKyzRV38YZKl+kUUsQgMwJYSvPWw4zk4H80FD/TxKJ
H/KVNVm8ZfLsxgygEwmF+OFgfgX+Xll9WLocOm5goweOhVXm4WVUSOovDDwR
O4fIByuOby8pUnp0mOl4Hq4tEfFfAhRzKipkYS8SMLUozTZZR1J8fXAI2IjS
TbD1BHZq8lb4UGs2yaqHokkqfUxghsQ62TGcVKIbgBvHaL225pwW1cPf9O5j
MEG9fFZz5Svbey5FZ+nZua46cqrJ15Vv9VDmbuSJ3dZHtOkZ59PjvT4iTOyN
4zoGcmWRQQZPgM8yEar5UpjrUni8S70DVkRXFKIPlnI2s/ewrUopEB0GVWIY
hvspt4TOBYD9tUIHKV/RXGXvOTHfWszFsh/m1b8v+4OIGP52OFbShD7D7oR7
ILRoGlXrhNrCw2DVievAJb6mCXIIz4UNLHw6r3K/tAK/RhMpMmga5HL5hCKi
JgWipU6tUEwEvANOUTwJ5VZG/oayQQELH/Z/w7IXZ2p9rssRgx1p03WQOLTd
WTVFEDJC1kycsYseXdv2Msk3WSnsEhb0wIaDcbsCjQ4CSG89NHxOG1nljzWA
Yw79QAJBEqk1krVAjJICTvIxRSRxFmYp08nv9P4MH/eoFFBfpzoM+BzHMHiR
TY9Ep5glCuZE3E16GPkQYy+0yefQQ/5W6cRTsWPY4ZhxmVTb4IGs9630Ncu+
LIAC+unt/b9fy8SSUKS9FemeLdcdasg+TLF6VmbHLMa4p9w9GK/9FEhkKpFD
3VtwQtGyLaL0lBBNnOhlaEaFtG3E3IEfldFevW0bmUVsYPsj/0815UPj4aE1
mnDHARkxqw1uv2Mu/gCESzVsyD1WcZSQp95nDTIeYf93hvvKfWhUIsu4hRX3
uEYXf1BomAATu+PMhNSE8EYoNrQYPFWzQt00eunzmmWAam7nTt8IpjenIZOC
uk2ExT1rtmSU22pSj3w2RpFEpeRkt/uX2KoUloK4c1J05sVuKiXrP9BgWjcg
KVfsPi900W7w/PYAM5J4CGbkGjf20AB+mKhyYBGb7cdAm0mlop425pA3iCFQ
rq16Te4AH3p+0+0pUpxhwmG726mQSbKADTyh+s961X7D58agwdTrgG1vRWcq
mzCHmFbNiT3PkAbLxxKCMGUdB6ksSuRJQxcmf/1SFzFuk0HcoMG+mn9OfltE
X21iJuNWMdrSvyUMeWwhpUVQopHRfy8Rf+T11wCJFDpWd8N79fBlu/zmyffE
VbJFH80sKKuoLOYZaUzKuCtPz+yY0MmUALFDGGw0tRyWbPiF1nnuE9HBUc/R
P8VAopsskr26rOOSeckh1wZ8jqMQCHNfLKe2Kt5kGDdHhbz7iQCnmG9pmqFc
VWD2JbxDSPFi1uipuIaoGIcX5Lg32U2zAzR900eZwwdnTKu+xT312V84W0bU
UWCnG5dcyLcjIYkh8R/sEZtOSutihGdlddMixx4CWfFq6A37byOLNlLndFRG
MsInWKmWDXntWzMBWT1dG7gzGCvaqhKs7/4uVNrhtKFpOjBwLBsyw1IiC8fH
MQeUrlX/s3eR6CrXMNYM3bJWZ9jqmrFer36ptYxKiMf4dPcHuoSHbkXx12Rg
KWX/x1dIND4mPdzVGSudYIndWmb+A04alcpikktrm8fEK+siy2Y0lNaBFWVE
gdGG4B9X7ZZF503Zo2H02BHJO2nm+IvmTTM2DhRtnw6eQ3m4M1JTQksHCmHD
MtcEAooVpAm5+bQro+wJH7ezPB87OI0PAfHtMM6KgUmPLv16Z8BzE3iWRM6H
9usCP7TUiL72fkGMN5lztz7ebHQY7YEXZYZK9IRurm5sckSUQ15xHSh9BUVT
/vv8IasvHNLFj+zJnVUlZlnG/YsZZWVh15AFyvglKoyPSySwitCW8CYgCEEQ
EAcNXeeSmfzUPws0imL5rNNXYz8zcgrLnSRZm4MlxAmhmSR51e8/9CaFFj2W
XHCQD9y9S9HcOfFb2bJ8dJO5qUOc6inBhJmGrRFaX3sPKFHfz5JEqUb/JCAi
DYSXlg78yfOsGdVqpyEoO1Xo5v+OuIRWE22O/997m9xALofQBSWA0/PNOfMX
YbYSwVARYLkS3U8wUK3f5dkCDoCIS/wjr3HCnAd/E3PdrcRnEq42aND2n9JA
9nYQiSLAYVHe2BPZqdOitKPdQScgaYHcr4renTUcJPMlsTsDSK0ROz9bCQTp
CwL7YdnqvT2HmXMTs0G/YIOtBNPx/INxtnJsj6304+BQq8yRNNc4xhsfkixL
b+jALCN/7xpaZ8N40++Gq4fxl5kl6lSk2UZ+4Ez0BB3iS6316Rledg9xaz5f
vqx28zMCqxdvGPo9AR3F9TtmPzSDYkBabdaBJUEMp4iZazQdm9uXxe1GLts2
5iFhbRSXuoB54ZSbLw6gkvTbBg1AzDY49h4FHDdTJO+MdcHPjbW4GjvQWLmX
osSBCh2YLOpzKd3Vy38LplLLN5KSNr6YqBMAk0LHPzpHdk2S50LKmvlsr/ci
6C5s3/u5zp+1aVjGxYR11tk2G5AkdfxYqTr8N2GdlGfgErDeRnJJi9S75Kwi
spIhfvN1pn0y/zbpZOLsqiVt5xyThG9P2VLooeaK0S0jUURYD7JQ562ku7t6
dVyXXW7GRhxor2XDRpLIKnf+X2SzOrgd+0jSh6RYVNxtuhwBBY9TEVCVqXys
Eqe/w1iN0+c4YKSRxnDQugcOtjDELXIx6Bz7bpiI7CEYgciex+vyAdSfZiz2
evFj9LDU35Y+QfyUgUouTP7XmXP5YcGF10vTDFHkl/1uN9BX7jil8m6H3Jk9
bWaiWKaWoqUOtVS6oRmAe6Aa9MXEbh0Bm1MXzmI9L3EgoCRQlYwGdQI6TUN1
q2MA2bxK45b3NaSE3lRbKH9nI7sE2Je0pmkZOQfPyuchmvxnN9V0wtOGyO/+
DqhLldrX6v6SDyiUTjwP1EuV/0f3lyyCKN6v9kWs03cNWXYZQ2Xf4Lh58BJk
g4BWhJvHs81FNqxMn/UaeaHsh+7Ng8Nv/M7ozv9MwdJ9UrCJqZ0b5rFZCz2Y
+zNN9VrflXRjGFkx/X8fOoX1TG/aBWaZGC3v9BPq3qRB42N4UkaUH2lv+646
up3Pqy8kL3yGWgypniVQdqqgTxvUO3pPtqcIAYsSLgy1WAeHux/cw9XOOvgi
IzMLuQv8NlD41wrG0YvCRKYjFYUx1iooP+Y+VmigHbfTH7Kr8pnusM/mHbSP
GdSLB5BSNCTSFvtblE7Wd2+cKorNe3RenbfccrwMIpOykn68LqqqIL/aSafS
P7hneTsc3yPj82CBqtMKtA0Y/AVIqjLEjfQ9JQp0NFW2ztSDy7Uy+Zjgyy7r
Hp8WU7ExjzQQ9QJSHpPmI8LqvQLbYovNY7ix/SS0ryQ4U0rTJHZycYbjaZNy
fjTELncCLt5ZyMTm6hFCRUpig6QRCPyLooA0sBbfcXPR4JUwJ8YyxZFbkVmu
O2Wpgk1VLT2e8Do1+LMQuHEZCBZwGIipUkpYIn3NTWsrdyUHjsiJcL2/w8yt
7LpdFfFo7JPh/p3VnCfhdzsFwvKHNQ+mAYaJ0Pxe0+FIryGY6E31Iifxio9g
kfuwoYtDZY+xuDXvcD3sO3NijWgLbfzzdmZXOLjKJnpgRaorQcVAYuJ8G1eR
n2DuO3NKULHmj315bLfQFioOyP96sy2DSKhJvr+Pb2AZxqyYEh83YBsQ+l62
hzHv+fOl9Ar5YOdQBranwLZ7EggxSLNY7+AK7PtpdFIIUj35uUTP/ftEr16Q
+pxD2L+FqoOL+R65q8Jxxrfj6jAbHmXrM17lb9ohNaH/gWWVA73+UMObM3z6
o5DwgJPPc4f9c6I/pdqmlTi08JMkyEMJdfaXQXY++c3zbEKZP5ZLFWCRI3FP
px+XU7G5IMJnenH8xv8kFmePguISoD1eBH6rPN2ZKwTIHFwykicqnc5sEdD0
AQeZ2lejSCkx2KLqE7DpkIjqy/bomnd5H63LYACK+cI5BUWmQxyYfRLYcFw/
0krGP97VHRXKDiXz+7VMv+EafwqCuJ80LoAnbNB1ogusDgrOicvEYlxm1sOD
llfC+ubs4Us6KEKB9vmG8xecU1VZgfbFJw2UvgJybZHhwPN+/qD2S9B949Ew
a22qPpdqRNETuvWJooe5tCrsvux2sDIr6yoMvVjONHPKuwQqHh1L26G0m8SG
SmtL3DG14DdlKqQHv5MA26vvvG5NKXQz0o6Yu8EunXLEdnw88NeqvUM/2LaQ
t/MH5wVCpg9rwXSTwv8OJDUnKUpUDmwlI/ozuOZJ6bd+cY9cqgHwu0GI6IMx
gqDiksP9K44Joyt7dc83A0h4toH/BmGejMpCS2kcxn4BXg7Z84dse5clZJRl
titTg/Q59Fg+kEhiSYvAKp4gxgEU5fWJKdYaMQIQIO7LQRvW9n1kaWfWHNiH
yV+UWPw/Vus2FupCyT/Q1iPr+KjGf17DvQ7kkyTk3NqGZiIwoRELrWXoZ0Ka
RZC87VkvJvwMGweXbzqwfyoplkOsj/R0Sb4UZFW7GDsNYzSvg+uGUGM5Gtq+
8HgomsF1xpEP6sXthDxglPgXCEr3BnnxwSxuo3Uc8h5GGaRDNryfgtCv/Ma6
w537ORDCwxRW2/fgN6lwejMYdZCPA0etrexlJeN90gYaqF1UGyVh9pqjYrgA
cKCU3RwCiWglWwC9T2e7cgvTmwxhC34nN6kwIktyCdHUSgigrv/gc6vRkEVU
F19QDpw3gGOnQN/iuZtScTF3YNdqDhMshYJWfuKj6mfx5GLTYZlcRhmobnIg
s7iSidf9/I66349ghyMjEBPr5HuhW7jUn6Gb/pkS64eTIJZ693ZxkN+/Nags
u4mogj8tjjQBbXsJTUc29p9RJPIGAqAE56eX/x3iq7CzFpz+4q7/LzSOIC8L
JCHDXqOGlJJZbWvL8vBvTGsO7NeAHIx1J3D02G5vNwzvhBDp7E6IAaugzxsA
lJPqZKEeSf2tv5SK9OgJ0JekY20unsJDgDZ1U/XCOBN71+XQ31Ft27fJ60Xo
e+Vu9WDYwiqhZnkOEeSoKgJxXfWIr13WCkuocTjgzv02UnSveOII6OsvRo1U
BuN1zxanvu5koRbcRtsPR3lSzIByO3uqMEv8tTRlsFziZ3uVH/QBGnOIkLHE
pYKAta+dlKITg/ehKRsfFgvEkndrecQjTwhzicP+CksKg/xYpp1qoYgPzfhb
r+kqXAzF72z2tDBjOjG3V7smhvbmF5wFWPFkwjZSpGARqU8SeC/zZEyuNLp5
8rnoQDcr9RTcthKnTcc/UDaqSKDkovolkcwIsfTsvym69H7dTyPEhj6lt9bZ
RxO1kbs0VidJhObdP25riDv+hWkX+JeD+wq4NFPkS93yw23N8DlQ7Jt3V4AH
8HxKGvSEFwuVe/FQ7/lDKntVMCd5+GcuoSIfumn5wIcEDwQDFmQmxJKdYuDl
Mn2VTY85IMnL6bRQaHiP0HQbRSSoj4AXO6BhfnIjmIyAHQQQ1lKwJ3WtYC31
6bn/+dLPjVzp0ysLsJ9UsO8BhHqGq9JNZPyk0/xKgQKxan+YCYipysjGDWAx
97ZEDUwimKZGn4jCvHMtM5JA/MhcfscRiZgBf1Duue5PuBnJ5t0jfI25TVRQ
9o6WP8s5XAiAwm3+FtVozWynPCqhG+NFKzepB47wsD98LtCotpcNdoQGznnN
6/yNp2dtxZ70D/7seIZSF/7miW739Km5cAFIepmhcC72l3h4+SARveBINa2U
1K5fqkXZlxnCZ3mTmzW50o+iPpgE5gsFq+k9q7z3tt/MmtZrhEbJFm3FaULU
JpzxORN2JjkpnD8GUgMfpYskbFwol7oPeCb5iwJWgp/cAAsGEgVCXYoFAuTa
lpMEHB7BshKDPd2XMB90O0GLIOmDJOTWe5NlCpInRbh0ByxYH0njU8wBtaC2
TTv1VIDT/ueSJtjiPQBcMPfF7HaqliALPsJw0ykrff8GB4PjJp2RjXjNZ59O
N92YWFH09HgifElG7w0UzR1KDG0An4+9npksA6bekxfQHt7Wt4QNFeWi6FFm
aYuwvNtl9VbLK2vPKot5dn9VTZZIhmChpTv/i+jJqr4JaqPNzROcQeATPvzn
+4UrxLjIKXhkZJsuxy+PMrsOsaLdQZBFBclneOXF1JnesDCw9VzZU8gxiZV/
fnv6kcpSerZBmB3aq4YzSj2nwCoJNrQch2yd9eRCeb/6kma9W9y6v1f9CVV2
+lZDOeWhf4Ff1duUt6ohrudzViJq+ok/+l5I75ARxgLKAWmOhxJ3rPWD4VaW
5wb+Qf9qmqSvW02PnJPcvl/9EC2VYKlAMhwl/87QNCe5bnC4ngKJtkuI5Xtp
Jr6E9mMQqWgHWQMTJR1xpkj9mq6AnlnBIXcSKPdvrmYMJWvsCcuf1Su8QIFk
xgYb4qSOWqJ7+hewoWcgbjydcS2MJ3iKizLktO+7s39AxTqWRCv8a7G/+hRq
0oA0AhyaRdO/L0sBtrnmbd/MaBdyecwp06lgbGxJoNkALEZdEPgGF1oyND/n
FVYiK4akRR3F87PU443zUmhB5W7teilP5cKqMqo0hycS0hiy+Hk9LG9FiI/O
RVr5vRs/0cmyTdr8/6upRgy511Bc3D0Vo8/GXULxwJoTwMlUQEXtX5Rvkvyf
nQiIkdfJ8DpHL8emqsUD10RoPx2hazH/J7htjdEweZ9nh9hjoye73RzRZInJ
hduRrhRdPG2kq5u2lkbNHiz504MzkH892xBe4gkjIxoAcmJ+4w4dgWYMI4na
lon8M1xLifb3w8/4Lglgn37av/12AQZ5i4SOUH6cRVdLlOXA/J7MccpSBvvL
fS4LA9TVkTXERexmpey8nAgk6wpGXPSn/bQSGg+fxyzO8TqJyYBCrDnFssG8
E6RiQervVorXlsfZt/fDdfttiv5rH8Wmew3NMfO4VMAfAyyQvASR0yeB0vHm
T7elDMLyvfkBjmcbs0oE0snUMo3fuJ2cGHjmxZmj/COoDfSi1KgWaVGx5a/u
/MMNHGxyT/Sh3gbqiftajUWAgW/z4vrgrTap/XXyD/7yQLjLZgN7Eno36wdQ
YZqTkWEhYyi+YGcGvSeckVUmptfybm5x37G0lHZ/F+GgTDNfkxv188gWZxoV
KONqn96an8SQjhvlPS+rhA6LGiNf3B0CUnJwq/G/23vZe23YsD6hnxbKZHig
Oh3G3f/CTBkSIYWxJ0w+jz1xVPjBtAuKOq+RWVyy1QZmcYPERa4uGBC2lafj
NrXsDSksJ23SkjwZUT2fGrUaf/vD3hENlqgXnltE9EP0VR3SX1OyCBy+aI1+
90as/Kzn0Zzf+1bve7KuevHA75xPyrObwHGi9zsbwDb1zQG7Y2dESg0+rxub
kVNZ0UxBvRT0pmlhviVwLegcO8MU0+b/7ep/lUhe7S2KehevN/seKEc7kY6e
QUBUu9DFoHYFywG1fn7KnF7P4sEc7NkVDr91oFbNA54mKZ6iUDVBbatAbSf0
RMoiEyeotbyFWs6rr+wt2UMc+qWBu4mcTbyNl9+FMqaZVd3flsD6aibwW1Tu
WrGMH60/5tKL/Vf7vt392O962fjUwwikD3ByzwSD2/VShZGZuVyId+/7RRgt
5h5+JzJRfnc9P7SNxtlxhjC+kvikhmBfi2LmS4z59rXC6z5Y9I25DYWguhdY
HQW7+dxGewgWQEKaOiQ8TfcXNOwsGVvtBeVY01iLtV1JGWCeYdCRs14WpF8P
CIIdfUJIcAmLBva2MOMPAa2q+/QCFDlsAKoCON2k3dUr6RxiXPMDeuVaqaKy
vC0tIkiGA8Mx+EgqkgNHwT+urp1NhVlR7cLpZ8foLq2cQQov9gY/SSW1NfFl
E4o39GHtWgNT8x2+JOI7Dt2RqGrF1pP2AhGyb/DASbI0pieiaGKAHNZWifCB
umesQSqqxye1jS9UbpfFnQHOie6v6bcJWoWzYB3QYBbtfs/HTbkkiA/A6l7l
dzljpMNVxlBbnhsoah8Osu8OYzMbUPGfEo3lvd8w3JGzcIod/T7fWHsN9y16
KibuI/0B9UY8f8NVlgbKGup9fYWK/y1W6+itBj64zejqxaYSf3Pmb4D3Sfad
h+3rABPdakxJeq31dgP4aEHE3nmPvFR/BBTZXm6dZi6oiYhLvHM0m8hFnQAL
c3fME873GK/8M4WiwN0JubbMUL86yXL4WF0ueiBYAPIuHBTmMC8m30lqpyTr
owpVcOIJNOtRXl5y2rZGgMQTkizzJCt6Mn25q0c5UQfG4s1JVUxyFcsHwwE9
cPI2YHKSJyC41VhmzPqw6xihZ+DQbJXeGrJX/TbsuGOOaxC99BZBhfPFfMGt
W+PuOw1lijwTxnTPJoJA/mml0zNqf1rQvH6R4kGOWqh/YeVm5P84A5ODdNdN
E0UkYPFdR/AQ74tUEh3vBIeGfnk964Q549ESg+5GdyD3H4uE0u6MYYsfEpRC
FhCv78tCTqRnPB8NeeM0aqHS7lb4gCS+f7zeLH4Yrbyuerix6GfN25j879yx
oOWoB83i8rCMaIDehkKyTt4vwxZejX4kHeoGdatIXKqXxeyeACYOGYCBfuEm
uW/EIEY4FKUEfj9dz2lZ6C8DJvN/LVdvP9jm3GLV9BZ41wgn3RWiRR385zgg
sddM3jIayQJHq/f5SJXt96u6PSGLPOR6sm50JnMhOGGyIKczAkB002D2R9np
Zs1FvT+DuF0uwLZSKvHwya/6jtrAKwkGoPkEEltqTYmYh2QPAw7f6YcUOjXb
fKw7mXnESOBkojPKeL2+b1gAQ2hYxJDs7AtqO3ob+ZwVC0ICilXptuPRKe2S
UGcENCZqhs83roeKWk50cBoVG6v0tRXy8eD06bVZXClLlA9RvshgTYn0Jzl7
ncalCvLQI9K5VkaL2+1OLpTwZqmFv/wgZUddbO6YFjNfixiCKvUNSgOqftDj
UITf+I4ygyvgOrR5I8aaJRNl7Vo/FlfuKImi3FrCFf39U7qfIWhKercWNaUb
r6fj62RJdEuG81365JqoD8jjMYwWdxZLScPdARMiG1fAlsOYUbPHyOIiNg+u
80o7naWy+jIg7ZDLhYr00ELgP03uGoA8CZk5mznI3J0wMwdmacw/ii88KkAv
ctavsGsj/ZVZ4O1wtEu/NgkL949xzz3J8whVgoJYfHpVrh5F23QyfXOyfJ6B
5iNjcWg6pVSHcCUz0pV0CVthtELH0hOymnA/BSTPpuI6mDsosAmKbUvzrbMe
3B2jXjYEdjZe2GmXCpzXf8FWRK8pYToiTlcPiWKFh8aSFdvl588AqMya8iT4
7e6shcC9fNDWzDKuk1ISKuSJ4oHzekYxYs06857rpkkpMiTrHGTpvW6LLCwi
B8D1zdasZ4LejoBwMxe4BlxBfqF4yIUWfMwkviNJzy7XuUT9x43i5Ak/nKso
F0w1CjCDblhM5lBxTP6IVSAOJr0yqXl66EzMe8j5EyURi65zb0C7Sjly488Y
sQoc6XODUs4tJR2emZsVRkOgekXXD4sSwFpY5cEw+3RAz8QNWQkuocVnqPTE
IwbtCSFj9Q9D9oITANcZDxOeLWd+Ys2OmhR6PlPnUAEm8lTHBeMJ9vsfU+Nj
HXr+VsGfqwFPExJKlhAVuh7HmIyavI3HVM/Z/dGnyOROlxs/UYFPiBpSlJhV
jq+MnbWnh10Ahpe9VVWmZ2RagNBj9ufKfOwmPj64mDW2orSc7OaRnTsWKL44
M1HfLZdk0kWzjWI4aAiOB+3OX1FVErth9f5wMLn+sRiCiFqtUYCYPTA5gBrX
+8RKIa59KwDFR1b6JeHI/Hd5vPaODnYa0CHhoAHxshTLIs21/1SLJGSQe5yO
BeTr3LhEhlWgq/daGI1PtcMiivwELET8Zd9QWygblrb9ujprB1GL/UKD8XnE
kJP+O36LGV00L8V9ra32gFa6ZGgm5Zk3LfMGRz0Q4+KIBp0/KgOrc5SqNr/3
fm3C0IWTw+nwc00zIKtjdB1kKdmiO9ZV1y46NCPZ09q3Cj+mh5zIU8eQQY7a
F7goz1geUYrbpe+7PKpfiHO9uyvchpxeyFYlBacZXX2U6/WOlz95OrohFV0G
4+zTkrIphlaMZwU65KBzelVDb5B4w/yI+DiVOf9t2YrARe/BB1Ahj14VWipb
lqua706RamdmsZIPvpepMVhPlPNV3c9u+i/s+eXT1y5rD+l90MdWD4lMyx4r
bMFLE8G5V/QVUHcBHM9MhqodOxBbqlE0bBRE8f5JGF2knDzhTwo6+g81IY38
JQ9KmZ1/AlMHDjklt1YwzJmCK5+rh89NqQhgbAuJopz/NnGZxkKut8v2Ij5B
/VGBVYmoW+pT+z5ZGDWXAT4Ia/spKYyDNbTRdctg73sXO9A5Bk4ExOBuP0ZF
g+WyqxeiNC0bWd+Q2fJhWqORG4rtCuTqVZTGPyrDDEXiY5P++M1GH2GyyTLU
vRDWZZeKsy/m0OQ3e+gw3jH78o/jWCt7Y8ueSWh6U1NPZpdzMJM3YalsLuRS
V3rW23ssP5im7whkPmM44ZkBkhDrwh6J7SBIiUiHhBIR/D+cDarc6Fo0ssia
Ty/WSfaMFwYCh6Fb7k5JHCruCAfWusPiQLqWUWpdLzzaBxtJJ3stRyPXThkf
GXCHw1JeMiJkiUbW/cc7FuqTthXIgC+1aHKlOSF+NpUwydw4hwwdczItusFn
haYBDHcmM/GIl2QIashI1au5bkiiL8oxI6yl7UI2O3ca2/mJPg4iIoheWgAH
pBUTMfM9TbhDTFrUJjMOm7EfOqDD8yAYm6m0fyDOH3NGRE3KKZ1cjTrQrpCW
L8XdeOlNRCcrzQkZlsezhFr1d9zfNhcjpVB1Q/4A40+rLuPXoEN3tLyLOF9+
/w1OMz8Ltn/Hs4AHV+I5058RNduInZfg8MvFPJoCr/m6iCGet0BNBfFJLFaz
YDYkOnc22C0cyOpJRd01pVRf2MPZPc51WBaqVwkVhnp3kQI885yJM7W14lk7
J1Nikyc35zo9DtDF0T0DcR+0z+eWOM6mb8XhG1+kn3v+n0F/+LCJq9lOBIYc
NHCLkc6SGAdgU2I9P1EI3NO3APSJCRBimNEvHUzK+7qI65AbbNZLVKE/NdXN
ilUrPxbH8BX2s0iCiXknFz4x1aA1Y7b9etQQIXUxYTlxEalnI69T6n5h/LQw
QgVXlfAkvddJkBvBaymiaKIt8jnvea56cqOhuwJGYovUMTB5Xd2ChUbZuZna
VSQWYW4S59OZ88fIBeTCYKGcZrg2E4/H81eyXNU/ic8n4bWLNW/c5o7DFcrh
5eQPncSr2DbP0KBSz1MTfVVn2ROY5iq+uk/ceU4su4BhAOzewfFZSXiNOewn
kdPVlemLwBX4D0xu+ZmyXherrSf1k5vQGRNJr9M2Hca0VeKT49O8pixVibHb
LAuumK85GhvY/4e22ly68Y23TqR8gUEraM+TAaVmVsuqrCyIGPo09LrKvkUx
YNea5oJulPEUdaukJtas1CTHyvVp+LhcIjd9UBt+mSd1WbWHWsZGKQQGFwPg
nuBxu8FX6iKiCYeeeVIYgo58qjOaGsxqSyNEH7+meUYsvENQHUA/XrJWbtJJ
k6mEGFNTTyoWImeIsZI03qt5321K8n5PEI+kfI9AxtwMVMsV21W1AdyWGC4W
PFimP+zKVtMT8pL+7pX88ywLS3yBrtSrMzoaOtW+B0EDPcLPlrzNaAZUCbam
NeEtpp/WlF3jsXrfxEQNtrSlIyCi8nMLrMCWkKXTCthVyMs0azOzP2d0Vo5W
hoBXK/dPcwzBXUtGThbrYFfB6FBRMCA/xCVUHhuhbxcIoVkORcr6qSeD9m9+
c4V48S0SFdOTBp3yToF3xXbyozJwZ27Eq2IZZBUFRHPrRgEHAJvnd8f//u4c
BGyyUxy2DiEpG7skrAnqGeBMfnGvWD5exE0mKmWy4DS/wSY1yYQaKqdTIsOk
T0OogayfENZmdGH4MeNjws+H5B9Z8CMpNnIRUjT63vyGTiskaIHuydEVSixB
jU1cesNOiC0wEO+FnGTACUWuZKaFClUYOAYegAgzYMhVndZWa1GLt0u/RYaq
IaOAErXbRCqebRbzZbcgSHh808WSAXRMRfi4L2zmqj1sb+5Cjf9ow5xYawF6
mcR7XqnHFe87bimWK69D+HYDKIibUzRxEGOsGJe3zM8MKX1AjyffuZ3ADluV
g+YZXZIcYyxCJVQ1ztOQ7c3Tvmcp0yazFaZ2mM1i2jXEjyln690LugD3h2fv
jNvK3/KO/eM+1BWY1/rNYKHyHVzo4zwiJ+Odp/Uzaq/lwa6/371OFChJ6ivY
DfEaOO1ar/h65pRVWU8Co0NabdxkjN48CUUG+5nvV8z1q6TMfgpD0VIx+6UR
NDfmB0WLrkAUSl9Z+tIxPAIEZKZHY0BZAxo7Apx7Z571q9Dy2Hfc0hBRYsUR
VIJAl3mou8GP8wU/Yp833WB9u3FeDm4RsvXLiU2Rda2xgVLRt+jK0dcMR4v2
/E5cz4PEFjEZksL5tZYytVxLAZdkiJEpvRJlwlIwSVvEB3A0xbECN4uzWo8g
EtGO+IBhq4DdQSSwFzZKRXe7zDjQSq+WBJ+4cjMi9o8y9YJSiMoKIhfFYjNC
fwB02lzpoKYgeP/yiGLpqdH73aW/wuS1ZcfPJFccxY33U2vK+wcBTPEHr6xZ
1ZFe7R5UyCPGXpI6rW+iOK/M9suxY43StyQ8IE2y9Du85DTyZKjbtcX4NIUo
G3ZEUbQGTlQ8Q6iBzrHd5Hl2cpbS3KpPoo+GP4eLuxEJikmjcVTw6UuTnCs0
GpLX0cwD1qsuOq1mtzU7Kz/DMJWw5ZWfJr5lnBbeRiYGgr4H9nLQqgBP711j
34niQa2OAy0fnzbY1FYrmcJonblvMMJ2/10oWYgnyQoWxW7SWDh22Ne9seA3
agDDMhvbrTWDiItFnKGWL6tAkNs8N+rLgWmHuyGiZxqwcvW93Imml2swJByq
KF7hHAOz2LgJM5Owsm8xzFVA4pEawoMcXXNwIugzYAmWpwc2E09QcNf31aBT
siLcIg9mhgClw/tvmVhmNTKeYW9EkqzUsTTXcRIQNVWiL3plf2yUP9Ybqqbt
c++kAz6QLz47Kck1jVo/UBJADE65zHXRTdTjLQyGCCfLOCZ494PoxmwQV3EH
4i8c0u1gAvpwCOlBDnRjtoaeV9qhtqqybId0nTvW9bj8JujsyEUGj8I8HXqn
eCYwTwubouhTVi7ShULS1GM1/3W+9Nsfn/sSB9+HSxtN5zL9iyJh+v5jEFrF
+i/ZHJgUr4U5IoImf4Nnq7gJBhSm0kJeWrH+Wu/TrIep8HIg2imKoMkU9Msq
+XSOBoUmCm5V1BmTYpu5BUO2EENHcrpiN8sNUlg9wEFdsbrgX+SiOJ0AxmBE
Lkt8GDITF86Lrx1XbtxePKIJLlXKcVvWh3oPFo6r98u34Glm1HjHbIAlMRV0
Dnl5pCXySaTpFKEhziTH3/H4IzU8HjAkWVur3ZUBanUls/gI9s9cTXVnBrUa
lim7tP8buGshQdX1RbaxqLfuOnhY2DH7y9FkgzGfZI5+0tBiGS2eoRivmifZ
gYn6MNjzDTQiwnZV4qmTf0JG6wxCtTfiFLu4QdzD5kQWRTSxXpuOmO2x+uSy
AUvQGjbVePpMl6oKX4lqMxlYW5TKxUvWWDqi/WuwKfXIYbQdtgDHAVxJ8aKH
gt7F31uBth+M16SsPkJTWORrsGM26DvZY2cW8kyoophHCtOgBaa50UVdYiE5
vfDHq4bt4AqB8A0E8Y/P8jrv12vBc4NEyCMmFtl/mGPHhubh1BazXnFhEhdo
uNwr5uFzWyGNlyvpE/fScjhg9RIwbumXB9W4d5VCt9RJ3CrXwsyOxZd6Kb3e
wGyPyCiJgBcAMi9JSmmSVGHkTGLare1Er+O+/LnotluW6uumfdheoHUwOFmp
oTHec+ZIsRbHTeyqCqtzI/kvsXe8kerb+SgwtXkyz9gKYnwwRIyQng+c61U9
TSDQ6c97bKPSO5viUVMQRfP7BChQnTeHYEzvpCOjQZ9ZxVkFb408UgO10rJJ
Z/clKBxXkueEFEojOZrQVDMIWjYIK8xl3OXOn87tHRtEXRTt69sqJRj6U3RP
MUzic0dK+ate30ROmLk8mLG8znp9/V+b1i/0ErIQZ5Tl95YH7Do1azTAXm0e
9s01wnacJV6QWNsfRmdmLC7+Um4aqG6Bdl2EmVIdWux7Ko1sOzCbTesMtj+p
okC0AmS3prka9MNRZ9ZKRVRBefeMbFE0f0l9i2/+OMSc8hkf0QqWfUaKrXk4
9cBZeBhL+kEA09uEwepdt1BYtD/JN4iH4FkfubY8Ms4mo0qCElCvYg9qjavg
cL0ScrbXfkWNLbjSXSm5LpEJRNcwDkFMolnvsrCZoe97IKBncZBYIDF9yMiA
wVZDAc43p+JtmlGtre43v+hd2kWHLMQJXyHtqJvqLm5bfMh466PD5aI5hWxH
j/w8aXnVNcVt4xkHuKU9assILZyTCt0bGRPmiYq5M0ci9QmjtKDEWqdH29Ph
h/BJXBLbEXhix5EZzWQzvlteHwvtf5ZvtTEcWLo6xY+Fuv1j+6rdbOhPPxul
MvQDLx5jVu2+1XUW4k8HN8UPTgclBWMiaP1zutD3EpaVnYY/DrDE5CAo4Jm7
BDBYEl5WND/PmDvBFLLgo69UUTrZwhc72d7sYiD5f8EC8mlcVHxvlHpF9tnE
2SW31GCU50/JemR4ctG4SzqpUGtmtI4siwJaCuBP2h5qJPNaj4euJMxNcxeJ
HunZKCAI2HU22VXBURlJD3FhfXoyAaZeNmM7ZXrO4zgABjYMZB9tjaqGMiwz
rGuU/+/jnpaNqTXGhbLFUPoT4q7xlck36JbSEnHIdvXq2qXPzUcPjvbgGnY7
UAuudbC+m6XFvPGBaJDrryQFbcddQTmnarW04BQHKqra9WYdslvvuyXjRAya
8rh7003VQvWCkg4rbFy6jBhqEaEhf3xB9g6n2BIaxbDPyLwg/xRe/U4EZXdw
AHT/JAQIEUxftbVqHu4vrilpqrVe6woe3WdIm4u9d/vbOLZgUekxdPALxLau
0lm+6VJRhcgsRkqcQ7ZgojZf2IaTRfwZvIkj1zUF5WeSqoQHsMnAhEOF+jGn
+IYhoxcvphZmHCk7vQfyS8ivRlaDgLeb6XOuT/ge33dFba7v3tGGuNtnPmHt
YG92NDRIaQzOkMM7IlEDejaCvOES9/vKIkWH/rLc7O3eMgl8UCKj9STMAKFu
i5WBO62oqTl0kx1z6iZAKVAFiGphRWywXUzwEbmPxJzJPMQDv4CT376MiM/d
VjAF5obc295S76mUph4hbDOmTxj1Kg76FeLz/F51Z1nCOinI46R0w/I3CegN
5akFYyRrtjWQFlDpvdeIRM1EhBXt+Gtin+yaQOlW3B4otrJvcNjn2j8on+d8
e8d8lFqjJRuNsjktdRN2nCr7cxBFeuz2srBSnKwfD4VV5ykq9v9+IurtSy82
RM/qWBt5tI8fctvNkcpF4i02dWPGDJKw3/eoRyrevW4sDn/4hDeZcAshyjas
wdRDlDnBJhgiLIZ2eNE1muacBqbZ1A/yJGHjIiNcG4KM/CIsn7c1FZKRdVlt
QSQLXXjOYKpA1rayQ9e8shPLfNHUsfpESiKWoJX4QySLIuS+GxEDfZRooEdK
QcTy0Rspe582JRmgPDNogM2SUifxJC195oaKBm3UIK7redMo0WI2o8rx6Iyj
DyT7FkxI0XRwo9+DE6qTyqcpMSPJsKW/LEHSMx5U24CpyTubY/v+Jp2bWFnC
m1CVh+cOw8hBg3R8vPrxW2K2+V6ezKwsO5REhPVfhIOD8P0LYgN4eZ6Leeyz
4xDnszmcJnimCB8iapoq3qOXFdcOTKQ9Enx1Uxmdwlb8B5T2YPSJNISGdIWm
tu4ZeUIv17BwFlGjNB83igaNHjRpGxYS9wb1mX6w/SXZiscUA8ovVUVjAH0N
3ZFmu5nW/WMJeZBIzuFBINgqQKK79AfO9xiycvgP/leOqjLSqbd+3n0jfeal
OiD+ueVY0colDBN0jkMTWgXYX1G2+zOSD019tUJ9n/vjjBSUdtedIw51fCHg
7PJRjjizqzGHBB/lYEAHpUnsghEyU8yoWxeElRmMrrM5Rnazdw7U6Odz3Ree
eZcsdCxW8muYYqirDpC34+nvtFu7gFH8np3ZnASKHkMPJTl9H5PMICPspb8z
e0EDmvMFHbX/X2OvYX5WX2Zan2ZKAQFOXe6/UWhANgmhjW4BdAWHL0CbJPP7
PJuQMrq+WSu3M8nePI3z7Mvay/GZ30TLNETmiUyGD0lwJJeFERS8MJBLYsqs
lsFtoCnnKNo68bFQSBwIDzr071GlzsJRQsvWDnLQPuPJlJw1dyg7XGaBNxNP
PYi48RT1qC9XlcJ8bnO/RAmiHpgKfPuSque8SQUFttvUIRgJh87a73J3Et0P
CTwBYsppzb/5+ZhOyyb01YjZjT/jEagPSTjHB22mL95jiQZ1WQIVRqZyg6em
pOzaqSbDyn4m+uA9vgcWSWP7Ik1QvlxrAz04jHpfwF0lbtag3iZqqgouynLo
wfIbbQTtbVMbAifAV/NgbwJK98bbseiLH0UsdDncsD03yWzl1JjBC9G9NitE
ODRo54JW8kyJHrJfW+EjmByIN5pwSZmQfPs7A0MNRSL7B4HoJsjcAdSmQSzm
2QHEzsIismtuPf9+s9aWtN03Oj4URqVTRflK8qtR0cKRbZrnnHrcop0ALzjG
t8R/VFGaye6NCUeb8Z5njOAhsw+rcwleoFOoVlwLNyd/wcZD79pcDt64CQy8
daqZvaPsNT/b1znXI2DUaatFaOmn3sGYobaFX3HpKTka9lmeYszcdhdB2sBu
Wsc/tIFVJpK14Drdjzg6gY+Zxfsa+XhvUYCKwwFmy2sNOGEYd96dcYr8ol0O
wBcXTOO6lzNJEG64LDCWdNdTsLCBCYNIStzemrNsMa84l3fqFlgOCWyI9c5g
bEfwA2LEbSoaOt+teYYAk4nSndEgEaiONXk6ke7KAUuG54KqJZsd3/qxytnm
KJ1P5kXgqHjC8lfGlEbVZpzBFHMnRvxM9CJjOzceFkScqtp8mmAk11Yr9OrZ
yC0p49Mwbrb6lwbz/CxAwUAnZBNnLADO+ODk9cCZpl5uoJSCCkezvrmqDjHX
VtdzBJKN8CuQRAMutJdLzOaCkG85smBv0cIPlTSlKf3yulsl7lNUk9rAALCL
i1ySACVUwFfVSf0dOY+ouiN1hz5AGRoAjgjFdHAMZO1iD0K2E/GUybKGnudH
zAjBbazEOJcDE1drsBcpFgaRAr4rbqnL7VxELy7+WAyTKU51ZiRGQzj6x3Vw
U4SLVBH2Zq3wocTiSuyHpeZI41PzQ0ofXGdn72q60CUn30+LfbQH67JnwdZJ
zDxuSVeWgF+jdqGYdt90bsFmCAgSLOgVZs06hrm0m4OHoOjbT4qL+GOGh1q2
chtoLs/CHHiDsfVaQWrKCQd7DO8EbIsuuAkPoeahYD6HjyldiXhXkHTYV6Ef
p/tZgnO3EKMbpstPf4NCmeo+m8Fx0PKsRbBD7Ii1SMmuJJu2CsWYQ3VuSDp/
ru71dWCe+BxyAUuFNJ797oDBYkebnoObiJBS8cPKxjMJflIFrAbWOTxbOOdm
AjAIVlLJ2QVKuYIw+jRnNgThGNz2JYyeBggixKPh5Qa2+1Qt9yg8h/V758Fj
Ud+FiSQpeXGc4mB4DN4zPFVPJ98i/g4RFKCDOK1KUGs6Al3nF3Uio9bP/1Be
oU5tdZCsx9kg7CGvN6e8ifbirfbbUMoizxfZqgVDRleYnnRLtyARvDDcddH5
JxDtIAGOacnQvocRygKO6OG/dmP6HPSBcLjbnb5zFHeWsmGC2k8xmu62/hGb
1STaSDuBeEruHrYXYAuQk2yuUWvDj5G2mYctAMh/JZCYOLdH6ZCE+gdoYZqF
nF/YG/qoVZdCl24kODBjtj2sIhv7mTZ1Cbk+EWCJ/P5DcUNlaVb6B6Gfhpse
vVqOVwBVFj2kFGoYxN1GgUibpvMTAGghjbz0MFwTS5bo9skFcD16DdOLV8hO
NJ8FGYN9/X5hUWUZKdIzq34rrbo2TgnAkseLIeAGQfY8SA0/0ZJPhzLsSZ8W
BkSa0pjgR/1rAhjFkF35ZB9yoIMABVMri/RbifiBT2cnlNIlo3m3Umd0vnZ2
rd94ccFPWuqD1x4+Mjf37JA2+FiDdl/DAbGGJHQNgI9pV/WdjEOHMXbpLfUA
7xOo2Svf1WPD7JlUUqmcmUNrLvJiB9AlavW4+PC7TLubBXHc0UvCZ0pZR89M
omhhficmFBAIVRjV8DmC5wBu8oaVT9cFWDWzQJd9y2VnvoThP+e6xqRIYUuM
99J+qR5wpp/QwJaHHauTLZRK2mpqvFe/BIfnYu55gwLWr1konhee4xhE19wU
I1HBxXP6ZmCVUT8MTKa+miFrkgGFgFpMMuMWAdQPIgE7yRdpdcK2KSj8pqDk
gXFAk4MAa4C7BVYUzPtzggste5+BnPArqdEmDK62ONKBRuR4hUeJ5w2GFFMa
rgtwBAKtH6/8cm2S0GTcPABXELcPBognhmDQ/7OfedjQiO0eTW2Y9cckxiJW
bNIF/A07Q8PG9W1RSNE2MyGKA63/9G4hRBngYIRo+jc9C6NK72ua+zn2BUra
umjNZBXdLsqrSEEH6jP/vaS7N2kKtEN50TjTuasmSa0dpyie+SGYjN21x0Gd
VGYDMfJIpI7GLQL0TaRJoEOJ+G0f4kPd0uimXVx3DIF30dM+8ML4PmS1VHCW
5rNVat3dHgg+HchRGqDnzkh3x72rUHoJJ9O8Q/ossst3AvvPQ5wItVHVT5pB
MVXgypOjYKF7yXqocOsQpVSrTWFp1IIuYHGec9zTVvJmjAIyn78sC7PZI8wD
Y+8m5zDSv26myPgwexx6Llin4ZzhnqOrTUqbWOV0ARhAYhtHBYpVoMPjYNLX
CVHCa+MUTfGMEZ1bBoMBA1c90u0HESN0T4AmgyH8InGSb5Fno6auHZKXA2b/
XjnKwvm3AdyhEfRdHgmxIK381g0wIN6+yg0YuHTDNRKLQT5oAe90BSSVrBhm
QhH1VtmKYo5OonnsVdjtLzT8SRfPK7rYwtCn8g/38XlJzjMGC14lb9VtNBH/
yZISBQQ7zmd77xiQzYOClOXalAtcJkDlRBZJ0p5yCK3YbARtNuquFDMihb4q
hH5lvdtTV1ibAipng/e1PwRbL2vrMOUfYF0uvF2wHeRl2qWIQbhoBzYVnVVX
taMN4m0SM8cy8y4gDTOhlwFk+PGai9YN1cMjqjp00239gHQx8v5gvgZt7P8C
5xw4x80LaJ9Rp0ykUXPvJH5rUXpd/42SYVQpnO2nJ1KH37GPcWGRggIF/0qC
ti7dNbSxaJ/b4dgXU2BIZBEmPDHtjs5/xBbTxpE7GUSDJk2iUFEHAf1Y0Sr2
7szwTqtByavtUR4tEbry7Oiqnd6t84e1uxRkPCqmcFD+1S+HRTOOW5SJWn3R
N2jCPDo0/L6JACLidfHCdfckuQvjbh7JbTr63EBIcUKB5XNVYmUOTEsZf2ux
6thFNEel0+l88SZb100rLVxUmjk4Ow0WGDiQR91chg9V4powp+Pk1xI9yrLm
FCJ4Fv3t8jXSN8Wsi/y47XSjXsAnnmVdXvVsIlv0mxtEctMdjDUnVK7iKdbv
xqb6RFjbUiuKvQOfbQu1+0O5h+0SzxGX0F2m/VdxyH0p/7WUdP590H0sySa7
uKB3sstpo2bl5et9Qu/+H0Y+AXzYdcMk+Sk7P87R1N03mFEqNs9aeJnCv7Ib
kHgOPoaKL2wPvMX78n/zMvYyj2d5tvlLPKcCpWEV4vWcLTBP4kxkVYC5Av9l
AkuFv8dl2wEF0593WtRcieALI9UnkIBTM1o6ogcuM/MOCYQQYfoM9tJvAeEN
h/KTrYs227XX9AOaq5RgyIxs9noCFM2D/ChKH/i8636h9AP52X79AEOIyPJ4
xqqdosJoZ9x0ZNW9JIiYj2p27ugQcXUqBDK6Fiux4hxzIHGOghARfb8Zu+fJ
1eW5CJ+auG/Z9EnbuvoMwTkFAkUibme+EmeTwVhEWsCtFZQIBRR1LeMXU+WC
aEpLTbf+FCnuxPw4LBnXLEVFUFctLZD2OCDtc/ELaw+i1RqFAcI/896k39eT
X+1DfjfqBqsI+RVO5pSQENZNCCVY+g7i+VJzTxrU9/VcMOyQxNog3kN8pKoy
kj92REkqn/xlMS4Ahu9wkukfnj71vB2B+GPEa+h69dHsiPN0E538Lwg7ITkJ
XZLthduJXccNMCEuym/MehVioGPcCGjeZtKPDwV+R1U1r7fyKq+Oooj0KrnU
hVP7qCGdNwnrZLx8GrDsealShvPl/jlMalELPMZL169n3nDOAxFeEjM+dQTI
SYuboAHFdMVHfBG0yq0R+qCw/2pIPgJ4Fqlu5vWIQRPMRHJtO/Ur6bbptmxo
kAF9QMX2GqCqS3D1KXmaF/z0rk8h+jkC9T0fUL1arXvaBS5ZhWjie7DCQtbT
WlWZ8SZEPiHjExHXafA/SAVvXWMCpZwGoeSMLPAFnTgVTRFEPNKMrSWQre98
nb9CVwDGeC3SmXfDl8tSrxInx5T6WHjh8fPWd1CgJsPqpWQ7yhBfacYcc28j
JIAYb+iRAihVKeNK08bmU6yP13RRdSy/nl9xR2ztGwhI7HGU2NiFWr5u/KFX
xftHWLRjqCzQLPUVsxkZLPYMVfjsja75vlvdy4T4I8Ilvf914klawCNfUH/z
6SEnYem7cNQr9y1XupTChmUPiaTpmNpnPcu9Vb+RXqM6c5/nFyOo4xg3nudN
UG67R/LsHK9BTB5ZLVdoSkNvVt2IURShdIWu7VzZvJmSaM5E8x1aS5z1N1jH
CrSpkeOcC892Juszh90Gyb3dVzZ/s7JIqdZj52LyT8y92pYdeB8Ei25Ez7pL
fWZSyWjGTQSiue8/fkuVk+/SzQnRdmYfuNdzsvar1CF/T7zQukjzgTVUIx2J
WAAE5Vf+ZoofjrI1jpMAOV3MYsoEDWqa8F85PB7O8dmRY7Mwk4DFopFE6JDN
Bwbru+kDye+AEjKkyOFE13LHLWrbdHoqgwJQv544yL1lWPr4Bx1CPmeec3mG
egazlEqa7rRiOik4lSkjD9Z4n/k8RMiYQcyjFMk85qMaBMnk+Wdx9XQuTd9L
qTumPWFs1h2tfFELos6ns1pxh+TbaiRyq8pYpOP9YT/DaNAexVaWIyLinuZu
uMVOvvT36MHE3a3CnsVAtKqiIwD3vtpQ4z2mgpypFdw4bLR6UlVkxkh+zt0O
YsBWkIJq39FE1FHQWQppTLNDbCCcvGpkivGGSrFBbVZQew2j2BrYU7rPKMdb
exDGmg6LtRpEmHvTAoPkFM8P8DVwem5Xuss3iAlvrEaUvcSsWeQ60G91IxJm
3vi2XST5+0e9Ffk3awZ2ENGvB6d0qap5ZN8tjb4VYJkqMsKyO43CzbNqTDQo
wKLW+h6bG/curbHV5tCLr7ctxfqItIetyraZpXAT9Dp42xB2VBlAuuVnHYrC
aSuQpOvyJBy3AduUBJILD9sL11/vgyzDZk2t/fLoZEsUveTFkk7qRsSh1NL6
KoMkelnYOebTKAkexVHEZg4mVORFCISE6E9UJmqQC6a4/K0fX3TUKRSRkhNl
zUEIuMl1hETGtGDk0gQiSSuV0hZcHMYH56Ez5vPoWCuXT71aPtOHrfwn/rqT
cUGRok/VY5hMLYXmsRyUCQTWpkEEB8mDwQtYTKOVSPlql8iGt3QTLE0RtAnT
xR9TU9zEd7FGMKU8lz/PxWk8jlwRNVm5Y38YPwqdH//y+rGYGAOs5aA0xfjG
oTF2mCuSQq2JSPXWLG2VhulPbGDieteDUVfyBss2rBbcTrgPhmJI97dqpePf
UTBl8o0WUdw1g/66Dn+bOYCAt0N6D6Ub0QUuIoVA6x9lHHcTJCfmN0IPOel2
HJqNWmMTtHU2f2jFqPc9tU3v3hm/oKcLChiG5AdG71jgGN6J859SnSXTXHf6
SR5jGwstb1pschDwuLHU/kiQ/2roU79vcHfz9R3qG88lzSSVj2k4N8P26wsC
i6eJskaIkQvo1rltz9Y7DbsteNA9at3ulNQ7AJDmqUxdBfrK1s3xIQQC0YiA
VYO689ONiF9unth+UJg1MusFHB/vGNdUW3OjFicA/VkdjB9iEh2yTJIKEOAN
s4VXb/PuHRR1aDNRmba5yMde5XkvfvELIqfInD+QnjILf5wPaCrmRsIUhL0r
DInZW6yWrpXLQVD6PScaFR69/FPjeHJ3vN8SyfIsQWl8BmjxSfj4n8+YhT+Y
nLJO17iPvBiZzttfUnWf2YLtMf0H0z+umS2h0HHndKInVtQcdqgWfABwHuaY
WmYj9C+aVsXOJSMJ/jxSh+ObBJRnwNy4ayvMFkEZivldCpRQWQWyGGRSHDeo
VvX10nc9YIBQ2uclOvyTFzWjx74ouAdRpOtkvSjJ2Zl5RDcg6/R5+XjKRgN2
1ek8kCtCxhv8yjN7LqE4DTafqGQ+xdk2JmuC5vUsP6wwdR+2Naxtng+SiVk7
CzaJKEi1fuLJmzQPShy9VcBVd0yZlND4DxSxKlTHsIgMqG6NTGq0Usr+Cd85
o6f3QjHg+HBaROTB3cVpe8J8LbPJqy+nCumcX3ow4HY/uOvdZ3xaU1ZX3Gey
G8Ws4zWxvSLCjjcQv1wAp3/kCGfYXhKgEKQrowQhwpqExAK+A8y82jaibio3
Hr1osY06yeDo2yChwBK0T6GeqD4d5qMLqdRhldLsgaOP+loTE2JQ+shueRsI
JUB1sUNTnE9/FVbvlgCa2Jv7mtT33EdKk6yH/Ql5LviMDRjniUaGPDDH3QOh
H/RdZMO9xEP4twZzUBn2+AknuwIWvR7sHA+n0T/1KtFBIJMjUplBB34hLkYO
ZB9/KCJLYI2my93rTnaMKb0HO6G2a7z7/MGlr2Eoy4JMsFbR94GYLKsnwLBp
eA5J/CFcghqWQ23djqTCC3FzhhYLPNDsFXC22BIiJ0YV4CbIicSr9oU8T0hg
JL9fVHj9//gFi7IjFajVZeqRhP3+PC8ZVeMca9ihMc+PNvFTZMtGGrm24n9Z
eAf6+7VaQrmroDoLgXBQfyEcSruu6+Uuhsv2R27yZFAuQ1hpSY3LMYpkvquO
k6VTwNtjcJNjczuUaq8sMxShOkx+ylCBx/+p3DdoglNRuw4xYaGNuPS4S3+f
HEOs/0G2daLqvQykb8XNmLdwzaCOhtC2zVaBiozpvd4h+LiUD37DqcjGhmMj
5B75D1VJukOhJI7NDThMToxonY7TcCTgQLSB8KVMSNSiWsB56QSfBkmoz2s0
IMZntLi+nQZ4ACabgM3riDETg24hc6F6gNqsecb2SLCT6f+2m5XCH1LJH4zh
Pc/UY4HlCndNGuYfVg+wICnBMz4Nr7lp30vwgy0w8NFsZdZ3BKytF32AE3OD
GNUinzkVKDK4beW166NmvDbUGc0eNeDg3xugKR5j37uAOvd59AZR3gqAgq+M
NXASwwR7zI5yiktS2kJcSLErOJrkwGcuyC9gg7uvXIgZmIBdndcfmG3XkGMD
mO6SH7mqmAutCcm3+ME3m5tbg//FrdV9Wo1NuY2zuT3P6YYNODTEIyq3JGYw
rlDJp12mkCFKNiYeVgW5Td+65cdU0F/+JnlcB1DWOTFzfUUkRvnax6RiFe6p
phIFijvMWhP34cEUpKhWhwPfzeT1MBUYnP7gKL1r2Hh1+x7/IJg8u4noYBfM
nH6rSh4pAtnS29rlZ6PsmG0ot7COek0N/eJXjCrJD7c9gqs18YUP4LNVcEpy
q+bB5b8HUKyvOU+4jU4FkhpWO6zorL//kXMzt16ISfS4EzLmBXvHtE4wnRvi
jGZpMP0dsnN/ryyYhW4mybv1IzGAI7m2cFo5EF6QQ9JyuaQ6KIeYwgd3FF8U
flQZY4qhWyuFm2gQu/eSAVcnkRL1FKYhJFUWvsPloXvvESYV3GB7m6GrrSAe
Tb3X/8TVFewu5v9hKV4fi3c8ZVP2mIAyyPXiyfK/pdy+ZRSps8FQHJakXRyb
Z1l6g8bawmmYg07IiEJbYsfuSSFaC2L0E50PXjPwk5Wr1A64qx9NwHwjGh95
3JNhw5laQhKAgScVJhrDRwGiqmvA3A+4Q+NGgIv8M7m/wEwC4B3vKXE6bh0Y
n7fEQjXlm45ylzJZc0VJmp0LPNZ6kaFsxhpJ1xJyaL4XCGn2fE9gwwlZP5pp
Z4VtF06opWgiNFUqxSXvmLe4q+XRHxV/ihKoJ7TqGgvulw6pXOhne10cFUL4
L26Xpffx6CLE0ajrI5fVa5cY6kEWhRouM5D/VMuoDtndylGuob1ZGi4T4UTg
8puOzvfOo4wTPVfElOH2rdFgjdM5zh9PpsgYEtDQgVAuEacW5WMoow82Oan7
ztx+8cNSDG5sqxlOz5vSr9nDDGa2hT79KE4H2w833QRFPil3Ls0ILMNJseIC
owLe2g1Q3ptLfMzsRTitgcONo9889fJnwvTBVrlKj8inydvP1VlMK5DIhi/8
AgFHT9onfTw15Zu2S2bsh53YON3J229PZfUMAnqRWp6lCgEDbKM3HmxD1L+s
Y+t4XTdDMLr0x8Ssk/Lg99F6njH9F08dMUzoIS/MKRo3ynJq30XlQgXC6N5q
0htPUuCFCAB8sSvLRC+4ttCousPyNDG+4mmBxgMpwf02f+F6+xbsDTVfD4VA
jhfOh6O/672mshsKNw0U5hIoyOGqYvNO6D1MPVim9pEivarEaUm7H4Tjs11b
OEC9dp6/yqfecVExnrjFFZflIq/wTW5cGR4yy0LClfRrGZH9EJGdSTVqmaH5
vI/fm+hTNPp8EZx9XeuPEWwIYCS1zPwECkAQVdXRusHSRh0CLiwvJh4fv9Zg
+w0ViGX865hHAYyQO7o68PISx136/Isr3ikbm7TxBhNSYKHUajb/UwK7RyeO
uzAYMGWQI35EYNCsHymUqNXJxGTgyj0yE6wX3to6o/+PNeEdZGJ7m/KkWXu+
hpj6EjQChX3u7vFN5/EdhbsgUSpQJH0P/lxwRtg17Mn7Bu9zO0DEdMKVkDJ/
w66dvSFJyu4N2vt4fgbtBsf7jz+2KH38uRgqkBs/jwOhEQ+H04WsaQN4buQe
UmghYohDw48+wQRSgiW1A418r/kaZP0+3nv//CvKPzLyHEGx6JzSJbn17+is
LkDIzIajrpcXz/tXsllbmOD1+icaXmJ/3VnF43d4PruPhYx/hCAWPE08H6lc
S5aaFDVkYujgbgBmutMi4Mj4+dR/r5vTMV0VFJLlLx3b6GezNRpMYo46Pym6
WWi7JC+XWB2JQv8trbW5R2bX+6vFZczKfXzgRjfW7AtzfceKqExAR7rFzxfJ
02GJEPHMkWZ+uzoXorcMkEjDQQYQHjeQ8xvDA+rFzWF2PUCW3Z29HD1gmGzN
pvfqVah6c6V9t7jr3WTgySv0PHF106PK5OkdlCczQR3WfaPFerW+DRNMP4sb
DPY+kUM4xHhwp3a06UP+forrC46triw8gGGbJqs6gk42p7VLrEeAu9J+j9qR
n1UE5LBUziKw9lO+QNXj7PkGR65jtvT/PTS4mhyFUr2I7W3Bf/HbPudyBbFc
bP4EvxMWyWiye6Hsi9HjL+R03HcoOv+yRCNLwsDl4h8bCimfS2/vd4Xv8Du3
lhDxntZexLUvRzUKDb4huS3627+8K4ZDXeEv/de0w6QnRy0csUJjH5S070C8
JDge+TIGoVdLHpprSPgVmRfXsU4uzVgaEH0ALQ6XvUz6uCBEm4GjX9zXLf5s
cL2f4xUooSvGFvmTOhsoIbZoh9lOVnYjLcRjoeiZe5ThOHhFKJeZkUOkr0K4
vKwO4F0flyGu6KCpJ/ZJVc6ZpnMpnNlxqoCLzr+P4xzAEhMu4F24gdL+XqEt
hQ3h4sXVa/OQVFx0MNs6G6i0WGApaId4TQz5rDxBhkqK3mifKsUEOKVP4xa1
rldWFziOi55hN60utp4CN6tNGTokxQCujeyqKvD8z3DTJlV9A4eCaWMUt881
UpHX8q9BNthStDmYJys1GzePVuxGgXdqE/KLmJqO/rjw4Bn6b8iUjODWASYs
HLw30K7bc1344iYIDkcKg3woIdWPNBU7zkcPBdu6uULY1aIoy3x3JKzrqg3R
oDpwGu1rLAdr+m4VfkXJCj+ST3lyGMRp3OTXZhmynua1j0Jr1c+qfp3cVcFv
76IATdDjIaOoXE6DQC0EKaSCBa094cOQnRg9NXN+lcQ9sX7zqNxkHJkrmTjQ
LH3Ey2bDoCOsX1jcyR4WEJLySbyrwcLXr9dPzv2fwNV3OPmbjA5eEKQAm9qr
7luJF8gO8ctwQNVjecC5gvc/6NIFrjxUSXl+YuKoiC8+d3eo27NvfZd5gGJZ
bDaHo4uzig9Jpbpkkn5wQGPdnnhUmLrmn/GZTckIqvX6yugC7hjhp6GSLaur
UrM2ve2zmuGkJWL8JrNqVq5Zh6Ijux8sscmub1wMYz2VLs9GCUsm6wq2GkSr
GB0T1YUP/S1p9Fqf21Pg05dgg0OCEjUYk99qh4k4M+I13eHU4VKccunVTF4W
+pvVBHU63mv0uHR5aZPkMm1fgrl6u8TFFGcpeOWE4zAom3SPmNftzlTVA1tq
gmDeXlL+MDK91Uw9wxON6xdMTdR0RXbdsUywzgdG2SKoybGDOQRif0r1HjM1
XgjfN4i5xLgNNf7RyY534vFIZgqqmcbYKziOytLXB9YftruCwCO36sldqKB6
pBTuRlFvueW6u3vb25s++njb+/k1oQ61+nJHo5+eA+CJUg7cNlcAGmlwGX0C
ksPodJwUYqcItGXaoqbsh47nVUJN6DyzIs6ljXy9z5hhVsTRzTVSGpy986Tf
jaO5f5qp++v9cE4/0KgVNjSLF0VdAl6DdBA6Z5trzngdWPcoJoWRrW/BPqea
atKzvLhAnut9ndB3QQcUiIn+jRhpB8Z44zywbNailq7SvYAeleOd4XuJ3i6I
RSjEEErYc6X1JRD5+OPCS0mukFkOYIfF4Cm4SkugjuPjXRvTHIkNOUoCXxMf
sOTrCOHyp4ReRTMyTK0w27sXJA1wM8ZVyWiA1tWWX+WZ+iRmaDbblzmwxCh8
VALf35IAqJyGZzWEEgXYoioDQXvHbF2ui2lodJwYAQnUF+HOFHRX4k37+3qI
Y3eWQusJC6mG6sIwrbinU4z4tONook3Og5Jwokzmvf2GKQnFJ1PKlK9eLuGf
5IiNhH6P00NqWRXw3eEZ17aAEq68s0P7v9sg9juGikK21fxJyKgzs3J4iMSw
QX5iFzgIu6/6QFZAFsPtMqSu/TQ8oM9Ii+aWMXVCZ9dqZ0wI0UFO6KGbN47h
wqA81D9kQK5MDvrhLen1WrAwJXCkuHx+D4yWQwU2HTqO9gzDVBJvsZznAxtP
doKzPmn8crcbNexOo30wzdVG79JHlk9hoGbpn4SEIeBEYO3VBcTL1YxG7qiX
Pf1Q8gqpcZCylrzOwJeEI3QD01B2QdQQUItWJclfQYxP5yQZkNwomZygSzxj
+ElGivQhIOKdnx9i8yOroWof+wXXGBJymE8Epz0UE0k3zLpcmuqEPZspU6KU
K73E2I2FU+BzOIgbnQWxMFiULEnBFte/l9p6r+gRq0sefAejHzmvV0OH9mhF
DwwhkdfIKeXSZOtKIm2Pk7Yb3Q7q3tuLyHgaBihWe/ObyjUxKNBb0UmyYkhG
KysE0ZGGPGLrzsg5sY4yhnSFbT7IFhknR5jsA+PFf7GrbKP0Q71YnN4Jc53k
+qDzja4IgdrbLV7VphB1WYAPyoAAxI8OR88Xde4FymBGGKwdWsozGyEEfZVw
Z1Hw9Fx7vK8d3QDvZ1zq/eO8+TzY5lVV37sSnp3jUdyJf2VzINLMyjFxGv6f
4TTdZAenbyLuypmPyIxFK+8k+fZuR7a+BP7I9GEaBRwvRx1g/1JYGD9bFC1N
JbtcYFb2YCtduGwc/hRBEJ8HGeKV0VKEkXY92ezRtafFjlKLoAuPjA7VFh+I
Z41d3e+COwff2aeAcnqFQVglbmIW2oSm32f3fVHMKo++Bu5k5HkSXUDQTicB
XUJbmS2a3mnzb+UvpqoBaPPor+4rurtWr3qth1geHEnq0Qy/eoshYlcyoG/7
qj3ZqxiSRYLXq04iUqBwu17EqliRWyOdK1jniaGZc3ZpqyBPYuLvITZhwQUA
4JyIud/YdgHoacpIuHnSN7OnZQCDy3buKdr1VvGLE+TVjW5WEbXSB5Sw9E3b
Z5qdV7szRcDW1wGtm3bu6H3/35+26T1QwUiXIx3o1zVl9CMQF7j5eB9ztr5w
5H0yK1iy6vXqfN66MQWxRj3XSpqUVedpIlDj404of12wa19z75QVx8BGyAHj
WyEy0xio4eIkfsudJpEAQZ7YbYDdFL8tsRE+mi3BpORlNlol1/Vwmy6sHHvi
Q7OudnHfbPesSfzSTZW+XGqtDlnasd8z7AptgfZ7QGhDwWLKRj3pSfPR7KhK
8ufdB1DPEqPH2PzrUevuw7GxxJFWLdpVlCB5PSwo3K6cXbtlkMQClbDvmkWV
Vfi6sM6iGoNGJ+7NfXPToZ5+5dKS/MxaBbhqhpsRkMXHWX8dXRL6oJi/fmRz
QeYCYyqqSzvBycXvJA14OflXUwH+LBqDq562ezltWOz7xkq82DMN0zy9Iwm0
32I0/FaeLw8aQLNFdXSkUzZiS5CfudKfXTOoXfufNZqFz2NyrN1rVbyb6QHy
85w4HVxMLPo/sV7eY8KtslBfxwu8IIOXkrq0FzeDdsgFjwl2GC8fuC+lGSpZ
dLv3+oN05yUPnGP6rUjkxgDJEkG+h7rKIuYd1uTFkVRH70mfLyu+VUfTba1O
3sfh0jCNrVk65beNQwp9jqIAGVGysvEntCo2/7N4DTtC4nG/hbQqKkKwPNuB
exA3yGOc8yiLUbGr+Cua+KL3JCCevXVaE7sQ9H3tJrW3wmp+PIFZAsuAzl4y
oVeOIhMa9VrfbNXNNX/jQ6DbHInrl7+rgehxXEa7HFvYGdrhyhTsTiDyiq65
UZZB5aBrcvw3xqJT5dUDohsVB4ypClryafYY8gRp+9UAPH5FTGgGA++nLqQF
ZDB6/ADTKIj38a58fatunMGFIe9acA/Yaa3V4ev8ym7Jdz8MxxuWcls+5ulC
o+JyS6JCZVushg04MxPKrR1x0XkIxFrWQS3Lhjll10o/03vJrV3i0hQm7sge
KZHGMTKHLMtijuh+UuCnM27S3mDl3Xd4Ne0qOyajk0JNwoKQriSmipVta1lR
EowR9P8OKOdbs0oRqf5lAFbo1ZiT5+YtKrj+54vpvqwYpOgtQ5XNkfC8aSsx
E0xa/NAXlWRVFstX8SsJIGZe9Ll8Tq4aIlQuNpja/SyRAhwa2PGeSxTlxCUl
IudMZDwDJdTEx2xJ8WW2TZvx56+k2VYPrP5tikBfh1M08RUzl/DZWyYQWxPm
qrV2va5bOhdDba2h7gpI5fGna0T/u+s2QtE+2RYzLiV3t0vm5+CYzIkdvRwr
kJJiw/avzOftWgeppTEWAhnDATRgp73PeeuA6TUbggsTgT8aIePMdWo0no7J
JLks+7GyLC4MhI7u7gAqpBZy7LcnxQL5WrYE9FLyliOIkuaCu3NtfpSnwoM+
exl81+Q+Dfhigz+Dzl4YxswxoqflxCpyUK3GNQRkiX4buEFoo4i5073dJ8gN
LXiR10rMSjsFIpD1G/EWhvoEeYzy4yNV5zRfMkDGyyjmhcuf8+uFw2jY9ijT
NvOjz1TRCknNIZoS7w2ANLuX9+hdPpW0kCQa34ldBxu/thQoK5DzL59RB8C9
AZ2xtd2+sEZ14X3ec9OHdkYMr/mBBAOtbP8YaOxI/bdkO4MyprFc2r4sDhOZ
paRtMi7OVDWelt2xznKy6kJ+O40oieoGcDnFLnlctQ5pRbW6witJdsbju+O9
lhjzZErD8R2OXQyXiVCAuQNJl6dmr+PGqMwQcyPYMHGF8KOnn5SEw1OViVET
umYxg0291de4xgfiFuJpKl1oBsbeudRD1v20CDkrXNVB9RsI2cPaqDPHyNM5
U2BVvzxk69G6fY0ln6hbljS77si/+9vxdPBpgA5f6/6azIZZikvZ7mble0qe
ojfZCw1YZMDbLJLOP7yswrJFSJ6FHX6oD4Jx0RpEM7fJDRYvZsLbRZv6MADY
KWWg8HVovHJLuvE1YzuqcTpvk+PPmbObqdtTs8kk2Y8fDhVrAtcOSTEDYMGh
pz1se5LrMgPWKKOji1EDSFuIdIP9elEqBv343SQUrCtGWjp1BoTtqi6IfHQA
8W+QXcVBc0MyBQr7FG57nDuv1c3qmEP2Wuz0sWdIsdtfFQAKBP9phyjXbhJP
fhulm/hOwgkzNq4+rW3mn0Oj/rQgX2EvvFBL9nXiz5N5AnAesNVVk76YZrIV
DYGob/O9MM2fAo95fOXKhrTZlS4+sm1POHSfGFnmMQcjnom0FoMaNzKiZyEZ
l6ofv88I+UHPo9fPgvpb9VOSFpQ36Byh89mnx6gOQPjbUlZ1b08Mp+NGJte9
fg5KaujkaVKKEIOQ7gx4QjVPG48TcNlN5j4OeN+UE+KgM2Kh2xNg8wvOhog0
NuKDs6raXM3eeZFJJFXxPBxnVHlhMreuMt5aYvwVdmQfYJG4lBJZr7lOgskH
Jl7oAMIE/yiHNW6PXLTiKzXpDBeWuZvCfm5hR488yiwrDTdCLhnSl4309XmQ
SwScFdhDdDZM3lHBwl0KezCxC0ziwGw/KIoUkU/hCx6RMgOdj7pTHi6nFmux
xTg5wKt7ABcEXpUuVsazRqgVnYlU6NGWtJQv9f+gk5fktrAuOUB3vSV5t1Mk
Mb967FRTMDSaLOQ8WYoJPg7lnvCDS6QXsDRM6EgnHE4RsoTmXmIxOROCc+HZ
l3kbc03m+M1U3sIR5Oiwe05nV+WUqfUFHh9G/e+PfnxWT9tDMUfGfihGTQaz
1Xd8z6Mlypphh7NQU9NaIBIhQCPKjb+nLCmUX23OXnOALCjmhA0LFSyOUC5J
ew51aJOkhiGEn9ErRsD9WdQlSniZE9WR893QzxCsf2/pz2g8KehRKh+ncLtR
iAM3hjw/q4cUDYIXL1elkDFHEATJjHibDS82/k9CyXI7kVF9ITCtT3E9CytH
Zd85y1YrYop8zHBQ8G9yCkwzGNE55J/DuEMcuPUFjYlbf9zaanl5DbmmVc3g
IJskKqTv/TFqqUdaMilrq2v4fVDbjBBqynM3HtpisSlh5Fc12/WJjmkhFjws
g2/N5w5FgYfde3zsw/nVxjmd/ojM9yoqKje+MRVm4aDaH+XT3jbEbav1HmzW
8/3FBJ4u43FRPnnM6cCeDX7tqxyAnLABn79wSak2JEqyr/qxmPRWOUCRuqee
/AZje05Pq7hqT1CsF3uGspEpRpyHAHckA7TqB3f5DScasac/PFJ0q1rGA8xq
5QyrmJXbibS0Ii0hY5lM/5GCKHVoK6l6MFYzlQk3RNR/KU/JFCgvtsTwmEjE
CBw/ktbdKG1u0QwmpI3yfgSpm6pQcfkUPZMR/oiYQAME2lDkGsBOzGeCJf8h
ADa9pI2Eg0rOd5PMvM0V4gDcp/uuKg2IXVwVYxzPqCP4FZiXX+3TZZUswG4P
vJtHHEBshYIFbx4LTWEKxtMl82NyJtTsLBrJnyQUprFpXk6fuOfuOmravH2b
ErIAtdAlbfQKJWnPst9vdz67Pfn/c887xUvwj7f2u6GTGmB9EVIVaB0Kn3jf
Cccxzd76oXFK2UOk6og+H1mXvbmDfzZ6jS2OtHzBSBTgalBSBikzasxm0ODY
ZFV9/s5v3BKQiOVQuO+tVb245a+sK+WCCAcapAWkrBrnQ41Apu+mp6wzUOx0
ILPyGbIaDwxgjwjz1CDSB03SBSYkfW9qiG8C5puGwv8DdFDXOxmhtiSOv4IF
zzxZGEZh71m6Vo/MxAIUAnMGzKdXITcLMYzcJDyHq55InvYP7sz2/yjJAKrz
+eROdlxhvdm78MHJE6oEtCSIVMVBKvUYMzyvv2zeSDKh/+hPargLdEiyTrnx
Hz2ff5EPg68osn1iq3cZNPy2kflNDAmgVuU+vO5eCzH0icWQwGv2yClasAf6
KlFd3wpTSM093FKrD3k8gp3EdfB52bnZptsu09MY+NrsNRC/WnuDX5BCxTNF
rpn+jRpa7JUA7XvbviJYimJBb41r97uUPyGCgwfrTSqOwRR2WvmgtIzHhv4h
TdvQXwLKD2v6GIUHQOeloNHJrDPrGcxWFY86zIbBJC04YBVsW0bUE2SNYk8g
NPU2KgLeZGetNYKqPgcpKKczafEKhgOj9T/moKAhdF3zx7rqQg9wAl0o4IzR
uaoU+D0is/tq7ChkIIxj0FRnvM1W+R+EZUDw5J6KuOqJ+zZe9oEw/qgoEAbe
wZpZLe3U2vQ6lXHO4D4Fv5rCwADID63orsf7O5KIsIvDkSpFydeNeS+XkwBK
l1dmM7ndbosXyLWWphnhVXSm25GIaGdH7vrtf67USMLWdTm4eaQtEtIRfcTt
dWcM5Z/GE0w0HUk6PA4QFsZ1MBnyrofaz/rE7ZQ8ol8Q6W+d+2/1E00iQlkM
coNjv65/lp5q2DTVMefN2YQ5Ao+7CoFoc8nfXdjFqcawFFWPYSEyjs7hlnKh
KsnDHcJux1MoLv8QqeOEMnz/Fs6LI27yduCw3ybAoXyzmfQNK2slx30bmVBb
1Fmt9Nq9kEtSYskkeSf6emT4F7bupTNiRgkL4XcgLsSwYqszDpgi2fr0Q/K2
xJsDbkhCKWDHALu3ur0lHwDZEMvwHFiGpZGJJ5bmMwbJbzdx2vfX8z2Ntu9p
YmyAFekiYUADvCAl2FavtLfbKs4ZL8bEmuNwaPakzdok6RdDSOzMrb1L5rV1
YNU8oIs/s0O+H5/bXw6me0zhOk/a/MWGJ0Luh/y+rLQ7RIgNC4jJ838J/xDx
y3Gzu6DO0FKVZ9fUs4X0b7+xBwlkUAhzjQtK6Z2F5V+0lJd2Tn0lTs6Is1U0
0yNO+rXdSi9E1YALqczoD8uSdivtSY/11i1Wd6VJsz34ltKCqJFqbv7hhNeo
QS9jw0rk6ePxyaP6yJAN1PQQYO6M15aDinUGCb0hj+3VOxemis79hNq/39KA
GwbGdcV+NED3w5I0u67/xQczGrq8WLDo9OznIzjmQ3IZIEeeMKz0SDwn9PhN
cWOE2UqzARRgrZ4JBMXs9B5Hmbhj8z/eL94DtRQGcLBAypaylRQq6HZaLSDl
qorXOgnR3HBqNu2ZPNXGsLQApAPeWcmH5ClX5POuVl6kHfEdkv/EHQ+qu7qw
jf4mz7SJFkyBi9UEhYzYRHtlynabzEzqlTNLuL3iQ+bCgY4oAN7Ddm2hnK1p
QljIoCoKirl7CMnlvZoRV8rEcLOv4sQ6DR0pU0hZ+ynDXYc37FfuWOzj2zEd
kyTD7fHf2ChNRNbYOZqwzhjZvSN1fdpHIg4k2wYZdoaOKO1Ibpdb87+sJs60
STA2pTtuteIfaGZoI/lxE/+GK1Afc8QW9IHJMVa/0XyGTg6gjLBAcq4A7Z9T
+SqX1C/6qU7FZHlPWr454oZfBXPmgsYEhyGSF5NbL18vy7AHv24pkdDcJH0F
XAphCh+aLsU7SGYE6FbYepWkPBCt8xghdiUscrPJfeuhvfbTAqtXgQc4UfmB
4ijDvHaH4jbNxvcw2BodGJji5+2ivJw6ZsT6noD3vWzVuULqw4jv1EwHRKOK
SxvnCc39JYeEh+vWwWta5Rn9l1JTuipZzdZPJaLflznIhX8VHz7JwVu8mbpO
S0AyG1heQVcyfiAHXt+kFYxOSqpgmY6C0QzyLmxXR5i5XvjqrGL75wMnesRU
MD5xG6u1h5av40p32zPC2xCzrBnYCEzb8/RFbKZad7l2PjTm1fg9RJx8fYDE
ZoqJTanYBAG2Oyr+ymeY6krJb89ME2i6q5pc/M8SGT6Cz0gLoKfl7SDYNb5V
Hv8Z2ywgld4VC2G10QZLl3GI/+pAl9JGJDulOyJxVIOA/fmpbAsI1U06WRSS
gfxgrBQ5S10tfmHmrli0s3LtlU3JbFtCKr4zR2bIo4/g8Pz++FDt1Q/2C4nF
eYH6s3dZwoeKkk+mp0oqaiqFum8SYOwY72vh1qlPL9yxGzGoBwQSUYGG4vLx
QN2G8uKXSy8I3HzVQSTll63M19ZSVw/XXbUYfL2o0q4cJ0aQlHn9OUVqNvee
5ioAPUln6g35LUZ0YPQ7fNsmfVDszA1qvmQH8gA7QaacmUreBuZQ3LxXw0Z7
lKLvqPCX/o+vsgcTuEw3SrIxjQ3naHoG3eeB8f0Al7MvZBX8wWfNIZJ30V/F
U94hn+iClMJvzkiTFDZY95uPBLLJtGEy5MIyAzHwgbLfky1UsH6bBaJNyjAu
rr3g+nbIFK0MFevxaJEbXmt/vXGSSDEl8ierVMMk1yfh97LMLvlPaJFS4VjR
9Z3BmcU6F0JRFuxGXov6lK5ShSBpxbcHkwo1VDxa/hd8sRNQzh6P7KP2Yl0t
9/RewKjvgHzK3d8ONGOk0KQso4a6PhlQ7yHWoICmsbqq1ovguvBnd4k5EQqP
vGkbpMZki0c6FdUf4R9/igdjAxCiPBJ4nOoaRpKlon/S7WZBdR+SXH3iO/12
ZgyeV0aFvy7vWzUuqnl4ApBLWBD1WXb8oqf+W1VNA3hgvZ8pmKUa+qgJN1A2
dXUIVywL4uSoOsfHaZ7ZmvXkR2i6YEd+sCE4Ubk42N/HCNAYS4KLIz1ngj/H
F1P0fvPUJiX0Xk7yw9jI+0aL0ZQ7UgKI8Mz+s7ltdkBmpw7PYwtNEKsXO3Xd
5i3golpF+809BBZ8gq+q4InOfqpNR68isUHYJSx0CUU2j69HTw8nbpyxgAvw
RdxOL+k43hUI2MHTVMHLZQA3kDXWeLGc32gmZGb25VGGKY967Yx9KU7mzLiz
0KJLfBHVQ3hvNKyprLv1tmGygcz5+kAEGbOv/myQaA4atwHibkAMdqy/0Ru6
DsHOt+ZMSvf6hvo+w/3ixh2NcIfGWpM3UNQIfjsQ8gh2s21g9F7/HLqo0lTU
ZGsutZT8pQZldr+krlCEh8cu02jV/3ekRLi76iRbUUAIZN57NSoosjrb3h3F
GqKnzkIr4ob2t8hf6O3otAUQ50EmuAdo43duwmJoqOvdv5Y2uWWJcAIuhkFx
2iJM3p1oRfCgFq/jPMMb9szOYL/0QMZuWjTGuLvJc9R05g0pHOlMefN3syf8
ZthY5WJDvBfejoBsGgpFAnY2gPFuTcREoaid8yblRVkb9hK3tPq0WoQJUasA
+cwGfnULwNHFaB8RAMw+xafuV3nSIM9LfOM8mZv1IDAiQYQBC/TJAZJZg7q6
CFtx9/02a88dgdF5c1fUELO2DHo83xcBVd/etvvm58vrlwfN3zgwlBQ2q48X
vpEysoYthbYFoNFK6Mvgiw5SoVlLvAPTapAiB6D19Q3WbCldHzVnb0DM22oY
Bj3NzzvFgD76rycL5j+f5VuS4bemnLyeOzljBZqP6buBY4QkXaho/uLGnYwg
yjEx8CI2lo/4ZW1CYVdyCEdQpgudXtLINSBVaiOkGctEUoH6fdolC55UEVOV
O1htQGXx22hn268CGMA7I704BSQRSGZuJLfSsCiDt50EpPgG+zbHbob1E0/Y
HokMXcPtZTgmY+ovAo7Sal0Ch3LRJnLd4JMtbE0QSO8aTorgi4Ky0XCIrMS2
YC2/tA2nWW2bTnelSb4i5cWMt9eYP88DRHhS2vbUWX8sid+mwMs27EY7coPC
n/Pyg+YNdKowgYYj45/qHjw+jaP5CAC8X+YRu8GQRL0imAbLeyhkPsRWEoyE
jCmJmT0mAgbGv5cIiX/ai+5P//Q7k9xjc2UXpM1UfbG2BqpdH0nUKaP+6n6w
mjxi2hqVjFjpKRqgo4xLec/6HfP4msD+5zRzWKXmeKg1xNTYswKiuehqXkic
eOkRT4rBvhdaCTUIMLf1h30ah+G8mL54HVbje2RbsThW9bPYFK1Oil6J+mKp
Zn15XFnknFIbcu67CAEvmFYSlivvub/kX0d6k4GQUAvDs/geQ2Jcrf3/8fSL
pY+nt1HD7TZDqRdi7T7m43SVcMaCxJoSBjTVR+2mBbolpim6h8IzKqVvdadk
fVyRAqJkPvdgk5Rv6Ap3jniqDe27Uth/364IJwzNBJWdHWZiUjemX9mYzPyH
wHnkKhkOSh+aPSPJ3mVwQsO1DeKaP0v5EeeEqSy2XBCzV1osBQFXhNvHCGmJ
iNaF5H6CfRrkdnilVQtW7T84IFTIOsLU1g48sgnNnsDmXKAViY7YezG2Cocp
nhTfGlVY7iGYmKRplnxugQpCPh612rslEMaQM8EqaB930dgmSEr5ecn1JRrr
iSJ3E+ohTM5FZvc0DOwuXZ0TldnJEJQLflu9YSWyB1mfmJgx9JaBj6SosWo6
mtEKhVhKNmc9UwGW5kSRaUx15Seoo+IZBUySpDLEr/SvJ2v29URk7AZD91Ao
3XSCglNvzjp8q+GHg5g1PsPV3IDjV7QZ2UMn6gDVte63s7CzyoFqNkd0VBMT
69psgvQzgosPY4MGMiJt1jjINSkdWD0P7DiiQ/bCx7DcY75ukNyawofwTtnv
t2gIbmJi6ws/YfSsC5wiPpoRFGjOmPJ6M/QeHqAko3g/KEZ4SKVYaKYlYyK3
xarVzW+ILihx6TmoSLBeZkgCk872c9LF0bCfDRAcUVF29q1MdvUOY1QlsB8v
fx5DHikkdoW5xXK0JbSSzHks3jhrUoOpjlfzhRCJBgdebCiOgggU66NmFB2k
TctQUFKR4e6HaxpHCJNndtjEEJwkdTDHOWJ9mCYVAUMo41xx8UodhLQ42itP
1cF3lJb1KMuJ5fSxgS0+jJ7O476UdJmMmryVjv7WDzJmOhMKH0+MHmhXXqmZ
yOpg5jCAvW4QYYLmekBuPrswsx9Ti9+Rspql9bIgNWedXowbqL5FBZLa+EQE
3vYQzbsRnwwoulL6Ym7W34HQFeqxubnUzUuk80PnUavpCcL7ljKvbRNbH1Yl
jmm3jPX4rm6JmmfHvdDPDIUBYQOXwDfwQHATuocgxkrlwFwBtPXRqXxJgqkE
5C9vIzdSv5ZJIilS/GnhXgs1eHD5JVdAJiq7wI3HBdPjfBfRjrJRQneSXE4X
Z+d05GKKrEGS+Invps/BkUTKNL+hxS3yWzs85gcLu5ECzXGjIzMIDKDYLu0F
6naLz8VLXlljFQkCggLtTmOfi21whHKJQab/kTChnBc7QadCuuX0o+xIPRmc
OJXRcpPTtiLBieCbfZegPIRfAWih0lEu6nQqWq0dvFSEUV9T2oKKgPhjOV+i
GuIpoSevF0Lx9Bmp85MOLh9jrrmGcnhdhe/MI0+d0O3MRl8qPHki43EHvE4i
2NFfyl83zWRfilciAP44WKnI7Cgz1SD8ypXcxhKROLJjP+fbDxtbwAfLlZLE
yGQ1osHt0GhtAQJycAWyGILv5i3f2sR/GJWIt3d1JWpRDCpF9qUwN1O4Qwdh
7WTeLkeMjZDGe8xmr8+nJz7iMjVeBdeMMIFa0bBFJ6+RKI2Rui7gGyAh09Lx
jp7t3bWHvJF/AKoMbKJkSY3ExplhUNK/z9ISWAllTgZNfhS73c0UnLcz3eIr
E88eaPIjjx1PEbVNrfvMDMt9Y803yqi+YTUaZJPmZqnlyV6SDppQ/B8sIc+q
wtvuSVMF+n25S8jSFqEWmUBqqa96mx4oZKSJiIxZPThVNeePCTCxfeQCpzmd
/h5fBwEwJX6o/GLZ45hHKKRaQJ96jLm1QSqlKPRyDFaRaj7JW9nFmzp5vDBa
V+13q6I9MLto0IWRFH9Koiq1TmGZmyvIbvMwdC5dfObzpTpsXwzWpRHPGBHw
+phc5y5jkOnz+h7VKIS+byiyaDkpu3LiWQnWKXXdYUge23ysCLZwBU0HLgmV
pt6apuYJdVBfERO8pBAC8HWBceNVak0CTJwDbGIWuDje843LOhNqW79jFiRz
s+e3onoXLHfIZj3xRomBq4LnuR7Msn7tfSSn8M2DqmHPNOnLKi60MegvpaAP
Mo57Juf4z5LKm8aDPx2g5gnzpjuHKq2tsoLHwcbyXs+pASe41xcgGgPrDvAz
btTxsk3/eY+s7q+55nZMGNAPyB5gQkMBK8z3pLTAlmspAGfOIWUO+i0AIk/F
qNDdN8uuo0F1eSQho80hIe8EBYlNVbis82QXAh46Xiy2tG3yfVxrgVTfI22d
SZF0I1uVTlcoBKPRSrGBbf/aD62T3hzfLsXcLTp+M+rOtmeiDHHm2lR/TRwo
FZmSOFjNwYrV2AwwiQmudI6dn8C+MYMYZTJWl6HeNxj4eN9ESxQ+xUhhPui8
bXrozr7OOHquK/CkFzotX+k0BIXNZfzyBbTz7YZ3xC/WSz+kxYZBRRwN9gfR
V6qxa50oW1cHmr7iE4J5VDEQDLsM7osihBlazfmmK+6Cf3sPZQ+gGlo2yWbU
1AS/nxkxdFzW0mbEhqSNEqy6q6Zih7sSrs6h569A5mZyU12S/MKYTwkgvkRD
SlMO1mQDpWCaK4DGSEdRe2QXD4Q9i4HcRhbHRKFIbUEQnWJ7dcjcwWdzy3LK
CPms6x64oj6n51RNsyIwydnM1CgF4dg86v1uwwhSyLX5kKlAzhhJ6VIjXX5j
s/6WnRIQSsLLhfNYtDRIAN893jJCqHBi9ha/1H/MtXYmqB8xIvRx0HdS7Utz
avTBBMml7sfOsEJIld9MgNfxCwzHPEIyz8y6ZzqT18P5hExSrbPSO1uGwwdI
kfpzoOQPrEkbyaXlYFm6h81CI6umnk2Im3JW8/Ngb9hzmWuV/nROdlE6v/iq
L5a7ERcsoI/ywnCXlkmCk6uto0J6D2zzWnOBF6y7xsO37UkdEcl9neUAdDNo
DS7vPNbWZvHg8CAuwbNWye58JSt7isBo6eEv80J97x20v0cOCVkj4JkyC37h
JuylaI6LaCP8m23XJrvFbNJUJzh8/5XnQQiHJ8ZEtwRe1+L2qhlP2hVpcYS4
y1xOo2Pde8/v0r/JcD8RfS5F46tbhkTP3Lr4F4KOGoBdA1flZ/NhfTJnbCxP
1XIyqxfa5yRE4CttLSW7hE0vmyItZW2bhj8Hid0LapN7xaprokJrsHEZXEDR
0XG2gVs9v2SUurQSSbQBgAd5/JWt6ru5q4EkUqudUd9V5dN3WdBDYGjaTj6a
++l1FL6mWvJIGk4BtjylxxdbzXrz0ohDvOjaroP0GYwQZA5MNgpkNGUDCPWF
/mULmD568+xOUitlRhZz+gDw5RM1JblSfYVaHO5F676oCMKcVd37E08hJZCm
WAZpVz+uvzS4uAvfcZk+q7A32WUTq0tFe2zLWiZuMgs8SZ84eQ3TRskZ+Q68
9H7gEL6K5508WH/y+2hIwYtLPEQFEWtHbfnZjiG3MyvpvxWGBMGTQB9mIC/a
PLoHlg85GQkT8dAF+WjXhW/yzg6g+OQiWyQ5G6tjQlO+qx6hOxStVibOWOuS
VHpP0f1GwESB3GwZKSSEH3GTnOu+vQTL1YvRG9+y6pq4lnYJmvFVZ2M2qtcB
Vg0PLJe/XZV2FWn6oybVqThxUiU8kxRZ6uvOGNRvFAa+m7GMhMOVGg44RwjE
wU+4hokF+zzr1Tz+IrlQ8CjqQD9RiSCHecIkockPrraP1bUmp1cnEtbYu9gT
t+mXQhbhsY4nxNKYSW50pLUAyoGMxe0r3hjejTqCErCYJ9fGqI4Xm90TdCVC
BCuludLOxfN/DTl69g5Z+tRbofBJFsTpw3LLVdkkCIbgpLfCGpe6f7D3oqCD
ZXDNSk0I2HmSILJNGRLJw/GxftAvutenKh8jKgg1bgVdjjRjj2OnVbKQWRnp
zS+O8fx0MMd76UQ+tNektypBTEt2O/lTBIF/P6xEtE/1ErVL+lUmyU9ksL8J
Eg8kEv+e1uWcYkVE4e6JRE96/gm1PUjL8VCOlE+O4PvsR7HFPorfnZTryUwM
b2ccwaDWjIk9kVEOGNgmthsI2e/y39rbJeA9ofb230ks/0yPkb9uGAtNXrqh
eFrC7CWltyhYfXA3fp6B6TH3xxQuUCfFwOowLbrm5b4wSnSRuZ5lvs6gkLsE
G3zlmcPfWZ7gOFgGCfnMdrAxPK737zykvUbFP8D2Zv5Uwd/YMUXBiw3kPYpq
1P+VsO0vd8DkDYviQNBVXDIQkD4Da+i8LDku+n1fl/gv3dpk6DTzkPcbRfXo
i147Ab/l0ZD7hyyX+iTEauP0DBv3vMU5CRZf0zIDDB6THDZZfcJ+QPoPU9gB
1q6oPxZH2Ejyp1nUdsE70JoIkj9rcrjvQCoSmU75LAstwFm8ChtEwGsxuQjQ
gPxCnaz92snOKunxrC256gQCGIJJPVa/+vOp3igalfknYqJuySA+43eLuUuh
fA+hsY2eHdL28ihNnyp2vKg3GuokTciyBa21DVhgzK3tF5nJ5y792T2W6axX
PjdXauzU84jpyI7O2UOvI+1ZGJQDjlTzptGY7jJbxEAcVbUhuoeHejjQIMk8
dMIV4iqC0CCF2rKluAlZjBuNoNxGD2f766zWYGPRGmPDOcV/k2oRmq9JIwKw
iXDdeyN9g68JSU5FDhsNA2mK4/el0LZfXh8CDFZZkRbgnC9KFo38Lgr/MsHX
h2QteBDxMW8s/Llp8r8FyckDVRm3gvEIx5G7Pp0lflpnWvnz5oXBLDaa/o8h
TdobH4eG77kJPvVIUJ+g+SWtm2dhm/O6XLgtR0cOdvX6Jcloyd67UbDgyorn
/V/a7uq9jQmy5udJY4DFrRnuTYTeWlEHPSqc330YQtgkdT9Jr+RwNrJ4uUPT
7hBEZuUfjA79CU9qR8cIXEt2siy7LsyJacCd1DQ03gVootmQ5qQPRS9cmS90
S54Yg+SeilHTOfal2GT92eNc+mDwVYmGsGdNM9PRn5PB13/vY/7/K+ISNXGL
hDlfxNZlavEC7PYRxgKJiJYacduRweJTCZl9HcxEpEQnYpRm7Ydj+7NMo1n3
4BEM2U0DG8cnh+R6uOCumxaU7oXozfjLRSwc3mFvz8O03XjGcq4/bjxP6AAq
pwP335tBJMf+I5Dn0OvjkWVfiQoqi7gcvQQ4aT3aUUcoCy8y/3QBXVdmvo0S
4XTdm6BvkINBrPkZL/ZeEVZpOTm0SMvK1LOtx6y1iorkrbszr9tKIGZvv0vI
TH7SPdsBDCXin3Vl2Pq2sX+WHOIcCoRaEoHhaM4UE46lHJUanNZHb+uWr9My
6sZ2h1gx9RKLeP0fuqGgzjapagasAqfpWHsvVeL9TEztJ8sA0/c5CoGO4Tke
1kbFbHmP3h77QsO6FzIu5hZiTQ5yaX3/N5wKP3koDy1e8T22b+C+j4vPMPnz
8B1+T6kOw2Op6vfI7h2zjy5fmAgRIu8YxryXuIsLI9KOpObbQkSULUY9nj6d
vQkCfBcMnFJK15XBEq6uoVuNl/sBgVIMNouWgmu58lyaHZoaKFTU9ZxuZmZL
uyuV1YzcONWi92RpfcKl2PeYZFX/N5syMtl5tWdXYrNjkApf99jFabDNormh
DimBrp9+rIGi+KdBaXr+IWijzrkEsrIYKJjNQB9OUxk/Q4zs7c523DDjzvNs
Ddyd4VXVegRT/VJwAvlDUzZ/qccHz2jNMPQUsB7cyUJOxjjvGpB1GMNabYzd
8RZ6nBwAsD0m7ZZbDcz8lep9ZWjRNgWNJURkuFCZ4w5b7k/PADr9DIlRUCOD
B/ZRtyaPiN9g1PpAwOpop03pqydrA+CX1iO+Q/tvLh5FtUvzXw9GEV3RESQx
6Bu3xJuhV3l+jEM5tt4EzCINvDH/eghYVm7UHZ6LHo/RKk+Eyf0jm/Q2ZtgE
6LW9N1ND3ueAfAP0paN8xR8VnZRfo1ugN/328DRTsm1yimdhlPfqjdNgIlbB
H+FKMxtMrjUyIzGigbz0yR3JIcphAbSLuhlH828PxBGW4QteJ907ZU/nlJR3
CK8hXx47QZs8gAbf8VaxhrKpgQViUvhUVkNeTyfc7VyfIwBqcsRlTKUM3mx3
j75u1Fpw9DUEHYvBe5Th5//fiPyvBnkhaR3IDhfwA4UWKdjRfqXs92Of7Ovi
thlIuJObvOnFC1BzLUTwao+0zAyrM8WhukeGVEod8zVRjM3kdmYPTf36HBB/
cMVfwF1NEo7odW8RMpQa9auCBtpJZFwmaElY6BsMD/cksPan59ptzQsiFDk7
1z00hOz4EuDHQCv3yeCkFfYa1ZVqUjrENWNMXie3iABa5GUJfh4jk/QJfelK
1FN1OzCjlSXH6NSM082coE3ncurE8FPTKF8ZpRt0DR0QzsK2xymXVEWMAfru
YjTBRzX61CSCnJhfUIF6Bd+yVDOFXe/SdoFAXnxPrbbkwNGblVvpggG/pzQ4
j1eQOuRgWruO+ZpJ4CT5FLZry4Pkjh8AeM/FqD4/8u6uazajVSFQT0tcZAoA
4tR+6uLRZNBDR1OnlM5c8PJtb8fFRhPXLGSTCS1VTobNBQw5tzOzaYj1f5A0
wJjh6MKtGNBDp/hdaOj5ObJNwnfcksj+1w2/c3R8a1cjEBSiQUJrlmYUKZXv
Zsv0sCgnzi8rwS9fnDaSAxYdjmzP4pZy1VVcqBAEqd1TGxuwpC/ijS+YpU9K
wugFwjQsu6dEglbd7hRf9K3Ll9iANW78CYu+cpWzBickrkTAIXAXlpikk5NV
jUJZBxKkSk6t75eSBrGv0+x760U0skcFNkS3c5/QEHvnw9JZsRoaGfggq67G
yYQZJCgZi82FXOJBpVOqzDrvrpuXxcD/qm/nzgyd9CITxSKXQg5nlgADp3u3
vILoo2eOeKaSUpdkLeZImsgsPRug/w24xh+ftpq5JJ3FiDpWAQhHjwrBqOLe
LjP1XbZNLmKyWm/F0x850HumvsPP+fL7h8cTrnHTmvYSxJdRYKbp2OKjILnn
A7frahSkFNjnKe81VkNCbQhfjLKmtq3F6MpMfBuj77OA8hMfi0VWqevje0As
NKaWcPjcIC4YjdEPNHph1mZ833K5omQQv7O/XVkd7UsREWZplNW4lBfNGTn3
DmwFlUnA0n1jWtponTJGaS1eq9UCvh2ktolApoih+TsHsGXMHVQVNF1tJBRa
ijl6NTJqQ+l4McHi50ZRKyZpZ/4ZG67lGDfKAl40G6/DmmHA6h/afHNZBHmf
jFvKQN4WQzkZpByKrJkqTkPvOlivmExpaMaiSYS1t6Dp+2l5iLai0R5quBv9
HhIY8ZZyPOz6lJi438fsqJOiRZTdIyYddXOuhbXqhPrP+bBaNDW86XxFzCfs
vWVAcxOn18lUT5mk7QJmZ0rCd6SQwp2ldOGDW+eBROQghJ5nhTTLIlUtoZIQ
bsCYaqBgxkMPGgm+W6JdG7vKieNrBla2X5S5BCYO2JxcZNThI/Fbx/rPS8V+
VfsHTKA87mrkwhNVSzT4lJcj6GM5QtaWDC6uj1oTB/282AoesuuukBNi1YdU
Sfd3J4qjaVPmrI0yHdBWGmWRgLc0Ozm5cLtiIgGlZduWgl0V5C7BExfy3cgm
ND0zvpp/VzSWyQDRb/dDSNjOczU/JyyfnFQx5zySpwLn9aVN4JV0dQv2KdqU
KxwNBA/3Avm3g0RDmaOSp9L3FfbEmwA/UO9iwkVBkgY4pMk698X7dAf2F0uL
2u6O56UAp9A93gIJj2es8uYRz3j/6f6P+M3HNxM9xYjk2QeYHIW2WnzfLzMn
jpqYLedKs/fATjCTQ2O3iSwft1FG6pc03n8JQFqZRIPc1iWVCnu9auz7CSKr
ZYrdgotO8WSqMV3aucI004i5W+q2EorHOvARQQyb4DfpWbyEEujk33GdkB4f
9DNQrdrLQVt4vvNZpET9HTFS1NctfpK8aIvhJOXYQkGQQsm5awvgmtfoFDYw
kpf2MvxKkCxGYujm4hdQJ41I4ScmFQiAPiI65L2Y5iEYGy0WfQozKBwgX9Rg
j8TbnL8ZyDo3TgZyN7UzEJOvP4mCVgCjs3pjTNbqTydY9pONQCMQrXDRx3sa
1sEbQ2YYmKvym5pToK89n1G/zfyGglhKw+zxZkqhk7aFO/VAl3BrwX3bUlXL
kL5e6QUCxDmWCbmOqpenHENrO99Pgkw2Rb/A3G0FaTCbfrEggeWaMVeDV4vo
8QVAfFIJyVtbJuDOXyRj+WaQOJSEsy81W+84Uc3xvnnsGeaCnccxVpAjy8er
Zoifr1oQrBz88MkenzbOId6j1s3KezovKNE2j+YVWpzfnhSOl2XvLxp8lWsU
ZjDmUpzDF6ii55QUmfywJ6Uu7TE/6HFffVcxIkN4LAZy8F9yVFQKlXLqordX
jziK+KfeLYFhCgVYmPFHg04V2eJsdufQBMCQfp9NOKEdUlk/eirWTPubdklI
Ez2dRrkTKYQXRknbyRhohF7Bu1+tR4yjSJUcCwJlSXOHYNFf/i84nm5DFq6n
ec+MexaZf7l04tZRuUP6bkXSuNRJJpG92RW6HZ5Km6BbZzCdp3EEptKnk4vC
7tdaEQubb2XiqvPS+7ILWRkGYbX5bHL7j4+g5qV6Yxou6lJTUy+u3XqNhp+/
JxzIzbIj44gV1RMRY7EW3OoBNql8uDlt7kuzlpW8zReG75dLQIHw/+PSsOS6
BxWXlkvinxN56wbEcn0DibK+0HV/IIOlVgZETa+PV84CzMe9l5TsYAXdI4kP
QlxF4xXlii8UMXYz5cbC+iGcYwFQFxtHxAyVLS91T0UyRwhhFdkJrqUzkERc
7e0AWNVw4o+6T7FFNaESnoPeYkMOy7TRplqv51ShLyXW3gkJZIeOk1kKuVip
p5feRNXWXUEsGmXOnkQ5DpnGM9r74eRl2PDsNjmwk/KEezxLZ4AuezwqwLz5
6wqKVmNR4wYfwEE50gZq/xHTGcRccBUk2aRAV49b6ie64Wj5v/NB8owQ8mlf
oKHfwalfFcEGsjbUBf9ePSvke9jvuGhyn3qlv+gA8XJCbowAyEHWvfcmkwjn
EZP7eh64+yerB989k0Qnb2gmy/MOJLUJKrSgvV+zPorc9v4QO7jL/KdeEYgE
pFJ/KiSHPo9aMtBMHaGzlz14PeJfeZP4Cix2PgUOqroKZyC+jhlWy+5BLZtN
9Ck+BGGribbmYY3LXQZLmNJu/00HnyC3TOSS+NlGjCilI7fybMwR0crX3fat
6H6d89RA1VL+n2HzfBf1rB38rnqpBgUt98EJacO53/G712sY+nzjp6h+SsFi
Z4YEl9phHYiD1gUTgLHL8KIvaaCBG3ycMTL+3HizUFH+ISZrA4/OyOUl240r
GROpe73XJKKWoUhfRmBl8nqPWMkyJX2RJ9Y9Y2TPFef0FWDB7q/fpWKd3m9S
s1uis/qYiRW9zS5ztCc8bEOXMZN9q3JmX3Z8MLTe4J4PuvoYedyo69H7FBr+
vLJwk6E+ZXWVxHc96zTJzMfrVuZkrmGQ4YI4Be2qDUtxfOA4EbTSjXQ8uKcY
HSBiemWghW8LU/evBATPdwfJLp56V73oD9pbToXSmg92Q6jeGFnroCE7i+p/
sqKLBLgJOnbLJLG9yoWDAaFQkfmJKDfOA/oIMBLTFyERPIlqfF41UdFdLcqS
dD9P6ePq3zMKnhYRiFeX/hZ0qn0sI6cqC189f+ljSvtCIQurZx2i88iyeuEt
qw5wlTSYjDhJvQsQXgUQ8JbpJXy8pL1tWzsiO67Lzbr5xwMLdcFuWT7+Kc7s
82at88GH0TaK4O3aueldCf+PKt3xWMGeKjWRcnngG6g0iglaB0aR0qzGHpJG
S1NerWzTNF4B8DIZ+a2Mt1NKbxhNpwDygHyVkqkjscMMGPN9/O7kjifkqQ0t
vVQs2tI5DZ5cCNuMPxDY7V7LjyfhZuIAY3jXHtpDLStQ4w3C2Psa3JR/SSqh
lxPbn2qIp7jupecHl/PJbCrTnZdYwLNzRupGfjHk8Vl6vR1IQZmRLjoVaafY
vlbcKsmAEB4/aVdvS2+65InligU0fiN7QZRv0gYRbC5mPJcikz53ienraeBJ
5bqlmoUwT7vcws1JN5bBMDr0JVouHC4yvWFysmG7rR+2jETb0yhs49JdaLG0
1c7xw5gtSEs9NB1u0qdsoe+3og9R9XydOmFnRZRtpp2T3GgbzglkZZmpkc/9
/Z2/dr0k+l2ngJZ3Q7W3C+kWkZiVMy+j1MBcSFxBwxKXsPxgqWUvEdhSSnmb
e50x9iOAiNjWNpYwU20w6UzkWtq9oZ1scC2d9ELuPJK/pPxF/7bjlQqchHsv
Qx2j4Aq0H/0J4OJxkFqgzyECO20yA9yBDfObhcgdOAVYQaJDBiV9TNHlLWPj
hqGPIWmeBU5aCllAjblFA7zHB/MW6ON63sN7YAD2KtI7JiitWMhBWN4Zxb9O
dcA0eLCYj+O5B0FKCkzO9DTR25MBu+C7fqa2b+B8WIeev2GqbaTN3o+62NhQ
MVSDSP+dSOhBUVQUtQzKFcqzh/sDK5MBZ5jfHW/mIehVbOh9zzFxYhvUkIet
zVyfKD+uN+MWvaC8Su3sv/V/vhCvCsiEJPeQKR8/8OAjM1aDl2IlaEMu+Ne9
uPPpvpBE3LVIi3STGsCgXTp9EudOSyvSPMfMK5coSJfrPGkKdUgu6HoVAr8T
w8R10zuPoys/crlrQtl3KGKDvzrPqzhiy3zCLHQ1pDEeZUME2gCs9pi8gPGs
SAHZUe4nB/MnDIrOTL/yDnC/cEtHY9QL7Tm2+dMkSZdnoQP6ynASTyILf2a+
gkbT3GgHcsGRrVloyD2UNI2JuhEL3S0eYkvKGQNO4vVWbM6d8x+Q2oNHdqd1
hB75JUg02Zd7XjjAiWMt50epMbqkpzeetg0bKdmWIihGkCIGdJ2YMc19Uyh7
gin7CwO2l8ceydLsdCFeotI+bENxDXb06wltZtBriIAZRfuys72CfN8bnMdA
fJdfnfzgXJjCZS5puFnH4iZkG5V7DjKVM0Lj5A1qbRluqz7nPVhs+zc3X3KV
dx76lkv/1Q9qbjZwM6dvWx4Yn0HuNfnHwlkHdzV/3hNtx8x+L+H/75Y1H3N5
U48j4EBtw0pIFvWYA4aKva6EKZW6PkKYm7iwyouGFG5EAxOtOGO0hUakgozt
9g+Uyg1N2jWuZk8+1AXqWTHxBlj2AncadxXM8M6IouHMg222UUrskiZna7Zz
jMi6zjHFVr5Hi1U0F8SIs5G3SnfSvIUkm+J/tMDMKGqwb1VOBZISdUnek6+C
1Gx2Uu5qwQUrMDCm9M8KwyRNioe6MvPn8s/TS6zjskoRDz2Y06yqr16q0/I7
udUz5nBTevcaA8FgCB4rsWJjx8AGSNBQkJjyKX+m6teN4To8aT8oHzVUXdUA
JoVlISaVMR+93H2r5BCyX4xjkQcbpsQsBl49cWLXzCIMMFZZACMRt+vS9Vri
QwKKxWeszOkhkM39dZJkWCXlJW/z23oVOJbAynSIA0aLH3vy2XVZ5jzOODz4
AfretYNK9WnFTCl9iHIq452SOnLlLzYl4LEMEXh8w9+3sfxYGeIuTIxj2Q2t
eb5Y4nnt0KWTdgZvtLodwOrixCvh6zXGRS5covtfgJWx0d12NlaWAESUArC+
/u3SsJG48r5zrh2aPd95ACWkSaXAF/LdPrJCjcvZVUlKAQ0nrniaPgLPzofO
gQn2oAAqrKK2grZvIohvgaf2p/Pu/97fnEzgeuxEngWWoxZxOJ9BElVIeU9+
hxHKzI54k7GgtLanGmz12wbwuT6uO+AXW9g2fPQMp7CxOZd68b9VOxh9mOOS
nDG4hGzhwW6tMJznC2cpQgOMpZCp7LIs6uPYPEuky7WCrGo9mqlLoMLiqNSS
LBfvHP95UA49FJfIrgvH70bOBP3qGXCqhpXXKRfrA1/FqpdTdFwQZjhEiJ1/
W5UWkwXwo+wOa6jscaeI5krzK9dX25JLlL4PeBQiJg5bU5VecmThX/moMtyA
duwPrJRU446GRR2cZ73ANSGxm07oidMMYJZW+Exd9J3p2oU2cfrNEYUUFiME
rh+Yy0OQHJfGyDea9AzQ74q++MUOY6uFaGvpfnDnld2aAs53hjuEF9GAQLGy
pnjHlBe91Fy8E1BBFG2cIagSTMhCSpx3aZ1GRv0ABEjVqAMObuo8wN/EIosz
4vUC9dA250qk4etKfMoT9XudX0g0ou12CVFvJEYmWeWOd8q7UroffhDclE37
YVCuC0fEC/y3rKke1gDtcpYwgdMZjGeEYJ+CVh3S4v/a5m/bDe1s74Q6PF9L
Zci+GthcpvfGyXX+ilB9PAji3AQaXPU94muXr7MO+51v8CzbISGxFRXYxyM9
+nyyrQZYYLJl0bD2sOGNXdpQR4JoXcM4408++1EJ8a973bmIphaJoexVeheE
mlmETqh6Wl8amYOuCpIbtCx6qmWpJrOEHPcIwOckGra9k0QIQepPmZnRDAPc
lYI4SvIvgtP1ZiXdlH+norGXi8yzFcaSBo3gpf0vXggRilBXMFLJJNgieTpD
O+sJV3/9l7QPqsOVwVu6CiU3rrVICjRiWHle4PzOScEDw7GpdQ2Ruof9vMk1
Z+QFQXLbJwhGhgBoFxggkRGHzgabNvkz4sFoxhZrRnwHLyTcLDWRTKOSTopR
EGvFZ1k8UmZVmBxXWDhqSLCniLdM76JdfzGQvOndvGvbzymKaKeuvPF9Q+Hj
ZRhopLXvnCXTvCyB61NcIMPrqqqPRs7UfWqjzgXKty/OzmQAKOxDa52521B8
DMoOkx0GjZD9YevCpnQ9ME+xrQm1ABzPsJFV4USTRwCqxp7Ro8lReqqJBIkU
rKiJm2u24GJWfMWSE/XUFk/LNdMvLCbkN424nP+BctsPoB8y3ERHzyc69oJh
qTfuwxcoEUyGm6H7A5w0tb2J2J2LtKAbKwBdIeyUIv5uBQ/x8Pa9wo32eaNp
IET3dzvGUZvkSOKLvA+4X73Pp+/N92go3Kg3zV9p/MBfQcKNoCj3YIwban5W
8Im9fBz8MaHvuV0BJ54/nwf9qiqI9xx5iy5PFhgFSzWY0ya1J3R849p0LC29
fZwchBNSmEjsMT2GP/sqWjUsJ1xkoAO72mMmDOvjNVVkOXNOYVOcz91ZyRoL
Q7FBSWSVW/xlefZS/Rlx9+n2ddiW7S6l0vOaI9JAb2Rlhr/s/HQpCq3Zkjao
vMzHQu/dXJAQKoWpUrnb6xkbWH8ayMeT8N9ZZxAihIsP8tby094iSytPFEXE
5rfAt7+w2+F6QMDmSebmSYIQQkaM6yP+bv014Vu/EUBTLU1kxf03GROEHZb9
29MDtS0MxQm0b/XJhPMPLjjF2BZB7ZBNYmzsmCWZYN6LpNODFPaOpSmqKsKC
M3/Lj6s6wknXR6TVywxU/wOVRKAgz7/H7pA5nNYwlwsYnRFQTz8JN6m1gRHR
Snf1EwEKRF5j9tH6Uj0w+w/um6zBXC3oyTPAtzjgJ+N3SHN5HmQHRS+F/qDg
s/ugHFExsj/U/1sucJOXQLf55GsnEi2QuRyWP0LRV5cLgGVIX6PPZvzAm23z
sNC+8q4xHEpMOy0zoNeTdo4XN5vI6xoYIukAgvMA+vtnKs6J/APN6BmUDUYU
FSOL99IbQXgDqij6LmuFMtuoj2DJMNPwG6sRvfpw7R7bNAy2ceYf0dHbi+vl
/8tj0Fm6uEdOQCQXupeDva7Ox+CmIPaE953zUgXUpNWIfOaKObqeaVD4qen+
66+o2KvXVsblZr3rs5LGCkdxczxbA6K3klaFQnx1hZTR5ogx6+fikq+ekg9T
dOpjWcaWzA6+aw95DTAOk2r5n2Of5ru+mhnkZBaLlHZV0rhe98SjcELjNUtJ
apwq8UQIGgMzlqIdZEFbx0jRT/gwyDMAU9rAXsHu3sDjgsmyCz9jk84FkvsS
7rHkhWY4SFi/X1/NQleHNAlpiVZZR7fuxKfOSZpmq06iZPiMY+x4vZmZKK+j
EXjcdgKRln0lZv/iuCCx0lqUCkgQHjm3l6Spg6yPQIwxXtN2y3b7iFynDefK
BOQmP1gS74X5/AVA0g86CHVRRHhe/t/KMS6BljJgV4aWZRisqMjWlYQvw4Vg
Kjuev4dibg8W0yWw41n8KMCmKWShOp6e8GlKgySxqlJOqhLZ+EmbgbKFkKzw
s/CRRWCICqlMVisMrnxm9M3z91AYZHipNyUALUJC2fDxJGYX8yOqFoFeeeuC
Bn8iCuPIiktCSgW8FG+F374ijI9FI550f7KishNuw4BEpcexLpAyE171HgZU
YWyHlOM3jpvlwYmxz1RkCOWcPMpDgFCNsPN7SGS/3z9LZPN+HlLLGvSfo3Rs
w4NhsOmgW4oCEsfz1uY+tjpQcbeNLGYkQCfDkbOggjVxU5pCQzTpF3CURB0+
aIywAwg10zta5U2RUDAErGKfcv9aobEazNFY7tEfRNCIGDDuJtFf8l122py2
pjgHtUi79/YChuK29v6izqHMMpSRPQdRSGv9n9nb179opznQCPSYsSdOSU+3
UYS6PZqiGmly0W+FL2mNkqS5vEHy+Z3tV/hrYauaF8BZNyPIksBwd1G7UiR1
ULWZ+//ByZH/LuYYMpb1+QU7xDrHoCCwf7nSaJI8Y2U0IYipJxgbAK4BPGtN
HU9d73fC7hrS94mBQma5DlAnWuG0W8cJYuPhksqXf1WXZWslxl8kC+vuvdAA
W1clO4i327L9HjAXY6nArKQZAPHfQzUleEaqi7ObF6E0FJzFUcaC8LEcy2Fu
k6hQI2vknn4lvza3NKUp0vmJ/4MHTB0SM3hqT/AtjDGMDCDCPa68cdxgALSm
pDQX5R7KrlwvMi7bSQMAF/NxiHQlQ53CgMuMjQeTjpNYOMfLIQL3Xe8xUR4l
FspW5oY2gbOsUFI9tY2b1sitVnwP8wUZ0LtP4UFF7d6cO5G4JJh/HQHruadZ
HET1vfmIkSiScEhi3oHKBYczMiDfxLAkRjQDhx1kFQzPTK18uVC2QHkym9cU
jQEZY1Z91M9F54Bv/B7fzSss7ZJk0N3G80FSfpxh5+VBb9LD2Rd7gLvmtzRh
/iUMK8sghH29efQA6J8ucViaODvR/e51+Umsrz+x4/tGeDeSyPy3AhrbN5iS
QdIEn1/+jaaOPyleGusfi/IRvgULs2/h6ogo6/5jW4ivGe6/e93MNgz/2TRo
+GuhbWTvr0yZuOU8ujSSYaokFdEEFQSbgRFiGlkGqS0fkxAUzxjPFZOFtLXc
DZsHvfvlNmY/9V5hCIvZqnKHbADf10SYS8wwd208XUXoGdclnxKNNlAwjVUN
4y+wz3ZT1oXOZAG8RwfAhdsuFDA4MWPFg0TVwqlXEi/MScChIc05CTa0JnQK
naVWPYRgQ6tVvJ5Q3X1gKGJCo4h0SIeLcfOL19o41Nb8656h9wiTBXAPgDfo
DaUwTePBbWYaQedTXQuSJFczVL69JX1HhzMTQs8AUlSLVKk4Iz/dDF1z1B17
96VYVNiNREC2HaMAtkjsE44r2qBdswGOq2fvKex1mfW2h/U4wwuam4g4RdUk
TG9Uyy6cX9dZB3urvHPlCvY0pE3Wlpmq93wa/xLu2oozN6MwQs2x5mwSmnvk
sTwhdSUl/EJJTQHAC+qm5Lv+j3xuXimKTpgYsBAYDMAzVFoK4dXr9Jsf2czI
+BvzsrGwQNZuvORoXsLFDdWuJ24WFGQOvMBVtZavnfC+V0Zccqj3V89RI6a9
l9VFxl8oHFaCiN4/wOmwNIrInZLvXpWoGXD1NLjZ0minc7wE9NHVFQMJm1r5
n023zc+byt3R6W0ObZharp2a8UQZcYUr2WvTdtjPQV9wwNzak0/pVljqppqW
7HDoaSlHTZLVt9bT8yQX/x4lAnFsvgCAMPHmg0albgjCvdjrPC/XSmVcPAYY
qMy/nw4KGPFqWRSdafznF8Cfk7Nw78uy+ipB5OzCSZ2tiUVP1TBPJKiMbHt3
Gdo1qa2DmPfN0ur2x+nAOT06+1cyDdAPobwJt3ZHC6/n1PZKaxYKhCAYemTG
vMEeJW+p9Cb73pvikHVyzL7Ee0RovEnjXGpS3cW1ZS/CjhObUuvAs8hnm1LE
8AK57P3gurH8RQp7gnalCJyxYMvBAIHYFnID9aIVvy6QW5L3KgZot/O9RNfX
l0uZtw7/4tyy9IQUZ36RZXkUNXybnH/z2AZRAfIB5WIrA+PoipTpYfCL92Pm
5o7xrRPADdZQGVx58yG5FD3NF3N0fmfsk3WYHPLGVfZ4KC1sxkEwJNB2mvgm
FUsfvJeCuCMva9msolvXHtpiJtcMrRrq+ZvwSDUY1qT/XkEPFTLRbBeyUJBR
FYsO+ztekBTC/DZdfSUafuBbYQ2P11EtyBTHTf+gS0YsLNcAZtjY5TZtzk1b
1YraYQOVUgp9YUX/9t76zmjEEwf/e5OzkFLW1oyjmQaIkOWqV7ZGf0uqRnUM
JZoYXKAO22dJ53XF6ymr+DTF4ATHGUdpCNLS8rDvBN01EYG/g8MuRHdHCtdd
rQyyxaxdLoDTx55jZaLfEvshATrBOf4Iy04IeeRjV/1vKR7UlAO2k6zrnunW
g9ELNfc7x3h5hn5GBGG8CfhINwml23FB+L1xpacF8QwKcBlCw54ucQiiHoT5
Is0FLaVy2doCVhiLywilyxQ5/kYvD8dVvn9rLM2afbxEPWWAUs0rw9PiMb23
CNvufveaO8AMjeUbVKxLCiaAFATfNFYKhMRTCBPGX0WsT6yg+rxT5Q5tLSWw
9vdldh2zFN2qwQH9jIFzZXk5zpCJ5xzLQIvbQsB3k60etjgiAxlJcunpf5BH
WdkLgvmnGiQToQrgTjQP9bC3SMIkqYj76jT4tYOXZu//cA4anYf4pH34JAFr
PKGnvnK7pJKiKXX/gsE1LmKlQHiAU24npkiHgYWHn5UMr3Uw4H72GIh2Wr+r
4Qnz5V52+UcmSATP0p943jfCFR2VR4/n6jY1JPzaJttH6t0RGF/BbPqHP4Xb
1964T37KIUYzV/bFxuaKvX0ptM+Umn/COUoICWj0JlgVI0L66ZcAk0i8374F
XUipakMi7QCuFAJa0rELDQyG8CashxDSdwIZm+jgHZUcG7bcMZJtYezGAafH
U8p4U48xQqmbwfvp51EGvkbXfouIsRFhxKoadnyfM4JFmiMSf10uI/bhlkun
2HheCyXNZ/EQUJJQmI5AeUW73p593G14EcBFjkRlUSoum8j1whalyustg84J
RpRDc1ft79YPs8IU1liTQHWDzZsl4En3YRroFsCoaXUTI1Ogs9YjWJE78dAo
mATeSvYcFGbiciGGyaaiMssn83gQ2cOoaI3Z12Y0xtpw3L4+xwTmo35xHleG
DCJYcAxac64VURLuZ5Adm+Bruz5xCt+jFWBb3ZqH70CVlVjDfgJashF0f0Yd
ypwKj8L1/boV6ATrZcFuoDOutldXJm8f4MFlxfZTk31IFbibxBYtWBUTvisJ
wFkYzYHIPo0ddCPJ/1BuRWcTs7fs3QQ+Zw39VmwPHZb96zucXP54zO3/jzS+
7ej9QIaFaGTeYZ+yNM7exxtRrvzEzxkwZnm0gwkQMh8t0k0M07jNZje6LFig
+XswWbqhHc068fjVBMg3ch7bOvOOCrWzN+H7LQ9gblqTCnFjFTf1lqVVKbFd
aOxNeB7ycsmPjiIAiicTW2qEIlovOjVBrzD+F5tOpnWzYRZJ4wHTRi/cv9P2
CiNzeqU0MEckKOPpxJTCB+zxyHwYWXKAx/HgNK1hcIV68m0oeJtbC1/pCjt2
0z3MoIdqLOWiRfbG8/CWhAtzq1qNGgxnB9/5aUOHwI3N+gBXh60e/sBdpxkW
gw7HzlMARpAC8f6xzNDPmD3m6qjljh5vxPLCpxRyk/q9oox2ZZmwCBSbEDCr
Lfl/R39UWACDDololHwoScpKGDurVH3j4hVa+N0wcHUC5Ge4eGcg9jH+ERsR
LUUIlROd0fRpEZdflxYvGvJboqS+yx1XsuE/qdnXA6W2Yqacq9RSrFvNgeVB
+E/Ex6SCEzMPlZQimfZrhrPkK/VJaMEDEnfgpkzF0Zwndrie0KDWSRexku0+
5cPyQZfhDWippwdK69DjY7yJUbntosuxWmLOWWsy7hkJGdqxAQi2xpr35SQx
TP4ov7GU7HEhVMsgaE45SUZka43Uc7g/NymdGDczNfFLX9RhPZUWh3V9ntpc
ieFe9CsdruWRkox63bv2O0oDeaJ3WTD4ItxvVpwYxaV1cTk5XkZOgmpz5d3+
zNUzuYUGJmz3QdyiZlcgZzv1mVwR6ld33U0STFbQEbGMQT7z0kg6kMuaCLun
cMN0G1ylxbI5esPVi79FMaIrZENh/59R3sGJZKF0TuNl85ItM1Yf+VGEsyhU
hKYiNLQqX6TmdFHmQzdvMIVAtQtbuvYrACdp/f8s5l0GgSqJuNtEkGlHROI0
NtvNVBwnT7Id0mqbvOCbQq7pL2z09R7OdoZB2p4T2rFsqFkFigJpP4tQytFI
xNhrMnyFYh522JFlm/uEYv0aVFoK/zSAhR/ikzoBLJ1PMbAiG4+DNufN1nd7
eAjIV6LrWbYpSFzmaheWVU4JfoQdxn0NdCqQdvOQMN54XHthKE+WkpeVa+1/
t7POPbRA7ovR+DmIP1yBkfyVUoHIP/PkOAlOtO8sVOhFoJQoxPqtjVcP43nt
xKAL7TegmJAAA7Q6RpUDMTZ5D/kif/EKAKw61XJfoUK4pLFxPRXw4DPK8Xp3
9fSdvi85wkQ3EaiK09nG2/bW0exyv5BlaPOA8N00pXXo0WEQilzKFqxo4gTj
ygnUhNGXaXJMGH3XAVXKhUPZ7YhMeUX4HZ1/4ms7zwoGefNY9rdG/YJoPRLW
aeZH+KjoD65YHIYC7wN8jPPjZp6PyQqSMn1K2WbHRt9fjNRRTjVJOtr+xKt/
1bj2lmJaPG00fXjZ55VgrOatdonnhb1ZuC1QnLijro+DxpoHeeKguYHvqesz
YmKav74ftnrULbXkPSUxQ/5/rWja6Lt3BFHcfIDkgYzThF2ga8qRFqlzwo97
Jf5oqLUKj/HGxWr/DVhBFWo72QGjCdK3I+c+4HJxdqXrb8e9UZqrb9FRPGAc
rufoaAb7aIV3F4vz9//Xtm+HRondGF6cekwAj5cgJj88CxdQxYwhbMFSjR4Q
g3ObYf3Z5qCj3Yd7npHoSwXs/Fhaq/p4pdOQ4DY6MgjDcDzGgoO4F3oYXSFE
0uAq0jNBlB+fHH74MTfJaPy2BkBvdJ6EAP5cfa4K5WIjrilDh3+A0L8glS+W
LLzTuGJcwcS5hHcmgx4+p1T83+RM8s40ZsEft34dTWrehi0vBlFHZJvDM0c7
VJxjd0yrxbDiQB9emgyGACTuqE7h1ZACuXP7+uyNodnburNFlNfcsKpZdynD
eWypwhlLO7IkeOpdfc8gKVXKeCT4quAP6IFsB1b636Gf77DMfF3BviUqVKkr
ZEAP5L+5fvklPVqR5EzrJK46gomWkuUwdlO6X4e3fjS7V0KEYUVYsVQbnpZq
a2zZLejkxm5mzlIunQrDbFo03HAWPI8fX45Ny/w9q9u8Pn00dEPhK6sHR2fr
ZJRKUCYegjctyAteUBSdrpE7I4RQnugjfkL68FdcDPQwhjVbl21Sw7RqELvv
rv4KHCCEw6piuwVSd73/KchbB8pN0tmgH7X+wsQRfpZWY/m7FaKgfHCPETsQ
U/67AqYSvkSdXrOhc/GN7YOp6gwBJhmsCmzlzhv/SWcPEqboxqihG4rbq0yf
2YIijwZRYzf/Vs2BP0I+oNU59Ba3rdhWTCysX47FGq00fNIpASFJDDAt4ZzD
e0B/zy5i9HDePscUuxBfQH5Orb8Wq9dgSSAXPo+tBi8q82yLhnxYu2P5JjpU
VKfAgtmIXobv5bwFuTgJvkXTPFPvkSC5Gv/x0W0gXWbBBSNdfT2epjcjxaWM
ZSYflo6ItkezNP5mlOqIWL9qPaZ+lWGw1e4TYBOeMVmrijg58iFXyZqhVUUS
xbek3il/gCtUf1eELTBZTwknP0s+5P7/JfKpVw4xNETT3trODGi7eCCpxaNz
isfr2/SOi4nwynqDzQ0pf508SV7Id+JBMncwYu2fKWCkc6bf2kUWWEip8ci1
RZjVxXYOsk8aklVvXDw+ULNh9l6q/4AabGoNXj+kdxWLzNkYzfRBkxYaFof+
jw88k9Ki6kvaEFAcAvI+xW4nu7TlnZx7Y3a2RMrwBCxl1T7X4TExA86tQ5qj
Dh6NoR316sfkzpoNRwLkv5Prs5869/S2Axa/Cc2FPiOFWEu1RL2RQ1nJIrVe
8Ab3iNWHb/MRq8eFlcsZdquWivxUcQ2VzbNPP88WK8JaM/3eBMvgK/zk74gC
YAGyTPnHkl1eEmPQVTJ3EsY6eKkvzlodYiVXYrzokQPcPOghh4H5Gv4UFurI
WKO1PTOJcbcY1Z3s5FE5LfjvFVjw9ZTmYFYEZf/woFwkwL0KGH2+aXjK9Wf7
8Ic7QSPsp324tiTeaRInUs50DOuaLsEYvtRl/4xy8LNmHwGQfu3ZuTG3rZL4
FWLDQc5eXYji9x8PzuhVMMI6FoycLj4e1Z1UdFktao35aHrjL67UB9vz/Vyk
5+LRyZCKGJlhjCIkHQAVMFSfA8SfQZuWSEnc6JL70Ol1V7jNbL+YPjG7pXLd
EYt+3uSW6LYbSmxgxoTrAY24OGqogE3A0Rqy7ZSnt9Ia5+TDO+b0c8JKgPBz
o/tQeY9CqTbZMctmRs9s+ABqWUWQjz7waLhb1ZQvo85SQLgkA6TOXOi+IoJ+
s5n1Y9z8SVecLAJO2QmFqifShE4uwGOx/13h1MK7rtcXCdB33RX/Qqse/8Na
yo3lMC1IVo8FHul69kRAop4ADaBlmIvSK6TLzsIFshjncBih8B7EhaeZj91e
TmbwUhi57Y4wmwwwYrDDiF8k70Y1WI8i1RwftcYmktyAXXM7wDfEB4Cvd+0o
qQ3I9bb53k9T8L8Zv/RNazanHoJ781ZvFoFmhbAk5qzi1y2cBfpg6yMW832m
PB7RW/4Ac/1h0O3J3r57MlzGPiZqi8lh1auR+XvrKSk7Yp9/+UHE9DkEQIMj
Lyg/ubzOBaYEAqjAaHouL2t+smxg5V+/IxV3w3irjSmR+iowvT4fTmj0nrVf
EISGa1PCXXc/je17orf9wduDEa+pV/JjZ0pnMq8MMc1aY17djlz26EGWUYwN
CmNx8L8oXPl1dUulMLahKVvZWmmRwU6b4tpoh+AgCchcpm0q8HdJrZiSgwFm
oiktz6OxXDMj5Wu6+7og0wUmLsiuIcm6F9sJvkyaqRGQTLV2ePx0c+BatL/p
jGe3Kovfh8ls4QzanSFjoBn7VSVEk2JpP+VniT50mMZJA4OPe4wBQKD4rhj9
4ug3KzBfS9wB1I1yvYIyR35cfE83t9ZXIjtVcjQFBLFTPQUnJn7kLNZVdihk
oCA9n0z+WKMoCeqmS01mwrJRHZ/Ze50SR126lX3XoChuG0tjToVZUG/nntY+
DmAW2nqmrjBcvFnpmJqyX7pVnlIwS9el9M+y/IswUBre0d1zjWcNibeSaYmM
Xn3dSSvP5ey6wiHBpecE/M3kZN6TN+dhLvv6rsdKYm22/YVilHwQ6V83/RC+
Xlj1g+dLfJAMrT88SHr4vcUWVt1+gKFGrbsQZDka4P8+Wj2nI+PSeHQTl1Cs
/RIcCXz2ajbDLuEaCeMB2gVT3EwDDeION9UlLIYHU+eK2Cnxw/LHraSfYKOv
oa5HV+1HQn8hRbST3yK3JHwF+tX1rZH+7gNXbvhsL4DY37233kffh8mJOvYP
6XLYR7i0+qlaTrwy2dIzYrGVncX9NDqGIOXpEf5IBJ5FszIg2PmY3B1ZSkKv
LnJ176A/ULTsRGnFbT+y+fyjk6XB46ryG6JPcMOi59b/2WorxcDsJc7YATmD
rn98+rcjO1LQm/cU7WAg6pmCaRDf25EbCWppiA2URBu8x7tGKTKZiV9bkeE/
BBzb0CFoRMKvbgVCyieoWtKU98kAcEx1XdnToowMOoNBEYU3e/9X2/VNcPe7
P1vgOsGUGmchtDE7qB8N/CnKRtlboalEID6NNQ8nc/MsBaA30tvvJmkIBEDC
mSgl8jdUJwTrC5Ths0Oz4DJGYZvmryTeRZGl/Gl8O6XWXdsl+0A+DRp7vusS
HEOxVIQRQq0AGLwgJik/zulCWwYT3Ff9KprYcpGQ1ZGyqz8885zAxEMm57kv
M8J1cXSNaubtvf+3J1qhKqbdYbeZ8qZ9lpmmjuq1wgztgXtfDsuFB9uhCRsD
zsEXBsIFWv7lKPXbUaG9SKdUQ8qxP4N1fikZvDf8O945Q3RIXxVAbtoxKdWu
aLfl3IswB8qPdp5ECIa1upf0n4KWukaU8hgzQ6Zc1wSNyO9pm/X7jZBrQ+Ip
Xp2RjBWVt1aYpuoUnylfBhQrpr2+MMpnFY8YG9kHfoyKNpu965Xcr+kWQ3xa
B1DUsUkp4w1DNHiHH8XnqMURybQHXyW0Mt7oPc6tTm5XSWo2+iftnDYQC3O+
5LTQm7RDN0PBdgnxgbVH9CeHq1IRD3sElNyT0yGDoPIXQgnHWgOvSwISidj6
3MNQNa/5YdqTLhJp3yy+xD9X2zGbQQHLsPJ6bI7Egxc73K6hHEwy79MzUxng
rE8LUSuGJEZUqs1yv2/YEmIdYLeJZP6vuSLPnRZELM6TNbfUg1vtgfCarOJi
74qdRDTgvtGY7htWgNERyerZ1/qfnb+X/0J090E0lcT8G26Ywy+Qhhmd95Sb
f/GgYZBjMUS6Sm7zdMjGUIWnRaN+/QebpQ8yBP7I7Q/XfE+0QRVVpcRixnJe
0GsDDb3HkHMHm7kyyfrmlK6fGhcuWYbSzC7CioZ/J4FukwAd5WvLxsZ3aClE
6LPISudxvaCNPm3cmWNraLSr+UrnIfuBVoGQVLC7/BObMkRonV4GfAHvSXby
XE6NkYnw3rX4W07aM4Zb7qVuTbK50/b3VHFXMHA+M/txQeTDsOfq0PYp8l7R
amBHKP3oIOnUxFf1ox2VoSQA7nItyQoeMyWFxrhWeAIzGZaMbczt1rKuAEb6
+/xKMUJJrOGixLpFIwdGrJ/JjypBHOEtuCwIppN/7iEe+uwg3LCUPUi8UDZM
Seaj8IdwS2PcviMAbjMoCFVlRdqGVTCzjRxyCct/fWvBtWMQET76JuWT1Vl/
31R01XAhJs84eG/SxANduNJIBToAwRFXq44YAMSf2PlgeIADLPxDgUL7eu68
E5Y77cOF67uZUFm37NR9SWF91d0Rj3N+0ix31alEgR4g2oATr5MurPtBhzWn
OhEm572qmab95bfCQwnhGFOWY2P4eFm3yyZlI4Sq7myif14fJnUfqrtG2xOR
WlDjCuLbH02zQ3DLp+2Ccxz300R9Fc3uhlv7/UctN1NUjYBUezLIpFMzAPRO
1j7frll8EONagNoGQEA+Bvfs7hJz3azCz3lGZUyP7pywvzQgF5eCncmkRXbr
HvCtXadMim1/RABIShBoBk89AF5J/8SlUS39i9WaX4JNSg8+hJ0agwRzP8Cx
VwudY14ZyH0k4i7yJzrW343Db7IyaEFsr10e01KPhP8aqAPlKjwwWoRl8BFg
FUFSLk07LfkBz++jpOcOjJ7fpOzt9Xec4dUg+iRrI43oJ6PU9n9bLLe33DxW
NHPecuKM6ZyMbiwevKNdWTJjZwbhGRdcgGzNKVbWAemL3F0ljGakJ4X8mXaa
IeItA2I7jU1Kd6fCjRfLErDuhiQIj1Gd8jkFtvocsZtkwTI1yyuzmlWdtaaL
CXLnncLc3l9dkN8qLoc1ahblN8doVETjEktmyE9FWCUPqJCDnHYGMHYcVvgy
mU/uzxbu3Rjtqr+XF7CWPduZ3SnQo+RcJuvVxLqx2KIY4Yk7Fd8U8uhX+I7n
Aej3NxTYDI71450qcr8od6N1hR84/ar+zLIVzYa/B3/jvHAfHBK/G+C71dXt
OqA1jsAmiLF9TqZ04hdYrVGbCbIl9nbuA4fAfYqdZITv2Rbn8Vb9FLWDLM/i
d+fKnC2EvdIpMEXUX2oqB78P7/ADCD4kuK9/pj0e66rAKYamnPta8eIDfGUp
5KAKCyZnEugaAtqC4soqyJciycn6W4Z/7/2MiEOwjn4yFIRjEhhD0nTDfTHT
EBAoVh5EHmGZZhmBmKWxyl4zrN+WkcUYOV9aSRpCYm/YCjNFgsbtkh60f6Ys
9ZoC+ESaRJjbvxZxBsD0QEK6gnxVXpoDXIS0uQtRxXILuIJ8kK05NW1M9Kqk
FUW7SsR9dznPzt1cwmmHFPEGG/wD9R4xWLvuibPLwIOKgQc73O1OA3cZ5ot/
rd7O2qYmPBmBlXpFArLm0M/CVt6s/JZd+NuqVr0idSdIEDWUudCl1oaMN8Ep
nULIm8A4U4guirZwDG9lOVupRg3R5dgBAIWlM5PFeEKiEirSqvPUVqHSkh2D
RLMMdPXp5OuEiaa4KHqgdYWRdzvlG1w0Cu88rqFg4Xk/2BHirAF/mw1+1xLl
qmalExiaxrTwdgvhokDMrCz5/dgDtP/tFXT0/RFv60vftidX7piuHH9rE8ZE
izZvm4VzZs0Q7W489lltTgHL4NusdQwcsFJ/Q0wIKEfbVag0U97rujnGA8UE
zPMQrKAOtTlP5YznXoUEq3l+x4Ufzl/8aUgjZErTyX/jyy1iiBvDBsSaGe9E
qX3X/8kdjL2i1ozTQBpqXw7/tXbJwJoB571GQlQCKWHxnyqDdhO0VXtWRoK0
F4PxH5MKoeuo0Gw0Gim0Kh/Ig1qFTGziR1Q0ZgP79xJRLuzhU4VI+fbPFPCu
Mu0v/fRqQEIQHsQuie7zQ9NIJCoaKFVF/4vqILV4nu5TUlCQOcCdgVtO4ZSw
o1gz7RS9NRnllZgadwMsTPKRJiwV0xzEiSxohAMkDwcgQDTbBkzLwSLpVK+6
dkPwgx4BU14/vtI60DItzD5wbOqE49nLKsVhXi9/BVnWw92p/t3GdmmJDLnP
pNjerksdskaFWqL3AUozwHjClfEddwTfegI9FHHK1W2LeZM1URt1w3PghGHJ
IBkT7IIllyZARQ/cK50537SD0AcBTAqjPjQ5aXdEg2CZERl2fwA8DGW3PgBp
nHyMv8OaA+z+sf8JxvF1FtQyiyFLA/QUBnP+lUeDiLUe05ks82bgHV+Sc/Xb
rhtihtit3mmCQCUt5nYouDau5BEFg9sCTHVL/Y6QGKVbWY4RGa3s2eqUWPQk
9him2IJFSBlrnJB/iSM8FsT5BlicQxpDQRGh4xzSiMvhLUhib1YdgMZHBC8M
8GdB0KYBVZcIGKLVz9+oh9PCIlz3SSoevU7Y1/m2e5A1aDB+3pK2fCrBzZ8m
/sRSlVObVc7POImXnbCa7UiCEcEDlslCDeSS4rkckk2KJqVdTKKrAiWD+Kpt
x1WAq8FGw39tOUx08ifNTK2knUA8dzjFxC5FTbMuEWIVZOD72ZaYZl5jRwk9
2tTPzuy9r68PTjtFPgEhTKzZosnww6Fkr5rwURg21u6OHBfd6csSHXXzaXX6
cfNvDTtdde5zWoLM98s3oL5xyUZzkrZmZcfY821PRxs1+PudW+Rt7cwgS+n5
lt/kOguPW58EZk1WzLggVmGcbHIh7V11P2zBjIGox9d/EagjnfPe9QUAAoc6
gLsjgNGHi+QVbGOh2YtBi0jDwrNGVTwj3PVDgDTZGBTZMZiPOO0HrL4PAoLR
njKg2gJYA1623w4Kxyvcl+pp3EkzInOKqIbh2plnVKVGDkGba65+4SZncE8T
U+aebovPe591WD6FWZGq4Nh3LbHAQNBnicZsHWLqFouWvmcA043PQtf7niun
rEZS+M7gouhuywspsYkTccK9H2cvJa7iLIwBaJS2kt0N2tZy1+uO19GRMX8u
sh2OMH1a7+t48vrYT/p7W4GqumtYLaY7A9wBygd+ip7HFUjRCIz03EPhlPHs
dHGDnKAA0Eqbo9S6yWucXaGVM2Hk9cvF2Y1KTbJlJpIGpgIHLPwp7kg30aey
YrO8jlwUeHFl34ZRjT16CoHJ5UG0WTrWKcYG0qVN2lL8XcnEFHQ/4NzBiafz
tyK5kRX+KuivxhBeyVeF2xI+12mK9JjLTq4aJVDnTDV8KuDZ7GDKKlaOV8eO
hSCj6qfJRwU/HhfXSHzRQpNflZt9pBQlKr2uL1VQzClOoHkh3thf+jABvpk6
Y4LSJx7EC0S+cnazJYysGNX3E6IyVIc7FQry/2FmwfQIiO4hmf4aMyXLbfKB
aQNuiYR6hImU5A/JzxvbvCupqeVtLFx1dcM1NBVG7v2Muqbs1MIZVRc7KE6S
ImU8em13YbXv9U0Ob8xXa8RFmTKqg19tgnVgwRYzfUI1bP62RNS1eqxZ462r
s9iTuRIPCojs2GWMsrQ1v7o+x6FZdQnybsfsKIJk+bJO+eU3+GIYaaAVeX+l
gNWLkQ5kIUwICbDNLlrqNnHX9pIcsmUFb5A45j6ImRyCodXr0ioxF3m+pM1S
sT7QL5RWRXkB5MZ4aDM2L2E4esu5wALQuYx+qMKecU3RRD+i+Zsax1qk7HDF
fK5hbIoa4q992eIuVtUN1RwYgbJJpR0YtO2FqNJZCWYgjqo8N0kq1ReFbIe7
3fw2azIZdEEg8QCcra2Yj2Sld/JOSAzctkDO/3kEq7ao65L9u8iA6k2QJF2+
+4OdtmH0ZRCit5X7IYmYX/sQ8+YZtbwncNECFZyQo9JJfJuimgDEEeCiuLYq
jPoTLK3RnZ1wBNw5+CBA6k90ytPmhppvNtSXeUKfsDR6/cAZ3lwJnwmygllo
+yNg+4Ris5lbVFPpv5t5+g8MyudfmFNAKOf9mkj7J1wQOrnPRfijoHYqpyQi
NQDfwoUN3R41rdzxlHFY6okw7sPsenCJiuERxzvfqYuUJZSL7sn81qbn4DXg
kSsU/r/lt+B7oL5u/PEEh7Ef0iaIcVf18b1XEmQ/fWMFwFGIjkBqudyxOHHC
G5LOWNok64uRqcTGPvKNrSnnpASlMSPnfLk+F2sNyM1DDMlebTjAfiDrvqOW
OhFEldUkHqkyeqoqCkHyNicCkn53pB3+7CNWgSFgT8sojOMOgR34peMjbQU6
RdArEfzM+MrtZgSHuz+5cebBgn6lfV6xTvaC2kfEqxJHtIxXpUXSROpP4Lde
fNLyEdReQFnUZUUd6SHHsXhiDewgBw0aASk5PSpiECgZo2LyG7ornmcLiFwU
7j9GC/ou4+ty/xDGZHPEA3puemEfKGfWBlkRET4GFS2I1sG4LCwMElZELfe0
M7+z4eu810o34o8YsiJxdkpS3YhGJFXpBPZ8pGBujXyZwcjW9mpANEBmf/hR
FbNCblGKujJbOh6ktq7gEEtPLcWpXda8EYsUycqfDVKzYTM9CiZ6AdGGZEpi
X8UGrtpaRr77JiOCEwXY7mfy8mt9AhcCr1ePOmrYeLWflF+qYaSN9/2kkGku
2EEOAtjXebIpbYbNL9zt9uLyfdgFw5LTTkDu1RcebCGCBMSrwKCiomB4qu8c
3MZmEo8NRltYLyJ9WPNs7kGTJXZKu9TfXyK7Lwma19f9hFhM0/X+Dpsejpsn
mlyvnbvvroHrcupWVbuzS8PmGXzb5/l0VrJrNbbbHoBSr5fY3gUWnCd2f7Gk
H7kzenTMLlUrxEiO+hkQVtlkfuzo7/6msiU0N1whY2Rm/SyUWOrpyH3hIeGY
aiQ5OlBP1eCUrBZTjK+jOO2xvtkeYoo1zIi99pwPmtQFxJQ3Ts12WnD3EZb7
nSeeG8DDFgI8muGww4UGhxOwb2ab4yWwltiEqjzm/0o4eiTRTReUo9U10ion
5pga8Lf7AYWCddT/CHKW4cq87Jl8l4jlt1r8z/iXTx5MjclITLnPetNKo9Fy
lQBI0ulFbwnXLIL9R97yWdShRzIo4KVsIT5wGRZeJy1JKlSLfQ0J2Ow2gYrZ
fFdz5OOwmvcFq3T/B9B6ytqKcKHQYnRcIym7J9cElrauouStZpqmY0f1xKNh
aZxjS6Xy7qKFlAZrbSKCqJOhJsJ9aIr0oGBEFhqm6K5qjUZOJuKQGHZ2vg1E
QSeOzg8/tT7KFmU06Qq6jyNKmM5TRUl36UuhFn/PFfE7KResgNRPTqKrdmYp
IPwl902nvc6fzmIUwYZG6VqTQ/+iSJt79cnfdK9F5MG8we2uFdeG7EkXe2wH
wKnArAcxpOT92tnOduD1ApsiphmYHp9YBAVJeKPf3mZ2FOOD2a6iT7GFoDVI
0QM3JL1Un5wX4UWQZ9baKuBRCJL1uRlg6Oq3EEeiXpSAu8F0q/umDuGOR/bu
E1gflRRhWpCnqcE4wsbwYZR9jR+kXY8E9iI2b9LLr+59bXLpqhAX5h1EHj8D
YlOj0vF3eL2/U8367CwRVntdyWgFAAB8NpVjpKHvk3EoVo8467NBhxfiNvph
BqYnaTzlJeQCPASh9LwsNRAQbUDlP6DTZIgBSyxgJ7iLFNjVrf6DF4ShNQaR
pfHLyHflLKaKUg0rpm4OpJweG7SMHR19qfpub+okkboPfn/QsILFuT+neIs+
HFVaiv9crOxw5d/J1z6x/u92UTBLCTS7ZALcDbx2DOCeYJraMQJ6FGcAsied
tVmjdMW5k8nZxhsl6VKt9sbe9XfEN7wvXSFUxHvE2zCbfx9zIlymMSMfaoFl
cRIZBbbWEnoN+wccAFKZDQ74yZ2d1ucrtCXLeV0MBGss7B7oHdOUzvw1pLXk
BQcvatZ5okWaNXjKnDJAUzBE3q12dvjh+1uch60k5UiQ5mKFpXZOMpXvAyp0
HY1qLIQ4TGLlQSLTpPvxCtyA5nFppc2DZKg4jeIbmoWDVLFsJ8TcenrT/kRd
vCNLsBKlDdTWn17u1ukwxYV2v4JaLVcT33jnMr32+5tfJAJiWdPtUbpBaDEd
n9La7nuS8h2Po1jUnalErD8iUME2Y6nSi51+WyP/l4wkcEy1ZeAT92togxfK
f3uZhmlcuodQBnmPU31R7khenlNtTrD3S95i4qcLatci9BqVYqX4UFCVQZ5J
J0L2Yx2tfyz9R4Fnc6l+vBZMTDUm6OAlrvBN7lKlt7uOlGR49b77ZF6XdkAw
1rIcUgnm10S1nTROpVDkS9GbahXJ8w9QLvVP+qK8rvk59F/3lcQSIwTYrl4Y
fxmL+z8TEx6Ad9XXWhqQEfodXVQCP9GHqXGinOChMfrGxc0Sb3Bw/8vcsgad
54FTWu/nR86gxWcts7dDUDOw7RPOMebTfPZCP1tp1wkL++RrzmC/4146gRU1
Q5llsaYpYPkuwaH3F869DO0p0bCHxahVAwYFZRlcCSx8YjzYRZUgJnE/r95j
0Or7aR2Aw+sWqhhqTvQco+mbkmka1ypj5sM58jt32HBLN04oZ8uOQ0/paNd7
1oiYrtqI5OWSrCUVwmzcQfYewNdJfhBQKOrJ8zf8o+Idx4n54dsOxak5S904
pmfrKCbDIGkfZRxtnkKiGv7LdOvN8HbQFlTbgXO4VsIRUVDTNU44Mp3E2zjo
Bx3Dm7F5x8geMUYPw+ZTzHOtAUUSIWbWrFyz2XdYxXnhSYZUN1kW3Kh3SSU2
gPWLCwdaAuYCx0E3UiOdd39HtSKftO4vyZ19DVCtUEm0Js09jHda3xkdH6ZK
8LmbY0dR6NT04qQqn7JwfERh69nkipOUYOLKC54evRFnIizTgpb+TftyRN9m
CnPQuaEntb2m/j+/wzkdnrpg5hO/NKtK/VE2+WysMdPZeMJXZkEbbncfIhhD
50pWBwxLcZL51cWPBpq7Se/owLoOfKD6XYUM9V2BDD4MIDFe72HM14Krktcz
NX3OJad55EA/8gyJMq0iOeDdynihxwYVi4f6AR9NqW637J2WZEe4ptKN5CRI
o9uZkLlze8VErX0sHDKPYBKz69vzm3nIsMLcbe6pWGObBhDOpslDW86vTA1T
xwyZRdgBrlwOI6td+NNAbwL+vrFOiv8aFpPSWBvbrk2E88QKLL/vW+zfnmUK
beNLiJxM04Gag5iSARTBa3FuaAPWCX0WI5wZgRpZXaZYPNWHJMHzxTPxMR8v
jhELZEmsoLmTXDTZm8xmFh5QGobvQKNuHhepajuVVRyVcsWYfRA42R4YSvyd
5uQsrHRQRP/OXC7R5ZPnPGKUyrj7XGZATKoem79sHLEJ7IxHZ6Jp85EThFEW
XtaRjCiMtoUxvTqHtu3IPCugF1ZtG1j2zvVvvaDkTV+LZm+8FEXVRUu8sqQe
t7woXNjCgn2XOqh4ixXJDhY/I+kGl44z7cWVKULEndBkn7G3UQy7F7x0xxjM
D3YuNA/MbA8pOnmFrETuT88Wtu5E4bQp91pJuSXcbApIfNBkeCngFjf878xO
FnARHDU4WVAZVzJc5ZwbF/IvQ040ye+iyf5AcHZqUqg1CwIrgw8XWdwr4je8
IqraC1KVjapiJI1dEfh3vCuzm7ve2DHhlmnqw7mf0rrqyvKBGKx8mlyhpKjJ
WQbE38zNQ7pqckpK35j4ouoG3Bl/56W0LE1J1TxHQPDrNFJwvkBeghlRiFdd
hWcsrWYivaRX10MOs2INEBC7RdFJCoG1J04ke0/tjBJl67vTVVClEG63yo9t
Wx7yHihLg5qG38T81xO40IvyoV3fOU1QsmO7jTCNO4J7sOwHqmmqCdfCYt0K
uSBRSgPcplH5n6GsvGT9HGD/MG48CMu92v06COclefWvkUSiYrEotDrPP7yu
R69iPLjnHXuqegVGmgQ3tYUi3gOqmfdhFZTVC0pDVz1gL07BUoHV1MgS56Zd
vMHDdjXBZKtl4Vzs8ImHaLzxIXuDj0YJ9F1YGYfB3Wdz9aEG0A5oSaXn9ll/
lRxI5gB3ssLHytiFHyKYcC1PwZ+Gz1t0VAlGLahtmgvK1/y6EsYzz4i9aYIZ
1n50jkHicSjxthm4FGuSn7NmRxy/Xoq7ltvBCufRS7O25kObwgYhJheMAlhS
eWkBn6GXrJdCpjWOqlvpvJdyMk7OUo5hxFwa94b6WObDTzDnWtvMz7PrFevI
8p0GEW+d9YhmWgppac8Oca0XbF2h1gO5JXhrgs7fpPAsDI7oJhE2r2cFAOON
COInGZ5KM7Ut5QAzBKOGE/Ep1rYw2vVyMpVBb8iheqN0Qj9W5inIYOdJPi1n
OqFr9+U8myJv0VOFJ4PU/rF8EKzJtXCZlJ0HhDUHQRBOjPfoi7xPJNvbUD70
EXQtXi6dqmseUPE+AyyN9kUoIrgApoUInsjBvhoymn1E8mPmAfMO18Fwr2b1
iNfQhU65SNxPMfBtuzDynsqvhDSbutrw8Axk49ry8Uv2LJHAr79LIFB4b+Gc
BKGG/W77fvCtsKvZQ9dO0PUk8Oso5q2WG+I9iImlg19bayn35Ordo6SDd0WP
8hM0yBKW87unHi1ovp/i9AsIv8ab6YFcwl2aAsn7C4HeMhGETFVcivhHUrKY
XUmb9ctv07b55xKpcyceNJqNZmf3nAiD/3BP4JkyQuvtHnnanY2Mk18o4cqL
q5cjVj7QCG0P7QCcOfyXFw+RuRARD0pFU4g3gcTlB8xhSWqBL4TW5Cf1YhX1
y+WU1KsIj10Cl1/C4zjTnu5Ks7V5G/t9b+O6H3Giix7lRzp219iDbSyGwQEO
mOJkxC+2dDQIVkx/mxIh2koFYEwwTjVkyToXx5kS+29ojS33LuMpOS2ohW7t
Rto7BcqVPEMUFypM9kCuigNcuijrCjUi6OERwPVhVniQncPUhiTft9NznMXL
5Fx/ej//ereg42t833unMMzzQrR/kp4NB6MPfZO/WOgKetnRrDXHp5uvrA1a
p/niHPNYMt/eEgtlP8qSA8ZxUV5sez8ojxu/pp9uGFStFhTIibObB9SAqa95
BHXKI36+cJz4+ovFvwQpqUANNw9jpr23Wy7mOGydXGvoZh1Xzn/LDFuoKCNu
z6kaZ98vIYEjIb18E1rcKYssvpYZ8dhdnNRbkoD6AuN1hpBjEV96IPc0QWek
ffnt8Xt/l6hHm4+0OYsV5zGYXzRY4DnZVNDONSNYdZws5EkDJcOAQa7P+F7S
Fo3+QRvnUG8Ar0/MKEAyfmWh+Fo/ZhCVKDqmbxLvZ/RbvOzEiZse9N3mZwJb
sG8L+7uaDXeFMMtsbXWI0ltAw1J6n/al23NM1AACb4AsgnWjfzpJbyflvFPM
zxU20uSNjF41NMqvBEs3Ovl1i4+D9xkRGVKtpoEtn/rcunRTm86mQynGCkyR
hIdLr/hCI2TAQMWNlpXAAqZrBCV4Uddm6CHIZFCa8zgaDXkOv7JwUk61NlyB
yQt7JfagVLC/YexUrcAvQ+8kEKtBISnCvWxtIaM4ys7be2wqqTHiNFvVOSvg
jBZZjsK0plrykDzuZHFMO+i37zm99+8yqBXeQnrgqibncPHbHYEbDmn4b4yz
MIgZGTvxd5RwOUH9wVsYr0IFNIJSTHcfCTeTE6q+SqyVQ7dAa2EtZArRgtL/
TWLaF2IfV7oSaMr13clfKtjf1MNzgW17hPkfVB+hwMr0ZmdtJKSW/x8p9RS2
BdGFmP/yJ/FC2U8+FGj3jzISspcZL7vFg/6InueHbSJelf5SF8ZS3VLJCZKF
/s7C08bQ+Gd+ZeDhAmyV1Xz2ECWkeuWWHGGHGg/2mT/W4VG0y4WjfaejkNyx
OuxWCn4aJp9oIBtFFW35G2p8QZzDrwCkzO2llT/whkJzyjurVyJ3+PkWR+u4
GRSdVfA5JMx78ty2ColJQ98GBxUWz2pHwKFJCT8i1wADLsKE3xjdxm+yq/hK
Ca+gVr5YuPoxxuRj/IPw3CQM4VMPY0VNACaixljVb7XKj6UcGxXgjY62McRs
LYSIFpmC4km/Z+BvuxeSXykc8IIWKKmbtcgrCueE+97HIkLobLXtqoSCcimN
IbdYXvu35Ncao38mEJk8U0ch0kW5kGOk1wBqm2nWPv+hcXojvvLV+6XLMV5+
94CyyhCLQFCGoqUCfXx6w8oCw9LizFsZFSqNczDnf8lMeEu9BjlB3F7O9iM1
nS8KDhdFwsEQ5GygwU3TFDGQuwLdB61+7gufKRyrkih1T8/7UuUeNk3Sl4CK
3wUcJMyCkdl3Z9NBp1FQf7z3M/WCAbRvaWjOcZgTrp3r1CiUIxAahY9LQuQj
LZabCk+cPvpdU+JKustpssDSyjgrSFjD1TCcjngo2vZ4zsxB7jkfXlXG2AVd
DumH9+4RmCoDiYqwGSEBOgukyMXJnaHc2Xhw4TQF85tDrrYzU1BHUIKqD+9x
imVNJ/OEm0iSBaePgWCKkD5MzveetfnlOAmStkbRj9jK/k0HJjS2PA5ZCJPJ
DGahtM01+MU497b1ekpMpiw9Ta+Uyr2CufbWS0nMPhpN1L/rmu0OTxMOJ8wd
Apwa2mJ6okl4AWgYfDDns2l47c3rZ/lB6HArgwQjD2QBy1+pQjMnqRyPDR3A
MgAfZulu7OoePr9/T5lK5QKYF1I+jWuBW+573R50+BIEpXvFMp7I1I9jaxYK
bWZ6bRb422+ILE6AKeMx9pGGzeLetvW447etMInZfQ9xRhF9Zp3UbtzJgrwE
AvsqqJx/Mm9b8/L9GyQxDXApb7Tz1HABFZpDei4k5AARwbV2ASS1azLl6cfN
0v65VIpdM2qdrOzLp2IpZNnchz712vn/8U8ZyqtIYQodWdF3SeOWmu8Dj7Kf
FJAESbuXuHIi95giOobgy+cTbDl2Rlg5O9FewQssuDEpgsBDrltkMrF12WTD
NMJ/rmHtPT0iDgsUGpyrBiG13Rl/mFoE+rvH2RWMMaowSRcFH4bTm6jNsIvb
/9QbCOwDMmn+YlavocEplTpGSvmMURwSjYCvsUKXymHJhQXdX3zV4TVvZzTt
ngWPPb4BdSfsJKA0LktZUFokZLGBqD2xKaPNC8C+M5xB4k0uMomOI0rARR+2
sqaOuATISDSlMWK3s3FBSIvb81ZBN6iCtJamPbM0F8liJhunlB4ZGmHrLUSP
2p8mwWdt8Cim+SMhRxG8yjP8k+npfbtPm9DI0FCSsyJNPU2K0HoGMTmY1qJ0
qRT9JGnCGrDpsGzu9W25Dp6MI00ibAlKieEJuUP10Z3o8qhf2zgsUzF2geN4
9RnSo0HY2wnH3kB0zpyHWhjSTd6/yDjY5Ax4816O9HDbmxfJhFwnDVQTEnmI
nKlLYV2QfV9CfkUkXsEauV64E9GTUJmmkTrry8tg6N1Y86I446ICw7f3Lb3J
VreMOp218Ir0m8VoHigSbMVqCIw6e0xb9eyUL1nKN6TzAqrPMqyue56Otpfz
Enhyd1PtTsxgK1SRcYwCoa+Mco1L6c6zTeo18gMDbGSoeA8ZcTjzCkbit+Z8
eNBNPE9/00HQCGz0mext10p8s7oUXbONdIYpkGzPJDMoDJt2lpkypKMyZE2J
OlRTqn67nPhYYK7ksyPCaRi9NzvYJbEuR0TK9Ts0ZgjkimbZnyLQBKCKHvRR
cxtNrtfTKMPOBDC6BEY/bUxcX0Q6adhUMv/Cgl++6MetK+UnB5ty2rCfz8ub
yMU5kZvAx7g72OJqUfd8hA3PZFqA91MxmfrwBtSPPD1qbXvz9AyiKE5+kJRx
AgK+XiVPwm/TLergGIWyBrQ6cYD0ZXs78JOUuJiDnUsNk/XJc/QeTnbYB+ZG
QfzwEFv1lN5N3a2pRDYFxgc4cnyOpGkaFYJ2EgbcvGdSKjTjQFBVdaAI9rC9
svb4A8LtmmAem1ZCTQR9sp9XYBoTtvab3HXSe/nQAomcw9FlDxiY0aVFt8b9
D4hzxbNfSR89yqldenx3TP5klX21hdYojHJsC9rXXo1nmBpfd9qdIihtvkgo
GP0ZDbzXMUYd42bIO9gM+HHGBYmTuIVP7Jp+6/+HpnGP2wt6jcOLJ3D9qJio
Qz9erUCFrkuUvnz6qaX/bA6msS8NkTIfl00UTuDv2Z7Rcb3aEkUhBV/8lCje
vmNVIq6wYWVq0S7taK4kjshXlg3XNomfFx03wbc3s6MrakoA2Dbo2PasUuXH
kHtL0x5AbaZbz03vMF1zHFxhrQGCGP44s0DYYZqYTsWtv5fnm4fQP27xZc0Q
vhtHJRfUY8PReDBB6hU2ezXQHmwjZlpEIAAekj0PG+OZhV8aSgoeX6VIiU8+
mTOpYLh4LI18232401IL/CnmMvbsPUHjifmsKT8v02U4Ij5By0Vgrp/Cg4qs
KPVXzNiC17culkO7oZyKXmK1i1/ORlv6oh+P6r+3CujK5DCAe1pB9D7wDlPK
FWf2+tX0Wmfx6dtz1ZMOBzB+UG+9Lxtc+/2iBvRtr9kqtwweTd1GRMpLXTRs
EBJw2iN7vebNZuj0JAa8JtpWTJDR7jViB6XMOogzLmnCHZh5UNMStF2qpRKa
f7+frhPBAsH8vhZirx/isvoO2H11o1d7a/ygvNBuz7V7i1Uii74oblKdloLS
c/uwa7N6DQke8ZmXk+Oxxa+AxMKCvrX7+GW6Lac9xZYov7IOkaJRpv9aPdx9
aNpJ/nBneVkf7kovPUjl3pcZhgtyDf2kEB+liCYz1nuBSXOmKpkdUo7+SiSJ
AR8xP6ChQGoXvpNhTkqvgMAY/8z6BKdUaTMRr3/XTsYN4TypenHogbFtVzLh
FGSO85SAcGgh18G+kPBT03rKDlNDcsVBcQUzTR2NIkt/wfWeux50w/K6XRx0
OQVWIwGGaq8Mh7PUCgo0CQ8SXrAy0cud/2IxtHI/VEq53UWj6GgxAuXBx/C9
klJIenZMX+nD+3mJvXxKMZXwuN2IG863PVcfLlqyOxb95udXORKfjuSWvX/9
CJWLWJqctVO46El5RMDA0tQIoCHjfj7UHwH8apdoljiZJu6rej8RL9hf79Rv
7+4wY6l/XbnnZomfq20VwsQ/wmPAnYzuvU+DPdzrYoz0LBQ+ywUjeRxWikEt
OOUElSjvglHzmbXX8c5qjV/Mhm52VwHbX8BZQIwyZ124b13IR3n+Jfgp9V8p
KK2fybmq8aS8gxv8k8Cg8EWieYGAMZAkj41ONPf7W9SFd1OvV08TYmrd5CVa
v9HtHq0V3+T0yQyyClxz+Z8sVJ0nIBIKSC+R79cPAnGpw/ybzXJlCGyteiTX
sAzN5ryJFiDO/GpBXusjvzwzwV7aJhhH6Y+WM38L/e6VhKtHLpakbHxW9h9R
m5muqB5Fg1aj9x9pv9UyZQXDPZQDU+oyT+s183aT4PVvkY+/OWEvFXMVQGBy
hnb+7bOq0uIs8CgGse7bzh54DD/o2AkrnGCPMDHq/xzEEcbQ++WQhS742F2u
zh7IY/fd11CDygmvwST+04fTG9wgvsqZYJUxRKyAQl184jfnX+OnfsAQfqbp
NQva47UnjUisUX6NDPDnQMC8dLQE5TLWLQb0vtgRsV0bP5n6Og2j8+rWg97l
3QaPzBf9Hlljj0wr4uJATYGjZHkejmg3CHcky4BVOW154bm4NBT4B7xKfQ22
UH6DoO1QXeRhLINVzZ5+bBaxcBvCwHwj5bKoI513onB0bMIsVauvEtNhhsxk
x/igWl1ckcu2gZPeRB/c3EEV0izGOayLXTIkGpIUTAe7EEja1VQTpPXxyMiC
YBn7qHv2XHkNsiFMkDkJk4t6HEwRry/L4KYitQZDPN0/Xm/6NFjwUIaW9Ier
YGdoiiHBbfPBTGVS6a4BZaT3Ydelk6TtdWBDprzEzocAMdfyQ4PFJQ9MzYjQ
TA70tVNivGOqFHcophaQdRqFqoQ8+0hmT8ksxNmzNYYZMVeXAF++tAnue4bB
14cTmHowQKdnMzJIbQwtVy6fXHaDF1tibMY99+o5bWJXLO0yj0O//8JuyQ5L
pVjmThJSIl18br6QN1CV5w0yPiJzB3So7Hjbj6TYdpcx501hquB3+LhUioHB
/8qPvYCych7MSi3BPV8VHhqwymxm4NpEapoX/1+teg7hqCS8mGwpNUi31ToZ
/pGWJILLRkQhWXnLgAa2dMi6oAxgYO1vMKOiaxnb53miuv/tiCUXs0Wkrwk9
KJ8Zu5raQCWqfa9jLi4GXcJNIFGxzOEymu6VVXay8vQ/ud163AItVCJ1VqPB
AeP5Qq8RCsTwocoMClhUbG+pIOcA77vGaHhfqnH+Pli56cA1ISEOImomAHH1
xaW4c05nofABTf6O6r1VSQX/ezWBDZxnd+X/4D0ZvXYgumyDOdmIY86sLp7f
rBngMvIjr/jj8xKqD14u7xpXdytUYQU1yNZi8Y1Oa4YcCYOrxut0Wyteknnx
Z3QB6Brcbo+cSevNLe/e3+USg/BhuMIP2DtGcCS0mUOEOxBOCtSbrWJMwQlD
+wfVSx6L1JqxgEuW9VeAcfMh5hIEXaSQjoqPHLsK52R70ohmR8APwdBOyABt
l4z9HDrp3MHXyIvbyXx9pdBwdzbOEcX8+a7bB1QXJp4w5ris2pgd2SRTsaJb
PKH3rypmcorrPhhNrmjSMBN1TZFys/drg/gxiWkN6dlJfGXqmRaK6lyKEC8L
jVVOmtE35IUSlz2XOMft/GpdU0b+J6UibL7e/AC2j8kgUBXBTj3JN6j7H16M
vuiovLM+W31hTB0wlAA85G0+hNrStX26YjyxXXlejEO3C9LyfjFIyi+0mYGS
V1AZNOE58dUY39gvBeWRcbKP61opvIqBWTpef+fuOoa9Y6OHgW8hPqHU1P3G
rc5FYP8tgLU2iAMr7LR7afVsB3tl2Z4EQ04jBHcxU4vTet4h4doCa4RIZu8t
3GHt6qC6sscJ9jDm/nUJQdL92vX0WNfz10u3M0VlIaRZjr4Q6e4TNWt0PqBO
PUxvOzl0VZHWMQm1LltdApJgK3SrEpjd2XhXrxZvcb9ntHPuD75UgeYBHFCc
BdkN+Yr++HcqI+0cCII7hPDmLx+lOPT9CBFFTJASRIal3kIFXG0oLT3zAjmp
8ic7kmv163lYFZS8WMaTqqFj3ldm1ktJHZv1b5JpEFRuR4Iiz1yLqJWhxvYc
BFyRAioz/sC2M8D2hCEQm4VDjh6XCfdxBwK77UbYtkbR4u+kV37eUKjSdoLM
MapED0WlY94e2JH8uHZGlalrkrZPikgsf/fZSlLv2m0SlnZgMDVmuJO9Dwij
gVW3DkLNfJs5KfbUo/FdSJoBzRG7I+yQxTcMAaatZinUqLGL7zP9/SqQUCzN
oA2S66POY86ViP24ohfWJZjTpcYf9/lD6OOj/HmqZrm3k/AVJTIP6lsVgWtB
LMcXIxVRoH8KwGZk+TX4nTpXkXC4QT8bxWvsw32H1SiIcTyoaoARGvZPAIxs
MGsu5tS8pLj35bl3Y+ZEGyeKs97fNVFMyv8YNiPP7R9ushW5E6fTNfTFrPRb
ChDXiF8Cy9di16GVSEDd2+CBxFY4SvfDwYzGa+ZPQMqJI4iR5c3/SY3I8nkP
coBoTOcqO7IOMG50fW5huwLpd+p6919U/XKAsmcbqj7E1+r9A4ozBQs3g/2E
I4ILryD4HRxpr6jNtMnAmLu8Kguq4vTkd51Tnrk/yo7k3gsVgCzH6BIOsDOs
u5oZRQMqF1N7Zt7V9p6PxCVf09WXRmQyd7FIapadKFpWCnSPM3mmDDPt0y0d
uhuRhnAsahu4itAZTUT7fDgGuDzw+97zY+MnHlUu21NePKWnhkk10LpbvSEw
B/PHLk3dBbyiOMxpQp+sxUCPLYdWA2wXapo0V2xlctOr+kqBj6BnGBpsFTP5
YbxlViWdN8v9rPuc91rI3pTkK0y+hJkTU4nTbKDEOcAYueK/iINeoMLezUP0
CUpCElixG9AegyaWLMka3bwR0ZcamrcbH+nBGTLELv/0BRTP9NOvfmpHvpbK
GxnGI9Lx+KYfGtijhMHE77r+E0AVbadAv8SSFxWqkiEh9HfVYSTp7eufhBDz
lAxveCIBsSq+C28vT/nZpERLx4Vpc4QopgiVPgTTBblLjKkNjGyHpEitMtEq
PwE2Wn28OPgBufsl4aKCSTpSVrqHxP8/P3o1t8e3FJDN3D/bjnDkMeg8FT+t
dVNPBVus00ZJ+sxEtM5VHcmGNKXiOQv5JlEIj4jH0UWDRHUrQ54I81fzh6hW
F1MNiZPCD1E6lYxQeSAW4tb3VQ9onnsAEL3MlmHXLSNrMjdVVEpuJNkNMQiI
y6hOgLlI5kuRWFWgv9CJ3gJHomOTLxRV30/MpJLVcUsYbsFSh9WwO5/iIUdB
CxBUv2lH77l14K7eaumxp1j9fpDABrwydvyiTzJd26ncPga6/JalJ1XO32Wn
IL8+7j69dykT2JiNcOLXnHFPZLEeFh4jjwOMDIpTFXYinjxEgbM6igTQua6S
hE3rZK2ryIT5cYKYyxDe+M9mScYK7HsFttZW9SomvOG2wCZGKGUeFgji9V77
KsB9x+/cuuWJ4ZL4tji6oS4/8OBtH5XEdEJJmU/Wdp+zPvn+YE9DLXpX6lvb
HpeLmJiI+d3V+ti+CNthWrsuUSTFal0I+xk4ewk9yweOIIujV9tKoDl3w/Ps
CPG/5hFmDb2n16M/b2IURCozyXa5PzAVNyGSyz4R1gX5IJBu1ETwQ4xoBjFx
tCmwV8DK0rJG8lxNfSi6LFqQ9+Yrv7orucf59ao3d7wYS/zCCz/p8AoBJnQq
cN0PBGejLOi/+2BJeMU9Y+fZ7qx4Nuiv64N++w48kNS1LiKCos37uLaMluSf
KbtqwezCdCo8QzZS0yBi8WRpXcgz32P6t0TtRhq13kk6/g9mKrsIh/m5w6Tb
w/R6X4eRZEztNeWHiU1EoD7PezapPCSvjBemm5A4OtWq/O2tNuLbiW2gLROJ
GfTzLKH65I84LD3bUQWerKVZvTUQBK6tQwR+hMgwkwiYNx4I5ZwPX974CSo+
81x+BmUF89fDT2snNeid93Ic1R3kG9zZXoU8aMgmWPeNvK5HOn1cRIZ1L5nc
6pa0I4nX1qZok9vtDBVeBNpGh+j905hP6vpM9iY60wz1B6TJ+Kv9LB+fiIhz
O08PcPYpUYn+zGvYd4n3rPgl/Ze9sVzNrdk393mMziw391voUbjsjnvGONYZ
heE7AvsNeCf/JJc32tPLAqadX+Fb137lW+L73IVwelMYTJo0/JPgwE/8Yixl
GOVWsj2uJtiQGsNLaOWQkbQzCOWAbPeUluWBmJczjGKVVQiTCPV+GtOxqgsN
1Uc83mLBho0gubrfD4nAKHYg2RHTZ2HviHowTYxVHWrhVyTNduHhYHXFRZGx
3JLb1JzWYPmMn8A69RA8NSQeJGwMlQ24hSD5QG9SVgITi+CbL7rbTt85LJZg
Yl2Pse6KVkc71UlUFO1ktBVYxR1KGhw/jJilsH4n5znFcL2LKJ4BsJ3fpKGJ
ZUwGON/Jbn3Qgvsw9XUKh0fKUKxXOBo528MBDFGxKaTcvOjinwWZi/0jw9hX
+9NiuBqiZHbI6lCmpg7z3PzOixNrWGkr8NN+jaDC0QtLHhGiwZGxQa4lNIam
LdkXyvu2X3wTHRRawxlvcKK40U0E99vTDRf5GwcdsZB1YIRWV3AA1nI80Esr
W7qk1Fjn7V2fbdGOA7zLAyybCOIAM2TqoeW3qF6MCrrzeltRJuUw521kfXXl
7gI1z2C+EhPzL8AGyJSM/9imMRT2ki8FKLX2r34iuRGyMmrMsji9ugUdN7J8
GFbyHc1BQYRcnhFInXwm3gnkA9J2B9nRV2APYy4CJ4FY1sHUdzXcXkus9aTp
m4FSeKmL8iuD/658K7QjIlUD5Vw7qDcDht4JnSfwIo/SP09B9wt9oRP9hxES
mHOy4eCYwqjLvcYittqVDePtQ/P5+/VQy5dJc/3BDIEAyw8kLxyL3tVURfrQ
dTgQ7oGISxEMVti/U5qsh6i0vjgmb4D8WGblI3vqXWxHEX/YMOvVGHx8bhEo
m2BPEEP40r6FK4MPaOs9/t+kufUNCZUsaFpCJC5XhD1sttth/APQA6Y0u/pE
dPKC5qzoNBVADPXoxLvfPi3NN5uEeq6hbJwBhmj0k4MLLMxtpSRXDKqlc0p2
3641iN1/yIomDa0HlKQZnDOVIII/xN8B8wdRVbtxaTWjt7/26crd5A4WpHq2
ZYuZ2PxsxJ1vGAqIVivbJo/1XwMoKaVmLgQd/MEquxycGLtsAy9Gt37woDkX
HhiGs9z8fPYBB3SqjVkeQYSDhyFjzTqLGb02h9FAW+wUZnKPEEPGQ/SNicmF
VHtYdDz/R9nlyd5zasrPhsTZA6wLjJpe9TNrEl25eu4b98livbJnjUcNF0lw
b9d8XXbNk0HS8IgTmSJhCTz5A/h09jE+6PUFPt2iGf1JI2v4V8bs7yLKC28n
RU7rezjqLj+SZl6sodz2R6wLUHPNIIA1435gcAeqfYkhgq1Jb25JTrx6+S7g
DNSfEbKl0flpQGktKPdxKgTt5j+C0ATXTPg/H81xGUghAexI4sMczxc9CtO+
bdiqd+PSZDcAv0ENhhG6mYgp5EQjmjn4WxmfrdXqKzeQgdE+PcK3ROEbK/9g
nxqNaFw3nq8x7CIX49Nt3byAokAsAefLtPtaAZKlvYC1eZe0hlSgs9ScCNJL
PggSyFt7i+aC0IDyf2ZTdfgnibH+tiWHGpUBq2rgsauO1IvuGiGIot3/tKDB
3C44F0IjMhpDTaEMaPRrPghcYfRbWFXIFBIUg1q0ysTH9MD3JzhXFrdjsjP4
M6tqnG0bFT5WL4Y/0iW2obQYL3Q7RA9xLDfj9X/qmPpsaP6vNcqlXKyQ5+Uz
OGvKwrC07fBVdtg/CeU5gLIjIQZf9ckkDFt0vOWgsUPHYZyMnKPasGywazzd
irHtIHpO1hsu4G0rU7vyZoq2vgK6brt3jkfcfld+/9zeP6ik4xRLdMFS3NX/
coj2wMT9tt1OIkvpfpNKWqLjmGTdE1ZCwHW+gaZzuxwDe7HHiDCm8rdpOSYX
XHr1wYuAfpNtNGssFlndMNNpBHXg8j332pmyKu5y4tVTwfD6I5YQVMP3AehN
nnWnDMsAn19ByzuvGqYsXeXLaZt1Z/wLTthrHKNpfzfm/g84ucH+KvGkA60J
EcYXLvqtMUjhl/lb04IBQk+aVs/M6q/4cczYgiyjRm0ua/0/YYqa8t7FG3JF
IMrpygBRsrCZaCaorMnDBzIM3JFKxBdeLsaqI/7tWHotVSBm6hUIMsQHQTD5
QZsX1tVxLGPYRU6meJMuZKwtU8USbnES3zBeGB4LgqwJDD1OvJOzVVvhymhs
5xrEQ7TL9CFvUtJpjPAlCxzm3xDjsMlhHef4wv7ZYD9nB6bTarSaJhCx91Ka
jS0fItzdsUsCkySKvel0TBFjPNbqByzkHYemepbok7+XCje0MZbadNueuPvN
ga/fsYeWVGrmi5IQn6w0I7o2H1WMmKO4rTOnqsDmNmkukVabSeEh+jrvDts7
5vbZj+6e0xVq9gtszdbg4LVfvewYuCm86vJyMgVE+CrPqjw/M/SlUUcnFgdq
iSHO1a4/0vhDwyUWgdxpH4WE6BKnhIwhw5FoChaLTGCcJFR70kvHN2PB5ExC
IBI40tqpGCKnR1F1ox4VX2tj6TDw41jMM7ryi2/uMtVhkmkFE+CZNUyp4oDI
4PFnnvBRowM91IahzrEtDvb+aQ9na32ng6O0UwBOuMLgDS18Io0Ru7HFP2ca
qfemNQO2ALAJQDmXLmKJ3cXu5mpBDDybjZaJMI96p1cMLYnX2sq/PE0cUQD+
GPlSHfrAlmVGEHvXDSkRPKQJCs/pz3qEbom12jBiJdE2upOuCmLQ8UoBTvjq
L0lqguGh6ZosZR4sr3ho9cQFlf/XgSXBLAfsC7mP014q6KeAzhhiNEKr7O+V
0XoDmL8Dbsq/aK/r6y8Dp38yIpHRDZzSdyMrI0uz0AutzPNWFsTGG8KEMDDB
3fDuyN6ndF8RaW42bR/lGf7qS7kRsl4AiDR1wjPbHLKF18E4c78oEMHSCyQC
8wpUYvr0kDIL73ylzlcmXlAlGjkPCehd3tA2+bdNpnWMuQkQxe1ooJabW63V
LNiXph3Tq+n9cMs7BxEWx07sirpOIBRHpsnDLegBDXjyCbbqWGy8ziX6Ojoo
MCEr3VZZFtyqQDlgv8s66wxsQ3z9Fnzr8smSU95fc3pS/8TDDfNLZiqCwIYX
OEQnxV8Pk00RxFvAUOvqQn9dDcxXwU4yNAr02ZTIY3mz/ZQcoXHq2oxXDgT/
yJQVhHRN2uEAzbf29aAn5NM4CMc1EN7uJn+qzFDPBbdX4j4gDP+qO8HrdDVj
4603JZZ/iPHHRE8bCY27oub2brlGB7Rh5O+B8TPORCvmcPIvhXkIla4QsgGY
U4DcTIqhdo6LjtUAAA83/enlQqCFBat96o1lAEP2FhGOuVVkCZeEZhMgCK4X
7CTe1bJIKnsufFDPxDgdpgorFBj0ETsEFT/q6WuQStTXqt/iHQbcg5yeplLW
0C+RCCMs4u7pgg0vXstDwbDB8vQZoKjTZCEDYp5vTDHSbiiqEQO/y8csphbJ
/6zKl5VzZoyq++0XYLAWdTJKZ1671i8tUkfM3Ho7Bqx1GkiaJKjsiEqxWJzd
bYghn8tDWrWo4sGugBO1A1aE+tJPb3jO3aflxKXiQVa9JCNveRyiMolK2g57
SC3ekmrpb3T6nc0rTaXxIWUubRCBXEIG55RWNiuKVpxdAwckTfkNC4ParXHD
r0W2/0rrE6jSt4Yq1r3WG0oJ8SjcJXVThmWSc8BPn5K5x7bY8reb76Rx8DvQ
/+ozTTX+158tYKmWM0Jq6fcSJR1FA3OBsyP7YQ/ssU8LTDh8FWWhgsQgUujQ
VUbJ7gaa0QTeuAoPyANBun0z62ELpZxvJmZwWTuFEL4ajw1K055urLaKv5xJ
FfuwG7k/fldhZyWt8jtSKy48sUzt1iMIX2uI4b60SgZTVcpIzaI47+cHayze
0JC8g7qYAJN+9XMrujLAemcp0jgJH0G7NPLukiToYEnAgrsoFMHHcGhV8Hj9
WHjdDTTDEKlOknB6V2EayT8Q331lFWUpe+lw2G2vdIMlKsL3w1qj/gGI8d9D
g4LGgzKqIyEU/TAjGkGVbA7D1YsQwE4NWpWBKYQeLvVHduRSBQISxMRtUOjo
Ir0ymx2b0cQdeHNKsMJV8Pr3ac422HQPkrWpZnAqjGJ5JDcijkpQSwWVsSUu
C1FHpCvj9K4fe7z2ylh8dd/icFNSX/gvaffqyz8VzDRSSlG4bP0CUN31gFRU
Wo9/KTPNb9gEebRXVP5YDBRolFqySBa30XAw/dgh4aoHQMep+YCuGeHD7YbU
eSeIXQoYRoxkv7e+6xkarEql3TG3FKKvPoDRqXk32i6MUwcdwrKmddHhqxt9
/Qvh5JQukplDq164hR08CZW4+kynKsdAxEnlsERVOGt7eg523E0UcSiCe5y5
/Dj8ciLxVc1huNJWyFhvfo5/rd6Lg0/RVxoo9QB3p/eY131AdJ7aHSt7/Up6
NFG8JcY2Q0X3emOBdy+N8KOZntqiqQm2lojr0O1nM/qMzMlCruG8g270gFD4
pgTi/33cJ62hhiwVhycK+P2GnNpYcTlK7AUR84VVbaYOQ4k+vg11GybUjJwN
e2OiO+Oe0KQf8v/AggoCvBaEcq7AgL4EfVcKYH2XTYLf+2vW47JcdcV3hOi6
malU5/OIhbL6OHEjfnlXNJF0ltD7tlxsRP+kGFKYMAykb+u1lE6SDknt4ubf
AaukfsiikAPuVZ1tWBd1nAYX/UWaml4nQlq0JUAqbpyWDYCKx8W6zqdFURgn
XwpZz1IOBNSsqdntOh7ktwGBncGFqWfwgffWKpsuRIG5Rk+F1JMnUJDB2d+5
t4If21kER/Eaa8j1P1RwzEcBuWEXcDJJhrD44IudcnZ69npT3REG6cEVd4D8
av/LWxniUea8V//RX17qULqOE3edEjB1iFTDdx7bImBkB3qNem7vJDkQB5+Z
6Q8POjAFWLT9eOV9vGPFX0FSglSvlUr0D/x1gyzodhZl726vlLEiIuD1nDU2
2YsK1zFmF2omHd8A6TZ3KX5Uf3TnGrByUOin6Ew6vHUlzKOr8yt0HpAgHQNu
ofWMfSfb4d4svGFMmfPShvAup06/ZUW/82rKn2nZSPQg1OuGtzUGrrI++YjA
d9smMOdREoGw0xTnLojzyHicWB1NjsIFFwbzvf4qpjjTHx2lGvVAKaQN4bmI
vj001gHCDRe83L3oOsFeBdc+j2KfxQtmaKNwlHCLLJIcnwMb4CTirVkEZnEL
DB+QV24jlXkquJL0vaZUav7/8qkx1NyM+dhgH4vOUGHCSjYuSsDcTDkbzR/4
8p2WVuYT8BsOMy8brAgB62Vx2diBMnoH6eyY3ruDkaNz4YIkw+SIfBoonJ0K
udcT61CHrl8koCGtH1+0Pbv55TqWteE24s3p46pZQ1nmITYu5sdz6aOsrv6O
Dipe15P+ZNcwQEz+0FOgKoibT9olzQxVWBv+d8HFscQKLSD+H3Dpd5N5hqBX
3lAxWbIMB8F3eW3q1PFkEQjfcUHQU9F3q7VmkzaE/QMsOFHRkIJ6laln+GQs
Iz6CEC+mUmRnAOtZdO4OPTGF+TdBotiu4KhBfXWHdanBGOduu53xQOsyrp38
jWgTVi8NIJF5GE5XXkD2gM2tg7P/OKHefgzcM0OE8yXgv+9Ugqb8xDwh2CdB
qpQfrBmnfRmq35r1Q8XVyXYKLLrEzsqVYoUG/4P+9KlwKide+I3fSAgHlb1I
g3Do5adx1E70K0yGGaciMwbtL4f3G1tW+RosaZk+dajQ5EV3BPYxo4sTLIqj
Y2EYYEd6JpIkwXaR0nlnAlSqkLWmPRKeQTJdqGASALv4+K0Ze6dVWh6JgC9o
OyA7ccJrlGK+1VLvq0hAuL5MA2yMgku78yuOcA2xE0AZXoxqnC5NCWudj6td
wpXT4/DtON1dYuvvopkFjFI/3VMS4sQ9lyIt5mH6WncQNUb0N3wiaEfUpuDd
vFggift0T11g0g9AF8Xqh5Qiyy/9F8cXzoJIkHIOmBmzEVt9yXz6GaP3j8Vj
9DMhMWHx1w6ASY89o/zlJv/UaQjXP+eqRvbvwrOR+/aZHQYNQ9d5LzaiYuMH
rr4ZImozjB4p6boKKk/8uwqnIQkXcj9ATHt3lyMn64txZpW5IuW7u9iOZO4L
R4/DEFX9AJLTB0ExCLsFuTh11LBDeVLEN7FLM33b9FFQC/8nrbugaFam6otB
2Lw5oX9bK7fYzT39hB4UrlSX755oztKvfWOR2AitU1oRJJSHbYat3zIzqeV/
VUPBLgqPlopEOFlUA5ZRNmBcllF8pRaeQajgi6oqJ4Q5QqW+DJxdKNk3Wzpu
fBc6fp1Kygroh9orWsWzGzutQmo1kSt17mSw5Yz3K4sga3bkeMktfT+N2NFN
7R+f26JgY66thLbLTA+MhBvDfz0EBUpkqAXLZI/3puA91sRQ2ud42cz38lxi
ZrAUzYP7d+Ithl40un6sGBEIcWQmvYV8xSyCWTgUdWMGjcym845NUPGG0gDM
JUpabBrhpAE9/iCeX3gnU1BnCDkOWv4bD/ZRPssZmS26lQ2HUw8LB9/zy0FL
FdyxfpkSdsFqAkkM79aYI08cECUN7nGeUqAAslI4lu7HAvyPVUeZ0VhS7HMg
Gze0ALuHiqmtIHvkUt9b4MhkFEgshcmLQmmiinGFJ6YEzl4GRPiuH/aKqtFW
GjPtIPwwxPd0s65wmJyMkVwQu23RjO7kdUMlw4WFI0iwqbM6/tR4EUnIYy/k
SoyrZ8tmXxDMmBkL8zwWh8XIPpKFPWz0aYLdtlJ33TFAPgX1AyrESRoM6c5Z
OgIiNzPofYZQLoToqBVt5kyIz9p73oMEfvkD45crsuu3lIHkFFahzXxk9EpD
M8defukRoqLFl93EEtjS+fQLeQfVKN7tuDEy1bJhC5B7cKQAoHkIiPb7NoKI
FFVrCZtrU8ogRPTH7NCvts0NXislGPzWDMCYcI6Bsm4AqdVy29Jn1oYOWFZI
pl4DLdD285hjKK/6Xg5c60ZQ2TKh4KYc/Ky7angTwNwhHGf7gD54P8YhrJOr
xpPTVIAyhHSHWLRWRuZWPS5Ef50BH8+t0myBI0NZjIALRrS7jBBTEZC5yMoB
UZ3IiEFPglSTYYQSfbqKmd0l2L6cCLw1cPiGJBXAyuLBZ2KJHwmYHvaBgJGN
rEgHJHJq0v2a3+1hle/rK5ptWr7Ac5oPchS97r5MWNfvj48FVql3jes1O3D0
q7jNTIZf6PR2bBi0IyR2Nob+4MJhohuRA+vLcHm6/98wKgdoPr11obQQqNaG
NYc02M78JHErHVwUKel9lwx42KuZIoH69AHfuuKzINM6Sd3QSBu32cDn5kcy
vYO9gWcXOGrU+HncsZaINjMEtof4w9MA62Pp9A+ydgxFlC+5wW9HtCktMcc9
wUGyMwevOYhkC8uXVhOysaJYZBv0X0QVIXQgcpFdfTaqT/rh0aPqPBKuszjm
h6q4y/o2LVlWg0qTVKMq3C8FFfCa6N9HekTa8PhKgl/7EQegCVHn0YM1rbx1
qttqrOPRwyq4MO4hI16cDBAsGb5w+11IN8B6masCN6Z8OHPh3Px7OzdGIGZ/
i3fP3YTRjqQjrBVlfRd/WrRm7MkYA63KG0+n7T27WBUQ+9pISVKgMwWMfM1h
aNCnjLBPJFUP46GMClvLX90b1eqDLULLQuZU7J038VHlacge15EP7Oq96WCY
LDNysjanrJIcxWcRDHGXdSnNBjQg0OtxSdFub8Qz8YlGl7mbLGEzP/7MPeuZ
c/A92jwkUW6zXZuSyQAKDloHBDX5e7f+7TLTKzaKL8EJAg+4UYHLXZ9tB9DK
yf8PoRhsyDK1BroEuHLFc9ery03rOslicmcizPmli0l/FU2PQe705TuCCGLZ
D9hSi30Ja5mo+GZvd1+HxKMq82+J0N6q5U1B4LxG6thbkfNUPCYk2UuuBXuQ
iGseD8ZmpHKT1BTyqQ72B+tTaaurNI45WDEmNEJRcfNKmupCeyNoEWUpIvWm
k/nL+nX73kKSz80yAr6B51dLBSVT0iakxcmfxGRXJi3IkQElBKWNe8KmSA9F
Nri8uja114gEw+CIQtjAEOJfJe4BiTFaVs/Oi5akROeclijImMGbWkdBhFTE
BY0YJoCu1h4VqohFdkdLR/tFOJFPQLCvUkVC2aOXq9mcPCACB1ORg1pdx/+l
TIEjmcYZ8tJl/MsZDNB4xJxFo91P+TtJj12cxWGgB4Eg1M7cDu85SdChPNmZ
NT1e1wINnddnFm+icc2ce1CyUtQJI58ZYzKndZkVSeBjmL7D1gZqi+Sxk/wY
eKG7Kk1/TNEhnw1wYEZeN8+XOQ5JX5D6rf1yzBfVeWBpEVWggA+YQy9zm7vv
2pWvkHaotd+ssWOexLFuuyTHXaA1zK3DIVLOLq0DA7qvSPeirXJ9OLoJtojq
yTMNd7jpozlh86bhXaWSLsL1Ct9CFOHqeJOyownGUFIqKmWEwaftzVtDobDD
fRYZmpDPCTeu8KBLd1gjdDOAKvdbKsIRHnvGIeTanT9rixP6JeU5Aid7z2ow
bRjFmmvoaBZ8uwMkBKOxsGdGvx5qh5656uA6qFaJpF0drJL8yzOnamUnJv71
6G/jliPOQr3bAgUPcQ5sJWCiRMt1PpW+iTnygPw936kzCYbvTQbGZPSiLkf7
f/vttzM4QxGmfS9PY96iICeigvx3r34fbRSor7u6GA8fcIIFEiW9Hf5XbXf3
ZsUJJCZifmtGcZf6aI9ZsxZz4GZ5L7zAlNpaoRvoAu6AHTyxGvHLp2WOHKhl
VqDjcclIEjE87tDmP9Ryx32rXghMEmEYeDHic18IZBXFqjAQ4pIU57rZm/3Y
4j2VK1ZJU6tSrkWyybu2Ajt2uMEjPHdFEWPJTNnDZwHsap60ruiZtYLmOfZs
B0Xdz/Fxe+R0URiYuYKRaiqh3eZvuWMdmLywkk62yUqv9Sv8FxzOXnHvFWfp
ujJIxWYpG5sXNURShjDNCrXF/DlcUt/0mX79fNnFmSVn/9nOMIA1gJ1GMsjP
2shni/FaIZBn5NbUR0Vq4mO5jIrsj2gA4AeEMwQOpMyq19NxvRvtJArSyYID
jsDkzKX8eZ2kqRCXRBgLcOKxq0cZPGpP3SJpq68n4jXDIWg1hkE6CZ7EOfNz
Ca2M+FF/GmzyNIXMFPQXWJiDJEVpHs3sWQewfrP3ODw1H0QObnHv0uVZ3eMg
wG6a8ja7rI365EbbHALQdV8dOZ7qPFCBXovvc6XeDz6RwgTmQ7X+vPVef0wK
MvqEjIcG9OWrssFywFFvEMPbqjizeVdRJODrqAylCoXdpiQ8kaH5VjyB4XKV
uMUVCvChIAUkvYDdYzbLyidnC0pIO4SLlz8X2xKqJEKZRvaXv6Z5lM2xGrSr
NtId1eHtHdLKlCO3eCzhj0ZkTfurw4lgidWl/OJ9LZoqVpMYOYbCNWBnDcqK
wCuURetc4zA9FIKZBjIMr/1VTlslzlI3H7HdFqXX/UJ4s0g6hZ5wPAG+ZsC8
4G5OwzA/q2a3ABEki7OUrAj8HrxzfybbLNFVelQ1yoJrsrAaQlNxgRXTCTCi
TXgMZVCuR+pagHQvMZdc06jXNW3LebCE+wZEeIBP+lf6CRHLuRqkpOibWVfZ
MTnK7Z5xXuNstlMigIBFhrqHRqP+0Dt0LFKyNByVXLZGZuBdVznNBVLRDMIp
Pa3/p/NSiHcsL3rjiZnBDEy/ABCyEUH+4fnJlmapG+o/iUQtCpOBV+sgcisN
Y3m6jgoOgEpeHUN4/eWbuRQyUDRjKaQfdlbzbNwMYVrpGVmkpQammSR404Vu
T4cYiLoC8LN2nuqbghv2jMlBmh6oQf08mEYgESUePBelKvyNuql2WvwzWG9V
ZVOA/OKt1BxOKf3WNt5eO3MVpENDa/YBKoZ7sHl8H7jMLp9IPHdZ4r56+Cl3
Ky/A0NQekt2UmYbYaIJlrhTglce84LCUfRULcbeK5THobtnyckZvL/u+S3tt
dRMWNF0EDmXnOlWiju+HEHJkVdNBade7AzOrrVAn+xzmo7LaUrjt+UtrUOBR
8ywoPMIZUTT83ea/MN4wcaz6H5cQNO0PNBPGKemFEZ+WqWksrQxg8XRoDSnR
LDs8rgP+xTAN9ra9VqCBiOe1RxXuimNIimem5Y9TuNQa89001coh3WIkmhgi
zXWnn2JsI+j456I1G6njBpi8VrfujbKXXbTw7Y7e14sySkMlIYjWL/QWEHK6
prKA6uyvIxoUamBjZOdXw6zw48N5SORhDBTmzDAieJC8QvJrcdFyxHzHoJDJ
eSec/spvEvPeiJz0P6/B0QHmVanQW88JhBWellZ7lAXps593qeAUrug0o/Ed
zwLwlcYk3s2RxHfCjnGv39edt2EIMKpg75ajlsCEOjG1Ubh73rJrRwcNbCjA
ajHmotH0gBOfDvNYsfQ7yC92GGNxnYddjw0Huk24CCPQEsJrKWS5bDMdz9ot
wmp8pxfMNW/tQBYFjGEDop64nZ+UmK7SBk3ezFZ/Z2//ruJqfv4iTXlkxN29
2U61TLKwjbDPfoR8T1Z7ufKI2V4QKnNO+EB01qCUOj7kI1L62f0pCHa7EQgb
V6xRQt3zmyDxpcAJjE4wSQn+HGw+xtmMTML/8G08YaAvGoy0UltGiSWWd32d
ib6W3H4+mH7VavxMFflBzQcX4m0YeZQtLDPYZyOwMXseZ7vcmj796WhHoIs8
w7fs7/Xpe2Vt/cB3gk06js255EFycD6HWPREiemcG7aO9wbiumfFsaCPu6i1
tiWpOl1tdZRluaQeb9ejvCrpdBQeNsatEAQdrCezfv0JsOZemRnk8I4fiQeQ
MG4zA1PESEgPJOndGZEgbYq/pzUcU79w+rWAjvKZ/6b2meXv1jVPgxEIvsLA
tBG//YO2fBY6m9bEcy0FBaSJsiN3qxj8y11KKvhMqneAKyPjy9BEwm8wzw6j
vtMrEF1MU8e9ERYFT3JzUrfzcp8tTIQRIgzpxO/XFTTNDnfpMhn3BMhqQw26
IiYpsLPDJli/EzWBI5bwurF2D290Uc8H6D01NuK2HZ7BHcToO5S4lFVx9neW
LigmjCNjRCMecmwIZqSfRfUvlEVLjy8RTfnWFCXjXamrWgCiHHa6jJb9bCQ+
zf332NSj3zMqNh+ouhX3zhVmgMS8lx78kBirYUCPkbN0whbXG8F432WpYgqz
vHMSAJryFsh0dqkY0kIAL7nW3ZOg61RQltqALWNJC6vvYU5Rfemx2ycgQMQx
9U4b29lRocRiUB5iR7EUAdhXeOjbVvQ2ik9qzcPy/BJlVc9DdYG3IMSt+YCm
TKXmc6seuXlQb4UE2eyLREBEYVTjBl3jh8ZvWUneW1zG902kJ0QQDIdhcNzS
UDCkcjnbaTruJzOI16naaF3PtuyM7cGWfq6WF9VVIX99vyyHadOG+d0sKSI2
/w5dPt6956wShVRv+V2R20ZCemUmmt9cVhkzzU+1sCuyZOcWiVlKi31mfqmh
cqb7WamdmD/mBtHi4jvghi4E3l8r8Bri2f2aOKd25Bb4lnngt+5LrTlWHyTP
GFoC2Am0J/Td7ywZgA2u+s20baSwdT8qYzJYghhU15NxL23KKRkfITx5tOcT
S7s31OJD7c+QhRnrHvcUjtC91qh0S6VCdtJkfPFQaUivUNsKj4+IoTkGFLJh
FkcnBGivKPO/7oxhoQk2D4O3Y1Nf1F50Nu6U1wxFASo4izEb5ZTSziRJVAL2
Q7bz1FZAlbVnWF90s0y3vH2nQtGPTjEmchbTe7kRhlYGE9Wtnnz9KzPrWKkT
mHmcFBSyOQfbcfpcAyjRoCzDcWRGxbXjmy7MJt1cd6gsKOtVGPfvFBEFDeZ4
Re4KK2YDmDJN6aa7vU3MJrVqDrCNLN2BhCndH2bUUBie75uBoEWedpbKGnSV
9pFbD1c73UuwkMh1Ydyk4QdiIHKTO4hmSNWOzI9OSQF0rqGXWEIRRPUP7+wN
27zvpmwR/DhL3sHjc88g1g1XiFTawL2ANGASRV/GXSFi25spwwERZb/SIw3R
Y8/leE9DchUD3EEjXhJ/9FO5Ga7paDM+4fIW77TTgk+rIt49JJXEPzroVLDq
zSBtObYtbypUmtX50aPrKXD2Fwi6rLy3/+3zezUeR8M/7HvuUVaocQaoqdvD
GnZCGolWpoLZM0MFBTKEdoyRPaphjz5WUEB4B3OvB+pcmSa4Si55JIQL10Vz
GAYrptGvKIRtevYNx27ePSZZnphjdJWwgbXSj6eg4+ZHgYujDZigTpNcKTuQ
m/LdIkpCHrbUZ47ab7VwDZK1fJ78Kjz7l+vLHG8y5+xcaLFV1pKYOIxR9iau
KvRscG7Xxza5DchGXPcDvnH4+B+jIe2ceTHnsl6VtMbBFnIsCzI/0AC2mg5o
UkzwtrzYorS+SlC0zc2xsBrzmQeDkIhl9UvpiJtCFupqYrz1PWj4jHal75gE
P5FdroorjWzqwfJxYCtgiBvKEQ/L2LPOPPrwIEYtYrGpxUjSZ7ioZN3yDYnp
KmV8jz5dd8rNsHXwfApkncKk8cm1zNliFCXdTzVqHhjcxW4oTGJQaOSnX/8Z
QG/5s3BEXs5K30N4RhI7VxVhG6Ala6lnixrJKjk42OmasFU8OfNUXc+/m74f
Tr9iIOv8Vlxzd7rtmXtFUY18NSr0BkMtJeGF1TnwMcshR0Vw2CKlYrN8HS02
LSO774pa0WYVW0Inwcwu6dw/CTkwZ9yZSYpsh1BPenRZu98ufcu7K7hIrvgM
iql736r7nlR2rgfXLKR2fi677txGivr2rhXXmBzLI7tX7k164ByUJ+Fx5Nro
wbw45mtpixM6gpV7qQF+WkCnwi7Wz+G/jNUG51nNjKuoRXP4miNH6LpSBnUS
zjXtticifP5Dxp5sXpi6bi0+pr1KsVWmcCmOm1jI7a4sqcCyhX5M9fUoiMWQ
Q9flULePaEXTYYAGKAhmHscl4obVEaGBnriwtsLpmVPlwCiUH6M/Q8Pir2rC
xHU6aMKKmCa8NH4vcqBElHC2tHCV4u5wb8I2yU3vsC5nPhnu+VO5fftWw2Bq
L5/9CbuwX3X4P6IFjSCNxO9Ud5oJQJvkBhZTJXtWyTmteaYvDIqCopVm4dpx
1tAjzTkxEMJlwN3SR3XvEihAr60pVRUtrlJ477jlMZC44GF2MHwKlzBSrIUg
+1byjUUgCr47Xc9hAdSh4IElMX9WkNJMA57b1UaE+2bPDsb2iDIQ+03cTvvj
FWpinjRfrrmv3GagotSuyH9A3yu7etHpAfSrjnmLSi3wWv12iHhIIc2c5SUZ
IzK2wzb3Q9NH/rAVtLSKBL9gYzKF7r8TT/sTwqG/MzsHQsQ1a5tYtC+uupKe
h3q0lcBXpaIMeWXjdpwzbl4V2sS9IeFAxXnveqBGoROTys2avFStzajMK/mU
vrHAFzVWJmfl/1MTgXZhYQ3OO6QQRoWOKkXaIGgS39IeZR+QbmqDQSCBTbBj
rPEc4gm3OI5mNGoxQa8fX0JFOqi+H3sKYSu4Nl3MqGzJlGd28nDQ9sjRbKTK
qP3eTgu6MM4uNzgzfrfelzA9n9ZxL0sI6c1RtAoGJ0w+jDEDdr6hszC/PQmE
m+aurFW3f3CAtCCdJ8rN25yCZZ+A4wBwGGdpGYKiEuMEUBM9CXbXPlvkW0gt
fCrBRvoKy4JHS5fym2N8vIeov+lIzGBcPliSfLFHKMYGBGqVcnDtOI0f/8YR
oZXpPsMRyfxnkbxK3Du3W9tqH1fBLPYbfIuy3tRABsK/mk+P2CoHvTjJ4KE9
GkH1zOb0xJf4oiuuCq+YSKiEUNdep6gyroQ1okOV3zgqnzT8ITb+RZkL5J5K
qaT+ITBhA+1v/Vi9+lpEg8vALyz/khcao8coUGjueSY5TkCECuEtDWVkqNjb
blJ7GOxnAkTfAk63EqjjshCc6nCwrNi3HSLcjj4ulaYmPuRfwyUJdMyxvRFm
eDWFrUC25ST3JTWZ0junKblHEYzbnMKIdSaR7z8C6j1iyZUa7wQXp3m11T6D
4/DEbxKiZHbCCov7aWSqqBU7e1eAxAKzlI0eaugEYn+h065fOwyq9U6+7GPW
kre7lsRqjPvbOvN98bPsYFUoGvw7kpK9WNVv1iofOV0Kb/3GhthHwJIy7kBT
ldIJGTjS8DRCpQYzoJcPSLuPN+BmPLDcLs7+5sL98yzAAc2dwFPlwIe9qjrp
9dIYxpciJhZ6lZIdUwhDq3qjmK7C+b6ca5l/WBWhbxg4LJgke3S48t4qbEDO
8/Z7mf61pTwITe2JCUnP6Lc6VTUhxcud2C986+xy2wkjUX+SiWns98wl/Fim
zTXbQ6RU40EOI4uORql2AIATNyEO5+wzroVyFQBxzzQUHZrKFcLHYXJrAsM0
TtWAvbzwy3YHB/sJH2Jt1eHekzr7BR9oGVIV/MhFuU3eprissu7b68HxuEKR
YZwHJr44VAp2kAabMH/1dSsyVJ4QWuVsCQ8Cv+nqFKawNboF8ZOjZxqyMk+E
aZsgbaL/QF3s+EFPNxFIYwCrSHvStoGTtFEfeEOv2sU7Oioh9gw9m+814A0P
no9AJHywMV/eXtszX9czuVxosRF9JOazc7OjhtpRrpfukMh0Kw1aFzcc6dJv
2o59kvDd84x1bPFo/CmIzrKLmV1DtL2LQZnwcobRifNw8pf3MnRQUd50li5f
CO40e/QZRRn4Akai8qv9ox3jS/LVS9n07AzXLsB/iyCr2HPGMq5MqbQ+Kw/G
WTkKYr7pMzC4CSKsrv9l8qOG17ND4YzCcGzm0mdYjLPbiBDLMZHfcKHfNqjc
RR1khz/NPCGbwwgPFvKTbQHTuueo6Nwbmcqc0N4xp9zX2byDBrn8wXo/iTEW
Q29Ve9shGMuYZZbG6KF11H154z/DF6XNCZ8sHbET5vMVYjWkYOqAYiCTHZ2q
UaE9wuxf41JC7wR5g19yquM8EqT/ng0QpMJ+9KN8xaQo8V4Ndze2ugUi7/TD
6zdXwmd8+cOWPXc9Sa8pbH1MSPd+VNDc+Ix2oscffBSj1wtt0fYl/RaKghcm
z8Kj/OpUHsixPaKkB9xrwy0PEOTPyiz3Uz1B+C9GrTFCIaA1C84z1Zq2Z/Z9
m2VkZwqXmelgLGUA8FIpKLplyykEdAtynbrcNO7L/yI4c6ZCSUdxEOUk9d4a
mf6XDoDsPtQBksmH+6X+vK4tT6g5unUMx6G0Oxy/iOoVcTMgpudRrPVHgYsO
t/3KJQi43I9LZPEkMbKsw6iOQQmz152YWdUzQReF1X0kWjfyOlSJEQvmAtt7
pT/FZpkCE3AX12cZn5E82/lfE/oiOqODtZtn1wbO1WAoVTIwjWOoWqi2uTeG
075uSaGACyYti5bANHxFta4M9awnRPByIcFb1e64RCboUthoG6JBd5JWlPnj
rEm7IDK55Z+4zre9jMp5z8PppyfI+GYKx/QyX6dM08p2PloQOxg0R/DXVx/L
+9eHWdVVTOibyUvnD1yQZRzCK1oChrC0XFRZ745iNg/AZA9aZjNvSQ4MW54q
RjVOBgm4G0wsYO6ig/DrLPjMntUlQkE2L28d5+XciPNTbf0DgoLHzoTz7Ntc
MyP0onmy2PZ1Mmn8j7LymM/OK4qxuWPHJRboZczTBViNfSnP90JX0x71vdlF
h9ohb8BGcLvozPipGzc1Gm3ZQOIKwumelDyBPkESMAcgrrIs2yj27pkIE99u
qDb6neZ526aQ7nYJdP1nJAA8nIJnLZbk3OigyaSvQ2yoF5bHR3a7Ni/SmRX3
pW5BRxXGZjU0f6QK/gGGjBrMlB+ROvy7ia2pmdMC8pX7xfJZLhZNCrx4Vlci
lbNl5DKPmJ3Dff4g3AHiJ1HNIwvnx6SU+Uq4AJP3Agq6Rht62b0yqHSEvI1U
GrZKJyOrHmEa5tScbRjL7MBPW5MWcfqr0I8obdmisw3b8QA+FaZPk3xuvPLC
JNDtiDwXFtzj/x2/UDQMB46y+xOzah33EJbktB1VVRFmHIriYTvegjj4i/uY
XoQZz37wJRMtO0hXAaPY0LziLus3xPCjGf6sw63QAk0aOxEb1QkMGqGrFRak
2bzZ7lugrY/u0p2RWGWIHosPYvxxgPQZKQL5fqaJ0MEA5OIbfyuw+0wtLpSV
40AkftqwkPNN/s4zKGKeYSD9gDgT0GMtACoVhVTr4CNXBE/Sp5s4N7ihAXia
dBLiQlTlRXSWDNVcokGvHtEvS2eYXdoicJu+mgMfQTtHp4K6Gt6vigc+blkv
mzaTINnyF6LzVe+v94RtB9MF/WwyYsK9Gc7f0gXk5wZyyrFPnbtCLC0futkc
8EUEfTCteFKs+o6qRqUIYeH/qJT2WJ61YdCDgjSihaPxuy3NhYNej7LngB+7
+zDMwCg4Ad1yQ30JfvVa6lx5av+0AkXc4Faz5jDiICDB5mgi71VK58CknGcL
nNpstOR4o1tHjjqIGq+TYXL653SW4SuBq3Cn8I5Je3D9Q3VLm12OF12oMcR8
H/q/OuqHYvKVsYcGZpVX+5F/Xj1gYvaIjw0pfPnoaUBY5k7QfLApQ9ljeepe
TNc6slKezr4WGco0QHuL0bI+nMA07UQDfMxLIyQzwqnwzAFv1VvpVd1uUNwv
37auzIUG7h86vWNUy5iDJQKKrdA16kBPyWe8iWMziAPyeAEe6iAXNyPWDcXc
NNAEZuDpP4eNDBXWCTNfyJ8vMqvhTcRhNY84/j6NCHH8ZGN7u+tuKMjOrXBF
UrhcHyfbo3osmeSDBhjtOQXtHSXib7S0+YGSv92BxNk0LwDSEbFh80nFpLH3
z/Wlec2vYVizmlFBeowa9QgvpNYYiJYqdk5RRq0OSa2V8eU15NxV4ewyx/B6
O42dlCN7Sj/b/QNbvc/NIXyn+ZZmpt+DH7A81aVouxZJOI5jkcSYm9xwPxJe
tKkw6B3IRT0IX6fTDfEfFYs5Dk+UxAxLEtWnzGehnWrphNqiNifWVheFjYfo
FH9ET3JShReJlbUrRjY4sROcGlOJX/jzCjQgomSQ487gzL+38+fzUSqOA1TF
7Scrk4wZAy4sFXMOyCLZQzy+6IPAfdLjYbDje15eyWVVm/wrSVk+Np2CXOUf
xN/vrSkCqOXKmrC5aKsUz0aUOGM3Iy0bhVvqNpoqE5cKjUAAKp8Qo6/0ZM4Y
wzEmL7mIWU5zXMZGQ8I7fCUocSGigV8e7crELMMVtyzYb46mc+VSUciFKe5/
RaB/jMZTSIJyXEvNUrV9Yp1zjGjrH4Dod/VHLccyyQgo6O8fOKko5F7VPIDg
Uc6dySnIQ0b+Wnss7YAmf1cCKFwKPrQC79q8sja69+yno7jqFfl+lJx2lGLv
EzK1apW1lfvIzMx58lWlG+4kj7luBsYAhh/fvLQ/hbtZF0T5LEdTevvOadfj
fhEgEBInjAyzQNZmqz/Xjl3ZXYf/hilKVW+NdjMCgxjuyC33FtAYBCyPsdoR
ZagQgRCpxWSEwwiojZnUqeBszB6UO5Y2GD/8vIoqlZJLZNUMyQRPy0I4pXd6
Qk1w27WLi3JSQQRqb4v/XVMH1qnjFXyUAGbUK0rqIfxOvAbZMOULNkTtaqjy
eNtMKVdgrQOQb6PA9F/ndjw/WjTrzWO/UKnEaYdAoFMXb/HstuyVI9FGksmx
pOJYO8+oiHLnAO+n6AedHalAe5kTtqOrLPSEc895J+5hV1lapF5KKhac8qyT
ezL3dBqALfPXddcSbsyWSS4J+NtEaAGEcC7IeUyx+Ng/8iHXccy83mWGvCLi
FwKZ24naIVPTxLDoGPgAY5+KgrLticUAK69pfU2/XDER6sI2cuiC8joaxRp9
l7NUsy3Qm80e/28VQknJ0UkfPLAmJ8olAHFcqC5aKoCi3eIxxc0f7V99GM8A
EqaKrI9IViQnb3xQbLL5Rr4v0bW7EtyswsRKojMmxadBrTujYm9rYS4zbR7+
2WE6WUivoSn1tSU7CR0uM9PLAalVS5sNcD292B7khpb9Iin91vfJcsPSwsrK
NhcWWEL4XiCSTvfFBLCU6BCsyvk5yM8SAh3UwsJHUPb8WdqdrujgraxHVKRx
XfLz30sOFkYFxxklzUBudwUn1v1lLZZCP7xsmJFmNiMQV8U1Za9rH+8ZLqPG
+DtksB4MUO1kXpq8c2SMCnO+7ovoaYLAX7pOSyCtY5VDsPv1CNjgWn3BUD8/
mDhqFJvU5gR+uWwxe4EaoMBzYneiUiMexV29V/kfIup1FijH7z9tEuqAnwCF
F7v/ZFdqwQFOBl0YXw7vlpn/zyaU9CyOVwxeTe4rq+FB4IcBpgFHJMwPtg6A
Kp+VQwfuzF8pAKHbjSELRuhpplBiRZaIl+zUMImIDUghXK3Tj/2wGCzOTWMX
O7PqeFRJpH75nBPA3UQ7ofymlp/6WXSQlzBkYys/Yq7REVXv2BtLXKwELbz1
rCZel/d5KyxgPrpum0Um94fPAkJHeSOsfaPKfDsUI9lWpTGPScWSTbr3lafI
GiKC8xFKuWZDMN80pYRn6dybufnRrs/A4Hh4N6YHf2uNBQhaQ/k/vMKN28Ll
QQZywllzPQb13MTXpMiNUzqH2DAfrai932cbiJWkFsRPw/YlLdNRURTr/MVG
HkwJJ3V+9z5FxWssrqKt5gfwiLjNMD14IcFNp0ubUNaF1rqe7nRtutmgOYOg
7e+GL+ypMXambzLrunmZgOG+K6ftwDPXvOVExyxFGUqwqWgmSfkQ2Rw2Tgu5
codhJVcar3xu1zLPv9WuvQDLyaZEzbTIfDC36wL+KJGR65fnN95NKkcM4hjm
CDhrirAUQrGzyqnYISYUXwlBx0CPLybMqiVM19/p3DpMoZOf8SCr8tZx82lv
NRo867obH0BOcl20gfarR9Bc27keeMBJmJ7BNH0B7JJF7ChL8c7sKfijF3xM
Yga8NmJy1d7GQSFU++rXM8l1i3oL0Sj7pa0v+L9Q91KhE1H2O1rbfzGWgT6d
BQ3AguS71xx7sgThsZ0GCIFsPJ3e44dxkBwKqQtw/4wQOaiTJQUrxEoMyL57
C47Zv2jqdSaZhmhiag0/19uzNK9f5AcCPvpXW1zVDxN4GL8jgYQlbgdfCQ6p
HqrrWXnZLobDBuyb9dG991Ovyl/yGmrPo3qj8f0Jwq9m59pbS2ZY11Xv7aWE
RSg4hSxj7grzvBESqz0wTWZltqPWrf961AZ6RT2vN1cdClYfpFNLXv+2xzfo
GRtSQRPolDMKNTgWX3W/4AXxcaSCBtxu0Vy7jBr6XXpE5FKRVSnxdQbojnl3
Lp2Fv7xFkD5M5aVz0bUlWZbea6lt7hchswRR4lRXK+wRL66OUq2/Zer9bD5Q
+YOPVJMhStTgQQHs6lwmxvtkE+pdTw7jyWt4UJjJnAgzDgo7LykrQ39S6cCD
NUWWKncpQ9UhoUXTZWvCJSvAlnlHqYiKMEYldr4HEjUeoxGqS1ANL1Cf2ZgQ
0ZMAUFbd24XI9v4jliQmK+GcsVkXWl62jfmHth3tXhcV7tY4q0JL6KiUwrQE
cFF2J1OHBf38S5Oo9+8NTRmjU6V983t2RPbdcFifISw6W5xfvwNFARuVYLRv
3AWhXerEM7Wdr2lWxxAASzFObyyZgriG1lkOqaoleq1VkoxBS0Nw7pyfey4N
UFuGjC7YELMDOJifKHzYAv+g0HVbARWvYXkv6qscwuMT1TW097pntakAhF9Z
MGY5YlMMQgaEdoztzN0MyJNmpIHgbmWBSU6xLlq2rPygafputqPLgEdBAh3g
r1f2AWj4G8pCDgabMiRZI0hD2x7Ln1z9Z6JC4WP46WBuiFnPtUKqT7V8FAcp
hh2YtnSj8GPHwuD6avUgdLJolrfqElBTJN+gVPgUbYTMCysvUNqaDfdErovY
NxlWRPggXnHaJ2lvTfi1rBdRRegs0xzUZiL3R7g9Cmz/W+yh1yC4xTeGCLLH
7axzK243yP28Td0hgpWdPS6otirjO8AnQ93YP5aue+G6+f2xuKNvYkOqKS6i
lpG4FfwO3Iet2y56z8M3NdEOEcrqUx3/TTMuiKG3ab0KPL6P92lOoXLtXKSa
b2D6o7po65hzQp0DONKMSVaOZzZFMZNkEqjLqluXEv6sPhMrqDxwoFycDNO6
DHCEYHaKh8p6SGN4iVTzgkkLClT3Mfzv+Pp+boNYS23e3oSIDMf6q9DijRkk
2bjm8LWR1wqeE3JC5Ki8WtAl2Slf6EcJ3BL1SFml1NjIlct3nY4uCYzOEDnp
vKws6keTYPkAd88f6q8eLrL4+sXX1U1yrN7VP1aXiO+tVYqO7XwoXV+l+/8v
+SCL00KQHJ9DM21/7ammD0N0bozi+DN0iVFUoMgNSBteGOGZKJApCR2RUMkU
TcGo7CuXgvjeQHFpICyOfGQZxZbUknhzVnmEqJP/yN8ejQsH4QkuIuBYW8Wm
83AEzCTT+DalLDOdqetdLTqX3bXgpB09cQqnNRLXgZAxr+Kp/CCKJ7Nfh8Fp
Y6EqmNgXSaUXDQ/3g2Et7ajlFmP5p8RWw0yqMRlPkZ3bdHbh2zPbYj00HspZ
i9KmrC+siKOFRIzH5YmggPHjr9Ka3vaHwjsmVx5bQspiYiO6FFQxIwCJgESe
AUKmt71rxWLOYkAGyWCOLrfONLpacQmk1Vk8Fpm3SHybmr4dN11PsiwZLcy5
EXR2Hr1D2V+MudCv1/YXtyCrcEx7/+fef75Z26e7jeiNNSapb4EjnVa0qfFo
2JZT1E0XWjBqphUT1tvqBENcWGH0EB0R/KbeBTSeJ5xK+KpihaQdeCbdKLdq
ZJIoK/B3XKpTHNQZmQUb1M6HNaA9WoKkjcsLeC4WrlLzP577+WMYFr9b2bzB
yonuVHe5lqWTA4aIYu9D9+M6jgq4GTpKt1Q/+WIPg9LpFbQ3Lqnghf6qKyyo
nahNRKY1x2PWDooksm8W5ITU3suv6qUeV6Ehwyy6n+1IAREscFXyffh+lsfc
Cv7a+QnnamCVtF641c8X5u5dNfKPVl1pef2WqfsScaooBhy8Xtgjtk3KM+Gh
qrUjGbjAdPrUMcTJ8QnRRsjwBXQM6mNUhj34EbN+dd/mg8EBQOWSlYrkVwxp
23MD5FivE4Bf13n12bfqFfhU8Y3hjhaR/mFQSIXqkP/mIkXWVa8Bj8CABHoN
R6r2P7PIvT2qSrBIUnus64nPRPnBJsiCkX6fm/DCyLk2UXi3GIXG8RIP08D4
CBM1dAAb8f4y/kWaRcK6XWr2GLILOKg9WgFTjt1JvqoW/Qf1qvXi+NsPz9r8
1AA9r6WfqiyZB5SOr+a2roFVmx3pVrJMsbldVxrRkDS6Fgfd82w/vNujDPBO
9LWM7PyGAtlFC+EeNDzgNj3J7YkcYNCkACaxP+IHXeRd14dXLP63LLazTzB5
U0YYpwI2BcgmMS2DR8Ddof4a+OnjkTrIgRdIyvkn+wxRq81F7/6wt8V0hQI2
MCl9ALi0D8iyWh1pzyIv1uGQ5dBN0sbuH8RPekH4hV3xP6shVc3+rawCPHuH
bUyBr+M0U8YcaKiFOHQZp+Tsu45hRgHGYTYIVMntkcJ2sES9dSu1m+CWVe2X
b6VA5pi0DI9CQFvN2aB/Wi89UnvXUqblUlcCVHox+gBBpmHdz5CwRj8lTfvp
o0OVw087coOpd3pn5ZP8q6GJPXb4G/sger8Icv6vnjoGnRsop9VJ5psAo0k0
fLINwdmVJCq2SoHWu2lyRD2RNckqwfoXhT/Ktok8cwkNnC4+HSHuPJMmMiTH
CSQtETGZ9V9CiADtqNhkl3XHEkWs18AJbfAe7p5uBSJ3P3Ig/ZbASioHcN8Q
05qH6i9MSfF5TTwcZVKwfY394g+KDoZGmELamKf7LDqcAQpURyrUzjXbImfR
Lace1oaH6iv9WZzZCK7H2ZHa6zcxjAdGIi2Siy6MoikhN9xnQnM4Pu8+aZDn
S0JFk3PACl0WDsq94RPxTgqRGl6YN2jm3LepnyZjOpevCkBUrqurOaEGfew+
VmlXNVqSEpZHZEXar+MEMBg6jLKrrOIET1oqBaQiDo/6M3JMN53tC2BL6DqC
F4EkDTLwI2/lTYZaDxVpz+GJgXt5A+AxEwbfhwI8zUbi7CibeJ4rTqYqVQ/J
g7w4fqFSoFs5AGfD87HRaQZP/1wQzyxyq41j7aoZ2d7bTYrnYuBxAfRvSZ9F
TeveGLSvY39p1jpb4Lwn/si5PVTTB8Vxw3kYUPvaNEuNT2rCORbwTXiiFkn9
cE/rxSatb5WDGYZ4ugHUbuwaoqY6wIVtgWg7nVGftfyVhxBNvtcxoZ2B/xX7
Ycjuoj3IMl7CKlVpmcQdkwVT9SsPkglFCUAgtGQt1IYSAG/u6vldYFp7N3hg
rQjbnLtDYIQ8AF2bS9lS47uyyX7rrgENDWaZjTU9kIYJTpbQ9yxCZHHG2zVr
R45RA427RUawTdSgigYUiNFgX9rB9+uHEyIc/qKAU4jxlJpCQymZ65a1L+SR
h6Ks8WkbGeRhg1d/hs1F59ngRGgcF2Zp4Y+ps8FRPNXdz9g7bzIBSxTk7H17
K2eqJaqTbgA9K0+ptTVUD3fK3gYYMMQoiLsCrRCthomJ03HrnOp54GxeHh7b
/5WRiL4D7yigqBvUcbEVXAt/N7m7cm0QsKM4Pjii72jsacexbrNCFeSu0m9f
BMuJQ/9TfvNaQwcB+QpVAVzBhe6nKBCIrI0vDsiScgo2Sw3Vvx/K5Nnj7kCI
fCsyYEqzt8EDe9+nKhReFSUu6VZvFsjly26PLqiQHkVwVz/HlbLVnXfNH5IZ
WMMgnH/ChuMEqZrAssXndDJb7diyht6nmj0+ilHY5jbSxic8oIuU+vNr9dDA
nGSSE6dMZ7zxR3BVS9um8xhCSsiSTl0IDSPNblCa4jMcZOLV/U5n2qIqqVmD
3Of2FPhaSSpaOY6QeFL/sN2fLaqJeaTZuEMls32XYrWyRVGy795NeJzJcZY+
u6rEPXSiuZTJaXG7swr6iirwr7kHTdG1YLnA6Ces7fSP4O3M4PdgKoVhoyNP
p0Mlt8fyqfK75nV3OHqlYuATnkGQtYMqq3LaL7Hsl8GzS7dH0oRTRvsfz992
YIJeeCAy7B57ERSL64A+f/BfMsX3iM9jaIOSK+NupRnz/S+rxrsGEFQq0gzb
hAOXq8Xus7pxr3TeZj6eLvSn8UFlcbzflmXnCndldqMpp0/OcQ4poOwHLaow
xBPX/afZgNfP+ENMiULA0CtGCUUhaAK9hfIyxeSa2jdxCnRMsFmlGBjlLr3S
j6cGCodtpwM7vyxnqbXx3Y21P58ruUhiZhY+DPkUdIr/k6bAEcOjFEl1Ybs8
GOT+/yRSLhYqmESk+5GnsWw+PQ7O3jFWOuIpnbc9ojskigNswCjU9+DQswv+
z02/Jonj4nTRFZH3hEpzzehB6JMyQVZiXc6HxDA0Wqfcnf6/FRmQKfsI6AQ4
9+zK/vG58em8l1FmhtHG+EJ8Tf/wMKBKGiWI+dRYu+839zK6ZHSuFqGXUnHq
lV8/sQPYzJNI6TKRamBZzb8wvVk3/qvfEFj1/YIlJCuirrhg6I4KZqKYLe7Q
CuEJ1a43ztKcy2pjFgPX9Uw6xhehwIGAtZjD5QKVjY7cA5AzqdMQ2AAueLlJ
GVzBdxswgHgKaA2GYMFXxOQjo6IiVJ4p4qR9D311Bq+G6HVxSLr3yL8odDZx
KWICGOVNrgE2MAyHlMEBWN9IaysrcjOu0Vl/EIlXMUa8qUqMm1TyJ4/xLRsi
bcufQ3PgH+xm92/n19lXOVEGA2tVElU8BpKddB1/ABvNYY2IHP70gpWTQBzK
uwL56sf0qvHbVPjMMCSwoMd/0mY4hJjxqA93oO2ESf6jdjC60lqSYZeW/Wo/
FyfLxDjipGxO55CxU/a8Df9zYN/tQNbwQboXs4GynSWUd/qgOU1IS7RQLeeO
C6LN5UV0JUza3RF1D872xHmuUDmSWr6E3srl9YeSMoToLnxzB0XOeJ5yeMvA
rbJkh6NEcUghpQYgnTzBLAYCVj5L4MRDTbdLnYRizOE2f+xTZ4DlAbn/zWOJ
TgSmn7enfkHNKD3JETTac6MP4wW3FlQV9JJ21JcyKJkRMC8zvy/U8X1gFtJd
dr4pxcka08gq9NAP9CjmexlYQP13RdOe+SknDGFVBWQHvzMx/Yyj7u1QxJdv
410b8OMJloT+h97zjzF0McVCaCG+vPQ6bHS//cb7XXy2xiWY1oiv851eoueA
TpS90DoTqePTILUYOd4F0gLnw62aANNZbkbGIwcK9c3swHYXhnNcaaa+KTfP
zpFhlvc9NjM2nChS+6iPlhoded5jtaWsChHbvKfM+HSpS9S7SSNGw1uyRLna
ugZs4UrTMwpMVa05p+KnDjke2Lopv0VWsqoiGvqIT5RvY+zS83sXnHNnKbqD
QoXiFWppvqN7gKg74HGi++BD3e4tXLJhpmnxYy7xPkXfrGh2VvFaRwJjwkfg
nSNBLW7UoVflJq0V2AIIpwnZMA7HGln00hwTb+XErQeVnHyuSL4Mn5soaV0W
gG/UTHkoVclOvyp8CJWNRxQY1EG8uoAyM7Gvg8nWDRKkO9nqVSi55KIda1BW
BfFpyGNeHOhbASfvhRbX2MoaoYuZ1cad4GzxDNHwKihlkFV+hQO8TUsjFpzf
kf1cmzCoN7qHZYdj7qOzUL1crnGHb64okDRW8vepPh34blvRP14kCKoEjm64
U+5ln4uU9TcQtyiFs/n3ANY/l+seYYA0UmlnTMT8FSNbA/qF2WWaEiiLLJkd
r/5vgTUbn4oD8C17+tXqItYAAgJPu1VosUjOnr3krjSROUqUrpkfU02zs0kq
mKLOvw/UWcB9LjY5cLIdymrD92uKYAEE4EYlqTLedcyC814KBFCDVgPdMySH
1dKMg+jotJN6t2mOu9O8vQbVepFDugRSPAL23w2hK0ZF87Rt5hkL3w0y9Uog
kL0R6EFWJETF04xNHFhLICgVcEz0tp1sy+5tgYLhoy/WmGJIws9C5V18EL0g
S6xHX0/n0oY9EnkGS3TcHPUzTiDJco6dfRW3LPTdsz3oHuxes1/UUAS0YYar
ZxxfoittUDyKp+1frXcMPW8oRM1cPqkAAZs1H1ToV3OTdDqVzeA8OI/AZgwj
2YL/08WYqKiaI/EZyng6aGbNNPWbbj71fyjNWe3udpaq5qiMLnU39XGYcjAI
OhzeLdUsvI3dvdfPezRqiJ+4EN0O8DENde/TQl4LYhw6fO0EYKJ1+SI1vNHY
eNcEP6ptvLvFwetMxzRa9FdY5ZtQRv20ZEHkI1FAbk/RWZKd8RbkfHY3Osyg
PhB0aCb9rpjuaPXJMch86ZWMZrMlR+Wx+HYT0iEjQ0CUUo5N7piY98PxNKoa
LkgR8otE2juJ7nRwnsGDxEl1Q4LoYSe704lpL7eIDL/tHK+oY4G9ggriPGmA
WDv+oUUnNX7zlIdW5WEumzuLyCM7XmksRdQTYfJ77If64BTlVLDd7GQBhlm0
gdizUwa1DCXCwp+K8nudlXvNKDLohWCT/7YHbvkbH6o9OTA3pEqZbm11s6Bo
x3N/xary4Xt+a5gvkEkzDcEM5lpZhoNgJTzZ7c8HFDzfzl6rVdrOefXfydMf
QDVD2annz2I51GS/1H9QrIVByYAUgWS7QuPfj5lonXNYX6W4yAfDQjKxzLEF
Jmu01pQQIjXV7VYfw5H8HsSmjbdic6VDMkqCsXGQ+k30TMAl/tXpEY//ivN/
QL5Ya87sZb2rsrPr60hmwFfd22a3x+4LQLeAM9OZJ5IIUPF2DVv37Ld7Y38W
tfRMJO71RFPUb7UCYQ5xF1LnU2Zv+idh5NyPyDVCXK6WJt8YftPLMwVziJUO
ebn2e4XD/Gv5j2Ez5QNkPpIM/z6Syit9ZUJKVL6Ds8LRjqMPfq4ijC2Wsjjr
pkjLrLihty8OjNRnF/42oHLkmU5wexf6rVT4uBdKMAo+yQHhYzpeJ4S0MFcd
ZUgmpOeQYWHrG3se/jcTl8vdmde91z7szAoin1hLN4Vofw47WUhJSFa4mqmD
3AIAPR4eSCdsefxJOcF27V/fGEvBzbUhr+GHp3QbwUoOK9o2bmCpjd5+a+ce
6iLKIH5iDFVqu6URh3Qdge7AZazjGSEJ0xNr4Ya0tEMZ+Ryi1n7Wl/xdW6n5
9BCZFb6ZaJ34BBYKQ0fUfvKI9wICFAi2fli5zi7+xd5AInt34zVJwFkCe1jW
dHjmF6/zYneeHfzGdLNGIl24Z4z55SAPVp5nVPZ53wzTNLEVF4kABUomWDJL
bnJEmlFFu9HgcPn69WmtrBsKtIsWHERY4I1G8RbassOm7TfFOMFemQbVfj2j
j0qml6Nar7C7CH5+CkItmnOA/hDkMgSxojwzylBA3XXLRqGJvbY1hCNjED1a
fxaBhtE3eFl0rf/fB3OPlMgbeDSjrYo+xUy3mx/IFCURWrqtaXvCnxTEcdLo
OC4Ob2ScSGLTKIcsjobJXPmN2aD/hU2x7bKM55AXdMDGiqdOLyjFuyM6xFFQ
SUqCSpKD7JOcTTZdNhYlIyMsRePmO0U8W4ruTRBuLutg26f1WJn8kk7rk7aE
CHEXSvYZwzQDH8QmxSq6IW9+wD5mHfmLb8jn8ueNlpyDLdB3NOFbei8ssaXk
W5xB1a1Dx7T4tQhrm44c6wj9Dyg7EOg/4BCdyX4b6ljmal7wDG2YDbA0KML+
9+Gi1IC48kh43V+qdgC6urLtznCdpHDBFyJbjfRAJsJors33AwjJ3wnsYZ0H
fYX9lJnN0G8AdThkvN1eRGU40epgNn3xkNs+biJc/ImzMw9If7k7e8J6W+ai
lbKXvid8hqLdergW8vx+oi2FBB6TjaWHBX7/d9ucWpDExnD1+ccAlZPVboLX
9OqJoL4kTRsuXD1M+dSK9BU0NXpnCzC89aNqA9Bp7WfaYPjlCwLBvulE8hWM
wiTyTKVZpeiIpnkpFYL2n8z3bmg47BL95byAPlrP4HSe6AlOr+ttiKBJdMce
gNLsUIRZNU2U9dkqINwH2xZ+4oWNQRZrxPS/YO/rHWNXb4m2n6XsG7H4ZTy9
be2y+HKjfr0wxXI1AVyoy8kJw93jJgQKtiFH5q69LHbhF8VnP2RvwwmlE3Nv
qanFmqNWB+gTDHWSKeZmwWQq61SJHbfHe4rLrLZwosrknKoWSBt1ILSzv0fW
3mmG9kFNxPYdju1C6aEMDNZPFTB1vOxT2JeutTb/k2R5l8jMx6B8mFrILRho
1d2SVs+vc158l7JCgtF9fEBkopboPCtFcZsYTWID7kI4KfE2d39lDdWfeAm4
BJNpOKITkI/lin1G0Pr6GBftXW5gEsRcD5t35phvrb6YGec52z6kFMpZUXWq
i1Z1pnRdpH8IdABEwpkBQ3wLowrOZWQ/kPipwDEHXp+q6vc/M1rLQVeW3zvr
JN2zwmBfmYGRCPB1VeXEKLiw62rZC9P2KXjsP6BtwCGDv2TybqGSQiHwmYbv
C/ebVlilmOCK/iUNxsXGcWVjwlKrurhMx70U3y8ZK5KzLfuEUGJXe+O67zlo
miwNPcY9ihkgXodPT30NgwSrjyjwb0zV5H/d/85lZXNoAAtza11q/X5EF3qd
JQQRmBrEKTgTe5pOzpJrYvPMtqx8uTT/NYHh+OVg6B4aFysNnZAQsbW1lb3u
eVBWq7hgTy1YtTV572uPN0t0sgrlNWdoIo+3XPqwnVxUjNJ91d+D73mDmy3d
ZUa8QOtiY7PoSP1OGhx896zXPYEsu8XR6Gkqm2zEXJqawU8YsV/TerGQp0o8
ZlW+aSKC7kThqHgyAlTGiriXWxTJz6yN3ANavc3YX3FiNSLW/u5UwaMx0YpD
VMA+9l3eLRhFaZhDfKgHk18Q5HXvY3Cgq61wGgbZX5zUjIQwKb1ub/Hrx4fX
CLUkjaEO1Wg7Hb+TXL2AO4aPnDv0/olwm6xguzHDbJ81q+s0yr2sov8w6A3m
r9Lmw5lj61KD8X9Lg5WAzIhdniutkPBvA8pDkVpOR0VuEmPrcs0pPLjrXdVl
Ew8BC0EgPi1HXRJNrz6HBTH3oC1NTszUDUe9vAGpm2E8yqYhNus8YuO29nKL
h5qd/aM/YWhhPiQfJt41dx0m1orS3flDQkfujIh0Fqv4YRXMYVpcpsi80HC3
Yk2U67SIcESsEdG9/OiHm3vVyAXABs3NaGk7HnnS4u+o4avJtfvQLD/gIsL3
pRiVabf3Dy4xjV2jesGrrCI76fnX1BS5kuE0Baw06VCOpw2wpYnyB5FXD2mm
i4GCIv/tCZ8UIGk96yFXOk3ycIiorU2V+XP1u0+Kt7xjXwebqtsKrAdwrwKr
okk4lEkCCLo6a6PLL0BREoZAGGgVuMMWGrUEx/lBg7q3du/PfI1tSs7KLVTx
QPSjPrhOeGk05C0mI2L9BggIGHRxVCj7meN5nDA+4oVIHeOJr8SQjAzC7rMp
nl0/f9gmn5LvYoxQhWBqbkD0P7SRe7w2VsFgTJfD7ykcawu4vSPA6El5iiQB
TC61Q92MU0gEI1tM5OCONFKV9pqmCfvDLRan3rFk88m1kFCcUFCSscgLP3tf
ypvQJeSzLciRQ0fz5LB3f75BHxatC9kASsNdQP27IYGrN29F5OXCl1jAeH5P
E6VdJcWDDLan9a3Km5QmmOFg2xAJw5r7Va+1VI8SNEkJXJW1a5wyj+jZ82PT
Tk0hM27cMTMuD8v9feBZ6p/F0FYO3A5U7MkuJqB0PuO+XI0MB8RduorcODk1
cblGnQjPUk5d9O3WDpY81yxpyUqaEtviTuHdJfN4/6/x7IM5eTcjrH5I6LAY
6atu5nsQ7pzkZ6y0eDX5oPVtBpvPoutaLIURSq4p9l1iuDbRA+K6yA/fQ2UB
WP8x0ZAjfjLsK9CanXLi1ZyvBVzwla2+ZCoHP2Q+7vZp7FVsmAwT3Udolm8X
2AAHzrTEGNb3g8mWLm+xMVK6962BSua8QjUf50fNLGLqjg92kwAmuiwm/EKp
fFgd35FAbGoxwjkqN/9nxdSWmU1RuvPFTZIWFD7Haqra9FhV1JuogO5lf3z5
c300qQW0pyeAYQMKMnHfAthIUASku/G5CSAvdQIToEF9rgZWOF+e1RrnMVXh
tUNDDVYcsAUXfruPoIfPufkBnt+nzhyuifiBu1FWlSBDgjseA83fISJlvz8M
QU4ZLkkyRFgUO00otw7oVr0/y9TqdNOg2THV6VABfPlHaWY0VLR/qGax4iGJ
b73zNb2WPQH/jimEnLNhhw39VDYV21fqZ+DnCI6pdAo1F3JHXukqOdFNn3Ao
QtBhMsiCdj4CQk1xbLNgoVwH/+NZjW12UcVZJawkrjxZGW76JGfJDnDV99uz
mwc50A6z1u90WxQlxPjG3O6YKXmYd8SZgWn1KoIeDnEMQWcG0UJ6D4R1SwKK
0NtNanWvmYYTvTHD0u0EUNSqnJzvtlxgQWjXPbXmsd3SKh4kqHZCfLompCaP
GI0pRqpTRtTKCSSOV/8GdcOpMQj/nKteTsf0BEaTmBporT8XdGtwbMEw6FDa
ijk2IsmBUsTJuiLwAw1VJU0SfxX5qxceTn58YXcFwaOP9N4VWbxAkPdJbe3g
XKAtmcz7CWeIbaBf3Q3CNIRK6ZDuXWGtOlld4ShCGfKTfawkR5i8F5TheYxM
tPu95l7js3K+JtOhzlWdot04WkMyVWNtrlBLSfy6cB7ICebiv8sUb2bGnMw7
bhM7vMZ8fHAFvH2mS6qXj0GSrxBoXCQfwZTDWq36dK+b0OBavO7lPDznnYdG
1qdB4SN7FKvjqiPzdqnHSjFRahCRV0txnLYiERjWYCf+X3gDsufvE9gcGZnL
g9SdP9DJeYuyVYKYTGYzDO+GOWEdVN/K1iVMcjqZ9HUmisTK6ywxPA8e0+gv
NdM5ciwH3vd2Bh/YupH3luEBTEv4r2vOI9BHtOW5SCZKPIh8QmDLZcJ2DzuX
BmrjYKlhB8yNctsaIZs5xPve/+Zcn82oH2PKrGp8dpqAGoXvrYcLBixwURiV
aTAubPuESBZlcxigBhI9fUE9xUX9fPepAilra3sy5EScAdjAyBfn+eP52PgP
DoTiDyCgKdUrnv2+rs1nkeK2Q6IcXpeZxKYQ6ar80WRSh2z1GPcjMc+f2K95
ljPGAfWaZSdbbe7HJ7I4c0+xoYF/gqDhi+qdBA3NFBM3GrrXuFrughBorjdG
vXid/dXPF21kRtvwgdoC2TIkX+K96Yh17lFokQ3rlOY66wRLWKxVfnJujXva
WpB9zUHy78oskmw+/r0MnXHpF8lSJf6frc3QdbNMkGYH6W3gUPiOp7rM/lpW
v8YdRqIloennX736yO12v1FD+YYC2qL4+X5AvENceEMo400Y3LqonE7PGvmU
+8PTMFBzLWHSIBs3JqoRhnR4zYvRAKDrE+I9eHtvvV7H9N5Xk1I1eBRXSOyd
gSRMGCWOiCPJ0tTjixpyk8x6B/5z1f+OTXB4mG0IiFo4dAvZsIyVUXZfjtTd
vr0kjB8z8JH2g/Gc1qJsdwwYt4zp55kH08V5pJeYuEnWjv3F/c202KebqlR0
0BCIhpjq8XO/u1LwCyZPE0ntn2jsqQQWiSt2gMK5V7jZ6ICZ6sgPJMYJzD0+
yve7wrLivl8SFkuwRgEGMu1dVq/UQ0LnM9N0mFq136fe3uptQ8cLsu26vXMz
1ZmV/PFHS17GPP2BfjDIIkp9s1ud0rzsvTvyiBtizgcPwlnU0K7YQ9xGDnBJ
HkDFhS4eT5UXaWiEh7Nx5u3UbHYBTxs2yqG1OsMp38OoDljLySs+fDBRjc45
9bCaXGyCcTip4W9VNW+JcLRQkc8Jazh6GOUF4pYS976NTBQEWpAjWtHILD9L
E/obtSTJ1/JCf9ISdqz5pVNA+CB26Ke7ibLOoC2byFjJGRCZyiUU4XueUh2J
SNij9MF+fgZArl/lVXlRQHV+NwWU5XoqcsVuLH9+RJkMNIfDKV5cAcJ3369z
HOoy2qjDI5p3c7c3Bze5nwrnzLLXQLDsqpBN5RZwryKMU8ugKkAS/ALuMhX/
4Xum5bDfNv7Q+8cqcAhAJADJbj5+S+ShxpNVTQrqoThKOrg1tVU4JNJa8xiK
tD4iJD9bhJkjueTRcSByoCkBTaDU77mBf+ZFZwgNcM4kaqiULa6GfgCdpUa/
xVIZaZRnfiSmc+fjHicY8w5B1MDrAYVocoDFN4ubpQ0xA7A2HAlM4CQv0sRk
u2cxWNZ0qo5EEQBsw+oDoTmtU2k04xLCNyDmjGcqmqRHc7BdiE+6hmjLQlIC
I0l3SR8u5SSNLeWDF92Ml6HZ+GAUWqXGmR1nbh2ytUBaSgMJj4/IStGkXfXV
SFO6ZpsVnkKSeuqslsqQlgzJeHriSIEU0NrFQUX/ap7XzfKq2O3/simqi116
Joeaq/+nTvknPhSNBx4u9wJ2dogZvMPsZJchVo0F8N65bv+7s/Yh5BjzLphY
ae7sOb6vWES8kjOP45LalClhkAaL7pMbwpPQTZjCaNLkD0bbFYIbt/L3oIkw
BdRWLddB3IfyEEjCPvMdmn2ArO75XB4mcDcWkkB1+o6d9LSMABXu09BCYH18
FMPFHuuL/PYtJ+95n4GcYAezHVVUsa6NywjDoJORkG/reUDZQTteyjeRJSWU
F/QvZeE4DC728c4HdfkuSbJONY7bfHqXYvx7qLYeQmHWUNjCoU1EghAPikfo
/NSE4UObKHBRRCAjMcFkkr4Mqa0r/FYvARvMrY7HdLRqvv0CVYrAMYWrNaAD
B1S73My1huHX+FjAkud6YSGbsoE7nra5q7QOfkZQBzZDCVrGGJOptjlBgy+E
skY8/Le0NE2PNLafmXfBxWG+Qosn0htdrxbnxulg3oNbskPvNu23GzLSCuI8
6SPxVZMRv8yjVEVzt4c86ttoh6hVd1cSaxWyxxBImttzzKgwIeNCOi/sbx2X
2Su9wflWbvEsNets/j0JhlhFoBV1Jx41p8a/aJ5MD9uZEICw3KEM0UvFLaB0
DUL8frUFC0RKK8COY1vEdAshbJo6YmSynNSBzXXx5j+thvgTAo89LaMLn6/H
5NrAlZ9Hp5Fi1U4fekzC7ZDpe0sBmwzhDp/fGbxLhocza3erBLLn2znDBwtV
Sqj799JeGHU0UJSJSLpMxz8kID5yezKlLP0ntiJF9s4ehj4RsfAVyxTrue5X
nyOenF4o9nYdf4ecK+s+XUeADecO9ilXsymGCvv6jVjLEvLg88TgQsEQgLVt
NUDstu0y1ic6+BtfXAPRz/gJGMUw7NvWZPgDgIKS6EhrA7Bcj0wsTA+vsld8
hONkrBX5c6IIMs3MQxx5yyjQt4JXm2rPNjFiOQHKqHLGX/2zSyLhfUrD46Ne
BpfbYN8GKLUribntKLPfX3weOtBpYVLFUt16NF2+V8SWXZBNFjHTLdIzi4t/
ddIUSpThq1PzTTWE5Eue5hV0J4fPafwsk66TSLQKyfua5HK/poZXdEtmHWEl
nb5XKsc+vqkgr7vWWLkkiN4rQU7SReGLwb+z87cCMM2Qe+vXnpSj6jLU08KA
ZrhxwFOJ5KmNpNMnAM+Q5G9SUnwSCcHqvFv1yESu5qrYMAnUnUTXMhtgOEpF
/AlvM8NRI0vqy7QFVlCRf+J4t12Bh660K4n8DiB/5YREgutuIxIt28k2WZcY
Thl9yKg6sEXdh4hzuaRtlO0fWaKa0km7KaSulkPjuSpVkC9w+oUyA6TJp7vG
ax9Zt88vC5tk9++ecXEzDqPi8qGG+1SH0wh1ZpF+rVIkzfzsHURFJWdJ7oKv
GMAh1Q6YcwJWdkECYeqXHWFz7/w9JnerbTGnNglfxARLFSYHExERW3oJpgjn
e57qPuZjuvPaZ1dbl+yTRqHgpG5UBcO44OGIcpqKv/XpzCAYucgEchf7z9Kc
2fbubnS1pUmQ2H7j7s3DxuHSrts31Xgw9twYkZ1xXQHYoJR/Mt76x/DDTmvD
uKGAcKFXEVcZ3B2BrOs6xJRiUtBhEzBmvlTuC39hn8jzjCBnsVE3lFv7gEhC
bo5HS1z+v4p1AIX5t5WPbXgYR3EhOYW31XPZK2ev6Qf4ZISMNO3zdykJkvR8
i4Fm6TFvk59+rgSsube5XRf0b0qIH0yCUQNNN62wnRQDnyRUnAjzztZFVRpz
vnbVqeJH3DTQ/gjVIuLOobs6wYbFnJFuemdSNkpkLTrttmzkmb8zZsNdXB9P
XfTEBYsSKg+F7e+9PMhQ+GeCnyOnOejonJjNFoMhFK7oilDaNVhSFfK3KHyB
kY28rHnLVJp1raz3R6MDVtAy7nizRv9a2QC2h+MpY99q2JHZroTBMIjqUlFA
7CmSS14xKolYhW9Ka1tDMvHIOQpiurxomv0z+QjDBdMZo7YjoqCc0NOaSoL1
WC18jtkNRzz+UcmE04Rary9eYre8C9TivaQGKQsjSTiyEag5TIrD36SBGF2b
uVERvih2CCplbJSpnj/9mlwZJmCwDLHNjYKJ9Qs+Qng2fmltc7UxkJ4iXuhn
3n9ixa7so3Mts5UW4pVC80OFTs0tJkt7ajWT4fHBBcJFenCcVVyRcCY3XlJc
fpnwCRkJu7RePyjqW1ZDZwM0MwP4QergObfM2DY28bPfhezELQwnOPSfKS8n
RjMaxPzWGQYiLubC/GEizhhaAwloSK1qnu0+CmG0b5Pmx7CtdGnnZ1qE7NeU
QprN5vuUsi7I0hEsOGc+YWx6/mYIcovPnspwX9WG6RErCgaWTX1LSQ8GZY1P
WnoRJ8aBKR++DM2QgXWlFe0tT9/SDuk8bLijB/AmTDQ2N2qoM7r1sYwaQu8H
FBNQbDbTvlpWCBOC6pTaW4hyig7Z6Mpzi4VFdpLbqx92WzzmvWoCjCAr6G/y
T93jzkMhRPoX7N5kuts+uHdDNObdPz7RxiS79UkfjCAphzpB2FwT0wEiDcO7
pBiU09WPR+HatvgYeHb8dm5/BqvLBZRj0wkL6garqAVxRiUco7AkzKtrVggy
cqNi3aHZm8xchtoPa7XWMcFecp+tQSPLn1wg7PXPKNZWyN1UIThGtN/X1K/m
K8eNmur/d9NeT8+ogjjv34YZam2MeodBfEWiYkqIPuToXxgjNLCFK/lKW2R6
1g3DO7UXbfVSHszSwiy01rc4pWFxoB0jfH06AlrixvVc95cedFLijWRvOCC4
4CHinY6Ym8qrQA1iLlIN2leLDHT5Rc37lhG1GftX9B+N4boVV42UE78WXMHQ
snHiJ8kXTCKLI7837OiYY7l4i3uWBFV1l6rO4T24WuVTOHTUfpb2UIkRPfNI
71+vrqPafnk5eMkCguh33Zksud2ENADqR63IbwIx+GxL/QL6ymlGv7jr/tgY
U8PMY1st4Tftb55QuxFf+eznozPEYBA9eFzjwpLWyLgXacrtKCOenB9r5erF
ysPtRk4OtRYMX+8O4BF09wPJdsAu8tOAj4LMTaBFIED0Omwiwfo25YRCOq/n
OpdEXu5T0p0WL9d/BQZyZyZG4FhFbjfxLkBvaZ0554YwTLfKi8zUc+cRZuFw
mAPfp9ldqEgf6aTUYXm3CrXjfrlXB1WjoQatbcIr8jnGyVKu0A4QUGfN5xAJ
hP62KeIQcXlEuLPS7KAaAEJAmXrptJJPhxZXgmf1MRcbmSanPswBKl578i5b
f6vqGyTJwKBlqbiBEYmBain99GnrTyLZXxefvetRlrQdQBvAo+oIaZ737CQT
IhhuEBBiKQE7LcfNpT6TPwQxIKL5uUKS5DgcOL3K7NeRTCJt6ksKDyAL4rYE
evmHav3VKawQv7eIWS8QX2seZdMrIPBgYKUeVzAN5FZHXT5BODA61T2gpYRM
zbRJFq2KPI/Ew1/1mKVtMDHvBPLw+YKbTTAByLDIIaq1L6ykHTCbO9tQiE5Z
BWkhSRAAStTepkXIVvzEFjSeh7P+uYvBk+G2+G8Ou62MVgpcNcHiN9L16MW5
54EqNC191NciNpd3k57EK+lPOnWHQr0rKI2/8WDHodIoMYTjUuUsT/0a27sU
tM0P6V9Az6T64jh/VpoPGFlybRCEJBSLZDhGapASus+8uc5/kUMO8zdFoaco
FxB5X3jQzbqlLNFeyr9vGb1yfcabx66MQugcVREnOnBVZ5ICfmZ7NrnK97d+
4B24f+Nf8vNXvAsTVlKXxXAJOur61eUYb/2+oZdwybVKCQc4HW16lJKc93d3
aCzwsY/PRNPSA/IONG0+5mXsUCH8MED7EZQjE23+47vx19yAdHHpmCfII/6E
PF2fuZMp6aL7Y4HToJioiTIjJv/TNmGGIEP6tj0asAoquoPwBwA/8F8JX4z8
zh6EGIrDd8mTUD6aZc5hq2CH2p8XSe8aRTCknBGBl4ptfvoCu3YdKoyF7DR3
zEiMVFeCXIJQbPGM7fXX8Ym1Tj9J7tjuJGDsPkfoDXuiOM474Hlekrso7/Gt
RhBd3luuIGS1bwYJr8iob0S+KXQNpCGsyI57MeOPE5Ay0l4GV7l98yV/b4Px
0N8tw07WS+8eymelScY08HT77jaTLlsZMzM/LU8mSlQbU3MRpQqAD289tEB8
Oezz3rGNMGqrygbjfgUDQPMRX+foL0ZxfZA88yz92xt9zWylelS0aeil+cPx
FJoj/QKUxb+9dme+7nrb9RBEkkHo9WYvEe0z0pC/v8bdVPWe+Exn0i278/K2
4Px9GaOLNjStR+3cMFFCo08B5xTNzLb5Qxi1Ug2KDJ9QyyEZc4mEijrUebwq
oAEHgv0doH9hvLR6MmUdkaEWCDBtoWGD+dz2miKh9+5HqfpxYsHAnV9QrluJ
kvXqAWYzqNzVsYNQKBvRRZ270GsTtqPvk41F/+XQ+ofssj6dATkJctlSBEwP
rorDtnN9axYUxffE8kUrbEJvlIQ4sBYLVXRY6c1RlFkZK0ZFpV0iqbfrKUMK
0rrcb+nIeykfeeHcEVkIAnR10RElDHyaCXSSQijnegOcSloljwmNYWMTtLSy
xV9zzAYbqWqfTjSMJEZnOHkRkSh3+oYNvjyGKPORqwyWF+H613N0nqZQfvkC
2yUuAFpEHI4Zo3V5U+GDz1XIBzwewzMLtTbs1rrcTqUKnFhdYPiIf/OEjbwE
CcLegiMGiBx34I/+YR+QUiPrXvAJcve4XUFw1J/tBRxBOgbDzKDd4gHkytNU
QjI+R0g0HJwJ2tqXvkBDWNtzYqLr9Lny/1LTBTFOPNe1A2/OuJxJUWug9Dgu
MNlGv0L5E/b7w/EVdcPMA8fQzh3X8R2vh+/aAChLenEDNWHUV2J+ViZ9LEIo
/FtmGTuZUrktLlF0EYxglUDFapPrhZjOnDbDO01/K3vJ1fKslFzEhSfUQY0Q
f4UGGAaecwvO4AAnwjinDW8k8LJxsVGNCh0W3X0XnN2z8dqV+wPJq7IBMZsY
Ki0SCFJy2Ak8wCQ5Ea6N8g7B9npFcVBD+otKRTun7yZJmLjkawoF6oWKp/W7
Ol/HKiIcn2yWntJzCXnC7t7l1y3/R/uh+1FGrzeg3NLQfbIOOmGz8jo+kdoB
P2Kf0t4rQ8qEtmSdKbFD1tblo8ZGR9Vy8y1l3i3MWybe5quZNsWPCQbEtgGr
snkJy3A8iWJcrTw6PNSg1qFykB9rNCTpt/B8RzSfTNE8fUniggv2YpX2TvH7
0+CS4kXOyIuSxU+En74fzmnpaD4nHP6cBem4G6NFT6QOjFxVc2J4MoQ0D5yF
DDTgUg0n1jQu92rnYkuBMZjm+zK9z6FlkODFeNyYgAZVDs/421RY+FJuzFwn
Ju7C8c+1IF73QcCmjt7l7mhxaCqwW+QFpjxCH1sg/KzqR3423Ymi8mavFq/W
Oql4r9pYfuggm06+Vl3qbLFjVkpN/roRJLF1jjf/ft3lQpB5UP3SRkp2QvlZ
vx+TrXLAPTyDQG7ecigOW+saVaixQi//UzX72OTZgicmOSup3kh+DzFFx42q
1zzYUzMGcMe32JaheFjGPTgapiQZHhjZREUtkeGDr9r2mBT/mqXmonWO91Gk
zNGLLJHRkCgrBkZpu2XB4dUDEiQbDh34bNmA6VPh7FuwsnxCeFSpTa7SSjl5
EvbWa1au6fajM0r5K0UrRb7CsftUGjN4r/CrKvzBKNPcoskGebTWez/xO0Yh
zrnq5ENxkkl3WxDDj9bpKTKv4BoGYh6GNjD/wGIVFbi36gLn9Q09MirlZPra
VeXPsIEvgoAU61ms/szKXXqw4G5q3Sz+RFYI0wnULjt64p4cIe9swvkQyRN2
jUHlrV+g33jgpXXJAifnbd7OOFoR0aFDfFFersvc+88XV/beCJ5mIfQIgLPE
95zLU4lE5mX36ZbpezE/XJgaqKo63ekfb+aV/+9H81oUfBKnDyQGiD65Xajb
CSstZuqjtqPl9W7U5FBkN85wrm2Ftaa/lwwph6XHS0MBKdxkcLQkv0ij6NBa
vp0d31FLEyaLpQ2VNg0EFibj0XPC2c3jgNs42NSICod7jr479JEqwlxFDEfM
qbE8HuOjqqlV6PRQMXU+oP+v7myPpm0oX8EEMqDWjEWosTP+XsEQKbtJUG6u
AkI6Pr1KWchsf0I79Ng5hRScvN/izVLo/TNzMw4sO7EJU7SibK641aYK10z8
P5bLxJQAFXgxqCKW2MPzwEbES2rjKKQOC3BWdDkvMpI3Q5qTeS7KFG/feUMl
XxCDj+51vrfBr0OwSV6CpgpmOkNVsWlMLaujgvr/VlD41Hp3/rLqNmC4Xg1x
oQC8kp9UCZa5sYe2Djo39oKFsTodrLrgVPa/hGhFf7bLqn3b8nlLz3sAVy+l
bBbBAEch2MVWXjqaM7OBQMisKcrybTZdSOUrg1dKrsDPgNrYNIBJ544c7Xwg
lnzCgQjpyOE8Uc4yz1DQjz85sSd9PgEpC3bnw/4u01/g2GOW4HoYY1pMvdDO
aBetc3cxYfYdDAzR0hpA1VVQLxx2u1LtJjfXIgeuvWdu8fZJQ1VnPueHHqB7
XMLdSoUJo6JxT66W8GNSa69JXwOhJ1WXaEaBspT/2d143JRz3d4KlHX/v/Q8
PWd2zydrbYZ53qCP0G4zpu9n7bHquoVTHjEG5ORXHQPMiRoCsUe5b5NaTx6r
kJ2GVDbUmeXKeE6bYADBmj5w4UTZxeZ3YI82cAK51IuZNVjkaFkbne8vkrtg
I/d7fLFCU1jWl/Ty697z4YT1EVAxoclVTer/qKR6bCn0JXbsNXOQnk16Xjkd
1rNLBRlHfUH9z/RVB/q4ZsewYqztEiLix7nUfYY5thwFmjU3BmGtNWKaIXD+
GHMuYKFGmI2ck2RE29obblCWSeg0aK2qxDPkq93GrqV7bv55R78ESsF+oiCq
HF6C9PXh/p/VE5wsGtv6VI1xTrVvTB+6TM3p3F9xszdEsSNCalo0hugcEJob
ElFMQbSiIW+1kaSzN9LfTvydcSjDAfiSs8pRfKUYelo3oXAiXP5s49HlE88w
neafvvnwIs5vuEnHvKS9rt92Zc1xCyJ5XXLXbvBZNS//H0lfPS20OcQrxGs7
cQuvlYj0swTHs1W8TNkW0P7yCLzjvL4OJoi1BfbrefkGQZSxikLK6o9uNF+x
N6KigFd0LGJts7uU3ftx5g5nHNr89UFS87+u5/2tw5F+NLpBK2hZnxf0IwwP
J9IdAUAyIQPoeIZN5NRvMYDW6JuYP7WCMYEOvy/IcfsBGgKNbFpqDjE2vOei
4XZKeJy263qrj6CpQ42RkOxe5X5BE5C4i/bm6q8P6GHELS91aNzU9HWvyB8G
H3yxkJgmZMvYeoSXcFR53vHxtRD7c3cZT+OKs71t8xh9keu5b/OGOq+OVmf5
QoTc2irCVuN8l5xFdyBec8X4lRmkZd4V3CR1D5dh7iWVNxdVA5rjmO5DO/zz
cBCkcsbZj96SSe4ZM6AJQIFO7DhGPmg+opkFz/lC8i7Gf/Q8yMtw3w/UDyRG
KgyMas/OOQ+/v/WzUhLiHwdKNPMZNsVCQX6g7NUmHe00KR4Zlkk7gbpWU7ZB
uB1sqlykPG0kR5OHkf4TuwyhfWfJU9hem+ngIqxhWqK+MVm0SsP75IVxOYrh
VjX9BrhGHGvnLErQ8itQ2BWhkoWjhIWIzHm11KKeb/bHAXbtkdTV+Bnrj/i3
YGlsJa5S8m5ZuUmT+X8bjP5AS0UkIMcs4S7IO+sv3wPnhuGW6FanPJL7jzV5
o4rDEYEGTGmPNUmXH71Z/kLJWYS+PvrX+lEMh6bOk3pH1Ojq7+SipgKlb4ga
KYxSE5DEdooDOKZ8311HjoFA5KtoXNAXyhbTh2aHprs0JiOqiEy2VdBao5wK
6q+xu6F0+7HV7mrWX4RDKj3uVReiRV3dmJPG3MxUjrFQPHo9mIdPGBF3KLSi
+nFrDEwG7ow8BVx7DG2SGEoJXdVh3m1mIDM/VreUeJWoNwW6lRmB6mlKMkaa
KpreTK4NgSDW0R6VM+u9U6OheAH6smMcoGhblvREzlQOB2GwFmrLcLY0ULX5
eAUVNSxgnzoO4r4meCqtS2KV/Qr6KbT49ujvAd2Z5mKeGSp/NPYKgIvS7mHi
0apf9IhKcux+0QHrpQBC9So6/N6mM9xuuxA35sJY73eR7NhpA1H95MtoEe+J
jsqT9+fMHedgju3osB+huctmsqw0FGZDb+A7OxeW7JaabKc15TDSHzJaWZmx
7JZl2i1eHxkzAsW0V+ncvfoMEwNleopguBhdrHtDk9qjgvY7IsLa1DHHtr8u
050HJaDQieC5zw9s7CgfM5wtxyZUm8eDAQmH8idnOY6JCxzcCl/7p58DnYvh
Z+SLUEqroJfexvifE9ZnrzQ/xMt3D8qjOdHdCqpN0DWlUtDvA7dE8Pwxjdp9
t900waPcW5l6exnM0/SS8r1SX3zOPjpwfXmDymEtyxoCjhuwSxlSksonkAPE
C2JjyajxmoKGzgs1SMgWr410WY2l7LkMjdUb8f7/0xkgrWqgQ7DFDnjXBqRT
QIzmCFLm2via+C+WJVwt6ksC1wUmL+zKVS82Ii51YPMg768S84ovUBGBSlLs
zQ5xdEOz0+lbHdUPJwsx4Is7o35LwVtGrJXadyGul9CuRlUQ+D27hGyyrTHy
kKOQXc5iWzLrOEsEibVy5S9I1Yesa8+FL3h3VcexLfrJ2Ezd3C1IeW88FW/e
gRBod9ayDq2vI+mbQZBgSfMNlngD25dOnE0KwKZvD8m2WsTPiFuJ+YsEetGy
uMI9Uc0dd0VNVCQGtfGOojH8+Ga6vGUVRk/VA8ML9bMX7FlD4UFnKvQki/qE
hPjth1+LMqpwCw52AMPUEfxFION+eqMXpJu73DEt1kfACqdT2/f+PzutCOsf
lSaJxsR1V/tvPTuryIlb3DTx2cqdc0IowFZqVIy/xNiNxfIhg95L7Y8Ul8k0
l09JCcumgT+C3nJPUTyXpHVGtMhXSVW10NGt+xyDJrBQ7zCb75hSgxDgfCx/
no8VRPOo7a5Y4QUojTz9jYuiqek4xyAJDPmI1ws+oH91xLGlfyFHZJKxWg8j
3XeE5iHjpxbHTBsyGZBPaRNVnFM3o/VA/OuuCt/oV6Md29+U4iwsjiUC1oJp
QevyQtdLWIWkK+enYloKqZ8zf3xqbuaL0XrfnRVMNRT0BrHlxVt8BBHE+K2a
8h8+fDWg+dkFmhqEbQBRO3kyWUJlfjUr615cHXSM3pgLDi2/Xv8z2rpu09T7
hABbqLaBQP5zmoWANKG0XRxVI12LShIrU1ITZVo3LARGXfjxqAsmH9/6uPvC
YPbp/65L08pqr9r6XnwLM5NbTiebFqbxOZcPkGLzxtJATvREcBN0eG0k9BoL
jRVItJ7yFIn7TSuBDigywWitLhusu5gNSt4vaLVQ0fTaw1gqMuloPf3BGkK6
KWsNRXVHRb7dP5H7sLYj1tjKiqNj8TGwCUo3YKqIC/+kXaS3RPigJnnBSpM2
R8j8w2cpDpjAJYZlMuZC32fU71FvdUICmDdqeV6M6ZPKn3TBRBblbqXP9XpQ
hUksW2v9jNoHZX+MOa5Q+znK+e3A5wDmMxSLA+YQm/d/eHsiHE41ZP9Clp5Z
nMdTanYeyxJHPZlrv98Yg9fN6XAkKutfrrMcXrpFwxRlYh7X0qEqwTB+Vtb1
l2hg9PtCg528o2aeB53fD/RdCS93qlh6ZxIKwtPWeaXE/5Tqc29+BdLydcgx
2fW4V5aIOTFe262yjKFKjJdo9Q75yfPUkFc4XUj6UhIp/uvNcTY1gBanX4yR
dvcFesgfjh1D4AW2s50rrvpQlKPl0EeAR77VNFhIMswbGkoKymIz4qajn5zl
Slmbbw1y/ahZFNVDtptKypcFNaulB9PgL6UuEPVa7YYBNr4/Id6zOG1YrYec
vbfyCVtCZnPrAZVm3NRPJ7vQ4k3WbMMeABmgzyaY8u3a3pmthQWqcplfIkEK
21XYreslep6l3EvWUEwSF7PCr6M31uV1h8JDom6vcT/xoaJTBPCCCGVsaPzi
916YwZ9aCaaDlyL3jB0um9hCzcmotB8SKtMw6q8tt8HHxNLQh8yePlXO+qh2
cm8ekgP2IFE5a/iVhMd0J/D/8adufyE82GSObaTFLksMfIAzB/Oag5OG/+6H
S5JF2GOdSZvqXbb35mA2JheWh/2GPzVlOOSipKnF0lAKMeU88Ja+jmeFvbJU
tM6GEZULFsZK9MnXINbsvpsIEJHEJNFgfMv1/3B/2rBhSSrI7YJ0NPd44PMk
2zI/SlR2u24p5K9oisNhZ7BTshvgf+A5NFDnPB5v0kPZSxoSPaX+HAjacm3P
UUljsgy+FROpt7odfPkPVoET0qUf+jqcsZva8Vf8WkIsEqvtMexcmgIh6HSY
w5fvhKyx/XVXp8UrE1aJ/rMOrUct10hvpoicYurRccLfAOh736KY5h6+xGMX
VfBwKSHgwPsaUKzcDBy87QvGp27PzI7BLtRHGiBke+0cN6M2kkiORHxVggiO
7aVd4K10HFHFNCA7VhhOshYN2DsUrjWBB3zYxuSV13gt4mDow9eIWYgFIIkh
77jDXx8H7oEN51C4Ytg+dfi6HvE3kNocIH06OF0F3Az6PlLBQkd4wPOLOiLg
HFPym+a82SAldJqRTW07bA0uUslZfcOtFKKnMBTgpCfllZ+l71VUwq/u9Bko
f9ICdoRgnkQgA+u4rTwlKP3IwMry9VbQl0/qHzIBgo6e9t9JsM+Rdn3P+uKW
iC96ENi8hxW4cedj7Pm51L5LNCS62ek3Ux6tEIN8OV1Nv2Dscq4so/C3/+TB
SLmaXnR066eC7VVPgn+Q5F9wHcNhK4MXkP8iXQrH365qdeBYZBE67Nd9DWVQ
VPYNmGtsKZqRHSrAdRe91Y1LMKdrnUVNp9IeSSBIgsrbUJ9wRi7MtP2ttxVO
7FFIplZ71tvf5Jxe/iD4FthJr7Cd2gIahd9m7LHU9xc9TD6MXrAcnqDkUeUu
NzrJQIiY5VfXQuHy4ihBeKgYcWbLbBDUcOhPu3qOxyEkd+gTjaohyeTZuNam
4yTBY/VXgVQvuGZsF1Rw15phI1iDA3LCyw4RiT03EPcXUhZQ1Kfo0jKHK9s6
jRbUXzW+5JvQhKlt4y4oOSpSFxhAvYQr6XcAVBKTKmlldQz+ZtMYTRAbBmXB
CD7obnJl9PnTkJci+aikFqHpj/tG6PW9AqTVXxlhzZDHp4RabOva7nXFTrIa
M2F3aZlarFmCJEIZxoo7GzERQUoOhiwgNE4+8az6fAiC1pNAfXRj7Vh26lXK
EOHYt+BaVChfjojp695JLTaPp7kuPEqiEFt7xLCf8zfaPgsRFIsEIXL5g4No
CoNPini4+g6SfNBKqP1r90R63EztLydMUCO69DKWUBzknJRCP5pUl1ZzM3U9
l8BBdsmVKdWXotTYPtdwrVWc6SKGs0PXWvvWX5Jd8Cd69Cr/4/yEB+21rIl/
cQHi8+KTP7NqJommeahyqeafZkKZ0tdy4Re8Q4CVo0WCxTJ9ikTguUhIGgKf
hcwdX5Vg02owNN/nYXv4DjbsUf8DdhpgPwI/SsWs06nwTTCPbiOR7zeZso2I
XNAxz40UhYJBTDvHQnajKqdSU8KUrtL01COsCIjaJKFhoQ5GojSx90DqEuMl
mvynXFm9oqG+3Q0LT5ftnrUkZxzWka1DNbqHiRdL4CMne6zHTzWAXIuKF1GD
k+9WHQuxX/l8dz/4qYCH/SspDzVB/1w70JfbLG0/O5wcSR6CvhGc4HZXkRPQ
113nNCel2+PljzsM2y8mbPCM7McPmr0tXasyF1w4S91RNmeCMzy7HN9fpfIN
5H05uc/8bnQJg9MfCqBVhjWXo8hbCOu3wtRIlkqC2btJH+urqHlfI0XTY8Qp
9YDMSMf0nSGtyIxDAXxydAyB/Pl75lZ43TdQRKjWo0rkdxRbwq1/a/hs0GBd
ogDaWuEgws/ti0EU40L1ot0vQmItv6jdrsQYEZCoO5ZGiP0iroMFVN2PYpXF
03RSS03M+LqqIbHwNsknRvjcpGA5Aqqq1RMBd6JaccTKeNb2KwzJ2KSry2ig
1PUBu5wr0KL6wUwjLt3A0FZD9rMqopaoL7QHBvPim9+SwyseEkTXQIzP0hS2
2ZamPCjU9Z5AwsKJmxBV0UI9rS7t1B3npDWBpDNBXip5X5qOlUPH5hg8rmpZ
fTNPWHXSfEHLroJF8xOW8h3LqRDGe6DpAMZvetvTPODnaEZF4BxeHG1HfCnw
ne1n6H4wxpESbgYRmNu5oxrvdHGPrHl5SLACsnnYUVU+HHWZT5UK4N16h8Xz
CyOTx+WdSbtqJfCf+WCZUJAY+YzNRgROiD0DQIFLyocaEhUNm1wzeYjYaqnJ
3LWoAyVef3PVpI0LiQX/+ivElrnx0n4x1HFbnoFTuKr5oPlpvQseSWDZCs3N
H+26HI4lefaeuFufDNl6XY0JZs6ts7G+lXwqxtMDf8gBleXGqnCr5CMmfqKK
C3iLS8U/A0gvjIgQw4pFp9YiN7cMADbhAtqzKWFGQd4hFcGjAF/Uk4C3Ifuk
ZmiTSw6rFG7sMeurBxaB/c01OdABZX6mOIQBzCbEbEFR///f5jHqYnmESVYP
LKYaDITAZ/XdVtSXAZUzba5A++xlpH/NpWF7xf84HMLWt2iY1SQCdLuSXljd
EHIp51wdRMXnKk2jj7TVL4CFMiIf3kN2C5eGmJ5CnhzJ3JqsfvkUNkBOgO2A
MDtWadWYmhbocrFijg3pHDhUa4kWzw6bctMYQ2k0cYlScE8VDR4IiLgj2O1f
yiED8l1l1dKD+3XdGUPE3B6Ew5QUorERG2NVlxLN4U8Ov5bR3TaVPSLbfx3X
LkCbs5T2LTFe2t4kOguCyXst0Sd9rKbgHhTnkwWZd2B/oo25Y28r8o4q1GR5
et0xP3SeW49ibUGObOxcg6XFs3Bt1Q3/xT/iSliV6g2SpDRsZ/q7jksKjtsc
VVhIvd4LBjHxvOQOwFCyhtkc55wfXCO2OrrN8XM0Vzi1zeXQ4yAqtn63xM8h
ts3ppcL9Py3NoCtSKSdowxwlhcQatzXlfZq1G1V5SAcNUuD1YwJk4Cv7zmvg
dA5DKL3vCHyne8DxO/Tubwz7Sq73henxV3K/vxJkP7yADJnlxT41iTo8u/Ih
WoHXOl9aS0qSs4RQXVI+ulR5r37tQ3nfhnUDKyu15yxrsW/bbvoyPg+dkDhh
I4ZVr7uXbzJfiGX8Bdpt/Dvf62FZj1P1SM2aFQkcbscnKkqWaKVQIJopuoIs
G2vs5vPh7efYhFEq562Gfk8wGHB7+GnslXULEeLfNADtVismb12xURD2otYW
8NR2aSgDc42bf9cU89XZs6iROqiFSYRIXauiBENG0kVlRN7nbh65H+A47i51
fBjm7Rkknnczne0KJMaZ3i2miCbVdZmQsYBAgfUq8HCjbXpkA2a2rdGXLY3S
1BRZNUoWOtF5w7PuY8qVgGE0Qlp8YE+iLFmePjcsswMqTf7Stdtu0tYs6DaA
8gaJDuzFOAWK3YQJ2uwx30yektIVc3qyy1lxRmt7wr/NI5N1pTuPXEjBB/ai
8tjVd3ISKuQPiCQSn2/ZLZnOVS+sJBF/Q/IkcDUxay6RbQm7RpSNrzIh99/E
YDOs3smQKwRqumd0Lq6HzkHfhR3u688sJ4R5AIzVc83fejwH7tCm3rJ4ZAJy
RNwvpUHSssCXsDufUNoY3hXCyO5p1FFzxlS3TYnkxBqA9WNxcn6T52wQJAsS
FeKIhNnPxvef6KAzbRbzfulo1uyduURh5IUYGIMShpI9HBBR094u3AvW/t+z
phwQydWBnkGHSfhqP1V+iRQEdDCPflxgOtPWTBsyxC822dAc6N5SI547bs50
6PV8S2GubbciJpAdAYsfaIx5T9Nkgj12UzX7Ixl5C+E8icEiIsUrSw4JPw3/
egEbPUgnBwJN35vaTro5seeL9KQ6XbPbm/FV25BCAlky5M47cHXXQkuk9ze2
waut8JSfZ55XUMvNQ7MH24Bak6g9fQiOafDOoYUkX2F6Vg0uA36lLfe5XYsq
C/4J2BzU3+u8p005v38vdY5NMj2rLOJqnCN4NA68tSVnIgFRkHxEWxsyk9N0
LxxMu/QNoSfHGjswB1zrynCb6uV1bEWOuq3NAXblATj6VQXIUySGJdi5cAxU
/wnUz/lA+Ka8pni1AFn94FRN3oZ4XXpo0y+y0nwYVNas4eALpUlvylvJrciM
5PI8TrzgAM+XUlRgPxLh4rB54ZrDq3/uyzZUzq3D6uOx8Zz5OdLIfM/vnExn
A4ax9faRtVnfyZFkt6REiyVaP0LBx3cV+mzb1lQRXzWkq7fHvt2eKgrxLpfF
9+BFXZpNtkpLmOFmV7fOylWSFUlkPs1ETcbim157ImXU9ubz5130A3Xx4Rr4
023Aqb59/mMXPyn/mnIDrs2x1C3A+LIUHVYAjo4/0Y8bkTicDrruNHcjqgN0
a5noErpwvhqpbQdJ8BiH9SOL9mT0y2Qq/AdJIdRPSilhMM4n4sXKQjlofjLQ
ui6iakEWzAZAn4Z8Sj9PYGdeulhzEITbi368NJtmRLy2bIzP5eGVd16+Uf/B
WPY8b++IUaCeysqv1A0PHzt8xM8BBs+c5dBbrwhidVHyXHLTMHgqP0mgypdJ
saT0lB7cGE5/BqbqcSrUXuzqLpBVvCiC7vTsgbQyqipcpy7OFJ4qCFjbBHsh
gx3JyyfdpRAp1nr5AeYVs4aDY74EYBXqFyboef0rU9wBawMLqHmKwIx1mBRh
iiOG6peFkrVOLkhD7C0YyTXTMAI0by6IUWe79j4FUPxpHhIAGD1plu5QFatr
EEVII/MRritJnEpaeW2Zn2cLYM41+qZ/jZf6p2y8yMzDMmyngOxgQVlqgZh2
0ohl6I1Q9zECphzgZnCxa0O6jP8l3ljy14mvvCUgZxPsaPuWbxGD5R4APLnh
XIw7pesOje6NWgtZN0E+4xOKBCy4ArmPuALovKndT1JVEIDc+6aDT8bvq09L
ghpLsb08npsZg1ep7eA9UhlInU66eC2LLtntcrOlL4J6NecSuIQfP7oMkTvi
zqWFqtG3ZtiasRZUM07jj9KrcI6QGzhuUzmXUOBDncb908jS8BWIXjL90LCX
u4AqfanGjQ1fLGxSfGmm1mOHkay1VtNUD333rfU00wJuacFN9S39aLIzil5M
pIsoz1FUAN/9FxbgzxeKaLfc9hI1lrOoY/sLJ+wBgPELPFwbP7Z86wDgybk+
hNAYT+HN+7ajkXyjsyVpWZqN5yAG5W2kCo3jV+HTHBWaN4JN5WNvKbUBUqj/
0t2aTwMogrQShGGds+2MYIp/5sW2eAfrklbRvQ/wRHkaLtOcfSRxh0DoCQUZ
dAUBDO1n/UvhzUTSkJxdU133xkZV6osuUFhCgk0YMaBX+mua0mgeumD/tht2
PLwvvh3uXeSyNcleC4eCMXLCABdHZA2ZGZrsrYysxGN6oFMK8fmoQ4ZLvAJj
v1YvrjBFI4gBCp4kqekI5z1E2wxz6+8PgBuCHtNR7Ltpc3XAws4BpUG3pgts
HeXCJ316lKW6GJdVYXSd/4o/IfpkaHVA2jYtr+CwY6fRTZvcF8mr2fpx8P++
WsdAo4tYFN9NfztHKqSO3/RO+6HDPWPJKHBtisCsp+pdITy0qkWJEGic3dsv
O6L0RGLRan/IAKOtN0+89pZQ3CxqAygavJJogbJUbcjvJGMjpLYbzDfLHB96
YUWFHtJDdWPzLckM46ECE/RHWLqsTa8MJN9BXpSD8uS5M6vOXpaMEU/KDGoi
TtshOtB0gk1E+e7R1WnfpB6XijIupsBfak6pnRVn3PsJVaMtsG0Hi7eq2Wrq
to3svgRSJyA26fzt9+gu1BOfAiaJUulT7D1HmbYAJVip3blMQZEksrGxu2rx
yJ+FnhUA/0hskDWEGIlV05EQI9ZYOXCAUBhj4juE0WQ4vkbh03oc/l0fzltq
NLAntGtvnQHiRPKCsvuOpWd7WAacmGrDjdmeO/oFKjW2z/QQQ2Yzm5jbz7Ka
xjPMTpw/cErXVTIFTv9x1rM9gMRA3xH2Z1irILDp3aRr2IABLjHpINECQ7Za
Scw0msOWSV5UD2irftEgKywDy8HW1j9fkwOxQ5c+SwcS4fSz3f9lV2wCIjHx
AA/SLoF20sXMybf1IZ9oaqq8Ngn0oL2x1dgI2KrvGErUTfcV6fosaDs6l0b7
Zc7H/LW10OaZ8Jv1dt/uC9eYqL0riQVIQ1BpZdebS3WfQJBuKRLTXQo8of+i
Ja9HBLu7+lI11XNgBfcK6veB17eaW05L+MilRvHdcxgaMBFI88550CDCoXFg
tI1yc9EVBLFpXZhWc1novyjzSeS5HZduljkRFoV1k54NED47sZwnwAj/vLLg
pJC+XCRHK1gDBQRBNf6vDfEsNevohLKk840okA8dBzkmE77JofnzkysR13Qp
ZDJcexqcu4XVafHZeutvoAlOr9UYxhWtRyRLG8fM7c5XOjEqiuqfAdB1OM/L
//ZgEpNbeclq+HvAkV3YGO7RWuIel6s8p43sUUO5AuiSXhKashZHyph/xTN+
DLYFK05GwlHupPO5tNLNExty2VQ1rDjIofz4n1lMw+4x+AY/ARwJQNSXjJ09
8cNvvHCTXtRRWuW+UIOs4T36mOqKjKUmX3na25bHWp15RKFmSX8tvqVmcVb6
6SgSaQpO2ES90+JyUt7ajDUHZpj2ExMgZG08ocFQTG1ZIswdlfoGUAO/8aO6
pQIICp8/TRZZFVTiFDKt1clZrmw6mJDTsFBtkEFl4AlzSVzRkY3nTWI3ar2Z
jhs0kTs03WcVjc+6qVUtNUqc94KXXEolK84JHfkRKUh71ofVVfwon6qyYt1e
R1GVoeFQfIaQ4slqtibh7lrqstXECoplvksA/QXef45D/+mm59KQVzuhN+Dn
BZxf2aTK61dnHbBoGMImkn3MnuYxk90q07eIglbmZ0bCEWnxJ5cykpnWXKpa
cs3pp5tWhlH+ZW0kZ4NelX6JvX3XV01GWd6/F+wkVfMHAarAwFbNuLpxFr6m
BC8dCKnIiubzRkEZlOkFZOKb104kmej99qwwcRyMaiaBZ1jOduvrmoz2yWaw
IAatJv1WrK5iqt65UG4o9Y5S0Vv8FmivQlAU34iI9Y7DVFwi/MOA5O3RJKEF
XCaBrt0BIDQUc3WYUKZRHIX86SExaB1qdkIuI0Vij8vHKVkeDFQAZ6r1MOLI
BKTKgOSs2j0ROuda9FcmPdHk0W/ZF4LZpSIvRlY2SAHG3VBGZ/8SSpq/6e9c
uZrlXhlmkRk7bNL0mTWnErW0SrZHsduoP6PH6B0ubusZUx8PMixeewAN2A/A
9Cp36NCw5cGaMAfO8hED7k0A3+FYrDUcGgMJsSWvJCYxQ4/892/7mTDtYm35
2Awxd7cguXpQQc8pQzBXx5qoQeVC12B2+CaxxpcuIw2xRCopl7BBVyDYtbBh
GghLW85Yov5fjjP3Rb8Iemc6zdcy3nNs6dYv3Hxa+g4S1l/0Nl4Fw8xUbk2L
56lFhvk4UO1ORuxmJ7KCEORAkFlk7HVwJPjJSdjIXNqxth7Ww/Y1kHP8Xtjf
cxDlgq2va/ssIr/9HijRaaevj8/1+ju2QRkzp6vvA7yOpcgITTcjt0ldTdrb
dJo2mHvxNkTOmHKQk7BESzP68sk87nyulia2qPEaUv4ce20+41GzRqIk2J7+
BK/mxvl3ee7SSXlsQy9ZQ1yvYlIpOyJyNFolAQjUOkOSyrMPnc/j/VLUU7me
RNEYP01wfdQn6+mcSizPhD+NDHQs2BQtFyovVEjZBjRQ0KDe6swvGi7DxmWh
iHvCbPIGBWuR91MywUSat205csb+RsAKxLNn9Tu3ravz9Xf0FswSMP1bCMPC
430suwSAVX2K+L6HcHkVsdOMXUO0gH8Bntn4eWV8Hdc2ueTCz0KvXCuFRk30
m1A5TZdJVnCP1h4sGZRdlGyI6Me5Sg7nn7yxZvLhi/2htojAslhZGZBSW/1d
KXAIFxTyEgArZLl5kaNNkwMEgeOBEnwETsN7h/LWNL4WE5aUg5XPmxCPuJBW
C7OwrRcpwgf7JzkALFBdV6roQml+y2/T99ZpsWBUxMssmDDT2PAezcQhfx9M
Wby+7w3bf6zmaTXZVxWLqWj4Di8w32+hmyxe2TOntIs/l3KZ37A1+IDNzX7y
jr9p1cKJFvFmWV1h6XMgrkrI3MkxJSclD08XJS70+ihwPaayh+BQQ+wPaoXJ
m1zy+YLYScXoLcOZN2AJnTce0hXKAeMhhDSLpc/2IL+2KQVvelrErwEnfe9o
fQFIeDVl+JKFp91CRupltjP56a+HrwuKdgLTY0X69ArCRJhSl36SQ4vYjFEX
aFhGiT+2rVEIUw8OUlDoPKxQmKF7eyVpToz46JJvNozqic2PlPN+lKFFR6Oz
Gt0EpZgYDY6l4IpujOIcHAoTFJrrWlB+PJGMrcI7keNQQHZoAQU5bFulHK71
+0D5j+tmshmV/P9DgfWFaRoCWe6uyIkG5tyVKLOR+CiP8pbnIn9jA7/TezHk
gDo5E6K80PzSjXXVLwyxjQWvYns8yW6Weay9AXpLOoTZnf1j1KXJ3n5vVjis
VtbDt3acltE7SZJ2Gy1R0df69V9+hAj+BD2DfLTP3dUqNB0RGiLe+ll8BsWL
cHsmekQK8xPuRqks6pzSqW61bdyRPbUy2CuK+vKZkTKXMEpU0QkW/om/ksd/
XlUbakmLTe+xrzPSHm8G17uGNV86nKu7vrCuoztmAaehfoi+v9KysLhOhqn2
PXnAcWEljZNrXLcPBvdlLaZhZmikARgwo7+SL1f/0ksoqEaW9gvqUXJ1itWv
HI0+3ppaZBN/1ZjR5kBEwQDhIexg7zPi6smdKjyIAMeUXi+tYBSIBOJYhKFP
MLiJamOk+CDVsNG4LZTZdTh7G484yEvkiPnmX5uEsC6dlv1eiqkKnboRaBOS
ZqU0zUory5HwTQV1SILGYrv1+Htb+DofOdsDBVfq11B2bX7mG35bR8nbmEd4
igBMcSA0vWkhu086GD3SYEUMVJP2OEHr3U9FahOkqjfCYcaYAeD77AWoiHDW
GRvViTCbS7XYzpIKwNo/ybxhCEsNBZYz1rzsOJ3r2/HuYtEqCmQG5hNT5r13
FrYHKbwAlQIkaHUskP/6M4xvTh8ds46QIHLlfMB4IicN0tvBw7ZIA76g0fcT
vNEDftXBk+hx+PjLWIkvjdZq6jra5ozcKWOJfogWJ2eWX1ANuE/oZjyHJnQa
rUkuWUT67S8zMq9doySJF/7UqWwLJtilR2P1XTtm1V6A9rHH8VkolYgL2QIB
qenE0OYmFqsG4KRj8r1kHcNHIWSCCpmtXeZWNCUvd/MhvY5IVSIpZbWbWRgO
OU+xpETPZBndGGXJygJSZrUMSTqGAfYQD0Y0k54GEKZoTH2VxTTgbWSo0g7A
SS56YbPYwojm/uHH1y4/6Lhtx9T50rZviEt0HbmLYps6tgHSqvyseOF4T6Zz
guDdZ3pB2VtSByhN0UHNsJYk2pONcksbe/JlGFdt2RROuKuvSLb7o3FCgVy7
66WA6rdMYAArAvwcz4pKV5qilaXmRyY4ssyb5niwKuGljsRv4EugAUOURR3A
ipXnYvJ7dVKS/MZM8I8jqAfHrHTvP0xpfeqMZ+KcE6TTQedQqZb/Tk7xIv9C
iaMr5emaZ24wIPB7DCG4wNnz+bahgWUdAp7GE0VG03w+f9UcOZXr07cHW+N5
78HGUASgqmF6LpilE0WZP0sAP4u0xxv8n31xQqTtaaVUPB/YnDk1jkOw/qfl
qvrkUmd8U3CiCVo267DRcTVLjRx05lA/UDq/G1YJLjuaVvrwg1szkdpOLPFZ
V2vnS4G+FIkBK2z7fLV59hfOI4Gi5XWN0BV2ZTeRVWzGbmaHD79mr5QAGThI
Cua2IwtfPQubIVNw/H4GH1D6JsUBnhckuTOL+NL35eQNPKIxhwc6au7d/AOZ
5evxE4qnRg+MbITHpXXGG4jhHdy8bbqzWNGDMy5l829BFl5NTQIA16KBUn9N
5/dR/45JXOlYQIErkYVvz3spJ3SNzifaZf5CqA7Cfg9TkzMOD6Dp6Zvvbqoe
cQ/ieprLbl7j4O28nFuhUL7/ZOpV3z/w8ErIhtTclMqM0K6BCgpQD78zLpXS
fl0nI87MVOrrixyJTTGjYFldGPQU+gid5ezjGerCM6zxXNEpfUV/G5YFZDmx
ZKMJJvPPz5eXpYTfXfSrmEhl30HO7XhN/fsziFVGEWZjaIJX+NhqkHFZivhS
WtkbtVxbgy5HzDXsrHEdOoTeXZUjy+EYpUbwyV4St5xCAx/sHVMPs5DAg8nA
oTPZZKW/hxPSRNKIJyFKHC5ajFqCq0jqQgShHgUJeYl0376qfm4Tam5Eywfo
O9pqFxMkIfdE80BzcWUbiPOUiRPK5jyrPp83fG5KKkZ6MrrmctHuJsSUOgu5
hFWTiNYz1M/ugTqDZqk4EnK7LN3V8fCyEVEPSiJjlFaea366oZwPPmDlssMe
Biyi1GpQCoYPaOj2Rj5wj4DUPApiEY/KYmgwdG6hAF3OCb3DqQ79iTNbeXRU
f2LkE8FMUtVebDg1Sq712aNaa/sSXQv+eyusGmzPB5PPdf+BbnlJosdWeoGn
+76Mxnc2OBURYUNeyAg8m/acyV50J9SjyF+i4Lsr+tQ77PVUqZWhOu7fxaO/
Vp9E8Megaw0wofzw+75MM2Xsm1MYsoWFOLSZUwFnbOA6k9J34AO+4R3/1+Zi
Md23xtaL4oKyNv34d681q5jOw6ua61h1BVSdXOG00sagbNwhoiAzcXuiSCr+
hZP7U1PXwdIW/Steemr/Yhkt68ECw6JzczMQf0PFdSfnSJUA2K1S7kK61ZEU
uNtiWyNbfEz6S6L++yroEGmsGBRiAAgx5GvqyQes1pQxssFvW7mavE2u7vjF
9OkLlUFzJFk5+KE3QZ4RRNJr//8rPFBF9Nw1TRnlEvSy9EY4tgZxKBzhdqMn
seDfAhb2LLZaOrfKnzZsO1gnAQGK651bEXTkFgVaQbieLWaSDi6EF9qtPYl/
OsckmuVLlREH5igtD8OHG1fjRzTDApJYKcMSErLkzMKXcsJSIntKcLp0rLOn
aZU3VEi8Ojn4PM+yWs/k8aur74Vf3/CPBJGAsCnItpIhS+yndleSmEt/MfMR
PF9kJc9QUSumz9Hp/ngFqQimkQsfCzUOup38bYDAZ8sCZiFTgE4gfMzAaVkt
8YrfWVDS2ZoYQyGFsvL+/o9tPEVC0QmPIN4Z4mcUkKq/3Z4g7ZfNB5qp0trP
4+IKOkVTQKFrfTekL65/eAMsSaYElgHanKQWlBHvS+vgEWlrnBPj76FZMVxK
QH6FHse9n8nNYd7z5KiJ6wCBXNzc20FlADftFiFkLGWJGdlZXIGaNi8np4en
dtd0iS8Apa/72aqGSWahy5u7H+MxfUAZ7YRlX/O3K8IAJRvuJaF17Okq3ixL
rBjoykZ8IEKcq0845Duajet5X3yH/J1wIAvL2EBcHEnfyCNiu8rKtjjgtzYI
KdW9qHneNduafX64Li1qObB9KViMRKxY6JRe+VxMSuVCiMF0qGfpL4KkqKxy
vjzNP82/kHGILYZf+VA62adhdCzan1Hubw+vuJ03G+c4Lig38TKmwQmIk1U4
ZgEL/MQfwhVTBhYJzWPK4hxwRF6H8V4qsT1bVASdyAJiPnKov7LYuFCW3SP4
n6pcp5OH4ngMqJEBfyPaf3iQhzBZnpACwG8FJ12ySnSELwQfA31YGwpnvZxO
e2dMHMn0JY2Xl3r9NHjuoxW/lQn0z0rqCHPAzYNEseItfFjsJ6OrD86fCLA9
vnHuB/ROCV6czz0qznXlbMSgbt/eppT9Pv/qzoUdipZDXg41pClIVCb4En05
hksQu163ku8O/NfhxA8pD7So76eZCvCjL3bd1SvCQYhQ3KglVFjjhsqdcBE2
gcxCdKsvG6SIbicMJwbJ8EbZ9qCfapFQwnam33eLitjQ/mxPbrImzcGaHMF2
S3TV3bPOHlVre0K9YEYvdAjyH7XperrSABZSkFqw2ShlL8u1gRSUFU+/Y5F6
3w5O8T8ahjigmdhJkIT2+5EqQIImbFWV6G7DavDAV2rhFL2Z6DBH6gamwfTe
wQjwLQBS4bOJrnlheFqxYn1yAwYg3N4iSDP4+S4nB6TjaJYEI95rG2C3R0wO
1cYoyx6uRTtXS8Z3c9hRFsghQnP2fJJC2eiihK90nYaFWP6/cUCTsQSd2BfL
Py27tX7hNyrqZ/9nOzOb8327Fi7r2fAR9AHku2eKUpj1EpTPP4zqDUNonzkF
4iLkO3vJGYVGIGuQx8lrIzTQ8kTwIpNJh1WWde6eIfV+XqLH2A6cxm9GAgPw
OXOZdbvqPyinq3WkuGcmbktSUaZvltmSuCL+csO8CsEWsmMVaE/aZF47lxht
wQ5AWMQ2Gc84n3RZ3igKgkPPyJOluAkM+weACWKvcLv0MJjCD7MXzG2fuTFi
r3qCkJvmHcyNnPfJj8belBvvNId77WQaOE+j7AtOb0ba1nWaqJA/KSkr6+As
U3CTuOF+oarAN5KvrHliMhKBMUDxTiLyrABpuK3MfXLOEB2ESu+eH+tTIPSi
CoiIvwJNiNHtJUtAEI4LL8mEqYkSXczWTRllfauD7wg0YrYYFBLmS8qI+vZZ
BYWYigrsA+avparSr0sJt9oL0I0cXXltQmZQb9REeWtxB2bknyORXlQ11c0e
Sk3p9s3R4Grn5zsfSupQwAEe5MO7OcsuM24XECVtl+B7njavrefxcnt8hTcG
B+vboid5yCQvrG15Z3w2C1JnITkdANCtaQOASq1yIXJkOuWCh1cWnmkAnLT6
TTAx2AYLS//9rK9oBFHZ9V1+P95EIeo0LciqNwkJWdSuo49cdecOmtA/ys2g
Z7te3qEBjHwDk+MoIpP+NUsDUFm6Du6pDY12CLasAXj+3Z2QU8UqXUPmM0JD
t4XjZbMeixqGF6GGwe7VjKYvS5CUr1MOtql2IFLMHmi2ibNlXdb/oi5chVjk
cBwWXlNAQPy+nn5AYH/9wu7ZuKUhJgPEnJzou1+7i+dpsxALfQAEsP85D3zn
BFCTxgKHdUDN73vC1kc8HtiTDUiUZE4mqTuIA2OvKG7Xc4t9anEfEy29i51r
CXEKYny7Dx3crc4Nn8Az/xtGOJWYqFgEIqM2ez+an/sj1VXDBFZsPoxyHbR7
KRigNzLZTLK5phbRcYyob9RaxoxjlcVQN9t1ZIk60rmtSGw/2p2nzKi5YEsA
F9QMaHg8OSSE5dPIKCX862+RtQYaY/GFc4890aBeMO8z5ROVCP7svIdhSz4k
xbvwQOUW83RGLB/qba02SYzDfzS+blsj4Lnxlil7RYK11u+OY3E4MvwVwCJh
onY8BnUF8QuChkUum117F5cbqbNIBnuX+qY/oNzEvJGCnKOGFyKBA3TiahnN
VlyMJ7CvwXJmQqRshdxq+RaaKBB3AAxPrxwbdX0J25ezebfguFk2dMmvE0IB
Mo6mek3DFgzfZ1YAx5Xk3TBAT/sO9TAGLGcIR065SyWIciC7btMwFVHFvWld
55/BjFmjbafx7cdhAXqbEisbW44vyKweEVCRyTHq1Rs1iPF6tWa+/Jy6EJUZ
nymY5Mn0jtaBqZYUHbXcx7x+Uj83Io6ievq64BYBBlJu8MKSLWBHDU0wQCbc
vYC5C/S+ppQRLlSQ0gK3ctz/yckgLj1FI0bCn2CKoQqGZQc4a7tFGWWsZYHK
uAcOLLeaQg0L42vg6LXuy7mfeyef+MX4CaDLDQ90gux2MrrzgJt88GRD9LwD
kLcW5e52k5GLi1bTJqBu0b8FUFjbaMLgt+gU30rmzl3mmta61HakwoSmeBTm
nwjUGgaNq6MeFxvI9AMWbE2pOHdb/GJTXilSvW5DGHLv90vmdHCAH9NyqzUW
x1Ev1PCYUaN690mA9oIzSk8u8VxMjY5AF+U16P5WE52zx9yc+4KoLZnN8eU7
TubzWxGT8ZNHru1n+hjxcfY1cjrZTEeL2eGzaLZVUbwmp4tX/SW4NI8IhHI3
xwBwtsdCsTXz1J5oCCDR/MoavmP2kdT7B1JBrsv/KbtyFUefbtbSZnLkAS/o
WslmaPk97dmerlWQ4j+i88fysrmiLYOSmmKYRHbYHQYiS3d5HCSDF/8hst3a
GJYZGY89CQEZk8f6hF9bKc9udS+0VUF1QWlmi+s9gmKHao6AXhe9QGbC40bV
cyEvHGQkxtVNAfuSVaOxnofoMaZJiZ2rA5P+XeWWGrQr09QfsmnQGwlKZkVn
uD7l1Sgq1Qa6XkVK4UM+SjZpCefyU78g9daOvfgdhWW71THjT2RWJucgcy7U
07zQyqqfhDjfy/FC+cH0N4UPM9mYgwqHB6AsKUyg6wDxFtZCkW1KCC5a6vP3
sfaTYhXtuXhlVa/eeaRgJlh5gvdiTglKatHO1Yfv68Fb7ref1sB4LNhrwiW7
J6MqJXzcVX1qSQLmsCp3SBviFUcfharp/8gprh8OnDjoSF9QcEJpOjLoOXc4
4qCSp+npl40fffO4J6j+D2AkTTTIZ0ZAIy06oDR2UgDyZK5ZuyDvBU5P90b5
rZ5QSU3IFODRZHOHsfx0wMRJZJj610uX+byWVZerL1DaQt5LfRYfmCGGc+ak
1kNkz5Ual8iKtCj0tpPEQO8Ja3O69RpwcDE7sbUdqoDHyjR8Q2bQtR3cOuqy
La5uYPCq0WuDSS7sNTF4nTcsBGzq1W6Sx6sK0rFgSa7GpC00mguvZ96me4ws
/5GGFojmn1RxFPnnKM/vTQuM25WI6/8Ih9vvfamx+ztCTHkFeEBkTDcOWSLm
VGE4VniKY+DGvJXBpu2fXBvQQ0oVcqxnDDCReBylsp6YBeSp04eMlza6JRwh
AcY5slRVBsjsp7b4VdZ+8I86ZjJyK6qqF46c5GBRVN+ssH9NOSK7L6iwKRsN
n58DbhChLFsdkaPOpoGLT7nQCMXVhJy87WZ/LOOOAbCNYvozHNy0aQKyJkcm
a7iVceqfza/wEQ+cYLuoC1MY+FBSCGIbH9Xsj2JkejAXDHzd1nV7bl+GQ55I
F91d2MPSEUoiMXY6Mvuowg2EviLp7RshNOXGObg3rZfOls5b0tHa+wCY3mHu
/N5sLJLgfHSSVIr48gIbMovlf9BKCrmMk9VKt4XblXqtx5YIPIbRgaXOmZoj
7uLtbnLnQkaiG1su4WAtnwMF9zXCrLKDczu15sXf32m2k61I5TYlrB28vxQk
H+VwrlXCPonY6zjt01kkAViGReSifQbXq1hnX5XDQrVN674OelaApSRBtuJT
sG9lF1T3HJVHWbwG/e9mSi24I1CvUDdQW4bPVgDVd3DVFOfYJubMmJ+NI3vh
YvPC3SX/ybXwg9b2kVcCORnCRgZwUGifWi78p+sHSFjaDUV/4X5XBgFq4wLw
t3JZgnt2isGk1uxWMRJwxnM26zCI0a1IHsoJdzHtd9v6X/s6dffVe7mbe4Jv
+ehr4OTEbrIE80CLihFhp2HnHqr2dc0VmgX3viqC3zOQJFxixt4hnxtPFu+s
PvVjz11yXI9a6jPwTX/Cs0nh3zD3NM/kh+bnIAkfYQhxq29O0Qyrv605Oj8G
b8XXaKJLRcarM3EQCkT/jjnTcjMDsU9RrnTg2RnIxWPhkSsu1b+uR/4CrA/y
y3U033qMsHPubs5rNYQcSGWSjZVQYveHcW7v5tCs3xQ9tL/YtZ2KokoeJVdV
tKogPomxyhDRIo6M5f9fGe7+azvVvfo42k3txkqpJSxV2yi/wO/nZExVasno
D0aqP0GLZ72k+4I2g1Afd4e/AEoGNcYtWRQWFX1VunyzAa8fV2sfVl4zWVW/
w8YyC3tvRawPAhbTf+CLwTAZ88ywR172dsP3MoL/N2G0RS+yL/06xlapFK8s
oRg4iouGP4GhXOlmSLVnHSHVOsEYxEntQdDdh277q4aK2riDuPcgC4eBY0x0
pvEZeAH/dRkmMfrhh3c2SynVFxrYYo14CyJLyUVVkHZc6rgCsjebJ6Oyx5eL
dv451jr0qb276OSApN3eo63kWPG+ANQei9TBtCUvuGnwBsupDpXVTYH6pqSv
jSiba1h0CRouv8PxYqif7YhusRjF60OY1gzgvzRQfdeI9NeP4p8bwXNzOUgR
NhSy4FgzV4LMQSdeza0zWqQXyTdOzt6lNsqFnYdoEIRLw/OUUv1vKSGX5ihO
FgJlSsBqq4SlF2zBDljCf6Fs6Y1Kmdt5si9s+rwtdNTpS5aje2HeP3A7wJq7
rjAR12jxVAXYrV8imp40LEGbNBktu1wY7QEWC5fI7AZU8nhaPGYNn083B7N3
iWPTIqR3GcUAqVo7KUY00U1H3MPEJCrdxzyg5HB54WUpBjeHAVKKY2UmlhR6
Gsn6rZepttgPaD8bG4X0wLm7AzbcfPFKDh+ugtDyZfnm7SRNQt/yLUVL20Fb
Y34+e3AIVWjptTBPgJLyfe5DYkqZloQvNoG1dU0UnRUdnIuHVPXUxvAuYMM3
kXLS0L2ngSpZ7wOVFyXrSW6V6+BTn4cmjxqxGuLLty0phv1TI6DXkKwE7RYX
fHIQn784gSIRSLX6xVFMCgfsmnFMwy8t9oHq7XLTJzV/2dQZ7O3ukU7s5bSw
54oWKI6XrYIgBVE0c4yf6HfaZVTROonVtBC41JugrBvXrWRd/5F9VNg2V9wy
JSXT9cWMGUCXNvrKqimD6WIssThTco3ZrjsZ476eIfKate2LPt5rPw+GoXPF
p10vOSz0GJF5MauRBbWID6v1YWJjpnmgjLivkL8HxQsgUpiLi95cT+bDrGit
VhYgYhLl2/FMinwR/JOPHNjC35POeZqxbNHJwLbw9zSAA4yDbfuz/YhfVSoT
FqlDIUJuoKLLukO6daiFfkWQmPaGBc+qIVv3/V7oxf3kSI1+nTZ7WVDMMA5y
3Ij3uJgs7zfY4laHmbE2BkzArPuNoUsA17Ii2EelZl6/bSG6s+fxvscKB8BR
x0IQb2GKDw+zpPfjU882H07fwZDZOqu2LbN1gXi5WQ+EiGGjfPyM+Tj4lx1P
uh9aMxuZequo621ZO1yP6oCQxMQP0++aO5So+FcG7zpkQodh84KaFEZrZqEg
wAzpsXuNtfhqaxE7KN8aNgoeA3jNVVGPAjX64g3WWmVQwQ5IOHHO5M3rx82N
xqYGvwgp77cyCGSMTM77skZSguA9YY9GB3MFkZndyZ5WdWiLFaXqtf4jt86V
6kv2HfHa4IKQAvVlGCY1iXcZUx5UEN1R5g+tevJpzvGZl6sWGEDRhevZ0z6A
uZalsCfp+JQRN1YHYSm+37MY63G/Nwf2rsBF//GqacPlkbYznQCMkQo8aTSF
vVWe5CcLoH+qnp7hQM9g4dUcQKMMBKkc7iYAXa+SRrFHI1gOZh4iEw/UY9cE
LqYAT+Go0BUj1yj5UAXbX52GvKKSHaXt7ELwMbYZw68zrCi2t1hFtQRCvjkv
SGB/V7FyCywl9tre4ImdOlyuRkd+RbWQVf+WdMI2zWD7KCRA584RqZDxm0Yr
/EQ7I2PJpToc584u+hmUidLTajZ501obtv8aRGAQtc9v+D2GsDygThvc0E+8
2icREw/Bd+cyau/KTXeSIu66+lU5qU0nZ3ijryK5Sb1Zcyq+dakgRQsFNfeW
HeTFe8RR5Y0QE8d6qP50JKSxIRkI+2TN5nJivmHx+9ofaHGqThrlFjPQGN1A
1ebn4i85OYqiFCBxiLP7KZgCbueBQHjJc159DTHR5udIk/hiD3EkmQql0dPN
euyZl/5ibH0rrvlDBT2Y+WxE4AJHBTN5UocmDghDH2pmEpCGg7P6EytK+x6f
y9cqh9xwC2B/YvywCcQ0lKtWlYjXfCzBrJT8jouSTaKvveU+0uUhAN0oIlBo
R7AOMr/OeeyNjZ8LI/fhGw3QuEnwo+GIV8YOqRMWWm6nWOC3oupSON/mMuda
H8S/4ng+9SKxB2i9FfprfXCZGlWQpwDwiRQ+/73VkrzkmGh7bOKtJDD4bW99
Da03TnAP1MqlZKsD+IlcDJAm/YyM8X5WHDECNo7cyHRQ8JQTPJUR7emcmNzk
cFhhZDOxvB/4hdcWZitsHNuB8PUTLXlxnBKm9yQToc67z9pvar2YQtXmNruD
FmTl1EKFn7nW1YDHuKepeep63ziQtiHezN4pCdhaVSdRXAscrlgc5rLiJh7N
xBxu3TzQdQyglU7Kb4tjaUJ16APj4gu02SBt1ubrR2hgUi5vS5ij28cBI+fR
BReWS7V1SOUk8ozVQ5P4/5jhBuTolAzJ1XR0pRhwcUZpr+WLP++TxQQtxcoE
+FDMRW85f4af/VCqFLm9Hh+52VIh9Uukqexfsrq4ayYheHkjpX8tzyWtTcJi
UBxEAjaTnC81ZpK2EMVOOorkFWgN1wQcJ55NN7+cEErH+aaJwx4KDj2zrtJe
0EiWYV0OQqKVvqmuEpIbv5nVR8rduWh6irGQJ/7Kn6FLY8C9uzH2Bs/HAqPW
QqzB0fJsyOOp16GqCk+/TDa07A/nHx8LozHX3coDO+XMu6JchXwLScBScFY2
fqjx7E68BEvW0EeEHCd/1Ypr1n46xOuOBvSmsbSP8f7ni7UOEvAwh4T8wR2r
RxQz5cqEjnMtGAz+LCpmMzro6M3A13K/1gZedOq/1PmlHnocBb9QeNSZkrVt
029DZoH2jVY1nvKNi/Cq2GpoPtsQls88EAiSdMZ6taIMNwviF6yOKd87og3q
0R2NyTOmwuorl5bAggYeObndmYiIsBTcRNA1JQCxPWAU8RVj1p3loAQhu3Km
orqmx04MEIN2l+8N1nF3fsGktPbYxseGuL/YcXjU8z4y0967UOOtezRxD63s
2b1J57wSU8LlLefxjf9Tr7e4Espq659nKBEyEuDs6IHHeuhb/DGSKYhCBM75
WPN9Cn48MX5yvPcEkU9/vAnBpl8Qq5PIk8vhsPzQSeR1o0VLon1TIwGnNQJs
+KD8D8tShGSoapeeo2zD4SLyGN0bLhFF3uxUG07zQROyJvVXsYmGinmvGX6q
WgeIZMlGQdW+9wHev/hvaqb6yg36O5hvkyA7Fsc3F3/RA5fM4qDtm0z/h4NY
qfW6qqFdW0QnZgJkVsUQ7l59fSBoAPyOyTuY/4MNfpR93qvsTIceh7gf4AAe
K3D+lgYRQgW4PR0RcLmzHvcxDoAShwrWVawNm1evSzM4/mbYXLIjQAbQNId5
mXR466t3J4I/Ow7xzf/P4yP5MQJAXZXCc9uQ4UI9HB6+xgj7PLqnNEJFERSL
t9ftgZPcQjSFceprF2TX3SJ2ZhB24+dBhd9chqtZUPB3W8xbqWdxJfkK/Ugc
DVDann34Czp3jMxCpPqz1HvwHL93sdcyWsCIf0/t4JqyE55wut/82WIGggRy
PoVpaIujMXrTxscbCaujOiTEkHl/X6WZtWpRXj9yhc9KGMl20vcYGH87wGIE
zZdr9OzP0C9sj16lR//UYOZw3HkNWVQRosIGziILFVJjqFRFhx6ZKnY9CZ0l
FbGgX6MsXOUf7wz0OCwh/rg5x9PKRtdmMcSjlFYl3UFFuhkMGSolGEbB6hRH
9GTp5DG44wuOPUIdFjNOOA/RD7JMuWyBt0S8t6XaES42iPECZgKO2R2DyqwE
vqhq8/YIZTYLgasMjSqPggNfMsfiKj9eXIOB+QXa/q3Hsk14kfecH3pz8res
xDklnbTaJ7I/wZTQJ3w1PWTcfwHuWILEMJXx2+sxvgPcs6i091FhW876NPbW
5n5FFrqd4wVo1CuHs6C5D0PKwH/6k07XFleMn9Q2tJ+VSZGHZ8D0e2W+iNE2
RcyFuG+tuw5Vle7CyvwIUoooJjz0bddwl71jdiIm6jpJiKpbNa1MuWTkmvMo
qp5Eac/AavS5U5dFSt4yK4JOWkFNkVRvnV6pxVropEJL39tOxhPOXhTDf7/2
w7fBC1vlpeHM2wLb+uRDnvgOfs3jad0zlK03Dhj8NQqAd7HGTh0qtFYMftYW
jtxXPb3OLrkx57A7n3uLhHP1WmKTKUSVQ7tduFs1gYQMmrrVOf7RwniSHQLh
VBs2p06Yiu/8L3BtiBDNWvdBOPXvLCg8Pc3+jm5dz2rN7qq3xnLEGEr/bvEN
f+5lHvh8rdLsUZx5crI38/2r7cxMF2MyjBtIeQhdcWKeyMc/VbmR3iqIXzOy
Povk/ggcqOV+AIJWq1U56CykBV2FoNpqQrRcLHUnptMXQvkruQ35BSig4J5N
XqIbgdYlRiW9iizyTgd30v0ZRmUV55a4k7+h3Snt4Mgqw30IxhP01+ulRznS
qOK7FIw9nMGxEVKzHgrL90JreIFtdcGiRIWH+T99Zk39r6w/YvBL6Hw88jnH
bVAQZWDo94Yd0kGXr9CFWSbogyuIPYMkv6pFUP+uq+Ebsf3XI5yrMQJOoSkK
Y/1s/aYwmUYw3hTfxldzTdgllm9IbUt33o9xIADD00e08Qqxdka0kAX8OyAw
Hc3yn868qO06Xd71MuZ7a49qRkUpV8aLoQWzyUiN5pASPqyHiW69Nlgn5k+8
QijZHooD1oewU1HjXiquFH5q4H+z7v396CBFklWVoKIALUOKJdgwq2qgUObZ
17MyZzl67/OHMgzUFPOk9as4XJuKkb/uIpGaOJuQi9PsrNx/TNOl0w54imTZ
b1Z7dJOH70pFAi7YZnwf2an2Wm9v0CwLtoQ/1eubQkdR8IcmllLuDO1sFqy0
wk4WTqonI4ZfIhzwBr3pINret98uJCcjX7GORLXCZ/zpj7efyWZadr06Fbe9
+xq3mnR4FgGpNmP9u7advqHpJzvw272aebhhzGgHgXwXsuDf4uF8l8+iSMyQ
LU0l2lEBPgChFWi0H4/RN8T73yzz3w592H7H9rop4jw2Hz4GtgtduQqu6a2H
21ngZ6L3iJvQ6cXa+8+RJ0o8IyetCNfPy4VB2qQSamCJeu/vhldJU957GXqc
Qiv9ujTnVvA+oMj1xoLQxypHjXkYeq3rpmcSKonUpvs2l0GpXNDONyI0wwRM
9wgAt4mbbbKL3tKwVqhkkPoQ99giHnJwUTlt98LB5/qqw0ZEvFgqOo8ZmM2f
JDZEA7owlQDHKP0AeHs5nLqHBtA2XQYqnI6qORgE9AfeOGmlO+li16L1gIjC
aOJbddKsMGWvE0kNS/a6/JHAPMDT+4LO8Hok1JvLDA2pSiXnl7mOQEYNIw/j
c/IeLeCaBjBw0Iitwp3HHpc5COubU4OfwyBmdpj4GTW5zM9t8cb3ML/AW1eS
YOZ7pTxmR0s4cwrDYSVPgUzhAmm6jflmhUi+BZUZ1wiNi8cIYUPQZB+Q07xn
bXuarsvqk34q3YHHx3mBd3eDesdmGK3noDg1EpgAeyOs/+XlC02NleTqGaw9
5bW7VE2NcRv/nt+YPeXnfJSXxF9mRQ7x7DGyJxYFLSzrjlB/7iMkCMx2JlPf
heJo3smUGmv3OyfHUCXoHl/BW6SiW/LlFbsZNHwPtPgCQUObHZor4MCs6kBD
3JxjCg+2h3es6pjt0SQPzLQtihh4brkpT4zuc92tbw/KBv6N8+2GD04X61ao
ail/xDXSSDOireBiRiz1S6KKB5l7isVSbt4qQQ5yvJd1DHTufaLy05QUiaiA
uiBcLcOmHlfhoOHnVA7PbzTKDRS5Z/ddzTXIV7a0rji0Ax1g27QjjpkskjsM
pJvkvaVDZeXTg1BZJ8Nl0w6g7vJ6Eda7Gr7lnGoGY2+wP+si3o09gITrKB9j
2fkKUYDXpYfWkPQ1qeh4+cSsiK1s/bDtOSsLtLFyh8OZ2D/YBjFl1pNmn6Xa
4PYT487RFJl6LOqBKGhVDbqsTfmA46+fn2kKcbpx0wUDsYgv+cjLcIp4uUIw
GdkYf1+sGh+1iBprXJ/dqMu0S83N2A+DzX35whadZcuiCbm2nF9yANEnXouX
XGe7KA/knymY9o6wdyU6UfOezILlyuCEhPrjO4LRpft3Wt1+pTPvvPbGqxRI
7CaVLOEoNw/G2auF1f9RWT4zCL/6iTaj0oTpCVP6eUmhizhceUtc2GjSKRri
06GuzHKikHZ9/6LsZcHtmhHXWcwuj4XYXE3oSJz9UoE2ee79zHlIJl7gxfqK
xoXVRzZAh6CySuHq12rI+CnUXCkAskKPQnBxTA1PfLuI5LWRbYcs7lBtcWeE
56HZJxKlmnk5O3SXhGi0cch8IBVVnYQwakJwUv3Ghzv9kqpngNszQPa/04vO
NWBWyeVGiz6HvtokPN43R1e9VRZrkBkXYaCAQO7GbSRqvHWJE74w/oh+UXpC
8OaYKxknjY4OXY48+r1RXMDXILONGqj0Y9ifhUHA0PHGXqvV3x7wDffzrIk2
SiK/ol2IoDza8MTle9AITkdLuqQoGoaSVDRNA/nqdQZdAZO/FWGztXtNgRfL
QodjSghVnIwz9gd55kMuW0qWpCM6Zg3r9s2ECqmBoG5n6kM2ha5zPD5BaJKs
VsL7CcPUBu7vgh8yr1nlBB5JojShNP9fyKlu/K8HhR8V8BGs90YaLV72s8nb
Huyj/3iknRGDTC2dk8xtWYEqBXACxU4I1wI3/uA8jBhjE8IDNAtY+zu2mQuK
Owp4TI6bVKmV8BKHOLVGsNwOcZmPkaLEteypaQpUcY7gF/imCbXhIG7FzEbZ
CHr+t+h6HwunO6eUjaEYNbquuRQ7gjr+2619m0gJLzK6+IyB0TuTrQ3NAg/5
Ovm1YiyG+NYU79EIBbx1heypLZQhREXP4b8TQtYsI2o7kaPvYwwhOgANOL++
2pJyffHUc4jitraKnLcsBxxMTwdtbBPwtS+/6t7CSXzTSrwtoM7z0xm0eMaz
uXtqsPYDrBHGT750O/eeygJnBbh5vY+uXyBH+Efqt9NTXlzRrLWAclRqFUhc
nSuw13pEWi1S9D1GX75xNBHgdDAU8qZQPMLxRSwCAq6X00HxR5W7ifQs0GMO
DzZZuZ9kE8jYJFcOD/khqTIr3HWTIXH2LvacDCUPwTUxdqvKbMxDAHqOj/46
kSQ0cuy10+cbG4qbLHcuOE3frTBOMSrckhbEx+8mBz7OYAt1H6cSTqmfRU5Y
W1l7H4dZUGRiPChElJx7t8Jtk18nI6BaJ8wwu5tXeRUOWBt5klNB/EEDfMnO
kcxsmzhBZvaqqVXQf3YHdGVZEW1kX2xH4WrCbdjSkkbFKrGRIefHS3xXJoYW
7j1vf0bfjLNON4IsCQfcueUEioQAqQDnetDmtoC7bHkNrrZXn8FlT5/YN95A
x3JVw6As1YiZ+WNizZ0oS8dbWAJatyLNcGwxu1thX8jPc2Q5Ru6X+NGHn5Yc
jFpU17opTKfG7no5a0JS0wtohtPBgy/tW/Y+XGKPCMakweIvpdLfAwf2XU1o
PplBzvkwa3zCdc9SWR7LpFBusI05EN722LdLaSekaQ9oosvFo4BVlxe3Xh84
J38ZDkyUYMjL0yRRMDagFNVQ2Uex8d9rlg1OBKX8s9j37Fp4oiEmG+TQTrOf
0StiVSj19VBq3NLNM45TLKcVDqedoXzk0MkqG90it1ufVE9Jcnw+yWwMEbEO
vR9g4T17n9cez2zJV39R/gYu6aEaMbqIxnfATgolDoK+ONnG0a3R7liN88mS
YkZQGMdEZp1zP2jcB33N71X8a7Dnx9fXoDy7u0U4+D0c286hrUnLUiuTzRge
QwYz3gIFiH5V3qE1IK8V9EI6/ZbW8cL54LZaLwPNHhquwAV4KR0SqeuhiN32
KbJLokAdWxN86H7DDbB0LkrZUQHybTZ1gag4f+XRm7GQppIWMMZLNEYXwvIh
KquZ45gcsb35/fbrECOzmmN8MvbvFaytys3dTgR4irZN/H9HqggaqyV9hKVs
SXHrFLtq02s5fBvxf2Keh9WY0/HeVJWPrMU/qJ6HMoEPKDBB3Cxb+mflqnry
TGCKC2gKQWGOKlBxmpzP3GtjeAVDC8EOnPeJmvlyydYZtDlYVCEln4TXLzOW
UxwmTAMmx/zS77aM5DhCyhsbM6lbZZZIBOUMstA0uB4OFcaqLqOcDM0iv5mJ
bNm5kCUpVWuZb9WHtk2thEqlbiMLivIOpSA1YqZfXvkuNtrf+3lZXNBzI22H
7YcjT+uNuCVGMWhFnPBDXNWGN05KMMkcfuV86LWxDza2LfVsBlXNQWyPyoE+
dQkjEUGTx9wFzG83f8jO/wVW9ld3TH1K7R2B1tqGlPRSCR89ZpOxsD8JKAm6
x0fcFW6DhaS+tOLDM6dqnLFldw7UchQfaQ37NJKwGjuj4Ek0LiboJQrq6+cI
fSUygLRoC+6S/iDc04dZucNweAvetyU9HZAmhW9lLKHvRsL/AMfSy1LQmDRS
mCj6fKFgpjB0wfgwXLMN6v8WZPv+U64fvd38SSKDIhTIMTVdMOWvBvnq9I4v
DcohUza3qqHh6KLLvxbxFJwUjo73VtxmnpHRKZGEPgo+Oer3DRKaPaBf7Bp5
mnks4WdCfpecH3ecxqDtb2vt8rfIFa1RoG60OypFRDFy8STs5gDQwCYDlTKa
HT8xf5Um4FtsqjMF/d9bSEM28YToV7oFM5zBZXeNolMDKK6Cxp/w7cxOt2eY
4F2fcjk16vK+GIGglwi9etA9NbCbAplsvab9n4his6pHZ/uPnRTUM08+433M
n8BHeza2fdqXanBMEL9m8+ONcmRFvjjnM2a57SqDhRoN6Y3gyWIU5Sex2hbw
2qVabOk0hnjL/LLZarq/gaEAnWjUnL4lm3eO/9n1YtgSmSCA1mDtYPnqJGG1
ZgTUaAz2Nteb0CL3qkdL6Xoo8x66XQDC5+xyt0GLdM5wB+f4U8iMeQ/Yn/om
Q3gA8UNHCsMrxBLtIZg0r0zwEsfMGXw0iwFeMknelESDQvtzynRojLwHRq6X
Z82xfWV2YuhojDxAIzvIlwDq3qCmsxw/yR/WT6D3dH7OuRnH8i0VG0Mz+Iu9
+ilCPcRim7BLta4b/V+gGYgwCnOhGKc5ONJHeSSUCQY1SIr+70YfVuoCKCvC
2G8OzgpWwSTueaCi0wVpKarONKtK9v2+Du/l4/0KBX0h3V09bEsjypgsM1aX
K6N220olFtIJm1epn/O6m3lOXBSzQ583o4zOkDJLku7mal72szh43T1wclPp
Aa02QfBa5I4twNgVlkT2FyE2bM8becxvVAxF8UIpaS7jd10diwIVwy8ACsPi
dpfFOsFn9ZOtBYXBELXFR0q/NF/BWWTPXlZsRWAvRnWWE5/6aHaXvEBqeBS+
DLR6i94R4pnfBDXAsHvyax+xjypCsV7fkUYNfBZfRDM7wiYd6Ccw3NHZBkU6
zTCHVHi/5Yf9d99J7sWcQy82mEB4jz7DisRescpV1TxuCUkSz6tv8+wg7AFU
4zDZ38OAdOhc84tWbOT7urrH0hKFHMKTLgGx/vQ/oXVWy2V4s3+RCmHHqaCc
IROo0sTWeujcRWXBRYqhqrNNPh4+vgUI0nSWNLTOFj11OQDGNTJStXkrZLti
HNNWvq3tD2DdIPmMOO28e2E+l09fowoMCGODAXmgSAROIl0tqUr18wcqgzDi
2iuCbA/7lYXA5pPeppjCcdQ42G+HlJCDYCWt1PHaZ2fWNEYa+U3kYh3f4BMi
ycUFNssQaCb+XJFHv9ZTxT8DhSAJ52OTUMo+qg3uAMizATQ7KRul2N5T/WB4
dedcv3uncFSNnLji2hce33KDhA62EwEjYf8caAE9Q6jny8mqk18BAyiO+Y8I
oV+cK7fJhfHI8ubQGgyxQQtTLz2+CLjUdjdLPX0yiSY6Zn2HN13bcUp8FfYJ
E2PdjEWUHgGfzTogVR3s3ovJWHZJzkU2Sp5TBbKSmOUjwk3y6Ytp7Hjm8kzD
X584yECUN1IIv5aH8POcsw9tx+C7+mE7arwMkBPnxWGHT3TVQ7Vi4ZyqTWU8
O15PldBFNih263tVhGcTErYu6vsHfjEUShAWHM2Mk5mOgF82j0qjds/O8Xhx
8NPytOt/PkkwBDNZuJYAK4HQPGw0AyeMHLFhD2cWjO1HyZ8ePuoK2hST6tY2
ZHXAiL6ZWBsZjTl6baypj/2AHDzvrUuuHE3ri08RR9YFZgG9FTJbPmPo4Gq1
P6xhKoZ9myI6b7dZf08oRf1VPVoKvfkaF11YJ/NTeoyJFijOWEgqJ8VaqQkZ
yzkloYhKTRjVB0VUdaKnOzX2G90ULfqNsydnIA1nncBfIvmNuXtkyfZB8PR6
+FsbK2I5KN3WfRoqT8KXG+MYfawVI8vGTSIlfriiiHaego/G6hqNu5kn9wqG
nOaQxWvIJSI2YCEbruDxefwrun9b42e/qZ/mPMFddSKB8x3GR0qVIfJKChpp
xm9WFjEA903UZayRjy+aMwzGXw6vlEiys4JQJF5dH+nkTWJN13rzGd/liRny
7vQRQsgW0uTeEPtXOVWFlgVw3Zrgb/JhLHFYV9sKjBW+i1NXLGaiRcv/Bia6
gpLzKWWpqmX9rlUSk0laz7P3odayarrg9ls9QMOjkpVeNRrhh1b675sWpKMj
wMuwWrZ4/On4RFRxiRFbmcnrJv9EQ8f/2Y0ENm8+n2kWb8Ub3vzufXxAOBMf
P4OL+Td+E145J2jtzpauOy4sgTnzc83w2vPD4n3gzV2ytOApT/fg4x6E6XBb
7ygdt+A21WQNE80YdF0AN9laLDk1tDPnaAUw928Lk0zQ8kkZjCDEKtBuTgWm
aCNgpJ04akVilOo6UMZZDJ8k9e5ApERnzDviyvbYzP7S2liF7SWlIVwcOVZz
Hth9b8XZ9s9DWtq2tSnDVXyGl4blwL7O4hM08G1WGNwn1DgEWPQ1Z+C6Behl
9ZcW0B68RM5HczpU1UL68QUfVnHTgj97yYIS9wxnHRJG+PxO856rqynOcqsY
yw5XbQ0ujMRvyGCvdsus6uAGXhSWaDbCY/3tCUxH3AL8OVBn1cwtfdcwO+1O
T/Mmr/q2Orkh2vGiRsWsFngWjcaJ9ps/5sYC3pwQxVfclH3zrvzPHhfFzKvF
dym0GGT5tQJEGdOz2KsFYmCtkCaiLXSRbenK//M49NeunyqAkE7+azyPrhj4
h1dqJEHxAt0uIlNxQ1fQ+KMhYeDRWPMJn0oqbmWkD5+qDKOQtxUfwU5E+ehy
MjeSvR4bnYM9QV6wKwDOoaQ235ZyTbzb3LEa1NGcC0SuVG6OdTPHujZgOpR/
WKY9ursEuFM5k9gctdVcPaw5jYbk9EKK25awdQagfa9cwAGiGuK9CoXrkrq+
2Zu+fi66wy7Dkf3t4ikKQg3GVecHtvb+UUzybtg4ag4dXxU3rWwC7lrhm8oE
pK+r3D/FXC+V3hnu1VEu+ECtm9iYEXBMVoUPPLX+WCTRY/kQzFe6rQ8yeBNy
aNl7lsMnSjDvkx8/jpQfiiXlYDRcrnSZQxVQQRnjvu+N+0ID8OKBO4Gl6OB3
kpL62ToG7r4MZJ9I0HcG4f6a067Y/AnmyJQueNgAJcZXHdoSBu3VPeSu/+OM
kSkb+L6W5iiKiwuXWX7JCNfkVHhDQoNBV1oO1kOO3RSVLMn2VDizTglmAvJ2
EZrqW3x0yGbxHtWKOCxxsq/69wn57C39uLEjMODHF+Pm97+sP+Sf4aw/m7H4
cVOlsbfdgN2n/mEs0aq/BXKalKqkGMnjj1FgcXaHKGh6lakZyJYncF+2iVRg
d9PdRKnVWJuUub9/wkM7XYUgwblyC6EnGeUVEGT7N7vRC5bTVmt+M59Ix53j
5bLxSO0MPS7o46C/Fr9YuOCNBDb+R6dKfSwZdX9lnYOptsRN/WEv9tJdMg35
0fPHB3uXCa2pVzsg4M7SoU1zBUIQynJYJSeYejOcVR9adURr6PniFsBJA82N
C+9LoRX9eKQ+KDw6F946sGNNuiUydB/9bUTgcXZKbBx67P3/MIFqxDz3ySrt
fsl3X9h7ZLFXP6YEj7UIaHVtRy2GRusxQRhnqdRe7+bL4HCLaT1hIgytu/0r
98Qjp+PqoSTU8SYuWtjqmvtVonqBZNaS8VwWy4e+G8bqkTOPs3ku5R9lYGqy
p9jyvqisIT/k6YjxCWHJgW0OEvyR/FApMBMvFWnEjVa1TeCS/lEKNUpA+aQs
Ttu1rvvay+xqw/q2k4u7KLHFjmvuVmjnu5rOH+p3H1JIfDDgWtmdPXVEPLz2
vvyCHm2ELBqoD/PbboeFLD/HUlAjiOe8UgphDj9rLMCmGDph7wArC8cEgSSs
tM7z/pdRDOD3FFx/n3aMjgCczs9lL8ZS+UlgLLN85NHtnbanSaSS5TyeEZru
mVh4LAgm429caZhR6XVs5UREnxIMZMY2mFz91Hgde2PqvCitIEXvis2RbNs2
E2cqIbqgPQtll5OlUnHfwrKFfedoF4/SA1G00QWhObDgyslC6tLnJ2ZEAaNA
RN/puHCVq2QY5plRC5Kom//IQbI0UKrKP58Lwwj0h19VY2XSLDOET6MYZH+V
QSzwEwFMLEMIyRUGyB/UTiif7lwkZNsz9Ls1tVgaGpQLkSEJTiIMnzanxW2+
FuIblm2hHx/SHvkKB2iJ6U52x+b4TBrst69U7YfGykXqc5N1yi60Jt6chGOV
4Rf/9iNorb+hCV5WKYrpIKeSFJ8hH3JtgEhsSCfPs58TFfIkS40c3Px4Qf5v
yOWpQ22E74pN/9DNKHdrgncGMxfzWDXZlJdRKfhRNO5+ra1lW27uaecZt01s
s7iZO3NSx2OxToVj6yVLF6nLQJQ74rmuOljfNfV1+1LmGrUnJ5+ZW+9tfkau
kI8/6cVBgeIFiGOMxIC6y+V1U/JkZ3PyP75O/GDRAxhwTDAH6P5OFetQB4iA
s2O6DO8wG7yMJMCGlvkUZg3pot9CVCBb0iavJuUZMfxqShDzgvNuV7wP3OTD
27IUWBEyRCvwR/LwUR+Ij7F9/Jth6izI/Qbu4EH0ZrVP0rYV5wiRMESDcx/s
ZqEOz3TlwRMWzZ3utwQ4xwaB8XamAufNVGrlBf3Nal+5zHXwptVKrX8vtsfC
WS3ySvrAlDQAV3HBVp4orgEVBwfaM/ztu+F0+k2/UKEaid4lKvnh0LyuaZdj
iEI8RQ/QjAoPePb7SzDHaCpc+Pc8Ys6yeTCsnbAioZddU31MqCHOJgFnKpKC
J4FAUQd1v/dIsOv3UXhgcmigXwgkheYupEnUxTFL+pkTNSI5o+nWOy1Zh0Ph
McbMAJAind+Mp+6qEBQgpA54A/IECGyE4xGTGtz7KpGJ9iv5IiP+TBZl5xFp
wfGCIDkn3xuAZvljTSSa6O1rHFHGBT1hY+1r3C8aKZdOZl6934g2zZtr44y+
v0flZnt3v8JYQmfUh2XXcf8Cp92ykGGpj9puOtNLr9LF1kctCMBUyJ9B5Fh3
i7W8SumCyICvXlJ/eAT1Ltq5hhbbImM8bpJrfDECYBff3LOX8apoWUKAF1XW
eeXkk7BLoUsaPu0szC+7fciH3PnVhK+xf+4CCUXNwQ9B7hzSj9x+niGa7lob
vwqArHbLClrDfBVciyPYDSsvuUE+xfKTC/Bo4Gzljb+wMayuc2/ua92fNWWD
kVLGo16cfo4RUnxiL+dbaEBqH+Qgd786JO+TPraZxoVUUjtNWc5m87E4TeUc
18NBx9qbDOckdRi4rXFYRJaynzmXsY2Ry2T1KXpaCTV7ckZ+RxxEDgXQrzzS
AgTHD3YgHs4nF13WQQYEY0hdAen6RmvxGlp3Nzlbmn5A0f1CzMfPDBtt0WDN
EPwcBgl26uJ4LLbRb5V/M68DpAzumGOiM7QYLknl79aiyqsKiDpNjTirbpcr
GbL3qjxEGsoOkfEqR4P5UZfqIh8EqnKfdy7/GnSwn/0li9zka6k0IrJIuP3f
ND5TLiOjgkWw8D4s7h37i5u9po+joai7MKkzZxdpVLeTE3UgoonqP46zMy4+
rWXZ8nCDWS5CPA7TpNmMeqHsnjxIb6pRypLxhEKmhp6UqekMstmd17SKYzNi
bsE6s7cM3bSMMkp5I55dZQQdVKcyYTJQSXJzJaiXEZOhKnmREiXXJtuxmBVO
xzmM6fuAolO/s+znNEq5DXijzAgYc1CiQtYLPkombmbr0DJxK5rQCL0LKG+S
wbLmr4eA0pfBHGJklnPe3WqEtbAakHBhOLzhaFnfbczO/eQkPimNwR8EVIDv
cZRuCMSBPzSzgQhHoLOO0WeE3a2/2LBlcAc32WGqZIHx9sDVMLpxfeavMA1n
USbuhOeVeIwVRKL4WcsrZuoxuSDpnBYiONxr+z8erTm2XdyOAhDOB+h+LlwS
ex5q/ZVaeq+n0suvhBDQ9N3AijRxh2hmeG4OVOHjAyAdC9998Q4JXrFgKFHW
t8qbjkKsPXq50c+I+XLssRXamhJFQwg6JF+8m19Q5ZxFvP11AeUqsVpeJcFj
HcVr1mymCcFkr3zFgcdmfXMBa2MY5DYRoevly/972vsyXJcC2dEILwXzWmIb
HorbsOSeOcenGDQF1b3kYByymqTZuxO9E3rn3bWDbksxRMiKUb95b3K75uti
ihlZTYYNiVgJrIQ0eCzVcy+bxv7/5fCnE9MXOkWWxRbhv0KNU5yb+JaF7doO
FQzcefYga4fBHLk++qm6jYsrl5rTbbKlqs6QQS0cFFeKbFSqmsKUQsuBR+8s
iSXlngcqMLauklYYswaTVHi7ad4iNPLLpnwnCbVjH6euWaQiRJJR9uaYwshx
joScNkACinPsfe+Yd/aZtSnTnRLLle2n1UALRy4vN0R34rK7TbZql7MMIIeA
rXvaE6r+xd/njMpLJPYg8O8OZp0zFViMyqKYJgWpmbmTC1XfJ4NRGUUQZFdO
/1AUafbWAIviYptvGGUKW4tCkoALf3+bL3C1SxQ7tqWnY2Cpme+QDDC7jM3h
A1RGIxI/+0kB/ITNIABVrouYcgcceHwxuF5fco+aJeSTgKbIZqLBGCIVd/Oo
k72bKwtTB7oxljfDxuYYVeuUs9FRqGJIzh4nHerfLsSCLYif+n7m64RhGUv8
9o2JWJBiJQE2KItGFL9kvvGNjmo1Ze2aT7T4jx7fl/J2PkM8Uim2lHifwHaC
xKi4UNI5flTl4MiL/hoHZvHPjMgfrIP7z8XzIbgzw0uHRtsAyFoe5OPbJhSl
21IG/Oi3JZ4Q4nV0BWBm+SnF2FcHgEGP6zPxuaKyNkEocqxsooy2BMayJP+M
kQM+DSSX5yKO0NC7OtMpJtkvI60EjcJH7FWiqo+VoOa0OLV/+Y24ZKasVFUW
qkaAxyZiaQli1YhSSIwcRdhEfW8EWsZH76YAWUdE4cyd1Gz/ZVehrmpPRKeh
AYEwTGKPGXZuYbME6PrZblhrgMEBG1BbXBWsK575GVnq+3rCscIt/QPbdYcZ
mGPpoIXycPjVv/1uuvL5vIjamBrIEqT7f+3QyzXMM2ON0NXnfc4WomsJngi6
mhi+zkD5Qc+NhRaK+cFfRZ01GYD4AStj1X3nsh6dwLcnvw+pBWp7C9uNDQNw
hlZxpQ1JRtsaswW20o5MqH2hDV37yz9MhOUV3pxdl3NuXifnDS37SOzg1Feg
ckQLR169oBAss8xanCBZde6TGHbHAzPc19IW2vXT9mGc7BcL1PUpkrceToxu
o6jyoP3Y0jlroejiAZ17COJIJw+ugc8rUjR6M0yR4IKhizWLtX7BEKwsVa7F
YtEvdt586yH21jp+ECNZ+FktseISlU6vqmXzK0YL8cG3aF2Exxmx9Ky22UFR
eaL4CicI5nyEYP5Ppa/PVjciuVqOGnObEOLNATaJit85/BxYnwsFtsj44yio
PijSFZZLCbxh6yZI8Fkj1fZQuIYFuLemeKfrCTvDfPgtNuyOaUK1oObi8KPw
mNQXExk45S2GJ51fmMQXYJ9PKFFO+S9qyFq602nREEsYK08nZx7ngu6DCXtB
UbO9ADQwY4xInZ/ez4OInGnk56jAtUe0PbXkdaQPYfU08+EikuuwtmKdaNgZ
dy5hb+SU8zU1Vl6kbuLk1/Bs6ewZc41mu9KliE3i50RiXQYzRy4wlwhqqS+H
/QLJt1BwadKLiluVFxBa/RcSYOGjMbhN6gvkKPcrty9BksUK7p1MiSoG1nlk
atqXQGUEfh8RyiAe0oi+kT60Io+FCpF69kJjiZkY5yvoZYV3tVGvHz1KJIOH
0//LeI0QSJ72ywiBdA0eT1PtDs9bVfPftX7axz920u3lqHjYNMymUiSdG6AP
v6mx2Z4BOWXOn2/ecsTzhP2R21Q4W8qO5qRrAcIVQiA8r8n5xGwiuRcFi4BX
uTEIsm8U15qWzQWtqWLmWAbT0O5sfFLI9Rw+YbxRsoYVjYjsWvAkXzdbisZ0
q6nki8yeZKc9YTFEVtA+adqAjV1Dgo90j1lvjHj5g7yyxCvnDnX+3ZUm2CC6
vu01IRCuqLvLOrtuX89upnMD/WqfVW+SmriSkM+mGTa2EO2I9CzOvrdLKJYn
9n9DEC1ca5KeBpUuOZnZcVO85WqA0TrOy+F1YvmhGIklxmBjZAgzfcFWbsUt
Dx/UyFtYp6u88/Jk6gTeZfSDmV7iHqW1Tqeuci/4JRWUiCpW/xWCSgFEu3A7
uDBaE/nWTZ1r994/Ag59c/J2MUy4AFqoUp+pp3fii5S2sMon0xJXeDm/oR+k
v/upzVN7FSP56usa7Vld849j0VpJcD1RatdH0Wrey+sLvikLYkn9vmnjleOw
XcF5x93p+a1DGcZuHIU+tliNWSCdoIav0ktFt4k172n0tl37C/L5jzb1XLm7
mSa7pPhuSBzB2OVINnboq2cZOQQd5GEewK6OmTObqDX0zjnjt552UstGJGR8
dsjVyMjG+kKYAnCKux9CqvLkTLkHK7MOn5V95e1XwtAiy+bDKQCCfS/8qW5O
Xdxyt+iDoV2iNUZbCIYoqNu2mPEyz04wbrlVu7l5luXEJZS8EJYMTmu3w5nV
TJ/OjYJBqF/9limMtIcm7nrfcJ9QgHvFCaPd52YuqsYmFCOBr2p8oCoAdvdt
jZQOWFCbNH/IzdTaorf5RQOI3DW8nGpkd7uEJ+m1FyIJEpfnmDPn52wCe6LS
k3W2N2OitVbG3Xk18ngWil8uYiOScVWZo6F74WJo4O5gQGRa5ICiaBQseR6l
ofQZVYI0LJ7GVcYHu2SI4IP1DGYRAfbwHQ9pwWornGk9s/LgrE/bjW6KndOo
1PFLH/Nees47dSSfieEOQ3xV/yVf3FSEUGW0QVK5i9POEUXfPYK6duAv4oHB
OXrjRcKMbFXyPvCsP4ZRb38o7+ZoUevVvJ3rbB3mnzrvM8+oZqWCQHjvHeKy
KpXtgnzqHJQze2yeyYJeY8CR6yq+BupbwMna7XtoqXO74Nz67hmoQq+TjyLb
+9xowN/0Q+wEwarv4n8drvM8P3q59IwCDl+pwVcEEwc+bY9mc41EV2v451yB
H76e1siisRtFFZN18o33TdbJ4SLhpnH6lDx1c+vG2eghSlAfpUtUDk8/eDl5
1CC+bATCV1BM32oYKiBzPrYOdbxmSiOsh75hh9AGhT4/toTd9RCxFvfyv7CS
dWNzZ6xljxuM80O4GeuhtgqZySI1I8sNpIX9fXVPgOx6TJtI5b1TS8mZgs1E
N8uzRNNFQKFpDN84yTvTVMvAxAGznYgfdiEYKV18IFVHHGg/QAhyQIgjJczg
bGjhswX7PytwOf6iy3aC/w0OvctAL0/WtNqdrAKykz6vSd9gFbu+N9SuKFoa
0FA9lUrcJJQT2tR8Iir4wf6BIB7Bd4D8hQ4R2mgLmNvywyoDojARAD0f+6VI
ZVecCvOONDrHPsEwhGfa4uqeszcYwd+7lYvCDOj2Ogcz6rNxYTzqOGlWhdKp
bdw9JkuLimT/cWLGnL7opzxSwMi/CWUiSGV+Dn0pWmvit6Ckrqb+QUfkfbI3
uSailiIoXzCKy5sHwBKavOGmdTI8J5YHnj4XhbfSkYvdRPQNp2nWba5SCL+P
MRELxI3IAEILX4POjfEfWgyB1MWxmXAxVKW0iwfzAu902vKR8YvB8ELFBqTn
hslqGgKJOC8pkwhkRpZKpHqBnKwv4M8Ljo+Sy3eJZKL5wvXxibfEutmvmWC3
fnV2bYe8y/cjgh6Pdz9S+cWRfODCT5D3ZMfrVil/0TAp7FNuQW0bK7KEdSoq
E5I7x6UmfQ0aXt4tT1PKTsut+/RPTfkGbmQQo7IAmmodXau/x8Hm0wLQHtj4
iXFiHYfn7ryOjxsdENmZbYgMJSHx8HsvASF3rV9JyG6GLwpsA/83y6nPzclu
OkscUgpD2H92v0Txx5IjkSDFVu/WDH5oiVoWeRAI0rQQ44ViNZB8hS1PsfCV
pZ1GTcyzRrduNm0IgKZNh0k7xIZ1V0zJEWIZuI1DhnvQMlxqoRpShl9Z1UHr
xjL65Nc033xSUHrDDg+73CQZdd5+xMiigcbPZWzOjnuUx+4AEmJgEzAPl+eH
3IhHgoi7JPjCScpdKN4Q+hVtab+b3alCC8RBN+BPPZegDNZxLLMgAiJu+P3A
LPmNA/5z2yU06jwoTc2SSM/vl/UtZFLgZ0lwRaCQofYg1qruNOoircbG2nNM
psDj7D8GVu/sBBIkSMwC8+a7sWhhJKbCqCwx2OjynNB6qOdD8YgURx03nXy/
zgXNNZr1ZVyL7MHl5kZrVqfkW9L7MJ2fDaOfwwzEs5eUs1sIvhIwG1x1JNJz
EVwiJQxi28rrG72NHeZZxelg07Stq8kN60byqln1DzOHT3gid6tqAkFXqzNV
OxSyNfAX8Q4XP8mk6GrnRhafq08fxXqia0+PRAbqj//BOcvyk29svr5bw4ni
jmP+OiUWCL6ZXXTHTA08SD+tKGskjb3Bvy8dmjE3+KYcQZGjK1irXynHG68b
c1vgiyLr7yMpwp9Lo37MMvIiS7r4wMrcCU+ujW3jeEe4KjgVAnVnBhVjVDOz
9+lXBdpcGpk42CHUnAkQNmccr2yWLCdYOV/fGxY2OvX/ta+2CKqolr0NmapB
XNNgkMTg8gsGjr3w/HBD/q19vP9xPT9po3QrjwijtBPS0YOm9sXtm7Z1/EUb
D32gfDPV9ZGw46wEyRgNm3JjfnNfxdSlJGRMDRY/xemaiGmfj8f0ZeBRHUGD
b/DpDBIPtc35FQqhJ1HWkgjEx75Om69aviMFzcJ/28At2US/6Ls9pAfah9qE
igNBFnwmXlx5d4y/bV7zBQNBHY46K3MGSwME8DWAa9KRXs3e08RZ9mbvTToH
vHXViW2HZ6KC0mMZPEhTj7EvgLVUDkVNiOMqjiUauF/qm06KyM/rW74Kfz6Y
rhVzofyi6KQHH/R6WUCvfAG3SUK2OFwuEUjqFQbEDlmBLs6QVd01oTvOOpQK
3RD/S3Q4qS17XWdjztosO6km6Q7mqApJnhtg6u3g2uy06mJQq4mFJ2PrmIAF
2hOjjz2/6j5K5LF39lmNyLrsn7oWI+0VouYyw+Xa4Px2z7s5FaIWXm7KapTJ
5NmBwvWOSEaWwa7LVnOM2rWpzgtAa2p7kQB9rVp4a3JxYMMACQCiokLJIw/t
PL9ebG4MxM0ZnUQg0D8F2PaUk28oKFDNAqjq41EldiUWu8UfeckTPAb/+PS3
mc2hfRcY5R8dlFRZnBTok1Nxb99QCeV5IYZ2tVDClM4zqL4HYEXVTgHzPItG
4dMc+KhsWSMjj/OBKIxW0xJjajjqbEjJOZnqA8APC4oVjVkcRkEp5tYWAKKL
yPZVvOVoLtiI8kBGp6gACrYGCVuote0yLVwTpue+BxTNTPQp1yRqMAUo7hsF
euky/RsPxmwVSAuJN2ZcWR/bWxPW6q6SnxzsHtyGiL1VGpB3xUSjCPoLf+9E
74j5JMx185MJ9nrjbzYMuw8i6VH0jefve5/ZCUxc2bZ1oR2qjG+RqXaakLBc
owGM5dg8/67UeJ9/+Hz8sJz4wwkDWj44OsNi8QWI87YgJA8A9jEXXlZuK4eh
QOiQGHhNHk8W5cr4qagjMxICYFnTeg7mlosJUkdfDTlyGVjEVTy5WQyEnlsB
ItjMeNzo72b/+uDH8ev+K/VfBTd+2BCIRi+uANGs2qERqcPGCXWjj4A+/kXJ
73awZ9AEhnynTkoo4UexMVDtPHjyo1VCVCVQ80r5GrCw00rRRjKti8lM4YnV
1cchEUgYZdz6crU9nr7bT+BYmxu/kNEJd250n7mcLPYtJtFoV826ZcRy0gBH
xHiRmSACkPSO9b3FiZOjeWD4nkkLRhTGgqEXlvg5aQgVK9pdSGpZHU2hNKT0
3V977YlkNYyBhDY1H5OqpPNZnzzOyoP66QQNrPdtoaFUZBK+g6NIFH5qqjvJ
SL1Itv0FsyXLiwXHe51heeVihx41PYGtzFgzFkAkPZGkjZ3JECIFb8+jLla3
7EMDYCET1r9urKW0V7aIzS5fZ0R5AbnhMMpfkbsd6C4tTBGVRoA0mMyheZ7h
VeCENwpNIp7xaHEo2VmbdJ9Hol9007GMxFlt73z3C1xhuguzjoz1uZ73ODrd
cA5jR52MciUJThh1vV3/OK5qBoPlvC1J5lzW4fp0lj7niJwXwxKy6K/rUKVU
esDtnvgL/bIFX0O0+Sb+DE76W9BkEinJcUm+e+IJ6YuDxa3T3KT+/+fkRaxm
OFzrqqQmDeWUzhsx6dQlX06x/PUeO0jtsmfpshZ+vjNNJNNJDtfnrvgcT0sp
Gn7O+VfdQ1oTKfORkAkpQRAji2ORNx2MwMdsWXNEtNHa8upui+2Y+NxvhXqz
+LI7mHPQbDdDw7pFO6PtwLvi5d1a0umzylEbDLSUghCsbCiZsUi5L3p4Hs7R
SO+HvW2ORD5U3YE+6cptDt4sxAoDdMGgnVsz9AT+6kfx/azTJiznZ0KakX6u
8rSB0/bhkgPh1jZF9uYZAli6KSq/in56TKaxuYEPV+Mo8BwGOJZM9yn+36wK
RMeZ9zq3zZvCxqQWT6g1DKp4eXV+wzfrXzvEuMHbINe6b7SKjZ0EkMJEGSUs
FDazIFlo0AsPPyeZVPMFv8/Rdzw2/b4wTpAg3HGGhgUMwachZFtXxEQ3BMUa
uDoMfuc6cga681IgBkr5JMdKyQDDlDcHGCoOfAwHAjb3N3VZ9DQgju2MXIkj
CrjRU+fG8GeX6cnk4uV54cb+zjFYD3uTM1/HNd161LmngohpMBeL/YRRqYaZ
96Ecz/+P8kGL4WzLaidFTGBNJQPUuvV6WAqTG7JlLac4aF+TH1a4bdo7+yL4
L1OQ62buIEXrd93bDzQx91mfNLHBndb0+9zBumGLt6CpElf4pTjs8FSG5EGb
W3AXAPmbP6CCOY6Y9jSd+L99vMWTDYMvHTnFn+2YZS54O5iGV5tSL0Rl/MHh
Yt/Wfqx7IrwX2OPoxtnY+MGJmLcTZImNUVm5wuJic5wfckVkRcdqHpXQcc3C
Zw5nVs5fFkOFQALLXeOGEeJzaGePHyqi2eisy+py7RW02jUF1pQ7X0QLKT7W
xQ2e0+1eiA0I58eZ2amwJL7VS3TZHUlvIvMJRw+kFQdTAGlGQnNw2dmWDzeQ
rGqlIqKfAhk3E4Kel1jucFvUyoI22lBdQBBzdLnEMvCBBoriwbk9RrBnqwNE
Ju7MK+nohTcgxsvfsApn9gSOA2IMDa5w1DLGiJFXmC0avEYlsAkouJFnE2dw
Jl15mWjgIoRamqKwt6144f0/WxZyAkUF09PW7jY3TNFGC53JRn3QKSMHp0Es
c2iL0+ko2e4i+Djeg1p+f3e8N52Jm22DGUhosvXeMVjdFAJ2/sSsub2v0Ar4
xlxAgkQZYV6ljFCCRViboErZZnMxRdHf9DVSpdXRFxTVYXcV4ePnAwFa+FoK
1qQql3ARHOwcX8oupQL03lyppQ+ISZUkl4okq363pl1U/mqI8WQAvgu/VQlN
Poi85qgXUWgidRjyoy+KP1RhiG1PVs5mrIgvxvSMfVdJ/5qTTtzIbpJVEb37
t+6QQMaL3GxsI1BEknvtrhbus+1bwzdGFlytLj9mijF+LIQyiDEeMPyfUrpL
2yCLQtZjAhZcpsJazzbFFGB0CKIPKGKi6SkoKQ/vc4vy1ywtLdg9R8TJOwSL
VJ/ruaZeKNxhN4W4HqoH+vGmN+XV9qH+brCkakiyiKQ/f1kHKcA5uGzq9HWJ
TkXwvWAhjuTZpfcCkp/VL/SRlyPdrQsXSrb+Hs/GyzGrU0RC5/GgaaxGhYR3
0WGYOdSKqMvo1vVfjvI70igg+oJ3xhRZaE7SPCQRPS6Nyw0M/f+G1JlIFeKS
BGjwr+RECqatb4axS4xpLPr+GdxLSFaDlEX4dzg84la7AhnuZGTIA6qdftaz
AZ4S7Ub0d7GzPE1IqjKKXQRosd2ccEbLeeJ9YjAxQhvpwwtihdHUgRDRc47O
QGc2GyL0RPQEFypgPuw9XfrKpb+5S+i/u4I961qAhS/duLdJDTLhsOAN3YPR
KvT2dyseirKSiq2+jL1LIWWMuWUNMetLQT2sJKSkDM0GTtqEh/AufRV0N87d
S/gZDG+woa4/1PDo+TaINfYRjon2hOUkGwbG6W2+ee/l3Cjx+W2foa1e3ALB
hfQshti4OcFn/2dgwdWMKZyizbVXGhIB+FbBz+nYc4sCOjLZWh3HTcnWFfc1
hNbsVNaHrml2nbHMTnW60Ewj9+ZgElu6lkCxeTOvH2px0ROTRmtP2TBrprrt
YqJZveoOAVkIk+3p+NYBxnKFG1oBlrj2ecFPCGxV7UeTUhYPAQCH0ide3/tm
eBtSjYFBKIYF3ze/+1rW3HMPhZy1g1kFg84DKBoR+Nx6KdwyQzGOQw2adwm/
2exAi8aLU51W7xBpHMu/XDJNRsLyGA9yoFcjOy8ixMoGQVXklx7OOeGffbqW
tkzIUdpYXfLB4/burpxPAaRB+QGfwgAlq6fvmyM7wnfCOPfBfWWOdjMRV9dO
l0V9vs+td9N9BkXDRtLDunqKMYmGNpUkZq2VGEvZ5c8qNI9Tn5eCnHyMUHLk
Xsm8sMCBZHUNTrtKxSSM+VWxfhjDrUefBCazZpHBZSIagZVogQ0A1BYgPww4
f6e6gnInxT0jXa3udCcsDvHK5+1DRcPSAEhg/tGvoX091NjoNSBnYPtLWSkZ
EDqhVLFwBkr4yGxw/rcCwEtmlZ8gZpi5waYNKclSxChcKGirQ3/6yXkfZI0U
A9HrwX5zNIyya2QMHf8MOdc1otB4FrWh0oKpzswjBf3r5j3RNbL015ti+nQW
CmbZ+VhbqWAImHkh8nIwuexDnsn1EwAPVC9mAftNyJsmiat6mavQ6Mlxwv7e
QjOMt/XA8MtR9PzPfhPHSkdHkDQQ6JhRmczKnuPRBH4zIYkZcIiBHHkvgddv
bZeh+VtluqWKAT5uQInmap+DbaEhBIVsB5iWOPHrgL5a0uQNZdn1oo4Qh+F4
GkWOiH5UkIKCuaQB6Ig00HyWvQPda9rPjxWXDPzEhq669VSoYO4euH9/wfVB
RCuhDzH+qglQyMRCkoYHKt5DWHSp29e3ayyIhsc8Z/t1xTS/9YyuBKrTiu/g
LrZvBnxeVwKW6ABBodv1Nzx0xE/WRS/XhihLHCz6l4D33GF7yj+hX2dRLo4f
fKKlpHqrpRyGhRGbL988XnI2Zjj+eJiyemYF7tHiIUO0AIykEUQnH2fq85Sy
KoPFb6CWaX4u9hK+tWn+O9hgu5ZNX5ReDPfiPVmHziFMJQOAygkxBqDTgxv/
3V2gaOaQzhjoMThfYinZtal54zZoCHXc4s3nziJ8SiCfuh9/i0H1SgYi3O7I
UK9gmFLowoSXI4BOfjd8ac1Bc1w47xT5qv1nPG2r3meoMZwwbZg1Jk4aqC1T
GjNZpbqAJ1JcQYp4Mv9T+EUKb5NJgP0kXRz11zc0TR1n6V3XQPponw4hKfwZ
h3NMAok0HN/Ml6UN1rW0XUgmiDSCg3kcHSY6WMw+Yn2p0EqFgbRa8gXeEsLO
qg0pOz/lsBImWWY0VSEY52pfkNtkw/Oo1wtrEY8CVXZG1uxVy9xhEjdhT3lv
sA1QkvieWZj+t+aaS8BuCTaxBzZ1KAChYzTfy+Kw5/yilsFgxBP3CR2Xc7Lo
pyQNb0uWDnOP4FsLukla8ft0z016+QfKqAuD+eCgeOb3LyzDGQvZ7VirNr20
xTKbBMhaPrH+KobJCkBdU7Aqmp94A1rnczOiaL10MYJPmRFeitHwFmbaoScu
p+lKQkEpnoKLq71Bt5OjVZ5ob7LMwVERVQoilXA2VQ3HGOiuFnA+aN1WZZzx
quu8pckNLQdPvgRO5wazjX9PUxB3Fpi9eXFkpFZiEY9reuccxkp96wKpqH2N
AdQ7tmnWGnZ17Quz95f0J3ZnjPTKV5Gh/QO5syj1thXlARyxYQg2pZlpKRiA
wGLChaY1tWHNMM5qOlBYwO1DW/blWEmZTJ/JSC5DPLOsmd1Xm643KIC56Srl
37QWctRfkkLT2WVpKLt+sdr1dGQSJ6t8l1c3EfkiT9tbRVJkHGBk5HJgfdI0
u9GjmIQB/j9G9/v72URVOAP9DODwfq66CbCEMq24ibso6Z0/IC1GpVDzHV9a
yjXeA2RdMVnDHQ3X2+CFT7HCv0R/ju0//iH9Ta20UnTd0SQL2ImV0fZyYkgJ
H2Nn6qo7kOMdrxLWNgWaFPx/rp0BsiaVNjUF1f2K9hgrztXp8J1DdRamtFPE
JtZm0gOGDLSs03pFR8GqcTK84tbpUAVsvHH8iI8olzEHiE6I5Y3xL5DNCvJl
jg0c4blZVhJcAZKgdn9+u13tsXIjYZGnbsuFxAzTjq3YbDaVAfLMDK0xKTyQ
pn9CKoBijoledQb5iNu3Daup9qiARZa3pf4uLo4wkK6dAIl4ItjoZqOVtKCL
+uHHFbAjTo53vBXozWQprLwYx1COlzEN2UZEht8Gl7EKzz1Q7j+18SsVN/FY
ZVflJRsa4jK7mhOaGAznsDaYBaY9iySYEreR+11r1fXTTH8v3UOhgfogE+iK
vdAKUtaWm6UV810C596IjyE/Wx1oZLK5DLkKp2Wkun1IOzOff0wNNUDkq+D2
iOLNPNs7+O0BheHHGJWfxQpW7tBStzaQ0ypfKnzlUHSzFl3LAZMQdXDKkL+H
JUZvV/R2M1FdMih+9Vcqmqo0PnR41N3jaF5yxquP8sx0no7Zv0QkI1u+iiME
vFgyfNb5KW20lhV2wFTlrK5IuY4RFf8NFTl0nrEeSkm0Oh5NqmJBSpw425mk
RVwiGzUm/QnV5rdNXL8jBIL0HVGveGZg2A/o95pwTyXXJM2/4hvOx7QnYEJH
MHstanS5LDShRCFoF+zpG7LHB2DTicpwDsXEs4xgD0guxSPtNWYrneH6P28a
zWK7K0NUYidIfmkOTlVFY+rJ82eYXHjIghv89NyKpQSPfbQUjDHhLs2OaWd4
QXNgetMe3cqVuzIw4iMVCDeuQi7rsadIyis+0QolB+QjyN+nfYuz9z+cYdXM
nA145QGnbjuvNehDlNTbmQfFToTYuv312/+aHhApSHVRiRS0o0p4b63muC4m
av/OSnEs99t053DGGAnuxrXsYe37t61GwQ7lWULa2oCJ36oWyV4ZELeAKqG9
jPuKpArpBtu3NzRHAEZdS4NLMqv2r4sLdCftCcPS2O63IuVzZaulaDYDlKGq
hMxH0eFvyTJGj3MhHdaF0QqjNiIV8Ci/ML0xhW643jnv8bB+fkAKqeAKQw5l
el9fVj660bAmeybFhz9h0SeaCtu55pZId7Wm7oVVCBETjAozSpaTyaOabDMe
hg5ApYrUKE1xthTX5MDQ4/ewxIJATgMw1giYBYVSVhI1d4jxPUy2rOb6C9ut
y8WoerCXH1k3L/zSSR94Arxyg07x4RMhmeb9fP8L8WwuD9SJcK/FptAkH8OL
MZ0KlrlQBPqgijUUrHGVRB7/nIynJXI7XtuXWY2GOh/F8/jPM2/79EHin97r
J8BhBDoRrSuh1ikYbRqp1DQ8q5dyGdOTHlzLuW1gC9tTP0vdiKIBH5sbsR6B
pyw1VjlQ2AFAuk3qyYa2y5krmtmvJFBj8B5H9dgeIrMvBKt/tItdV2xc9+i+
1V5uuTJeRJGZcAuGXNwR2+JHkgSx/4PMnzUttVO5Rp9OJtSRmuk9KFmknuYk
pC76vzJa4Bfmv6uPUQoZSBtRZS0wVvtzyisJLfmJNfzfPCuLF5OkDLlq/Za4
DCs+C4NNy4VlNUe6McVRvIskBgD9bSpdChbi3yI0SbD19gSD6Ykp5xNqvxyW
b6WJI8TQ1yNdclH2BLfrGsJ5uvQA/GcsmZKsSypD4LootNq0ZAT9UgtMD8LV
3srjWSiqbDnGqXtDi6z4IfhxC9cczgAZM92Jtvd0kebD3KEuDk2ceUoNgzUv
7RPlf1oF27lFlPP3rbYgTgqc2mFv2apXPkxAIOzHCor68rC05r5bg1c2Isvw
396mTQ1Qn1bVNHi/3iSDMrPmwNqS+d5aqwhU6YB5VPHVfooXRIAmRGtFzfCn
Q5Zh77Z5cjSl4cxBVFkeNmK2E6DIQKMmRz7zHEvbvIhR6DXHTRwxwwImBwPV
QYz4+5aW4IaO4jWjIi0P3fF19ZMaKcPMSI7hiA3WgDzIR6Q5TRQKa+fhwHYz
XpNj9xOubpzF2jw7ohRh6SnMtr2DerWb3NcuY2/8rnQl4QLieDwBFex+4eta
UyxsAQmNaV7D6llHIPhuBDlFmvEwOQeDu6JH9MwIknEMNMgktHRqn/SxngPE
Kp7t8gxTqVLPyJ0aiNH8zHPd5h7TZGE+eYaACqy/JG9iCD7B6QFcpFixKtE4
ujOS8zaUrTppvTY0UJperz1oheet0zMdJdv6AmA50Lk9rRO/haNQDvt5Q0G6
eUccI4wrAbqv/f2t975uJSD50rTQmNlri0yUMbfY9gn+pQx8YiXwFM2W5BE8
jwXlN62Gr5RO0b62bbXylG4R6vxivYxyWilMYsdWkMxHWZ7n+HSHnsEeLIVB
c+XBpRjBJx7awYpjbW2Rw/Fyx85muU6uwEB1xbiUL67tXRtTrO324Wx2DGdm
C/D5VLcijXniYHi0AKOl7vSB2c5dqXs7NdAHKQ/+Z4qW018qDEN6Vqvs984Y
XY3IaJTM4YuERG09V1OgODLoknLJsPWF0zv6Mn4xwo1B8XECsbQIA/m5kYkI
VsuF6IVXQUCPo0H0ddt3Lane+zMryX3T8HDpbMNEd3MDhlWNQfG4ypZSKIsQ
EzIEn6vPytvlf4Uzp9zPbrK1uLS36adtSb7hzo7ahnihya+rYdhB6q7X1o3m
aYZPjHbUPcGe8MW4ON4hOSBi2TM51iOiVv7F8MIzCx/l3s5ubLF4DYSktNrS
wzyb8kbT/ZLT5P+/+TZ1L0NIU62PtQHiyGa2DrJEJS4cfITntGhLffRHW+J5
LeEx91jBnSZx9iMEUxs59Kb0lw5AOwYwmHjy3Zm1R/QP8GMqHUia5HACDbyq
z7G0nzPVxY25KBdJAGK83c/Hqb7G7oBctjMeMqiv20tkDX7FqfKWZ6xkiya5
1elvCZc2LlfuwwNBDQfzJHWUREj2lyPW5QC2AoY+D1cIVJ790mY/uXYGCrL7
2Owr+0SVXquZ4b9LFkFBD9F9YJJ8UbDvBaUR8ARVRSiTGl7pCvbMTO/WosZC
QH+kCOOrnW0C8aMtcMBgGhLXexq3pIPgO3Slfv5u8KmGMV5JKAF5G8PjGpzf
M6j4nKAJC0+1H+RQ5lyrn/V4apusFUc2gY2HS6Je77XV2hS+kYS1jkW8YNro
u/BIrMPUrtuK1JTHMrYap+kuaAZfeGXTrAVEohJnNJKRgbT4pfOL5CPr0pOe
4Q19REBvQT8ottWeMEpwzd8GD/GLCnNx3mQtWmWO9gGHXHLmeMaV9D6pvi7p
VQRWmK1CXk3UwG+hrrVyUr44zQW9IR0KVEoaUXhFDuY5EVG43Aoaw36oOJzE
ttldWhnvRuf0+7+UWOpAkQve9R+8kDcmbSCnsbQU+5HZlX9fEPTIBlhaTfE2
+wLPW4mF8veeIw06wo6HKwE/pTireK2lQwi8isa/sbovP/n/C3/X73ANBkhy
jFO/qjl28dutJZ0OAfHo2qUNDo9pLZ9lNIPDYJ04FQ72t6G0w8Oqa9kcDM/c
FAefJw/l8D9AVjyFQs83HfuvFMugXnDU+ruFPQnU1FuzyPbNgvXX9ynEEGTq
WpqD/HX4vWt+bkxa1uaXPPE5a7hPq4eTKozsozvqTsNaKgj/b3globwy9dAz
VsOF1U55whev5GtorzfHeM6zwwYzf2nDgfssKrqKV9jBzoXJSd0qYiVqUUk7
Ef0X8bWHHnaeFJw3bxZvZhE5Qn5fxPi3Y0DeUh8CxEMFvTaGmukjrtcfk8rK
3kIQ1aZWX7JZ594LzOax6tdBTXndrvLFQCmg956vCVWijM7nOKwgbfISqVAD
L//KxWssHZJ6PhsJMD0qvVPeaLJoT6kZM9wEU30OA6YsOUNa7tdWLduv47HE
dFWEsJy6bIx87NSkI1lDgANoYQpJoSgJSjiQvkNrw+IudvGMZl2MOeoGPEl8
K46PHCCGWEVwSSVj5jto2uaad0bVy18yfkvMfXqQJWRPFVSjqjSx6MeWzECu
Mly+K/1eNRAyLqiLv/yCUPR/jzuPAjPX1Oohfd6XWGJpszF/T4BnHukTicP2
oQb3PfO7aagHsagikJPkbYoXfJVN/mm1W2PQ+TSGi8Dd5gjWCcYJbZEfzatv
K7ufTmMXkXbmrE0kg64pwGfiy1c30qkujQw8awZlmdWvdcdo5FE7h4zNKBvL
TnN7sZm1XoKltWeTZItQmNX4QNC2mS8fVkWyVSugtiIrxgDuJ29EF1FYxy8S
bZJ49i1I354BBU8PQRzlDWazzXu00MwE0QrL4CAnE7Fd0SBLJNy2KA8Y2zqH
BJrEl5/etj3ZrWTVNXd/B+710cG9XFApF8Q+hh2jE8NJYkK2oDjD6j6omVPo
kcHQNyAnhfOYCDAB65rYtEp5gRz54GKL8f+Dg99XruEoPvNNvJfliE5Gseir
haWJ0qQ1BpTupO2gB8N3i7w85s3QjLKMJIOKf/6udm8R6ZhvBB93EundmJRY
D7V4BQF87SO4tR7ANipoevdvNUSBeppW226YGN0MTp80PPeJ3J7qTeb2oYV4
mUReRszX9JtyfHcNjBWdaAS7E88J0J685c6mMxwNyE1fEECT7Si6CRiszTci
jYiPMK2L9hBKVk6Q93H5+drTxe9XvpB9ZiSEt2GRANhfPk0144CMu7oVr498
fTnSHoRcJo9MA2ATnGKx7Q+QL7f2OwGeQeemkRGTm4Qv7AmEiztgOQ5MkxGo
3+AwtafX+BMPGrUGFpgjx+0Daf7lojurVPx4Z33e4Yw7ePCUtDc0qEcJK672
ZMe3TxtKPKDsNiRFNU3346vKxQQHCw97Ch5Zpsevm3c6uRgkjMgxNc3smmud
4UX6UBYlXdXwh3NEBAJvLpaaA2eKo/4sAy1tD3kYyqUmmPwBhXpTdjkyFuVD
4nyxteat8yEEJ5+KnZRjKfJogXNeBofU6+FDvFs211etcYbQwdewpL/4bkBd
aDxWqeTv9o/jrioPKTL7/5opfGuAQNquj41a61TVzTnpiJtfTdnTosLQX4RI
8cyh01Ryo9/GjM7zFds9oin9Q6E+MfwfO1mP+Kdg99yU3IzBgyDiyoXMCFqO
3tIfEjHM98YkUquuIfWwS0GdI6M8gbpYZNcQxhclF3R/6oh/Gwg2wcoxQF61
9JsRea9Mn0rnH/b2rjLdrSsyTVRSvAlpp/+I4vFXUQq6fzeyODKk53qmxImh
4koMt+B18JMrKxh3mn/s8M3l/Ur8U+vj0XbaA21+uT2BWysC+aNeFCcJuPnd
C9OJSNhpxT1tI0qsmp2W4QGdryksjl8u0V/1rkpPdmFGBWoGjpxCmJYK5rRO
Om9fPiteb0cja3Kdiidtg6ULU+0+H9eSYEsVac/SsoL07pHxTFM0NLrVs8Xv
NA54deguwE/eB/6h5Gq1IAQmq9Vm7AlAjxccqSGUpjUsPGMbQfb9PJ/TYX2h
ElG/TSiFOGZYcQx3sbC8bPSKwUfPMRfFJq9NmHC/N/ny0mh+n8jQKl6jx3od
ph4jkeNlILhW5aFs8fdUibOTEFLEY61JVrq88p3KTj9j0IudRDc14GQCKF2v
ySnrbRvlegIgLl2HQaqPhWxwUXp59lLRtqmWSYknJ8QIFq5NiawnbNn3xuVY
xPSAlkae4Q8NJO63pbe4nGo4npoXTDRhovre7XE9m6o3fcZTaF9N3U5wqYTu
xQMCBvl4qMMgx87T/6PWgunu8hpKUKSmogUKOOM9nfNwHYc8WtGkSp1KCx04
/+YCPl1c8C7X7ZSWh+GdEP9TqnyABk0FwHXzVxrpEli0+Mw37npy6hipHvXj
26Ow/YfNbzNaOUtbef96zz3Izw/y1C/Dr4iBLMY+jN0EIuzKSpfLr73SjwKf
inxXGIuuiYSX91TGJWGYpxYT3Hpp8QYotBXzDFzV0kUEWSm5aGW5TW3Ncjr6
BccqwaRI4LYGvdcImnnOi6CSppLyelH2BqDfLy9pTVuIsbCmXQdqz36Y4JA+
TI5qXGquxC8gQ/hfkoRcT2f9MEoRr5ayq7CkOlmc9wRe/el1/3GTZoDmgcQt
eBYNDWytXJUm1WgYwvn3wvNZ2omTzkz+oD/qsldo7cVlGmNOngSdu1yCvM/g
ebfV+gxDtqfbXuWAQH8luJrqWkHn0KvLYewWPabv6H8LR7CW5U7r7kZ3GnSX
Tj6i1nGL8nFUPsLBAN147cEaGgpC/8AWLbtxij1hRcU+kWlezmS9IYO8Z934
qp/l1RwDLKcP8CoAOtwNnXnehpgCrZe+tXdqsx5sxmVye11PdiKZ4Tk1eDNF
Dr0z+fS0JGF1vP7gzSDj4b8mqYlcm8nznzsYFh9eHh3CXao5/QZKeE+E6K+D
VH4RUbp7qg8Yo9AX3V9ZtMiNU1pYTbzakXLET2gAVkLKabGUR1QToMGYPw80
2Fn6uQAlpoxJFoJ57nrDF7jOvP+fCKwZXe8lfrfrmUMKLplvr4Bw0nEDoS3m
N/7/XWm+81SAhCnPfUZxrkdUsXYOY4mF9Uj0X5jzmbPaAf93l3p00+E6YduL
EwsqR5616oxR9HzgNsjHonFZjuMYHxPIatJPGMJ48nOma7eJJxCEqkVQvKRL
sU7+Tu1e6nKskC4lze3+fFQbU3Lfn+gM6/mIlVZQ9HeGo1xyQ5gc3x47OJOG
vN4HK+G7WyXcaH44UiLfxZ5cOGJpyWUNtnVNNaZME6qEsxqC6F+j1lrSDUot
UK1iVmKIXrB3bDkI59FQa2MQ/v46Pnogct4M8YjKWiqcKYsvSZI7qbLSikME
7eBSyp4xPyKVv8afg5ct+GZEJgIoh30S8HZt9JsrAP1atNs2kFiN4ReZWWQT
Lak7nhOmm8vvhPiaiTMQHYzeMssD0KggdsynhpjCfwdHn81/Ath/W8CAdpaQ
JcK1OPBu6UOJ8LEoRSE9oqSh4CmfSWOBWIpiQlXAfqnD4SchWWPYgbJD8Iq2
Qou2/CA6I+7XSE+Oj6J/nBRniY5vZ5Mn3pe+ln3JbbKXDEuLP1pWfjc48C60
GL3S5LFr0dWDCkaWlDTFGp0+pqz3e9glOd1k1rnDNZVv64NTGm0XZKGPobt+
iFtockKGztx2a4IVFkutm/ZZ2REweBCN0JzRqWvjrQo9mu+GuxpGDxRoDzub
//v/+BBoPBAqNZqukcIvEExT4FmzWK0OIMHXbyjX0CwujVnHZkBv9nlpa5TZ
xQjJ6wX7oVVRxMYhhagMw8YK4PlhKvMSSI47QxmzP7xA4IePJjCp753clovK
G4T9KbRjdWdvcyb67FjkxYlzDa5R0BpwcFHb3JKwuepBh6meXu14KlMLR3+z
+zQCGCVLl6sxA++TgYTwAo9NYp2+Ep7NcnRic8l+55FCXdZM3trIUDZzNTKh
FD7UnFMulif/ZVe9y6RB2c1TC0jxJKCkSZBoYA7JKQ2M30nvMT+V6tYKiVT2
Lok6rUAszwswL5f7bbc4cmef1X2CkUKMMlIlEv35CiT/zWKBDpvTpseYTq4l
Q7CjeYeZ6KBYpuUYE+5touhg0jq5FO1T6DAwcCia9LxCWEMyl+dscJe3LxNP
wkr368BvuT+VMNCNgJbR5at6YOAjLd3hUlbQ4fXDMm8iG5eSHpDWgNL9Yqmv
0JW0qCc27SHCySTtf1Z79NtXrbp9MPafXxDfUfsp5b00drNYTI8k4QzgtIA1
ha4fcBZpzOG8zkGuyLCQL2khZLr8J1J0tniVt0JXHKnJ4hmhcj5sXX1Krbf1
te8sE/072EkSFcoVTenPhJKFN3BKiTrn5PKj8t+gPhjQpWLG98KL9MBfxMGi
EQHzjOK3RFnU7JzAjnJYUZi5lf1dyR/r5atTgIOfJnaQ54VMTMncTd+craPo
Ltf2rGe44JjKogWHzwbt6TLfhg1KgMOHhBLFSogsvlh6YtsE9Lgs581qy4oi
uw6qa+yXEz0fCYKxtb/kl43ftHw5PqlWxiMC7XoFzB3NZsoGENNkH2OjrhZo
1FYIAFlMB3mEgKQLqp3Z9OykLEcyXu7jS0qsAo2D1aD4ZjpPoP/f/bsSCwG8
xfp6ipfGEvN7PnkPIg6rU5vqqKjT+yn++smnvMO1iorm9nQOt1PooG1RPXmx
6LRXmW/N2WkrkzCMPozbVCmdPfUDzgRoZ1co7fGTCyiZjhcq/GYX7FDqC7oW
17xigd+kXKeQVhT+znowHuzGMSRQ4b2s4W/Rg21ygVArwbTAz8RdLJwX+VQO
FL3MpPnzWwG5clTiWB/aBq754YUMiSt3gs3hJpRkzKgowhPvNsm7HVA/9JeP
xI1MVXMuQiUXPyXwI65EGI62x5KJ4BOPEBHnK/hMv5ZyFgYuQFFeHvfYn923
L6pf/8VlCOSIh555cpN92qaIINLxS/7tT2m/x6nCVlCfHKg0VY988gBg7YFt
s91QrG/b/Ll0uwUNYgOC4dJKbQL9rHFyQu8HrrKoFhrFVSPtuYD5wb8uj8/p
75o9nPgLqfK6j1s/ZjdE7+P5SdXAn05Pykcq87HKmWfFisygvulX07chdac8
AQZIleIGn4G3sn7iBGIh0es7Dn4q8E8PB1YCdcPFRvQCLKJw4P804W3pvuMn
dS4hCwByD/q73FyMFX5A5IceeXEz0+yAKx7KTUhRMmbl4e4aczLm729gU350
e0zn1PdJAZlkRqrCxDtzktM0WfxKzoG5yjMDfcJjX02ouI7VT5ZNDkq+IdUN
VA+cEB9yicRZI5Mc7rq/jUQ53sC3bkmPbaBVp9GbD39tbH+HSVoxh7DD7V1/
o9PIj1EeeJcxZBmne1OFR2BhKZTZc14cbd35wORvqXlOqbbMsLMWAe9b1l1Z
HRZLc5DpaV3+jJTu3+ptMD0vWCfDsMELTXIUM2iNMI4GOex05qc+zmDytT/b
F7qmZxDv2ZmAYqI3C1c67yk3b9tJGKPqXiQI0O8LQMw8RV9ztWyHmIjIhU4N
uzwrqOSTI0YfO7L7Vj+azxVW/qoCy9e+3a7MxTU0aK0iZa4Gw8wetB0Dx3TJ
hB6cR8Lvmwbs3jS26pL+zeX6kLBmenqSfjuJ7vuWUwW6FY5qQl8qo4rlw5vs
Q23iTTxyF9MdIUUtPUjeN+4Js6oPYfLelyBcyRAYfvNJkbXWpyKq4lyjoizq
XugyB4QuHDDYMX2GJLeVlECLp2cbNzUuZLtvaQtI6mMEpThu0ud6XXGWfpiC
3a71FR8yBUvsSx6Ynq/KTSeDmJIJLJe8pvvGJKY2kslwOqHmbLQK4uJe/8Lu
2+eDLXJ4N6wNXzJcdbtFCDv7biNCuDjRp8mHzmEIcDf8RfibdYbU0iI00Qh3
M3d75w5baSAp2/qH+jPoN6YU9Qv1ylEqgbkdIR5bmM4+/0dG8ywRAeg7xuye
+9oGi1hX2e5Rw+sQv5llju6Qr5j6kRQ+j4arOqLPvDJQBqulGFSzKdhJIgzL
M/919AGM3/lHDaBnW3mOszOKJf50PgKKaZPuVN77Huz3rvhUUbwPz5ibbRR+
oS5syW+EYkT9P/TLf6oSKV9BKrG7JnByyaRThv6Lt3zVWOumlVA+Jchv+pcN
PjQkBdOZevfktbsF4zsRDOcPTBHg5NjEYmR9trvqcGCvqYNS9VPlZ0zEUUrD
PpE9ZqFJobS4d6v0fBpgeChPEEkeWWm3/ZDZulQ1tJgkZ92KfolMeKuGV+Pl
rDOEVrVXVcUwDdT+l8heD7Uzvr660NCA1F2cHiEDreBBFGKZpIBAQFtCPByW
b1uuaLAgH4c0MtVL9xDYfhjHBTNMTXapJxNImFA1epRh+y6uw74cpuAwGoPN
Iwgx2wMRHiYWYlTDm1Op5ZPGiWgmssWb801+GfVn3Fvb8KMt7tK5cKu+NBYA
RNW7sW3KJus4qSC4mxY3A2dTvnXCWNPvcZVOpo5V/mb6Iih2WAL+45gB9LDu
5ezm3xBD/rQP7KnAMxPoR3kuHA6E51R9UKYYIuTS05VFKWJ0usOkt5owbcTL
bRhiE9gjt4MJCjbpHue/Al3rsBmfNwQy1j94wn4jwgsU+7HO9df1g1UQk+S2
8a5K9UPS0CrRm0EC56vMlK0xxrf+LJn4Jpd5yUrNMEVRY6nPJokxE8TVINqW
3kWkVoWMqHNRoGs/l3QRqLJYhg9pTM/TV8gQtpjySV8xbIIEL5KCi2LLI52M
uSF5rD9aYft/4aROvOnUckUheCuy+k9tY5qIvK+Exfwh5KheN8TEa7jWlcoy
B4hGdASZM2uq4yr36xDNxYP9OzRMX1GXiI/eNjOSqbISFdo6SXPrmobvU8Ip
uT9Kd56YzHcF7GyoCkvh26o82KJAqJrjnUjUF2QmNzmSWJKx/PBB0mKgxadj
aXNGeERLG/5KZlGLZrDcD8BSs3vYj9+2sJthwILHnBbNGlm3ugg8F/Fxi9Sg
anO2jn9GPRftTmI9rKfWsGoNLFOSoeUoSDuBL5pVz0hHObTYqmcyXQ9fOnlq
VnKCHHP+USWxYXXiHAdZ91lh1mehDZ1E+ZlKZwKgssd3wHm+I59h/oS1pFuf
GTyiVIX2FGCSKHx5Dv2v6/cap44GXWkSPqqbFBQXwfHpWeezF2fC3A4GAbxP
T5F88+qmd2dtr/XKQoSuBeylqoF1gyN5zn3u1alQ/3I4Rlp+1EjnfwjG5IVx
P99InmYGVp7FoFnHKXOASe4TXIaTKkgacJHv9bYAW8AK2bMpmyB0rvKNN0iv
YkB/sZNisZ3Id6mvdlTdmfjSbWfmdNboOn/AEv7xP/3hvwU7ziM9JUhiljmV
QFvHrUZp7goxmFrXpskPnP4eQrQC0ppFMDjMSgJ2EcEHaLcjdk69k/aBLejV
H99Uht1hbd+yYRTNKkS9ORi0y0itA45c7tq4bblfV2Af15I1gcbduXs6uiB7
Q52rYbKvdh3WypCnpjkUgSgLuQGVH70UA/3SNj5A2VnQgjSWb6Fq2s0bN2Tq
3z8F7QskqEOD3Kq2AHtnKc5i40SRHEfTkyG14TA0jnOws55yPREupbVAEn11
ZDv6+005BVjQsI59o++QFOSBmXIsllxY4C9QpLl6Ur3CjU/o4VeLEkoCl3D/
gligGRHOFff+z36pKfe4r1uEi9/l2bShqMhyr9/O9ZTEpWltrSq3ZhQJI6G9
5dz90OLLcpXBGL/3o7JjaqysdpAoJYw6mh1UyfEUh7iPAeV0rLsSFTY+G0u9
Zn8f9ZDwPKm+2Xs8+/sed+WQPF2dHY+hpfPqX4kbydUC1Dgih5rd80959KjD
Fr6R/fKEeiRSpHUAS8gHIchbvwqrE0GgbQ0WCSNAiTM+u668bktX2zS5V/cp
u8GSsiplX5e59ihDJqSUjxixgJVUZbS7rdyHRr9FfktsbA8ebyQz3E3XseD4
DVhRQeLG3EkFKkg+ktLA4zEqsYQfSWgXmubKA2rtOBoiwiz//4SvvczqpeMt
9LBMfIcGc3TTCabhmGwzP5+c643WZ6H9HPKeXtQL9Yzqe5G6EZ124siCt6Mu
KVeCHWPm1q24uvGKYg9nbjSFI8ObeaxZBler+mks5ro20yv/2+NcGHeDH9U5
8O+2EtHsG9R2+HzdxFBoxjk6zZaX6gHPxBei7hCUwcQwW6uqeTGM9lyvOzSy
PPy78ToDnxZt9bCakanI6gmmAdElzwsqpYRcqn0UEqSJI4J+mBFX+TJuGFgx
QOdUAW0WgYAGWj55cYrIOOfqpf0cjgBO1/MHcvcrtY/LA51R04/v6jG1e7JD
TAX4WrGjlISKJfQxXyYjiSULI0dirbIyfMA+oGvhd+Xt4KXWSMLxHPVq9JjQ
DXCeNHGLF0Vx+JkdKWkLht7aVRyk0NciFpkQm+M76OHOOD1iqwpOrMY3HfKv
uFwLl+R2xd/aZ1GmG6zjsqh4Q0OpQq0EdIppM3vJo57YRm98110QUiYTxfbN
nK9ayOY805MIwFa9ZRYymolM7m+EbLFAP51xxbogm21Wt+7JQTbI7safvOS5
kQWx54KCqaVppiHmu3r24S5+VMPu9xvBGwpa66smRTF2UF++FTph7so4x7nD
NnPzjQoa0TWq3F08OA210MZxcGNAx/Di4NHJiEm12dw7lKMoZL9Oa/BJluU3
nLOlFNEjxo7Mfj+QxIsEOhaBPBu1ODGsYtiipeR+uTEcYigmKJu34zikNJej
Lb4EEqr1srl/2LL8/RhFora+qPQIwrQ1jajhbYuAL3lC1zBo1eJj+jhAdrWl
Mso+7RgX5+jGsEtmnZXAIJd4dsoI3AhkvmpacIT/AoJMi1xS6LuKSqMSOmWY
XngJrG80vCerz02x2aptbPcXvIWTiCLbUUhxTaH44XtbDKT/Baliyp8nCAbT
9tZG3Qdm0CY4Lpghjmq9W+JjFFsJfdxkxVHnfk00Nj1j5RdEzQ5448+E6eaR
UWM2OVEN1j5lIMWoAi8ZNcP/UQis10lUrfYzIr3YyFb5kM4cdOp1of6pdSFD
hqbuu+n1ssVBF3ZQGAWUxr4pxSz9PXrJ+VP3kriGVkMkxc3jxf8LOsIqhbx2
I5ZafGZnxH+AtsjNPbCBtgAdCXQ3n+yI9LHQd5LA9E/PIoqQOcmDTia4FDNF
tNbfSvCGiq/65iwkTBga7LCHN0x4LO1MV5XcIylhpL6WQVHPk1JOpm0ZDdAO
nYSsGaVKLXX32yZJoSn5hcqUdUtsvql79JDAoURST3DyagjmaVb+8ugXDQ9m
8gSLQfjXO0erIW4WrqV1rvpxmHo4J5Hq6Dayu7pdjQLKUBG/NaIubq7IO9KJ
667j2eUr4lo8timPZwb/GCcZTnIQhJcUJbo8H6EpGnz/iTg5Ku3CGJkNSWHb
1zYDfQUvafR3JcX9f/YYkKvQnA54YycG84Eplx8x42SZzloeWztd1AGmJNtp
3FTT9F3ZAx+NpzzZNngC2jIuq+B/ATItG5Zsq0N8V6G6tIVsyUuS+zGo8gZC
awPk7hB/6otEpivrF8iYOEWvuNl8nO5xfE18RDY41e6mhZGCs19ffAJ5r/7C
U9aO33gAyXY82YkS7rilDGfcuN0j9TXuvqNAPb9ikd8q4QIGZ6NBXjhCvu20
cvNnobf/4W21oBL4mxN/5vr3H05KPKkBZK4wb82uj/uuxZlUze9/QZGtF5G1
eVWWpdBXo99p3i18+IkZwpg0G4jC94qbfc7Mq9dHSeUqotpyMrRQkV0lmIWh
mpIokXvVHOglyPpCks6OBDLmTSy/KKElZ8ldR0yHt5Qu8uRhi14y7Si8wmZv
jUt5wyKnImwfP5Siq9HDnTFpQtAZjdYDKdfOcJWL6MVA9mqiKsiIzjY6/Rrb
xbz85ukOsdnzl+6XRdGTcrKfZsylO71Ggj9A7UCh5GWFy2Jmams0shuJbKIV
ybFDIhejZAkSDXISkCOKOT8gAW7r/cW3wiE5yohBmcIPm+tUOIshDf0ZbZsF
Wz4M2tvEy6pxu7SAVwn7hNrP9b6h66CvmnGstf54XIAvbL1UUT8eyNSzgUjj
sBztYfw5GyGQlR3hFqV2syL+7DbYlqFsGxv57b/CpCRNBD4Ko0zaUIxcbGrL
Ddbj/pMiwXR6l1kiGujfv2/4DMWXXx4bAMOLD4af3KVT+By5v2YR25ZfLGQ7
Phe6yEVuuhH/nCv5S7hSWq1hv/mcZw5/beqxe+af4HRb5alj5YETbGddvgkY
mwHpdD90K6SaYQgl0UjSr1ZJmBtU+zY9W1c/6o1RSPvu5W0B/vSBa1acYN5W
EMh5T10/YmcvXRbJRBTAC55lrRZVWmNCLYYV1+tVQDKhebLUY68cflukx7oH
qvjM3ry1sgvmO7p/1FkvMbycg8DheqJaxNBVl6yymBO6nHYB4/mlB1qtTkOj
ysniLuXHdm6UEWaikpYKM1UEIMN5TtZwlg6JvoDj2WFCchVTBvxFUfxs+fps
pP3S3FnSDp3Tp6lg2AXuV4+EL/eMocY2iMCQ/h2wu6rKsPFUozRrmDAeNagS
/QsCbAzBK570RS7fVT4JSxcIFYFqNgEbscy3jukU9sfgth9/0T+JU6xYdBXy
x+1hEwLX3FTBNORiedaFPF0dDNi+Y/MbZO03pezmwr44NUWRl4CNyIvSoSEw
R3ZTUSLyy0K3mkme9frig+3TBGOAAEgmbf3SDcHqasgaUCbt1xp6ie3/fEfS
FKiewA6S80/He1AK5kBwj0PT9+X/Pn3y0vqVEoW/3nnvsdpNj85CtcvSfFyO
/TTm5bWRFM/WqS3T4e7r4vY05QyOPnCvx7JpRRpK/Rpkx+dlPkL2gvz+NnOX
WI4ft/8P4IfPNKSNq5XoWyq5j7rsmUfp3/M5JGzasWiqlgGCYsoTcjxkl/wF
oiWm01wagaoTwK2mwpKMfrVcnYTnkNyWHRXM4jXGZIver8NOowEJR3zNQj8E
jjXqyme6v6z13yWBLQU+ZWabYHWdVwR45hZ5Q2niT9ZfS7FSmau4rWm03Gc6
QiwnLKNyX4xnF4o8NJBm3fAowv3avyWD9n4/2dzzpUdRBXSrivAaKY6EShdP
COG3HvXVWFf4/dt23r8rcP+/Uzcdd2X9h5hRTTNnW4LBqymUWv1ifIAR2bOY
ge8MPJldIVVx5KBgVieda8hDIQ3ylRF4UleufcDp05t9tNHGc0SvsI2kZmCD
TGCoHnTdi9uLgJlKWuDu9B3tF7WyBGyN+Nh7NJcJgq7WsuuBaQ05xalDspzy
7w1XyUx0Vdde+PZPOLC2hUv0eyxgvSzAkv+cuKSGIsho/MT8RmUiobuvfjNf
n5Hxww0CFlZ8h4ncgDKFEwYPoIHCT4tnW6X+kmk5tellN97fip+CT/tK2IPN
fd6rwGIIgqzmWWmRgo95C0eUQOxcFxdn7nXIZ1OnEz9E4VkZkTUghQ/3qEnG
VpMju1/OMJYqlmjphRGV+If0u9P/gyMIMHu2PH34CdsnvsiDqPRnVMREy3Gm
TesxNCY47YLnyQt+px1DOXSKHZdHkpLn+wtugR1L5Li2RwjZ5TsXYnGQFxAT
9UU3rIDJfWAQas58e02bkz6i8CK8FRYQe1n3x2RtPK1GMg0gB0UjmaZBxvu+
mNer1p7VFBhD9rZa7PUal4Cs8vzUgv//EE1pH0oH68uKj7jwQ1QkPusIwjr9
0L91AtQI+f/uY3thIBbErk9tQq+Ojy8fP8Im7W64D8KiihzZhd8vwbsycNJz
0L61aPO2vSlT4pFPAsntYRzOaTrVuE7i2uZpIy+CdBUy639kcW7OC9bwmvfZ
xVGW9KbTo4koW3xrv1RF4M0Q45NLqVgllcXOHNgUKV64xuEF1ZEOGlF6lbsa
P77N7GXj/zGJJ+D6gc57cyYFz4WFZ5yu9/VALcIC9yusNfD4USjb325vU4+9
mHm5cc6jEwPWd1IqvmxuRo2/S91vqilNwqixnrsFnv6UBcyHJR06p1Xe3/fP
+gjCkwslsedAxp22H7MbbwR/P+gboWHLYt3PVSiVjtHOF/F10SDOIIN6y5tH
t+d4eOODut4TU78ifF0oMvUhiSd7wR9NiIrmVJAE1OIbDmGso/y9WDnu4BJR
nLmaf9Xi84DNXRI8IcirvOZBOALrXzifjpiup1W/iSyeD/lfh6BiQhvZRQ+i
CoplzwPrs2tg7sVtuyh4306Fhsl8tcb4ANxTGf5qEOJIFsOQXvdU7TKUmzbm
YKtl5KUvNntWf1FQDFJuO5+tmmrYmQGw+kXfg1Hx4ZgavFK1AtCiIKYPIlw1
3d32nTSkiWSPBo112+wyA1w3wtoAe3Q53M5dZc2QXogGb9pzhqXosucz/y/x
8Cl8+MvpPCiBcFOUAaIYTOL/kcJt0lZ3j06ZyYWy4AaWk2cDhJtWQb64DZU1
fGalbVC5KohA38Fp4BXgVh0mqCOkAM1ZYqlBvX/OiMHdfDEduuZkUDTY45xU
rspKqxE5V5IEZoGFe/RChVtYBNm0Xdy6JMBiY2EqbZff65NqFVDhjMA0IUpw
BOM8lSqMl5OWAQZu2jdq9MUTRtzNihAdqKFFd59gheo9Plq6Ju2/WlhdXr+o
0RhKHcJscQO1bfKovOgnppfU0JAQCwoJcA1AS4AWKRqfow0KYGp3pFa35qIM
hgoOuOFrwp+q/a8Ld7iJAsOVXHC64yQG0IsGFlN4Jk5khRMYj/8PV7AADrNR
kupHUSkeK3J4+7o39oNtfAnBml5Jbjf++shvds7XGMZTRfVojqz1oip4mM2M
DftpRMrg4T4bImBWDkH9n++BwPvzTWoSn9T/yOVHFXhDt6evW6qxO31nn1QN
3YZTv4sS2qowKylI5xTWFVhogbndlWUB4DL31TRuRpAss/ZL0XYXLPqGlbOX
tYpcKsWpK/GFZgWb7jEgbSb6U1uhf9MEUW6PiDU0vW/wm2lBofXXeWidjGaQ
+QY/OCv4VMP02bzF//riCEoV/Cn7r4xwNltQPovAKa1JVfrE1AzW4CaJkuFW
VBc+e3r0oWw1E9iTAWYrOzWWK52dFVxrTFaHEE8RFbd5l+LAPOhNtmqZNHyC
Wo0xhhRluplLr9vndvfQhe+nuC48wsG97L9v/jkHZXqLuHaxKmdevWBM7Zcz
s/4N1/v8pAu0P9eFkybjUIz6bs0XuOqFi5WKZbS/gJBJTQQfz9QEVGVLnsMF
sEq4uZy4ghRqUHIYtAMzkexk+wz0W9hYS/q4kGf0/U24BFZ0/IuOgNqYRLkE
cPyOl8dhiZhzxZl6QdUNPgj4z6nLfW7+KcpP3ib6UteCn8v4vAsPID+uTGXP
AlpbHO9apZa5mApZZ2d0mMGqA22zTIvXWGWdu139bOT75PPHs2J+kih9/VFA
qsY7r5j0do2yKAgCo+9cwbdM8OJhD5+ZjuETv1XODsh+o6LDx5GrWhpz5UzH
+lmZCduA9RgVfzfbM5kcjdUjV50sM7jwCNh/7QP71i40+kJ8NxZodLw/dGYO
sCuVpFlyZhNiuNKejVQqzL4k7Bf6g93TtSdAnkEuvUdtqIGd/b64UKU8RDH2
FL9YzQrssE59pWNbNVOmjazgAk+WmwEiYt3uGMpTvUlfhb8pAvPKIUZp1tjo
g27fgd2J0K3HR8d6KNWGy96QjbeZ/Qn+VjBI1UfXCLQS+v73LEociiLW8a16
DYPbL+NvNiexkw+Da7/PliIAAZwT5YUdBcs/TPzc/cQVlCw9+lSf4Y6iNmZf
xiESt+a0QjK8VxGxpNZULwTW/roWmnmjKatuhuucHszmHu/RgMZMHvK8Hp1s
ME1jv9X3aBpkYdnJ8pR9XuXJH48yFtXcyfQ8LqM6YIFbLADZKb3LKw2Gtpa4
0Ub6Z2y0SClb8tY4Goc5fRV8CAaJ0SMZ660tGE/V2h2FUfS2c+yeLT3Ys1Yy
tshnA5C1+4TsLqppRWytj121TVXWASqZWFrDg/VjnrrlDwNxutUGgt5su8kq
aLRimkrwa7hedp0n+ZHdM2ZqaboHMZUMojr3UJBL316nGk7xTSS1D7F5Ib8C
E2GMeXoCz+p1FL1w4c7F3MPja+H2jmCNPL6F2agQR4p607CeSguA009JKaTs
IVezFmJV+ZxLPI8CQUy8Vn3bD3TI7ut7ZgU19t/zo+PsaPiCrzfB/RCUnNmS
NN3lnDpDkYX7EXrgVZQ0z/CMSvIjtDeW8vIbApg5ExkoHvUPT12AfWq/wrSX
FgxCSEhuVbrUiG2qZUq0/8Tzzx7cZTT9hrwad/+LJ560ggbekEKeDfySjjCB
EKZ9tG/Jd+AmoAxYpHeamkxih2MR+IsIDkxSJQf4j4bWOJILQyDMtrCLuWsN
q8Cp85Npe6YqtldZNeLVtdH5liI/aJAvsbPzyKkkJ1AcXs/rIeYbneQ/kmZ4
vNxRo/pS/Mws9dtYP72HCJb6k7JgtInECZT/2k1+frAL0hoVJNtS+yrondyf
nmyr6jsoPSdNjIfxHd1+e8is/hUPnZwpaTOTqoddA22lM+IyAa66fWcA420w
iEyX7ezolPcWM1L9ltlohx4/+5/PiY9qc23PdyjVAFU6guDxSynzocrQ1GRr
UNcwrVoTP7sg/kIcg1lLpzAoNvjRfJx5CXTPEnC/gmNuYu3kkg/YfMoLRi72
kt/rFZYKsEaY7ncyyE7z3slhQduPQyREpd+YrNQopLYoj4qXb/wT+ctLB1KE
u/DOcvH/DbnQsyohDSmUZyiOkb87Sb4vJ5F+3wUuxBlUDW68JZz6difEvKM2
FVpJ7L6OK5fbpLbpM284hXJNIYy+thlsbPVrwXUO6x3hy436c4DUFAnXA9r7
t28fAvwKf5li6Ok9Vv+vTuMQch5RQ6JGGutbuGe5+tCTWoqqAbkEEjJuBRcZ
jlZkRFUes+R21vrl3HtXzqXYgdR97HnjleFu+ItN8JCAN166rN0q2mKahUnU
JjbaVbmTx97fBeeMUbF8i9e29ITifMV6+u1m+OQ3TRMvQCX1B4pRGo1I3DS5
D6HOleSQB7i5BfxP8bdFg8c+sFUd0wBOoroFsdt2sXmlUoI6HG3KLojVgwYd
YRrSXkBuLQ9tfZsrK8dVYwsCTjHn72eF/dDHnTVfZFxVj5uvnl8RT8bDuqcT
bd2cd/ZxAsmuCCLZzssTpBx1ROR1uy7zmnlSRtyfSFueR7Q3lxtBVRWsbfG4
bHW7+Q1PfMAH+pscRILMIhfYFYmFgfx335oPbJio9ZMNhxFbkd17FWe5LQzQ
UqNFa518SiUGfWVyMhwjSITShwEgQrWrux2S4Ix2vo6LhL29NzAVURk+tgf5
uh1IYQ4hTmEEQ933+NZ/LGDejmLrj852IieUMma8jaP0bD+bDIyK8mg/S/nK
gb4NJcA+oHvUNjkf84+uN3qhEYlBX4ajWleVexIsYhbRjlrZRBlUQA04J1Gv
RLvsA9EVscMKPiIt/rzftwoJp6nOykF72DxXHuBeGJovJ6AqW7V1KsXSEr5q
xj6NbSxfiL4KAp280gDh6D6PkwsSVpzp+5Pj0/Yix7OS78J7ZkwWSk1SMJsV
ZNQ5QVVkZgqmVpVZ3TsfxG0ZhpvxYwUD0JWt7DQ7Iif/vVjRD84ZAS476c5t
dF2ZioV6FypIDQaYoB+DzaIPLz1R6OttUy8Ysn4zhjeSdL8hY9zmSh1mGpBk
UaR1j2U13SBfeZ+1IgKqson1D2fC8tPvofMvHqASgPkyb6yjHUp+96PSeBfU
uuoJ/Qx45ROhKQDjdiD/ov480e0J20QH1FuONUKn+lKFbpRbJKm5b0aGbUXn
o4t/zo0JHDnNUV2iT5x8xTx350j46aaNxbAPvO8rB2wJBNTsBKyvgPN1OHtF
kPkJ8WmR8hvXJqdHC9bguRa09EhsMlVJ4EkCHHx6q3FYGXYFG5Gkvg/03XOU
eUQzz09nYKaDL0XOcUcKufN7gZiAW0oj+raAJmLzB4K3nQsM5Slq1xR+4qjV
0G3/7C3dXxcuwaIKiSx4QzWDqDsuX1M8ghHC8J/yUmmPWJ1z7TtjFnEnoI6d
C4KfArWM0J4Vy/llIFjx5sjQlFBon52aDIWJl/h15oGyMvBE0Op8ar0ogNQL
7U8+ElURV69RzEfTKeIvI/Mv/3VE6K3VpwYe0EfB+nz8UVsjy+kDXMTpUJqe
p+J9H1W3zz0DeaSXECf3DzcptDIKpi2jUrKEgtx6DAKE6ghioeLku9jhbHPa
duxz5nfqJR8juLHebUeIRkGcd6OyiGoSccTjr2LeDqQRAwgZMjr3JqHOgl0n
KgAqPYKOauWNoU1Kt/2LOV1983p4S6F7ZFQ0rHN6EQsPZLaRorJLMoVHK+Ek
DDRktxqLsKBBf2+9y1fq0m9Riq4g/UHSX3ZUO/la05xpFhmycMatPewZckin
s2eWRPeMbZUUHnFD8SMQkHIPzaz+QqDlbOIhA4C/4wib+CDZUE3DSeGnt8Jt
X4AlyVxviWAs7in/5jbp6Z8WgNCYNhB76apuKA2aL9vxZAYewll4wvwRe5nX
UFpz8j1AQXjja1JdKhMrYOC3rUMNFb8fSutUOHTLdCfLEbdmYvpl1LYIluGB
iY7ShzZJ/Wyc4dSlXt9EjtpamXVdQOG4yFTPndSPKbovPAK9avdB1C981zxx
HnqJ3sU8ub8q2MgCOHjyAq+3xdZn7BR3oxnfc+K5vT8SXtfcJ/k4sdpPxJK7
2NVJ4MR1WkhswZrIeH6Q7jeDEH/a1IIY4tnFJVMyxbcIJ4kMuQNuDrCzCI2Q
cgH1KhV9L7/v+6T5ZUcqQmyjXds6Z9WlSb9lr43fzZzGYKb2PAfT2BdjepeC
pQutvAvPjsS8sp0HMZNA2fQOAT/I7IYV52mgafbLOFmZUfwh3mCktyLaY4h/
GfGdQGxNexRY9uODWyyf1prR/fAYeRG2Kwu4G78wQtr6aDv328mphSOXFcVo
/AuYa+nFyOMVVvHAqIxc08L6hBy/a6vxArbSs25lwNhum992+2s5dDQekwXP
Onx+MM3V/ysOV3dvxal1vTD1dN8OGGmGJYylF0LuIVcWOx+17JrR5EX2FUUG
vF60zPnxnxtLzXAWR3yADiFg1gTgQpTannvXcrePgfJjmvBt8sE/Xm7ROLbh
pcdPLBZNFHY+Uc/zid01ybl/9p+4NtXGyxXRt3Pf+q7VEbotA176HVDqypC+
aGNN2Q3Cd3uyE3TENEotUWbUoRUYMGMyiW5cxCZCKlHpon2qPQV86xac5jkp
7zVX/HHwg3sUH1iqvdAX0kDSnhVxRN5fPKHUgx5SwgiPbGAO0qgov1S6l6NC
Dr6gazh5HNwAyrFUlV4VDQOG3d5XlR79Do/KwCsAm3RI00C7RqPq3qCbVxeq
z47EJiY05oVLtatvUI1JmZBmmIuYVK1uOFkTCFSYUrCTUnqxgAnH1vqpHVpC
GzpnIktEaZ+eyYLGqWyQT6y6aOQu8dONKIijDVBlN702wya+5/VNw2d96Q9x
2QccBl3TF68W5CmKDCQPkPnu6bxv6WSc5X6gW8gB750Dj4NOk2NpJ4CumnLw
eYz2CEggBm7kd9yksD21bqxwvGnegiqH2U2lYEmv8iYx+OYzeawJICdEnmSX
RPJpw0qpuuPEKoMLsjhlTaRuESq3lLpxj9KwQeSJi7evaB0S8Qwsl5eKQtco
0yVZKwofKtYmPVNUzPJJp/HEiNZ/NgkjV+Uf0YM4pxpx8FwjkID0ereZaWT4
/WeE+kklqvpPypNUs9bnU0Ql7PG2FuE/GrvMGCpaABaRWSDsY/IBdMNW7BZJ
tlW9SOs6+PUK8UyAFxGA9QQbUW6gguZTZV7HWz1fIW7awx0yHMHXyx8HWOQ3
uT6lUCtRZFjrUr6rUHlbUqXAZ1e1Leu7JG4TE8Pm3/rq0c4ya9fnTikXBDKX
CfM38gjsQ0zFzXUAg2oubs+3hU1WPTozJu3Vd3zQWRML8ApvgvUVhtkTYKq5
Cxt5OhIVgvGPHgsYMBPhApUQ82nAufWw6VmR6/zMs+OZe+ZJGdkauC0yavUn
tWN6upxyc0IwRCVLATinVkcD2SLdoTeYWh9+2hz96DFqA1+wPWfccIwSkopD
zxVBnWUc5glykAjxhBG3gwyvwbXEqXUHgtSOn/+u1V90HIwP/LGGlsunXFFI
lM9wCW+LrRvUqUpjT/SrIH5KHN5OT+PULR2aMeL5GBL4kZefZ5VBdAIYBvKP
3f7qajyGYmFYnUNkN+cZ3Mm7aPD1J+OYsMUUB2Im+ElQwkC58XwGGPvLJtMu
2+wV/iJcN0suRGZnEBSFoZfoONWlOUX26kvdOQ43XgF7bhxlpjHbL6pROHHs
EeI7tUVa8bmPld0MQcgIBFfGObnhg909EOBKjVsYb3OMoTjB7DhiCDCPCSDv
f6QkM97ugL3Y2loc7qeDyztxytBZBmCh4OHrx/Pv5C2oZmqA5ds37IP1DJjN
+7g0TFAEKMLfn1KSl7JLyzqEWWKchf9v2m8ZDd1SLaSjui3JDeJvH7hAOh7q
nuYOvlOZ9VSofJEZu8BGUi7fS+UOtbbQzU6lh9tBQPDg24f1eSdsF3l6h72x
DmZW5aFuyJRSpbpiw+EBbMgUU2K/koIfKz/QgE7LrrVQKjDoLsAiuTBGaErc
t0mY0U3GpUFRhdGx9CKEhkvGR37b/RmnSKIHF3TtEBtb4yr/aIw/GLFW9rcE
Mb41sR3wAem4WMq57jntqEH+bAiZhbFrnmTDrM9B+WvBJUsk/Fol6cmRmATe
gic3nTRgCGg+xzSQSXhEXfUXfwFU4kfTOn2X36DUfoq6bX/rVJb9AEGU9B5E
y0LJSf6ulPtaeozEDC3KpW0g35+l974HgGgGqFO3KJK93nC+G29Tz628kzY3
oQkubPeei3DwkObVTX3saQAhPpIYEklNHYEh9Z1fdrf4DNm4aER70pKvmj7F
qcIqMPPx+zUA0tvqHDWTShc2Of6CX92CZKepIGcfHZPoHpPrNXWsZOctT882
kGC4gjpuEQvYwArQ2dayBxrZpTFG5yVL0Gb4ujcX20W1xBAV1yZ+GfqjxMJL
TkqYkgMvJSyMbKYHJBeL+l+Zk2KT+niesd5GO8fUzI2dI9ePSwObz/zGqoM3
/mvyoKfYJtqc3iQr0I+Kw+fJcRys/uGFNjUIP4OlA9ySy9SagL+/4+X/G3R3
DpTjLZTAaEAqT6n/6Xqtt6UFj6NE5OJNi++EtWtrKDhsRYpd/1D2oBHhG0pM
SP4zjJc4O8ew5WW2NvdFq/NpdFbS7gpAGANXSnQ4c80UioDWuRyIyrhHcV8M
O+0+9e9U+EKWQmzonjeU4e8ZPcTfHV/fWN9Zkl4soMKpqKHGW9wrHXn51N6q
MNIqW+Y9B8hn8+tE/BbNinFxiGK+ydOdiuY4bxhC2wzvRqCO4ApNG4Laal8i
sIXCKubGT+6xKi+qdsbkdHU9Uj761WyOBFdKXk3CEhOy3TsVNx0BxQBEvcPV
jJDv0XkTc+o3d8qlWJBmRn0ISvAnthbZ7XzhIe5qbbjexeOHKZOnnENIG6GR
w8IuZxpwDg3ARqnUTHIpRaqO+X1wM2cmDSWSjQEu+9sxcXpZIRNRUwuSG0FW
I4BcMP4vVkzfne+EpxHtdGREHduRTg3vrCWrWScIdmwbWx21gPhveIfy0jrt
itlMYszEI41o+iIOrPJObVZqpksfDzFg+eskXSEdS5SR7NIDEjFgnBTF2EJz
2ff+j+iG1sf8n9ijAc39nce8ba7htxt5ObAJ2AzKesw7r0dUMfaCfL/YRriT
1ycXbJWjYGitSiJR5t3MI8rxCNAZv4P8RQ85uCr53yjwDbdII1ieW3NTsNEZ
VyjDm2AK2DdyyhWo35WSm8F6CjNUbjATE6xNq7oIE5XP8Zlax9fDd1KxamRZ
BU1tNbS55KzUYuXG5M1XO6SC/lwOVMyEDPa28iyLdBKX+wVmTTzvZb4H+tAZ
w2varfdSMhvOetsqG/LgzRbaWz7gfa4T50G1l1x6N+WBJA7L9QCtYT+L9tVe
NfOngXwYF2NcMHErzTF58MA3pFbYTS1vYUB9vVSTqpHHjoJ5jfdhuGFDq7zU
ixbrNLFwizZqKFHHwvXPcFSKLP/S5pXom5XJWNniw/7Enu1q/+BuabfYtHsn
79c1uKmjX0HE+AuT3el0i2kz/ewWcKE/G4goVHY6b8kcmJ1Flyuy3KfK30ST
I5qCUSTwtUYBa5ny+Vnz7HJKrkqs+ny01DPRZ+hkxSyby02gXDb9wlbBvI60
3j4JSqftAs/ATjsR3+80FmHzfrm3VDva04fT0ebjU9Wzzge4yr+pYWU1jXHT
025AY3SN6M22vsowheVD7bnhgsuuNVXnwStf0cXOMIErXjjHlJCpWZMXNC5B
FABO8IdXOsM2CAIXSnIiGOV7Y9QY45EOdFjDFtBV6PMD1WG/5UTL1G9Hd9LV
85cKbtKw89AL48fQB1AmKBMMfeIpPjMa9iPyxS+UCPpJmYTh/QPsTi5O1fez
E5EzVcUbup1+YASUIt5VqxX5ITlGQPActpMo78Xl/l1k8owrc0l8CDVtyRck
jqmnpvyO19YDEdHATvEAyos7xw2pW/HCaAWIbhVualcy8nJc6yIYXrYVN+4Y
/PZrXBpxd+O5L35/YKWjnd7tcu7uE4XmYTc4XVOCXnfp/KkEo7CWLsJy8H98
mtJPa01/Zw0RS748qmll3j2201LqXDQTchd1CxTGMmdHyFUtP7L7/BChUNn8
r6TZ6G87wXGun1j152IkAQHeVL6TQwoQ/J8fViVHkgFyT/igghidobjfmIff
25uEqYsMteNDRnvlIG35zxqRXW4fygH6PAbibYxdCeKVz4MpbMMdOdIbK7p4
WK+2t5KkDGvjQjoCTrKdb5PRJjoawAh6gpco8jDMnoftd54otw+TVXXuESaO
TNG9BSrRHiGby9Gt4D9YSRguQG8erm2TaWV9Lc67VC3QcL4E+z3+y/OYDqlI
FxQJ88cnD5fj/y68Nnl895vuzsj4t2lv0XvP+UAW+sr0Dk43gMxdGeQ03WHT
HGlb3w5RMj8ClcCPVRa2Ja5HvTPwhyy8HwuK8jbQEvcPnHADvvf6SSLf3/br
b+fWxKflENYHntc8FQuppNqivxdv3v8qRKW81dK2kJFVyv2pyEH6WvWIfswV
LEvHEEmdrQg9c85SSEM9KQyJlJ3ePjzoKtQo+Knwl7EGbUMjHP2TzrQiXkuc
gpBNwRxm9yp7CSKoN/Sq6A6V12vSib5ejNmVtsTu7M5M6UK0PAPnl4GkymRf
do/elWGKJLB6jZXhiPnh6bFJclR4kCrYSsPGp2C0Aw7VogTpVf+oaJfBXcvX
zuk2TgXbZfl8Z22vTLoXcm1suQ4aXoke06xDgX9Bj7RgXDpV9zA/EokZ+qPn
jNL9KqgVZwvE7c8UCP6McmTQ7FJGsFFa7pIIbY1dMQtk9wGOQjh3UbQ7jXMH
zec0TvUmjgpZTSdUp7ZPQgy0fGPqN3xfSqgVColUQGfLXEMBApjJ44Xlxb0p
xcInlKQv5BLT6NOvJCngnCtZoIz9SPXrd3Ku7PsXkwp61+yzhbsgFgxtWre4
XWz6eciYyy5ChYEn/BPT/1LyfPB+tfeoECAFGZdEUQRpDfgAX8lZYU3A0Beg
IsWsuMCg0rxpxLKC3Cx4NRNxOrwLuY+aSVxSBYcq4kJk67Oc/Lyjtts6+MjH
79qPOdCAbP9l0c9HnQLYQWCF+EVq1VSZ8NZijQbF+4TQWFXG7BnBNDenWroY
RCpf3GxbxZMnK/yMq1z8ZpalJFkVzV5vtTzMAx/5KGqZ9FH9L8qfdb8KwtVZ
ljafjZIxDrS3uKowavoDBd0tkqyIyUq4efFerObXl4NtfYBej+v/fit8497+
8LfBK+31XU60JyjI+6rWjt1qaD9JTbVO7l3UW4ZKTMgCI3/TPsa8+3so+ezR
4/mnHF8JCfbS2fd5CHdSafB46Hn2AjmODh7E2CfKJhzO9e7uiRZbMHOTv0G6
M97VQv1zIP9uiHFd1RaSGzZO1DTmvlYi+j3JZNg4C1JSxswi+5CDFGSbNXCK
+yEt5/jWdKE1PpSQUVH85FxNWHo5L7yJEHx2l9Du/FjewzIJjdy7ooi/akQZ
ufM8FADLgdCTjc0G2ewXOIvalTPvwdG5rUiHZk1/ae+FkS0Lg+olobktpEbU
a5Jd3NxNtAUGj3XokpbYNgKj/BbXz+fKdGxfx7VsXpkohX9ddJG8btA2WsTg
B9HLPeImUX6IdN3qu4DbDnHn1QpGbRq3wKSZ4/sQSBCCFdUyCG2c2/gySKdg
NzgQNAEeO3ACJUNC/gwJSM6MFBJnqKT/eUV0RIb/TFxU0AUFBkJULIiXlGB1
UAVjr3yw1xO6koOOWUbxdV3rl+m+uUYOxNBAUR976lbWnUKAAEDOD82TI84q
kb8acoSEuOomme+x1qEBY1h3qjfM7SV6WkCAYGZLbvawXObrsOzdZPoyISbg
j/xsLbPPInT17flWrHPouK/TnyLhokFy1Pxx1RJUrRxWCm0YqYbzZoZ3r9aj
5dnsf8oT01ORD9bjcoF1R2cAgaN/5tQWbhNuNUhmZSB8i2bCK1WogorJEQ4H
d9MQSq6i6aRrzV4PC1PLqyh5kTRi2ozoChUwDwLwFh40x7QdxmHByJAq7kyJ
pDyvE+8dWqbPi2P/CbyiI49UetcVSal7PF+mPz219FyinI2mEU8SG/uR58Dc
JrC9A2sVT68oV+Sra4gm27VgJ10P78N0Vr69dU+IO5214ESth2VRpwrilspj
yDilWSpCVvSjpKlZ9/Pkv2S/4VcQx5Xv+iI1BuQN2H6XhFxOIChA7vgD4Mn0
fLxTpfSIx7trU2SuOdiexcbjnI6O4cuMP45Gpi8B3Mc+i7vObnniDAcU/nO2
nzEYNyQQ40gH1MfSe8riCtK0ypbJlynkC6waN02N/+omREdy6FpP3747OS7Y
xtmGBpzTZ3OJ/6Jyb6uNxHpwH7gI8+URvDuNOxyWZ4gOEK+nDT6Enmi4B1JI
M2TFRufvVsQ3HX5ampy4PtZ4C/CwrP+wbFuVf6MJRcWqgXTuJG8Fy4BLF+6N
5kiq2/Ty8vIEX2QhCw6ylkpK77E/DQ5rVGFHX7VfugxIIgQrRaXvtMBbc/GU
Y/zrx4t83HYmGwPJAxqAdDE4lyBkWns9PQdD4fAlmgOtGMWHmsfE3jwFjw1N
x7KZYagoh9MHovT5i43VIVsduYM+Y4MBUZxXMEdwm2gMfhcwuLlig6yIxOCK
SxY19J9BCmDYM5yKmUfstpcDuaPqElUavFgtcBv9WyX2dwLyrM10dBBtL3NT
OImtDTSZkAmbVUBZvQPP9LLrF8zW54sDihXskOPvPDDe9dvBQunCIIZJVzvp
OtbS7XR2xyBytvpRDr4eOG5V6tMalygcEdRgfWMdxJe/yoPioXfo/Ob3HzVG
USmCQiJEjUQsx9iwvJZZi3exeZq7GvGRaIGko2oif/IEoL+fuwq+fk7cLYtn
G7pr9yq3Mz+wG89jxeIbuMZ+D4wS9wU4VTuD+7TAxhWWfyHrWRyAXMiiWPVs
4YaOUEiGHbyJY7iVGTKHX+QZ5X859i39509nLk6YpQWlvDReAsQ/dREFH/ry
rv/z2lZoub7Qb/AP0qvB+cJ1Yp4OFsncZ96Ls+FmFJ19+Uk1pqIveRvaQSQx
qdyvpAgm9ZEMQgakbfK4L7DF665PTybchzUKjcPoWvttbuaHig15PFTzhjla
7kxb44IuTD/jt+FrvIhO0NtgddQqZ8u9IvF62ZuwRAmfuxaZP6gUSkn30sXl
0snECeaZ/Y2g3YiMCB68MTdSGYkA3v9ix5wAB/xj3kKwSgrPwTNbdcj/DvdJ
ta3B+pPvvorJFoLvhOVTRGg6e5sS2T8F3a6hz4RJlbwKNiCOuDEx4jY/tMuT
MT6F8ueSf4gnH5p7IntJo8ZG0kfdMEodbOv6sG5yswC1coqCAh4nzDhHgHos
UJlZP/eRu0QOYfX8aRyamkVKqZEYD9QcMigJbyV7nDd/WXmZ3Nr62FMpcabl
utDZfFsXyDTJMMqp9NS9t8Prpex/X5gFLUQInMsT1uBZQycV7+r8LjBVpOwi
zmj4pw6yX89Vc3NMB6JoPylYNVKHtnebhV/DjvV9Uxzka12G56fDDEyDmB6N
WR0LBmNjy6+ksyTO4UZhA+SaMN9583QUu0BbaT7tjXolG2Jb6bH09gSuskep
/+8avDJ13x8iCV1QcNBijo69cYRu2g0ckKUeJSi4451umGjDH47G/RtLyNzv
N9PNo31y7Vx8iMMY1iiwxe6lZsTQW4+XJBhSL/DFdKHv2pERLUWu4eCFbyQ9
xYEyXU8lIjqKG4LKnzKIdz6XFyEYYMIx6p9/ZE/UOm53e/KH1emU5EQilqzi
5UEcXR+gCZ+s5OuZvxtoGJtl4XJ+lJ/g5Ozhvt+J3f2cb84zwKDVQqq7uk+2
z4KNWZzE8OFBTWMK0SSyHESRqB/Ks8hi65TP5fjOtgrJQAjVzIZF85U0qMJK
sSflxXtlhaooqwtLcEe3CIwmk9PrPLMyAopcsbEcFYIcnkqsYdlSSfbco4F7
V1vyn3fEE7TasSslQEX2XeY7wDdDuV19B8eKUGBbFNelgtKh0YBDatIgJwnK
8OPNddiC52hFEzRVkqmc8SLZGumK9525wsVLX/TcLPbcX1vBPLQCe9MaLZx1
pftoWoG7gieg7Yl/LMCg9q4u5blCuRQaCzGZljRprIZRXQoho8BcSWv4w/43
GkHG5XpuDGa35ScR5cRo+TXQm6NyUQ6AVNd7GbGBd4mnDcj+AjUu4IupS66l
R/ZabopsZbgJWtcB00k6EEdP5maqqoG2YXi81QTdDAeFUmiu3pYz7xqEXtek
rqfaMxAaU4x1yMfj8uVknkpDAotYY7Haehy8RzuGBqnS83wvu4rDGUh4zb8C
PKJMMeOnZEPEcdkCVVTKF0glHpd+UPEITkLw/AqkhWxAEHLKrp/nHGsx89MH
N5D2myay/grOi/xFeYfqmoiJ4RliArxURrwE+8YwdCSxbZBGdYZNTbtmUVr1
psWGtkmR8nqrs9o1+cof2zLSVPvy2H6VJlpey0K5bfIZ/jGrprl4NtBJe5xl
kspiNmh8HCNZxmHML9cA73RI08m6Ff9p56wr2BKI9buh0FiC5DLV+cnboYRk
xBLFcV0ufzNXYhCmT8q7HDIMVu24m+x+9o+7n2lTsszVteDHlNKVmk0qYEFl
oRqszdQvWFBGpNeIaHpEBrec4jebAweFfDMzjLyENNN+O12ow87cUJzNjrzp
v+v8n/iy6y4cFoEoOfJMYt6pXc93cUBHyaWOtd+LEAfcJkD6ksI8Bg3S2WnW
gMa/Q1kvPGrQGnszv5K4FuyMQUIbuzEVySJQyrPRuTC0TUbs1FkxurRs9Obb
b8vzzsDga+Q1t/b02qEgYcmw/PtPx4rChddWRWe0XRpmUD7eVcFw6GJ0Burf
ElA8aJyM1ovKzqLq8Khm+nITZz1UNrW5sseDyOY0Cn7o1YGvVv+1+i2TLav1
HaZnCLOkHn/CvDbSxdgChKm347fn2BGEAnVJp8bgNgQ2kTwYdLpqPA8Upgh5
zr/Dx+TSjtyuLKPRekNu776KEf8HkuUd0Vn0Gfw6dgInkSeZV+eNDhVelP3K
96GbqAuAfCWdKDDR+qI6ddh6T3wqrCEBNvNfHGSSkJGzrGXdy/qbZUV0DAhp
f99EHwOeDTP6dp5PP9kbVIFd8MXH4JiGD71xU3+4qhTgiVQGp9TlOMxJRkCq
1XdENgcTwzCrN9TSjGHKQj+e2C+N3EMiOEhrLfQ9yI+sJoSvmQ1OZA206S3b
VHnZ6Z+3nblMkes4tHB/MszIMOFMtcKT1QrSi6c9cER8iZeICkl9tLzWwLy0
0+2uHcS4+zWSnB7+IvYq3XAgOM6Rjpwgjrrp5hCb39pn+R4siB3ZR9W4+GNk
Fdk4YzrdqXrlcXcJM9iGmz6GiF5LtEk5KtQLd6/Z1WXfKIW+qTJtZJF7zv9L
1hmUdmBbtBS7NNt8/KW9LBBBZDsrY+F4rsRjye5c2ImCWNAzzZ0fo0p8sEeO
74saqVut86RBIq0raj+RLh/nsmLTcHYQsorBgMEW/Gjz8asyp68UPV9IFtEc
l/BwATzLtFWtdcgMDf5kASjhX6rSavhKlE4fbihC+pTol8Q60exigzXUp0y7
Y/6mdaY+w7IxGXPj1WQo1Rmo6BnnhKZ1SwzN9auZFZ1vcEn31KN+3FifC3xv
l7pyyjXmpLjIjYi4GU0l9qinIzdG0ciM7uDTXgg2CUQuI9FwQQXG6c1Yncro
HOLMSvtqZ9xHnr2RbJuuR1reOSCKHlk5qsq2qREeN53oclukW+FVuOsfLNdX
AbAhMrse+++D+K/YhOQtYxIFlts9cp6ZVSe8+MH9/aZRLQvIm0dGwKejkpLL
Z4QdRpsGUwQuRbb4s1Syf/USDQCvSoN35KElJSzCiNhMYnwb/pciV3cNWm9I
wBJpg3DkNOEztMvoe17zfPIvzl3/u93/s+IuXeErDR+BcE4zd0crHfARQdNn
tQYIm60MZytIZkiCYstV/wVsoAq4hhltrrHjOZwoxL8Yirr99Y4xHLblSipI
tp+1EKXfAkEOddizT0KETo7iXLpmpXuR0EGmKR5Nvee6Ujdyf4FIBDDkdzAQ
U4eeUvGsowZybgoTp7RRYv/+YPQoWMoQbt/lQrRAzonisFL5kRHOJHgJJr2H
DwKA72XykdmjtDd4uvkXn/qMAyVH/9nlcXgGPZD5I3iAFfBkc/YeglnpMOdO
VNGAzI6tY85YTCP8rHXTXP0DCQyQWI4a0r3l5KvTdfevhxheENxo8qVxzsY2
k3YhaNFrpvtvOh+NeZ5xcIjnO0Y0O4T5mLbPO6WOYU0X0REo3qqwc3U66qF9
+0SFjAskjl9mhNnyJJEaFymkhT5AKuJcfCPHx/R7HIjKbLIDxtQDFUPqsTgB
VXdWe13TVNiP/E16TXdl2gEpuj2IOgxO2sc64tXN+Icbl3SKEI6k56gvXkK2
2TjrKAlk+aTijxIQ+Ymra82gghoCuwieX8XLcBzA8Ammchu5tOff/u1ziv6n
qvatYzFlp/GGLNhAxPAwSUV2c19Q8yN+AbFkuEz2wP9Uiube8Mb1fLMQw5yv
5KDJJLH/48fyrC17+YZwLWdx/WCLWFPVFMI204VZYY9onz7yR9IJcnRHG+SM
lKvU6u8asFQB+wxS53839rfVGsGFfAKkgQh++gVn4dd/ilzVtYdSZ0DxBwJO
ptTqowYMrZ11xIRg/HYbKx1mlNBI0Plj/peJo47gLdUCSaG4ILvvRLOh8Qwf
ikzAM21OEWg1sX/TMCftnXErgzMxejdDtmQ+wbXVp1SgyI2MHjagrAT1pPij
XBma0a/maoHcXmq6Th9Fl+c26atmDzLrGqqHDtNO7G0+DF3yc2UcMc7O20UV
znankOvlONbOqjijA5WNYpfzaAwkPZOq1Pd1/blO8ZKnMqIWYoVIMoKKFw8Z
WalRImZFT5Y4ewBO4Fs21yrZOV96oXGdb9IonT8p0OqBesrIUY0aMTin4s3D
8iXXesfOs2YsdAIXqpz/x4JCPiiRgfJOxvPchrJxEtK4jdHAvWYumLPadBzA
QsQXrceUBl+8pVaV4qb2Mm70Afunudi5VYd5/6KuqnEU2evGIMRwg6kKaMro
mBqujDhXpYpDsLfWB7q0+eWaAInHPj9vycMrxN8PabD1NoqqwsdLDP5tSuv+
LHEYy84qhfyK/q/VP3qnQTEe1BPJKP2xuoBJT02QE+pK+6jN2v0/J1a2XKi2
X4Yuhiqzwfiij4pzh1UYE3D/6jIBM5m+2auvmk2f/Jv+SstBPfRrShio4gKZ
Foi+q71i75pKHJ4cFPgVQkETyKjNxV3wHPjsK2WrjwWmWMmcf4lUiq+XRv9f
wuekyVnUc6T9C6LFOVFczDhGvErUKmQqiraBQC0B1l0fAamdKtfiuOcRP254
0QLeQWx4445sWrT7fe805hlDOhXj7TTYsUBKTe8ORLy3lWtUfkjQSEwwM2ok
dZVseoq1h0EN8g9j4CD9wgDGGl84AqHXIsnjOQWoNmZ69uIP+Kh1U8Mbk3o/
WJs0RuHh1WhiVw/IrtWon6RwR+h1mWiQYKcIIZDhe+iWW6tbJzDBP1S6M6nb
snDc5RDGmNIYFo79E1Pz2VVLmz5CPlJ3gCYMu4IudgruRjYDeH/DaqmHPUn0
XSioSIOuuWLKYagbi+rTKcZNT4BTaD99ID85eI7Umcqyidn/3WKKDDFXLcwB
5THrXMMsc2PTobadvlAQvky0zcrr3AMCj2J1jouQCqvETmy7qpEDpwJC/sjo
kXa/R9bD+z2JMsHgYHG2pZW+5k9YJwf71xW8VO45b3taIi9MXek4KXBodZpF
nh9AHn9XCLYeFmpuTfdRsfCKeRaxE63U06GaF0XewI5Q/UENsg2NNo3XelRD
D3aDHZv69QutAM3XDObRZn6Nq1f5VEe798J76TekK+a9ymzvXxul435pPucj
rGlSdIrht/1XF6Bh/nOxSYHWuggtYl4gH34upK1GAHBirROQH/OKq4A+qcF4
IaSgLksrvfrABxGWD1aS3uUVzpWXciJagVj/2ZObHVSZA2yPdJWBqAS+SGKc
YaoIXQnCqM1a1wEx6r38LKBHnxIkOK8+Hh9EvWB/2Fira4bXP9G1vp8qwlDB
58sYShMeGq5sUboCRlCJZNzdsIeJlpgHUST2/pskHEQ6zq3BlhUXw6sch7ph
LesJk5uPqoj0XKcDE44uLyHvNZ91ZLk5Y+XkkjNsi9ULkUo3a7WJbsuzw4wZ
H9o35xM+GeLzrDTq47IpW9XL06XB67mC0/HMqKKpfy/9KXyl0wfH+Wi0EVc1
eE1xPALmriH0v6/yZDX2SihfudktXicnQjJIDYNPnmxxNzNiSGJ2QbYdqpgK
BilFRNK9kHN2XucG7E389abbJVcYY99jQT1WdLMco6nd8IhakRIW/bSWRMLI
jn9C6kFNPMOpgOmyraq8tzMRM0ett9g4619DmhF25XZnkQeAKjEcSuVkXOH8
HOa1eHY3YSLleXtIEfAzDo1MKm/taICwuR9jCrUyr4kbwnjQVoR1bVfxRMfQ
5bbWBc9JlKopprsMDloX98YFkiG2M7IhJtcLqg+NUUZae2cwoB31KqMvNLCB
BfiLo9tjwuOyAvVAv8fE8pKXWvUi3wEli2kuFapuvF79KEGoRLw9d4fJB2x6
hlvmuMA/Q0r5nTZKmUa7Xig0ABBcWgEZeYfyocIjeXiCR8fPR+XZW0vWdA6s
I5emHNa7dzsdvexNsX8jlu+10U4o0QX8kXpCrQbT5bOL1V8QkfnBSNkblmFp
gnpfKSM+CZmd9iJPphRplZtl/2qzqzU6qyZ1Y2vqp4f3wpl88pBiZdW2obvN
7TP5oAqXDsN3/5mR4HLIbDvtyfHlcb9Kczd0qRlCGI352b1sUIhSyQa0xnn1
RB14dyyvWsk4lOqpSp6MVtxWOVKJSaaMffwkIrivh+qta7Ntv/XXEXuP4SMY
r2mGUqGdtmjhOPVTbLN8T3QcAhTTo0O+I/r8fIDlrxhZmh40idvKIti1l0JM
bzzrq0LiwsvYJvDjke7N/MkUodycBB1McW/ONO8dhCPqtFdfH25V7NLgaZeG
RY1a86xi1dij42PSuBYsHKdV8WJNgH/djxt256I6Ganp4R/rgYjO8eFElb7d
/qZ4CpAq8ieqrkXhMY4H4/THsmmsLJ0F1ScDxxTcab3T56c+FXP/9Pp+efLT
hm+oe9vJlxhDxIqiudabR0eEemW1KZAtEB+Hcvue9HrR4THQ2CVIvC+5h5tI
OUQhYP9cady6jbzkNL96wPpubqoorRW4XbRi+RoPNONekfB9KtXYLRG4jvs2
dExmr1g8A6RY0JCYAmDr1IccDbqmlk1lZcFk/EtKcmFM8ypaKVBMEqG6gTVl
mDy002bD2PZ9ciK9B+C3faPcou30aN6GbJePLIbtkhYIyv0IHCEl3QTYMN36
5zfaFm4PFwho1kb6PBUJCdB9fgixEJXO2eokOl5L5th4/Bxe0qrmkP295QEU
xA86v4ofWg8cHbpYYn/hzGOudlLgxnB6RlwGUwHLB3yasullgG4PmehHMp+S
3oGrT1Q5rmms8ytAmN0nfqN0viD+H+X98BO74KA4ROAhwOX+LgrE21OjPkA2
w6dfXJyYYdUvvi3soiQzQ6UFIJA8yaU53obiPpzUFJg+SliTvSQEvqsV5N9C
fQEtPjW92bh4y+Od5i6cSBVtAbasLHxGMchygcEEEsFU0iFf1afXCDfu5x7i
ekl52C7pcdXbeWauY8TeRxP1Q+YBx5NSlAFtK/e8XjA9t1mmn/8mTdGZnBas
EtiwvczVPt9TMwqADsIUgOES29WdTvUQ5kpj0LLhVcmuNqZEaQHfpF2Vo2lx
yNQLboszy+kz8bZaV5Nu8AdtaBzkPZijmw3N8fFpIHn55a0M6KjBF+sxfv05
V6RamazSTGpI8Tet5ZVJJ9DYGkc/AWynoOin3oMdSDlKPvEmnhx583uCq1IW
hlkImC7i62aV1ek1lvla2uvdcPw6xYY6VbWl71Bn1xgomC9L+wBZVtuKdnI5
iOcEUQEVgb10uDrXC8quLiudhMO+AKeJE1EDQI9aXwkmYIqAZmnopbYX90kq
hU/epKEkDwG94+z03wm5BmbtlXiSgSGaC4iElK2vw2S26an8l54dUQbRmUSP
oPdNaPMtq8RFKNKwqQ95FI8XE6rZYTEryqDB8zenLjlnYnE7DfHlJdzzay3n
GrH/I6QHxAVMgdnHqB4cNtg2Qp6nVFimH+VKWb0DQlMEWVf5TIv2JHTo9bDy
ac54TlGZEr/jKQMG4Fv+PfrlCO4Sniuzt/3wn9eyxSYT7Iil/0+41f8aX10H
hCH2UQ/qvOGa7TCzQrdyh1A9sng3QlMjFYANrTaMFSUKi7aJ/yjNgkP1jKl7
0VliHTihV9WIY/RPUTgSjU7octiR2cxTowAJojFnToW6K/3ToKI7tZe5QjX1
stOBRG4IzIqwgcLb27pD1VFHUcRVDh2I8FaSwipmOgo/cHi9wBPX4nZqIYya
QAXwubJszbZYaojgu8qtjCjHubztNN7xtFyeXQjAraB15blHQuUvkpxkwEz7
PDSr6RC6Yu6+STiO9GSG0j4Vt2C698Ey/DjkcULurOY/ATeJqRn9RhKM8JHq
ZidxtpmMJDRlWXp6WcmeYNrb5RWhewLajO8Y0q/ysqL55BTZOxuCQtlh3VSH
APiqJQW3dJEVza2r0LA66/IkP5ucnAbyBw12lrUU2LRr+nCcj6L1T88wuQ30
hH7rPUitvKcjMAeXZpMvb0Cv8F3oyIpN+XgDUW3Vr1zQ/awZW00VBqNdjBqE
zxH7no0MYlCDcF6b/UR7E68+o5QQrzXzYzkE2cm8Z0DEeBcSu3fVUP5mUkAo
32B5aovKBL0ZKHxap8XgKQN1e9jhAj8ulToBS/vrobRzJoT1AQ7mi7iccOpU
+lpaGF7p/q3VD3j62/ou7NjNMcnaDqe+zveAlXoPFBxPM/rFQV8OIAEkwpCm
1mtEzbih+OhaMtA6RdfJFjVaInvSMUVSMOXDvbUagMnLL7sB56F6eXDCZ8rI
phzy9gn2rB8Wd9Wu1ywqdKTNQMLvzqeYyUTyG3CNOlWcG8CqLsRSNKqA9y8I
WVa5o1oaBFUsV4NkAy0HLycUkOstZQz4643WtY7jYZ8iU6AGFzKgJAQdl3XJ
qi44YIigaeCKBREGv8b/7jmAPmz3SrysJFdMduEEVuAcR+UWFTUnERGSu28K
uZ5QgjFVKlv6B4YZFgcIBIsb+IR6hwvvStFqr9Bs4dtVX3zy4mDrW0dh/r6/
S7Y4P9ssPqMQnXK18il7JZ3KmwAakpRBiJ2oZib9/ls5sh+IKCQ1bClA+b5L
pxA1JCuXNBAFWAiW5C8AV2RA8OrvqQXh9nW/2oborPYvKF4dOrbpJD2zi+CF
YaO0JBnKS3ZF45kgu2JFLSygTbw5hn7NQSVxY2yH0GY0TaoobhWfiIdlyynW
ui72cFYQa73XSlwB8zm11mOmvuvieFfZGJYQVx2CGcFFjI7zGMuom2BX8wed
86dPT5kDaXwgdXGVLsW9w0kTkZIc/clYg6Guojd72cOPs6ugc2aNlIlGlgzA
xveb5wUzZY7r3+I6Bd3M40dV/G5aHyOMuhBpoytkBaeDC/KfLUgC55Es5Zcx
v9QVbwJxS6w4p8iQSGFyulo0dooqIcf2KnJ4LzmB24aqiipg9ZVuiU6ZuPoN
ioa3AoLp+ZWvygys+UmQcjqceY2VMgO+i1aHmV44YBxlqvQzW1+PQ9yaK9pA
Q797CqiFTrQH1QCJAqQEjMW6FE6ZtRd0cKtFNTT0XbZ8TUuPntFrw8vquCYZ
lBuFU+T+f1RyeYxtJbDZbib3DLyU+Vgg4k/hw0gMeyC1s3nvvB2QwZZQxE4J
RG56M4hRqs5tqwlldqgdqnTD240KXQkvI0cT1jA4p4D+Lpc8GgwOi2b+Pnzt
yVeBpqyUcswg0MyNIhv0C9tit3k36JaereAuEFVE4coMFI9v3J8QKUwK6kVO
QIydLJLyHCheOHW+Fja6aEKuOaMmgrH23Y67V+0/O4Fv+tTo4h/YB6c3hrzQ
ChP+uCgSntSZ6Vijq0RYRfQd0CFFac2LevARKo3S9INKk4/KCIv+YCYOTN+a
gUg2btJ4EAlVJ2bbG5zUlyAzx4igvVTY6G0iQrZoAyhX01CyM84Q0UFjbZX+
xGV7aVS6DzLu5yFxlrGFlTv3b5XPHR3kL0GicwR8jXIw7aSosBCR99xk/Fay
PqN3LVZE1/Adp9RumVsnx3OMr+XHEXuZ4jJQeT8JO47tBkFJ2ajHsz+mTkqv
fTFM2APUGTmKpft/7wSgqqqbvJqIa+bnG5GuFuTIPYe1jBDS2J/6APnxDQbw
RGh7BGs6lhicTl5ysTePvgHN5qzgDRgv4XkGbrmNxw9z8qOpHsVtGmlJlhiK
M08UGuc4wP0yrfpL7jQgERtQdZgg6MtOEUN0yUvq/pFn0xSOteYOG9Sn1SqA
b9ElWlI0UQYn+LsEcJW64hw8J31073Lxg1TkM3V3qaqtz3qx6HVaUo92yie3
8m2UzaLokgKFJHCFGvHGgkjYLgx4YqqYzYzzNAPPZjNx4g4z89gcMM+iVNqo
wLm8FiWQAwXJFo2+IsJCprNhkDq8loItTtuXNcH5d9gZ2QuYs1rnu9k1do5q
Z5CWldNWLjfLT5Er5S2guZcab4J5Dw6JvNYo/gav1400vBDyk8+H9B86L11r
ddQM4D47XHDuU6it9HsP0AB13at84e03PDAWglvbPos42skd59y6OieIuDlH
dK9vnt/ndeZPgc5gTU7joJaTqjHKwfI8pBSZolS1zXvJ7wX0KpELOo8NYLMJ
jR59SC6N+ayoGT/ySx1VhZZy0QZot9+cF1zhCyvymL42g/BhUMGmY9P1HGvM
C+LDFzBBEDjDUqN1ZuvKB12wE1A36C7wdXuUFWBblzg812nr9y65+Ej56SPY
9FJR9RhkKkjERADGIV1ifn7CmS4FVpWmvSLjiIZyf17d5XxRsf8r4JYXovg1
2nETTyaO2z0TPQUxozrNOWbd4ll61WFI7kbe3xJdaT424ym07fTCKeHXuwrp
HxXCpVpk6vf7+ksoTGVLW4VYuDC3b0dKhQpLFaApO8iMOTokIQclN80+LodT
JbOZ8Pr/nKIIX2X9LXvmk75D48EKATF2AnK/F7Mv3gM5dnwV1pEN/dzMGday
b6gkiSc2RqaCi1DaJefsRNS7kTPkzJvedY+LQQHQOZQox6E2t/XiXivhJ+SV
wY6WO9NZX8SdbqxOxHpfyp1zhIGzpIdFArwM8DBOPeOsEgqeyjXmMa9oumvt
4F/Wq/SEEeaLZ3qxsrOEa6OoF14sZlDAJQcyWd/ZL+iW1qdz4CMVWB1OZkUx
FEUjk29wkcvI+5F9Rgu3RjTKqc11Hz86OCz+YKFLdN5Xfk8jIq5ErGAh75MF
KxWufJ6pKizmTS9pH3GIj74zKWVD2bF/lz1e1/VnLtM+eqfFR8bjEkmM9Itn
OV7tN3Ts4HcJbt5EXG5u5AMUZ/r+htyKaOPJOLIwuq8jVV62qZ0XDe7gSpwL
taG3SRPIrtnY+CxQTJNLutzu/fvWL8pPhH2FylaTKU1e5woK9/Ry0YAIA0Fu
mYiRiXOjAyv6ImEsyEdA35W8hI1UBdCrermGAvvmQVlftLsr5yo5XoYt7QRQ
eVNKD3ogpawSXcBtPSR0LdO6WC4m5qqOCbJxJzXQIQLl0WOaW9b6c+P8kWoX
cRRFyTWEj8Pt2oyRmZ/oWKyjQMZQdW9++PYT2b6f8P9xnm3GC2ZFovJP2bLZ
q+efzNSnIix1EyIobaH3nEEgbG+CjjtOaoo/clNjY5FKHUEaxAUvG+F2APtB
9h/ZqGtb1uUnbpnNOgx302pNPt+NTwd22b8TvpiBxvopMzp58XIdTZeVvlI7
9ld0qpKUvjNGjlfU5IG+NM/X5jFeFDVmzdjveiuHKDff20a8Y747Wbk9ypRw
3ijlWjyYvuKb0yYD1oKqhR5NrtG4W1LDZYqOOX+NN028hgtDr8tpePtfl46P
xyfWemf2Omgk5ywMLX9yJHy6PJ8j4cO1z7yw1hiLJ4CCaS6kKqs8CsMNRJIn
WgocUa5HXexRs6ESU86UG2Ew8iIxXQIAgvWrtKunaPc8iFRy0YkKT5K8IuPk
9K5+ov/tgAJ83bVrKT1Bew3DtyToDbF1Lv+hw1I8A4/2hxb8hTS6GK9+Y1yz
FcJS9pr9vIev7gcH8Evkts8kXAhZL3Lzb0xWhq+YBRxzH0Nt63lkcE+intzK
fY6ljOe2V+qhFaLJTKPcsmYBN/Pc9P94YQMRz3o1pQvi6/Hn6eVnTPoDlC9M
mZexOwrI/fbBGB/xfTAibbrcmLXMWTrzEkHn4X4Gw92O2ttyc0KDwOcVeO1W
gUNWRMNv1/lynbvQ4D8+SVrmj2VlGIJZs7U0ymb68+jlZd+1Y1rC16rtpOQh
nRb+l2qJYGgmnPsELtd4OIP2a+giNU6WeEXIIWB8tvD9iLdCKmqRHyETtv5h
Sgk+LBehgnMUl31JmlBYhnOkME1/9xwH5ROTIc1bHYNUBDwUFInjcvXX4KMN
+mF1U+tpZ+jWfDO+cA1+jf0JHy7B1I1Qro9FpkJv/7OSBFyE51tsmVqluYP+
lF1LU84KJruH3lgEfD3FDG7bkb6XzysNTAcvi3+iVMRCky7YG40vr04rn472
zwx4C3uos6VQ2gGaMdWyXP4GLEjEuXuh5d2kncuHRS91JnIyqBknPRKtMIpL
LDQggC4EWJuETPeb2W0cGOIOVg2nj52O2dZM0c9Dxqhxmvi0ahuZRyx5pbz9
Xnu6pC4+67LrIe/1zlNx6WonkZ1VA2WvEcdWOTmMYiDGbdccAO/zZneHFNd9
cHKPSyAxlopnUZ8MmnMypMcPb1DxlyxneYB9ieRnUOFRZf5HEVcesOCI/1JX
w4xZiwPWR7oxTg67v7KIzzKBIYjPzf4ZEIYDE7e4I7X8YK0+hpNX2ICngJd0
GcIM7YYlKaypJZaFwAhhqdJyY15WPOEmGkFkETBZBVpewaAmPMkt/EFgk2ef
vLeoc1a69XRqxDXsUeqy+IAV49Gt79wkuOdY4op9tI0QPtCbgpZADPuRkOgn
SWrWQXFGfzAsvk73vWrlBka5ugVWOoEmEemPRxe4/lGNvYna60Wr38Mj7USz
iBCsmBZdpXscw8IflOWK9Ls39fQ6xZOZuCVj6+Q9cBmdm1nuDai+IR/qlKwn
1H4TxL4qc+s1YMUFeiNccCgBiaacLdzo/oA5mmu1IF9R3qquC+0r0I1sQvjq
uM5HjfYew2Rlbs7kkG/ZcxzHT4bRhNfBhm2J6Aw6jM502EW7oKKaPHP7bg8a
ljLAS51Ux3clAqO8P5qo4a4krvpporH2fnCW67jQ93+cHUqiXjK2YZOKwDpB
W2OaLPCUVIGuKjP6aCMCHj9fC99OZQXTxq7aoynnXPoaPv8eLpXuvxMujywt
2r0vqStY2dbbTohvDqjgmzYger5tevO1Jcb4wEDvKsD/WWGJe8zesbasjIYw
qbKTLrCtHj3B4Bk5DKKV0tkateiUTyttC3rd5TB0/t2P2LDrkSq7CNMkahiV
p9xMGmkY1CIIA8qmpEnMYYic5Qj+ANgGInFVKJ52eseqfZld0AGd8mn6m8R4
uRFPvoy8WCMoBojgGF1/4OeCjAK/6I03AhZuauZcDvIDL7Y9scIovTfMO4ev
eexb4h3as/xgA38RxUw+503841rlL8jTUaKdNpBWmyNvyihdScijbSK9IXma
0r/hcbezKX8Dyzb1IYrlw93U2rpmdft0xMPOQuCUe+IZZTb8pGk+23NviMol
NP6w/ggIZsqLkc8dfjGkG55J3bOcevaYeUVKqpijysyAQvUkx6bs3SIffGBr
QLdmmBzhTFhqxY1MlaHL7NCD7MLoJxJ7ZaEvKg0I4tAZ2W1h1Mbkh0u8FaN9
QPJhHCy7lkVjrn4N5hrtQa3u/I4g6XT/7uArR7iFr11k7KdUPXFvAAB4E5cn
t3p8/GTEa6jnJZnU8kso7luLMwo7vxLeRea4kq8D+487Aqyo5zm1rBspnVv8
O4ZIcdALsbu8Tfo6Am8IPbz+6NN8VWP6YcwQvwLiKsykpPuo8QPBt2F7Wofi
47++DCFyKZUAmSSu19ik1JNRxCJY+UwqcQPA26EsOKZDC+BW6oq/r/TUExBc
LzWYMlx5ULSghKAtvXxeps01QI1/n7XbCNYZMyhXyrEx8jk1pu0UCf4EB8Pw
kE9EBayHQSISaeCY5zIiHgLAlgs/eNfc21mhrFzqXq1uG/H96dFhsPfzAQ9t
aZnpNqjDyCtUK6Jq8l4egrIZjknpF6DV/nmtWDUfSQbbpftAPCV1LxmVbRn3
av918Tc+jlol1wtUEMjo1wlYNmRGCjZcj1D5XO4/kL5oWeyRE9ELqiTYnJ6c
W8gi2M0007j+ldGQ7IY7MiF0prEboJRV9dmYJNWLtNnp0YhGTS5JebTikWue
l2p58dIpnKcHfaj36F2sRlMlXqK8lWVjTzfJSOAnaN0dv3vo9CjTzY8AmeLi
HFp/GE5DSfWD+/lqSZnYJl87psXDtS90d4H81GCXDh4k8PVMCIqoNKe/KKVI
NDVurRq4X17e1EPUMv8apVuRXJPhR5ApdH4G+uQjVfSGiYgW0EydmYxYMNSM
tujNUuNGfHojqfqR3v2garHqTb9/H8dG/E9QPoUxyuAOjpPh2n47a80qbiaW
a4bJUN7jT2THOHXyQ1Y70qFJnk8Ezxt5+QPM8Uym4ZPRbo88j1moFmI/MKRp
NUTmi8608tRzyHBOhtJAGoJEi9mc0jf/n8GV6vM9JZEfxjbM1NZrrYoaB5Ns
/7a2rKwv7gi8NDuHoI5Gnlp+DuB9rm9ZCUyvZp9lU/Pd5P6z171Xi2WdZRdT
o9KfbtHxB6jrDP+XI7Y/7/DvlugppjlAWgurzctv6rE+zKgaUa5mF+apnoZ0
B+9XZY3irdYQ/YYRXQk12+/dibafcTv9yNN24KFuZxLJ3XgQSH0gt5BFwEUy
38RqDxxEkhSEsZBfNWGkpFktzyE/H551N0ORveJezahL1Up13Zf4TJozvIKn
NJ1PIJ1y+wL9iZzYiw3v4Lp9/wv49/YW39QWXqJvPcNR6jG7Er+PxjahZF/H
FdbC6jRlMDXzdCMJD4NeLNxl0kJJ2nYbPEUzqY71oo3AVddUm1b2N0WEP2tZ
3iAd1Q7Tx08OGKtelP82SA4iEF0knA58FiAvSzYSNDmojycxpzpyFX/UF2Jq
yeBriaVpsE4sjyV1q/MxOm+Q/3Ivl0vxA40rjOsb7jzJrrPe637ebTs6fYoO
aRhi3x8gaz9+jW8HSt8/rcGtJWwYMxZph3dpbtIB43WLlCHMVmwxPOBXIdWe
+mOttefUbueCQp8/zlhwnHC9RVs2weA4YKDrZtFyzvd9H/Yy6yUjgxPH6Uyk
aP6AHSmJZAqFMlVi1IkQo24qUh2/W9dD17rHYgXzBsyg/vUwQEyo4ubz/Dc2
UUwmBoR7QrfOlaKZRUf8iAWjxQ90mJtciYwx4WHqR3i1+WNvX28SVaEyIADe
6xzczTm4yXir0crFEvQOAkGL8Xvfdt4Go/QCEDi5c+38bz+v1iJHk3NY6WEY
WLk6GsuVIoJ3dwtQ6HKCL30kQHcCECKUgPfAN+Nl3ZRpELJw/R65j/nHp1mS
gitTKuyJG6k38vjPUgpIYg/IhiHtLA04/LNgqGHMXtiOdab4o9qW7zc4z8nt
qTgFSQmfyriXey2UW6wPxuqoBQQpF5FjkWaeFqhIaLOoyA+8SKAVeb1jZVqH
Gd1eD+89zOJHGjOYpileUCRSkO8E26o7UssNtPWAtEgs63cZH3ayWqtrnxcZ
GvFk5Un5ZgNQJMmhHdqeIeFnG8MLBxbD5fF7XwrunVa3/27jIz/+BHCF+7kl
KN2RjeiAZw+g3VOgH2BzJC4TOUmrjkwXlDF7GT+TdZ0MftiWHlWRkbeqHjOZ
dt1bYW0MMBOLJUL76kIrRi928yeJIy/o/LvxWFMh6f4XTWk0Y28nKnRooWv3
6aP1zjkk9gotafgwpWTjUDWjd8LAKsEtfEOW9S/c0s4/pUrUy0h5/cLN1OIP
13htoeScGRmYMNYezGanmNsC56ru8fjshaQ/RgHShAylzw5YwF9o1ajUXMyo
qs3NsPKcSMaze737GMg3s78Z17SakyQXw6I3B/zC2zYd5pJ2LMpUinO9HwgQ
nvA2uCvSACAzU1/Zt667QVSbwVDbwIoWbXH62LIen2DImRkZdyW4NzFZeJOY
PKNSqTD4T61zm6dAAVRThk5/saBgIupjcakVIna0Q1YYpdT6AOR513XTd1dY
xO2QFI9M15EP82nmBNHo9RKar9YC98bRQ3I4W5DxFXELpAFDpFsMdHwH6BZY
b5ogBQRuT3DdGSNq7vCNwHAhfxgs9BQli2+2JLAVGo3gR1Zk7NvDRBTspWjN
CLb4wG8XY01IumlvPH6XUlwqHB6UHznbrBkdWDnVF7HhtkR/JvAQaUb5Cu7n
nYqsplm3xb3Zp77d9HkNvnHP3hah1rnRNKjOz1EYtWTIX/Hjph35qF22iMKb
+bvlv6eWdUVKt0sashGYqyj/1Nwtitv00KYJg5rGKfxMzJzbMNzqvP8Y6E5B
tcc58BvrlJA9/UHqmoxwd/Pyq010Mg/Kuq/lhaFSPpRDpHXn/p2HueaGYrGR
GwT2LzoX1Odd4XHlBjzUbgBr4cbep/DaDgQRPlez0qI2YQyERtcapFuIoTG9
T5pfclxls8BxpmWaSCVcP0JiQwF5kvLkWFn2ns9e8adE+Ck96jbw7Q7yPDxS
yI+SSFneb8tSlO40crF4kcIWlh55xTdMOOcqIT7SrZqQol9wP9V1guxq3WoJ
VMs9VebpKJ2szUQ0bFzndYyOKFix2JrGkEe478BmjOQCLxhSh72xkI3X9mzP
RLegJCVA4fbJhk6/VnMa23KUEarFRq4lOzG1hzM3N0tjyxjnS/rO10W7ESyy
in6Nn3rsP8N/QCDz5VTC4Krl7Ara1QEEUQfIsWVq8SSTexmb11+usqG5Mdbf
rPKwd4jbBdDOrmVMq22KaZMyc4oB0Seup1YI49bU0X+IaGDvNwdjLK2F5rJv
/xm4+GwJqRMG357X8mHUl496LKF1XJfbrjKZQQm6Fik/DMMQIVU29L5DrMnU
+7fhUYA2CYkbOMysI9bWsDMMGRjgJF1DvYVxx6lvNU8Npevk6pc76kg2e72e
Zqa/aJwx4nLVeBES66axs8dYQTQ6YthnSzJqk0VZ5Fkh3kfiFojwWNLi7z6T
2hIVBtCsQdh2zV/R/lA+cXDjKxS07HJZRNuPcNDNnBY6lNw4HvNiTndkUDjg
QeTcbA6Gc5d85DyqLRjzvP9MgjegeEgwBcz6WDFBK9EkeD3EV0gmr1U7ihNl
fWSfFsgoVKZtqgieLfs+/SF5eSFrQtLIUTDkdRRO0EctorKY0yHnRy04Im8B
74xkUrQujsMqVuZwSwrxG08rKTavXo9cxdaRebwVM+oc5zrj+SUg/XkwIyq9
FTA/xc1w/2fzrCtMkXgXv1IvF3O9TVTun6MA6Ep+Md4bT0dSVGT9mJN30NjE
DWCP/OKSGbePhz/kAG9shAT4yP/0pU1CcZyuZ+6p5m6LaiGVPwrNCTB9+nC6
iH3XFyPme+ZWswIFUXrxs7xOH2+QS2LkoNj7UAucsH1MJpnPZ3Tr4HKY0AVV
CBsjB2j6SdOotyFK0uBM71rW1kfpfj4wdAqDjmi1t1BzHs2ckoXd9Zxg5tKP
TEz6h2TBZoY14u8L4UJJ+GE7MuFzn3RF3jBJiHXUgIgcb1Cx5rCRWedHZeRY
k/vaD5Q7FXq1oPCebUidQQriP3DU9m3BQRr8lLcLoyRV1f0w0GTVDS1k0BjQ
PXMLHwxz0CI1TO0ED6XioH8gl/kyLkZv4dJgQFmzX77NSizmAhQOsxbUh1ek
UCZxvS/U8rNyZaUi7inx4i6R0OlCZQOk5u6B1iWX/JiHrHBAQROeZowz1Zoa
Ou1Ln8x8Hok88t93gEn82Ps2M952+HWdoJz7OlvqI65ocufTzsEziKipDS2l
du22Gl5kCjiVHPplDzZwtkHXFqhQ+SHBK4KzQf8fTnJVkDE9pUTQQHVNtmE4
QMPG9groKrw36SCmYA4XT5AA7I/Ze+rASIlSWx7xe6Jd0Im7t1NrK+NLv8gj
OBBN7uB3qu4H/7XrTcahhRAsWXZlNwpFlt99BRc1gbdpxUJa/nX2bwoaZyaQ
PZz6be6YeV9gHHAY5ZAXQdXQtsXc5D0DYwITWB5KKDBd2OBoWoZflTpKHi5S
aWXeTr2VVSzHThP/xRDTem3DqRsUqXmmb91hsCZn3l/lHarPA5MM9P+r/Nbw
6Qu7GONtTzE3GVb2fAcaZ2baZSEnOu/VkILbYhAY1h6IEgFfUZu74LyO01G0
jW6UNMH/kCouyx2httZtQ7IFGQoth1kaIad8i5MwBv5+oX/McNrbTnPGVNnm
+bRr53m6i/trD5PbbjMhzQzC9nBVau1njAUozB8Y/HS+aTwyBMEHsHgN1y5V
NB75ni3InvlhVOxxvsSUJZi1aC+itBo5peWdErDR3YZ29Jrfcp+g6XkSAdD4
iv4+NTu/B/k0E49piwr2okL21exRG9UWDEh9d4DypcsdPC7CB6M1EBjhs8dt
CPGVDxgL0om+rWM6D4JrEVVeIgG7y42dBGf+y+bQE6PAuzSzQte5hvsddCkB
EPjbpIIAZuzgGw5Q2mbB3KWyNUHV1bjSIpnunR85VW2ePrE+DaqmCyvQRIB+
PRBnYOaAcdfkRTLy4QDaXGwlrJ4aBXdkhofTiGvUnI0wrlQ9iWBYOK0a3ENv
U7CYbvjsN0w69tBES3487m0AuJAbpMrm7cwJB6bREHCJg1IqhCWGes/ONvbG
fnVqBNo8n3OdFsnh/DeYwYyP+DWvLgGMsSJPJObmhTkM6GOQsE4IA1z+VBzL
VdNWY9itps3xH3YJS0cb0UGRV/vSiLH79Xzs/d3xxerpDjtuzYTeRnUce8+U
uWcVWYAx2Zt8C7AEqGpBG34l72P7Pv1EG52pEX7UaRHh3eoTNcpvh1aJVkTM
tkTFfrWBP/YKWrxKMno7cmyTOYtjoYyp7gJnE/Aw0cligyW0YuuqfSyrB+Gh
6opOrVW8yQZByDWGnQqbUzwCf23GsvW5E8V4VUdgLLkQKruIb2CKKV8boUEr
KXWK0jIdxYp9j7bHqSopiLnsNDmz/9lSNG5WVtZLFsme8Z98r4J/omRDlf3T
VmO7+Th9EE/kKekjV5AZQM22QqVYBSR8xMjyXN57rUjJeBEwm0rKs81Yu9DV
5FQhIJvDIEmJ/Z8zoJMpidHuu6TsfwLdbqPFqR2CqyUk1613RWLdHYzWWh+z
MaH6IaWRHZkDTji63qigt+UnB8HFLgOmqLNEd6LohkrzNHLBHQZgzfeCET1d
XPBmNvhkaZDM014+M27yDG7OYw6N6VhR983b+w97itESFuSdeNjWPoLkqwvu
iomxHJnbHwxY8q3oDqHtL0+iqTGYQKTbNc4TWiJYI0G67igNL+wQ8Uu4TqNe
sszP5DorrEwSxRe+JheiTdD8P5WDRuKdT6oEtSqujlnbRI27EZSCUhI9Odj1
6r3v8ETJ5t7tkoTFPloVwanwCjjKmSONBahqNLdXM3EuDUTh95uyKaDKz/Xk
srHaVQS6rkVaUtqymmJDXMUHTYI3lRnXkcSFYMsOgSmsfETtXCDDNvZKloj6
6CLAZSEt5sLR/h1BM0zuJ4+IUN6fLIri4u+ScC/EO9qExPRIiHWBtNAjW3zm
2qVzQ7pXJ2NvoSIT5wgifbl116nTabSIW/a6s+CMcbKCKuPeeruZuiUiB5Ym
KXTV3bJLeCp5eK+VFKKC1FelQA2RJLNdn87b47V4M4PDmg3B+w4co4cOlvT7
j4YKQLSc8VAbzG3sbXk1jGJH4aCdVUu9At0zUyfoHf9nKP14B3gWmw/8HXw4
Wy/3ELOkQ8xeini8mecAn9aYV4I0ZmYIKMbh/bLytjtYOfQWUJUDvTE4r6+n
LHKk0yX1PzCz2F0TP67QiOtqhyCwmvlpxUNhvTOQelFx+W4VT1sDEF4hMe9J
u3AmIG1lrNg7jQcoUIevdGY5W329FgYIBYM1niI0p8rKIgUtHRU0pX6j6I6/
+T7/OKFuaFPvbU5EWf7Ay0fqF2UWuj8K+M+qUXUCieKKRZ3OH7GyQpp1GMHI
2ssq2I2O499aXnJIJI8WLklSRBBo1NxjpYa3JBF2YYpGH20MOY+pXJ9N2Rm1
xxuWxAxhna15I3slOuM9Dqf3VSLQMXE1zurbQKBK4Uj34K0qXGcFvCE1sF61
R27nrZtQHXB9S9kvCwNmdWrTpOWG3mQT6q76zwkyc/tPGyiCyP7NxvEm4FHV
v0m8UF3Eq14PZizM8QeESjrgLfCNXVpwi4kr8+r7jEIgX35nQKU4W1y5RSvp
hjQRY5gCeeIX5v2k5UbVGk/liBJFayDQjuKy7ZdecPLpFF9DYwVh/EAJF86Z
vI3yKYF2yVI0Rkimkcwcec9wA+vbDhRbNJ4Dqg8YlOprgP0PnQT9Km3GmZ3p
xxSV79//TNYbhX6+ZDUDs9YghX4nSMjonX0O5jkhD1kTB/8NOZZ/VPeWKZOU
uvivMMZB66b1vCnXgNEfuKK7NJC1eI0nNTSUtav5Zx8EGwxjF9Rtbb48yS6p
9UL/D8euD8F5BKIp6s3iD4wnb8mHsuHEPn0TRe3Lv6rKEh+3GbvfedgmMILH
yv2rqUGx8JFYXLIKCs4nLNucZXiFPjArOG3lZGBuD7FGWsF7rpO0Z6mzeZqJ
XGqtAk+nFNmQlpNWTJKoEFlJ7KehU1H55J+9FkXkFIUoi0bHzHX5xPxvanYb
LVfBu58pxKYrH6xTPFDV6KhR2nFiiswqMvz3Ygh3XNk/0/2A7t3rxqYzieV9
RAzGA0zJGdj1KYDRs293VY+CiUEhcbsNdI8IDAmygGrGid8uRmWGni8eC4qW
naOeB4EseJDvTT1P6R4WTNinUqaXimVsu7vN+rdXkvbQq/WRA4wNqzFzfSlR
+vD6hL2x7LSqkB2czhuHt3Iuwze4YtWXV1/Zht14qk/tom1rsvgxYgUAXodU
OjnInnB/l9B7QenbCkFgR3zWyiMQAB6kq5Tb1/EUC1bRMqf/o/FwQZ2MPN+N
3s8wflY4M3xDTF+tZFCAhR8E9/rxzRpfUQ8FKDbGehgkKUn29vuhVzBYRLgr
2w27jYRs5ABF89cwG+yr6pFrvzVm+UgZR/QsiI2zg4eWZkc65BaaIdhHNzG3
5JZi3dAUJCWEvZNaPYOefwcl3Omn9pY/YGQfY5OwVKu+B3m2D58HlNHtKwaD
BaVj0SWNFfzz+oQvb76O5Ryss264lNEEbVLfsuAR28pGz1lw8YPDIj79gpUJ
+2g58hrgThso+j8a1kDoqMyPl8ThuQfBL1MAFZsMOqBf8a7tY45VClUHrMHX
qhhob9DQWf1Cd5G+RhgK8b3hCCTMGdksY9cD+vzBHbJvA9Q9pKSw0yTyYaAK
yrMyq1YFH7MAUVriaAr4Ltt2LkuFf92emZue95xYjb7bmMF2Si9hhSU/U8HS
C36QyNHVTbX9xA879ARXsL7BPuKMPbFrNzGLgBl/snMnAEUACYmqD+gwePWC
8Jr7PXs+OGl51mFgN0RXIbhEeJEcQiUttElaZWssdSShwqr3ajtjpFNyvVrR
2ewPr5xiXB/0ZuWrkWEBZ6q+u/KNwjB+QzvHZe9hrQxRbdp1kLVBTfQZFtz7
lYzTDXFmm64cddErBS9YLl31i2oTVzO76z6+UcCG0F7ahQRZjVTUKtlpHet5
2vQi3xWfBnpKZlxyjpRWsWc70wsfaWP/gyDU1pcFROk/PsOnIQHqdwv+MhLO
nAhSTkVuXY8mdoAyrOdOCrRZ8e4kw6fkSalrRf3D3BYkWLO+1pNeGcaEpGNV
QmMYYWYRuVTxghewoxbaV8Zr72czNT+lg4dc4sUyPro7q6UibwiWaRDiyTpQ
JwTR+39QQQdJnDvsRNLlN40upOaa3ExOdSjKtMHZ70/IMiHbMCicLGpytQ6J
e5goFGknjgvPCATV7C9I2u5gYQGHZygFIIY7uN/RXVVxbvmqag0u7FopIASL
zKWQO7btnIVQH4N01pmC6ZaWRHzdEP2ggRu3yTIv3EfVtBP/aK/4Me/i323U
4UaJ7pGDbWigMJ+NvucL4CJsMUxrPEXCQR3zS3T+oq1tiuI6UOix7TmG/ipa
QRQW9S1q99J6FMc7veVAwpZyMCe8RYOF4bMW289rRwDR9hcHg/CetrizPUUk
6u33kO5mlb7rpv80nM2ZHFQRy96MP3HxAP2WSz6gnh4lPdYo9d4zrEMDgxOo
sSwAH3Eh7EGqgUoEi81VrR5Wy55T5yY5KWRI7b4Hft4mGckGQOJnytOuwhOK
Z2dtMFQBNy+macaCaT9EJV50CsQgLmXopOtoPRI7PauujBzH64P5i1W+TI2Z
urvYLQoMRtK567TLsXdJ9cFzAZdQ8jFujvi28gLZo0yX2to0LsJjiV7U27P2
MJhvUfml1gBwwaTD+hAFIhML93cXYL2yCe+6FnWk2StiqtteuWWVWEn+o6zi
x/xSLbvcI+PHG6Xxph1n9qdQVkJD65JrDHolUmZY0hBwmxZYhTku2T9WZO/L
6UgyEYdCT4MnI3vBsRuE5xID4q6pczJjU7MR4e1ablhk8yl03E1ik8WOxPGT
c5p22CAvO+nrZAymSCCKw1moBqJjNyoNyGahcPHVLeMykvxv6+05m2fH8dZd
VM+zq8F9+gY2JLzL2qoOcKzt1WXSLwWqqmvpAp1MnPXPV2pQrP7ErShF0Cpu
YJGr4eBKZYFVLgMSMxYBlcCQVgK6oc5iHBfhO9+kVa3UwIJlQTqSA0feL5Ko
HGTak+dC3Ok5AwlvnfEWjIATTKlplqVq3lW2ZDuqxctzt7sWloUjBa/cFNtN
SnGSf7R4BZFHlk8sQpFZNKbaCcysmg9VqJV25EucnMq+Lwxe4nsxUO68S4Lo
Uij5Pic4s1zvqVypYqWBDIaU67k/u4FPJgjqoDERdn6nvaKAtf35saDoETwo
Ip2aPrf6yH4r9jR/qMhaaNoInvO5o1z6ld5WkgHWcNPg3yA4m8vYkBP3xxdl
NW0sccQfIaX4XGESBxn+5IaIg93AJmEBbZBV7FEekdiYP9w+Sjyk6F66ks31
SEXigb77h3n/+lXnx/6JTWk1tUvno94NTnVMuLYsjbsITHfx1HYQ1Em/qqPi
eYTvWzmYfi1nQFxx72U4mDybjtjmRXs0CahlGZ4ymtkkSQ1t5lbF1bur+X6O
OyVYGveqzvZVp/Wutkt4SxiLKctnPx+nFbu3QgUUC+QQHDXuq/mQ+gak6Teh
VO9TO74JHBfxoOZWssAK6D1KB5RP7QLmDcWPx75Qzgc3JMobCKazM21FzwBk
LJJSvYld4Sc8WCNX9mKsjcf4b82dsjidK9IQP+lzSYAggzb8qd33NAqFAhij
I3E6bRqZPiSysMr6Cvi7feKQ2Z66zIkZKujiC1Q7aimfVINAD9brvL/1suNu
jm/LpWgjEjLnCmAmMRs5c3slxuNjJYdiRzoGxAUmZojp3dDektqg/v/Oci3Q
oWtwq3guHSmr4+yCV0yRfmldVt0Gco93iwaijvI0KiuS7ZX5zl+l8kLWQo5s
9dUyBzMhyOL2VbUow4qPuqhaE8+ynLPrP2XZi3IvPDsLyJ+RMIBDSMZpn+rK
QF2nFiMI6U5VOK6EekU3qgCHa6CKx9CWNcUP6loVXhEi264IAbPJEufGSNDu
1w+el7whCuCunvWu9cSphMBD/Qai9NrRbx4oYeJzXMeeubHyId/LCjBT0zTj
xZhnFUn4SyCJ08rICnn3/nWdCXOErB/woith3qtwpW+VHHWIl4zodWQLRIda
93UMo6s5ZcZaszbCWwlQq49Qd+p1FSmoPKuWaLZ+A8Me79vzqK0sXUTlaauM
h1wIo0tXaheO032/0uEpi5mUG5zn4mSNZRp/Ifr6ln0AeVJPbbxGDJ3PpyQG
42J0kW3ygsQAOih5OTEpaW4e9I2JRN9R+SVo6ZV4/keqF64BFN3dNBEu0Ua6
aNQPQlAZuJ3I+9G07yuixKztSdUd9yDMP/vXA3EImIs2ruuLTSLWjXYtFRds
fK5N65RoHxSxEbiduUwuarWednyDx+2xkbNdf6k3T2lwms++DMfJ8FhIl1Rt
RMnE4oVnwNzGwyq8WCYNX3j9tMR0PT91jZ6yb4B2moiOhB49sL+NbxU07bux
Nbvtobq3Vsw25WF3w5ey597O/W2Js2fyyy0OCJbLatRDm7eM1Vx1TjPaFBe6
jg2OGbI5VaaSr6aGObn6bttF22/S46L4HK5TInyfi6mAtcO6UlUtRvkZINSV
KJeX9CRrKv00EMMn4pZ6ikeFyRLv2NISNj3hPMGw+sTwXJxOCC6ODMRCUF8G
QpyaTiDFijz88kA/14Y02wUSp6E+1J5mx0YeRJnHa0R2RPdD+Pteje7R3bDU
x2dm5If0NHGHugBcJjjyGYQ7OcSzM8P+saEWgoQfqKIZr+/IlbQJr1EmeZ5/
qq/nOtFn9MzMknO/Oigb91ZObetXG5bEbV+iElhsq+sXDbKj0eFv0L0qqXRt
hiS5LRBe0aHVS5FYCI8ode0tVdQYBzaLfxgmULfCNVhavOBK1rct4jf09qJb
ZxLLT03cOZnOo4DR7xD5VgS+BP6F6FfJ5H4erwyAIeEzCIFf+phbRflvbaCY
L8glWwFqGVUm9vMLmHeidePXsb2M+He5LbZAWCc54EDHSQ2yl0cf4a/hcp5t
e2TvfHwQ9XoFKv82fOOv2jztIP1cwl02m8b25wQllTe8/x/A8nEmdqmngsk1
fhr4mokhceOJouoWBUXXlRj+kLkv/dt8vO2tve8SDlQIX2GDoBO0+tVYpFpO
0xO8LZEi9S9XIqvDcgrRtV/w/s9aKk6Br4h//CE+tI6IZ8n+qqc0y9S/nnqn
AsB/TE+tYnBDKYiuA+ZTBSpZmUac53n6pvRChEcUnu5DBXPAPNC9AXdAT2Jy
GfPtSjSvrhvBmUee/j667x9S9rsjyqMdmnuTqo/TWT34Fv2NLy4WKoRSEHPr
cbSCTnEUVpv73RnaqdbNVad4MGxiRfi8ZGdbPDdH4ww5qVh9Aln+gP1B13Ni
B34FkgOPsbpLerfoFAMr1zNNzI7zy8NRvaiaMIKmMIB1IT5kvVssYCB9mB8N
VQEzHp0Gdwo4CR+uPD/inXCpd+COEkLdrfN2yXtoKGodAjOnA5POO/qigzv5
tq7RLbHy1upjF/xsT4CNgmnoTzagmHX7pbzmkImvnLxZ+6W8YRIrVvKrsoZS
zGqwgXND3Gpf3Kl5ID3jxx7gGLdTW5tpLUTxV0OZWtmu3oiSviZ/d3yuB6us
/8yYzhVeQ/UaoLXxzuVZ6YqsMZN91bQM2HgCGch8mirTSjHE32OzpS2VrsTb
MgSDfGC9uAvAPpENwznolKzaWSVNjZXqvum2nHGaNTvVlE0Z9xLM47/tR+dp
m+6i/uFGi/GFdkWWw/UUPigWM05eNf+/0G7wWJnV7WNLDgCuomTYyXODbrpY
/iWwLl8LxSw4lyCbSrMVY1hEIlI5so/hNu8W2Ve1kAaIzO2uQm5SWk3XzQOk
AiMJpSOKNDT+ByBErraDxBC3cDEP0OO7CTnEDRNxp2JKGNx2fDHyyFPwj6sU
im9JgjvwxQe92YchhLpQ2rcBKPeSbbONQJWZ66UduoEo97m2yJ0DBPtsF8SX
FmRODQ/cUkTZqRcaxsqiQlq90LUTvG5AyK4cdZp2hHe3rByBGcD9QsQz1JGm
tcsVrKn79y+Ozs+yRRYmVfv/VxKcEX+crKrZE5FdG+N0PZH+enSXFFFJ5xpj
e7bVFeJtJuFJcpC1jqDMJS4id8jsdFDFlSno8+bBfpogOl8cTKaAHAU54tB3
Rveojtu3kgeGZMFoC4E8ldf5hRvVVC8BLJFuev4HLFkr6VhMPclS8O+l/dHJ
80DedLY6n+7errA7N+GFdIR42++tRN9c40SAxMSUe0xJ8eaT5UF5Radalao9
FN5e2NOZt/Yr+F2QerGhOHWBbT6pRbflTbBQrS7nAfkZxpC3b+f+e20SgYMq
RIG2XcQemHGQzd+gaReZiQLZmKVWBeDT4XB1u57vRvLOFr85B6QHzGc42yaX
MzNGCUJfGDIVbxaft+SlRb2+aFAz0xp+ZY8z1smxED4R4kuU2kptoFdiwbBn
qpIjaJ7F46RMf7jUlTTzkLHxz5l+c5btSyyrMk9kNmI5R63JRClQ4EJlJCq0
J0lgAi1FaocG8xJmuP4odkXZYuoNHtSsG+XNgE0NGHDJY0qLyX7/1WTOE2Pe
hZC7XTpLfwq8SKCADZZpR1hso4sDCC9iBN+NzOFSD34AATc5ksxIuJhbXSmn
SE7r/41eDFQAsojyn5TKBQSKMDNUGJxkIPOM+UMGX8r1Ou9ijetzT1/uXBwC
c7ZcaZCnwTk/bmJIFEHE6XchKCZhCM+2cooCzjxFhhtVyY4SXzcUHCY60Z3A
66h4tbhiG2+h1E5C0MHhbzg7pvrnAXRfgeGqrnh3re4H7PUOAYA1wSdAeosi
kUlajsHR5F3TQD9GImvTM1u1tBfL0+ro2AmMqzIvu7hmIobByNC16wQ9mDW9
x0CUjl871Uipq8cnLBy/CGoy5i3HcOGUfk0tPHskKYNWejKePQqJHtUhAfPc
H4xqQdrPY52bQvimsJBxJUzfs8H2hACD8xQaCTiPUECMNvT1I+AEBqAIN1RI
ZYLDmw8cd5fA59SG69ZbD/w4XhqmefkAjLqcM/E9Qt0qHUkj6pahzLqxKpHR
/L5FuuE54a2h+CQ6AzlRv0am7IyKunlPYkGSw4pYivj9elnMOpvbqXoWZUW6
4P94LNmObx7b4Cw7RuypkgDmGRsKjgASMBWr1PS1ex1ZldANt6yxbRJYZFeB
rPb4jllytn8cKDrith6+l7QZQO3K1Vvbg4EvQ+ygXBuniPceYGUdY9jJynXr
TBU329IulHMcR8OtxgDwo+JcPifV5D4hdfDOEWxGUW+B4Hbp1p8YT6fgc/X4
9R6cOPWfmcgSbNxocCtJknxPGWkNh6mCc4+5QjoLEcNnULEIhBRkSCutdNBW
q5hoyoY8JHenE7mz1vWFsP9jfkwT+B1tBGoq72YO+rkK1nlJ2gldV5a43OXg
2ODPjkPd4BPL03W3131G7/geAWnVP6imqjlGj83lpGNU/Sc4N8kKSR33fyXw
MXl1Cp8V6NwVAhGVAEbXYnkj/YoBKfcwEmxvw+LgK1Cfo/48RhbKWEdrS2/s
ng7gYShFnDuaiOjiB4LIc89GfKO95If5fbO6XT7CFxZRjEbhx0/fTeEwMkzd
eNbPKZeD8SRBnK97mzeTuq2T6TETgS0E+kVEgyEDta0bp4EYNgpexaQ9EGOE
w1r5WbAJbovpCW52ExWl5lgH4+buATnRG8oH1YyNslSHgel5L/0UPyAdJ4LW
XCeMYtPKNoGFyPniDGMlfvcdTeTrO8befw41C/LqPgJpZdVm2p0VRNqeFbC4
nAEH+vX/wc/xO6AecCvoP01hGTRIlhMiUgH+sTIMJ/do2AIkPe1IOxW1Hg6w
I4c31nbxSnHz6PEjPgPrFg5ZXbiW1R8+LDuENuru4MnIRGHZkhQv6XArbkRp
I129YdTcvvF+THKuq1ZkjM1UcQGcemYrTYEBRG9Os1A0U/CE4gptFAG+ONYf
krZK91eHirvhrltCzFVtaUAYg+HprDccp2xZi8cExkH/+FDp5+rSibYkh616
xC+VHz90eEpWix9O90HmG06lpRYHLUop4Hsn3j/pqdhL+Sg5lLmuRF/E6y7/
c/MNdQ/gJe+3AnxpyPSwtAi7Xh1Ha6Fc2qOIHP5l/5ohtpwJiuW7SjHwQj8g
qyJaZuU3lwSx/edZwWR/2rzN6AXdPMQcbJJPicE+TKmnMvL+2JZ2q18MO6Rk
4+dKKwzndyTWXr8XdAa929QGNfrZx31Ue4nWdGgaB7F8pUIxPCdbYT3s4pcb
e1+0D1v585l55mxqKUrzKSbstzTrKCo28JPd+Vrbwo+asKiu+Nsxn9MXNN7n
SlwhDHo2pD2EgVdAy+eYdM3xEIJDUsaHjXd2e6xiHovtBIolUubETFNG0ldC
N2t2OtQy00arrkrhqapk3DclUUdldzn/Y9gQ67HZYQK4bPpWrUzaewrcD+xg
GAkxlf5SpHmC2SUYB/Zztn50SVGJHOceTytNx3qniaCQMCHyiAFHgUskGfhm
XGDD6CglyZv5u2/2VccTTb1eQBYCdML6VhHw9g0nnPyo+hSI+avBY8gTdvDY
v7aRyeoljyxoo7sy+8SP3O3+MMy9ZU3fVurSnyCZYclU58lo8mIWJvhle8xU
gAeWg8s1tZrJUdP4UdXFuQF69k8IbSmUK9LKuDLvNLsd1/vyP3qnzO5Z0OTH
YCoFMPZR941DN47LMqYaygdVbaqd5ASKMs9L+KhPWAlwUtYvkQ1ySXVPBIl9
MCXNmWuND/ppQ0yxOy/WZ75+FudI8vdiHmlpKxsZzrT0xzbUk9L9WHx2MI9o
qSyQqyRwWJLcEgkCY9kXwlgjsvGFpFDDfrRf73z/1Edy4KsAo0q+G1lRvakM
z4feuVggKo8EJZ+EwFZg1OzgFIL1Di97tKDZzO/1VbDH9dwogh3rntL6HIQY
uqdw1MfXDmua8V4xlp/FqUTjyXEo5cNbWCXVhR3dEqx9nzUOqhLT3lPtnnW3
nSertaGg+3VrW4rEoTJT3CWz/9lC0ecMSojwlC6oy+phR+4YSp+oTt1ptXdA
8PT/K+LzzGZs+HFwj3eacu8gV2MdETceL+qOZYyfv9xt2rEinPnYMfcj/v4L
a6Cb52CPkSRjVk/zLCZsC8juLuKwcxx8T5OPA69nT6pU0fO/ICj0AynlS5P8
H7F6GjsA7PjSw1f8oKKK0jAsPxlxlwUFDdRBYWvBd6VwvjUR4hGnTsUXG7i1
cDPhNgj8jY23k2UH1fOTFBLwraRMnrcb8vCIv6QxM43tdq1R0ubQppGeywuJ
IF+wRTaF8W9DDrD+wwvJykEaR+unAQ62d53+oLiDh4ylzQoiIvWdt4O+0sQr
i1RU9RQSp0Jd/AljsNGISgo3u/iGaTKpcpDD/s4ZSA/HMn145KuvR7f21UKz
fvWxltM0eQng7O0TJST+LswRPTwhizkZbu91fQ4wTWuXviuYEOoP4QJndN70
soPpxSwEUvYD0deJp9ZZZvXcxVJxHJRH3iUSvAllVw6/JJ9LRY5J/PcZk6GH
e6cPqdEJ0b/Gx2xcf3I4BIeYKSGkfBFX1Rn0uqoAiT5PrhT6WhIocNwUanl1
0wQXjlHpsEwj7Y8+3MG4f977k7YPeFlNZ4QC1y0CwVMK45obdoXRTswrn12P
UAwSrba/Nu1cDiLLGKN+WMJ47Ph0Y0fZzEG1X3/PD2vV3PZ+61Xw9sE4PcHd
CBeqCNocWA1HAauA0csa6GsEcis+tzJbrb389Gvrvh6RnUIcDzDRXlfOq/52
bFYqI1SUJvpBS+Xe/Un2fshcYrVNWjBiNImglt4MubMUkwWAGVlFf/Xvpu2K
LddSJBejahG5MFSynE3SpWUEk0W3WC2emOxNSIL+Ekc4zW2HakuCNADdezFW
VLMRZ0UQyaPXdUsXjb6gy0H0hVCNqtrKZqL/yrPtdEBnUt7CmyHAXxz4jGIl
FRA0AVGvNMGb4O620aaI0nvuG4Klm0/TEJr+fpLeb6ieR4VBHJUcOqlPalN1
gxgxvFv6fXc46NllzJ3be15MHKO8OZhR95OKk35c5oA6fS0SMBOrmUEKX1Go
4TBbuYpYvenQs8Qaaiv1jqg5EcqEVGIcd7fTDh3Mu3m13JG+AgtGJ/hkOIO4
9c/yWvdOaA3/OddE9ZkyRMw+hcVBQTUY0wodGC9OiEislA45MyA5Fv0nVzxS
ZCKKbqR8cnEHWEZm729M7547IaR0WlLx7NyTg5cNBmtbaKIg+DWmbmu4XZfy
sqqDx8FtxuWxkG8JnrdtqgzkGnPpFWAx/NVGep50K8RdDW263Cl08kjT48+2
T/pj6pRCfvkw5MJ/yNGM/Sf4a8jHo2O8WAtLiC8uFbuc8ybBFLy8w4R4RsKJ
5swm2iApj1kXQXTp9dNnYM38mhLX55DKmPDkPTDh/O6tPxUL8keRNTlmN5yD
UEkbvHskzXdMmWduO9zlrWqj26fWnrssKEP1NZAynwYmastBzIPXup9JMUjT
ARLRWIa2PT4zttYwafchCO9I3qK8X1UobKpd7Lw6nWQ7RS22E9JOZO2E9SiF
gZpWyedF9oZQxAYA3aKqELBfdWuxMVjiT8OUYPt+X7t9sz1xg/hFFPFAaRCX
XaPxxA4cER964dLyM2l7hCGGAaDzVuo3bENFL9l3Z1ySqXwIUugJdp2i6czG
W5fcUn8m5TEqIW1x/MHLSNmF7UWl4XYQmgROPr3ImND6AotGK7SkjMpjVTeT
VZOumtuR1mjlevbOYJYYrDJbOUsfAKe9RkPD4lKFku22xk+koMof702Xd1ty
p85hyiZvRhwPPYMPUi2+fMREuisEBGOzXJP7+AxeQfGjaibYX3iO5soNIJdc
PWr86bOzvN4nNqRna+9ZvpwDBlfVLKYEb9x/qrHRfwuf/FDaDIuk+98HqLwm
OTif9Tji00wgOw+AnGIWz26ospP7IZ/pP4fXXvi9QA4yVxBs1FNjHZ15hXgS
Y2bzWKP9RhdSqfId+gPjWzrrtsSNu1cGEAwTVuhx2lenSoxSKoPp9h/PY/v6
C6dB/TKQdgaV1jskasPkHAMkNiyvXJke4Zh8jLuRpGG29tgARG7lSDvBGFO/
BMnO0Ql0jfs3eyNeD3ieX1KSULZJz7fjINPtSklXvJ59Zs81tbb1iLX8F0re
hQQNO+fKKmts2WN6oh638p8QFmSBs9fEaYCwjcdY+pPVL+QboJscSSWtjwL3
/zTYKj4ygcel2U6FYvoM7uune1NPxdbx7toGIrY8rP3v8HMauDMKnJItXqlw
UIKkVym/k83/CMToVWvhPCzwpkF8IUO0tcY73Qd1sidJbHo9Hr1TfK63CmGn
3Xy3mubCkjviPLAoUhtVi/CQxeKUXBbZ2OzWCXCfBNeF0SGf3ibNNwoGZVbJ
r/iXWGl8laHllp9g2DXzdBwcOqCzYLNdumByV6IQHZTzlZyGaL7ps+/Wa0cU
oKP9/vzVksHkTxthBnhqC7AbxKNytfaZ+9sZf+W2eKRviB76kt9SJ3D6nwXH
h9wfU9OPzbaS+5Z4+tY1+OCOIi5kzMkKv00j5duWAQ5HA07JKJalGbWenax3
ikuZZ7OP2okwkCrRtbEZuvavBmxHD5iguf4D6yD0R0EztCQnGPMZ8IfYVX0L
K3/dznyZabrx6D1kGLrSAJGiGtavfC/p/7SB/VrqtxPJzxiPQRXWMYT/ncqz
flxdEN3WqTMax/ANXqDzjKE+l87+jbZD948BZkQs4kQWaNGjkLsaQuIeA7ZY
EQvjh92WjKrDR18AsW4lQcRgPAQn1TWKa/ikNSKlJSO1iUtxZkAFEdUutZGb
3aU8Ik7ZAp2XQ81VQCb9125eOh5t5+MfGgSnIlzRtz6dFeIiydgPW7m85Eec
bkIbu+mAVQpYMHaAOEsvtoP4FiAu2/IPkd06M8QT1YPdZHU9rYoNxTYI0OMP
ah9+NDEmVHzxZ3bgh3nPIowk6qdk/jD4HjIYU//YR8ZZ5sVjHWP5Wjjwfac5
QtHxvBq5/J1f3Uc1bwmT9Na41hSjRrQ0IeCj83FY3Yozol25UMMTVwAMgMQq
tg4Wh4XzjkYtuVbC6r2MZp2/gkQNed1n7n4bhDunYcEN/9y/VfTOxrDTFHih
hjHiSWN81NLO2Z0xXXg5gfOcbkZMfc1rVuE6lbPxxlX2Jb/lSP2WXyQXtgTn
w0LVsbqwuf+VPeng84TdOyIWZnTa1LnHC8boOrrnBKTJJfvRBWX8oCkAJXmW
e0mbikZHDDOMLYQGnKnGJcZ2xhkrBszJssiOMoD/aK0bcCWNfgAQhZnEBpSs
lFQgTCjax317Kh1R44kZldvSvvktn8pyUawBFGirWhSSPEEetxY/LmHBcFtQ
c5im+BOgdcX2h4xvWWtawRTJKzV6EHvzhm96ayMjWXkXGLBE5BjT8Mv0QE96
VjYKcufaPmezkqUUjrMCJW1R8/tQ9K0bYY2sxzoauV9aWcxrhmcxXCSawZL5
EHnHzVfugYpsFE9H+Ar5SFR/k3bUnATUYlB1nTPHMC5zyvN3AmMhkZuw1ADO
P1rIp0InzXWBYciPtHzHBYFTuj6ZxX6GDZ6OVDenhYShm+Da2bcnI+zZ7ee/
UlU60ihaep69g5pdEPElupT6DyToLXIceIWqr3NmzqoWreOAVDO0NjdG9GDw
d0XRBVjrUaiLoymyiCKjs8EiCc36xrHhTRaBPn+2dTBXd9kE3oC6s3EnJ/wd
QJU+UsjUL9s+1+B//tIA5pt8SR4KScZP9KU3t3lj3l/l6GIaoeZ+CZqO3FTl
dqGomOUG6es6eT6T6FXlXZDCWLNJmiT2zCTU8O19eE5TJsAv4RA/z2BFAJms
UNQg55PjqC6MadXE6EC+daafMMEhw177Zl6CLurT8Fucb7HrEe5/EeMYjdfx
dxhJrZZi82850jndVP/hPoJ4JDsX0CgUt/e/I4Gd1PLCWhW1x5Xm6yIytHSC
QUCXrka6fPyPCZf/czkp/7EW4CbfAnMc1Gt+ehNVlhaVhtdJ/OOn06E5atMZ
8Z0g5mGiAt479afe5vutAisZVr6amFLjmmPzo58lJhT/YhzVDqYeWMOorMZR
kS6+92fe1sSsVVVlWICKVkmaPw+LljC72NRxBV+kEsD3vlYwo+bCgwFvCtlA
U3mxn09sHKO5howFBXV4DY+PbRgz0YYoaYCX8UEgT6ccaPIO7LZx/vPpt9sh
BvSS+dN0RYfKMEBg2p1Pj/QlmXPufpZ2NduJShf41j67aVjO8C4MPmf5lwAi
b+O/eKgjszWsr4j6tQeGk7W6pFkEo+BWYLNYV/O3xdn/pOPptgXkPfQ4dsfU
S5xbG4szC3++ZN0EZLQrVWkScwiA5uUmJQODlyIQ3byqqBE4da2ijUaQwn9y
c1wyXyshkugqRRiHpha9N+y/kqnyfgPpyll2jyqZAUlRaTw5hTSIIjlyYznp
pgcr1bmDRJkcn+fol+qNi4cUiOwsF3Q1+tNivc8V3IYeX3zHl6yQmkAwV/Wo
CbVunZxQFMJPwh1IwRhfaCbzPwU4vHZb/GPx7m+5nX2UOV95kSTjVn/Dadjq
XoA4Vp5o7G3wfrhhxoXkfLvqoC+3V+3cr3Mo995RM82bre5Q5Xutw2F8JEtA
TzJAwvWNhkg8VMlZZ6CA8W2q4wLk1CNw1/lbx+ux5YHA/BGTJ/em23zf4H0/
H6Cn5lsmSoidRISm2SNnBWkWBfy/nKVuY46rU0KQs1bBTV3Am/2m9c16oGVh
DYgxSm5QLgJOaXPE4Rnnz5Jouv+m0pDYov3j6HpAOCSfre4SjFJQGo2NXq+H
VMo7t+2SYY6OFzGgkXDMlojytfWAB34BwFYGZovkxaqZpOV9wEkvCbWAo5oC
q2dR4tDoNd7xquirw6ohOCfltfjg7mkj6EVFVMLQYGE1bvFsYFWvfPmhqnmK
pRsyZjlfz62320wC1dM5HnHChxP8lNjHjV6XIfrnjsjjHA/JxzFHJjSyrfeZ
OKY3UcJQt91nupieU56EnhFJewf1H37Xyt4yZsWX9euVrfbzOB2yz0nYeAfi
h0WZoxEcTcZgkFkYt1KDkxZMwLVeYD3i88AedZ2NJ4sHSc5fxignx28aCP2H
5/LWzpVGpp0Yq2w+0PKT3/6m1MGk1Oz9eVGwbDQ1RddstV7HsD3LVNKCt12T
psktfZCgO+NKJ5KakOBriDeGLxLoLmD1bKz3kuOAd60ezMMI93B7KrlNePAT
daJhW88nR2b2jsV5ooKuHY2R63qxXWrIQRB1c48AU2mXQgJKCs8tMel/aMzs
kg7e8E3RpmHAyJmfRc9WT+DjQ9/wNE1C/60R7PTacrdi6Nx1j3yailM5P0zY
lGPtzLEBCbRbguRfyA2TMjIsRY4PrM81p+0lShio5X7DHJKIBk/CvOvnmTFF
uVgRM2b8Xu0qYuHXoNwslQ1EYHYWDgTsrYNXqjPgmZcrl8Pb/0WYzd00psni
By80y3JDqWK5NjwfWXcvlfCbUlRnmhCoHFpHy6tizVDUhamWkRRQGcY9nQ9q
jwMXNd2mVb4D+G8fVBFIJn+GJNeipTyXEYXdUGTsORzbanbVZVnYwlix7VjC
vUpeYjDZAgJF0h0+4gAqYcoF6UBC6T3kFh0q4T4Oft5+ErRN354Vl6T8+Eai
Cy5wpwP/M9112AWhzW7YINPoNCBOubd8MNPwSV6d/bsO0X6x68gmyXGdAx1y
XwcDBp4oDo9Rzx282VI1EPZpfM/xaJxDhj4Fl5gzf2iW4ihjrg++AsnyC6B7
nVALexSi6DEADG5BWke6VB9GTEJ0ns5iEgxAw0yjW9fbgt73KU1Tcef25zIH
OBspJ1H5FuSrJb6xnXI9eXlp7inJC/FEqpT3V5fJ9q7DYcZGvgXU1VFGEYl1
kOEfQqOL2SCTxAj4E9L9yxawDXb5IIBN68KpAxHq86K5pJ62Jtgm6xxcrVYM
7F/jHmHXN8I3JRAWRlVLYhWs2p6/fbJYkMaxq7hq9bIJysYSTNo9mHRx0kyU
hjUek/tcT0ZZOF4DbKp17F8bHmHojRuC419Iab7UJoNkpqz71wsfrwuMOu0J
Ql6yC8YJRt7kDE/O6q7T1QENNBEdV2ADzwU2oH1604+fUmqZzgarW02NVUwf
xnphkyEPSx2nBgjwAdarqWug4UrJEbOkKsyGhldMCAoQboaw+k8/Sv2awK07
G08EGABw66sAZrxmO7EksMGlIWTzK3xubGGYxKYCyznAgnFOizpvYTayyH0g
e77rF84p+l5+956IhGkyRZbW1EqgXtVxV+fCzpOSolMp3vntkFRBZLqZLEz+
bbS5BHnQAKfG8dih6TDbpYdmQ0WvoZZLfa9K588JXaNXvgpy/p32ammSXO83
/4lurm+GcQC8Ntofe7Qnd9tf1MxIk+UBRGbyf7xVFE3gNKnkZWefSQvjXHrs
etepOmUdfJBrWFSp/sL14QNr16nIyAc00yjQKeI/RYPAce29QHeuRi/v5NWk
Lbsa5Pr9dgMbJwD2lUAkaCPfi5Wv6DcIGbUxUoW8XUXai/9kapaUQp07h7b3
DhyQdTFw2K0dTOaNg39du7ELdaY4RSNGS7yatlnIqHMQK8DbG/6xYe5/lln0
fCIUqciv0UFtrSP21Q74p30JyPw01RdXvmaBstCErkmQ/QxO/UklFKw2hMfi
wK35KW+W2QMcMnVSF3OaU79UPJcaafyZO/8ph74x0i321dCmMUuxOQqawuAo
izc1usC9l/MyXvrrrqlaDajzSFd4ksfo/YSwtWe+p4vGuZuJGoGy4XbeAumv
nB06EIQfRhOjIrSdeyWnUuY9WnD91hJlfkljppN61itCt157cjNH/nDWNqSc
h9GSflDz6Yq94WahiKFRmJ5N8idFDC7q4DsNKSsQe6k0AQwad/oC8pFQkxUx
VQOUxMvAZBWEV6rB5/zoGebfwKrMxz3qrQDPRrqpwlj07IogmaqmQcC1kdmv
nDGLHnZ5k1DX0ot/+9q0ANIRN0WXTSZGmu1giR4lwW2liBKZzSD0xJBFvsnt
yS5/NAFIJwVsMgiW2iX7FTjvbUmOgBpd40li9YRxtAnSc/1BDRLIrIPlGNnj
svSXm0Mwoonv0t1NhqMnr/RFJfEQTCD+ftxGkuInZDBy9UGNur1Ai/KBqRey
IEc5L/B4JVLnURTI0gKk8dvWfhdnm7N6CYmiPLwsOnyoZbMi4NPIIEqIHIEE
/L/RqD42vliCoq7x7ILBCdgIYNBm/VkzQ+toYcw9BuwoqWPf3qHVFNbJG+Z8
QL2g/tQWdXZocZ9EdK3ty2bF6R28WIKcPtczauYXsH9/VYbL1NISsHAWRNn3
JyDrO/P4OAUZ8FwYVkd5UzkLzE2/XLOFSyRNCYzKs90xdOKffhDhFgjMluMx
K0yNFTK3PfYc9Sp/zCU0m8IuRx3NlOdbmgM2VWuXHBux21YT3/8VIkw7i3xR
Duk5lgiy2SeY33tWzIVO4UIt8ozqi/nglvnt7fa312b3IKEFsv+5b4Y2ypTO
GPvQFW9QxSgAqM8QQBf9gdG4xyUMixWZ3e4Ab8rtq/1v4HKYE7U+fNyJ/ht8
MS977pFbKCEnQN+P90MV75m/rnJTmH5FfbwwaX5GOGvkkkgcyMVuGQCs+aGe
4oh/NSkGu8euxN4cKCQO/xmW/yD1bRZ9tt3qYn8UxTuKwLQEGbq9MwycPcnT
JsGKrN3ZglESgFLfJoP0wMb32/hATZDqapcZOaY0vvAeKdZ1r3cJi3wHfZDN
KvKBz2N5/G+ePqof9mgGvWLysED+0zp/5MulvgzntJtJibDwpROMHadSm+lI
1145u8jArCLNHG7bj8rBuu1EUFVKjgrBk3JKpFpia551aL/Y6qBHuCZUZW3f
LivVv30NXAWk2kFCRAFu3O1fj3e8bv2UhqEbLYyJ66quURtcju9zBrJZPVLb
sBtIexK93rNQrs5qN1YZVn1++pNfKcMuFA7GPBfnieuBx4l+yRYpD56HvRzy
qw+t8m+TZ+VdaS3z9qXlwwG+MFwBx868rFqsenpeTNW5b2kMDaK6CcX2FGEt
k6lySa+qGdRr4eJOwoEx2xelGh7OzlRdeXr4h7LGMHVAkGZ5xJZ/ajq0U8Sj
zFsoSZr2ZaNKUpbkEWbAOffBZHKwZoAlCL+uhL4w+/0pOCg8vJ2BQ1nH+Ytc
DX+rk0gcCjUBbeUqAO13677T40YvqXZQOQpbML5/fukS9lFc96mzbwEFJBOg
NIPy0T1UjU/VYcUvLlvwlqgAnFjGjf82r+FI3l8fxOCkxYu6A66Xhzbd9foX
i1sj3ypt/69Nqe6Qlrjfsh+Qn9TPnxFH56avlImIHfFeBqo5kSn0f61EWuzs
7YGG3zUl+0dKuhVPDP7E1LM3miFpo41zTgFsbPQ2bgoaK2RZ/S86tO2G+FeG
8F3rrTpVRE1BqavtvYfXzR36MO4IXZv5p7pFK3ZNSFaX5G+1Lq7KKS+lzAz8
qHF8rB9PJ4jCVBiFNkkVIsr8peYEc9zjjRSSeqyW5FAnzdIEXF7sugI3GWEB
xe6RxkOZFcwpZHzZ7v/gN2dgB5FYjhznyfDBHNj0k0zYa+5l4LWlRjZczkCK
uToSz5mTWCkYh468NtBql+UYkHtTQpMgnFQlpkJyTD+7fdisHNlXdCMDLwdL
/5XlZzsRbROblgIS1DSKMyd58X20/3/ir240frHBkrfJr4CzNCqxCgHOLonL
vhFMOdQNQpXzLR93g6wR35NWW4Y3UTS89zlj8bVQinUbIlLMtg8Tvai65J71
1AfO5kUFu4aHcyrPlnUgi9vu9NTqEh66fvvB5kvnMOGaQ9TcClP5FYZbMrWo
hK6xQiegfez0pHj1xxdsT+SouTpjgG1sPbXvvVihAoudK45qOudXqiXM3qzj
Y9j5N5xGDUM6j9rUJMLiJD23ZG6iwYj8260i8pAI1SE6O+789glexpsJPtqx
RT80XjKeq7j9/cONBB+u/whhOMdWooqaTqtnaeHndhX99QYriQ/TrFCOORxl
XrlpPT6H+99SSDUYRva44t085xpjfF1S8SJUuTc3skemgsSSfyp73clWTOhe
c0Zr8SJVeMlMJxFYivpEYrfukpaof+67VbuDqQLAS1/y2q0Z6+pqMqyh9qB8
4F1g615jzVTNGlowx5Cfbv4sTsMrq3GkbyNMWhE1ZONSOCyG6UQIp94VOc+t
33cKE6mHj+Wr1UKrDpZHlCeGXJIzlN/M3x2YAa8NLSm1rQ/8iTNRDLqpWgLM
R31P8+8+KP4HKPxMiUyHcJKkl8KE75jYPwh6htUtWlXvuRH9l36EtWLRdROu
drv1B2W2fHbsEtMCcrDZp3JThk9YxcUf3JZ40pxyZn75efHf7TvEP57/uadz
jDPH6YoSKjbDlh/w5IHt69AkPDrJZ4JWXiQ1Xpd2N/owxpXl+vArMjooV0j9
QWR0Z9kA3DqEwYnsXjMiShNIuZsy1aL0/a9LfbwxXW02aimFWRt4k0Qut1I8
JHGMqZjN3qNp/Hg1z496DdA/l/V5QpKMDYp5MSL8uUzYs/mEWH/Q84Rl2hOR
U8gtDaVSAscwIaw0mvwN2SCcFOZ42SXT+p+25QRAKHsdcQXQkP9gkmwOAuBy
l7V3oexqErvjgMPaVzsZhJc/ELg1AFFBsv4t3V0Sps4pYjIouSUtH+VX3tC4
Se/PV4DYm6rmKjsMw0H7vYfp2U7EidWYueKDKt400yZgfKWPyJS/D7xJx2b4
Hp+4mbTddXP42UhUTVBKRGXjnSHMRQex0FXfk43Re8KU8l+yDXgJ2U6VUjKq
rXK5nXL1BV0ZEj/rb0ynVMtCslt1jO2B83C9WijQ4ZuxHLItLjmw2deOL4sm
qyktw2/43QzvxxBoCMQAzoCTJvVKVHXd2OJ/9wuE+gZa/rR4VqY9ouvigyRK
lYyKXoIR9aS/+QlnAH7qu7KN+rtTF0QQmomehNl5I+pdalttLTGcnZMb9hmo
iNMmILjOt6oyST0Gv2+0awA9VBtkXmyuCWocUz7eAOsSBFmt+YLPQFUy668f
Z7Hwo5DTAxse8QNrpS8Bt/YwSoTLqBpNaV5wvlguLWtcsvLQ9TgQMHwRGA0h
PMQBGF/7L7rdfIZOfgHDwRVQqQBZw0F0HyV63FUPex6bGSF4WWDRIn/u/4Ls
t2bFR1HhxGgQecdUx3G15ZqayjiBnp1FImpmk2RRbdgf2nwG62PiymGN+HkT
hfSxL4X3DTHbm3bXJJ/Rudlelu7DsgEQWlkhuy3VbMxHAmr/IwCSPnmIztED
pkdbYhE9VHAe293Yu5u2KQD4+wTKn2yMD2eX67t9ixzNT0GhClZu1EFzJkvN
JaH3Jk76L+D9MuiEi5oNMN7ULuQrKu/zcU+wCenpvVAeJvXUPNFWXz1H+mIr
E7hY1qexZaoSk48XDV3XdZcjGmxTXyU4Wu97W/YKhI4k4DyvNHKs1MKiLkrM
5Sa5KwZDNCmtkaR12xhMhSgizvdt8YSyaJjagGijVDGeJF4bJx+MaZVeq3el
bnsXzsYHfi2LGWJM2h9JePGHRyj98nkuHtztVjOmoJE7SNezGbDOMQ6U/SqQ
MZRzDDev8ubPvRbowGgf4+7aYCqNkvsxPYgdcLyaQyfzkrB6fuVgTYUOJXzq
B48kFV0EQlvM5QGOAGhTmckEPzQIFcJboC0KxIwuzSpDbY05ua8LP9YBsSgZ
7SX9Q6fjSqsDut/E7Ymhb9/8ce9mTn0WGZtOYneSawyQc1bKKU/22k+0d/mw
S1NQ3JgPPdA47VsX4SdbU0APQ/Nai6UXCzmAYGllHipA3obcYkIE7/bWmyHX
pHrMcSJa5jrezRpqkm4v0Fa6ZQ3YoTDpGra1dwRJ1RPjeEIv4Enepc3/9v0Q
Co3p3Lz1+cm+hFxmYCOZNW+jc9RMP/KIFnGUWNSYr1+UYBuyFnpvoflex8ON
JTJOIoFvdbVfMHhhU2hZReoSwHEzs+mhR03oOl3GHeBzAlIYBIMoJPrNfv5H
mL6qSWdDpFRG7mRoD+s2L/Md6zc4JYW3XPQeIoQetR4CbTAsm2D+5MH60K4C
QR42CjC2FqGe6q5i/0/RYzJMOx1tdeSO6k4tLvdmI5tnvrW2xz9MetVMOpaC
hJ4Ko+5ZMuHTl1YtHkuZHd2ZDr+A5Shqy4qWN5i1DDzEnikefUuvkixinSdS
AnZILvN6O6/GhJoSqk+JIH9aaun3GlmuLW1oKwMHLzU3wiBlZv2A3lkMD6cW
+OgaWB3eMZ/G280PiIBjvjfVM7A3DcTYLa/f+78FdEmXiLXSYei6xUiG2Vdc
j65BvO/9Dt2R18qgyrif1wDppojjNnjnmanWiWcninYsvH7HhEx17eu4F1qZ
z9N7aKX8zuZ1AhwAGX5fXaY8GwE21peFC0vwCeAnrOACUi2NouwatS4W7IRC
JpSXU1gFMPRzxSdvjCdJQ8aiN6Cjej7VXRpXUoyr+IyXQvwTISfqBh7V5Arg
8m9wbhlFxTxZTFaUfQqDn4daNAknnfNHT4rdIb46TiJzY0eNOFlqso6CpBdd
8sQWp+ZAkkLz2dFZwPH+DS8cSy9DdXo9b8VpBQU4zhe7JmgEwp59ho6fasXo
I+wvG2ihBCfXe+GghvbxLfw8tUpQvbjf9UZ+IsraryqvpOetmTkYJcoUD6Df
Jk84nVE+Ec0+EBOEpS1lCUiU0ioaCoCFhaxMfL9g4mL9oSv9bjzIocYeA70c
103NK/RSxUfFtWzyFlO8rNvWdOkoBH6EJgrXkoRU1yr534eIRcstMG9wWOhc
xs0E6dtB3pgyqTdvgdTCK8KFYBA2xGV50pPZEdU54lL1EwAWcNZbi+wru0bu
MtZnKtrehGqIE3feBClD+4TGiujYvCfPordH1xQOu3YOREvaVDQ3O5w3jy81
vGdq57eiR3PPYS/gxxDum4lCYKv6+R25cw2FtqypvIlGPJq73HeWKBts1XJK
WOukq78Vqx4JNQyvW2qV31/VN8F+gi+1TIeanCPmJxFu8SMUIFiQgjCTMqef
SzLs4cH9ft5TjPG4xFZGf+zWsMdWpnSISemNYTDeDSmrkRfti7DQS8dOsYt4
LMeDhBPUdBqEGcO//Cs5e8IF/h6qFXKFqPcO3VXaiFsJDZQuGHzPtq822TNH
9x4r6JzLBfbnY9dsA0zjILL0ojdNCXeQ7HZCE/d28gQUKdgOmL7Jand4AuUi
IwEJAJeJYTC7zGSVSBCCfVCQwYlSFex2aYYCxFx+A+DlGotw7f6ipTXlPO1I
bW+YIsXoeGIKD/SXZ72PmDBvgpUNuC6YVT9LjS3zU81DyZy5jG4ik1lEymXo
uPQf8TySuHsDSladaJANxTPbevxOZMbICJS7QpOJy9OoXG4YVL7nDDRodCuW
4J3UdMMvDAy0bruE7DfNrGTjGigP3YA48904JHJadOPhyz2hIqpfu/OpPAa7
J/tESNLYp637Yz+1pKFVCWlg3dLNXMV9C6IWOJgSKeozGb1H7kmE+Q3itOvU
B7kmnWDLH5i5BXlWjpDLWQcTk9Npgq2JvkLpLCE/OS+EffOf7TWTpezIcTd4
2sRHckcfdfUTz7YDGcBNhx6nTeB2JnfSMu+byC8QT2UdRkzlnVBZwH4T62yQ
zdd2EZVNuMjuxDLkUL9Y08C5KWSkSgPCBYIH9Sa7zribiXWsBxd3gj8PryCf
64ZSoAo2jP4OAqcfc7TNFXkfKORVNN0dVhI1yrGRWFzY+gLhj8NpcjQt0JM2
AHCabfce0Z+suFNqUWCIBwwBgaVymHEETDdY6Fup8gJrmCyaQ90uFRcalKrK
g/8oAeIcG9YDEFE0d3aOTV3p1cU+Z/a8W+PYF3/ivkjJjvtCwsVq4DzGoiI0
Eb712VW0GinRdYGWUvJ9ap9uGcLDvlAe4XF2+6q0S/mIjNcBEjO/ORQUMSQW
+y/Zdw0hu7mVl2WbssT5r0DgfpHBVrKGAWDGlq6t5KQ0R+CSl9SiGxaAwkTj
2YCz5ayNg5sxTyqlvG/NaMHzmqjMExzAOVaXIwjaZfGKSSwJG316pTZG4fU8
2eOEqXt0WQp3As7rBpJ9/nT6/Yf/bVBeZlm7qy+Tnxg7DUPi8msrGLN6+5YD
FZ2EwVoZxdB29jgb9NHMPZlR5AiZt4vOjXMjr6wn9Fr0Mws1j4Pr8ylNb8O+
FHgflZQ8k2fU5S9+V/aidMESDUgsNTj5QvTYQcZHGBOJNozx5z/GuecACmGo
hR8TwldaEtSUVZw4xODxx302r+uKtQBN/jrvvVnr9s3A0dAOXnHN3d26Auto
Rp4MOTd5RIuuyUmP7nG/vk4aUDRJ9jVtJQ7dUxZi9rp3sD/3d7kdQWMTeRax
6nKe3WvY/vq+yjt3wWAj1KK4Q5aVi1lBynCyeLEXmpSyptDfDQsySHkkqR5W
EZsPeP4Ejxv1wtr1Fb7AH/OtOyHTAbxf0FkZjkCo3ziQjgcUvNjFqpFcDa8x
9nzCuDuTzWRnotxMXhNYT2eK0SN0RTzJWDW7Ph2/RCx0Pj84gsH4KefbN+YR
C6Jm+BZF2QUgsIXGQ6e4aPqGsU3Z7t7DhDQoZ+zT+y7Pqyti7mdBisDDA6/K
QhnKeUym//vO+R8B6GXHOak6gCs/Twe50IEQn3xJ5kmi+jdmEeu1nmkS8Jcn
UzEy7jg82JxTjxECJoMbxzbPnPot9FzU5m3rrK3m9c5RvrtuPXVxpwH8hk1D
PInJ9AsK88Z/sodU3x6IQ+K8wx7ougKNciBxvX8YoRaC0XLuMD3a4a9PUVGk
1VoXvkZFl3xgBtNXXkmG9tdtqTSeiH5uYWOe4qE6itdjRaJo2QAHzEOAicrA
A3aMWLC5aXexoowqpDbkxPOaYmvMOE/WpbpSdWupbYzw1goDu29oMqMNPCpv
BPhTdj1wd/9m9qxFHensJbHs1Zoq00G96sKhnoA2tZXYVLx6/6l9/9A+li2l
CzYp9iY2kBeTUN6yX922ZGZepTIa2DPBohwB2fzhhUuJ1tSDqVLuWHNCLbiz
n1ze0HcNiUuu8rxsw8fUBRkoGdgL7TR5gL9Cx6hAMem2fNWiBpldCmqd38aW
Pjp5Uwzhex/K+P1SkG0X4i5aI6xDYUqkxWTI1hRryoiLrhQaPzSvOk9waKkV
RP5iPmOINl23GB5/1P1u5xsdr7Mwm97JkN79KzrXbd7l2Ro3N0Ml6Dv4lSAB
iCMGfLVlJdrX87C/6CEEzlfxQPfxsxAqW6bOyI9J6ECGYE4kKZoyYEmsrvE3
nTXCTDn4fFIIwe2PtVhmHc4tB07REwPPF9QocnU/SGRFSxp4SEIuysbgOL4S
1DCgh98/Lz2fR0fHYNeYxj/7Xvnl/LgiTAJI2zWkiTTl0D8+bwiNlfOI0PU5
j0MlIoajCttob0vB3cm5RHFqGWFYzUZsFhhXg60twsq58Rxwh1AY5zFkGtuo
tKuKpuyBtswympZ6j9fFnojFfhZEYdT6v0WQqvzxelYpTtmcxFC4+Nay+IWw
BUD8uh9/TmBr4JEdmNbEU0IESdZHfX8X3i0zMCdRuUAlyMZde8g7daP0CuNe
fntUnMzbQ8ZfLsjJ5O9o6ROSlvEq9Z9wR4eQ/cYHTDCoYTeBYqMsdzoy879f
wYhr2rFpII3vs1S/lVIaLmExbannre4yO77tsOjzKnH/M8BdM2ybZnWClihw
iDsfWsFk1iLB2wWYHux0OSwBFPDgeV0Co7rHbO8+PQlpQZ7WM9HnvlI9cI6X
qY6pTTfffUavhueHsPCLh9T9dWTpy4Ovbw/8ceVy3BaQqp3eaVoD6NXdPLdw
U0Ork4YFqdomiI05FencklvJE/MCY6Ury0bVFZR95Z8tVUz5lTmtSqu1vWdJ
6IwTEsbW8xV2RptEo+IDfTvxy8IAvqsGq0sHxH9xB9rFvQm8R6948MIpUNFp
M/tr6xICscVkCx6aBWIf8h35fPTtIbxMxvcbciObCdJeeGC3tf5PPN0GqfVX
1Tn9w7pI6o3XLDa4Kax1lq1gJeEBO/MNraAKkJER6x4U2TBHNXjttfkWamiw
9mYzuix8lh5ssXoF2wO3V9449r0Zi9PJVsrtVjexMyJF3h863OS5j8fgHnGl
yG0Ojb8xx2joZNQfddLsMTJYa4wkjBr7AwfabSMFfNNdwbepjuw/Cvfr2bxw
Q+eEvJr8RUbxRgZ5W9DYLt2vRTnDd29uPEKTpILfgG+zWXfonC/MhRivRSgf
qieFc9Oy02wWpMrtfE+wKBQS14rtKCoXS/wqDOqGp6EqNwVTu71J578hPuuc
wSjP44O0COwpMWbgPApSMVA49vq+RVYO95Yg563NtfKUt1yYB3szTirChWqW
w9q5suV/Gg2huQ/UE7UAKl1oTBuk5ZgQRncOFgderx1ntt/vM5jjcTgz4/DO
cItXgQKDOr9GE8rudiLn73W60bi2UFPsBMCllGtRMGdP1VDfIMMDu+bL+9LK
q8e0aIy9HnNWhHBvQhykLFj4eblBr7uG5qJKtzUP7YZXiQsv5jiN8eaj93uy
aF8Yj81uWTKyF3uvE4kW8T26i3mLoBVPYc6Nmy0hyyHdtXmyfCgkvrTPovXm
ZL2RfmEwjyCvF2YeHCPHWtE6ophd8sT1rpE51KZ/VTUI5gD4hgmraEgxjdcy
iG4DnFhgYr5LTI2kkNpDuAvS0GJG9a/HviogOxobAwlS7gH+nBqJ2EpTdmg1
D0A/MNOphXcN4YkiR//sei9n1Qh/RjZR6Ag2q+A0uPP/GCGt4rLWbmiwa7hW
87mBcGeLcYjcx4vTWGrbqJj16yPtLLoRytss13QFGmKwNQaJVadgkyXA+fLd
JtPKnd3MBbbdnX2jmAaE5WEM4vVXUuq8rwmmHtxRLe6GRpnCuPnDfx4xwp4D
xcfmczdl5qFFyPI7Fk5AWg08SQtOp1OF8bWABZbQfhp/9pB3ZtaPVro11VnL
yU1FfT+2icNoUDbbveh5A4kOSYC2l4SwPyd374V71G9Ph4hZUIYBejqwJgon
Gqqfl2KDZFCItOmGV/7DBvElHIJ9LwnkwPpM/g01kJHe3akralIG5AFQ/0ZE
ehum6ZdJkqn38WRXvvq/fX5LLJqQqJelB7f94iY3u5GQjNBh+cmXh0h9pm1C
xwERuBb122p/0YVm0Qp3sgPhhFflTCkDlO2Hr5LsraQZzvCaEHKZxKYwxC35
hLoS9WptMLNgCP+scYbE2j5T55Gxowdgj+cdvLcIdkTGHHt/CZP30uIsVgPD
dmo35WzhwUVVK1eJ5XdalKbf9elMEkFIS/BA9yTlPZbpJHijFA6PhqHn3hfn
9HtRzXp/phG3Q9qNxA5njTE6By37ngUwfOi6gKhd8lCiQ75Yye8N+vi1kCyp
0dV8FGECPh+RiJ2juH2Lt5xb9rQWhsIywZgvoLpk6vihU28amBcLOk4aRJb3
OfkjhT3BA37h19z6SGD9FBoWlvHk18rQOD6PgFCAtvqAuiBT+1hLrsx5cOTB
lgW7dzpjZX7o1dNxZWStrNwh6jiNEIE06+TkRmxMwrwctCt/LptI0wwlytZO
A8kdKJsDlRcCvBz6fCybwW/nhoZHbuEYVzrGy0cP8c8M9wKc4dKENz7EeWLJ
CS/7CK7L6oU34AlhgfKDi5FCWUdXIpyBiu9u79wTcdvDZAzW0YH8PboGos4i
Z5f3sLR0LEG99xHvjjKy26VytvVUq5t5CcYFkPm5lew6tsmu0iBy3ZZi/KjQ
QrneUkyIieLnv5QV4HS4ukMb836vZkMbp19HAaVPfHh2nFzApB5YJwwhVxen
IrUP2JAJjL6T5XTBKd2xovnA+kA8lXBdel51bHVL3ai3QEb2HVqxqc3Lpt7/
Xi2k20AFDq+Jhj9bLDGsBm0lASXLzI1BpPineOJfhIrcdMk7HFLfC6iV7U62
bLSjrOWNYgOLFJRS/YDyo0ySmHH6J31oap2B6oQpD/InifeCUUp6DhEILK1h
OnoD77H7wT44HxqD2R4MQiiCH79+Jd41N+wi2uXMOd5eVJwlP831GGz0Mxuw
XLZE23QEcceyafGy6Q8EBO/ajXSabW/w5RZbKgcL/nY6kQyt4X7vIfZx9Mx8
u92AT/1XXZPu/J0+QKHbBcFUP4yMCs7kEMClPBGmMEeMMhW2Cf8fC7QPi6VI
BJ+iWL3Pu2TRaeS+IxRcOPyozDpdGeT+yF/+iTQZcEINLG7UZqvqYoNv+WEy
IvEjbxukQ9thjtCOZ8KhOw9aUWCBXqhiP/rQ2u75ENIUFToUo7x440+4YLHy
jOe5bOQsY8rb4V+gMyLinssXAl7c1uTx1C51AQgbYq7zNadBD+ok8mN7GxZB
krCsq9GG7mIRIleZV5fKpA9xaHhgMIbkQ0G/knNy5uncaP3dk6uP98PeMeTA
VOJJri9rOkGQUwJZu8MILib8u5+mAeMYZ60rRE9+no2oI4ss+BA9Zcssk8Nd
u23JKcjg94VgTxGjYJxHIvUIg/K4rtrlhRlKxPjFeS+5b/jzypuS6xk+ZsaE
SI4axAkdumMbyyGBO23jIF63L1HJ+oLQY1Iubca3UV7H6W9JQsKrr6aSiKeb
yJlER1GOx47thZiBl6BXyxFv5ju0bYoVV+AZunISGlsUGJ9NNzBE1QSSQAiV
3ZxTuySZMQqulhgmkJgSXVEF9W66NlReqP0uDJJzGB4ruosqGANgq+dWtKHd
G28S4XsV9UEKVGeQ3Zxs4X379qEwPizbxOyckSbhgwLsu8rYr/zslNhjCgof
7EP2/o6O4qzP69O62BTg3bnIMYZ/ASu7tFYOmRbGHa9DHxSQn3P6aOLO4AP1
TgHJXh3fdYbHzIKHpLOnUhN6rdG4Qkg2Qtj/nAx7hc0UUe1Kj6kP63WcTq7b
NCafbhn6yciQGoIyS3gbVdWhZfLLRXpXGnFNiIol53DTpBbKpKo5XCO85MnN
7CDAbtbIuHekv/SzK9ygND1OdTtuhwbHawakLfwzkfe6NKR8S08ajL8k4Awu
hEoev/6msJ8sNIbkudwY6KXxdWixxnOzP5cY0Cq4GwV+wcIlzxVkIGwcxnxb
7r6p1ukoZ+sOlvqLfnyxMkMsYe6vc9Afo6JFdKHljq5y1Y6m022XROxKKkYD
dZCZ0oCwKS320W4W+5u1tRBhXwXT+x3S8Hq6kfJVoCBkN6HKwdHbRtrc+xdh
xlG5o8jdpWDEJJ5dOGk6JDBVoDNzm1DY/g0uVxbdiBbDOJbNgern1NjlyrTd
GNsBvN9g32P+8B54PalT62GF8Kd6bilq4se0U5vgVUX3yAWaWuzThsqwEhD1
G0cFnVuhDk5g4qJiIddpy6mSgdW9zJxj7ovPjL/lELiVe2rBRCCcT73Otrjy
3cThSkL/ipPfNp1/DpRGbGFhKwhhdnH5xgZorIbkNVdHVia+Bsu/BRwFUCw2
yCCLr02SkkJIsWYxADuS3idExGGdiS4Cwae4mp7ZUxFzD9pLmP4uNJZM85Bo
btqE1yaPHwTCfbfy7TfT1Af+lf9o42lmKwkKIWvFnca+ew3qs0omsqvn6RNx
Td0V5wbfv6Hs+zj8GKyDt83w2c9vO6beAddui1CsJNNDd7ra6OvBLrgZjwtJ
5nM/TjxD8AKmBjd1UEqEqo4HMkqBgbDx8Gn3G39DRnX5q09m/kTtx6U0CgMT
7KMJ4GyreueVlXDGEB/yfgLVPoz+JD0yqZb0pxO33zdi3iPZpNr15/ZDt3cP
kH/lktoILR0IeeWLx0VL0sWiETf4FXO5h3jmiUqj94WiPgFIfO8XCkvLTIWq
Go6sA/zo6yeqFKscrjWfOJRYyMeR6IXo7qz8ADcFM0ouCn/CwZ4doPdnH26k
MkXzJYloGNThLTWWj1H9XAEDWrhc2p2DUNdpMFO61xd9//he3aZ34lacvzoz
L6R9c31tyS8xygYUtDR5XKXp+G+OpXumH+aZ3S+OqDzbyY3tL2siiMEaLBip
FBAc0yTK/u6O0eAI4aP52mLmmgHOp9+PU4jpAwbTTHFa2mW9xKSJWqCSahi+
GneHfUJgiN3cK4QNnu80LGHq1MMMmcUUZpjWJcverhgoSI6DpFjCA8aBz1Ox
MTtXCPa9JG6lfYxrhSs5e8pIR4qhl/XobmzTS+YkOpYpr1VkDXaXhr+luGCh
P0Egii/QcwRtsoGGUmZ06lWv6D7G4rCj16/8ZaxXYy+5ida7gGzTwvznBJXA
w69AR4tjq/EwNHXo3Z0xHt1s488YjL5m+a8IN1qL2EQ/HQ3SAybAFS7tmVMe
toEgSBKuuqDnSe8+2wzmAdNaV8WfKo2eKurzg+jixLYMgUZmz7iD+uNYpOa5
+kbTvW0bLfQtyHQ/+0rJTaUUQrFcyG96WyHPJ3yXvym03GgmNyBtup5GMgC+
mkg4ny8NNsgmthFJSSBtMwxQMA5zSWDTRAVOPOUYGZsXLtKi0G7I1PaNzLeN
1IaBaE5Uh5sqyApUpTtYoPRBsmQfVe/tQQqRswHf8F+tvrZv2RaBDj7K3jT2
95l7nyvNd3UoxG/Uf8Kojq1QdQYeuRuhYXuyc7yR0Xg3L5n3LlQFyYQ2awgp
jnrhNCF/hh0xeIu3mqA3du8Ef7lD+tPVNIKlajbMrX56Vsvo1gb6FzixaMdd
RRk4p/jvT7OGHeKKsVSXPPvcZ9aCLUUZR9aQUqove2y4D/M/ZBx7lTs2yXFW
thxY4h0291nLZXo9c7R5OkleRxMK/vO5rcMY/evrQDx/7INxooa/f1ZwuTmQ
mmrWEuovhGYcq2Xtf11S6m1vasUZfAkrKsQ08G6LChyy4Sm84KxtJ2/iTqMh
33PRdSEZPr+AL4B9TjIoc2GruDQdvo0DtanB/aPU6FQQQVmuW2l2QVedX7wb
Ewhys7hWLhMZL+itmOy49/uCKFsErRRgRXKrRBLGlYX0uorcBGtTYGrDvsWg
BZRVNPCtKa94BBrsr8zN/XP1OKwkpd+9JsJ+Ufp0HLUaGbtZrErs3Ntbf2Aa
+tKvEdP0f+YeejASg3jfMbPmPxAr8ahKCOyycDsbLpAiLGkj84k/aLPiN31L
wGadKmJj4WojztE6HNy33a0q143UqAqF/v26kK5ELVqY0jk8pdHgzBuDV6cy
wx0s9BoXfRXZv8xjwGdw1qpu/hN7KfhM/i7P7gjVT/0hKMynSK8CHHJQ447Z
jMKBh6IeZupphg17agZMIrgwXVJn4vt2YTQIvyea1VPnlwjDopilgmhmpa0f
64Wl9qq9vHXxjRT2d1ozHIVJlV13nMphM5Lg0vrx06EgC9t9tUMtmt2Awmwo
VYM+fnf0Sv8oKbMimxVnk6R+U9FQ412tdTVMcsDhQmaOc/zDL4t08koKm78j
bXEzAwpcTZbPyR62zeKjEziFOVWrd24JTIzW/yvl0QrXjIo5DMS+/8/xMMKT
DRz4S0i9HFwGIoNLRBDjLK2Hs9g/L672JvpTcy9wWSkZ3MiT2RYaxcvMV6ES
ICYp8JsrygxvLE7yKpbC+1vnKMCOR8Lx0uYqzGV1clsk/rnhzGOMPM/yUuI9
MN7PRGdKjX95N+5ezgMb4eLPDZggSo3WWmtzIg607qDrJPQDgVNdlzsh7S2V
QVsXKzUbgYLgT331hb+fbTwpVADifeb2712lzZAyXSJXwnmj3AfRXKt9qqiC
pHiWQ//+Bz8fu/P1fWYuqmBT05l/hCGYkTwCQr6zMpOS47c8dkpvs9x/de5+
nt08MUZL6h+Q57pRm28+cNc9HIk8R5uukWRKxFfb9rnuxDkDTAcqSD/Ls+58
cNhd57f022Vi0yCyfSWrg+abO7ZrLwKCwPGELvsGedS/v8lpVaq8MkrCoEAX
LYl1QISkJb+fxnDTJfSeWeCtya2f5I8u1K5R00z37xNNYAgtZP18RR+sEvf8
cuVC0JL2XVBOPG91TzY8pWzuAvxBzmbykvUWjojG8Vjug7p+ZoqzW4KjZrfi
y9zekhFTS8a2xYnkbU2BwtYlLx8eGu2GTZrpETkKC77FDCPVMvOPYDY12mdr
7yjuItWcdvPZ/nZLWUGvqtdsLSHxPHK6N2E2a1Q9GdSpbhwIII0FPTdFQcLx
0Zt3jAuY9mV6+bCJso0ysFkZsXOYJ2/tG15r7wbhv9oRC3nlkh8TbFxgIMB/
qLt5H0dtx8gVnqwk4dkMBpMlaabfNvnOZ6/hw89wrI90H8CNBYgYrd30ah31
NcDvilRGo18CKWtO84aFEHoTxlPOdEGNgBX+x0n4TFx+5ARdZqtDV6AhRxNo
h2ULuLyzBcCVwW8XeyLlkt+2psDijvK+5F089I/fmEvcxBCr3yPyIKX+5d3k
YekodeXxSvF/WyAwlp50WgYGjvQMW/YBGG68a5pUOWJ7fltr0/SNrLaRgW93
4waDOTJQiarOlvKwPJ+MeLYCUPyDkGDNv0KMjyhwuto1YfpGOD4+GWC+4/t1
7hDPnztOc9kHnp7W4otlP5/d7yWMQkFYfixatDuSL7oI6SXBH9JTZg4uWGaA
ilHGGQn8uiBqAUUw0rMGMZUFS9uKQnpIV/ZybSmG3Owazy1Pcd7aSt7btXID
GrM/6EY+MAztdWuCpWr8QL6ac1cBkGBsGuEKy95K8es6bVpm4KGGt2IE4B4j
pX8lKx2ID//mu464cnW7CeCcFwgI7PY9+uR3PkYm7/B1gO73B9u01/wQL+/u
9oQsp26ik6ocPJwpkNDPfoqqr3gZlwvmMuXOexWCyAZ3mMfWKwIYoRpjbFhV
xWBaZ9W80xbv2CchJmcYUxHhM1BNkbtdEr59AiYWafXjcGISM+RUv54lwKE3
tUdOiAyP0BwYuuKM2v7UvPlu7Hq9c+EJZ8sgucCM9Ya2g6DUZbzisRuVio+e
gzKIfdIDyFQzsRPzrKF7RwwM3edwuVluw4/rtswPDf66gO9nJpTGfqxFs9Ge
mh5JM4GNTwXfuW0cy0zxkVe1GX8PzIW+X2CCRq0HmA2urOHHLvHHfAXVLsHk
tYnhdQudAdasflIpIOOekqEQG869dEogseDymYUaXOZK0mUUdoqryzm7YG5/
XBnuj/3kJSlw84njfH41fk1NSqauuAD6NYOVe8Dv/2wXmnZamtJ0Ph6z4rDH
2u7rcL3BEAyM1hoZhIQmjnUPxv1BIGLg5/YWK8pmIEIJ+BUBdihCU2VH+dq5
ccyLWzj2zjlkKzkfuTmjfZ1dHUyVRJ3Sdk7QmAMkGRPUAOKPYumbOI6+2A5K
O3liYayus0/JyMMyasE7nAFgM6fD2H0iHAvwDYLaNQl/uvSpgzjAQOjKS5bL
/BCJFWPbt1a80/+yUakMqMcaG8eI16jm5QkBfKnNDJraKpaBr9KijRTjlK/y
y3VXlDhUJwwdOod/A3GWV/QGZ6kVoFjQZDX0P+YxiS9UIiUK3INmHelh1bSB
/gEPXS7H0zB/IQsxWKn/HvmhKAczHszBoz41ydmh0o4syDaH1K+b5AIDZJy+
lLfirflLDHRvWTI9KyPVzDy7QJUvMs93CbfAP/5Y6yRLCwOK+ve7BJ7SrjvT
bhi+7VrC8mUsZYeYY7CI8H8/OQnHHaoSd3GLQ0mR0D0MpuE7mOXnZaQGhgUy
Kjld03TnNSV8SkWAwvRqVfC9OM1ohSb00mMztrJN3Dir3/0d/CHFfPaWbagh
TzX+bjEBKDrrNOxgQpvlJcJKq4FN+nb+ABJ+0vNAERwb352/g5eVc4CXsoYr
OQy8pgzT4ejr8kEmonmvYE53hBGE3nUKqeduqWOQ9bhntrN5Wmh7f69OaKZR
NST7P0CXgKhfX4cV7RBq7ukg9rnK8Fl/o3vLuexFl7ksPMrjgjmrX7UAgfkj
chsK3vjTELhRaCNRnHD4u0rwGQMyfVJr1mIvIAX0ybRYP4z5g5jkWKatSsZw
tP2mmYDXks9zDBPm2gxhNZ1PSuz1jWdCQG+TzRYHHp+bKbfwJ81r8cJoQCA/
CHSEkn4pkvmK4N8DSwzkkR+3oS6KESeRmfaIus1MwvUexHn7SaLdwuylgizB
V6LfaOvD9T4mT44ClS+dJQaZkp5doFzvFRAbNVOoawPIRVlnboygOmpyF1zW
esYnV20OSGJSI3z/OrIPsZUTGG9Iz/JdRiwTMeI4jo8aVZ0+9n8LG1PQyx0A
6tZ5FYAjUVeVryNuI7NHI4NJ0k84ctk5Ou9Tdalv7buGB9SYPBzXUkDcSZ0+
7txYK5pXrXJzLSD+gmcJQcTWNG1HQcJjiFL3wTFuSRBFoeQBFxZd0wjBU4T0
qZPG4u7l8dYdO2TdVrHqgvT91jTKOavd5qY504dj3HbuM+qPshHluU+oAups
vosjGj4Seq9LuTt+ta/Xt7veDVqyO4OPWOMcKNe21xcjlpP4xmIGoWwmVWAH
+svvREBaSl8doelkukFUNMT2sF+G4wbtlKC5aiJ+iG55KJPq7sIN0IdAYd3I
86QWGa/YqsZAc98Ms4SgOR+bBiqIj5uvX1V+kduOkRBVR9um90BUjFJxW4KL
lPiZFvKu2kImB1laIpKq1M21+/sVWegGskf+8RGyfcFIuJyLh1XZJxrSyI1y
enzT7Jb0ucyWUGJX04e2HtFFrSgt35w6kinOLQ7jIn7lgS45kJQdZmiAAwFV
gkk7OdQOX4lu0PFjFzKAzDxialOwyIEoxoVPSfykjlPy+ElBgiOW4o+GIDrd
Qiv0Nl7jMng03lRkDo0VxBzGmOMPDPeXR8R9DagKPGNedH5mMQoPrzMmWojb
2ENCmazRflKsGdiuwO7ZcLDl+OWyHC5hKQoDlyrGa6Roq51T24q/wB4XwiBq
C0zG/KVpUcjvHbh8y2PsTNPnwkNcTgIe6Gd5gPOcf2vru8HNXc9SkZZZRVjc
10caMqMxstITDcnJDcVnEjEHSaQt9qIc+wi0Kkq7LXdm9xqd6eYgqnTXI1Wa
TrQOcjRwMdKNGtJo1cZitoeHP42yWBMMFQmHb5gFx2kEq0LfcrDSbUSV964U
X3uleszBphzCf+VQ/XvuMZQAPjdoFIQp/44vHky7ew0y7kb55pop1ngrf70g
Qj7/w4BUl6dN3QK/Fx31Cm437LAWqKTxBW3Ch7pA++N3Dzp95ZykOEFEQlkI
vBzRYkKzEXc1VcbLOIqSpQTwuXZoEX2fE/f+Vd8pjpFLg3gAdAVP9VrIOdiH
tnHnMQ9fL9mOnYU83jVuo97oz2wu7v7ae8wSlPsKcKD1HxcrP3eU3yZwExEM
9g3G526lxXunTXq9R4cqGInTS4rUCuJAVkzGpem8rWg4ufLnuBgWDsUc9TvI
QpDrEZf70q5Fn3gPU07yjes5cIN5HXlkBI9sjMdUviQ95rGe7N7vU2hD5odv
5764QTvuC8G5G8+8ew5UxeuKd7w+SUHanjv8nGOOXDNzbUNcndU55IOl01ji
fVwneMS0qi1S6gAQMi231O5jd7QB8cdhS4xMk4vwskIwu5j0gxEi2Kiuy56m
kCgzDfeAlk+AqtzrBeIMmrz+xE9ThxN18atYd16PRY+HE3jCa5OxQkDl7vt9
s8CHmSNcyMA4g6uiqcryQShdo9nj1nQENNV+FD953eCNncxNgYXF/u7VjasY
TlHferhZOo1+Y90kcxUa8vJfQ2mmBWPsixS/eNc6eq7SVb/64sbvRA35/NvG
q+8n/uLuta3bVDgDvjvCAGNjGLPiFPrqGoiIWOiOtFxidTFAyr3YJdgM9aZF
Cy2YJ4AojunLu8XMqfzqmUTNiG+Q0Eg86/hH6xNqNTsmkD/yY3qIxZytiHru
Y3suUIRL5UE57XiEHcSRa8JTUbnwWJNXI12VX18wY9Jelrp11NAMjql81RBI
R76K1YPsDfYu6gk1dqOFQEAevsLvu/5CP+pi9lKQALeDtYqwVe82lIFKoMBI
Obiaa7hybHezbjlAbBbXH9OjCUddSyrAXaczHc7nurZNkhYQiDRH2kpHSIZW
EMckddB+M14basIXz6dfe+8EScF+afFoORReB8ZiHQ60/elnypGUSVM6iGMu
Zz3XQrub433j+ixMuhHQ/33397uyIW2IVHFXCpViNsk+XDkKkK5Tq96K/1L9
cgPM5yME9M80dYdEEaB0BsZ44Q88JAMK6U08LndPB/vA5RCNBLGAFQCMOqai
AgdkgQ9Iq8Q9Bnusvz6CLqaUSiBQ52PSCq13eF7ruUnzdy6TNjeWOjxUS0LT
bCXEVaI8R5isi1eQ+xp9f4olo2tW7SyuX/mDTeeBTO/H/Jxz0PC0Rwgr5qcT
7gd7cr19P/ktxo8ILblmz6/UYSj8RKE3nLi64Az8nhAo5azdH6mBzFTyMUMI
h6Nue/5nlH591JQbKT7vV84zOlnEtV3fUPo4LWChy0frDShqpypQNera4Uoc
trXYd29vKCtRZ8P5PP5pZbDvii5MndGXiyTqEhIXZi2CaWM5rchOeZVUkfS3
UmEBnNmxK3kTaJ6PvPEHWzcYni8ghDzaYIiPn2KBt+F4t3OlpYTSXH/dqsTe
qOjlLFPAP2G5jiwGsEAABXbDKXYscX5jgfuiOrI5f2M4QGe+YD0Dgn7ZaeZD
pS8o0+34RlRqoYCOJtL6RJGA9Ll73HatLQQ9XALWmroYHwM3Q1loxfVu6o3t
T/rQ+TP5tKA/vouk3okhLP/z+Gc5KvVWn0LZLBT3YGzSub3rFvS9ptjJhA/a
z93O5HMXSKYtLe5NzDQCk8VKMe+y1jGzL1aIcnqEffP1wiR2TV5Qyy3Urvqw
UnKq9JR937VzW24pRQWTG1xmrserHX3akLSiRhbihR4IP4NaBmm2ylVj0fUN
2ORkNAi43Y1P+VltX2MrfQ2yMtaXuSnlSxyOsMMQxz+IJ5z3ptbooHge57gM
l4gMTtMluOsJkUdFum2rwGmsnnB6ivPnv9zTge2ngp6FDx1VTamlEwsns738
SkuIiHgPIZteIt/1G+xxyW3wpXddQCMDY6DTXNLZ23BOG+HWr5RH+ZySrW3+
miP0+kN6FwZKminYiCFz2/KZsNATlbxTg9lq8WyjgeO2k3/RvLKvoZ4b2jNm
7TdLSNTDZkA7pdR8dDThSIN98lSRMFLhK1RTm3h1GJ4x+T9FhjNvAYHq+zSu
+Q/PsxJjwtTsE9es5k7tCtx49YJp97H4lJn8KBCHB+NHuKCA6Ky2as+sOTGI
O7nkPc/r4Rp6FkzcORuhSsQfJ2DXOZseHF2+98+uGG3lNTwNG0Gugi266sz4
60Ln8RUyiKl8YN/HxSdaLt8kHSOHEFkD1uhtDYYYk9BCkaxdnwbbE0GlLQZy
DC51ZkBk3X1IvK7z6mD8kgu0LeUiaL7c/hbtqf7B7qOKAJu07YubJJXRekfS
cNC2j1/h3Ixs8JeYpD9XT0OPGrHe8/GT05ihW/KOoe55cgC6H9EP9OOVeim5
4riYwtUTWPGZtMDVYYYNgkmk1GxeMjhCjvvBNce2DyEIHe043PK7ipqEhooV
lwA0CzHr67oQFwDWVJl76626rLwQGgPodGA1RCSSMM/6Q7N5vJtucxBUjAWM
AvBTbFLLdTTuM9AThUhnLDbKjQrRSl5ojIQbjd+zP8MKUQ5I6Mzm+qZCornG
MtgLU9q7nXEwl3hFnoYryDzcQMhOynq2YgowHVIs1wbM2D5W+jHDDURchVIb
D+GATbBTkoHwZ4YPT5Ry7C1tPEw3u7DkOeZhCtby0hE8sefRXyDtF1DydFmW
AZd5/u6t+V45Ix2utpI6UoWkg7J3XsH92QdwkauzALJksIOzd8qh8PoOG80a
gCOMOpg44qwJ42gdhgHgZsygcWh42D6QLyZORE0Gbt8LTn0K8VTTPcs2nJ1Q
mB31wCYmquEEMOn+HrsCN09l9Eu+3hF29qthP2XxNzrN7gQJT5G/WnPR2EGM
/rAfobG52Gbfhoi+GLiqf2hgrd7t9TDhQQhZCj3pp/EhuHwhGsTbruDUNmpD
tozSVlhGDrq51cvyR05vkqcGuiczcvSa+ZSwexJAiBodXBFOp8wdfstsK8e+
s1BVhXmGZ9/rkXKbN6+JKGhyO0ZbHnm/N1egeaUQLjAF69HGPRDBM55FzRCL
/iBGbZnr7rdFDRqRHR11gr5nffVTvDqSvdXPTbfzKUKJpMtv2sfoyIeR55Y9
I2t+PbFYcYREgrbaglPCBYjVvJHc5LdXi26LOGm+glJkeU9ckdYE0f9EcmzY
6m9J9i9yf1apd3VPF5w7slpfzzwtgHUyTIF7nTvM8WHOppsi72Y8QUwIwFyI
Q+/Uv+TJJjFhQ31vwROL8DdJdaNQg+xUlwHzid3X4EcauY12nZWv+pYP7Q+z
24TH4fiKQINU01PmbbK6QsXGMOLsuEgtEGus7dtqxQQMQhe1Ebd7r5Bc6301
GQvD+ifINly3Zol4LdRzhaUay1bbO09FOM0FsWhurclXZBtrg7eo0F5O5v9S
nlgbFsBAWzRt0X6yM+Qv8zJnITP6wY/iF1mhVOvPFT13PcpZqG7RjPjlTxXa
rmDF+eUh3QUMOpgJ5vQTygwFPOGXtxtEfZ4e6iQNXZudfykfFIuROuq4Ga/A
gZawl5rGNU4/+/yioaDnd7RMUz/6Sj20mhToXxb1xZHlk5nj09IeQLqDa9/g
ymvOvhSf/M8CLtrWRiH+uLdyP/NkYbEqk12UI8dOl7ZrliZvMtuJDpvK+Fts
cDiwramKJomhLEnoOkU58FgYbeTuvuDABZ/Y4un+uO6IOov/KQc7luNK+aAQ
pe5n4I7/ZY6OY5ZmBlKaPcAx1MONsuFVzd5MkDbi5RIewdk6VJ+mX3RSCjBE
XPr63GCKp7zQXM5FUXFyP4GDB6Lfh4XsnD84hCvdtrgj6CK82x0sXB0C7Y5w
w3NXY5rSGlYyqq3yCBdljSrV7xMEubkBSPhZPzDhheDSAzeGgfvZY9/ngXOk
4j5BFl0oNQBpuoQckeSc5pyha30jzjjHdZYTtCyC1wcIN3ur32V5giJVU842
HrAZNC9nlykqw4qMeOAs0MeejP2cYiJFLNTm49y17vFTNSx9cp4XzM73a0qu
mRJOTEDnEdCEzIwWig9VDNCCklNeBwhaZ9heLjVOr5qNq2F/tc4vPIWYWmeW
aTrfp0ghcmm/FmFne+COETQhs4l18Gds5p8PWbRd2wbJohJs688kpMxcRai0
OowN3yJ9z3q6Yvzz2NvgxiYty5eOb5v6eIAdA43PSNsA14BfsfiXXhUdZwXN
BlUSIfzRBWwepb87uesWKDCN9Zbo1dws8IDLxQxMb7fuFjl/DVk27lnsFIBl
ae1r/gArCBAb5VJVGICfNtYiqJtwiEPXtktDPKwpiOgYyx/vTLah6fR+4CHI
F0vxfIE0jfGTCKgeqUk/JCsgOX1fc1g3tvcDHHN0O1PEsQcuxqgyxi/prCW3
A7moOO5UVZxJQnGSgHjMkKRMl1d6xuMjBP+7V/IYGUy9kRLDJ9d3/TnYi6ls
VvWTl3Q1GTwoXqUC/6AeoXfTTM7SkAoLu4vQ1OrmMS7Dxaixx2kTINtTfvCe
Lb4lutraF6WpnyZFsqbc6/yUXjEgMww/RhoapzLpSFDXtPr8Jb6GkIBsC07e
prQOLcgNuML6diGEY561G7YP5ElOygfU2a+J+2FKj7eio8x2aQIhDY7gbzfF
ocsluNMk2b56lHIBm8oN1aDmh9wBgX9aOTyDH/IO0LmOkWW5UZsjER1EXSP2
1RTe3vDtDZn3aFHLOpw6nIugZdokNp5QW2zoQe10KXijdpYvrrUcWSxc7cPf
qBEV0qjZkTio90XVb8kPxdSDoBHWqiAnILP3E43l8arnQeRdh1izHmW+JZVr
oRUKSeBLrzLMmWux9iEwDNlmVDgBYZTQb5rF2p4ycvtWdo2hN5x2FPyg1hqO
bPMjENaWd2vzqAUO7HaAQPxPS6TmRGjbhNoySlxsyQptihd1rWgo/nhYDKWD
/X2D+LCiJOcK3Q/6hJwkcvoi9tLv/QavOjxqMv+OegzPvdxzar2P7usriays
mMu+6a1X/P4porg+17L+DLXOEv/PMvLwVSnISeAUW/sMB5PVqDxWHXEZQwXu
o39rI/OAc5gGRRooWiHHH35YBYEIjNsZZrBE2JPIeHYNLUBiz44fCM/te7Y5
D5B8No8ebK/k1DyjbLyUrO8ezlvudJvCr6zx0wQ7iBkyv5tQs7HSUWfZp5YW
AldNt/rt5fWar46bav+NKhUDUjOYJsiBzqQ02S50WnYUgyyWdahYrbe9O4uJ
mNkd2gfKZTQxrFfibNoOwhLdr3Hb4fYC2581qvUKXfPsTeuLdSf+AaOUVyrL
6ylOb6INRDXXBRHCXAYUdfeNwMcjnnSm/H59nvF1CLLkS+0cYLXPAidchWs4
l5ImAXKPveUZZkWbhTl5UJ+Jgq73QQvxntFGQuQvo/gqUyMJHLh5HRTS+pOs
gIqg6aA4Oy8c9M36P72t7P8V6vBZB3CEEEVg6co7/oVjSiikiOW381i5uVRI
MVGumkdiGRmyMLHCtHdRTbqTchEBgABpbpU2tbxKa/sls9fxC2s1Mu+nDA2E
S1YzwXU9zQg+K7EJLFMmbhLoiq/+R3f/ewk5mH+SSOUIVTPSoTuo1KrK8q67
CsXf6XO/6SjMzS/4gKXvNd2ynBHOpe6WUDnGuHBoSM6T6OeoViy79Gqle/M4
wDkRCBZ/rtxBTh8Fu+o7hvAh1VOymgxf3FygDXVu54pZ0AU1Cm8D+1XQHata
9y3klp5VlG2cQHI137DVqkxIaHtO5g86ucUlwZw7Y88QBI64r9vWZ4LvTuLU
ZIdEOAqLLP+OGNzLAs32N4H7YOTG8BTzSkLL5H5MHpXKLchSfkmQ17XaakHi
8lmfPSYu9RLa9w0nuqVare8leYNh3dxGXqHP7nopdv8Ua7URFSWVkqA7c36/
NbMFrC9lfBZRV5WB5pqjovqEXcK0U1nnSoJSXNlFwVrKSvGqpRJT7PXCxv6H
+vV6IbuG0/wbCZH2k2teoHpatknMRxUPaJj7i270UCLRahlOAhOZOfVmXtLQ
ACc3+1uercUm5FCVS77BPvBh5XjlzcDaygAgRGnBaKBU7Yx5szv4m6Ju3pwf
eEFrgpvnOQ3fhIhikD3xYYiCUQ0P14pJY8CkOQN2ReKMxynYGhELKJTyIEtG
KsiEZaEOy698uDzNUxL3EFywctrqC6MpbJjYzRIG7LWwvtry8Za3sFCIOuYx
Giuxt1Xy1n1JXtJk9aTBEP9TOynzG6Bm9j25UHbqgIoFmb/YdN9hQFDW3pAQ
DFa2hyf5pOXKJ59hSQZmsHDewt2bUoMRofMdxdweEuWv+pUriVUM8QAiLV2m
+tDofDKcvAsPWe3LL6BI9f4HNclVz3FkIRDFNpPncZup6DJ9a7vFT9s8Py24
2FqyNbjGzonM1NoTZwYgOrt3feD1W4HUSmiTmXMlZ7/h6XAZBFtq9/eaFHvQ
H45VTeBYZMnAhF9N3IbZ7Xjuorbhc44t+2KEOFF9aOmel+DoveKCHnhqILXQ
pkSsI5t4JfiiTZ3BMSA+l7TjYyqM4l5WY7mm4CTqJoI2HAv+C07uPU/4S+aq
eBgCBbhy0jIWFKUSxBG8niwv0l1y80BvHQsCfPZp7hLZBC5aYHHmHWqchFZb
w9oBbek1VqpWfoifj1ULBsgeimJnqu1gs5L4eyAgLoHzGVwY5nzo07zv+l6+
bU7TzF7FwRQzT8xyvMe5Sa/T0SMwPJEU38W0gLL2D0nXz+2+QEqCgO2x+QIc
vNbqexChH3xaLMN5jZznmk1H6z3hPhd4ibdxYTg59ZtCE77u26Ys6D4KwU1Y
4JteKvXCqzMs54kqE+K4Dh5ENp+vJ5w4pIMVnd0rN6uylGlkoLscZX939+G/
EYDoIdHQiOBI+cE3S5iykENfhPGTUNwq/B+iG9jCX6Lz6WnKNlGgM2efuI4W
L6EHoYdE2PmG3if5uSXplMyVr1bVFR/GufJMCnTK/d2t6GlHwDzkDYvklnSx
dNQ6+yXzH57+pQNKcrqwvvPkyePtNBFBxSRquGvzCXesliPqCnL/mP99wiso
U+zCbh8xJZt5H6Fz+C60DJcnCiz/9iSzedA60mTymmQ+/u2NlV6r7hixYFTf
TuFRtOlnqiDnGsB/rKPd76tEM8nD2+ji1o4iZZV6hOh+56DlNG2VMyxrNJVq
lufa019O0DDP67bj2Lw9lYRXhe6v8EwynzgynaYlAkrnhNhOnqrBlv0q5KOk
uKKJqQ/uVW0RuOrZk3O4AzLsYuS7UAk9TVVukQjFkmykdIDTUm4gPyWzqvbx
2KcSH8TBsUCRMCYzlpxrTR2P/RY5Xn1/tIJoMfx7yuPRU70U1E6RGl4lLH5Y
g5jgJDNk1+6MGntPbbnVwEfU3fhr9kWIlQxa2/gShFub1O73B59TJAGDER4Q
rYEDvu0MK+kvxUbQ9Pmls2P5SlHGHi+HSJn/5cByRh7jlymcTXZU+p9Gg/S+
qnQnRyxCqMrLs0pxLrOYV/uaQ/AHkKtGSj0RUC8kC+QV1YkdiXYb/U/7rppx
PMwdkS4KdwqyL5rmENunAIXBy30/Ix136W/QHS4OSLhYHEaQ4ZGZxsUUPIAl
igTO+SQdStaSjDQ4KD1W5lwlh8/ncQw7ZmQK/iAna9lBOJfKFIdafib+2lmh
G20WOAoNKl1hUMjAcpyjFcmSub851Pj445uOx30tBg3tj0YnGkqgZICoWTiW
R8mWxLPQzuEU1yFs2LfMiM2F/wMFFA4aQU8cnZnubxJo5dctnKRT71W92Ffm
c1XgOv80fq+3v4+5E/BNzMb1YJVCgHWR55+lm1chepcyQdDULeipZQtqDc9E
6SCe0U+JQlbho93Wz0bnf9pLNR9yNcqb3m4TxipHBx8wFSMXaYSVgfy/UFg5
Twu8YnhwQ7nuDhB4LZ9trHJ1TAq8SLmjeFWr89zAvX0Ne4Fc2SL/6xdLk9eb
aEg6dL3+5leiriKe4Hoh+Sli0Kxz14YxXSHWVHrZ2DRYS+aT6nDE1k3LIIsL
j4x2BFvmLgepCmtKrYiz4zIZCnTwcGiIjct5o6XLAiQYLYqco3LiJAwiqzsC
gELlenrrJVUvrSLHlb2um/b9vPut7qc3YcJE4nao5i0o5I4pVVIFUZqogZ9p
IHYxZcP5fmZ9LLHq1nYZnI2HnAoMTNSvHR+JvGCUaMxT81ehBn7iUgOltrY4
7ombatGJxm45PK9a4FaqJGHiaf8NtMvHNO0KgRuIv+DSS8uoSveA+OOJQfLS
C0vbslMYk3gDJSR9oItDKva1GwIL+o8zmJN/XbSySYWNwlKLvG30rNUvXXP4
1XR5YuM7YNSqdxiV95FpwVBqRg8i9E+ZqsPgi8VhGwlKpApMW6AXk8P9HrD0
YNRbuX1IR2pnIZu5ozVU4LAw492lWI9NYLKirRelGV7CkpMRc3bJ4yk49SZB
2tEAHT21zy2PtOCuWNBgYPBfzxHTc/I4CpJZd7KkSWwZodSFah1WEVIQ6bXW
iUH0sPs2Rt9ffj/Fv2Xqr/0cKqrbeDJvZHetTjg4R+57GpDin9pKPWjsj9t6
Zzl3VRVrk48LcpJUsik9AUfXcOSbR3/nrvHtFjfFMW6WZQmqDjjVvZxAcFtw
NowEasLRSOiNCqrpF/DsdNigrGz8WghBBdIdQXp65WK67hU9CrzLsU2nmjKq
GiGM65qAAbBng2ZcRtaCD5owBffuF+jNQ2UEsMUpfkB/u0W38H5WvkZ1EDyS
PyA5C9e424BIPDX6GVHPIWehegXoJ8EglRRJvDKGve7+vQ8X1HefEO4K4uvY
OG6bBTYQG5Q9Lpm5oIaIUgrBstts69W4UxHVr8q5bxNe0Dwb5EPbe3h4S6su
+RQfZg/N5TW7/rkw3tIEyGWMoeVcTJXMfJQw4UmesTtPGJXBAcKC8pBpiiN2
Nqt5tMYozyTePrxiK78raLQT5lPYMm/sR+cJs5ZGz73fQS5jvC2Yk/a390Te
MV+xM+RlA43p2AWyDaufQPJeAkU7EmkJqbDtk66nZsRa4lf49SMDDzCK97qS
uRR5s0paBOemSQOc5BL7+p7L+0JeQ/8SIXt1ft8X4TAa2S6PyjJZ4KwAO8oV
G7Yvy2VU1uSR2OQDesbE2BvVDreD50JWk5uvJeKfa/ur7Yrmm/mXHsYu7jpK
FEgLn5/7mq+dSVBpg4KLEa0EKV13nnnDRp3TmdrMxT0nUnytTY4OHXZb5/Jx
W4DJg2YlJ4uYrFFNGOkupVi0OEdjGlazfN++LTZpYN6kKhyx63mdCgmBEECG
GqrLxhZrH8iuKSuvO0jEwk3WY7dIzkP6ykpXSv7/n9Z/9NRuibxvmSYjLXwS
lbigF4GP0ykeYMOX/tkiSYnU5Lut+bp546c0FQz3VQqogfmSj8qfDR4vaIne
hGH+KrLe0vqUPgMV53MAC/FrMH6FgQY5JHZFqVCQzyzN+BjtrFfgjXQfR/vR
NIp5Pt82CtWARr/CSnW5tYtNcSxBk1mtnAZw6epf98o11KPmNtM3Uwx5M++c
KIvRIf7/DsEVYc4dt7kfF6lslDL1NnY+zd23ikyhOtRun9U2i0S4lYnrrKCg
+cRZLBbnaACREUx6oEvDaXu7s4OON7eeQTunpruMeDSofHkZE3bygxUJEi5S
pxewkUJexq/v9uszE3fiN4nkfnhyfw5MC2EbcqR7T+1GO5Raao9QQlTPx3oN
GWdPSWpF/FjPKrPwUdF3PbdabDCFJz9RH2Ga5aRnEUSHDLVxogKLb64UnkKi
NKuvNCOnWHsRqF64FTmp00/J6zKMzCVand/JzBu6N9bH/st+6wDJheXHU90/
jws5SOSKK61h7YhDfZBz31ZzIkrm/TXf4SP3ihy0Jy6eUxYJ1tHMHc/gcxkL
euXSjj4cX3DTlH5ZwRtNP3SmI3c5Uz8HWv4qY8i9T+DPWQ9CZg20wAywSSzL
YbRqZbcMBYCi+nTPU0TyVSO8068RMVC3yEjpYSHZFLRhD92EP1NQTNqgDoEQ
nfCld6R5KvqpmnFzTVH+Ql6xYLXc8rGUJ0RwoNjBZvtuJ5JouShSw0Z7dEJ9
k6vERvdFhmt8JQVkX5W9i0tO16zJYSf0+Ul+uWcoKoeERs/YsZ2BJJdg652u
989/r8wuOYr50QBRtp/n1iZ9RGcsD0/H+JwriOyPnKkgPQzC884bqRM+4s0L
16tw+eLSXMJnxGsH9K/ikP/3/+Ii7xH7rJaJvxE1C9YOyE4i50b+9TcybdPV
HibB3WLIOgBg1Qw05K2PXDWBEoGcRx8oRxFFJICivgouym8c5QJ65MoDLihi
y7l5PcodBC1cDYgQJ9VOfoVAcv7KLtpAE5K5/vcJ6bC+M2TiPfUWjDY49JhV
9+eXyvw/mD52PTLUf+i3LnEw3GFvUEDsTc4ikb4w/A5NFYDKzy0QOK4yxzDm
nucjsfzRz7bxg1m8FqPxjoW7uIwy+d84dVY8gYVZPbqKtQEHNFl53yFhkLaj
dh8DZ2QImXVmAyFjN8/wHrEMBDYSUhK6IgpHDLpZGvKM95mNK/gPOM9AHvSs
nlyRwgMNMuNBv4mh/NFBXwZxtcBRr7e2rB2gS8OQVcT4C9QjQuFKFTn8lCUt
xHZHgvGg3zg7DIegQ7EVzkfNjnlAbUFF+0LubGx5XOIbQp+3GUxbzjywHcQZ
sAayrAGVE3N/HGrcjRSuotGmgI62ce4SLKio6p2bSzE6QXV+7OInFUOT3E2J
p2WrAxf+WfOQJBAUz5QobsdKdfB9EFD/Vc+3CypR4vXXTYJ+WDXlAQTNjfga
J8ikBjmy8Ke6/qIkJ4Rdxo3ui2F88nVpsfuyyiSgHbg0an8BqbmpvLKFZPN6
j6bqjuChLJgYcOiH6VO+90fqcvmgbKoboTgTZPU9M/2fsGJYUROQgfLw3sVB
GY0FxLxygFoD8d/AT9Ld2oX5Rw0Muim+Fvu3K5x2a7UEGCwhzqEomU/emmFb
XyZgWD2yZdrBBmEJM7/lg8+a+NLjCKtoOsUcYmPO+9+Kl6DlY2PZ7gf8F09R
xer3hTIh/MnxYLzRDZ0pTY/NiIFZJZT5zvGahN+kYAF+8s9P4DaccIgxLEkN
eG1TnFFpk3jg20V/6W/Hf7KJ5rSeuF7HxAyp7fzyZ2dpvLNt5FH0X4vVeiIR
CFKnBXEQVqqt6VEOUv7ee8y0lUbiY8TWsC2vPGYkgZEC7kwANEVXD4YItjLX
RtziK9Iija9wJhYm0H9sfp2P/H/xfVMyqsT1Jh1LtnHySy46+p4Yy0mcDhjY
YzPZ+EpsB77CoWAbL/m0STwA8/Sh0iRqwHHbDNI9a5+ae2wP3M0ByxKNZStI
1m3KeMzL2GcChNOf1JtDVSsrPGs9eDeFXq0fZuSzkwKTTVLAGOuv+xQVyTDw
04JLXPl+nQWYVTOwp8/2CKiOjA78hEohbDKVl/LGOdt1KyQhS9+VnaEHMBaI
ZQEVRmGYT304vlVYeWBQj0wl9lx8kbfFmicQEU3gUijhsyDiNdsJO7n+m7+I
q/wVzXctCIAt1bIl07hG8YooqDu5sKCLKlgX5xj+VkPr09GKsrqLV1wBcqjo
M7bT6n3PHDAePze0J2L9RBXnJBnPvnUilePXLhZkp9B4/tlYm3bpllGUfEOF
umO02cGVlrLOspUWkJGjTESqXXTdkbQMjyIeK+FrwgSUVO2PZNdLMuegYZ+x
XH5piPEmdbcCm0hvPGfll+f25TW3efU3nDXwQJm9MuoVcUNwPnmDgsN8jMl2
P6L1B/TpiP/X9Jyi6LsFAm7i/NKX3UiDcIpqcY+J521xIPd4MbC2SuR2T6y1
lsRidNv575Qbo+F7jMs7FfMMa2paP0DUqUJsjnVo8fF4PfdqOPu9ThV/f2OO
UjipuS6/FRy6KJtUblxp0DhNV2P78TOThwdJr2El9Tv40ubb2TCp+gMcK9ys
1tQcNJA9mUBuXTl6cC1n8JHIWFTt4EVnM9z1KtmSsKi7sqr0y8buC5p/Kvps
cNNfn88temuoItZmKpyKMZC8ugOu7v9AOcVbp3CV/ekD/nAXHCYcdEYn0SKu
ecNY5xSb2Gup8DY8/PVfTSPCXoII++cZ3qoIy89gHsuHzQIKdrcpzofIWC9W
GpvtnrtpZLnFTJv6WTFGqAFZbC+Mvyr5gcrAWEgRdKboj6BzxL+kZtJ02+AQ
UeS8GMyDhQQ12aBVEKARDGKPBav+99uv2WAuDq0sviwVW5LETFMD3OvZDC5t
6aTEryh0VVHJCV2HVGQWRWzNI+J+cLolGJ4aVd5bCD+22UY5YZqaSI9tLZKC
50j4wAo9W9vpiPEYu7SbkVsjx94JsH+bhOLK79M6jYfJ/sctBH1WPxPy2sbh
zNxu87OqWtv5N/3Tr7PZnTbX+0PICRnWx56xV8eaRBHZIRLau96ZVMbKa/wp
CN0iswH58bhBfBFkDp2jT3Kx/odiHHC3RCBizKfftNpoMXL7Rm1+Q96OFobI
EwyZZlzBbnk4HcPFx/mE8WicE6J6o5T7ym2LSV7ZPOt0rL8sUMIVotSMqiN9
pcQPCFErGQdTtVw3qTl1nOI3L3YRQcpbUCo4LgNZIPHLqBcqA/HUfp25oLC2
uMcW+PHe8woxelVrsL05L4EGo5EFpJIjLPMaH3DqNNQPCdUTrLLCmx2rzjfm
zjxN+n3jB4rYwQLSWjmKwYiLWZ3hZeXcTZpuqp+gZj5R3amspWKTgiKugH/E
Ublzx0Jn409sBH+ljXVWe9MNlagI/QAuJ44rGwbuQSLfft3y8fjP/2hFAWvt
V5FAbI4X8sK+5gR4QAmTj/El5L+syOPpXymEB3WKYOD6fi5zO+3ih19bi9H5
klhzFOt8ratUBkinZbXfM299/NJDZfQSQWnmqY+3uIT1OLUWloMd7P823Uxs
ITo7h/IinQTdJyg6WsC41kg9sDQ2xcMTlB0laIXyUPr/k0q2widTReCjF79z
LkM0qANaIQDKWTGALRggcLrvmBOApi2foW5TYawvyXFUxqOnVsZk9KXnbHtQ
P/2lmneLLU1fiLc+DaUDYcty2dTRPh+NiAHcasDK9nDKMzCzW8V6Kj9jXDBZ
jnyI+HLaggIRs1RxW0rPzIi4UCcGL38UrSSUeMUGrmlXTr8Q92MioHHjxLI1
/Xo7YAnC+XcJ4YG2+4HnZzH7yF0KHLVI+CfCf+jVTQKwozpvUolCjTMrNM/9
JLH1llhhzahg/NxJNZrKHrk0baPEg1dcmvFYdjOKb0LI1iEqeDc9ngemBbvi
GoZvduAHzoKBZUdRESvEzy9ZFz0+VniqtSeNneaby52I4jXzRxL14MH2ZIT8
PnMdKuy5qiba7ocTTbmtWjj/ObvfHwigTCQlYdi7SmrJajNvpjtt07zcrdmB
TzZ/RD78Y5x9kAzcjexDkI+YPbDT2dsuXDHe1Wk/GquH8wmU24bkLfc9heIh
7Ou7g8iJtAZU25oDlkkZroc33zHrfmBfXCZ7w4IekDXViMUwvjaKlpjzQ0Xu
2FoddbQlmj12g2YPuQN9aTCQM31r11zZjrQYQaRsaxQk7BfsAi90cEUJ9QO3
EaYqmsUBdvvqnlsTbbK87f2KMRQrFV3xSdoQ2EUFjw6QoNlmsZINu7qaVNAj
hPAjJYcDN+OkFl2iaUO2sfbx4h/Ncoqsk9BbP+qecwhglFvcmAg1anc1HVpO
uFY4rEsdkpZjnxrw+QTGNAdSsgPGbGKzDUumR4QoWHAGQRpOe62FILOTJSw/
cILtq8UJUaO/a+OZgq2CFcE2TQUrvmNmJedoibUpIGTwEhccSVje6O9yesZp
ID8QOJbtIbmm2EISOMxLYgcUXfbhnY8Bj34VFz39oLBFy4Y0OMu19dGy0/w8
RSFzcbmqecd0zpwFYm7UMKe0rDjmG7UVhxJOXMklFZILoBlBiVOIqeJCPP9f
QaOsQ8t26vJdJ8ee5YJS+I8SXK3d6t7yyB3Kg55S6L9mrV4Wdg+jSUVvTTii
hFhdzQhcrS8Vn3g3TkRonokaL96DV37BzvKPq1UZx4rVPh4+Y5Onqlzo/IVI
TRF4iP3k0GaCXT/vfNViKdQ68BdIJmMGJ35Ogs9JYWb/+FYey7ufD4p0e/D8
0rdD5x2XKWW19xbHT1xNL9g5fpHomlc7FkyTU8DyRE8AUe7gggp5flBMqOrg
QTBOurbugIbLEdc3nKBR4YjwrNWwsHFl1gwn2sLgHKFqEYoVC+P4gzEpYCKW
s70ajyBFU2JbpYQ/3mjsJqxlrd3Sp4f5PawMasmFzIEB8B+COXAehjJQPiYn
lhoaqw8Gr/cpQei9VNF27keFkoBxv6EuHs+Ak5ymCiNfZGkvseZJIf79hdHS
IWg89ZG0jM0O9Jd1u+WSWxDpQPehEi9t3ISUCUkZwp1+IY/d2VN3moZ/u9hB
UEluK2vI+ui0PtWOwYlCmSNcckdTsB8v2U2B6rADX1cj2rxyvVVXLLOZ0Nr1
MOTW/xKexkdwskoJP/j9FgovxIIPJxHzKrbLkGO0b/XQ+BTCbPyfqrazVyST
wgipTSDsS/EX/BgqtmJXyUff71a/GhTbCW0o1iGVTAcIg2ne3lSFBUR/0s8W
XBxQC2zR0WDe5wS07FHTFX5Q5Qz9iI4MWulGru1sRYdUOplVfnHsvPGnjADg
O20wUkALmGTVuQXxvpofT0bzt/8UOoVOLiZPBaXbv4tLvvxOVjUcigjca8QF
1+bPVp6wEBmvYTlOdFZYru2bdwaxHhxdJp+qsxM+IVpEEnAAqLWjxC2VTIin
6g35IkGdOICd9HTgEHTlEazCXxpjokWd/L28GipSdn4np6RnJwlo58xcBuzs
mOHQ6efubr1NgEuq3alFs2xYB+LDMjvr17J8hitCaGD1TcdVvla+Yl3crcHT
luL68QuFLOaiOUgvSfQDMqe7NCpq8HUsDnzPD+6b/3ET9R5XHsmWogXy48Iz
7U5REYoR6/eSE6v3ldGO2rfKtn41Ue1yjDVwMh7HChrx1qy+hXiy2P497gNA
1qlAoZxrll6vOLZRyXhK1hwxOMq8VrQV0bKcoY26E2Cvz9lrVUGydHfsz9RH
ZQlIabLOIJaAjwuZa/HHOX8fhtXecLvCiXlqE7s254TJ1epxmxrowJbIkZEK
e2mwLggYAxkcZ3rCNe5PF0p+Bjg7+N+D8a18RCleV+ZhNR/krDrARa414463
IicoO0giTPuTuYmAY+KFA835nzuhjDHs5l57hnQLO9ivzaKKYSeNdbQsgJzb
/OPr+vYX4rCqqDXPdIaSH1JJAYXi6FmizJrENELoGQBhjJvnmiWEClPmrxG8
0FjtKFl+1S5lTGQVz1M7uSEP35gKDZVS4gHo7gtl+Mgr4rVYre98M2BdMkQz
D95pt/PU113/yBM6xPXObf4CChQ+YlrsGW80gR5r7TGz80gxpzmWPa47Hw7N
GYCtThqxXwM0vNAo8KNtXsFgowNgsU0o5QlesTnOBkgmU/XPkNKLQnkEd3aM
RLyoOZTW+S+Gb3LAYrH4hMANauY1nPDsoNnuwFvvpXqyZIYFvpeYDJGFj7br
00tw3p9i8AiTP/ulfj66F9vTLKZHoJZM6CXgtQ9gk2ziBm/STlo0YCDXHijq
ADxRbIDSJuFGbhI3KZAn8HmQCZ0Vc6d963xx676yhhWIOPVxmGhgBa8V5LRn
6qHEOwkXyEunDU2RklygTfGl5Xg2HOFdhTJ/kPZ1HyyI0lJaWag2NEeg77Kn
KJJ2oIwPLppB8DRts6ygwoCTsgBTRPJJmF1fXrOh2JZ7emgSItfXkQb/GqOJ
eAdZpqKa4yJxEQWGFSPP1JtztdgDpeCUXXFJlzkv5bdHJvnXkCrj8Aw5B2pF
BwhLz/zuXVFZvSjlMsa46L5ljuMjVWEIY4hgj963P0DuCAEn8jfcoWo6hQ+U
n+ukY7Gu69AHgVRx8ceaezmjL9HogQpqyX3tzVjwU/pdfwIkv9zpQA2qS85P
JizmeiWH2ShTt0FYKz94UEbDXz1ycz7g6oSaYJsA8iJCvRzjsSslGEE2QFri
HLGlpKI0wj2MKE8YT3WDB8cxB51f67DjFfGEBvdiKHQudAuAR+SCgB3174NV
SW7GjLt8KEYw/hSvXWekhoJp06cjTAU95u0+Nk4uoGhD/nu1f0aedq2q/K1Z
rcGnryxy30025wk2AelSOi6Nd9B5PRo9Rp4h/g0pv8fPqnduFkOgohpMI7ey
XCdgumCG60IPJ6qCvwSjBoBlaUrOlmLuQ6dBDZQqm9yJ0uBNYspi2ldkoMW9
aivuaG/p4RMptCK1wKRJO+6lPWJ7vs+cuTY4aIXgAvtyQ5hKQ6BBKMfAH5wQ
OEPB+Lx38fHnbVsPIS0UB0DPKO4XcQXPb580NXPfw4ciiStpvazabTIEO0g0
52x7Bx//zfFZQifzMen3t4tQ/Ti5eDWym3XRoVtZEG4eH/zfscmFcY+8HjpL
sJYn9WMfuZ9x5XS75jVmxQTOFciys0gP/FYn26X5aWGeqTy8e8NvlpiSoc9f
qVTKFRWOk7nI7F42yS0GDg5y1K/S0qzWf71Cpn038ob/RWoQvtupymZ+n1ED
RxubcGEhHeVB5VnRZBeBXkmrFDq8C8xxFrFW59Jd/+frr+cC6ejMqnYVtEYD
PhX5VTnuPFAQcOFI4Nder49kA5Kteu01QhalSdzvZd+8Pc5RvFel9Ilom8k5
cwJs4xgI7EVLh1MZhmlr3vDzkoaFXOpSmBAqtc8s0PGoEPwFIxyC9N3lKX7m
IVRcgegybhOaEpn/ShkvIaX7iDbxTZ6nvtiGXN1sO6BH+PBRWmK8PZ2PzaBr
KoD8bzgYpFYNepo5oAztTcuckAL7cBRgPVDdXQIyo0F33/SiQCyT2C1W/ERl
htmOIS4jJ0g2PmuaDwZ7w/pMVeDgDOoLQHbSs+QMy1PIjOqQ+Tn4KaGma1MX
zlwxV6FXBRJpPZkZSz4bBeoFEwUlZ/+pk6OCvMvRQze2XN8pkp0K8TDTEzEb
uOOsaHtWVKxbYmteSmk2oQX24M+UfWXNoFhQv4gOqAJ685dqclyIJirejAaQ
os49JEfUqHN5DFk47yx1i7pC/ZU76me29pPJalat73WPu2PSkT0PWEhzM1hr
vacBGyRP/NUC+UOZp/RIBKMWzyOdMPd60UC7kz4XXlxAFFjXzPCpKAkWNbJy
uSSDotTViMksmzK4Tvpb7FYD8zeV51OpybmIHYJdQIRONLtIDuv51Ct7xF0/
Y2J24nc+4xoCU1PLAQ8+//m0pFJafgyghacrINGQFIYENUa1CHPDQFmzZIOG
EqOhBKFxY+KJ14fANEGUxKNyL3qJ+XG+77JjRTSU6i+Nkj+AQdfQF+G0IYnK
MdaAt/jP7bkTB1dyCQzaro2jVjZd+vR7KjKfoqOrQHaNYPZZAsk5w4/RNXK7
R8l6s1KxVSiHlPy6bpT4bY2syvxvqqhOmEi4TegaW87n8vynUPvcY2+QI1mQ
cCJnDXLqwbaAfD1ZVrsWaVvv8GamkTGzlDBXS4ch8nwMZHuWYoRbL8tmtyfY
4z+sURaVO6Qr+dpRsGkU9QvHANj5s/fhPZPBndKMIjesxElZplqzAoTsnzWc
GsTSAfYarXuK+eH/Et+ApSAwvugPQnrDJ0tZ4yqQz5NfAJIeNHJ6xg004IR2
c3VxltptEXxUWGs6lGdifshm8bw3ttefMBvChZ1E/9lGceEFWjMeBQecIaxq
KqEH+y1ZqT+G8n+m66qq9bDbdcx+E9F1ZYHgLtVBuTEwTBmxSfCA5bc60ZjZ
dwcIcsofAEU+M2xIIEmv6eilmi0z03Q/fppmiYSYOsN/X1/Yxkd98f4RDA2P
9AsN0hjL0RfSIb2/fqN/prCYo5u9GpfmxliJMHHvegUqrz4td5nbfWIleMXB
AcX4Ej7kE+YrtNh1BlBJTiiuJjwTaamdfZIDx3X4B7pqpo1Yv+ok9kX3qqdj
LEqcFQCg55J7ylg4jnkchydRCnQ1ZHkpYIBEqoVRHGunW1f/8XA1QdO6iS1s
d7Yf4bcKMXJXLFVK8Tw7ymfgodtrbpF6dA8YyYSbxTTcEC00+2hHTnBBNI7y
DjiURSlym3lqmDk/Hewqb/InfDtmdax5AMnTrv5zuGXH2B6gy5peCZ9mrhUK
PDvxdWtYcPOp0i+Q1c8AUs29N1jZm2Gu5Aes9KfHqUmriaT2iCCtX31iBNai
lkFE9L2E65DlEdKZV83LSwAhpnnvS9aePnl4ddA2TTakrL/N5qc3u6McOd/Y
pyKL/OqSKl8T/uvU9Ri9SJoqAGG2TX9ieotYH3elpl2S+2cS0Tcg+/HDvgKS
gYnBfuHvOWm4re2a5O02W2aA8w4b90S0TJAnbx1w3woyWqRXHoaIHMoz1dFr
SPbLjLfFmb2yy+Ii8AFUMBtM8+yVy32iUq11cPw1sMvjhIHjW24rPnWIS95b
iTSir7yG/cQJ3NqwlUxeUqs9eFWtv+mRuyDrbxL5wt0SWbflpT+G1FQxQQ3r
wZeRu3+BOfVapqbiJ/6uaFCGdqjselAYBK1X0sCEbz7ssl4UzitiSDO4ifzw
OsV3lf2IBio3sXRmuZFIWhfehcbFb87h6S9AbO275dJKTOIu2nLlxPDG7ZWj
VUR44BFe43osxrmb3zkbQbA5yTpHqJatDyAyCFKwOH1V6Db9URxZ3YsTxOcb
X1CsIwWp+f4L8wscqB7Y6kNJ02wGAMMmPxrZDkrbEpPUpJF5QYxCJiSjIqH0
CXeCGYBIt7lo3V32p8KSw96nrqdnLKueQhsKfGLKdiUX00YptUkx1Wu77K1/
PmbnCEzE2lpF9DoNoh7WtehxhHOMoyB+OYVySKT8TmiydOVv3SfqOK2hCeUX
Sgh9OD85qQazD5JFRRv537PpRJ2xwop9fKeOu1lotbAumYF5kl2y8LVbX4o6
7b6YCBsZda/On8tYJyAgrT/hTXbd/Rc3ZIn6kqZ79ozXxnLMUns96ngozuWD
yug1tJWQR+GyrZDlRvpFDSQiLffu5kjOz0qwSYtpyZncUdNXVaSYMdOEgOnk
DnV/7ue+ayODWa8DBx9jvTyCqhwZh3y0tdz/XaHLc5QZuCzR/08GTUMSSQxL
gkk7esd0U14x10n8XLBMGyzWpwdLUb6N5mWrwZ8d/EcXxynkYhKU31oouFtj
k9HHxjIseHZ10qI4DH6qFxHzHO1lrXVyCk0C+VlAEfWuFJtxi8I0rabjc0HK
BzJY8siBEkzaCs3tL/Uz/MXH6/KrEAt9u8ErRHbo5IHciIMR60KmIUJJpbAH
3x6i0tv30YmPJ4ifx4IPoycCxuaOb4tbX2VHfeXOhb4bAB9BqcIsfNvQK677
tglZwHjMJvA59Z1I4zWZMFZ1zhYXBubbpfaP1LIA7rbGCvOosMJhhZHOBqBC
xwFIR8X0fyRaU+ybDMfY2jXzeLRhZYyWskTuHxhFsIFGIwFtvbgtKxDXwwiP
f/wUVSz9yEJ1InMYiVJvIkuX8eFYkv4sW3tIAGWvhVxpL+mGk1A8qYYtQmgD
L7JqFtzjCM9l1kKgiJCjN5hw26pOI2gHXtBC3Q0v6KKpvGx3U/EX0rQV+cYc
YvutZkenouAYWdhGr+Dww/3p5V0rInP0Ewt2qve+FZwGa2XWQM34IHuhfzPP
qqvvvNGePWa8rKVsMylmBYyV1Roke2o93rNpUUeI2tOsBT/r4D/JVVwIu3lD
gqjnvo4zJXB+cE+DF4G2gQ4ON2DcOHESDX7CJG+q5baVSx/uA9Dx2IXm7Ib/
O7MoIbJnm0LaIo3RdoFplOgWgGbvDNb0i9YwjYrksqN17JrILib8egf2WrBQ
jUB7xo+XbowbnPOpdE5mklHXKfrhdOf/+j8k7vZuSiKnb8/D+2MPQ5uw7HEf
NmsFzO6GasC7dkPx8sNtUgBRK087LxmmATZEsUpS66iGa+IH3oF2jm/OMuMD
xb6nO0OcFMcHnDWFdXoQsgIbyd56X4EUhVpBbNvnyz1wrcG/kNtonfcoOcKI
w5CqX8aH47zeX/O5iK0kS2s1TI9bEW9c0aEAtwHkwrD0W3rlub/l0nRDcsvZ
PlUcXtDh1wD2ochcJ+tNjtOeziE6+kVm33Ir4IPNkgVt3QbetOPojmSHHsjJ
O232j+gFk1fSKzQi0j4ZC78XJnV6h2HdSQFOZ7q5OdEtnAb3dENR5VlYMk8I
qhdNXsuj1M/nmlkMqVAnjVLBclee86CY1sVPIBet+L9LMJP6Vdu0qeQjrGsd
vEPax+hHgwizBhDgb+XUk8Of9RqqEo4F55gMhWh5H+0EiGPYzxEOLcL1LLkc
6uOcBNqM6svX9t405mwUF55oOdMgp46OaEn00ouAqVQNw+6S9nLYKTnO4EVQ
r3Jg/7VUTHNK64mU0DjYjcsJ4SS/UW5Hhz3Z/fO5ZzH4zh2TZDOvcg0e1qKu
pYnbA5p1Vak8iEXeERgM4ShLkJB5t5RTBMO9k6fntOC+2Dvw1MNi4he+dx7z
0orQ84Yg3am+fDAuGHmSlRqjfl3VonscLnR3FFIQz5ycyrsUKpoDRUUKRz9v
3QYwWuHQBEGH/MKfqZGwYlNUwL8Ub+UMRCe74R6Izgav9sxOGlZ7F9H28RYK
1onJTH74i8z0yYrCWV5XDmwM18c7YPuClM6rZt+iO9UUBr7lHKVpzENdEvhw
ldBqRyaryWLxY1llGYyAcVXY18+IaWJ8wQPjgN+2xnXA1Z2nlwSL4yPHrW2W
kp8ZJAUeoEoZ2XOKYC+FV5BO5xP+fxG2WfpuWjRVpfcamBpn2Mkq0+XmvrIv
zplV16fpaIM28YFoUE1SsgQZeSHCng3Rs1nXe49feiPshbEIsXPPm/0PSz3Y
t9jUexKZ09+m12E/nNqyO1WnTGQuQ5Rmgg850+0D+JZsxweMB0zArzG0QDwl
9czvy2kFYHakg0ks0QJXi6kZutW9PQdeioxzW7HrJhR2+igQRStZPkfU3Msp
ybaztTlDuUp1bC8MeoZC/BKt+EDtNMPIy1B0nmq6pbPXZ9El5DmMiKzQcPGZ
riv4u7/DvEsOZPpsdNiqS/k8W65+kFrzAq5ouW6nG5SFkTK5F98op4rv3Q5k
WYZg8f9+LaAIGUXT5XSvgLEErVvIC8ViuXKq+aPVxeOqdVRocX2AqmFBCRtP
NBV4p68TRu08HPvId8hjfgaXSB99rWPFj85a8BTjooCfwnnRqACw+f/R4C8J
kEUhHG2klsIVLOsO7GedlUFbOmwMIH08FUGkYBH1O7MdJI16CgxJpVvNKnUQ
PU9M1LTb8aw0Rho/22Cr0fsd5DUOZvkVKQLKfF8ONqXGQ5xAFSyMAH1apfua
tmw0hVYv1r3ddzwt5BPrFIuLYSSkINE6nL/kjlEtffN3GTI11UVXanrziP6S
Rc92Wg/cvKL0NR+Y89ORBwB8eR7UaVjsZ+ppVx4nZ9b7qC7xZes18HfW/AJz
YNw90eVguft9qToTn9Yp4kuOZD7qeR9/2VOxwom9H0Bu6h3v/bJPJTPkbV9n
dv4csNPlFHCy1C6sMVu8eh4JsXxQKMOt2UCwZwRgJpCBDQcDRR7Dz72Xt7i4
7HkJkQQfqW7YakjS8tJnYrj2qZ5o7lZyp2R69kxjLO/p4DQRX8fn7A8fmx6G
RNqpkuWEyb/uTDYEmbaakRPtN0eilcYaA4CKl+zlPGMc+gBOMspuTN5aGZhj
swNOk0LKq9NK/F/PcEcy7znQMEq71qFHqqDqtdOR5CZDoigrCYR5F6N6Qt+6
Sl3jpcf5Cfbs4CLF+QteYVtwm9s3mrvOKnXn4REjnR3RCT6ptal0JVwt9Za1
rUBZjodnf2Tm7DU5ZgA8PhPoMZ3q1QuX1Vr9iIYQNxI6n79n2eBbV6FOUY8i
SeLVxGVx84+92N6C1/M9z9nZEu63JLEugXjArpF6diomfn8mFlN9TmY+iGzr
TcmwxjZDzoa296z9QvXIkiRqr+n3ew+3EeLhei/QzG5brnBW1P7n8dVW3BRb
0vNGLv2pFQBlR/f2I86Bvu7FccbE15uX0df5PIVAlGHWcVS1dPlRoNbKyg4c
Y2vzy/5y3AGUIc2xB3GakVTy43HiJc2w3UDGeN6r8Jh2A9KvSIJZW5FYzWWQ
qAlxK8CsTb8kshE99yNQwYhom1D/nIGYXbO7/mNyZ4a9zTM5WgDL0f0XDq9T
xr36l0QwA82Xsel5nUeps95DVxWqgVZWbXY0P7m1lrlsf0DoDipdrscax6aC
VjKlNpjL7e3yjlwqE+GYtaTyFlEADtcJiyHp0lay+DCcD597/p8pZVq3ABoy
Ku+ozobAC4lG3RTEwVmn9S64wZWm8wjB6Nqeaf4PO+qtUrlqxXqTdOHjSwLM
+RK8hNlfIceFu2eNOYxPHuZW1busMzvkrvUb3Yrj9GMQLDdVntnd/ITOjpHg
JIRLFPt0CgwaQPunC1nVYytfHFa/6hTjmzIERBM91va73z+5dkFMOUXMxsEv
U70H3tMs6iHKT7d6E3nLVvOQfXZORDmonx+9Sd+yNNe2a1rjFECwgO5Ajp97
u7OVUJuRiparv4osonzPf1o/pzS96On1I08d6mAtB2FP7ihSlu3KFkPbqMz/
pNJ7e3WrS6NG5PETpxGIYf2L/Ev1xL0kQZuvAcN983Wv7s5iI5f6TNjVvLBn
zHQ1TlovqZ5zmct3o15ZHgSUpR5zaMCziJtmdDGgfdsmP8lVnhIWR91Ikvo2
0hJ380xNBE3wI7MS2RzKdZB9V5rqb/AQ77wtmc1KoZ+YZWU4OnxSxmCprRKh
ranSBf5F8f5S/elOmfPejM1sVDVelasF1zdAIEWxV8Cc3Mw8VgcGY+02QFEh
qOtzmVWKi93huNStPlDCY/JFRPKrKAUv9b97BVwcYgLMiNEQXAMWZ6RLI5oY
asFGP0fevaC0ZtMmzj+1JbOMic/ePy+kjUzCfq0BlMhBWHzOsUS6XTI9VMj+
rG51iqo0fnoVUmZFqbYOAYUy6+egZhtfOwUGbK26RmHr1u5obL6SN8AvfPdx
qnIKjgLfbxNH+rQxspzHupU4QX2v+ynTSCgw0OW1ghONPYmqL9RsmGGTKIBA
wHLHI+hoC+G4XG/STH2Q7E+JEOT8HPJvcUzENv/x7VdlOlAt/7YXKtyFaZl3
V3tQaIGtLH0gJOKarIgGG1MNN/YXQv0QclBIiRQGx/3VSxvF1I2a3FyJxH5h
bvuelhsA3Cgmlvp9OVjiDpqzfusvEynBDLCZPaevDXt+Gis4b8dwbc7/3JpK
t2WRssuhLZCZ/CAzCSPk1LQ3G40WZvNJtEvEx/Bl1BOD1zGi6BFjE7JQgZgz
1e77daAc2aOW270r51l0IkUfdwkCpt3IjmXijP6IxX7rsx4mSquZsOQ5DBmS
PSgT8pp2qVSpjre6t+RM0wTs5SkJYwUwnbb5yESOvv0hKXGpqB4/dIQ/0c24
iEjtyjKPo6Pb3nOYAbr5A3+1xhhSk0MynSxLquWmDhyMUza80wHaodgJC0h9
IGeBfj09Efy92eDrd/1Dx5YbJkR5PFRy7yf+kqm7GghkoHU6nyXWJF1HWVbb
MlOtGUd7p2fNC1Kgacr/gALl7n1vN5B0iOUi+V27Ue6idh9JgJoQGNi+kpOG
HaLh2m2jYd2476hONRctwZu2mveffPXtIH09pp2l7qmWLEafWR3CiSUDAwHR
MtCQAFY6IzxB8bgOS+FRQac/9Smrg8vcL1KCSTAXgFXP7zh6ifll35w/RhSc
frQwLIZH/3XOOqTh8oux3R+aIV7TwrjS9xPDJntTDgEKj2foR+tkUaIl/GtA
oZGAhgqzHY71paatLokP4Tvn/Fh9j3VmBMAyhxVXROeKQ8aMwpFD3b3dFg9B
63m0Tc0dY9yvnblm08pUEB14xS9QnuYyVU1PjaIeOBY0E7bi2D1/mpvUtghk
gpGr1jk/rbBLiT4rNAbd84sk5hSmiIG+QXjWMFS8w2R+phvXyBskGCIcEeD9
X0H8e77gxv1H6Oti2qucZZv100/wXKgyoiJMMkyCcQFvL+vL7gP2zP25TV0F
166Qn5983TrDsn9J4bZNS+6q7EdRQpRB0Lky4PW34oGHxI5Ei3Egjni+zUTy
lk5idMSGGHggecmkPRJfb6KENb92akAevNWDCLQBmSZ5UdCAcf8lmnxNBQ0J
5FMMJurSt+akrVXxWXhFn7j3xGbeDCC4EHArFncZDBYmQS+1GTVQqDNtsuAo
CxMRbbO6vxJaaJixOZNFXEHqvXjpJ7BsBQXb+TNgmBYe5WdjcPhlDx0MAhob
T2W+LDzkGSIkrx/IKevVDFdu0opE0J1CxMon3XfDpYJbfhaIq0V30UPFuUbv
pltK6fECxW/9nTXmGnAjM4sLUTF045yy+M+q4cJ6AlUPElZ3fkhl67ssfI1Z
gGcFqU2HfTadpX1XMYLZhanDFTw/fgXLxeSivuxEVrCW66viGqHKrD5KvHg5
kTaIsDQxFpS4OoVwk71R54T1bt94P78tEOMBGC/B+zGV9mImQCEgExW0t+8F
vMUmwj+HrZ/U0XWap7d/SgI/L7O40fzlOV0bGStN+wduI3KwdgvC7qV9DbBp
iqYfqM7cLE5NQGj8qJ8c1eRYXU3ZS7xo6k/BP/whjRVnZMz7r6FBh/gGyKlN
yYQjd3/Hu9tr1pFhLg2Ibhan0yU4ujtVP3lW+wnU/ilstHIMwzRdAYaP082Y
Bk3hyCU5ApowEDiU+M3+G/79RtBoUt/QJRkNdHhUpfMCLxwQUUIpvoZFEE+8
MtRBv7HcKdOsJ4PMt6z3Sein4Sg+PtcNaNpXvn0nXjKP9fwnoR2YpVOP0Ejo
4NCipSg5J5Twr3eShcmYtjIWX71neXrtNaFBAILOZnUbTZz+ADG351s4mjoq
QGOs/LjkpL2J0GoFjaOl5ucTIBhBp458aOVhdtSn2rG8Tay5fSV0znAl2b0N
/OMvM9COg1IOUx+RWtkZ0rndCWGSk6Le23+EPbJXQ6WF+WSACrxz1h8PLRWU
V+lmmJQ526QOZ66Q48b/unadWwXfqLpxAy/hN5V8iULaZQbEuVHwe22v2GZG
k89XGUxu9Vvk9RXw4/b/fSkKPjNBeFpiu+2FhKtUkT5xgrZV74D0HoYQQOlw
WbZn9UJE1uwphaLelQ+4Il+bfgLtxhMT6WY+YtLmAuHCY4p2epdjAScPPDr3
I1CmFAC1CtWywPnCz04Q0d7iLqU25yrc+2kC1SMZfnWaEsQhAKjh+Ot1RWZh
Grun7CHQkzgr8OsCXr02CldPW9Njrw02hQRwvaNPwo9+7Ki6lPPwnPyHP3Qj
olkPg7owHhw4lPm9FjnzTh2LunHKlKqK+wxsuQwjzm9Bpji6Oobtv9ieMxky
52MLoCFlLSSCm0z139f8QowIgpDdXrte3a/o8vShvIn6OOTPP6xs2+QvckiC
AqifdZmPMrjkfbt617+KMIUPw5I5+cdbwxngKg9nfu4Om/f7XPfJm805848f
3x2v9ww1luR9p2lVIk97SPJBX2R0xwQrZ4acOQkKKbZOADcji5E1TbstO+Mh
i8nQ2i8/ak3s1++XHvdGr7rG1Y716/uxTeEA2G37bfOiL/fZRQoZGejGdkrV
iCyGSm9G3xYdRqX4YKZlJnsSoJnGAq2mKdM2QVbSTVRnI4Ch2pUygKBYN7Ei
anQV30lzcgXt9au+Dub3fdbtkGZgBR1p5pEIfGZ63yYZvRdW/PSomRZuTtkW
pcDftNHMwurx/rFqY6g005gEE5HqEy0dB1OZGOKPDTizDCMHhBh1e6cmiZow
YpdzYDe1C21h6ortpN4kWlSaquZHCEHTZBqZ0WiG4+jCalphTcKaK1BN4G5t
s3VM4O0wFX97RZtloqSZussm1bwQPQHxqLqIfs12f9puySfNwYFwK36GV9wZ
aG5HIBYEwDc+/0PjElQe0N09tf/chRe6paQis1eOG8LMkiPOSj2NPgcogfqA
PtUftP5OYhiOTghY2uCQCVQUaOMQ3xddx1oknkq9tlXpto+Gag+KMerVAyo2
MCpjYAYkMF6L6LSzQdV8gktdPzgir19F28Xwlk9/HkWoS5SRy59nwFqNdrL+
ehZ8xxud7KveSs0w2P6XUkhmVtE0ZGi76KLBS0yvjTXDUFCq9lleoeUt9KAp
1cgxyetJn1zB7lfvJxTBUOf8SkTz3Wf2g6k3+kMPzZ8AZdZZABFctzOD5SRr
FSNj+ikEh47UUZFn5uQeNk6+ICwcuYHCKrawHFZ+xjKV3+i3yx/D/vlCZVGI
VfYSVRiG3U8Q9qEYTAuKFgZpd4KAqGWy0ikolo+zf0QKlHRb9Lr+FllaWEVz
84bWOPncQjIKygfifYun7h/m/b9T0KfmtuyxzAwv+ldTZC1vxM4fY9NLCk4P
fYx2VBb18OdEmFwmvSWRnin+LfEgMqatImBcRu8gXIgK68Ka0tulxurO5u41
0v8KCpaJWUIcLhcY7gkmjyR0skFf6u1cVW/9Q2AJpDr6F5oMZfpA7Zsbvea9
vJiUIu73uObV/uIIAm9/PYZsH+20lB5nL7qUo8law1tP5k4f3vl3WCAih0o/
vgauqeMr4psSfYTKPUGqS8gdwwA9qAb662DWaidbuIYkEiNNBpyxoBy7ER28
7raB9iekHlH2+2dSGQIk1z0p9ZB67/y56KaFWw6evybDr+67wGqOhE2B0/D8
/JEHY2rXvfxkC4Ect3LQCd7T05HBj+5bYAuzb1oT2swbJX4VGhYeYnYd58LZ
u7dNLI4QMx4LfyxAy3OD+Ld3FM68MGHPz27E153kZ01MXErFNCR6Iy+yrN6R
z1pDA/vYU1E7pjYjZ7uJy0n4IqxcLtHwnzxNrKKHqRLaK4srK3J6fwhRaltN
syFERTDpW3p08PQE9laXyhhP/cduDkpt6WqVO05qgp560G4LdGoN59bAmfoP
kPX2AkIPm+zRoMF2B5Hs0MqdFXGlUS0mSI3qZmEOv2O7DsTebGnfMWvr9/ch
arAL4FMIP40URSrm2t9kuBGy4iUOIuAyTCo0cQ28Q8UwTZETAGmcYGe6fMsf
bf11UBLirVaiO3PPneM++w1XD4SbtSZLN3QWnOV6mvmMHxbLoSDrzJEqT/DV
Eb+ltGwAHtVlwd2krQBO1jZoczpXFACTn3/TBZ1qQvueZNQywg7/3x22GzW4
ZYnctff8fSiCx5f7zAwquzjkwi8YeA8KH/erKwELcwuth5gGS+QJW93ajGx0
PCzYEgFvpwES2eEZw65JP56eypaPRe+ADuKWdXLd75oKTBrDBDW0FqT8oHCn
3mNXcrUpHkJbkk2lISYfcPNm0vBiTp4X3PH+GA90RP+2UVh4WG7gs9CayV6N
ItMY1UdE6IlIMTsD5f+oFQre37t5FkUJFMI5GTzADJ3Smn7ha+Zzy1dVV36g
9Nf7CdEyVdVQyLfO+z9O1J4H+4PrODWs7CZ2oQ7FOAGbsZCXFNKA2I3gHSer
AWNEH++k0vB21TsQ+1LSmIZIPzA41uxkJE/+w/iQhtasSe5rNwz/mlIYjkrr
IUVYOGoLVXw6KBLUgOAiceWdO4Dk94t89M2bna5yi8JkQ3Jx9CRo/2k1k9J1
Vpl+xG1KriDosyGt7ALDCcGmQfMnMoEBn9AwJgotUBX5PuKzs3wQjBwTptZb
hILe6hYg8XgZ+slDkB0F0ljUka0xe4gfEcyB7uNyzOeMjx3AVVLKNHYY3DtJ
MH9rxXLNvxTxZCj5f3WsR5V7FrSCKn7MMyjiflcXwA3XVTRx1PqrNckiDxsX
hvivAAOZ1GO8tXiw0jqa97ozw9796lhTLKU9/GTlXaOM4yyC1pGpqiyttw9Z
o2VufspdyvME+4vOIAUw4BpLqSSNrT5Z2MHzYJa1j5HoaeJlblx+9Gi5EmSj
4dOobZl9nOqaFcgbdMQF565gNVsZpNzvcU9J8CU55HFpYk1AovApT4xntNJd
k7c1OBUDJQ7cNmMFxD35bym6Bm6vFtLi3XrmPH6bXBPPntvBvxWSYVU3pu7U
RZsnNaA/MQ1OQNZjwInXTbRvyk+kiDj1ddXpBiQ3vG8f5jMBt/P5T5UUURKq
JHgP8+xLuCLaUFT1e6SxKS/qAYbvB5Du58EnMC8/DF7mlloTu34KFHhNOwt2
2l9mHVv0UzArmcWr7bPqYwsL9Ca+HtFc5xII/nCSmlEcGVEACFpjz7h5zjFt
KjXpm9ff8FxjF3wHwsK2ZnJZ7adVRSNKOlfhHwnDIa+HxQbWr+yrEsmSd4Z3
ONSsaq+mKRz5ipzFS1iPLF8z7FqfjGl+4KEGS+TFHkzTVic7ydobULK0UdgA
uHFnBZCy1HXjqD+9RoVOP7p73i17fDFroYEreFyE1jXyiSkYU5SR6zkLZIPC
NxVauvtpEQWV/gEJAcAeH9azbSsRQJiAnh/kDdbQES7jUpYtOk1synNAGcYe
tJTZBJjlTDh6wseCoXsTp3eLaAceiDdOVJ0TndnnXf8lAdpnQj43zIYZ5rtA
pop9u11QkEVODfPudrkeeqNd+p3OZ1DBco0Yf0tMo95BR/MswbKXZnBgInGG
evY9s+Iw4NQF4qTSbNupnyJo+V+faYfTCgYreoVe+FOKw5BpBCw5mLJuLStK
Eml3ZmgouuS4A79syFa9Tdt0b+ti9fz175E8r4zumTc5ZrnKyzn0FD9K5ZCv
3JwtCxPHxNyb1xc3qxuXfptarAmQd1G0W7l4/C+N5u0WgOjM9C9+MpB8tiLO
orrhAqFmkx+rGYzkUcD2Mv3emPWYRntKBJ/gpt/5u7ZkLljixADGS+DK62QY
7XXzQZM9slYgLS4s5mD6vs16REG9tsA/AvJQ0ZgxXlJy5vAkf5Cqek8ufvtE
8+HdFAin+Hyw7LRUXjxD22/vQk1yQN1VShDX2nYTkpSSQaB5xgV/Fk3m4wjM
9qkRk5+CU5LcvI8t9X7+c5Z35wjr0HoqP4XdT0KWvGFcujapECSDPt/wUkdW
t4hujAYXyldc/Oc6N888RD/vn0+SVcoxLW/qjU7krU7K3T+Uy4ZHMwOMutmI
XK69+GTUFNdKcJO8IXOZQAfyJIxaWasGiUVqS1q/sG92jUVAcZheyl1oBsHe
JFXuM6T67CrA6YdkC+/Cy0mP5u31bOF0FoDC1Xx4Rh0WSm5WbqT9uKVlqU/V
1Nyc3yWEEW8veRIB7WaXD/xtxhx01JPWREvnLd3wlKERi87RZ/yyMiMqhYGs
MhGb7Dooaz0KNriJ867L47ioKH9iCv+fS6GaOKoN7sFW+hWg/8LqUuoMv/1n
5kSXZOAX+jg967KnDEX+hPCIch4DviQ065W9Vh/Oo/nOSK9wrmfwQCTo8vsn
3o8ZlHTyCP9kP3lltL2OeWcQipyBQevWQGBm6a/zlxEMVSVpVKi0V7GM12UA
9mrI+rr86wiQOZwQffQo75bDqIilVwVmotQmrP5LyRlLVmFO0Hid+ZVAnQTc
3GOs8D1vo6BEYsOSbU3VP9RIthJ4M241201kk6HAVWlxCwZlrTzgBEu7k+J/
t7miiCv6v3nZUbEMAoPb+EoZT1w7fU9D6mQxAuP6wB7Bb/EVeLI/B4WtBN9n
g7HJFwcU77JA8rTy8gUgMIlbI5BB+0TKEKZZLlHUXqaZExqtZRxBm/xJSPMe
0pyegXSgldNmYYlzqLmciET+DT0MB2gn51atY8Wfvg2Xef23un3jKUnB5Ryh
OAh+QT9/QY04kMzoUnWLwzunFuyOnOed6HegvpOb29lpmQbdQh0KhgGuZGM4
9kWg3QeTsMYlwkKa2Ux7R9cZeAiBtjHxXcArX8smDJIuHyBGIzcyNWGaxuyB
X9PZv/HtKoLYCxvO/7Mx84jy4p9ugOMmoTK956haromRmZhQYVxCx0DHaMPy
mg4ijvXNgremuSGeimw7x55gCrw++MUwj/A3f3C/iqyTJWEoxZf2d0uYghag
RaXtCQIXI0AKDezYQKeKNLt3yh7A2QSgFJRSRsqW8Md9eIM288SRx6l+nLiN
YtMqpGMu3I7aUA9YuPfLG8xGOE0UVvtsIB+aTqmQpjB2a1YRfvG3Xd0pcvdp
ElSwhTHvbGlmA3bIUY49+32bOxcsxFdLmywRKPGRwEAJsPFTRkLjUHHUX+0b
Cwk+7InDLrqnDHqLLTOeYwEHwES34JKQzpkruFV+XA7eNtFwNU0+07uhU6tU
WL16HdehnlMGmiprbtuQcB1YP7jLl0P/hm9e38wvMNVVKpCoOpXFYA02+O52
gU8yFz2o/JyfcbnD/CseONJuXkQJVftx1wFypCixFOMR4ijqPGlKbutdeK0X
nvGurzqpXTJbZZc5d+mSry0FDU0eliQAODf7b9gOX6hZm2M8FjWNrx29P3t2
rDA42EFxAi/4tSZn6IEH2awHl36yAD6noeYRwVjg8kYtZ6XBsoAnHTjIru56
1l/yjHwBQnFuWOZR8/63pbBJNHKbqcVBiCdxTRBurrBG+3jDpSkKCrsiNG81
BagMgrcxPdINcFkQ8xFDXjmmU4qD0evAtptEzri2t4JMqlhA4yHWDCpNspnV
zNc335MIlRyaPsNw/aJBIakwkTHOliqc50+c7hlBOy0pvOGb/ZzMTFDnJimg
A8nBPklYU5QqzBieuN2qd4VUZDDzePc8HVlC4XaLzABnvsLElDnFUvI96shE
IXGw3lsJN1mnZuHUEGm50c0nfJfdMvOrBvro79NsaKW/o9wnoveZeGbDmhGu
VyLk+C1BU+V8wYDz1h5fxxMtVUzCZbq3HYdJFnTtkFtMMpS7EvLzPzhJ5qCi
cRLWCuDhxoR3HVc44UTH46zRVU7KFXYcburEKEkq10uNK9saPoC/Go4A05/0
QJiXrmQCeKddqNB6jzz80vd81Pt5PyIMqDR3szCvBy2BKBn5Mwk+kkkGEBIX
XvPA/7RWaLIno3smCWmQbosMj4FXwXKEf6+1IbxE2O1HDBM4bh8F/R8H2U+f
Lc/Db5Sgvxk+6+O17QEYlfNC9t5/+TMjUZiDhNMbMu+CrMCX7Ym4tkJh6E3e
51bW5dCw0wJADxmnRfym0PksiGdyySkZxd7+fD5+fjbvm46OowzCTHkRz+fw
Fq4Rhljl1S6rd0eBIllpmrntWjfThVrGaiPjO1QDTjn/9JrwuzBxe7iQUIoe
KPTqbEGNGQ9Nvzn3stJMZ4JZCRLytan8FGpl+6US3xZzOXc+4aYeLGGipMQW
GMJjDumLSwSs1A/qU32uxbzEBolLwcL3eEdnMbEUFmeh70lJZsOvcboXR2B6
QrNNQ28EZIy0t8u+VSVbTmAEUA/x5SZuafVbreoMgJaO6/19jb1qXhPWbxRU
fa05JJ8bLl06IXlxHxKmx8gpB6bQSKlXBM69JIQWfnFWd8Tv2IjSqSC2DQjb
Lt1mYJ2Z0OmPLXUKChCB1AU06zKjzlt/6Nuitldn+Q/0zn0ZuxwPGV27efPS
jm2OdBpiDReKpslDCnXEIZHV8l4iSCOORiyjBQ7zZQQEs7mZXFnHHl3FQPK4
eZbb7s6WH2CeluNeWNKrj6oryunjiEAepGjL5EL8H3UHQ2y4VktUswpMKW2X
GFN+SAtAeify6r5zYa7OWp/spYAus/8Ll6S2mxc333IZJWxMLfMLyLXMXQ8S
TL+w2Nz26m71tF/kYQqdOJR8xFOcTHLvOd7SwopF5pszcZtkCViJ1k+20KgY
UHZEBhsePPItyPWUUldzirymepMV3sxWOGZZueON0ZiFksI9KO7H7v7hAsoi
pYN2t4Q4mu1Go+x6xI5fFwvB5Ytl0srpPjCMiaQXpi4L9nfoT3cBj0J9YiUc
eS/6wPDBs0d0OkkdIeKZ5Of9bygyXnAhNBCIpT9fGZG16KUg8aETJUOopJrv
/UdkPGUmPgD6hDmAiRdFG5wOjw6j4BIV9asFkyV3ObxOG1BBYRhZ0rDReSX5
TZN2Iut8ibtmJFRNr8K6FVpixWddPGITlW61dLbJVgcd3tGZ6JDwUl+oH6CD
pkiy9etzgUdzOUiB7szubBx37ToeFZ262kG9mGxnSmDyPBTaPC5d2Zas2eYG
L/2qN/X6/NtMxEYhP50/TmxMgrqRleqNfhsCBzJXW7ps+nk/+3sP7iUf1CCb
0rdVvzpf3jXRDQ8525AWdcF4aGQFtsODekv1c3Z2iKLata2SPqJI2RPdR9at
PBXXuYvounsiPLFJOiutnRmEDuQVlpXDd/XC+dGptLZuHumzdg0ibjPgRF+G
NgOFpbMJV3BnDuv/eGQZNG4f42FFFN0tkJR4+6HKlg+gVPNnUWaCv73YPjyK
NdR542PL5/HvI7i6R+ZQL8kPd6qVIwTEobDbcAA3peSHXU5gmjuyDmTVneJO
bVd3DGuRyMH86Z5dU/lEu2+fZ0eQ0T36jRJQ4DOxmrj07EE0mO3pWRbrtbm0
w60EL2HisDboTd/GjCvNFFa1KPBisl/ry7JNob9dKV1md2T+Zv9hl+DkKsjz
VA5h8YZXx2327vH+Bp4VAHaAD8jpQKZvQBZhCP5bSNFvtLB/m71E8QeoddDK
AK/gjYeQwa41YFpkSviZ5BGWGgd/7qabMLkhOMhS2TmLct/lWXeI/2wa9D6G
xjtVKpBPh7DRa6r7bii8GV6NjpvOwha/PIsHZceNCL46bfQdXqUDqBng3Y7M
7nvkxyfGL8WeKOXhqaJvrLedepHjJXkQfRTMSQIe7+c3lyuY30UJyWL2mGiP
Uc0bojgXDTIOC+sDgp+KriDl5Rro8Rtf7Mt1Zz7Iosk7JhmEj9wloPDbskOy
KwDqP5aX9GGzhI8kCmh1qFGu3V0M2wMCsfismT/BLeyYg8MpH7KhsObOp43J
yQMGyH9YZ4Y+Sy388iDDt06qJX9oLk9Sq3QW4n8lwVV7VUpo68sEe6kYRxdN
01YoZB6XRCr+YmJ+RPsDOi/KDCXbHrqkJA2NmttToXQOk1Jkfd9z6XD5ATUu
iLyct0asz+b7qDMH8K5owN+THaJVRSH3yI9+lI3PjGicK1un3nRdcWuESslN
DCLreIfFW2ihvCLVx3zG7PU7S20NaoutiEKy4ErCvl5KhWs/ZHODCpICjb+0
3wAvbnzcepThsCr5L418G8FSMVdWOPg7CR2M/m6aIz/Ug9Su/8Y0s2OLJ3zY
Sr7pvCxf/oKFY0SU+KDlJtTnEtXDk+2DE59wsRcBolr8KfHl5xYSoOdDBRjQ
q0YgzJR+QsWdapPKp513oL20BaZ7W36CENLN24KkbT3rQYAHaWOqSQeDcRFb
gcO9xdsMdYD0HgMSqcVJ3cIcYH3DQPYr8NhB2qdLpX4obnuikT1XTymcb2Cc
Juf2nPoZWx9i8XOWhHoLLAk2hzuni+JdNLtscscCLniSSqIbKXyhIcxNYQhv
lcpY9BSZjSFa/0Pug2zXV7GHw7W65wY4jHLVE4eS5ES7R5TXAA0Orl2D8KUb
U7Cfwc39GaE1I5cs2kajMrZLK8Scdg2fut7P3RQDNbfs7hMJWMRK3ZTuVUmS
LdFmwpHIYE09YnekzikwLbh1SqPaycrr1CWPW9i1Rq/VPC1p+FdCDprvk9UY
isjXaz4E0cg8vxKXod3/NUQANEpznJhvsMIu7TQyPsnCkQ0W8pNBgj6BUpIX
0/1VKwB/vn10WhUcZN0KUzSbTv2oMiKBPYBr/OqjtysUdMshgemu3kYqeabd
QqGps7tpwhqi6Mf7VOZe6YlDg0pHog7pGEBDv1daputqHK19fyTQqdX8m43p
Q4mth/jFDPLiDEfRWifRs8gnV9zK79U3NYLlTuOizUyDTxs33e5YXDjakcnJ
jPcZBl5XiKh6I3F84AQfgIIje0LUrP0zTccq1WkMUyjJfIRd3s960q9YsdK/
QAPJ2ivdjohrxlf8NH50EPZpwewvhMTRcZV3tECOLtl5OKYor0aQD+JypGrb
JsaHjxgmF980frCmnAb3XwrzxvFjtr787vn9WdY10xS0rHxgxoO6A8dDOQnM
As6HlDsep4ykZFvFa0woMBsWNjLX8jZk59lOLKzhJzVMef705HH5d8p4ej7c
qdgieTPPOsH+p6L543Jgqo83Dhku1hbM3qOQSNyuJ2Z99/HlG0SPUIZTKlQs
cKm1DB+cdhXq1JWOGzv3FUxJAsFMN1NE/X8BAukgDqeJA1rJ6G+azReSvXlc
9NHNh5Ud/G4aEKW+X4G0XVoOrdj86+cA9Z29FILtjoFGUHsEgDmPZVM23CEK
fT90PwAp8E9sRO1zmcJjYTQQG3vYQ0fmngPK5/zqsi+o9EuD81vce9ZvPToB
yYwuVNlNGPkz5Fp/qfEoK/MIaWj8cj9M6SOD3ZRst2WBEJQmMehDF1dAvT8A
pLclWKG3USna3gDVlBoc38YJfxKIv3OUG3GxpM8CHnM7ZS+feR+vgmgIkRiS
x5Xa0FnQmpfrXO4/tzbYdDurysBOJbfSys59Ra31xYsPH9FK0qz7ss1zebxR
otFejJsB0P73qqzwQjEyjVaYJB5VuVWEt7Gg+6ofCkVYLwJcaOA9U5ZCPGFx
b3oKGxRMQDmy82f512Vnt68aqJdxxm20PB7kVTlmR97tBoOx17jH6Zbjj6Qq
QmUgYWAPhiYrAd0a8Zgfq8H46Nfj6tjxPkuSWfN32UIgfXQs3SpzQVlf0xuv
uT2tVlVCAFqD5nfhsBftNObrijEIugR9ZuwY11zGLbmcKJ2RQfe7u2iaYmRr
Q3Oad8YwQVuXqMa59knvrxuoLyMdL1PWEQq3GTs0spknrr4Mp5EbW8uM+lyZ
Uc1rlDKfyoIO5PP+700HeYh0asH1+FbP3GV6yLsswhZeX9olSzjQE3UmzrvV
kTE3TAGewVoMhnIBQebwHLsdLccNd6grE1h8dHnBmUDZZ4i6li7y5ms/vyuo
/HMI2DD7qhqa4uYUUVGNMv6PLJYQB6J0jA70Z2tRIvMDuehWBbAwcEZAysPY
V8o9cXqPa4ee9USnyr8+t47TiO56bCY6D9x5WapLzQs/TJQldJzb2YZDSLMp
/ZdOyvzDzD4y7YXO16SGvZj+id/fGHCyreOri2Wok0xDoA9SKhsMST/e683H
cJDnIIvqeTpoeSxZZQuxBmtITGAzL8Aej/cHzIRP/mhx+8MQGUikTC8rb6j7
UHTRrqeQih47nRGqfzoZT5W8TR3LAIZJ7Rx/1M8XiQJSPs8ZdyCVk+ks5Qpa
A2iOOVms3SzgOiut/Jes0FZiZsnCNE4/6TQL9V+1lo4jhGZ9U97L65yxs7Gb
JlwKP86jvapM/ra7MuGnGomwx8ca24lUcO4qcbhsY13RDuJiYD2txeg6bsWF
i6V9O9KkJxXh9vNwYTSifAlL0UK9H4LReCLRnsDuHJMOhbrbrMOZdqfFaAXr
6BNs8x3ohYymYDWUgI4qMATRIEEKFddOTeDEJsU3GPSrnFze4KbYU/FQXTbw
Sgo4BzYFsiGlv8F4wr5WxKsKNuzD8g7b3Te+VT45xOJoK/Whd5DE1wQcNqX/
b9jDW/gLufvX8TNtTLth9/GzCDof4sfOiQimY5Nk1ayoo44o8fhW9iIXVDpV
K6IWwPutz8LoxNxcp6vJ59HWXJGHmgKU5uMzU99Vn371yYS9fDlhCbd0K/9Y
a/YLBpwwjSzdbt5NQ2fQTzps7HrEn29hT7dAfY5bFLXbx7rSMZUUJCzqJSaS
C+3/JSb72gPuY1e1OvRn4V1vRaAXv4fwHgyyLY40vHuKmBqAUHxqyR6ICeAk
y1wR8YPr2Y16pL4abe6Q8yiPtFCcywOkaUfseTw4LjdcXT6jEz7IMqMWvwJd
mqkOgPzgATcxD1RdxUaIhnN/3MYAFKIKvZhwAd8ut29RNZoo1lr/8cGGrbtW
7PhlbLU1V9FHTGh5it2I528X7qKe3LMTa30TWvdqMfD9FT4K84YHjqtOSn9B
9jTY1p7U4ThwJ56zGAIGwUfzcD56rhAKZk7h37yRlpHTNOYpT3+B7+rQVDow
WG5VO1ZGoh3iKPN0MPQE3kZcci809x57UYdWg+XWtj+ZP98nWagq5QWentBK
uOXQyRKVzHbPdJkEaPb9fjtBa8HBNJXgwnwdyzrBdWcWfbII9PQltwOuhup5
b5/YgVb8KUFhF/zPpugt4p1FaTNOPcjStCyMSATFyDHYZxF9wc4gguq9fDJ+
a0TXC3/Ag72bvgfBBPXMauMdMf1PbxKl2B1YJld5tDYTlmQM0FCBTLfbF1GM
QPqAHXE77tKY7sFMbL2ZK1odz9MLNB9/cGixh95lNHdnUt8bKQgD0PSFqocn
HZ+HRcjZUdXHs3dvrf2Ga+z3afdmwpe49ut7poXyJo8QvJJLR+MLCGMPQcz0
zjJwjy0C+LJ90/Ohpm1qNmho02CbmlF9CNmpNjUIQ6HvCxl6OKh8Eg5nUfVc
obKnrimncPv6+ixzBRdyGG0Q8mjZ6CU51iFxLqUWUCPTtdMtIW4q/IaEkB3U
CjnchG2gIWCeA0Bbgo6Yidsii8R7Pfx82rw4z4NQwPMuUaHuwiVXQ3cYbGC7
+HdUrXACljMaIS6QhRS8aVKRzjVT7va4SX7cQ3i66Q82231lwyblqnW4BIu9
GPvJjNi0NOlupUllk0+asukJW3wi7WGvexTtA66mCFVeBClQulqHQ+gFTHRi
x2aXJFkU0L0hhVuGSiT6JNM25YIzPRtaMPj/h1v79dHjQQAQPCrTNN443xji
0ywM5OVdlnLqZQbFg9fnacdxKCjcD59o51pAflrBO+Odb9lLO5fACdOyLBNr
Kk8qySahy3B5e5o0zt17uem1yiH/qq1EzoldaDgw6ONBSjL/7e2YSAkRQGPe
2wPx1/4Qj2T+JXc4EPxifyECK5IeMr2XCyLGhVCmJpXSD19ECNri663fuENu
Qz5/rDx1JX/Crw9B+V5agEuaJ/z55/ax5MnDEaBoqSyGVU6alcQB2+DC3c/K
ooJunISuWokEHymiKvCi6lNwntjbxB0Dr7VMkoFHYlfu/KcUex0aSW3d5MoJ
slvMy/sVvCnq9KQ83SL/IOT+qTk+5I1Ubi9QqW6aiuSLDypppaEbsUbKfJ7f
V8r8nZzXgncYIGI1Mg5bIXpF62OfwrGUW/SJ4V4+QCKLh8/DsDTp0GiELbr6
rTPQxq1rvQS0g3G8RRct9h+wJ8TC1qW+Z06IC6iI7svIqiKVfp2Q6y4MWCoE
RDdjn+EyOQ8mt8vfNFvoqi7MkFMfA6UASzFmJuzb8lgxvR9czYvQbbahiC7l
EFuQ5Y6RxtRLL//tolACtForKfH2Tva6JZrHqOHYgzBN5zPVfuPPGoKfqIJW
9C8SlPumd6mxkeGugVtHRRQ6ekNVUIMKINNZsMBb1NE5OVv7/uklgpDgqM+M
FHlEUwhsztnInCYYy5nhFDRTO09pN9B2wLXxwltJb8t22tlgqTdhdBtntCit
uIdKsQs+IDV7bNj5n7JwfyM4gVcPn9U/D7K/X8xJ1ybgN34D23dRpamlptjZ
J76h9FEwql9vXOr36rZtts2RA+88Khmapu9QWn5BcVbWL856FCwVRU8EOdbn
ZdP40wjCg2/BvLLlAyeAR7hUnLJWpH8tFIKjN516J59B+gQMmJe7t1SU440H
zvSNuC5EP3MLkpUuit7WBYhDZZHWN2cYDSgT/FvPLqjm/6OW9kObJK1mWk2S
BwRtgwcc8ty3aet/dc8x1LrNnA78gUOFcyj43lLXr6ud2Ha94X50I0u3NbHS
dH7SWILzzwbqnhLKn8i8asf50t0+pM8AHuiORQnQRv+giqWQb0X0qjbtWU2M
yQh6Wzj9wIsaC6BHR1ILiNs0m1K9KxH1FRlIY8DI9wqsxylMyiyl3KlbtiEI
olVseLBa0EHgUVBlZBBzvD/63P0xoUEYuzo/zlwJ73Yn2t8sOBI+rCbvqLGE
k5Ba60jq2gozyAGazoWmJXfqO2/5YxH+2DjSE7eD9geFxFPws3x4LOR3+iCl
lrIXqeyTO1bPNvDXs4XTGD5MPiIaVdQWwOfPmkvAHFxaER0ki2+QrwSFcJ+U
oE8PL+p0jHFKzAwfbUTRUixUdEc489KNDjTPCuqMQ4qJAD/jgWpQfvaw6YVM
32CMAdQlK65Wdani52GDCunQcCkyUsbQXhHm+lGrmJtmW0AIbyhr3HaEn/YE
WWHdzuqKU4kFvyMYcdhwPWnO5KtxJQwlLjs8dSyMsQBf1FdV5J0hMIBAsQeQ
d41ZFgyDsJOjo8s+VCh4Le+skYWT5UXTYKMOuLCRe3qxB1VpHS7Z8NHjUks/
lxL4o6E/emcUOXotfB5+inPkJ5TEFc02Gva12imM1sC7g9KtVG7UY9/D+L8l
VPM1RBU/sG2QpVM8v9fuYDEP9EdofAYHjUfDGtOAD0tLI871HH2VhovRW0S7
LBwuYAP1upZmOXV1KC27ywk/BKWwd773lwvldzRANmypwhjAzUIkg3rDX+f0
49VSZBDtbe5B7PZcJ1DZFKLKHt/p1utEJ9Kz61PK+RE/reAxhlw7J/lg+t2z
5adPl8u0bJdDr/gkdjbo4wrxXk63rpASMs9jp2pihLIK7KqagIf9zvEFEvy2
B0Wm074RgZZVBWEeiU+QjqlEVvcBinr1RCgOoExPmTCVEbnxDIIgla3HnNGh
GyVb17OTp/KE1cA8lV/MGfmw+l+7xj84GQElEyevfomk/LGI4aBRQFi/T7HQ
Z5zgDmL8c4drDiscNf7EruKm1ThyLZfAKwVv1Ldws0h0gkL0TZUuN9wTA68Z
w7vWBAEMvyGBVMje1ZViw8Llt3P4VbSnDpjuH5fjaTkPkFYVoItC89s/e5MA
Y/9R3J8DYvoHvD3QU785BhnV44RHmUF/nxEhecsvjDTRMCnKyVK8BeLrPdMO
K2y3z94kDS9W3LrlcsGk3RuV4KxcIPZZ8w12iD5Tx/nZHjK5H3qXFXiX6WH5
/q2EINtkYx6GZHUgOtJJaOlhl49P5cM06jIvUyKQToEvPFdsyq/0rUVI83Eh
fvn4SLlz++ljk5JA/Cr5mrPS2+/8pKh4fDPigKo+R8PjtBw629PnDhMriRJz
ZGqfaK+DgMkPHfppdDaPdJ+cVQCJJj96aYsibPlozJot5cwUkCunsRfxKfj7
ZeHJKYng4nqV6zjYe4gfgMap4aGYlSqsWzGc30RKws3vAoei3tvwix28W1Mh
x5+RwVr8cuX1ONvmvznQgJuGbXtAvNyFO7JHvoqEqD8WJbFsjBsDSCk6Phas
jJ/UfrZD06gGhUHvoYw5eWftmL1xly5l5A0RLIc2K/w0hSzNVOqiMAjV9gNp
V36VJgdS7ywDhRePBOX0CGsDS5u1OqamJ33eVhxRbn7L9U7raYEZACBkUcMt
h+al+WiINOy4Sgj7LNwu+IzqzUf5KWviHAdWo8NOcmqYoL/3GpFFqkHvYtl+
IfGs8lSL2OIsYz5d5rexhYyjII2G7JXgJwIZlTsjXHYRwlnSfd9pHDHh2L4D
HxymtuL5XUnEbIFUM3RKMbnW5g+M9MvhH6sf3swixEgV7y2TYf5L1ZdLgGBQ
C1Pf9yeDNaqiP8xGtKmFez+poSGzT7C01WdVNXo6EBngPokdLa4Tov1Hlwek
iwTrfijy9jjS3hp9nfjJjKlMO5N1iwSzPuME78w3O/utV+BwbXfpzUTU7A+D
YHU+yj+xEqd2tDuTMptWHYhKS8dkJdv4xR89AmFY5BLjwjIfYmOy3mZxn0o2
IdMZAkXlZgXXj8K5Wy1b6L5iglaD8FpKSmVR1j73HJo3dz9iqfLhZJVxytsP
PlEb93/QAWA/DPSmqvQL4xaOXXu9O0GyIUJE7gFgtN83t421L4ooQ6mGToAf
NhBJWGLnIFiyZUBtBS04dmzQbGEN1eD6g1irFVSiQB//xpOlaLrdJJCZx0Rl
B2NnuAQ7lqPHD3DE0o5w+b+m+ZtuDJre+BPfCe3JJYgod/z4Rj5SUSuFNwuS
Pv9kysZ5y4/IbJzOG4BjTx2WXD2N2o3hAQD6+4vMvYwdQb0HaOZ3l/OPqKuK
h5c2c5st0gi1pdJ31Xy4vMbH94WiXqFmQXJ7VFC/0rRYTtPtQEMbXJarPutF
wfpq3dA3dEpjIsSBrXNrpV//4192sR/H8pYOWgapzZnnk17i++KNgDdBHRvn
eFWD6SHxagO5w/ey7oJpBTz8jMKXAEiPq6Ibb8esBBbXy6uVlQfomTimr12m
WhvS8Ha/QX3gm4wjlb1C2/rvkPIR4A54o3uyWrPdP/QtAYuS1Ko5PbuoGSvr
JHDAfjgH5MfNMM/gzZ25DMoFPt8WZeDDXRMZ1yWuF26mCZYCa1FYQU9kk16r
IoBk8FlyySUQpT9W6aRWb4pLsScDsH8an2zd15LtBigy2FHnlt7YkeKh63uN
q04+luMRmpczXkKjw6M/1T9VEdzyGWYxDATVa8WhDGWVo/E2y99ndYOS697e
xhwodRDeO31Xd4Ul36e/JKYz2KnkefbElIp2uDwdqgNILgXwhPQZuBXVqDze
+SfsRRfoFPcOC34xXwP0OJygYAQ8r89OwrzR9ppXh1u9foYmyRNZFe4o2UQA
MhqTk85cRG+KdboFZOTRnUMUk2SpxtDxdvvn9uTI3diTOkjSEBZqPJxWqpz/
fXBeN1Dp/Otb692kns1HErcuMsoq+bqeYIDv+wqdQc1lz014mmWAYBU3Z03N
B0oDONgafDoHztfF/OL913D5Wx2zaK4GFHx7fTfdyfXPkdOpJpPpOeCuNmQI
c8up/vOH3ZpQ3Pn5S2RGQJ0WlPx18lhOqbyEZdrMBLUM9s60qMG69sbVDT/M
XhG69Atp2iU7wr1Z0nKlAHigd/d5JxcT/bn59V3EZrUt8NBGKKBK8u6oIwU4
ShtarCZJi+jVspPLP3iWqzrmlbTp6RFT+akUWefcMXFhPZZB4dGnnTE8WoIL
XelRW52Ima8UOBAytpIJbVKzkGlmxXML4ueC1k3NML3PYfOkq8haN5ribKeX
99MoczdQ31K+cmY/HmuPFTDS1YKEx7B24Lp2gPoOCxcOEkCKHl1Gmudruw8R
b8T5xcm/bIUb5xw+IaLsEXOczbYsOHmTugXZC+962C7W/CvqSbEbGFfIFKIn
jFe6aQo2FAlha0cidyEo6R/2yY7oxdTyLh43lp/rUHEnWqwidTg0BzwsECXT
8frHN3du7hnoav4YSxsZgtulBP+3vPaLwcIymk6JmYEfk4t62JBkMapHmFf/
05sBUvU3t8fMKUCUq0N4r/IqzypiFesJG7cBHCLQHvgLbo4k+wvY+OwAoXs1
qQQAtYoZDzwRNrzD2ClKKJGwp50Nk8D+KuAmxYX2mGufu+Lr3SyN/0ZDmbUK
8ZWfGvYyA3MUHYwhiaR9GvhveuMiPdUSs4Bd/3YuZguJ0D4bMAsFlvf1gKnd
RX1J32OOPUTTgZqHSWx81mrpQdG9RUgCLr0EKM1b/szPjsGGTaIKH1lWwdjg
ePrCM39nHe6sjdtati8+sY3zVBacyQACahEEx+UUlFmSvAhf1lEFQ7b6KvWs
rSb/UXGkrCn5Txf1FlEAWFjzYJuQ57w5d7xXr78qw7VE+J9x5kAOH4Ju6IHc
IkqNS8prYFNMJlPobaAJ0prCHR1iJbUE4UXbDWSn6fyJVOLIoCMe1f7EwITi
SGZ33atbEgUu1n+9KOYFubKlmynvEbs9Wdyn2B+8m+sUs/L1UYB9UbwkiO/D
Teg5QTQjGKAC34eLGmPrsAoQax9e16LEaVjEdb0BnEXLGCIMgw94cGXx51D6
DvYZxB7oiIZCiMRoifHZfJ76lGwlHuY9YvDjqHQpGlGz5K7Kx2+DAst8A4HK
DNbeBqKH+BuroyxStDbKGlTGNjP0aB9YDylSFt8SslJbusCZAeKrHPFho/dI
X5CZijF6R0N1ioN2OCvp1cH2giMe5hOcYvDsLSzHZm0zOsSO6BN6rlVzyaeQ
EWlh6NwaevbRz4nvBKt7OTWyeWBkXvEDAw2Jmjwzh4/pGOc/8DJV+xP3j54B
H7aINPiztKX/XJxtZ3NNPoj2mbOrtUhAOZ3n0mAHgTpWfCjWlG1ab0y77LsM
QuP/decDLrikFgv33qUC1ed3VMRIZBL5/3DqpGirMzPeLsau0xMVai4AbmyZ
domqtPHcU9393ONBK068uyZ+hKvn8n1ncfcQAeKuTC7GGUMo1RfCeem/e3Hy
WxJxKyo5dkNnsruYOZEJtapxkExq/pUwMcZxb7WlZsNGapzzZWutdKy8pykn
kKeKCPbqzZpsRzC8zFdVAYMWnnVq2S6qZ3PbxDWRrVaGQlfhgDfkdyN2l+/r
WFLDmoNY/AZw42qkkuHjL9XdKHuGpCjPhQw+Grw70LU0z4w+Bi1wJxW8vYOs
o6AIOVSIKGcg86aVcqLM+4TwnDoePhIH8u7eOoOWoKTSSfDd2XrlQqiwhCE6
+WyIv74G/0OalQD5CY2VKCnoIsfVbrMwwm1nNCgBGMDF3GuqJGW+BV9gtt/r
VNEsCvoi/JQSLvYGRTZWJ/xfOncSM2fEiP5ySnVgcnZHdyb6igNcIJ+6YOB6
WQeUt7GxcfIl4S38ppOfbN1VwPzmg4IkDpjnqCr6u8hz7tD1oW0t4sXsDri6
6E9uJeTm8VwoUr+H0O9BX19kt2ywWBFtTHbPaGyfEL1RRj3sUBaLQWlDxmIM
F/mPDQ1hWZofbxJLt5fsAtfWaenfo+NrCh+qliLVdWBSDn02uhBDnoGUBt5R
S63Gg7lyJLXs0ClHjvZxFH2iSjsb3kpeQMZswja2fxrTJhgHwvoMO36jdCIy
w4npMCVqXAaR0woUE3eC8Bs2VJ+7pfZdx/ED7xRdqNvcq3pR5FOkvEfwfwUw
CaXIT6isVF+4UDNZskW+0tPQjhCtKJWOkCOJdFZ0guRCfzPJBKpNqxAWvyaL
9D0uVcubdF10Kw73wtj7pHuJtSJkkSRp+XJNW36I7JHTNeqc5sUssryBrNNf
IMpy4mpppIXcUOrUHcbSs8gXCr8QqclFbkDkxExk5RGH+nk9v//yFiPJ7wq0
p4nqZtyYKL/ED/lMX3xXa/zlLbUdZZjJgx+G7QJH2eiI+tXhyrlE+xoGZMIq
xRNmpMq0WIvJLZrQY0BI5PEvEHUJ2kdnmoTEYTlKfz/wRI3SU0N5U6ysOoSB
xCElje2wAWw7jC4v3i3xt31B8nZ/2K9qLhwTqj57w9Fyqyvl3i/82VynROT0
Wkkvtfjzung1KfkIOskYBHNm8Q++ItJEY0QDUav9OuLg6ylJpv4TH27vzzZQ
rOBgTTlCBPfhOPsvgr1eJnteOwuFZcipcKVUcPagbeIEwMUX54RnT0IAi2Ue
GANHese2tGRuSqsqaOcWbxeSp/Ew6gqcgrjvUUNiAPAlGAiMidjgFZhlFiDe
VLiWdEoDUqlnC7+ihIRXxdswSeVeCsfkQ0EiD5KbygA0TtllcMK5aP27/1uq
X6LEdrjuuyNMUe2z1I6WCBdE2y63X+07ChyPnVZwC9RKMnKzgJa0nE7a5PNN
iF0XWFGmvTLWw3qnPZNYBmCoLAVBxq1aZ3H8Moc2zI6oawUC8dfGGkkUFALk
UlPRbvy4hSwepwnduCdv509SQSCtYLurOTzroG1jbeqW5U7RzH9ptRQ4SspL
asLgI5Ae8TAfV6EbWFd8z+1q76wAx4ZuDJU3o4+5u/OjevlxzV5U7XLHm1u7
iO+jPlTNdOU2DNVbUjaOffLsl87y4Zb8KpA0JecziIGOgUWaPp314Y2VD+D9
prdTHxrvs08REc2DTEaQSjkSpkgSTuuldjRw3HKtMb5Q+xW5oYuSOnfqcqVt
LkoFozMAETcL92mS/wGtc9DdC/3hmCgpn6bo/Y8r6UX74WtmW3PEVIjHCTsc
skNBVqvDhWJG+cOtDTvcZxexHz3S2mFwlJb+xLy0BAJeyg/eOpbtMyygWI5x
MRlaYLKxtnaEfjRbjS2H3/a89ORvpYtn26fTi1sPWl8TTJFM8AC+oO3Vwvyd
IwKiBiL5VRiakPUFRNQVmEwQADIgX8WHl8NYWBfH7GgAND3TahNO78RLqeiP
Hx19ENqaZo5Zdn7rHkTAXXgY7W6aSfizu3JN7Zp/KQ5kwgnnYyMM04DM1swe
4TWoE59iKsckN13dslaBQwKf/P5AsmWDKKlF7d8YSkhYqVYRquEp18VaxPbU
njD4KLfUppR6Ye19IWTRC6r6RT0Zh7i/PSH/xsCxwUcNyrlREJUY8mRu+MNv
9Ev2zirHZ6Xw7nzn2APYbu6lb1sbspqvVzW3X+hUsKGLGWCWaO7o7/MqbGKX
89vULimqJYa1C0qLW3R7bbT4XkZhZxv+4O7MTCS4jo3B5R85h2Gn7qfzETxj
lkhchoXnLWLlqTaCKoFTfUV/Dz6kjvLEjAJXegK6G3ko+fc+sexexQYkPTYP
IJv8KWO2kDgrFHXsVK5zEQeTPg8PugJgdvVjs9c54xjOGGsqAu2FHQ231BxR
5Rv0KbKogVSuaAj9lEf2EStfzWhhxsnGaM5KhfLtE7YSVo6PsjA/Db87VtMc
3XrnbgZFxAQra5g4OD1HLtL1d9Epb4owk0BPrU4bTuCoBxIwJQZF76m7jgBc
2RxNQlgNlF768i7SPCVTkgQi5Uka9H2Qfn0E0XZBFM0HoweES5IB2RNtz938
tm77h5x11JdlsIhsRXZ7QJCc28gOYxQUEXAzzRK6QNUtegxCY2Hb2l2ZdR8o
a+sPWfur2VOMI9Qp7DjuaM1rQjdBKGhsyb1/Y/3fwaVxZjJv+yEvvqibWdZb
/XCkJ5Oopo3iXuT3At+r3nhGv6oEu2kvBPAzVayUQIGDeIO9Zi8O1lFladNs
AI+lnSt3qdUTutKUZGdvJPGulujgMhaVknSMOEeWwSE5HG18z0/Yhr6l3ceB
/1WT4WnQ3iee4hrzzR7zkzCDwBXOTQ4Y/ahOvRN37EIKh8FZXgSEYUzpDfF8
PtUr+M+cBwiSmK53yuzgjB1O4co1jIArcUXvETfyXtvqwxRxE9HQT0NFyzAG
Ef3x6j4M60j/EvJ6mYTjw/820Y83XbDg9aNP1vGCJj6wzgMMhbkU+GRmEkji
HS9q9RxyWT/d7mUJwI4pKcp9RGrJt1mNMgwiLUs/umAulua5rTHE6BcHunci
RE0l9fru793KGs85X4bBa/+919FkkIYH0SAaDXVqHgerr69bXk5qDVYLNqys
4mCyGUZvOwdF12plSMpRUtXBJhZ6AJH1CbvZHIcfsx1Nsch/m+nmd2Fyc9DF
JvJu19pwbAGMdfFn9e5IqCJYz/TKI3OeBVijtThsGt5IglhT/GbZsk4zL2IF
WtKeJvxgc9ooetmBi+TPirdmJwguzPdh0jqvpSVX+lVvlP9AIDS46wiyiqXI
sjidOnAqOQ84K1xmosIBLrgIywQXO/B7OVuFyX9rnXB9ZUHpvDwCS8ucZaqh
exvJiiZBGFyTepvWDYezOD58dPFEz+XR0Z4COgqtrlDy2exQSTNH9/5DzkC8
SO80FD39WtHxZP080HQwwGqU/Mqg27AR7hgxkf4RWLAPGcVHKf8OXY0WGJm8
r0y/GOaS6i/G0Xc24Mb8nV5Ja5Yo/Fu5C8ULUjgfFS2ZkT4QuC3sn+VAn3Kb
8+KONEQjDzHO0Acnw/I5sy9s4N50pHakUmqUWX+srQ+uHLO38O0K5qnx8WQJ
YnbP44N/q88oDFY8Evibn4WP052iGXgYN2bgAbjd7SGPhjgL7eO1C9FpVU6P
9RROkbDzKZcUzsW/AwKuilD/E1yRsk4oFZWmUpRl2d0hvvMC3v9R9ftIdu7Q
tAHT8h0LxLzlMQSKfxK0TAiU0mhZh3CNV7EyY1wcj+r5zc9U1gPiZ41Ww4ae
0NTqIEsI/abjyu89Rya0aI9UK1YxxWHswQOumhknrVV5m2CnA60XYP3DTMr2
ELrImBxJnW/JEEDNnnb+rdKQhJinQB+jpbARoTvkRJTpU8gzr8dZ81Sprwbh
+Qso9tSceh/fkSkim/XFbRZJwOLpK734qlbetE7rSb5pvOX3wVwNNErzDuTN
8+mhIVQ4N9vvsS4Ilvf0WWRSxwB/+mUfEHX3hKmbepkY2MxCQLD/LpBej95h
y6B9IP8qdcrVVumHs0/qm554c6B7vhc1O9DPs5XEAsfY69ojegpD1MV0015o
JgN10yeii4LVJrK7muknqYAlZ/hYIHkXOiJkamZln9sRjjhNHmaTEyH9T2an
YMMaMJdaxGFE/aFDVruKcj6sIn9oDwub79l2sW6LUO8EqtsWBvGnbV194s9b
C4PtpD32ezblrkaeU3fRxhlsSLyB01/qYN6f043hIYY26CcphJykQ9tncC54
fAoTJgsNUxJgGWWUVtwLKprrV0+2ue3kxe8X/XPaIuC2ADBe4479gP0qcc9u
ejwz6skUwhw2rVgFyKp1OKiLTtzPNfNkxU9/dMASCG7rXGaj6wV2X2gTnRFm
hGVwSi+e8tIZH5+vhDloXy1e1fEk+pnnYuCc61rHDbI3WkOjxu8jwFxkOUOt
fgdNyGa286FeV0dBxgX2G6tyE6yIkEV67NRhu2u1xbXMqI3zubFlwadcW57X
Bk33D8OjxFiMqIGUV36XG9Z/6H8Jpb2Pyho1PhAfbCa01T0B8wdtnsEEweoy
JNYQy7Y/HLbeaV/YcyAzeNuZMA8A5Z0v/095ReyNQSsO4zIA53Obu6V/F15Y
bVZ1Yfl7X3AO9Zac30nKxuXi5kgscgX+7pMzo8rCQX8tY7FeFyIbKC7Vswjs
Ejr/eJ+ZblU9v9L+RLMJLnwSvoyj/qvzaUgz9ciqqAKhM2dIvVZSBu4K2pBt
WUeiBKADlSKmDO4XDbExPrLb8W2UbmI2dVclNgUZuJ+VcyTP/cny9Bv0xYQv
32lhA06s3Hx7avnEH3Rp6QGD/0tVX6UPKzPfndEwFStoh3i8gLnzowvCcXJq
mSaDcyar3HM+H8E1lyAX6TU+tt7dwBKQeJh+JsGUTFnFiC5bhNPQ2hMEUI3E
H2J+He1N58MV6vHlAtjWlItTTpY/KeHX8JBMbCFQRXTC2dGkwYB1cNhlm8Lo
FnQTaMZXNpT2S3lz/vdviTVwgyy/5m4VfworfgDI016EOYEO86Zj5EcV9X6u
Ud3RLx7XMcHdu14vAnxBXkXT2wTwN2GT3niHOSbZVl/spU+JC2TiQW43GYdc
OvAbRSoQbjIqp3ubbvb6+v8V8EFFfVZbC99sKBhjgUIahBDp64P9ameu4hhy
IwRhDTp+LBZ8lNniAuuZDTiu3eSoNBeRb7Vvd3NtmK72L7iHpCbHjoIvpehJ
g94hmpiw8q5usZxYvtqBmlXesnZgH9LU3jnooJ6za5QdOr6EPrWBgfzF7o8E
xTLqa3sUN0pawgxioF8Rua6pNVBMtQm0q/qVU14Yh24u0PTkYXeufgk4ucj/
8xZyFL2yPrzC65jvTZawhDe/vmhFxujlhcAYJDmn0L2HKLNDQX9tuwfwBI62
hiAhRW/p3YMBIvzv2mY1symGUpTGa9O1jDE8zgkCc234D829lrBzFvOCXF8a
Hw5d6iBp/9+o7oPzTQB2v0Ceqn/v7Px2u6LhZ4BUXJQ9l0CY4NwMaBTmigxF
gXkWscnSBqde2dGJHJkVMh4j1uOTH6VFguIiEUBkYkdObfyuMj+pivZrUTHt
WIUR+7EOmrmhFIy91TN0bRKbgGaLktz25bo3uIMGLEsI5x2guHC1EL6CZe+P
0OOn9rrokIPBeUDf7oKotLo2+XhnqgyAtKhcVlNH04C1J59LRkHPf00PmNtA
L6PnQ8LxLK+0P6y6Eg0CCWSSwp3sGXHiF+wPQBCR6xFvh9cWrRdksmz8A4Wb
YrcbkvhU0qv9OQ7g9nlQc+9Rd6snZl3+gdaHeTnYfqPQuVgKlrcodKFog+Eb
ekrnGWG/BDkNs2BZPCMKXisA5py7oI7pb8aCGLnNAC0lbhivUHGzVQfHAeQT
aGXlICYf1YdhIq497R9UaEQt5uXIX9F5bQjKnLM+LHeyITDpkayk6nCF+gfW
CeHgaL9So/q5ie1fOzv7NjWVklLbM+LkduTf0eXftqMLR2Z2P6BdLWXH9slB
dhRqrdNY1DqCKf7OgFoPUtrLzcrEah31fhaopMgBqTksUJq9wou3k4gRClSR
vwd08hgYtC4gH+Ouu8miPoZwx8sSWm1KzAXTQ4T3sViZVxkbkSftjLbdXNv0
jjo1eWhwC8vFnoXuepK3neYGNPE0jDJCC73fnDanr2ewxIFAgXet1IWJP5cG
mV7S32tfrrhShz9eLf2eksa7HXZiWlye6ORdcE2i7l7rUDeVuV4ZAmMF8gxK
QrQNm0gcbvhhJkElJkl1vR5VZS/0n86h0VLurbIty/CjlRiWhBAFWdVVC0UV
6f6L5zqtqH63s1segortYwm/+P93nBAFqoFHDGDvm/sSYSWeQwRbpc01sLCC
Gr/mCgnoEynWv3FaPnMujwfS9E4msHMtmn64vFJLnmnmgc6ewvm+Gms5ri2c
ejmTzaeUClJuO48px+I6Qdubjs1of1Zywyk2snaOxCNGUUvKYMJsyPEnPQ+D
gAEo7kjdB3e72cBw/wMkn5Qh7jm307Lmy1rqTg0dtWqLkCGCUc1TKMBCRFGw
djrgASjBCoVM+PMUFUqzTQjooQ5lxMUrO20BIOT+sKvxQ/OGb4neNIYbD7NO
/v8Q3KOOQUwwDtQbA7gdEB2Gb6tWe+TgN9+/RgM752E4/Q39FXN8QUijBXSM
X7RYL8lu25kjB3SlLYNDcijP+McqdSnanIRYhm4HQnP3lvZKUgYEuBj2iPMX
CyXKjAMaVm/W1OSTkWN3/9t36lb78N7eNkIhhdHkPkJQMlP+ym0KmJ/2Ruz+
YXEEdKQvwbs8JIfux46InFf5R0JJ0gA7Wh68ewThOGcuZvFKPBI0Lw8IR6tt
AAu+edW4nYJNu+rAcnhaG5GJZbw1W1nnZ2nUP6ePHjKZ3la8u0GrrViBrmX6
L469zlHnkLOvnjO0HGJA0oIuu061eZb57hpfqXEceSCg2QR7VDnTdhaY2/VK
vHzsoAcyDXOhbRwahl+6yvayh+gGgh6LHZtPTfZLA47/M9RT3RPIzrQnuG5a
rDmJxkHwkwLRzAlBH9A6DXkDCl93AFTIhANBeLcYFZeyZIM7dZjpe19jv3EC
hZjMXx9sbI/YT1rNYTEPjGTZG2we0jMEzsfmHltTygtzgKpU2p5GzUNn8xGA
r4YBHhiS/ldn47M0TgPPPpB5bPnn627K+QN6QzCSdyvds9qLnST9FoN/diMF
899YtQLl37jQVvA/aUwyjkXsKhuqD7dyulspD8juVKjYZmZN5SaGRURIMTNM
sx54mnCfiM5Ghw5koTfR2Tf76VUR1s/aF0dRLj+EFO+LT0GPr9kadtKd5aQt
b04PNCHlVQTcSW5KmZ/A89Xt5Xn5ugjr0Oz3BuvJUFfE6DoVcD/hzB56ZXTs
1W8kaUiQg0G4NxAy93M0Uv5y2Gap0rY6sGwxYgP3p5+KoPg71d+2ANagouyu
RuAc14UfIwsRo02dqXzHtGwZRym3UWOyq2r+ue072/6IGjBH8jCrJAW2HsgB
cZj5pWU1oyQjcZET+6HVLFAvt2NWJBeOP9tdHN9rPLBr/pE+UhNL3ra28y7B
WtgAD5Td9brqT69aedLCwWjm3CBQtykcG/OJEZHJ+V+LY8zM7fUmH54A5nwT
5nVewZmmmFAhZz1zUJwxWqg/1lDOwM8JcP0m2QldKpZGPdnOQIkB0S18nDQg
rRFSP9FyJ8/hQYxTVXqlirphGpSBVwoNuqy1aY8JX0fsceNoHpxLzuSgmxiS
Y8WKcqKnchVepRVVorUhwfsd63anvKbzaJk38pBDqM22qDylilnkNAx3I8+T
KDAokdHqAp53mMHGJPDcn71qLiEA7v1imwDlAYQ3oaYEb1TFUirhiwkujuP3
N4X95agPjmi8xfYWX7PxHUjuwxDlU8ab8+X8Otwzczu+Vhxv2YA66XZR1beV
XBAUjHLxd2QGQJ/wE3oWJd7SlQyAe1mWvbJAoaRvz7Hu+dsGIb4giEohLkd/
I/+aciKL0wiVtbcIQYuW5hM5RmpHdIcWgytd43auDK3ldNnPRvUnqTLKpvjY
HWq9aM84SxPeTKjVfeb7xqViV9cMY61UdIs/RJkGU2h6p39lt+ycaJBa7v5r
Tus4xN4gpU3s6jnDpiwhPer8Ds5dqWnjHeWvJniRu6GgeWPoQuu/fCiEQ7TN
rPbpkC7Y8sLrD29rNYWjHFcZSzVJyLldh1NT47a2X3p4wCfhQWcveGYs0FT1
qazGvKc8fD6q6rnY3Ojc28RqCPv/8IDfdp7sf84XMYZYusFFKmgQpwV26+Sy
s87T88LA22R9erwVgY/hnQhfSo6DQTlOpivn1rnqLzR7ZzQMetrQRJXTD3vu
XIbeVZHa9pU0D5WhNcddQHhmgtzK0ZB8YeRhfkK676PxH1aW+W/O8lDN+Nei
3OEq4hKoreIoatGRyTrwlvkZmAmclcadxky30DcWJH01ROeot3bdWUHVdBye
jQJuy99Rs+AYAqI9slHXMLK5B0jKY+P1MivzSdcbzUEaQmoBp34quEbR6b1C
0jeIaHcmoWCNAd/b0hP9WzLz4nvQmvf33uMatCNqxgW31R7AR1qRWpwy72XG
tgyP7Ue+JfDKgSV3j1FI77cXlXx152wbj5bZ5Q4AO2/a0GD27X9cC2QXbaBH
juO5w8SEmw1NeWUp7ozeOdFYzDnBH82oUNoI1ynHJoYOj0QWq4bMdw7ErQdu
E+lByPYwDT1fYx+Ck8f7Dvxp9aZGw39f4F9K/MDGvWN7ITcm925EfCkLeBDK
yMJ9ZKprSSI8Qn79EFOJEdROSJp6FDb3MGyzmDBRg0aqZeubVrY1LI2MktD6
fqs7mf6sLhTy30/w9GOpU4bBtDiy5Qnpq0ApxOH2VXjrYV2ECXSao4Vq5AaQ
/dsJLYsQsxiJWjDebhScgYU6F/l3WNwlY7ow6Pypb05algacVMA0I1dyJ24Y
KUPsPaB0+TK6ZYtH8Naxw6O1PXd4aFD0GpU1z9O6aLbg31vIx8+EVR2N7MgR
zPnVZgKtlmvHKzkZajRspdu3/6X7dTIsfWoStDWQGXON3yKIR7cfbSzPObsG
A+8OPeguvCWvu/8pLHannMxJy1/8m8K/yq/Y3VCYwFoxu/rvQ1cgF63l2OuJ
Ug2Qt+LOyhyjnFrDXfeIvzgXTsJgz9amJ9JV19RS/OSbmrJaZPDxOme3BkpP
KNnS9nbQ9XKC9+6tc5/SglPrExHkWCnmhecmN9EtNQp1TD2vnusvPo+BwFp8
Zg6PyPLqWlI/IRQyRrxg+f/YucBJibxzrg3gPiogrTeL7w5nrH/YLrJXwCDG
kFPLJH4IA9Yi+Wy9dWwRKTm6Yga5KcHaul7//AV7km5TjiFKVHMKfxW9Kv6X
vXK9XdOKT0nbREUxxlljR/nOCnLEHw5tqGt+ie49ppJ410Qn534k7xtQPd7D
9x35fVJWQiCfMdTffMqzcxx+Q8hf+T32gSYQVQQBo33Lc/AtxLRqGdB6C3s1
hi0MD11NE3KDW1f5KIOZdJf3Cl3Vm5EijVdXWCbgGuY/dTZaZJ4NMnIVjKlc
PQnFKxblEXMfF3iuvcB2Qkqsht1ZoB/rZQf4jiateZH5+MLlr/6dc2mkQ3Li
4UN8m4XdPkKD4V9Nm3SOckLGKqiP0muRgFuOefScx9o8CiEGl18ZRfhvYO5w
UKXm8PfOoJu5kkIy/Qa3MWoe/asmkmvFMpoV2ELqJ1s3XcIEUEvOswY3nBM9
Iso0ZmHJ2BOrhSSkFMyg5DBuU8c0at/jhp/T0UZVREtdS38Q3vNPGTvxEGl3
UbJCQNJ2ZfwbI2cHZG3G4RxWOzbtmt0SWVyH+Qyh00iQlzCzHp8/R0C4IbJ7
/eLf4NhN3W6uFUuQj4uMSnf5/a0kqYSKTQZTBfBbG7Cf7h5xEdiSC/0IzQ2/
izQpIesj9a/cjC3JxsMOaRvEScks8yrQnFq4kInzgkRKhulzAWY1wUpTHeoj
WaSHDzcZCJ4Iasg2xK/jLPFwXFSEBaBxWJhRK9AVrwdoj8WhbXBsTEufflNv
Vepm9XiTFav6GN7s4w/klz38InRTvlgT5uJ37NLKr3ToVWAOsjuIZdWwxZc5
mzNgwT+pTJnDOWiiLA/x1W9LnCylcP3p2ALLX9594/Oe34gXBYVKVGg8skGf
K0ft6sO0vjXxIOQXqLFwgfmaiaWnxBXogRlyQAEikBiSUGSiCXerk9Vylu5g
Z77euoTK4OE6587SO1uEUAe5/GYvqFQEbb6wvVRxdKJVLTFLxqcexhYxoDVa
OHR54nfRbTxxNT5pP10pH95BXZYVk8qFHDN3SdW3mN07L2jE7VVbCR0iHWVe
l712t/gmWRhtq091k8eA09R3LwfwxYlWczXc7vPIIWPUst+uSMqYfgk1cCCp
O/Ly62qEZB1MT1Iw+ckBkRezTJ92zijYdNvyCTK39VyE4f9gprdkQQi62tjE
oFTcZjcX152n/5tulnyk64BAl2Ny08bcL7GF2yzN5qNr4Y6zog6e1Jy5LOh8
yfzNF0l3/VPYeSc+gZ2Dy5BBy64F06qG6jAsPr+ibOGoZxLQFxkqQG8PLtZF
XSwhVpWAMzjGerRU71mAfA8Ab3YWR8Ukx3fcLZHO3uqTFmKDSNsVBmPUaKtn
qgxYm53Smv4zNQmRqScnU4rE+BqjhUmVYxw1o7xPN8zQRw2QgMvNgnbAWWvR
v8hluF0RPWZI77PaWUc2G1+OvL1kAVzO4OUoMSgJU7Bxtisjd50LYvi1TfSS
ky4QI0oUUOGrXV3HFue9duwf8YT0oqd6nyCYpjQ5eoAuy9k8Er8Wg9poNJ86
rsmUwviPnksUjq9NNB+2WvDmghKcOpCK03InRWAVeu4RMWVL+5hgdodPY/o6
LFB5eOF0L4h0PbuzHyHSIYOKH2f9p/jwEsJDS/Ldtk4JsXyOX0aIgy1zd+Ag
iujMViKGD0P8muMMnEp7+PHSu+zmrpPJmG52NK4PrvXiTuHDJ7QH2KV2Xmr4
7cBwFFIq+GYlbL/9E6NXfHk59yaemKFXzKd9c/rw8xm+qR2zBENp+yMkMhNp
nCUrlk6CWILjIkcQU0BSvlsjB7xSMtIgzsbKs+CXzq+Om4/4xeXoEIwmN3Uu
bwP+5f08yjvuLaQeec9JMmRgB+crWZAi1CEtfuR4gHX3NBo8t3Cn+ou6Me1m
ahlKa6tMzhbEIj8OTEuAlaXYzkNKYOIaajxe2IfQpLYUnOzH1HZ0nyYZkEIK
BcBWlh2Gp86wSP3gM45EXt7+8i+EijOseNXv+4pMBVgbc8AaDKHMQ4E0vPlX
S5r1olPhV2oWy4022D6aKg1nB2zqWPIh45JZhpCz/UWdi9Dc6+rnOnpCci/4
8aERVafkYqeXa5D29QB50sZodnKby0IakASG7ewIITzSwWFRelE7TtTTsnYa
/Kujpgq+aYUwmIxp7drsZhS2g8pweS0VAW+2v8odcaOJEUrDnXDpaIvp4HFr
MydsmAGyDDE5ZWedxc8ns0eJY/hYCmUVL3BapkVDKiXZ+jzf1EwqFoLZARKl
/IApWJChCmbXGF73Y2nZs7cyKbld1i229c5Xucr7WOW4BnG5Tp0KdqUBaMd2
6xw9TMGYUQNxCeXsC8/vORST/v2OZmYRudFhRZmiWwiKoKBBHvkFB4Vxj2oF
FiOPMLv1uc3yXHTcXx5RKBjSNto1HAMp3pTd7V0ZiwcZDhxFAAj+wqwU/nXw
bRGFWA2CHpDJ25PYRHBtEx2LUSbkoIZF3xERhi5oFEy017v1yXzgk8Kxiygh
J1E/w4ssA12Fo1cj8pddWWw0bi4cNdv0rzIv0rLc+9rb/3We5VN0VEcaVuLO
QX/WfCdNATj1sXtE7hcKElkOD+gWifUvSoIbJAiyyd0JJwbNr9Bl0Z+uWRsb
WPQGlS4ndfGTbHa/9qCbv8c2w/P+ViASvFCi+g7+f49mxEzGujFIf7IVtvXQ
pCmGwZ86B8bPikTGtabkgXHt9rACJsq8g49zjwKB6JprTSWSmxWZan1Khx6e
qiqfF3MIGcxwythmwqLQcjwthbU7qIYmW9vcTNBVJkjnBt1G14yr7u1VrLZM
h2tPcXABO1c3f/nL+dCe+j8OFAq+VmpagTMPs+IpiT1/+PJeR0IiiMw5YvrG
nvQwOGQ5d6PKCxeHIRslrvMcfeevIPNGShjgkP4HFc0T4JVl7t5BDSaba+f7
YYlulQKUlGstOMO3kZEUBo7+6M5pqAgosbko2XzrbTP+tAv2rHx1SoR7nllk
9ALQhlZ//oXWRWO6GTTIpWod3QynDREojoDrlX0Hjji3uCaLm0wAoOo+1dq9
irxCg7GTYBPyHs5s06fG76xypNdJ/fRJAsKg3k6wF4TcpbT6i5wLZkHscjDc
ytJ4Lv1RvRJKTY43EBqqsRyaSIWoWnpsl7Mb7Zdh6olt6pHNc8nzmXP5Ialf
GSAoTm/NaWxNaaEzaMHdt1t9jjKtOyjlc+3MpQp5Bsn8awnCyX8kESwObmJm
MgxfnbJgdyolaPRhNl0C+noMeuhz6vm+NhHBqVFxlUnijhnU13Rw9EFwwl0o
OKPSWGzZ2SN3eYWsIrnWChzrndwJTZZtGZjN2oDagv4+ySZYcOpbMciu35UE
cyeBN+YXu4U2lpV/yBInPeymt0fdp/HQ6sG95Cfw21yerH3ml2sAgH95BDZD
j5eBoGbN+b+kJbII0TkvaEKpaLuS1UzEr7ZuEexX19O+7RGOxxQZ8wf0urap
eXUt2stx8fDjwb/3PsOIjtMh8194vThTSNVr7R0+91mqZ4EnoitqrYVcgfJV
mzrO46ypHix1x2e+jen21OJiJ4CcKUMLJgojnPoFTLj/yNz+z+D1aSjBASYa
dEtSBMxpgoqtk0fy7x9z/Ou0+8+RtOyVQ13Pkc+W3eauNUwh6y9CaCP1F8wh
UNulU7nsSBjMOXVIUtTKtL5e46+X6RvPTRygkfyv+bMob3iuSqxbEP+U0XF+
ghC6sgpcO/TxXwL7PRBBpRnKjAnnmpTkU3wUbc+HkcKuUapSW0ErIz+Lf3g9
goKfe6rDzahYvmdCeiekux1v+Jwdb3HyOdVBVzXt8wLFZkhd3jhSB++2+NNs
qb4l2IfRIGu1UMXEjDwYtj/Vl/Vy4Licc5oSB9DB8bqYi2ONLjHhkgr/BRXH
3LNBBwhmdr0cL1ri4WwVvO5Edgg/CUiXWZPnSfdW8yGbKEXskP/3j00Filmg
rLUJUsHPeE1Q/B2UIc2PR06eJ/B3KrCrAmIiEW2rX0zI9ZLXBJK7/pEun9Qs
7BKOCrlBIRRbkug3tiImU+3vtRPhOBhLBob0gi+P33ETTk06vd9H87PC9YTS
Xgk963qvGwqOByFG/KbXYKSs94OTDZtKHcX+CC5jBfwnHWBVKR0dSZ6jB507
IEVL/It9WtVtXJSIf3xalyUpvfQ+Bj/3GovW5aTtPA0IGjobq7fOFZjl5Obh
aKmbbB8o4hGxeosPKjBu/kvgE2GpENE83X5A0bEEFj4mgce0AYGQ9NIBPw0l
i1dw7CNxdEZrYmOqyzJhjmpFjkugX3TAjasgYph7WT8x7j/mzllXAkFX7mhf
Z1WQM5ODIxiskgGB3Cp/l7DPAPkHQ88fAs3wrp4PzN/lT0n5GRSFlTJloxng
5K3n+KEycRoG7NLIZ5LwT3bOGrlMbyEhNfRsJh2DxNKLzL83aPB7EpjJpYfq
hAO/Ob38I1ww3l8v0qJNp97F/E7d6Uc85s/1fmz9NtHsM70XWFcIA7z9lETQ
ihVI06i7cR6ZaDZ6T3sQxiwa79KmPkOQT+WZxttKVuKZoOgAcfWdwebxSLha
Bh+vwR/D9KXgipWBtz+rTlOfj8Mv/2puaw67lzLrTX7ezqnk6kA4Cv54Mm//
tw8JJY0l0h9jQ0SZr7gkwXv9rfW91dvelD/skw1xb9jgFpRNj4oT7mIXZDgy
UymnyDKCu3+x0AHXARaeHCdGbNCavh56i2tG3PoYsD2JQbFdzX97n21P9W06
8/M15dfYWj2Ee1PDlQf99ibcxGo+CSULVfHD/QmGhNybqFFa3vYTphc3zKGn
KplE8NBinYLpAQHSY7BpIgW5qTaDq6se8REeX4YAmTQbE3yCQIdwdq7frXij
esRnN9whbI5MJynP6i3BVTC/Z2OCDU/pZcHuOpwbwN0gHV0X+NQ/O5YQS5r0
2q3D0ZThZC4CzSf52G69RYjrBhIuo4pHWz7QwSnBX/sYwy8zRtWo57LG3eb3
e+mjgU8givrJJ/BVghshCenQfLPuISkXU6E7Jxqlxsy+7OcXD8fKOJso8Dao
HJuEchsQh7HeZIOF9jezOAeFHOlj9j8JTFYK6bPoK3NDB0s5aoXjcbPCGvhj
FEDwoZWAj7P3WtxXWiWPcqeA+ijTM7gnf0GDCSy1IwMtHZwdfasjvQTP1K3s
2UjMojCNQ062MSFLEekpFPMIm7WuDuhLBiX+y8xQDxwdFW+40rwdJVoYL6Q2
XxOvECSAB0HFoA/MAFRyGaec+5ELmYm1SI7CAcaaUk08Zhm6y1ZXL2KuCMsZ
FSdt1lomytZpA6QwbD10Txmslz7eWx7bv8T+hysiALzFTM44dxLy5yesswQW
zYYF6iGU+sFEC+VQh6qDoCibncIG0gJtctRSIEgdDX8IAGj8KI/NRBNcckEy
4U3Wrr3xEVEi/5KNhBh7BfxIhigs7t1LfLyaX2Xn9LAQVSFVa4GLZpkX0xso
bFczJkxSisH9+3R/1WjnO2bzP/5sU9p3QEvrNpVSB+g2FsuXPHjx5vFGX+HC
jRaLOr9wAxYBRn0BoZRpNMUzyEvMsd4p2qekA2x+IhB1dSajFKqTTKwl3J+2
czaqPAbgVYl/sDrU0jKazOozKDSXYWVevIYtyQV0h97OBsNU+xunpUKWfuQc
5H6VPy3oHG85dlQ9p/dHeYMlHJE22NsXPpzuBBcFGj2zAQwWXI1YCErv8c/B
3TjQKdoS1FT7XJR3hq1uZPMj0S9adoOxTmRs+bmfeNdjzeCBhj1xUS13Rz4V
oC2qCcqIFb63MNofpeJ68+5giyFe7UpoVCL2EXZ4B+abfRg1ZBHMhhbBSxfK
8ZsRwtXVs8o6KCrvWcyLYkFq6T4fWPJGozBG68o25nhSDquJq5gyVWX5Cl1H
E/z6ad5honC23nh9/6SHx39gmYsdN2ElYpVE9I23CRYHA9Mf5H9jEiVpEsxl
of3XBkBk/i0vjlSCq1sG2E5/+h25A641Hun+AbF5+AbpzKtDMuZcd1PCYRDX
bSe4s5DVPDD2w8tvUAIOH25NfhCs12B9RVWHFe2dGDCeKDUob6nn07Jocdqi
g2hgsnv5ZvCT7H1wUOy3UcJWF5IPNN5LUlDt/Pv90KQh2Lg1hagm8aDixkGW
hsXfoLJbL3FIA77Yn11bMnot4UNJhfGZX31UrQLmYDGwLgVClJvdW2c0H/4G
v8s0zS0vKqrfXlwGBPr4iq8ggRvQZWpUXX9pp8O15UH7uw8wkMp12HA13FkE
HKPeN35G3OcCxwopXtknxNWteyH17k25ayled0AYaN8/IMZZ+gItscoA/50a
fosJFXQv5jpI6RzsdIyto40mNsS6v9+hTxKU96axU/kb34RWun74HKkz5Z+R
BRDBrY0vD3QoWioj7VvmQm64GM5VcH4aax0DbhlEI05ZIcea1c5j7NCQee4i
8j+axycRY5UTZJnUstd/wFFtNuqrgePx5pMhb9PD9+FEfNeTZUQ2C3u9/ssE
XwvPKti//+0bXPTPWBBeat3C7gB6jgZ+VogUVdSOdL1bGZ89Bzfm38vqy62c
fmp1itesMp6Wte4DPs520XBnRlWS6r1eSKiWKRkNxaDB71eot70CcauTxWEX
QvUxJk/ZzlrShnyXAmJhfz5kQtXPGoZR8Am96WOy9F0togp78rR9a0MNh8+n
/pO6OcXthR6RUFWFZv8hGT2wmnVGMefJikdPTo64BO9bpUkXniS33cOI7eIj
z49iGaV1EAKSsccx99+0hkQ/Zmd7WOBBw9HQy8/3LL0jxrXTiVwymK3ohz6b
So1jAFdH4SSihOcQU5e+zmVPJ9V0MXXDtpzBNFH51g12Mtf6q9ZoOzXG6Ae5
lFgrWs5Aavr0KuNtm+I7O8TS3Qv1Q4205D7uWNdNdtvlA7TZYkVfvgb8N7Js
EYfVBr/BWxq9M5bd8kDq0jpTaoUPjgq5Gawpokb/aFJh4meBIYLowQgTrzbL
z50D3IhZKJGl6hK8pnBOL0Msx4bi1RMO26GenCSkwuvosGYUIR701APit6bE
+wMkcxL8Bx8LQRFgcUjEbNkw6nPE4rWqVIO31d6Z9AITGsN4qZveBkVVGu2A
uqrvvcbkBzbpfC/plkHNnD0KWW64iW4TqW9paN/iVcXAuzCncdCEjfEjoyT0
r9GFoFc/1pnxy36VEHBnyV0lJfqW3D/Ic5CtHa+0yj3d1VuYfT/1EyDBrxeL
KyWFt2qpeRw4URrcOQPk/+XNfcmYnp2Y2W0R5mAj+oitt5vrnmfZWyq+I8q0
/aWdx54l7PioHibaSGDj41mZs1fyrWMqZl11RPhpaxS1jT+qKl9tPbYf3GLs
81PBvH985UkxT7NJcf/0BjbgCO2V71OOXgsdEA5zPUTWaaFr0oi6ssYuBcdL
H/stEbGWbwK6k9hAqQs33EzRpfv42LHc8MqdVK7/djDgOCn1NS4ZNUJ+t1QX
B1MH/KJpFepErrI5CLHHxpITPZx0kxzELU16DQ6QdnpZin097PUUCRgsiW8C
EtsztNG0tKRDYZH+AnDhOH87BHM/wE3oZ5QJL91LE71p8ndogKk9a1Yx3zj7
M18GxasmeuyeGrAvFQJHIK0+mUmjI2lORQudz17ddILnnomBmmVdoHUdqyg0
D8NAijNpri/79zUooyvtPcbjsjcF9QjfD1+vTFeuHUWQGKl0At5n6KhJWsj6
Uo1g0scmjkRO62EHbaAFgkJl+745CG5CcTi1t/8PVE54J+ZnxkbX66cGzR9i
4e4BkIc/n2zZvX3YdeLV3av7EuzHR8kD0XpDJ6gI51Q6IYJOlC/kdMTKbLvH
ZMmxV1f1jMxgg5Xwy22xOfxGhJyY5RqHjIgMAHNiVKjCtpDjZrPIpJu/1oyn
gg4KjipXXbRBmupRw6y7MWYj+NZYk/icIwGiC5eG8Pn7AVve7d/cF/7nP/lI
SEaOI44TOk94mduNRolWRPONOsASseSdNYYAFlxb8/CczVdZa0mDkZnI8uQY
Ju9P7OsY98f0UuxKP3Kq/oOA4e4ghtruTDdjt1C0UJqNhIyobRpI6Qr8QMBs
rX4itkJLgeBwO+Vl8ubnsvf1F2xyEAYpuhWbvGFOiojiWflyh/bSJKoQAcWJ
5p0b2EjrL2mVFxW4c/BKVcDKOyNQUPqLUFvlXwe08JKsnU19Vm+2j8lzzE8Z
j1Ecc7yA3gnKhtZDynihWv+OEr3oGUMhAx0hSVIZKlMxR8XXKYSxTcjYFkIn
OYaHtiIW5h/5uXzY8QouIXHJN9k+2YXHplokelnavElRkuQE72pcxkaOqoDD
1HNlPBmBX5udCr9Dy35BXCFCc70tFGxwfypiFbdY8v56FXLpFBqELPMJqLXt
fFL5XMRfA+BedNXizT9u8lYc7kDN4B7nR6zgyL+jO33/yFgU8ImybojAeY9C
tM+xWDQxZ0Y0jJVwprWwqQRQQkS36VIZLiJb445JdqwWlLaUbH0fxEifqEYD
4Bs2camZ0OdeuW0uaMT/oGsj69yXJEcWAjxQrytcLLuALieo/UmTRtCnckjt
jDbuJiUOvBz9O5Hf+Cfi43i7cO96B/LCPM8uk+ZYl0EzymVv/b/SIpsmvSfX
KFhmnji175DuFCorvzvyL2P6pv9h+8odELvxgWW//SMIoli4iz4iPjc4CQs+
a7YSKM4WtPw7ZA6pEXCatDHhunMB2sPEUmUgOcnL8aItAMMLLHlQo5y9PrKl
NFjvHrVZhWV9Qr7CTod9QiSqSm9ULXyCRAIk+0utgfDoEjmq69Wud2Ewko+T
yf2JMMQ/J7MTYMgxXTS3zjWpiaDrfMjQBbp0Jgtj2Xo/g8CIHkY1XqNSOIvP
b32W5oPjJsqEh1b5BDD9pyUu5qoTft8rFrCqWFV4V9dQrnbhJ1/80L4QsL3Q
qRG/j8nReBZFqb1wqJOfsxUVlnAB4WUxkh6xjn3bzwf3KKhKyaPneqAWFtyn
RuH/36dTytGKvMGiFYz+VtUxEvFj0XvXZv5lcBDvTUwe2sAv8+zFZuAraTsB
Hj+jGx+KpjAWrvWuXx1Dzb7zTjuEdu1Yqh+8N3VCUvUgs036s2QMnHaMrmHl
Oes3hf2w+llHG3WqOaIcJtTFTRuBTY6TrAb5LWkW08Z0RD0czalSywMfDBWK
1An08oXsvBWRySnqYuiZx+xRS66RlO5/W4WZG67kJFV4WQF6izQcIjM0ycYX
ALbmUDp1f/NZZvEubYlTJA8bP1vzSAVlQ19mwStKKfY90aWoggQPMnMdDE0l
+a5iQclA1THxFzs/74rkrUXdzgdi0CLLa358P6VhmDQ42NofiNNeSI/3PyZe
21qA4eGpxyXJH0C2XIpPp4n3PSYiJgWHMmXuCJX4/PXhvmoLdzQRjkbhq25Z
N/jTl6hPV37mQEVQ4E2SUHu5g7TZLc1llqZnfm3Mn14Tr4n20SAZwtEn8KfD
opN2nLe86MuQ41UB1ykknBPkzUW/3knUtzN0oWaP3dzrBZqPPGXRyVp7HLNo
voyYp1DmAzn2MNUnwh32M3umh6Apm06CwE3O3Ii7elRqTSQZ5MA9m4PN0vwi
EDrLUulJLTawTylw8yRerAmTVaLsjNcnV11Yn7wkHzmHr8f8BY6avOfgECI+
TEzOj2aD+3pxJ2NMtA0RuvvRbOzJDZS3mHoyzbgGF+Hk4EoojfrkWG+Fwc9L
bmsISGw23InkUhRGVsYnI8rzWqzPo7UcjdRjlag7PgcEPErfLeCe1/5vu0qP
Ftf9sG9Jb9Zty0EvxBID3v/KxOQ0KvrzPe84HKnlYVMkE5gexkXLStOEgTML
5BPNbdseKnN/1gKhLfYKEHCWbHok6yJUzrZzalDNtGQR/rtxU+f6LOI8zILe
ldRAB/x8WP+D9zpE4lk69e4Oux9WOwCRMS9gJiLUNRTcaWTE1pDXD7HUULN0
L8Yc8ms3MhV+/pF3rRl3EeS0d3PJyCrH1cmVhWvmOu4c9QtbAJjFuge047IZ
LslZ2rSojXe8yy0anYBTRk9qc7YbKnhhHJTWd9ajz0CQyz6JfOeQ6j5hjy88
u/bcHQF/6Np38WzYNIbs2yNwCcmcMjJnZKqu3Rntpwrq6SWLKqR+5H8DUQ6j
XtGWALR+IPE5stZfnyb+9FdiWHpqZYM2jYBl2o2EFF4tSs6NpuaJw3suv26u
JEqcT/tHnlAklH/agC7TUkfFEBBIC6gJokJX6WP3D+9jgB7RUhetxWHP3MVd
s/25oMYHq4Q+Gj8TPY3gcdqgNXUpk4bFp3JQaOKn8LmT0mEZ3mIRnzvcUA8p
AQKTw/uqVNmJX+gr/FZaW5hZUc3AUNoahtwJpRgvqs27F3BGJKGd1ONIFg/4
Ul5r6r+wW6tP2T+RdAx7Mz5PxVszGuz237LhAJP4haVAibJKrPIYIkeeN+Cu
Ek0yHvJ/lTaPUrSo34nJgFNoeR+Y5V42EKRJvt+Np/hcGe0YcFjqNZWLpIV+
xDqH74MNZCJ1mArAyT1EDLMijdBJEu4Rq2LcwBbr9AoDv9BFTDxgA+Aj0w4x
eoMqlJxL0wZ8HwrEfTz/DdA+lPTMsx/9pIBHfi3qlLLlOWeOg/ERY0/4ZfXf
ykM3CA0UIk97BN0qQlNgXiNaQ2e5nOn3OhGHskUvZByx8rHAM5WXDgtY/VCO
sGB8kRaO4ITHO2rKHqdBsxyGfXZH2eqWk5gRnC8Z7bputRMTiXPhUWhth6Rw
FA3hu29r4mvai8ZLmWVnksKMjFodk/mZZ8e5VfWstg+2hu3qkgZ9MyHIqAXS
dlcaUw8ZlpXd8Zj7T0DeR5JX5tdnEhZ0r2H6weDElQqh0Xadl2MRYAUY54I7
W0mzJ/wUW7rcpqlnkKOlHR3R1ZUZVMW/5LpvcKTO9j5N9Y5wHD0v2RRcKTlx
r6xI0ywJMXUqPG8CtW1AznBu/qtQPBOZDPS+uSV2hK2/BHKKd/dl1Bu3397m
xdBvkh/5g17iBoGBE0zuCxrBGeSnYlfJeN+QLwpDJwpbBz2ZsKyN84JTXBcB
snf8SJtq+36Xyr0GIniXuAuh5UX9h3MgZRMh2fbEcxUiigFibb9dQ6vv/c3x
m89misKpy1ZKB9pqPD92cCibZVxOEMe9EuAUKH2gMtA/E4aVn74tKmWp3Mi9
seXEAHu1b6kKXzv7UciUwpYluStFmz6WBh1ePExmsENpIQkCVlGVA354WlHg
kr4SMIR+SRtNQyzsbC1Ki+P6lZx5IdEVWJ9upGX0FW+l2RjgTa2BD3EykXEh
wfSP+iDGur8hKjJBiuT0rvGLxWy3b1bRXGMsOsAfKrSU7QLOrOGfNK/8zoC/
cQAw7O9c1LgUGdQd/EYg69BG+gUhcUxtU8cI6VbT7xRVD2qJXQlq4gEF/kuK
jbQLZxpgr5K4Q4gQwNpe3YGnLzGk9vk23uI2wNdouh5JZS5WACp1MY85XM4S
UGIe4P8JhE8VQnNDYFcPMZN6WLtI5jCZgyiNNqSsvm6Nu58fL40XrHm0NFag
nnEToYlbPUktBAP/BwZQyBJmPYZqsyrKfWV4P8gZf1AYWIWuaXBmWzCd0dJ8
fmGP7eEpM6mhWEXPN/jQ9XaiUNMLbS/0N3ZBO2D0JDtR4h0iarBXh/dde7tl
Op4cyQpKiUXp5j9zcF23xJkFRhEquqS5i6f2hkIzE5syJ9NjDS71EIb/1H9A
TFegWbL2/xZVlzNIz2UT5C2lh1aWQFdd7XYPtzOhHw7vlwl+C+EzH5ug9Lbb
rJdhS8tgd0qWv8wq87EHH20RSv7Vn1ogg+izmmJxU9dV/TK8zPDnM05/84/G
XvGCpKFwwReIEAp/qh5onZj0fi1cUMpL1MRLb3KszjnVCJc/D+BfOLhljiF/
f8WnRpFJPefsNVnQfZ46SzT0YyMXsArg72JG8cn2SVyGJN3Jj0GcyXnScQhc
6PgDoU6Ao8Mp6oBCo6WIZPG5K+85C6XKQ6Bp77cW/IQII0KwmRJdlpL1xxax
/Okq221PhoUDk8VMH7C9aQRRt/YsUPPG4kP0hCbDndATR9/LaCaHBcMFX2a1
nJLa3OPzYeY2LtniDvIC4dLM4iHYTyn8CMmSQiOOh5S87OlngKAeY7+14UAb
d6n8LP2T13OAJR5quYR4uzVw1Q8/I5T5ZQwMSBOM0C2TnCYSlswJgHg5Kx3s
S6E11Pkp3lfbfnvYtdonNXzNF2oUVIhyVNF0dJMrIVLDy6EHK6cjF0nh8UGQ
w6gbaPFsu4tjENCMkfo0umZ5P3bfGUfdoHi3MlyxrWZWFbNJGrCgx3+5+WkJ
jpz8K7+uflB1bpj+sps0kluoyjHcUxf5fFC/AOjqZ640E9rB8Z5gNFMhCsj+
bkBnXhiEbnb6j01S2JsigjmtgTB9dUHli85hWra3P/6ZVczLYj+2I7AbdTcI
WU4WOVPEK9Pt+RuVUGD6uOVTBDa7SJsRuigA8lbON/k8Fng5OBIfW/gFOb1U
hRPADp9rF7qUylG34yzZTFqO4iw9qh1xqT8mnefNnJeMVoKH3sT0KnP/2dvn
ss2ahLtMRmPO7yg7kjkS6u1FClP/SZj7DrGsnxhHUTaa69NqpSnN7ULgkLWY
MO1pJgLhCQKRDxFZ1xMTdLd4jwpEEsiF9/Dpv8lTLyBDVDFBw4Q66PXkmiME
lKOCDoK3N7PEAN8saA8VtIEM8UPrY8Waqss2wvayaK0ia8qrteGd7ywQTbUu
gO20dS7khKXQQyRYl4h4eTnF0W6VFYhl5WjEMM7i4A/mXzGH/D7HOQViVXd8
jbUC1WVNUQyN+U71NqW9geL+QO4hAOyUhwKa6XWCocWtJD3WQeBLa+b1/wxK
9bZVgFiIFTgtijSOFdlxFhn8ABm4SVq92HkPWyGCl7LCpOSZuZJI9NwUL1uA
aeRFCPxU++WgZtZjOH62dMe7jqvC1PvynsjoLPUyqccTFJwUUhleanz6Gh2d
+PVlqeq1WHnKqOxz3EI/fh3nbkBYi5HdaCsNvkNyOuMTEgfH4Dr3fyA0nYUt
ycimcFvEES0KEFpP8eVievON2z9HyPTwJynhlNyK+HqZIQ3abGeeEW7TfJlI
T1By/PgEaewKQJUAKnehAz5FTeJtpegO+MdcgTOmTjrkc6sS0uSBvPMQnRHQ
mqSWMH/XuXMnBUKsGCMTEFZmTvOzsHwWgT7ArkFW1wr3qy1G8/7NrU0u8TSi
kZlHodC5rhryNfeZmSXGOf4z9TW8AiVTF16PdUqet3sxU1LlD225mDCyxu4Q
I+niQr4HohqaIs7VAPB6VJ9R+Yf8Y3G/64/3tuHhHAMzjPCpv6iEqCWpOBIp
y2gW7jL4rM360alxwjbq9W2JmqFb86jwanOYnH1Jg9e1k9L51kWOe4uWF1tZ
6vw+p7JjNICW4JAW0CY4qP/SovnLBifJPSDa6Q71QxUH1mkraiZpm5iM6DOh
R5GoMWmEwNU/GPFGmo+/wPHmHekAgKIqtvrjmRqv9T8MTYkovhsqZG70KTuf
pTdbZfKwpIPgroBACb920VsqOm4Y6y6VO5a7sAqjJrH8lVQuopWUuN4EM98T
8opOJ5n25OK6P4cc+L5mTQPr2kdAUPUI+1ri2bVR9ZKppDplvDi+LzyPKsff
JS8ZjYjwklLKihAWHXC+wKG+E3wN9tkF6+o0SltoR1KP00nTjSy5x46yRUgY
baKlz9l/gFYL16CPVd5dSDdmhZ3O8ouDoPQ2KMK/CBjSK9L68aIRo1h5cBWX
wz0p/SKcT0WrdZwyfLHzme4GF7HvLQEGeT2tbexGGV8KxQBEytZHySKF5sAR
K1OUWyTywtwh8SOcdZiCLPluonBomYH34tsUAqgPGvIrKtQR2EaRhPODrq5C
ru1dkCBcLhCxi2aw2NW9LQFGzGBJzag7dojYI0HeSCjbjf7SghKUKSOS+Vic
4eGn5Ld3hClceL/FmIayMIohIqv0/h4BMp6j6+mip+vJWCplYL05aVJSZrAg
jx2WMjlELofF3JR9dxPVbSYH5ntvRIhkgUQV1SE201vyVZPEHJ7wvMRNva79
HMmGJW8sd/JATUiSnMbKPbITfnycZmx2YCO92u5jKKnY9MnsKLjRr/xHD4x9
3UemzwCVjfJlCeTf8k/TDlcIQA/fOpguc+lzIOS8FrE9ADSM4QNzU/f1TsPa
rir4UYxcKYIB0OJuF+LJ0R8J9uz58+/a57oXDPqmNSBkGD90ws5It+UO+BUH
Yc1npj9IMPBfkSYeWjb4Zzgtj3CUi44p+iPoOG8snBBKgHE/jqPCHmqxiTd6
70m0hQYRhRj4RsEQclad5QRr2KuQxdho8rbU9NqZzJG1xroF/nCZivAVTWHH
L0zdsEDm8zWJJA9yf52KT5ytW1PLhsMYlR+50y10jC3RrQoHzkcv7TP9I75S
zWhd2ubL8Ce5nwzM7s116JcFVzxPQl1O8KLNhb/fgtVnUlU/Y7kO5bffsFjp
+wq9O1BAMtRu99Puip48HeGK/NSi6+W3gEa6XKzrIY6H9vgUAxaA+/SGxzv+
LSC7LYdIgqsr2lwUHBYIl+vMZc1pL2Dv1SrAqV0s+9ggviuAl3v/r8AiTLw0
zIJ2H0dY38Bwke5eNLQK4hZlD5XqtUKlQ6YAcBbw5o1iE2lha1p33SS8e7nh
nv2MH5MSAIgK+Hx3NnpZ/YBDU3jccCVkHMzMPvstnIq8OZJC7HmbinII58k4
yRLM+UEAX8NNOod1IamQyJ8DUqUufyzOi78h5DE2yqjnX6qzZlvJbEnxrmYf
WLUYT3XA/KqygwFXp2ENdo+CvZ0msY+BvfTkvgNYgrQW/dIs/HhMH1qjDWto
MZw0XqowEAXtAKI/CHcBSA/214n/6rM4zBGdPLVIwld8OL6JKyN9PtlO9r0V
Ae1bZqtXU47JwGmGsfMqmAp13Hh0h8F4vaucM5b2Cswl6zvZ0gihqt/0yW6A
LKnI8/3DbE8euLxY6DQKLhTL3VaD1NQrfMESGoeXirBCsBLygLADP9RrBqMO
ROCwxUGjciFYlni49x5+5obwjn+zIhuTeoRCRqIO5WptqjQHTGV5wL15d7/s
Y0ZYUz5+HTzjBHWXdQ2ganQ8UK3yZ8xSpM85o5MsEnRqWRplQ2YCxAhVjbwx
F4lSzVs9D1GUXs83W9LhQhmqKb5L4ro3O5Ru/rktBKDTCMNVfkKlQ8Fo6p8R
jRuWd0owMp5vs/52KsUtnuyJl35FFCfqOzXy+YMkeRJX/K4zkTbqW1QAyk9z
R+n6IQ4HxIH9eBJDw1vCyzd+evTma3WCbkYg1ZGMdLdLZUuiC8xCaewZYRmN
BSnx79KcZlhe4VxRXZqZECLInQEQWB5qN7aCgHwRm7tTN6CNLBhVN0jiTkWy
K8DmnHPo/ScoWit4XrPXtMe9corphqL9ChdTpNKxovCbnFJqgJ8fMkYzC0jy
/rz2Ac8aZWMrtvdHjAnfHMGYkY6Llz8jtdYKa9RaeemsDLalQLiKuewuDhi5
uqELYxKPCVYTtNBa7H5aH0r4uPLb+BRUXi01G+eCkNOvS9sEDJe7iZtG66SC
Mup7Kd4NWEx3cNxbddkDePZ7RZZeNmAKZWU4KbZx++8QvNXPKT+E1O1Jgffj
HMe1FKuF4/mHvHHw0u2Z+PKfnhkNNU+ykq50y5Yn37l//7G0UArXy4jk/kjY
1/YqkvcDOuJP9Lemoe7lPqOzY7nWHunBxe+zswMrTFzPOC3Kop8ecwCi4b3p
wGqWWbbv0YdP6kVLeQ+DOdV1g4HWij35cXKZjX6hvqJFzg9YRNowX4GMrlxw
exvV+UgLDUXR+Q0jLfO22TocKDtW6CH1eT5FZ24WqoZZOs/7gBRdQR4M1LCx
J10dA/NI/yMcYfxX9ICU+kzbvJvcREK335mTBAMwCc6JIRbxJZzUjaEeDknt
e/iIXKTox8aK0YsO8bdRC7f6ngBbV5B66HAnJwRVihpYK2iatA8C4q6ykAYH
311ROH3Fxb6XSxxqueuoWiP/Fry1FDdAVxDIc+4pYxaz2yxaZd4PGiVUDwRO
3upjeJ4CrPgQ5M8Asd830Ljnx4Pdf+FQFuHVgtDlXYTYOJnniKQFfm04u60p
ZDYX7pDkIl8F3kzPDMVVOT17DsK11M47Kb/piszWVuolYTzWLw4Jq4Rbx1eo
7lTb150WausaOcZyzj9NcI5OsH5PqaQ9H+dRXUFYJTp0m+19RG3+OWusqEcy
P4QhMG6EfgAtXtnrYYczTWIzyoP8fs1UdSIxU2lW1Ptn3HpeaNYQANd0l41c
9KPYEkKxTOaFWa/1j7VdZ/2qZFVqFRdcr/4zkNPgSyGKbD1RkE8KzNvX5JTm
TNis+f+/hDGwXTQD6CfPhmxhkOOW1HrJAM5dIgICnks7M0rRSUWhTKpS9kF+
QcksZaEwO/UQj/REscuYZxJEJC3kZQIf39JiY1F9LC34EmPhowg5L9lTRGIl
7g9KIts/+dKZsvKkp4vcE8KajXZf8XcFikSTIkLW/u/1XLUN/MY+iGX7UMlP
HCqiZEuXB0ynLXyG0AS00EJ7AfNOlMBb15IFCceaBn8PcfMXVYTmU/wAaH1W
6gkhgGCMdv891Lp8R0KRHZrZEJbyY1TnUccxsg5/Cj9IZRdTgnHQioswxEIB
XjniKP3YTn0G0ZAfnIxZAROCvWgQfqbe3IgkuRNnscLRqBrRjjfYT9XWeGr8
oPGFleLEyvcTE85ETgzGW7j2R5UbIRZdIaROT9duNksH1rI96Q97sjBBaYy1
mwKATdVhl0AbmPxzkfl9nua9TctAQvmc/9qA7mAVxtlDjjSnSy63pLJuNvXZ
HWjFWskv951t2gM02URwzbE/JVWGZ0g+Z29iV3qCKvbcRnqkpTIyi4UpV8sK
CkIQZUg+KLWUY0gQHz3aAFxr2JzovkPtbX1kzzYfeGmesDbqujqXNvAFPrtX
MKgzx5OCRRgu0TKdu28ai21gX5aXm0enVdt9HV2yiHoH7a847SSbntvlqA0O
J1OV5XZG/iyJP24oXUjA7IXHaJFsVVaJLGlKkANOa0hIzPK89pzcd1+1/Mvg
Uuirdu+9fBoB+7fAo6uiT2/Ryo+jtc8K0CegHFTRH20RoOkWmjtgo2Y+05+Z
Phs92N1ACjNl6GnEdeG31O9HHKHgJunatfwX54Ngob+uY/j6PITgPuPAZuvG
wm/zkpB5oX3QtULwOOjvettsIsLmKyllSnWFyNlv2uktHggTTEQ27OXZGkh5
QmxzkhVvq7yhLQQP8u0SrJ4t6Tc4Tx7MJEucB04o5AMJEIzx0e2hnZpoMVTT
BeLSCmqATFekZuA11tKF85HYkPb41JZp5AC3WbNldlqcE5ybf846hBi90/3n
99lJO8Yw77mkpK6SVuQzzEuvNLAysMaLR1zQMLEqkpFyhBle5Kfoc47zgOco
nPmxpi5SFtX/5JYpMm1S/QoGSeW0hO+qcjHPIXUJdKfsETmAW6rU1CGfAwTa
KnpvJusOLEQ7hUi4CO8KnDF+MJLq9YlxrMNENW7gqLO1t0zxPNRmYEjPeoI/
0FFfDtZ2LgVYUpmlvpxecIWrvx4rSGHCmMhidj4If5dsabV1O8uezxrj8yzJ
ff332gPb3IeY/A9/aGJmbQxNycy5oAbiCrYJNy7wdBmv5+cJvPAcuAz72EYf
6wEHVceEVZXcQPVd/fZsn3Qtec3KftS7K+tDoyDltsbBqMTw3vAuroNvyv0M
9t7NGFoU5C0yqTVDF9OCLLOuHg53ZhoBHjHz7vy87TquSMbWvrcP03XkV7ts
4Pymm4XK2VFV/eXJFY2jMb1vMgXcldKbTahLE6hajNtOCub8K+Eg2P0uTj3g
7HY3ikKSJC60BUxdrgFduoMj3LJbbT/NhUFuRuREqPe+jYW6mEunGeTBEo9W
gRB01u+pDQEKEPe1kfMZeGN01eit1LSMwXc8OFDu4krC7lE6advaZgRQ5a61
xDrkSFln57B7ZPsiavQ7jqPgsI5zqtsuFVKjHBfdMl2eQhcO9U2cN0wnPuJc
47eYr1QdJY+AW9ImciK1ENjTaCboo0d8Kdl/o7WvbEjct2siSrzv7gsNFjJz
OKDcZNiJkvf613W+wWZZa4kKxcokoGzw0TPLrtH91QJmq5u28TPDuce1BoCK
UEupEbuLEUWvqeBLm9KQYL0iOsja/symZfwFGBL9kAEPBrIu0wXJEU+wSgqr
5QmQxSzPVwCuiU2fpL8k5Xbl7nbYfg5zJgSzitBQYyInyTMebDz999xeOafu
zKvjxBfplcPEXTyj4IcmtnUBUeSmJv9wTbjHOq/1iBojpQx3g+RVLEmYcwMk
oe28pjxsa6l2R6g2GWTxXrh2O/QetF3Yff+mLp1Ha6WOEF0jQggaqrttiJl4
/DokePBl5Yty0FqnX5e3DDq+M9i9b7fDyql2SmeNE6xc9dl5oWR/NU2GdPbu
bZl13+DstzHeud6HE9SSM+QfK0wRoq25d0Oo7M3cMm5rxoLBg2fzbexpIA/W
9e+kf2gxZUhIdHp9curVPzWBaYV0WjI+bGLOXJ56+gLGZmEwRVEb/O8h8KBt
9aeE/vnATfd/SWrCGLpmk1YXSvsG5vbZdoCI7jcZmaUI2JxYTIDSRQjgKJ9L
xjFjpYE+AcDVGTNgouAu/lIlMJ/oKkIGzBVH+CyEBelqpnAPcwHVuaWimwjW
cj+RlVjEV0xlmv7ze642KES4FPBX9IM9GFJ197jY3/PkN5TYnZ6yHQS3qe7Q
scchg/Z/s7qzPnz3ZAKEx9cpWdrbW/4QDlBJbCKuMKwP+VkSj7iHoq9UBMXs
sfGNzbkbk3+OpZE6t0NPhzCOy5E6nji/HdD6WMZOljksCgo/7g7OV9Sb1vqT
Sb6Yi9DZN9T5cxHd63VuQZiwt1cvtR+xK9ys94YjhV4MBZCt2lFE+cBl6PB9
4mdNpLrk3D1QROWMmZdMVf0puCZsI8mJ0lJ8gvPLKUki4jo/pKYfHIMRhWTr
M5q/ICWtgkKlT3RX/GiykiKfxcRIZYBC5gDzJp72CZllMeMw54fTlwB7OCVH
e8kQOio72CDqLNVj1HMF2qhcmXfjpTYM99+6AI2fS6f3qEzeLxB6NP9a3Q9k
FIc13h2RvDodld57rgQye6MNbURvfjTj9aMAwbUPjmGHwuhOb/5C39XtSFtb
kr/x3mBbQeDSQehcNhxpblsTtulMyrmXK3xota5CoHd7Wr4+j5MkFL3/HD7c
S89k10waoQJD4yNLEFi0PTPBFzuKRcXMXoa0GC+Owtg4gk6jPBeNLLUjw8t+
CvoVZiOPY5VyeCfXWBoagwHg23coVjt5KhFTLQBVU5G/NV0/9YjArCQLsym4
ULxgnB9HIebOly/F+TXUAe/fzNKkZkCJkMjN7fJv3rSsuSwGNAGUG1Pdih2W
nrKu7ainwGHLXDGrD8NSv/ZaTYzAH0H0TxFNcGiObUpzUscaNyO2G9kPFtlD
eFAHi95oZAclywlY7awNoc4umOnZeW+Yc67sJkDPyd57rT5u5bm7LS1FmiI2
LbpDakqxav8nmHqaUe6i95ZTo6eZ9X/mq24nq0anexPJn6j5S9cjEuG07mck
8Pxp1mORUjvWKl9OW1LskqqlRjIYnCru9GfqxFI1dAYoUEMHLwS1r86oh76c
0McACZiLBgnoS6YxpYgkD4ZEivaT0LD9eSJeChMIYHONXs0U7fuS25hBS/+b
tk0C3l4d6LqzAUkRLF7nz90b9KeT9jQIHmHqekolI94JZuZhoRlMSOhsPtXI
va57QJZFM63vkuX4uNr+m2d+E6NADhs2sAJpotdSOEMaCyY6nRNlKvaCwV1e
A87aramCBTij7WgQonmvVQk3YjZKtJlQPWMP/g4H3NujFgKy8cUJYAjvV+Cn
J935JzxD1FG6CT9p3Pq+SvnPaBs2lnRlhGFDwZd38Gzbg0NCJOkhzokZ5Q3o
7JHAfzEicshTWykASg5jORLbitD6S2mJWzJaKZ6SjB+DgGE0klKrFxl9cdM0
CxuVI2+DBsa2fXaqX3xyUe11CZmuluIo0VHLcVg6VSPhJjq2eI83tED+G1Ls
0EZqjUdIFKg23T7MoKVTaAuzz++1dkBDu7QjswROsysaDF7HEPvMQmyh5OaG
/yIMjj6db9oiZw9TslJv2MZ4BJNAlFru0Urp8r/25h0o7lm71y5wNXSHGm7W
wW3HaJ1tKOYdo7RBXLXoux4hCgi7rn74k1pKJM9fF8M/LlN4Ph1IPp11IzjH
BciMpYhsRdgjBZLSzajxZbdtFvb4mbLSnhSnoC6irFlAX5JSBBeh3sVrHJEi
eYtOAV1JKMIlpoDd78TMU64ifsrefrkY2iM7dbmwhctEpRcH3MTB83WRhalw
QMn+oRvZgeRnklXS0yXvZ220mq+rc1N+YvEeVVDgZdpnu4B0gHPWkl4jZC86
IIxMPCNaGeZm8Mnms1w3i0doTaLMjuCxl38xYU5JuW0ILVszMU0MtPSBguSc
GbbacBg6n43hWYg/V9eAvtfWJsZY3y3/LFtbR+B6K/7fRCQHwPdlFEBmHECP
dN8fMpHR4nKVSP24ryVec6GvZG7haiEWWMVssgjnVyQKaa2oYdIbIHnFe9Uj
+3+/gDo+PwXJNHfXQtGlD0oTgbnGuI3jdcCdTXGyKIY/xS1052yflbL1BIO1
pF1GPXqL1YGkV0Vv+FyhzdjxNAorjoI5s8GP48JKBUBPF3PHM7Bhdz10Jrqq
LyHELZt3AOvCuTifXAKnHtEckgSgFR7JAup1Nv1L4lmRKFOYtAZq+j45KGJ5
2E93JCG5JmZssFm4zrcOiZTyW2CbK7FaMnHidu3lGQDISvSLTz5DcNVAdO5A
e/UI7O66sxOeJlfT+NYKRFqY1xXj2/7YVr9d/t4aAs1z5bHjQipjy5x+8uuq
eqGgJu45wVfiHzZWJ5vKiqQUlVj11RvuiWhQqWruLFNGUnvZ/MHhUOa7VTQ3
4H2Xzh+/uBzsnTum6Y+1r1yUUn0TYJQeR3SevGgVrGo3xNBEeoKuXim/OwE/
Is2pBEDa9n6txVVQSiFiJVRg/01IF0oBeI+i1Z6PHuXqIVzp1Zxp4OzOcFft
g4yZa74b+YIAF+XqYd4SClzRShCxdAKmnRhEmpg++PI04JEBCEb7NWexnYP0
gA/nPdznlf4wZLegqJJK5MrP33gQnQeSxMIw7hWIDTULMkEY3wqQVxyAJgUo
lzjs35e+EBk0aFFHpUJ+3gHwybgmhxHRZdAnQoXdfYqKiDe7zTQWpkTC+onn
KqanXgmOoxyinzkDMye/CLcUKihX/fRMY+xbwU+w9x1rjpZYf0yRxrrX8rLw
Ch9zvOMEtzN8aFJ50uwgnCXPhULfEaQik8n6YkzgM1syxsBo2AjQ4mvUYxW+
8PZ5UebouI7F3GOvuOP630/FgkGzUR4ofUDqjqfD07G6xg20MaVlJ2H1kJG7
fQeZw5RFz2VYZ3Q6lvHxB+FffKVxt6GH/PbpvWRXi3e3b9NAe6XDzfX0xlp+
w4Cs0IFKQea8qg9OgA3XMfBAsAsHXcrbCiSyjCZ64TDknU4c/GmQkAjjYfRc
IbPc3sWkwKlKEJZgx0y5W6iJUYZ20KO/3pQd07qqSPzgCo5uNZF59x/xxiOK
ek03SFqF31s0RRLxfRo5cx/hIEnel7vFllmVJRJgbTq+6hYDiQa60lAXSPBo
A9AsZ/mqiMLf7mygIHrNY5Givkb7GFox5z/jg8CAG7WUGGwmBtDYaoo+DWHl
NB4jcIY1/P8R5MejmoJEE4Tn8SpYgO04MOPO0edN0sHti4/YaZ1jSOTBMDQM
D7MmLCyCcm9KORrPjh00Jl/75Ur2aZj6kFl+YDzIAF7WQP0KCnWZNXwqCOBg
QgAqsiD/Q4/nMvCOgkXw6DMc/KiwSSsEW1QSXA8JELmAs+D5vi2OnWdmMLDs
GIt2Z3wgErxbuLZLJHM6juCuL9KzZKHDhWcqxQOdGGjximx7z76yBprmCQcb
vJPIEa6i1CUVpuFbDZAK1odJKsm8L5xQtLt/yfTSrLUg1J3fj5yTPkulLs5N
et+Tf/MLT63VTBpdnWMZ6fKZz65Ecd88qgOQ6nE0ioOLJGwsO0dcauF1jM/i
yjMT7ROnd3fUkb/PHeQoIEtzA/N99bD8htJqj3zAqUHW7AqCuimT3WbXWIiK
+aAFuQiwZ1scVW4WtCtk1oWqacdzYobfcpUQdhd9PX57RWRLGxAn2rgwELb6
zkDTVqWKQr+IEguQzPzUP3yEbBs3U+0+KTzNsn6yGnP5qORqVHd82SPiO9bM
nn4igb/31w/UyFVepFpr7q+8RlmeDNm2VXUgbnHp5mkXF5d51bZ6wG2pVgvX
Yw6a3XKIvZvvt1vEIJ/i4TVf0DJ4K3MUNwbGQLMQDfKPO6ZGyCFHnR1X91t8
LCbgEeKC/nlAK5RC04rKoERTjfmPPVVqzv0j6BNXAHJC7dUqAOoSC1zjb0Al
jK0dFstZVntVVScMeRXFO0SbabvTxm/g1CN8WPTI69Sp9IKLCvXmho7WiDFX
wqChZM9qD+ynQD9/yyMh6wmRSGw1NUDYjRAvO1V/Y14qYlj8lF5hivd1hXh8
rFTYsLr9SFBh3Lf14BllYD5jXcUw6zyquKaFso5D/cGEHDj+1Hg+CsMRw++g
p8844EndVNp1PxPBa6/XwlIne31AWO4+3cUlGm9dF4i4llxpWgyaxsxt1ORV
be8G/iAyNA0XCcMQABlVaxsZV6IIPyVT4XM7WvxRLrChWxBOpinRd30ire0j
RWpk5YNQplDtxXXHUbj+23V9wtkcECcWkHUzOQaG19Gl84lHfwaT2Uqdm/5C
mdvmnTA9dtCkUheAT+1lh6OkTtCLG0yc8F/4nkfuW6EzDRRt8R92n3+UaYtC
HA+pZnjK1zaayei9Iz+k7X5ax5uLuTTqW+GSxjfeTo4v4xPEVL845DEh4pi9
AW4GIl48NQFAuJscxwbzOGoAC6RTNfaGT6Ef+grqO6HCLcrfQCRz0Ff2Gxw2
A19eaFs2mk1SzRHC2Wh8rrNirh897do6UROzhPn+Arvf8qhCGGHpXAjsGhYF
Kq/Cw6lEbdFzBoBDQMOx620nYWT/s2yLm8zYtyC1DGKcIaMLm6ieG03hmUil
Z656douTrkNiU0D44DlcOxDk6xpfL3jlQf5RrRvg8abJo/Bk/mnkgPOCEMe6
KrVEhRt6c1lbFw+5UrGwQdHd2hvtKGgQDGbYBWVh9eBPHOuJvXCpZquP9Nw0
0ooaPnk0uq8FBoMNMxam2kHM5ZzAzy+Hu2F7iVW/4DqFcDnZyltQZrzSrvhl
uBNgYsnxG1Nys9Hm9xUwhdVi4eKk6qrGdka7HwtKyUeN1hlfpVnZTEuPgPoj
0m6sRo2diLG1qQo6Eqmp9AYrV4r2CvfphAHtT97sahAyYO3jBFjAZi8pc6nN
HXcOUWxAFT4Y0k1bvnyuiDjHcuGVKvstJtNwfpBLevsRIjcd2X0M23iV5kCr
BL9EkMG+5qVXACyCN4yw6KBbdRHpppUFm3K9S/oPRqAtyFuI1CqcW7uIoYd6
9ULECLpo9TfvdyMSUaNropnhrb8J+2bFeyJRE1JdGFpBZTK2Eo013TOtiBvP
OKevMghheOhJ9n+MugIYBtad7CvMRdP+Yjq3VoJ+aZD6vXCYvIbvqW/Fz/xN
q8W3knaLLe8fGL1hKEWJznso46QmuKOFY124trTQkmjiVoHvPBw+ak8RcG5l
aeXPSQkOyDA7y9IG2V7TkdGMjRaUrqI6l3vH6y+q03OkgAFVg661wFJCUZi8
AqYfnfQBDb4llw6BNJHsdy4rRXHC3m3DhP6aB4n2zvw1jnvGkRYwcEabddoZ
PgY4aoMBxiiUSj0JnuEZRcJdJBeC/4etS9BdxtHzYJ2NqlhHt70Mu/699HGR
7uIX9Y8HM69Jwo0TP3EFbC3LWlZboYpFymvyiVaO10LLYYAVuGR761eNwACp
r4wCexjrMpHaXIrPmvvexMqOe2/zsRpIWo1QilfRRX5d0u0XfI/Q+wlQC0nc
mA7vRqjehsyiTBa70175NC5M1NIwpH5UXT8SPqxOmJeTFaBoUsFoCc47wbmP
618U2L+PSHR0AvfBtqntyrZVsUNYfuLDx+lnks3UIg9GUAR7q9fOd0eLW/o3
rgXpy+8S3l5pUh/Za0oxrHvDF0ug0AD8MIa9bHysyEM2ClHdIiv5p8Utr9sB
iow1OEtxO4+8+s047JR9qGOAvcNt/TJ7MORaP1FhJk4WLKNqeyebCyeMFIcm
v4yJLMcs8JZ2dl3XvSksQ6f1vd8AVexd+RNJS/jy5iffN2+rLy6uIpPEKfZR
bfq601h4nT0Axv8JL5BeuPing3iVCIXjsnAvHSup33Sgdqr+MYStmfmlc4uZ
fV1KB2P3X361oHL6e81RlGePyAdf87TBzwUCNsgK3//avIQuLnAj3OcZOG2n
BJB5pThWWy4EwG/LJbdDaqeYYkNUwvU74WgtzTUNdV7qsoOotckJE2Ectt9F
zC0wLQ2r6j232o7jHbqVMky1ztT6dWdAGG7vb3+NQX+iXoMvq9+1i0LJz2c8
XroXyTWe62aJe6uJMQA6bAqRnSQjKh+bIzYzFcv/vZqQGWhvJzCF2sprx/W/
wsMSCb9jQWI5dWndXp688SKe4gX+ccbArAwFJlVa1p4lHFaeopN95rf5lxCs
Qae8MpRY5laW8zRRQ4wHrbdyoalSVnircaq5dI308d+6Hqaz3pgk9fBOWrhA
fo8mmAwFvO3GPihX+fICf64yXXuyoBuNx530xHz5arhCfHHsYi/UJGmevpmI
scna6egyFtUcw5sMgnZAE+PAODBAAejUwsuLbzdpznagLhXYggHQKNxc2Cxu
61TPwA1aWuw2sDlpuGmdFPdbsQZ6rFsGov/xJh2sZ/mgyB4exceHRt3ZHhFR
9n7ueMRoREicbpGqHQh0sdgs8+GtTnJXR4wHCSNXvBSraRzYyyesbSZVY2sj
1+NtiZu1yXKDoSq5rmF/0HcDXNqsdKZfVGJKuqjuSBgw4t5mHVB3Gv3RFohw
vHOzRb8F0zgugjqW6fx41kDcB8XRlQCzNVkS/sKbD/VhZA7qSHrv60byoYuq
ewWDcyiFSlmT5qp2hZBvzSEJFZMTVJfmSia3jr2tnGKGXcACg1089vsRepn2
tsyI6XrDnFTwzh5ZQXxK+G4bPCWBZbHtFuvfigVDIBrh3ekbgkOr9Fk0p8yh
lNZo+fJqec6RT9coV5lquKJwq7DePKOtWhqHZzpYrsczsSMpgW0fKC9dxoCk
2E/iTg/wd4GVyXRxwp0RtUJ9/E34h3IWhpsmjzmxTVYY6fUhVXbPFDmVQSmr
GuelTdsfImrjS1DSs5kAHf3kDwXsbqBJ1a90XSlTJtQFBV7j0KQCxX+V21eZ
A27IPszwi+Up/OZyBHAlCuG+gGi2xVYDMEk42NoVMdDgvmqzA22dfJDtALuY
1yuCFMbp5qLjXlu2aZlPcoxFOwC7F7PEuo6e17uKBfUXgZYRwa4QCBDggzXP
ehVkzoHenRsS4xHIcCwSuVew0o6GKx3kyZ4YSWPFXBS4KqwI5afuybskOzX8
Ayr9mphlVeS4AW7ORg5zHbuKvJy6OI/yiOv6/da3OvC97aFFvuRI3qs0i5H8
pL9XRfdR1EeKut7c4Ed1mvLzun2dVrOyVXnHFjcf4G7bSl5h5u72KHdmY297
gUkQJf/WQCJFV41lrBWCFpZeXQ6p9CW9n/rFlGgHqM5oUoDctbnQkCCvRcsc
bgk5eWhBTKAbF+tcinWDg0Kql2AoN8zmwrLPHGZDHVO9YHygX7CubPgebh9D
7Yp1uOJaEj9Q5mhcSLduXHcIOQgcLUACHjfG8GgO7MeA8PxzyBvX/ZKNHQ52
r16i2cghVT+q93M6McuKa1dYAZuklqCfzf161ZuLmXT9NqhJYnHK86BuRMVA
GEMo6M3JKrG7Igsnkow1LeGSSY/T5Vh746jzj5+9Wq61DRvAKrLO/wy5ZUeE
50hLXa/OOM4aK5o2fsGbk9sKEzDl+ODrzJH4ZNbQy9fAKEUmK5FhyLx5RaVY
59LIKWa/c0GaEInkIERQF+Y8y8I6Tp+fJROHhx+2kzmRIo2e/ZW32HjY6iFV
Oh319WzLGWCMQa3kdtuswH1ERVHPfvPay5SKku9bYsXJfSVn2c2B/VfPdaSC
CdGClAT7myfqSHRv83MIKgBkHDmFnxTJFHNCdBIIka05DE1NVLF3CBls22mY
AqXxu0QBEJ2RYlBW/LfyYIbvivsZGIN8VwB54HyNFNsjFSxAfeTjNt2r7r52
8PSt4Q0d5tXz0B4L9JhO75tr9EebSGlCF0Mg7uqAeyTzZ38HkuQoAW38AbOb
3lO+DoRDSLjCu9H4jOCWKH+OlRj1qBsh59VlswO38Q4N/pRk7maKrrnt0tZz
QzsGaFSIJAlgL3Oo/FfTOCqeemIpq1bTqW1G3ICoyEfnaboJi32s7ep3/t6G
rMU9zGj14fQKCj2H27nBxQDVP3Yvgzrq73Fj/iytJH2EVhnh98USDS3O+LeC
zK2LKEgko5xvzeROZKtDGe0sMZqG9Ii+G2I44dLNJGqWd6e0GQU1+fuyboV/
TEKNrC+HXho0/2en3CIkX5ZgC0GhunanvUSGoC7k7+aPk2CvtVI3L75ImVRm
H2YpXQ2Q+naweDaXilDnNNaWfXK0E0W5OTZXKzRViPHjuIgmCnturFY4vgNp
797HbSi/O651ebTX0kBAJCEve6PjA7l3lNTwjid5kPct2B9/eKQV9PrvSes5
GEDxXJYLwRW6ae5qijPMhBmvZ+tEoV3JXS5LwNRh9LdC6Jn0dbnbB/cBP5j8
ospPCjSIbSmnsHGMknX8dEahQ1ovk+l38cRDitm2w/bgP4G6Ckp3DAHKKggJ
fdDC9IhYYaYjv6jutdcf+tXxhtl9eXb6p9CFO1O3ahzAF6qOVYMwqtiZXSk1
VLtRCy9gF2CjgyxJXErV/wnvjdtsd3YVqiX4tkKDk7qYhQuzgiAc3+m/AdMe
//E1y3vJcsl8v8IEX9+K7/hvhGQV1c1Dn1KljszPKLEvKo28XWkHCZ84TzLj
zu15ZfIBckTZPXFeevuRYwOU/atbIB7dJynRslwIPCUspBKU6TBzoq6clHbR
JeLTl/eHzXvabYzR5RLFhy1+F1BurYUsbX+PEuJbOXO/O3ZGLRzl5WuACbeB
XxQDHncJmI+u8E1cRAB50MBpE99s/5hZQxWQUmA/seXg8+l3frLCglY0luC6
EBvY66xdsSK7sRm4ItVasLnCOiWdXhku24gZPr1H7vuVaFYi2lTVt/2xvCkz
pmoSy7uDpJ5JMdS0MRK8FIGKDwRfsUut7wRh/iUCZssZQSmaRCQ/xWvsyCGG
xU+GNilAILnROavW4hLnvuPaGzRLMjczPCOP+RYKL7yRdLfuXywUXmafhccZ
qLbzqz54EV2MBIeebTf95VObW16ZKaW8Y5lu0jozHK39nSaLNqpljT8JsJ/6
YPZiwapCWrRjvUrsU45/sM8S5VA2ATO/j3m1YrEnGZ1Ez5PhL9z0W++w//nG
5LNlQw8mgQEhvD/ZcZZ99tLKIsk5bHH4ju7N7JRpyRckdzq/CFriw8euH7r/
1Wq2gDg03QWJbvHSq2Hiu+psxQEJHa6deOT6HYtoWK8bkKnmujsW481gZR1V
IX7ngYepU0zHmpfae0fDIoC9I2liV5MnKsXjqCSNDrJXmetH1ftPfCR3GO5k
ibofO8gW9oxkk0eDXojg9T+AqmcefaOeopNq7gkQ3Q/aIgcdPgpzXUvfd3he
Yaelh9F7CoZjEmzdJL0t3F+4fyhP6RLY0mPiTHIAMhVrLYtz5Rd/86IweAT3
RW6XG/i0WrjhlTM7TJ9aibNJkuhWxuhz+JisR6/yWGvY70ci+LIzOxrBSVMd
OIFEWGt8/QkY+tZw6/U4UwAGjY69ECQXcVsXp3zyzmWmWQOfNgPyqpoIZrYd
2d8U/r21TZFKU6Tb4WZQgXjIHv/z1tTwIxzehjeIx5ocw+rrO6PwE8dhBujn
614zvZWgPLVPPh/C8BUs0X1pdlx3bSDsZ3SIud4C7l69zJDw+8/13ywHTBWX
YTRgVqcHpyK+nsuvMkL96Gt4lE7Ty5oiyLQ699nD3b7CB6DV+J2k6q/8eXPI
5YPU4khq4DBmdrcQgL94JjpQxcA3DMcGj65I6vFweCybeGfIlGYvwcatlWbX
jfKBLfj4khsRQ5gh/MzK/Qc5D9c1+/jZ9xubgz0GGBfoazmFsYb6bNLUv6uv
s4HLgG/RIGiWGWcMrZZNEkdrvPQ0333Kr+2EZ/LTp3nz92e0eKBSrinpPzZs
8Dp77CTX0KDl3ZWasRqI59EGjw+7EdlK3fGiAQ95U2UR0JIunTzOAwGVsrIb
Miy+IGwB3T1oEDTzyRHy3s+2OO6HFV0LUDP3IE7d2ZjR4oxrZgCJw9zcq6A+
1X0XB4mEaseyLYbZrYNWuZtDL3EsA9snSJv1HpDL47ZupTw+ikWQcpmOuoEQ
Rdm795er3WjudBkGpPybVbQuj43TEQdNAFPqjvxuCPrnrQarP3CL8FQZOK9u
x3gE7N39Xvar11m/qpvYa2VnXggrC3pbib2LcAkx+91xAPJiw0SSckL0W3V3
yrJA2Z8p1SQVY2HabZkW8OuNEAFbmltvmuhDHmLO186xp/PwYDevRYRq+CU4
7gBFhVJBiroKjCZUZX5GRkv2HNHlvODPr1cNLoFZtenvlBn1N8sBPZWA1fha
IrY/ResuIxeNvTImKXE1bA0mEQIVDT0ahKjOM5o+Pdqj66MHsBjNK1fw5VZv
qxhzvS8j37BPFORx1G+aA/w0Kifzg68FpIYFfGSvffaGFbzpV5R6THj7hiMb
sg3IawFaOhZAqR3t0eQpII2mlpTOkxCfLuWpK45vc5QTIeTNsx6kRphjik10
VBdKMBYv48WQ82SYqA2I1rU9dwUNrBCSEPJpE+AMi/vPkJlFP1bzie7Rt9yd
Af1QXYtsWyrXH5FqW3Kzxjm1QQNsy1xrlK+NHoBqYBEI+eWlG8DrfQ3M7xkx
LZj/1fuYZtuWXyD4C81CZtQVIV/Tjy5cqKv++BHcAGiDPoBOW+vNpcBVvnCr
SyfOIAmAMww+Qz/FPt4G5XtUizy2tJa5nWkB+sx2ixjEWpMAp0GObV7iCLym
57Ve1xRsY+9bNabmtDXC2NJ2W1kORjq9k9k2PsmCV+qKoLvElSH/3X8SliAd
CQW9ECtL15wzQ3o2mE0qUhXrWM7nKMhh0kYSe7QmLK6HQPeAiaX8nnXhug3V
ir/rSaB4HauWeW++5kNSHfh0uhCdfec4+oasxUortUck/J3u/9UeNSzItOoh
h0zbOYV5DMMa0DkoRyPjIm9kH/ezDfpI1WYhu/1lhshadB27HPVbWgWAJ1kT
+1DAY+O/3xmBbB/+DKy52v3GfQnR+8NkIPvfcn64zPlo73GrAP5nEluLXy8D
FOdpMr8CMEyPcbtwrM9xJnB60rx6uTIXLycUWrdl1fcvqRmWBVPshaDAxJMq
IYTNFFEYu5E/iiO678EeF2EqvMuY+tbt3PxxjgecK+ezuKm5fheXGtU2dGtL
w+Wt21mz1y7IW7SGaiYMIuujF7zBMkYB7yjgu/BITWxhUisGakIkzQAyqxAC
t0Gy/2e5kShXUYgy0SDVU59F3LtCO99VXy1GNj6flBP/UYL8cK1BIy+kEA7W
0JWXdyrHyvSK0xFbYF0zHjDUFFabHO5pjRU1gS5w8jMrcnnvaJ/3zvaM66ib
kOQs1eizCX8GmQfDjWtQ6YkNqGFMAeLaz4Q9U8WmTAXeKEsybuNnNQojqf9Z
NwsZSg7SAyZV08y3y29GWWuFJwAK6JHKR5cMu9KRm2vEtomeyRlxs+xfnl9x
mylhgFZ1qV8KY6GFcBGWIuqUJbXYH1KhymztOy+q9DR13daQ9MDCr7awgih8
GdfdXZ5rvDQ0hsWbvabdBxzqQl9J4e6bLtdlZ3NbkI2md22X1dlI1jdVsjjD
jUzE1Q+vvJ2tiaZZnEmnZNsGoF7t1zcsHw9h4WMmS/cjNsZe8GmDKdA7hOuf
oh+vuY6/uxRcZttzbJAmtHnDU17ekxOa2Nxtb8AhxKNLzKkSWmoLPEZ33nJU
ZQftu+Dhocp3SGc/k9yU7TBBYHAiwrh4zsnA/xRibkesFfSgFziQu6LW9MI5
6i1E/91v/PqPn07HYIL/sU1mEBNTPSQ0QjWnSMvQtvam1w6GFTV8TG69fvgo
e6Ty/j4RPYXjwGFV8WrO6S0AuIdbrbaRu6xV4Egolu+ScWVYgCwrTWreT5RA
ZT8MBbA2lMGHw4zsHuKJut4UME4LlyKhTeJI6zj/XlYKA0TkDsPboEM85ElS
P6Epio/nbjuvhJpbcotJRo+SY2HSctVWC/rgdKeX1rTQF0s6b/UXfAfwD5aS
WycmuSvdSSCzQgTV9fm2ZYTDUzyqaefGkLonjbgD08YN7j1JoMosxTxNKhqb
pxj/+wYFyifEEt/tAzRc8Qm4fw76U+x99Nq9uwUJLTlF2DwT6LJG5vcn5K/9
uGnZqb2D/06MkBie4qhQL8wPymGzeoVrxINBcuv6fgd07MipAufsd8CSG0xz
3lSJL+d1gtO2YW6gkrC4ssK+shE9CbsGLQ/GcyEo1zI0WYN10wRoFseAFBQR
2yUKmxyz9w/+8cKfX0iGQQ/S52FuVfSdSKzBeaKhfyVq6mhAmktwGrV9r7Qr
n8grdFIKJrE0Nbpa0/2nxOdyHhR3obIQY6RALP1v7Hzwl2iA4Jc0M/j6WXEr
H+2xAeFwQUae33+zKBLRxZk/RaV3wh8Y0NgF0qJgt/3eyL9bstEutbeUB2xb
SEM1Ep/tCjiFUxpV5bcYpkd2j0w86/cFk1fPw+l1dhsxs0h0WqGV95P3VZ4P
pUI1pRZzajDujDNyTcZ9xTOS5U/F3p7HB/EQtTxV3lUe0/oyOhHFp/AUwNd7
dmy9/xvSbToWh7kn8vnZSCauVbyjrwWfHB/J/qsKGEUSNqOgXX5jI6e+7Jui
UiJN6Dl5+jkqitNAtYbI26ecus36jCvhzUSEwruop5AdePlesmIDgkuHaFy2
edVxzS/fmpnF5jaihYXdUfbKE349xYtHfH+LcUaKsENkdM1+LqIIYA5rBM9f
Ql81HVy87iaLLF6JYO0JS01SdDCSBjHfDQZirU3IPLI0/gW73slLsj5JCZGy
21uUPVOWaUGjZ5YRGbrModgpP5l0DAALFCBRikJZLVw1m6BrF1pXMGzPnZz9
b4Nbfa5uEETmNHI6Q/dD/8TR9hVIdTjRwHflDy1Q6Re7eSjNSE7RYvuISC4s
3Yw9xneMvo1QnXHdRRPG7cRFisjGe4a877JRC62MRJWAfGd2q+QMsURmlNDO
DTXZaAA7jyfJ9WiNGwC8APt7zKNDRO3slVWzgDxN2NjaxW+vTGy20eUMqMqI
tak0N0Y3Ki9/2jPl2FIQ/mSn4sWgIcylnA1hRxLD0dUV2J5EoG8azGJMTWBx
jJuVeW7aXOCf+CMq6pbI+MjaNki6tlsyNGT4CCKYDQmHPzbYhsKBiHFPLlpF
UfJrlcq25NbmfXB9D8JRl0uH3QFT9oNy1n4ZoIJPkSbXVptRxnwHJUzn79DZ
arYH8YKjn5GqXxgznfPbBZvaBEstU2bcV1Uv7cLlDPyPYA+T2LWSO+2txQ20
KY5bHN/ptIK/91z56eSjIVSrBVgamo0W8EkiNVF9UaLB+uiDRZZ6CbF6alwL
VmnS33zi76Q28fW0JiMqY3Lbo4CKKxpIIYLxOwqXIqWXhPDghzbzMJPf0NcO
c+SjNpsAXSPjQ6s0/omAHS26IGQsv+S2b4tqxme7VfrwvODWxZyh5p7oplJD
16Moho/A773Drt/rAIwPSoj5GYCHKENWoPXCje8tQjKt7wArmmdnGwvikCJP
x/lOizY4z7czUGcegYfAn35VNmClagZVrfevIue1dzkEhGzrgujF0VmINd2O
9XyHYYo7IGQpp4lufdes7W0a3OPlZelk+9/89wPSytD41MdL+3WgUvlV9+/n
fP9Jgr5ay+s95B1cx6F6AWazbjmDSqnAoB/de/EqsdeLlNtYXyjW2neCQ0sM
EvyprzBWtA1g4IIPG/1fdlo4IaU2CTtl4lYIms1jQqX+9eFGOmmVbELOYNAP
1qZ9sBtz8V3ZpGmiMAvLkaoVX3IYySE3HY//4zbWGkrDPay65tEPh01EzoQp
JSfAYSH5bmYdkcDwl3YFdjPhkftUMoogkhVnEgiWe1spR0WJ5UXDIjUFvDzy
svlsaoDE4RFxQG0RwHh4cd9efkgMdNaJOLhoU7NtkLK9CVa6v/kPKHp82aEa
oSdk7l5UQQxzjSzyMWRS+N/2VFoNWWiclyGSR5/5gVkZbrIPsTH+1e9QRhz+
quyvA5lIg2r6x5sxwBmH3ePy+pVlVkvkpocS2NJE2pC7svRnEd7fMSPu8D9l
01nxwIrIBQqtNbY/VelKnR58OFang8pBZVps3VbIR564l9g77FIzbf9hp80E
xjvvdUHxd2S7iuqaKvhKctNmQmXVk5Inf65PlhjNc+NfEAMeTwmJSBQOrl6m
+0DSlkV2S/V69DQutr2v+CQtFmWMEdm4MvWyt6hg8n929M06lO+MnF0X9mMX
jqq6bso52itOcJF3Teo0jLkFJUgX/TuxOiLtFIVKC5ZjjrosbVq7+dy8X5nZ
QTSNBm+iP4zWqOGJrp5lKtnoq1VKhKbVDoqF4xertZPOfD5QF4Kdm3uU2adv
GEVcevDzpXc/zSLG98iCM2ExQ67aCFP1qrY1ZnQh1531Y+Kv+nhHfQFjofBq
M/auqN6yOPR2mf3fpJS2K0rS9Rd1yMhAQDbkGEGX4EiCXZzIuKnhfhoJ+HF2
uTwy1H5qtqI9miYhZig1qoZLx1hT2uCc1BKdHTuxuT0mBUABQsMubMXlZ2SD
NPuwnwMS3KFqQqdqcyxjvHn7vWzWQ6JnxiJyjH6YboBxXGo3KwwdhFc/qP2u
TLshDovZQiE7sOsj09KyMSTddChulnxE/7GKyy0q2i+ReXEUAPliI2ySYTHi
oducsZvCcXksU1IkAH2RuedtzsjOsluIiXmItwEdpzJx8vkTYfRS5oy+EpvA
ECptsE3zt6berz8f33ErG4WRaK9HgYHJvCTR1FzP2OoZkkEBEiZ8miBgC+cM
us3peO3xA25xo77jjApGUKP4R42gsBqIMYtKnF3YyZyDKqrM5B/BzRBlq0Kb
ispM2P4+GmxoOg5fuait6sKKGDBjnIZuB8t2vdiG2HoIkZgR3u6XZA+rNaF9
/eTniStwWNRl4dXnUHmygys0lomaPYff5fDYF3PbOE6/9lGxfPpXsWpJh9//
Kr5fzdjJaOLhh/HQNcS9ceNQk+HgtYAhCaFUxxiwARbmzdegSgP5kkD7/mvY
9ngTpTCWSeeByKf0kdQx0yF6cSGEIULZ5g65yQpkODuGhWejbGpbIJwpgQU6
I4mQNWW1aKm8IfmZP9n+2pcfvVdrxolUWKmfsYGXUKSvn/cYQS7Zt6n7OH9e
gXVHxWE23B6Ifg2LOXvnw5J2lLhU/HLznjHeFfrfeDG3GAg91bdSG7/MQpoV
hVTB1XWXcydyyFrvwz9nGZ7J6lWZA7nDe8P32VWAs9zrV6hk1iHkzKCdOU8K
wcAOzdr2nKeX8dfcHWrNmqcbxCX+48uSgO5dSuzXFnCYMGEvJGLWXl+LHTf4
hLo1PX9lc+T/gfhkHrVBhJLg3fuuw5M8dreRtLuQSkCQUGU+VVQZ2JtQF+KT
nqChYUzqyGf6gkNI7GgClzgN3j1gGu/h3JVS5Vep+e6KfAItyVyIvr1g3OeY
PsAJLCAWUGzmFdq/VGP9Z3/gCkC4dFnsHDOyJzP7GIDHFDAAVhj/BUxbMv/P
0oO8oJmu7rYuHzNmVUmnNbro86zmR6knOV+Giz2X7VsxYHYGbv7Hc6JvUIHg
Hmu9TFs6s/6E7DRRHsrH1v3TUOmz4353yqClIzum4mPXhKPnDuw9fRCo6lQ/
ZSc2dA8qhXRnBTJt50jsKYEpZXzbTMeAJyiSxbLer5Gwy9kF3pDNqVksydJm
nxPc3gnNNfrnvk++Q6E8meXMAi80BDUb3Rr16S0SM3ZHCKBdXZZOXN4yBNgx
0KHwug9FcxRitn9sECkS0g3ydhpYHOVblHONklbf0xxd4e1cCN+gto6yKKky
2NEjcFJX9f5YdLQoGUQOETZTshHJQgElrniWHsx1OhwI/6jqN+kXyVJWGoJq
eKllwHBr+E8Qd68hGAiXbp/6jIKdVblLoI/fhZoAwks5M5iLqUajokdN04OC
QymGylTmbqSfqGE4wKd3Go7zTBvObGoP1s0nK8OhUjR7zlQy29RrUT6LDlta
rrlohvrPQF7uC/jfuogGF7kSijnSWBC8NU6Muyc1JOAxrZPH/oFdEmcPi8+A
gykIzj+0huobn4XsjO/afyNDjoPfwMST2LwWeFAfF7wvvBpTlMiiAl5X+j/P
96WGmPge1ad8lL71r9DGkhTQ2HQMHms3UlMv7FQnjDaIVavISEqI0WESbwFB
hLK+9Dx9PtHMNrEzIOnUJ5YZS9RagelfBgGDbIllT7/Xc8laGI8OlHoZ0dLn
ur5MqeHA9agsKARcl0DDRTIEgL7Tgr55l8J84Me/ROqI86Gmsxi51FpthlTy
WzsyX+NmnjmRfCiPG/cM7P56+A5vTAKN2XXGH1U+2LGEiDYV6ZHRUVhjB6oL
XNeHt9sVTdngoKCUzYw3JNW3cjpy18GpwdUi2LWI/gecijPXxOcakeOSmSCi
+hEM7pEHBbRMBo+mp3NChz3O3jFpbyirwmgFZ2NpFdsqc21J3FJe8KQZpvMT
Yxmw64AFNsaZuq01yd+4UzEFF+ll/HtHE3xC1biLz11nDOyJ7asm3SwhTJmf
4JY1K+wqft+KvITkeaq0lwmOkm3DFaqDD2VaXKyAOvy3Qpt/6TYr9jL3ouCH
fmPaUsdXh01AWihxmM0N0/hipcsIiHEhkR8PktOtN3NATbQFT8HJxy3RZoGg
zKmnEmPZdsa+KAdiL7sfE9zli4Lgm+FHwMCrjo+DfjG2jmWrV/33bXf6vS+x
rkugSmEFnV09p6MBEdxmZTUpvkxunCTeWo0v3XHTv2TfpmhL5jpMhQ3LD4O4
uPEUlnrxeVimtLxsmJs99PL1Jk7lGkiD50rgpx2Fon+3hnKDUb3ChtPj5wNZ
TUaL8IqUGRZR63XpNz4MtcmHE1T5dAOtF0WY+H1kn16LRagYJyELPxa4R9cE
3Rd6kIoYDpjTt5+OHlp1OZTX1HvdxyJ48TPRm54D9rqeeJyv1PfAcPNBREV8
d8oudOUYTRtSZHCTflFP8QfrxaUbB17pA5tkl/Pq3YWDz5r+W3T+xijJb7H6
xvjQrqP/Al4REF7US79OxlQVQCvJgb/ny0fTBYf1lUvic1UmZFWPhxjiMSxZ
Gu9uUgw5Rbuwu9S8Yl8/NyZUskyZ425VRP+ekX3CTSlLSmAbQjac6U7FyndD
fX8EkWBMGVux7BIMI66sY+Lg/Yu65vBDG7IpUs4TUo7o0Edsp2gzOu3YkyeI
zP2rMN7Eyk3zKzhIe+RXIbI2FBaHJr3yWHtxv1PiZRXzROj3F4uzBt6X5LC6
92FJ9VtzM9cAaf0Liwn3fTVkYRHY5+8nIPh6sXHR5te7pWZCATuwH7H+Y4bv
Xbl0kOQwkn7b+/nZjot6RqBVxH6T4fYu73jYlnr1bpe9L/s45FwEwkhJ/Es/
aM9Qy1kpLK6eHM5NdztRQaCztP34ItV+jYzu7X8SVgDlG18Pc9Pg0I2nfjtL
/RjOW2z8PrJsRZN44hNsly0sNIOE0bzx0zAxHe/X9Jr97aKyfHE7PjE+UGFY
2mz7Ztr5IHzN7jwPM00gKvO2DHHUH+0tFLbxXoSkGzc7qBbjzg800gcxnhig
435Yy5XRsThx41Pnrt0fm+dPwgeJPLUzr+4GRKEKO4k132ZrFYBNgZuvYApe
wGF8y8YHzunfrbz4Iwux9coXLQpgY3nmDw945VWOgGCzov7yc7SV+XO+HfR3
p7qv/Qkz3uRSrC8PWinOCbHu9BNdhRqQ+SgZkJguF/SNSyAd7OJqVotiN3dB
LpBTtmGSIU5gCqk7BhekF55yxICySqckukH29PWulEdi2xaudwmrVmgw37Hc
VnFtusYfFE+Rr/vy8t5Uw9xS//TGm6zvHXe93dYxii/VYH1IV4GVOPi+D77D
qvHoZDTVZRe4KqheuDPYyDSqD+KpMJ/rplvvRLSui//TrBuSw4EU4RPPfkDt
h1TTgRXGbMaUkwEVB2gSdKafZkM39kBl/PhFti8WK4HT6RX1nhD3LN8nY5p6
ZXCZw239CsNtXKav7lPusUwkdHdytS3byhhEZ1yVKw1wYqZCgBZd46LDuXAL
LYdLS+lOmYd1og8XAA/TgDjjFm+Bf9VPxYciArWUP0JaCOjOADNWiL1N1nDn
a/QkIdUidJ5lbaC0JvUJw3gQOFdUtrc2aR9JOh+e5QdwYDj38aaVR4FmaZ0/
uVgdr2dOB1QYASP5vodH802dvZu0ax0/Y+50z//pFdoVa07Fxs03yAtpyYoE
sO6LpAeNueTeE02klppCbb4hY0+hFyE8p2tTlKtUCUfkWJyUKTX7rnTqpcdB
HzA6K4AozY4K6o6KgEAeFiCJEPkZ5wwkhdgRCx/0xL4lC/Ui0dWuUT5LU68l
vHL37C9TO+h26YY2i/ZlaY7APq8FJl8gGAEiMNSnLpMQOL+IQaQE/f1KQenz
XK9zYpINTYN4yryiIFHr07zRNei+/G9R7w8tERxge30XolFHTIT8flEHom1I
bjGKwMCEYudGj33mPo9y1WfcizdnaXHpewkeuk1AF59RdTlZcN7c49jKouaI
EM6F22zYV5E8ontj+dASNkY5qopkKaSA/JLFTlPHxZMzkjJ9bzbfz9lh7f1T
3K5irIAjZEl+8CRq8J2WKE+7zxQmLQPlYDZWxJjHcgSS7q0rMMrsMWLiRhfA
wlL4n33grcbkqAIiebE0ta14xZyhkTVbCbUDhpPhbUxPYpSw0W/DUsAygLUu
JqiKD5sBPes+0iAJycWcfWGQhsqj7paLQehROBKGLUngLsgYmlcbbrZqS8Kj
sKlGVPmq1WXb/b98zkR9P6nmV6CYXIPkOs9y22TCOrTGHjJuIq7peXioX0Qa
lGyAccvtlNxN1FeINXYmm1ARcrYkmcS/UBgOu7Bkv5+VLTJ62OjIMAgDnhja
aP/Mq4279hQlGf18m2mtHl4CKr4XAjKCR0nN7p8UY+puL2ln7qz3/OfH8YEf
vZH0+UHP0AVbi68ZG66+82LHzhsAR4vtDMwTM0Qelu5zfvKGkBU6Iii7+w6r
ytQJikt8ddFKF7ooj2Lg3UeDLYdNC9AgjVqcU9CkN1DibT2ve+gcch1OUSyC
YZpoXqLHonTDQiBpGZxBCMxS4h+69jXCXsQnf6YDZ0Ix5iCEEEtWZRCXSpip
2evYn77laaxwa+HA1lQNjwSfcAFfnunAsFgWCE/qssQaTAoL1W8lpid8q8Og
JoUVN//TUdxhQwnz43JSvv2IdvyJNILLvZhsilgx2Uz2R7FB37KI8tTCDEZu
y8t29gWIzpsof81Vs61FChB0pAEgmFyk9Yz9dHvssvBdJscNy7W2USA6Eg1d
TfVjfIRHhxvvAbUU6VTfCs41vQTtPfaBe5QBIypsK6DTdz/OrPXBvLaQdJDB
QQCac03D2pzKX2/9Zx5TmsmOZY2DLm3Q9xnfO/sqV1Ihwmwkho+XOB98QUpw
W/i85evr/nv6p/g9sl5dPxtiuClC4Y6Pb86etAKC9H+ot1cMV2nVqKz29c9F
72XhbBhThM6Oyw33at6Y9UnAoVmw+pjzK0Bh3wimUn7hw92ktK9DMNVti0wJ
yX0FqsAYz6jfFbh5CuW1r1mVKwtohVdj6tmBkToQuawFsS988WRfPIdZ4kgT
3n9n855UGlX0F101b088hstoBVTZGJ84zXsyWQ2+SQwRi0SZRY/W8aVZek2a
vi59sKdVokd+UIBikEgHS2dyk32TIUYbQ1/W4F8rYlLDjdVRrMTa1JveDJ5P
3l0/8Q0rK6SXpcg+A9gnNQiBOuJlxrh9BE6p8tfDOzPhH+MqTd3/f/Gs99uY
z0YUv0WgOd2bX0PGrIWGGUEM3Sl9LijnTgAdv1DHOuKcjptEpM/1c5hkFTad
EQdkxlgd1iUd6zoyCc70r9QpYy3LB5XNZN2TkaNETW9xZBnDnw8t2nS+x9lJ
5BXK8e5WPi5VGjIz6iO2DryvWI/MwTBIakbTG67+EhuyavowhDox9eZTUJsY
t/7S6JZgguc3ZgDh91PbFjMNU3SdrcwMLRKaRGEvILWOmxmRZd7Y2THpJ67y
7I+S5kuqIVMvnmfSb7JCIKL7THFpbJ1mfpaEqfR4m+4v1iElQ2ynfXgjrnhk
LyXcYlswPtEFubQj7tC/TezWNKGs6ph882VxFdCPKJqf5x5zaxaLIdUHSbYL
N6tCR0dCCX6SOYWSkBVuMEH1AiWShfNlGB/vHjillsH2578G0wtkBPdMfIc6
CeSu8Gi/iLaWpmiSX0N9ZYC1b9M0mVY1GRwCAMV9ikh/piIX9OzcOFXrnyT6
usAbZiAXyOViLJVw4V0QI08RN+p+x3mghFSeK2JO65WX1QmAlwudOOygOIm6
czdCkpFr1EL5OoTQeAl7xikvz1ZIfODZ7As8GXPak9gfx+I8Uuq/6yPvo4hz
MjesuXxOy1wfHplVp0pte7JG8PA3MpY5RiG3tJIiJ4keBbh8zFYOF+Obio2t
CxpUlvihwxMg2hEC8jJ7sjUx2f7aL5wmX41fBAV70ajDhtFRIL19NzQ5A70r
Th4L1l5wlNO7oVTYIoZxsf0Ndr0gEB2PlHUrVzZeJ9ZigyPb1u7yDEnCnBQv
1Ht3zrEk18Hc5/q7fKQvD10KTHDPXVq+SCSWK/+p/LiUKeROSgvmUwgJuAHO
Q0ak6nRF5VuwUgBaJpL5NKy+tr3EAiBCkhXgE0g3y37AXZP2Xf7VtlbL5E4n
TgpeA3CjwPvBv4A9N3OelnILJcwhtqNeWw1HPOS2K7Ga4Fiz6yAG5OW/cCWf
c2wr+TVFjtg3sWBXkOSvGICVkdrARwHogSDnCpH7ThLyD1aCOMp7H9RtZ8kS
HfplwHaUS+oQecGPYOX5e9Ch9X4D2M9Rwl6GHDxPJ/gzkUoCi4a8wbrtYCMD
wVQZV+HetgSYA+fcFGnKs2XtOFs4Ns9/+mXR/NMXsC0o6aOEm8k36XCpat46
7nwSZcdlYOrkKwMtwa6cSa3E/UTJd5Xe6xUyLS/zmqKctUmZqFAAIZXdDjaE
DnVdwt8XKVpk18z/CUn7bEdvsYhEwf2o0Dlw/QddSiNMLj7knSwdYxe0MOZP
N4of4jMZexejI2LWBN6Q+Uzrbewmc+3fOOTKcXE13PJ4Wa0QZupt9jRBCUbE
Rcl/0OccvT5UzcL4X2ATfpOSqGofJv2EWtlccHi7evPT/pSPs72alreDLAy5
VUQsAsd0Fu2VUZRTHiIlgr7hhR6crCtxmxofS/guoyaJHIxodwzeyYhOt51/
1bknlPTrclp/JVpnAU3gmBxO1y3zzA5QFUxYPXVpITpnIBAEMhaF4FGlPMQa
Gwg55lEl2eMdEoJlDlEwLoYDv/qgLLVKMPLsiU0kbrgtVWeAEZoYPtMWINrP
ReD3aWJhAWz2E3i6Fj9cBSiV9Od13VG/ZSHkqlGftpz+IEE5PeLU585eC0us
5u4CV1BdVfU495+MrBN6ocKpL76/Gdwr16YDAwMYZmF9EkdktwXh9RFjTLAu
2lq3VO5JxWEO3Bi0NOcM8TEDUocVEq/nzK5vsjYH4amhr9CnWFlyLgKoChbT
DjHwpOMy149qGBAXdEBswbrNS/akZtfIvhCp0Elsnai30l2dKL74fAx4rOyc
yPUudpoXND8yj9T2qj13x9PV/6so54ng9SZqhgM4lelz/Y8P582NfMrUbIjg
zFILTwwvTsZr2HWYLpjPnRDq+sxNgN+HSzYQ75QvEwCDdSVn6pvOYNaskM0W
iZXpF2ZwAbs/cregev+qGn1ZpsUQywSfujyTXPVAXZcv5ZNFe6M3O9wL15Lm
KXEs75fy1Pdhp93u/Rwk3daSZSXCcXJ22fwPe5MtXGwzMK53DLnigaBPbFnM
iYNAHXj4ReHtKYYfIn4Kp0hGbwlU8eqBPv14cYb385jHeLxGGHoFVGd6iLOO
/w+RM1UhYhulfSBDc31s5eWCgausaMKOH9ZZFPQCsCtkwjQ1qSF8kYfB5i+H
fVYfN43zjJdgR9O2gSDQQOs25wOjg+KOkYAjczw8XztK6wq7OA0vgfBkWkE/
oVefzeXwHZaMdYjID1jxDbEK7zUltupGnujSsIZmjP/VZFRF9YGBE2EyOgGx
iWNc7NaJWXeRJYQV0pp4nOw8//Q0vOOicXnKM7t9IlDZ99WL6Ray/zt3yNgs
CNH8NdSRAuQMQ8KnehcsV45wBp21+NkA8o+Z76PnzTDjMRmyLZXP/vNAeIAo
ACFTGPpCi6E/a1n0onpRuoxXzWwLmBAhJDd/FNnRmV3xEWh1a8OdE4jGM2KF
FYedJEwOi4dt/CIQdZhUf6KOpgV4YnJaUmfxdxTjsZjMCfM+mQP8IvUlN7Pl
w/WO252vdB6WXrTbc/l6LqR1okVzDQ2EH9qs3zuaCCFHTQxogZ08nzNNAFh0
vNd0HntUOVNieJnU+Wk17qqmdnoxFWo3m2Zugv5cUmpSSNBFDR0wgVcD4zAN
8TrybQLU5NEQoMmoGeHcUG7QhH4VDT3ZJ8mnpSGEojlg5peuuVC1dfPfZDW4
g3kNfAUqkSu2MPHb3Eq0BPm3u35tacXi8RcLPBR4dyzh4bMyu6JGsj81VZOG
p43QMW0NWQS4NC+vrwVXt5lKFSKgYWEuVQ0MR7+um6cPN/gV4jHu68P4B89y
/BnH9u1SZZ8kbCY4Zzoie1j9Pyk/QbYFo+rZlalWA8wzcjzYFHFtK+TsbJkX
J2EFShtBYgw6kVCwVUYeyLOjm7RENByVx9J20NRRfBwkd9u3DO+AuoaS+2LN
S7iodaEdtS0TaDz66RtaIZBxQs93onXpMa+/EG7sNZylVVOCX4w+XuAWGLAq
EQC0+weBr36IQ+TyOIGf+ks1KGFDyu2vQ2Zb19Gu2BZ4grXPLZUkYkCfnqYG
7TBg/fRCJRCoZtkzxOgfCEciNnvhIV2n0jz/K4X66FLOnG15qcq9X1Aiymrt
1+prdHVNm5QjcxPb0dZwBMDcvWyNJamlUzxmVPfmQeTHvH5zuXnmflJTj1OD
I8T8Xh+mMmUT5vyw9o5s6fCzKzfaMIX4bj49GeHyLuq4JswXBSvPmwgOine/
/bktVcrlATE6zbmP1m86kSBgShVbkQZexQgbKTkNBMo0+JAXstotUwSpzyck
pvHeQO5rZqlkWUqfTtNjdnEuvTgGM9NbK7jzoFtpknEsqgVz+fT6Q4OvL+IL
5rEtMCPvj47rfzhqFbNbaz7PZeOs1e4okuFxxkr1VXCbhD79wX21Ra7CqGke
hMRAsbz6edIoNRV9PPcp43ecRRWY3InyK9+o1P0fNX1h9cuen5sXja9f3mxQ
qbBQqhZXM8FLwu7Yc/v+BHfeS1abKbs1pOtPjWwTseyFrFDXoYfFwNic6oVg
1lMQnX/EhQgFBhDr1cByJreuEuH2gvnrSrLXkFAbQgzF4Rxp8kpEbe9LeAlb
N5RSS0KEvs9vnLk96pMwt8dKvl6VziFJyqWHlDuD07+YjI2O2BtNPax7YXyp
0LVuLG4GQw71/y16lDNsuQCe1Bk8YEzK2xWzJ6TREWDnh2I4TKcxpMVWRBDC
bMqp6ELNyu+N/SJScfrA6PEecUhevdiwY2nN2+49Fzqour2maO+hs9ld7f4y
IaK3G2yFoSTHnM9icZV1ZJiXxfS4XMM4qGDPVlwQHMntBY7OLmxB+BL1Rnfu
RGiUpNQRzgaVLRMEBKXlVAL5f0YXqLomeaVpFtQ9c4HM3drS5ghIIqKOqn3B
QtONuYuY60jvfvaSuNOya1e7UKgx2YLzjqk/X4kQlyE/bodrRU/IEWhjqfQC
QP7c4/F38tLaXilq8BIxmLRFmVJUYGaGq3R7+B+G8gGnR83ofunKRKy/A1zd
cDze6Jx278UJImY/nMN/XfCqCX5h/h6LMHpCE2dkTobL/gcJVuVw1aw2ApnB
1O0Swq75IlcUQr2cXxndTlUQsSfcgzmqgL1Q0MKbAiXIIQTO6+JADix2dQW3
F0X5rrXsRDvBvnRx0zKbvSY2ydY2O1KaFM9TjeiTCdomKLrwleE/ZpVT78Zy
c7CZEe3bi2wEwme24CDvHo/pt0ph2Ukiys/rJ8qGCzIDKmtpE4yW9RalRpB5
0DB5qvk82Unrhcezk2aQv6Hx9v7+CMIny3vEsq3PEyQCew+zH3TgixafMfau
BPxTnS2ydN4NmrZY97Jr1+4VEpBjbcXJYrrAQycxjOJMNHy6KzRg93ONkBrI
8LWNSYPxJDSdj5AfudRygxtRhqkF5iKrY48yx8YWKkivmt+u2ZEJhbOhthOA
cmEgcCV+P/DsxdorvoVJeZ6mrGROM+BNjV42QdfkaD8LxyAxyst5cQR+o3f8
G0ZkSAImnyig9sqHV19quiC4s++DGlK8TXV4s0OQubh22S/Se64dNZZ9ohEk
HMPnbn+136sMI1AFLlz35SFR0V7LoTvd2l5jIA8YCYCOQMTQfb2FE+YYXww+
gp3CZpb8cp5fG3onYpJdahD5QXuEDpTjBcPbxilMw9kyQXImMfrUp3FDZope
UqrVucwROPXC3IrPqPv9EcFZBjwtCZCSAOaCVqScvHWYXEPLSG84ffIaNJAo
7cneTbQBMwXcVBUrbByI26//545DrQo+xZ2Mas3Y4ACuqPSFagXXl5LlncFq
QUc+Xhdx/9oRoHLbhPMkNqQATCfYCiRrMr4YExXjeYeb49XcBfua2X6UnNc+
NVdJ92Pzkc3S+EkYZ+ATEXIlJC50Ifbm+AklLpIiFPu7aTBc2PMHytTm70+N
QtAA77uD7FXkX+2v+185sS8pDgof7rAbuQYVQoudeRmonUuWFTJsYnPmIYNO
HX5aaaVGul/ZGb46wQqfhFbO8xFuMCa74pI7fAGktNBjWCqfUEzKo6bookai
TdCbzTI1Gn6pbopAKi87fFSrEEP/MgGOkM0ZVsPzQd2cUyI4W/gUMF2fCdP2
xt8GucvSUqMxeRLWMAfU9+KZ4nd3w+1X44bF7snhMvSvBkbfgUW8LP1HAwjR
KFFymAP/RB2g+J/bBL6OeeRXp5RYTES7MDVC6c4roTka/GawQIBNV+tUQ95k
cIbpVNlUapWd4iH2G3B0/CM6Erlquu2dh+o3FgeoDVw/skyMVee7V+vzvbDP
znoFbxEnPNsVhstbfWjw/3uTasALA2pEmwo+eCb5tD1hzrOi9Dh3yBHjBqzr
a25Gz98ir3JBaoAwJECQ26n+C8ZNhV+Wubya9UPEFQa72bWSCEvgiBRxrN77
sGX8wY+UMk+fZ+Br59kViz/5gdb0R+Q34Tq+0i86lzDscBDRA2VuSLgdfF9R
ILQd9meTLCAwUiwj+7CR37c6joH269emYgPPwaSXvu5Ln7WMzKs+vVCF5OrO
3y63P36AwHiqYNx9iG3C+HIO1mvSlscvapaEQYNr6gYql1mdCXn2i4J67NBo
/JFXD39uqnkONq3gT5jB/cFBXmjlx80LVsfyluLsiDjG1mrcZtfdtBr4w8Sc
qObA8hltggahqDNDOW0F74EVPGh1YCSW+xKmxFLZe+iOWLHa93Ysbngq+m49
RwvVGNCM2vEi0ctAHKNP6KQphq111V+hlqjWZ08ZJ8eTGH5ruCDnV216pRv5
6273pUOaKG022jmBeaBkExUz/1UiiKiaAdj1f28fTKdVx/FPp/rbfc8v6G/+
arl1GMy/B5sWmhZrpjbxXCRn/PxrAL7ts56ZlSGC0BdqS6gKBXZSFbc1k9iA
ifTud4y2sCVGl9mIMEiBC7g56/pprjtTJrdL4pLVJ5hhSpRVbtUmuxjT5AQU
ovosEfUAtM6hYHFWenFBQlsgWLZzZcB2Xuf3zBexS0C+iToAW3BuRJZpToZi
a/3VhonP0PNmUC47huGqF9KI4Vf1RBXn32VcEELOAJuFjt0aWBnVuXi4txru
k3qmbAxn/Xj16IF4GyHq/7PFcVaNNUfhpbKGlobxvhazlgXfswgIG8FXypga
qBA9JsAIz2oY4m7JNNk5BLT/FQ6TTNeN6xE94mKjNvKT6CeYG+fwtpOeK35h
ksqT1YAZNjMkdgWKnJWVX0pVKV9NLJLFZWU2mtUiOH0LeUefa7pM5eJYbEUe
OvQhTaa1Njb1mJaNR7/gK5UMgUDAZ+pV7w3ODAh8iKmqcVIcySqP5zNqZckZ
vubQbMqzO3ubukdwTdT9xbyN3zjzs4sBpnCBYeCArtLAxMOEfsktpUzX9KDl
tjrrB+02heFprRQsGy+JFN510U/ltNx7OvHYKdCFpdCdTX7rw0yq+/cstPkr
SK1EWLXxwWKeU1GP0nyLTU6+TeygPk9R01XDq2l81Becnv/JIlooYNmxoi0/
bJLggShvsmUs68/h5BbBGh6KC28QdsOPW+58stBqJfVSmacPdZJdQm66Za/r
cBnL181twifjTtH29E3qDdb1+CimHiEd3gcrC7OAjU+TnPgzPZ0SM+FoZzhL
7Dyp9nD3ghIm8hoDpzQP3TBudznyoQu2WnlaTndrPWh1nv+EXU87rLIxuBhu
z32JfnSlcxzlnn5cTS6CSSp9hDDcj2NZRjV7VV9jG9FBB4yIkhD7SgAtyw89
zxOF1ZYPDFShSFV2bqZ9baNrd0fJnKf24fBSIX05KERAxDhnsDLttNwRCdr+
DiFhmmPP4Zg03dk2BIzdrfeW2pvk0G+taffLJV3MqU7LoJ6zFXI+QjqWH0P9
jqMwy67d2fxw7/Ar9RfwUIC//E/OxiHbl8Rz04IqQsrEmu0588d+AD04OosA
QrMO9JKDYUup0vZOO41MxMpeSuw9T2tTH/3HACnRt3Rdd0l973b/V9oz25CN
EtEnsDfeIMlquC2ZEZen7HJ2bhsx30lFo6aDZZWPeXM/lNDuAWCEEUwq0Wu4
x5ppPSDTPQks4DiNIMQvELaHJi2Pd1Au0doKcERNjDPkrloCw6WZiniysGpx
YX0t2azKzlW4DrmkOYHCfXH6Xqfl6meRbP+i+jCbkHswKtsJItHzjag4YygG
pYZptf/01LhcVhzhCj6GiXzyhqFiq533BtKO95Wix5W3i7GVzM1nZPasPRSG
yZo3LS4t0Qr1yzLI6pq7aDpsS8fhazBZirR8Yu+nXxGPwa+cgA/QhZhqdQtJ
Iqs86LYIHgshxgGiIkr1uuJX6kI1OHcmPAe2lfpnVqFYxnspzMAQJRFzW6tC
5GRK5kJ5tig79BeaXnHoCkczqpSngnJbcq1WTpnBtIlf31TUjsDtZ3/NpNdn
dHvL9Y0KhIxZy9Gb+5ufV8PwkGeMjrqH6ZHeyBosrPVy9oatECIT/v4HmBDi
2EQBQKydZREy1r2oiF7e1GP299JdvAAA1I+IN2FV/7ycfASwZiX7GN4pA7eO
Fo0oOYJZ0gzP3GTvAAcTspjPiTlN+Xx9uR+eLXFZeYF5uo7J02u082Kyf3Nl
PcSGWGiTNbedL7Nc9smZGis3OtxQAn5LvlyHl7V2gtnmG3XdeQ5aPZck6xG9
np03SL6XpFJUQZKv0+gWBxW/W95dg4ckkibgt5W4iFRNJhgTAnVaSDcTHVFg
C4Mr7g8zLM6//vncO0zBNOiXmrB19kdTy8b0iTBFsOKGE8Bbe17aA4V0mP33
7q3Be7HjKKWkyiZGnbBNy8AcYnTFd1MQdDvhEIPdrlokAXDKovGkomPCQ8je
cLPTXagOWD459wc1/2K2f1RHqM0E+7W3Ji5VAKJAUrqWWskGwVrASokOiemG
nPpGK9BdhIMyuC42ul1KGczhX20+OMEyrlIBiUBnYYFOryrqgjA93Dm2+YcR
7VtCXYJZfzYDu1rFLoXZrRT4/xex54o9PgBuQrRxqYSnl81IhXlPiC5iPtKf
P2qcG3eg4BQaaEcX7u86hPNm8Coi18lBfyGfGuHCphVcE66VzWPbOireTR/W
12kpJrSQGBDfNGQqdykYE+i2V9++QdAPOaTiISJiwcCDcj7tRrHfq8LImmTm
JXJVIQwxBkrrS9tKjsNTVvg51i+JIk9sAnyYWTZ5LpqqDrJDxV7eMM8+CuBR
h2z5rMHSpPDpnS7aBpCCXFSl1Y0tQd9tHe/qfvWBkt7YYrwCODhVmBQATMvJ
a581V/T6TzyfIbDf8Bo0L0H/JyuVvW5nwrcT7WbPsIpe8hUcN3XJWAJcYw8o
VNVF7UKA1YHi6bBC98/4nr0FzrIe9jl1eb6iV2iuwZxnkxJxLITdE1u6GD5f
OWkEkXqRv7uKxwI3cNvNQDTKP3gFvEfxug/92DYb4mBG5jIElfem0KrYAh1Y
0SDmQMqelevVZtZ22Jyb2qt+Te83f3o3+ef2Y7NczhReUS4xjXP+jFbPJZCe
RM1eS2Ro8cb/vrcJA5qSm+odplh4keE/nsdJEde+VM+S+s91Zkjwp/WV9bZb
whJ90+QB09Iw0HineOJjuQhWFdgIm1e/UAX5psekykoZdxreUwlk4NxUXhl2
RvEDPnCbKHbSBjcbMy7dQnLRzXc8PQkfLpuRE76EtXI67jeNjywb6B4Fmsvm
jJxmv1uXmQnFz0kw3wVCA27mZSIbYJzrh/66+N7BnkYTBJp8zHhttyEa4thQ
18lLBGVz8taoobCEIXX9VnHUkPZibh6k55w5XUTMNF+pWNk/FK23TEvOhaLJ
wG+0AtY/KGIr7KRfNuYqDi79aDuinwCS4cHXN/4drAaVs9oUSQ/9PUih6IrC
1+50fdB0jxYNa16mkGlkEETTaVRP3g12yhy+ig55dHw2+Dhfnc4uuuXl3l0o
rEmvwZJXzZIwPfYpEl7U0VeBE6Z2uBFlMW47N2iNDwVgy0zyIdpKf8YJOd4s
aVPTNYNzYq7L0nmsXrkHI3P2DPTaP2d0rEVCliXKXiqPlCSGchvYcDaGjC0t
ZqFMT782b+DIv26fGxg0eq51RhEtabvW4kwmZWNI8Zxybewgu7dbsQEKV0a3
m5ta0fcXBTEmDfmL7prSDNTnAxRrTw0skOYZlm8ZudxPsVOu745uWLwj9dGx
a9KoBCgt+XFnBn1XgalVUNoCpZ8vgJji9PEUyIARYRDxyfU9mlc1PaFWnwBr
dlVv6bobpTyFX2Qo26IPCoMrcLxJkDCCC4290ck9uw6cLx4Sp2Xtnf9+HQh1
mfnBrb0Ufwp4m2/7iG/bSmGhj999VShlFJbBVFbpySp1uvGav8R02LCNBmEj
ms/AIhti9AlvgwoUtB2vZvu7dqU1JUx0XHolEbRngJ0vEl8hazRNie7RqD/0
+BgNpoZjg1hSNl/kNzp8r1sU8fUnLLBaBcl/9TZP4yFu4CEnvZSf3z2i0msh
RPxca9LjDxkZCbag+5ysv2YH0I24XtXi2lJTQa2chVjOtGy9Eba1+vIomkmY
mB92Gcq1rHZmsOvCrue1w7Iar8t7wG1AHlmIyBeG4jEB4jalbhooi7KQM1QW
LuoF8NI7oM/z/bBGMv4UtNY9GHIk/Ccwr0DEqa+Xr3x2GBOI+CmEAqlAoDiW
p4GOGM1YxOT6e/oMcPZnRTIR7SRKnSQFMQclq5Z5VpvtwveVNEoIqOqpUoTV
rNfcrubrb7TMoDqttmC3wiZ1qhFev4z0O5CNf2nxpKMN+Yryq0x+1Zgz8zUX
m1xDNhgZCi8ogkkTBMJfE2b3YbHm+ZOHkv4ylMevMFAVmuNcBYLwQq5v5M/S
gqsdcIhewqYSxCPPB1MYwnzP8S9RtN3QRa9ZweQT1+R4cZ213CUj/OszWckV
mSoXnM5a/heMOUW6KauEZprpKi5AquYN0wOwVqvoOWMv0IiPq/Qcd+GCAX5w
cjYkFe0XXbZ0A49zXrMdsXgsjBrrHM7+/norxAutslWJxG66V3DvgMQzSDRM
xaIyz6VvRMSAdIjCK5XveKnDfjeCkrSpoZOhm/ggRiUiPLMtaJhkOhVwauw5
kUc3dtMzEGwI05KHmF8kLIaf+kgKd9EV6Utnwyp7PgGQdYIijESbLQ8wuArU
fQMcfuv1t65jRRCEGw54Mo2IoPpxc8QGC2pzFecQNGnwYD7P3Vog+NYm/TAw
rn1OBBVOBZsg5LHdeLSoz46RefqPlcd3XysdnPgIZea4/CwyDhpz8vrkm6Zg
UhUEtqidydaqbWJdTkIjUHejll2VbDXdbFrE9Egsv/XuGcsAo6kFatjAxPpp
pEhbG4tVNxM2XZsKgIOJuyIUSqDoEyB6ncpg5V0TDvskC/P7zrywn1FIywh8
J9FXoIwBVdVBXvnfNjAmKFVXU7m7eiMgw6ILWw7dI02RH+xQFwoQ160yWad5
FugD33VhMiDKUEGKlc9QYGzG9PFvDXBj+OP0E8kqqyhm78Z+EZMqobS0WIn8
Vs+xjh83D2gAdmAXDepDyvzKgqNctvtASYYNVUBNA+ntgwiC1XTEDm0EyrOX
dCb+wkQYVN6tzFo/QVkMRf5KiA5Ysr+/o3y+ZdiePZgq9hRX/kj7Q5MnF5FR
eWQyidUb8zqP3EbnujU2I8cEXWp2sA8nKs07Nq2EJbgTDf9A/PNkx69eScjW
EDDXgtCyTGz6VwxxShUXCuGENsJEgv+qOgxtFatYFPwJybQKX5X/h5PYVla+
PvtNKk9iR0cXe2Y2u78j6ci7Qwh/TSwUMuEcL1XLtnC0+85BV65I+HKkGi5J
mXZnI9g+r/aDuKadnsxV38dwNgCLkzinsYwzG1Ausn/f6ZOcb39ZpHd/VonO
Xe7wzHIO8yChtIO7F5/CaH76w2w4W9wB+dd/ZH0jVkbpn5AEC2hVM3/6/4VG
H0YJkl/V/J7NlZy3Gs2FFAe1s4dGm8Bd/a3z6rW9ervKPLKg+SC8OCKXGW4p
rM8fJ3AqAiLNMiXagfRibogcOKuSRmL/McWFbFOI0YkUK9I1ZiTV1AY/cfDi
vJRZzmspj6TKnUoLWdCSCfVsW81c0m/WpkZWM8bCHIQvTOShD62MeV/ixeK7
FhW2w0rGOx0wwSjpry7poLY2GDRTBGcEPkAvk53Fnq2Qei6paKmCCctcEx4R
UTvx3Kd5HUvdN4RSbI0zZIP8c/Zo76F9xcZofOK275Lt79BXII/RhTKpNyq4
8sjoriZ4ge1ce5Izfcc9DNreSaRH5E+gi7V0FrWYgZlK0asscM6nqr5yrk3G
gHkF1e6TmLwryLsNLp4llJnuy8U4D2opaZPFafwsQeqHciCYs1zVHYAjuu6n
EkGY6dhh4zaeC6FkihTNf9ImnzvJpLo6fOtYcz/Rq0GaV/x3eLp2JyvGrQ35
iTQdRpc1xC7jdz884Trbh93vYO9yEbL57QF3hWP3nlSS6BoH0SaPMOTAUyiK
1HAXpG3dS/TdZQz1uai8InLuRxInm9T9VAKkqUqVmStdoVnGOtcV9tqz0XiI
B7gKf4dRiGXccRZalZUQTQKB8AJF3JJAGSYYkUAFjfNcSkOU5EKGWOdaE7c2
dNpsZ1HDu298ZfagvOAomLmT/4dtzKJ2YG0HSz2ov+V3r2ttgR9W8vmo1ivb
ernui4D8ZqF436ORB8qiz/d3s+F/P+UYOaVyngcXe7JbaBcD5wFBFZnsYV7k
GmwVJUu7xfgcAf0fsep+umH4lTw13GaNxgX019RilqfbQwSwP9ubuUQjOf/o
9jtoRhIZr1Wa4hm5LpOS3Ch//z5JvP7easrSlVbPz0qFMgaz3U/LIPR9p4TD
VVu1Cj8zJwLiza3XFp1zbPw+DAs9CK3TBNVtKAvo3OwbryTO7jxd2WflQOLe
VofNlk5lQdw6dpfcTBk1YobouOIrBWVZu/uOuRbYV2cvA9Hl4cN64OAwvaTV
QN6dl8PzyQYUQbm1PSfpeUJUh2fgSNPh8YJkvOXOeGe4RltnwAiQZgYz2+Hd
eIT1WhQvLiZC06Q7BiioG7rk9Ho9DArP356Aei3BN5LUl4j3A4K4m1XNYrJ7
AnSe2XJoDWvogmRxZDbIerHnlWSBosN4cDxv2MQ307DAs+w7+p3M4Xa5Z/XJ
GhYzkRpirhAMUmOjGqO58QUuxzYqLJeS9lfbEpNVJx9qzooYVgRq0M9WCt9t
vP9S1yEt2pEU69Hw1eqCWrtE0DydALFtlwXr4HR7eUdHAB3jpUT6WEJt2E8X
QGirhUbxN0id9fwSnPwpthITrxWDWvFpl8S6gjcVQgQXHq5g+W8PySXxHjaX
PG9dhqDs+lQ28CUqE4g7C8N5cnNUqfxVeSHolvTA0JKeFyjP9SKajpjptiGI
zbkzw5Sh5pHVWWAtxI1E7km2Ub4GGOaYK6PP5XiUPcfVO8YcLk6ohlPOiA3S
3P8v4bHPaHPpRZxnlU7YqHSTRCun5Jdq/rMNlZlRep6oaBMuuUb0LsX9aGOI
hynvlKuaAD59plGIX0Z/oo7Ak+FUaXX4iyltrxpnVFwG9za+ZWdIUgOfArae
21fUGzjWYScL4CsvzyTVeVv6YwJ9t6qWajwAYJLjcu6cT5eJKfhWIs9MpejM
LfGTxBRKgg8PgDhkPVZVkFhJkL2q4MXEMOt6AvkCN78C26PRwukp3asIfV09
l0EoEeOwFOwoLi4cF/Q8vMhGXKVAOYmUsvIhRaShHq9q0niLrC0QfyZ5YbeP
4Wb5nsCLdCCszes4EHbIOC7bGj8IJEVMmEnjGwPHyoGySpnxDcZQluyVm6xx
6EaGIk+lwNqf+2AnoZn5LvOWJA04IhuVjPGJpMLFATSSgD2oQxCnL2KONzpr
7SP7sZ/ScNBCpvEAMWxhOJDEtWviZDG3jhhlzOpmOYHnwPc82K7Ox5v9wlqR
tViMKPo6uXlG9jqAtu3CAA4oSyOfhm9s2Xxpy7KFWeWCEh+zKY2EcjyoB2cs
iVrDucgLgCRgxtyJFutM68vje4BOEdENOKfRQm/0OoKiO6wXK2PM+iSWBzBW
Qv2wSNojGYAhOJI4KYZ8z0EVumvotujS4lPsQA6/yxKAV5YgXbgd26/IwAYj
NKnQFgpqig/vrW9Qw60iKjA5DI4Tvydfia9S6MTK8ekMxKXyz+zlyKAQx1wK
xumr4arHaZgnpaLO5lVF68PanpX+wnzjcBI+LgsEYA6jpYHoAxTfdzV28Z/m
N14uyWGOXgDS5edsqkQd/EHJzix9jgeWXPzfx99DAMjD20fXlm5VLiUkSBkG
N0BCGXEPfUYpUJw+k+08pOEI1Lnp8V87MZCjTU8mxBmjwMYsY3af/kK2aASZ
KvaKLSiO5g6LPTxGcPcu6lrGwMYs+eRp91efJEA+cQjeKwmDnffkMISibZiV
+QO1iY/4Ss+mfmATgHaeeNYFGAVvn4J3eGWyXSriNhNI0SZ0FrhzeKNR7H8I
2Wt1d1CiXlHd9JEEA8o5EuDyJFQRcWh9hkQpqFKAJE0BFVzOa/dOstXwXNBb
w1IsqD29qGMXEaBV3OQ9B7WdvBycs31et2jm7dsQjYZb4FJAE9cSMY28jKO8
IvmanJ3ugqvgos77F1nqqW+C+3yro48RXdbWi8XdNnjerq9331dXnJLLipfi
bTUX/vVq6nexVP8yaK7U+baj7vyUkzz2SPqUMlIMg1DJ5ny6NpMCHSuF4NB7
4aLFQFgLkbCXpOZYM3oU95tI8d+IhEysR3/zk1nEDXHOK97KgMJvzTthuKEP
PDPRvDfwky6V/WrUDHuG5PLAW3Jdqt0Tz0+UBf1IMRH7WPiEBLbp813tC/9n
rCJSStQbwO+2f3cTRzBjMZGO9iTXYrigw1fxnKU+qLDOkX6PA8qy4hgzQgP6
BBggwvstLDXTTwoGJzx7ofgkUmXjgyAV5jySpCP2w8AgL7/LHV1c4t58XxMm
XdYSYm3pWJdIbFRLn1oRSimwEX4B+bQvdaFGVcWBfdfB/uw9dzNn9ZlPzgI3
sIqGhYXyOh9BaAG7w3qoLX97Mz2M8iGf7nFZWzxSLZz+11dUtqy30xgiEyPG
hGmHUqzkDj7zo6BQF+AHdblt8zjTP2mdsPWb1a7nYGRMm3TC1H2I6n2/KZyx
ohK4Dh9KzYO1kWPSAj7Ud5De3H7goEYnBtEi161WQUtluIsbnBz7dh23bkGS
mDn3+BtFsCty5/9J/ndgQ4UXaEfYZrP8IvFs6rjy+za1xtK4n4tftcb/caVc
ZPrQ4bahY+XpBid45Pz6w9l2XLdTeIetN6/VFppgXG31kCfEMcFXB7fT1H/1
lV4ULe/CKZPbQQMSUOB78JdnkDlzICPduGoTBumxGZoyuWQg+/2apWntWinV
OJuixLtq+bp8GvUhPRzLLLIP5AwuzVPy5z3q0aAUZrSYvo6XlBgZPYtHZvXx
N58bLWeczX7D/F5hAeZR4EfzsmSakmPfsBcrJgLwvc+UNGmsVqxUwdD8Y0e8
4UMDPiqBFyLalWSb2wygYwLTONDuB+5zNn6OFDvjC29CmawAhosCaAgHdLQK
QPoQPIw59bx1U7QF3jae4XFQNLkJcUNLaUbHiXBfp2r44665WZ3JZYe1EKUL
31yrF9lWTRhg3gVBX4nuLp7OUSf3lO5c3il0EUD2hB/dsc480SsTmOwujM2U
kqKEhVyDiA7nANsYuz+unxoQCAiaHfJvQLiiglNHGTsG/qfDW0dsLPqTD4KV
HHOINVallDIaemIhoBVJ3jQNbRluo+d3Ywbbwpg3YCXXfEnWVuzMA5Hrgq3m
/XZwa6tLVHVS01MdfPxOXCtWw0mUwVF2ZE1DbjXcyRXxMo6ZZIb3JOrb/Sp2
iE0w9Gb/6AHPEGxCddgTvyit3+NCb3OSw42N8ZkTQbS5/14+gljoroAn25MB
kkIu21zM8ZUsf30f8psfKY13vru9o3O9jzFq0htRRtBIyA00CJuvvMbB9OB1
JoSmJ5n0hw8aNEU0ynbhjS9G21f/i6C/sti1FwS/rtIFZ2TuLtfhRArZUV7D
iiuxUbFBoQIZSgwCN6u5Sx9lWe0PEaXLgAy3yMIVgZ5w49V69qY8ByCnyJYh
383An+YfJjdfnJ2pSMG0BqysXe4t29sypcqrv+lxvTa6cMc+IQChyPNxJKyv
YSE5Ob1aKco15JWL0K/xum0DBHqxv5MyxMiegMtbywe0e5ioz6jW0IR3mW1M
vvG5vfzPncYaJjVuthFuc9jnTjdxK+Aqy0xg9uj7Uwl4uC9RU3s5J/J4LAd/
tYThdrf2FVLzswSFJ9bjY8FoCFfCqF140npohBB1XZZ9hJoU2xt3vV77bpyE
X5t3GJmDA3DiZUTqK1iUC6ARYvLQf75LoW3uBv/IUGYCiXBYq7/FW3EeEvZg
XTPyexA54Huau26PxLTImls2xo/98Ce9AJm4fOnPbxsE0PB+piwK6gCWA239
atDykrzGoxe53cblTENREWgi3kjlXIcYx0y6HqgC9cQKlO8SzJO7iEht+9uo
pIwlvWSnz0K3oikFNuOXOxZk8aR0IbJpd/IQqYVJjL2xsfGrCYU3UFKQf6Yn
lmLvizhwU/XZsT0aNL+2ivKVLXywNVLTx7DpTepxLfFLBlNi7NS6tViU4sfL
kRpxfeXXemv+2y3LBapyTX//7d+m5+/VF7Xfhe7F/GtTFbH7YXIhWMBmneEk
y6fYV11rl1gUIduuDLQtsSr688sWUp5Awrp+vvpHP+lVmOY3kHl6EI3Ka/Lk
dekqqdx+1VSJMOlcuH07zbtSEl+zI1GrjtlC37s2hbKWJb/6WlIwvVBuWa6Z
k1TSXenc0pYUPRQdd+SDsvy6j+ts/3LsxKUE+wib5DtUE70FXxwMIoU65DtX
w64rwAR4g2QcpH1WBVdztJtdoLAT4nSHWiP3tLilyhFkLHKsAL5C052uiwMA
d3Y/mIPB8aK4/z+QRq6Cnb0aI9cmYxk4ExH/fn2j8y2nB8AYpn+U4DMaKV3O
PQ10gFEAiOapQgXfRZlZBCL1hBipFGfkNVlcklcf2eX/3FyvUOIRpMOic6aG
BgjqCi5jk8OiHINnjs3m1XG4UlJYEvdjlyPugqSbjNlxfWSOCgr2DAzhjcf2
nB39i1Jz0+M6DjtTYd7BTW8EgEG8NTKfeRWIejrH8wa4cF/N67N53tQq+u59
2bHGqJGxDzi5Z3izedmfMh3HBnKnucPSQkAGf+tVvkpteyd1qw7O1GcPqsf0
1tWGN4TCptmI5R7ExiBSGv1vpuJKoDt7vSjjw29PvSzlRb0vTgmWEut39q/z
yAgYtI2PCxyyqOGxAgHFIuZxnGEHc9aCzp0ajmE9LkbDFIUtk/m/OAWWo87k
aguFAdfexHW+POH+g4dTtFWLn0AFhaPs/390QYeT72O7y117TSmW40VLcYfW
7n+19nP2g+Q/T/OjuoX5HVmSUigQjHMI9WWvaskU0Mur5jQ8vvHfmWbJhzjH
4HOKmxCmHoORIrecq5HtVdZW8TsJA2KmN++AxahCdtP9/HaGvExtd8lID8H8
9BRXWzhPCcZgGjFkXnqvBYRAOV8RMZbvTAONUE+JCiNUJbpdodzelLNj9+yB
PB4c7jvytf9CwXfB4qioX7h9tTkI9WKfVmuu4DsiGgE5egWmcJZWENIp7RSd
T2VaRT+2mdtrXsI5/62BteMXlXq1YXBn3IVTYjZlprstgB6LykzU28mLzxcE
hNtoHx7+ktDoYe7r3C/+pDkKcDzyUlp88YHPVhTXPcEBGnlw+ZUpf9QovdrQ
sAOk7OGwvcKXve61ZYfCAJfnJy6KIo6ClV8ElEMg494vv5BpZpLqhV1B7fNp
Geh6H3Z5ejsze9JYjUryssCdR5T559zbAKrGIQPbN8yavgtcTKUo4JvjhQvT
CM1c8FJSMKcmEDARPPkxmMLSypffUSgxV5/4z5NJOJaVm7qGfvPPDLyypJ26
nHDhCG06JHsgxz4I+/PQrasiC4UkY6CmrlyWT6iL+8aRQ8kcNniIgnQQb9ti
6Ooay12PZ1T5zYKMQttC/eNtJ47KiJnrv0JDFnTQa20sQdglfFVhcx/67EQL
7XEbyoJXwQLERyvFYFIvhcQA8Qla+X2D5H7bk7z5xgk6yLkGwmkSQdEZ76wf
SQUAafyzlXRFAiSqZXPV6pW05re72M+qRfa5zREvqb6f7Brqcq7IlUr8xGIl
VGxe9rt4qKLGq5vMK4qo8pvyYTx4lQ5BRblKQgASTvS1yWuY0xTInKcnf45T
DbA181EGjtBRsenthvjVFVUIgZv4dUwjxnCYvcgkMN89PVv7xwrGfrPMRFlk
dGClhfIFy1lPdWJpXN37v4WE+uUPxpRYFuj1fIVK/lFvEHbzR82yrsEB0gZo
fhT3k+SRHDKcJjWE4cR/3PbdOJbENHNtgoZqyHCQkFAHBHqzrzLmzdihX4Jc
tg3m2AnMwZwwo1LK6sjhAe8vdI/uEg+ly5q+rFFOnE5LKc/xfklVDb41VNQ+
v9eaP+pyGcs0rAOEpSPk5zE/v5TuGI049WteoCliuPkTutW0gFC/YTS42hI5
PMFxHK+ZbrjhE41LFbuIhObtTnBuNx0E+kyc5Gnzlrn7blig0sRa9py9Ulgj
vXHUjsOTwsODVUkvsxTR1796R90qS9NXWWHiCTNWbf/fpW8MVMQvUjSHxk+P
vh6At7SGkbAYzCAZUlVQjLjkx9wwC83RLIOErOYw3lnFEmG2U8DSNeGSi1Dg
5yJRD0zqXsFnFO56/E/mZOeCpbna2AwP3nmYH4O+AoiC5YVc5HHyLAndNCc8
RPp9htrbl9/Tdyz2fIzvEVwBacdRG3e42qM1Gv6s6diWmTgnRd25BQ+VSNkP
AsLOobqSfVbA1jajR27k+X8VHTe3YpHbIzsRH/CJn1+ZX6PZ3sFjuBV7hnPB
xTm5ALvkTvKceJeKa2T5wUdRTnro2WCrd6COWP4QJe0L2GUs19GpjQY8DUjt
bxsxK27hN4N20DdXGmLKVcY7JTZQH+H+r1W2nlTGCM+iVpRj5bxsC5Z9hc7K
8hgHrduQlSv81MIZEsKK5cbrPQGpt80WX+2pyCSJiOAtyRMJWa+7lHasXgRR
6yWFF2oQsTwyO/2Lv7IFV8oqCou3oE6SZwPaAXl5D2TKu0TR1EXGEH7RS8Vh
l/NmzYrVyLwN0Nc4mHo/Bor0hcJBfe3IsIlMUgcT9rTMaXdOTsUlzcIiqll4
QW8he1UQkvEBR5UXRgARH4ZWNNP3TU1IQ+3Z4jPRPN5imHsABhd6U97KdkHH
WyqbOaKKcUfcbL/f3GxkfFaovavyGs6W3/FeWLjFtf5YTFHMpkUjZO+eBjYp
9d8RUy/Y9xvpy66NWHk/Lp7iE4H+3oO8pEF05a9RytVFY9pUWy0ojsb14Yj+
Rzf8sLdnjvejhq35RzItD1R7AgFxQC4DM0EmyJ5WxxYjpGLD5VqHWmUupTcV
34AWNhP5+1JF/7RV3zMS5/eZ69fCVIZt/y6aY+8ph6vStLVJ/kCPuj51Ns3H
7XWiKSxriIhy9IJpGTxOT3Dl0miMIbeu1uZFfcxFJyQmswrcr0ExQMYjLeuu
ALv7mGKsV6Ybq5TeNQovBAEhiNkgrXzS50B5DhCtJhb+SV10gGdo1qc3H5jL
T0QhClIFlGPU7zlc8xpQTC1Ju6CWR9BE1aQQ21KYVaBptAkdIh5QsnmGNQrE
7T/tdK+MiUPPJ03hqF3/n8uWbukRmAd1CsDciDnZrCgDolsUmOGvj7p7pJc/
iFmHtD1O1UPCceG16ogZK8mUo6NfzKsTl8wRFzUet7RSLbYGnBQ9F+F99xWj
430Y8UTz/Lme75zbNJismcC03IvqmQ8tLeAxWISQlH0bE8HbiTQx795cXgBy
q0w2kzysgZZBGKYbXiZX1honTtPpKTfW35TUnug871p2sr+G7d+ecJQpsIN0
XPRXy1M8zK8ZT/secYB9sCAyU7UTuP1Eis4AhoxcMT3vNFYGEbUp3bF52X7s
F+dVAyw2e88nKgU60oX1OqQvoOFtc/KZT72QTyy+ER4MqinzMG/QEHLvauqY
vkWZaxDfoLKnuUEMtXs9V/85ul+dVYa586JFiElzZaIfYAcyWN7r/lITBzv+
kZJV21R8SBltH2JfizS1Nzzbz8cmTvwO3DdunKPcGm5TI9CntD6Iu/6Gr9Gq
pXY4aYM2JXLMV7APwRi6/ZBIPKpi88MXH36TF64a8rgGuB0Fhq2k8BZ0R8PY
Paeg5RL2rHkTfb0CUsR/KmF4lrP1EwlEkFAREoXCej+mSTQWf5AKjtGukXE1
1jzfxKNj9pTMX01jPMM9YOmMoyETuzWHrBWOTk8dwytFE/iACF0NYEhP599q
01SSPBVR0MdtgDtep3jvcHinA1ZuKRzY+t0b5Vh8xKl7gEEmA3HtqBVGBaM2
xuIAsEKBRyCgBdrhAGOpJ06XqMSOQTRRiw/xb1jMlg6fGyBfciM9kPLA6QPG
VjSJMJSQfO1dELsQzyz19AzjxihvEFC1hRvtjyPl3DAu4Y43E6vNMdN88Klx
FPp1YAyXQFeAoyomMEcr7ULBSpMziBAVh6lT5c+UKVVpwqjRvllpvibhwhA8
SBYvFpOYWZ8xbw1rJxGa9LriFN5bpSxgymnIoe/2++bu6mB0ZAoHnRipM7Ih
vcpNUuXgON/kmSolUY7Msm6HbNsQhtuSN3U1HX8jH03QQtFtbRiQX6I4+NIe
u6j1T7WvTDKAbPA5U4zP9QqPy45E1/LM3bRppdKqm1WSycagLvr3rj7e/fuP
VtShbO5UzMb5HeRhwSmD+Gzy20YUvzgCLD/H84b7yCUZ6IEVgJB1NyDv2lcC
86kyaaAo1qtI/uesIdUBYvoxhnGbm303zCZb0LtK15FUrVdRwyJUNvhzwHb3
uiXCNAe/JqPB3T+zFkOf3KNcjv0a+UTCAKzc86d7PPc33RdUdU4369jMLORS
iq0XFc7vvGlpfIC7wPn8r40/fE7f8PVVw0160H7oTcO284z4F472xy7OBEWK
8PrkwW0HtfyeqIEKf9FC+aYqAGuAUKGGdg0nFO9I9Wi7+L0OKY3uz0z7IVo9
9FkfEYlKSn0VBMCICQFBN+lRL6kyof9Uzgp6yfUtgh0RzkFsOgBcu0i/8hLZ
4mOFpDXEDWavaGDbE8LOnkYOKimb42KTHHIw6GG76UbYnoPIJiqaP8WDQR3r
PB0JdCO1A1jELHG89TKZLTHram+4aLHMwTKJGN28mRYlUnf13J8BUVYS8iKE
HHLvHHfmylTgKebT6i4RHUaTev8+9lHhlCVRvGpsQ5vwPVs1IkT4FdhOPqRf
GoE8vvU1MT4ajvaL7aQSjQvE0SAwui0CFDJO8fmVnlQb0qgPkpk/ZFeV5Kr4
KCT9OOS+vsj14gVeVCqQQwJsKnWhBLiBtYBB706NWyw+tDjpI9MfvKKJg6bU
gH9TPChRBM9jBpilsFWl/PMdXrcIkzwCjKtWHCOM/NxH3XHJy9okuhmD7L10
4DAwF/eO62ki6ShsCxekCvK2HdQV33tBPwKbEVIFFWn7gQVQSa17T0Q2dcMr
1jrxzGBy1z43ia9BKuryM0ha7ZrQgBlTIpEctzREeMqZVPFbn68MyFCzL6IE
C2LaHfdmc225YfZkzmHqoitlpSRykkNipdk1x8XxO8lvOBf924ptMCDRVgmQ
lGgm9zAlaIF7xF4a5RBaG8j35bMwnO7r5250wOIdD6lT8QnJa1eAkbSDkgdz
Oh34yI6HPkqr1riP9ywpyTzlm4F4kfID4bHMGZ/mDu9eQ2OMLm0iyz2VACen
lZP0KVXBe50+LzJv5cgCozY0WducHTolI9m70O5D1RhQYMrlEkypoRPrTFej
di1aHLkrmlRrWYtLCMuXKLheGvZuETeoZRpdOAmBBPCEEH2j6iuP2lIxNnL5
VYwmZODYy2GsUp0RflnaajgMkgJRKhxYxzdnI/0D+uBplAki9FVL+1ru4P6i
GnlQuOAP0N4S6pyGdWtuZbUw53Wrnb/2p+04Gof9bYIp1nNNTHdTYFYDJ5lx
3ziICBy6s0DY2zhVVQmwqewkkAouE1xtLYK17UmkEt3JSPZgODkMAYP4B1s+
oAwmBW7LLn1PkLO3SGN5VT2TUTmz6uU87A/SthqUumOkI2FgXTPawULkEHam
IoR3OnPGOi1/NeKuxlGSLxNZXMlzCtmhAleCUo7SKJ4VTg0bWEtpt24aRX1F
V0hZ2+uRoWML/boKGwaEbs4OLQju11gA3ySv1RaG50NkmhuSGglpidkB1u15
HAvLUQfMTPhiSJPlP3u7/kq9AHvrnokSykk+0nHpw4ERGpJJyPmtdVsWWNcM
/FcLtWnxSeOcm7jE+kOHWcOkPLMQ6R3Lmakjl8vlgkyrT/DuSgKc9Cp1h7Kf
/mpNycmhms9yLtWxAlbpJ+Miem6RiLcN8sqzQjcUNwRErfj9w1SrAj62Hb0j
srlEHz6mnwW/FnyxalTAcb6qitPt6GLjwvUUigHWiKT+Q8s6QchxNhGoM3hN
+0Qwjxcgq5Y/FSCphrjb0HHLAvpGsf5DGUbOAxsc9761u1wDwnGmRxUhhTbO
+oQ0CxBFmVIm8zyZmTBgVfD+Cm/1JQdldInv4aIq3XDO35ceIOgvqVEUPPYZ
iuxfw49rQO49V2nAb0TGvaEU4QeeZM/t9WoGIu6pi/U9MkHQS5Br0rBS2N8m
X/drO2umQWSi1QvbccO8u/sCPq3jNr3VTj6Fz4+oBOO8YjshsIGiKWsvfFp1
28wwky38iN9ywdUGu9doYgm8T9slXKnNkOqGEKTI8ccSyV7lh1x1FVMCT/iG
eL034UwAVrkididJ5rOfP0c/chDBS2Exv4Gzw1/7Axq+lBVQ2UefN/DNn9aj
nGlXN5EMKT9R/CxeYidId0Tl3TYGLsQKM/YqBns+Q8ipOkW0jXa/KjV5bp4S
DVgtuYWc6ZkXdv/YnYT5bG7XMuPe5oSKXqSARUPVPjsAnWp5cwtDLpK+huz+
rvdKTADEbpNdvkJIEN255wEKpmeNBvOi/QUCJ+hsK9WPPBjfiTTaXKKmPSOW
oqXdRW/stXUTm/38SdUDBe2h7WLc5cReLNsU+RkhVdF6zYKcTANPGM6AZDw6
gyc1CTKu056fFvmy3FmAqNTutVlEMISBQF1/rFTVEOsTOsb2/pVVWjC+qgLJ
2ZikRXIMFTbBocbI+M7cG8V4rv/UFGQXtInm6KG7zZ/+kC5IRvXhUIF1Qyc3
/VsboIKdZ9gIOmDZ/QoZUecvLO6A84o6luJI2sKd98Lpj99n431Gj0oAev6B
5oy43Keqj+9lIwVV2RuKaFD8b5EW7yL32XGLquglJAjkhqUpfgsZLVXOkK29
CeWH1lDF68KKc9tuex46R2RwoFEdyU7ZR5ItS+YjfrhjJYwf29bQhCmU3rl6
XXo9NTMIYAFCmXGxKcU7heNu6yrflkED2w03BWQvUSAcOh5rBlobWDQtNMyR
DLtPadpMnKjE2nSHHILTnrn6I9vvd3f4uLKGO9Sw1l+4OhOnPeGDD0Y7JkUn
56GMGekfu1c33s+9M8QVvTefG7fgOIvbjHO5zk+FDilCFulk/bQ1bfqVEO6c
3zlC3ONTIecmK1VmvVoO/M+z+H8Er8R24+aQTeyag7jJASFrhstbwO7IVW5F
BtWzkIVdNuXtFzBQDXRBUk1AjZHhZKaqTqRlbgqH4gS2x8WocIMZsapqwNY9
TAaNqPXD57bIWlcLbiq8UwYkCEneb+jDVjCME+l47nlEjrddJ6TQo/I7fXsP
uaeCTKm7MOJtQjwIWH3fk1zBnc+oJJDfo7lPCRnqGtfl/ROYAzj20KB0wXLj
VnxDdkrw/WkXY8eoWZps3UVsrafNmlkpwLnBi8n8xEDG5pAletKzDieQmFI6
SPpqTYrIyAHscK2NZjHbUh7PckQESuA/SL0Ol2Ib4IzKJKcaucxAsG0rXSgC
p76Rup04zw/WzWkYK8v14DLnsqzuKJS8szPYzhB9ux+e6vTAv5wh7uOcFc3Y
sPGQBEpMVj6wJb0ucqFaIuVI2Oox9gwCW1Ank/5L0gv4cxpikZDreQ5WAXtV
CM8BhywQZST08ZOxPhXOYOkgHoIe/0vjkZH3xXB52AaAWdqITnMzQy0/Krlx
geU6fztJZN4y1IZHQvHtYIM5jgPp5KvndAr0EEIasc5ZZvkPDT/sSZWxqDeL
3iafbt2bwhRGfP+NsLRGpMlHn5O9P5C0pOztBf4FmUpwmjDq1IMrQoM8yEy1
EQiYtIlrkKm5jeJJlQZvLRsm9AJMf7BFhW0KD8XmZ7ZMfGNjX1fiFKLazY5h
Im9YOdrFdAeE6Xn942Z8ya94xaQiiGaVH4EGeLvXtYkPPbbku93JENNVZ0ZW
ZH0wbCY9zG/4LnagoORTRFv1II8e686tzhsSmQPDdwFytXcUMpelnfMXynnD
IyUtN1iGyc9R+17sQjQjMjzyRfd6yrQUZhq7R8NqT+w//GWZW4vqUUTb9B2H
QbGxbzuaBun4v1NCR/hblDEkHHCp9ke1cN5NEPThxnyYLSR1++1P6JJDqRe7
QokgdvIlQIHSlYE4BsbKP13doFwROeE4DcKTdrJowIYXXdQomjlmhl9zLWk3
a6Kr2nNzfNCif7b/D5AiqpmE3vdZSQIBS96cDSKf9RsXZkyKJf2v4q0HCVpA
/HUYgH/eGP3ucku3a2NwAoPRX9J8vAmCCE3C4BdBQNckr9oucz9hkwlFQFZ+
LrOKevwMt0A8Ko18jEPYdgIm12SGlO8535r3T+vNjabwBhPy2f31PCvXt1zn
OTTbZIa4CQEAYGxTIX/KTZ9sQLAhZBbSuRndhzH3sslh0jAALFwaBehT6mYq
4E139fEIlLEhRJMmCKFOItpRg9EtP45EcZrI/wUTAZv8w59F4GAKJ6m9ZQwr
jM8a0/p6iOKO+Z3ObjkKmnvT3PosRuSownIjCA7CpJJe+4obJA+RDfPmk65P
FTvGmUQbb3ItdNfkCVUnAN6XTSj3WlEuMzBjVI8YaliaR+vrMXJTPJQxkuyO
sfOsf7Tktsp0xWT8phOam532a7m8YyitFZifdCZAu3WejPMLT6rj2fnSUBuA
CV78IYY/+S2NLnH+nuq0v3y4gzBkjJGzVQGyUHDrbXSr5JlIE+N9FNdz1QJN
LtKTVapw/fx4ZllTH/UkYVTnufwBSPw4I/Y3Mz+VH10LbL3PiEMb2D9iwBEe
UclAsXbCfeB3bUs7YqCXoMsxTEKMJ5pUTDR9ikVGUMa/2nEjhYgDQPsYnuYZ
LGuEww7FgtRAynfxNrnuJ21FOdkbrJRok/wi8t6qwrO2C1BOKLOXFAE7gUNZ
i3LnJSCLklyJ4StA95OwFH6XiOznMLdqX2MlcZZNLOjB6uLgDdxVbVrWuawt
zERRPogFHm75BZmFB/MauGJ/Bc31P0Xv26/lHEaQm6ZwK4rmySPJZiFwbiti
2ChDU/PpA3Q5MKFU4GSxWmfEhYzqHUVtObijDn6Z9FF8cJw24mVUH0ECqpQ7
YrCkS/exoB35l1vKuKYUI5nufpvj9NDSU8ayZp6e/F1b6eLD+mviy3EZ5/Oa
WyGU8BjVN0hfsZOamyRuf+cT+jivpG02hkqIarT80qMMiU2OBgupuD0qU002
lGBC8uFph9ZJi8InSYy85abuX6IWe6W4SScmzzgwk2ry3iiODzPucIRB4Vd2
HJ1Oy5kwIX57BI+IVxrbG3HvPmA6QQ6jP6Eg0A+uiHNzQnSYET3T880DDmMk
MObxdM5WGJsya/ugtgNi2s9hpX4ERN57IW+k+1YVRqnZUXM/EJHn6I+C4aC0
Jpsg96kxsbiHln03YYIAy1GXHwI03R8unNQiAYBJCp39R1bkR2QMiVuaevK0
EQ7N+bdVzVK+yadQfKCU+g0uGX4q+B4JhnpL6gipG8QxCkbSEk37Wg0A/2Tq
zDmL5AORXe6iwP/URfO4MHO4zH615GZKKLthKFcs0pW/eXh9FuozFx1FQJR8
CXWF5tFmqLrClgIn+KnZlo8486rH9uU3GWHN/R1KLWXtsvSQbQQ0Pgrr0fQR
QtgT31+0gOqiQQlMBNzCAG6LUIAs+/1IMYKM/B4OztuESkU/QzBgVoGr6kNo
+Lxado3fDIcqcHfHBU1dSwkhVMeSUTBgzomz/7wlHXn0MA0KFTpkFoGEgyk/
gsdzJJeQfahn6DXZeuIIY21Z8I738Ssb9r6qKAmcQkqNyYG//etL8kkM4Nyw
kVpoeVCJV5euOUBR+5dUSqJx4jkDpW6D0yeeN3KrlX75FA8xNgKJwkVyM/6w
+7W4RJszHNllEkm5NsyKhEMtseYhQAug725qJ+OqlRtrM4YeIQMwcL2hTCt7
wwEzgLZttVu9Vn9XaN278p68zo/lXojv2gw/WvSZGIWcMBGYIwxqvYKYRruo
E9nXl8XxWsBJOaS17dVS5Y+F+iQBOG+urPpPzql1XjIUdU422kQjGwSlhlWE
kn2L93NcadD5yDO1KSHtlgC+h4vPIo0jWVfp6pLCoOA6fZOVZSFo36kELzis
+28gp/KtxqgUnSeKaX7HKeuqJXG/JW2GhdmQFnEhRxC0A/OW089ZL0/oECjB
lcUuLbKxq3IFO4W+h5EEx2Xb8f7710AURTws5+MEnikDrZq5bTssxTnhuizY
O9/bVjnCRo4apKCNfbJ/ySiW9GTs4wDYIkr8AWJGO+QNTxIvIz3jgTlC8qdz
rF5BEerR6kWgFPNZh6UEy5YX43s+eAMyZ3lTgJdG75ak6c/GEHiChxIaES9X
pd147tYO0pkxT6IC9JOhYV4jObz7wTsfWZZrtnYTcuyTAwpeCWuyjDDdwqAy
o4Rk4S8p+BrnlohLjD4SsPpdXuJqyQ5soFBZfZdaXw86o0brY1OTPRGtwON2
xLtJLrUexuaiZinzJxnQdzxrRzOTnobG0ay0ZM5Ef/rSfLukv9lN4mFlN3LZ
HhjaWk/6CMiGANiOia7kU2iZQ7XX5pwP9nF6jHBfumejtMqPV2rk1cwO/440
itkXDMRnHYsh3MwCX40l+naEWTbYd79ZcIc3ArtLOVwnMYEjWcu+ffPuoxcK
hjRciyYx8hhbCfHCO8w0Psf1sIyExez6xtJR+DTfwKijC1PsAPtt3U+vLo2P
Uo1B1BsGnWZJn4q0WGPU/seDTR770r+LXB9zr/t9yy09NdeWSiQLdtTv1Hqj
SoyfKlUvWfA4jzs+2xEA2HwtNZTAKa29NgRkvskXH8p3YdGucJSj9IlwKEhb
bF/GvUpBgOa9HszcjTYPSc698xlw7ackp9ZJViN6Gz9JXm+aOsGsfI2X1v+o
ql29KIJU9Z9w2DrodAWVey1k/W0mvuBkJ6ij6ccEViUBpsuLdPPZ8rCydgK5
3H2ZmYrfzISiX38tnYNGfbFPBPcbmUE/u5XW7TUQFC8o+dyENu8hNAeORuqf
1IbZBrnHN4kfexdWD+byyD5jVF4acGyLF/XNOovowDaxQPFWEmGOzbeK+Al6
LvYfxaBS0Tv2LJx/LB6j8bjPaVnFk2JbQ99QmNdYEJOQzVXUvC15nyBSUviZ
RpnPHEf/O7rroujkDkCaEg6tvLyXY9NShCPOZyVRJnT1+j/05IIfBDW32e4s
OEOwKV4LVtDSzTJRDVUhQCXa7GnDqb+XYjplpskv3LpTBpAVbpUl9NXmem3D
o3fxPLdxorLc/5q3rddNddNn5yDEgvFpI30ril3XMrbS+DZfWDCACR9mt+Go
9WvUBXNzb+LtdZOt3dFey6BAVvr4rrhpqIO3sVHzqf0gCpVGx0bm4M6j3WHM
CBn9Oge2wc46rvtcDZeVOwMzemBn2d2IgtbTeVTUfF2M+ywwEo82SSDPScwH
1z4FHiYmjVWikFPaeMNrrCTtH6qzmWM3l0IEOZBs/ZeWWBRVUkFBiZ9m/Ki1
aTtGj0JY04UZiwj3h3fCUysA9dukDcGdPJrnjGtzYd7/RtLgaMHbVl+GyX3c
3KQFvrg6cExBt1ACSrOGpl0fWvi2J+0JpUXdNF5Yxhw9v1/jrKOr1FINSMWX
g0bvhW7DQxaPsxxBz3/nv4lyRAb10XhVSMeNTefd4KbgrJM8AvZuEr511aCf
u5Rdw+bIIXknNb7P4IpiCi5JWJJzeNP6leLVt5g0u5Aq7uEL8M3F2JF7DoMw
j5HDAwLEj+pbWh4tTaBbI3+58m1vVc6jcLSvilbPbE8nKZMpMpHUnwDiPhpM
RedZh/mEopA88hrsZu3zNklQsPH0W82iwdY9v8tayFI4kWPRujK50w3hb4Sv
9hpdir7rPxAeyazr304NiFxEG1X4MO0jb/snwpTr3C00zqrQsHrCPFyD9noQ
DEk1zZubc/dXcqI7JJ8GRcTz1t/6oNIpnB5rO/LArFbXJioEInoDfP220h3I
CR0JWE3JApQP+ZTgddKUq38KvurHCdpOT72OxFP2bPFMLMpsnj2Nui7PyeKh
+4La+YnYP+lu+FPVxtd+BXi2g/6F9d/JiCXiNIONFyje2ahRVNnLw4HyBqO4
giDRqtgEEDqJrCKw0Vs1hNcoHXM9TTyhjqwo5KKW+3g8c4YXbQvcMDtFT6Fz
zZm8n1WkydVCwpe43c+Pyxe8O+89V4K193Ln/YnCFsrTcqyS7zz9t1tPNNGw
kX1doVp0e1CKtBhitcaJC1MCKrSMwFE+H4UZmG6aWnKSXnyKytCFDrXrXO4b
fcE+VAtBeEsFvfYBYVPlkPgdx/5K9dmHszZVLJ38XWpppZVVrnNmDPPWQnKw
3O92RLS9nogDUIX04yrMqhpdTV0zpwjmu8CnojEaY0xqC+Ygnsx8wAbEtNoD
RPLxS+Sxs5UsT+cT2l2FtaMd9jv1QAmjMED1rvcpAaCKV5yNMyYwedLMWZLh
zj4qJ76UpKppQ/3lbzIiKQexvOsvtHmFty9xNJ+HJP+0sE11jZP5gxNFyYus
IeDL7os5hbg4DXQP2q7LJsWrgpPGdUgjUY83B+bFpuCPeDQxBAze1TJmmj8H
ZOxSprcuCYj1yjykFk8ef509FO10+ugxeakfOCWqUUV1C9BXbIWKk2VxEept
cXV7WfYPaIQXcMAJEkNPVsha427cz+R1CyuDW033ChKFGYxJMn0jBIcuilt9
QBaC8GJ0NeG0fT2oMBZTUxTofGVTUXLgzHsAP50y3v2B3q1vO9DVB/K8NOvs
aqmTEna6P1HjcQCtVfMMOuxjcp6fEhU0AXBpGIEnFcwkfBKcdBcY4Qo3UE4u
M9CCeUhS3ZUIk/FgxywwoaZ9aHx5ejSYdWIiX5ZvTU/XV8I1hM9Di/QN9c+I
8MGHXbwlBpqx9G83f0tQurI/NWhxWYwyYkVDUgHJeYvrIHSFHwOo6X+Auh9+
/7Pp9KHOWj+fRHuXX+A+NAIgkbYwZxbd9ONNRbvkfZEDUxxDoS44PMzHxdIT
mW/Ij5XGMvd4Fmdjni3LRFew06VdzD5vgDccpWEhp+af37roi7QvPyD1cGHB
N6tQfwgSnn3/N1ZtZ1C8RNePEDFaFjdHbZy1FJ+XgauTuIM6NBnTvBWOnizp
5iepCRd46Z46oq5E9EalvAALk7kmn2GstvP0ZCENDM/E3FBfB7MPQgjsQ23N
gCY0jz5D9iDWQBcTVFwuz9xh/q6DUCYbAOmA3fuct+1nmBpwhS0nwrPWF6iz
+vwwaYxgGm7NgHbrwHwzU4+SyafZFVWc9DgIPlQ6LV9w287oqnc1Y1EMCTvr
ngad4Ye8KtHg0Usd/M+lt9YKnhJ1DWn8Fw+MgiunHIqtZRN0erxCjFM4+wFM
wNtTz048ntIP0UTGLqVgPSPsRbf9H89ftdy0T9xfaEPsYq7EKrlWs+HFahvI
FjwgYvYzbYIxsi/a8XngcM8hsHuBNThH6WvFRPc7P85bVxKh7wx4nrtp3HTP
GwA9U5xiZ1lP5vJ4/OfNp+bL30qQ9u7V1Ph4izFb5f6nPlKzoKoNEiibyDiF
ntcITbpc6DtRsdHW72hpKMi8rsFEsKd7aW8wH5VE35oOvXiL+GUBiaDEVgxI
oHhY1Rps9voijbzzSnIpw9LPU9oA/Lb1i4frjxtljViepABGxsiOhNAS6S8l
q9D9/7lUcdy5SbeDHJO3hTjSw1fN+J/8df0nvF0Z8fY6nATxom38+r7kiqfg
4gDHe08TU4ip+6aGd5OKeycxJylbZaABfiqd66OMtJnJ2KptPvop1MIMX2ai
HxTcUeRAM7bOJWF5ZTnFeO5vmQC9tqdKeN6/E9I/Dw0a4ebPRL+tYx4Z3oVL
YO351nhSimcSyzb8wlP+e0aDqqeiolJmhmFO2sejHL8GEtahcpZK70HMkv2P
9yrgkNXzkVjaw89w84po4Qd7Bjr+JQadqxKmLLcYCkylW7xnnelNyEOKvzyn
MqLAqVSugOBgmfSn6eJrG1nlSVi2ylNmDl4Jyvs6bvWKKgAmFyySQQs13JEA
I3dZINwT2fllWFfifY0UthayUBr3ne0hJJ7pkcM6rZLPYrqeAkOEmqm/0+du
ZOFCx8qlZuOjRO5j1urpSUN8x15pQnGWjXZzM5BvXPOPgmBilTGRItUCZeGP
xkZQ3/FEIEN3BpYceYWCFMKpJoLsy2v4SFm0nxvC+QnzIVioz6brhEedux+0
C44da4fO0HJhTq1R7LthO2tKottkid+6z8NlO0L3r/ojedlDNP6+86aIZtyo
PilE5XPcconRoPSByXE+gK+9WY7jZ275PKojKoQZgHleVeJ9xKVKHnreBOmR
qjqdo/N1zqO2S3d/kh9DT6xi2VclZLwGx5C18ICB78X/3/6Pm736FPv3zzxg
IFLH8BDMw4yZdtvRMNH1IVdCzdmxDFKie//SQf5nea67wNe1ra+aXaK3LvEO
bQ1YZb74O2so6Ur45WpY3oq3qOybqjCx8z23FST00AInz/bupC8JAdPm7IuN
2NwsJF2GY/zaIMGpIAo92RDHA2FB+KGAS5ckTpnb5eBRnUwu6NN5PNC+H9bh
gJhjufIVWyqCBdyxOgIQKXd2KYNp7Aim37ltKI8MHy2Bg4JjJjBse4LgYNk+
i9kwSFGKbP0BsJCGn1YvqQ5rI89SgbiF3bnRY1FUxuzMZ6YFOlQet0Z1bYbI
Z6b7Lg3AlnqtTYgDOni9ug9aJrTsBIWPY0NSPZ/hibUnk21bN+gGuNOK8FjE
uvf9ZANeuA59hgQ21juOm47tAvskudUMEDGoj08XCwb0RT/tGMKJUx9zLCpH
hAIaVSN/j70snkLzMxaNt92yBjHFium3uFXUAZSo1s8a7zeVBvf7NBTeHue7
oqlXJCuxw4IIFHAN0JuxBIkRkOveOH4K1ch+AdD5V69ennRGlBJHx+Yd/4db
wZHRn1P6/cTuRTMPF5q3nweaMjwwbxlvrVQdupAhpsdBzzhbSkQnu8KM5+M5
lEXAEz+Gd+xGNlTz1xQQylOVHKuegd55Nq0D9tEOwxwvRbkzz5LFcwAnHw0N
HCv5D3pkA9TmbhFZn1yB+q63SO/BcrYxApln3R0e2juwtitvCAJjD+CF02Fs
Ap+v1RH/8e7XLjIYnHTB9ALXb8pGDwxFsUyGNxk+pk806PDCwfHpZvoPA3gc
EXISJExfLkWA6MyEOuEDKCGUxeB5BtLj6DAbZCb5WcJWhHZIVddrGD72eDdR
jTAhG8qE77B4goqMG+zHvtn9fpjRFUW7xoGGwcL5Od/BZKsoa2p6fUhh81/3
FOtDK3wcu15LoLuAGCEZaFS7A6azcB4Cw89qmqt+XzUdvveMXYGNjxN3jN2F
XPhE8U2dou8G12AParsstLqQ7tmNevhgjM7sH8LU9+aACvjL8r6XMj7PPTyb
VyUSIR8eEca8IGbXy4VGiSMygZyktVE/INBhKu97MwVVN24YBOaJuHPuS69r
g+Vb4iMXDJt5y7gBtyUeOgq0DJARyeGH60en2W2RZ33SxX47sLjIMw42b7Hj
+wi7a3TsW58r7C17DLkTu8YLnx1x5I2/cmRP/0kip3AqeKoQiDXD0hIxe5bB
sN2YAiCglHMWBjxDfp2BpQakiR89YtbSXQ7sVd98tYfOzqlKz1JmE4ltzhPz
zG5tm7DSLn5kw7bVwWPPc6GZITBJ42oV5VvIKCu2313YSGk8fCN8qt7EBkHV
sK2HW7WB9uU/tiFf9LcH9tGhQAc99ePOPRcWqyhRbFL72cbzSQahPvRNccYD
qndP0/PJgLe5CJy2ck3aZMj3pEVMICafl/LoGvbDPcM4QozM67gdVZj9WgDb
g56TTH6IpzGbufXe2ocHH3L1ndA/2HBRogxMWoqUUwVbgY60Lw5YtRfg8W6V
O6NYYUJc2PjqsYxUfxY2QBvN5lFJ7YbFAVqXB87ejGhQN02gTIUhiR0zV8jU
u0a2kZo95CyT2BBLB064Fgf8fchfuc/SESl1PNiOiWcuW99ogGwZ9DBH3oPW
XAvqD0wLy1leiHoZ7iDmIaCT7iQOzU/t7TtqBWWOJAACujVuOt/J+5IccdwD
mWVALtiwih/cf/jwfka4viJpa93XU58+sZ6NQHE/14q6HmQK7zhbplorEyDZ
eqhVG86KZfgj1FkXEQp4mCcf8OxdfmMU3m9o62wKUNfynEL8YuGBP/SInWbn
OdPOu+cOJK5K9YjRS8/FJq626/iSO56m7R7P9SYCp38CyuOJZ0b6Rv+Mqk7C
d2u7hO4lOS5W4qW/KDphgFN3u5M0FFca7BAK8wxbx4+5Mr4oCmoAvTR9vAoR
lkHz3VpG20oIiTE59gpdo8deB0wCLtT0QMzNT96nq5CRBTr2Q2/21nfCsw4w
QP7YlEGMLUTbFuBhdH669uE7xmoN1psUImGED6hCGdy8e6K2wzvFvQESq4ND
IbQLVcOzNHH0cZtduI/ld8KrOfbEjeMyW1ONUiLAq6ZWRrWIM3WYa0bHrgNt
5thX3R/4fhqwSh9JoAjYT8UUXERpKHTXMpZpkCawiK7XHZI3Q5x7uGlVQEai
vm32w5XMkvZjuBx+ipBtmtKRtJpiBOpUgHgDPtklN/twqNYcypGDR1Euu9jC
P60rIfV7iwrbcAKykp3tZM5AUQoopSaED7toimeiZX6khYfudZyLkMSa/s9+
wDOyuOKq/IVDB9p77uwF2oPcZzfuW31JvmLnzbdBB5K7sADnq547V9GcglOj
SV8eYOaXyecbZVBhtGJz28lp7ljzsXnqYTVBF5LT66HxSUpw+F3otVxIeNR2
f1UkS2KGKnMA+0+O4G4PqkV47uWF/F4X1bnjUlF0xMICw4d60B6ZBqJmjvzj
fO1YgIv8CvLTZOHiIRpUOwKYCAAwvIMmOU/KWQlCtVjD7gmk5fT6h4avVziR
8/hdYlkpISKBV151Yr1LQ1Ni0cOlX6BT+AM6ReHEDvpKWTkf4jk21KAAkXJW
iwOthjcu4o6pMr7EEVc+UlZjqLXm3uD9VtMJEk8p7bOwMmAizuTXBpGBv9qO
fzb3iovOvreeSRxiNMFA5M7cQfT2DHeJ5k4PkOT/uarGhXNawZZFnUgX2LRC
A7P/JZmX7oTUG5YvztAz9b2yKKL7K4HscjCvol8EDiwRxc9Ip2Px3xwnGIt0
ySWXsAOfpcJSZtvhWLwSP5jM3tRil1l2NVtvZ3SbL2T33vtYKZ4iiTDmH8aY
B5LZMXbq/G3MKzOwjBfMGCUuje9SZ2zVeNUXLTNpjCxu6rH9/sVWp5X78Acs
sCFVR1EUzSrHWKb9Xy2St2gjYdw7+YRhatY1Ph7F2mxjuuptGyqgA/ZdosZY
5a+XnDNaTnMtTN2uJNzO8hrpuunvBdid4ixuJy6UzmXuQUSLxlwvVIV0Wjan
BLuleE+cM82dS3R9vGIbqZhmMJTF4RJABIMuqczU3ps2w4e7NBd5nQMjH0sp
bAMRA61A754gVq2vPpielKjNF+Cg6WMh6vlmHy30jpe4oRLRWek8aJGiGPkw
SDqFM/SyDUGK82etMJdteHL6sjfWZNHgVAoA6w9tS5hO+ioNQYAh9xox2bE5
ngutFolbxzPDa2Zsc/sAiA2P0u4jDc5xUev7+6Bx27GNl7rOSXmK23/SEAVA
RjAxgjh4aHvDDyuuf6zdnzWfLUwhACTtHeGkfF74tMM2xgt45HxctXvIwgNd
yAwsm3arBp2e7RduDzS5ESRzDYA6pkTrHFiQBNB0laao9fkRrgc6lcSHonel
rXOKQWyJrumqfrGdgdc617vFK/XEnRYu2aSVPxnbp8rkE0UglEnUkgNC9R9d
YAxWhfnxdIuHAFko6QnZqtcZTro/CLre+MamSNhjYACv9SU1EdmErsZ6FO37
f0cE48nr8ZYpBaxzo3LIU8OtQKVZSlKXOCYL8qVGTYrC5gsuhXIUG+Voh/tq
/M30vzR3Wnd3QL9S4vSByjVtH7alZmdBAFy01wqjnvFWTRRX1GHsOO4yJCua
PSwWsmUYivsxHlNcY8tMzmfwnJTvpoCRPXcrKKBz2pd7JmIX6xKfO6ScHSQi
Q/K5urqdst9OpLFaYXMy0OEzLRLTPzY4DFZaob1NKWw3Lm8GogdbqHkqr9y3
T2NJSVg9UHyZNZ5Wp3XApthQVHFwgwqgPUQAUQf/jvbhyoVPSuqMf/Wl6mEC
QOKihxa6y0l9O5lQOQo/OV4A74fD1h9QZt1KUukLXj3MjmXKG9gMNSmUDg8s
I0jQNScLw5do9wmi6vn0l6qACUCTZsoNfJ8FBqe4NVdL/OtF1hU3kGv49NOn
FHlRp8+HIDWsynVdtHAlzvq73d6BWJ6u67yKXtvFGn+TLSfZEjVMjbX8GZoK
0hZr6yrdyCK4tRh5vX0yfQg+gIiZtLBevdOsOPVPEb8qrwXbVd7M+FltBHLa
ybKboOFV0kPK7RMbO3LfwTANBjvi5tKoh69b7ev+qsjMNfX8u5yd2pt/bPRV
V2W/0tAKIwkGVot5uDegIjYI2MbWm9tY4hU8XbM4wuLtXzno2ek3ZaRHcYSL
BjlQ7LP7Woy9da3UodNUfk55teoi9pLjeefVxzOHAJp4e4P5Y7JlJNP3KWPK
CFmDRZNihp0dsGQ5CYEmb+z24ej6sv+NuDRGOEKeNggfUCYtmNMUSPNeftg3
lyJpw0F07ZxUeWdU7vCt+gXweDrR2gMu/sCudX5lc07ox7H3CCBkQJyEtMt5
CoNrknqYgZTYlJLbitH0tcFt1sNxAEL+k5Rmwwqpp0abTaeJGGswMeOt8LCd
UcP9JalQzbCNfhotFbGxWE/TkgeLD26mmJyVsQuQnyik/a3FtfESiBt6jpqA
9bZeYBUTSByhCrdFb+ep/ELzXEKqQRbc9XSobdgl1iXioJQeVrawkpBV55nk
8ZGcPGSusnacb6q4nFQ2fOynf1r1O3+ktW9wheYJl6PR3zSJPwESEmM2CpUs
iF7nXKuMYtKc+vsEdrQoZcIqYBflWtEhp1A8Uyq9H8MHCr6T59YQJVHgfFwi
giqkKN1rgK0T8aqBElDcv86Qdb51Y4g1PvhjK0UsLn1H764ekMjmQGs2UVFd
fjXGeilmk8yx5fzwUV80mjGDuVvPlTy6FEdfoomzuoM3lxv4zGe/A2kKVvGr
JsYG/I6NFnCaRKkqgnX9WZUBnoSijyHikm58AqmhXryKFldcZ1xHy0iB20+V
DUiv3z/Y5V+JLswaz7P7BiuK234iz0z6sdM1sYnhqeUMajBfOgMXid3zReQ8
3wpEExBpOIVnBV24XE4I/e5xASKB5la5FmruaJO4MXMlyNpsqq+6GezyX6Fq
zMvIrgXmlLXBtXaD3TQclfiSAFDG/Y6cAiydcpOVpFtl6NfwU8vKpkl8Jj5p
Nrh8uxLpjbzHfUri4DZ1NX7AzRLobOx544GmBZx5qveXcimp8iqIIRxhuwCq
2Mt9s2H+6+zBiZXNl34g5iZjkfAecJv7+hcFtD2MUDAGTdhQPXHPsY9+BBye
liPSxdx6gvhfG5RcvFlxlymnvvhaWbfkiXRdOKOpB+/4jcVi2LadKB8FKnzs
wF4wMTlFtt+c6N1E/yIzK5JLyQYqsNJcb6yQN7NoSqjKWCvqXBL6AxyRhGHZ
aHakFAczmJ6p2Gc5s4WKmqDY3aqrRRTizDeTZ98trVpwR+Tkemy7Rh1P89Jj
K60gU9j2dcDcBxlGdxk4KA8KTtxiZl3MkV/GESTTENKjyPCl3j4cCdqa/rJz
laKIGeKc/7tpl+8GKmvXHBGX2da1sa9whUrYCozr9AB8Nyz8cR93/7m4Nu/a
znz/HJrnPsR+T9BFGlx2tXE10sx+sxnpDkvewgtEPiPRVyVhrZgxbCQ3VHAB
2x/CXrVRHqzxzKi05457OmYu/fDa9hidWGId1iXSvO7KWIE5E5FKWYZ/4Tmn
3891NURLJcz/hsf0ESoc8W5fZrya8wy7HwE5L0Djhj2G7T6nAoc8UQi8hkkk
/UWQiZy3E55uhXbm5yZL2Izs4TeR/V/FDqFMBfbT6NwZYzOC9vtjOPevZGgV
zbXFb5VPdy2CwzkCzFtBbW+V6fBRcHks+epIfreCxmsiWaCO2CK/Yb0a+5nN
syRLr1Czl1J/B+iOI1V7O/ZGQ2RusKA1LqFTfgedZby3/E5mqh0dou7mUgAI
b4ZM6Y2nN1/064a1Z+QazwtVVcRpp1Bl1car1HN3e32SfB05/8gikaCeFzSw
poGeDiUcmkx0+sSqkwMwpaETx6q1h9ZehD/h3+z+o0nohr15O6K66ESGMxkb
1871XEKUbNN/S9hVcGpY7Nmvmy+pOc9keoPzt4zDCMBlOY7Cm5J8T+EfdnMB
8DaRGD6QGRgJKS5DpPBUu7oaGGTf4H1OQt8LqkeU3i//BXzn9Tp1W4QLNZqc
SOa5/OXTxnJSKkC2dxmojamILNPWObyrGGjjZXOhjBSACimgNS5moBFM3KV3
tSPtouxJe/x8NDWhOQc6ncKMBDWJcoAA7CWCrtjvxSvnc3rWvnhA3y9Ky6KQ
kSfPfkkC2P21xNdeT/plrx3eW9LCpxriC+HXWtsX7x+//f8yvDVY8w2VETlF
lbX+gi6ZLI2W4ouvbMTky+zjGkHeddzG8TSK/QazHlfib/dR9QZEd5BI7/LQ
nZZposquWd1qBYjlGIV1wI9KcBmoaA5EgOgMWEFswE1TGBWf+reMwTiN/e/h
DrIm4gohfWvNrhd2QPU5lElWqYZ5SvIqPkeDxGVmCfYW+7bHBzkOP+OvqC36
Yb7b8T3szAXk3F2WBLpF1gnikAJgyYJVf5UMu0INbpze+q52YPO87xTTTD7i
qPwyu8CqhvIsWxYxz2vVCZz7Niymt8LnlWWjOU/rE1eKqIsIH91GbHuVTx8K
8SV+6PdKI10LScMvMgH0VoOIkZ5SVMC/E4Ogicvy0Ut+FW7octcC48rtqo7F
diH3bRzbfP59gRo0AxLa6BEO++BleAyKrJgUwxh4TYs+TxWW6IVHIAuJISaA
yEqI/Mm/bvVKWxo/Zug8IaefJSn1F0rr9cM2LT4qV8sSutBGIT+LIT29SidG
D4ecJJ181zSBT+TuTiIPmko6M7EQLQHw96KEzzIR3BPODTHKBAW34VsKRCm4
w7xpbuKHMuNFqIk67ZtdmvS2ai7KY7A7FibyIURF423Rv97Hr/YcEGalQzNQ
SjPnnx3TAmPJ6Vfqeym0u9gpFhUw6cwH4oIqKNb8zJ6M48caP0wnVD25A9vM
7neYWeLHxezdsfKGlvhQgqUWKvZFJWw0soWLOYTrKTD7gSY3Wbjk9B393bq1
Se17j/3unmoZxyu8P1SHSCIeTx/260wVDwRJBxLUQy+etDjfUQwtjjamn1rM
MEUIRxWjBG1qiKiBokXv6c8s/wnx7TpVKF77BvG1dI9KVk1yL4yvG08VSNWu
2uIAFmD1ki8OO70TfR05RNLz8nBy5BxNFpjw9h7LLUfgT552qsnovxX6EVtX
tzN1SgIboUmiYbRfuz18qwMLh+RqC55T+97AJurt4/W5gBouQg5xsm1CwJbl
wN0v6OgyqWZekMDil21h6pjVT8HR54rF8yaTh9D4hS98FtztBdQg48iQrk4r
pBfgwzx7ETrJnjkmL3mnmkGZfWvSBxhHsof9IlWzU+1ioIX3oiDXQc1QEcnd
H91Dc5YOS5uKft6m4ROXkFXrvc2Y7u3BalEeYtmZV6p09RIHU6nKRjpal45j
ejkt4rpVB0L6/nLrBNlVBzMXqsKl2b83y6gseMKK/uVQygn9bJiuT4hXAlor
FM0eR4Y8xOXDttLt/UyEsq8JiQ+gp6sNUD5YZ1EwennM1bHz7YnVcPSaH64b
d2p1jFow8VQ4QSxQN9NKtk/BLVKXi5MLHh6I3g1K7hWGFSUweWg+jYIW9XES
FpZrR2i8nDt/5IGFG9zex79YFyJYNcl2Q1inQsdDBIlYHZev1tnRhEIaXwp3
8OMRwRbP8dmcJR9awMDz+N85UpY19wUTThb0PyFS6+zUdDfVkJ4ISZRyGr26
MiLxngkDy2TkPJXFjwTkMnvewc6TagScBNml+U7gmIutWrYeMtLXKD5MfAgE
S8uIhKUWC/Csxyf0HxySxALpJCOuxuUYWXLLhdgz/Toe2IurEy6GxZQdWRPw
Gbj8CFcgT/T7EKDC2SPiQ/XgoKWtiISzfPnXbJI2t1Q3yZM0ubzsIJYGhjvc
qtZreuesYrneIJTMtVh/shoTZUi07d5iv04IAXlqYLap1lByrqrTA37HZvrO
P2/WBsu9pxOadKW4j7q2WykBWhe0JNY03dgm2B65dlxg+mPJFJ8+4PHW8mKt
ZepuVPsBuv+oYjki4kH9u+OlEjbCe8fLxQH95DKWOY3mKs4oAXu9iMte6ej4
AtfvmNwEtIBTjktJ00s0ZvGE08G7lUhCrnQR4eWA1nVUwqr7CBTBYNiC0g6N
W/WPtJ83iaJZL5c07D2Nt5ENm4zJX8Z0ftwWc7UAS9V+Vu/zXzJQasHMIiGA
3ehSFUN3x3eHqBs8U5WzFrtPoKyLdmpg1Rnl1qnEyuxpc2IQCp6yc2/ByvNt
inUz6tqLOzdIkFu7hWgKc2BQZdefZlTq4VsHP7ZjqRn6o+CT29ZRMdlTpGGH
vQyWM+KDsaed1hLrJPKbRIx2gFecWXcYuyagj3lXQmO2RgqOFD5cwFUUz/NK
YZCp+6weDNm+l6Mhf6B0Ma8onqV4MpkT8APD03riWoUa2Rc34hnEG+s8KLD0
N6rtFPUX74CNT4ElFR9+IKAWVHr9Ky+3hsIB0YxdrlvCXIMmK3G19Q4Rg86E
x64qIBfZ7haX1dD7ZvYlf+0WPIIDmhVCTcXX0FCquQDiLXjw3qWuY1sWbb8o
qoGHsi7dwA8a5sKKUnU5CFF8NBBRlwCse84dg41uWHn6s3IMonbQmNwyGBVU
jt2qTaXaGmcdgJXv6QGCqpwvyIwL1kxUD6snIq+NqwF6fi68Wyi+PInqXIwH
wDb8qKicxs7A3tRmIWETzEA89eqN15sQp7czmmboSmalaMc9xR2wvZH4bUm1
fOyUFTTRkp5R/HtW+XRqE3Z7imRDYGUP5Cx1Yki8cpPmRxFe6qqt9seNa/4L
4MI/GjpC3xtAhNxpn089Pt0wmydJ+E4VHUCaDWVTcZvwZAie8rZacw8h1zDG
1W7px1HTA8Sqb0Qp6fwLulI8qMfRsAbf5RVzM3X4y9b6OSHfZRnjjugV3jfi
XxyDJbueECzfKx0GLm42TDQfJGlCwh4ZehJzEJzN2CnohxL1E1KZNF9c+0/b
3w7v1zHVIV7FgCSyohaWQG1U+y/15DC9+uvkU/IGWsHZpOCrd65BJrUnzKdg
ZOpkCwc3HuVX3Ex1XvkhMSaX3EhFiJWrep0d0aFOTsk6GRoJeDUDgNfEQUOH
c/Baq/OgTBugB39NhyebSN/u+J0oHmB6U370r4IPe8hiUs/Grcky1Q+6gMpk
GK1CEGewGa01b0t3YLYX5kH4ZSY8nt/ncqLyITPHBHCLwzZFmZaZ+1PZIlXP
16vtShpMYJRJwxdpShFU7mt2tJG7SdMbsUVzOLTSM3aRyXkkMFFzG7ftxjEA
Iz45UH5PRo1EZMuMWb3j04pPsLTq6j+FXPA6Wp1DCxMb761UF7Z1zlok921g
n89OJseLpWVNGbQzDPcJRLdEdV+B9Icc8lX0ih5sh07RkSrWyKFkXVUnlbPT
liXYH6AXu/GburDOt+IvTnaIh5I/FHf99/ORzyCCla9/knLZpyVUCG2/RUFj
SpQMttGg85ppaJbjWWv9QrKCtxD8pMptpo0AiZ3fvWQUaQvRrVuF1/GV4NIH
kJ3EgffKUd393+lDiW2QnoBWLDYf70uJhdAUWdkrn4sr3TUJStcBXXFbieMk
aCCf2vtYZBx5gVSrsVCmADzPb9FSdz6nNrsn36DpQ+cRVF7QiLK7srs0a2oP
fQO0Sd7tzel08CU/CQKjqVo63yb7wP0Oe8xaRZK9vP93vGPPhBwLTcYHWN5W
SXisHYnj0VdZdO5QrmCknInW1mWSHt3Y+uvoEzNKTtNoQDlevbnqAbxLP779
FL1bEPBB4+B6DGTCFgWTd+b3ES2p1tiewhoZU7ly9Mb3qcwsDc1yOVARNOjw
YHqH2afILv6BaETnF6PAga01KdVLoK5Jtd49PaHQu7tVQrFpyLqls9iG/+PF
5fSbJWmMmEsgc70BQ8gXjvFGJPcKwY2Rqmmjwjm9nKKPhfycn8rEtahVWhwy
4BGG7MKoHqtGidBFr5d7xfp2gMqK+noeRZcgWSTVOHvsyJKM7J7ewdcl6hJM
DAOBpoxL7B7uicXV27NR44AU24hqM1ADTzR9LukGszwZY9E7mGcZBhSbfr36
5+Ay3JnN25CV298NRb10/Wu9G1xzr71p2kP1XwbKlIgsQDdNAtVqx0AHNm7M
lF2g+wJgygPKCD6Wu6M+5QSrX6jVld4y/6k6tM8HL7hAArGH3B0PtxKJwRXf
OokIyZ6BNV9GoP63z6bpFpGar+vgWWbbjDnHk+lk6z2sRrEd3JfqGhP2tscO
655HSveUg7RAsxnGOawwAMPml4lMe+yecY08rXbI52A8EHug/xR5Q0fHRv2i
19s85kqysmha3soR9OSyJe7IL5MDhjJO//hWNEf5yjC3BFu+3eYANbI+KdiQ
Bf0rinaU8sEIR9fshIWxMdwqSFYHS/Mu4c9dPg6Fww1MEPdVPKC2nOLjqKNA
2ja6Ds71akImjIbnHQlRI67/+EMNztUCNoWpHzLniLuG4swpOpIh5jA+UhKb
RBYZEo/lSuNDN3pkbF730OhEG+LL4Fciqbiq/HIp504HePmAXf66FLfGzRrp
bOQqAnaexST8P0ECxMpIgDkd7JWn+HjUw3Y/oNxUP/FST/7FvpGBAarS7iIU
yjUfuwFe6uJezgNfeZ6y2LjkaImnASBMklc0YcWGwEC42SvDJZWi707uPvZJ
yEFlTYoESidp+6nGX3MsKzXBpIkWNCmA7ynPBDSnf6xFIxtTgwj/f65wHnHE
fnzhwPSJ26aiNsDV+Txuz3YFarBtnMT5Z2XtPV6sPsXoCWTnG3XNNvzuzjkt
LLo3V29lb1B6xWX2rlA+dpYZkAKpZTTidd1w6iOmWDW0dWojpXdhVbmUQPLo
sYXtsCaf5nbakhPHG1mwhJ5fk3QrXJi/42e1i832TGsf0mGaU/5VN58bwcmo
VyN61uodvKBTYT+/B25Roy8NUpT+XNt0BzEHDgNuhQRN3Jjw2w1Dud5W70ZB
JbrAJGFhi9mnv3QRr0kFASSE++KDGavn8WxwPLVJMuW7LsaZzT00KsMuqiS9
KgmMhpChWmDM2m2QPK0tHuB8Wn3mQmZSiuvOowdAZaQQjMreETcm8BPIPOTi
9f9Nm5+q4SP6sNh4ALOJRnSSx77S5g5bCJZqVpzIBkkVRmbtYkWN24TicAI+
YRBkwa3cRxTsnu3MPh10kCt7fLIQd46n0Gnz0zKEdN0kr+9cNa1a3t4cpjep
JgV3ytUHbs03qTwHj/AE6By/H3gWInjTMj1AvlYKyD1mFfHojppnPLHGJLcx
3Ud2jMetjDwbIkemnn5j0mX+a9IPLXI5wx3HYb2mwSgK2oXGMGowW9/8FaVk
bCQNzu/Zmul2O03qnIllVk6jebtp//rWdEWUrfxlwxwfyjdXD+rnv07LRAC2
bv7Sn75qkk3fJvmSUdfm0L+xUW/fIYbVthFryKX7g7lzUiriP0zjA+xazzX7
ZPVamNs+aB8QKyOwkZgZbR7XnvnhrNKrM+UeV1VerjhltczEJ1m0OoI3vA6d
KM4NZ9fF2RTA5bQNvCC4pI3snGhCf7htQDeDy2vEKaE3te2PqnScFwnUt8o1
Xi/IeZcWFkLiWDLfz4Qjd1Wb3pjInqI5CzcNfk0FNz402V/4E7YUIizHC7Ng
EYm48IYwzjAP0UgHuR6+WMyKm8OZQ3Gx+8Vpgr1nc5QKuzpyCYx+A54g8K53
6c+8mWBsi2pnAfX+0NRGxQzKQaIqWDOdTRduIDANvsCmfwCHN3ZccyGsQU+t
2Ltb0sWcikJt1QZoMYFDeDxbQjTfnEpbmbUDC9QI9Iio6+3irujx6n2f1xUE
NwuWeAMMSFrR7mrH7SgYyGTVsHOX3aijOwOKz0fhZiI5/Dq9nCv3Na0rNgbl
A0DkyUDkMPuHpXwAruWHDhHugdfkcbFNPWtBcY3e4UIqKFJGCVzPTfBBPP+b
j9lRG6q1NUFD5DeE8VYWe3DQZlqtdi4NMtollluzYVwie0ir+w1Ym3AkZf5c
lhch5+gKFczRykmKfdEENUzpvNfotRdbHjMrORSCp7uEj0WaHKuIeAzP9UJg
lJli+zYHzlJ+/Pqy4KsNN/TUZUQC2exGJTtk1yBuJvZgGhcs9Bg87cz93SXL
GY0r3sJDIIL3B7nXX8UjLrpY4cPqcL2wzMvE3E2b0B3XuPD5oaBKJAExln/g
wfWSN4Ab4TXVc3skUfRMnI0h4TD1A5OJNCo3OupHNYB2QjXwu6j6jn9+ZwUJ
T9b3Nm4z34ohgOSyFb4BI2hIs+J8Gq/qC4YUVApN/8hjcDCCIrfyEHmKYZL3
SE6XWlPX3QGMs/3ctT4Mz7tsZKbR2nj6PTfQPK3BO/tQKwFkruRtoS5Bnb0N
RZQpfYbtUf3Q2g9Z54J4bc+5gokHsfgEGV1SAbu/PgtD+q9cD/vLFcuyvoP0
b2f11MwRQSyYBZTIRwTKwMG304PvglkaybXM5rF2OubEoIUmWkJAOOm9ZWLu
VsvxuKuVOSful4cLeR/Vv1xjfulQqL5VcuMFWjmtRmEBGXq3HhZPAH7WFPhC
gOFshgdhYDFc1fj+/j8niezgmzp+OB7G8K86vd6bPMEDHkf92siRovSiJSIy
Oi2br3/yn3ZLlebuQGt70GYLPqPHDCFE98jmS+3NbGHEqLPFHN7Gnf9Szaq1
YpBHuNGRPDy8CYAk4dI621S6TnWHF7M7eASTVSx/n4Kx+xS8or+BAx+t2Ea1
Ya5Z5Y38bg1FyagyYyxHi4ghmPY5hn0djXtuph65QDV90+c1uTK9RUhodtP6
ef4XrtcxsiHHkEmoIlDYH07z1PC43tUDSreCP3EOs4sixeFqtAez6Dg/vnhC
K7WLnUYJsazkM2+EexaeMnS0Jbg0lOluQfStl2O47NKDV1dTz3jTcIZRVQ2H
K1NBonzKluVSLVtgaKgXzF6OxIeOzshP6ey/zBQgTEEeI9Yad9bsqZFNOTaF
Wjuoy3RxMcxNv1y4WjDI4VjXflf12jAnBM3r1TbGIJ5NTO2le3Nd1eSQogQ/
wDceXC2+fl7KrNXSKjqhQUoYYepVWJxTTaun+RKfgly+QD1yNO02GtiPvZFF
W29ogkMf6d3B68Lv43xEPbz4885dnGzQfkQG+IJ/Ap6oLKOKaNOcXg+3r5mv
VVMBobE0nZOZr3tR+TOBmucJknuIHNtXWK5fPV/QVy4rmwLwPUQwe5w877Kt
ZZSX0Vxe4QvizLYTlYx4xV7skf0aneiu8iGonVMzyznYR9YtLhA0odga+oLN
tnqtYWvRMoFAVeIR16bi1RIy+R/NEQseRU+/W8JoLQMUUwYmyMCc/t1a/Myt
maZ1SXelPbHX1SPb3nR/x6HRzwRsIK0tiyrf6H/drDuRHEEgeDU46WvCO/Xo
/mz5otAYUlrMsVMAYFrAyIYW7VcN/e6WAUD3bPdiSHi6X6dDqb5qha3I65ft
Mo2CsxgW8dpKgejxANFdZstHu/Bmx9TwQNipxKv/TpGaW0Xb8fARK5BKP3hC
Tc+K/o/rFVwbfF6slp+yWn4w7MS7CGGyHwL7fPVi2UvM1v5qX+UyxTYs+6YF
TaplFftansX2MIootCJ8wZFgrT9F5X9YLTPGfv1sJ9U7eYS29PnDnq42Mc+Y
o3TYgPQ62ZYyG/0FRTe1L2rLUYME5deMUIcIzxtfkoHRROs6dZOyFxTgeq7b
2ya3CBHGrNAlB29LF5JjeltofOAFi+Q5R5YKHDopXciT2HK9ZCqb/ymhgKTy
A5ZFyfu8aFYgwupLkgjG1EDXA9M/8JSgnvRb7jZ6uQn1TDq+FABB0eJ4nxP9
QR3heOYYMrgj9nFy5HurTqB2M5uDHUo7ixX28m70iXy+7txhO0x1IPlMivtg
TT3e7l8KCWKkIGJ1qvnONXgaVJJZpwW23WM3Xzgv7tziSzUFbE+yvjvDY67c
VmDaDwzuhhIZwZ8497KejpFC6qUVQTY6tf6YpdzoIN2YEveCG9+0QTyKlZu7
hNDLyS9KF592YTRRJAspj2Z4D7coLCbyIEujq8NSoBoMOYG9YxL5sIobRDvr
XmaMKs50xVZWHSoBc4OAj213lbmSmVVVf9R8neVL0xHrZA/YlKm6HpCMuOj3
7/mOlPnea7hNXP8WqVbYUZZHCiYWqV+yW4ADcy80xVA0zF2xh1LddaESw49S
9CnVszB8ToHfJVfBpOocgmo2PBWYYJWrSSLhpoD4a/J9wCQjTPilgPCHnvNe
5kHVi5qruS6EwyoTT+nBPMxchdbP1kegaHvYmR8dmSRSzyBhe0/IeT3eFih2
FixIEVFTe9X1NHtX0o+cnkh65nIQ3t1Kn7g9dn06H4Byzcl2p0QMwcR8C+28
HB/ijzTCLpZ7PaRzsCEVq/oQTFI+1ACcHNyAeW080e7eizOnydFDvMZVK1R6
1pWCC5abAti/1CJ43PevYXUq+fyosAHSKkU6B0TwKdtGFhmkSD9RE9G2iG5f
X6zLf+MH6mDeUF5XYs5z/RCEKgb8PZ5wnrRmXJnfZZfeYDa7GIaIsf3saH5e
U6CEPmCCDPWi7A7fd9ND5fVoMip/h/NWAojrAcx6sqNWmV9lewnapJS+A57a
oOF6CDm3mwfRAu+NSfa3CZfXF122tJos/7KrE7dtI4jP8zeFmdLzf1uKV1Rs
2IUZskoRdGIOmLdo/Z+Ph90KYfHnYYYPaFV6fJ7h2oYq6OVYhWcRKCpqaxkI
2eo6kwdb5WhM+o2bd47N1yNU2JX/nzTrR1SU4sXw57G+FpDYCWehU1kIlyuS
qXHD4mpMI3O9BQaVcQF2mUeM64CqkdzCheGSkUQ4073b8NhVJ3bkLNaTmqJQ
YJAcEO6qivLf7XbeszFHaQaF1i2Nno1TFjDemy42uU8S5nK3IlePlvY71jp3
RQaeHsinKnEWfto4CcbVxIlPIx/arpE7nRU3YasXu8bKENLZFuBESVIiABOS
IFJXFoBDNNsV40AcfOlWuWgpyXmL2p00sAc5NhzF8RlzpEmETscH8IrClxDL
v4j9PKRlodADU37DI2Dyin2elRpI3EsWoPc8qpG8yu39MyKEcXAT9LwzvV7a
f47vU1FPV44+VN6ws/3qNTAM/6HtfZAIikuhEfIg6VadCfAJooQAqv+7l726
AyBNGMXsasPECbFsQtKwhulWtNK5kJOdL19R6wxHpXArhvnOEcjCknFpRe8J
dbEltamh/OPjZ7vVZq5MUZozLsLskRkuvsgmB1+qJEBkLw90qKKvF23IsISu
Fu2sO3QFs/5JiU/toH5+OzjWpq0wVgavtzVMUEgyhcx4X0FJ0rCqEgIUIZlU
SHyggCwdIhRpxz2N2pyHKA1uTT5MqPwbq7qrJEOveQpxxYyJLLFPIHynkbjh
Z9p/p0GlFHgV1wtJtJlmQankqpCdZ5DP5/t9svjqLXji9Q023q2oFOeqkye4
JxSTmTEMtwl9LlHperZuZtMoTZ0ZJgn+YfOpLWQpjBGB7LveV2mpxJagDAlZ
0sTATFr8VPfw06QRmQueAmawzKC+QAznIj714OIcAK5DhoKR1DRhOM9zMtBL
60tBTNrdc0wwM6Ee6BzImbIceZyMv8rNebpgWCacfGk7DoJUp/gvX6x1kgM9
okNXH0MHSthXWK7MtISw6SRj3B45TOvfDob0S003DyI0IXtV4EhCO0CH8NDu
3dS5CRSgmCWBvbbYlw0kJ+BwlkT9k0lT+nr0wYFd0hV90KFkP0ef/YKNP9rQ
UT/Iuqoz+sGkzm3UnlSCvVDuE05bnWSTsM+QPc9+e9hbBs9CI8k4Ju2JhZAr
PTd/pv2vnohyjn2RErSH2B6u427U/7JcmvnqjLduIUhoMWvb8CqUmQ7lsT4e
pu6iqdQ3FUmNFdGjKbpDmPb6qbSCcaAi10U5f24+VmMCIRuW8upy2hLFo5KJ
/tyHb6ifwHK2jG55CoouXUEvvTDSn6qlh/EZyrgREI1Tjh6bo8/lWKYM4zxz
zo45kqLOqIb7QbBuKZ9qRk65NKcXlFirVUTTn6OAgDITD5khmsFSpybLLf3i
HYDKBib/PKyL455ecEHoJFejbUJAI/sW8eS03H0CqZvoadPFx7/vEdVou0pC
atZAy2TvQdT0liVtKAeu6eOtx7Hnnl60VlX78419SlPSduTWHj83nUoCJHDc
2r2GdjseN8oiFx7jUPA91o7eEWlNN1C2TFuMcgQTbgpMk+tpfi0D8ncgE9ID
shhk6Jx4gWgKvLU0wRYNfNeBYMxUdI+VK3gQODQZcvlMUNPv7Mr7o0AnEzfw
+VjcTxlwAnQRWFYYuGjFcRBOM3+uOjLsqHfkoTeWOphJwgC+PRvp/R0jg8Sf
KWtdPGhpW9K/14Vp89QpY6scanQbmyexeofhIEXx8Z8njH6ZocKNKhSYB3V7
KNzQ3M4f6QjNHe9soPdo/Be8uZ0Z9Bf+sm+sgTVwPUGRMZCQ1ZfhP8WC+ihs
cJiV3q75hSlt0UQCQi409dP+p4wrZg2Wy3Kf+v2dX/RPnM9sEM4y5GZ2CQlk
t9MvhR/TCokmy9YUeLJgG1/cKO5XCGn/e6wk4cCV9aCJrfkQESH3gTM/kptD
R5fuqNvnhmG5gXvhB3I83Xl1gvX8LCQSxJBqkBSTfF1g9PBsYZ1mwmZtCPsR
4fSI5A2GhEltBtO3Okcsih5JcDU1W4Ta66bJcvkwkSEnqGD5k0oqnqZGHTED
nO0/b34MK4i2RB/Oaz0oC/cLu5shIAuKDgEFlmLYEUZehf0iqEB/kRTyNb1r
GMXRYp11cooNT0ImKxhNCy2iuiXRZBEhJ+YNS0jOsG/QAFEEQurSgyuNuw+O
Ke2AtSzIDwuHDC+7T4mk/5lYoQ7ySmxkTPI+QK3mLtviZrxX4Sc8GRNpldJC
NEYe7lu2eYyDoJG7DjbzXjHkmrtLfQ+KvSIF8HmkekUqqb7s3rGDLQ/nBtVG
kUS2gthP/rKggo1+hUvpTQrHamJtAMe/7QOYGOwClXgAyaVMJNybjcHgZEWe
MJM3XAirnxL6/dFkuo4NEV7ArgMhmigfjR/1zGxNNSoiujs7jEYZ9Malqd9C
aoWlB5cF3uHzEa1yookQMCanbX26x/qLPthIgtMhrbcb+LCLtbBgCFELs7cY
jNjHAHY7KP8b9d1FvDQ2oBFqkvY2nwc0+4zMmmsHk8+DZWDyG7iDbcO4afBu
teY9B1CVIZKHMYh36ochx9k0o2rWHeMHKrhZqlOdQxr//wDsEqHciHNwmxPM
zo+/NagRmmQBqxt5IfTtt9rFVVQpL8x8x+Grib/MpZQL7PWukznh5DEIvIM9
33h/fP1xcGY3VhodtUu5k1aoccLLw2GCDKb1uq/WJl5RA4SFZeCufnIYA9oe
XhW90FUH265t8VA19LwhRHD0GD/eeB279oDITB421R+JCk7AOEg+ukuaCTBb
+RkCsv3AIBkd3G+rvJvWN34Jb5QsTr2dePZBJJoh2iDngxDmWTABB2cYIFgT
AH5czpJdVxq0IBhrTLd+gzdv68Bk+DznXvDmyKzf6ldrzIfa6MTWSGFXJNdJ
5ueVrb9JmIHq2pnqoNuL5x1ablEXavBQrs3/PID16SoCJ5ye4pixjN1b1HTG
wYVDcrIEfBnM10Ov40pluVdASarFwKFBmI7uTK0aTOZL1fp912emt/XftiXs
Cpkt6/mL/ZDFhYBpHXvUzlOQEF7U7JV/QV+D8tFVoYCkaDr/HLl/XtOQJy4V
kXrR08DcVQNnJQv0oIsr1+kINU/wvyDr7dSRBl/kS4C+s/SirWnMkYkCIUoW
zKGyM6zMkjdy+02/cnTZk1bK7RIpCHbpQKZo8Gy7ZqzBor9iaNYCEukzNlKc
DwFsfMd9vkYQNDgLQM0w/IM28BseSScJmm+gzeuZGTPK/jo2QYZYOWwCfrDG
F8uQP2TFjz/ZEX+HNjptOPGYccsOzJqdEqBru4pZ3n3R9dNeva7Ur4oaq2OB
jMLl9CMsFr92iWlcyHOYs50ClxGOv+gD34FyLXO1y8V7GEIBgFzYuaEdZ+22
G8PWgUloGmp4xeja/qsC2vTyoEg0vYctxuNpdjCZWFhpOoq4v99dBtsH+RH/
j+a5y5iNMUPfGq5i29/F/PW8ipUjyHbm/1IE3Ig6TVNuJP2lT+D6yAMoXxQo
J073sqEIBck1aI4017GWflOzq6EMiMGzgKXDNmmQjmTkEKa/UVcEtsY1Mu6c
lA2FaLIScJqtmKZNpsccwvSe+CIXBF5FiKX3xpEAmisrqzDY9SZ68IdAd6VR
Oz2Z+cTIYpwmenOUF2+UkNJ6Saf4gzJ+fglwARl/2TQVK5MZLktHWj6fZSZe
n+u3njJBiLcEVsqHm2n0ZqgYyb7FI2XNojQ98YYncxuDn7hJKd2DCTnqJcXn
VNZOLgTRlCchmSenXu+lVz9IZTWICIOa5TLe7ZsB/2U7X6K0RDYGCnMIV3vD
sRK/rYznTJBXomatClXzR3FrdHGXIbAJJ2X7oLHMkOGxeQmzzV9UvZ2Ui39/
Ynqx8nX3tItNHL94JLjNZNQbxeuAW9EeTHPGUQum/vaFu9czfRck1jmfIUuu
FQjUs6jhf8na0pZox1TN1RcA3cJCHawd/SuxFAkDWKpNuW8UImIruguxF3K6
t0RTe2Q7Hq6WGHeHDCjfQqmAMUwDrvrn92+oYWL5qBbbm6+TV6oAvj/nSF5D
iANEfQhT0AvyF2EC/ND81tJSEAf/1ET+pO1oLkjWwFc1pjupI+3ywPGjS1eY
wAUF6k/V/tJEXIGTNrHxpRKoulVweXIk0CoYSpaMipmyp3mYYhUU093UjUD+
bOY3ZlRksobfR7dPjQH1DJlRzZZR4VsI3AIfdBJrSODwXbZy5qmSnP19uPuV
628sEi427k1b8ByAoWwtavsSK0jPQjnFSyeprjR8yIibKdTKrX2I58XqEwuz
bYIY/QwdCSmDnmj3N7UNQfUS2MFBEzu1cOPgbLM9pn7frCaW6l7TfrtiELNs
DjykAHyYM/ek4XFw+YU554GGyvefG+PRQkpo2e/WfEj9WIXXBg/yXXWcZaMb
7JBSgNleOkxtGz19GFlj9GLdQQEuXOBDA8O5epQsDliSjFDD3+wCjbWkNypA
oCpDz7XocrX2aUptSl0J6NyHVNBNRg/+kux5faPv9fgEk0Fm57fbfOo3Q8vW
Czfr/Bdu7D4WmqkLjAuaij2sIZGakGsTe4+vgOkYp5IEnqYpdeh7FeHAITDR
MDVdjHzpNXVAa2yiPrdNXhSSaBhxfjcIT86aBx04rcoARSuDR4pr/CEJo+ix
n9dA94P+QMDz5BtYl7k5oKE/2YZPO5eNPagfIfgUamuQyqHS8Fc/1aePR859
0RzvIlalUBJ9O6K0SUSksmZj65dWqnQapWZavUrP18DhkKnOHeHjN2STqdAo
6PwDL0A610HH7VjVLupRKwk25RrcJml4tZ3NnfWrTESjcSeYxKpDr18Jb4ta
bs35AY+Doz9mxE9KqA4vWZOe8bqDqQ1+Y6tt6NRqujq/12WrP6rghCroTYT7
IL0sQrj4VqlnFZF7A0mpqq0auAMtxON9JJ6tolZhV1HVO9Cgcacea8Ld4WIY
OsOnlDCZtXVuyUqCVqD0NqBou7kkNjuKP+3436dF2Nn8gSo9LnVlDwPfk6nX
f4U8zozFWZJfE1hpMKwX09wV4xmRkPA75jebiIepHTmOsqP86Kvd/mQat3fz
gOvuVe/05I+hAXpAeENoZRJo9sAK5C0XD8kd1O+5h8FZDDm4o1ktF15s556/
Ptyx55fFbQ1MHg5vxWOLtt8jIuUZsmifMsWXV0x8Xi2r/OXatdjaThZTDg2H
Rx/JMbUDJCzTUP0N5w5TEUdCA8cq4hqJQQh1KNcrpmEKnOrA2jUh9Xva62EZ
1uUnpxNNBNy56/ObBTcDvr16cWvXDGXh+d5hVcw/+FQ+90dgPl83lZEhP78N
G4102VWExFy089e4awRcADnJ7qbzILsyPb8bBXUzbbutzg03RU33qJIeJHjk
R1n6vQwzXpBgyjlZa8NtTvW/mhUz/OvxE6qOzlawh/iNnpNWk+8QKLbRBaeI
VWGeCRUrBJ4u4gwoxRt4y0HN0lyLZ2lWF+WOVMi8g3RhJRYEfNIknL6tdYVF
GIBi2tGunRN6kRRsIb2VatIht+J3wKXq4C4Z6FJBXJVlfzojjkex8uBARQhP
mdgqApItADhqGM5hujgjg0X5pZAWaM9gnfaPG1C5rhR3sEkHydBm8RwoE3B5
QcgMTKjCv8EVH411dwflqksd+HlZeDkh9jQyb/O7lG4cEtrP3+JkIyIP594P
Y8TDMU6OW56ZT52DTLDKVCO53cug5jPp3hClFeESP0qxJyjJ2+0KdPk0xLym
p5uLUsM75g3U43KEeL+80XPVuyi/RJimJAqLXH6ixKBiXYJ5G8d+AzbwXUMK
joQJ8CcbzrMqvsQtjb3+ioiZnuJVD0/XPH6uqy0Y1giH16FDvuIwwyyZ6o9G
Lm/tJ3cK6Kq1cyA605cmHZBP/QkawikYhcQkw3gqVxnffySzwfqnP9Gy6ti/
lwJDUXdsu8oWjzTJsQVB0g3SWQLWrIMGcQo+F7GryS03dzlyd/UAIeIwd3IY
0wm10rkGmSxdRdEYQhhnl/TkZeJOOrwKF+aFQalGx54t7YanxshM2ajjA0Jw
eoibW3rxGIdUu9C1XmK2aw8pvj6j82TCKVSh86mXA58ZeHX+jXJ4OIUGRQBY
kxlAsKnGdXgfnuCHKFHPjWv0tty6RRHnVOUJfh28KCF3JsVcPnD+Xml9lRqx
Ahska1qWQCJ0KtagImzGksJw7yToN/m3gTrNxc5R2rmq1NaqY8O5kbmvo4+C
qzjO0PFDfmc4onolTQVNFmh2MRHs/l3nj80J0391LUKNj0Y4DZT+qzhBHnXV
dyphpCFcwiQrB+cyhDhGL6pTp/Fjds2RiZmJ4aQF17AkkMG2tdEbaTV0kGKP
VUOLRUpF2NmxP/WvpOQ+jixIaEU1GWCVgywx9nde0tB4Q0B2Z886aA6RrIfy
UeasDOAq96rrJTNk82URrXz8pEEVRQsb2KE3hy1ifu0KkjwjHp5EyylVg/bl
bw67rEAKFS33z5MgFwZ6gmet/4EN1EL1zlUOHwp++FkW+/lJ67PrmoBQ/xmp
0eCfVUHiAXgH8YzeiE+XXa5eIX0DfBLPAQQYj6Xn0pAqQiXUjUk0YspNRmEl
Nj+a0RCHh6efslOSaXuzoX9iitDXKyQ5F2ssbDr8WjhBXpLCXTCMDqdee6av
Igs6UKz6OvLXlgNbRJY+oEW3Bi8pbUEOly8C3ZvtuIAp7eiP7EPVOJP5aB1u
Oi28MoeOhDblwi/l23G+GNvHIMrFWAyVlxd/r0NsAYbhHJN1AI0GzJ9SNFRB
0B628+xbOb0gOrm8YxQb/8F2/AJCgk3cKmvW90LgXRsV/d74/noPzB8dgFt3
OZz22SAAqC1qVEDMRWPBgGd16BYMEqPy6r4LiOlz4F6niubQ/G1MbzgtB4ka
egwLPGBL9G9v+8Vuu/Oy8cHpAtEDVuZUpMizMqigI1YINXZp/22OKljYyF+G
y6AGdIc2E+kDcT9ATaYydWP/VmobH0wguGeC38rAk0Pku0HtTG9cXqTzKsgM
nT081lM7v3yA01soyAvjLz/SwP+clfgccxP5dI2Uvwv5joOzHhhaR7xEydrY
JhiymuNf8GOU1GBOWRKU8ubczF64FWy1AwWhuoktignthtNyoSk3jcZ/r3du
ICtDOSnLzQQCki3QykBNCuBX6XQ0HLl0/xAIdshIAXz9ff7xmn+b7GdQfd9W
9TpylrS54JgswyxKSTnkulNYn2pllzBqiFLC8IqdYg72i993E4BvdoFAlpLN
UdUgxjRIG8rn0RhqH712NbqDjCgQIi2ebHxYqz4EiwDNH61LdjEA9YCxhuf/
1TuNYLBXxp87/FPtKzLr1d6x0PEY7EGMcYfBqr4i6i4x6VbJu4S+dlp6Vapy
/+YfCPf4T9H8IRChQzCQNitXhv4R1JkJn9MsHbuVsdqIsmG57Mb1ckxJn4xL
PHNiEUG4xVOSnpOwefHTvR+1zCiNRHGtoP4ndsd4q6cv21dNtv/mVQyt87Fz
KBw+uXNq0cAImrb1WeFaFf7Pt53gkPqK+LYoqLZTFr2Ozq8Y5mDRNKDxDsPr
pw1r6ij/dXlSqpME/yAwReemra6x7LLn++bILhL9c9IYstJUmEp56s5WU8RD
VnZwWvgv29jZGZyZvuzko0XHD4uqJMRNrnH5bjnvYbRhAkfLcvLYA2tSYkqd
LWPCZjgyfv9aKJY/0ghZEvF1mC8LnQSLUQKGwIcof24L5ExGoA8qsV0gLGIK
QqcX7W2Ore47sBy7IrsIRJNBoRv1XZkCph097TfwEMLFyL/JkhnoUcqvSGFu
1N0BxOsZXl01Zuqognko4m1y70hfLflz+RGzqCa3rHHf96nazgH0ecy+aUcS
BbdwrAfkRA4zD10PFfX/aqnk8AFYqfBMFjdeurHkXHTCA0JyAR8eCJtYl9Se
nYMzx1gNi47Xadfl9K9jRVyjotOAXleUtB97s+qKZkhmOztjaqBQ70Ej7wkq
AaLOAlD7rbOLyggIlpl/gaaiwPB6xPvWzkVL8oSruNLV6tiiq82SUXRcATlU
xcSBvLmONAPqTifNtI1C2wMCAzRqs33qlmeOKl/pJgamhdSSYkKb+/uffhbA
i0DBqPipYe/zUcu5efQCyeePX7o6B3GszUVum67Noh/ovHXdzAm200iAPrXd
OB5RH+FhTXTDog/dflDoeg1g0UFA7TrkOG8/Nup0i3f615PagHjS56ppOTD1
/k7G5foKbhpHWq51p0po//5V2Xvaq6F6XbXT1MaaQ/HXv9MrH7vRr7zRkHee
dQlDF7j4SHup2fk4rA+DDYIyWyqNurfaVQyl6QB9n1bHeYOAdfJlSvI7rBV9
9F8vn2d1eHdjwRhbQ1jFBiA7aTLgUfkKKcboAkG0G1uDzl5OhMVwiKzD/QYq
9OdESktp8ebaDuBbNGir9FdWga3jScRPlNZOx62VzGr7gk3KgH3Xk+qyXaOG
U9FEZ6nm/MgZCB/VvysX6mJm3/lPWcEl54eEE+Y4vf+bEYBtjxXJZ0WBmiQL
4LB7Y46N71w40lNdwHvQrL+f2lxjZybt4vm00pbPJFuFDNyck3l3XF+rsFJa
Z84YaPW3tmWr+9MZIykBC6NZIk7Ek7aCYyiRlTuiv1cdFExdODU5OdrhPgAu
b8VHdbvOEQHzzeL6HtC4mNv/Frx7Tf3eRJXwrSh6E3qjlMXOwaHJIilUeMHl
79mzuq3nY75wbJ3qMf7/bKZTERV9hCsLW3zZthce/ohUnBeGhss0GolfPODN
ADvZfdaxSErrZfNJyW2lVbOsN8xD86HunTf6LCP9zOix32GjNxf7KqFN24jF
43QX3++/moV7gXkhgWZkoFIR5TylgrQCvNeL8b3+/8UzYr4XhiM142myTNYA
AtCCdK0aTStOFt4o0GLbfe6/+jvK21WIxiPduGkOnbgxbJGKdC8vQK/mwJwO
8W9J8nenMwZIDKA0tMtCcO8YDcZoAm1V6gTzoI/RC4unfI4824oGUHQ0PB7B
W66zQmfCPLi0eXNj6hq6TScLQKScAR3laCeS5RXFoGFgpYZzeww2eiw7SMeC
yyr/2BFPtMpKN8bhh7minOyE2HuffyLUecCJYBF1jl+tTbd+j/6wEvKgLNoN
zzMsWyvbLBQG7yxMKRpY1yrTr/Xs9FJYs9Wp57JDYrZYYju+H7TJ21ym9AEO
KPuxwU1JcO8pZaM72bt1NWujMmYKK5M8XP9SUhHKj2peqE8UKfkbj65BCJJV
/eJO2M6ZAXRH+RxvWFRllr0H4Y+0Xq3Q4AVX1Bq0GG8Z8i/d/UDWpGn76S79
9wQmWYUkBGHscoBlU9Fjd6PoAKAgTzJJVrOuogX/Wsm5YmG8LPFaFjLPilI6
qZZBVVLk6QEUf0SPO++x5t8xX5qfHFvs535qlJO16SxEvQjuiJqfknNru3jN
cWcvMqYjCw1Hb2FAEJeO+Ea04yzCTCXLHRQsnL2A8TdGPPh5IlA/y0HcH27y
qIIOAlloAp/EedmGSCODjZwimmCw+EkxknnXAnEZXk3XqSTGMagYkyghm89E
DnB6CAxNEdP0Zdc0d8BIUUPAzh1AdgjTJq7kT57BBT2leVZNkWJPn/P5LmoD
hxeduPMzCXpPZTVOdvGwGC7UX7uuTW5sXg3k9GHp1JgbDrYmRLwUcuSpgq4h
1ovKH3VxCK9wzpK94apIWziwW0bkCMkhEHjx7V616yZuudU5jqS/k/+SZazR
xNSUO9YkdfXRU4sMephFR75Axg0rKBuhCNxA8L+/OiktGFhdJy1EPnUqxi62
YZIwA1YcVoIgCNWGiNUlEEjtwiyNAW4XS+yzmax6p4gbdv8U+mP+CXAYR5rb
CNVOXGlMuvsJmqAWUdTMQDKgLE8s/PK1H3mjNTwWWUsG7IH5ZlVH485d0YGj
rZkNyx+wRtPdn7SG+ZT+L/gewC4HCMmcZUN3fV+kJ6DFKJoqiO/G6MtlVczs
f61uTna+nsOpDFf7dIcKiF1AUZtUob/XrQTCvFhhtacDN/9FR8+p6cbLYZy5
RXlX0nJuuZQ2KkGMf0GWxG5LkLyffAI00lfwYBVxOpph++UcPxKe1TGRsREy
uCifE+U0pZWsHe4tFdML3PwrRWZVENpvfoDyrDnVINXoBaWnxx3bEAXncc2R
/hGZAVa7okZNEOCfe+O7wHwz3VUhLUBrb28xI+g1fbJtJkEYh2ETvoKDOUBO
fbxlQO5dUK1HbdQp3v3rEAzrG4s2LOrqoezBLh6gWT9JCT/y11kMh6XdX/t1
qlEhmtTqO0WBTzZrLViwVbvTcaIBl/NkJwjQ4VM8rkl9Zn59C7Yf8SK1Ssl3
LLM85NpUUCJBFdlTdxLzvq7LoHxYQdCgTVR5eXaqyUqimRdoyj6yiFX5fNWS
NcjaOV2XQYFdyFHjAqASKmgALCCBnHHiI1ElDeHQFsSoyNN5Y/ABtRhq/QYz
HVOG70tLy2JhIQIofui7kE7QAHuTBsv+EFhkpGvRa0Yg80GY/Poz7SD6PMoU
1U67FFJEMh7OVCjfGFvocb/uRL90nbWRqJc79OxVzq4wmi2fV8BaKUsV5MXS
2udhhrMFfNghk/FrcLyTgeb37Pp6oHJe0tupRW47lbwb447umYMcePRmdIAp
rtK+KTQyyV0nfQOW6DliSRHanHOKX42M5KsZbVXwJQq+SeQjYcY4m/j5/xs9
PZlrqwWw3QA1yjDBcvvuHPPyPfG3WN6Ml4HDd/dVOdGO6BCgIbsCncAg/z8K
bHzB8+dBnmBK1+BR4UcOJPfmMPRvNOqs6n4hpNo7ZJW6QhVy2vCF5/gE6uXm
u8E7l7hMKCzcBmmVBORFvGy3s/ZuOY/ZVLhiZGW0Wxp2u9wKrWiJczWPxc93
0Wn/gCUqFv8nnbcqVOIZllc/vm0QUCrt2m49m04dwiFtPIEJfOuIPWQsElaR
YraDmnHhS6FoxpwExpIv/7x1bGppDL+xa9YsEDeGrP1hZAgZZuWj+X+tubWh
oQd9CwzZNrFHAEoVKdqdnBclZENwZkYEvM8hPCh7tXgH0TfCdyWUsWdL3aZx
pEdyw9ZvxPoQHau00KNAR08K7Np/BEq+RCQum+Tthsbe59uy/cDEXa+o6w4H
XM9P6+RBAYCHw/bmiEXDYWwfF6myC1LXD1b2fMMSRAEWvDJdxVjfKH2OyTOM
Wq9pUjhhoVGfOuL2Nsxtc90oM6WQBlNZYLXPIcoZJ2VCUGsxHxxc2WgDwEoG
A25FnyzNhdIA9yDoht+mjzsy+ulp5nZ2ocwQx/wx5SLczUofOoYEyNMOhDfI
Zp3aAi1wyW+c0PY3ohjPtHMSEx7bSM4RyA1sbVIFKnTASbyZpqbJQCn1pxcU
IJQBNwugTxRNcO4Ren9GMn9x4Pza2357Qu2zXu2nmZnBOZH7j14lvMLX4rHy
uefVTGO0CX7+O6UgY9lw++r1BEktbcAlL7gqpe7UtHxt5FtFxfcd3s+vf79n
L2aVr0Y6XAQcFnK/xT0Vr7YkMgTdIavZZb+G4Ya0utKbRhxBRhnEkbd4pwww
M2pIMiRWf34xqv5iUPeAz6ODk2n8b5kiaIiJLNWaYfl5mszwIToyAVMuHupF
LLCKrSR0TLKzFTE1gIvIjpM4lOTbEkM17r7DlkHcudHGPDH0VipwLDM9mCX2
2i3bjKnemSK/VdAaAe3qY7TP2uMn56cXTaQzPb80gWT5Hg2+ZyrE1llrlaZp
lQBsp2863G1nYMDlMDvYf42Lg4nst3qI568buONjM6w8vtDVYRFAd5NRiLYJ
+1chmJMuB213lxpQcq6muPv7wkL2xGfnUhvY8r87u3spI5YQ0IF9QIrSM5vy
f+ZL0R6uU9dDL0/igWUuH8vRHQIPTnDaSnrBVCPgCdQOTiCtLQkeXO63S203
5enzs1H/muFuW5KLydi5vuhW6Jz3pKTXnXzQiGkpju3tAgrqyop8aEV5HlG6
/WwhfpSnLUEOedYidTFg1q0V2/Z9Gv2MyQHG/Sn5wr5PL91ztWGfDPGlv7jR
qrd+H1c//OmEQPtF+zuSV6k5v3la14tD7WqXZNS4QoXPmgJi4/Fj5hBxY8LA
hQ20o+1rv1wvgLKGE2pmqoMEOh6ktAQhWCgySSiG6DAE8bLnhjGEP7dCYZWO
O4cLEMJ63u9znfC2sd2Lq52eQJDAI25l/AfDCTjghwVFufSoYywe6A1o/ssC
jUX9U02ZD8r5bpCoX210bv8JfZAklpQvi4HP3QfTc7+7iGgB9n00GPBy/03s
4agu8uQcX+tF7FkZiloVtUdpPLc6XBSYQADUDr1K2nNJBRSzfGbD4KaDTEDE
fhIBNcJLV3NLjjW5t1Aj02QUTAbghz/PNwBDFbWU3mfYBC+nWhTNGYgCn80E
P5H2VoXwLVKqeENoGlLSJBTVJJqt75Ivi2EbWmFDTeeo/MAakTc4y1LPwdtM
q9AM4+wIf7U0mxv3ObY5SQk9VGFT8Oe8sl1m3MqAFhjNKoncSc5R6y3j+SAb
kdajA/+zlUs4zYJH+ueCnWpKuKB0CqZd6lAoWhVRE7kFIYL2no8IhiNnWyAw
7klNXaHgr3W2CIm/AJCSFhMyOOVjIGhC8S5GhBvS71aeMaDgdSLwcs+uTlHo
hvyAXZOAhXd0rxVoeGEl8C6DmbugZciW3QVzH1ogyVK+TXhVWoc+S/ZJzHhX
nX5b6BCBaRxlMvhmFZS0bSuFyvPZEvSo9fGquQ8VTSweKY8VccMRNAP9Gf0n
albdG4t02F0qitI5T/OlrwASGSDXqEdPkBoTfkJUgrTjSVBRtnXQDKuxdPDL
/ht8+/d+fQeI+r+yulq6aiUM8D+a9Scl3muGgUsrkKmXeLqALIQPYW6CGBue
qgjSk6t5RtB9PkVOTxW2XnLkjdcTnmIGLJsdX5PJ2sqkdVK/Q7rhcbabbun5
P0XH/TIW0bbCDu99YNzCK3VS7JWQDqImdtIaZXLFmOZk6dU7bRNhOQL0ArLq
2K2sXeo8CK3+CX1jgltOmkrtYqZbi9OA3MBfXiI133W6sRSBX/O9jYSz4fPi
+0uYY0TDcQUvRyQjPfcumSqNFl9faG6CoZFsHXtS+OJCRBb5EkjUyL5/9Jrq
LS+1myOu1fDXai+IBQhmKG7dZdbYSFUxI5f3YalI00N9QWvCNtb7+9sNgtnY
4JbMNcmZ4SG6fXV/B5blBpCW/rUb01k5NOwz9Aaxx2zydB3poQsohRxUSfdf
p5WBq6dA0BZocvHXhnOJjXCLBX5aWwmMDuL20PmORFCkNGs5Rp27MWUxjJTe
ikE6Z2hEW0aXYikakanGx6ybHXOH8ELUkmzdVeD6uyO1sygLrZMMgvitl4Bg
p6g1ByzlgUtzTRY+3tMrN6ILJEuW2B2lESP/6leUsJ4E9fk4uHHHJ+mnF4Vh
yVdabxfjAxS6Re+5PSlL/MI2URpSnXyCLN/w296ejWOUDZBPsCBBEMF7EhBD
Q79/vFpUI5emmIoKgyxpAre5lWt5xbB2wg1jE/5ojVALVWD/o05gRzhpIQb1
z44laCj28e4HOIVCc2Z6jRdhmlrkvqrrBaZnMiHOnHvmTs8Jy8QdMpt5TPUz
9YZsr+pcUfS1/P5h+BpnFDen6mABCm6sjemlFxgnJHzC15OBGjiNiGiJ35Oq
hWfjzHS4MxlGt2KhGK/E/VaeItyb3aNojQm2gECtBTaBuL1l1NORnzllsDIu
zn/sFHYP2tQYPIzIBxjnPogUJlS7/MpW1/Cxl2osnE6qo1b6BodwG9fHAZB+
81XJmUN2pxbg/TLblyyGNA+HTvsx46hqe+luj7WeDQwgukpPX6qm5yKvznH5
/RzFleedu9fSoN+XOUSgob8vv1Y+s6Mono38sZBcPZZl20X+PP27UeI4C7IR
13D7dHpEePy1vQpJeui2u31YJHzttq45hgtcv/V5gCcYWzAbZesEhA9D4Us2
3K9O4Gk3BF0Wb+hv2tzcnHNDLXZUH27LvTs+pxFdbSDJjAltAMvKW7bVpE6q
96H0MQiltvODc04sF+mA27g343tLrNEr6eRV2fI2xZMpTMi5WHPc8MK4tftN
5wUaPsaOW0VlmWWu+VU8I7h4R8T+0H+V/d6J3TspAYwniTGY6qL4d59mbcJx
1D9blOWOmKNeOiEQ94i1cCaxOm5LiRGn9cuid44wtO00kqXzjHywbyUedbcQ
PtZpFhQVPDr69lrSsv44Gvtx0ZGi6M+qbIXyHJ6K9P9wYpvAWGD5XR1uk0rR
rHYQv7FPtJd7jTsTRTxWeA3F7TKMh+BQkfaKwtaF9bM1qyH31VETs72E1qY6
1zfsEuPNu2ajisurrkClufKJ0wj78QI6yPiS9yx6jwHZaNvjlvSoA1s7Akyq
uzAZswaIazqxGvEnAzRnRiG+QXhDa8ZTJ5ki77QEcMZtIPoO9T5wEIy85Q1v
prB9ZEiAF/Qlc/TOrb8nO06kOMxo00hshyIYqvcWu7RTp9c2MoyLhgKLelE1
9CDRBzqdW/5l2rvlOucolZpbsNGwxi0Pp1YxPi4PU8aSiZdpb7BqaN58MXMU
YZ6lFxCQELuIR7gJnDP4EGcmEcbXqPjIveQJfanlprDaLZoSMXfOZqsgabik
uS7vO189EPPri/m64zBKceSlKH4h2IKiwR4NVimbmNJABaZxWyr1owkS8idF
SH4dqO4iBOF1U5mDLpcqX/X6ITkmJdiePFsr5IbLtA0jM5/4iFl1cB3DPt8V
RyxDcMEFAUa4nkTjr8BgaGilXhwngmP22JR3dVB/WdTtpAS49tz0I4g3RQ6G
MLZMbcuFadkiOWaymRmtAEtq0+ppUQ+odXp08rMA8yy7x6/vqRPwRLIgBgQx
7HsEr5QK2AfeTgPFikFWnJM18PMJIj8KU78NtkHhjrHpMOfOdxzkhIwfpAoD
Jkcftnr87Tbi555MdyYXgIbgo84HpvxVRaB2fvCQI5uq1ypDEKuWMbe0LETF
P9lyI1K4kUSxy0ynXybg5oinYUgDt35WVPJlpa3AvCVkvGBdOfmfnrbvngm+
Z5m5x7h46j/tTF98ZE+pAMLOgHa8JYtRa/OOjUWAVDDs0J00hBVwGf6MtSMo
suki1UIMH2X8Q5nSwHUhjkedRq5jxNAGuUYlPJdm16JoMNmWW6rC/baS/HAw
WQFDzIOG2DxANNGpVERDhjBpAu++B9Lq8QvhqCUtxt67uSV6f8Wv0gIBRFU0
mph6mYhFS4oRWwHVRA5lCqULQ2P+z/UKkZArIVqBHZHCGPgnRPFd/O5nG2Sp
JaYEnuTcytgwP+5srSpnwmkaQVzir5N1aBDE1aSztWQZd5iaUpggcSt6zpr9
RYbncTHznySnodiZqllnCwpIdISPg2Ii/txqCjf4mZtFARxzOirgzicvPno2
sU0s6F3m8zGh16h7bebNGPyck5RFbuFSLSogiiIii3Q6QlSDr4jHkvQuRkOA
fj7CojUZysKyJDRTFwyakuDSLu3aV4vam+EZ9uNjD9HGgYUByF7pOsTR293K
5ROXxuf8ikwt3EsSzsZ2vkyCjAxDPWyMiXRplorC7jbWZTp3QXDSEVXmZhsX
ji2w1JbYI93qX5APSTls4nK0qSt2kf61V9yzhCBjSD8mh+wPOkXZQtveZip6
NbhVcDiF4f6mfzB5TEknOzW8rPSXoz1Bjhkd03iFNR4K6EowILm+Rm3YRXY9
Aiul+UGKXlgFyRykmNQbJ9xGiIINUf2FC6jebig4rzv7bcVVgfNUJsmJNTqp
OEj4nAZx6zkqeEs8DC5/8daTuMHLpxkznjjBRkk1hPdp0TT+y5GXyy9OxBw7
rxk+6p0Toz9kpAP2agWTps9B1HDGB4KQ8w3Q2R/bwtzkly5yT/zdLjWD2w31
0f69x4pKjRe+yQ40HAvBlQN9PKNKhWQ8c51tug7kaPzOt41/DtRwNNqrCCXX
fhLbrYJtG8+TW/Nl9qw7KcgO7EEU0tLGwcaxKjdzyLVCQgbLqz+77hrusqDo
hEt9IaslrVMoU/eFIbV1+UbW284FW/6SMa+ovd7jTQQFXdy7E+c/DOobWKpA
374FJ68wMbyfDizhyQt3JMfdqXtb8uIcojua9idhGqyIe2kiLPtqwiFDjIl4
udXouxWG+YhUE3e2oo+8Xf93NzUWZJKNrh6pDQLn+LMEXXbk8oDAgY7FnKUt
tYfc+6B0d2teUBg4+zNRWeJUiry2IduqYar/14x2vU8CQo1qNf3pcR+Xj//k
WH5dEbIwjZAbHxigZBoiEzgxMgF8dbcBCw+7cnf1mdAZDgRUoDBg6yhlOraH
Z8oJIHtBKiuIlMxMX3g4ueENZZLvEVMS8sR8iYLUn1GM9napWRwN96kNjTPF
aiwSkuY4aKxAw0NoX/jygFYa1pwj0prXUxHiivmw6PIsIXJ/qiH3YH7ud1g4
wqbJfrIGVJPFGmsCDE1HsvXihVS/zUXR6QvAcfvWomjJonwny1sKFhydCNcq
tdxDPgjOH2qi/cwWfWJFwSYOJmZvNQCSYLjSWCOxhBK3akhHFu9WU+mtJudB
k/8lHmobwzs8ZFoIwM5tEg2d7fDb3B2cxJAOTn72lsmGL8swcOfX09VxLuAb
3H7ycy7IOLwzuovtJi9eUzB4FT7rZRh4pbOqBiEqLxocY5JVI1hAduTMOaPz
9ZaaSWi9Rq0Nb2nn5l/2jLV9PLF2fXyl1WQE/1N60ycGWtmXGCL1a5K14M2A
5mNICXrxZzSsL+VZbW9f6YcUnHwmn+Sm9BT1/3ODUbYp33MbT0arG+qEf0Cy
soI3JKEKAT02MP6QK0X2Q0lkNIoT0mKcc8LcQ1QbvMQT5Ss3C7agrzDbaHaG
6hvSTO8x69/fpevowr9y8VRcvFWDkQSIPgrCroDRXL/Cg+ftRqh+U76jr1Zu
a7LEDDxLaAMzUJiUdGGnRgy+nFeiSgMHfdKEehZtapqRN1LBCIfWNoiBX8rU
lWZCCSKAYccRCasRGzqWnC12j5bxni4LawsmRO7131+/yiO98vTSOajeSt+9
D2JJuq4E5tqV3gU1lUjCwqQnJ3pDsizOr8nJ6yxuCdqOQG9UkyJSaDvjAGPt
fMk9GJw2cM22SIimreKiu+KulzyMlINA8ep2aTQD3FXDvK6ZfTv9WTXEw08s
Sl+y+0r7otlD/8Jnhu+Ehpe+aMo5W6hfqx843xUqx2QjUNjuXR0jpiFNzwbC
v8LsoTvUCBh0n2Ry3jA/KlHX2lLS+WfnoZpPAp40zjfbqzHRQ5q54XNAEd7T
bsxJ1mLnZaq/wBg7AHKJUFBXIgq6b/CkaQQ1Bt5Hiy1f+1YC0DbqXwAgW17S
w7OO6qm8xwS6ix6cJQd/hh9QNP/B0v4qeQKCeA1Wut5QU2FqNTCWPTyULY3n
PuImSM59pKuyK/09kjhE+rDjOd+n4MLJkgVPMgeMJuD68aIkn+ecx1SooP+R
LSugKlPn+6MqsRNDyeFsDnGme4UZUjNN8fTiamE3PfvZbNtUdDG9he9XFGnO
iilsF7N/KqXjpf61F+mKrrlF2dZbeGDIV28PYh1rKKjY0LeVsvKjuM1n3TK9
oV5t9qvcF7YZIRwnpRQsCJEO4FZgQMgO5o34kXTWtjDLBYDxwpSXF9jVpirk
vKVVUBc4CUkGuXLtfJhOzQAT/1lhh0yTRvGqQdUz76pLz8qK57enA7f/n0n4
0lsRBA+Wni/oRMPsmNnL6DI3zoozsilfEcQnK9wK0lzCrS5GkoyvLaGQt+Q1
N/8Ck9sHMk6Xwcu5GAc8KAGbeKoS3uGshvoOk+aOYsYQgcSp6ESrEC4rgjBm
rctdW+8clxkBwi+Cq8Y1Ay363rg8DouYoAgNwgEZj99282OhAVAGgALOjqfO
uwLWc89tKGm1KcIIiJRRCzHHev8AkSGTZ5ApWUWeDMEdsBtXwZDg2GTrZRv/
7EkKaEcLO2egCOZmCPnFztU4UWNJWk4DDcWOxm7cAVNeYZ5t5Z2ZSmUGRuIz
dXvAE8/QL57K0/Q2ZDT6owQfKVFTl9VPxi4YKdWUlubNMATKKMkBbNbSdJkz
vRoW2sRngSu54e1ciJSXWDRfibEIc2hna1EhyAU1B9o0PO7EO1btvRsULcOl
r5qny6IGCZVNyqzDlwdJs1a2OBfc+ZDeoj6WNTrVVOz5wdUZBpGF3wFXLrCD
hbyiFPZUSvpbdkjdLc3cMJcjlHWR71ggB9NCQYs24xuFpt3Ow1o7BbYUfCxW
mOF9P4u3AfclZdJUzna/mYtXxWWGkisrGunTz2lyDPiRn0QgxxJ+/rlcC5R+
rkGiLhambq754BKKmA0gFxOxs1wb6lGqTsbQihjxRZdxei6wY7C6FWrqoQxM
WPEBk5DZcDnb+0gZUg6zZ6SU0ZPMR560mFYZloBL2RFk9b1d8iKYsWhNleJt
D+TJXyvGRZ1Dopx37vXfypzBvqu44YcuKRH1v9j2M8Z5mzB6xxOY2xqxUO52
R/Aty1YcoDBRCCXg+dk86oecCsFutD//wQdWLPQBXqooveW+NxKEiqJu28RW
OlElad7vYwMdEVZNt6WWBjyC625lMgCeNd9Qdoos47J0Dd9QeZNUqT027eQZ
aYmi4trSNqpagYLMpRHYc0iS/hl3rQV8JHadUroANzEhcVauv25+NBhGO/vf
T6fXCwZvBzb0X44Cenh6+ClyRJ2f4GpvutEXCSWiFcJyB1GiK9xcneuvSJOP
OTEaViuBa+pRi4esOZeYFPk7D6npNQ19va+7twjoK2OlGG/avR6LQYyNsVSE
ARIlxMI5A7M7ORm3dHtN3S71ESjc1K0sFJ9ylfix2u2XJvDaJsYrGzHVKxT2
YlpS+PYgfjwr7F2gzqGM9Nm/k2XnTBFLZC7KPSSvSozKGVomXBLnovE99p2M
Zdi1ZAB1ZbOBa5kFAF+BzqhjZcYFgCs/zpbMjU4xjo530IbWwBu7n+Do0n3Z
+AnQeu3rC5uTOWq5YnTDK2ymCAjocPtBm/hbzUW/7iofMHvXCuyPRiT84IJ+
Jq3Bf3hOhZWkn1VPilst01Ams5A68UOh9jMGSAw0G49PCFIGVCyoUzzc1cO+
GDnDKzrIH+auQoVv89Yz2yFk9A8937G7IIWVVRLFd9etWv7hvsLQnux958Wd
cKe+rY88pfG/D4U1UDn1R0TQFT52yubDYBkuLRr4rBKCG8KAMuvIdrKqPLmG
c2S95UF0JzKtglsPc5XWea+qOFzkgNBwq/+iEBoOpC8AXylhPNAj32hWMniH
gr8XGAZa38EJPtvQ+S6YmcBaoYc5kbdJUyrMiNraMmyvF1XclgVl4YT/Zicq
61wa6n+V85/qFzK6ko6kt8BU4gifVCcjbDxuJob18WHC0oXJ2RKfhvH5Srip
fvX17u8KwPd8mW4h2XF9GfKmEiC778P8SH5weSiUz/0CVPxe73NYdM9LNHJV
QmBtmzjPbWbvChP3JXd3xDYyrwtZ4npTG85JpYkH60VYRi14bZyUfCAHpL0R
7XwvXQj1VBaLjsUQhhNX2ZZbvZqI3XuKyJYmiEBIuUyoiz6XZ2TssaLi5n2D
rXeGGYXxPND8FZ9OAwX52sPlXBo5bb/ueBL8FN4hRTsv4nbCCHiH3uCr/pRZ
ORKGGuZlLsXWaaOvI9VK9kpZALEfGR3Mmz+uZZ9mQlv3df8D73CAtTqxY5jZ
Kd8QHpRMjEbLCteSK44Qd03uxr13ZqwMY3p8W3jskeAAuX+Uqk0NIVwC9LO2
d2bgpZh2h8VOAfR2OeeyNmGALshLaoq4vPB44eSSB0s+6Vic5kxbSWuKheUA
8qA7EF3FeSJk8FXUQMh3oR0TxwKSaW7fTzkiLEnB7o0dI+2LEw+U4ZtF8WR3
x6q4IYwZy0gmLerWZunNK6+dFt4/3jnpOBW8AHay/mmJ8o2OLUdrHbTHnf8u
MxqLdcjnWPtMSI/ngC/GcHV3T+5hSRQEgRQKPrJFqWXlU11Nds0NfyXhIlVO
ul2nUPvZKWeRVpAoIjXYPpLMmO44JKwS+0l27zR7WGB4sCqHOY0RNvVhyaNe
Q54AcRy7u+MLRhlfpMDVaMf7X2KcpLPmd1otji0IEUq6qRePRfU6NqM+2aOL
UkItubRePEKCPQ4uQWzKGZ4mc+9/aR1JBgVaVGcLMNRuTw5cwbJ+B9FlkRgX
frAFuHbOp5akD/RJWP9mkeLImKq5OUPbidbprdH5LNSLm9e06CStn3eETrIP
o3meNiV+55KVoH8wb/lA9q+UneQ6ewLUTupizdpj8NnMbHL4YM6O+EDU0ZJF
9W5poq/fJCwewNrpWFM8YxJ7UjuDwUBYyRKdItvPLhMQUhpVClZD4iR+JPIF
/dufNDkhdfw1vSCSIP/v5zrWCKKKmo+tNnEhTCyKo3zfdOpvEsrUoBbmJuKA
XYJB8pGy4VQmcNMYV2MQDRJjS61Xg5D9p+PA5mdFBCksoMK3ncFsZlqsD6WP
YbaFEzCjZEk6/LRFeI+6MiNQIjtLHGL/3WB2/G1ZvCkJWZfIidbbvsLvdrrR
gA2P+vsNejjuUmexPZ6nzTjwhJes/iOGhhADzFmSrUC0TpNcK6ELnE5TppVX
gSRRH7ZN67FrzLWgIX1btbimJvsVax8j0+3zSYyFV2q9Y7mye+3p4u+Q1H2W
lgAtE3l2258JZzvmSnaZMd5XpQcGtyFt5jcgbB/hHICs1OOKNerERdH7/CAy
19+RMtVxlR62uM7On7/lfx+QhMNw4YryCyvxKKuNlfeR4CFyIavUIZGpNxEA
xPL7Qx/fjRoLWHqWvHeuS/zpLg5SDETftm5XJej7HQCYg6BGqBUOnoBc6XwT
dhgC3sVKIDYVGqniqG+5aaTYbbp2QNIK79v+R3Qkn1KPfz/PxXR28OpEDgbP
AVz1mjN1RqqxFOfkMJM99EzydRX/USFWA7pkqA6JDpwLX/BFPkD7UnEuyukf
ROu5xxLM4fH0GC1QG1kCGwf786jnq7qfrxyThbf5af/CsiqD5u3v7xIZ/ZUX
+QtJpzc3VqVck49c504/nUZ49MUa2AroIcGf/cppX6uDj0b4QifvRHyekhKh
OlhE6VRDyOgu5b7tp+mB2LIKxegfZsDF9gnT2XwSGwZfE2l0Y9S5Cut4e5O8
FJAiATknfuvU5k6bKWO8lHuaGYbuEXw6xCpz2Ne8BAwA0MY6S6eJVu3A7AbM
Z85GRNtMw2SW7uCnV5aV/l/JN/pNE66k3gLJG3x5wqk1IgDX32g1bJYVzkPf
IV7g/Xysr8MYnLFgR9zaaP5jETvOfx1HNls8T3VZV8XWFxi4S+B4yro6fyGS
3bi3Ta0rpSWNczaZTnj/n6ow+uCBgwiHhHIM+zTrzxjWjJ93aEg35aFY+rrc
IIPuCBod4dh2VeUKKGQwuG+1PE9ThqyQeJi5Weu2XUOW6gGBE5jpQ8z7rNec
NBSo0mC7+XJVCGtq3WZgzG1WBaQVXixge+J+3BIxLSnhKHcsy+8uuAY1NBej
6GSaoYGIpaB1FjPNmW6g1hUC46md5SseylMmucI1JbMWCMMbRUoxm48nu/sM
5VtEXbF64fczfoWsznIn0w0K5fSD4vYnnbudeYBC4KMCcao7lBDNoehdbWoV
a1Raq0KEfyMdHsmxL0fAwZob6vrfSF6wQSiSHzLGAfyYbGo5EaO0O47p6wri
W2PLz37iT4lKXiR3Fw+2v3NKdDnnZ9pehaQ4a9/MUlXie2t369MIsTN7vjBl
W8YjAktyVn4/6b9uSgYCta6dALJZjSz7HMCvTtMK7qqM30xm7Pch77fWgFki
87+gsfFauQqef1/+exlgkqUDulVRbOsyWdTtWAnPtAbtQawHcSebaJO0B++Q
gPt/MoeS7M9ASqT6JEaTMDJpHJf6rEDP3zch6xW1zxtfyO+pO1roWlwqvItJ
8Z5GnuJLBEIMFJhkS1cFyBbS13UDDMdH8SJEl2vTVRSveub1bXvpnZFawVhi
gC0QebGlb5HZWYGi38N9m+euPmV4nqkJeh2MBHxcymV/MeNRt+P14gXE+YhG
zasr6sg8dx3hMAnF91j5Ksd+tGcWwk0CQSlvILwUYL0rU3y7skmzj+09I0t7
oiGxVDcl0i9z0LFUX1v1QAmSFZE8cnlwN53a7K12G7xtx8/+ZBro3hPNmHUQ
FLASV+RILb5kk9N6H+qlXoPbgtviUvGM6AHlPS1upYF0ysGMUFzbGjnuI0M4
Bj3+Sr/SX/XKPObIrKeonPKe8Phi39ppfTiQV63HM7de/2NN7qaUXI2WzJrs
gHhXJYGX6WOBaeKOtnkf+CmJ5+xPUBSZUL662WTXyL58LcG3auOo+1nay4r6
e4FuWy+dqljvEJHy8YAZIZFvH914+RtKtbPDp/vXXuQESHBqjW9tpojhOwrw
cKXKz+F2eB1QDNKehxibmNa89fMj8kESxHkeHgqJrF6UbhosVYNatIfCf1fH
j9P13oYuAcUGCs6o0chni3dMqvmNH5HDmFvNrmQ80Cv0+3NmbDG3sRc/WMrC
EzVJg49LzlN11zFDqT28+baKmFUnpo291icTB3GCgPIhRcxnvY+xLq2g2tm5
32RL63UZ65NJZtKk1sLvZlAi1qlbPb8ODeP7toi2W3JuAHzQBmRMhZecVWHq
ga2er1dyY6e4Ej3IPtgnJWRnR96RFvn0s7Bx18UwTNv5SLE+0axNdon4UV2M
DR347nxsfTH9Ma10Th+tluNbNesbksb28ZP0rWbF5HfbuN+/Zx9JE1i5D35M
8AdbtKol4ZBRmJexSiAMLG94Yxhww09OJ9KX8APH7QcBU6lFBAhup/7IcsKU
NgXcYeZ5u6TlH1I6C1vrwOEhJgbsxft+5lJEusKtC30kqaejJxgJhRnMkPfB
epFHHXyJvwKtwd5CBcaeX2A5xt/R1tc6r9HW96FN0dSDGy5zGqRAOCCi1qzV
LM/gPesdi9TOnk2DLANlVf9P5vK8P82511aSMCTy9LMEkizOjcT8at5vETJZ
pMyxCxXqg2uaJIq5y4oDuvhKxZHwXJFCE85Z7pEsAphnHmQRwQQKLE5JE8zb
6M8lMustQK32MIPmV6l8324lBCTMTjpcb089lpOrxqzL7zlZmILxwFq172eu
R2aUhUkpd5BHvmlGgZR8BbgLY/PRW2aWkbAqI2/Iq2eNc1XYtTirCV9zH+5g
gyKc1oCc92a/bF0rVptbmKEUz/ACr2mxC2YQqJWGfyIWq+AwZ9+6bDQ9C3uq
broKUEqBndGDiDzHYJrY2VxE64g+DvYeBn/fRB1hYHXwPfwvR+QtuKsXyujU
Ztea9UmsidxK8W5h6E3qACUKmaaz5qHfJqYZfumoAoLru8Vly3U/N5bHbZjA
ugVkKgHcWuXMGYvsBgPCZl09PiNlBBbLjl6fhKgWp2rPJLBLm5RVylrkxhHD
AlpmFTalIlYrCC36mKugmwSUy2aiX63jOgQ1m+oEuVtYYdr3UBMxbFRzXMYB
3zfYYZwEjjQE0VCwMjL9wVBklI8fn9nzdjC/rZxHvk6xjXaVxakY3u3Z1YUz
bIEzHLGO4emtzfWILqRdiMRZ7W5S/oV018LJf9phdpTax43sMkZXj+zv0O68
ou11XYbYtYlTaKuotMZQBaWE7zISF8i3FS5H+zPCb840qDP2flt8dDDg3yao
16xaKfu/SYeNgNlTWTFzIaO7AkDRnL1uQlI92xhGhcjYc6bgX+hgQlAYpLYs
4FLM5ovbDRBfK2nt6aYCd2JAV0HVqbwjLJtMD9HXljlUlxLX5fB6vRQydsBD
j7wCPT2flhfEbgVppm1f288LAUV3kRj9VMN2JaDGq1T1SkckcwZxRONwp1X1
f9VSqssz5mJqQCzVfOoEGE8lov4/CZmXy+vwRVulUW1Z9u2J5CSVK10eCFgp
3/ALeNvuD+XK75EwNJRv/2fh1i7KZgYrt0M/6UfAhiFnZCHbG3BRf6+SLuE4
U8Z3LCyYwghBKPw9U5fUj8waRMBVxIMU1ZjqSM+Pp3xSA4mN+sEbN6lW1bbv
5TXGkMWJAVGTUGB2F/EdBnzcsGdYmMK3UM3AW2eZqZRcIieMNTNRwFQDZh/1
Qrqko6IMeufVPCvK4w81NCbZGv3h+CGY2bd9Wvl7OJb73dhKO1AFkRC+fCUQ
9pHn3uQZXs1wYyHooDWTkwJI8Tjz2fGXxcUW8zQS/6NwqHfUHaG1HrKFSXXR
bDqu4f9bQD6G8bC28R5C8cOGLala8db0kGrtao5qN+to+KrSbsbCtbzDEHtv
6XbZgoUK7KHxLZROQAOPIXrfSPNsO8ncD1VJBwzpG0GeUA6w1NysWWi8RIgH
fo+3TWDfm0J6UF46o8NNXuIUZGmcooJx1Hk/XgratdQfMpfOFXB0ILgtPBy0
UU9RwpMVo7yPoxxdvUoglHajxSmLCgVzOfktoqssnVMdH0DB0PvWKz2AHTaG
S9HusrjHfTGLAjAs2vbfs5Yww0bRtdPn1uPNZFjubkfymDGnCoje06IR2ncp
XeDFsG/utxrzCmGI7fWw0NPWI0kJ/gupwxt7ogkng1BMIATgTSyC3KuFq4Ou
JIAKYedjvNIqt1W0mMrm9e41x8prgLckOg7Ad9UmrB2Yol9r4jw6x7HAfduh
WLdYdiwMoCr5YRwKqbCGQp9YpdS4Fd/KfGuTXizlPb4PAcBRt1x5+9SQ8NJq
Ua0+eTfoXMLAuzhWujGlENd0C9of1+eqwMSHEPZy+mmYMR+15XYpA9NB1+F5
iiaO7Xz/xqj1ZsNt5l4osgiG8lndFTc/+PFBIARSxdooI3RJiX/iOyDAVb3n
QwPPEGddDhFX0dX9AKU2bPifM60/P3gLw2alv1AnJTuV/OsxW7XzBY3F9L7v
J3EM5Xtm6W4w7dSOFe4nWMYQBSAiB/1pFMlMwYq0Rw+uQ8a126r9cSIYtUwE
rUiz85IzKr5eP7omGJFfhNvEHNwKWU+MdADJKlU1X1BgR58C3xzWVsORjmx+
YxnTuDgRpzWcxqzc9NGdtv/2K30m3O+vpYclRzZGok89hm529wWtce3Yjr7k
xYcrgkIZKZaiJqMNtnlMa6dR96BcABb0wsPzApr1bMiD2D4abSgJGst05dGK
qgw5AmKCJwa3RZNFqWEOhru08A9YbOnJx6jvq/bpUnqX6oNJskGNue9ckKQI
N0vuVrJnhmC9jCEKjwzTHUATpd4fAbpqTbI9prbnfAnUkl5MfMOdC3SH5Ncw
LuAKxFCcbRud4kDHFnmHXQ9vwPwz/6PcVp4ZZ1t+yisXz8eGp3cXRGNt2qSD
98D+SAvqSPXsJiHIs/uyfcj2IyLeNLhjideBIAiPeXKjTKkvSHMAQBLjIo0+
LC/ozcrdQscqBWm69/Kd3jv//WQHa5kHk/tLNcSBS8FtZ9+XibOpR4B7O29/
00wJeVnXwAKekRGhFIMzMbTbJ+YdcIqynAY1XoYgbhPfHKjQPtCxUcSrcpC2
4LnLSpYxaUPA/YsQUs3wUdfsQVfQjHMja6Ib//A8QPA29M/tGjVASMbeJoOg
bxQUXnroDjSRHx9QzNqoCmtwt7Ts1DAXEKAiQm9vYfqkRnbl2xR8SePklTb5
FWq/0j8odoS3NzUIas8itiFLCS8Gt2KBQfSDAdukaprWUnsu3ALmh9oDpv/f
CpSspoBB9FUuxvVH9XCmzoSkaDJPoEZDDv3B0XAX8KdGcUaZZCipvwwZWOP7
BxIkN4vq85OuazqWBn2OUuGR2/m7qKRErKNX+roTSgHow4AZr7itU0qHm/0N
kYrGO4g3spnTmuJgSa7J3VrnU6B9r2l73jSIlbB+rp/TWgc+wVFgvXqkiBCR
YDQSL7rOH3KBIPeiPl/0C4J8IjD4uNfQyXLFDqbRzlGiQ4OPm7BvKvPF0U77
/mG+XJXmPGFKMhdPr9HK4g/5zcDukwvLhcoJXXqm8PyG2gVPNvMRRZF4aU0K
pvGH4kL94w/rMEHbk1oAUKXOB/nLuHt7KjMJm4raiKNCJOVXCcru6FZFOvBd
WLCDksuxN10MyXXh9uJAyT3C7t05H64b+WpoOdbeKbaA44DfuVj6wrNYFWBM
WSvo2AT2ofYfD+TQ1x7GoG5feIOfxuu8oxP9WwE0i2AY0ShveZD+utpc+7E7
sh3VCiZ5pmWCXc6GOY7AIbjOZqENThcyqFk5TRludabDkrnT5JI0RIaYrsa6
0yQJUphFu2xkrwdlXJe9v4BQ9U/a77o74U548ju+hk7Tw2TdTos1JiPMVg4Q
uai8ZljkNxMkGY21PalaAZCpAP8xurf/lXF64+wvOhK1K78GW4/HX7JwTRP9
/3BCu6qctqxG7M7ylRnZTMQ6X6b/VHnAKx/7Yz8HNLyV8aEmEJRh3ZzO66UR
dglrcvZthvbivsACCDUfnHZwiTTZ1aE+hVvjd3GoJVnTDujik6zmggz5W0ta
UYU+OmWEiy+lnTs8NY7cBd4/vXrPSaddWg6ZbFd2yDDP7fTwlTZ8nlitqyx7
bpzsUCOtTDbOZ6FcQpXXkiQ3tOLGDyrSz21QC96edEifD3cShg2NskBC9rJf
PgUnkEkb4GqY08v6DVGr2n8KfjnTWl0D+7d4QBo35OQXCEvTpLf5+ZaAArB5
Gw90CDO1tj19hRkPJJO9qCtQWXvBAbROBGlx1H12nXvnfQwDpJCucvas4jen
KXLYTVeVFdamh6BxKXs9sx5ho+jaTpNiz7HWBJ1bnpT5JYK0bPNdfDKHWLGF
Kdt3W4qSP2Btmdy35HZvwA51qoEenjJu946rHjezvXfI1oTsGa1acdx5zhbf
e0puOBw25KvYCMsBeJO0Q3LOzc5ippilhvHu9gDbUNrFNW9lET2jBWt1tZ8W
vrJ67dqmWejgx72uN3AC90gDrCqLT7J89VRPFctJsvSJmwa3G1ZeLU3Pi+Cp
1YonVoKO83mOMrvqE/SsiCtZKgtjkt1Rua5eyV9giEaUkaCaQRWHJEO/+4Vu
ryLtit1pHwtyfn+0tnc+XTYsyN+VvkWDZjNxSvZFnb2JfgYHPj92cfSHVaSc
jHyrK/7+auzrlr0KUg221XuJhAHxbnv+yPIPlthvMXKYckf0NF7/I2Qrlgzw
7IIweh3YhePLo3PzM+vOlIuOeRuQ9P8wQ2/sJEwxDbvQStah5pM6hLEkzHET
Yyy2apxKhg+jBQIzCeD5pQdGhiq6k6U51r3HSS0HtUxgdQM8vcQ4ikdwDtsT
xiucTTI/E97l5eEuOatkLPHq2EIej8L8t3UG2+QTi5WepJ0JUAx0tbSIogkx
PPsuVnq627pM2U9yeS16wQ12oNYHCTYdb+eANUn7Pm3yv2bbUVdgPVHo1F+7
tVvAn2+Gb4Smo+MUOQlPHnhJZ8NvoCK+sonRYft2yDZ4a5l4D0gfhz4wymyF
ELaiuKH9THtG9v5CIy4xe8W8cM3184MLhOg1KJ7t0PxgcPzI9P5EUCTnmC1b
QgtoYO7Ulvk1LJrhsPUTnRsJS6KwozbTW7GE6s0v75Z6IyBs18rjgwTt9lxq
3MfnbRfnWAnRndX4hebxFx3gImS5G184b+IVjjT+qrzD7I3gd6g6Hd98inu4
L9nCONPI2OkoSkFhsPTJHGa5BbDMa5zSF9mOUrcgFmil9HdyJWHY7LUaaQb8
MgyRs+R57qDCXruoKL5Fedb9yW1vFZ66meNI2/HyhvMRTb/saQQ77cEuiFMP
OTgLjfPJMn8FKcxQsqu/l7wF1HmBaaG0gJKtbhOEDznXcLKOESjJTClPgCbb
suTjlc64U7/tIdbT28+MzMyl611uvqHIuOjQbmFm1Zm7AngSE//mIf1RrGVA
NIT1HyUrpnY8260W1n+DuXPPk3r9aAq1CtLx6IFunP9MeNxFHw05eQnXQIf6
MCqkoQwXXSUPdwzVtAhks+jt9uIkG06rqCUEObNmm14xI/WvmR8/7CqLsFPt
xe7rRLjqG0fCsO0BoEZjRS4KUXfilzuXCoSrVTT7bmTJeBtQAeCkdCl1pRcS
wu+hotP0ImuWSUn2i6y0L0i07p+QysIz69Oz4KBRLgzJc+VyXo1tzn0IYSc/
UWMVxpkv0iHc6iFTe1Mpuz3FKKZf6soXfyaeHum/N7M/yeP+cnI387mnYYeb
n8FtQMuaLSu0pIu4TjTt6VQW+KrRXMshIY+peBqYr2vWJJD/N65PXD/wbk5u
iLTjEyp1DsiYWWs8bGHr1wO2BhcDl2+dc1n/aHll6cAy3s7hKFxCbUv5Hr7a
1yHr1HOyEDDCCa4ZJFGJo4cHr9FF5KQoHZ62hzdrvvB4CafppZW2kHx7cdpJ
KFpp2C5eoJcu3gYhI+Q8gHUD/zO0UTjtRAdBPUvAHJYt1I+GEW9sVqxZZcZM
oHrBfhV8qJPyU7gMtGxZIMccW4aTxMysPDKhRP3fzKPAgMseX8ixm7qbIwHA
zfGPmOS1NgYiXuEi4z2zQRE16DjIi0vi2RVrppBdTWYFjjTLJUW3knIsYLMC
jWToZ/aCGUg1xJ4TMmreOl9a0zkKBWk6WZgyKEqIk6auCGTYVkxIDSkLGdZq
qDqv4M6SQAJA2rCHmMOZIDeGq+tggMBfCHtAJvqWyEJoswreXR8FOmgC4wRb
XE4MBO1vivhA296rUCKwEkZdvnO/z1BYwu6XUWw/rEiijFbL5lstTn9n5+mQ
EAphlOiUK8d0tLZPdZ6F+/UYDiKBjDVDhHqgDhv1HZDWfvpfA87MdRbyFHCj
Sdkz1oAu7mmqHU3WZMc4P3qz1ltahgAnhJNxAVeLUORN3rt6qTv2khJe1q6M
03K0/usN7jtAKWOS69an6+mZ0HbL8vw5BghzWC0UwLcht2gBtc+hv5mY47nU
7v33eUSpe7dMH6O/lGGVGeyHZUThRdINOfbE4h7xH8AgYt6ru31eiWmOy5pM
mL5Rg5MpAwDeasUALCTe4xC1dvDEsD/JbtQsKGmydrQKwW8EowcpWkcRg+W5
gCNT4x4igmgjMkuBKGYL8COYfQe64R7LgqULROezvLCNXPB42u7fTd/5DK3u
LuROipWZzOKJsUrI63mD5GgCwx+saUgNJWikBPkXu/m+llHLR1RlC6/l7csR
Cv0Bh+hEnv5qB2BYQQyUuK8QM+lgelVIv1ZmbrPSGr1VmwIZs8ZZmPFbN3yO
lG/Mr7f6MPMTQYFAkrsyinxg17E2NUuWaF2sqt6VAJZyx0cOwWF4YkhJO3/8
J7OjYm2WjdQiq5SlBShqCk0oPR9B9I6lPGl3VXbv1tPdwumm3F2Y9U5grCqZ
vQ8TWWY+vgJSyZN4CcEhthHaNmWFlaLQyTPvUarX1TRXrGmJoPcYZaeyxM5r
zcaISa180cDqr+KP5pdgt4NIsH7XV18ETF55gDYBnPF2n6G53USznucdkUrh
wnGobs9rgZgzhAJnpvd69ZqyVPlgbiM05ETPW4ssCCt08wLQMIFqy7HnxT6j
XPM5bt6Y41YnAOPdBLf6ClgaPcnHW1Wcmuck2iABE5HVzkFf2+81+WveFkhG
vq+Qf2k+uZG0WmgrCxndgsnQ+rlnMmh3j7jcwfMAcFHQwFp3M2O5/QyXlGCT
di/jFuo4rhXb4rr64xwaqZ8CQFTMPj/330MYK2kfoV5zMf9/igH7QummbzSe
I8zdLmYW362SJyUujmSacaL98dqNjgWUNrl8lCLWo6iQcVm/93loFvdgYXyP
cwOhLQPXETNLF9j9NAyZ2oIHvTGasUqvhyTq2Jm31qsLNlLsjrSW0GC9zB6h
SYKSrY4Xre7V8CLuLLL8yyD+ouQNdVxJVS20eJGGwaU3wrBwogQW8DnwFpz1
KBugpka7qxhKm0l6J44SPxn6Rig2Vu36efYelw24OpesFDVbKhY5oWJfJFz+
zMkuO5X5Kf7kvnv39TJzoHPOBq7qq/w/Ssq1CpI1JBO8qvnOlaKhge6RPBUH
hfy8rSRV1wxk6KDh38Lm620MwSxNwr0u5QiM/Tm37K70EMeEAV335kYzVoTl
GiRjE6wGFCDA6nRc6ggezXqd08yUu2Ps/p1muzS23X4YQORqeNAiD53MWnPm
6aaLeUNI5IASfWEcEJ+6EnKwZYE4YcpLBKFNXBy/MZFxI9n3TnM1qG2L4JKw
8O4QJVzThi7IvnSrC8hGUmIaGuvnIyN2UdNVDc7eqqCHQ69E/l8Sa57khFMN
6z1QYUwMl0AYRV5gVYV/AlJlylSGf1NpXEakWCLRpqhg96zSgpXgHvsgwJ31
aadR5wpyBtHY1jlc1LBf4YmijnRhwrRTWVS4YwCpgGewhoQBDSBGAGE3GXYi
NFG1R2uPUbjPpBSwOXcGnuDHbYEARaNr18EJkOSy90zk7ebGh2ufrs6jobkv
n0Ig1z64SHjKrp9d4jw8b1i6oMwoXA2HTRZfHX0i9L4l1/u+rQB5TE+Iph+L
pkpFpzMW5U2OlCfqKXFTW6i/zL3mbJpMaC8X1CO64mgsVc8S9zBDznjF/Ub0
0x65uhswnYdUjmcr0cg8xgXkEEUKgbRbGYnLGOHAk/K8EXxDghruJKnvINBv
XCK6VcWF/svZxpT+jWkSboZdtxcOqIjaxVfziL5PHBCZZCEylKWQjtesP+0Q
FQlzFu3uNxLdzATBOCl3ZnxZU5fJ3nkRBihwxvUc/rseBCP+41WlGghWH+Kx
4cPaKHbRLQvmfmk2gvj1Wh92ew5piLxJvEnhIqUCH4yPRlhNvlRZDIwSa61y
aJWfKpfD1EAi9wZFkdY4fl553kDB55RRs2pyYNq9+bn8WtZ8/WVAjbvPl8EW
uoZZHRR7K2/tYGXqlQP8lG2UPG3QSavF/xKIq4fTczTK3UZMBli+ODK9uY2y
CboJZeCHa9U0Jd3w40+dED3Eb4cpIBydJGVof2ENLzuAHnh9FPuRjq3MqLye
+ta+g1n7GErvbsv6AzLStHdjM7QMrntnh4PUlsgdUzlWSLR1GITtgdjsCCZd
hH2bNj0l1D0MCiJrP51vwaxTYFTwjdyWcPTLfOMI4GDW+bZOgsMsS7ExDAq6
bv0xN5NBJhKRiVAVf8WmUa8f8IBD87teWyzon54JJG/rOQVlwl6nabWOkZfA
nxGcLocTLHksEd/OnEIlbXDM+iSQDfxqY5sCDYlFYr0YjsWKbM5MYgDwUA3b
h6SNW1wkw8+IzeZB39vqwTOjRC/ReefjJpoeG0DW935+BiNge2gEB24b9A2v
1QmFuehDiKO1iwOpIKJfpRlIERLoFJEKCEuw25Pb10/Nz09VDtDOs9iQyZMJ
R5zi1VVrSNOiJcYvVJxa5ElY0Sb5E0b2Bgge+cLVFjzMhXxEvLl9lvNEIoTu
218HJQbaEoAlkg23T9ANPuERFepQrLibkTGJ7BXNLNGu4038PsWh3zvi3Z0I
Yc1RB/8xKLLrEPri61V4HI5LjoZIYdrsIAPQWkS50Uwx9FjNPe748Kf0NCpf
U3SnGRD9S0fvOuYu8qzPVXhhBYDgn8FO0t54ySXqskezub2TPRkQ4jaWYnsy
Jmx9U1RJEbIjuxaM4xCSuZxHLLbYJgqwXTzHlgUhXYo/JWeME4zTvoyqzS5t
gagyaIQj1XgAqbZtWI8ly7k+Plqq08N0/MDw+39W7fjf1Nvo8QKVHhQP/W5F
zkmMccoLc8k5JMmA0mafb5dttVLoMDMeWCK5Jrav25mR3Bl4ozt2pnH6I3eQ
b4ayDLqbzvf7vKcFhU1ZCbagqtWRqtMTdI7kK64XfpCrtZ3edspF0q9MuJtK
AqKSZgODoadYYQQMb2NI8OZwV1OuWAHT/1DFhy31odXif+xXwe502Ur+hNxk
q07mZhNgMEMy2XtJuBmcQNkSkxMPyvMp7V7RO4yHs9DqRtpAh+VkaCcdFlWx
YzBH5rjiJ9YF7Ccjj2A6pcGk0Okdlh4jXOUPipWEJ3NQn+u+rH7l3XVNS+rA
6lEKImMq8zXkuJrtMNv9ndKdXwVD+KEk/VV4+xW180kzLUQwe18sjFP4zOcb
XgLf9FEv7C3A8mwMc4KcspMhOW2CkgGpRN60RPfrCAE9wTXk2Le+ChR52/Be
Zp5+w4F8qICftkphSKEsfdV566MlBMnVkHBdL0NPwVFqA8p/+Ik2gmvcy35m
WisE4+D8kSrlsSSFy/6EqWalxTaYJDJDnUksaRZitEowVV7vNYHoL+qPkPZ2
g0FZv/fHijUZvZlJQ+Sf1/PYcB8E/Ry3CN5m04jIma2xM5i1FIqD0aL8SDRV
+Y89eRoaEbApQ5lqPvm74cVVAmdpmStqhIG0J7n9hZnpexYSMLy0Kn8iiDO2
545IqkybcdkS8w0GAvnuNp0QtrUK7mVhwDEMOeqWtw10CEj3qt/ANxnKjNoA
TzQLWWqvPLdGZGJ3VVw8RS3ADX9wkHM+e9QJMsC1h0FcrjOFbMrWJxbgc+st
m5HAcv0hXCIFi+N336Wuzhv6/dzTffoAVd6htgbbFaw7mhWaufiHjXppz4VF
MbMxJDHb8vCQcvuMggAyefV45ORFuAwRywUGlZMAF7RDLDIKLBiXYXYe3to7
4rSqU11lwebTtJNIFT07RgCm1gVAmYdQ5TL+vFxbze9LixJfL+YVq+UtoXZd
q+C5VZXN/6sf/CfUn1DycoY+Pq4yrfXtVBYGy+r5Bx0On5+GZKfEGWnWdTHe
aFjYtGdQQ4KolHE/pEd7mY92WgTNc37wbtvJhhQiL3hSnIByLDVa9ShHNYvr
WIROjs7Sn2SLFKnuL+o2cB0s8DHbLnlgUhFyHtuFRTtq3RcniN0wrBS36DSU
1H3+UHdUkpAa/406PRUbYXjkdPx1UA1RNW1JghNg98Cfjw53RvyDIEEHETW6
xJm79XPDAA2x5TxrsSYtVdOMe36YiQe+gum468g7Q+U3KgVG0qmJiHlnaxfL
j6a1WuQEsVf7oJySDOTocOt1RpEcPx3X3pvOoy/16bMZhohBfPzIx/X6o8b4
0f7WopJ4/Lvahp/y/KSV+qNlSLfSfoGUQy+MEzZzxY58Nsr0jsDpqPOguEZy
ZL5cFb/dbJ8aL/2bzXwoBOgHyCR1ytoQC4SBJ0f65O5ljPJIXrCQLIwSvLL7
rYXIxvaOR5E+c+dJ/vSY0j5/WYKXZm4OW+/Nhz9n3f3gHw5DTzQuQIqjAEee
1cBI4N8SWXru918ZfyLvbOztCCxXADFSYIs8RJNpoZAMT6ikA3uI6QpkWVai
wtf1aBA2AEWWPV5xWFlqgnGJaqMhaLxnsCvsUoTo4sUyyWBUj1bxou3wv3bM
MRyk48YGvL6j1DPk+EQQngP8Bz6wgfwSS6+WQTjsl2xKqs8BNpAcMQDauC3p
K9B6TcmAW7iDZgPBXfywECkFCvP5QhS5ItEXBKD5t24PwTRHItAmM2ScoyN6
teqLppBMyQFaFIeD7lwPPgoZLjN3W+4rtlqIJPEsZPjgZxqbIGwolUNSuuYj
TLkD8NNxG+5VzOua/F6Q4TetLPnLOgJ2F+Su20WJpwNGbj0GPG4Jrw1vknhO
tZ6GCcgwzrQHPO6vCReYO2Wxtisg5fsBr9C0xcGQsjjzcV8+8ZosKgTg/bD4
ptzrHC/NeapAB7W7R4I9W8zoHpifBZAtn/o34Ry8+y4J7yDTEd2p/QvZuxEO
tMgZ4T1cg9/U7wE3mcNO+7Qn+R7xjp8ZMWfHu23rOyfS0tcKveLAT6YILsD/
c/RuVyCM1T03yYR5gX4c1dF/in/7qU1bWraVI+SeDvAXNjt8N4fkUBbZIuKC
vj3xPhd0ekXclvdN5eUmCnrtKY1GlVaeQdnbcDlxL9nYmoY/v0IdnCA6dcU/
sAu3OwUrW+eNTKOUaQ93yuiDdQDlL5o/pfs7p01RYHqJrDO+xrK4L4ARQIBZ
2sGHqXQFdheVGxpMo+EbE9L5gLotMBgtabfQDwlxj5q7YCuXe+s9kA/I0pQN
u80hkLbJ/lB5kkRHKPFCuxmTs/ErRyJ3j/EAVnEKuGLG1KvQm5PKwRsVKHKV
qERAlQUrJPLg7t/yMhhP8OS+chwxkbLx7V+inu37EOt4PhqnaaKMNgullmnp
V8oB/0O6y/FSnF05+j6qdr9XKcaUSMOz+HxwDfLsyf6xq+zRW8yiPk+JUc83
FPsx48bwe6gIGC2YUKoSVPPbzhODSxTxXMevyMSafpPD/7HDqJB7OAfMzyA9
d+0R9kos12nCvZcESrdjsJQX+xFGzlOa1gsKW7ZYy3OVw9aRdeI2Q8qg9W+G
r3B1BuHtHLXQZqnFAp7wMYicsgyS8VfP5QnW5o/eEiFy4Yb4CNATvLgOrzki
QmDcK1EZ0UzHMbm1jcf4y5ZpVmG4ewy3xtRzfk7wOZATf16Z9C9mIZTAaqtz
ZhpMqlEtxqYsAErPkrJiTeaRjnHG3rOEIgHNChnscZTYYSHr62KxuLzdMRhM
NWMkMAQx8HCWWwq7l0+X7+gW75v47Rnayp8dw9TUDwj/4d+1NPFBn2V8QFp4
Zkf5ND6O7BXtgf4BdPALZgbiWeMzZaP577WGT+jBD+SWVHrxrRFA12jifpmv
a6Aqm3O4zO35o9qrQHuobitQhDB6fibjgRUohngD2DQN5zXIOQe+B1nU4Hpn
9k6DnP6IksKQ3PHqnzLWJMIkZUvwDCJ5Jwj28kkVvD6yRcaMgzP6HoIL+35y
b1OhVWA+YaB8Z9YqKIOEaUVBanPXFo1C1trw4JVxYwDPc3I1iGeCGxLySHCf
Zfw0HlNuygWnuym4HOq4mrmUZoE/0NqT8rJuyDZb9Z/5A14Uzy8a5HARACAd
G2GRvQ0/cFXNSIENYVgY2SKGZABtlZpMZc3Mom+LPj33UyYRWFiWYu9zbzx8
1rO3p4R4CbRbC3l/ki844oVgfOnLuN2NopMUlYfiOBfW+68cpstUN6pqhA8f
CfX2OGY0u/sgBkS7ebmCUkd5ZYzz3Z1lef9nEme/9vUpdswcdQZr7fg6+6SL
8MdRj60nrUvBE8imhIpeizhppFxzxWOVZiSS4KpFX6nC7XZHZDRr1G4x0Xj5
4lPcCVj4HZpz/awon3jTYhPkOES3WVyCdkLPSKYV6mewMLugjkqAiZnw8Hx8
aVnzG4Kpo6f2BfnCdJxqhgpnD9dVlX531rjP78XreXQNwg5p0RqA5eCctsB8
ldNnBGgLUcl7OjL4rV4CmpsMRVuAIa2DbhDeyC+8CHCuN8EWXBfByveuuAu8
ujx/V7HsvUS5+KzMpXb6/OJuiEJPRx6RXJguPcYV35LmVgWVacTJ5BXrS8c3
rkiYeF6lMvt7Da2/hC5MKDTmGCSJurEuTdlFSftxjqOAGJxPJS4zjoPH0qer
haUJBt9wslwa+znYTMs5GqhlHNllR039XVdBCWtuw5xgiXQBqpSjxrHDFCW6
maqDeb+efSuI/g2Pf9jnFtvqRZa7UDReyoeqKSUD98/95TzRccNHEyp+/2bf
5dH7IsxzxkahMZy3FqwwnV886dd49N+bUrzFH6QhJ8PGTy6w68BEiA5iR6/1
ihlGXvRnmbIzCWpD1z/Omvjnz2H3czDNqrT9WPkCyqpIzTyhKY8p2rQ6fncH
PdF5x0ADzPGmbbr1xW2EYdT/lrTO+OUk9z0QR4iIYeIRalssQ20WEIe700G0
hsHe37OckBe3QflEn5rx04CFXGjd0hNQZM6yzRlL3q4O/dYDOtauDZfRz9D/
o5C2vlq5/xffVTnnz1oMtN7IIBoC1QZAhOJH2T4yWkMQyzE6OUDKCb2rcLb1
QeGQrS3Qo9Gb8sg5TNrwOPsVdwaThCYzwAfXNoV4aw0zGWiRHqHErf+cEpps
3JLwrgLnI3ySdZl92z6J0toUL/zhDQskauU9wiOi8I0WmencBizxk6SURLh5
3r+KYF3HR6u9i4ZeKUbJyixoEZiooNhc5nQmHomVwq66YK0rirCTL0miDcIo
DKqMPeUPOs+0w3mJMIfVAIZuz8iIZ76DWeQhN5lCAMtWukY1g7qN5U0iGQ6i
rwRBkRDLVtG1el/3zQKDy0xlH9aIjB2I9Sw7cpkRFIBp3OxYZ3RtcyADPMk0
fQp+LV8t+VyEmDzPiReQ6KqW5sSYoD7LL//vJoaS0FcmyhtLRUd51OpcP/Ec
OUUCmclwNq7el7T0KV3zaDLzSF+7Ehd39H6epf6Xf3EwoVsSnI7001VYyU1J
UpzD0pDIMNu6T2rVVQ9wF72Lzp0ybMNA8fpYegH3DLRJqtJI0et/CS2zseqs
ZmLWdUrNcT0c5WJBbtly3JkgZlEoONOCqMV8uyq+gIPFGi3vUbMSXOgyTxE9
xnOwDb34MhuYlowJrDuBnEJ/ibEaeIgGfjtp9CHs5eIXwmw07vhsNS7dIE+u
Lo6Q4zQtTIuwY8I0bhJ9487tqCv2M9KlDG+ObuAhLvgr6izUP6tN0XRgM0I+
ZnFsJTStGdEJeSj0Y/aHGK/HMx3LtdqGw51/lLSJi7DhZXdUrA5TkkPmUMdF
ay9t/+41ru96toM/12S5rWyKX+U5oRCubQJvZLZUY5vJ5Y1eL8LIdas4eFTi
+q0GJEjoRirf6mknZ8D+L10kYQEXN6sVC30pnhOvox2A21Igs/xw9ZHZKgiR
BhiaG+7U8wVx+NEnfXiX5UgutG2/NmBMHQqbtoMleinNXVKx8iCKROIU7AXj
DfCphCmwmvexeuwffiSLXf9Vz7PDQSnlUYoOMp1sDKqkg4dLfBqfSBIo9Bhf
XaH7XGltpddW+d2oiTdtOqvbyM1cfPz3aaqC+qzvr+yyqaLkOKjNaQMMOkv0
lbcStFBN2p2oEonAGw1ikFbiNeVF9pN/FLrGyFQkmsyzdHby11G+QleSpzYU
p/VpLPmtzXyRYdEQkB0bRRE5o26SNbxcDDzvRpbPlTZowKn6QoN2+PbuV+0Y
PNFeO7lpwR1k2IcAytv2K+Nq5nSmiGYKFCfOucBEbgtBa2HrPWVtgo5aFmvH
YJBmMMzx2C+LreFE1mz57jS2ifS9ACBWYwJbsbZnVc+ApUvadUDfKBAWr+bY
C1rkvMLWjhT1a56Hale14KcXa6VqLySl54fWKww+JV03sFWwmfDfmdFMhjyR
kxYs9C6GzBv6T2X1Fc3vYiHN5OIa4PqnMhAH4CzpXB+JCKz0V1rOs6I/qzMa
O7TkqADCD5vV+OTVxgEpP3Yn6KCG0VI7UPXNQGIw1KQrQ9nB6fMtUSoefenD
2Wek4clyyBZ93BdH1KG2A2Pl9q3UgA/dO+h4kcFFP3Rl7anzuRuVhwnHGJdg
Hi2ApmaBY/hGPCaAoHViKJK5x5TYa1UyIj4wnYId4lRBCaHXJYjFZPVSSoti
Dq8njraqRvOXYldRHAV7gflVHwQGz4Qgt4vbj0fTWa8qRoBHml2Q3kjLad+2
ueUpFCCq0SRGzyUFaFkEJUTeZzj1KGurMh3iizE3Ziil4Sm0oxOFof3vgRg8
8q00ZqrANgL5MNfTBlhmMXhsIWC2R4BJYk9vtnUAuh1O7nYWODyIxWr8Tdsf
xenpvYrf1M/et8HAoi61j6APmaMcV1ZM2R4nR7jOkA7rz6Yp8FWyc6MvBwYJ
dWsccjkCag7KQFVYocDE6kp5NANLLDUqb2lwWR+TvJwaETmaSVD8G+/rhThx
E4ysW7zdzXaY55xNvzyEslDqnl97Z1Z97R46Y58LJhdxkxCNiEtk3hiVld5z
hYuM0FwtKPez+ajqYvtjFmdHVINi+8aYpy+82S35Rx+J4WQVCcMg9e/5spfB
CS2sd2MLRckv9Pkcx8lzO47SLs7P+/cQTSOmGEQukV1FJDdbPggKUW09kB+i
qztcxrM505VtT7QbcND4wGK40bOnyIRkyJ0rT0EuL8FWJmat2JLIMY2IgYlz
yoeJ+5mdDLun9DsAVOBQ/wNhqeY8VF7Qszdsr9s/9Y7UBza5do86rpzQ1Fv2
m92G6Vr99vxiEfXIT95+6SfS1cN4987RhJt1FdBwO/7qp/uu3x/nYDFLeZSi
o+Oarfv35D8dw6lVtgptiBaP88z5+GxrWLE98AmByqDF547JkgRQ7IS59/N1
7uqUZAVJE6YTxvMWCm/QPDpZMbVj9v/U0uGfp7X2TWGPp/jGKiw3/Tix9Mpv
QiA6vMCfpg+ZM0TYm4eP+H1GChSfYLz0EakD0p0EGWTLs3RFAoHm8HjAqVhJ
hi1vDokcIRr6rr7Mpw76wx0StalKMx3qxSMTyE0UXiKwr9HcSBtplJZ3Bx++
lN7uKJZwMQsmnQ1lVTNQ7tM1yyfuP/Ki+J1jZ/UU5RO9pkeDBdXOsDOgaYoR
2GPFBcVAoCVFuRQzSo3kxFvUS+dtdFM8xt1/eVwuC7/R6Wh0Sv0+WwLy9Qy+
TXkt6NYk1IVvqqpAcJ7q/HbSmwTXWwqU6lkETLvBgvl6waa/ye3CfmjObdmB
gwbdChBy/DzhAb6H7vA06twSiGsETSW4wJzciLDhFaTRG+XOUNH0tzYKI/6G
GA+29gY0e2/MmBwBvk/ApLKnpZlBJtof8zJyMCCPPWeSZblvfmtvZITSmdY/
w3vv/lHf1rp90IWviYMr4xv5oUu24mrOqnqjVeNziR/02v707gNNyT6L3DLm
NJNVx23O0F3jqHfDteyUDd5MO1TRA7N5z3EfWu2j4Oy9ZaKbZ3Etkdm1IcK/
J2SCNd0b3VlWUQEKtd06cfozCPZDGgnJn1Pb0+y50TTowHdpMUdWaOdPTyPV
aTlO/B/49Smjj5ZiPm+Ia2ZrPhrtgfDeKvnagcQ+xoiHc5yup94eoYh0uUP/
dnKTVmqkE3qvPg4nnMW/BLNHDVSVbo5A9Qhqw2Lv9pWH8tD33nbiN7cdKYP6
y+RFK+qwVK6AAfRQx0C52C3Z7aqpz9J6WcmJ5vT8QWLNGf6p20aeYwcONm3N
qHin1v42Gxt1xpPCsfszBDR5mSTZ6DR2hkXJD7iFmj1ZS89bDCeb2ee/5/MZ
2oajZMYLnCrqI4WQQ4OQzevv15+xJ9cw0QM9IvcC0JXeYFJIafOyWHfAYGw6
gNn+lbQQvmDfX3NRvvJa9P5nKAplGRsaeDu/kQUaUxQAzTenEZKudMcE/jdx
6YoCGczNDx1wzclKWekdKBfVBTIfidEvRLWjlQ+Nune7usoKwscAoQoJGV1f
Rh9eMjMj9W7jDYOD1eBr6OU3Tb2PLIob7f0zndwt6y8E94ZhsBOVOikSRfoJ
I6mXU8g7rHcg+uwjrOwDHJ3p7ILuEzjSbTk1GAXFxBYavr8Sosn1JpUxvO9C
FACPH9FBxE+v/L3Qv5kSrM/SoiHRrbbbKlf2ElUwE6WgtIiLP9XEqnadbTgv
cd9fGTah1umgPOTAdgKu/9eEdrlJDHtF0F0A141GpyucMQK4M/G+J78koHcy
bYD2+cMn6oECrOxPXyDRAghvsaTDUB8ZiSfUYTMZB2Qm9sRIPBv8KyBSjxWG
qOCRAFl10fImP6ljLNI34wly7Qv4NoOcvGDskg0p2IK0D+uWMmq0/rphyV0c
nLPq18+bdRPyRF3wVUDiafkXC4sFFcjvXD37fJocQqNsf/PSUZ9rfJLCFYRU
eig9YxbGFhRmWBuCJw8sPLLEAFrxcwkVDQy6qqcZyw2PTxli/IQ7QZ26umcw
qQpJEhU53eBqqKS2AYqFyM+anc5KpznaD5Oq+/E+x4BSOWcdT/XzEWCWQ7km
iqirSpbnAuuvfI23kj88H3kpghWogDXzmdsgHmfM5nq5owgB1zcROTi4h1cw
uX0oj8KbLPjIbTFg59MTRx2/jQaPt3BfXUM8nCr4PeLvZhpJg6Fv/HvTRNm5
eatylrpWVyRD+o6t9Fm5FBX/rh06WMo/Rs9QqYZVTG7j6BxHzEKRNGGyIS1A
+aQWfb6Jf6ksfBKtQDhzWdqmzg0SIVZTUbNsWq+CXDc2A/RKyD+62P9WurnV
rLDDo3buqLjfpsObgJFBIEQa8UpHuDqi+XfK0WFIngmpYwEHMSrboPUIKOZV
MsFLWxB0yxs6RsYLQc9vEqPgVK48MKeeR1JfBqv6r/APDY0GYruy9MBdnKp3
dP6ZPX3d/qOIBfcKKJWn9CY4++U6uxx0NKJ1/8CnmAI4Gno0x7SSHXk/6DZy
ClcbLNXr7lFFcwJR6c94GXUac9fRAAkUaVJv4phfOC8Lup1Y/cfimqJVa05X
89G0VJSH/VMPsH1vV0i0kY3Iqsw36xGZ6OCvsKHUA6noIrwcRE5JnPA2WA2X
Kv8gefCB1pMcYPhw0AgIyccqtlJy6HVe+85yyoqVZPCgMPombMBWG2OMf1J4
VXQ1Gi+RnykNbJjwdE/ItkDQ6fPShQVXCP7lPYBT4g5c5y2OHZqJJEErHjVN
gp9LwTc3Z0o6EYjTpbo/c/3YMRuLfWlzhY43NwcVtqppsGLP0SLdljYjOE2i
QZlRZF4/eicNxbszfWdUvNIl0Y/98e1UVPTMQDMUracVbTMUbaZj3VwbtP/v
uGuYps4CI62JbGykNtYqdo3QfzdJ7ALFziwuLIBx8G7IRoxTPws8N8YsbODH
L/2RStgHyoB3DxTEfhUXJxW+rmrVTSDojnG88Tf1wyVGJmOtGic5nde1rY7m
ZoKZoDsrNTmENPFzGU9t/PQHcNaC5rlDQh0eOCNpSLYQpCrORq4iSTgXN5zx
i2JfMIMoB7iU8UYjdpYxdoMFw/EqJ4ZCRD62qzAV2eCrlK4LuLzvSsAh94Go
Ozp6cL7FVVh1eJpaR8J9s4kFSaJiBQCTUUzH2YeE7oWcQS0Vnxk0p74FkciP
k30aS97tEMsgRcqcfueQnaeRhBvRUt/l/+I29KdbGmLOq1M7v2IOtfG+iB9q
Q5Z4IIkQKdEwaHBAImFO3iaYWVv7EWN5vob6bflIch+09UDPXDJu9i/ZMMc/
Uo+TlwG6peE7XoGbkv/sXcObdvyEFm9ADstURNtqnaX+EE+uAvcXk4prOv4f
Rf51xTBnKtxGTYlZU2Bv3JNvqwQhV8fs4j9sjJ8w0YclTcf4BTQqUGq8Oveg
bv7jmFputwC/er54CP9GaHBr7dNqR4xNxlWLSnnlDV1890A3DJiernL/Ehl4
yOkEZ2su1Ae4uSeI7eyQYQT0VnVSUsctYOhDqkL2CQ12T/BJPn67zQsQln0g
TQTFr+FT9/83MdeAlvSSjDA6BB1CmtivK4nTqYBahh72kiQQZ8gZNUSHjjY1
KwDSZD85asmQZvJfE8ZIxZfSD6fccApgRGzg7KTHgAmMMOCANJFuZdrwK1yT
nDuk3SBms1nWUMla2abSUy+IZQ9LI6NFmBbIsCgv8uN+i3HcZYk0Zt0g+La3
s95c2QcF/zY81/zPIdXBj5WMSYmK70SedffZjKg842esNTMMB/t7budWlyST
b6qT6eCA46AfGuPONuYnhU4plre1MXGuZZJE/sss0Ht5xkja42wKyOvZZsJX
2PAra7zYZdCooOPei6yBD9ongRPP4urv/kOv5LyLwQUNzBex/Idr/xh3jein
IBFrr3gsANLw0S+eRrfemG7lIQRQu2jVoZvR8ecNn6fX3665N78QgO5afyAI
hG1FyBxu6BRgYbSc0scplADf5Q0URqTcxJ+d5zy8KPLD6DUWlfKH5WLC5MGh
X7V76i6u9UUYy2Y4QMjIZKMOqzW6en3gZOLrEC8r9XTxNEjpVIF+p0GXmCTn
9+1LteiWCu4E0WNDu4L2ZwtWqePEoFI4iFAOLngdPpFLe53OVGX66dcmODJr
tGyQu9bpkyYOl0Cj16J8P/auwCY3LcohKb3VOGIZQRh0JY+V69lABh+CVtB+
iCs866HnMspfeSX0gkaKKwVTbNCLohqeVd0h/OQjCBlWn0GgaYTCwnMjPVL9
SoLlzFXcO34RPWB4xPOTjnaieHxIOlTESDeqTVSZsX/gyb2HEFzzfED4oh/n
s5afHqcKXxtlnaRA+et30a1+W5ZzYtOBI0qyQ8SRUZ6vxkzPqofB93NFSFuO
f0VFU9YG8k5B2lSNeRQs8vkNOBrGm4dMHXX12jPDEKirjwIucCg2w8wsKinj
fD6UBsTpQpldckAofZ32n6pI75AGiG8kmd/fqZTyuTLrDYGoaz/mf5pSpEQo
kIdlPSmqkl+CL6mEEl6FpSvkBQ/UwNsvTUkclYpbCnHgcIRjbfPwR4l0zmFI
ZmuRB3SaZfXBScJGSEuNXKYVxmsTeg+lu69gsZpTMTtA+/kiIRppxsAdJWeE
52Iyi+yGVSWhQFCoNa6/7dqsYV5kjNvKsk3po+7jKd33IGagg8JYk+PwkgFj
Puvua2qSGZvD4kbBtb4ct45TLrMbjaBpkqaFwqDA/ZInAo27mHcX6SQVyuZm
Dn1oloBE3w3Tuum9ZxvMEpoeNrrAsJ8CsGhyxQFOCKsinRzFIaCLcDmH18op
4JAQ5BE69+1amIL0zG0bItXJSNC9ZjacmA3Esawask2i0MeSF8dZzJ+KnweO
IfJemNKq73Fy2sVPSSb97+GOtbu0PA/38GgVa62hx4A72jtcQ9ur6uuXBJHX
En63sGS+NWFk2hjl5M/sfkClk5pePi/JyjWa6kepq6X8EPxWef0RLhor2xg4
8yyYAOiMacPuuz8q8EZEjJWi9qte/FARUvy9YPsmqqIWSeLKLGpr8wb5iEaa
0+GURCB9LG3srPer+Q3Rw6nmfA1G/Lpb01IWYpRoCwcP+IO44n6Pad+78t+b
oE4pw8f93Fp2qOps3vGGGq1PMudOmyIE9lTSuc71R96lMwavWW326IfomrDg
ZTofKZOI5C0skcM6laumd52EqXUlI/YVo+M/xfA1csA6pNBBgKAriPi+wY00
jT9lb6g/NYDpAu92u8h0VpqCYQ2L9RNv2yNA8pANpt9i9bAfuwg+YheMDgf+
wSjslixpNDpMQLTD95+tvoGKKXSKssPmzp//ZlMBnRfsF+WPqbz+GXcbA7Co
0UcC+3lYf76lW04Ee67mGQ8Q+T9pxQW+KHVYmix6qz6s0qq4VEmXfgT2FrqE
1bIer0TAl9PxV/jF3qZ6Bqg4xHHJoBYezhlatv6VpaCxOxyBPibYRzlmapaw
AJS7FIoJKeDBBAAsZbXhgqmCe+ziyIunniyJTRRdAGsoTY+6cjNFwqbKNQxc
VCnCjq5/QxCfvN2AnSdyJ/bMikA0Jcwvuiwjt1oaEYIZJ7oeXYY8kw/P07Tf
Knoh3BwD5rKUUr4HyLfLQpBFIJkQeBshOfsOhPvKELMt8ia/MTDpapYaaJ6c
U0cFQypxjf70WMM6DqNesAJaU41zeFSI/uEHSjRNSvdBcO45+m+O0WcGAQpU
iDdLvi5by0I2NA7x6tViPBxQ8h72OOdkElfGdCAAkLQ9FBg2rRuWcSqH3vZf
DDnscyP3TYpO/h52lUbfO2FmlIoOLTZqP0PCLt+Un3UTo0aaQWmp8kydexhj
tNc0IxXGhB4P4viz1UVTR5xmlr+c6l85YBm59oTXAEIZHYeYnCLGna8VT4RF
/zhEIeVv5HQXOopE8g2+zcFTlm6VTRvSL2iNjWfgtmYupshthxnPu4EkLwPK
FUkxXkb4dKM9cJg4W3hGEVlLVxO8GhYyjNOf6yqoPFROoKNVgLq8tsov04YN
BpLRgPiaOGteXC+r07dSOlzaebOms7s80Rznsh1SnoJYx/2ab7gy6bxvXa8w
3weoUvQrbIc5K5gKTasYa1oegZvxWQ2FuXUL8OlfvmrewYeX4N7PwfSoJf66
K1CJAxNnOy7VNXV7Rxkci7RjNkQAfi1zVV4TRDfSlu1QqQsdVioytANibTlS
xBSrxJUbns9jwmVUiqk7MbKiyAwEuRhju1sAAOiMl7v7CYR/9tPT0hC3BhO8
8xiOKDpOvSw4y0fm1Q/D9wsMPO4nyAKJ3IAgAU7AiXSsiD+6rX2NEns3MRFg
uUwE5zTomhQIIAmEsgKFnrgJYBdpw1//6OL1O2pWUrDfv8RFB0Sh8FesKcfi
d5TzCeccE+Xpx4ufbEA4UZaQeEQuwhoXeXVC5KktOM3MjngBf6zQJWqOdqye
8UsTYt+xmp9VUG8ZwQuw+cXG8Ba8Uwu0TRFgVlfQJ5f1AMmt4yVKrVqq9plg
pkhO20Lvov+WkbPHxNe4YM+nl6F+GqfuSjIxe9lul0imaM5OwUMjfS54ecNa
/DG/EwRf58KT0EN1Svhl8NGb2GJqfdE6huj07+xskdB5ZkRHr67tQpsOIu0Q
tymLqp1Y6RIgBQIp/LADrmLjw+LX+5PjKTqLI6s7inQK45JBr/hXQE0SUKeO
ldCNG4Ve7XlPxOrgH5u7cQtbnvH6x1p/IOBE2rfpnYFQ2JRDjWvfNNuO4Wik
N3Dv6dOu+bo7Wp1uPvdrUAzhXcpCkO2j2yK/mvp3n7r9Hig9ZPoMstIK+aYn
YQPPW3YYoIVKcWAokTVYokpeKVkvCLYkfCdQiGY349b6fczP6jZxO3maouNl
U00+7rhjDbeM/IIsG0AfyGTu1eeaDJXvZ8TfQ3hZBHevCS+fe0fIwJ+N5UAu
zGKWu9GcU9rkRnOGgDhENw1ngyhamfUz+3PMRYwUc/OyqyAh3fmoK41GV/M4
hemB0/MWrWC7MtJfSQXVnKZ1JeLu9ek5s7Rs+SoQNv/sQVLGqN0rnEQVBDcx
aO8STukFZbEfd8+FPupfF0HMtwqphPxUulMwS4Tn+fgj1IUp47sXQiv1gT7H
ysxp2ODwO5mV4haz8xWpljZ6YkXAxcC4LS3cZkrHcYpXBWTfvlzzyySi6sCD
Q14sbJHAGtUrBL1qRetrUkhw7gmuR7+b1RgWjNHHzquV431F2Qu1JYFiBlVH
ryssMi7yL9ff/qQ7Hh6Y7c5TuVEkBU+EeJYwUOvXmA8+jJv+k/y8LwWR1yN7
i9/mvGNO7A9bnyCVlJ/4qOfvkqxZpvjSt1Nvq46ZdiKzZRjDsT5c6Wd4X+hL
HX5f94pWBEpbBUlbSGl4KVvzxb8NDICnAW2bQzaJKKIIkzCNtZc29h3UpoQM
rPGed6gP+XLFRrwnwrvDaZz4gVmLtRwOhSn9oABmxxkxfbz0645BZWUxM7Ir
+6rFfJqtyVvxgA4MYNv1syHtIKPapiPJxyF3bWQg4ZBImBIFSCGVrSA18J3+
242Ld1+5s5zGTqXG1es/x18p8Pp7Kkb4V3TvY6AJAuSiHQ2zjvTEddIhWSLh
7EYIDxSzshY7xWXBZJMFyFY3DHhxZAgFKXQQq9ncWt/m7WgJJVXOu6IQDGsI
Yfg9njX31z/AeuHIZwGLtqMGBnAxPuewXr8GdF+17E3IQM1f3goyMxUS8EyP
7CB8/dRrYfYQdC4eE1Dw/YjgVOwrHMouGLEGxjBvHvJbu2lsUgCXDf9+TszI
IYMsDhKUiT7PmChpA4skQKYz4jFRPcXxjYwrSC1aUYAu9xvEg383lTVTqJiw
lIQWoy3VhqeAFv/7zI77/GDDWLk/yV01LnqJW5tyeaAXb0JmORb5RRjJgVD4
yk0FRUVM3jdpR4SJDQM6LnYLg3iFv11xU00r2zJhRaHaaeQC574hvrAmMbc0
wHg8mWxXM1PWjuVXWSQ2BmDo5q7hzDT0+ybtSmkXYLyNdUZkoZlz78QU1Hv+
PkaoBTLBgUnV4Q4CYyeWsbJ0UpTd+McL8bJSz8VAcGATaRcesgo/A4AQyZPZ
PYPBMw5LcaW6ELgx5V03vTyjpv2iq1ANh2F9cRGo7Xw5OA1fjvlj3K9y4ZDU
GrBWqnr5Eyab8sCwng+uSSyq4sHy4vl5Uzcud7HVgxJimP+69YZigmj34cKI
MmyBdp2Nj6q1I9N/Jc7/IEqNkSAdbQIVUnuwjzYWERFJO3HUD71rvxHDGLnU
2ZqXNWf1+YUz9HtskGhSeO3RdHL1VPsX8LQxku3LNdReRvvcDPosUpZHXeRt
pR/4vveZyAJHm9dGmOxizv0Fx3Awmk57vvbwgoAKL2PrSTgotdgSnk2B+JPg
IJT38c4270q8d5U51oZ98M9a9gVRiPlB1L9WCzORJbEFW9baSKaa7oeUwmsk
pbUWUZStp7GYEhXaUKAs1d2MWwuv3v8kJfdSTuhtJ6ZxnFtVJ0D7i0ONYAIs
LYCuSktoiXTAKi/Fl3r7toMr19I0hAO+Z5i1sG+vlPyw+VI9uqABeDR+9rVh
CePidpaKl0XZfEaPx/pcrE+8Uu0lqU5XxXLCjDTRcYNMXxQRT07n7/tN/LBc
giB15tjMbtXijdH3A95zcA6rr+nHxUziB5lxP7HnPcgIxBHoPsABzOguPvHn
rPtRfm3QVtHebaxCWLTsFbix3OBvU+0dO3KvXljpQNLee016hingaLdqV6cc
jnmvJJVG9048UMIykuiLOE46+85+JE3fLDbmV4Gf8KO8SyWwktNCDP9Pl8wW
n1rxuBmrHKTflbLwRvHHUl1s7UJJ1y6wwhDdKQ1th74V4eDYVpMVH5LWfgn7
VlhmW8hsbYjzs6IfsT24sXHipOX8vgfuLe7U6/2t3A03J5I/oDVeuaRxiPmK
y4/8MDp9oO/kb+VEcVDT+1OQtnjvtQ4Z1NZE4jmmGZ3Dd9w4IfbW7v/rKIh+
X4PQlFVbF1Gd3IUnGDLchouaAqjw5ayHR2JDqq0R3ZfbzteMv3YNRvvRv+Eg
6ytf6QzlC1ehcEKqoNP8CaJXMh9jOPVZOISt/lPODjxXYzYMEo+dR/ZnpHHb
vJ+S4HQ/TyjdaJo2wYtWxBz68WSJIumc18rFG5nRSMUl8KMGiWhgkjEK0c5c
Db2ThmvpjkmekmeygUJtjOQY4fFnMDRAwW4U+LhmZz/nKCJpr6CU8iir6Cw6
ztWqpLc1FHIiP6LoDmRbtagagWqYlLiOqV/dCWdo9rKLbgJlMh4u3pyZAt76
dPzSSYGKVUNn1V3325cNNG6UIXw7PyeTOxcbnxjbtyWo9aVSwkfDPBlo09n+
Fzs9P0A0ltEx/XGwycMRCm0tM+sCmKZDSHfoFwtv2HrIvPmEXAgOBdaZ0Xnr
LHvxG7RigL/mmnKfLzTb6RZMnZN1n0mghcAZ0csrjG67+8v3Dgqv1txv6iEQ
baiykyokOp1vjyFDzxbHMlaRzi6nn6VV4J6cKW+2lsCSu10GJWDQetVlJFG3
NgY6UDQ+oyxvUu6jM0NVgjnKR5lI9L3R3iyxSE68YAvqArLs48N8uq1b+Gt1
P6sR2882DEkLbwV8W4XxBNBcAJxc0XnTdAiCKI4mPRCqUwKFAk18Dw4qIxLE
FcgF3e88cQjikWea0EzskhivrgIJgLQo0TGv/k3KXBklrd2dQOD1jUSTz+DI
JqU0T4zL58eYPel2NODgTFa+b8NyPPhY44it0DPsHqadUEX47oyk39DjmiCz
ZkjA19L6o6dFex3NBZpmSiz3OiwENjdVDMGbMhRFVvH3nb9vWaNcAVU05c+n
XaBVWZLbIwhFx49+ZWaNoGKyemsaaCRQOUfXW13aIESpgEgdNC47qQrWtUQO
Gg/ZNeciXHmM+GtTdvbXdF/ZNclOn6qboqudZzjmy/zm1+xskAloIWRZVdoV
D/lYLu+9PU7ivJRqjCElPVX2NW5u92cIxiZ9kEDEIKpT4RdKeL1nqDjFHIQg
/7v4YaSwecJgv90QYG6JTU7JJ1GyZCZtUQ9Q8rZJWSViAKZmwwEyDHPAy3kR
HWyZ6To4BLloG0LhowJFx+AeGSJp3VSYyUNYaeSU/Z8IaqlFD1/DROiXPZiF
XZgG8+BZga+YWioVZlvPrmylMg2wv3mP980XlR9zogspeTkA1tFtc+mS0nyR
5Y7WGrittBGf2cK8yM3x5bLn8yZDDCCUrKUGHdVaV9ALo92lG7fyKtTrsOb5
lD7vLVmLjV2mtRLO652Fp4nh+p+JnlYPKod2/gUyPlQ8vm/+bB+B0ulszFds
ChoRMOakNQzBky+6j14ymS7TKEPp+tzCHI1cYH7eu/yNH/vFrk0V4Ry2WklL
+dxnjxJ+rAbtwme3TMm2Hc35TvEozsFI5wMlK3YZ9NO/qOLk451A68VQ3kKv
dtLd+A9T47Jn/qz7gsUKm6vNXTS5ar/cxWggkPgBQDQQJfMHqTJt7wPquWNN
z08ZCf06itPG+jNerwF9EKS9AxV9yFFvGAeS4mDF8YOHyOpZPxx4uhvlvV03
1TH3htabMuQ2DtTMrHTAcszk4oEpUGZgIY3s/GBMQVzqwILq88U80jaMjkPy
pt3SZKQpOE6j/GvKo/Hsr7m6YDqQRpUy19xdiD5WgVdoOxTOag1xYkqA25E6
Zym+QOnoHGeBQz2Hcfa6vwR8g3O4tzw73ejmKS4N4rc6pSv3Bc359xIYzBrp
HdIPMKCakILrFlRL0VfH6mltDEG4WBJx+uxIWiHwxCa9+Bey9X/rlm7ezdgT
INSljsOGDtWcNuw1BHnxdKgZIyMSJUh5cAnsbmqRpcDD3+ichSLvWuxppxiZ
EXGo8LKHvuFpRyqhoHVyvNT5Wv7hpGeokj3gFpIdV7CWj5yE3iYaTgj4OzhT
Gp5LhcN7wxOU1x6HTUZ+EentANflxCMFLG9jiJ4+FuR26dAIEAqxyN4aGuNa
TRTgzTO4zIaOktRPxypGr7smX7kIDjO4MOypnMjknyOM/Z90g7+8j1Y94XKI
6oRK6Z/gJbc4OHi+fwtuQx5s7Gbp4dUmSSM6E7XLyH4N7TA2CnLCbhsDQWlt
2Ixz1fx0IZUGXsGVcr6bZ+CzsRQxO+uizfWSTcgRXk9DJzdddJD0eFS9TYzk
vLPL7R+Q8uktAYVOKTIUOJbOyfe/LycoQFkOcu/js4hrh5ipWUGynXb1am7a
njOUs4PcSRT47+uL1Rl16Ltu7t6ZBBgnVfNNGOKEiIHK7t+BYVbmDTD6zA9Q
Zgrn9+33ryr42Yb3iBjBXo+XdiOatFLvU56ledfURwaGPa1IQBIJDQx5mcQB
KPZraZ8JtBSG+/S9ZbcQjd4+2BBCinZ/280WDIF9vPsPbLlz0Cj5gRh6OxPV
SejCrFl+Y5p+u2/Ne4e2S5io5jxEPvMCZbJC5Ru46V501oHbFP1PVHB1FQ0N
8n50a+gsztsoDwjI8Boo5QZmRwDXHUngjy6HkevVQD4nRe2NKupdS5iAP37J
ZHFSY6gEtsJX9FxJDWPpwrtI6r4ab46CdEoUCrwiYOmw/G8T+eOLKIPihFZq
GbF2rA/zLnI/++62r1Sqvb00F1kD8F4wwZIMgnBiniEUWK4IMJ/ujz8XQOcG
nNup1aTvxMtCrr1AaxOke7YAlqwUppwWonfEId2wvXn0iurXB21usd7cOgmv
uQlT0wqSHU52HjyEDc/2MhXZtzQrt+Cv+wqlkszZYj9BZv4kgAT3ja8pIFJp
+pE4+auripNark7fAXm6+v59idvnWV1vno+5lM1iXw3NdDXxnrCPcL9ZgQYP
TMpvcwJ6xPtTpGg9Ay0LoTazRZgzUlGBmzDu+sIAXGcCilt8A6fony8Sqgel
WcntWY3Pe6V2D9UwqWBHl4Si8j9lOpAsZPYijCuQjf12ox4Y6q6i8njq6M/V
ZSjmjEn2pTCcyGKYYcERFZe4f9+EGktA6rjOWaM6hULNDYZgAxyVSAWB5Y0U
QdukVu5NDpUsNDMajtTseK2ezrPiBktQ4KfypIKcE0N7sWkDAXEjJisuTsVQ
c2iZ1bXaH0BL8va1/uO06dFyv+UjV8umzpQa7fWnBovo7HFo9EU/EovY53dY
2OZ8d4Eu/P+rF7XBExPblw6uIrD6GibeN/8NIm9ytIv2M0sOJktDv3GanXdB
dRpVDWtrLtYpcFnAjz2nXdi5ffSBsEcdsDjO49O0qFLRIjRq8eYaeJQbUe8i
Ny2gZ7hWgc2xNCpCYwKAUMmkE7++1/CzLLDOoDbMHh3yE8iD0TpEnsz0Cs2H
nQnbmbmt7qUEfZVpLvkLtNJ5kRgCV5p14bOmrxv9zoPLYAzZ4z7JAVcUFWyM
myk6Vllobt0RAWL3i0wIV+2XE1PiC/KDYU99OCFkhvMgcEt5sfDgv8fKt6Nw
9k6Z2duoQYzaijol2DFdZikGgbO0SUOukgGS4l5pXEyg2CSDJKEg59iZFJAf
qSBt1FQfUOadkfS8DVcNlYW0jMxKsWpW/a6ekVQC53BwmfnZrxmQ3iRxswKk
JqGhoFDwceReS2fsk+Kgk+f9BTmByPc8SupZcfwU2EnzeWnAvpX53OBcX3ps
o70EFUK5QEuZlPZvv38mp9FpuSRErezIbcYCYajJx4jTyQsl1F/eRj6MEogm
WCRbL7AWoR9zSutE438CHZOTAcD/icxDCTrZuc3DMY0ffqaMFO4i+Ac8k5+g
ak1U7kmcwqA58RWUaXpH/8K95MsY+HwgRaAkBGaRFJrVyd8pX7joi0S07cN2
FYpp6UArj6n9ILVZLcbQ/97LDXIWe+eZDYFE6QXTnvg0H+GTvvW5BrM+DVMm
kYr5eTojr9zwDpHpHLmpGaYb1L3Nt/zv3AVTQ7ChFt7JuF0GioxthLczMQkP
EXnFA9bNO0kACQrHnBU7KKlrzcuXknPKUAmPAvy9fTcdoEBoH5nJtARzI0QK
LOKJ4twVhzK9pbCCrfq30W3xLKC5IjMHGohKsV5uKbN5MVo5mEe2tz8oEpOf
HiR3oW9XLVabPfRnIVnE08+g5xiBm+fU/pwe4FQ5uO8Qah6iUq9vVLasa/Fb
YV3CjNiXlfGnKfLEcwsmzyLVah8/aCCbjmx3HPJsV5dX5KCF8FS78GFuMMvn
e38vSwu6RH3fmmyxNyaivtIrKsjLdvtwIj4RMzu9m/okqqnEfmKf3N3oZ/Zx
/EbGrINTKWzaumRlSLzjZFUvAueu39ZVztIE3+lL49v2jV5gaX6UQdCqWpbO
9vJiiKJ/3PtjVegfKecz8WWuEg+eVNKghQrsccTaU2z6n19hW+Vl/PUzO6Rt
xS3ArFhU5vRIPDp1jpSSz95I93LVWXI1LBr5LcqCu2ASqvAP4WYyjeS/vJKp
SaWAzbeKABoryiNcPX4KrTcwzcCaTnsTO0E5HqEJEXwdqLJL+bK+2fRonAj2
FPFSjO1XkWkRzZyB/vfDEBDxgSzH9uwZmI5TrlHtaYDeQkty+Uo6152Vboaj
3QZ5DAMCl3k5m8wyfo26SowCKc567Vu8vgm88j1KR0xMfeBIs25y0F1qqrRf
NOdD7c4qDQm8UhSN4kMhObbcT2Nr/aasGss1H2i2MlNevMCajaPVXfIDBf2e
NkWBjE7/T17kOGEFc76zqkrSHCw1h5xPinY0DbxaCaptf5tbs2eCAwaBaA2n
LpBmwCq8IOZjp8jbAj8CaTb3qQ5jkk2X0H/m8X/QAF+yUYSjz7AfnJCr7anV
SYffQ5m3MW4x8x6Y/skBpKEdYC7Aax+QgqoTGYP2X0zCaPFr1cI4Qg7nwm1g
Y9joTcTQG2aWEm99QVV3PzhkEvccQYz8id5xCTQ/xapKwtVgzYs7Em9U3edj
wiWPyJ7gOSPhs4Tn6EX7/Nm2Xe+XsA8ud5YI7FjL6n3cODK2PRs4YkiLa3cD
W8/kUAEediwh+Moys35PEieC2cZSs7PaE1iDXYypIo9hO0CCa4tcxXikePuX
IxmWva2WENTBGDJKXANbXYR9zPzMzFSNQx8b+Pqt7Su/ewmHCMFEnVMTohPP
OGd3yI/E7x7ziNMGtG0mtMLIG2BBV+6DlKnklUG67hz1dPExFgd2dIMbWQrn
rYTRbgtvVd1lv5mt8gR/s73Kx6x95RQyBHbt7vUPZIEFZnVALgMPZFODkDq+
6UeGPvgdxfJxhBEHQFc78Bw74tyiLbBnPmb4m1ykSbx/a4xkfhXZEUEPvKgm
uVQzlZSRJ/T7ufSpvvc6Z7YIOM8ThQToe7fl9nsDwr8mMU8PY5C3C4wTRcB/
c3mpdBjblYzV+urKZyl99Z3fw3H2q7Yx58ofntHNhcNasBC9Efn4FzD43Ebk
Sc3S99VYKDz5zN9EoE+1VgKFCzJeHBGyv8EdoojUQzzh/yPorHqEecxvtLLL
TxGwH5oTkn9Wkq6gaS73/e6hIFyIseDjoINcjEa11AcMHfVSE88txCczXZ8o
TQLPyVG2CEBAEL+YivgnkxdFkhoeikWH7RLMh22vyYIczoemDwmA2YX/4Jyz
3+1eDkOIdcr1U2DKpC2cOrJOPgdVPurQOYAwRdZEzkdULY1hqK67YJ7bjeHv
k7leUmgeLteN/fdFDgkjOwd6wR6y0CqSNpeHVegcJPhGBtKPxRtmYHlH0o07
gMHIyXfFPriar8ThLoyrGZ0OyNsugjY8JbI7BpP3jeghCF1dPgvcA0G2xBoD
/xbexMXRm0F1VeliLdh6mky9WR33QdNsRq1ILI1mwumy+HF6HUBjW505IWy3
TpERdG1TCZ2gyrzii0+32JBBCX+iwNg1QzijVsVKFGygQKPYMvjSwowFF4fw
jE8IolYVARqabltNDhTVC0/QkVrzbmxT60Zlc0+1lLy4X9jBbdj/4pAl0Q8q
4Dqcj9w+dHrP0d0by2MWbSD8YoCLU06YByICg8Oa7OLhUOKvKq72K5cP4nkr
7BZ3ASLSlqn+1wxUsjCImAsD8ROWuDQwm0wJRh9qN9nsP4ljM9CQ/Z+hSD0S
j/VZy1ImH4nk9hl0k6a747nYZxKefGvfN276GnwKnlJg+ARPUswRwIO9oIgs
hn3SxYnFVRyTRyVzHKGEhIIAZc7ufHRnNN5NQnOvmXBOkggT9BMltPYnzk17
YZsgrGtnk/JRQ7lFSxRTSeSt86IANY8tTvH4gy2SN3ug7b9Za2WOm+CSVWay
DPM2Mblt4JiEZk0AfpSInwFK4Pnr4sHoHh8Ae6Jh+YsBF+3UQTBdmJlKwmHz
nWVRA2nTrj6qzvcCRgmLtysQy83rtba+go2f2nAF7yMEpQ/eEpgpr+uI5jj/
Ap6935yfPLy3rL2+e2b91AhtjCSR6H+VF1Re/JKDBldOREJhA2gGS+GjGg6f
NOGJa9yI2Gprsh3P9Th/Q7vfF9ytqfiJWbuGZQ3fCsLYd+56oK5/qWCDExl0
W8Ty9YAkUIWcJ0avWLrLoQgOKEIh+1rZ1FOP9wWk9giRlVZpySV+1u3ylRwr
fAVeQMlkT8RjkgssW+Va/Tavc0tBjIax222r9ROBwsi+TKCBQscTs2o/Oozq
nXv6UtiK9Pw2K8yJu9gvNk+hFQtX8TNPPQnHPzNlLZtrc0TRGls85kAKq+h5
QDw5zVrwFdBoly8SZA4z/TNGnc+wsjdboVpQ3mnj6S56ELyb35wVSWL487KF
95oTcp4LLmP2q30jlZzQ7RAq7tsY462yWJJqVBmYAO4xf2AbE+ppUFrJuqdN
HJRJgrukLOJp0Hi4obDKqVGX9gFysstIekSqq6v4hp2iQLdTxNz9+uHqluaw
Y3WMPfar3KSCRZDKTJ0Nuhmf88GJ9zanbhuvqQZ87eLRbwofKEy36udO8N3E
We1VuJQV6k+iJ34qKu3USZ7CWG978lrNDEB1sjUetR4KIQGm9uMOI6RFsCmp
njL18fEYgCWvP3vMsB3lhqoPP1kTJ7CwI+r62jgsBTv5aKH/4NRHZ+9UfN08
CaDRWvYQFRjWpiPAMFo9jJdQiGu38a9VrreMjpRThMVTGzJFuDSQWy5XTa5j
fTVEWITRnmjCFroPNstr49Zx5whnQgw9V5skILrH/rv/TsMcrIhLChuUUa9a
/XEDTzW2+tXBh81tVIKbtrtkLQsyNkt31dYPSSyuJK5TtZFFgely6I1BeDtU
sbohz/OD2tKU7oLt48+MGTMEefwoCwbc5H4J5RSev4K8X0l3rVQtVeTso3a0
BQzDGIRDaHIe5hSYhCNhXIlKfihtNNyOfzf1Gab+DFo6nX9hNCpgN3Qj7Cqn
eh5/IrTcM2Ct46fZpRxyKh0tjoW7K3pMa2wnIViyP9T5KeXke8zOr0NDdnzx
rlyXVbbZ2f5JmbMR7C16Cklo3S5BxHgRtJF2/P7cLDQJSEsg8/Qxk3wP67VT
SmI1ZSJ+SwSH4pCIKrJbx4AADiTOKpGRWzJT+0bZkMoiS0BSPuu5t8PSt6mC
tz1QSw1WgAp1y3EEy1QZxNRvZrDcralqOi3ieAMB9t51fN3zlVIVVYSsmggO
QVgwp+FffxdHYOC8380zkyJqGPgAjCK4X7HKCQmphkg5U94QzhHMTNgdmIlx
4rjSqT//elfWt/HIpOFpvO4E9svI7h0Indhm1XRoeG8Q1x7fUiJaNw/aiQFM
G4rEgTB7IcWjGXB+jHtyjObG2xtCeTOP7vGys3TsusDsmwPU50AD9HOcDqQQ
VFPZAxwPs5XJu6nr5f+TUYl4Htc9ZbyQiFpb91v892XiXZoOYrRUUO9VCCOS
XJHpYetkhqALUg//3qjAtNSIvL34iRASfQrnZesKimgn7iaSX16kuTu0Uy8Z
Qpb1JVSlGIqp8MyZsTuqD3SKo6ve8eu9xCuxZZ8R+i/r7YdgZvtrYUqd0r0z
jTELbLzBapDBLXT2JK8eIg/tBH8ZO5gWqIixf/2joS4NiqYu3LSNXIjxHSKK
wvktrunaZ8NnI27HP9B7RooMV4PWmuFQ2+2QVHeNVXE9NBoxATnLTRmUk749
2y/5He18LEFlce8s0et8cCTI2ByuBPrazogeL8pscR4p8+u40GAMr8RaB9BB
aF3N7aETBnaQa1dnBmXZGr4tM56z2IC8ZwT583uW5B8YT2eUMju/8R72Zvs1
cFsy2YBb8qhHGehJD6+R1nEkZhFObJhFyWH5zqq6F/MB/guLpp28vChH6Yh5
K80jpg8J6K33rfEaedzW2A8y5wFd7Iem0jKLS1fQ+lyE1pV6rnlgUkfZH7G6
/fVk7+7ziBT2AMyttQm2C53DBCSr+NVkuKEgGJR8q/vTX5+/oH3/APXuq6Bi
Hs/kno3j7rUMSMWQ02ABmDZHxL/wfmwEKDQZ8I4sGDGuNKEyhTWnxpC+ZYVN
zm7fTs8BnRLuL4bT+Yl9YgxXLUT5fe350cK1SZH2/XStjUP3R8sIcEEr+4FC
ncgw78ejX0GjkxX1JlUjOndXU2tBOO/mFZpQbIOKalPvgzhX69YNRSJ/P97A
iN+2/r9vbYXlyWSbbGx2YdQSimeCOnIn4/ORNEpk4U8dZPOYmtSfvX+jmGO6
vJ02YrWmF8aeQAM23jmtwxW1CGWpijb7fwWIhOBf6CFfEzYX03gjg1eXTPpd
bggNaaF6gcl68hUhRvBpHczO8f0FtQy/Hvs89BadXsULwPvxXMqyTavl3NmY
BqrEWsTUYzoJgoP1HG5/0Yk7nuX9vqy/kfvSX0ra8Dw30OaRik1xg9gkuDnH
BgNp3mVOZLZCCLto50F0MawY66R1VSSdSRbGjnl0XiH183aZHanXGAyAJB3h
FQVuphUqkS1wMV8Pw49A3vW6ti+G/vbm7mHUI0OTi7xQf/svUE55FMSHseou
3YZN7jW/UeveCGTAtnSmZYmPEeS0jJMSiL5lK0XlxPhGPdIAxVq/0md0gPfz
OyBG5iaVsy7JDiOUqPW/KCgOIL+yUjQmDqqLvf3QsKOWnAfnQMmcw2tN1538
JDNjLOVte4sEpyVqoaQuewBrYs0++8PSvyJnT/IEpptWCXAyXpG1Bt4T5mB7
QkKHcuDgpDcYtxb8gCWfqhHqa6mORWKdjIwZuTzm7febNxyQM4jBUQV6HBlB
M+EMz0AZN8PUm4wKihb6sij0r571U8VyQ0vJ2xDw7I0Lie7BCnjzre5dST1m
3uB1aKDA6YPDB3fGmd7ZPRemLPctbLaaeTmwKI/+45hs0ZkPkPPQulG8RZYB
QLPz6HkjeGPfGB4Pi0ccqljioDlIp3z8wuYUKdHjd/8r18T4i/yVMM169wV6
2lEPVUwqbh0SAO0vvkfxVpSfo5Fk/HCKJQGSiqojrxXtO47MA8DejLiAEtGm
5+G4q6bonVVdbOOtY4LXKFXZeXcv/l094pyUGim9hAxqf3AH4f+Jo4GnCZOh
l3ywr+czCem2rUk/xYV280MQCr6+p+3OkxoTNAprgBb49iY9PWjRWqn1nK4e
eiht2bacbH2RDIwsM9IzoyQN7BMw19caUhrT4NUvYQLAbkdlds843LWYOvG/
R1ioFzRDYuiEGzl6vo4fr5pgQGNTTMGdjOHmQqGfKR+/DzQsUanccSuYabrA
+avSDJOICUJoQtzPJBKEgFHbg6MgUX35Is7ZQkWIsj2mQKsY8O9ydt1aXG63
Wnyryg6kDsqHgA4qfq7vG5KAo28sObe0HrCVHw1x7L3MTonupRmjotrzDH6M
cb5SQ0fspi4zxXYxBdvUgUIaLEj+znDs/doxm2hMZ6qT7xjQJ4jISMFxiOZz
seZ5rBnOs/R8en9P8nY3L+MjMBR5BEXquDL6lUnXMtoxt4UrnajGpZMKgkBF
elR33636vuThGu2HBokGzTNp1bwqAyYjN16p6vs4+VZW5nVorh6v3NSwUwcl
oaSPLe/W2Vh8W7wGV9CyhR1ew//ptTbKFYeH29xl5KqjO0yFGRkC42dwXfj4
CufK44KuKqNQ6VgpOpNp9LpIFas0EAn2Mhz9iVFe/MphV//dXgZ2pVF8jZdU
jS/LCMoZTzWtMzshp0dR20otPTFZQC0kcU7jyh2h6yLsbgXDlCmIaxBe0iNY
gOw+MtD6S5Hy15t428k8Z5aeKbpzpPip2ZhUrI17QDk/SLqU8TrUnUKraSkH
APHrQYvXhNFCtO8cQk+na+GKGuKl9RA/LV41Lv0q/M6NNme4g6bZH/7C5mzo
WLEbL8xMr6VGiNm3iQA4/G4IjyfJ8XtpM/7hK42Om4UQMRJsY64H0oUFRgeN
VVbrclYoSeHryGdoKDj/lGfCO4CxNYgI+pFWXNhPOIL4msWo1xfhb3zCJt3f
MYVK3GKv06rqfjLUxLyexakoPVJkkclHGye9b6BgbLuQuukhc5fsOb5T0210
oKE6OQjIfFgGRApd0cBoUnTJV6HE3DncSYhBAIsYJA0iPgdmvjmmhCzYISfg
gBpojrQfC0OsSxg5H3MysNNXK3lKkkHBnsf6bovU45sa+mmA8mkL8Gsa/DMh
67cc8EeZcw09yEvUyHFfOAgRQbXSDmTYl/oshhzmx/lrS8VZaggyisgLyLe5
h0qHPPhvb5EwuaUeg5daSusYuJ/iLOKBjOQX57Zkh8laC5dfE1ck96+s3HqC
Cnc/MK5pPxCDRY+cdLV9dQZIy3ZwLjSlPIKgMLHltcMAHOjDRh8WVWc33AQt
v30u6Ei+9aXdqQrlm92ByR8AMmeZnRnPO1NMu0DoYUV2t+qRkCM+rco1mXYd
ILPwP81Mpg43phNoRtMVPOW9hGCvXGfGv5ONOxCGUXutbzW9NxOvV6CdicQM
97acx5jUmd2rryKK9ZFCj0rCL3e2RAPpuhEtJ02YhcE5nA9n1JOItqyVf1ig
AmABQtZG6EcBwBhnUOeKAtvvhdK5gZyeFCcfxbBwV+OSZRuYYVb/0rYV9ibG
Sq71Vxm5mHGFpANobdQZ2BmuO6473gzp4dfzWtBGk9PfvA4wYUAYlfA+0dgo
tHUNs4kYSNdG4h8ubkHm3DhnWgpabfDCfXv0ExmvYjTX6+vSoRRjDRlb+4I4
U+TlgLPbAU6pK0Z0AvNMEqq2kIJJpkHjVJs5Jx5Nv5wIXNHKyRum8/R4vnUF
p8ztGYH24IZxVdRphHiVvEfut0ISm+xk1l3ySEAGlLFB0UU8JouMr127UhZS
4pJKznAgZ/liki3UXRluDgKg2J5xLrx7a7M/9r5ZSM9ifu0tTxPc2Pagild9
WB0nbrnsGgaOB9SSgdKfbb7y+dFQYdPfkFhKusaZoaPIWuHQ40PpCp6sw+2y
9KyUBmSXdaIpeXX6RZD9ULTx8o1vr00XD+o7Yr1v/T6KwOFIQiG0cNnzb2C+
kKYI3kS8FiBPAxQrTxHDElqXB29hlizP65gYtHfzv1MYGSQeu8h9wofQv7Zf
yiOxaSdwPAiibRt5Tn6l+9Z1pwA0z/rtGam4ZgEi1pKDGuF/dYK7nnUIUlbk
Q9pTBZczTiKZ0nl58PgIPzqAL6I50PVFiLejKZtVuX73utMz9tn7/om688nA
V3BuMb2y9F0qI0m2NoMA2OPCCIz/A+AJj2bJv3HPR4Q00OUgc4qIALNwp9Wc
dV1LEkcbulBjO4JxE9PiZxTZD+Uh6vtz417EHAL7SDdZvYpnjM+FVGNq4PiV
4AFftvveMsMmnJJiL/QcY07YsN6g/Es3UJbUp936djJBodIWZwBGBxTWy+cT
ZOmVvr3FEtMKEYjPGSSmfRPRxR8TvzCWoKI+hvHLI7fy+7vqfS6QlkLTuDTU
Sml13G97E7KGVsY6j2xjtLtlNa34s75P5Os0FS5VSmvJOdX3KXS5U/kV0f8d
21gSUyaTpEC78QXmjFoDvW6AqfQp48QDAr1TIeb72qy4XGbgveG/JbaX4HRg
JTFL3lk/p1Tj99efjpXS6U1h19VbJKaNDYdA8ZXphB46TrHbpuwHM8SJVRph
YHK/h6bI7Kt4me0KweT5VndB7JAHdYHVBymYuCcFS9XIWphQqjQoGVSawyU6
iy4kk1vBr7/AgnZ7wwQxcxgi46IwJWWhsj4LMD2aEKG9JSFdCspTE1xSPQiA
lUo84+yh/CIxlyIX2hJoQ1oXOSbllOIJnoUW/IZwMRb4g/VrcutHwFb3lqQf
0z22rbe6KjYH9mZ+VVdeR9OWerGZ/8ilcwNlzecJ59ncmldJKaN+2GIBpd+p
erSbi07d6UgPjk8xSPLngCJkCfA536WuKaitV/JoknHW8yE5pHecuOSQ6Qt2
mZnmucF3j0iujDUuf9b1dWIW1y1z2EotEcrmRExZVVLSMdMYc7GwHIyX6idy
xr3Q0lnl9QcfJ2Dwkb1pFJLucvxZJhIBNfLwzY+WXli6tv0rVk+OafDpL9GD
QKilpphZ/3dfMWd3yy1j5z0beMWXXBpTFmxP+HQ9tiqIFm1P9QXHKXqTCQbJ
c/Of1syqC9CYMsXD0eNYTFYBa9bcb9MYjxr8rylAL15U2tR/TfB9YW0y6DSY
AksE912dQMcqqGgo4JUBgzZdsAdIQ2scxdFLthQj0Rc12Kiy4oUFilsncWbx
8ao4odUzvpdl37EThAUiTD5yvrSGUmsBVahr7BltZDxMOVtQt9yK+rXiVewk
hwjRAmUHIYrphjfA4/76ctb+9hwDA0W3K23ZEQs12DYsDky2Z9s3DCDwSYsj
Xl1eBUZtB7TJvnfPeXAZCp27tc6twpYzYooGhjVg+Zpv2PkH7Ho2WknMeIV3
XhiVOBoKGbjKsDjBUCUcQ22Fopexjb+ADkx53IHSRJ7Ir1cFPwT/6BOl2aWo
TUqigMS9YPScQOrDeO7ZGKBGxA0CfmKSi9chof+t7DyIU1XSNjVzlURG9LE6
y5EhSCf+Xo1hVNM5wUirCCkP6FuACfaNK5AQ5u4esjZqgIRmPxgCror1D6Sk
wui+4UvKvbHTtzvE9BsfsMo4ch3sCcHoUetFNBZB9vXKJrZ9f3u4y9BQVbf+
ngu2RzDI9mdyfqm21KU40DyMMK1swuujRtI2+sFBnboh/sXDDW41oiu4y+ZC
z9o//j71CinyGhOapJOnRgLFv1fHyB1Y+t8gwsGOS+Tvwj6IN/T0f1cnFo5l
hWsyOhy42fJP0dldzWF4DMkHgfm5fKKFTLaccYBQE3Fc8SvXr1h0TrHt0eXl
JEYCjvtvW9nFF8ASpmXILYDgFDtGWv/QFWIHrvdrI5DHA+sGAj46GVxPA9oi
lNgt79zzkeb2gru4AO6jqKZbepzld/1avrZXslyvei60fsFkOFE3SR7f+eZo
Zvzg45Isx9iMgN/JSE6aczU29ftabiKDK4ZCAmUyWRNrfL/BSOtaSSCCvUmU
SdiOt1l3qTClfBdWrdODO7nysDfwhwEUaNX/CeK7qOqPh3JdBmJbyr9J7WlU
djM8q1Sc+/J4Qjv24np4RXIEbxwJZtBm8Uy39tt7anbLoUcPf8RNRJlJYCmW
trRzLHfOZxtr7pvBKDPgKdEyZ/tds41nO6FtpaufL/FpQJnc9XxcUzU+jXPK
fXUM6TOnnWiJqrT82uPyM0mq1kFEQMpgizj691qUnAJ37T+dQjI3ie5jcQQm
wq/afHsu9P85zz0DDFViRXOdlQ/z40WVmVZj87pgT1nHxRJSzmQjWHkRDQqs
tGU+WkP9TN5giIObVadupfjOaeJIfQsic4Lf54VrCJ6COv+dGqLaraLHahsT
hgn11TnDGrkWbC75hPy7+gQR5POvmxBD2iYHyIyv1rNr66s6JfAfIX3f2m54
KYtHUG0COHwzFmTQXykTZ6I/Ua40fvxJDMgbkGanC/cFfQiFrL7L94FXS5Vm
Kb26Om1nYnAOAKuK6oidbw4pjhGmPLL2vDb0THMRkKDBJwqaETEifYSXiE+w
f1SSVjfripI7ucfnYlkYzCBcizfxDFhgkMuKbvMT3fpP/TXn7bsUSdnZoDoH
wG6KRudabxS1SdYwVOQL3uWrbC5fQ4bCnwU9FUTT7Sx6gFYQHb3mFcTnbnZR
IFmjHSFrUEn+O/ef0E3L8o3NUzRmAONXoJQoCXD6nTLJ1buiUGetuMPk9znH
h7Yne6TNoDX2f/Ri+EsPf1qvv4YhDsp8i/4TKHB8FpCIWioL8EtHJHOZq4t3
uyKyJ15u/RntE5Bq+iIX5he7hvBcUfmXvQZVxUmJPSLgjUk26kfOgLAEX1Ku
BZgV+4jiq50+SRWSPy4venBXFPvjTQ2k6lnUjhAZTTxotZbE6vxjrmkt4W27
KvaakOp5Mc4gUbyRA8QjWoRbml4hmI8sfeWD+fnDj/BtJfls0JagpO+pwg0y
0ptuhzcudLYbMgHHxlZHnLNHrnyjgFc8GglTXN30XJNe2dMfGVe7Qwu8+Ky+
zfPrOjITQ6r48IiaQBiGhsAQdLqbHGFiTgzOj48zbin0JEz9Ifb/xpAxZqtm
+3mxGBfH1PRCmE0F0e1UavaWljnvbejAxTLmPkFsVEFkd5yFl786BHhcRKNq
yL57Rrp/BTv7tKI55MrOoNqZLfuWisJK9pVMdAPjeqdA3T3NF5bu75poaIGq
CW51Di+4F4639w9FOwbMRil3WclITw7vij9e01vWXCxC1HeleU3iD4ZPIwQV
QgjVE4tb/Swr3WyKxJMrbjmqo1EH0LMFUmoJey4pglUOQpQaazacZl7V97oM
HTTm3MrlDmvJ3z6XtpUOmUiPAi/0+uNYDjQeKRU03Fym2ogHX3fcr+bzEha3
tjpTb604PbU5fC63xm+Cf3UNTcoJWRbxONFDMopqM+10L0PPvKrlY3FTtaIL
ILt+C1S8TjXyXXS8xYBW+Gt6DS2/seUwEDNYgqxw4Wn50N/oBVP4fa+INNGU
QTB9acfgGIJoUuM/A9nslGHGHAZwWcNmJUeGe2lMVgEHMFyBOgKYDcfD29cu
bTfi/182HCP8HXs7HgSX5RYvAWSPbX81KalWNXZQxYOShqb3dscaZE9YnLjl
4ZQ5WKz3YlqE2u3jMsOcVvac9kVbTjUwCnyE344le2pLulmxoc5ShajZIq7Z
ju1hC8rJz1H5eKQRmB4czSlB1Avlp7/K931mZtzLwrviC1nGncpcRXsFwjws
3hs3v+WmhTkksr4ceQxWcdJ9dpKiLGdV63DgGwAZb6R/RV1jqhfu0nDnCVI0
adwHvaJbTy14slIv9m3a+BbfkUHsv86GB0q73K0nltXducUQcQoeMcPFRF80
ItRgbiiMx+Qs+Gst1/ZxE2rIMqsIlSBkmhwEjGNfk+LHr3o4OtgJ44xwjqdh
Uo2GGrwRrWTtWauhSWTJKI82q/rWn82YLIj2RpsrehYTvWSvqSWFp1kZwKa3
HRjvKIhIuNr7F/BFuIiCKwRkMA6RcfzdpW6Jqaao3C81btIWnH5vV9GL2tW/
6ctZ4HmHD5h7nUPRL91keGRpyqlVNzh2jMhuZKoMvSSpTWZAOTh1LDpbv/S/
uW+9/n2bzMqUC5Dzl71lid91lBiY8EL2LjukWVOJfWkAHSGUQw1TmmUdeEVj
gVatlJxTxdZOYimD3odZURLgwVCJe90np6zjbdJfL4tkAaYsLiTes0rURiSQ
9apu3czXJkNmEb6emopVS8UM7QqV6d8yVlQxUmGH79moXiZCob6+k9ViwhgI
qMI4QxjFOOc+yXLWroGZmOeeLQ9usxw8m/FqBRjncDtQRWGghL0wmqrCPvXm
U1a9QqeW7ursI1Hn+VRxLvPPySwpn3M6zyVTIPnJPActdr3m6hfwtV8rtArC
/23LG3A58xsYBvt9R5uI2bm3b7zpZx7MdytSxSEtIsiI+Ju4sUy1TMWVkt90
M+u9VR9W4vaNs29LG6mhCU2GRabDtmF3u/ElgKpT3e1VXwmLsWEGFk+b2EGd
VkzBSvc2ZxnbqdyWCWkQCS47YNtBn93fzdLFoxEpNr9KAcluzluTkbvy7xjd
98SUc/mCGio8MYL+7xptQcxFuJ/OzwBksHhPvVQucCipxIh/i3AzurGIpHim
qxZe/gO1Qv8OIsHBszKXSqaZpX/IPzqYFUIycuKvLDTmpQ8q1lgn0xP28+7y
6h9FkeKnTe37o9PmDQpCT1FwS9wZ/B/A2WGdrTHi4o4TmT3Vxkav3gk4szpV
hVmEr6ktfnStbXj0fui6lUlHtpEMyWJ7YfAnnser3hlKjCUiZDYpqtxwpAeQ
TgZzs709iIzE1xCfqivZHZeZAwuco9AaFPEGgRc7NBHk2zrj3QqVvfJ6sChU
1V45uVTB7R7P+/FqwpsLQUugXf0YVeep/cw0WpX1h4P8Mb73Z3UlKjiO6KR2
IxK/AfYT8iQLwHZuQxYxJLuJJU2xT+mZ9ZUQKE21/asQHvt1kgPcK3RoHgaW
WOAM6KoHOH1nYaxv2io6kb6B40di1/b6TtDWEwOYzWrnz/a9PbwNaGXTKBJB
hfrpjcg8uxUQ09sX8pkZV7I028Or1uFhW1GcVPsvXNYf/j641XQFy5J08Yp9
ouBVn72FNLEZCRMrJWkKMBjh5wuB6zIqAE/CiVIWWXoIGvdIidtu2nVbuyBb
/4rbqGnF3O+btiHCCkHHUp3H5p5d2rKJlXHfp2kMejNEdxKhAaFzFOxGFQl3
aB09eapfGx1yXx8liMCSujCE26H7hNJyMouDC7glGIF73Z9bUTOibtCGs4Jz
H7ylNeJ5+QivjGwHiXxG1dgsGJM+wKt1OWD7lk46ODg6mrdrC7U0J7QFf4tr
R9tcmUnEqAae8njYkJT/bAnVEz6YN8rulPtQre1rHw4pSm7ki4Gvp2MV1Tcb
gOEJcnxVyD/xmSbUlIipxfxz494Bp2J+BMgrZFL+0yzGVP8sMHdJsk155Ch9
Du0Xew56KJykky4cqOcg9ZtWBIlpuM1a0NKA1StgZcC4YufXoR6F16QXqBUG
AH/3AbF0bXNwflW3P6G3sGWNIqH4Thylme2+M8PAPfg/rMr854Z+IdU2Zg2k
xrxqvRSCZULWhYf5pWey0pcJz32w8V/LUsDTyUPNeIa7L2l8SrnDK9ufKEGB
+niVKDigxZfDiWHklob1WHVf4YIHyVM+6NUiAaAG8MsFLj8uk5xguKVZBZSA
iTpcq18uc9M0e6vUeCHaaYKRc5fTbuZA7rpzwt6ddKXmAgr8WiT7nRvb83ti
bg4FP++HymtBzQ+yLytK5PV12mADbPPSyYQg1rg8uUNwx/I2n5xIpN3aulpl
iSWPIsyO6QNFAwh2tWQ3B7LzGoAXGs8asVsEJ1ssUOCqm0b12d5n+arr76c1
j+fFlnBcP+BmC+cn4zaeT35qGt1l3QrnMRH2WltwzGbFzZjhT29F/JiOZff9
McT9V7vL9XEjgHycwGHDi8W2c6DcI5hbdmFRz8jc2qbYsqqQ73aP/x2HIF5c
vKy0jQRLqrhayfy0IyIrbQTsBuYpH5eTvAEGBh2G6NkzVusuiUMxBWTcncR9
i4/Hom++1guh4C73jjocVGxuBqywZbviZ5CFFaSBtUu4/GhGPmH5sOLFg0mJ
2l98MhPnzTPA6P/frhyX5BerSe7njus6RrWIMsQAtt1B4tr2CR+l07y5htCz
3C1o/yJ6OzmY9gv6LSfSnytzE/qmV9Jwj1MZ3ttJ+21DDzrLV5vUUd0qS606
L0TErLZahx91QXtcFtPORbWr0QIeb5egZdbtmobUR3VuDRNwnrXsmRW19Dc/
X2ozmfH5ansHxg/oeeTTnCAToWNJZkxtZNTHb4Xsfk7cIlwOTQBZW3MgeGPj
pSS2jPYes14adzGp/sSovVGmzzvSVo1596hXWBFSGAd4tE+k7pszb/+cP+1c
3172KENqTsSOg66Wyx+yaBdbMxr/cC4XJ8P6Ap7o9iPOWDfuut03rvot/2EF
MYAmOSK+ZIMaVTrp0dtlFnEAVjF82LzAMOEVyVxCwiO7qspowld5rmG4yWk6
EST+HDpqWrVs7yKeN+gT0+vJRQsEP+stYUCYCqqAQPsHDmtcczQ9PhlMqiVb
Lr8U9aKF/88WRTmj1mpEYiaCfjsYn05ZpPOb//dpMgfyXBI/+iKRfw4l+ref
z3mRgt0p2w6X2QQ2nPfH7GsJrtBN1FWOSIW3hgAgO/mFAYQuIEvreMB4wUXA
UPzT+pGNpyGPABnIr9YrYykAWcSWdMZ/SDmlGqFQ9ix88HML7XjTUIE75gcd
KvXi9O3NOIKM2FZhi1Pt461riWQz1qywuYJdl6fgRVdAcJoUHykp3y0fv8cx
0fZqjWoPfVuIpksXL5proVlGE9FFijQIXo0O4l1O8ndbO7RuiChOuPz6cL8k
DhFuZ142uJgJg2DmUoJKdj2JMthKC7cILTO/vTqJMj/SoUE872JioKZAqRBj
22aEJW0e4Eo5Y0l4/M6KVG0Z7md1bHNBKMgOyODqZknnNAyjUO3sGmqA4Hn1
os7+cJOhozozp2so6f/LEaj0S8/NUrVVaL5Efm6HRtpwrjQnRnPUgCzxZP9S
R/I06kzhMSKCMzDfwKjYwuW3cHDL945VnGd9DRfPVDA95bq9e5Dx39sfGIqF
dQAtQUQ7/ekvaXlKblCmSO0JuDZxjkJeIFVgU6BsZLUYJANKmp86GOiYYgtK
fSHw/PPQ4HKkZ5VO6emvavXmmV5m84EWr0cnOGgHV8ISAE6zWPBuXd4KO1mr
nyw8SpTbwZRlDnAshi0+Got13nZVOpwTB/0j/wJ6BDMWLAKBaE+YSuw5oBI6
oUh8AVQ4EnCXn9TK0rfJDteNYt0TAPK3Gawe049H7k5D1afDgY0ER4OjXFe0
706hbBFJBI2TpAr+nc9QXPVJstzuVSpy8FoQhccsxbLu/IPr2V/GTiG7Qsxl
eJyEqy5kQtyxDjL6MwLcHyXp9pz3qF9ilovxLapXp+pYd9BMBKO6MldWUGSx
5jIzptPt3ZfZUfV9N5n0ao/xPRlo8IFlY/gqtCqjWFQx9Fo3E/1qG/sibC2F
6Vq0IjPcolf91eHTOGq/Rwn11CWwS8zWWnPqVDirbZhmKI26JQsXgUijbqHI
+P1I7AwpGINSZGBLBqRPliGtRwqqU95yMAEFeHUW4N3lIYYiye2HTof3NeXJ
zTNByC/SVUOesGbziuLoYxsvt5wVm7YxFl+0xwQ6Bfy84/m88uE9eeJZ6xlH
PI+0WFWxDKfm20UDQg1yq1Gv9vbzhoaUAZR6r++sf1sd9uPsm6iP6hB9csEt
Ir4kWpAfyCno09ooKPDDx+ttD1hADeJciCKmcWxtsoJc1kXyzl7HSm9MQBpV
EJPxBBw4R/rcNj9YFl5gjy1YCXmPr2GwlNU8g+pe/+YTkz4QcTJ7KHUw4Frx
aL6RsfTMU8aNzZOKG/i/Ql/C5PwbnlFS7+p3sQHJu2hgLGVOOOfX7kelBCW/
eO7kr17lTYnReOsyuzv8AY/dGa3d7Efw3328ABwYPZKT7UX1MgX2mmSmZeoZ
btSaPmu28MWVVpp75W5CMUPibEs1/+SsTda5jiKXlTeagnMoPVbhdgHxn/2Y
vHVkMRZG5tH9OxbJ4hcDcZvaCQfd2faxx7rucjZZdj5O0FEiYesmPReJBeO/
l5fiucbFLapNSt6plqRLz7YrY5hm7Bjv3FC4V7ofXxavsp5cXBiVmekLjO9F
3lTJYPAi4ctoEZgdUKuW1Mn2S7udREieeZ9GYOkncoQzh5bYbyw9k2ir3QOB
qkLDb0ks0thrpA9Gtt60bq6DdW07ZQNBVH4DotLrBYlMvsT9XYFdJ0z8zSr/
rQpI8l7gUzDS5+uSU7rkkKMMGOJ/7s3uOVJPksPiwxaooIW8qpHnPJi7yGsr
JkY9ortQlbxvvk5kvWgSsbs62u13dCo6qRaafAmCom8G2mJa5UuV7oCVZr2+
R1Nkn9VqiRVoifhvKywQiO74gjI0iZsH7wFaOunNnj9G2HLRGqVAq769xmmz
eMPqoBqcGymjcdUVS3TzPSqjd1UpLitZjScZulRN1mhdK2iCjR76DowIw4ah
9KD0ycquUplkxSn3RLJaDqPTlBNR7nyGfPXqiI3ibjvEt4Kvuj1uehGsJImk
MSSf1vOAoJn0BYfuHgu29UU4ZTmL+9Lr/gpV9rvYmNQu/HrZb7VoMt2cwo0g
XHk+NktKUsvAp2qLb2GI87w+gHHCTZd6TUbubv6uVTZfbFCUBE/gxNaDMehS
0yNy5GLBjM+sYEeM4PBnseMU4IlG4EgMwN/k4m5pNuePCjFrdIKsWQaE54Ln
s7GZ0DvKOtsrUnDegugLjj5TyU+lWSS5n3VHXnx2psZ+MGFoHRPOSUMyEv7E
9uJoqkLpOb58qN88FNrmAc0UpgYk/VJBM/USa9yJmuEkkR2Fs+Qs4MomDbvT
Sl88Hw0phtowazhZLIIufN60abFi9WScdN19ixcYCk9dkshO9T1C9uUb6CwF
ztYHycCQjM2skgQUMAOebQXMwZKCNHeDUNA0Wou1TLstMCx3ug/dhsuDiLKj
o2NJn0chcGPXvrIbwKWv00/OuipB7cPi9aNSL2Ew1wEiXk3QPdKTj1CWKPKK
/u7oHHqVkf6goelYImgUppwxKBwbfhg88q8pcmeu9gN4pj6KyTPsVDoKojTn
ulrxn0ToSydSRSQ6nYASlkOZuEtTAHSBgOpGfkscCSmEv51X8rGML7Hu3Cs6
p8/YqxHLgTyhffOgdScqiQ8vDbzrwyePDb+Xo4BPvEPtpEU6DZKtq8AUm549
8tlu9p3q20m700Fi6QdWr2PmGK9wdsYhwoEcReKvAMNH2Z18uhNwaOiMqmCx
l4iVjChdErtqvDtKQ9IwqEwYw2vp+KCsDjQLtf+DLTVdWGptc2RXSrXkBPTv
bhYtaKAvMzz5fSB+YQZvnbGGp9+GCG7vQ40ATq31Nakt8DQGzd0rYDTGmEYs
gDCXZPW4QpLuAe1Ptq/efVNy356N+uCW/jE4f0g1pKz8/f8I0RtIbGmZdW2u
FtzUiga0UsWVRC8TiXHXBgfC4NMDUptP6xDJUvsIB+FQD6yoUJqiHTwKYg8e
7dmCWKt2qgmsFISAPxPLLqAReWdnhFcFGj3HIyhJegJXddTyc5bXWYQmyMiF
ft/SHt5cFWhcB3DShym/4q2R7U3QxfJai6KZneXkVJ/Q2RYuNq+eWoE4o4XQ
KUQ9Yhe9PWj2KU3qjxv9g7EbThSYSu7InbKTdTFO36Ls5cGuypydzDpCr/kP
8pDU75IXpwUuzOhwC9FLsK1oqQBLx0lyvb0a/N1JDq676y1NT90VKP6Te9g3
dpxJkrfO6xuyfup6wLql23CGr13pgQ2RnBffpYfq6bet+YRgTYZF79xsu6Vl
7uF/jRwtg6J1hvyWWTw+MzJRABaU2MwhJT/nX7SLMSI9Nlfad/DHfhxRXaQL
B02tfFabyLuTB2/DTYgons9utpbRP0Wt3WXL7Jhg8vDUvhLhwScfEu8sfK9/
gObIPZnpf5zo3zXEJa+28dwnKedOV1FtZ4hWYL/EaprpeaHbwtFg9EvF8eaU
SkUR4mTAvsf/Q1pC7xVe/VZ8arKW/8oY7/FDz4C5lNLBYURnMPKA1dowpKUx
2LHXnl91BsFW8zwiCPmfw9Na1zugVmA0xLQjNmexsxXO7xg8JtfdxR9sb+0c
1W92B9W9JtOlMqMU/ADRtVQCI1AajT2WttOOv0iC6RUf/Qz8agu3ZlchoBmH
c8I9vKUpI7pUGMseq+6wObD4p+ZTkHHjnr7r513E2lltVtuvN6DGfs6mkCFV
0gn3ByvVszHdAA57GExyxlLSosA6Rcn8soKTS91TeoI6O/ZbWZJqO+YqvMiM
hHYkcCpV5t1GlwVb5xCo8vGrp4+fyzUXAOSrCrW8dCwse8VusUXkF719gno9
tUZiyxdvWgv7yjuwfllSHc8nNXmg9H/oRQrNvVZUxAx0bOxIL6i+pMCYEl5m
LAzb9z2CscyCATgIQygL1XV2N2JC6WQ/aHPRPwGWWq1H0wGJipNA4m93ziUV
CNRFNzPFqTh+JTwoy0Ievvvt6mlQWzFPN3qm4Fff0l/Edrap29Ybu4tq9gbA
rXnNqdP3dd2nk7W9kUlaS0EA8Sbtg/aUbT+Y8xYoq+YUJNf6LV7eYjAqZ53z
PyfyawXCk8ILdKswWbrD8bENVZB53OThR7VMK1Mlh2S1oEQ/VG2duB3HkXYr
cvq5w4ib98aoyXvOxB7aJRdh5AriiZbsynB0aTcQ0c5d5/h+Nt3iZ5VinzvN
Y5N2oHIiawNl/SQGLXrRgqava9QGEaACDqZGARC1d+SI4JZfkbXJtHk49A0r
Rg+XhnN7axBNp1kdqJ16P+fxMs4f3+TkT2EH5b8V/dHBoSFj683DWRhKwIxK
/DfBVhU75YOgulRpJrID/U2fxtoMKLdkNDgcWInecbs9ivY6ELPV34rscdGb
bh5DahtkjWWCEItRyhalelyDfV0sbYqMmF2dmEQC2yHnxi6VOKmswJQPRMFx
5VuwSqk0xpg8iUKFIyB9c6yMO3DztWjdbYFc2PODc1F+oRuwjcO7Cksq4M4q
33ZYBJzgvjmF2uHc/s9UFBsOSvUtajfdpIPj0CV1AfW4rIAED5TCPRxTKQ1Q
5WMKrHaoJvq4Bt7dECJqnXJsJx9Q77Onz3kuMyQfTHPhh3AiJmVsRw82P5w+
zEO7+Ff5tZrO13/iwr0HjbqCZ/UIf0+d9gP9aV8VSOJfQLL49Kz8j/l+CJ4B
rudjCMaT1VdyibQFZbiEqn864++4JZ6GAQDBqMdGgXZ/6p7KNiPbRICfN17u
+XbfKyYERKEWku9gWvxJyAZ7xKNcNydzNOvDn/S9KuCaEsSU2tyJKxqw1vYV
tM/qNgxSvTjllE7p4HifdTTeC6UzZAg3sw6ayhnYvFdvXEUZ58dgl1ZZBq7Q
Qr1soAqKUPpHxH8zmQudXBLO8wC2c1XXHGguABC3c5D01CjExnscsO+rXS5O
VDTNbCd1OAB+RLy+GBlP9zr6gkXd6+FTV0n8oiirD9PwpXKmNrrr86QACiue
nq5efSKFPU6Cs7CP1HG2KeACwPSWCG5/erLs76nf6dQHtb0BX6S2GHmbrGLI
qrkqQ6ini01sI1Ln3wWFJ4AqARzL9v6pg5Ap3jMMHZg2mMYI0DQs9NiAFMmT
j+8G/dM8D7rcd69y49sKWER7h/tXLjMgYOUDgw4FlFM4i9jvrvcVRjRNO/+C
vTG6q3pueMvOvZY65ePcYUGUWamZcU/eAKToMHTsIEQ173IE9OlSHDpUYJ7x
1+AuKMCDt9+ZtPcKdp/+VC+5pBOfiBFIvhaE2lyY+TrsOWZSZR6HSRAXSBNP
C+t4zzKB87vbCNrPSqUKTxczPP4kWTM1DHRuhCMKyOpiMeG6LBqvLhyci2kO
wgb3hm4A6bFZXZwxy+0GNTMj+ZexQ2idml41EvwL4O0ad+k9NXpP/EfiN9SS
01fajA+9xo6HbzR/Am6QgxwNaxmTTXj3IKemqj99VUTwBg+6n1WXv34dG2sP
T59jIVSmv26Q7ARC3sznirYfTSezDXBtXnxFab/tSDXe/U+F53Qdz6zLT+0d
4hHJG1+n4Xnusv1tocvDoghN05awB2tYTuV/jXkNcQCTU2eqoxIlgHArU60f
y0cQ0kk9dw0ozF0x6Z1T7WS756/58s1FHB7hGECupyHb1afgUAbVs33hwq+o
MCa1GI7XcaXtr6Ys578tcLFu9ItFG1Yq8jmsl9O888NjA2rfVOV8uZYAOme7
b5vspa81IymMWj6GYEpcVjqI8W/xgNUX2kbHXM72QrddXgXTzTWiATuLmpvS
62tPcG7zPrwkVZr3pFgKprigGs8bqnDihlynwrPW2k9nBgP4y1Sk+edjU+6u
Ph6E+p9KdN4MiB4a/zU9sqbWLDU/+UPwL3P+BB2F/AfzX/KrXBDayqs1S7a/
1SRQ/9Y4MawJ79oq0VvwS6ibxENJrnWLEtQW9rZKPVsWXSZFtI8r53IDQyTA
RDmk+P9F1M/5pHx0ZsYYW+x2lc+tnnZZZznAlRLafWvTGXlJ5cr4tMNG8Ewm
whXJvPuYKpZ4bH/Lf8KYqYimwY22lUsqJmnYcOjFQOHDSAdgTvNXKJP/uM+W
78g81G9h7PiTmnND+9szwP72zMmR9v+Qb9IYK00VFS+M4jnSlibkC0//fKyP
VpV1bwLxNDT60N7ycNZhUw9WkuTvWlRX7+1mYCRlL3jxgGP/zNBL4IIMbEWa
0iAtMcEhd7T6BZ2Jxx+ujhmtAE8RyMoSyRd1igXtGAK5HNYdLwlXz1/N1+hE
/BIOy76FgeKxN5Qq77rJ8FJudloVbbpHQWbJy3b5zWNMMbz6WZRKbUVM9nEy
Es6KRSHMMiaRnoBn6mzgrF+X01L8HfWV5NMhN7c/6JgKX1GeXWv1kYgOvry3
hYMjNqFU6vdsptaoBR6I2jJyTijUR07OToyC20eAr5sIdA9MJo0vCTFjsRHJ
v1S9LMD3sftDYXULRYzM8G9hz3+OWLlxPKZdmEWmNvsSLTwvC/3ZqhO6CG1x
QZiOK1JwE8UcuCm3eo2dQw1ZU3rF6Tsz4gL2DLyKB5PWnoizzZbcJ4pmMlO/
97XtrnyUdd7CePCJsYaKhh66bigXIeE/qEhwNJS6nhWJOFTZ0EmVCiHxpX6z
2UopohEsXtDf874aMx2QZHoVmd3gcAJzJIwghPsAjFGNr82uF6va+UdN3iBY
s33F8qK1jJEzsT8wKVOpRBkQ8swd6SoBpjgvpF8oozXX4eWr/h72qpgqiAtA
P4b0HzbQwLZDqU8eUSASfPcxJPgFQImX7rkNQKWFlXHk7aIrqfdwMq0bdxtw
1rnZ9Sj76UcR+EuzIT+dN//AIgkOJTRX/awwIsmKxbU2G9z7o2NaGUz75xv4
nrSEMlozz3YDS0e7eZgw/ixxJz8Xjt4iL+bA1p1itGY555v3nikE5R8nLi+k
5KcgaNVZnQlWLwMYyQG9Fa20gWAUXkCfZocdMu5T2zJQeK/eQ5OGu2GKY0Un
GSFAgpaFw/1xpAEnhOOaSC+XG9I6spond83gDAkREnAl2/6gJVd1N5ZAgGO8
7sz2lP1asnK5M1gPjTD+Ip7VTueH0xB5hBEMvesKTnDNpzr0aEuu5NKwx0GQ
FWxOz3kPDxriqqBbUJGvzmPyGtOPjkmMjteUFqrtZ+NvNZVkOTZQr/m+kEL0
70a3SBlQiR9Q4VF28eNi+x4vYcPiarB9YoILEuTai20M/2I7FWyXkdIPjlPG
lucIm5Vkoo/+hYS+sl65vabLvKqHfhwG3ScWWOBlroCvqT6DJPdRt9vC66wU
n0JAuWRboWZ/R3k8Kv8BxelkVYIX9Wd/oPDjCUDRxXzx5co6BoXKXWY7FsXN
BIaaYPU59EllglFfsm2Xyq6Me9UI2ni/HrG2c9TqcSg0qYPMxLuHzBWi6LEt
IOTx5jcl0X1SqhJgCjDr1ITCTrQwJPA9S8dbQ1ijwhYm6xYaZ2kNjBZ76kaL
ZXqJYq6UAbmzsdvvMyiTK+Jrlyl7hv6Fk3GxuSAVOc3UI98gm3iEm5AvdIhD
bkSj+RHnKa/+4//OW/GNIv9PVJC3FEZGD9W9L/Gfxxmi4fwVtfnqnYeUZVNa
bgdqBW2jCglwdFfkDNKNmnAc8yzJSIaGiVYCfIz98/Pjd5Bfwj1N4Kr+dXMa
kC7kvpbcENaoXsKyIBr4Ef44wTyUhPBW5WZjrBuMVzznTRfSBTpy2RDyVBMn
cfFOv6Ff9upW5AUZ16pPUTLjXGEaSJbYCMIsQcCG6RG6l2axfoMRctdjTMVE
7Nqr4UJIbSu2ax0/7074W9edSQZKzNi7yaT7dpaYMz5E2GoAOnfCZHipjDsa
Ar6zZy6riC4156p1xN1rSOTDqyvkuEpGm36B6UovoakeAtU7ri9ggBGvZCOZ
0qjjIXOmlGHSgKYS21mDLSXKgF54C/LhOw1bnyYVmxCGO0hU/ixKWHN44y46
EqgInft1pEnvsYc8UXIiC1f/hyC3jh3jg3A7VCWcnf5FET1hXZAShbNhyIdZ
F4zYrBGo20iQSUJhBRwSUgG5kT47E3tQyqcsogaTFEfvHZ2gs/3L48wzcvVG
GMufvCmcjHBu9zZ906pVP/r0jbiXa/HJ9QHZYa7bbtMW0sXt+NJJWEj+AGRR
Lfu9ZELoWDLScsu8co170QF6Rvqld1ZldljvDk2+JhKIgyw0RoFoHq1WkfwQ
yUW6FFw108eBzyWIOcP1E3FZnxhPIvvhg6HxW1+CcPrkJkPBIuNsMJqLg0Qw
QJAhZKeokvmDokyujs9wG45/abQe5+ImFmqzLp0w3+nUP0cio2SCfdpsu2jz
0ImZAgIE+mJwfro/F3SSp6hFs6Klamj561+ot8vJj1CIHMklMM5+ksbkyKXF
SCN3LFVizvTyDCFsqy4ESiw1V8RhOepSZKi+nvt5Kc17O8yPQqwAYYOzzNXx
90UPhrG6wyDWlWlNKJYxiUhLfwcOo4XYb4jRg/3YjshsHfgW5Lt1meL4coIC
RhGRHC/fcNKJTDGmQdpWLYttviCzSSapvsbP6b492LhEIfgqwukYVkk/jkoD
iFhrKe+Ne8UyFjJsr2bwaRwV6yMOU2l9SIvQCHqZnG5XlEMZKttLApG6Z07m
PTFiNZG8rJr/xptt0kUIsIB1maLTwVS2yHVDx3ftwdQvYhENR3EMSL9S2Eq0
+vKF4T8fXN5mLgyx8gGfNHVeGlPbp92YCQGoOEwjrSPOyp5DThUiq1lT5ClQ
a+zO9YgACBknNxLrAEFONfDAQ8l/qnt1THdH111M5jZmRyAYQnFweSVdrYkk
Hf1V29MBfmkwiBvEeaxG1oOTj/xW2W+mUgl8PWpEKFU72B8cfdC4Qax3y6ew
CsZGUtxNwZOh28+c5Pu+M4w+XUCftNgZTBK468UHwxcxIMPNWAFOxetWCqgP
6N3gzEW9yLIhnokasECCsHLnsIeJeQ6DzRliQS7nxNw7pbz5RmatQvNidopc
68syDQzZtchJWqtU7YWC8BJgSqvKGvg2+KbI+eoNjHT7JLKR1mqvKvOzD+CE
fY61Vw+M6xJ/KHxD8hJ6h3AIDv6h3hPBrNKrrgEgDC3nlJ2HgZ8QaXHIE1Dd
FtQZtFpggoeQ/JND4oo9lyYmNferUCWhRYps+H0OYxJnF34BK7i002WaKq4f
OI3lilpampYd1apV0CCuk34EkU4Rjn+8Fa336JscDocEAQMSuKg8Dx1tjw+0
zJ2NGUJjA6vEY2xb4HBKAvEcOK9czRhbeltoFHA62ert6kK49q296YdXje8k
Yl8xkFCKwml0WKzvhSFgSDA36wb7jVKi+d+pbFZvDyyxrMDCrfmRY5Ysb7Ez
29CRRSPQUF0UWbWU1IXU0fZG1iuuEZxG2wPi4lxoweSDtZh04lzN2DRFIb1h
r6/PdIV0Hh9ceB3d1p9AYHeDEhRfMhRtCjzDqyQ5Pn4mP4A/aJZg2T69zRxP
q9M+1kJfYnmm9UmLXLoX2CAAd8KfJsO8k84E9g01ljuavw00CAfv6fVm7QD0
iuAKkdEnkyCw2Qu+SfHyV7Es1VJuk2m3P8xKART8VpNZcxXUuLbq+BvvkvNe
e2ms9ZXcniAidP67SgaZJamjpDeyw8tg48uHSbKQKIIkl0uzk5LcbZf9MxnA
z89JpvWJ0bOlt7PLl5/++ta73btM2HSGe1lCby0bW1tOxFuslEAVxjssm3km
cQhmtgzcjghZaHnasVqcpeKagJVYPMzzqYpSp1b/LNjTJpXnCmPlzK7nkRAR
w7UvBtsIVcv/thMa1a+bc9oLtdiRNJZb6qyLppI5l/AQ8aUVH0TZ8x71rQFr
7csUj5lYiA+OxP2VsFciXXZPlWcZnycYw7oUNdTWNGiPrWff8A6L3LUSTNWJ
JfM9u6cTAHa0iCGy+SgDkgnxdkd0X5fCCc76BVw6RozE7L1NhiNvv4QWyck0
vnvSbCYmEXvMTaXtTlA1vwu7u7FsjXEvN05LEVjGS6haI2r4UVdDfRtb88eO
NPXip20PbuAYXQutbql2qZxlkPlfkIKaS1HqDDIT4t/qM8BzVZxPbFG551mg
ts4UVXVyOJGfotsG4wuFv1vMO7+VWYPN0CdukDmjFzsDy6QHMlq3VR74BvZS
o+Zg1v4HEGlBMG9gHiOKQX2LqAZTF9TpVCBd5S0J1d+QSVjimgSiAm8E0j9S
ro2WNjLtyO/7LqmYSs/T/9fdhgWEqSp/wpYXdCagt4vM2KH89nijN1wOVaXG
txyP597/P0o6gjwTKNo8027qmyqBMaEq6IArU7YiB4swI6IlCmHhWZy4va53
izc0s0vW26DHM+gIzHi7OOj/iPUU8ugTTWY7694vHbmnYr4+LEYfxMcUQA1o
gTQ9Tstut3z+47BOvAsR236LCb3LFkI3sks47KBSLMGvzfO/QgTC2WrXAOR8
V+lj3rtQhyZ4Bi65Dclj5Y/s+ZH9IQwf7alp4CHGxa9w3yIF65x66VgRQsz4
ea68c847p3Yv1oeM5OEO2xAF257rB+LRrsgFHajWtQLou+wbmALsZDaU6JH+
U8WJUOPjExP5RaBj5NNRJaIFl5v2O529qxHFpciy7mCoGEMvMxerNywMVuJI
x7XlqpvEVwULnLVKwV3qen6gn+1+NAGr/o1DEQt1uj15ycfw+vZcyIAj1yY4
gJNfLGyEz8BKYTP6LD+qfoRQAHk3HsMA1duuxDA3DVaI9PqelXE35DeleBZY
SNYbdqCxs2pytMjoaQEuLPdYlB//+Gg1ALCALo2y02SnKF21dICgEv4UAqqP
0W6YDKhwR9cFFyM7mgMOojo6qaEWjq3ZtCY5wx0aQRMCn7BV23ZjHorlkOtW
d0qvl+Sfdg7XDYmlGb+H/U+T9odVOAMlts2LOz7n13aS8tSugByVSevAgoOq
1xCkdbF0HaL6gUBt2P8DnnP/UGpJvVs3P315MtKA9/UxIJ/DfBAanG7+fYEW
kxdIqWdVScN+og7GNRsxbi9BjgQuX66X0mPzhqmWY/I+RohLZWLjR91e/dCZ
F96rfEyhWjBKjzkI1JUVZ4CFrRexsY3n3aeX4ChfIijnnCoXUIjcuQHqmHCL
o9wciJuFX10FoS+skswB/tkiNmNMC40M/GhfgBe1+TbyGfzz7447TGiPrIPI
2Bc+eOGomTCEiUmqqaCYI1PIHfDDGIZvB5qu5vQqtLS9BZuJ4wZxFjoSGflS
9YWhQmrrWXFYu/QRhOdQTAKrEQomvsf3n3nO7NkMyJZ/skwPKrIf6c3bsdMz
HeZF4RkL5Xw4SDYddf14t8Jbe+CA3GME8q80ZTHQGe4SKKWzQNVCeP2hqNeq
9omcTLOwjkDbpjaKbGc+M3j7zJB62nx6o3A7LmIYpmnwpWBQRSZsUEKl+lpi
gsM3139OBu9P/YH4ODT4OmxhVwZcoCTbi3IR2ppnugk8/uUJBo1aQI7Jl3nV
Fx9DnSnW2zXWDO7Vtb/28Q1rLO4DOcVVSR/KcDqRV9ebdHTyPCtOtrIaNREU
JN00xBSshk+p1n1hwEw+SFuYMnpFBgko4mGNXwHirDCO4lH/ruLq5ihdJ7zd
DlSmRiBqo9mR8BM+bZ/s325de6xCOTlrh9Z1HpjwTq0g7rb+JcqhEYtjTD7h
68eAv1Buz92FlTOepMDsdq791Hk5+INynHfH6apoNDPSxwkNDRgR/0B0cDal
ki6xI6UWHg6kXA2DXmZIFUW0YWaU53+p4YIFx6BO+AMAbCt8qZ4/KxuduySp
MylUCDMGYBzBqEig3CAI4iiPfTX2tCoM+fKxZvLAUDya0kpoYq8cCtFgONIU
visfGSDKCVG09rOZFnsvusbRQVCerFeOnbG6Ov6MTeHJuLkQDCnV7kCPeela
vtDiDWaZ4/Utr+l7dTahZFLkPpiOFS9YB2BVdwps54YT8M25hTcBDZksiIuy
bZ1m4fuEH17vBNu1sYfGLzKZN++JubmZBIFhVM9uUkqffBrlMxGx1Ttl3aYH
pTIk7xcxiFdT7/dlP1C19pxgN5o528Kd+wQ9wBDFsTx2H/qVMalUPPtNGqaZ
a2DC3asLcVyMO13crgNonWtGxJgje0YAnx75BT8FWK0e9a1lSKNSrymKBrPb
RMweT4nZ1hIj5Bfve8aZpyJ+w44AUjIJC6oogeTKiALaW4x/xD2LhOrDUZcD
nDsvEuwck9u95VMerVCvBL6mbPM4W+yWpj2kBiqTXimtUJ3cov+/QG+S7kMv
JI/2td9smNWYyPG2IYomN5tDKn3bVqmYcubBk+Ev+IoPTsBfcJjBAti1So5t
ous9G4T60h3M6lXBHAlhCOVfhlxAxD1wrJH99c0sNPaRzyRkQsJIUW+pSHth
DxUiQ1EHYLGPDpybvlmdGNe4S/b1Iw/UBT3T1DsnzAuC85hhnLX4HAK/kd+o
8CFlM5MR/XePsHplBHA4SCHiDzApWB1sNN9KMt82AlchtEhoPIyUT/sWBnY7
FDbMX0sRf/YX3363yb+iaB4ap4Bimr/2Z3N8exCvoY98Q5mFtXevQoFuSOML
hvls4tLeY1PKGkTgoM7ctvfvGE1QCoglYB+0OuE4r+EgOqpFtV/1/WMEwLqg
j4fMXBz0ei+NM79vJpv+SZNtB6giEPKH6ZolBfLNiolb0Y0jSYRqcxCEr62e
F/xr9n/u/nZEqrbxyZaTage03g8lCkL+gxTjqDp3Dgyd3+1YpTuLplowRpzJ
gfmprpHWGyhg3yNzc4clRT1a7Oq37VsgCDIWbJBbViWve5lbkoHxi1DNIXba
79zlCm3zgQYQc9g6/83AxuFIRcOmdbjdLsRWlKjhq1g7swmC/npnZt0VKxWq
z2Al0U1IoriBFyPrDLv82sOY6BqIXb+Rrrh9OPBw6tN8QyYI/VOuXadioA8s
JIQSiWl5dmnFU3fdaVCca9Vo48DXiLn/PK4d38hT7XbBuEWRT6ohxgiL/OiE
z77yUbHwJr1jdlACUtU5H7SADHh3BaA7zfOn37i/5617cDQHZ9e7ixYmqwLs
Oi4h2H0tI/XQkjvZC9jPnSDJZd3Ok01DOQHlHFh6HzlcZLuVyeOMp54lTZtR
1cr09GeiQBmbTt0h20cnr7CCFas9AauLbVSYg8hmBSh5x0xf8CiUdg60u/oo
0LsXMSbgh3T+Lyrhd8Pa9kcs9ZPwo5YC3Ab70rTh8BEXH5MCDCOn54h9w1rV
0Jdz/a3knKWyeEk5uSRUXjEReRS1BImIlRDYw4w5MYocGT+Xfw1+qpWuvO1Q
Q35kcacvkVXsVLYk3Pdx5UGprU6hSQQcZsjMTU+8dCvKygj78EnY45zJ67oN
V3WWlq6wwX28XyjE/mE5lTU6qwxCA/YKA6Aa15dVW/t3EcVnx0I5wUjggOnk
B7+3XuI0kr68DxAthY2M0ICq+FtcqdflAQkAX67dUybZ8piyT4JA6hDiNoLO
Dl2eNlB/uBlvL0txVRPRsVvl3kcUg7V8GFacbV+ddjxCS4rgcAlC2oA30Vks
gN2yiWZxPSzFlGMMoZJ374a6mlZjyN5JaFDJ9q+pTMXQaXM4j7m3saNA4SP8
SBC7cTOjKRZzUfM0szbS0bA6V+bKqDhbzkbGFwgIGfvMTaSA2ojSvc5WyU0T
IG3+S0oT3kUD+awvUZSgVxE5gnoqIxK1Ld/8lSfFoPoO0o1+dejAPDRnbJ9/
smo3GS8fpShDfWs7TWS3TmjX5pfZ6k+Bq2QxOa5PZXq2PSWPaBcNc46Bgv66
Z6FeWjXyBk1hbqWVvgG/5PPdPbnHwtwyPFu7X2qbQHi7gQqH+LGkS/8++tn1
EWXmWWnLa6ISIQJPhMS0qAY339rXq0HhabPziXzLuc66V5ZCkIno/VFdSxPB
H45lo+h4PJ2OWu4vpS5hZk5hX4kqfqRc32XAIN7nXz4CWjtT3eoCfR9eaYeV
w2qPamxqzt9e3HKH0gaD9IV+AwkRPQezmo4Z2hpToYpQgry7ggN+oxjhF+ns
1VSHU+YEMcxmcAbotlOahGxCgJ1oVv12FqBFsRjnHirork1oFg2Ir2Cw78Bt
1UaxAPODRAMbAu0U6ngSuQOJqu9SEjKrf9V5MQOLGYWEDRRkxXNqZRE8SVVj
2rci0mw2GzDPcK/ooCk0NHXp24Jj0ypXgOD1fq9VLSTx497/Dqbc7tchz8Mk
lujdj+StDv/NFQapFOIHwYY/ceA8KI60ddHFuFydIpL2fcqQeOTtfJDUkyLv
4pO5EeM0SYtqYQIQfP9UMlzn4ciKdOmXC94MtQsu7zCZCqkoooYktCS3a2/w
/hmhvPQBXXDvt7CsdzFnnQ7QpSTqog7tbFNoq6X/rRCE3D1kJOatwD1+MrH5
0/tvSU6zQj3+aewvqjjyrLvAsO/ypD7jU+cuKAQCSQYLkmMut9nKcHiUd0E2
M1UhCGzwNxK27LdgG8+pWehfTw1eoVxS3pedG2oy82Vp0JZGv36b1acbpNgr
eeLWMJeqCMElkvUrUC9Fx5uHWVryaiqY+BSePTpgu9wtDMWx5zg+SQUmUw9H
e3ieY7KM2r7zLW9zuFQFKmzj0t+dJzk2TELXo+nh9Zso04IV77DbG8SR7IZO
SXcR1um9Ztfqw32umVEpoY4V4ydNfgnu1qD8NGnuN4pdOCagwSyzlh8RvWpP
0k7ktQhW4CwtfpfB/+eyTddAqiOuNYrJCzf1pIiUiRyEPYnoYGdXu1nU3xKW
MFNuHAUvMkDPgbJ7BuwJp7Qgg7sCryolS/07gDCKGO8A85jDR+MJSxfWDsal
GXPP2jWh7GY4aWKr5rk5uppJtoeiDenpsaqntlaMHKUzILoEpML/uGM52MXX
NM2eOCKePXmq1f+2oP9RFNpby+2KBheb/RHwCspJhaitDmXgcX6lt+65zQU9
54VsoXcoq22oPhi2M3oMcrL0pgsxOP9ny5FVqT0LrMemLhjyH2ZNt1GIV4Gs
enhnFnyfA7zpe+1zwDW3W1QxVl/55Nv8v61wsaCVx9dVqESQP2MHhy+riZL6
Q6cUKqcNTt6KQAZk1qIivzBAaC+QJ2b4NqsVyD3lYO99Cruz8kW5yqz0c9hw
2pCfqmM1odR3woiPJB4+tU5j06wCmAeRbQLRfreCYYsH4HKtnvzxxLjTvUK+
IpAoi4jRZawHJp53JxKA7/38OLhU1qPBCQiVh+4n3FcKEruwUfz+oEherY9F
h9kyhKQItMBOE08xfdoazj0BfQPXgWbLg4Icg+RplM97ikn+iLTqYNdf4GIQ
a2ZQa7WbgquaxRefhJ5MVXWrasEqsN1Ed2MIuAVPQLz6Wuf2ml6apUU6jo7j
JMYxUszDZg51CP4qBnmhbjCIX8gvusIHGgI0tko5rqaooJEcYRzM7tdh83YH
1FMoVzKHiN30UaZpW/yOu1dXINLDligWJTgFX5sR1v8zlFKQf9KKBE9rqTSL
wS5cRTdn84qk9yj97JIgEof6SV25ytpr8r08xgNozLb9mF+D9mWLySLSCXqP
7BOQozHf4r2J8bQcjydMaAaLETUFAFtA6L/+eEXrDnKd1IXLJHnH98UNA/fC
WcSM82pyp9XhyFE7qezQRKmWuGHbMNO2JJy942qT4QIuwuU5zwlxUleTkMx7
VXpiRCR7Lh1CgCjclSbfNnsQjcIX/rxKAdF3eSxJoyKRigWOHhxm+VsOq09S
mPJO+ltSN4ZPRNqY58MZ5TJqUEtG+yLUdm8DpTHLiG7qMkzkRTR7oe6kF7j6
GBpYKz4yXAxZN2cxWsyu5Q8Vu7oMc0pZXGW9cXvlb8ZiKEgc/HurQzb+RoZ/
sBVu+rVi+DT8KWc9/4i/yfLIxCPnhnXvHJUrXjPo068aL0Whl7HcL4tTnCfm
EuPHfcU/fo1cWDedp2GbkVxC/BRp+QL8MCaWnmG0EIKPUWqkZ+aLk4vvcu7S
9l4hSKXZQ/bgqmzlIxBWU2BjsqnKUyOhM2lM4aPT4zZN8ZwNXZEU5zCm7DWy
djUgwIn+9ICfEHbTsTENu7iSIcnltw0iojCq3Xg/JLSJd82t9RV9+2gqCnGa
vfM9HUGyFWwrM+CsyNsAJWozvQ9y9skvRJCaWDOwpw2u5Ok5C1Yt4ENAndgL
72gDbEFVCLghRWNG2m8goO9CokkCXzvH0UQOllJ8fnSMvrjYrFfmfwTUfLh8
Yv71LQDtqDi5+Y6jxSpOnR13qlJ38BQSD9TpmVUJlZebA3NUbfm889wEJNxo
b8o/lj8e8WhHZGHtsIpsTqUc44qx5G9o386auzamECgg/uN0GPPM4iqyScBr
OFOzuOK89q73nd0JmdtFV6pB4fZ/T6p1K+j/t7P7gxSPOWLWHrVL6qmc9FPl
fiZuwEoS6JQKcL20f9eTkuik80I3fOLsgHmePVrqC2qkWBt7SOv3j0rIXIJg
H1/anj8tWgPR8K2eCGiE1emC5nTcG8KUT0hWz+kWe9j0+4zpgQsD4e+wjeSi
9/oOx1xv5vBKXT4u6HzU3NTnGaxoTn/amWBq0XiA/dcId4cm92iOuqTz4bWq
eYGP7RCEHypb0kNAidE/QU1EZJoSqLXLKohjWHCWVEizuoHJXMyxNI2K3Jit
5tiN/sNxJY8yBbWssRK4ctwqxakhHquImze/Gg4PnhLy/tAwL/zTzBZLxBMy
gAV1K0c+OWY11pXGsRQcDFD9Fwpp8frXZ1602rRmfTv8s3uP1gF+9Wwbh/Gi
YrIlt94MfuFgxcJAFSQjJH4Ov+H2sHWkkQbeI0evIYPHjCYVPmw1H+guRLoX
VVGSMfr2R7eyPllJXkmWsmf8OW6YXUVJvs6f1dW5m9U3giv6j/gGFKO0R7b5
Sb/elwjlMbmhCdsvz2ibWKu2TdzKU790+9tzIgOHxMWPBgeSlFGgpeXOz8vf
JEcisP4YGday/xMhUqInFdjXMba0Ilt8H5UXNDui/90DT4ezDXDs/zsSDnyB
SYZDL33RId4HA5bX66GtlFRm8NXhn6NQe9424VD67Vpf18zluK/uHLaIfsSj
fc2HxB5LjrSuVF+ElNFrjwnExspRBIN8KF+Pb6rFyK92H8JDNNlB8Gs7mrM8
zGmla16/5iFKrycrRy2jVPzqtVU5GOSZo94/ePdEJmQGSeaRe0n88yJ+5g2c
FV3Fk0e4f1qM15Hfmg5i7jxbN69xom3CFfiPwPWSezbLTDh8p6nUOZruBhKX
6Cq8ZfXSE5Sr9TEKRPqVltDxEAjjIidbwmHo+ZfM64tdtTwv+5ucD2Biux7o
wksIadTN8yE04FQCfTtUgFKVI2K0/HOCEK+3le0Omt16T06oc7QD8AxIzVEg
oXmaiaMwQOLUatsivh6TUFGsx78YP2LyYGGEzy+br62LJ0CT2ydnmqKSIzMp
mmHXzAzrEYu2xh1tZKt/fMfEtIXaZLggf8Mks/3Ve4+fQlTR8CqTynrafEBY
xOtucXVLHfnp2+svcsnl/MGiV0tTikba3yFNp21Vf1Lla6RhLhRShPWSUVIq
1io+H3Djnjce3hWI1ozeMb6nHeNFVpmd4W0ryrcxH0QpHC4nNR+GbqX0TVmT
p0ez9eyYCvwEbcwAeoEbhDk+6LWWTFtP9fhBRdMNrcPnAPez+TWnuEHgoy6u
uq6yU6u5aEf+QsVGBBmYFf2KaTlFvt1K0BlUpVqk7lFp7XjNS4BUnrLehBBL
pq328yzEwv0quVFSJU5jkHTuugxZAQoIvsVxCggNtRF6Pfcp+V75bfDNKgCz
tAs0KesMR/V8jIrdKeE6lPxBZWRtMU6SoKPe4mL9r4sr0ry05h9A0ENsayba
9QJkGWBCH4pGfNIdLJFHE2A+QBN/OW7QoSjFDYE98Ck6vMY46HbipH1tC0iC
h6Pgwz/gHiXCfnG/jrnlgmjyzO48SKYOyhoYdjDczCF8DVlDmM1oBLeB2FoT
LQjrN3AC0W1G+es80PIEzjZVVS/3XOavVogG3ODAaU7qXeYb3fY3j5j3doJs
7RH/97wqjR7xWqgnmFkAQqxfYa0/po5hTMsrQsP1BXiUwYCe3oI+rCBHvgpz
pQRQwFmIuFFR+Dnq8iZhxxHARzBsjeYTukqIo4fLF2qe2p5M7lSXgnvPU2Jk
hfIfHdNqNkPejh1DOo7sY0bdByKDCj5a+iUdsJHv+mr7jO7IOX2FsrCyKv/F
IbEOLEfcywDtVvYnXG4HjVnZYEoSpKLdHY/heEHR5LsUR69chv6PImN4qe/t
v042iXPwSjarA7OxTfuHHIICCbXBf0Vfl0HIBYvitppWhs8XGro6HyUdzT03
vC9fbI7L7ZupFZtPJ1+inWDXOnIun08gHi1fHuAHmJuZyDUKNiclmydC4KzI
MgI5w6lsn2vp6rJoYjRxBPkF9qY7LqbFP6G1eYl9nrEe6aDGGSYN0YMNYI+C
ROy486Wx57xffbMOVnGkuSpch5qmQmMAzoW5zowkWH8iOOAsgI+7o15zhwK2
xIan4iXKYsGt/KTpaBsIP0CCH+MIMFLng7xvhD+gtF51yS3peN0KSE3wWZYS
PlExLgaVSg/h0kJfATDw1JZSsA6K3Xk1XstfU9IQ3iIfRLFYx9fPnL400/cl
/j9NpQ1h39vnT8VaiZXSqdTl5rkSD0k32tXUxB1a8nL8TwsVCwPDRqwtMcaV
a0SIh+pM7z02AaHQWoCMxkcxZJUzZT79fCjsgfarR8ybWrPaqHEKYc1SGD8r
HQCMw7ZBZO8Yeiyvbd9eOX8rnnKD2mi8jzN/W8rMwihsuiltixzGmwSXuaaN
rf0FlzOf5n99aomlKs/0/Jsu6BctYL2NlkzE4IjoSNMiHI3RQEYht94GP3zK
7Er9+gkQA1HwtPd7FzxE+AhNy/vtxNNpfW5fEGmZEbxbwvjxmRWpQS6uEhZD
nffFYA3Py42NwrDSTbqHGdQSAp9jnN3nyOUqOvyzZMXVl4vI897Cs6IA4bWa
MA/30TVxwECxiW0mJvqNWnPpAYmnAo9xLPziv6RayWhn804cxw1sWE6gqZqH
BJ01ZY+cjPuuxn9D/Vvc8T/aT+2U3c/u/oNedLT3K5iVSkqZy08W32Ni9uX5
EonN6uea7QgtDb2/aPweVXfbdwNX4gNHNTb9Z0SvFiKiFU4iwbfmEP/XLZGn
GsB/N8Q9qPF855E5IYT5agg3cUJvXANUHg9KtN8LZeKxhgR0jLGydqtF2IjH
VT0cBmHKtE1XicUb70F2sWAp047E6Hfh4PGpT89tLsOeHpMp5RaB2bXzewDa
BlX1TjJ77rQgg5FYEZV6AofQK4lI1xeN4py1jOS9DUMsJIx/pV62b/flBCdO
YZLqeU9uMBPtKdhaU5XVdaNf/SDTOF8W8Gr17Ppi9r2Bry354qJ9BuXeF4SK
RRjvt6/GWsGt0dlESYNxVrjeqpbR6ywQBpexWYUaYk0IWxDMbVYkdUEbE2+x
PuBydkQb52Gsrm+gHHhQciCJfblVjdEeYHhGZkxo/AYo3eDqwR+XSsgs9Pn+
tmWlvLS/uTdxRjB0ujdLrZFcdXQlgZE1ZpQMn44HcPGFghEFuxPeGSy/LmRv
+O1Sfja297298BBIo2GVywFL778ytdBkhOKyQulbsIctU4u48dH/M/Y8TYgG
DZkqYeLpt7FbwnhghGlTKGJBq+q3DtqnHXMuungChJartbGyvvU2gJYhyefw
1K/u4TNbKEgB0JAe6kRJbDpgR28aySlPaPp3XUDKB9ilhkEGlvo8gFMoaTlA
cF/PEYI7l0F8jtHPIPk9HKCxpRpGfaLRrSOL6/keg6c0eehxBoSHhiyDMYtK
Uwx46BCwjjd4ANVewR2A1okD2Cjw/DbJSl2fISs1eYzXjRxa93D/Q2FoHFH+
Nu+IYp/UMiQ2tjYj9rZAZ20wq0brVccRVUskxhsbI6QF7U0Trg+o6jzR+Jg5
2sQPXR31ESEitOZ4lUEZK+hxKEmuuNKx9RiQbw9kGZavBrYxoqC3UU1G/wL5
Ah3gD49ohdh6z+OEuqFNF8MpC6c+J0vjgO5gyay7FmcAog7buWmZoXUzaatY
GxbTi+fQSHkeBimT0qU8w1uIHYS0EV/4gv+Bx+QxxeokUkBb+k0gIyGMnPhq
f9iBT7V+Xq5XZKLwr12SFn8kZkTb7O3Yx9b0BS95a/D0X7M5pZ6jjN9opZFy
5C0rcXT20hR44EJgZIcUuW8nQMl83q9VihZv1Oi/QWBegQDYUFRdJNuQCHFC
nddxsycXvevKCXbdLEaQr4Ofo1d+bLp88L0ris/cd+n/RWhVmvJR9dOw/l/7
m85VQj26nJFxZ2tKtO97tfAi8KUxg3PgLXS2+a6QpDDJSKw/ewGELjuu1qGi
P5yn127ZTzkuu2LawqjIi0IMj5ms6tbqa4wMFEcnuqCSJySQaX8abE4JumWD
aTSr6ZFDyMLoM0yCy4iWh5PBfEGgp/Pim67+j4DPSRERTG9qkzj52YtwQvcz
F9D2iLo8Wdb4ulsxQIdEzPB/PMOjrb9vRPKJ7HD6NgqBNNmHK6xXw7jsrsCx
otzZxt+Ifv2ZDyWKQl8RDaXbeTOSMTgCslhZBXU3upIs1wsV/jxwscFYZg4I
Ra+EttqbHSSJGubtZaJd1qERM+GyYRq+iwdgn5zPAoT3vCisM35hLmzs5FnO
Bu2ML+y9YQeiDudPKH78XwAgZcqME1+AscxZe5mRGvZIfMmpvIlwokqFAHPZ
+QRLIrgv7MCWaWTl7CwsdzBvjn1l94qS7L7nXNws4YZbzAMGxJqCLllscWTM
1rDBtYdWogp213b7GFw383xrrpCfYytvayJp7LNahnMzDC7Zzz2J8m+Jx9nc
0+H3XcTBK1b0QRo3og2G8qzqnGOF8Hmh3voJF+tdCKb7IjQSPXuvjuuJ44ul
b1DFt8igKZHk5WY9ZemUVjo5T9H/BUK0QwPwSaNIACQNaeMlT8Byheao1Ei3
HUE4yaUoSCIKzTXv00zkvx+Ea1An8VJZ3hpBN2Nbl2vzLJs56UHTEZ9yb6Pi
r/RRPgA7/LU2De6hNQ0Anm3CAVPvJWOC4GYtLld9OskBV5dYdiGyIeZuO93P
uZ0S6WhgHSxWK7oxH+8tjPgmPiZZ978sytuJGcm8LEDM9RF/G+Z2Qjvkzn9r
lYtrX18DuytFStx+fecAXkFPyLE9BO/RuotZ8h7ANFj3GeT01lDRtKskbqnq
FQxBgtHM3Xv7HC9Kkt/bTVwyTfzJPNT8CKZDkKl1YofbCtzzELKwd4nWy7qm
7N+KJMzA7P2MKyqNFun68AyAIIbtuyuPG4cg2zL4QlibteWULTmiQiLlyuxS
wX9Q/pjEiDCClt0Zn8QPdQIValHBTmRNxGTDlt1Io89wynWxAWMkviqCJ0GW
zEugb+PXAO42vmp1quAAJXJyFMC6shnPB10i8Nv1PFITtICCBhsZOtyNjBmw
PYR4VAOkPZe4D6y7+sIvDikQvLn4UDeyyo516K/HFwI2nClNN7jSgnLznKU2
kYf7K+708iSNMouE1qCB+yFLjwSoUZ7JuGDLkrJMu0BSfPBWX34qMKIWhqlA
860VlG7131vHdagZG6T24AojEHFnUv8p+jl/LDKxHHcOsdah1ItBuGJEXNcN
hOoz9ZgC7c8g5ZgZfnjWHZhN5Jd1iJSgrM0gCKi2E+wjAFyJyUyq9QyaJpDS
/+9pk02QmKX4EmJ+VYm19aJOA9288I4yi5Vep4BuJDPIqTtQwZ/6V32gr3SI
iBog/ur9nKZknsMHyVFIcB9Kldzao+nMQadqtxTUco8W4PjzV5MNcO459uK2
TzLnzFfQhon9mZ8P55QBtvN7s4RgcGbuewRrgY38tN7XRYQT9dlW42svpogR
/5n9BUmRRr1jVZ4+cTuL2xlWgSG4AAhEMwiLYRz1zAjAzhBEURV9l4LxuDWM
9it63RyHvinF2cnVgewY127zsRMwia539MYqMThhyTjxtGW7gxG5ZGqENwC1
7rSDHylv8gfGHomq4RSrvJaa+R3JIekjGvCGkTIhnEy/UzDA86cw8qrjfcH3
4BoHU5hhUTrjOuCUWq3CJOs2UT1XU0qf0I/i2VV4Fk241UB5l8lJokCWkAJ0
BZ9NKK7MPB/qHhn8uPcgT+Mt+jVxVD2iskEnqGPyGDEFdUldM+HW3EQg35S4
UCxnsI6SY6FW1BWuhbswthzBxby7b3lbRh6/8Pj9QKPNhxRegvuagxkcxlie
k8QJ9uOWY4Jy/K1ZuCXn1oApAn5VEanWuIMynup9j49JDIDUbKVQ+O2zHcT/
i/KL/XNsfbwg+hy8gSuOrjA5drXRzINqnRuSUCuXteH3la8Xzk8QgJVdqQjq
pgRenjg1YRntRk+Sul76xtWolDkwWSSYeDuBKNKJ1iqt95+0kWKcfbxsnFkQ
Qjc1Jxt1RXe7R8MU56RG9jmFM+wX3Wa/6LVJIerdzcgeu/MF1YEvOH+/akKw
YrQHqKZqkvIDu1MqpugaGOYjUUJa6Q7fvNDUoH7nvS9DRsF1p4i87pNj3OUA
9Tg8FPTMayAYYtr+uFilV+MWv43T94oLbDxQrUbY0th0ZeqXNRWDOoFSeWnF
wPopq7SkXtA++N3JMaIQmdcpZOOcrtQU6h2pDTGp1Nvm1G5wsUGt3l/eB09r
/K9dpkeIlTrpbjxbyV1ahPOw2n+052blvcKRRDKZ2GxlO6eJ+/gXrGP4VOI1
tHNHwNCIuLhiYAgf+ikMQLF7iddX6vaCAlfBVXqVd+xNbK4pd0TTL0LRTHkQ
uehuHzyHqfsFlQKBQqiErZEDzRaeCKG7mHcMiAVkbnt9eo9bMrHVsnyZndxY
JlZ/p+Z6Cx9PKPNRSMfkXVQnSkvmI9KEhCnZV0Bd6nbr+BMddibr3Zc710d9
xB6QntYyjWpmNEIpB+q9MMYwNw51aWVVJJg+IxvoZOlK1P3cmq6zcjU+GyNl
uZhEsgUt4NZyzPydybQPig+PvExf6jCgxdBSoinMuL55phEJEFUoZ++TGkMe
XBBnm6ADPKn6JcQhX+XdY/9g83C+WJh/p/D9QdifN+BoA4g9rhoTRHPmB10G
hVaCc9ujMRohmyYfQ6McRy48o3UZivK1EVe5DZkO0l83lRQRELl/XEdKO4Sv
aFXhShbRIxjspb0jDf6rKEXDLUDacrdkmOwVBizhAWyVfrdMI8LsJpCxSkiw
prPD8n9AVed6X1RvT+WoZMZxdDZ/90l0pOfYR59qTgTRyHnfj7+mq66AtoPk
Yt2w8zhYc2CBTnCm0XvyB7ib3e+CUty/Ajl5VTfXg9mQQC++wWOnS/lV6ydS
m33IPMRkP3Y2a8kSax/mnOwclwGBIzJFAqPVqnndtXXj/nvLqsVMH5z6J8Fn
pRr8cVMTdIzRxnpE1JfoP9gtLquib6AzoJ9PxGZEBfYa0Pn0OvxGeEdo9PUs
nD1dfGOG0UBlYPIld7h59whEs+NaXcQMIgc4zGRI8BuAnD6qlgCSxwrFxwtK
BRkKRYFIUd7+7V+WhpfS7gjwPmvuTdftvSU9NCEbYgIrYQ9Syw1ghJUON03B
zUbCualcPqwr6Dt5BB78L77TaZMbpkimjx7ga6JeRidjYHKO0D5zrl2pw1kN
xf05EDh5MuRhRuJthT6ZUZkOkfsAxtn92Q6lk0XT4Lvx46z7KqMehZzoZPXD
/o7q2l6Gq+ivXGw0ZcT8nX0M6zvHNaVAFajhW1B0GAVXYLPH302D4I2NNv/t
qBYWBv3U3+3yt8ensu1334PNpxA+EqEguUhEz0lrNen71DZ35UK+wI1jeq4S
X8bVzjpvQuirc+gTYZ0ndojMXmVdtKqfIolkl2vwOFCM2IRhkJzAxlxckPvO
xiZG7efdjjOG/0OenV+LvEBl5ewgsoCdkyTMJmwIdzxiHIrBMbjFelPMxgfc
Vqp1Iovddhz0vmH7DRdbz9oSUH/Mth3XCU6WON3hehS5l5DQdvWAzjfUXbau
feh6sxiWj0eGcIVXwqYF2K2BYgF9VlUqgVZEy9y6K7gP35l54SV1msyn6lx9
YMtdlsev4ea+xMCgXCj8l3n4r/N863Ic2nxrNa6fyi8GMIuenTH47Y+LtPw9
GllftVf/ZaOb7n1iiiUoJYEu8g7QhuFyYUmugcRRQ3VJqErn1j0lUOB2J7YG
4Uz3Es9iC+hb2QsIhuHslQX8dS+rIZo8j6IvJ/K22ZAAYfGcN4RADY5egpUY
pRJSimbaMTWSfHDn28/JekqI6mLI+pnQ6Bxe55gVdsMzzCNnSIw69xifvGFi
eP5Tpjq4uESjiPav8Z+9vOchSI53lVeSJueUVz6YrteLSu/8QPFLabJZSHCN
Skrj/JnuJrugnHic5XQv6mx4NQUYxC1A6fU8KEuS2zPUwN16eT2wyf8j6QSI
3C7LPJR1AwT0/mWXzQg6PRW3lZNQ6lM98in2Ez653QZnr81GOjDZ9L0IhvTN
AG9nD3CoSQaSrQMoiKG4N9qSipUWg5HvCpHLxVoegUW5oV4GBy4//g3l/Xgc
/CZj8m/8wLLuuPNgY6252VCQQncmN28uPlN6/ZGqLKO5stS1iCzKba6rvF0L
GxItLBwePRKao1ToVHtKldqGCOTeV6KD0CenBPWr2oPxqnLvBDQSadJumQ78
xuBi8/GWq7Mbpx2NH8Wsptw23GKoBa9R94DaoVqPGyDYONGCIxxnRLLmrWBm
oltVM11DJaRTtJQWbRQLxFpH2muKvDaqXGpGxX/0Xv4uHu6dRp2c2rqrSKg4
gaMmMQADEhXGxWg8pBMLoHGs+0h2odiAa2ez8mogrrbqJ1alnNgFIbKjpEG/
xW3g6tv/QaV/pO38kPaFAaDEa/3GcBeWv8CQmX999AH/AbvOPgUnWsy7bY5f
iNz/gbRmfLEpdGvFgbyw+ggcsaAuisxF6zIMyDrJhLodWwI1t/YqbV6KHyOe
yZf2y284675aOL4I5ypu8hElLu6qUMcTH78BufygCqtieFWq+g3orMN4PgDi
wbNKddZ46a11fFLUoPe7gkeQn8zRX3Osjgcu6ZTFnAZTGyHfO91n/92uvdYm
jVuTILaCoxjMNrkzIxD97F76Svf5aNRxvjPbEEItj+makBWBJXbPwUqWjbwb
BMMEP1Xlwv20++6D7yco7NzmRmAMzfl6bQOWZAQqsIUHpMpQCapRHauNhaY8
PvRWGbzGRh5wloUVOJDYPdqL0ZVWHwje2cUBRVBieingp0drtkzGLx09MFOp
JhzuZ7Pjq3kKq9LdwdC8IVM18ewx5waunahbbmzzayir5k7hx7pywFPGkkuY
dGo2Ctlilwu2aA88Ba6zKhwOC4u2D4MgeUlCTub3MbD8w/88YUjClm3UQUip
Ec4mhUcxkxciFZ5D33GNhG8rCo8KLBgWHgCWSMZeAqPl48ecfaMJ1+mFlCV3
d1KPwsEN5iXJwg9Ow2Pvrvx5NdVTnx/HENJwxtYQF3fVdMfSP6RDe+S/sVpV
b9DeJglQCuhPt3yc28clmubiZGfKso1c+tptJjTQEghj4pY5T8/08Nu1VwkI
ta3zIi+958f3sjmZl3o0ri3Vr2isMIvA9yujybthglQwTUf8/gByPB6WOfDv
dFMeS0SSbQUAVZEHimo5O5dv/BjoOj4au2d1gMqwzsE7Yxewq2AjR0y/HwKt
y5CjJHFVhqsWYgXRTrcOAmbtu0O7t3BYwGBDMUeIcQvgZAG5n6toFfpMYxFj
uGVz0oxLSayU54nhlDm5Amw+FDIDeBOtr9Y6wkmuTv5Kz1JQaeLEVv/vO6bo
kaLyCzy44rEzIlK/fOAGoTQNLzCkUQMsNV9BsqFQOuIgpQLKfY/cdpsnSoLN
p9t6ci7VoAeSBfiuDWTfdq21Y13n/4wlLHoa8nP0/3JBrcjBpOG6912PBZhi
oNzXIdWqETSvaBhvw7KZd+xpBW12I9orbZh+aVK6EQ7+eTG2T2qqZ0zmn4Fp
tCmY/+Wtd7loqp9DYCIrpUr4CabH9H1Ufwg2n5Z1JXuS/1PFFXTMV9hqYjMG
uDiOijE1WdiEp4DAjotxzQVAP3Xm6PtQZ1F3p8q5fdypwao04E60DpTdK+6Y
cXiKe0jM4KO7q+MQrMm+kLho7AXE3cFnmpRY7jiCD0mKaabbIXzDm6B9uZlJ
chUg69PspEz7v9BN4cWRIFBhEEc3XjjLPsG7Kft2iZzElKLyDlY91alW1w9i
gO3N+udJ4giiL9vYNeNU26GAx2glNnMvqVvWFdq/yzGbrrf0tCMJSuLyP8X2
Gh2hr36rMm35X75y0TlHLYg+vgb7kQ7vtG8Sc6ILRpKzyienMV24VZ7tmQvl
ZYOBKrJ+3v1NdIaDWx0n5f/T7niHfkrs/Gq9qRMBg8PZM79iDO9V3gM8603C
YuTsirM+PcvWGtGWmGiKnaC6MgCGirYG10PzvgbMVrKWskFRi35lT3mD8J4W
9G5Kc5/44DLnVOytyl9JxplllysSX7h5OBieD5ww/54bPjHuO3b0cGYIVJ4D
OR0ZX/VhCzXYkGhOfVFGj5WKFB53rBgskzmXSE64417qAmp2j/xb2d81KMQE
rs9VqNHa7DntLlsi+uo3plSiq01H1JYqk9xRrfUKSGOomt7l8T3KjNH7ZIQS
Wfbsym2ANs4x1pepK/XbQ9Pm/PDL/iaDh94MJQE2eT+RsR2cA80VcNGChzU2
3uVcnJrH5m6Ki7+Nj30wCQxX+flNJdevbiCiCcZi8SVLa6j2pYt8TdscDNn0
urzqTDf89QrxMMgKLuv4vzwzkUAW1T9pd5hHMI1p1FW0APZIy4/rUpNyrxZ6
pqCkWyVDiH0kiKNlFpKJ30wmgqSCwapwR8t9Z/C54U9ftf3aUGFKWxYXPuAz
43l7PT+dKYsfyxK+4ziP1AaiaphmhQM9U2w2ogP5tHxKC0YEwL6wIM5k/mez
1i7mwv0JNB4khPcNvlwWTzMoG3DjpYsSYA+csEcE2zP9chtliSeOZcFXqeZt
5Smjm0NaUKXUSpnJVg3GjJrN9v+wyIfDKOCI68ZI/IyHy8GdcYV2hgW8Ng+C
HSExmXxyLXysl3FGqzR588DSairHKn0cJ1Vxw2nAOjc2e4X0nn+964aAVR4r
tO9wDZPWg9F9x34suKourlFxFvpYiQzgLSJ/woPAmq/A3yXNpZHbOz0TkxYI
xxqeT+mYQyJ7ZzuWaiRB3k+eWHF3OIvc1FrldIGeRue9TFOeFyIT1F65mtdf
ODjRJrRPnzxCl4+B/JtvhbLz7m8iX8KhdiDr2YJobWtp8smN5UdCFOyA89UR
R9RcLQD+uN3qYDebvHBFmTLTYmZQ37MXzS41DMzDdMMv0JvBfoVMmNIex5/y
GMeAMyyapH9lgpDtO+hUp4wofr/gIgqYpcOvDguQG5iOAKeFtIyzq+Jtt6hc
uZEkz7lDrjeTpcc58Ttqpl7gahHRNMeQ+sWv13rjWEGyHPtaDdYDcepeV+zw
NyeUlWidw1s8e/BTc8qgVmttWSipcj4G1UWIZyqWJ6hQ2DqtFRg0wr8O0cv+
um7gMqZFYOeijGbmFqioZN1tZ+1IdjPO+iyqCIkKCgDGBWsVw03t2HofP6fm
3Hj6HhsLhkzIdeaOxMm1NXWGsMTdzkgnca4QKpUaz0L+ppmToDeBEOg2AdU/
ZdHJFhyUvALVR9vBJDIGEmH+WFTO7Bx9ETn4UHzvxdI2yfxMF0JZVfH7vA+V
a3k09DJ68xLIYE47/gnsW5hg9KZMQK+BoRZF3YPnN0v8o1vmkQeyM8btw0KO
vy3zIjbiP+64qKk4zXnI5i6ffs/7pzVh1oW1gzo1kWOO6v+Ln3ZuDNKja5vZ
GNnBYW5gisxvGUI9ujMNEOLPMncvs9KnLyKKiIihhu/7vhb42O1ii40N4i3A
54sY7gHmuyLLo2t+/5AQGj6Xmc4wjzTMVitAuhuAZUHh0S5QuBCJpHFUdDVz
9Aw/T0xOI/WjCTn8phrww5/JTWdYb5HPX3YVDoxNZvRA1LV2cMgy/Q3bVLlb
ye+VdbD3fsTqWAYvssCkqegyDa5nmYxzmzOjFsHCmbLp+vH9lMalhqBUzn8d
ilGoC1nwNeSDwd467jhHrbWwNw/yz/0IPiyYt4mCKH8dbl3LHgDcA3yUFJ40
pCDRdLaQOu7hIwA/j399CDtYKnjmAYT6lLAGjVoY4yvCg5xvf1bjqwuHYLiX
/RNuvGdfcS/R8yzkR9LBU5LOr6fTccAdTrShe77ih2Wrh/jKWYXFvF9C4H0c
pwf2xziNXsYVGA3soDLSAYdZWk0k98oTZjYbKUBGaYbTtz+GLRyl3mpmfUP/
CmVDFS6SQ/bAAOgTQpf4tjWMKBPZUYyAbQrMZkV2spOcoVQFlW4ii+vPirEG
c6s3tTc0VOt/vVc9lhF7YNQIP9tl31roCsa4I8xt+IobmDyZvz/nZl2LxTBq
rE5PpGrMc25lxskdrd4+sM3C8I7MDBeFwMl6GqVTfy3iSy6/DkkXdkJN9otY
GjtHo1iqPq8UhuzRO83/xYht2R85bgVt3niVm8+/eq/arECcORab3muM/3W0
OGiiq0N1+hjgwFbPu97jQsz3zmEnG4xxTYhnBA6ZwTzQwKi/5s4d6Sc5WlKm
BPkyA1JUpEKpR9x/gTVKcWXHOvjaVD9TfuwE2hLvAeRjOXKW6TdEBPIEKLyg
Ylwpr1CgIn0v+HZuI2Nn388+YJ3l3KTWgcreOELG5L2Y8rI58HKdEFABvSrF
HAjT5urkDGpkSMQrf7nPAHgzT4RT1C11se2N1dY38PlvUaAN84kGNeoMa8Iy
Xwyi2p4J8sTMFABaFseyORzDfxvmvay2NE5tXajtHMgiMi4gt9MELIwuZg/P
YipYtKI6IwjSUBzJLf86LLQgwB+cLt+ww9VugeITIDxSi43PRxmIjZge3xWs
1jd23JaAIIs1ayjFscTOxhwHN+K6Dyg0cG9Yj64TrZMGz4F0p3l2Sm1VvLK6
tjr8NJlxuIyrlkhf/TS/o8Q9hk4TWWUYGtYfNiYypCKhp9sSU4NXBgPXfBq/
tnNRF3eYfB4JnUgmLtX3VDC4nAwrzm2uLNKV12f7pDFzrOjauTJzcHTtSiyL
u0tBwtMx8SX4MvZckOAF+lxywM3x0++1d0efF5nJEywZKy4CdYwFAm5OUi0U
fGk9anlB2HXTRwY9WDUTR2dT5Xmqsp5tHgOjlOTcKB4TneS/y4q4Qsc4OVwd
2SSSriVRtWehTKkJRFMi/op1+d/rRSVl9xdoG7ri07yuKSb3bb63a5D+Gfok
goAq8l23/Hhnxem+L5AKWERW1mi53YEDUPrhZgh21mDuSnS3JpDfZXBJWZkH
jaliG+r19SRTkX7NAoJ8pxgeoZ7SrQ0JwHIwW07xHOAdg64VimYZxobn5BTZ
BM4KKCfSJxLAmzqIbdC77aY4DSM8j0Uxi0Hw1jMiJB9aAFetJN9Rlm+aLXLh
DTRs0K4vXxhYmdvYuO8JlFAIMwRshRY0NCt97tfksOPIm1oQPppXTNKmh73s
bdXdv362NhaqTf4UG+Fen/kLOWEoVm4PIkxDjXq6sngGSbLbY/FwJD/YY4fT
9YYDax2Bpprhbw508uIKK+wNqsl01dhgf6k90oWUjLkyA7BuWhBqHtBdDBEJ
AKViLkxe5+yZADgpn61srR0dEw0SXaz40TkwZlnpgXg8MRVtPByxQXqs1APr
jBORhiAEZ0WlZZ5YP941DxcdKKoLcN1SKt+KRgl38NmJ7Pq/3ACnI0JBFt1w
W3hXWBc4u4Fy9ZYaOW0Yh3A/hKU7C75R+y59i9qw5ISRg0qa18K4/ZKzgo1F
/s+WfV0yJmTFFrA4xvv61Xlhx1Ia9g7tu8tInNDnPZKwHN+GSTxggJe84pHt
3Nyx71syKOo+zmyRlVjb/9fzUZP3QUXuzM/8d1YyupNSi9uw6Hhw3UfrgMMZ
XBCY/vScvf0gx++rjBV278h9JJNFEVWBSjcY/saALs48J2xrJiKBYM4nbHA6
asyJLwSqpl7BuDlH0IPCMNU7nKvjUcDvowl85ShL+lS3t5+VeUDI0tIBMXiO
2LGDFlJ1Ku6w8vr/1TYtSC0ty0IFag4MfLJFGvSbNeLghZpy9Zsq+D24Aznl
CfIkMeqaHjFl8XrH8MqZMKtpiqSoiw4XoVInIwP7zao3OdE3yt7H/nhICH3W
COs+d29MUkabHRVAICMGr5FCnXENGCVT7qoCeJVwpSdWXTmHxiJwHG/TwjWy
iWv0loN8zxjjUfbzrTReV1c05VsGkjJoz/V/WW+5INM/xq985nv8heOrYv3Z
tV4OmzzixM6Dj5fMSEp7DsIcg48rHE7IWNeQZWkjydkkzjYcKu0s4jGiksuZ
azy19QFUf2CGXHOgOqNr45fDNmJk92i3jz1YnPT9uPjWbtl/PYFxhBScMxDr
6NkmpjRjKGY3D27qXuyiPghRPNopiA83T/8El87FnuLFlcZ1uwNtNhBb8CfG
TkLZ0PO8FgxQQIugmQ/Mlesc9x//UgEdDKYxo4bKoquRehGOzzDTXmEFMwYO
cCpVlSyR/tMdij4LK/1kQdHEqOXYOPYbFuJhvrMgffS3gOHvI/ElvACo8HKD
SZOyi0cm8L9PVlGVdlHSlaAhYyJ/UxtasWEhWFWfA7q1mNS7cAeld9Zc1lOO
zN1Q7ydHThrkag9QBVvmBA1Gps0gBVtyBE7eWPdHzOPmfaC09iTjOecZGoHX
WQjjdoL6JfDDUuG6E77NI83LPOwkaABjTzIHljwIiY877RjPdHKDFFmQ7FTv
XA7lDLZxWjy9vFi5LaXdcImRiAct22LXZSGmA4Q0YLMkv093efDHz6rG5i7h
OFqbwhP26sMCmpjiA66Ij+B7XmZRaz4IEKrbIzJAQLZ/5IFv8DyqW/RCWtSh
nTjnaNPhPTilKaayNKhBj2KYzLWrlzcvCdDdGcJFlwJWlhmxpd7kJNKBPbyS
aghPgzN65/HC0ZUPJ/6lzBqwlUoEZwiEnTegJZpfnLDTrVuimg0BRACwBYMf
IcrSfRaQm/nwgf7vmn2ycVUykRcycnbz2OJqxD+NTnONP+Q5wsrdYd3motoo
mm8GpAlaanOu3rDo3biEZdkF6+V+rSwHtSjL2orlblKBFeINwrKpXu/2HFzQ
O12NmKYuGXcAePvvbtI7sS+Q73GEC5s8M35S6C0724ki/OBWYpjoKHjRvBeQ
mqvrIBVHE/VI8GGq9t4iGbF95IfV91Ioa8367DrP69DtAeeKiVi+eyeYAh4R
rDMSKzg4hepoK2Th37hpnFw0M+ISCBm2XeXjrhL+vtvu519fqk6j13ODPwRY
VedFsvTefU0BQeKlR1X/FdD2LgsU6Q/svqD/BGpe+GBFBn2JX+KSNWwDTqKY
FSzvHLC+dm4e6Nor9EzNd9YhNTbn2t2tQlrEEabTI9l1R7zw0QLDekIl1U/e
G8IDNvHpoou5ON3R943e0mgA/7I8yIozRGsnTTAjBAob4DjWJBZ1TLB3fTFy
eQHkC1f5w8diSJ1ib9jFdWu8RiaoAIfGt5YZy6XPD0KETzGd8S6uqUzgJ4a5
udBPEH79OHj3Zg5ZvZwH0e6aVkJIheNZzMRDzxSzWct+Y49YBpeTXE4Y2Gr6
XAWjgMxzI9ChNuerAee4rStllIzENLshXkWm08BT6QodJpUhN1wRWe03TR+w
XK7+rvooaM6WiFO9/7GB5P4ZF3p7FY2iQyXSoSuQtPko9yfrAKMtMlAmzLoi
Ww4XE9chHhq5hPJtNAvjRhxifS+b+xTfwxTLldW6WiiGBSrXBZYFpMIdmYyb
zx6SFv1L7SY7xVzDb7Srz8POOeLptkza0X8n4xBPebMffd8hzTLKVBFZfP+K
enk3EjswvXLYwWMlw0DweAgp+pYBj8vIrFived7Y2MmfNNY8O/xQcBmZeA+j
ocEx6W8tw+Wcv+eawSkAkmgsVuoSRhrIqyQwRMCG049N4vYvB4krj9ckNgch
lCY6VYRjNxHLw0bnm23OQ/7v4BPbyj83pRAVmNdH7fgxZM0ojQX4PBYCdM6Z
0AXxlFs3pAj976ohWCsgu7JNHyeTlRJg0Vae2iwbM4oEz/gCh4ll2kT4Yzrx
Tux4CfBIJ9XUyS0ZXJo/jqC8indQZc9olsd6D+oiMChC3ISSnL8Xw/LZX+IP
9kIlRtM5grF860xFKYjbyGrX10rIRdoN/E2/yeST+xMoGe1gkaiE3xl5kO5o
IbCqFgz4H474myMhDG3gU8h/r7mrVoUYt1RMDRBnJ6tbo4MaQfzaq/pyTZWK
Pph1f848Wotylbnk3cqSNcQO7ZfDB0lWelK1Yvg+P5ju3ztlu/cmdUSDG6nY
3HW1low9W67tjDiNVxCyvwbKI7RYkYJEhrs2ThCD4qXv6mfxJ1zvPLComh9r
VmAx0UNBummIthAePWNqGzwpmXSjeyoLaEumrcrMR6Db7hwXcSX0BbqPdrYj
Tky6kGvsEIBkOSCr8jcVsgaItOhWAGFOpMmkkMpfU5Rt9EmKg6sFNfCQsiRJ
oMv0QxK8gSCpSQg9+Krvtl+8W8QqCd2ON51zsFPE8Rc8oF1/kujaZ3pEdQ6p
oiCR4GSZYB1jIIV1SwwfCZ+eVtTYDNVzSDymAd/VWg6Os0WEdJJAMkFQzY6L
QtsfjfxNfXWPDUon6yIMA9fxUmaDZlm5bpJhBuV7Y09oOomJYuFPXz04R1mc
JJKnqEukxKZ9x4R5DAA2byV9JbWLGt643qeEv/2To4m5T2BJWUOdmqYrP3Zi
M0u48d4/xlXK/nNSNXpT1P5e3uCplqXs1Njtq2EzMTXCQg40PoZwGlAIQ0LQ
QTMvb7GqyBBYaW29MUX/KZDw9zCKbuTzqcZcmetTwyPkfhnO2gEFPsWwbF9R
90Ws4PDnSENKLZcHkQkIwyeq7ageR8vSuStRTMEBi66Ohw6qZZNFAyZjYZop
d/ngQ2SIf6OfdR9y/ZoQukuYSGeAcDJzGbLY8a82C0uqH8jgsjQBn25v7XZO
nMLt0PlQ7W/1TvlwB8euEA0BH6oOfHRzDZ8vknbYkuJsKTkPQLJpjl2MNCTV
rPyoNw9qkOlznPRW+JR5mzTMr+idinVVN4hRhSLkXTxk0L60XmfJV4OCA8xv
i6QxZ2VINDaVptF6uUzs1qoep17ADjAooDxHpufWcy7HKAQyWl1fB+bO84dH
2ZOTrZIVHiMI8PTTu6qxLy6qDo6gEw+VzdBgiG8tU607TF6n1ioGlIsfem4w
cfOxUl0MRWpDuencrgVC0jQ4THkyLkjtY9bqnMW43Z+19W3Z1N3dAekown1F
sYTTFrUNtkPV79MXITGQWmVL5dKEWBjSM+MafVnS+IhZZ3ap8W6qQ9cRgvUT
yzMreK856k8jWSTp5cynRCijKrasFpA5jrl3o2owz43oVg6L4fcFOXnuxo4R
/jkuhd/YHZX3qw3pqWV0pue6W+0mc6mFESq7bgM7cS/ldp8qynBUMwGxJw6S
rX04J4ef7JAJa7Gh1R39+9qatI4frkWmVcqQMjhZQAQbqHuNuMjcLJoTtAV0
8KMS7uNnChfq4acygTTRD2k3d9Y8bczaQMk/G2EIDsmlSdJUDrDxqeN1beNh
6WkmZ9G+qhqvJS14LSKPD92r6ZIRWM7oi42OACn6zjkdP4ScBLvIS3Bttu34
I/4CQ+C6gfECHz59X8Dwya1GWJsd1u21TkLLiQKt/uEMLRG3MvsDO2b9orjc
iaj46z3tC//OMCrif2I7SNgthaH5dPWdB5+KFLsnFE6GZm9eCoaXPeGAZfje
Z24G7n84XJDAJlsENKJ4LfbjRnThgLTDmf//JAM1RG+jI45j3fdm7w9WGbHY
I7MfbkIf7KUljMpLF/BiKro+SAlZ1V2YgXZ0QPAWDDzY2xuAweAIAf1sBvpe
Sqh1UfO81tJiUOgk0dGQPHsZ7lNMteFQvrv7lbxIxAH42kf0+Q4tY7tha4EX
Hz2rAPjbYLYg30ixMGraNeDBWW0khPkPABRAf04YN0BSu6axy8s+MBNWFf9k
MFBHtKqjSUmx1Bqo/AfvGxA4/JL3vArV0A4o6AruyhbkcWWbbnGswrbPiM3g
VYa7M1ejqfy5HCyB9Ucl4vcytJITI86Re2eei3d9UW25jhXHHRebOYgghEWK
JtFjWWyw6DvEKn1vfa2h3WNNV16d06Jt5Bq1H9kfUMk/K6ggxUBX05v17toz
6JYRMpEi+w+JYziJCPFp+XP9qNy2F+LJZN8vNhFw4+EfqQ8BAWkLZPz/QnrV
y6/MUR3p8xbgCwCV2nUdpFH+YxYK14/Yo+XJksWh108Y2ASGA3aLewHvQ6eA
8mKeSn7auTWCUQEQcyEBZghG9ZBRo0II1LxnPLQq0XrjHc+gj10LMYJvL+5S
xJl1o0cO2CFDvVnmkBcHRcd7+RBc2hZ94wzll+9F+p41YCC49CHYk5O1NqyF
bzDXhRGGhL4xkof+Y5fMUOCoe4GL224gXBlOc5x1/WLuE1qoXU0Q0DiZkFjg
iPL8Z3ZSYMS20q5vnnBCT/2h9nwn2AM9K7s3x/lfjp/vX4qdzJco+cBPQpP2
aOVo82lXKSth2k0e0lmj9Ez6M3J/TuhEvDxNxojRYJNY57Ax6MWs3IM3DbbD
NRIa/bOwL32UBt1tu1PnQO8OmlmoeN7GKNdc7vwqjWjFSVmHG2roWdS1hf5k
/BDRn7C1QPcj5YfXkf+2qieSHJ+nVcSx1KmM+DYsYUNGETxsys0A4B9YeaCB
fKmLxytuHiQ+qlUIMN4nFV5hzCAnbFR/VffUh0u2io/g0fNtV01HX4yaeLlw
y/BNMZCb9vOEAM78DnKHXevbJSZRTfJ+NeQTmB2NHHOs8dB1Pv5uCUdvOY1R
dTMadnTdAqBsaTRzsTxbMXRPNkL9C9Oy16ogLEw6BYHVbLVYAsS4ymrbF4A8
aFKzEFgSkAMXBqV093ICC3t4o6IJoZ5koJxZyWmaMqKA9TxF94o1v318rs60
gQF6q/NVCchAvxR95wXgKqzPFzFHrIzNy3rFyjqFB9vF35pwU8qDUW7NN/oz
cg36hrHdAFYPP2SuC1yoyHDzmy6wTFUaTZLNTmSV3SMMZxqvhRuyYyyDh3ki
xy7C5TmQHPfddc/QU7MdoXBQCLV13GhY1lDMubX07w5GVQ5BnRTKimUaarnN
uqxshVKSCDGWXWc5J/apVZkYSKe4195vBtoJfQs85ye9U3dR+VzTOpVyAU65
naJy/3Odbq+qEFl+ePzgmxdsoykWNu/HVNtrS+KT1g16FfPixVjoyH7EwE9V
+8domeUKAW5swBYTKhnYpb8+uoBHZvZblBJwdq5ibLXeXPz74J91x6tJuYej
U0w2w3aiDvvBmtpLxxRPGRPlP34dUZ0p6Dkg8SUxvohWxwP5O/AsicDOtEEL
oVetyjt9USukZC9K+crweXZP5/jlFSQSvKI/c0Dl2saHlAHwowcjHoPfmTTL
gpVeOVopBmTi8bEAC1M13JQRWPc1JrOKEonAdLEcx2yA9spG6SZ6FVI8ufbd
JWWKxUpYeD0OukalOK35jwzwtOIcZBR8x5ARgmc0pTQbBiUkP2ZCZpGgJV2D
wWlRnai6/wO3odz+Ewya8euEDuQLirfsnZH8YVrxSbtP/QT3gGOrLS4iUlB8
QdYtDdRgOTq7jMo1RWn0MJPwxxjy2zcIggNxbmE2n53AVdBjHng/Sbrko39G
wq6sBPBHmR/1owL1gc/+3+rUAiXdhefmfsa6L+VElUILV1DoCDQ0LRCda7kC
sd09v4JiTMQ1Uzuvy87d0nkpUPwnGZQsFi76sqKWD5bJiTS2kGosg/x25BI2
jr2fXyjieQwDCXk6iYQsa3ZhJuheihi1e+AxBVYa5O+19mskdrBO9OCsDBPx
Dfn7r/fJZ8BYs+5rz/6NqLiRogfBeZKYcPVClT7kSAOsOevlMfhQoVPTvI3E
DLnzofN7YEVToAYW0DdV067X6Ly+IE2cKttu10hX41YQCFouPU5+5Gb5pkJc
3t2uHjIr0xJ3NsR1X8YTlE/MHAPaqQhrIG6zFQDemWOHNbfaqOHZuFtF8Vus
cfCX8p94s0wGK4Cg5zmuSHsCz+yDPFXIbVVo6URpyUCddXsN1io6M2sP8OoS
LiIgiwlB3YJE4WN80SWowtsjglh5cu7tMOxghmvGzemZf83gjhIIst7L9uU+
q5LvhtbLpSskHM+tY527N647kX0TD7z2HpSOP3UWLiGZZH4MYXWjxI8AT72D
UnHDUrgRfvV35/VTOoAlNqSMjsCzyRnKCzHAoaB26jkQMiuAoN7tVt/3sjIn
2nUm/FYOP01oM9Hb9QnTtey0E9Ze1dG6JiEumCPiY8Qm7TKVr5qOf/JvMBnd
hXu/zjOAwb9BWOvuYKB2mh66Rr3Ic/S083bKQeE+jIsGB1YYsuzMSPAimBr3
pfhITvxHeEuFenRArqbYKovXV+YbHdI6puqFufuK7lMrH2kL6GVEE3Cjw10n
lbnIS406uS/uoDtBnP5U9Qm++PU3V0XebdJa3ypMbw9QN0sjPIlyeXQ1DOy3
AC+hTDnkT/wSJk89d/fUlAP3rW1tcum7pujFOHGn00so0EsFyNaHu1RV/Wn/
MbsYJGWyqj0F6PwEiAcw86lRgphU6XsaiwN2H42cpp66i5Vu+GsaHlqd/NYL
H25j5TQO1uYlfRn2Mr9m9VEMZ5LX23M+7KJMsawRaBYGZMd1EyUkbpGGXzyD
W+3IbafM2939brqbW+VPVE0ouYfnHYQ7G8W4Wq3Ye9HCRcDjRjlN/x2/L0U9
Em8PBrmwMXHTsoIWFFL93TPUuhBCjat7d31jPVpEi7X1wANEd/AJOvdRgHQu
NgzwqOf3Y7tErTjXgIuGGhL3EiFgcS0ToT4kV/POrxVFjNI1HvxoNErpBM9X
QmaetDSs+0+yO5vE9c9oJqDCBlM18W7l5gCkGKe17cOeVrdKLwJVSxw25Z5P
IDi196TTv3D2B9DyjaEMeoyFlZs5X+SZXyAlxVK1oOzboRtQ5AyaxhuXKE9O
QXzP4vDhHl/3SPcBr8y0pVleVNbBHTFiovMWWdXRJPgsmoUv9+IWXGbRT4WF
meGhOW1pcXxTREyOwS39X/7fDUBze6EACOaTLgI2Zninpl0co9ZpZOXJbu2G
Bo+G4wTJukiXlz6VTHvgeuMM7uGwkHatnmfhisXf8LOzId47vlbOiyv3WRaD
eygefuZi+0M1vuNYVdOtaMLVPyPoRVJpJsvFt7xd17+brSY+h0BNf0zBu8DR
TF4tKbepR5uYubY2Yq67cnMqRwFtN9kpwNo4aJejl9fDfBHM9KKaVezcSZiV
hSACFXg32iglhmTLCrbl7LL+YmAdcGyamP8y7ZrehAQFVLkzC03/3s/e85B+
hdVz1fy28TRaKu2Pkflbe9S08O2ar4sCmxlMKFKT0NmN3BA/EZfmrzNwflf+
ZLya5Im1mU27xbyNmdndr7H90Z8ync6Szj7KdA448EU4Tv+B5Gj5P6Ha7+nj
LPLBdVwv5ehkIn3fMGEi19joOhrhq+EHSddfxdmK8tjOE/pW+TzizQDs7jYy
+RoyRLuJ5erEjV+h6l9TlZ7S7JWLICRs92IvGzJu7f2GWdja0E1lZ6Ep5rvR
bo7AHwMSPAvNTktb5WGLtehPLLaP+nSTJY5kqjJtU5YqKENIwap2ec4ZEEP6
RwZLbG5ZY0mibJI8nIFU6IQmiUbBeKkKgps7fdYaXuEUz4ehfXjUKqaXadbd
fHUWdoUC59zRj748kquucds3cCnq6b4SMAszUAU1a1fAkb14eGro3R4S4XUw
TEEVrhtnNrK8iNQplLkkwIcRiEIcdh+daHdk3tZLShL/hx4Gcs4bAhdqvn8c
dw+buGg1t0sUogPly4jPOrDSN3uPvfsvuozdL4X5bzOtixlZav1ZVXuoZ7Xw
z9cQaNLyeuA81wqPbtdOP8M57B6WVRsvgbcpsdf62FiICfcSRYSeoQkQPSXA
rYENdcF2td/CdRLQ/ruKkHetzG5jmQclrEh5MbqGrlGEf/naMjFIKrH5pFkj
gONxAubix+BiyVMbV9L6DgwpfgliewtrvXffwV4VwkQOqT2i7pubDDygteGR
k6PztKEDk89WwPe5fl+diIVgkXuYX0F0UD7GI9bTF2VHp37yzGNwIho0D5YE
uXeSywQlRSvm/ubDXSX8HcfM3yYGLwL7FUZwuSNzn7GhST3NeF57/9FFA5Iz
NQ+lLDTD4Jd9BlglaZdroyt7Ub1zV4pfb3PHQRzTpWxD9ErD7+rs/kC6Rk6E
Q0IilwwB1tt/J4zjhesceiFB4ExVvvfstKBSS4s1bRNrbyEIbVJVsj2tDOt1
secdgbphFQ16HVZgYAxx19VSXqvpi5zPeAtMs8DIM0cvFyuo6OU2pl5kezbv
nFJJdKz0SO/AmXSaG3br8aAyFKeZ9caP/BMaogu79OIG8w4gSrzPECidMry3
kDaLBKzLey/v9+LlrmIcbPsAAgEUzqWsdxYejGjuiVeD4BDceqPGO5nX964D
RNQEppmLMXsDzYO9VD5dfywlUB8EeIu9ctOn1xkqpvIst78+Aa9knzmOMfuc
bkzK2GxLYt3CAjZbPnvTMiR5fYMwh8HQC49ZIzlJoBxXvqqsqFzu22CMMqH6
Wgp15rpyCDaSC1TqAmH6vcAeOSogmRZSak6C1/xgy3im58y23MrYKKgVRn7v
MkXXwR/H5SWzPLqsABjfjebzla7No9LsSwhJXWpNGuSjhQ5QD8t2XAw05ayU
4NJtu3Hf946HApJB4JsyQWRnhoedV9hgRU1OMdcDt11VQbkwBGzL3ivFgRwG
GsYAyfnwz/wDfS60BTMlpyicBvB1CjpIeeYR+04IaPvQU0uzdN/knZHnAJkh
wunB/NrhwcXZPyp5b9LuOgg3Nx8LQKx1fInK8J9CmAsnAeR+G0IjLn8atsq8
8juR3BVNL6awY8XikHuAj6jsMXH6Df8c4KVSExEmnA/+kDWWxqxQJ2JfZkjf
wKQbL5+mnklRdfVK6V9MriI7gWieC016OtWA2/YQGgmZGNgpqg4Q4qflFtB4
qTOan//EIb3giPSAnGFlhoobPf0WBHHdrNRRa67bfG3mL4MQScM1g4zSBi7i
xGCznhzMqg4k0kK4F6DQXlXRhHVsKhvQ0NbDsQFyBHYBOW1aaTUFhlOPkRYo
BXr+QzGDFa4RICe7/ay7/0E8eunwo8DyfdSV+1B5/dY/KZedSPCKYpFLTI+N
qXFbWFp8hiz5pm5OmIxfv6YkwHbThggH5sAWWJhJX00f62PKC6SVfJA3Tthx
uygLxBUkdPgOgoUkJ7KqUAoIrlwvPE0J6IDlM+VsO/g7M3XaGTgfgYfhBK+H
i1OzlGVIb3u92bHsePyAbuLzxRD5+TByFdkV6JWpr8qTWwq/MgfLcWxv+phA
ik30vfNeJBiZ3O3WuNStDJqZTC06+y/STWZY4OpyZNz8I5NiWdIPQobSCHUW
h57yF2zjLcW/XKzY9fmC4tXyTKO05j2YK0sF2gS3nIZrU3rpFkNTXHbTgICU
LMb+J/VqcKYrXsQQ2mc2dEhfkaoY6YQ0UB2OxFIZSI6nzA6J+TQoJ7D+Z/6O
kdae9Uwrg7WnkopsXlQGZuf5194wH3LQXubBCu/iElYpvV5aav/qkmW8StPa
21YcFkOqv8PZ0rV6VDi6aZtFnAunrqtg+B0L7KDCxox2OBGtrfbVnHujmc6q
je8QepujCU9I+13jnmO4BnGPlXvUooadwJU9urQLqAnxo2souAhWOP17jEL4
ZoCK3Tza/1Y9Hn2unJYgsOu7wf0HZJvHlU47Dz9JimAV+DnpAm1kGMNoP8zk
mVR73SoWcq5YjVsR74nkT7VocbaUVAbYSQVtBogefaI+IgfWmkLcTrkSTGsm
g0+0pwdVfFD7k6CrlCaDBP4E7VKGwgITHmuYVc55PyqBZNe0rf4HyHw6xgSW
50TBTpAveVs5HnXh9saNfBzqAkbaLIVPfaigCGh6OMGJotGqJYkFypXWXa0s
KDVfx/Z4QfO0svMqZxRglxlXtiFJNGYzBHGOnyoo96wZe86Kpsnqh8AbyoiC
iRL4AoKqN9TOiWv0oiX1SkS+lJRXreAO0QBwKa6Dcw4fh+Jml4wvbGBbTeZ6
1OvytvJDe7p/S2KOSkfvQPEqRuP9iHLMVYNX6hJkcvjPsIZICgfueNP2Ty3J
Wrh3zFuIH5itflAvFSI6QpXMWvI6RrVSNRyJrLFbKcx2TpACqwKTS6D4WV63
/S7mZzg4mnD5Qr93CqwDPJJWCQQwwEeDRglweU5a64kRpOjmOVwMzTaAdC8r
7X7ZxCT3AUDwH2RExqvxY++OEvTx63Qd9EMmKlTlb0y/ECHKCAEa4cG3xfhG
EI6LPu5rcp03LG4Juo6cTMQgVd3U1XqUKWBgqhbkXlNIlwwNe2TFSP+GOEpf
I2Zh5MlUAiCVfa9AEq4+dzr9h0U+fh9Z9uSmbgkStuyo1nl9rvQWdJ8EHtjO
hemySaa5jmt0p7N9OWqj6brKkf8MGhOyY27NoR/+GZk/DrgoSZogLiQ47p1I
8bPvt7xhZlxPkA75qkJEawMQlpJsFdwEfehrBcj2kmTLRk53JESadx7q4SQv
rvedFcLuRVrMurhY5HwjVS9ntwI4UEgU8O9YPDljs760OQlias7JHwBAWkdY
8S7YEOGHLKbM7kY057qeGaXkUN0rYi9MOGNOXDZsfujd0tNgTy2tU6munfKg
tR7eYUvg7gEazPMK7nnU7gVN7P801piFuFAM38JJ8GHVUTsRnIux5JwSSe2d
FXicJ0RQiQEKtpoo4ia+QWUl9Ifziq6wg6I+SSI584hDT+0QNwSZXhi6SnJk
/TWoTapjqxK0o1BBqep7Ef/3/0wfHnMXHnrNsZZuhLoFa88AR/SR+CXb/pLC
SVBnmcStI3ctllRSuWc+74XV3MVTWR/aBJyyvEfCcNKAqC12u8BTOY/Dd3rj
fOG64gFoKbC2gtRuvKXXESTqhLBA2uTL5BLXeiTwXeG3NT9yKiMF67wgCJMa
57djRHjJzAv/B6y+sAB+4ccw6/756ZzfZlU89uuuqHf/UPqbdkzI0T53TpsS
3mr0f1m//TBep8Yo9HJkHs/yovjBcFivaUkWFp8pY09Nhoiy4wN2srepaXLd
1JipYFYd/wgxW+R0V9CPEtqahr5116R52lgjvKdSsRXMRmeEnaA2G87d3PGa
I6akSOIutKX7PJ+yJgtJghWWxQZ6NhBVbOUgZFEPl59syd8muVZKxNk184FN
ZPGZfAlMpPMIBNqBXbESdbR4nL95dSHX53FOXFZcq0NJPt37JeCl49+ySAgv
cDURO3wF/7JcTIHgDTB3MPaJchj2vVPvlJh9FcI+O7pPpawBg8ILS1B5epfK
vrIGFcNomNTPos65lFor3ECBw71cQsXl9IRAYxBWh89xa4QD0RuCGuPJDVR5
7eV4hbrjnCRyWUODqIT6Xj+JRqCGO0iVwF99BhhfGLvJhyFS/MlrdAmHB2yy
WUd9+AABOZG058h17r8JCaEV787i0aPR5Wmeca4H5f+j1z1vDknGlLptCDj1
y1UEOeOthVFl1PofVo9tyy4fae1pR2Zvlbtcq7o5nTQIGydeS6dGBH2WbQTZ
77VL0CuXITX/7i8ZQOhCTj6o50sZtmBVauFTH9PhcfHR3h9N7KPUK8JxRvfU
ear/9nb5iVQ5XInEWe/D9ACZ96YvoiWdw7+u5hEVaHkXrDJWHLmfEK9G8Pgh
lvg10rI4mEvQ7q/RYIdSWtQ1ruwp3hfOc/u4fY7bNjxsIUjDYumDMlX0OdFm
4oJ+BRAs/KLt9EOMwKEYqzNHDt51OG7F2GJXGsFLtKbMvE6QhnmO/uE1d8Gg
47oO0FM0sRAay84HSveNmwO8TkQwn7DJximYG0CvM8Jusl/+v9SJ0RgSPRbs
rRSImPtPAzFJ/Rr7TMKueOYp3AnzXkD/n0qea/Gm7s03yZ+FVKM9XTPIl1xE
RjzHfJHqVEY/d13jGaJJU5F2IqJmY5cwg7DT5CU/CnjZdlSd4S9NU3nn24OK
h/h9ZIokn+xyE4wd08/fqeP5sXz7c9Bwr6+OVjItxZehgygY4GxxNM0IHwMx
KMBsK8mMyi3mg0t+YvBuQJyLF0S/B0qTJeUWJ5Db5jxrTYxNZPrEQ5VQB7Xb
L9hxlWIu/WBmXNxV+jSfnCrR7n7ncBoUFHg895U91WlHKIC3MrBqwZEFKKOC
GTumloGMfb7f07jcsrwxS5uc4HTgD7JYAVf4yC2RoPqtSub3eXGetvTyI73n
e9Fn76bGP4lIYvXUd7h908vb678qmEdtvNMIh66g/62RlSZd+U4GUqgMFw5x
dAOrdtzgL2zzT7+3oMh4LYH1vGhrH+g3yHprvZLBZ6ASenKAF6RuX4lyzsrt
wImXIBgsv7ve4+whoQ3B/kkw0PMAUYhW1DbzIHzA1c+h9OM4/EAD+4PRPRmQ
Kq6YTUOsbMicMz4Bxl7Ivcp3kLDUKtxfrotlCB5e5YX+mhYT6Y+dilB5dzyU
1lEbdmidkOvFZgufnJillP3lLGwzj2crIuqgFRWeSrUwHTSUhieV3XvGkiYE
C5TXbZdyMXoE/n2p9uqZ62vUmM+ab5Kivl3z6oFt1nLE7BrpNfP+CAhaxUaB
L2Hp1ens4lcyGwxEWKQgvn06Me7KGmGYdsAtSHcPU19KJ/iLEQ2tD+w/BmOy
ENnHJyjxVUpFT9gxQKcOcX6ONYa4/W6e8VaEHPbPpfMu7dTks2CjkihuhX4o
skb2TbhZc43UVcvQHbTcw3IgtR8jCldukKMqbiQoEy/zYFFbf9F0ST9u/1MF
UB9bJ0XDdRzi7ynQJ9Ne+VgOOlUvqzqrMtEwUrcWbHGmBtWYsuD9wOY0aU8j
5hPp5JE1tDbYc7nDxO0uLQbS+lxf7jF4om1FtT/2qiN/6uROd+hME8kN1/oY
XWPTJhJXSzHuK7zgF7qOvX2S5Cul9ngWXohDDBN3ZbPcUBvcQ3P3I+yG86Fb
sUwCFFrQPkXBFpGs1ksfZtJfRNjQyoNtEntnbnjSvkol+4sZ42VPk+C7IFot
iqrVPgvqcpUFELpH/eJj6sn69Dpl1Ljf7EU9IPBvtlbt4VJr0ZjJwpojBekR
cu2PNYX8yakEMjG+Nj3nrGniNRqwor/HtTpgA2nSZC4BoZN+NxyP7/6ZLnPZ
8tJdZ24HHIfUk4Hx9UhAL5GkEHpEFytyViOjsDcNz7PjlUArhfWp/ZQbmSub
BNeNxRRoWzF68zwMaVAq7SRWUJ/Nlwcz58KzYeBFx5QFBV8DqXMZcN+j7OcR
ozaBQxJZaX8gsiaYCYxDRxka8UPOxTF8TqPdONiQ3vOy0NV2A549t6ZQOaEA
RBtMPhFroBsnnuiHZxxl2/IkMvwyDojOGPTojqtheyNzGvJYKmtU+zcGCcrd
ENpYxLB+EHQKAmdh2C+8aOtDCI41o4/A+vqxyouHz2OAlv3naILLC7ypi9IE
d8H1BZWMkz7wAsP6BR2+zzieOUFH1CWJdiQCRx5wGZqzpRr+HAdHfWzIgEsq
jOcNXxYAppVx2EKQVaeNsBr3IpdqKx/brUvrMl1APddtlu0HSc3a80wCwy80
F36yxxUq6tWSU0HB9g09X+aPdPqq0RIrk1U3hGv+jg4H0cjD/yPzdgxuWE96
MrnR2AygrnazW2QajExaqt6z/woQKj9U+0W33Bi08q9/aVrULMEegnKlbTUv
8mLK43xE9v4T2Q8opmVgg0tgupCRkuo3zsVDRuGWFv7MndTq8ZJ31N0aG7mO
+CsOE0HNVVtTPW5F6rqEjK9ZqUhKWZfxIU60vECQYEcqGISiuLbIJy2n2ovD
wpaNuEMBZ7/ndeT4+867vDuVasP4T6neZVgHKso/F0CQTggwY2ufDjYEw3Z0
IRjCD1SynJCxMI4w+1yZ0K2oPEzMyWU64dSmQIMUb0Bo+ovBGKlWGiOXwfwt
0nR21D/7J2/59FL3bhB2+PXmG5aVwr9vd3p/cySxfPTghO8zzAVmSSvchJ+m
3nLTlCiQs9LnhzZMa2aDNeTf6UgGcsP6q3UOwmsbljRZ9ut/do5sgFB7oOuJ
vvacG7p8v/JOEP+T2qQXC92eerp2GMdI8pITlUUHcf/1TGX/AJN4DCUaUmIo
B9W0GS27UZefaKJh9PmKc2qdOFwTpd7M366PnBEGwN5hjFt0rLro7JOh7bkC
ZdG3BBHYu3ZaiNL1d1x8oAfxqPzq2yE/ur7vpgCBKFZHWHTBNRznRhzkRvkq
FSvokGnHD2jHZ1AyC1girQ57KR3E/oehdHWfHSYeLVPAid9QnhiZg2IrJUun
M0U7nRckpzGyrLKqTICOyz1JLv4E/384fbAhQQQo54A4xvafCyTjk3YP1nYv
UlfDHIchOGL+vf7c7g2YYPuxPQ1JlHrxEdGQ8Lmg+0kE7bQj51F/2gH8qKmv
wmdScX23qtU5gbtgtcjhCDgwU/xCkiZZloUF4USJXvLDWM2reTQggUKA6aP2
gUtpBdHuihJYn8n0AvJjo+eXfqocvTLsG/QyRXtmUa8TZK6jh6Abz5QuzFvC
okvagTXiWl7EnRuN0FG0I8ZWvY6nZ69qQ1UJDx9BdBcI/9XLPHw5oRdZYuKU
L6A/da979bpXO/yMJDIgNLXFYQSjrg4l0yDJ050MeREXkUv2Yz7ca3ulVi+t
I6XqiVeT+E1XCRYNUqqnpV/USH4TZRDMbHJhj3W6iBr8hP8RHF+b67gV7ISA
TfotYGcxHcpnWeWtzKWPXFFyn5mnvP56jn0RtUpNW733i4xIse/7mC26nkTo
JMjXukmmDuXhc9wPWJGOuLOmhhCr4eTqe4s+1SSbI0843Mb1B8Poyarndo9X
y/5VHD9EdbO2kyxHJCbsV6vHSn76q89r4jHYIYHP9KXOng9KKGFl7nDPR/bN
uGtMqj0trPGfffh+t2gWQpJudJ61BFGwJrq4Vc0uyK1OpmdAbfZJIhGN1qDo
9i/Sq7/25uZZVjhynYbfottEqD1ecp8yibm+J0Q6ZdCNM2HVfSYW7iKxqhhs
gRdv7SoSiIZnAMppLsdUDUY7pCFfEHBSAzTXSx71zx1M/kEpHEQ5vBR+r9dF
mnSvyar6NbUgTQv+1spbt4LoWAotwdYttEBaWP4QDDcnD7oKvSwyJyCjPMIL
iJAYyxZ2v0dXKsf9tuHdczrCDSKOmZOx0/sOjQQblBmgVG+QDa9Fh0O2NKHE
dY7hrfFUhQCuWYNZ6CkvG9v7xCaq5BTGUx+4+0VD3/mQnZYgvS1uA3JELiy2
vjW6w31L+CCNIB/9t1wudNuzQpL2joTjNYhc/HHc6b87/XcH1+F3GA5KRu4V
K6thmLOcFtqcf4xrFMzwEj/tfbT0iBw6e8zdeVH3bUmQ5VOCGsRLiX24awza
wxXUK2CJCDJqU5o6Li1AWFLVFRo8ooJVaLJGs/nJHXOTU0uQHxU51QrLrOir
SZSpJktvDBq7aeabd6acIaBbeN3gVXXcfac/NUM2dCPEERJCyTEA79dQid6N
1b9MDcxLyFwRGaA/TFyA8Dw5n45IyxAymfPbpHGEsneoezV3DLm/yWjzxat/
3+As/OljuiVWf+7xF85d+dExG5U+TIcENoGrQT7yL34XNYCCb7826zc7mCDc
LJg1lUfKjtz9h02S0Rkaw93A6WkfyHGYp4LYwBCv+SW8Y5ps5gxuPC0t2oPR
TjFomvfUUwFmDbp8czno3/x3CRa1syM3D9os5ilWtZrHSn0fbboqyYbY4F6y
23iWuExgPNlC+8xpwtp6ABBnCycmHwUMGqk4Y5F05bOgQk+rLCRAIVLjvQFt
5hY10jzTtcZLeYiaLnBGoJim4BvC+BVk08hb23dqAjifFmZLPVecBPj8epHm
56IA0QQkyBvlrG0hDqtmuYaw1e2SiYICwuuxIWwIBkw5rZDkl9nkQxQLyNR4
Sm+P2n3m+GtRSzap9UzTzgKhnBsumpSRQsABMWrpS47+ZJdWwEy6u8wEJT89
JnTGHvuZp4gFFOlqHKYNzlcOxqFXj8IBoeXK2TQSAV3nA4asG2Je7QYUs5ZW
7K/v7CY0YykHYpJu5n51cg1VWrz0hjJNJgSOQ9ULGWVEliQkoFI+3TUZ3FTC
GnyJIkh2y2SWlv4uXB82a6WCrYEQnAPKMuSdtmouceDMQ1VpAD515ww+ilyE
VCPNpG58UR9Zcb2h4YLgmfjkxirjC+yCSEqiBKw2dSJRfF8n/i5oJc4kywmN
f2yjbZu0nj1H/xdNLB2rpQBVCEZeCVjDwbEJ81tzMb83M9XD5ArSa7J07477
7wp7YikWtFS+64u9tC7jvr9tYy2qPbgqFHHn8/+FuL1/txxxM5EuFYw9YTdZ
kZzZft0xJ3oj7l3GEytM9Tp41KLeJPxkZ0OHm5GuVVqxsWzzvkhX0mXAZMdI
sFeO+77bSOiUrOQEHXwvauWzjb1S/s0LehQWtQwANTtO3m1hFvgJlPS0lcgT
ymmBqdqXuCrr2LQQt5+Ikf45fI+b//0ZdK5dIwwcAMxR4hDXiHZkYvSoxGmQ
J3vEZp56iecneqcO1lI7lAMVn+FUnDrHN8M2KSaVT3r/OfQ4zHbSLEfkTX2V
/8Q33JbE4VpA0WHC+R5NhPoXzO7PUuZy81BWKhmjil4jDh45vmkj38NmccZF
tFdFybNVi75LgcpoNRRuQvprhtKHVWFJHy9525RIu9lRL4COlaEAuM+CQghJ
94+mrZxIdhvprvwJkk7sAEgAuEMXXWsmtbnFRfpq5gWJwSNPXsceBWYD++Kh
NlXE7khkM7raj9Q3P99Mv3V7AqYWkWOEbsVNZdZc/h/kxwmK861d1WjfbvSu
F3RwM1LEQk6Iw2oyXzfXZiTzG3f1lGFfk/FkA01FJCGotKelCF6AfDqTTrQT
7gucZIF/blQGmd2DvQJdKDqgTd2P2nhx/gJcMlrAcIi0QgTFWNvZu/IqEKK1
2XiRhAz0cJRwLbhXz46mmKzqt2ZbXbnVdu3ZTThtctDXeJeuMPRgpUrMxwhw
tt7vCu9arz7WMc6mxVjOT8HRoB36/aXuexlurKAUVJvgHoB2/R4v5n11gCvS
qjAV9r2DMU5L1W/8MMI9OW3WwWwiTmKG4WTRp0pPNS8tIUrPpS5FGEV893EB
xjVNrdOw4pz1D6weiBTj2/XP1Qu+igxrD2oslZXe7sRBcd8G2t0vQVkV5kXP
wLEx+IiMj0Rg31DZGN4c7+AJ3O3dcW7csS0MgJvkxNdMEn5H6I65Yk8UXkO5
Gqgkqv6xU4wXbq9WXQxsk7o43pRnYFTcvI2iB4/MjidYhcCD2a8Sy3vZSQ+O
DM7DFfUvFsib/CIxK02EySkZCc7fQqpg3FAgLbImINO0os0gyOhulyJ6pmcM
2n7tcOJqnkxeemZJ1fYRFB2TmUW1Q+Xxh4dBfi5gYMUK2sne9UlCoIKM3YGZ
DiBIwWas9BTY2OrobpiMgVU7So4NJX8JKE8VOF+bRp1uHXDfmAocQAwOEnTP
PGXWn4TCjYeEzcf5SZkd/81We5hhpEAB9M4xZ8L6spDStwfbMqC2/lwsB+hS
P31bSsI1KEDYd1YbbvZa1X82aa8R8EPVjD0X2BrntRROrURQ10eV3jTCfMck
a1d/WHhsPvlmTsUdRiAZvim4/d9m12JVwUBoXe6NqugeAkxgdlorl0mzJCs9
Y8K9zeMQtrnjpDE3/LZaHioyg/ITXrrW5y9MlCRVKDMNdzYVHR1T7TDZ/EFr
tUbU38ba+qz/jPO0wJquKmGBfMk7G3j9rKr2k4iyuoyT9WUAjt2Y1UxO8V8q
c3XUVZgHUrNojZjpfTw/ZkTUmJyt1w/e53FbFsWLE7DlJRv+FKp0CcWYiuho
0UuLWN/fIKMPa1XD651UCti1HWck/2i9N2qn36cQVAxkUNKx3G7S9CAmHUF3
LFF5TJ4prPc4pyuqST8AmeCnJnqIyCwN7+3A66rpEpaWIeq01WDcYSi9wXD8
LO5HHdSeFmIV4lSDylrtNltsxpWIoGWnMlnPzDzOrw8cZzzbzNEpzh2Qv0pc
Ha2A1x7zwYEoaMPZd3BU4nBKKHId6hfB8CzLZtQJFa7b8ZCY5Id+uURSnmUF
r1f/fS3YhYc80RKwnvRR4gYY2M5HhbEuPS1IlVzKLZnWuDxL5DdLhCXITB52
dPThCL3EFz+w3QiglptGvLIlj7rBDc2a++EVgV8B4JyxuRQOGqxwkwTI+EU8
r50c8Pyl9JvQ/mlW+QWrEisUr3vAmmzucfiKqdH3TQOLtNfxWGY13UciygbP
rDlt8kF5AlNd1Htjoz4j3Ce7hswdJWf9uUeskDUvci2heeb0WS99qzfbbBMO
6ObaenYEfyBXAWvJpOOojcAapXK2XX7ZDJvPLzpeVD2tWujYBJk03hjiQ2rP
NoYH9mSJqIPWFPbVE4rZRNUK5bn6lgi2kv3m6PfKWjNXnKarUp5qNWiIVj3k
OuP/akTda5moLajCkT/GAxvFJKq7zkIdtlC/4kkHTZbGat0mSU3xAit/+JlZ
B03ZyXKOv8EE7b1WSdBFM5J8SKW8oGnEZ2+FAc22MUU7XWo7IJBlAONj4W9f
s3w5kx0Ca3lBbPXRP8KL+YMe6MlYdjkl/AIDKkC5hPA5srd9bCu5w2nNS/nS
qedUhWjOeecX/VGnjmPcBBX+eMiibgvx+HlSwJDZx9ZPJ+3vbi1GVoOIGocN
FH7Gz5KBtPnH0YLDHP70xAnApc6zPTw4+3XXh0Lm1a3tkV2Hjhj0jI9TErpZ
DhE56g4quznS6YRvsx7ykMIejOwgnkNFl6PN92aSC9bW+lw2WdD4Y6eB6ykq
Y0fABYdMsMMYBgsK41NFx0BrDLnaQNAsPeYiwAPLOGGyCTPm3XsvajWTO4Mq
mi4Z5pHW2zURnDADrUZmYGGWu8aqCH5NWcannWZWiublzBH0Z95oL4nXE9CK
mPmsDp/1IHxM4nM/t9EIEs0SEGKUIxIHCldirGrTbUgThA6SOh4Su4jervo2
RyUSm54JJd/Qd7+u15Y7xaqHIEQIPP6KZOnPWtLS+BinXJP3PemTXf22K5xs
zYsYdUD3rCoJo4NAd4UGSPbrLgZN9QvbJmPYXxddWvO+kkXiCkweCXj5y6Zr
vg6A1SLqIJrJ4HB4wbsihOLoGlcY997IB1yigfYUlJZY/kd0MwoLKlfTCzfX
nE7H8KEn84Wg9kF1OdR9d5ceMaz7MH5DsfV8Jwa8fi4maq/Qh6cZWuSSU6w8
6lMN5S1lRZ+s2EoQsZVAbj+gS5aTkRyf7EcBYemndfOLMi3TiagMg1oU2Jso
SdqmUDbP4eyV4tTw0QCf76c7MZlLQovF75MnFw0QqejaSf7dIAXsRyPgnCKQ
Qyk24x/5lGh7IVUxwSd5RCmPWsJRIWt7l9deeNjFxzBVT0mk9KOvLIogalXV
YU+v19s8G54UKiQ4yxohJoYT1tg1blwMmuQytGrsmtio94qW7cLokbjAhfGs
v/zoHSWhYnVwxtSJ1rl7/6L4ScZEzWZaj1gpFqigZkBbxNY6rtMQCD5SLIcr
D/0LRel3D2t9RFw9VGGe4BlPYoiLj7o0ONZUxl17dEg6PGuu5OO+QiSs3d4u
RMKiLn4eFWXBzV2Av2mcgkg5OzzunohzCH9UiN+3I6EXMDsKLltqXCq7Ao+5
t7ezPCp4SMVPvc5b/jgdiHtle6SJMmc0RXSPcWhz4JU0BJbaA+kjlQLSG8M5
d75X+ya7v5qhCiLWr/OnZU3QOa4JWaDnsCLFCCy0qrO1zROXT0hFPDpUa4L9
FReqzCclt0FSb7dKOV/r0sqa3k1m5XtG1irpgTP4JrVBbL5vQ3r6WwmYAibZ
obKXHVmbdx5xfvNZeaB9blJmx6hEldDb6j/mWq/JBRlAMpA1AZ7miUvwvjjc
ntgdIlvbPJfnV65OlH/8E8Ul066ijej5tYsER7s3nYpV0Zskms1SjMkAddEd
GDVy+PO3rkmGSxKidwWpANVofY05InxLAbu8NcEnBSTe9ytreIp8NnUbUqKS
xY7AAIAlSGq0THk1JnDF0PVbJc3ztZ1bo8+QyWOWSMnOS3L0j9CH0mW3b+ki
v0SLKhqK01lgUSva4iVqDHH2Ggvvr8ryh9npSBtUEtpgeB7EFxm6KIt4VHGz
ZI1/RhAix4yX43F4oRc2YKvWeQJEfVjjc7T2wIOoQBKLjx1O6xGecUXMooW0
RYo4xnBTau6GibeKGm1eyNckYZcr28aWAQr3dviGVfsUydbBvVf6bd4xJn80
BEdPZ2QmqM0bGM4Je0C9FhOfDLzWuBLofOcocWsXYTlxFYEGTqDSPGmrFYf/
FnOhsd4pi4O0t4pOby1ayfk2ArLCqBU6nf+KT1lj6SpJoKLReDCOxfMXdrbT
+ZIHvZ32mH6EZ0WxaXB2xNaaME7XrrIpccT1bD9V9A07k/WslWH5MCDXNWkr
QpCyrJQH0PFsj4EsdYsD4SkS1jYKS06czJ6h5HbuacUumLPLhL+o5S1ssyEV
7QiYYOpO/6ZikD3dyDvPur39BUkLiIEeX4Ak/gDMZb7kvtfZGnxfQniIa5XO
p8v1MPF+pWjwgaEdw+YbbLJ197hBedGRlmWKWtO2xIIUwMW2MCc99waQA6gn
hiI3dmRnYzMLA9GWWkJD1+EczBAQ5GE7knUZaQSFlKenERw7PWB4aD+Kou1E
ITglGhl0xiwUzoSZorGOEykxW9y6GK23XHzgTiRgvZsiTXBg7w7xsbx+bH56
Uaap0/8tr8SwyJAbj9gIRezbB9HkbC/pCZkW6lbUngTXbf2F5RgqrnevKvBj
ICR+KNCz3XEVq5pFYuKzPuFThrFAVFj+1xB3mjqcZApangkDl2vbzDusdOmM
2OLTFNlaNgs6q/9aiOYv7uf0ZzHMCwBlibk8akXnRVLPZetSQAhaP2vjuDmw
vmMJs4lQksMxr+6TcaoQ4NoQ/EjBgxh/Wwrx/MpGteLO2QHs0m2F/sO7mPS/
/zT1BOkmvvM1+l8tmeUu0heSvDL+rHajEpPWex/J/RNnf3lnr6r1vh98w5uw
8VPb4iHZEVIsrhRyomp8gwgGC0SN4cdVwZ3hxTirtfJXqi7KDQVL4JYsr7vk
WooIUP88LqHSzWc+CGy/qIeXeEK0jDn5x/jYTHGvHlTNLM0QTGZWQQoy31iJ
VUwtawdDAvQvnaGs5dh2avSWMxRSG0TBZJpHlRX8Fzu/sSsMQ096OUiHn3pP
3YkpMGajiXZQMQ8iUaaox0C162jNOUXPFGFVBQkihmJL3udV0zjE+pzWoWbl
0jndqmQGU0qiK3gahjb/TjKBt+CAvrLBMPBuX+lk7M2ABF9KGKbAm9RgqTe0
sWPT+fOh+9iqXtCwwUEEZAc4V+/ndPRDTePoVJGZXl7PfDuLa7IrK+PYNXE8
LT0MeaaDo7yE+cDvcM49fkSvU9dft/TU6FNQMSNxJInrWj8X9OjfzNVhFUbw
fosl45qa4e/NuBPQSAQ+5y7asRRQqROoQKCGeRsWzUhzJcdW0epB5FLAg4pd
9qvWiW9xT4L3Tw5Q9fYZtEDmbO32sGA77qg66A90FFH+RW5rAVbSiVcQYhm+
0lSj/u98cUQZTr8wL48Bgckgw885QdG26uziIWe5DaOruk6jj7A4OpUH5z81
9uJeIITj8T3CrHaarjLQ8Z+2lP83cPbNcdy3xvZ8CiFGk8+5bUK56hSOKrS2
bwTZkQh3phvGRx5Lu7gunnkFeNbhAsWENL/Qxf7IreWU0VCFfcgu2Qfu+HJr
lXd/8BNXc4AIoOgSZP7NHdouG3QvVb5Ext/HfhEg+O6LKYin0W4U8boxh1Hu
4Bl8vXLdRJF29s/nnab5kNMfp2kuDLQ+rwpzWV6FicbZ0Sfqiyw9Q9RnuaHk
puf9LqgVo4InncJ1fJRCf6N7TsjkgDqZpr93ZZvijtFUjMlLqDHy9owouORg
X85lBfFHBblh4tK3Eyn5S4xXZn5NnstHrihwBEekw4JB8CI4Z2fewquFPrmW
OaNDD5+awEFNSJyVJuFKFndDcRwr71wm7ek65ZM2KUIQ8DW5vi6IfXMC8w4c
68Z8FtFQT7uK6LvGHlIk4VX5TNAWp4ZsLPJm4Ad4DFq3dmiLLrSvywPQ7XNe
DJivSgZOQ53Anvvj3k725J3rBLLlu4s5iKPJPJUGBk/yCp+lHDBo/n0aY81I
AWU+2aOHe3TmpHZ9Mv1GrWMWPIdWPKK0TnUnPtJSiII6J1aU7elcjOdtL3m2
JVibPAZJiOjC3mFTCqytHS7a7z0MUabj75buWiBKFY6KhLRyQ/rRJVLzHQ7a
An4vPIrSpy2/1s8B2AnjfFcc3pCxBSz8KsMc5kiIDAaKazX2ONuGpeUx1VZ8
HNqyTVSiBbImRcsBpiwg4faTDwe802BtwrrbUIa16nf6f9G8YMbCCeozesEH
3XwxlC4tILkQwopVW9b5Q1REi0sZLsgCht+roWUPrfEKKIBJ26GfHKvMREtS
74XI/GFf8PMh9jb8k13vdEUXMdkfF9chngQa1mcQ/bhHUWUqFfvF5Xxrmgk9
9Ka+q+fpc1nK6Nb//eV2RZKrbWRTRVSLqmMU4H0S2F6luE/fHB+NHbKKnIBc
PwjfDqVx/OSOCNZhVWPTlr16th4+wIxecCMZuGC7lLz+BjTcOBdsPjo7T+bb
ddOR8TlFCOIU3ftOC2234BBmsOaNJpZLT4uqFuYS2FcHUgxnkBLKWSc3thg8
V4h3AGUjmLRwQze9/fUR/fZ6eAaOSglXAu2tsDiD1i35Ayk9KUlqkLZKIQLR
UuSodShxKBBrBA5PhVA9isekMTRcQLnViOVwN7Yb+e929RdQd2LqquRKo8Rb
/om7sNqKyNDHUpjdFARlAQrDZPn6LUU4Df5b6saN4iKB2DGiwxeLw9pWxIiF
+ivA09BoxZszGm6Qc8IwqF27dJwy8a/1D6m0kHb/05dOmlaVGI18n06LamtX
YBLIL4jL0JmVfUhVTWWQvtSU67AuiG3f62ooEIHMx3hOaluO5ANl5J5kbYDY
+xRphqcKWM1lwoQFBaIQiOc0frmLA+j/nd2kKDA96j1Qos1B8vSLx4rJZwFM
20Ti71+7KixpOU2qzdmsLM0Fsh8TixxzCHe85omw30uZ6nw4Jp8IHpS+3RRx
omZUyWywRe0/YNDj7MpSkSVNqnixS6XLr35UyKGJ1A9ozQItjCHe6XoS4Er7
76VivX5nAJs2faGXepxiWDGZCcxUa6IWLPcLj+cxhmeZx/T2NG87ptqwQagA
mu5dzPwrVSU8nMWjUTBNl7i60PA2Ss2kMr7Q1iYBh3sPspQEOgVrE9qPS5hi
MOLj1IFyryEqczEe9hyru9F/mfTvuF5m7ExugmRS0AnjabAXPGG19VC2h+GP
oBACKcuJ9Y1llEHQo1Sq9706OgJVViDN6eiyGRInYMAXssW2YSRGCixSprEj
nAUtAwPr3aKLARO9toFa8UxPpkae+iWN1E/cUPewO2djE/ivCkojQTEGzsKa
1XSzACj9qhZnB5RN9efjS5RluiJ8o+4x2CCP6wMPWBn2c2YKhes9eWQzMVCH
ysZKP886I1mPYR3+fs+g5aA8UmLx051xKo+b8Mq82NunI4tMOcjBek+i7slB
wX6QrIPBJ+S/R4HOXfuKYVez7NEzncqPT2vOUvG2hfGv8a0ryK2aIXMRl/eN
x1oRHN9q6MfQAyZClNvgZvCX4T60rRU+sESQSeZS4e+aw3YPR7tFK0sUJzGP
4ZM+4epYIKyqaPgj22Af+7th1nHOxJ0P2G3Txg86SuwMps8y3OeEUigRIIL/
XGF3yXjUmRTE1tRcACxTSU4Al4CpOvvzjHXqqHWpE1fzWai/Umg+ve+flTqE
YddXkvyht6mC06dQ4nNFVU1Zz+FyVnszsq5JgaWewf/LUolsfOXenwdsV5Yg
r5bGU9GQrFCXnUhVl0p35O/b+jhuiSBs5BvTPKhWvCu/e8ri+kSOy/JOvIe2
P8h2VVn7Omo89O85NuNvGjIbDND7ONQuRu6bicrLVllK6/lo0jmKVJBpmGo1
2FVJRuAaXlRQTZ4rASEyST/ZpGV8xZtIFCJF3CBQrr45Un8zt/8/CR6fzJnS
WikyYXJUZiHuQ4fH1bK34eoMrXmZ/6KTl8zHZzm1TBM0V1+afydxfa/kk+kp
uDRVZsi3J0Ofq2UxuiCny5ne/4iYmVLxiOr14tm8YEn+bdgtXmxYEg1CO1sM
cpzq1T7/xGKQYqxo6vtC3lghVZtEm+ngut8iEQsps8vuaoTbZUb3Ab6/iKTn
XWA9IDfgiFk/ffskoejTwB83JkTPIE/9PLO+oD/qihF8MToRiuuq6syZnRKO
I23/SWtiXzVwyJLkza1LCMjaXr2m4dMQ1xQMWen/eSr6dGV5Nita4rWlUQkg
OjZhQu9ZKOrW3eMcWZGKRZPIXMiVSWkCwQ1EH8JcxIyln39Fu0tQWvKrReJz
ZZs9EQwPyp3GEteu7XccErn/COE0Xl5etT4e2O5/r2dZ0YJM/2EMSSO9E20b
isX5k0gIfiVlqWGW6Idx2y6qwv9kb7jXSh7dMTEvQYLbVVhxcDp6IfaghZNf
42H5abzizL+N7Bg140yaOMGSbQ74LIXA7QOVSYbsGVCKb8y2u65ouRfQ9YQ3
GnL3Zg+oRjSY9GPIGK+uv/FT4PaANL2t1UNYCneVGtJuA7FjnfizGjIdEqae
QKHPeU9dpgbb7d4kx3devJcD/zbxucl/z3PVFg6kDFkrWUYpXiQA/No81r/c
tUXxte+EcFmSfi9QhjmVL407Xd/IYAJHnFw0djL0hfc6Tk2rru8dESCD1mfX
JF8mEZZKDbDS2dgiNNfFZsuiDyZYXcrNM9f7mBljoCvIy6taGKKLQL7bgt/n
fB0ENjqCw9RhhsY0exR4uawKzG0lfrpVw+6+4s+8P0pfHRSGgUa4fdUiUGbu
YESQPXNLXCKl60FuahUSxf4nKxHa7Dx2A97k9KRadU+MufkTDLaW/PEZ4lUs
i987/HMKzvNFI/5/QrGf47IV2LqI0OmWr0QC5bQPv6+K1RtL/8F0yyiDNvP4
i7+7azMYQXK5lLAPgI19giqm+AL6OdxCVSvLSydIxEVL0dlU6T0jFkKhh3n3
zlCiIWCPcFjCDEJ9PN3CQ5yLzSF8LazEdk80O/chOnGt8EA3duvDjXzPhI84
FKbNxvCb4DHVdI27Imfz1A4nWzngRte8Pz6mulJBeLcnfEbGYvGe9d9LiWE8
l0d2ZaxVwiUi5a1HSKZre1LXkSg/0E95YDBFaX2f2LYY7LIXI2jQiZ5dDxey
achgB/5KwDOXsx2PVXpdslJRzRb3d8Ufe8TjhTKfGWkZ16BO76emAxgNI40F
PGVOnMB3mBPzPF0tT3ve9PaSS6KS+wmqirZc5BI2P4UHZnFMJkb+8L6oxe96
4CVzLgsPWKNW9iuNN9+1Ll19+esGm90hKdzYQVhUoFZquaNN8pdrofIf+vFj
2K6fwlxEHZNt1v4I1jHkJE3iEcaBTPRz52ENFgKnycVg/9NAsv4PwRPveWrU
q1ScQM5SaEab2yTNuq03Vepxcq+JmwsjcY/Dygy2W3yqFsPDi+WbmvUTRnet
L3t204kSy1cxhXiUIMLZtYPUpPGhYTMJV3hGXmeibg/ic3nSE153CYIIr0PU
6S8tYWNfwpyqnT6Vq1RrUMcFpXPR+WjAtwEBZ0TVLft/bzF3GSgkQUzU+BO5
yofpWkVsd7E6rRjfhl51YQrL5BxIRy0xVszaPZ1KZzDani5IPdy2438ZhBhs
CUmnWJhS0N3AiRRjawPd8wczcso9IMSLiS5mID+xkA/oVk8rUgiqximu23Bq
+4Q9jtcqp+s9IRtHIKuVCRNI92BUjhfj1wHb+mw71Y0SdRXhGAH4jZESsEeR
WfwgtO60pG3g3pZhlC0RmyUpVp0SO9Zu/TgAmstsI9Oxa08JZDQiGbYfcg4l
Mg3OPxnGqNqXekbwVtB7COguSqVPYvDzOCcTzIKx/V1Lk7aSmpjmgo80K7fC
tUK6bnqjaF3k7vh4OMVXKtAFK9Q61QPRLmbR48lqCEBUG9iWyK1P5GL7Xaj7
aqHab/KcyorAnOyhLTMEVN19oElZNBL/loWf900QRwrIC5KoVv9XhL+9Tr7Q
celxVSaokTYRwy/MNC6M7WRFd5O8qHhHmqZXbSSCL0WC4GRU4V0pc2SpM/as
IFRRPawifSKWsoTj9nV51Uno4TKE+0irAQzghIH5nr2Y5ZC8dYorGAm0RdOZ
WdiKGDsoqWHhGOlNHAHOEYTKqsUBimf25HJ8VSO6cxvykEVfHwrKG0vFAd9k
W37m7fVIqwlkv3hHr5TSWRPecuJCOOEtzDMNfDw9akTffd7/70l1ywuJwyFM
XxVePCo8W7yUuT1l2XcMvd510mGcbNqvgYrcuk5LAIJRWrSOJJqHq7+EPqlO
lhl7rhUn9mc98yxx3LirH23RRNsDLpaoPPvk3ItaCMCT/AHwc2D4KeeSk5Sp
rfOD9WJ3FzN0AKTbXdoj2AgtgSw6+TP/hJvW4TP+5vb1A8FQiSQZk9RSf8cM
w9sj5oOhOKYSvE1YRD/nCVyufYXNchbbw/PovKhtliEjShYrGP94gJHxh9u5
Uh0NUIrkNmtQo9JMGo/0ByJnPvLc27PBo5n7nEKc52E3ke/hDi8sMH/ixLjG
faCk0rzIoaN/fm2fpIFAuonF5llkFEpqvWWVBy5CSyES0lIf0MtytYJWBsG0
pvOZE9P85BiLzCIas+dRrJgXamuGMyebMGb4yVWI6McOmJsOcjzFY3ZCkFSo
uLkDTchH8i3Oab5xHuBXq6khxj7uPExaevxDUb8K1NMkDb81DTS+K3BN5c/7
3tHvab4GpXJlih5WkP+DBobz0pHWFxLhLx64pLtO/Qj7ari8Aq6rAwaJgmzj
OGRuac2urgaskQeQE1fND6teocVGpwm+XwTqfM4TV7Px16ulcHi8tcnE1VuU
LuDFxrlnrqpCmwiWNNfzBnRrm+u9/i5AMhk9/V4sFwe4KWjcU/EZnslsR9rj
xFcl+7EHtCCFSPAYVjgP6zNsFwqFOytNChuoqgz6lKb1YI6aY4k2QuREgGA3
ZDFsw4j10rG7H5ccIgy8NQBGvis66rfFXWjl4ZU7pKVjNM9XVN/eTeCLtvtZ
BMRJmEK0rFrI+WvtBwHiwzDNxb3mGSZjfvu6BE9K0G1Pdbafwew2B9kVSslF
e0B+YP5G4qSb4fpXpH8l366UIj5sIlX0Z73HVWRoWe1MrI3J4nSxBQL82FNB
ECVwStpxV02rVunE0P536bcZCtelTVL84xtU62w7GIas/X2bwMbOUj6RhAc4
bppnKcIIgMF6rRXID+nImVya9wLcE0VErRkP5uUjVLtBe+bRipf44THWZio4
VZsiPGiQTHeD4oG8Wv7KPrNEY8HQYBB6EnsnTAsucSiL83wN0yq1WVTOu+d8
cnxoqQI+rNvYC+db3gp0HPGqEREogj79oc1I4FNkBUSGTel9Ihxz+Gy1WAb1
RR2EJMPXN3P7a9pMlUlGO4+VK6F/nmBsl5uWCCezp1qKZ39fBkqn+1wUdVEi
nmJKym2tbTY+K1m0KnkHsh4qxSViw0KjKQtnjkiQuX0c/n2ufYLaNNhJTDKQ
xDZkUGrDiwRKJXvNXa3iKJFj8e06dRkP3Mpvxi3W/h7xOzlIQVxEvIwp8wH6
vI6n2i/dkdHme/FGSlpm5H8xSkONTpOUF5EigkJBPMIh7dtpsYdOVJQAB3UP
8vrp4/JjAJddp5UpN8z1O24NsapqQzic9fsdbb7LjfV10Co5D0TB/F1lTArP
s3bvhWWQD3Feq2ftKJ20sj2SSJNPOC/5Zqftu6uIcSB2I9J650vFmmj6hNwh
hXlImzwRA/eIJBrU09Fkeh2PWp2XaIw3/3pCQLfI84Qij6MdcqtkLJzPHOT3
N2OMRBdAaHhtjcmRqovbbQpFUGRAVYU+8TvSeuGimwErkR8hnwQC1z0eRoAH
8QLwB8UeG/hfVe79BTmQgZRxpCVrmvpwtNl4Nt9N/nIB53ENp0hQ/MprM3N6
KeWR5BRbnd3CeX3+GSg7ThMoE4wM1s7Qm9/5qpzC0czBiGdWMfJuvZoq/sYC
8YjR+Al64HBQSwyv/c3nrrfSuRstNqJoi2Gm3cTrVRwU6+62Slu7nfLwVBIp
K2gCD1q5oc2FxHS7jZ82xDTF5JJ48H7KRTXu3OcVfuNyQ07KiCB/XY0EJMBU
428NPQA8OgXtDv8XJNZr5fOIURl4FqdoiS/FvNk4HNEUH1zqA62BezMV3tem
GkDoopgSjNFb6A0W6AYeDykQdvE8lEeOu3gVDqleL6SXj4cWZLgf/dRTfFj3
pnRzCmvRE+JQOShR57BRPn6WGk36tUjG8AaEbD5l7AZ4+zg3YmFWQjHV4oBE
kSOZq35bbTGRb7yMYRnvxUnrtlQnPOqgFWcl/E1qDWfdBL+rSIMHsdS0JAec
Ro61y1nJjs0mQbyC+gzB18YbBsLJsTYGNEPgLV+JxmM8TgJtLw/94Lkr5kb/
qIP5NMpe00hlFuCvciJlx8vhIQ0rlCmF8WtQ439LzXc0GhsAfABMA9uxpSvK
RM/innPCA/ZmpnQ9bWaMLIETqAHDx3CeezdDzsbRKWNNvO47ctlE9joc1JZe
6vcdSjTMIjs+fecy6WwcTlGPQvNh3XABHViGReq1UqGwga4e54Rh5PWChx2Z
vlKO/+iMqb6BBXyc39kwXpzszPoVcksUKI1+GoL4jisCUd86ySAbZJpYfshi
7csmuJvQHT5NZZEk1gV2CM3S+aKnUln3St3QL/d5UHairHh4B5NqQKv4stNo
Z8Dt5skCI8I4R2UwVidsgXRji3WJlQHtt4dOhf4xGr32znxuFVVY/x87xwp3
lXG6NDEftkeZWP0PzMU6/FpSztfWmqgBG7XM2lczSzKBqpWEX055bnx03pQw
GPYl5y1ZMuVfgovOfYx84q7JPGS/6NdLxBUClrp3pnWvPW3SAyvPsKbws/vW
3mgk/WXraSwNWn/+wUXBOJI949Z0w5rxDVaJDs6hc07rPLqDeJMqF1DvJ04D
JrmteZYcaByCjKs3Vh3AyMU5GotT2kA3aZq7e1tjg0URrhw5NgrjRvMUzAyb
WPGDbcp584Wrh/UrwVWu6clbQsAW0wtgYfbnhqmQeGsPRfoKIG1gx0p1GcV+
VLh7iGJ4trmTXUuMo7hFn4VQpKdaSp7F5rvXcOkCCnIxCqCYDhLnLDzQx9Aw
Tbp+xYwUU/0BlnpbrQXBtCJ2K5PTGS8abqEF5rPJqjyQXHyViKYOx9UO7FCS
8v8gdVktYOBgThvj1Vd2DbKn4sQ40UZcBN9Q5N7LNl/G3bP+eBuvdgxLscvH
gemmg7mz5AcgWHC8xk7fSxqy/ZQxF/9TTu/LS/J+l4xg8XL8E3PGT0qotF6Y
OPvBZHvorOQWxMj1/VBwRtP8KDIecxFCmAmU34gtQ0xotZv89glwdtQrA4L0
MQot6howuJf7SCjtyoCCeYX9gCsjZrnJkF0fl3LvwOlKGGgTx5MgESkk6p6j
sW/5xQA9JqcYDgCQSuEo9MDLH914T/X7fDYRHvHM9/zprOOKt+Iuguvks8FN
sWXQTykfIZwM5LovJpRpP0RwpmMGSAq1W8i50nkRxjUcgwPIMntA2prkWQFV
FCCjSDAK3GALHvLPKKnsEd6UDlhTwbqSrgiZU9DYNnXf9RO1E7G81KRGMeOX
1Mlag8e6yBbjKeJ35Z3OlTBObDq3tBOZc43btLRDueW3TjuIR+BmbIGM/LJx
TKrK3atLpfl4FXjUDGM0VsWSkJfDDfLnPa+OPmVbqXuQMxZAqCQAPgrfvHBo
K0W5DU45ra4ZEbzNIkuP7IX+a9n1VPMRfESy/NyDGNU92o7bU4UeL8WBnKW4
Xpl/OfWTnEiy+e4DlQjmpc38B1XqUgxMYbJyY/tg4mEjNE8k+RxmD9DrVoW+
zptBEN5rAFm/PZZ6cz8TvCEjftsjOTr6iMHpha4ZMy08uX82+yr23w4ORZ3B
8kcFfXXYFnpZ9zzK6n6yw/zv6i8ASS7yGI9j+ruynJ+9GDoa0tAJi22VjDN7
+DV9xTrtr0yP77u1/QMhalvSRkO6EGum574sPhYoLUJ27ryk67PWPhhGwY4t
+/0OpaIxc1T1F08MPdI55ei7/z+pyfbxkph/S4X3/1TEY+6m1viOVSDupeAd
lzzWVpxVw4qzJnjx8Ui3V8KYTrK/WhkMzvFYiy/8uREUuYhF5CVo2Mf/GajD
ilC+LkQl5gGAZzQJDD0ZV3Slvmj0gzy3queX5SJgNd8Se8RJVz/u3e6oVnc3
ooBmXvTYQMyAvG5cbdj/jGkIqQRsFsbLbwJRab7iJIDxWm1MT1LxNfJUt5eb
t40WBilqnwuCdOs/Gkp40ndHjUgtdh8gsUOZ8Ov4ZYdjh7R/3pEdsyzc3wZs
KM+TdlreD4VQUC4ucGFhdAiZ3UtnWkxRSnAGotyXAT2BJjzSlRjk3zbqALiW
kshibSlv5MThXxpRYrLSJO4SIwhilNACrDa53CLnD7gvaWwGmlI6wm/DGw7i
kqXwe+kDwnnT6fUPnqJ+YF/3PCgB49UDdxhWQbK3d1wZBoVVWadBkkBVop7q
rDqBnN+NmJzrY3QIUs99LO5KYCAXnQ1ljQ7C06HsbMEmls8lY7RgU4rzSlAV
nBVHeHJ/lz+ktukA+ikS84rrhSqS1wSnmGIwcKm3ONtIIsD9WRNCNgIBdtyu
Y3WviS5C9yruLTURIdH7nCkqiURUyL5Unu6tHHymprxv3y59zMo9ZB4LldMW
JxpyS4F0wHaTyge8mpGmn6NSPolMKJftNQxt/eQDtb+jvb7J3AUV4E+/HJz/
0BYNLRp9BzWM+0RwMXcmj/4HktRv+uL6lqYbM+qMylcmgtCB5YOVA4UlOUWE
Q3wrjsJAVY7AKVWPytrC/LKuxvcBJcLU0cw+AZsVqxK3Yuqk2V8s35rpJIr4
6xaVZ8y7/m2oV0Xz9qDHBH0JMfTp7BuI/V8BX9SXsV9bk8hI3D6ExPN5iS2P
KhRgqJCIhAf3wAK4MDD/N7n1NzADSvDFlUl8aydH7HS3lkxOgLJj3/z+B/br
zx2xeBKGW9hSZfnoFA5PXLaK8nk7OrWTyCHRlqhA/wZI1jHYlVxc8BMfUHf8
MZxeSgfyLzLXesX6dKDb8RD8VVoCSJBGWhIfsYHpab4eRDthiLng9j+NFe15
l+m86MVJR+tkpnSgT0AT8TKXE+U55joAwSFkruFnLesIHMPL9G+jMw2IlueF
Nj3Vk+LyU/y94HjsBMaJEkcOM6vAbNdcxyzxtgXxJ9lEooGGh/7KmHyAkR0r
oenjFsgsaO4kaTCEk74EiMa58LFRVTia/T6bEfuIxwMHAiIZjsL2IBUM/MAw
40GoE1M95gFIjHMiYj8uf77OYj5d/TEPrnl4Ep7RCNIsqW0qVS4Q74hWMXzU
AzQLyyou8gR9XT7ihZT1rVlWehbNB5JxZxuBW4PyM5Hb2Qj0UYuUyNcyAVhn
jqf3zRO900H87+pjcVsR1tbeW2MvW0aFRmrs0CnPP9r0LiDDaFAUzZQznNrm
vIVLdOq2ezpDV1GSFstTCbYdTqb7wYTqQ6gN5zeDn5fqpq9iZqJD0ZZ5Fob9
ezgYWt1BJrzF5eCaeoUDSIq8OcaypjqZo6vsjGuz6k/qOCr5/BwhFbwpZ7E4
ZC6e/PrGWCZTGE7kdB2d/Zaw939sGuIgr1fh6VXsYoWFK/mu4p9fP8afrIHu
8xD69km/3PTOJ+PHBwKnFxRcafp1gviztFoMRk/3Wm8X5wEb1pYQXOyUAuGd
1foFd3CEYgF19a4lazUTBF28dCMrz+7H5BZDgOYiFE1uYhA4PEZjpD6izNdL
rJR9WU6Cs+0smNmbJP+ZAXeudzLV+za/cGhi9zbo+09NSHC3QnaNQ8n0RSUz
D/f0TGYxOt/tJH9GyNwHklbtk9JtQGrbiYA/Mvx4r1clZY+HZMm8mBMADFCc
E5yZ71HWbGyy3hdDQgcFEbgbumCuEDkG0MyWxPUFYwtO7c/CD+oMgju9NPDs
mkZybUMcm1Zg0cCTJukoofxPEXgQrzzU6XcIInah+ti9vmx34zhLHzafyL/D
vFVCjRl/y0W9lf2MNcoUgN75EXypbhzeG1XWvWDEWLiDOhBNm68o2+Uh1Jwb
uT0Sz7N85MbH++kqgFUWo4Ic9RuCKDsVZZQ9KwNCOXWdEOfR7g+W/YRfA01u
izU/xGfC+QYgptQdlirP7oONHfQxW9IbsO6F7vynZKAnlT0r4hQXrF6TQ+aL
a1gl1abz9NH4Hw3g62oJoq/Fj8GVGaC/9wF/ojdkZaqabMKpnwx3RFrxLsRN
H4vIiRkMYLOnXHCVUBoKtn7eqCu0Yc0lntU9b7qvjbw1qkHWZ6EvAJwDJ4LN
8v6/DzDvsUw27vaThpcCZQhHtD3KI0fLslsrmgmmL9n1k66gfo2JCLns6veF
kxD4X33dzWqOjPob6ySNX9bqweMBwsMwJ8rYjkJGBz9zbuoMCDQvMXrrB+0z
we3c9moJTbGgW/lvX3dQuGDHo5LR6wbyAG+raaIs2Oe1V1oOdzL6gHOk9/Jl
p0QSdc/mNVufThGOpNtHYwhszJnFVubvh+m8T0eMgF/8RkahcT0DToHwpp/8
APCzIh5f+3inFHGrE75j+bSZ9XOO4Q1GDohrFEjTkzlh2T/IoMMiPBdIZ3K8
yOSAZlcgfzhQ0r6u+E3mbYKzO0/4Wb9xWc/Nl112Q5VK/1SOVnvLdVnuuf4h
Ch15P7nWxaiflbwfMY4SdY6pMtBbH6aDowPXwWeb0+orDh7fCSDY63HMPlt1
+IkLADyGSga7GtnMu/C5L7Qr9bzuIOU2pfXZAIGEOs3z5MXVc8L1YqjyU3V9
dyGOkBCxAAF+YVeK9D4SZuBeAJF1j01Z9nXjT/Vj7h9tXoKDLVoUTG72vO/Y
QsCG0GX5FXJHD5UVD39tzS1TKRfbOnVEowBLcERA6MdZAZ2Cim5eOFGAaER9
MrMh4g7B5sDsuZ0QFztOFFXAEc3mBWmQJATmoBHe5xl2uDEIrdZfOVlCZuFV
8h/gUbMUCJYsbIyc23xkMnF/qW/Hhp6wSPsc9z6uD9A+itXPfjeNdxtgNaCm
KjlYLKrlpAZsz/a2f+8rXDU02fKYMDqBjOWvFbCi+TaD4RpiRgxqdCft+/w9
Gh3IeeMdWuYs2OeBDvsRDsaBI8DpD5624DMQwkJ5iHzVZY2KBW4OQ9vSEIge
uTOiZhqWw4Ze+IVaH1+QbmJd3uS+HuzyFrG4tS69VuKWvulCkCRHnWcjcfTW
CXQ6NlQmOM59EjqhKQcBH5QXFSkfR0zp3or5h2huafo+6VtX46nhUnZfxA7p
s2NTIF7kO0fEkT0hOlH+omhX8fjJq34TMcIDfO1HXWAvF4BKCM9GV7qbw/v7
izemAb+RW7gZycTxVacCiZcqRMdNauMJDlxV3ox0SL+iyudxzxTPSKReIyAN
7qjooLfyGqHVntPgyPTpbOmUfnfih7qKPzIsh9hJkNTlONX7UWN7TkXUE0B1
n6t7O9M3fbl9dleyO/ONFRNymOIOiRjz+Wj+h6tMB8r0DqfbQkrFjUXcSUzy
6LeLbq7Q2qzyepkN4cJrnN76v+dE1VB6W3e4C3GpEUnSjxwRbEidzWV9o5LT
5OEx73RQZ+UjJV18I2dIcrEatdPkc9vzxPlIb8DYe6daMXAByiP+rDD4DJKZ
+TnjO8CQkn7OHdcgVPOSYoocAHr5uDW0srB3ChiyUimIea3LANSfVyJnEeRu
oEmmEvPWnAoQ/v3IomBxd2i57SUkz18aXD5XXtk1Vun1WA7joax3PXRnuZf+
awAecqH5oqbnaDudnnfIx5aiv7HBFNMgsJ8s9SPRvRTyUAjfkiJfjGiKnpzZ
InbxzZu3S5DR6LeHATyy3OvPIaxKGDxeNk2cO7Gn2LqwNFFOqNkU8ief/tFJ
oXFFLDNwa43+9/lvPIATMvYevj8HV+lhWvyJr02Bj8bRTtkFolbUoBoTQ2BK
gfpyhh0jXI3SsMpCjILUp06iAap5ayQKM4Ea8oiYZnP91Cbxp3Qwe39bWFvQ
oidLIR0cbkjsaOsrpVHF3w6tag1jVOtKIV2lIzKV3bsvCOBKzAJluRXwCx1E
+xznVuZEhAjF/awO9URCsvW9Ju6j9VUze0jw7q++/8/1tnmjN+FSvx3LvE7/
howepn7DrInFVuqa2jxzyWE2fiXZx2jljfMQHMK7a8EHxOlcyIZhjmm3B+d9
eH/ytHH3hwGsYu82yf3sOlh4nrPulRQYxawY6wQgLbmaH0w2Wo5ivcG3o+GQ
V77z7cG2oBSgnnuD2drGqJvjAMJs5a7jQBoWDhyu4C99SdHyDP84q94gcjgo
MRSPFSZCIR3lRHnOzaSIEaQiAnels5m3w9pPSo77O7dumvNhhgn6VJH8HKEm
cnQd7jZBgqjrlDGnewA0J6HnHiN0xTi+CAWi4r2qhlA+oWZO+shp+qKZK5qH
Q7if33eOVI5gN8aGN0zcPeivzoFjLzqwbwSccGTuHwzttNs2E3PRQflg6Ayz
sCuDBocaONe/4K6/15aR69y+TIcZZm/9E+o+5ZAVGgWUAPUwLQ49vQZ02Q2N
QTK5XvW/nUh3x8E/qHMIZUyByGoUFvoAR5doJ/iIC7vH8qkPIuejcdZ5KoqN
QaMqPw80LAGiPKtn855CsbsiKhJ/dzj2T12T694Uoob+2pm/brwJqUyZJSGp
Y1QPocz/mARmM0fKK9ZuLY4hLxWtBxWZDI9CKKbqg2Fsu39R1i0t/I7+xlA6
hpFEFHRQHxxFiQn+FGttLCN6X4IPIT/TBdFO2AvUKSaIPplGhJnpPvJuMrVw
5vImWE0GunvZMXIJh+0mbuTXxHdGMMedGqfiKwtfDwMWBGtRosdC9hnxAZZ3
NHppF/0UEDa1LD3Ts2P/GARJjuxx391LQdRqVvDpoFHaRS13cYda74T9maBN
H+kiKQflbitlDLD3LQWHwe4FVsC6BNQQKkV2/8l/CU96rbld1OzDAsyInG6D
d2aBEX2R6Nuk8+Li7NldTFBfB1ASDTYJ6HhBxna5IMjvA3bxn1BP3xKtFUzj
LYTytkq6R2ZIeG56QDv37ihhaDjaCXJPxq7k9k1AXnggZofqI+ebyDC5WArr
yyHPAzPe1h9ixktqtgM6Q7QMBBXCNj3OMyGqmFMR7LkgmYhGbK8fj+MIvHAO
0/7LEILfO5JU7t0wQ3PoZYnqprqbzPKv6abPqqJDcK/1DChgo2MsQp5mTC9y
WAaVOg8pa0AmvQUY+qHLlxK030P6YO7begRYRR/OheXgLB4uCIOcwCDcMZ2W
Uw6vuocApBdQ02336cWXSZfv1AmxxGtJD97yOfpxbX8/UISXpBpJxEi2u3D8
2sQirzXOo2ZvaaLijsU+k2oDHeoQDNTpyH2RQiRUQ21i10jf1k5cYFbt2jZR
biS2liAmah5OZkJ92bdO/t2Z8DZSl445FE5sCmSLjof/wJ2Qq0BNTCDUjm8U
A0g4BcTf1BAd24XFVcF1OYHJGdkMQBiX9Ysd4fJYmi52UL2AVeUdWtDN8Pre
XPncINeLaOlJgjpdpQRe70FzuPuKUlX2xL+lYh/dO+phiyLpt04LcXegfLMr
kOn7obgHrizgdOv4EaXgaKNJJAusI4qI3q0azU2l6zC6EUk9Ghs25WV3E8A3
rlDC/EkbT95IlS36432LpdN1V1BsZvRQVn30HAf6C/+ZhhNatNzKTyn8TSpk
kCDiX+Afd2tqU1f9HLRrdhBEAwbA77cwS+FFIN3JgcZM79eYTo7blnqEp/p6
il+rxk0tN/MzFJKyRfL12S2FloJY7SnjkBZ1PnQP4qutH5TDGaP+nXuruaVn
vw8voeHg4IXU1MbCgUH9c9+u9ZHHGJhqElMW4JQtm3CwAuhrciXqH+Ji3H1y
aOimW6W+EOsz2uGyu1l/PtyC0RK9k7Defjl/F+mKUz2jiOm5p49xsufeLoZd
ndyMddCkfDZgvnBxm8kB9/Z0K951l2ijhG7ILLFXEwOWHyxUw+/DIVGbcVJW
sQXmgEUXuyzreKvcA3ReS8tLi+/wdd2935GLLPLl986OIR3EFEeTmZVOWwG8
W1EHfzTB/K3TlHRvf4F+kX/udwllxvbTiTAxZj3/aq0Y/gV8KitTnJB3pn/G
z15n3X3IC0x9N9ifAdOKQA6c+KCNyxzffhRB0uesjGP8T6IjmCABsyEXcklC
yayWdF+iQ3b+WFvzJmRvMNoI8LR/5FPImsIJgjH4TLVva1Xkq9Mxx2AobPl4
ePfPTKYZmNcEij2ATNXMym3Nn5CN7dxfjDSXy0WwnVUZopCt2HF70oqFVI/6
lhosgDg6bhbsHtC728Mvts9tQv9qJ4X8ndlDXqLKAlDWi7YRAMP5PQ2LAUea
PoHdfCq9kjHeInWf3ke/zVbhLj6XRyoRyR6CZTRNsv0tZXwSlcp2Q2rsgTJV
lZWbjhc2eNw0PQH6vHE9FmtrARtxkb5hDM2Rfek4b/QWZT44HEGKVtMz+TMG
VtFlw/9rJY1uOCGn6XnrTPTlVstA7txBW+ANxLfLlehlwj5gOnUPRjQ/wQj4
zp49vA8pPuBQnEmM2Po/cFWVK/6m2E1Rq8efB+yb72SCFz1dvBD62dpB3Oe1
rfME7HTTOX+TheFvLSl3FbMvV8tsshEFxANsAZcm7xcqdtujQg22aem11mBQ
tn4fGQwOenfL2pPll4V5sBXlxv1zw7SFupScb7hRPmYChwb0SBlYH6gHS3tn
7NgF8sDMuaKMSawdvFj2VnL26nm78YO+Omflk7VwK5XJ7Cc7XhaKrHWTcxH3
Of9BnMjpo8hh6sn3rehHzD3Xl7L1gsn6Or0YmkBF+NZuzltW/s/W+iU0ZWjU
hiUNqGN34XpecBHEDq8vcRLB03Q5v07WKmfR9FKAMpWDUi4+Z1bJ6Ia84NG8
cAubwqqcfq6F7seOwRPy+3HbWkpUNrf1AxJY4PYh9nMuycGMtWRffuMJhJam
UErK/xPMOWdhuWrlWDqfaNZ59moMhnN9ncC1F//kHCReMEh/dadNTBoZQLUA
eiTYk7KbRsCBuY6lmC5JeB5bMc+2goqVhHjkkPls37dwXA6UAH99QXPnS5Da
CehTI3FENmLVSIs5/RCc8dJkfcNq2SysdxRgF+MDO27JVWMk966K5X9SZL9k
I/VYXiWkhFKJyjIIRproD6ZU0kBdW0ku5Eza3PXITVcR5MI3L2VZe8vbzq5S
KQV6uLHUgOWQFzpgbbgc9E/QLbQXLvtYWeQmRzICiQNZGuRXv8cZx1HvT7ZH
1XejcdzLBlMnJifH69VjYzrch3bHpRQl7tystI0YgjVIuTO58T/7SOADqYPo
0ZaufWRbS9HFJBragE1/RxUxe/Bxe/0/U++B4r3dRVGI5YjddGk8snguLa7+
82KTQ3KfjxZhurVedstmaCcuUqS5Z4TIT0hP5NVeip34RSdjycDDJcpJGYJq
tdG2jPKFZOxVCBTkX8ZWejoFzD73pWh5FD7jzkuoyPT7Xb+bOtEl4JFplPdX
hBQtr3diSv8uN29vGGYaZe2ROz7fgWLvdbSGRYY19I9z4eMh/HIKDU6myY4C
UOXfLK5SHHi8cSC55s3/u9FrhEHfMx1dMhm04K3cJm39w5mBY6MUN2M93V6K
x6k0c4qkPxd7Wif1BsjRdOQh7ByhRgfvslePxI2wqiZqNnGXhIxgfhEyzPc6
szp7lvpIS4vWUch2p70y2mCzh2+N1b7X6ivBS85ymTHWx1vs+uUgd98/P499
6wTe9kkMf1gk/4GVMJrpHoHNacKGtcAuWEE6tC7gFm/2Ah/Ybg45+MfOhPW8
mRvfs2cMtqbPsLD8EQNsX0wgOO0UMe8SRX82aX+8lbhibF91qWlsM6oQVREZ
sdqBk4D0TlCTMuSX91Oqe08LR//lPFELnuoaj+jUQ1e/xKbainCNN33y8V75
A1ZxrmiDJDfxm9MI+Gdh1ou9SKzeSF9KxCdp9hGiVhVukVZJiXiQ7rsVcwJ8
IYR8je8kUXfsntTDuxYrI+lukCcJR7Py5V24Vy19TvqNjBAwyL1HfA04bJbY
m2RsxnnFakpQ25WLWT6VKI2+gLZddQpNJ361Jk6Vkn1mTo/HNq9T3oiUrnWX
Jxq38uuJ4V0JoSQ+Bh9sIELWbyPJGJaNjmUdQOs9jNiQDK/+HAl6boe+uhcR
8coH3RUdd21vsazE4t7dHgZB3UsyyHEAn7B1Ip921eyIZToySSC8uJBhRWrP
9WXofBznAeyyx8IP3MvIsyixsKrvCdYZ4Fz3mjEB+GFmGa7P9JL3YrDxoZYp
rt/owxsDNn6cBWUFF2B7J7qhcxCiylHDILBe7bhkdUuq3XFvYBbnlkTFzIfv
oI7DDOgVWhfIIjP45kGK335dXHY3UFgkDXhB2qOGcEZ9L8UTWC8J7IOh374d
p5aIB7tTTt1y5+rZQxJrycXTQ0wJm5GNvcNAEbwlRU/F6T41SYbeuEICJ9Kk
/KMbJbChUpmZLnQsKRjKHJk2fawx5SfV3wTRV01NLZswSqkyonBf1peG4zNm
bXEKCmyJ0CoXEzTCHPNtsL+wDlGAAEtDvDxSgULCnC1hzvqZmJfyzQOv+f4z
n/+PemkeWDfcKB9vjAQA4iUE3bZcatU/5LGiNs/GATLXzi8/9jRtYMhuF+o/
sm1tqwpWkMwlB+c8wMiW44eiBAXQ5cuN9hpo4yMHcY2YBteRQ4grMU6c7IXM
BYBLoOPBxV3s3/9LIte+OZQG/UYEvfCSeNDsgfcNYC2v4aONaz0fPEft6gBe
sTBL1k+6gaVTBNEKfAu3g5FuRVAus3bsaBDR7BorqCDzsnxN8Uk3thRSX7rN
ZAA0Sr6QbpgwhkKZiSTn24opR5cqYOhsRd7CCXpKqT0RkybvigLtYYph/Exn
ZJS1GnwIAGfh3A2nWVIGos5P94BUCUNxcnYJuqsBPCic8E9tgy9ZMRm6YhpE
Jua1aLlqcSaVqRVJRU0VlZ+d1lXUkBo2kMR6kjp3pT82R7qa964jjdX9sqsB
Awqi0QcX3sAkxDUbNStAZRGEpBj7jbghhccbStu75De1cwBlJgPBAcLHy2ZW
qoBhZ1vVGEtUuByMWtXU/zZdOu1na4+ab+puiGSwLQbveo4AQyAhk62yuhj3
An5VdWTz/F+bvhLa7vKmehU4nsqU/6R8AC1NaNJMMpHoPOS7b8nT3ydaLwnf
x2xlU9DbGniFb3ZjfdmuQAXu3R0baaa0tjxypC5L2fh7b4f4SA3LWjVk+0Zv
TOCPLe8dyAEUuFOeMvMbvRWwAhmC1qIKvHEfgvZI7kkbIbruZ0QY1SNw4zlf
xv7R7OhIBKyLzIt4nrE/Qwul0wV3ZllWamkXfjMFRZ0E2X/bKksgZ8pHEUGG
dsKSpXa9VZxTKCKrdnFEh6W0/MvgbJIHZe1+R1rRldPGnPZg053ju0C4Zc35
uc0sK9bi/urC2vuRAJQ2eT/pDpwK7kCCmLJcLS5at9qMh0rlC3oxwgP+Bjxx
GN8UZMTELx+ZYQWlMkG4B3jSD8CQq4MUsSLUuNlz0dIv0T/iUO1OeNZzsmZl
tCJOtKbJ2MxF4QkknUVy5c5efT2eYhsYpJnX+VvAphh0WL+56JkhGcT02IkT
XSiQ+GSA5jqtW0yBZch7vN0rZhtJVEcn0mi2yXMePvSo6n8Vxnvt0EjXIsf9
Pg4qHiO+KyUvWhu8VBokMWDBksHYDKVqDO6WzyQW8QHasg9vDij5k1B4XWjf
2vDocNobT5A9hM6t9fN0EfO4yqFdqBcGWLOOaoYwSpcAOUftB+EEDsxV5UGY
nqNOYLbfnkLbQ5JP14ihCN54rcnvtufC3KzzfT6AUxkS8VH1m3NSIOq2Csip
hF9axL3k7NeYXwfN80uIrIZTvnAdlPCxE4q8zfjPp4Lab/y9QlYNCl+rDn8a
Hgm91WebYaAg0xsPnxanbYwSjJm3fhfRoDh6lWDWSOVfXZtHkJX58DKkN2yy
A95c7SHliyVXviPfcwcDJ0y7T3bdIwBdGySVLeFT3z9cG8hK1LrfwNUw2wYs
WC1SfFrVacmf9jtmpE/HJJ2fbjvrKUYTtqMpzl5Zh6LOWGmsEwGMb7CrdimN
90d4WJoatWlJuB+JXux7uCag2mCwGWm2GMmOKPDLjamP2MHCE7VFz7+4YhrE
ZymNZx4RQDMxXgmyoqmN2AE9zy2+Gex/K1kYCxwNL4MxjKA6U9q8IJXInKUc
Aci8dPza0V+/Kjrv5UjWr7EmsTZPqIAbjM8HYJwSEBO6GrZsh5ubNsbZ4lv/
lzx6/EkugVP/MjNmqctQcWbVQCwr+nxsEl60rgq/NP5V+6LeghCxshEu7FjA
0fLrVFlllDegeNH4T1c17IfmHicSGAqKDPa8lDfCFguR0fYk9NV9ZNoj63ac
LgCj45HDL7g2DZD7Pej5kuJBqyt8X+hlvO2OGn5okcwpQXhHRrlhHYBgf8/O
QFyRfE1EAAhf06/F6aVAraGxXS0SfJhmNoSVg1tF2g5xggBMNWeE/PJkuI2f
AoAx8B34m0MycXUBsuFrXzeaIMVe3qxgIe6W3Ytgz94KCocVftvYCDfDAzhc
G7lgnLuPSAfDFlO4BNX4cbvePb1+TaFRCKQb4DsIObQZD8/RKMh/Zqe6sMHX
s4jPDgVllprDMAbGpqRT0NnoQ3qVtIw04VDsDevHfJ6fty5gE1LcGqzo20vT
jzqEILijA3HAK0L+c9xU8W+0wNWLWj5VMV5T39JyhrQzFaJd+5IdwMldotGS
taecrrN1wTmaygkbpT58ABumvpoRZBr0ZrqyhJPyIbI/L/vQykMfr50JcrZi
Xp+/qk4/tfQ38zBhVn7oiqgDbFWFHFMsW1gDjw7jtcpTrsjch57CCTwSdJ40
pz1e4OJGFVlgwAYloi23WbRmhqM3BGAxcT3ZhLI6PscR3bPQgjAo0dOWaz8s
Fav66QzAulywmKUwI6hSDCSd+E8snQ4YTYq3GDDG8g0grPpoUSmHGEKHL3rK
YpMPnxyuzPz7Gj3Kz6oBXCRi33iQvdahBOeKVRXkTKcXRrqYT9lHLHM3wWk9
QvpfJvg7DkCWd3YZzKFBXMCSJKqBiDL7qmODCY2hpm3P03b3JEQaMWjyP1Ri
q8gKnkSdHx9DZZzRf+uojFw6bwVYrykXoLFTRoe866Rxk3uxRSal6RAEasxb
vTBJi8GqOT2Ud02qI4cBc8gpAalyjMDPu8/geqaO16C2aHnx5yVVL8FILFTA
493sIcH/AL8OZ/cBBpF/UkmYmgLpTn/UCUanRmIx/GJBgCJqqZKcaKN5DqSj
50hqlg6R0JfriKwtu26mVKFkrDBMnGbVSrogfGsWvZ1c4vBpqg3tMNjT6q9M
ZOI9vy8C6PAI1PGeLGfKQInADQqrwEixXc4kX1PFDWKCpnFzrP1r2556Jxj0
BxsX4+/22VYxdj5dgLa1+FobvHjiVIwf3bHXCfX+LXdrUWXXgDgJ7GLnAYxu
FF/Zb4qbk8zedsH+t+cDSc83ylq4IKUs6WAAi4lP0L1uZYrLPY980sU6M58G
TT3G6itEkMhlK/ZX5aHjx27hU2gYaOn01k12SFSo3SGTfQEJecf/h89w5Zxq
vAzORAiO1kp7b/RlZlUrVUzsFPs4Nj2E0rLp0HJPjjwmWQNRW943ITPBxWzu
mABHZpGolUmGRnxHeOxLWstRSNC58Pw8qlG1LRHB/iCatCwtd+kIZFHCZusq
VQZX91SrJcFV1+xCD4yiSIFs3N4SmVxTcFkTHJE1ZOgoInHwWRuDkkPeCVbT
EU8Doto9jWhjVb+Xp9jJw5Muj+24rFu5vCXzFbUoHY9S5FAPwc98HfcoeYZw
3SinYOFZuUyRsZxh8MSoZV9riOqxA4nBqORnIsYSAYLXWchnZNBWz8fK1s7j
ctxsG4jeZ9RvQZL/u0EAuIBNZhrIm1uDaPB0h7RmMUraK3CkwbDqJzt0To/c
uZAUOZh6weRmtSqmLZHszsK7SPOwWWhccjqyK3H7ov9edHFPQkaG5crUPX9V
vjPbENmCEUPlp35QtBGhRrsTm37paW9kS1o1nkW33LL9wHK0LN4ADaXg/HSc
Ng6p/UIijvxy3ngCSN7SKESVd2amXbwNJaS8eievkeR+HFO7+2FUEPrGoGr4
z8G4QqhWJ7eGvuO0vhTQ136kfJp5Nk+MlC18NJUNkSpUrtcMGwFsiAcC9OkU
tnjAuL5xcFpO04gBdkY+zyqMHYf/4sYwySIaXLHficz4Wq9GwSxsv45Aktyo
YIVaGV8ym3lKDH2sO1HieTcciPGcwEC8CKXROdyWV26aiUtq0e0tKWMOGp2k
PnujzpkrDCpAeudGexSs/UPCRsyASVQ8wRKtErjpKXtirn4MfT38v9jqILp0
2MYkgKzuvRc0j38/MOc+g5v6KCbWEjZ1iN4EUA3iWQAx5ZgZEo/a9q5nQuqv
oxlBXGAOq5lktFv1BolNlVLvSZzpVow0cxGbrGiF3ls+4+6hbGtv6DTVS3i6
Uuoe/Q9hR79WUMtfXmz8y66kk6LVt/p2lk7GGyScgl02tUlwpEUx51XjWn3d
u96T90Kvo+80L02Nc8fVSZz87eQzDHUfQmgjQTwRsNvb3wzwqPKAcjwezDpm
E7nizKbbwfCIouAZf4eM0CmHKxeddJgoOh3U+nzubXZL+Kk2O0AYlKnJpKS5
CohCRGlgI4f4jzrPSwiT/sjS+l/VgBKUbdQYcllNkfU6w0ug9UhaLeXBjK39
t/lMJGd5Bkq9IG0LVabrAact9GdMlU3cX49+bF0IO+kJm4IWOsx/oCtSqPju
75AitUMZQQ5KYl3drnZqK0DGQOaerUSQ2gY1JAvVA9YyahwdFqTB+lMkizz/
SfzS/EHfos0ZSKInJiCC1NvN1hdoW5hHht5mPPFDjCCAIw1VFgGCOI2PuNqp
xVt9EJPxK6IGQpHdokKtPId2G+jUVVGyW50LxpmuCiTnrOuWyC1qU77/icm+
DczblX5Ses1LV+TTnjCjBPjqqAIQ0UybzyNX9sMxYGXziJExB+Ef23Hv1iFR
PsztEtQ4ICk/qXGTUh5Yqv9nQKkhq8N2VqiidBeph+U12fUvS4fCFmIgDGhT
pwXbt0CQhIZvledXOsW0bdxVtGsaODjWPlhxcJfXV91LRWBeFx0p5FXjOvjY
m0rDN6DRYudtfOpo/vTzlbLn4KHGxiY4fJJSLWuMrBPEIcr7iszFaYiz0zzg
O+fqu1w+DUN2LFwnTJdQb7JlhTOPpk8ReuQseEhTLsvWIRPakLAhY2af8kuF
LonrmmIMncSnQRhuYLEjxddm4Flo3khOK1ZSvobziTADc6dGKFFWN1NAOjlC
C1DEXJM6hGIYGwE0byqfXFZKj3IJmbu6SGqGyYXv3CjyGKLry6b0bj72S6In
f8A9zLikhb6r7FugnN9AlStWkmYBaZb+VQPmLREihC4JaJA+uJ051yAAGHiW
89dfXhj5Feal7/xabDZTB6NBc82Z7bw2H2wLknSYxu7Sg4X3ePBdmKFwSfwO
Gr3GE3DUFcrOK0ZSBCsK+QFVlmUCZ7bE0OQU3t3g5hr0b8FoFlRFrOBafBz+
NlVJ/CewFSj/nxVeaf+9pRqXT8zIGABASO8ePQmbYjYMWB842WQhBpO3KvNn
fSBgs2K6ZrYWpq+bqg7a11atWvbnoNcdcZrNYyIPvaboB1K/pzDAgZ201kGG
bLy4MZdDki2jKkigF18L4buoHbnMIPT0uAWQqpXG8C4mPJrD1hrT894e5jzp
Ix2xmekycwvjkB81ZZenAof12ESkrApXVMk+CB/rrin8d8s8E+G23QBVi8Xg
WL9I5PLOPrikjyZnlYLqSkgss/12i1MLHbnwct08qHHo832BGAnWaYLaW16T
albIJiywXbq/dNPyycM3WHmph1yBrm+dsNurHjcGriZ9CLFfatxzoyFqUE3h
MNgId5W9HVmuDERUjOM6CUkyRRUopSnql3FnO0MtxhI3o+zb6ptNRat66EUr
V/9mULUeqqhFLenxtvREkPJYFFY9D1Oe4XxawDa9d/k9NTlQxi5JzYBf9Si7
qr7CXeU5L+WvC4pHacw5R1Xe0aCivYCfzblabwdYAwkwnxhVPbS5RLlBJlHL
3zrwQ32ekhaPUYcJeg6xqZz/tHo8swJlYGfXKpoeza3pn5dPDTh0hVMXyM9X
YuSVc9bZ3FZioSeUfHTv11zcbNUNoViygcosKxHLs/qYMiEHmzHNuQwK/4Kr
B5LMIqCyOKRBu8EaZ0Q3UupO1kyQ/Z3mI07wyvBZH4SsxDtFwYbdBkENjtNJ
5OtTA0E5rLbAvGpSqWKHYO8UUb/QU6KBoNaWPrTuyNa2xdInot47Jff2SP1A
MuaFmW4j0NbWL89+A8kl/Rp4AagGDi/YcPgOuMBd8jTHjcp8DLGc4Kcx/gf1
pWe5N0WgRkMwZI41heKAoa+moV/uZbtWxd2mO/5skzsOXBiZaNDDBUfTb1kg
FG4Pdtq5l9QGNlJ9hhvGV6scUSAG53gdZESpSBsE+rNK6mPh1PouV+q35gUn
k0R+tHOhHFRyrGC55Wpng7hxqTrweSE/SK+yuKOSmnUgo6ZKtmMOjT5tKtsn
ziOB3ufcIDrXtw/aiSm2TOHv/rhcL+BRhc2b3D3lw6G2WVG5ABFwsGpp0gHl
M4nQ5NDOZ3BDpQelAfLTI6gEdjNK2Y5AYLeEakZkxtFscLSeQ7P/QcLLEcPu
qquJ1ycDLidYHvT0iR5eCv+llJuUV8Ho1RUnpxYdvjXP4an5Ij/NBgyHqHNo
r3F5hmy9BP5Nw9SbnSfBz7hBrUUEvOhuIFRJb9qUvYdNpoxKI0shTKr5P4DY
J8U3qIYTBeJeM84536ORkb43DvPWQiSIaE4mG2bA4H/OMhqwLGEJ3KjU9B4n
5DXtGdb8zenaeXBL/mYr8Y2PqQ2ww/jTq/jusgtbEmxYOblq23D8Sl3B4KQ0
PTsj/GXd880xyXHRhJExWaTdLwM7Didn7LLKYQG2tC9qgQksVzEVeUoMOV2o
6fr2GP6nS6JjozaZmyujEixV5SegpIrg2ONywFyP7mPG4PA/NnJWZuW4mXul
k0BYh/jmlVAZqFYRdcrMAXEbdXsqrqRRchnGadKIaDaZ4E/PYEicrx2OZViB
JGx7kfcINQDEDCTDEzMS5tZm9cQE/S39a1wr3WJx1o8the9/W86Zi3RzGKmX
NjGLzC4c4epgfX6MqxBylIOhEF+yVAVw5kbqepng9NvVFCHk0prOnl4kq+D5
3U1vawuTWA/LNXEkoNFoV5GZn3+Cjp3m1Wh++uT8tvcSxx98qDVBNFPrqKro
NvMeSmZ1evC9jw5K1uDb+GkjfAZkuUBXJfA3LXZnHZyAuq9nqrK0Q7saC1c+
vS6VZ7+I2+tcnQVa0aQanxAD02ooRdU4zKQ74GC2+xN9ByyKiNnNbWmS6Olh
zm0aXxxajvS4PixAv0ciJU8bkDLlpmP81IoQUMxoHwmKtR9lE/vXd4+90oO1
5Q1SbVfO+XwoVI/B7bX2805X4HMmlc5FRTW1rCcH+qbiI8woh0ZVtJJ8xvpl
pY4YTJrVWeHBZR0VxvwrhPV8P++1nxpQwRXdmoGK67HMn18G9qOL6EcDOIty
ZB0LA35UXt0YEwREMeO1nr+5fYecH3GAR7R8ttVtarwwpQv2JysKX2M90041
VBA/V2Of0i9CXW5PKLzv/BRgvxBKJy0pCMqtxGYBp/hhaF6LstZJvlueArhu
QOCdiWIcBDR848b5H3E76VX6AajhCta6zeco9ViK8ivSzBSxYO+E9gzsgUxd
1Dx+RtG7biPm0ualdbk3gl2gXjN6+3+xgeWxc221UTzrQPCG/zEGE7pHDkbt
8ihb1FzGYBd+eyMWjFwXbPvXA73C4fajXAA0uiYYOxNbPSUOPt6BLyRpMhSh
Mbl+fGRx8uuZcKVJwUlUw1p1IksBble9lShS55DpNxh+vJrc6kqYxOTbejQ7
vc38F3TH1/FKH1OA+XocuyC8q/NGmaieInInEk/b2naLrzttRWgxm9gGO/Kc
RGjeTfg/ppPJLqkOAgKhPqr6dooqwuIin0rILn7SsVMFA8wqTO1sQbI5p7IN
CATb/Dk+J0caoCdO0/CX8aN3KTjUZvOZ1HDzLsvVLQhstA4Xv68+Ud3GLvK6
A0M17guo0lVtdzmCFXRCnQCDg0+y4ov+N//wew7/nCYLxOAtqbr9tq7Hre7c
ngv7w5vLxEP/47b/GqgcGH3y7zuENQKDIqH56FwhEDWE+Cs21OG57V9Z6Zjn
T6sTMFD6Q1t+5JiAjmVEPcNQqXRtkD4l5P2jF/nqiZnSEhIB5dwbSH/ws4n8
XcGOuK5IZIUYhFC4OokWn9zgKrU1EKjI6whauGR+VLurjBC6qvPJDkONy3z3
kBmrD4A+qwFCKijpVXTL5oQSBtw0nhZCnuLCzs3YPUP33vDF8PgHyXS5Bb1e
hOFb8U+boll9FwQqLDrBnWXW2PuqY0TYtnETzr8ZU0uoI30X+GSVCdf4iIW/
1vCOiPZVhupJSLsyIiVgqzW0fPRT+cJa4xuXTloSgw7Vz9K6Vp47BEaxGI6d
o7kunL+Rkbu7KM0LW0jq+hND4aX0W4KhLroHGvChA7uX3ESrkyz0Meho55KR
4CaUnjXBdPjLlX0OypIqqcyVeLfyMGcJzEGf85rI81NNWgd5sNH30xO6ciNu
WtBf3B7DncVUHFh8Ev0u011xW9B/2VgwvTlvnC9Tx3DoPfpWq/MMNU9tf0mq
Ra9G5uYK1mb7aN06sggvqmpgbCTl+En5JU3biAWKP+2aiG4GYwYjKn5abtlx
EnH0iVK7FqnEU1ZeHjrqlunbfMpIy0/zkpQTDjO8e1FWGXn3Ops4Di/6cnLW
SxpNCRMBZapSN218UWJCEVdJUw9TX7sppID7LsxS4RLdX14i8NshmpN3jzHO
2LV/fUmzBSy/X7mZGMUATuvS9348d45ndLgiiERHOU0NL9IH5Ly0/kTjlBON
Pgw/3+aO3UZA3X3XS5rsuP5BYLjxu3PAlO9ZgNoHr2cHLlSpWWQobr3V+zs8
7KXbX7AOEPV6S5cgbyBPSh4rtZlWM/vu2KE63tOWbsrc3HpPUbTkOZIeI2l/
kaksTDRHJ3JoVYEC0QNDA5/WRIuLYtqrYDqCEocUhh9/Hjb4XZZXwBG9qYwL
RU7MdGlwxoV/1JIM46XfBoKzi6sG2pqojenTmy2kpaGoivO7HCievFB0LVSQ
2rO44zm6xJ7adw8Z0yijsqgPX/d7h2n8ldX694srAaUE/CiisTgwzmtRHO+H
1vldWY5TuIpt9Ys6MSM4EnyeKcZNtdBKmB57iP+q2LVwA6Yc+4yBq7dNUvE/
HnXYibU9UE+iQbVJJnFKNLN7IOM7d/AVXjxtEfNxjMQsd7n61WYebpjKvFCA
EQnKWXA+8FdmdxV3Epm+DcKZ/hitCKKz8tc6b5T1E6d1F+PUfqpXti6bkiD2
91cG3FjUL3uj4eX0gOSTtTrIxSpaP3BQWayW7KSJ1+ZIMk3NLs8jHrq9JcYS
4oPcQUbKfTtScvBjC5KIXJaKffX649mtu/T9ezmOSzcjliEglCMC/FkJZPd5
KbXNHjtFZZkUc5VXf4Q0kEGeEthsJ0ONdSmrgh25fZcnPLseeF9Smi7PLe7C
0lqH7YzdCFO7hyjyEmrOLOaIYfRGogxQfaqmNB+QUvs1yMi2BjR5HjVLpRzL
kQNlctTHrE73UNBwmuxvTPGAuIyCb6LCicmNNNQ4/tgls+NiKu+oZbD3e7n2
4Rb5NFp02/ZroaO/SITQ4q2gYKNHaSugIiC+K0PewAAnzIKz/nb1RBYMpDAM
HIU1mtW+5ymEEhRHBwiEkygYyZf6c6b5q862XKrp77c1fz9A+rNZAaACWepK
Ny6SSf8+RXfnDBkLUQg0gqZ7RRY9KnfzbQKAR2Zk5UJtlDMwuXsciOxjLHeq
kr1FZMg48zk+PB4C5VNSckdJYMQflaCGJBmyVDqb2LgqWyU5bDekNRatAO9s
0FrW5fCwdlYuh/6pZUWjl6AUY9CRqswQtgfVFRRfwo7YeAsBXCn64FRCizy+
yPzyYXR/t7bz2rxxw6CMwPqHtwAjF6LHEVMDlDLfTXnhQC/Njy7G1Cg5yteX
957OVap9Db6Swy7Ocq8/8oLAs6uHANjDYLZb76mZoz58AghbDk6Pd14Aekje
tlslWAC0B9xobRUKksiBkPmT+vz1dRm0sbalcgpDGbCOIw8cI+viADh3oLjW
FmfRUcxu3sKOJsRtgni/YVeAN/CnOfNVd6Edbd445Fk6e5WLeUA01wW7EdsQ
RoAxv4TXa5JJvhwy4Qdwvz3HIB6bwcraaPqN6KB1lPlZZSmXavUyjRvUEc2u
v5C0OxEeuGyY6HQWeU6SLyHgt9U4u34gpR4xR4Zde7H4shUPOzD/Lqo9njub
3E+qttsLdEn47v55jardGIaM2aG6sR4Xz7p7jkmusO9B+Fi8owbILJH0M6Xe
c43DPdazOD378jS59Pnm0HfFjBFNktpzJYL/R/NkSUuHvA6eSNFIuBBk9wys
Q174S4QECHFlLfiXB8myYFlT/1dA0V8VTOwohzmWYrRUINhcGOu7rypLAOMy
M4KAxsRr/g/cwlO6NPhydygJZI2nGzSSMZCE68ZQdLYT9Uc/ExqrSAaOWCUM
/yUZk4OG0wE6QyBo4Rh4X+Q428O59WMJMwEJjrzJGsCAr4Gsp1p/q4kM5EzO
luwjcJv0E1Pb1LMkpyRFE2BxCqseUxAYGHgiLNileKcM06v67aD0UZG2WX7J
g3pAY+piVV1cqW4iP1eRkjoLhVsbpD2UsCPhGGdf5jYqSdvXIMX6ZbR4+2A4
Oy+8/WhSpNKzNX/0EhCvWuyFEiOzACu5/aFXg8KlqfYaX/DHCHcASENTEVT0
1D8BDErS4Rp0StnwLaUqQD9Os0rT/47y8FnlA4HBhE9jnA+iYMK5QUIga0nD
fNQ2LbHCfQ0CnCq5XlMccF5cmEeEbfijfvihcMEXVao5XD96XVFku2MITpwz
HniFgXvugGRD+T+qbDCeSH5n93pntQL+hzEKAxT7ZCeee6qvbWbFfU4O31TI
in8Qn6ikY0B+HzIkqypuVEvULqjcPMUthONJ5MWvpepNcScxSVliYp3Wb+5g
o+zV/savGuAVMM98LTiUBKT1Dqh6kuwbhJSunz9ijiF/OPTx33KRSR7LdH3u
BfTJSNLUJdbOb/VPJcS6Xqxv7pqgDW3K7Z3wgykmSp+coC5sZFgY49z0IORo
eRsMLSJmea/i1+/+aUO+iR640DvuiAchd34dt/NtkanOepom+TtCAjBAA2XE
yeOnKf4XQGRJZbtomqpGn54Y01JFxEQamnsxDwHqAg/PbTK5CdbRvZ+1ugvt
BtMCTkOX+fo58ss6THZtJ9iLZ3FUwnuLMksEm+m/DjhzvqHo/wffdJxUPvoD
NOWfqWzOdfb8ybmMHQ+69UVp62I+0qSjr4r1lmbCBIFVL/PZYIaWhhaItX3e
c6zFx0w9vzwo/7dbjYDKhW6G4iZXOV0WttsgBtEwI/Q4/RksAjnBzxt7CCD5
dc0vX2Cb7MYsuKpjywMwnqNUVs9TCD0VhZWf+XGVS4AS7i3nFoDae10vsAj/
nEdYveh5ov11Ytk2s+4vJ1f579Bb6L7MtcQ3gvJRNCqhYq5Ly0yOKOXlSdVw
OQF6cxl8lV9uxj3OLUNClUq3OVWHPSWy2OfAuPt0VFWOsvcQWZgPBZLEnF/X
zu4k5VrHZ1kbh01czr2dGm9u+AnVqAOAor8Ns6mB7oILOV+VCNsQ1zZrAGVF
sEQwgAP+XbCYob7nJ4wAqR+u0dOBvdJR3VAgdqDQGysmA1IkwsOwHUd6yMYp
ujPXY2htC77yQXivPS9mlyVMHQBqlcfBFGiSQo3IRH+sEQ/cH+Ol+RNyJ9qa
vV8k53BtbhYAif9cy/12prRrgy5sVSMJRgeGU/22dugovaAPnZBcu+BcjxtG
nMSG6ZencH227DKYw+njBf6vbZ5f8wUhbhetzFtLkwLwwfnf2XG/HX2tZp3C
FH0dRtSWfifbURkVX4sTClIlun3tMSxkbUNhv9IajywUjYDgj56Oosk1G2za
lrfpbMC/2mbZLYm7nI7m695VD2U8B2JgZrzCXyNbTDKLN8CTvU7E6y18TeQe
rQSBW9utubp7LD42HIl2fS/XLQDNBNjMOqYRoCGfDfjDRD2WtI0QT1EjFei+
rhVnNo8qo180SUr3OSl/xI5qul6UXheR6xaQPUzIu+B1evNWdLnHHXCAgS04
+s0ChHhm/sl123klq/1yUKx+B6skDRDRoK5xNVfEyHFUwqN4Egt0MvcorSdO
ajuwJthtd88sYd69usIoQCG6F2Ah1NUxLtFOESLwuWHCfp21JEoUPiIrCeZ1
Is2SBJSRoqc4INPH8f0ktPbjg+uv2LU2JrOLOCzXHUmFescXy+j4eMoT1iyB
OnGMkelKu24KV+i3aPd0MRvHLSPqKG7QjKoUAWCzVxiUPgjgVVe3bk+Qs0D4
eEONP2BPt4EZ0xSS/hGSe+U7SraHvGILJj+M26dqZH6e9BByCUP3jPUlBERl
l7lMxXoqi1TPL/WIOb55xj7RLhz3i5MyfG0fUwiAT9bFcduzjWapKgH7zkmc
9pcIb3H/vctztE/NT5xgpWM2RdKdACivcJWaMIX+EJG7zEPSnryiF5WtOBEK
E6gzxogvF6y3pBTlwHvJgRj54eqBDHdlzB1NesOM7m6e6StxiwSjkdNu9lJr
+pDzpua8StE1HdQZFXvglYElf8WpsG3D6ms+1TvbXY8qoB61dnSCnxcYQpsb
rFQ4oll+qP+ouyBiLDmCtMgtFLXgQM//+9iOQvDVbAdCRCrhtIWVKKTePQvl
hGD4Eamic5Zlvk5G0J1OMcyQHsXkikJZT9QV8Zgg68KN/QytFJk5ebEP/kCb
ZA7Do7PXWB0B0sRpEFgWV+TzOx29lyZMpiP71asW+9CM2yWPlkk6ysx/QxW4
lKOPxYYWyCiSacTCF6CCxFUQJPigEuKuCybc0lBS1VySIpxMti2M3GLAt2is
Ksw83KhlWsmvFQ9dmkqWs/SZos1nrLXUP1v7X1OZO5z+N7B6MuF9iyI3CVLg
w9Lk1PZGdHq9Q6hwdZY0VxrGM9qGQXLAoUBLClKKw4YJoB5xGB8e6gTDraJ8
36WR042iIfwheaok2YDK6H1kXsLQUkighmYVYFPywybx6Va42B0T/+B7Nju8
LFVHFt22A9zS0u2ZxfTdoXzhtj/CyzOyExX49fALidgsCPYlZ0/1o+k8zRUq
dgXg2L0nPw0fqZOEPyKEOci+7lo5qUCHSpUBmFLIM2Z1eouh9dM3M+EieCz3
Q//f0GOEUagT839pVZkaRT0s1GeZ+Soi2KT8P6Q/BgPlNWD+U8eDs+ZBD5DO
tjNYg+A7tUH4H/iNhpAfuFmi0xlItGRuNCJ1y7rg9vrS0fONV4+HJ0X3gZ+6
i5r1aAmwyCtYcUW+D3TUhv7touOXUNhXHApPAnd+/iaOdH8OR5QCOp5/WK2f
vdDwMrdxEXiY5tE180w13Y11/J4oLho3mjP7kqyptwiqDQzlq8MruKXXOFEs
Yq+nv567MZ/AYwGabkubsgpfKin31iFd/p/UKG/1t1fvfQeQgpjzbCk2IYgg
a3vzitfKjIuK99ZrUfdypdcRuf1tp7JqGsJc3EJ4R5ZjG5fLf8zY1ruG8gHn
1traa3R+gYQ8r4JRTdi9JYu5ctC349Kjsnt0JIaubx7Er5XVkJYrhoRrnhXv
PGCQb8aiNFnfpmFJL/ersdgidGhIfJzfTCL4K1KxwoceaqCyNMryAtqCzlh3
bBIgYw1eO+iIuunEnKbhd66e1gl6BHRLXcjnGWqVeaPjLm31M1UEHeVSccD8
TooyN/d9bjNObxF+GGoDCObsUBTiQJvHrH/vxx9vNRtdWowvp+winZYhZeoi
OGG/JiW9jbyox9hrESo4bq+zY96fiyrefoCXFpYk8CM98okzb5BGRacUC8lU
E0sHKFM6zgHQJPjGdTM+vgGxPl4Zk5lVwh2HmFpZtT4bYNVJ7A7hIdlc/U0w
vcFdfcnCrZ6Mctm1+XvmcarMAEYh2GWR0BYGpkgWUQMOPYEF+uqK8kVTTmHY
r6NrrNeOe/yxS2+W0oDz/ySBfkFgBZDICB+QALMHvVwgBSFA92QBUq+EQRJy
l97XgPTc6hS5jKZsoTfZe8828Sv2lkw8Gm9zxHTicjD5XKsSarSUe25ScRLw
C9ai3F5AUBL/BSvk3BjrU9TUiqhaCxHUpaKkT/MuWVbtDvvjSDqJT6ZfHYsO
plcLcYycALd3TEZFW886HuULAmaPskP8bqZGgqQO5hTkAfto/vwdGhbu5vzr
e1+GRGjTvLALSiiHRxaapDum1heYkYiUdKGXvsG/YUT0hUdgafuufmLI0jtj
vPVmePUrHFs2JFXXX1amJfmJ/u7d4T9WnukjWeZ1VhYkqj8ijqMsxKcfni+8
rvRLfTmi80RQkWMFvqfw8BbapliQNun/gEZE82xeVmlT7siPmNG/rMpCZFzi
MGfxX9r6l7CybabfOttk1ZnZHTRE+3t1Jey3GlllO7iq2x2vfZ20YiOYEmm7
R5THNZzYTYc4DT4/0o2z5inwPNUDmR8jb7lw/Y9fdm9wkWSKrhFORzeqkY3n
wcsPt95jtO8YWzMsjYiz982u3rnjoXWF+jIMBp5vVzBVQ74L58culu23x694
Q9hqJzk+qsPw9FSi7/sGsqdAIYdBfkf+9SYVHQgBdGmOGFobnOg4cKbn02vM
ZUvCGIMormLlba24v6kXEHgjJO2lTO26AkOkpHhxuKmvLh8cN1nnSx6V74KD
fFF7Mtd5mZCLhg/1yFgYnHYT41xiKsSlmEcw2WrhTxHQXOaGYWy3ZW7aO5v9
OLOzenX1NlipFIQknFAVRQ0X/tqH2UadLVSQuCBnFY9+71ZnM/o/+8SwmMGh
xZXOGUl84nE9e1n4aFaS/6wLmWMkKD2ZYBI7VNnx7+gfO/O2IfJNqow2imZ7
AZyj0ySwAIOATugwz6BeJ63rH8XvEtNUv7wlDRB01oKuYzVYQGmIVf2h0ufl
YyGkFC+LhLAMpmiGAjsMSyOTM8KuQMqgS0rksfTeWBZ5u7dV6VTdZEUmofRD
YKiqeG7b56iI+d6XZ4oQgOkwvX/393NaqELcGL16TFpCw+egNQfhS3F+QL6m
jGTjmqbiyQUUH+9byX5adzJjK4a35oGfDLoVkwPZ1aZKC+VTfDV5sFiv7CGx
BzSi53ny2l/mtEq2ODtEBb7tkAxvCQ2e/VTEJjuMQXWcsBjjOuwc37tiHIhw
C3JTxYJGnGFrV53L8yxLF8BvYr6qEXvulTd3N0RIvHfuykWUu4hdXLF0ETKS
vZk9RjSghyqKBuGciNPICXY+4pZI76VBAxyN8YqSA/YmSdDI9T3v2e8A8e4p
whKHNRbixs2m/QQ/3duXyvxkWbZOWhEHLPitfe7TKnGerxuDZyWMB8axsqhL
Ro9M/9ESZTrsJOGQZecr1b5/tu7MwZp/ZHeWsJpjH7kUyjmrUiPSlRpS2mko
Q0BFxKbTOKmORITBqgeCBkJOY3mduE5pSEBec+bZ/f9FEl5IyC287YForUd+
jTwzPLHXd8dX1ikstpUOCDxoLfXRjHdaxMe32ngjlmSAQvyxCSCDab0Ff5Zt
CYdR/uhuoRldfmtrPOok+6ZiH/MhlMLy5pvlFEEKGm5aiJRYECtNPwTCPrBD
Wc7j8tE/gQtpsgalKQ7r3s5cZiXOgQckmin3eKq4qJoLhrB+DEcRJssxEED9
M8GGHW6lVl/fz0Y/fwk9o8PQ9pwvxvITAW/nibesZBs/S2c7oiff7FjO2ZgZ
RSyd8zeO/xA4LoXlDAJPN44ClNdsYlVK7q2yArmZejKNU2Qz8/WQqTKifoog
rFaNK4YJXiSWHPsvUn2+qtR8oL+HoBUWGWDDO6/XbEoE+r6bkQ3I4X5TYcgZ
v48pwAch508Of99fUWK1NE/0jEYVpzlZxgyQOF0sZh833Z3A6DQ1m9lco4+y
QgKYs3Nvj/G189QFPP7FB0dNYqneQCo7g1/+QbvofE8ZQICityOiL7Uu3fJq
04ORYcg9GiV+VSkEjOzgFkwLmSfpVVGc2eD8YR0fF09MNV2h4+Qs2Wa0RKpu
Qu/8X3ySiaq60AdRbXnp2GhmikFbYzh+g9WuV+tlhaVcUFdY3SFCBzHhK0r0
wFxvso6SloPdyfTz2u7BaFLEjKWwXSWelYku2AipXLOzfeixouTIYIOJlF3m
qlACMmelKP2Bt0k/vjMLVZ8fn7xejoJpTzU1wPT1wzcy39CwAoK+0zYVgzT3
AWDMZGBgTxAMTf9TJbECbIldcq4sv3yXPwsAcHqZaDGhzal+AvzNNt0/APNR
WwjW+wrFL2XMKoW65jUqDYHGKLK23oEnRAkgQyVbao/23sis+1mSD78xYThI
aTeBMmV2ZZxdGiR2HRFivoMKwn2CRYH2Btk9TRXm02WzSBR6KUa+1CNp26ns
tn/p3MgpzqobO8zyn9+rFirb8ulTkg/Mk4KkIUKmlRRkJhzO5ujI00ypf0xR
NyJPRKoA79Yjv7Gi+Q9wz2PXPcBjvvz/cx4TLtHpDRmHFqtx1fP9NO1JFM09
OxlidnywxP5Rrj++nJq0d4kc7kO1qrEI1v9TELMXCFtWxBY3WRUmUiLpFoyO
vW7PeW3UuMUfQj1e38t9EkNPfB46qSRRGSBoisZT/CvnuYThnfJmdWiXhM+a
fYH48FXwH19bIKo8zn+zxee9yBOcRAYYwdHaBEs4+qtNrZrIOe+6KOA19jxi
hpNlpB09JScNoOEblEYdgiFOww7D0vb67JbfOZrv3QUk8FLr05ZtMR7CpzxD
2rtgKlsLIlgIO7tDyqCL0AgrgcUsJcWNIQ2v6RXeaUDMcD31ZnooSJ0zfwsL
wl3alGQpMTzy7B5Y7Jfa9H8gO2MVwuMT09rlPrIFnsF7F4YDnodjpqCqIg6t
nwknTa7ZrVnQ77TVHrje2gm75L9LLwos/0nYRjeV6dvDpBsOjQZnNMB9z8RJ
MyEP1UyguV9eaFpR69AWfhYIRGKyP1nJsYGZJBv9kJUlzwSBGvc2ihZiDiXw
MBjyTo9PaB3XDfF55rXUKldZESKaegfMRvf2Itv1B74gLDINFPrTEDgrukBD
Au0LS3QKNTuYMXSs3+y2DIRay3vdCp/Bd0H1q75kaSnAgBwvl4WMv8C5Ab2Z
0ELiLSN1Pxx8a7jsGnaDzkgPuZH5/rfpc6iTF7j0kyaqxUtjzt81o/c19uyE
WzIYaMlKNUHGbJtybPrLLDXnadT0poUPSBiKjz9/KI6wtNB0Ya1tGq8eltZ4
AyJdc0/mdrVDaJHal+AHoOvr8JxJYCPnN18Bl5pn6AtYpR2hTEcHY/87GVe8
j9mKFMiQ/ac9fVrRlGTVxNIY1qmZmC5/fyGv/UiI1snsxqwiTVay58aiMSJ+
TW0hT098aMkw/m7a4ZtQvXQvVzpm0EponzUih4rpshnXL1deGHe+cdxQCdzt
x8z7aZJoLHqXR5gkQ92MQP7VQsFTDyKa4vJNuBj2OO8dKpiMYN80HU0v8zJ5
DvxCLcaWQdSQU6jeRMFTYIPSPfi9VuiMZ5e1dQbphtqBLhL/cdNFboCfAsd7
G99wbpBJG0jW6/za0f+1h7cZo+2+4MtIRHctcCIXuB/PzkHKUPqg+RArjquC
k7RPXD7mIu7jQFxm8ttTgi7GG6f9mvEilyLBCIDsL0Vrv3N5hH69tAPzY0aw
zE9f4wjXjSbREneYJGDoygnS5n8qBNL6K1FGTpcW3SiVQ8uMnUbmOymvDR/G
l3ouCrfDNgKryRdCZntuQEQriBFtMJO7bOwC6o5DntLqAdRrzyOFq+ShK/p+
OaIHNvzIgXDTSkykdNtopCEB9IPm6Nt3ibz8N3XcwLDZHcY3LZeOHM05RvAl
19HwZA2uGAtmT+keqhOAna2OIj2UfKxuc6no8zgcy9I/+I789WP2M9u0NaAw
DaXm1YhTs3CelYH6TcMUt/do/Vx3IEjzk/UZTH13gIrrnaIl8BK9OP+LbnNP
sEJ5rGaO3ByyxrrujZyITH9M44mLxtzf2k+2tJjJ1Z1CMcTln+Hh3f5tIR9g
6/797cVQ4F1gFUT1OHzKKPrtMhGI0c2/Km2sIdgMNCE2PRYjbVUOiToNwdWZ
okDgL8PgaYsFFiQM1m5FJNx1aqnmNE6qom6dy4djNZxYLx+ju3iP5EDRJeVs
Wx+KCkb9FpN/hZfoI+nLxxAjhrRacpvmC59EzDkBvfdMWOv1uXHJbJUfPY2Z
2/zXV13/7fEICrm9N/6i3mmif/XsV8tlZTdag0jb/WEF3OUiM7XPVtIsaFIC
e0VUzwjR+Z2N1vackPKrtgf16Jr/KUA0U6oP0cyFFrSHQb6N/q+8j4hVUnwf
4SIQxiE/L3irIxs4NKRBist8jzBbLsRcK0c7ArUM31aiaWR/0KuC3kvQ/+lJ
Em6BoBeN31jHE1LzwRE6IGJ7DCMq47uV9B/tN9kBACb6f5g/n53sMz7PPdBa
ztF69ntZBgqouNp5MIgN6ibYQCjVWQJ1hXyXbNCTRbPzwraRN7YBnA8u9nFN
Xqt69e9ghKoJ2qv3EB81kFa4rT8NezRy/BzOYpoa0ni1qfWEdAgu7Lfd2QOM
Twkdtx5iuQamU0ST/Bg88yW9LaAlAZKR7/2DS4h4sUOQ5lH9RyUcFhuOo8L0
b6CNlKP6YvxZfn8wFkj72q1aJPCd6X/MqxxIClSayDh65Kd5DkGGjkstD4ps
cNU8DwiZH0UifW4Cg6nxQ4LuA4pJbVdzWncOG5RZxwEVJrtT3JzH4DWmXIqY
1JpBzdlBZZ4LcyTDfluIlh5O8SaNuaUwYEkA8BZ+Sg5q0dwjhB0v78G5I+lT
bFArdgc6/gdbXl/p9yvmE3vi45wCFioQD1KTGQjspLN20mBud+2fuUWDxi3+
vKRu8TUIdkEw4Lm5LN401Q3HG7Ad4hjHcyFUigtkOELJodj1qR0RgMNl5X+M
Yw5iuV6D0OyJaolcAQksrAhMpURLtK7NzbQcFEmiEPhLibMxQs75n6IAmjE4
Obl9BYhvuMytnZrCVDDHSTAXb8mD6K9LpgkVWw6lin4T+8iDBuRt8OambgfN
wHDda/npCfNBeqNWUpcp0PwMJWwfSuK712Hrk9RazVMDuJbIs7UPJctQ/fsW
3PrecwKueiMpYq8tw0xVe3l1BDWbfxBVqLdobTT/k3q/ISKt1OSRLpLHMwwX
9kB/igBD68PH5MqMmFCBH0J4yZEluF0vGwRcs5pgx2vTC6+Sxyb6C6NTyrFl
7yyoNz8S/fGGhuiUuobLdYu2VJRc0P+YzMnjXDOGLbOw0WS4UrUhJvRCJCez
SJgAuplL1uOLqU+ZEeIocmGbbPanYnavmz/KPkXeEoaBJWHpXUGgiyTZn/S8
HkeV4+D4rcvW7hBJMb9qQToMTBXzLxnjI7dnelrPmbpMUdlF6wsKpPIJTKP4
KAf/DgHPdgwZhEMfLrTwBcH444JdonmwzFznFYga/xUJkcE+DITZwI/611TD
hZvb4L0yACgl5r87pOz2H+lqEcD1pmkgdo5zanexcvEgwWXerfRooAUvhB9Y
Z1hR+PUbQVLhDdbUltyhZu78FqAlWVpaJMMFS5Uz2mNzr8MhfuiXsMAYPSo2
JB3xU7xPc3OH7hiTAfDrmNjADvckiaUDUVrV71NR3vRyxExiiGCgUXm3DP6N
/6NVBQuS9YGKC1AHCyD9R2ulrPWvUbQFFq65+z2QGWXhwbCv8osHcG/K0J2z
E/Q400O2OchxY5ZStryrOfd9o7g+ydQ9/QstvO2hXeqV0j7013JvPTk8rYC6
XXuTY0IKQBTQPmC4UPUPHkkSmv808G+0dMGaaG4shSxwed7Yr3dmMSAqZ2Rv
fyoIsgmuwB1chjcaOlZ4Jbb9vFzVs/0NjTfLLeuQww1F4n5LxXj5tUmQhQA/
OyYiYTleApneNCGw773wDo5FTD2YITJR5BXimQwALgpaFTyhr+kKFqZxii9p
7WnsgupdIaHC9I3PBAzKDHXvbYvH+Gm1+tmEek48t5CD2wn6+wosR10c/b0G
iW7TcWz04c1NvdSxK+bYot5P512Aq46cdmEvx3SJtXdf8+qfDb8jliF+qOK4
b+8NAZvZ5ddpSXmGoQJ7BQkoS7HwQL72OmCxkfgT4zdGlplcnHuGfoD7IeKk
Ri1W+/ThHdK8XV17zd26ST6BFh1hw0gBLO25i67VPnhhQHCMGz4G854iq22x
7gtkrl7rq5dyv/c7E9WMOdwmjZq1VbrmAafCl9uL6kzgzbNcAbG+Ssk5wdcL
wievjLBSEr+SlZ3wfLZTztQvEGDBBDEGwRO3hV0/5bTWMDiNfkDxiOOkkmvr
9Jqa0LCOstU1Yh2aifRuqIUimQ585vTmb64Al+xUjTwvItvBQYRb6Gf0nk2B
EOkTL318/vmxw2BNAx+8Nk/zVnpIa6OoR110IPYeJc9Ji9kPF1Ozz34/rtgl
MrQP3JFRe8TV3uB9/P93oVy2tNXDrxPDP0ac+sp6/B2zI44dgdsjJHnljAaV
28gcKm0PRow9bcLXlQJ/6ux+aElPEAi/vZpbhZTPJjaaYzeAlmeN2TxU9rCO
D+Z7J9dVQ4Dd3IXNKZO+4ejGVPIY0TFgWRc8UowFzcOT8vssFxuhSKEmG5dR
mgMHk7MpcZp7U9ESSuElHscyHqCQzK771pn/I8Fab018RMWSb1qNEBL4ZDDt
eKJVupxtoYyWIscX+KOz4/aDq1MXg12DvfRqL2tkl5CqZqJi6NPXvDgT879e
JqETkxyRODQLbkTfXXGL6m03heSA+arYXUU4iBsATWE7t/0mhgOew07UFGoO
07ymehCvkdE174/9BLxCDlhTLTOWyG89PV4gczECrbZLKQol2LoUwLkf4sA9
TKGgcgaRc5IA/+v4xsuJGri6jWpfXiHCY4Zeg01YjgtGKcz/IH+6wCcI8Dyu
PXMQcTeMXYNlkROQqHCfwuirzEwuFDpKqyax/CdKxi6eG11su5aAZu7J2c+K
bU/ykKcJ8uuV4hllkkBsKkEb9346AtPJT8lz/t+1BGvqrRgl0/hZtZzzdFKS
KPlhWhgYrgtueSjK9mzT+YZ0jUJG0c9ZGmN0JQhJLlqu9l7zR8IS6MdX8UCV
zKTXNLKmDLYZwxilUb4bJGZp2umdfGfLqvzA96XirH/KVzP27h+XZBiznRUN
D0qtXxEtWY7qK4qPVKKle+nXM0rK+H68imzAqhIj0S+9awgSpJo6GmuK5AWv
obDv6LYeLbfbKlWqdW357RMdramOgw4E1tDMLA7vYU7P/TSyX6eEw5nC774b
ZQ+kT8q36NhOOwlsJ176d5SUwL9T7h62rS2Kde7vnrcjavcgUZOqck+TfzLx
6EF/masD6jhlDsH02hXVXlLdpctYxfp34G7WFNp3Nu3/3qeFF/Cl8QrJQuQu
h+2fDtgsQppbRGSQsA/VUtRvK8FMfV8zXzfj1bFDJva/FBttsmTYH9JZSjnu
Tp3O0pRkifQYvFEs2+SyYzAnZZ/gsAilj/nYvKXMeEyA9iGjJq8cMRJNCS66
a9Ic7axAyE7wc1lcvZ3X6sbGo3jvoKexdhEN90ymG3vTIRa8Bpa3lQuTt4JQ
KCdmnVAH/DnlFVy1J/xHRKpQwRscavvPOFNZ8IlrJ+RCy3w2byREEmEhb0NL
fBvAKp0ENZJ0nNTzIm364HxFZbCDGR8GkOj10OdDb8T6Z9gXKJosb9l3tUxY
DfcIe6cTN1dzMgdCX8LCKWW7WBLvhLGHppMzieCh6SyF3Xz0kfmt8l1w0LXq
0m1LmVV6GzWrV8w6RCO9+KydkQ4r/j7kR/5SvXK753LbKrmqnrRWs/Q5gimH
qQWfcxEfXOshXx5lILjma+QGhNqgth6MxwKGHrVJ8rn5J0Feht+G5oUZ0qX6
/xo1FaYMtkdpR9P02ieJy9kiAKY/xemFkdoznfWFgOgDXn5pf3U24GkjqEzY
C+MSRLg1ZzKs8l2GZoYL2Zh0YNz0UFELh39eUGtibbRDGRcz5VBbxZT0+O0s
7rXrwCRbL59dEU/hsV5dlZq6gNL22B4aKHzqelSDn9pxGwQIZGGmMJXRUll2
kcbNGAlrFZQY1blnGPBui+IoYv8R2nM6dKU2jyByqHg/e4J07FO3ctEQ6bQ5
z0b2Mvs6AWe/4qBV68xU8p6A9sySQc4eePsXYQRew7K1tB7NNxtfmk4IubZF
elCfI2NXc1T+FxoJhfFarE9dia7ooN0Yd1a0NQKeCU2n9GJrlRSPXk5Acepe
70TFu94f5KSMPNfOJay6gk/xW0osqCDZnLHPmb9capPe1H1Nc1R/z7zxuIbi
Eq4kAnoO2ym54QCiqrlJfbMHF1AUg6eshW9dg9CIH2jiq64XxrgArTdlmfnf
KFZjzhmSnU5iOdUzv7B+igmJ68K69YAZ8UpWjh1N92T441pDNMCmpKsLg08K
4weHhhKMPi3O+UZ9ULdK8wsgNDtkZavBB+LI7cNaHNSCjZWo9z/FRzoWv52T
r9tliiRwwhBoSSmSzGPPkdzO3l+glRWnRVSv9WA+YPXOg1e1gqzIG4Rlgbt/
eugiMcQdMqcS3trx9neuIFWWYOvMIaJhPkIdhcxR2AsTeRY+N8IC7Voi9d2h
K9u8Q/oOcmv0xUQQ4WJFPJR0FuEp5E9Q9TZ7DtGe3DxBEU+wtnyTQgcOo4wf
mMDyIkq8rvDPebZgaZ3gONdbKh+9ApKmSGKjLgPi3OE1jpZ/Crc00aK5ovam
5ZrZgVgXrXNILopr1UUMicnWSj7mczWSr2Kfa0j+kCIuL4AQuxZR3stWA+bt
JbcotayqFlf1NcLtOrL9HcVWlOLJhr+mrp/uDIG6zpQEDP2llRhxKIocgq4q
XTKN6MFbgDEAlAjmGN1gSvmZnfop69A7Lg5NjzOBe6kZ9SIYsN3N5pihAlGm
Ip2wI5UNz6VuwRw7aBxLIui4F+/ibIB2YvtFyF2v+z95BURsv06CmtxFONT7
ZdHPxV+IB6G3i9eocDfM9unug9fi2hyQxlFVGzuuaExq5gDgpeUuFlgcG2a7
SDxOHndjcGPd1CAUKsgPnw1iNTG8VoKaUNRIVQt9cwkYtadYZa30n/Gofe27
+wYS62wkyGxbokXtaX6yol4tTp2lWxDOZYYI6kxehh8i6njIxQJx/pz9q1e7
C7LxH/SJ6Py5ej+IyTQqNFxX50GLcOBDzGYK/6Ml4IyAv5+IOkoxFkuGTWXE
hfFsHyZzQk2hLaL8srOPeCXHdUp+hJPPYXOFrKlkkE9mC1f3h5GcAUeJynyX
PZp35HcQPOUcTWIcMKPIv5t9aD2Jf/imN5SlbrH1QUm0xKKTgPeb0W2Z3ziP
SW9XsdH+q5MnK2Lle1nLxJhH5o1Soig5idP2KA/yjaWHbEswgmOJlXPNgLms
fAw7cZNXU5eGls/t227XgTQKWZYkZJDQyMLVEoMEM65AgAnOWxntS1xwq7ay
Rws81BaoCrPS+C4MEezQgHi92TGm3HfGHWReuFxGy260Ioaygj2tiuMKENMU
8FprQfEb0Jgkzl1UTanTxe8sdjGNrwn456fZ+o9yFIXCiS9erLW5YVXE1HJg
HopNdw3iJMi3a9cQ7k+AOCYLPn0MNxi0ksy+4eCQwBVRcuGw5cgKFR7Um8z0
OjC/Pc66zwnu8/nfazo+onTtY/KwxjvpNrhv+IcG1e6qaVsBFnqByMmBqEv0
dpsTiTW4Tg83svHaZaIpytBdd0Ox9yKz/TvXWlXuZDS1WP/FkehS4zQT2Zz1
G7IAdWNpCrepz9IW7NDgg8kkfNCJmwiwN2zqJdS7XPxVbd00GrnR8jgJfgxg
mYjcQuzRA/flN/hn61Zkg8IlWmBp3aG8sDquCG22yY+YhTdmjX5mCXOnIst1
vBYubzqaViQGqVmGVvg4d8G2cFVCp2BSVvzbegfLey3C4rP9mlzClLyd8vtt
LpFHa/92jdvErsJ7s6mkDlHUdAcZFltdSMTWZ4D1iybGCx6sqNOR/tCXp5J9
HEMJ4v2+VPzzknwKU9CvfqHa7HwWI9aKrakQaBJMM7RbWEE4zRHTEHOCWbur
QrwxKkoGrcdSdMTt4lgzzKiuK1/YBpw7ppAlSQvVCmQrH4t3RJHPYB6DLxWf
28MTj8ImPwlkRkVijg4B5MYemRDgl/FmNJUpFIosYYMPAVgeSQAecjhIt/EG
NCKO0v9o6NC1bM5bvlZSDLtxIqvJmQadftKZynSEfIrBmHVaXSbtCBnABzYf
qxt5knptPwpkGl2S2d/v0aJFgf9feoQpGv+QjLIo2unR/Mjujl+j82DCicMs
V5DF4QbSyK6NPdk2e9B9MjukHiLWKVpqBDJInWDlJEdpPxxjdxLe72dp+sWH
B1YWVT0ziaA2ZAfc0k0KDcVahjAmivHsvBxuzsQrQX44KIh4AItYS2SI60ij
HimmX1ruzvoKkYwvTWoC5p4CwukijY+LCS8GflUjgPGOdipIkwV4sXX3x5wx
vyHIGTAQmbLsGNPZ6jeIGGPHpUvFmJ21D/XiVlCGrnq0kJ/RFuLRiQY3gxZr
T6ueT/DNy5ACAb5f7f8K96pCiy4Dv+nie3Rv5uSIRS2t6groXaBgImMnwIs3
rOdneSSQjLVACxYenwIbAECCK+EBQZLouPFUuDd/xqo8b/8CrF99WkmQP8Gc
bNUlgCjNi0myaJrHHMCfNYO4UqFTzGPEi+u5d+V3IVRqzmoJg6eKZoo6dAbh
nabkCkXTRKkkc9c/FybX6H3JuEUDDPH8pBo2inZCeN7SZoO0BxQykNZOwjNP
Rg6zY/9BRGc1IYcobEiT2AOUNJhhKlB4bnX2ONQ2S+DINAIA+M8gYjNp6vyM
QDqkxiSHIwHrmKneSk+F8qrXPnQtZyKF4qBQhgHQOcKraTDFY0adEidd5yTG
LfkLXZFtrVvMZ9e+YWhD48UPiCsAPcUv4uxvwLWGKAQxtZESF/nXnHDh75v4
7QvoNV3jLodXWd83d+FnrgOoGilH1nFtkYgfKkYh6wrEiqkOxt/sHm1LJQ0x
GXWWjc6CSwhdPYILO29iCXStQJVKEPf64OdQnhVDFJooDexZbs2VLNS/8ev6
Se06WZPVezdIWwzKpkoxnv1TDGcRc6Cd04JOOYlOCCSe3PZm1H1X+qq89XNR
uJQKDeM4mLAeScgJDt0HWiFt/g/WJ5AX50CJeHCw9iokt/9SCwYzZEfsyEwR
PKUANOw/l89CjP74m82VMmGbPiPXwtaHYQzsp7aWfLiziki2Fcvg6UK64IkE
zu5WgjREuHWDJDSNcgEg5R1r4D6zaEuO3x6aCJL5CmDKQBwsVrIY15jowXjz
qmdTpjed/KigWIrG01FfIIzXAZM6FniY5tJE8GHl1ToAxVlZVkXKqjd2qRnd
yCqmOZcGJYc5yLiJiESRa4LMI6drxr7bUGgcrnfkyZ0PLYql1ddmr1jBGQLK
8UJlVa8k0gi8rlJ844l08+hv/DLBCUaRr4dyRRZbCFiqQsdkxU1XvfxXjzU+
WaLOnVVPZsUbXEVnV6cHytE3Y1cV6hTA7EwL0XrIKtPjSwKnhqq3x4PmCD2+
XWP00W1m/M75Di0RMJczfGJtHTbg/Cc1R9cry/7SZFcu96QFS5aXVKXnuSLy
gU1i7JyIyeZUqv2EesXVRy5EujhQCJXbd66myhMwNJ+oqTkVTL3qTvgnITpO
gPwJHDhUWQaM0BVFM0mPQFtRTlFZr+4IS5DN2YKjrxQ96XIi8pY2FcaLnqVh
jamPuUiT4jO6zH0uq+ZNfsQY2b3ELJO44lr3mfDW9f/ELZ1CVyZp2KwAu0XW
Tm0gQo575Tczm5edOR8z/CLOJu5taMcYBM2cvwlh+wGanSlff12Pupxb2vkL
2KLcil89zUrKxvfFMP+9m2ufIVbuiiQdimsWr+jRK3eOEz4QHIHdLbOgtla4
mZqetKFHtMUN6LekW9EpN0N3ecE1AGspt6WGCUhqX1kK8/L0HKde7BI1dvCf
AQtlGH1QmPwN5x7Lt6oqz+75YY7M+3qJk6El9oXiB3RsmP4gDvayCTuZjAga
823QcIxzejS5C0f12UUvj8SM+DkGrcn4pVNDn/vpwOyNMe5WWSMsxgyzi5sI
jwcGk6Zi+Z5n/LW+9tHxrzgliDn+oqh3CgBnT/Y8tpTnDKdivZwpnLOapCrc
tRBB1s03DVyZxaTir1rG0HfLkbq/CKU7YIeHYQUKf6+lDrWj2rIs3RIoSRfD
FcF8RsvgU/XxChmVe6SHnwvwMipTi8wZJaaPvFyRSkdHLgD9L+PoxYIq5lf+
1fbDABgritZDhWFSLktmevStkvu/Cg65aSo3M+outCrAK340ZgOA8jX93bDO
++bDgHgfZCvZDMK1xsqJyrLvSOJ8+DyNEc08v9xH25GHxn3gMQu2qdqUTkeN
iDCl0jmmRi4wo/c7pRoEbIjR7X/fSbtTn34gPWLAO/ZCwrNmJRu6ZOCnaYzE
GQVa6nT7+TRTTmCISjay2FNCioHowmE+RDJpYm/ryn9zb6q9dMa/pBNF2t99
op0TtJRK/46fBqS0zNns/BmXByKSt4CJjtvtuKzcEDoQ8wGSNUrAQVJLDy+3
ITka8qtpII0plXVsQx+p4eyMqy16L6Xa84ft7ZYswHXJfLd1mVBcgph2lIoz
WU3w8uHsvmiPOiWI4UJ9x82aUnejKRHnlI6aoIvP4adtTC7txu5LXKVt3/zy
e858pmKIuhKJKTogYLVK0gtRbFuMjY8uIjzL3wl4kD70P36KlNN6jIWAaEdh
vVKoeG4QamB6Rw5274Bx3BpgPLVIh7p0F1mH0Q+7UP4gufu+S6mfkP7Zu3y1
cXIASYLJQH6q1LiQJlQ8Ir9OZBhUMUbyIJCj0wdams7+CCO9dARfIuTnvxeD
2RUI+H/wqw0NqbnukFpZH0qr0Iwfj7DrOD4y3T7xbwOvABQuGCUSrnxDaMf7
QFKgZ4cevv818WjflRglqUjFQKIrWSTitRhzwcIJ+D9+a/YffT13uUfMYlaH
/OqPTFmD4sNTWfePsGHSCqoaaCUWQl5SM7WTCd9qjfl0NpamKyDUxvjO3GNr
OV0vtIa5wfIvMhVxZjotsW1IJyXtxKkODAtL3lGo1lWBT6M7gpKSgVpiyRDQ
V+kaIp+CddiIusfw+tBggW+214tB1ir1MJrMvS1or/GptxZMQ8xMgOThTtQw
EqaoItCNWVfoizU7iYgB7RsMOGwKyaEs28XnsjJ6i7eQ+G8UxJx5oHzTuf//
NjUNgxFvjxOuV0tXOPJMloU4jMCldRrYprEExOA0vWihfKjpfndEyPXosPn9
74GR6JIuL7IhZeFGbQcQo450wuYSFWvubhQ9NWhl2JYX/loCeEJgu9zQTxoy
by92abLDsbQ8diwWxKs9Ofw4Lv2J0HuRYIpBG8vE8JN4skbrj4Q2CN701NkM
/xPhMOTqCbDiyTkF7HkYGsOS4gFeMTElV3NoDkXx1A/Ox/d7ro0L+3H39n78
a3KMnkTQXW5+kLszciaXkzOY08gHJxkBuA90BdynQZJv8F5/3yJMohMrPpgP
sqrHWe+RdYsd4XuXsOKbKUfPIzBixl5+qmvF6pE9hw8+Mx9knaFa/oxUwN0o
JYnjs9BPX/MSLPioOnGfn1dyoEc3+RKf0qxnf2PSx44Ak/zFE4ZG7BK4/hql
Hwhwmzb3KnEGngK74tl0mT3mNTDL/H4KubMaLjUi46YqiDAFC8fBBSoQxctJ
psalgxVQUzAN2TgJa4fO5jvPoTR111qS6BC5WHHwav3Vv317/b9azfCyjfpN
kSgvk6tZpVITaRJUrCQrjXoTSo2tFKAgppry35pXyvcI/ft6XmHY3q5rljQS
6sPc9kFsFgHL2DbKxdPSTn1oVEmVkfCiuuSwCUnG7MXA9vBILQYW+xsMoTts
SYRpSrx1P4W9gzJMCR0ytE1ddA7r+yZlP0LEehNDlU7phX2NIaqiPNm41J5T
jdOaoojpKe6FUpMU+Z6QkQaXtmHyOLh0EMgGcXPKmM2r0Owlq7aOoMg7E503
yeIO1KP2JGa2yj+nN29+Py9EIuL9Y9AFiMsFrW6h/1m4XjAnUSjxGK5nTimA
aMwX3KgEqTkAAQmxKdwa8YC8hZaUY7EnXJELJVUVJD3QFZzTbmLjqA0RcU6i
RwYVNuYKcKt+sNr8+EKoYz9SfgsKKzaV6Ko2o2J/v7k8mhwqf8SHwv5ChTa4
UOSY83GhvEPpDfd/mHms9n95u6joxe5VGaS8QkTVw/nRtcLquKGLw9IsyVoJ
0+ZbXvy3GEBMJu4W8l3fGIi1G/4mfmrppuAXP0rNbxwvhE0sVXjLppVu3Jw+
HOHvoelAVcLIV2BoTQCjZ98IICEHu0usesQEmH0TzeQrmCLSyRnwbyuz1+4i
VTreRsXSLKfa3ohQBmJ/DUhZN7aiU8aaqmiVMdPHs8oaKNwUm/4crB+b3+QB
nJcx7ZyrLZblEjaOhzsl/uLtLtzXOcHCj+H3HLqArAmoKMoQBo6PpjtCPiIv
w5IIu1ePBiRltbvrEqqBFTnUZj9zmpWXftLsPUGqamDTKX5rY863ATiOk9+4
0pSLCj2/k8F3XnWTzbfeqRAMnRlxIZ1lJ6xwUvisArc7rKW2XxXTcbDR6Uaf
KR/dJ1aSoz6GZjj5U/BXph7yfFgNfXvNjIuUO24Gcdq7AvwVWFrv3u4vCscL
URRYtlcXXl8O9vfwGDDX3GMmrh/gJUGwuYUJ0cr9xfq7G18evC4U4OcMm5qO
O1DjgYj7jHL+5cgDTgfwzDWEmYEIhp4IhIReTUUW8WKWlJ9sMWF45/WDoy+/
xSK+wJxj51wAsVKap7MsICyOng8Bg7Er/O4+2B1nGAxq82WfuvFiqldO1cb0
ynxx5cTCXk8WcuMVAKWZjWd5vR9NCUkrtVztlLIQd0aP/b1SCb9fO1TwqUN1
7rj/ZAcy9uliuPZCFJ7x+sL0IM2Vfti8Va8/vWA4M1xBIbl6ewrK21JwMnhn
+HyGzywE1uZ+fvlPB0j/w2u9cB3pEuNmE6TyXwvVShT9ZPZN2RLXUF2aKZsr
nQEUAXnyS9vDCf/UEvLvgI1LLu2HEIVgc4PilkkEdhcXJVZd7rKM0KgbCSfy
g/xOkkzU9l/qkRSeHDtuhPV6l+XHp8s12bfl6INSVJ+q1531cToQgP05Axe+
W4T+QGAYnZdTJY8NSUgycq5868Z01CnyjGlTUQic4F5XPszyhJYL/Mo32/ng
KaLRDZPVw917VfkeotWVZp5hwVwupg0sBEMZuPCWJvrnAsW2G7C2/lA86GH7
YuocaPdg3eFYj/ISaZfyvox2CDJ85A1+E2SmDkoEyXbo7Y1P/BDQfokxFESb
GuLq2Wm/JD9ePYEm39bbd3zkBrha87AIFN4Za8SfpFBH6fJzXZsNv+7stpKN
mvaJnF2ZzDoPY1TcrG5oQLL2ggGMf803IS7yjMMKNs11G06H1BrRR1mVII4F
bTW+iUkcExQM+O1WfSJo/Isp7bVz4JazFPerqsOXkufSr+qEs0dDBbUUdxIQ
X/r2/7GQlsY5B7SRvfVbkj/1qTqqzOSvZ59NFFbsD/RkwHnyuMzdrmBEhaUY
+lkslgIXptMrxooPnRUghkG+HbY9vYNNowopoFuuV/7ffivgrR7VkrYDyQK7
Uc6At49TL2snVAn7lxgpQXwe4RcNHpPmM1eA+Kot4ZEE4qO7fkBCcq01R7ED
bbDeRF2yoKHOKjeSsQdhtXRs615RAFeobDwruSzzcWsziTB3WRrDus/qqFKs
tp9ZXQdnMLi9FOzfNVQ8DSNjtVCl1eOrpBk+BDktS3qH9uWBlOf3EhPUbyvs
0N8BU4IlUtPVWrRuvHaPz8rwBhqFDFihTp2N/5Axr73YC5lxRQlyW9LkYDMf
AFosh+9gWYygdfQtoPaJs8FlZMmm7JhgSUyQig6SopzeeKMPPgRyiYQsRHma
u+VX64yVm6Z2GNktamxj75q12Te6Bwhf1G+fv84J9TaJe6ZGs0GLgexfz4/N
/vFjeio+J9qsgaB5F2WDuuGG5uV3q5Vz0O9Xo5C1AOrBjTJ95mdfPU2wq/Wa
9+BMOJ8TKYRO1n1L0IzOift6akxRsaSH/o8+f+xXaaQr2GpMZDHdfwDf/3B6
KDgSXstOs4Kant6OAlk8ipnGJapKu9DLZhfNEkgVeGGh/+Ywpzn8zdIknjEe
29OlkGNJ3azLazhNCvsS9z/vrQZhBniie9Sw/xmk0JLgf1Kg48kasXPhFH6T
XR22vgvgMCyMCDXVf0lUsOFoXHEEWbp/lanfusAITUwM/Ny2gF2jxTwbIkEG
9WjmmLsQLtEPK0vR/Z8YosdMbEmbpz7HS6U0z/Bv/N58qFKoVGv1aDv9MAC/
h95io1JIerT5BQETB9g4A9HMnc78IkG9AYhTul7udD+DETs7kuNFmKVCLZSR
3IkhvChfaZoW+u0HRPUWUx7klOLsy+ypHcYuGMXohATI4NIDldy62A36PGAy
PR38jaIPbwr52K5e4YYxP0KkgB9hQALiyfkBWSvXdacaa64a/agn8Q/UuS/x
w0Y4l0kbKM6ip0/R1tQpc++3fcdlsoP1WEbEV0fggIWP706Do3o17hEKkRxe
5lQfmMZDrVSIL+Cee/gN3p/efK/p0DXiCSKS0ifU3NbpGa5dDUKLEBKLiN8i
fJCoOrzmOapss9Y8Dwqp1li9Sr/4Tro3C3b+i4slWZxkO/QBqNuugq/A0MBn
LdhUro6LaDi+pG20WsgnTiYpH4qEeKB+cfituujsv9LmoT994UPeR3ol8yZf
U3TPCTdGeM7QO9riij3MbkA10+3RSB8ZTps1YXmFIX83qcG5VRy4VctRkbVB
HgjIe9e3fAOWb1wEL+AmjrHbB1U2hTo2NsmezwpxHwrXG+8I7HmaBvXY9JeZ
SvEVNQrxQgfhsZV0C53vaXd0CpXlbKXfTPxwAEXeKRX5PkkGZmgH7FVrKl9s
hm5kVdGgI5AC11AiIdhBe+SQDmhp4rnmlq7l9bmgPfJak6N0fEKLpX6sgyS8
iid5K6oVs8foe9iezo9ILvvswwYdDOP8whHyv5N+layShWWtBRlUpRXleeyB
eBLco0CR+TOHhIhhRZdv6a18G281A/o+Ia3ogwjgBZDOcKO4yrdGYCCpGoPu
YI0i2cJBug2Cd8FEXZXBMopPhdUqGU1YsRZ/SRaUKMq/Ind6WOn5NkPFB77/
HgWaT050GW5fSF6wo7FFMVRaD3IRGHhxnkxdZmXTawjKZAilEBXAQWIKOGM/
B1B7pfBYFW7jg45TY9qqBS30ATP0j9aw2lg20BcAXddt1dMTmG5pGcv4w/wy
pPqme6rhA7+HXHR2mfyzUUho2fHLYd9utTC8szAPGktgXsU5VjBNH35S/gTk
eSsW1TgpEr8wbmu+aossBxkMYwASBLGtYTLHINLhakwC333BEubGbcQG164u
oBzgZEPQTNyUTQ/f3n4ZhlUHDen4w3fr4HRcEZX671XH9kRj7h+lm4+1pIBp
1Gl+D5Z80lJOq1J95S83lwCAtGfV0Po3C+ynW5vVcbGjliNVVlvafE9MQDlk
XGgy8J1fy91d/WsLmA9amebSGU9qS7eLzmfgmlS38NkWgU9n+Dvvysiue+RU
JznzRtTvFl9NRdJ/BLWidTgS5tK4yMHaO7oyNhn6tMKfk/VnbnRHnCfL9HO0
BMrq9HMo3vxJWh3bGfxPSEYkGl+YWv8xkq9WHUthu4m8cfnNQ4fUb7Jq0QJ4
0lNSFriEa5DTcZ1axrh9QTkfPMgHRnKoiN5NoS5be70udV9Dv4gLRoAmIRH3
u0AZHegc+ap4Per3mfnFGegaZVwnp3Au/VjQrsHBWt4/j+Kgc4mwcOMHF9NI
rjSPm/fw95j7J+uHKkVTOXTCE7f6WbAAMIApLUfi2hS5wTMZsFHkrPjJq5GD
g1wbhdXDo43vQEvHPFg7+5GT7Tr1x8sKEZC61F0cwWG4L6/j8v9Rgm99SzMI
gHXD8OCj0cEelLX4pLQvNJ2Inn5qyL6Zf0WgYo8mWnSUTsz5RBHBb6c5Amah
jAmBeRmGPyiu1EONnHNpH/YK5aRm4ULh511YsL61fz3daq7liAZ7AGp72wJ1
6Rw9E8K9FeecQU0KSf2l3iT4iupepM26Vr17JiYTyPUYkicYSNsAC5IxGhid
CQF2G7GPZ4nlUJNj+LzNnF7kx+CgvzkpeDqqKzYRuuJy74inYJV8cQK3Kebh
ZYYKl2W44XZ6KY9cj/zXcw0EbICJLZnlE7ji/LcgZHiUladdZQmD/uX/0ML8
QS6Bw1A82c6h3qu1RP8rtiiNwg5jI7ijIp4n5o4AONj0lzsH6Bzl6BE908jS
fly7BxCmYNjXfF7UhxYrMdlQZY1vdmXD+5NHWWKBk/lN13OlC/g9jX6ies3i
Q/9Z/g2yCmTuVWiyYEtbvIG2QzF2ia9jfqEupQYd1yi+VUyMklo9JqRJexgi
ZTlOV+X67eFpPPE8d4JWEOdNF/eXCBoJVJuYw6JBiFQVYCRSBdrDXCWLkwVX
H8RxfHZ9ntjfsN75IcXWJ2tNbnCxsTI5ABYzqEj4QeF2eRcHqhJMOsdgND7L
QnK12YZuMnk1odhGQqGQJR+JaKzzIo4v25y5XnFYJ1s98twxmTgsYKrTVhkv
GNzcZ211H4mBd7L0llDc6cOLmCDkcus5xehmcsGLybYztsDWRTlsWmrr6Xw6
raUVAs6JSuJZr5a+OH7b4zqeSK/7L+c7MhHZ+r9wGt+2ZgBvXWS3BpODAiK+
sUaUTDC7Mz4tM17yN9vvcJS38fGlc9vzR/hjn/ubO0iSvF5NTjFca4LRFwpP
cYUkZkYPj7R+HXN4iFlOXNHV+vEId711NhXu+v8E46zcFhXp3uF23prKeDVt
sq97AqCuR5LqL74Llzx/9h1kOVYYA9HLRoQR3lgEc74lrdVtNU0Qwph1iOUa
gxAc2zkwJMkfPIvhWj6AfKMkZUAf3QRaH1K0eAyhjGWMmx3+ck+Cs3FxfWFg
TOp9vwZxvHAbSPi6ErkVGj7//uaund7gXwkfuF2eqi4TgXbJ254tq8ccHBUj
qdT5DQOpNHLOL+xM6r2C/RYPggIv/EUfLyocTyOq725Tq0i5h+BK8BfkGpC5
dJMtxvITBo+Xpno+y0WxWFZv08CWkj5+HZtVpHCHVA/20amqC6tf73szhuXi
duSN66/PC9rKqroNQwD3S79CuRK/NmgAKiD0UNLuYSjbVvVoBko22vl4fexd
g5RZin0Uodu0X/XDTPEXhbTkY4Ty3DBIHJKy79PNTm1AJhwDP7/0/DkYgDNr
4iupNfrEelWs26KJs0BbxSi/h9jX4fk7x5lT+FgSNpltkvs8hHFUiQrOD7+Q
kAwlC5CgBNM8cpyowf4jB2RoYDOzsr7YKkMvNjURyKW0I4PMhjR6YbbTo0+8
tIok7/xMhpQfaNRqNX+T19AOHVqS44qkSJbHvdolAk8T719qr9h+geWRTaHz
gd/NqGk3eHUum7avbGIh1WmulpcV5u2Pj1mGWyGzcnwTJ/bGosp/gLUQQrnO
prE17DC1Ofucg9om5fe7gP1ITCkebnoRoPmMy3CcsasXhVFOQRaZYV5rJwzI
etfIsxo5RXoLK90s2+9a+pWOFCymwEmSFlL7Kt1k7asUsyjVlPKNQN/HMY9u
CKH9RLGV0MNe3ZJdN3u0n7Ogp56P/1C9mK54a+Zo72wFA8v46NpxldFI8Riw
bsV8GMWm0Vh2DZYHPWzPxw5lxJUKAI3GXZ6KYpr/bd13gJpPIRxq35UzuMgL
gQwL1qu6sI6qaW8s1yL4gdgNJVkg5PcWomdoU1SIciXEqSEfsRHWiUXfKIV7
t3woH3N1yGB1JlUUbGokzX/h+3kolyfvBqyhRsY04AAKmRpY/fVba7IlrarH
3HSKdvsJaRq268HDhTvOgduhLXDG60vl+2EM1/JaiOGKR39aR7D8aCjEB1DT
VKLjD6aKSEOKvHbqvKyFXErVJmMUvtRqoQDlLDqAvs1Ix/v6maI40zgkc6MO
yHjZb3CXW9FYH8VD9+92QqoZ/QHhXm0ZEnuP8N7ddZFwyasW1uaUm+jLLIn5
A4wOjjEs9lTj6tBvPSaWBqhae+FdrBNj5C/0Eqb1iOev70E+VaA729uWYlkb
fxmOJJX09yYGIVSW94rlD2ryNdd9sgmJM4yAykQI/eRwk152p3ROCDZRtvWT
7lhQ4DWO5pXPs8IzKkDr6lvTownehJWfUGP1dMWXhFNucAuqBp3hX7+iAW9d
l332iiBgP5AvgIF7Dygch7Kv/CGCHvpsnKdrCiyvEl0bMTzPWnkvW15fJZmY
hGIlwQzsxI/9/rOtUpRzOTFaJ9FTRPlxQfOreHkayZSKOcALn2kEl6BUgoFQ
eDGTOh/ZUZMSf0A8NENLmgesMsqU89kb2F6Tg91dl9WYL9O5sho53B3Slgjo
DifzD6zKthGjvOOzX8wktWUBVwA/Nz6TYYeYYMDTNFAfOMVgzvvqFq/VzVoy
yMBDNMcBkafUfuGXH/OnMNYdWhNxaM141CrDkgNA0EvS3uiGW4O5xzuJgY/S
kprQ2dT2o5bBYbdYSERvMpTe41UCyaJ6Tl0BJZmN6DkN86LzHbEyPOUcOjyM
1SWs4rmW8Lz1iiH02uSJN9HES7vIZnUdg9QaIOuZ6+/pybBtz2b5bPCcmpib
q9xTBzG4paxA8UChOvVKda+4f538mGeZwr/VBAfAq3sIV5R8GsMS+rX88lBD
6qNUAdQztXPXLbuF1iU4okHJRSmCkkyupqAdzwChyjA7ujigzOoFy1s9ZiNd
5Q6eJDwkaNfudswnsITuPxmM5WKdsirosLtzuXFo2eyWCEZ+nnadIUfQwFHA
7CVidmKFBwyTbE9aXdCBgyTYiT4nDOC2es88HKILy+84mWwv6yn4DPUOr5+t
5zFaHbxrDcZzlhzJnuB2fFo0X3d2ihX7QsLRQxypvzj8bTGBRTBArSqB+qzj
X+hmm2zQY6qBW9TIpAiCnJMaOvdf/8iU0VEt1eNrFcb4gn7V3aX1for0Db9b
br0d8ycnZ592nIiFhUk/N00KemN74DYWJb/nIUA++Puu+DfLoKuNoiNL5iRI
bXX7JbHuOvd+M4Hl77BJja2h6s16u99QU7MzBwbieYpMSeUv/Go4XT2eXS+i
a8J+FymLpvOithPBseuxj5N5ViUsaI/it+2gyGy2EMWdIXMwPvDc6pg3Bunk
wT7MSskVAH1zWGVZjKyCetx0gDupTJRBd+BGmSuIeDZ76/hA8j9GHIgbSBOe
KtUwvYmmS2fE7Ku0pdoW3RJ2n2DigCfMHd+aSrO810axk6LKac1vSIgH7vo/
T1em3wn4bb8iqamu5uEha0jgEqNTXePMFMOpYHr21RIA6J/1Es+yvNT/drS/
vgB/Q7UNFOALGz3A6Z98wjzF/1EzWeUiHPWFYYtMuhSRuEl1CGNwpP01rfaz
Hodo8w/9q81JDcwVvHbHBJuPlKwdnhpTNGjjwnAc5SBFp4VTNOKwCu1vFpDl
9mofLpTFdRyJWRNpWmPSlr6X5yPqyvqnqKzPJV3qODXfOg8OzaTteP2Nhmy+
bJ622e9GoBU/Z9UkAsu7S9lfqhwvQYZmuEd2jLCgWAcYW9/MOqqrOzf8fgnj
KWgGU8v50VMTk2IHPy/ihXdGTmZdXj9ilVjgk4A9FVm4RDIcd2buVI9wa0p9
3qPVxLtiFfOIIt05MBlK80GlK/GoW/h3NIPdmvCPazT2HylfmimyoDOQjvyO
g5GstKTGoT1s0j13RH9lqwgQtCJNyGu+RuSiv+KmZJcjuOPfUZ+E8n/RzYJB
GTrT8JSsN2TGmJ1cXPISr3CZSiXRoO/llbZ8WSb3wjymPmwuL7ANVTkSzScS
5Twr1jay7gnUbqfJ58sZvxJ2wx4kifX7q/spCMQ16f2Ky02H6i0i6wtptAbq
7d+ogyeYUffuecwIOcoD0J/ehR3Xxb8nQ0kZNA79Ev30CJhaZ+AUIEWxqSap
NHwSZLUuC0pN6m/PXjkuz5AECIGSKOlSVJpPurmXv854YEgiR+rEmHz2nae2
t4pEWTRjiWCfSjnzQnFjvlqGS6W6+wtKJv/UaCYe6KMUVN3lDcgoLvkqTYFh
O5dmzuR9hMFKOZQnqwwpDVNHC3FC1070VOgs8tlb0K1LOpIaQsPnAXbi9yBY
QUKIhzytm4wSyO0f92viUnYX2qzA99EazfRb00CxUn8GugYiqfn9ulvyYJn4
5lUzNfzJYD/42NP75oxSR9FyxdYzWoGfweT0X7wRUbR3yqE2RY5+jsU4Ze10
337JuIy8ZdDKMyZaH7RAgLl2TLaLpu5Q008igCIO6dXgTRLqas8f5Hzj1jyj
HMRx/5u2scqY0wh1XYhmRHRB8U942lTDLxKD5vUqRN5XkiygM56ohLvPccVl
Z9hKgB2t6qmWCc+iKfnP52Umsp7VLDvw0ZF0z/u1avICRlKkjmdnhrbgQmGd
zmAr8uULC3oomYg383mG1ZfPi2zopm0tgZnTYg63AcLGhCdUH5znTY86MWjw
hW4TEPnu/HzwLhAI7+colMa3k6MDiVoUY8FpCTDOZPYAia0r0kjIszWS1Lvo
dvpSsV0RdZXQNkbHgtxInjZP0Es19zFTngGY970+FsaFWHk2V3YnkmLu85im
r7iCdZO/8Heu052Owy9s9gYGUxfTLVHxS8pL8z/2ecoqJ/r0aHdvw03dDSTj
8z03HMU745Zq1ysNPc3lKkRPzzhIBRd2ta/9Yyjem8phd8/I1MgAQJNIdIrJ
NREafSgCW08Z4nWjq35BcEcJlr8snSB0g/jHP4sTpa09qATbhZwuEijK1GvE
6gV0p5hpfk8WdoTaB65g8048KEsiHD2fjYk1UPV1ul+LkJENjMGYKHNaDYK7
HPSou32750opCGB8tJ/co19W1ifuFS8VyketlNyQTCE+Y1JnHb0BWi9JbF1F
p3Zy1r+Ue/Dd1WbMBDH9L0BecZcB4P4igrvXTBj5ml2+Sgk1LnNHUkz3mIPN
benvcUXj0b0BsRoPox7xzPDwUlRBRAeP/vT5oMc3gSWPP+vQKlYst7nU9CNK
3s00K7Ij2B63UKqOA6N+AdqFSz+y3jERlHEWGqoUOGFV1Ofr0eXvmUCXHAe7
803W5PJwtT9GnDyzuk9fZEyg023oBUh3m90lV/ZdvGBlaFAEYKcfKi1X1PVX
VOrA0L2UrIbcHli2NSyxKFxbqfEkHbedNmlZcMhKZ3GuRF120EmDsqn4JQcW
32cduA4RRoqBhobSPhOoRJsKXSbC0hOHXGRhePBIQfk+ZzshnEn4l8O+9uDy
G3nYnazQ5OqfrLFC2U2VzYtbc2x5zM5/GgGce2R4DcCbPINGYu9inf0lw9vp
OFcoXYKOAwidHDL3c7Yk9ws8SCD/ibP2AD/rPlK//5iXur+bbWxJCAJ6VHyQ
VkrU0rBv2ZHFC76Kt6X8C/N/qodGoywpyP31o8ScvZMO18kPYx9FcoLoZf7U
ZBXKBrGhSYW9vUPtyIH5Lgmqe8DYgl+oY5u7pY/+gc1EANVD8vipNx2frDh/
mgo/2PTYgzWFWe0NUqsDGr1qzMi+WOwkkOyK7GlgYcezncN5SQ1SdqQbqs+u
FFxreUYqXAU49UpTEKwf7oR2pex2K9VCe26HwPxmL8oMSl6p1g/Kd4/NrLfC
uh03TXqA7Ubkf+LaCiIvPNaOXqSBLUotipvtiiBp3B2NnMMiI1I6runikqff
LTAkILVztEe28dEv2ZtbTskHLxdpdkB/V3weQH6BXNKJvjtpXWCDk7P0J13T
GCqBrKtdIV7PjCYKTF5YJ+jGyMTaR3hTleaY3jC7rbMYcykipsF/Sj6KDW74
nD3Nwlvicyjxpywl6zb9v5WZbp1wRtbnf8JDzLlPxNiIRVlreZYlxzWBr8uc
Q9ucQWHghzU2pKOvX0GZswDFB+71oJfLnK2xYyETezhDRxIPNVPiSlZUM/Yn
TRrNwvYocBewHb0AXY13UdS7nntHfEShcWGi9jdoUJxxLcbD1oRQ841wTnAj
8bEGOhIqBRzCM2s5K9encFDfvnOWhc9Z7QuULeYx48hwtjMHtce8HfFXcEbe
mMhsJ4ajyRfbULeOIyFRJnrP0i03Y90TkOVp1dYq9v+lL8FaMdK9cZTESt0q
ugIHYVinljKzLnkPfM80/tat5RfF3sS056U9RvFE8CdXR0x6FgoXjyv+0wxQ
FjKj1SR5B1qfKlxdj8FTdwYlXUxsZp/0jVhZiB3T7fJqAWkjVREAPMFOcXce
w3uiDHVr2moSsq91whGG5ljYt4+8sJSF9qDBmMq317etVbm7IRiJf4JfRIGo
FpvPdn+H5tFMYgLjQM+38q/PqAP2mTn0ZDe4kcklWtKTJXl9DakNslQDBm1j
CK6BDScR8Pbuz3uXLt16UYZno/cI0gaG3ayK5EzJsTtVsykdy4lmOz5GYU6G
lynvNdoix5EYTKvYjal+bCq7BHw3gMBOduadLHOL9K3qp9WVgcE8YfZqTQwD
8wyNo8VMV1Dz1PE16qQgJ+mfSWhw/r5mm3zRqjC50L8HCsHm2VYZD/6X8t/N
yNzEFBnKbu0afFRhTTfk+0WULFqg+v17q8nIi3uJtq2eOV651PGQ/UNDIlnQ
meI3gEHIC7OhPuVrZRfGIKfFzztWsFvbWAs/YWtH3JmGAGhthJwfPAPFy1nS
bQPCt7Vhd+Y59X7l0ysXbnaN5828errketQt9HOfGsYr72tkdYQ2bLzxP7fd
eJBJjA+luF0ObVQnmIml0oI5T2YvIzw19Di3xWXwvGpmMTtCiIe1NhNemaUP
gu5/kwcXyQvBj/6xecBH5vk1CKi0Uz7fA8IZf1jJbZ0/ABxx9dspECzS3dRT
IiKjykAhv393MGG8ycp6H/ur+yGqCFj7+dtsDXfHcItahyawPl9C+5YprbjE
W8dkQPyZFP1Mt+WLJ4fk0MjXquwOE/2Obixp9TAfSw8hSKBHCeFuBfkyUcRt
arHvQwriFDYvtUih+LyMnDq6nBYXazToRzeGCUF7MXQPN0ZkC9DbTHc99M+1
x2QWSDBDy45cgnLC6UwsjFTaafvy0F2Tq1qtg1Z8Zz6xvio2JpiB4RUx5L36
qDTAVTYo+MD7I0bjYDoYZBCMTDd+H6hkbhDg++6OV1d2rGcEth04CDR5/6NR
y2tAGr/DVHFgK8xERzqj5ZCV6NbZiWxnmmxxhZCXXh+AMmCmvKlTcM4Hd6ny
N7DUqu9KxWw46j4nX/VkHDJ8qH6mvXXXDG/cN2YrQ7akQEyO8Gx4lh4ja2Sz
W5GbZCS0dKSPIKmol3xZMV/MR/Tw4cJ7nfr3eW9t1ENk9zcqp8+loJxvX5Ll
KI2ENqCEUyTkKPVM6J4jmaw2J/OJ+L/vDTcL9NJ3ZKR9k3M35PW2cSy3wTZI
9sqxkYwA+uXi9KnQQce+6n+V+CbylYHhT4SoCiCH+bAJfft4ZMQOatWEG+/9
p+RFEAVl6jHptZAlPDGk4FxbWsy31h7hP//AlOlB9oHUueX971whq5Xl1s6x
wCmcYXpMrOtLNBV0UBbE5Eb5YTaEwRZsSBR4no7q2k1rXXME2rB3mYEdqEPh
wN+dVxWnPTL9Ag707vBrqwsoO6rLt0RBv9eZ2OTjtAfEs/e+xzrt5ylKvo9f
DkZCJfXBlBp8f4gr7c5zAJq7IyudgABsbSxSFbR9Jwm7DT7CCDlXXtE2NXxh
nkUQs5yrWxkRGppmdOSZLZGpJC8ItkINwIqlx8yvnMDFjr+FA5DlXZZ6AioL
GsVrdKaaYepL8iNRxDfxNhCdboHVfzqtX0M+upCdVo3uCp3eHNHHnrizVeuz
+UgDA4ocGfWgSiXP3b1ylpJGsE6hHtbUQv3O2F5EC92ArfQTUbWgrqEWKVxe
2aR2/s/gHAAp5zIpncfJHg6SOGaDWvPnwkzQLOtdWjhvXRIgrHujtn4UVbp1
/ne+nYwqJxcgM970coAM3pjyf7j84CLRLRlvHrpEKZGKFJqjyKgO1UxJ5FLX
ojBDQPyzpr+RXKOC/3h+SWIp3fWFjX4CBjeNuiVQ6GWHNulwoNKsd+wooBSM
EXXwFjRDr12riPNJwt7+wKMcIrpRvQWNVJKj9B6hb2gIpJJ0sB8/D0QKjv9a
RqRAerZiInbWllsxM7WHZSfB4hcJMu6+3iq/pR/8MD7oA/mzWZewZxLba/gb
0zjw+p7r/+Pkp9UXZqRJOfjvC/yS5kbTdV/99aVVkWaEysYZcYGS205Viiu4
7YsaNHUFtpLBjgy1f8/VoEYPUqFn3A+Jxgv454FMFPy5AH/eM3mxrbkoSQIY
jP3NTLbx9UluYy22HW7N5hdK3p6KHnA0pCF/f6bSj/9WAF9AQk/nAzz+PfdJ
DFQ9+9QgkbnWFdfa1h+URX9tT2hXEUn5h2jdEFcqJ0/sS9dUNj7JQCUf+1UD
AhROwQezw26wBpWiVPAyG8qaYg+zFJjiMBy9En4VzBteBdU8kihX2qq2V3zq
t+ZG5e4C/265xGDfrXd55rPRXg3eCcvOLO+e0OzWBuFI4UcKjLfEeLltF8s9
xeCJIanLkvQ4/XW6s5BQEv3tukJEKdbe4DpFnZMWsqMA6Z4R5sN/LVHUXTXx
5wkBXkAti9k8SP2n9XVhBPdW+jTBnky8LYDw2qACmggNOvyOU1dth6ssrzZM
1SMZJxehJ1G3G6t/pgBu2p439wRKZrc4dL5OGtlC3fbGE4i5Kz7F+Al4pXtJ
rdP8vuBvkTekS45jbibINuSIxFElQj+LpUiLOFexNeTTJG9nWofTuCSsm+iB
7pnVsCBkYbBhgw5r5hAfDY+72a1x4xi6qLiIVgojiJ0A/NUlFb6NvnTfEQcL
x+qShd0FiwqG/it3EC9Co4FG2waKr+0ddVOZ9HY9A6SOg9/y1dx/VX5xr0HE
BXdlZBpL8mNAYNcN4bmNVWa918peHPnNZBYZUkfo/6V282t4h1psqQqKj8Fp
9E6BUcG4JfbUVsOnMoUobTI1g9qSUyABgeU/BFG6GEgvXphBxARjW9UxcqVm
b0tU43oU/anC+pJ9nhUkJIQDnV76hCpuySgYVkNbkyZqMy/zIFousZ5PkVoI
Ki9ES2kpFaGtmXOXN/tzZlvphBt+T8+19cuHhi6YXeabHkMhmXArcxLKA17O
Rvoy3KE+7S5UEt/kh24aKtXxujL31AKVCI78Kz5Vt5mkaJwq/QeYWM0OHsqL
t9oDhXxUdKud6K3++k3cYFPKESy3F2tl37ql1JX07HXv4t78/UmC8Xlm1rLP
3SaE3URWJcD9/M2ua7kYv6qBZX3hYnuX7K7dp/agSVOL9brElceMHLnr2e+S
uYPumbA6luR0mED1cVRaaZVSbDOUr4Ctv7C5Wl8dg57tXP+WRAPRY/9FYyqZ
2UsEOB3dOC7FrNtijY2WMS92Bb5XJN9j8lUi9hWETmE4acyr3MaPATEGkecg
roJo/iHJwVuOxrEJoWkREW5FaF/SJLvOdC+qT6ACCqzh8/Ft7i93Q0K3Ii0Q
/bqghtYeZC1PwZi1xW19iZQjLWwTfKsub/F+ETREqk/EGHzxF1+vCaL2lcXz
gRwco5O6zIxtNps96KDWxFhQfZEAE3sbgdkfAOjIpZBlRiZNmFt3/WPNlDi0
qaSBQzbCjHTKYSSMPi+9dJcrmcW9toT4HYC4GN5D1CPQni1daeXb0LdJklRc
Yz12TFdAJAULq4auYbcHGO/jwEdG43puC+5YvF+yyAro4ulN86SQVq5aYbxa
1JhDD26PaJRRyEbLkghUoCTV4OAC5aDwpCCrmQ1Cfs6YHga+jHEpaLDS77Dq
1UfTOYQTaHV/vLXBIXdOupUYPAzuXJh7FwHtWAJ5OT3dUrM2+zVY2ESlMFs7
ANJs9o0jJdolmsOPQpmMoM4CZ1CtidFyQBsCn2E0g3HM1MBr1dQDQrT7fU2b
CUpdvHO7lHVvispqkkMAtx5QEadzbrJmIFACzqh8w0/aH9bp/DvAC9m+5n6Z
+ZoLMuupFbAoYSpxCKNKjGO5tYshGeMNXTWAr4COzv8SgDv8B1J319p+mDDI
pXYnnRpaqlYqtZU9r/KVicEYRkRi+h+wqHbbwOJeLk+N+giGtD1/o06WkPba
7HWkcXSY2Y1et/Urqc2yAIxg77t2I1N5dxXt/5v6GtS/Qxr1RS14P85n6fl5
h8QJwb4aon6WJDn7/CVrogXhQSbaIFnQd0pLMvr28Z8mTSlXSReGeYi0e+KY
AdPn/YXRxX7hgRuOCtkvXBOiTQ/JU08lqPwenrtK6Zzw3rFiIGRt1CYPNM8G
XrF/bV76ihfZ4fUmuJS4+LGCiz3GJqPvYnR69uIYwIQejjmYGaewrHfXvYZN
NH0MFPonx4np5qGbRR0yd6+d44/ART4Eh1CY37X4MYBvyRkfxIluyv4TOPEy
+bzvLJuNbN5WxqmXxp1SV2yAakXDPDLtI05ZNDrp7hLCs1eJPqEkljKWvdlm
Lu3urf3Fpbwsyx1YrcudcXsG3L1rh38k6R7OUoRWX+sds7mSt90tASXwd4Db
FR6PNH9kAks9LdG7CJxE4xdi10EyrQaujXeVSys2bRP+oMEovmDMuGylb0tg
eu7bXkdkXslK8ZSsq5WThV/rdh3PpYgz54G0exmkqeJNkk6titDeqkGN35VA
pCcJ4Gbmn1d3zdaqpJgeQszRsJUUEGk8HALMF0EdHPfCYkX4FLXyVwWBCvJ2
xwGGxiadkBg4f8McTapcPw+fW8/KhImhpy4efAJOgIH9l0/1e+T5/Q4Pwki4
ZPLoU2D+DKpduopL5wL2i1dh1T801xzylsd6TM9kM4U29RaHZW3ogQOoVzYh
GVCisDyMBXd6pvMzW2reyEa2cq0OYm7SB/zoJGk5OajGmEtONA+24UzXMjXd
qdGASa4Gb4cnCBOAFbvd+nC12+PlsKGVGO1rSiyozSByDEPXe1VqTU5mli1l
cx32bp5frUWzfncuctcEtsjxJ+oa5bUZwTMvd1HrCQkb2+ecqK4pVLHb6Wg7
Phmy3/koG+1FB5AIZnf9tNdUsNQ7HT2YTJgdsokfuXZjc1KqiJfu5VJhoUBq
/w58rbxhObHxfbdjTt/pq0pnWPrsHlsTZCoj6TN/om9XwFU8iR1LdUJJ89WA
2SrqiQ6dGxuQU7HxMQqrNDJAKxVIQz3nwnd0lcUfGcyrVY+N6BqaOM5EAPV5
wOqvcfO/6Zv3nWwxXoc2hwXWg1PHSNWZmCS0O/ZQRuGaeFpa6sWLmgRl3/6p
rvEJReh/cPe/RQSFUzpHv3ABnZXa1PexYFC3QyoA/4PSa2orEaaEXF79xMUX
WpbLa/wLqFaYKn9v3uTie1fQm4/62L4mcMGwrrbKlc6i0KHdDRA04DZybnAa
GplK6O5qnb6CWF9XfBHvd3m3D+ASHMbGElUy4bNoHjOxIUkxcOL5n2+CMWvC
GHoygQKeDSarWpjaj5DLZCdWlImk5m72TlMEPSI5hI/jVoi1b5rjGTsVr594
+bNPTX6s9psMCmaAXkZfnK6NuunPP9OltdNAyWI8aVoxCjsLmSzSfob0p4h2
eh/lrsKnhf/uawHrbrF4aDbCrI3Ir4g0h3gXSVtAe890uYCJzpHeNbY2nkrZ
rQ5cUuk9yEkaHeLGGQCuHRkHRM1YnJBhMhtuCJPL7ZnwChbBfbgPHTTk/jSI
DaX0/588XLCkjpd6xXMj+sEXQOj41SaMBYMyH0XsX0Q0M3ifZNI3G9JkjZCq
fsQuGQbIhHmbx/x0khauyYlruoMD0TK4x81iQP30YtPCL5AZFZWqlZP8vq36
0kEwfbWf2IAodymLMWBeaAwTG4UTsX/EktlDV1/Hjqz+c4IzCFa2acIL6ccM
WKTG2qYLyBaBuq7uOx/DT/7+sEiQa2mk2w9gmN/89Y28ilYPHtjWs50Rz0vp
PU73I/E1h2UcqoArN5ZTJ7kdrWaBAAc3DKx58a9YFZ4djpeQxt1FcuCAFiCJ
giM+LZ/YG1d42LQ8qfKeK6WgkqlYm2hlKwE1vWw2W+lepKH9A7MWKZ/NHoyg
UayyVeOn/kXH7gYFpk2uKDZAyM/IwNFSkrWvRc49HozrbgtjiFF87ROEz+GU
63cbkPmBSDTW5SFULZKmNvdodOw6m+EU2Yv3MGw/30rcY6xEuDjOmZkeeZMq
YwrkI2ZLYg5lto74vFOD5Z5L0b0fbxPJb1nUZUudujz25893u/+fyjzQeeYu
Bi0k+1ShVajidd6uFXgkBH2q4IY5g7j2o6GV+Qk9uL0yjEV/qx2JNXwHjlEG
DX508FyJK8y2FF/RIB0eYARrnMGVuqWLXHzb03Qzapeo/k3UkhdIJOdjS18j
iXg+a533iWjoFQoPVQYpFqeSwbEaATmki3PKYD1Mn1BYo9wLA2O5YhhfAsom
t0RnlWmtWoBE2gF1zg7eu/uA4gRZEFzE0BFrZQLvQtPvjWqD/paGiG1HOJ93
9ZP9k3gWbdmP+T2Mv+XQvRJlfF58zDz3ayu2PDHTh6LBsj1Jwu3dSRkLbqTh
ZeekPjbOWknhemqYuBqWSwLiXLqTlcBaN5Gijw8vyoHPXUJWa5H+R50zElFg
8uZLq13SWHe6LCzds7021iIz6eFl7Z2TjkhqMwEQbHr8Fq7BlWAVUnav/+Tp
D1Wmu3HmxMehVxyUCpuug4Phm/GBLfQXiQ0mjgkRlAdhqYwAaSZfJskhuFHg
tutvU4PaHgz7MQBV4eng9zP8FddZCU5DJN2KadGjWQf5U8pOAP7c2+9lAFP0
bdR84oJCzk3jKSTC9BPZ+9qssTaPXTS8zVIMB1B93viSQFR+cMyhjUm9EAYz
d00jPAJcpB71YhGB9HLZjfvfpH7CCJJKDqcSD7lrVeERPXl8Dox20E4zHKgA
aLfpVVfSMLSO8okfUuvXtdF37zSdwZ+F2MoxZgfAr9MQDnJIW3yijmwwEQQc
NoXF7j0yDhBn7K24AqNYZwkoSeAwd9tx50eakweKUrxdZvgEc1pCh952oszf
MpQ0fx/WjQ6E2nLzLIrj8rCwgN6ZA8ya+ckUTXI2aKGn1Labrq83oh781y8T
W8hmNBVNZnBw3VNXH13yBAw1n4cM65sD+UXft+xG0L55Fnu4mLtixE8NmSah
ZnsYG8xW91fiw+QsYOBUUiHyNJiWVK/i/tYcOKa/iccZ47lwT9+Lh5YlGT84
XqcaHsleWkivDU/G8iwpJkTTqnCqKu4Yr9TCLDwCzEQEGDXHg7TFL/v0YQz8
RUoqqxIz9djsmwGzzyws0uSbpEETx8j0vfcTKFBxr0DjCshvy3ctvQI7wrqY
FBYuHKygxV8CLk6wIoLqD/kJ166VAbxOK3JgGdf7ByYtfn+/t7pjx8YkVJh6
YKL3SH3QWtSfCpeCBdg1LQgSIELtoAqkYOfZftd0qeOujhs3YYxWgOFzDoG2
EBXD/TTB8botChUUz+u2cQCdEqGHKo8tMk1Qyt/iKtJS7FWQMTKh27UUnWCa
2i+B/pTyulNy3vpPqeQm6GOZ7icoVEdAITbKFsn0kUwujvlygKY+L5TnCf0l
JCc66oQtMREJQB727P9noT/IgK0ElLHIUS3Ki+coLchnFYIbzFDoS4kqIXPx
+1Mk5X+/KlIfGheyKlSIFz8RWL1HhvALzrqqeRoDbdGanjNwsTFVaYFV3QL+
WUuXgaWZ2nBvi6Ro+Hztsk2NWxwCdayzGE2uqaeFEys4UFTxJ6QUeCnqkxFg
skDwnKK2IGccAOTHD0J9z0wi15VWdqvENGmDumxp9on0rYfLdxUlcvq7loZH
CNLoNyLZxiwlLJmB7vYR0KYUTtb3XiaAxAc6YiV3GGEtDQCrh8fsNrANBVZr
RDJsNV72/wGdKZyIk8RQg5eqkLH40lfQX5A512NM7nLfR7KGXr7pUrFhSC+D
tnNxOmF9xvyDyTBTrU/OyQSg8TXV3Rl13rhk0j75TOVjs3maPOVQZDpskwQf
LA7TQPVBgaYFiMLMKKFlxYvAeOXj855ZaQni/+ubldEq13MfE24HzKiWcSUi
e6Vo2vOVWKZZj2ZuoGKpJ4C1Kz+HtkOEVzVP8DpZbTtvk3TWGwSlWYkkzA59
rHEUcvQmzmQZUVOJtcRDx0WGS+JBDXBRpTlES/rBguEoHZpJOlEqxG2EWKjm
IJau1itmFIVkut3o9nIeqBDs37Gc0Tb+Cg/yNuEWy7kGGVVGD/lFJ6VJpYMV
O/WZXmXpoIhR/lELamT2gxlJx02nKs0dKtm7oWJp24TVr1nugYLnTUTKsTwS
qAGDxRLIkr6emd7HJUPGsHWp/ds+x3DWvJg2e5wPoL9exVg2VqZTacXrkvlZ
A3OZDwhq5SpOQwCKOrDPNnMibJFZkkAbiDjK+aON/p3V7hKLKPX/CzKNgUmy
NJdY9DqU6M1dUn8Qw2uIxgimDQd+07rnYBnbF2pKvpF5egEn5zIXpMqEbpoQ
kApYdQXkpQL52osp0WzpqgJ4L4EOX0M7zNFwtS987KENHCLgfEYNpl21qCX8
gP/gEEqNWbzMU9eg8nM48LXjOMz9I7ga+nTdfxf8eCXI3620089q/Tyb6S0f
qyfPtVKOjpMtlf2B1c0ZviWVtUqvseFKgDfhdGf6yX/o+LnPlNTc9A7jMakN
JwxEQa3m460Wy2lr5N8vIunNEd+Xrso6Dy3uu0f1FSWNxE5ezOyamIcZ+Zhg
u3LfF79Bm3ag0lDEb0pHnijEBjzYRGIgh2LVHZTl1bGV2tZhJudlnV+9meOV
8g+yYY7y9GbqF0qfExqUjEctMeWUZax+4FPcfFYw/EpkrpxZBCqZs6ZrsSOw
pPDmf/D5ZZ62zHRtDcYZsBlJ380lVvkfzCJQ5D7JLjjEk1hp6mu4789SiRJo
E9WP72hgreGQhPyaSnB8CHVGD20qwxskbtvWlJxakvCUM4VX2jKFyx8xu9WY
cC1GGCcJWJlcvrGoXFIJkA05BD5DsemAF8LnT70T2QkaJjFYdXtOsHtT3GC4
k6WEKLEb5KUDLLSAjtc04Ev7EhwlDqSUVldLxf5YLjMjRjrb2l0fXokD94G6
nZc4VGqhcw6F4eLRiQxVBd1L6+z6Q7VZ9wZnp7JKKSiIIcfWptT/8HxEU0aQ
kxLqFPQNNllnSJgRSXyUonVNVdg1q18jQYAb35D7Paz/wPc8VqK9be/dqolJ
UrBq3MiiiggUX3K2DqJpjhxszacny/aKfSCa5BrUP1/NMeXpid0UIVKBDCPp
kDKfspZ1Sw0hsHv4Mwz9I9af+eq6OXg73iZHzeI4O0R8daKXy1xZ/vfTd4x3
GxAhWsCc0oyD4G6gakN4w5xjptpWN96XofDRlM8CjiihBWT35lHiBLWoPHi3
63EWJxPiRRdSOjfCXkB6Py0s6NcJmAW2/7utBzhFbPq168oSVV9rpSteezsY
bhEay3TuMZJfKxiCRowp4c68bIN33bZXdd+dQswCg2he4pP8xp56RIBEPX6G
TkD78+Kg3uR3TaIZ9d+JYqOaq4M17xDr7mMmIJ5VYe0Vng6ijsAFJfhzHWvw
4UydTxRh4lsY79k+v2CNydrK1Be5EEtZw0cCZDv4eevzqynL1nZMqc+JEVBs
jlPKBVEnxVoPdjJT3GnSxFtCwt1hWtwlolLQHcSIpLFEbbXZ4mWswFsu/cYm
J5mLEMVAfUgvhJWTYEgw634np0eqR2tFRnXlqPgi66EFFsRbtylpDII5LuMh
OoISfWOtTf+Yse4If2mYHW+es9I608VJL8nw1XM14P+GBlPrae55JYIuvSt4
TdARnALq+XC2IrnOku+5z6Fd0c9XT0JaSr13rzAVMs9d/YEugD5Z23+Nh2qE
duL0GqkZjPhzFf4tek4AtQCpSVaAV8twlLY81JPxez0GZHZ5fIm8uw8D8F8u
8Ly62mmPA9BnMjmvRwvnBrOkd90klF0Mhje2CH8TKyBTC/ErivLOm7pZWbTe
/9y4Wey/GMGluRuR//4Eb8J2yDuKyS5Gqn7JS1aGIaKtqCLuhmE56BIWihc0
ZqgwiuRbkvAUs9YMjR8yZUwFqA62NLIntbY33X0Se5fHi0WXlhrAj0JdnLsK
0V7HIGrtSSqxSpgczl01qME/6kg2tYWQpV/3l74EdPT5xh+tooYPPk8FqWv+
vnd1arngSlnK0vAVfuu9/IFgDqeeVZ9D2rdVfJakH/MxViB2dg0+L3HydswX
u85IqyCaMq0VKBVlR2RusqXEHh+Y5LM9plFN9rK5MYJAKZSXp9QiApE82BeW
fRqYEhyN2/AdwB5tHJalOEkztsExZ/ikShXCvll6efEwQMBGoo5oodnvPhes
ExEe7o79VsJL7r+tuC0xQLhdaF8O3M5CLefqm7VJx6ieBLCzq3jPpt60eoQq
lehDoOBp32Qm2Xy4765JLEhMl5dEWOWDX3ZVudTwXr5qpkfGX9Inh5M3HzXU
3rqXgfv/Q3a4Oaaf7BHm0R3cmi/zbDJ+P3eHvboFduFC7JIPRFwy2uNJmhfy
SfM2CWw1jefzEsXEqtXIyQQZ9NOh9ZYYLdysiYRUzOpUk/zqUs3j1OjOqB3i
G5hNAcPRvENioiQPX3U1PZPBq4rJVyO5vB++IL6qPHUpYYwb5OX4u2XLW0sJ
nEoHKrBnQoAbQPC0HccmhOtVci/mclliU+5SBhgcneLd/UlPu5kKOiC9CU25
iUwiLchh2fSki7PEB/BEkA0yGq9oLNAJLrgHCW9CzKnWqzX/wWdu/mkh45JY
hY3cDvP6kFsLJoPsxXLfSEOkD/gw+8dHjP5ovBh0v9iroo0s8VPp14YIBgDS
9vtM6AL0EhbqpKl+L4zh63FO2oUpQifVbvoBjUDz26TAXkJ+15DsCWxDHo6Y
kZHYcJdNvh5P3YC0X+oI5QXjPjtHBI4KO5ERDCK3lQqxq9gJGcmwpUwZgvBj
MUnE71UHhXfDG9vsG9BAdTArjh6aObLQ0+SZQ9rjtRAWXZvxmXCIc2o0TlBd
1FR3Nv+Hd2zHDAt7TV/zgI+GzTsqZRG5svO0NSedX9J7IFS7daptYHhh0Rjh
DKPp8Zp08krQW+bpJM+FWV1Y+era2EnG1aG3Zj9uHQw6NEUVvQcfTip310RB
om3e6537PtwO/j2YEM3b4NnDIrvbn8b9IXoZZD34YeH6dklVfqBNyWME3yVe
S6r3yUrja6kVCSsyrW/X+Mqkbn4taa22wdkHCtWcjM3T40G8EZMhjpp3pKRW
qCgPZGqOtQGD97Zni6fy+R5H+lTQNXk2/NIjO6Hm/5JiQxgg+8NmtrtmZsDR
Lm0zXOgcVH4sAQAjRw4OwCR049FNZzjGfUTrBLlo8UiH+RpSjBwvYZ3T0h8K
+kkFIvSrppfkbjlt/MgOuDYDKQNF7o/wfb6cAWVyIDXJUtMHGYAoC5zm/FNI
4UgU+ZKPmzTRpi3trEupYQZLWhU6ENb2SSoB4441CoPWhJzAJ4f6NcoJ2WN0
f4hiVQqVsan2pv8IpWjKW3Ws5Wqg2KKSetl1k7FZg9onmvjGX1fBVuxeyHOM
GLrl3Lvmj6V2NapHuAFXcIMD1gqs9K5yGA//ubttLLX8lwtyfnmZGHARrFOp
Z8hDesf7EALe7uxX43g2Y2Y0rOHWbTyXHpKHOwBOuPPLuyg7mH5yOLe09ohm
zscgbexEmxf6Mylv1SY0YeYW7abzsSRFy6Vc8t/T9f/KFmecio4f9tXjhQu9
PFw66LKkSe/oZMSE1YJAua/laA+r4rkkwG63uxeP48lL8wP7TAXhNN+HotAH
IhpZBYM9I9WzoHrFbVnOughZWtGVKnJ2TboqvVWP2UuUggu+0t21trYPHpCv
bbMkm0q/b8vaWWgkX+foa+cjm1RaRe8NY3T2aphbb1Np8ahf1ENrujHAObGh
hzG9JgFJ0rc/XokkRBHw5OoXDVTbox4xqlpS8sck2oT5q818Sh8yUECScgFa
UMAu1Cnefo9EudBKUqDjujkgTKexwonqb8/sX5l75UaRYfUT2bW/qfVxoryg
FlCrLV50vadXSScBhcCeIr/tApeth623T66C4bkf/HFtt0D3ifl/VcO59v0h
dkzrHkkLXo7/gV+DTlz0OqM4ADtWvyAFrbY+OulfO24T+lfoyAh167E6y6RF
89BSedfjDN0WwDI5yBs526ABrR13lRhb4T/rn3bV8NDfwenRW+DAx8ZwFq+r
MhcQV86Tjr+yzGrUbaIIn4zZXBaG22Ju/5Y5Vg8JvcfzfBDHIW1k8HFzAAFn
JvtozDzqo4gvRMzAVaHIuJaU/SdSt5QHwNh8FuBn/z8G4neuYbl8tPzKCBlc
VXxic+/F7mnYrH10kghdTRgZBu/qpjD7oPsExtKed+Vj0TImqBlWcgm7EJQN
33HojgxDuO3OTfuQ9PMwd47N9SaMQFosgva9tSDb4Fr6isni+r4r9HFGUwO8
4FOiR3T+MZASuLuG4F30ghFmSJksKve4kQQhyRi52J+LxngKyzYw0TQ7+pAw
Ydk8mXIq0ASI2jrt+9CblUYRN8R/eYhsBNoPDNX4e3Pc/NMqiZaHvEe2Y3H2
zm69laXFFF54vl5RXIfyEIINqEo8Xr60noh/sSyOwYnAzS4ysqKBVx0/uagg
mw/Y/P619Hwf8aUl4d4Njiw/ELW4NBPjoSJPMfrh7lDY+dI9ADNA3EyIvNjN
bx2XM5HwTW8kkTjvmRJ3+hxyjBmAlenSsCB6mdEBWHQ6rD8UVNFyPmJf4+ti
1+599uRv3QiIs+lKAd9GFsA81Z3+gr1EpzQ2GzW+4vY9XmWxIbZkgNcCZRXr
8xWh+2C+3tMRDhG88SlCAOjTgMuntqkn9oTnMstpxA8d7jp6s8XvAlfzxetU
ZxYWlVyLCQ48dSIggz30wyu3oRMIRpcW7/o/xrxeHQWljB8bKNo2UgeO/pVv
1ka8gTIjn1CdQSJ7Ip2Hq++vzBNiVsPH860HxwbeQtGo+RTnt7i/62mYZna7
D5LU67My3KxApFt+ZYeKUSrpls3Kzi79+QFSztVIDFdgm77nEAZTzn4FE2p5
K0TA/L9L3qVQIhxJbE2hEbc39nvaMWQDlLE98CzQRGt6mFADLnwxIsicbXF5
DbaPLxqiIF2E32MA6xbBpsAN3AkoB8vxUU98H1786WdfOOFiVcypVqeMT+QR
L049SiAIYVFuW3GoKqp+Y8H79FeWe3sHeksxjY8GAJL7HwlhQEBpnoCF5YaE
6R3owx8XS97PxNEngGHdSf1D2z0xex98GBYgnvljfCvYnqSyEApt2rB6ggyy
6UqOfrqPqFFyXFb+ayYAM/nT50YWpQDKoLxPZ4F6+499AlVggGZdEr2v0GYi
hYHqo+Px3OqepFs+tcpendyRn70HLrMotoLKWj/u2AIR4NTxTVu/CgVJ3mL9
nsCBuMjJqqe/fBQNAD+Pj1HQ+jC3SR/pXIGMvCF2Dv4tJfQbZZtUMxhM5F4z
PUHfsYx1NJHSgHlShBzzT0C1keOLQRDiR2LW5h56Pl1xwpun0tc+bRfpXuof
jmzozaRjS9vjEWrhOS4wigkYOM9KalMxc0ehmIGzx+YoJuIqsknYW4G3Huch
OuNYF/NHfaeQyAJvg8S/UxeQBcXAiXgjWdgbwB6AABP6FKw2Br2pOp7oGTw+
ukTXsX9ITEPeSU+ZX8J3t0mHXRbH+Mcr0yVNH5X1paiwAB/3P2wLi40MGxBG
y48WummNja7lBHGcaRhCILKifTvhoYgAdO2Ee4u4dQweNyWOYhv7t69fhQfD
us/oCMRfFaOrupyOBjuUm0Rjp/Mdg8g2VM0wkWZfXfkR+BDfn8cBktZ+jfly
0Hf9B6yEGCiSbwwvy3gWcAWlNc1ClEqwuExuTrEICvoRIC44IEqvYXY9+PF2
T5lHqu/rRJ6C68u8ab679W1qeQKIyU4A2RbR1zzx5numAIm/GfDqPiubu7hw
nDoErzb3dx5/h42aExmsZWDHymjFdBjOZBkQnuJ7Sd6aitW4hcJWO73imEA8
Zvsc0suGAg7AdYE9U0L5ZsvD/JAukeqTLLeH7rDG1OexUVJjE+Z0UGdZ7JyI
HYr5bsl0QKZiUFQFnjemKGYNX6nH3IM66lWztTmWA6lYgsmp7js753RzV/QJ
4wC8qu1w/cc5gxGjJhcvaaAw3MH0GL5Uvl4GmGyzSmBHV1AbyVE/iH8wwmzy
Tl1hJohtl+6TsUgf99BMFoXcfnxjFP9KX75sMZyNiYVQC3z1chA+XIC9x4HY
1eqIK3l5dYltkIK49uXP5UCdRYMFFfQWTkMUC5qXDs9y863mHzhfOnwbXz+D
6bSxVn1GeJ1Lsf5xnH98KMvYekYG59FNBp6LTKZmybjibswEvMkppjL9q5Dc
SGcjfS2lFxIEljjc/EEDVr9qIcAF702ZLiAHtmcT1o2Agc/258pNY2sFW1Z5
A7ME+oZrhGv1t+a75Y2+mn5PwlzP+rkUy4hjj8mm7TGr3jw7Q3kF9EGb1TKT
5MJrQ7BljYoG4z5v8/QLomfw1Nkb3IF068UiBTZFAHwSxqhdVbkjv+urfi7V
x2bEsFXYNF7EelAF3hMMvPrCTpDy5rpBvtJKO+3j6UgGoriKGhglSs55M//B
bbjIRQ4ffHWs8DXkmrKeLs89jt2mZ57zYvyZIdu/++7OsfzBDvGODueUm1/C
TZ5cnAOnawehq0xHpPOl7SNY5BGLOLl+ZGvrinJC+Kbvs88mFUGm050iFLcm
axHsG4g1yHH8Xpe5I/9tmqACkXYV0NkKpOryiFQtDvpX8nc6LeR/HcKE1W92
TMDj0FgaoopnzaP6WKqqOu0Iy2txSPfJULBjlzxX9p0B0EQTmdG7ozEuMhP0
Mc2c7VGBt2liNZ9CdZcdG3KCgdx0ySwcKP3K7e9Xugl3p4geKLJYHLrDyaAl
skE9mmxh/Jq2h+Sq4aKTOLlYIDyA8MPUdxxx8TrFws7ba2Viq03M8xyYXfaw
Rw4y86wJx1R3ww2bnK7uxx5xlAeYREIz/mN7iycwynJ9vD1CCgG6+9W6l/WE
ljtfupCmbzO751CnjloVzZ78NpKSI3fF7cMIx9C1xxg0zxTryt4e5UtVV/1G
kqyZJgYYGqQKg4uNPIo0UM8ShhkR7G0XGSkx8TMXWdvhlvciFpD5mcTDtLaH
h2UVeOeRUgAzbCkp49KQTkf2mLkCpWo1Rt90wrjDbtBlyZYtppp/LqEKBtGE
+2XEtfTyaJ/qxAu9Efl0q7daJ47ltMyyUSg+tALUsJXgWOQ8+rx55af3sEMy
4oOw/c37XX06B3ogwVQMCwdje1DLTlQ1IVAz24Nv+a7HskOHADHY7S2d2QZe
Pzj0MqCbe/gM7Ca0fNaHNchZdTuLokXLSwiucjB1zUJFxB28sGBj1dXB/c+a
N+M/Al9CeDA8Xjhd/W1W6ju1MSixP3KBYnP9jiOUGLKFfGvcFoNfeBQZB26s
NDb63lZVW4M9DeEisqqI8FkZ6t0eODTzQ7dvISz+tPux2ZunvDRjk/Cu9FQs
ucVhuWCBLHLOoqzfQ+QnWqcyLRFh/DpJEyCTKx6uStZvLG8N30ykP4ZIAscn
X2GDxsXLWghtMQwm+99SPZGG5IRYtfab+0l6dLpuSOSiUbs9RvPHjnN97mBZ
591rGtPQhXz1Mlkl9QLTHb2ZS+yqq50c3M97JZD7rv4iDBq7giGjXbRoM4J0
ZkKaPqwmB9Nl8aL3bljGeIkoPzoXZLS4HhF8SwLwfu60UW3Hpw8Q+ib4Z8Qt
dqWo+zK7Unjs/KaHhP5yz1ftaL523qwzG14nYAfqco0eOjqme1ZLukyp3b6m
sBwz1xxuQvF9Dg2eZVfc3yvZnE0eBazxaGIh+bvULxJGgqCvL1bIHrgNw/8E
I0Q8oevl6TLIMYyWDnxNRtftnlhK8iPLkKDi/NxL87bXpdMsXXeksA/BEye2
gA5xH18P4n2cEaJk7qP+Y9rB93xvMxtgLbGLl+hImBJh6y8PlV4f42o0q+xB
T6zhVUfgVXWbQv2ZGq8/WrPIdgS+rQSweohIHN1ncQMIxopjUU6smiviGLqW
TFiMiwg7otJwVmA7D+G+vJ7u+w5sbCp4cGZNWxS1vIgKMEfxb50INfjRz3GX
B/TB9owN0k5yY2MRTCV4E4exHYLBrXYV66OkREqzviW86d0B/soroUigQUCy
zAQwA4e722o9gKZspcLpHL4Fg3ugXpEwz574obCYUno1tdWkAPw4oa+AErBk
0hu91nvYDIFElaAagQdc3hqFiyjv30OPy3yinrudI2HWawm24Y2kabUmfGo4
MIM7eecv+OHK9uJMRNKoegp1yKDDR4xYOWg4ynJSpzQ123F5OhcBSgiaVeQw
b365fi7WD/d5JfZSQ4AgEYBooBiooZVPCZ8JDbIjaNkgvolZXJeMuQ9RgeAX
n70jfckiNqQG9qxJ2WTO67FcWliZLDn9I1xbP7APni3DQ6/CdfohFzabQtJ0
v3GYFiHsw5X/8EzHnjlqIGclCGJ8IZhSj2cHljhWefmdjsZNwxbpQRentERR
V1Dbs9/9O24Sjlri502ptMrOzheh8PwnuFQoXiQVxQze1GplJzcnzkvAolmH
16ocXn80s8kbtrc5cPnTxig70PQutrE8RR5LD8x4/TTahS27FYOFe/Ze1jty
A8su2h/YoAAY5OfkgAJwF5gMQ/AxW6G5YbQS5US1a3oC0mbm2764jkb2kiC/
dFf78rB5lLFVcfEJCnYg3x2DELzXQlYp3BTeGtjVVyBJ7ExmD03q2ngzoRLD
gK6JjJ0zfO0m1zO78fQsbNGjRSIPqwE/LYRisc20nvhpd1xJSLoZQpo+viYv
n9CXVusaTpiQgHRXbFbCHs+C4qaxMDHt03E5nVYmz7LG4KlCss8Lp9tMnGhq
oc/MlZggnM2NsIQm+OVSjeOFEasN0nXfEnRc5R6MlbBBk3VtW9sdFH1I3pKs
ha3dOpezsXQ1cKXs7bYpDYhx1JBJSpmnipPc5U/US0iLfFdf129zrgyJzKbM
0P4xpS+dV9WbfMEnJsLmfgZb/9SSeXweHeJ2AJBizHg6JuVt4NTOUaqdu+oh
MV42W1H08Bs/AP8Himu735EUTKD4idnSrM9d8vMCqaDndVUvwe3kGI3phIw1
AezAQhMC797rY50sHrUrNo7e1Xl296Q9IGhvJKUA4JzjHiOGqOy8QL8amjrC
bohsh8kyaHBSs8ulrgkLo4chX5dGKmSLxag6gLm+4eVDBYPyli7o4ojUEYQQ
AlW+NpINWvXTBCwlR/HfdIKPLAGQU8Vt6MK99Y5UETh5O0/5B+Eypna+e8ZP
eh6Mhfjxjigi7MdFZ3URpJUKKJ68GegrVgIno6wff96h6bbJ+WA3bO0LoIfs
17EhUAojqZn10O/XNWmptrngELov264v4zow4kKl9bWRrtCLz0SERoVkh3bO
K8HvNa8XJps640VUgCWKlWX68wcrPb4d2QPJRO8iX5NJXQ8AyYv0cUVW+Uv1
HobLYEda24sp1fVVaLPNs3Z2kLlkBNW9XBLVRuKtt4mUQtNH9A4J0JyO86+x
pLFenRx9//H2qp0uqLKWnEZtO0FMGhJXXEcVSViU/zamDWn4/zgF5tVHkd7v
RuEzuFl0+fDlbWwcU5QMkBNrBgdRuxBlpDaaOV+rsqg43ZTnNg+bfjl9q+7o
QfbWxOKqsu1hLRDRZ8smuwQcmo7yDctdBe+mcUWBBBZyZKOTqwyOXHpBmtZB
1P/eZkul7v6muGTP9WFifa3KPCoXlN9TmSQRvmQoOSLru6nan1LQCjkHbUj4
ESglhfyVFwsQNquGfgxJ+JCEGEvqV7j32vx5s78plzmPjIfrLdAZkUpxVQqA
EnuMlzsP9Eb5aSLg4oZyyOMbBRT63loHI2Vh+FPr+7PBTsNuhqKpkbIzwbC5
eEjQ6JgbjIm1d3ZOi013bzXI/1S4jtVf0eUoT/fOdrb10Y+NT1CcO7HirK8b
BlpyGqR/FM/1w4abSdK3caRuAKSuDDK6xABcqoVbf6wmHJrEp/Awk2dR1D1f
aAlxx15xJfiHrmyeLaDnC3O1ynwwIWAat880NmPDSF6R0QYSbqhR5h8/K1uK
ygaz6tPIQDWL/lg/0st1E1rGz4v4ANWGHdnODKryM25eaV0oiTrWQhgpPvN3
wDtBmKkarai4dhcG8L2/5qMfbRgAXWwyyP8cmWVsc05BAYJ+J5d1hrmcMDVS
i8JEtkqh39Pukv6uyUBRNeZxki0mLDNUK6o+aEgJKMIb16vQlNQUiQw8qQmZ
46NFFQE4v7pmRridilUe3v3GoXV6oTELhyMOlndGIM5Q3xxuXauPJTukLz+H
8OzyExcUDrzXl3hxAidn+gJpNcfblTvo2xrio2xRl0lD7yVMoLltqWgZdEJo
iFjux6aRkDO3Wf5m8OloxS4NwgwcrO9lJk4GcRF0DVONlQ9tAKHOnNZPKNf9
akuX1j5H7J/IHQLHSSLm0tsvLAkVUTwIIkNWcUpqfITZrBVvkZanSD+Bv2ak
HFg7o4tn9UUp0fia27QkCFWelymRBeRDYvEqkHYLAfSV/KQjtj2CMjBuHwlJ
T1uOZp8ERLVwdCFR4dqathUgMtvAqruQXasVAs8ipFo7fIDknKzx0eIOTNjA
5YBIBHXJMhRkRwz+rk2oYzsytD0piIrSf5veTZ7sMjwXECnDO6eF9F5nSYH8
XUCc1E8nt838UPDYtNA+LNWlk/g3AWTgBCzAQP2HqLprovkbuQJA6/WWBq8l
efIR8BhTE2ACcqO078maOJsf5x0gdVgz+EDe7CHCNp0OdjHv8Tq2KTvzmrHH
RB4DNDi3PHfkZXVnBN9uDkoIU7qB1rP6bNY5CJ/jI2BI0/WIQo2abAOfKvkd
JnWRBqQY0ZbjyMlq4VpXvDEFR9dTjcsXGC544Wzd67WfYwxgy8tPs950Slu3
mVES0exyo2UAS/hMThxkn8GwwHlVvmIm6JslPgERHk8ZMLZC2gC18NUaYGOy
r/ydHVyGx+abgpHx/7vEv5bBfMfHYJ7sIeop1aanEJffT6mcr18kmLf61apj
gYb91fnnNPhT7IGquh/mvK+fXfnkYP0YYYR1p5mzCIoLYngXoDpATf4j7sO+
zdPImBWuzi0SKwlq04WjNmEssCybOkJVboJsRzFYERNzh+qCOm4AMD4nhTa5
Lh9aonQ7swOS/kuEw3vZkJa+Ee1M/joEw1YB8lwXGq7iilA5c0KxWqOrxMEe
oI9haIuSraGEkrDoxOrUWNP5yAMWjZuntOQXIDEC6pfL+BrOWq+FKGqwkMlh
/cKC1OVFsIDVc/C6hL5UzhPhDVVVMsWE/HuJM37xyMtllCvan55W9hn43gvE
ZvVAGDJAG6H93wSnMHGyrDXsQLp3zXORNgQq1RmFekoSjhrz93U7/RAM+PCN
PVeeRq8u302uG5H9Pqfw9ryTNZnopZFky8p6AdDBmZ2O1Gz6KcyDxojOAvUE
xpxey+YWPLu4neCdgzd0E4P/ha9cgFGorXD6oDUKdgDfQDKG5TNQUndI9Gpy
DYzyS2kp8vfRKFromEI0QPEcdJWSI8KD64mop/5KxjjIOwUIRmdwpzWdGGyp
SfzY4L2b8SEHyyJ5/EqeXg71XepgBR2RRaevv8HkQs9XHkV7v2DXZSogXIVO
rP4o7SuyIdYxxHspeeraoJTL6dbmQNobnDWLU8imj6iPrNl3OEtPIeVpiMh8
CRVR/n4Nsmcqhy2BYAn7yhiLcNaNsaGX1+MAvnphwAteWf8s+fMu0/ZWiRYJ
06c9FgOci7ffpI0SdhIXVGPtsRalUVcXYJLHo/0ODU1QngflyJeDP8IHlCrP
BgS0AtsXPobecom0gQSJf4mFDbucEd6s/hC75+PSHKFH+VZ5wWICKj9DEK38
jgyUIaBYYgOw/i8kvYB8+9isal8Q425crMAL+Y74Xm0dDagVk3kHVBDz9zCM
8HpYqdLAtH25wscEEibhRX6+jWCPWItGJewk8HsF8qxATdAwTn021B0lPI3o
/vSw8/C3F8ac4R/Qhsots4Zte9dT9UJH4ejrFv5YFogtF+I9CzEObSrAMaPL
fMS0A9AHaeE6BIkQIzQZK99J6Lue1BQD2LgeHn4Xj1VPJJGuCLT6i3MOO6BB
p9oQGObal+fkrRPhuvyhpjXtqDsqUPSYxAlwUT2xlJVZBGhIoLiMU9DbJlO0
i2eDzC+laaLGWlAAyVKbHnoSkCBrluux0OXWsRxSJkW1A6/JuDV4CvoIylql
3oxvBZhFwj5lz/0r56RotZfwSFs9ojYZhEX3V0RuH7FVTDBszOCJBlZ0qvDB
KvMX5sHHYgwzFh31nY6jjMiIhlbEDC5C+e5J/s4BGNN4Y73vAzQyigWqiMPs
qLWyoEomQs+bVZfFkrSm9AQBkgCDy2W4WK7AXPbgFrjOT7Jgb5Q1b24ZgNch
8ENX5zLz6EzuarrAoaAa4rhlfn8DzqnxP5rUPdHvxyRcWRNOQOrROElRyRVD
9xNx8IC5jHKDZKTT2Fw/cpiL1AkoszTWuGPx2yptULJMsGc2C2fXQPUnAOZf
5w44FvkqZJF4hR1RZtndcPLwotPfrjQXghes67Jx0/GfZUcnYinYz0taPv4P
gvwO1DkxoAL2XvPbo7zBOO5lg3T7Ml2SCMdlvSyycYOfdPMjdBscyT+oLl3t
1k3ub0jmkJjdRJrUPP27Ue5lH0lr2DSRhHDg6vRwHq/I7tlfzA2n8Q3ggFbq
AEr6qe/oyVOKtyVKFjOgDBsdGC05rQP7eEfanVJ1fAXspJ0RQWjZr4z7caK2
fjnU+L2FmHJtjj7ME/lv7WqFHec3ytLSgR93KdzI+mlj0DxtU5ZcTslWYClX
c9WbNEiq610V9dMHIxx+6yu6qiiaeJv0xySCb91Nt304dX89iv/mE4OsVgZs
Vq8+s3zr61wZjW92sLsv94OAs3GSDC0cXihZopK9lMvhxRL29ysIPcKVSfPB
lrpGZO8BLzz/YuJAn37lNvyWD8Vg86FTgxFIehdDrE3M7SOj04rnWX4D8CC9
VMKT1hYg9lVBIGj7cYbFO+LeYCsmsFBQAB8WpHSpcrJZd1qzWgNFqp5gMlOT
xKZUYImDWSnaxPjqxbOaUztJq8HvEeHPTQrdWS33yWcxkpIfKZ4yI4pTuFUU
4JWDpz9yyQYtxNQao8syUw1LhFfHROlVm41amwCISYyeV7EOB3VJMqNUp7Jj
wOTUTCvKxROvEYjcR4g7lhyUkWV1KPwkgveyrqDyeyXGaSjniJdZNTB5QT//
LuirLk3htdA35R3ZOraTE5h+lBNDyH5mOVYJF8R9KWRvZfmOqQTdZHEQ06IX
ytJ/B4PeDYuITdIRyOpd3q1Va9GcEo7OxTqH2fOIeDSNT8zaf+3h0+mfSBdn
+Uc6kFU4/iZDJSufwxAlYRRChg/0aXrPhObQUACDA0MzDL0XK/vswCApV9+U
tsj9PXzvoJA8qV9DtR0INlHtbZwOZGGJv7sF/axW3P5sBIlaKEBwrgxKCle8
TK9gD4H3EkCA4SztDBJZL0HPc4WGFOiivMu1B+sUmkjle4KzhDMPhhzuWBXL
MGQaIEbK9fdfGxVUOr0cLeKsPFD/eIj0tsP+aENGZ28KBXbrW5rLBsVRnPqN
qpP/Jj/5p/MLkHBbGTDlGl0uMS/PIhf5VYnigLNbisBRHgFT51r1yXquR2/Y
6PLBseQ9j2mKzLoGtIauh9ED8P0700SG0bxKwNzT0cvaGE4O+b1s1uAIBSR1
/Ec9izIICOy7wgNSqmzj1Xm5GKzt2T1SjeRYiVyy1/TqAEtE5/jMOPPQ09f1
yGyqfAbWVEVWHUKvfeL/sRXUnProo+JeNyXjqR6QISEfEUdb1FKiBE37Kk6n
K3n3GdqPEXlcTfIr0EW6cp+CvA+pWodr/1toMWu4Vk41qtlWR6Y6sjMYub20
SSaG3Zi141y8pRag2b4LV18O3XOPkIXF8ETcDUWTr+MnUYK9vSRjs86xKv/F
T0NyHGJPsDLnBFgENvsUq/Mxv6CCLqo4gGWLUrNjyjvboDwNWs+uQpf7g7C0
kCNP3z07hqwLEOguY10K9CBnj/kxZZqKau+FY8h0SwZCWsGf209UYtGg0YcJ
oM7slhndVcFIefvh+9e5b7kBlO14a1mmCbHjUIupyGZZMwzILwa4Mv1bWWxp
K5uUwQQFO1CSv/gSHKMNK4sm3old0n5j/ZikiiM53AdZGNM1SgyXHoqVUi+C
2Kj5ZDtMTbqOhMm+lU+P1JGOBZeVvsono1zDgoI+HTC0bNV4w8Si5depFen3
850eLyORP3J3R31ZzJQ7nVBZ5eMHeDuEli1FxgF82bJHGjW/43kRcer+JhPK
S1mxRM61l8St6rQvOJxOvb3GYQ5lJkojE3CaCsL0GhSmQkIcsDamTzjRPP6j
tgEiaA2gOzM9BUwBTu6l5wtgNssg5UMxy/xMVFnxDe5CRoyVNLGd/MeXwHWO
2fnM04vSfobStHcucdlE+m79PTjqWz3KCGboUuDmrolKBIWxilNZlEtXtqkz
5F2/iMSALvtuGgebWLh0/pQijfmDjUTcLbwrPmeDUljI8KH/ejGAFRAm6sge
KE+ja+BjDL62M83/EFAav+crz/j/A7wrD2RLZU/xS2Y3Aw2McumcuWsCbYIj
ueGLXXKgzqHUO2iKmJnjCaPz1FRnSUEEMyL3jFBJsND+M3e1x5wmdTpt4LAW
WKPEfGytS/1gCNXsXSopillfUyvkGH15jugl80NmtQ0wxIh/KnCXdCsg0FIN
Ngwga7JCNcO3R522JoVnKSNiEsjfRgJnREH3eyJMkDQDh70HeOZMxDiGMqwU
EgHrOB3wj5UCdpl1HtwwZ8308aJngxcqqQFbgJ+WMvj3tdpHSqHv1G9RqmIQ
wSRdb4GZsGphAwl0E+cLiVI3jqcZ1G4hvnahKpFHR6G3Fy6BJZW+qg2ReFyO
75/CXzzQ6IN3cQyGBQA+ZWAV2mG8iPssQyRAjQIvEn6UyWQ+nVqyJAAGtKlO
mTqBozg9oWxOIrqUCfrQiaodVWUKeETPeYWiT5wdIKtx3JEjkemjH33tDsbh
d6EMI/eXiRuzR4qm7vaeqHJbcPFqHtwyfVB7CjV9cBlkD3PCStZRSgXpGk4w
KfPEhAiGrm+yL+GrylnqBylDwIO0lJ3IqDbvCD9nRiCUNRpMURjiw9crQjzk
Y2vqW4P6+/i1TbktALSgmUw5/Ncov0TAsnV8DqAMoX6hb7tDvdebOA0s1zCy
XyHnyM6aFw7neipeof5/NS6kEQzJugeoyjb+AsDb4BO50si8l8Ij1KAiQdnk
cYl/IZpZlo4r+jStX7OH5ZvvDVg0tlOOIil23oAorMh6jcTAC+6SWX+FuIP3
aoObKpwf7KzumWDssR6QAdTPQzCc4q3n8QuAv3RXHcHwXsc1W2RN+vc65CS5
l8E/qtg4m5fqDuVsJOE+syOEPuLfFBOE2UpyN84lRRY6r3og+rYFOwzsPzi6
szdQDXjivRDyt5+oXmQjISclTzJqJlp3JCLUpECmc1tT68RviAex4GpEHZBe
MSiJB4CyQvp7w6gkv2vi6lbILX7ElJnmrJHQee5drsNC+i+7tPRTkHvWVOxr
6SneaPb7XyUn2zZqv7dY57r2Ww5B5fi4NkcusgkDO06Ba85n2lQF0KvM4bpV
ySPud/oha0pglibnQdcv3OQ5e11LOKVogSHFcaRawBXzlie+TUsJ5FcoTFMR
DyGtqRtJmYvtLj2ZWYt9bo8rMOCaQV7Z5gitEobQ+gPjBaSk/u1oMgdQ9N52
r3+m6jgJKVKZ/8ErF/UGN5EiHs78dCQym23EmxU4SMJk9awIYzIBFkKohexC
twUonzRhj1S04r+SSIC0q8/P5kPcSSMvGrcd3Bt7gkbSLRu/Ku/es47GzkLR
Dh+rWzD9euXmTFT942IgTcI1KyymLtDMRLHQxJiMnCt3U7etnK1AJCbuTpBG
IVMYyWQY8vTVnugPWP6qYQQfCG78oZrki8Tk+KUCy+Q00ztSVnLjjxvEHAC8
aBAw5mJrTiJ/5djWrfMd76iKDUBDTkDiWfnYot6TMVlyazl6y/ZVwDSqx57C
Gvme0CSZTNSBSPivaTbeKJc1O4U3NPQBkfwyha/Vjp8Vrd+9DkYUMslQvC3p
9l4d0xRMqMz0XTKkEKgp8in+aiKsd9QTFHIjfU9BRydcTWhAeMU3gh6OMUEy
lYZjwaRgBa2Ct6E34AyJNk/lx7qk3YvnNovRznT3Jw4VOryBp9+zv4TD/+9G
D5t4kRts85rQ6ILfvdRLC/Nn3+HAs8D0I8UmzdxNk/N5E74MN8X+uY5Ykx1U
5f4qMb6w0G2mKeFHpQ89yYAl6qelUb3Ydr4HMq6UsgSLYPL1O5RCK0ox4d3V
oJyOzgC41qyKIcO8YkGYHITrcy46mLmGsUSm4Upm0oN3WcSpGT6BxMgfrpJw
6PPCbikD9OfaA8bQre3zHti1GbOJ1dXDSbSmRoyb0STMtCGHIhRjK/+LsNm7
I/ktVJlL/2KFx4PpieOoM4ubnBJipQ32NOxR/pmJaJnHR1SKbt5IMU5RfWRl
RjA+nTPjqf/MXBvv+RHeftnfjTtXLssUQUpDxuSPrDKpHC1fOlr00yA5t2Vc
svPiDW+Qlazx/ztGJH807QuzSypWNM58MMiNsU+Q+i1CZaIc0SL8RJu4rsqi
YqrrXyVa14jfJaKzeOXCA2JgTT8HYs6QABunmQdclcAheIIunEoam4F2h2LL
jG+GqIdG171K2QP30Yvvj/i1oKImeg3WL72nDCyOODzPgqB55Zf6PG/c9R2e
FsjboppqOQgt6aoQumUn4ul+HBLg8ZkmH1pWIYuPM96qOwyo0SLerFbcpULD
OuEfyWgJrkVGButfaspilXyWj3BczgST8PJOiB3xmvzVarJMlMbI1q8tGcwk
VmCtAJqBcmdpU7btBwIsDEhQy10rD+XMlcV6NuisDnkhm/bFJOcx4dLzALQv
rid8UVrPczSK3SVV506+X6cwFlvvvpMviIjWncWeYL9hqs8Q1jrLPRU7tv2X
sKCdKWdxIkF7LmjYIF/K5n2VrsnQ2VKvOxJY3HvmpWIT+dDZDAGJDNdg5Bs0
uU8jvLMdATwdQ8g49g0WForJTq6b9n/mz1dyoOGgg+Ez+ua8kCFsS3TVFan1
HUjYlq1dc01tbbRwAMaxf3Fw0VbX/8EXUY6Vr2V15dxAuTRMM17D+1T2dQ4n
Pn1/z9YrM7tt1w5Lbp07SXYxd3qxcm34l+ORj4J8SUeaPp8OsG9sjCgwARuE
1ss6dC0wcpkugxjEqS4odM//YjlnXgl9T7XWgU4BwhdWNedtOVzI1XsxJi3d
EAFKMzx8CjdhXzTv8i7w0NUgimzOmDkXklBg54Qp4nmHx9KsxCFbG36QIB/0
zrjkV5IIXUYvGrBKg3mKwf4cwVMBtWOXE5Bpa22+tiZIBLxI7o5GZX01rqKB
Gnw2Wpl6XT+JPGRn0BMyMzos135xLdj+4JeUYQDSm9mdLGAKMRgjBBH5sgi9
yhAuuiD8e2Mn/75Mmz0nYNAbZNhgAhRdPdOvO/IX54uvQZ7A4sRW4L6kgD3W
9MkPd7Mi9wQ2m3ZqaBAGPo9JNdlqb8xSAhTYMwoUD+UqHm76gNJM1LtEGk4O
6+8vHTx6yo6gc1OtumI26lZtE73oXoTJHDXuyiq6vqrqwrbtF4drR9HDzkyL
Wn7s/sWLdOfaBY5Sn/bWBRasXaOvVarxFdkwpMIxX6Lf7dbUmkN8UbaWp94h
BYpak8EZnEdGknVoDR04Ww8iRO8qRYL4+RNiT6YXa5E1T2/5UcT2WUod9C6A
KoeynDhT7R8TcJ57YLAuUUJGjnPfgoC8QKuWKH/cd8nkTzOlWZNyb0bGAGKx
vOaHb7KrN5IUCuGPKWrkLcX8RGEy+YU9CJSmRFNFNo44jDjnxf8qj0Oqeq49
tdUmwgzOWl7RIbWq0gORtgCJR+jfxX3tpk12A74mFxiW4kdiuomyhmLoPZi0
Fs8kNCoo2ht4K1xoKVJ2JMsoIwvCV1q//yabCPgiCnTCuvgJ8QhVDQBoO79o
KO0Z0w7m40qaA3uUyPpKiRFWqT6Z/OZkw+wwnQM8joxl7cPm+ZTbWYNUsr3T
ukNQhl55G007SWirkhqkg8mJSUUa9QLKL2gZ8COwZeEk9KrxmfndJuOLI8Oq
2UxC4g1KtofMn0xxFJWm9MONsGdz2H24eQKBGS6a14RPkI0670Uszg+Bk727
Sm4WIcIh/CX+2acdoKFT+L0DzzCGnZn2Q6Rzas2XTBMIt9QX88ERDSCwRC04
KLKckEHaOS9mzjh6riGMW32RSLnSz1HlRjJ5QiKqiXhzMLYB3g1J+KOGDaYL
lNsK8fhB2Xo97QHt7nvGMRJkObQ7Bfg7EYqEu3E6aKlt8q4P1SI/eD/s3IiE
baJ6QBpFVh78b2wHRaYQ962BFb84c+SbDPuBn5+qdJMIcAjFbVqYhAGeslLh
GKuZLCcLpoDlDldVZHubCv3V8H5WqGXekn+XdhqeE/e4Gm+3CwSPhTilEu4c
bfGSYar9HWum8ag/AnuoN7OrUnfPzOcXT6xD3OpV5u/jUk7FCHWyP4ifbw+j
KZnhU3e8bFREvqvEOFragI/Z7TM0dA5y7SsAFzld0Q9Ga4griE2KbTuScZPg
+mAW3urPt9YRSIunR2Dn/bQ0iOWdrNDjDQ1sWrIX404D6nvwDBACD771UWdM
4XXIeBn6drF3lRCTSseRMDYYx/el0R3vZhslgajGFyolJcWL+7ggNIBm0EbE
zMglfHos31z/Bxd0+9WqcTwc4uQ/2atkgETkkVRYx3vC5XKisl/o4tepExYC
TOa2CyghFeKgLYXB5R4+EFEITI9oWGjBIRXGQ0KJ/eIwS9m9VKA2rHnQGfA9
mGn4bnJL82Rb+OmvxZDQAVUahlotfc76/+WQ7qZkdZh0MtlhCA+btVbzGWA9
KhAwHSYUHejsxCdwJN04NkFIEXfmUQB49LNlUrUk0OSe4C1ULGpzSpiBhxjX
60HjWsL2yS6Ur673M1C3rsKD3Gd19x/aH8AevOnm3g4lI8AGgyEmN8xL6pZ3
wYjVnw1k1fxVT/7BVY+2Ni7746rBf1awIUTFS5Kn9SKqR+6HQ5OJZ/0zm9r0
Wcwm2zGcXKWla7Cj9ZVOmNd/i9wje7b5JLryINFR3f0/bLvcwsUMR1utboYq
Im47jxl0J7GS7cLa45WYhTIy2jr4+kiAX6AwHndKg2bQLxtw/hFt/Zb9OTFc
IonBxAoz7kIh4RO6aWr9zLgT/b602cqu2WIbLIdS35gsJRw33vFz1yeQc3Tg
F8EdCWL1sNZ/8zqb8/g9StH8miuHjwOqVrJDOLAY+KIy1vqgzOrlyY8UoCsV
qv+wBOOHf9hxMgpu8ZfRlZppYtHXb2cNo17AJsWWwUqZNaOUui9/kwtewbVM
VQIxoB8lh+iXY7ILLNDeZGanvvrfy4N3Xat1H0v/3OPaLk9xlYLiNC41voO+
esyXNnhwAPvNHnxT55nH5udS1UBoLiODSYtdxYZWtBIThxcvXMH4l28hDwkm
bqILkeMurjhkJuSpS/PkGQ/l+vd7Lsg3Gbx8HWo+4X0GTyYVBgUEFpGpQLfP
UDKjqymhUcpR0aP+M5v7eihzZC+g+wvL50lsg69jDd+bbdpCzbljUQBaHIPx
Uas3EDIfxeop3QCS0a46t4U8UM4BcQJ4Im2CQX0/E3Oe4HlqWeReRib0svRY
XDTr1YNTEmyswrBF7+h2Nzug4B9kbNPIT1xgE27CcZuoEQT1i1HQLyAMX8z6
T3tOCY3Rz1bcDQnPvrNXJycIAJolcGEpI5dOoGk64AzVfa4dj5b30JcQ+MwW
U+av1ZruMzZ15X4MEOhmXYL9TazzZ4eSGBgn8B+tBmzgxX1TP/mPK9KsuYKI
Vm7yWG99U4LKIbSFYFS37bEU8nbsN+sAFh21ksoytb2BJxU7pRZaRWNw6b5o
ua/69/2LnCC7sQSZCVhOhAK8N9AXfxPvYKr5s73UgUCU1es3XIL9v7n89WOm
QvO3Z3q5e6Z0re03sEqbn+swRjj0gxCW65HadeehakDQsZFIILK+AP1t/zZk
G4iWB27B/89z3+kZ/cSknV6zeRFEzrqgc4V6FmQyNiNUGK+zK3srpmSrJeoY
d8IieFI84NrnzMsct+Sz3QYZHcUK1Q5QMsGeW2LEOzmsqmv9AgQahBMQxPqT
MjxhXqsWEJJFzxnSUiX+bquWedbB+chCPxJ0lt5ahPbGdccjfXgzgGhKMDJ9
DYpvfb1L78Pc9jX78qacVfDMbglW8PDeaF7+t6/RWsKMH3RoPWndtrPykPXP
v6Nkwe3cyWQFFe4DBxb0BANJHBKTP1HagqAgfKOF6p4mPDWOcVBqheBTGL/P
gGUOnzUUfX0sQirNpBLH+CncDeb88IE/Ubx84lsXhdGKEv5wR4wswrh2u41X
b9lis6QRx/bLrsPCU+oxLI5GT0W6+Pc5mpTe45fPCQ5kBzTAU8oHkGYh5aGc
DxP5AypdxJcQxo1Lk35kDXnhjc1GwPdqNUdw0dkayXCMq2kK1SS6xNx7xK8b
FT+A/BJhjlyyag3PxiYbxEIfo24xWNkF03yt2ov9hgIO5Wgmx3niva0Q/rKh
3HRjPfpLqKrH1M8nxzz/wX9C4u8LCmtjXVtK/9eSYDgUcCkfOyRTOA54tUKB
ektQoqwDUX3GJgqEkPi7TJVS/jMlTpJNjd6wzaCuWZ71jowG4GN7/Y8pP+IH
u7Cw3+5wQ8lIzf2swgBz38Bgyu3dHX3yk3lWq/8TZvyWr6tF0xYH7nT4yigr
jXAJvQXuhGymT0VV4CfRIpvDiw2KG1z/o7YkQSCxDo++zC3tgY9anOLxOQ67
rhTXZ3pRs69QN29iR4jxV0zu6e2xh9qikU8PGziI7LgRFXdV8j+QXdm3nuvY
npAw3sAYdzNQ/djKXH//4jnRSyKF8vbMZF/4ktjqbm+LotAaqce1+OjHWd8x
XCjRZJLvjQhexwAtNCjwqhPp+QbBT2+Ggq/6qyD+vZZgMIaOnImwJeOwxcZz
+dZbuijsgE7f2n/cNhzzOPP5WLTrw5soTYRzvlSMaKo3JwpwYUh7oGh6KUXT
Bt5puMqBZkYIZQesBAhRx+oEWU9tCshrhGxl6VHQ+N2wmjnY+xQAz9Y1QDxk
U7ikC/GyUDTCqCDbkTCIYousTYuq7z7NAoLGCzscZrMg2xDxmbBDCwQvjRjq
/F7+tKrnOkDWYLRGtOd0e9ClZ/Z9JJX6aelMIW4G1KTuWnphDwjdwAmCoTY0
RGMepjUayg20yrZjNT7/CBe8HUNHr0W9pWekIEwjla55fRp5pYAPGl77/pq/
v5jm5+Odl84K6hZUuWIVxFN/tSi3g5MBj4YRh85A6L4+fEkuj09XBMMN55ig
2oJ6rnG9Lch8dVELZAuVd9PrjsPJn5N+mQaZxxtSrK5N6jKdFH9Bw9YUboJ7
E1nCRqBo0DwPOVVEKpzDpIZSabfrKJpTa6oklMGS5nwDYI5nUx8d4agjZKvI
OpH0b7sSmsXFV7YDqLyoxjW1WLHy+lMZsZyav8qMcrE2nUcT/U2HywSOfm3w
YmT2sGzhhde4qoZZuIpH37Ti0K8HGokHNgWtw8bqdvd736QFKN21XxlqRa2W
hv3bOgPR0bxsWcbokjUbIytkM4w1UvrbZwvmCfWSYqVNAH99a45REEt8M/jJ
gW2yYzvQGCaHkypDeZAfD3Tmu1uzLJIUSObKttTPFUzKBdWNpA+zwizn6yWW
V8sS+jcRpW3weFYSX915zgkBfeY1pfbbjdSN50rixOvCQjRwEnPzAS/MdAcq
kWd4ZHJrMugLuo1Xedrn8A3jEceiDaE3lqjFrmOVWnbJvxrOBdIPw65mbvK+
tnlnRa0/o3q5DZdOposZfiX7Lxyx3SxI+ay5e1jVwINjV4uv/dZTivBDOr+h
HZCLIUdBfYjUsTQknuzis5BtO0ZmER7uurx6fT0d8n/bmuFCMFJs3n17wgXJ
b3PKQB3G3Ucm40R+rLs1pQ++WBgJpPN6Nr7kV5EsRXMNM4FDivKms73kJrFS
VpQY8Q9OG3XB5hD15N/yOtVvC2fwNrGSD2FwmZAFWPu7JXRSaKsOrlRbHX7l
mN6FMbZBxrFLVX6niUU7eeWJERD+HVeojRuGDIqHQHGi2SjQGCBO1ygdYD8r
CfvyOxhuErc96Cr5ctKaGbNEQZrfm9GIMhS5hVzldEODw0wkneNPcx+P96WL
xhE1uPjD9xtBfeJNVIwezMDn42s84uKnR2D4tHvpnCTFs6GKENdYGLDK30cF
4G3+PqbhaDO3P6QkqT2nwXej9oF+uITAk0Mya+G7y09+Wr8WDZHJdSow4JZH
3n60r+BuozfXq5hRME2EjfFIxhKbXzDtsDn92RZEC2wEWMN4mBGwSaQNumOu
9LgPXUDXPC2P9i7NZC2ac1HMiQupPFCvxhfPapCfpoDoqt3XNi7YonQdq8H8
ggGgiiQpdSIzpRad9VSsZvzfe3ul/nqWBOmmthwJcnvoIEo4hzdkOtQkwj5+
jES9TYj+6XonZ/v+76hAe+iRLgdPbTi/zkl3AfHhZe2SGq+K6/zxPhXn8TLQ
s5pC/8OlXVRo097YiW1eToOjwhfgD71KVdzqRe3fnwNCUtgaVFRgsqmppR0h
PHzQDSFRYqlMV+1QYa0N8yHDvEYMCG6HACIodtxqraoj3SyULXmVU21vKJ4U
e5qZ1V5K9FUfpcga6WoAwaAEoMmfuU86uT5+L8gfnwZ9/R7K/rCHxaZVknan
KxSNscYTwbNFIr4PIoUJ7DGAfRmFOfCfizChe9el2kjv0TLSCq9ucXcqPKXW
vfA07/J3C8RX6XIBVqEIEX/ioc5/tOZRtcygkE4f1N99cb0q6CR69OSwGJ9J
HNpO3yREURu91ShYkqO4AvkX8Ufcft3C8d4IJdCNPplJlpO24S4+j1SO13xy
/n/1apuRSPlyOoN5qYk5oySi4/L8jYyacRWGirVbrEdsPdsWj+pea5Q5+EAO
QAuGofQ6FUAW7lUHiqhAmr/R46kxuvrV3y/kTT+NtNZvFl18sHaglMfK+syG
pVgNpCZ6a/ucbX+BqOhbLhvzkG4WV9c7AkEFu1WFXqBXvYO6/9ZlB9Q+Rg0c
oUoEsDxG5VRKjWMwWf9h9Z5rhtvyUL7IXcROshIguc7yQI57SL6Vqid3L3ay
sAqzU1hGSlVrK2YFpDMggROSoVmhLqy9sE/j1eZsdz66a+Ef4wrudJVzqbDc
FoHa3Mj8IShRtbqui/ph1/YNpNRIFA5KEPko610ah+ZBEslC5aTeD0TMP+dV
Mw6I8HfKXZTL9tWKdtfRtwyyVKfss/PYCoPuE4mJ/H22AwXHSdOejmWbeCr7
a3ncB17QS1ebmy6ivc/jQ2OiPAE/QcaUcptklq5JXGo5pO8fFGRrU1OHQxLt
1T6WxiF1EFIY8Z7akRXVSVkFH4ax1vtRsIekIOHNmdpRfAOWfUyOqTxq2gEA
V5LuMZXhe98YX0HfVAkxPC7yLzeeyMaZScv7awBI8KNJlDNgnYjUpElqXAVn
gQThiaweAk1p88Sb9I8RlhOYRZ5ih9x+j3TytBx7GuQhFoO/+mr8yUPC9mLX
+wvVmwO8L+ZHjmZiSBpvC2CRw12DnmpFCX+ukL4gw1aVCuIGvxtSLCyj0vs5
G882rFuaUJLzQR5vDLJcDNHtHrYdyI8a6EPXF6ZFN6u6Taa2/GC+KCf6sKbA
Kc4CFObeHn0EvE1HFNL4IOrV4dF1jL6b1vA7Z2LF0JmOLdjqR5vr9kKP1yv+
TArPPOOrRIH8W1XHb65mO6/31ZQIc4RZqCh+Fj9OOpL/ztC+MGbSmrAQ6+cS
gTON05Eqi5iIwNSjYp0bIW0VJP4kIZWBCXilJDaNfgxsOQBKXVx2U2W7W0r3
YMTCKPy0Wo1BlOxfSkYCcD4tKTXWD0cwsurUmeK3nNrfZYF7Uv16d205Jc2v
HS+hzGbaSZTibudz6Drv0QCMZFjFA0PMNDokTlkiSRPxVVmPOm++cnF2lO9h
i+UiwcUuoV22pW5zILgyRfjqTzOXB6/0jFj3IrKAuw7ieTylRgx0ZAbJmHO0
SeCnOySrhjzJ1esGitOwMO0fdmtgh4e2eL+RTX6JvIfkwHzrpjmbVzsJfQuD
yEbTY6XD3X9Cg2jHejJtbZdv4M3m916Gy4+iFMRRDKklQPR0QC5FqJtT0zOC
FQaGd9fs10DxVENv15ipE1CIXlKglIuFvpmEOjSgW2z4ZEslq6l523UO6cLn
/E2AOp845amFkTDHWeKfl9FoV04LgCvbiuIXFAoYqeIUpUcJSNeYVLg8mETB
AdNG5wKb0GbLbqvI/T3W6ziDN8o2NFggaB+ZqbppohU4dE2oF1R+d37j2+Oh
02RRFd3FOAq6eH1Sm9X0EJjen2Qi4Dmd+Ppqe0l838A2+rzM7ti8jDsabSo4
mvTK8d/2KSc5+PGcxLbG2y4qTNOI7qEfzUNSgDavZW4m4R0eMd1itYdRdX31
FOc49PWfgen9tyCdweS95UDubndhyvoNq7AZ8m25O5H/hbvORFFHTvdfzFPk
B2zEiYk1FSV8K/f3NSb3iXHTVGlnMck6QjV6i6+RbgitIv/AdzrlB7BH65Li
8pCNLkmsfETXEFStq6T0hE27HiG7CncEmh21MjLr1vCvLJsgn5lsd14vgaT4
zd4QAVN0xGK8FJ5cpu4noBCAeQOW6uwES8SJn8P/L6lvcIz2LyqOduuwpmvn
Q5IQ5WBP9c5UW6t++sb/iGPXKJ3Lbj2Ix8Gq7Adb3OHXxHXGkchOQMiLS2nm
QF8mS8rVInNTUW1f1XxCybGkiz4U5WjN47WNPhoKslrKob+7qSt6yAgYW+Ee
4VHZ/BqQrE/FE+TRaSt5fSVYMVz9dchoJr5LAocw12F2sirK9/ZbEffGCJ53
8saC7Fq1tjnOk9lHrNz1gwG3AIjECYf6aK5GviU5oBJXxhsrA9v4w8cJQ5/R
TELYigFBLz+Az2r+7wQHFVrjxqvz6fF+A26tTVSBYsqIbDyCBIYHVJ6u99Fu
y4fnl2WZ7yrKshY/nxvw8uwEJcXj5By5OVREQyjDMUFWbThPqz0VwaT/WeiH
yKKCENtGZKHic3pEFrvzjybYtUxZ8OsrRZBPCPkDwaUik0l5Y1Mw+x1zCrWB
g3ddQ9+UC5Xjgx4HZzrXN8nr3xQazmg57wDCIrg+iHgd10fPpVOKK9Ueyg5H
s8E2XiB0/7R4mydARC3tAsQAVAgBn0hOcxCFZLyVeBojU1pjMbg/oy44R0RI
j/cCXJYhTwIDIwDAe9wJIoI8ln866AwRZ/WXtc6vnczm7qPLo1IJ+m/6Hgc3
sp3/JHWwupOodvlFU2uWEfLeDhQIplBg8LR8AdvxmaXX10QBp9EhLpDstdgC
yDFsF6K8sqHe3FyrX7xagJSinDpcWQHJh3LjQwZMF66kCxicSXJHYHy7h6yt
tL+yWPJu7NftNhl5kCIRDjdcDun1kQMatmKOVuyxzcThbYNwWrvg+gDdsemA
7c+ldrBvALV/gWe5gsGuhq30Y8eOvXbRapu8HCXPI0t2Kil8z3XwRnHsEX66
2osoNi0CewkKLJ4VOPTdCqsyPAD5Tujik8+SKtkYmvxnZddzStQZW+ClpXtX
tQYv8eO2U0kc6bURbA9yTQ3PWfmvlZhGiLHY+fAhoxvf2zFa1z/Hk3204Cd/
hOl4au3ov26Ih9V0MMz0CbAE/xDLOoCFGI5ML/METSFmCFS+Dmxe/f+XLbCh
FqSo8BBOphElUF0d/JR/qWRfHxx5yrJWrFI3LVT8NqFsu7SkKd+SY2ELl6mY
HAWmiClfkZuBo/zVY1SObGXQL6Mt1j0LxL+Xooz1SFdFvg4o8zi0VC+HRyu6
sSWtEVprXnWaztm8NC/pT1Jm80lShBv+x8eb+bc+JJEvKA97VUmlA3fEw282
IkPobJMgS/3jwU6lZrznk8EHSi92Q47wHcrrjepMB/W4se9MpknIiwYFkH9X
lfCr5H84VDAUzRhoGASwg9vDc4yqnMoQlYDrweLLxQb1HmYNTkWnN+PrCxGj
8F/1o4WReQQ3Mr+NSIrnMuYzjJ2vUTdwxiLX5U/vcB3pAUHFMjE3lKP5etCp
+aMjEdgjKaWD1ynH+LTA9/yg1I2CKmGyf6VTMn8dTSoUrS6QnsXEf2gOBinW
KNBUQzmg74Py5MQpFblIMVrNp5RWz4oCmn5pytVzwEoqHua34kE0gZPpBoRW
XkloVqViKoQGQTzxyHCqwMat9GOPbOnQPA/vMnYiOLYkSI6CCff6uDgsTYpt
oRhOsfklWmK3xtRYJHcZCUu9JdrMAAMzyISigUkHinPzsBQ0w3r5CNuclzfk
FEf4KPVBOMMIdAI2/ODWyftocizUGSGBmE7CpNI8Gwwgc1MR7gAhSK+AVoGR
/hmh0Zr7NIqWcxmESJyxLjxOLKCGqzriatGMf2omRjd6imLhVBcauwveqgjO
tmUlGVaHTs+mLA41ncyGN9VpNloYpyo73+HlBOSPK/OrzJiHdyVZWwnvCcCG
o6Mc9WFG5gRDliRvfca5sXLJlxCO3Kva3GxWca9FUOBxHWfK3Z3259wmZbxf
5GpSLq0YUzf8dtlhbayRjOBC0/e5GSqw9Hfyf+CHctvYls2Npm14cqyTMZlc
MBxihl/BQ0XlAwjs/tZSaRXBlujjeFXHqFRlcxvZu9k/zxbRlS9MZw0/lgue
0rTw4em3nCRno4fBVL6kmQqCcNTiVGLR81hJ6pthafuz6Y3ct664mIYIRNWq
pYfSFT/5RMElsaru60hqxzmNhn+ycVU1poh2irufsvzHyWlFblE5U9pU5DXX
KOyTfKdUAjnfv4tsxrV5cAfE9yTBpf8JY+RLaHYytJwUUnUtu/KQtWpViIlY
AIPRVQCRQg+e0ii5aEgCsmpCM391NvCNmo3Ub3gk1s1WNH6+xuaRvXeKMkta
3R8alSOqtzEBvRyJUL2TzS9zFS9KSLfrOBtFtdsR5AhNx3t1da9duEAGe6p2
8rU8XMZFeOFBgjKihh2T0CrLhQMpVFHGiVEFqXHB5WRQyi8qkUO5buwuLfd4
hLFnFDy/pjf4AptPrFkWbt+dmLSdW2UTZX3FhALDBk+JW8GfUpik7CrhOjBR
TBnYk0oHU3nrpfqSQogBvQGLXmSWJThYbqlqm3bp+i6qxZ2pkOgH5SdqxeaV
hptkqQ9MJuK8KBxb8usyeKHcRBeZm3fmlea/6OAAEG7d10vPBqa8PDwacRRc
x8NsJ4uksrG/QCKBjEJ+5zAVGQ4Zlu/oP74D6WRLdyVDpVLzZyhmD7m/wNVf
v7I95RUcuwJu+M740emTpnciwnJalyU4i1IgglJYkzTsR51NKbfmpj2ag9aV
fycljII72Xr+M/P/9C5E+LjgXaM6QdLkncFM4C9yYjg8luaIBjAMpePod7xA
hxYCr5pFSKSxFw4B0x911rUaNMtirL5QkZE1TN5d7etd2H91jnjn453OR5Ns
8MsXUZNHrp7OttpJNjZg0mxenvOODQQlcufziAkXcTeBdZkrG7r2sjjgtwsf
EvFq8nzoIsLvxZ/CIdcHxGoZF6/kbxH4kAn2G6GCrDRfGLNsm7udXcelg2HL
CuGHoDTjqiOyvcfMEuD7R8kGb1UBc8epuSI7eQWn2DTJNsRK6QtWkNTF8NjZ
uqs+qm/V/opw/XEhh8pLkF2AlYo/K/1s/og7SyCgA669eA5r20bG8VUJrks9
FnDzFovsTZKmNJSdL+DydiQEc+gIfs+22j+kfiqdQzxvsH5XEtSv4lEEdCl/
JCFdI+MGPsazxc8GPz/yInIVQ9i5hgvoKnucw851HHktZbUhmLUUcyxbAyx7
K/bdAPCFq0dcRMsiOtBeQxvYonQ/nFBwDqpPYjk/N2te8NHZAadolYNWQfJB
9WaARh4sxUPqYEfYblYOC69BBwzBkMASr5uNW6o5yfimrh3sQmILZ9FxySoa
rSczpQ2sUl7tlhKKNYw015ZQ/azWiBEI/TIZE0sfKMwxXjVLZJdyTWpjgH18
U5Vv2p7Z+8tPLGyPBiyK2sOfmXd/QlKZb4Vvprbnl3E+mPyyQEmBlWwwXilA
QTL4OevL3PAtshnTHOWO9FlHWabGE6sJ9EDMyXOOdbfP0o62PO8CpK2mQ5+4
jZsf5G3KCEnDpE/rVChX0SGYmW9gNTXto7NpFAt2XrDF7y11llPnYQsk2tpm
ABdmd/yCA90Sc9F4zjgR9CV9HV0S1gZ72dRyuQjouIakqD0mSJcZ/xss5ygM
qaiT/Plx2hPdFKanuRgn9rm+mOdUTTcsnMipyHCjaxmKZSH6on5G9qXRd4JZ
Uk7QcaKQixpkSi3J2Itk8Uyt3moi6KVKuLtQ/ljC7xHgvbotsgPWLxlXU9Jg
IKEbNKnk52L0DjaiHL9ziiiWz7c3hAKL9WRimTZB3eWLTXlD2O253vLAA6VO
1AVEN6u9IvSreRUqagn2HPg9CaFhACZQ5oTYB0JIRe2L1wvsGSJ0kBmCqisJ
P0VVS6YzyQXanzyGncBw2IA4Lg9OJEGni6J+L6YUoi3p8UfvDgI3Kt158y2W
JSk3NLS6qchWt6qVfrMe+1jc7akSs+HZcD2IkdAPvP0IsbNVRdsxVRmtE0G0
GcWR2Y7YH7NDmLtPRUIARur1ya7O6AbusSMpi6qbUQ5luMtbXEJIK83Vg0bS
aC8/jDu5SGX1vad6oT+7et/0kHnkdcgkSZWXNfHQ2MxDkoMfF7cFUuFFFHjk
xMkdnrWgfQV+eOx2K6cceqHZfv1F9SPltfxoPRVMp1ie7xLHwaFstHlG5tMm
vUXMMXDeHUZp+xPoDEqzA1D7VEXD8pGfjkfW0W3ZhyP//h2vIKSFyWkJXRvU
snz11zgEdFTliJsrYfJQszQf1rVAy/uNUYTlLE7emHpjGCBt4YiR/GFWAKKg
WYY3y1N7une/VGCe5pKvDQqU1IQsJUgxXAFVAsZ5vYymgNnXURc4LJTDO2ur
8eaNbTjZxcAmQKmvdbVovbahkprv2ACUe/nt4YoNq0DixcsPWDnyPUJuFoud
w4N6C66O0oQdI+E9Jbo6LgtgpMs4MTXQmsVP8YUgvQmOyBFYyeoCRfZ6i697
TfwC1ChNpjJ2WuKjrEvBFf2u1/rijaWN4WB8sTQjyS9mD3CONXcW7E3eLW+X
S60GCPjy8PLCJbt3Plh/K0clTQ2i0CvmZFDAAQi2QUObBuUJDQKp8Id7brSH
SfSoyQvYhRN1G2I5ldvU0lZQ1Urzzg/vYzbQln4r2evYMNR9ievGfnat7fWh
TShfABhj7vjkRX2fNuc6yo0jKb2uKWXvcyFYOsxkO8fwW4xHsWujeqV9xg/O
P19plzS+0eePROb3yBF+T6jZGTcQ63UW7bjiuqE07hs7WsdcvRr8uHVae7Cm
RG3XH+NM5Nam1sRe4GSolIfQkOt4/JSjt6zAEdwYl2FRHILbr/bPescy0zqA
zQTgQ92gr0M9h9jyFU9RL1U2NJaiCAVQ94ggeMpzTbxaMqcGRCNd9+9aV1yL
9fjprNkJ7WFxME/goNh6xDey5ZcwDcjXrTEiaftikabl99w7Ysp/JXpSHSDT
plU2NQxqK+80loVa4RmhHaDidu5dsvbFM5+gU/MogE7g6BKA/QtvxgmF2w6b
Z1n/FgV0FjeHoUQaBcQKHP8AktMNr0xmahHv/XBBz+eIgiYXqPDZr5fwHREu
+gAsZhEaDO9dqb4t5E118yaTLpU26bfPzjiFiNf6ocLFsEmUGIT1zsyYIBEq
ZhxJ76Feq39+jjrAAXJ52Uat89XjMWOqPjLOw8evSP2JwmT7ulF/aQzcSJoZ
8199f+8dpQB4sCwDsG7bC+23G9m6bofH4XnNMrGj/iSRPKVAZmTUil+8s3nU
2GYo6tOejSuSjhfafjF1kMSA2+PVYlDBJ04jDDtCGtGZTwzE2v4ulS7sVpno
QoVMtN8dw/lxkPm1A1pQ+Ap9oS2pQ2K+dFj2bdqJ9GplISsSF8K2yXGnzksX
Mxsus6/AlYKIahv3D66UYzIYtB7b9GqgJ6prnQfM6oGkWfp5QcGHV/23FPWP
fc07uqM8cf58i08b7ifDqMo/210m78fv697F+D9wdk0P7yetEdLJ4wzP2q0w
ezLLBh97bzKhtkxeZc5RQyq9LyiAWln+Bg35PwkjxGw2p8kJ9o+NllD3fHSm
qdnaWg/kkh/hSXkRC1sRvhXMi7NnoS2FFT/QTdBNFaJ0NZQqhnbAYI3vNRt+
sUEvUxk7h6OuzH5VsP92cx0oyFtkef0aLF479+KCPahGv+FtdmtqAiUUHqBo
tnHf6pZ7oVercl+W1alVXDGEkCKeO6gl0dw+xNeAIT8aw8/Pm7ZIXgojR9Po
RJQ3eor5D/OWkDsa5zfBTXrmFO3U7olYMCFFUYlOIf+kwGUDRSykw87e/aXw
2p2EIS+y1cgFext+oLT9JKhAnN/jQxr5V0ehA4br41QZ6CRy6+7DCzLqymfN
0/CBSHyH5WKYSMQkEqNenqcI1oRhdmENXH26nF5LlTXGi8/LDHCGPiImCggC
rsH8AL1RBSTujP/CaIb8ITFSmD68dn7gwqxwipMfkMuvwl3oqCL9mHRsVm3i
w139me5+bum2n7EE/Y/KDdJLp6D7LRb/Ug2AGfdBOrp9hxcUCd56YWm7ywCE
Dp+cuDPajfi/KnNe1BUvAVJlrXQKWqWG+8sAaR7urYkrHGFdiCbz5UMMrNzO
yNJi9r5hSugjoHSYfuIzxMRCp7o/7KgR8lfbr887O69cNEQX/xKtPgbY0eKm
8ItxDCnim98zNRvRSlJ1LbXW/OUBS4tvN4ZyUfQeunJvrJpPkV/pn99bFKak
f/RdQjd5QDSV/uqtEKqu+nuGvEd9tpCEkP4R4rrEDZOTHTLNvUhTGepAWRoE
nvP7Fqe/c5PZkDAEzyYxhfcx5ScCcrcgQ4BkZEMW8JGnOzUql9dHc/rzdQbI
EPlzBTfEEU2JOz1nqqZZEuUlhqj6oc/oRiELvswJPr4ZitWu1IgmpselOwyY
ykWwcR0nxzAVKPl03WCtLaSF4Ows4cEKN4an2pW0yRVPXz/F1S98Dlo32TtK
4dm9NUMffMxLEGeB9XhvY6dzK2p3Ve1sTNjOj1GS/s8Qv1r6qwpZkIOrIJOO
Ve+gfQ6WBWkDrbQUt6aoOPqmojMk8M3xaybbfuNqemkE67aQFOd6cPzW3RlJ
kFil8VYwOVQ1G4WMblVAr8pqwszH6J8WWs70lY+xC6VeJrbBk++X/BX+9xSU
LjAHcRxoq4sE/KM7utkynS/o9hQPnqr16KF4tLYRVQOq8ZJDs8cRnK/u6Xdo
E6sy1SvudtTu/kaBS3ySWLXTSxEy6Zqz5HdVyldslxreN0r33GOIX+feRVF4
7b15RfnBpWFlokihUEP3VJlV/U9pk96QvuEAu229I0bmO++JjVvWTU2P1ZlM
FQ8W+FoBz570rQe02difEGTO4LjDEp2qoUFAUN9QGFPJmNWuU90iWQEL/zhn
0OGpKZWw3qxi5Gik0EgMg2jB7gWjBjYejJDDHK2caL/XrVM2eBEyCj6+sMzX
ptie+A9vN1IymEvrHLqyU7vexKAoFUIvH9lJxV9ErNNJZz4iPZUeDDLv0hLE
FZQ4kncOXsICTegjq0fpNL6WCuq7Xgc3kyrSGYQ8Rg1YKGVHLpf4idVo2RoY
6WIHs+5CT5ga2kqoDYSVN85SuasDOqe9BdmTZX8tXgynC4/0D9ark1OhjLxP
6+CN5Ti6bJKIOWX6+pyeIWhG6e+jeZG+oQWS/26LFfDT/Ez9vY+KL7YDsuyS
EuI9EPGD/8KAAkFJGX0JBzGibQDBjVCpsXTOhCE0bgRzMMJQzo+mLi5Pvh4H
9fH5baxGK7WX2CfdDH373bO8+XSJ7BOyVClbsUVK+KqpN/j+OPowaMBcZ7os
Tpzp2PU8O7gfh+ulIz8pFR76g6Dg6Zqs5rjHVqyjDmWqc5z+Ya/PP0XiaVJS
iYMtLZ6R0MwW/oPLQRWGbXLbf4VnxkIIUQJkp7PIaHdqV4xUCtZ90qR8BtAJ
gt8tFS1fd2Oyu9g/v5+i3xfnB+YwYy1ixogYaiRug5P8R6GSAAXsvjAnHcpb
9SFiRuJgkxBjpYPusMVZZ/BePMW/30N3XaVbnHdtpeUDW49yyzNNj0d6CQtq
NYjP/VSvpcnY/E6geGewvupfculssS7lPid9wvPKOdPCcG0IgPe/UrvClcLi
ifXbgwsN+kfFwgv8Fgsmd3GcpiAJtVbOd5mqQa8Q8aAW89DbLxRRdaBRT2f3
o8++8oe3yeyYyiE6sgR4kc7dWrpe80w9cIb8MzB8H8QOpxVioiKVilnAOK3m
qRn62kSnM6Fo4TTBeq49AHExZHfZZTwxvH+MyEz0VV2W3yN0lVsw4z6GvENj
dx2kveSDnrkwTimXEhJteuMYl/5xJ/LSt2xbWlQnP/cniR4YymyFEChws2/D
KFKoVbrxi6FMkcMQ5FhJWiuOINY41gR1kymXGVCykJgEdoh248+Ohz5beoXu
XvqU4rEmII7tJqxpXFUY/SQjbfywTPpu9wOYRTTjLxXPLFV935LbP9b88lXh
GLqsqZqjtY8rGFoj4ocJ4scpG1xSSw1jfDybUABPpVjUbLsvDnIm3zY69w8m
oEdunp8oMXFlvC/Ql+XpFADWA/jSQdjoIBWrdgQOYRCFHaf/PipM1aJ8Qq5A
8axcY2L2ruSsRLJk53ThavHnfY4lCSZimcZ3HteuX6NPw/iL0+8vJSBIGnu1
pmvApfj986/dltKLSQk3+hfDbFat57VtkrKc5KHQOEW/Yy30vMsGYxCZS9be
YayzB9TpPOzlRexMXwXOe579FiL3ldazjqLExz2RFLRpd+2Sw1zobHyLmmEM
cuNMzEwjqGus3rdKLVaE8KpaeRvBS1qzovapcENaMQi2fEz4MFlJ1vuBCFap
OaMiCMsJuHtaZYNx/9KWf94XfWRM6g4OzBsZ7kbN/TCk0Q57PkGUktbO+s5o
FkKKYHAEOFnuIrvgu//NfwesS8ERfiEyvdwuSgHnYncjWRwwZO+Axh/2cJhv
XawGsQ6N9VNuA94gmw5MZb/dBLvvrwR9kB/fukw2TpMY6lknbRTLsuJYWTgu
GQKGdRYTghg8mansfeppJDI47nYiFIkZoEHu5nvHE79QLV12B+fBTLSbkhnO
0fZm2b3pZFbZ4cUM/r8vR+z+rFUraL5+jC8Vjm7s182MP8SKSLXwJl+Noae2
N1UsDnm7Qim7Tjly5MmA0RC6C/el12nzoEuY91QilaBm9VpECYD38KZGWHhZ
HHaOHi1Tr1vHK03k5W10anafbDzI7hftvfkT0XMZxa3SEijRgGbkYGE9BqRG
iVuZIXvtc6+BKfvxIop+wWN0u7AAElUQIRq+mei/MhyFYPOZ4YN99kBkoAvO
sKU0f3Pn6xh0E+iOnXZOEyL/JcpLq4n2WrTf7OXbMisQopzFl/uzh/uQLc99
J4LG30+MvDDEGPp4+YYX0Z9CZqu6AQvQx+Rm86BoGnQXJWt2EN/ZjB2bsAv7
V7wefmEtVr/cA6UuzYlxh2f15OXnImmHSdy4HvvtgkXNhQZpHplGjq16eZRw
RXbQJVAH4EikE1+3qYC3a4Vk+1GJhsp3FZWtH1V6egETZgSPL0AoUsr2rpN+
JkhCp5wL68LHMf6ABa0C6AguvO9lew5vBvLahCpxNnbC13hQVtBvkiYtzG22
QV1qMKfe/BiKNIRjcwjrWo9qW1aC5TedP5dNE/Orq8g21sWkTBEYqqPfIeqr
Ydt4WMoJpiZNMNp8ZFFuFMk0t1yHxi83hSP/WPyX6QOVAOy2+m6jXCwLfNFD
0KRYUJeYW90VV3FI/MoVE2wkTFblFnHvOnBlD0oSm2zLh4/aW9q/eMlzHyl3
j9Th0iqnaj59gSCSCt0I7+Ncj87i5l3oYfqV3zjM+d9QPdJSFjZPJDrACUdX
DrSmgWOnuFb9moJ+oKCMgEg2EDpDbilwlYnSH3gReHLi1UbcN36KkKA+fjLk
Dr0NNsR7R5ZRqgHmbnO4NFGrqOgGKSN2wKzm9uEgJGE/S8OIz+4BXacjbDpZ
85rpAhLE62QZcmYGNakIPYElif2XpaDTvFsX23c6nQvL2v4zRJAZnfrlgXK5
QJKRPmEUx7MSICKuLVYsvH2LenqZ/N1wVQ8s6IA/LJRK+6UmocWcymXqVZh1
FvbnRZJnWLr1/2kTsIzKDCPzI9W+m+VXpn6RtTiahadrLyvx79LUfOvDxmXM
ZFh54KRL9k7tC7tJkruN18YmtqG46EEYjBPZ7DBcIgQaztn1r2UaJwB8hgkg
XTy+nFCQVCHXraTKiwQEorLvjsRiBz7brtJRuR8Q511I5O88/FI0TKtMO9br
Ab/jZzxcZIAlTFJ7TKAhRTZfiF1/DCOQNhYF1G9OBYcdj6W2uLzejZpcN0d2
NXRB5eKx3DeAN6u+geV2zokJZsjUjXwDewcqCbtARn/d9axkFNVl4FZV5MD6
STkmy7vC1htSb+pKtNiwz/8X7qQw9S3S50imMk8d2fIPk0RBibWFsv7UzgGA
5OSqj5/WxpJLtN5Q2I0BxosQe7bekQkqnSJ5vHs0X3DJYaAwuKPePg8bC/tp
GvVQMNCgf1L4NF045IklYpIYANWO5tcKNye4es4xLxw/mEtk0gk55/IzMQdb
m5RUt390Uu8YqN4nH2g6fLYrx9S9a0RwsycmjGnS9d2KbsTcca4WqN4RCFzZ
/PjIvKzJ/5FqF7V8KX4Y8NGKp9OGDRYOBfCEG9R8Gkhjq8BPnLpQ6oJqi/mC
ik51W6hIYnvrpxfEKNxCaa0C7DiS84JFRvqgR/prXbxbFSOsVPets81xTurb
WOVm7Qu0ApzWIydRHsIHopvDXVYJZ/J3BBgbFa9ZElrI5ApHASDKPuBEsAf7
LxE36CLTW/8RctFbc72/96XBi75VuvL5ZKgWW05K/ns9SPemVB1i/FytNcR7
oim+yoxSO38+WLx9aqOiPwXk0TpasK3mC2qv2I826DcY0pJ1aUAc7uxtbgXk
TYnARp50Xp7cdtDY7s4VqgJZruQF8sszpqiIAEu726oVITZgLp0omEa4e9wN
rYz57zVG/RMiaYD7G0RTKgAOa+dtvZQDHdWeRDARB9X3EFm2Zfsj3sznUk96
gg+hFijP6EpI55Q8aFZ5jMGQ8wa7bvtpdWNXhwtyic9+7EaX7PGYArTwSZEd
wtuyiyqEqhkyF/1wPkVRZKIIYGkIrOFjLWT4ySzwi7JII7vHN7IUg77kgPuB
qu7mHcv3SnCyohaD/YxbRZ4NoI7VOUTykhxIabu2Tx6eCyrJ20ADgH6ld4tY
tOZotCD8ztzQVEPmNd3Qu7g2N/qs0PXRKwsB0dG4iqUQStDmuuP80wi6PueU
aOA7UgWDvIigfXM9VTJ787kkArwEVcMKQNlgu+X4W71aPdG+mbW4xNTFpO+H
vYNTNpP6F7+BlI50hGyUAdWPCW0fStHaTX03u+2UaduA9Pw7zYtB0oYeFlSZ
zymr11YmnZyLtq0oZHY29k9xA2QsR91s7fX/WcAgiV8cKp+81ygT3NkvAmlv
7+8F724+iru+jh6pa3c8eSrJz9unuJZ5dX+8dYxnUA1Id2p8ZSNsRo4i4hq5
9rDPW9eIC0mD4qMwob8A3/hrLr6eWyuU2KOG2eGkEImdXCNK87A056YVe4+I
eidflBCFiBmlcK8hu2BjanoSQUn94F23vPPJi/WeawxX/tTZYpTktyCnRpFa
K5BFaDdYTh+gZB0OGnAijXugsHN6Wqynze/StbNsbXrBshrihKktV8Aqh6rE
IDg2nP6X2Z4d5m47EtcAdBP0vF1EJNuRYh+ZTlJE6fyjDpcOUFVtaxBy+tP9
RXw72G7pPUIFzJ34ahmjpcEc2lPUCzit1JICVFVqgS4ZN4eRrq4xqKL3Q4WT
QK0dT3V5UujW4XKUmvXLNGAbTmcjMy7T7QKt+ZfA9KMOUWcu3ANHxey/JOwL
XD7HAaTEJ7mA61KEtoE/81A+QIjR0iiFbZsAbxZ4KOk/JBXXnibWbMx/7G7E
55EmP1TaWBpLMk6LtrMciLK3/GP+hFm2XQnLzasE6VOKKUOibxVTF2HnvTGS
e1Z4UGcuRxVwm+WBJ2B47mIPVBeLsY4GJo5s+9nm/QCNRn8wpyn748YQX7gd
2jUzjI4/wYtp5QWtOeaP/nufoLBQBwbo3xi/nbntznE6+nViHXoeOQgUD7bh
lFqFxZPCIZ84MPBqCh3re4KT1CirZznfJSkJwaxpU+G1bRIsIdNYABlVh310
70Q4GOYTWDZYqf2iF9pNzH738qi04/BHPZdT1coG8VR6pN0uWfr90eWODRDP
gf9IBUtjG/vGnauXnocQsGLz9GQcJLVmlZ/p4PK/gFOFyYviyhjSc+JjO6mT
8i+DinfI9U4znIkeQpDI78DmmzF9KLkTOgoauc3AGz5c1Y2tgv532C9suWpX
ib6fIQXlrYBHp4GXwby+PESC5OEU9tIO2OAIh21OpW92F/mriTxQcDiccb+u
XZFsvmzjYo23cIAGocZ8pu6h1UXetssPD5v5yZT32t7tua3qOEqSBlKWFQyy
TI5bK8Q6axLq8HEh7wViijj5VOXQLBURAnaAaV9IpTDTCvcnVJJnCdidNpy0
H31HbELevpKQcxf2+QieRzjQtXz4XBDl6Ki7KXiNbpX1JJDfU3Co8tIU4Rdr
oIe/iRw7hfwG5tR29f3HHKNLJbl1YKyG7COm1RhIAZKUv/8xq9hoR1o7Y76C
a6q2BUjev+2t9ru2st7/kZbk9OyB4SHalOXMiMS1rZgZo3iOJCtc4wBQ1bXb
vHrwF30doeYmUnWixVua+HIKTSKe9brOLY0ZEGeQ5PEmniaB3h3nsluedlms
p8keG0lsuO8IyzU8k9BM+V7Qh+m3b6g94rElV2V+YpnFks/fISQEukp6WEfD
ORDlWzigBbGzKU1fZwl1XvVr3++78OWaOHp72FacrIhFxu/IsxEoQ9Dh1E6e
m/7fghwN1F3VSf0kU/s3o/pRYhWl++QCbH2U0wnpaP8+mFx5B/TTn3P5G+ze
1XZJOlNgEKn6D0TfLzKjCrRRn3WY2UE1ZJmnav6wJMSK7xqq++62JP5quFln
a+zpv9krax1br8Ku2E//SQAZ29lUx1uYATUyfxOWQU+7OIlogQbn8ckZfOmj
1b4fqNVMdYRDXBJZMHgashDl34Ky2w35h4K/sLC0OEHrA566iz2/DjxsLvdo
imUon0bFoREJfiviP0vrs80y6nx+cyf6GEm6zmS2HVFrM8BtvFZ7fCaZJCb2
jXcZBy5NplxeJoFjDxcJ0Vu/qFRlD28IrKi1flrTsbgARa0hO3B/XN6Wu6hF
kK8EIC3axW8NmOjvI09LGhyxo0Wj1lj4eB5h6ma6NysBgpfWfszf6oCul3pg
Rk8C4fI3t4zoQgJGpkpfMa7jqqXCKBZiEE3JqQMjnJz07W1Yff70aNBAtTj7
nQrATS8Vz35NJ0+Yimr/SllCnB6c+osy15d1mhvxtKnnPWsq0BDPPm0oit6j
yWS4OlV3f/q+SgdT+sPEwUpUN1QJYYS0ArmnydHtMjCoQa66EVCerVLWPOdM
p/6glA7+arKXif/XPbBqtnmggOktC+ySTg/Tkw5zRKnp15uXA4WIZM0KASwq
9R7Sgh6bP8WYkulzklZMAs2wXL1KskNvKDkspXZbhtN0SMlzues6l1Y0dkqm
PWJEx8942y0AN8pVcc8CDhR3EqaPqnTUjtOpaQdu0mvVKL6wEws0IF+Bmifd
Po67FxK1l43GfS0WxtrBJQJB6oKYnrYXaii13oZyw5nTmgEDHUrtzyM5M1Cq
PsN83ErUIUnVm8DNr6forHkTwbWRA8484uPSKo5UKca8ffz7aYhtGt+Sb3Bb
vwYltLCCWXVhdcQWJRbTqXO29eS6WUDb/ci1GBoIfZ2b8co231qBmW2tdvVY
M8s5jp/iHB4EU0KcTzL4RXmWnGwACi+DPSAxpItNEQX9rO0bcqMJHGqZqpv6
b0kUvx4HrJQKGie+wNlhSWytmBMYIJ/lyKvti8jnJgq6ghDg7oMExIZPNTho
4H34eJ0OENL5tBst+UmpNAv7/BhKfkR/VtKMOOGDtpgL0RzJch2gM2jmGA7+
G04Swxo92mTk/Ll6x33UZy1RHM9kwf+OmcwNBJIoc5iQg3w/K/1vzlzErRDG
2MHCoihN2Hf3CS6DVjSv5DyG51SjOJ56uaZiGTCRpmk7p+J7EAbbyMwfpsbD
H6Vsss4U/VtzSWAUdKRCPaaMK7rWduiXpAJpKLzclDL6czYQQbeN2ZZB5Hld
e+ZxWta0gYG/M3rAV9u8QAigvvZbZ8qKNDj9whf3oibMwvIjM4W2KR1pbpvg
nAXgVAMPXRXMBND4uT+knFiIlJFYwB8hoLebhjfMf1l/N6XipEpk8TsscDGY
Dvdw1M8JI2nlV9t2Jmmn8T9Yb7Re594LWiM8jT/WBUr+35pxjhIy+E7xjPLA
esIsPJON7jcCSHKO4ctHLGb16IE1Tg4AlTuIRrrZ8zXT0VtSkhdaEGPQUVBh
jUNdbd4j/2PK2oB8AQWKqSDmEhVRD+gmOydckXWAiZfrVoAx3DSXj1z8hMCX
VYehfPHPszTgaCxMazMWmT0m5fC3SodPVg/YHahnr88Fyp1QAfvTDB62NPlr
OSxfbubt7qE5TM2lbvvrrAPlFvD1PTWoss3d689FhTAGhwnaNfGrzo2am92r
mHGUFW1yhBPuRF27LJdWbUzAqsvjMZptJj1CMvFsyYAPzHdp6/FWagAN1wyh
GihJFXhfV3KWTzdETOmTii/iHGs6BpJr0pQWL+yCWztczrg+YLg+5HMo+fF3
zJk+SjIovY2pT8wSImTIg989t4Yv3c2SQFOb2irzlJcAkhoOpeCNwSaJsaFP
Ka4nwPiIcZHZx3GjjdzPCnyE2EoKey4SU2jfso8SISK0ogNbEiVn8fpsJQkl
ID5gVP+0QalWMOQobS4ItMo966DMzMdUvRg064roYU6W8YPyTBEN1GhWVxK3
DUYn11mRFedHo8ISjK0dh6NEaqLzkB8Hb27n7tLGnLQXmDC68LUsbKAIRbBJ
HHkGurCdILyGFfITxLssmjbg9cN0v9k4XBYitSI9N4JOiJMhlolPoAaS9KZq
PgsCDVPtuPZQANlXM9rpBJe6QBGWPz/7fyzNVu8zc89K9AfiTTU7JKr7SWQ7
IxRf8TAW54r41Z+HY9E1HO9IssUMVEs5v+sxA1vkFysyRBZKJ0XZvbOKzK/Q
PehIL/BEvKhNxxCpnUEZ/oaO7dui4LUai19mrPHfC7Ewv5gWSJHOeajAa21u
psNA9tMWGOcXvKiTQVrEZVFP5jz1pPbTqj/P20Sma3+6wNaQMz1fPiPxLqXn
ctwC3DgyGTfTr/EetdKkh+8AX+1YmjHVGxovQouTdbe3Umr5UXLNJP1L9Fv8
w9Vgq8U3kdk5HnlYQXeDzzm00R+2yU9HHiQgZGj5jDuwaa2M9yM1fGU11nQ0
I1tC1vwbuUra2rmXzgdXwBnE9riBiJkUfLm5yj+x33s3sxlQHm0cvuCR1CU4
TYjmcTLYM8Pgodtkq8U3/tFYigw8YDUTQMbOnK1CBoJMZD8cFge/WL9sedPG
cpeK9dQlMijDfylhVhKBhtIeVl6EFOItDts2C+bLJluKNGepK4LvgVX7t7Sd
B8Jd81HqvtEXJgLzSDhhxBN0odrqcPeHawM7ciy3umVyiMtkjAnB48TkeyIZ
4uXzasnkwRQkEPDkWWRL9rtsu7sHnd5mmDtEyb6pWC8uSD150DcC5Um/5RzH
RnG2ZgnS4Nmx7WdD8D+jsF0DsGc1yOF9DIip6H2UL9gWVIv7OowUi1LSgbNj
Pg01soJ5Kgbg3MGorabs2v5NRLt/DHlYoAlOZXs+OqEi9XJVwggSGMBJ9zIx
VKjtsto2/ztxXdqSkrYrnF5HE6ezHGh2FUsXHDLtuAmU9jikV/pcDt9h/VAR
zkyAoKpWhFXCnQipZKMTdnJf3qKEhC6r9JkyRCRZgF+SznFgCtKfbYh322dj
vB1HIeFMo0r/funo4SspsipYbxCaTwbLSNFSzscQsJICvcm2fK5ufh1d4Dbn
zSpTRW1dZi2IcaReSuhNgwhFixmpIgpBNEQhtw8GJ1DCKACtSDa5wnfhIkyK
w0yoQxLO71CM7qt/eaHpD16cINSwaIHW2vNLcnAz3rsJiG/60Tlfs/w001Tp
6BidHU9nFGVbayUYniTloiQgcEjg/UzueXHqWpnaMzf8aD4hxABaIBsfOL0z
KPdQlDSvnPAPDXdH4kLUmTqgmU+nzy8DskyDZelMdTYeJIdHojGE5JFKtLPf
c/nX7z4GFA6wB1ywrb1N3uEAaV3X7xaz3zQnTWAaBJ0elDfGZwDrmQTFUtwP
1nvt8mlrUSOh+0uj+hkuzmhMaA3bfjLAEqFyG1fJWOD8NXAjQBNz/H47uanj
oTDNr7XKl+WHYFzPZPu6wQ38r3qB9l1k65P+GjPk1T0CvNs7JsDChBoyIM2N
67F5oiQomlkROqXmroNqtnC5gSckz2FifGGyBpHYTBVz1kznwPBQsaPhx4I7
lLe7avzVnTbS5TsBmnYAdF/MpByzcr9PbyDawHR64RS/I/sLEJToHdQb5Aq2
bnac16Trn3VYK/J836QXWqVk0OU2yiHbIALt2wirFQ6kg07Bp6REVQfh6J6h
oXN7MIlQIM4SZBM+D4HtEKctRmfe3E1j3/u8oC9Qay8mIdqJTsMP92RlZHZE
G18tK1e+rthAkydorKc5711Eo+2Vl76hoyufZFJaB1UBOwjcY97sp8B8NHge
AiC9T7wYSTQ0lRhi8cz1s1zzvA2nk+TtdZkkiiiVOFmL0q/6aBPGNbuRRObb
Ii8BwgoOU1KRwv9T0DNCEpcg6nnKmm5O2Um5FMTlpLh3Z3r0GQmHLGT7vtFx
lyzS/dd+N9PupiXa3OcZP0Mf9a/itlPNfMPQaRfgVy5UlsQ5/ba7OgRwRKYy
SaoQKKNacotOGV2VIzR0rndrCfR4CTUbQs8Omn/TVXXd2qd3Yy+63OtUjiPR
t6GSN74ORvqUPe2znwUfDs30OjFR6vlQA++RIbFrjF49gsBrpXmvrJddliXl
Sx1+KPx1w4LrhJR84WdRR42jqxwMrOneCi/kwqXMgZ65S50ppCqdLIAIbm7S
Y4UQIYjwkTxIiH08tG1EKcYOUz/dID6jqNtb/vfqeZAfc8jeuFyV+w5OJgF4
ljqbEaEt6hLrc5OdUEDQ2IeKGvsnKcNQ5Qr0XuLMMq6HvDB3ZyMCl0jr13Rr
zSmyufPBML490vFCwsN3rBmDD5r9CDQP5Y9vQHW0jkixgTpTWhqedrLucuxr
edDt8SWrLNzoHwn3OeN2/NIP6eXDGuHJ1B7EXcZAfgRzMD2W9BQ/zKAtMrfe
WBUC1EYCb4GRKQGlEIfmHMSxke6dClVqwbSrrTXvbxjwLvrFu+NPPmUYx2Hu
YgRLSGK3Qwge0X9nn7DPq7Z5BYECN6cSKRFH9D3FSEjlhV82t8wzkv0I858A
7yEKauhXMD80QMlsrGMPCgu4Xo5/QsZiPSolGZBvUZFe3Zezk9ZSr1Ea9RgG
kJDuiJefzCCv6p94VFEk+uNak+exRMCLFz823E7/RxsmqEJMeBp4hANqQgYO
d6WxtI1s303HDr6OL5OJCFwe96rcPfOiqsRvGKsxVgq6V1KZDFUGhWMrih+E
fhsNF/FnlC+/xmNLekVnzPfohgW+9KHEHFPMAsBtxvpepla0B44aHIlCDt5b
XQ/eqGulcOD5oAd/oVZSgZ24I2VO0FOe44YOVCGfWYqYJOrqCchIW+V/jE7m
TBHTt5ayuOU3/7VITUQ+1tEd/EnzJy/dCsK1RjiDuDKN6ERcz2UF1ShnKJ+8
jcFXk7SJQohk+QXcVtloRXrlrTSH4ofkVory4A7IIP2wt+fX7wdymXtAIF4x
EFPS9xRync6SMVq53jq4L9xsX3nGMMPVFiraPYEQXrafxiNZTu1cgVUfWImj
x/v0UMqYBi5gIm4EIEqmrx/ErWRfaS/+4nxuHueLRBYDRJBKuU29JNrhFlY9
L/jumgy2PC8gOzRZ2gc6XQQWHmfQhd9pSNxmH5EGcOYZiR/2A4vM44+TRyOr
tknJEI6bRyCzS9tJzFMbAJuOTwIP2IAJOwTFu9GqczFUO+JDyKphcYw75si3
md6wFksFPPmnQ/lYDFxxklqt4PKDIcJlhsYWhh6GxYttAKWFlyRK/zQGkg/3
jFXGyngcKJ4dd/2a55McfR4PeTwqXLZySW7JH4A3KVtVNnl5G3kZEzABfLMJ
T//vJmO76yb5C7Ydy9xVHbALS6veBZERLdrnQA2FGnwDIE6ROHndu+GzinuG
0z1P61TrwIrJ3xszpy3JXnEpMwfCpgl6TE0fW+YzGp/w5lmithLN2Gjjugb5
US4SUz1O8BAgkpAgL5GiHEfw4OyGb1R9HL/vrnBtzAvUeOCewiGtKwleymAR
cWqq6I9bJIumTFv9nnvmsPtLxEzBImkj/uYAcAjEWSmZNaCUbqnxkzVZAwu1
EV1KtBrJ1ezBtn+p61fMerk/mmXFqEw+P3M//4IIDKVXkWcHVHxC74YkaYNz
lcKf4/ViE7wBUZ0NTCJqK2WoVAd0q5CTqGSRsdk5QvqrggYrmyfYdPUr+ulH
SWzMaYusbvlcg33+ROPhPTmzTjd6mhQfPZmnv16mB2p6FtMZez3eVASPVez+
/uZM1D7KE5zAu2Bc3GiPwnS+nARoQtRo64HWVAjSY1V0IGvDb4MdJ/f7zD0D
FqMy4kzrskAo4iXJ49phJV5FT04rPs99q1ulQ3Rs5fykcjQWqkn/58JaxwHZ
yBlFNa8XYiTHgs1tQfaZYbLcGTVKDBk1FTFEEsSvcnKGaJLeUoN6TQpg99Kb
lIgdFaSiKWDu1Eix1KdIuo7CXLfixpF5iEap3d61K4l3PBKkR4EIspd5L8cH
2IfeqpegG37BOW8oHN3VwiqSd8pLA9dG5zeYvsjX5lGby1ssLGkYHA4YN5Bc
C9auMrzhQFd1W1xAAgY0qONMp5PsxuxU0InoBYqX5w4Gnrtib2ybPPfDe1Ii
kAVn7LMRuw0Ke5IcPYUEwRMhW1TE6UAMHOyIcnKFlSlvAqqHcFI9GCb3HfFz
xkbe7nfcZLH1NHfe04DHhdT2/+SQUk0j2cUAHLes/I7hf7Ixs7RzOc7eaI85
LLpKZrhtAugLfJg8scCZAbR00M5+6q+4uT7ss5iNJ52h0wkTbakD6XjFl0Mz
zbBJKoa0gWy6LAZYpVJgzVu7cEBdMkPXk6sYrE1sD3ssR+FgecmS45nSZeTU
QHP9f2WoNHqSRpnUiUzdORlpyYOLVLNXIMylW+3uUQEIIQTseAnJUIjlNxAJ
FunSs0UgZFnqAqlKbJWvCrTCMkiFW5DqQPWHKc/W9gbJ6R95llcPdYW/qmja
hX+VASFqxgf/1exeuCbdl6OWKZ+LMmP0xjTzLkR+LwtRAX3xoSnmYCNM5qcB
CW6V4RyqeQCo6QTAEAeUMgEcPvU2ZRNqwXKs+K2hMyBqBxGCORkTw3Q7vY2R
UN1Ceb7AGDBYjqztIaAJkwiFx9qhnTowQgDBMUjlPk8WA7qgHL07LESdm0xU
PjX/gs+NVv3nCVgzzn/ilO7/MntLY5676ekNNCsdausIl77SB47GJ/3HZf77
0nmwhpUcgi0OJQuhJXIzfTzabZhKA2L2pWAHamx9mWF+lbDdvApVK9HI5kag
Eru8haePrH+/+SlbF9xM606n6avacKM69H6eRMwacxodJ4PFCBPPcOTXt5tf
acLB1e0lUQjQ5q3WuKv++HSLIab17jKsYNNIubiymSXZtgwYm1eS8+Isw2kM
VmrVXUzMX2fvpCw5IP+PKwhz2lmNRYfLZ9smwrJiZE4Je0XQwHHg0Mp2pxGJ
U8/odNJLAc2q3OL6HmibB9zJVFlkf60xjwMzfWDoomMbZ5FuPY7S7uUHvSYc
RlNIn1RkKA+EGkCqH9MyLWZAYWxxb9mZkuG++kmKbGicSY8kyresEv0BLgkz
luSKt4myIfpHJtihxBTjiWZi3saN7jPb5A6MSjTmnlAfcCwsvGstDDIXY8+o
NhCycFe9yjSfUAtaAttZu2bYsvePFVk87rO4zeSQ8X/UoPt+/5cLvo+QPe53
gK6RDXZFi3xik1G38rJqx+Aoo+x+9fDIfR5IlXp7H5UgucxzwzrzjjqpNxG7
x2aS1vCqj6wwSgyngfzA4XrSU8KMiTeEenLpYBl8t0Mi1tvp0ZMy6XWUPtGb
ZxMiCC+2caMvVdJgDXRAYf0bY+a+ii0zcl+K8coQxQihkBDiMatGK45EUQv/
S62dKkXlt4wb6ezOeiLpPYxN5Baj8swqfWVKS7PU9IGsYZnQ1bQvEJQOOkUL
RP6z/SAC0/RtyWEg+pHMEpFg4xzQ1T/7ZPmjsuW5Ok1LpZy2pDNSCCIg2zp0
syULRoqGJu/PxZ+EsDkfzeVZXmpda38nnCyC5oq6pkL3QvLtgpYU7XmCWZGi
oWn2Pbz7h1uFK7+LYvyUw0Kl3SimqFyMx3Be2EWuNPbvvxZTw2vjeYGFfXV0
Hp0mzXqrDHR+Oaj7XZ6JLUFbkiakIMsSE+/fIVpbHOzYOxt9gS0cUndLhyfw
W3+guTqKVRyvmHHBvb46lMLFHwRhvxlmvtneZgbWHnMJhCmhMsVVcsqQ/WCd
0L07HwKkxigEB354IelBCA4FNPQNe5f0mtNngbxDdwiUZqbRs1QXFwMxwrxj
LtQoqAbTVxjBt7SBL1mxo8JcH8UuHpRpb+vSMiP+ahneUB8bXrEVIGf+EfU+
v3NPRJLuHXF5mt/nYZqfBQKUhmNbM8+Ntn1UM6Z0BVrP/PRFr/qS8O7AOtP0
gnoTsTB3gRtUTnRv6FbfMZn9hhnilKOMtoUdS8Uo0I1Ng/4ZOWItaMqoBABS
SQfsTQ9dX9K1nxKSETfjlGBy3n+26rqyJ8y+ZmdTnhsQ0eQKO6sQiOh/Q2sR
jpV2s9i0Mfn0/GbOLCK4xjUemMNgVOx+0LmmMf2kxC9hgDybYQIMnN196vfG
FWyT/36giLLFMaoRm3hajPJRJtbe2EGh45hyPcTpDnEACTAiXch4anmXUl+E
9kxExpwpTrpzkMeDYhftTy94mNBHJekBTB6dBoO/mGYH+T/xWYfG2aArCEap
2K2hS5pBJRLXDqXUKMSTUrW/BjML6ufndJaP7LZpZebZA4wZdpvztFPk2RrS
rTBWh7i4/st6HXkFh8HVqnJFJRbaAMeFlvECVhHDbI/5wBQe0oDFbYLzsEtx
vBjxExRw7wJalSyI25YKDvJI5pTwzJpwcYswYptAu0GY4hSySVYrYQLRp0o/
v42XHdyuszcSAtMQf/OJpwdcJdzNVOx8ELI+BUTOYMo/9oEqbvC6To1lEp8b
LEFjkcr4wl08Ol1sz3jBuwI7cztCpc/txUXWXleKBdSIraqqWfp8SELe1ph9
6YpJFR1xBqM9NHJWFrrh4XDMdB9v4kNGDEtAcLQZwJQsTCWBDB8cLCxPdnDD
a0sRHOsiVyJxYClRMGINdGmobqMGv44Bf18zE6NWre9eDc7I6OZw7LkaXM8L
vLLMOC0Mx5+NoYg2ptNZKB/d/W0yRniyU4lpoGjK2oIl0ROxLrCREHHytQCy
28cC/Hi2bBjmiE5HmCO/d6N4Ibg2SRT37oEeNgl2SZYRKp7MGY/+GNrQjWk+
qyYe9E3+vt3J22wKbOH8Ephl0ItUFa97YmMmLi6jU5h/j/Dm4rxB5nDmrWDE
6lqIbE2Q/7rCaGlhZkW/7pd/Cllw4BUqXn8wcDXbL9incXKlrnZBepb3Armo
lPVqdUxHvcVbHRKFPMmtdJ1dvvDVRk8Y6a/5+0LLyujFy1xXV+ckEvDM9iYZ
rmwkq9iE5apgqeSXQTKol6HCwFE6s0D0MS33fCQmH2Grq0y4VVFF8eo/hDu7
A8TrFTsD47z8gbtuLVNH85Dz+wbidMdH6gEN0oRoyxbPfDSeiXpbCBB3Y/5C
lnIepgXjPyUfi//YLiDuQdZ8V3Dx78S2MamW7f7TGRgQcU75MSAaWoOH1Gch
fNjhuDZAk4k6XWl3DYkyOLee6ApQ+29dNwxOvbrYZ4fjrNwU9PMMCy5gCIJm
TBUkPu9Pp/QZgDHkQFMa74h2NXXeQFkyceI4HvnU20eWKVOB7mb4mLZTzNHx
rcytHkRluk3fGHJnS6lB5qCM7N4Isx3+bJ3+3g9meBDYJE28EtorhMeXqGRt
XA3wtOjTT0ZzSTNObhlxBQT534/sg0Mkg+cadZ57BTfQjVP1f91WPuVzP/FG
pRe8FSDcASrSlRI0GELKxDYbmkJtZpi9yOo08ib8B7rOgfePpyjIjeyao/AY
/a/qAjqnISx/edUCl/EO1tPQWlqKNlnrRAa2uLM5PfRiTcdpyXmmDJuHgIYc
iNn3qmuvsdFk3RXd/7ZCyMK3KTSm+RgZEncsHgZqTShDVJmOGZXjwiPxHmcI
NZ6cqF6p91w8c/NmsjvaVetNvF6j13TSpVGAEBLworxfE4jVGMfjJJ3AXma8
zRHdZCwMwVhr+4CvSMk5sdz0DtequuhmwbCBLbfhuyxD2FQxedr0XRTCwEUV
eMComP/PGMv1sczQEjaGJks8yoVRgjclpMqyTqe4hlb8Aa5Fi6P6XU/n43z3
kSV83Y2io73W/xDvRptv0cR07rCTq5EtcGZDUFYh3xJ1lQru3gq1uOJ05cZ6
uVgwPkgxUHI6r/HSbgHOZgEwImfi3Rptd1TNt6bC6cUWuSINUiyHlBLR5I4d
vRV5t7tXnhR+dY1IkCRDSlXu0U5wj+rbO9lcynksKPRm7s1Ejvah3pmMIdKm
HkNu8L41849i28+LTdOtPASZrIHuKAD8P9i2AQ7bYa1+cmcMiLQSiDpuyyxR
FbBTwm4gyNYbBoMELGwk/NGT73u6DkZpxAlgfkROswp92fss+v/ts8+jmiKl
59wfTIhEsS4LC/LTfL4YmxE/PMnCW629g7GmWWYrbTQPH/jZciMvwrso7XrX
hn0dqqqA8+J7GU2adFeCwMJFH+RuwqNJDjThB8U9gU08WyGt4pQtID8Optvb
7Afdkt+GHnzB25e0Gt6LcbPKkH9qag884Pe5ClqkoV9tzBACnLsz0BtyslWl
dGNKu7wYlb9sNMa5SG7m3QwT5AHadF93oV2gn+GEWd4d/uwS8MA0F4UXpIyt
LyAhkDYIh/PjjItEuMP8ss0QPCeyaUXsx6fgZnck3qDCH7nQk1XNIzB6UKiY
DIdKGi7IRDiVGW5ZiCmaMDs0tD430T661va27cRQQUPMVt5ZtozfZMio/T//
7N5KnG5rlH8JjxfnTl4Zgk7eC5rs7+PzCCbQnHEDjFwxPgifhwyiA6qoM3yc
w6VxHzyPTuLcRYtgTk/5fgqZrZ2ru/pllAmU9M3498GKuznRjStrlXylnUPu
KI1F9bybPRgUJAIyccAUnj1YvKquKNxRnMqnXsFV3g8n+KI0kofmcSfcQAwQ
chrt54aoXY/Mr1oUWiL2ZMYyUN5VU+VqyqiP59or/oLBaSfVFpiKdvCm6pyB
OmphNxOQuiEIEBe2JotTFpXdkar2jDAuqT+Xsh3HrkxR/gRUJnYM3GAkL4bz
TSVueC/LJjTxd18IytP6LX2+pk0VgquSOLKXg17tHqEj3gU9EXa7nPMUD+iq
EG/kSR0FTMG06LXiCW+UN3bZ0SpHic2WmU7jCdtBrFFf+qHbpJfWtlqDlWyt
VqB4uQrgsUZ8VCa8i67kDzBGuMuIoSCPwklE4+D6CCgxedqw+UA/fUruZcoR
KohSoRKF1r4G2TDy2EMK5dGoKDVWA1VoGtDoiDFyMNvPBIB4chFmbCVQ32fD
1t83BizEGhHvwyCjrX85VZwrizPnlxO9Q5/et8J4LO+TkldxJgcUVtaK6pjn
fukcv6oabL/PtiVUOOAxPQdxpvFwQfkRO8cqDJoHfjmXvMaZbdyJK5G0J7p8
AC984BnOWdssGprMXB6uTGWvedUN0mRyLcYTd/+v1VHGxGA/wwBH5HSGFBPF
9nYIkAq9zHrx6TszDFU/PaLbGl/UQQK1NZ1VocOcj4HXT59NY19DyNcYOhXJ
yJhnqngaIDGeisKpx/lbCtJ3Xqm9gpG7FLfuS3bMxfexiUl/lS1aGjK6uWwQ
8DYsQ0VxHKYiZOI1De8sVwvEzGU/AO/rrgUbSp3kzwZTyipSy0DMdtjq/n1j
keiJiPBCEpAHOmz2wOsWV3uqBDf7DGimo8gHrAJxjTCoQRxDi/ixdaQwASD+
USwVKllGMIX/+phh/83ghkwlnly+6VyErAsaJZkKG10UrkVQhYr7QloZu+Fc
6NlNZU9x/SldSCZ++HuqNKAj7wNSyFGKrV0/N7IePIXwAQ5fjX0hsfGaT57Q
W2LM7ztrKZGV+2sKrSxRTZ5HDK2SZR1E0tmkkuUElFlKgRLCI8492q+1A7Z5
axWHa8mvKHEv7TviFJYAeXHRNiHcBiLsG3McS/91RVKVKTrsv1+wS0e8USuN
LPbwrONKeQ2ypdJH9tWYCng8KR2KYkh/eCP/ZVS1Z7o+MwXIXOCi7Myox/YR
fW+14mxEwFWckBfYUtSP/bVZKOQtQ1qdpDazS83CK9zwJXeIfIKssEzx+/WA
Z+hN6nAwL6OmZmecym0VU4CwNo7Qj8MNWiUaKHxVfalbw28n1ChEze+PTOOk
8BsB72CHhOO5Grgd1/YE7+1RPj7XQYivsthbD88oEmoqUyGHWDnU3NXauFMT
LZC9z/UcA/7JEpgoSfMt7829WGxxRHS8NzKlKiYKRKGN6A1V76l+d+/1uODS
cJsFc6RfRxfkmbq5oHYZANZk4ojpnRQaURTIteAvFGyPNOUaqh/O5QZuk0dV
t9c+PxNA9cLznGxxgUR72KXNdbpwx1SYFiW69T0ATIt0FEB7LDWrI5IK14UO
dPAnoNKaby5nme0bjqS/EQHL0rP1WLyRjrhr7C8DO7KC45a1st9/c+Gx/18A
VCazRcPZKqYslZAXNG2DRCjRYnG/3gpitj1PnL1SI1Akr3GtOb9fzmdvII86
UPVAsX4z4UKDnCBcGC+/9Yj7vKlJ8oTRdCEqXfGFUFghoBH6vOxTiEVyhQYP
QdxYEUBhDh2Vj2rYM2NXi5vFycDd/YyAS/NEn5SL3e8clizIif2aLOhtdl7h
cfSMOCL3rg4LVXJ3Q5atzgtE+RbcXIidiLeT2O5fZSiUdijtWQF4fgbP/6Wm
kX8oBx8n94qIb978LC7mUpeCOX5xj4VY+XRJ2k8scPO4B/j+QPOfpI1Xg7KC
ravCIqEzMnLBMftz86CJn+QcPxAzN8m49kXA7o2/kYi8KHCCTRo71AB2QotR
400W3WIcAvUAotskknuTLZ23c7cUk4dt0J/zyEXTeEbS0K5yQgM5CJfuZ+v+
1rlr8elsFV19vKHw2ATS3Bw5kX75wZCt5aI203GKax58LFQckaLyQpyORQVg
Vu4ZgpLrOU7DDLpM/+TxCBWuMGxKYANo2QTx921VTiBYqRPN9Gjs2DGDDE23
2fvlSEQ1G27xW1og7DNdMhNUyQnyy4EjBedmy/tMkFs8JVpC3nkkD5Vha/8i
3pxdFlmTBuQLv0gj7SZJLJDV5h/XncDmBopGkSMuv6Xv+WvFEsOeIgITOy+V
dMWMmgXfOLzlX6+h1PhlyyZvISrQlMuTxO8dFfh9r2xMpIuPJz/As3k5aGGv
NpjbDUhTxRXep1Fgrjt3VMMg0iigmqziRVPmzI8MJbajRVFejqcn6lYah7P2
8nB3XNIpcTxtIDDaVWbrnYbdZ9hI9lsFH4Ido2mTvb5u/wZaiso6Mlmigjpm
qFjWSz5NqkPGOwAn95y0+ZnzMHgiH7U6pxKs2/V4Eov695g9z8gwuNdAt8ft
AwIy7C+HWuf3Vid86BfSd8Vm+TYemE0f5qe/6LAP+g5QAM8NvSUE16SFN5w2
GJuohrMOqKKDtJ0CQZRSl5LdtSXx7DQv7JtQEXgBG7DS5mkBKerNtyO+SA4K
oitIiKGTWeuY/EwjPmIYsC1I6ZMXgl1P4BELOTKd/DeeRQbWi4+Dg4uL+qcJ
986W3q2GhubtKZuQeFw1/dy2aspA5xoUmWarbqJmpFDSehjmIOIlpEIQHK+E
kAPjdYBh2AbnBPeXI7Ms0Bk0CfXHzhtgCtRt8AVpSSFG4ykGRPPubpdFqrq4
xw/mpi0UhqZYyOmAzWnUokhMngk2WDd6cE9R5Y1mPBTTPCpjBrMKrRXRjfSG
7GgFxOFdAe2zDsW7I92VuVO0RkWNpHA9bR2zKeGGgxm7BMRIEyXct4Iu+qr+
e6CRn3zhKON0S3XBIj/egoBeSw7xtCjdFFtsubQQeQoDV+bUpAdA2avxgnle
w/WeoKN6lntnAOIUgH6ar7Duzx6tVvmd1W/YFhwPTt72CxosLvq5L+RqOdmF
rUna3X6FC9tcMWgLM9qyIshC62TRij2jD15nKPkfTVpsMwQ7keUFl4xPWj4c
koQSDVXQlnmrPvQUL16+oGbnw6AmxLNL1Ks9ibCi2boDoWOZfd3WW5ATSePr
EUf93Ft9k6fItFUo76KQh7l0FLvBBfP+vkoagJRQbaOh/TPIhHz9QHIvuNNC
QXrRsFl41uIh6o6+U+KjduLttcmEqID/3jiC4dhrl3Xt4ugSEpZa7tRJxsdK
y4Bd6+ZlWoLEiCIZrwHdsBq+3O593fdCX+mzs7yR3++4Vv8rQ65Ar2KNPHds
RIaMOeerhdQhVyUZmXYZEXWG0vFDrkvpzDhXxhdWz5wvAxoZBEigCc4e86bh
qSNH3NrvKT0duNaUuPgd6hB0Z8+WJdz5p/4XyZpf6m7bQttCl+JiM3KcEWgl
zKXVfwdqm+HKfMtwT+TO0co5GlNfLHeElmfMdPvQCuYCSdUGJBtqj9Rx8Isl
AXHqLNylBUAlQV0tmyEtfP/H/2nVS/qFywuK1iAniC0NB9NabdogSrzGYdbb
Uo/NkQoXsTd1ycVOGu2iyVqGbUXQkQlVtOz7LqAcEMvNhgQD/jZYMh3Ov0qY
LVB7TNo4i7sxyxQ9J2mgjwQG87Pv2Q/c8CacnagOS9AcvbmC/6QJWRPXp2Fp
vlUUWDbzKfHtLL6F6bvhwzEKFUP2+UfuR9pz6eYuLokDSkEpbT9nuKUC8FRH
av1kq98w/fCJME3me2CD66PRm6WPAp2DyHtS4ZcjlGVtSRzNmUAG2e4Xr6uT
qNCUYajIAuRvrzzjMYHaqzPcfKfQUkyIqzu6DVhxVnEcGLKgttj1tQy48Urz
8sBnsMQ971phuK7tJN/QnNq+D9fs9yvBIjkziw3EmhaHjThIq+mX6EPCzqms
gaJ39lsxZHqr6uEOqZx5IsyBvLyi0X5gghv0o8DdUjPfvkiXBnP8ifFhknJh
AKqVxLwu0jrO1CVTWcDEL+nsOPZg10z2kgESklrDxsG9SCr0421t4xefmzVn
I8kfpNoNGr2wlLcKx2UIbHTPKdI0s4MDMoJMAqI2D8o9D1SYzdDsuKiW8Ylz
tatY+zrrfXSItk3hwOQt3M+cakioWVoOWTa3pE495EykeMM8xlJq9qViB5a6
kBHqClOOIc/nsrsP08brb+iE2lisJRMHVrVxitWmSTZ90bX2wQZ0z1f6Ky6i
iVNj88KMALI6j+j7OUkKuC4k59od7cTCYSXxVxWL7xONGX2uF91baz1haRLo
ju+ngp+kL2eCoLsgwj4M+wCU7ZwMOUw3WKzVFgbMnLDe6lMIS9q3GySKcFc3
ane2bvF+WYn4vHaqES9PY4IaDuD9TdKYWlJwV04GrM30aQ1RuZ+axeq8PtoI
1JLQTeI7LOhT+IVqwANZSxxa2KHTq7sYfBo8BGyIV5coP/X2LrFb4RN734dw
zZ/KGjX2iRlP5jnK/ejTJBYSd2HBmqzvNl2c6dVoB6mSP92OZhChAHMNPX5q
b+LtwtnWXv3hdNkEQvKBbGjC5yEBcVexDZE61Cxh+p6jz/Qzs7cDsQW61jCo
KmGCSKfSMMinPgN6Foees80w11PK8zSSemsOyBAIJF+gVijizQs6VCyHKcVW
uo+6pg6x7pXlOXgbH/+5L1d92FiesVBJ2/mua6gso40/m88V5CCw5hjM+1i3
MVI1/KYfdNIZjbpfPxQtTH0ail79rRZUazjkJYE2gRsn5rWGP1Y8wH0K1eGQ
5EHnFulishPeFNPbkXJAQsX5iGPRf/qzLxOYs4TXc7GoRJPsCPKBA1gbMot6
WSHduDbVCOdovi5zXlrNKbtU7tG5Qkzgzij7j2Ovq1TPxwUk8mT8BUYBqC6u
URJz34W2J7zYqg0GXb1rjwpO+j4Cy+g28KSggt9FzfB9dOH3bFfCWdmJHb5+
lMaRLMCtl0ugzX+iL3oU7aGAixW6sMMCZfldzGVpUP5No2RyRqXktREmcOij
RXy625EIbxvsIHzEA+P13thmmTwqCOf1mbHKApejODUfTc2Dnyf4aphLtWku
cLMOjAvk9xOPAJ4BzjG9A8Vt16ZW6/yZ4Uwo+XerS90FLzqzDYzAe5BtokZR
f4hHD6q5wrUwPdeejv9cFOE585KY/9QYBBZSMEGZ1V8s1l8ZjWvm2qdiyhAg
h/xzVbTW+GqCSsSj4LEKCX055ks/d9LkHBN5bN90DgEqGwdM1M1HPzwQKVBd
9ycpXMwWzAtB1KtshxUZu+tK+Tkgj1TArEIcCDBvPMNDxf/SV1PLf4k5y0Cf
sa74xkcdf+xgiHgN1rKzGa8xAefhS4Max2QWfc5wV5SJWTCtAho2w0SGYVIC
wsAMzpE8eSuUjDQVt+V1MeNeYya1WP6fATewwfQGBMHeHT6tVc9c5RPluvDK
U9LbgHs8ehK79IeE6eIkwwsqXgRYjHj6tmxLEDL7Kc5bMv0y+1Z6jwDFOOZ9
55An0qEDODhcOgsB0rGgyGbyJNZUzqY8t2dR64xqU/XFFSHxjDOjM0oFW062
DLb0ddscPu2m0/KUXn/++NPrLjs4xB2u4Xydfj1ZlZbz12dav+qwJLI6IXNY
OBs5BnBQ+rURjPNuq6wiLO/EAJinI+6zS9jm6R3gJUeNMAc8inE+TLfAEG52
Om//rFkH9IYMSgJuuHFHr0GirPbaBVdJsglbXgSj3S59HJAOkRVNFRjGyKdp
rJaDmcVlv5XrREJQIWpLyKn7SlG1hIuoqpGJyIwab7TyMVx2Rk5BJ0xB4jPO
iJkbH7vz8jqV6Tq8AffsyRX2DWt6vXeOKUWaHCrSfjgY9s/9bbubyoOPhVDX
7AqWQbmcsuApnvKkxBXPQokiufe4R+Expb5qjwy5Vr2ZG41aAdJPS6ZleqRN
Vk/F34yhNEVAE6FsQiyaU6YWYKNoweFWoW81EaMm0d+o0H7vMXEeIvBkqZoT
69Z/0LK3q2dZPhpWqf4EWz6X2t0v5uaypYAZl2lNxcUAGBw6MeW1AQB8pK4q
SKG4E5CIHZADNyOLCx92724tH8vMt9gA4Ns0D+9+IXoMqKIC89aVLoK1DQ94
GnhNXqNcpaG4OPRPC+k4JXPqxKPKscIzFUCic9K4Beft1xuXDf5vDIkK6sDR
Zw/8nCxm/vXXNVt4L1mxxxePQGNoTBin150xEWmwdDeTWM9ixGx9mJ7lBSWT
DUand7j4fqdGWvs+p547SHNrPKy+WBWmnOonYBaBTzLv8s2VVhaKHQNUFIHi
wxfaWa97s/0wBMfksN7qF2mGdaX2WD7Ztv7E2+6nygr+maWEDUrkMYRnLiUp
wNMSWBMYgBtrcuFUopNMg8bK4bLCwYUbG93YFFa5xDs74Id5DJDULq6jou7a
HnMIYzeyEDcQkHI4Zq/MhO1k+X7smFnytrASfC9OV4ycWOqf1cjQEqHVwjog
f9sjPcj4NKUl+jp9M54vohVTX4LNbI5pyrPZM1tCratAz1XyXY1P7hK1XEQX
lgBINH1K9PFd8hj7jX4a15IlDel69gB99ge06Kn5xTUv1Ho0Tjlf021MtsAa
GnNAiTq/rMPK+aHxEk9cXzdC5zZA3JlV9PmjNZZkrHDZXhPTCvh2+Wg3Nx7+
Xszok9G5tsirWETUXcBVHunS0/U9RcFL/wFLOdFKoO3tuAVZDzdVTr/amTZg
v1cC7tGzT0jiuyVxe8x9mcnfhFuN6aQ3NXSqMkD1N1Xb4HGU9dDkj9TDRV5H
aW15nhXv6Okx1xLWNum881nE5kKj2AuVhV8hiL+vZR1mMYlMwtfgGVFfBAMO
cbdy0oeyn0SuJmYFEEi7ODqcotn31ACD+yeS7QefN50rM2iq9MAiZ39r7q6o
Wu6KDXH1LjQpnuUbmbngFGl/qLBxxzG8Fkyw4R2D+hJIGEH+zcufZqVZOaOa
E1ascLAf5droxdjEAyaPtKBRofRhNV8ucUG6u7u7b/HiH8sLKKYHgo9SQLcT
ko15Y6sI5MEGo8w6jNVRZXeEEEvaxJdR+3F+nfmEbaqPpMcryQtYl8nWrAY9
9tB304+nfg4C+jY5Mltq+RBPPsg9IA3Q3nnd5/rQTjPxegoLhTDZPDQP6MHy
oJyAtvuKp+2U0ThYehNSw+gv3gebWs1GFFmRqXh+zYpeMwAXzvYI+nEeSpUP
oM8wFNEcRjrKOmfTUkjOJoF0Q0nLoXjFzY9QviW3/9QHqqUuIndgIS07PuDl
F5ogKkmfVtuIbdxAyhBoMTKXTZctN4WIhQkG9SkBvo55pe9Md17g9cD342ad
B0oqLFzPzTjkBzcI0zSEa9mXsG/tukYjUMNiqRemkchySdLmjPjPUEybQonv
t8FIXCS3OyJC8I5Muq5xe+rLoAiU2S6kHibddC72B4uzOZHKky4g+oinE1I4
JfjequQNHUql2Y60X1ltd32sUkMBvGv7NVDpRICmn+1aUkY02OX7z+gDxxio
B0S+dFhMqLIlKgGE3/qSkw50C6xxEY08gXnBjhq7hajYnPaFJ5YTy4/VrNti
d7Kr99FcNCgedx1Bunrfii9XA2C/arqxIGjxfGtX68RWTbWhLabUIngPyZ03
bwqpxrJEM2ZQDLvpDgZslEyuUiSBqh6p/LWfRIe4Mw7TAWtHPwSVF0Spmc35
AhU/hzb11JJhq6k4qOilJULd/EfofAHjZuXRzW/WOyrCxUZT539v8OYoo8Uv
YB+cAl1lQqT0ao6UMmoBOUVyySEC4kEllNjBu7W0V8pqQnB8jxrKaAbhMMXy
5FyWGyALTABqrTHgCoCxXOJR6XxVuD7rmXHZanMBQ9x4we8M6jMSZOA2CJNR
mcjESkSHJ9XZJP/XYxfcT/3fT47CLUxd1nnzHFbBfhQJiJIoDBKxduUv9ysr
hi8viP8ExIwQVLeOp0Yjnyh8zf1jbysIOsyhOptkACDylF9a8OKYTA3DopAY
/oE7VdC0gEzMJQOHX8J5tDg6gQbTGVF3soO22Xq81IRbOZhLsXo88UnwHKUx
wzUUGgDSQapINT+gpRwjApk0x1D2HSoVLS+fnEEyBjj8PJPv81c0GRzfzP5k
nolj+Si56R4ulMLFcO+k2KiQCyXYBRUG2i4bbXJasdhvMaLJ3a3Pptpr+gBt
Ot058NUvVCP0KLsQ2OAbeoNezrfamp2AIUYaFlsbBPtwfE82icQiBB+dVGeK
EM4iSrNwcOGHIYGMMVqlqD0FIHKbKzOX8V3iMyLXiS9CQe5oGQCuADn11SyM
s0j9G/99uolHC6FYwaFqCWXpuIjP688VF8UO74u1E4JhSXZsmRqNE7Bv4joq
Wo9WwpaSUTs1FfgBCnUM82okKkU6UO79eBFr9Y5FY0ZOdaL3PzR8KLHI8Fkt
SRsfd6CifaFnmugijEi5oOndpRsY6GcxiPS4XlQdUC9SY0qDMysU2nhB44/m
cspkLkwtPfMnPbQLMK4WjcNW1AE0i42I3LbP9OmECg4fTDrcWIaioA9A/oHY
TM+D0jaeC85jid9G+N3KpKdhYR8U7tDo3QcvXSGzMxTjsjYqkhB1OpT8hNXB
znc+8L+rx5w87ZkjhJWB/Gb7g1yGUoNlgjxPKcOgwiLjGqWJNlmMZoKoqF7+
06Fghe2YILFe247bobq4kyGioUlROgUnk3/Yufo+5H22oujGuJUg525kzkvw
CDF1En5ChyCP7ijT6IT2oyJrcx/li03BaO5br3cBVBWw1vhjpYbwErLDpkWC
0Cmgr26o0aqwqAUaAZHCt3s74585vVAhiQ9utkYaHGg2iMrYteILSVxNTEjC
4p9GIZVddsJdikdfve71iPpyTKXIewcKHK92pHdkuOoW3QWIKFYJ7gM2jSKC
Nw+nHGhoRaPYN7PMJHTwMsYKkqKxEgBmEKgiNp0lgmwz0QbxWGIDsbdIq/zU
D9aFewdNk+P8ljeQPpklkT3e3jikkesi+FYyKESVmRZ56VyOUIgneVS+mVnV
zdj8S741Dg7mh6PNolskF5iCWwACrGs7cqJzEQDvWmeFuiQ/dR1lWGgnt+qw
r34QpTwQfl5G8ZLW5lfxjzbg/UUY+hnT4sZUPIdtZcSeNiwpPx01MT6fjNc2
WkvdyYZqTTayDbEjBpbQCMdld11DyiPo6A4B6w+IRAowkjtxPkXM8Loh86Hs
yYPlcOnDGRVau2qT5emULiAeUYBK9trGaO8a4h0HRbsfuhyC7OjJ+XKU/x+J
yhb27KNkSvRJGEPn8gE/wH/hOqPBAsTGSH6BDoelH7xbpmcEJEOvNO1AKjUt
Rsa9/Ei2OHqZM7Lc9PUKswlCWVw0/sCx0EYDOojOlT7QOLkErV6SIxnZjAUI
Z6nFjdV3mvMlACtpNA7cok8Xye+98EKfRGj7U+4NzBvnImYVoc33k3ybEe6x
ubk10jVEagTSiB6tncSICVEzZ1JUkJ1n9xaiW+hL1R9Gdn/y9H7lFQu9eHMX
6I8RcbECyFSk3vFtri32RFRwSlO7E+62cexXuCmxJaR4AXT0NHSwXxvQ7b+r
W/znW5ZiZMRW9sANxH9irDpEf1/DM28+LPRUoc8ITnhjoIme/vxOwtCTa88i
zci6MX9AjPDIGUs1WsQVAzp0b3ZwARuanXI8R1jXmjhoqHkR4LVdt/pRFCwr
fMYUoFlmJMbJy6Q3cb2zn5smfb7pq82wVnJm7iwdNBeBvJwISk5RO9iWa5KX
OvHZo8v7EHypPDIa3zr6PWNMWyTAHzp/7siJRI5O85GZgwLaLK6USxzJc0y3
DfADogbTeKBN4b5g5d1YUU3oIjRNtAEhkgr3CUoTaCqGKdcOKuO1BQWofTzQ
2Uv7H1vaAlOyxR6+27HSn9CcGtGr1JoPSg4stG1O3f9KswjFScfE0w1IoxHw
aT5YIAa96No0B2UNmEpnsaKOrrTq6sbdCJ16uyfqMT+MhaZrR89qepWkF3tl
IgQvfMCqP11829jY7vmJYnVyymFlSmUftWbNirwmzR1v7lGyEsRlZZ3IGz0/
ytim+Uz5Qb8PMPnVz5oFIPg5/ExlnJvi7WkzTdGzwpgqn5GaS+WQIVOxJmWD
k7KbThzB/WHu94zJzHYy9Zdx0ZmIHR278O93lBLbLtDa5BAKIDKWwSq5VOgo
PXtJav4lKgU0U08IuTmN2448QzsW3Oap69JdaOb+gkyjrtCsFvWVeYxT6kmO
Qa7N0TM+2YL/9FpaHhmb5gtOARtNgnUGZdZS6jvPB9DBVTMoE3t+w90tYzub
UXu0SCDD/4pMJZ5eBvJQ+dZR/rUQJsHEW5WIprQ6CJOT2vCS6mYe10x7EnpH
FhFURCwSbhiyMbVsN4L1bACnalQx4DaKFAYmbPPjbxFmuaBzwd0dnQpLUw+o
/DgVc/3Alhzo2IAnAF89yRR/7qxYxFS2crCsuU0hy7dExtpsgAsTyL5SVM9j
aEjf3eabF84+rUezijYMf1cvpfQeMHMBzNeXnzVGLSKhd8XrRKBKJfHCHm9R
t7FBNfpXkt9TacLAQ9K5mEQnjx5Ta2O7voVqk7RTE1DS2wrmbiQOp/v3sAKh
KZDDCmHjgoWWZJufRS+uoKmUgWSUfwIlZVXKRaGXz6Qo0nofgc9M0TnI7993
JFvOvnws1sAc6OJKq2zHiX9C8kOductBg4ItXoKVlTgVsDcql/eyHt64h0ry
FyKnVvagpw60rczMaxI7vTVFU/VYQZVWTEAl4UxyyAPTsJ7byX8vjqFbsy9u
00IWZhA7thyy0uPhg+beejVxM1R2It/h9zTOTch8yHLLk2gKX5VNGRuhCQ9s
Z1gEYMnktcbLXPIdLPh+SDWGbPxxDJ44PAgWLm6eImp8P1pPmGKQE8mdUHp6
ljZ/X83ZiIaroP2XlgFT4qgRxY9PUtu/VXewu5vc4/KVXvTYE3+tAZAIgNOY
yvr9uPkPzRDvWm0WOZe52y+818RK6wuXAYLiiNZ2703VKRJSEzosC7YjC7e5
AYudoiBiQPmdxW3/Kh1Z+VPlPBcgGqXgylBKl7VtrbSlbhsppWSAoElQOtEv
P8LJMUSIAgVpQHidLWkwSfA8z1p5G99A/ABpt7H1ryhnj8w3RI0VBizEdz1R
tqx1xtNS5DOYTEH3tpRwlyPOrtxp+LPJ2l6UgKVB8zLIA0cDVRd0bv7TBtJh
CNYe8+YXOu+YkV7QRA5iixOUMAcpDmSfKN/RkhkRB48LibcrW0Pehl8Zbphm
EtNPLldnP1AdorGMDlbFyaZ1oM25aMjIS4VOIWV16nhNq14EUo2CZKxT1G3y
7PlU8a8lojU1Vd3qhShgZBXcXtnfphJSmsZaLVDTnLpVRYf00TL06jc+KRUW
EgcuDKz0RytVHmDXZrqttQikidY66vYWvuz73dN8/0IDO98tI+MxZCgDXDcO
XHX2lm3bG8XsP7DTaZhA6wrvwXA9Y+nmJPtJnv5kArJGGvCvRarTdlfdMR6X
qARB6s1hV0y7I9xj+v9lb/ynuFRtvixXsnlEsKLsXuBTPmf2jTTUWWJUi1rk
HSugXB2A2AVjEp82nPR25HXxTkhzWBLHa9TYuhu0Pya4TXesN0y67A5PD7jk
aCo6mPByrtqmDznxJVQDFULEdIcmWUFSjjZdgh6Vu3A2czjyioNGjf6NB5GU
IoRvtqEPDWRlH5qzB0qqpKqPk3ohEJ+EN9ijuOtBV/o5/3hOGuyLD7/rLDup
J6o5i5KrSv2COTJqzCMKQiS9dSmnPR9VaBs8s8pydi97Ay8NgO8fukrtI1a0
G/6xd5QjLEP7FNrFHfxR4rtqryKmMQHZAA8PFlSNMR1VGUV+4XSAcEif28FJ
DHfTpk44sDcaWIC4Qb7kiRfSS1Y4XS9Ak54HsPkX3pa7RSo0kL9pswGOB/53
f2bP2EnDhVx99GoWUn9UgG7ykiND+sIjT69fTSc/skxBoVBHh160Qc80wg1t
U9uxVguo5MilKscFroFOiNAeZ85HfWt7EM1s7k27Es9Ca5MCwPHyPQ1/oaSd
YqpWs7VdCEspD2ha8Zvvpig3qJp6al3965Ipb1BTFU9C8zqew7fhpppRCwLt
BqIRX1X82Yqku3vhdomWSI3ktrSIgjbuj1j3g+zEPsfFVd9QzIxr+bVZAXau
RPwFNa/UKY9L3EQxwkCdFYPrB4V8YjEB0FpL8feYdRZSBP0LXnBQTwfK9nuJ
dgmM4jENw0ZUQXzFBSmdsKGidKG841VpCHneS9OIZTyXJftUzeD1H48JqLsy
75M9feqcEQD99iqWeSXr2PgxnBHDIYkEzv+HMnUxq9GJcat3pmWnDx5WM+UY
j08jjkFS+AiEcWO/djB9UACTDDljxLSmhLt690RGobFFOAb8ZvylxkC+DdRF
qwSdbGTkgZMPbLrQCMifbMzRNqgKc8STEDZc13oFilxRQ1K4YZUUEgg1LM2H
ctif0OkAC/LkunYB8d9icK7pS80RS5Hk2GpVSTpf4S8Wqu03LH9C1XMj+3wh
Jg7Su4jUhkma8VAqfyzeXRVVf6PjrFqLOKIDC2WU4YymKkG4hzWGcHFi4o8H
vwucThru59uCP9jdoMJ88SmqqgZsop6bNI6FqzLn/AKOy0gdIVOxtmP25BJ1
MyOa5oD4grDV3t1gB0GHOxiCv9g/AqKxqCJAnwJFUn8nDaznf2RIa78g+nLk
MFoycRNwinoo14E1NhNMv5bYYeflpVeBj68AW7K3gFgPMnFjesWnefGxCHxR
uuiIjS8w2oIxbFDXJ1qQ5dYptfKrQv2bxi5auPRFn/W+YX+8R0e2qW8/yzTu
C0YQlkBhFmGLSF0AiCJHA0lZhZ/H0FqD+kjj6C1EGQDOE3sT22S3IpqeXWP3
KXADYxkZSH4z1BlCZsHkGE+Iy9jbAA0328bABm2OkOfpuLAfNZf0rqn9BT8d
vksHGPwLbz3ifhgCqu8z4FcAGaiegy76VItAEbhSbvmir7dI1eD94Qna5VqN
TDZoJTzRlHAbp4sqxYiBZROXegy1QSMPZbf6e2To2TIsiC+PCGUu2+2jYy0p
IvOSqJ0YpqsP+j6Z9CK22++YTRR+LgkBaSnWNvNS0iRVaVtm8jkaPBnIwlWg
cLkv2GgrfPlSJ/8fibGU7eTmZC8xXf0+XJYNywzbyiLAyfLHhsUM0VLgYy9l
6AR0F7z375eNfNscB7ggkzG3kD4Ajj62tsi+QakKYpJQtr5GQhXaNPcKLLmO
VUkJ9O52RzhwVO4XJMXFIbPVZnsyQtLp5qinEqHUei2/u6XGU0FrOJEaCmR+
LGsl5QtUUoX6muiBLzjSUpWKUatJsaieM6sCd1M9cPuDBNbDb5+2b5ZwDj/U
Bo8YU8aFNO6nKPthiRddp7XuoCZBjX3L83G9reAfzo1o8eo+HrZC9sgh3leE
O9tUCYOOqc7YTWMmAC3re+eSyyC87/IGZ4gTnS3dCmjFXxiXcraxXHjzZF9r
LAjang+hLsFgY4fDEmm4BESnUT7JgTjH4N6YyaK3cR4ojIvnTcsz3Rp3CJ+X
Dak5VYvUoQpHbNKuP37IC1LkGa1sqaSR1YCpRg9ZP7zOqGN8f/Ts4qtyfHtu
wUvc/6xbDbLe6FLMGRL8XwK+oMDQ+JUhSPqBM2aAcaylETas3qWy+opjMTZB
1+pRXfhwi1nuv3BcWKM0fMydYlUegCe7aIhAQ9YNp50VXKYr3SSFgHNSsPCm
hR4l6b7kqJatIGK3qYGdC3Gwv0FRU4vifh5iWx7z4QtO73Kmi/jCx5Y8eNul
OGucNlIu0SLNWvWj8aj6oXWbCSO55IBNvhsIz72IFGBaHoxXDwY+XBHS66GE
a4gKJwlVqNBqHMiPi5p9KaEe2BFj0NZKhy6WcoaV7OdtJkjdF6l2HxEV/AvZ
cH4OMg73wtcwADcvkupweBrJRJUiAwzk959OSLnIGmjhNSII7gs+Db3PAOJK
HBnPKJ1HW/M90g+/LBHKva83NbKYkwrbKiiDDaUgPlb0GY+6Ihav5gcecd4U
6Udxf4qgzsKKB56uSG5RbL4cQG1k74lHQIhyTCQOLyWcMSG1/D0qqopGbsvi
D3xeL0VKyOSoq/+G+kVDNP7XQ94cV7F+kbUs055JjtmSDprDDqTWzpwJawHD
0yxesMATL2jpXVlsvqt5EQL1pME9UlR/rLZq/9koWiB+8r8+w0bCMPZXiWzm
w6SSovGet24V7B9UubrIG0v+cbFeHf6BJnwbIeak5DdNUd0jHTNwZrruj+M9
xS4mUxeisL3Xl42lKMN3toaiGUozQiWc+NtmTL0YnHus+2FtLZt8R5Gmael2
hAmFkeGQZgaUudcAzmVJm0i0WBSERxqBXsMEji2FpKzTzwYtDGPHFBIUA/2p
eu8BeA69psf5oNwGebyhSoYH+vCXx/LDtJH/Wo4nskgo/s4NygvzsZeJCOlT
umilRe49Me5nHLpEQ1qnOFyEw7C6yK3mr+6T/QoxOezNOlClhNfPuo7kHnRI
/ztf/bQbIJIpKKkn8hABQkIwcC1XGZrr4as/16bRH84eCMZ3I2W0xvUs8i4R
16OcwuV4brWD9Z/MApGRzWS+MIAYqRdPSI2TgQRmAWBbRJK8cKJYKthmaAdK
uZjRzdqgEiX84bi8PilLsm9NWwUEsmwhHHYJnC5rwFn5OTh2uBSlYiOqwTdd
jWoBB++Zn57Ed3aprzwL5BzWxwCzQ5GOChMl5Lvu15TTOyaCVDXS0XwvG0aM
SNBgZTGqjG+dLGvet8nd6cI4g9yWosteC3xG53BPlqwHDox5DEIuLq0ExVtR
Cn8eYdG2w7CZs60iq1vIBrE14q4wOtrzqSODMqNP2gTqq7IipGo1DXxA096P
KtdBQgWWg/73RGjHN+0jLExCnmjlaGu+0vP9O8Ux+h6ll/B1aQuivv1swCrV
+Xy9ycOfSFw4M4pMAiQFdrSWboU7iy2k37dFBd5Ef2Q2h68Q/H7bj+FckXZG
wjNACd2Iduo71Fc08hmBK7jOZ660Nsn0oe8yc5A5KuM3gONoulS4t4eCVW4N
LoEaPtNug14OQxOtUUPHIKQxZVx6UBp8RVDEMnkA2I8jBkMiDkBM20wjBNSA
1wo7QKznFnWTqaeTpHHvdVEYEU+CHW2PIjmCAQFX95P1Vo9f+RCWy84CGJ9a
EsmHDxZO+PJz9sR+Ls7iUeUbCa97QA7ufua2EjKFHparpRfsUZDA1+KvH2AE
bXGohCgQtN5o9BSY56OiGsucw0uyhk2hskNU8A0s8KOjAFGd+i1eAzxcWlPA
jKLlWm+GVymzj8i6bIfYBWoUPX4spz2QWSYQ2iV3a/5jWiNxziH901k8s2j0
JET9MI1CrWh8fxQ8ZEfyx/xjvwmbXfxeW0ENrbB9LVrU+rak1t17eNSg2tQv
xFjHt5f3Jn78Yb64gx4/7Ph9mcS/zANDcjTSYvBsPdjF1tGsM29bMz+qe50y
RaEQZqNCr817dxFs3TYlykFkpPCZ76oGHcjrMADHxPcy5h1czObUS8oK9qNQ
gdJ0ekOFzPaPTOzCTssqvS7oh8Mar7kw0onABDPDT7FbtDHStLmeaFd9B90X
II+hunftQPE7OyEoZsKIBOINXvPaD9V8nrTw7y0BVWvAGn9OWbFwMtTSolHs
6f0q3XBu/I5CNrI6Ueh5wCsuUBmtf/IoKZBgJ43SsXtBpPelaFnI9hUma9jX
eQ+hjChW0f1r43RpV0k95Eb5pwgHf8wzotHn1WVrLpIzziTSp4CDHARrjssX
h8S5hSfjeoU44XctJ8BPSgytW7PXRfK2DuF0K0K8fyxtSO1V1hk+uaMByqDZ
JWP+wonwf8IkvRRHT3c0W677bXvPNsVc+uhZfBhtObzvWolJK7+2iSOGBUsb
Li0d1rep8mUYkyiEuKXJtx7Y50jPEzfJQMGgRYxLLK2jdolw1ogdLzcbUVAo
HcgAGYxwqXGGfzmfntIGrADN6yATKAevUHVyi7JToxuLMZ0DU8qQ8s14SbFL
vFIy6y9Aly/yW+tFFY/kifsqE5+b9UAgLI2nLaeowMwEqkA8oX+vECATsZlr
z0idEw5iEyR4GbM4nGDXV4unxBGGda+dRhyHoSMaZTZOkK0lI6p70D6NGVY7
wKKqkMpgSwhedMAszv2cplEqT7D1Uh7/BK82pgPCejWLj9Z9EBfhv0LaFoRY
yRL1MyNgZ2+YyuQhoZMLoH77UMHpyuNnTXxLUxf3tTTuZjRr1fDFL/fqOQpk
64tQno0hgVI2aIO1ZLu60ekDNYzJQqpZekGMGHNQrfRhrdNM0SZf21bGJKVF
brjizQyHOZ+5TwGcIyJeTtxFrydBjkyuYeSA42a1jGOjanspov046GoISxRD
JBJf4BPAJ2PWAoBF7Dd6dkGcsNxYanoGbCzxHLAHGvGjJXJ+hBNSTCukkn/4
mCI949BxVzobqVupTIjL5J28GnRfk/QwPf87VBe/s2KGzdOvb7B9ctle1ixG
oty0R3nVMvzJp/NTrLScFtC55rVV4RyOQ+bqHJzflG8R8NgNGXXi/RUfywE8
LfpK/k7p5wGgsNx0C5V9M8FGSwvRrxr6y5URKgO5G7/bHlc+bozJEWz9h9H5
EYghbyanp0aVKD20VokeJmYkfyf9Mz0J8hveGqghn3G/n+D652eSpUxJ78LG
vHYVFdy/tEXt458QMcR5os74kx9frkzheoluwzvfbwfTX2mfmA9zR3NZl/m6
Mrjk71ubQYKGd9KBL78D0nWqOSL3HL8UWPdpNsZbv5T8txDo3liV0ZumdcLg
diJPaUsRmWgUnoti/hzhTs2T8GTBit7wLtBTSWSY2nWPSBZF1B+RxgRDiagX
V8JkdIFOOHi4DT0hmyEANW4qjgdfovAZ5n64eMMxgzBNqX5tphxJG7AiCXLb
XKgdzuugmSR/D6zDxzLFjec1h5/nD0WhBS0MtzqStK00O3aXuWvhDt1BOR75
C+ja3v0Dimf/cd40sABv+FljFfJU924KZfcUuhOQljCWRpyWqH7xDyoW2i06
maACVWRFqEUelbXdN5kyr998XF9vbw6Jp+tHZct6AkC5zhuaneCka2W0qfy7
QzbW2HUybMrYYCl3vBdlnZmvzM+DrWhpHvw2BVjo/33bSgyk0okrY3kekzMU
1VolOAm7QWyj9EXgMd+WiLAUMG6WWpSkfivzrisHfZvk4TpKSLkx90tXDh5N
Tzot5wytNKfewqiQvNl8XBgt7ivV0LoVhx+KbsjXcQeTqexvwdX/J/buQBCE
D8pXmSAXDd6U4syOIcSyggGjCma5XqCZI0O0cYEQG0HTO5xF6SvuEVllH511
A4PZ+SDTRIXbDvtUHi9DCuhB2msrv8jBabu3fzwV+4dhEZwkq4MYhduEHneC
lBO1QERtLii6G8a/MSYFhNVDQYsBRHMZb9783Qi3YCGEuGzolT7Rop+aiMrz
I9vAZyoGsnN7ZV1Tv7JxPJj+ZrokpS0qkoicDnxxV8oVq9EUl6abTXmO9+sN
dc5J2msFnELAXKPseY+Yv2FIdHRRQIkpxsiIuXYqXaqoPVV+wDQPeSnAVg9Y
ywfH8tacR/Gcaenbcuq3tVJwOJ7of7z4pemlZcEd6zJtkExzRryT0+WwfGXn
Hs5akTy1m8YNipWegKCrq65um2dbuBHrpl5Iq7oZNZptrn7zMgB5H2ihSzvb
bbm9vTyE66OTp1HFqveIIabU6vqnu5cVKtqO1l6Ls+OiVnUiiCv3ToYmEQeq
HgXeVJcYUP+balgXWzf/78V4tY0pQ1f8iE5idP8oRea4VmDoCCLYQ5gVTqVQ
Nae3HtIbLoKtDxFJYX7kB3ZgLC0O5rXdThk2nQ/CdqQ/AT1ynZv0oC4tN34N
JTrh0A/7aOMn7m1TEcWyFe02l9QpniOU6KJUeUTAwfkFzoglb92jPh9fMD0a
xhGu8ClbH0Q+lrGt8qAvQ+svz+w+YNYD1fxF8YW1k9jM2zv13i6FL6QkyHwV
yHLz+EaQm58GuRzbx3G2kIQq8thWA+K8LnaIB1hyr5+2Rx3CCQ9MkVZTTQF/
naGhJPfBk885P0zKq/bcn/X7k7sRcuDMJdRgSzsleKcAaEqAEjF3Ojt48IT/
39lgd9HrGCHaH1WErv6BN6hrKc1+ySC3XkT0KO8e2NrvbqzdECY4AcWIG8oX
m4RiUc1b+GRy9Ap6lFbaxPTzeS3OY600Z2uH/Ll7XQgCe+CTx1okY0WkOFv2
g9SH/WdhWrAZ79AWKC+gd1Pgv5Ik/YfHCmCf51jSjMUiAvj/wpoi71xoO8a+
dfxsRN4YIdiD7VJq0ANjOSZYNiiivt2FsS7JcrBE3pNuUSPLkBQLEa+QnBGu
DM71lbM6j9e27sj3XwyWGPB3t9QuFVf8mOBan5+Zm334VOGqb9WMkeBaf/5u
9isKC7W3FvdvY4BeVcbNqS3lWezprm8pVbu9yq+xficn3NfeqEALloXkPLwD
Vasl7hRggK9RGg5DCM7rZ92hbudvX/id2qMdgFs0v3PlX/qoK1OR9QzPdnL0
MUeWnAM9EmDIZCVkBA1O29XCo0MLBoasScXYZLtlsukkQoLr+iKAvoOyallD
eHIJMKevBlpGu326ElV5YK2kRYuoNHsN5V+AbcO1XTwFHPv8W4wkyc48SbcG
usDZlrTheRA9HjrTJE+/vQnuC2QA0TWWrg3GfX/gjGOc7W5Tv3iXsvEt8jlB
eAyCExQGRqIoiI6ZNGhlR0yXlcUTf30RQYVXR1Go4wb2Lj0RkLz0kdiT6Rlm
cWMDeB6nFYV6MlrlA6AC+9kzKZBdPO4p868fKb62kp26V9UET3fWCJ9I4MY4
orKR0/BF7rZeZLbiU5LR3+N19CHeaLv5mXsNzizioIUkq3vK1/dDX+tEU3Ki
XmmI4UKkFXVXCPFRB6QT5+U91qHAUmVOuQVwiRKN7Bf5x7fTVXRSteEIcsYn
SgnVsXKbtDE7mnAZCkk8iwgGYDXNoakNnKtj/BYpNWf6X1WpzdrGtAtVYMMp
75QdEEerGrwkh9DnFTvgw8TJwePscQ0LlbA5kKRAaErg9N0n/wsv99Q1VyDE
dqqQ6oW/hQbiUcrIjFpJTVQyeuSFiQ1goZ3jGNRevV+ktI8GD23ukV1FipvZ
jXUENLccryxUkG+q2XczaQvuN8VI/cuuB7Fdkhn08MJoxIqf40wCZFtaz2JY
llzOwxmLDKoBB62pgGMPYMnCZEtaadC8A+pdtowUUH054cFE/fOflzSkyUUi
gb38PLpDrZjQUVyPOhV3dyDuWCa26DyLeIaiYnZTYOO/H9wCboIBKPsZKxh0
gMe+ah5VOS0GtYSDcdN28wIvUcJO4Bc5NrZVLkHCd8bvHb+G0qzbz6y4uVI6
/hvUGLL4s/61d2CWo26gzC+eSMKhQaQufTEmI29sZ2M7dZGJYvSama9v1WtO
zx8Ly6BANv0YQAqzW9oL4AfpnpRndYO5gyDT7cVggSHYnGIuCNdmaW0I4hgo
5gwTEw6Lp2Malmp7CsF5w0PQaS49QgtjlMi/hcnDE3ZdXVvpodufaq+0EGci
oK2eCTd+zhYuBW2adisx9Ku4K/AIv95zF4T5SKUZhhZISmZ3rb3O+fSH5wAQ
3gTntHUzUQkUhIPo2xWga3Q6YmkXcuv/020T9zS1f4HhzXzsRZs7BM7zh8e9
zxrFj/FloXD9NJJL45fbMf3eCqWTJrzU069gAzqenT66zO6nFTFK01eo0ydY
tdg+ByhCeIEDnM2V9hPjKYCdA4eip9aNN1skpMfzydk3CwjompRtf4l9czOH
ACcu/yt81Lv8I9hGNZi7av33b51FEDQdA6RYwqoTkv1snv6uq6I1gSvhCXS7
6/TfntNGNQNpbL2YSugPwjJyYizDrfGvm4961VZYYdhXs+nlgGPpNzkoNpiZ
4QgidfI56sgstKMZpodi/KF3XwcQtH0C6fwcgsifN27g+VEG4MJeEne4PNRy
v7p0ZAzZiSP54ypCSAslMSCpjRkfV4TnzTUuj9FtQyIuTuT9Z1wl1KtgbIZT
QqzGVAgyIY+Ebh8b/9iu5RIfLi0qMlbLQuSefX9q0lMOlzXfxUN2UAfHoNrG
J68Q32h82cNrD7rUW6897x3rIBz+M9ThSWeIhhVPzoth2SNrMyUz8k9gorJ+
iPBm7xJcYlwttK3vFWwsqubMt41k6DmxyIhBGgJPMeGKgC+eIJ6247EoW/t2
f5CM+imoRfd7/hyIGuZqSCMc1zI7htuDqyyivzVvuHGOBn5W1xrvtIBA9yR1
PQuOAxHYBEdbvTSYcpPkidtGGcid61C7IcjPaC6+7qaj/p0pjJOwtOgB9/09
lw2HwZosjhCMsiqEZYpDPyiFDDILlXIAv1211pwa/zFT1XKe6JC7h8xHQXtN
v1yLBDWhwtFfqLemps4w911TflMcaB1BMpkquvam4H55F3+7kwGpdxlzX5TS
d3nHH4JUvrF38lPAZWmUbnRRZ8Xy8pVNdTHB73KRS/5eHmC5hJV74Y6P0gqb
3XIXH2ngSF/zyI4TQ0VrhkGvIERpXKWXOMz9LSfD5QK1CYVNhXFMFvzfaoN1
q6JQGzJahOmxTeKV2voal+Sgoxvn/s7Cls5N2ExVELEnrl9ee2pSUW8AaIdb
7Omil1/3dDQgkhrMyXJr8+UynfskD8tq2QrEFRThVNcy4huJqDiun5A0RrzK
dZRPDUt2VMV89ghc2MvfbQMi7YrzVcKIK3mxXFIJZi+XeGBIjcXSl3cormEA
yP0xTg865LanDdRR+3Mm48agzCPxEo+FRoh8Nq8r9eo6RgjWMHKu/3MVRqq3
x4u6T6oLKY3a4x5jGJ01aTPnRj7gMM+SIDShc5xkVypzJhHDl4vkCFMfSts+
KLFC3th5jq40K9McHqM9ID/MhVl3icQrV09ipJywIjmXlNzTTgy8bmKtu09g
C/T8ncPofxbTmEIXLn1PobSr3tMRWzI3MwZ0JLwiIBspE2w+YK9RWRUZGieJ
TmIdNzt9Uu4vd530u7hNpmiC3UKWMONIoucncHVrkun3zEyeqkOMu1zVqAA8
14gA6L6RNoUiePpWei4j+MNQmZ37/Ty9g1Wt01tI8SU1KYdFQtIzfgS91Any
q4M/5xfd2FePTQjd1OayZGJlloKxKiv/jOiVfvbDkyVbUCbj/9SmSKWAwx/f
BUbKNS7xsNrlykS91hzxQVWrtidAfLYRVl38ELv45htEMSQfalQ8iMfnyNe8
wgmuG2n58WRb2nIR2JKF4HR/8Tu1/wqrXoRw+yH1gjwV3yf3xMcaUZIe/E/b
YZWChzxk6+6VJ9jP4Q8sJbXsyXu9vRl4pi9M7IzqhVwEdb2bce60Rek1ob12
fRjNKnaikEszFkflrc+CfqfhgmTI/fw6y1IaqN+Q4vtWrdyIgahPmRtNp4Pt
2TVDIgZgPQp0bTkQ59hb4KKFQ3CuExqiwNZpBuHAHcb3TiH9BmXEkP5L8DuO
dR6ZVek1Q7KlhxXX9k+n2Uj6sQXtLqwe5DMYeWF/ejUYjcKzdFQtgZLgx+r3
KIqDgCWkZ0J5/w5iKsXtK/D8V8dI8ZWSESHXOwhShK9SVndA0/YXMike0Xas
q7/sSHwxOE/o2TGBsIysgkERwkYJei9WIU7CbJiZ7vixy0vp0WZV60OIGNTk
m2zO8kzVMg2RzQFqQwzqMo6N32+akBFqNQiVdtVIOnhqVAATqT11DnyqohyV
jcP3cCrGYLilMDBQ1GHVvgSOYZ2SESWXzWJ4UiKBK4aR/V5BDaWkThCugT99
kRGXFblHhGUKwDh5DN4tY5W9GC7LarK9smfTcQGdVUyL2ZWvbFAjNB+0juhz
5R0FtWjKsWB9YkcLI9Yq50Td4mups3+w4iL3NxMYY4Xbwi2SlXP96Ii5UnFu
jROJng8hkIMlf0ERWwyO6p3CqXeXcQoeCP9tLoWq/3NdmdhrR8T9P5w84vqP
6TEPnN+li7z0zZnp6o6m0BSpvBIF5t/F09+4Clw3Ozk/1zfWsIj5a7+6B3JJ
Fm8cq6MqBZ5xXFcrDGRuPb+kJv/2TDuAvfVkEJixDCievpYlnClsHGBck8u4
CyYceC+KV5IaBZdXUEOdc4Iyu34SeUOWravSO/ASlZqTXLemhp4DNtUhOQRN
8OOb1b13v3vvnJa/CBop9Fox2GabD37aCiR+GcPSPcDX1vMuMUJ8dv04DFwg
MOyfbgLO3pzY6lBbAd7z2896rRzbxwutrsK+9WZvokqfQ73YkWPVDzRfVN25
dYO9y8TT0QFhgQOPU0tXeJM52xBwn5bMOCxEJh24Cf0IClSaaq2S9xkPVScK
kR/hOcRBwVaN2J32GuqQtXmCNJ9XoEdH4mSc7jEbj0G+bIBDt0xfEcM6slQI
4Cq3f+FslhU5Cuz0ZqecSPk4W+9FXonmq8vXgDnxRPpPfm/r3ikVZ+3Pm73f
0kD8WYvnIZuQJNRenMML4rSkXrqGmgYmfS6JrLkbDkVhlOcqTDi1AjB1OGYj
y/+N6fNdFf1Ri/pwuScunztqzxq/ICO2naHz/Dcn1hbqeQnadpKCT9QRGQyr
dSVcQgr9Tkn73xwx8hDumOd8mFcvM79m3+TRjvncHNSduysYt3rCZ/ICnpIK
rYFu6l5ssE/Ch2RHAXrp0+b3L6GIrKT1rhne3RbOypSJGsBlB03mRaGjG2AY
/EK88mdagUwfARCBsKWMZHMoy1pN0+W421rUVucuaaIpP2TQvbumDcnZJ38j
pUYEMnRYFwEJ8CqFCw5LnwsK8Ay+y9cQiDBXa92zWYx6EcRDSFFz4Yxj38El
A27DXvcV5P6u60DwtXicXP7iNb9b2JyUHTEjr7xd65bKjy3ZJRwQvSjXW5HN
+tTlkIUr38PxLpI/ElSQ8TSsYkcDf8G3yWmo6cbKu0vU3JV1PDutrNsmiq6X
R1BP5K8VoX1UMp8ldkIu9F6qLiDG5rAhz7q9xhwsNOzd0Z1zF1m/WXhJN3V9
ZvN/g4FKrcXZ0yKaG59XzzkjfCtR6CP5hHH2gdgIf8yX+T+xq0IJyFSmnbNA
7WvHqNk2jOBt7ERymigH5amY1VkNvxF3iC4iEByJ9CUxA0dTPLcP8zEVc4S7
bjH0PQV0NDQXs90H6W1UgMdzIRneCuT3rmaiSPe1Sxuooz2QKFhasxrQ9ejB
qTjnBz2n1VADt3awzMzMKtMzRZqKtAfnPyruDPr/SdNubyIo8Hyz89StinH6
R3j0+K6Ze8vkFcQCQ+Rp2UQy/a2t2n7N1343AGjj5DRZH6mYnEiQZobsq1gc
dpOBdQeyy7ovJfM9x8/75ZcDg8/a5/aKULq+tuMJHdRXUQEBeRIFaRpL9Nle
pOAHIP+4Y+o+wlhG0fcNnCY5SKuBtS0J1nO+x6oGplyb84X0t5rY0aZYNi+s
K10Z/AX3PO4tMnPCUaWNitdrKfNbCZjIZbZ31AvneDd8EPcJc77Ecm41K/RQ
2iZrPBMprRquASjxV5VobQJSVgl6PfRTjW5ss5iz4hKnG8//E5EewGG1W7Kj
7f4/9TxU01nL2o4Hb3Kl5FJ9x70nJw0GRvGYzZ3z3RpkGuzkPocfBPKdwVLq
MF4rvTXKfXOj945lv9SvYFL/igMbqAMn4OEo9uPg9GD98inbvl7QbRnFIfaI
ZJh84/aVmBIxLO7P+7dJvpHupFFYIuNRpEHLOffJKb0QZo2wiBHF+eXvgLN3
6gCybKR2sqRYTCbEguVqCaA0N/6nnDI4o1EbZ+cm7Lyfs8mknE8WXY/i+pSd
1CDEfx5gcWkeroSXyPYOoS7NcMWrzicFsHI7Qpv6i5lGCDoGfVCWI+1zYwoD
/HLHjwXYRaVoeTHPsa+NQqd4eKujuALCqaWH9crbUTCuk5NVJWHUlaExyOkC
K8/cDamANfHcSx7z/NdekZy6CQUpRKSbLiz8W9S50Lrou5iabwL/sR8m1l/F
zkYiEUN+ljdBbGW7aNy/eClwLoFFclP7/KpH0MZggbkcL9gdweaGzkwKcdzD
lzcUNq4QPOuKAVrUSjKEQHHyNIvVtjdLh5/U/Ld0B5YgpfaKp2m6Gqcp6KnA
kjYpaDk6q1tqsS1Ij6StODLmKbUa5gDPJ1a9KEM/38xJP5g9h33lnA9u4EXX
kZdwinlHTCr9J2GUf0AGm4Nx36Lh6/6fi+4m3S+VuI0IFfEvQoJPl6wm3Q6S
a0cGJ3WmY974VZJxSiMLIxGHbanLhItx2XXdRd940O43AZ/HySrlIziz3Hcr
90YnFM62ONjuL0WHqN5QUG4blqWjEluLLFAM+UdS9p59vrDC1JS5N2TCq6I1
tSGpva4SUVmXM0ODxsliGxe8RcIZ98SGQDYI/p12AVOgBOIYGxlP6lUc5TEV
QHPqqRbCayBSaZnl54ugpVO75mvdUmCXGHizO0LlEAUSAD8rnLRkzWh+Uc8X
tIFCgs9R9VlaTJEOQRPxfmshi+n+SH/dCYDlDYKViAfE40cYji6PpjUrWX/v
uKAa4HkNdbNFdsgWGm4ypz393dIrGG4nBBVOHdBleYrx0PBR6ko+tEoGmctf
QTFmmm6LlnpZYz0Y8LoSzInAnLxZHQNObf27axQIocjb2gesUsi1nSo58+qb
2n6HIPkfclt/gzrA/Isvpb7p6vKEkbpwSGVQX6ahuYtCsrOlDDdoVNATZxbp
x1NauPkcW4/pbk6aVYcIhFjGoJUw1ie+50HVErxVi6UYAFhCqOc/MOIgikLe
CwnZsBu3tE+JaP7RK8eQ4dt2geHuoZtX4Mpc4Ll51w/IEM5njQpgvHj2h55I
1ao4olszqSe8jTH3Oklj/8rH/k3b6swSrLicr4pVg6GY2tbzbk+7JmXcTl5t
TBPLkYOVa+dVcGbwtm2EaA7XibuTNzDdHdddDt1UBSJgUVBw2fIAZ7dcNuH3
lRVrY2KR1gD82ROrElkjc3xot5hEwsbsMDx6DhSlRs0pys+6CrbUjpONWOyZ
Y9FFZApukw4fhZUxOv1LcD1kh+H5XBqO7PxMzLvCjfjLmOl77DmxiW/qbeZi
i54ZzQOd66gEqkzlrkNhuD6e1GVhJQlc5g1g+ObZ1LPXOALUEqDMXpX8evT9
0lgP1LVfQo5cPRX5jMFRyOP/mS4IJdUgBWn2Se3ywXPFWJbQ5CDEzIvncw0U
2UnT1jQGcs26OEq8u/HHrL4TKiSNHgPtaZxchAhBFPug1FIYYlwR9fdsO+dS
dIWicCjLTNhp8TBbL/REifbJylCDVvPewd61d9JwxVqcBITltbjIuYXPMYUQ
BMuHm9mj+l9zg3cxI5I74PgH/7UShMO4enhcaSUV0Lk5J1r9CgRtiyhVa1M4
Pycp5Njw/JyttHWnxDedR4+9r472R+vIYGQfA+hRH067xvomAdP5qpFJO5PF
+ki3Sv3dM3MoOf0z0QZGpmWdfNeiUjqRNdwolw4vGs/+1ZfhstJ0tUgp6W1X
iGZAOOTkfWn3DubjVPYkFI8haM0Oi7M12GcXYWnWSj208EcB9YbMOpuUHCt3
DrHjoERv0dPH5jW374PAe0gvJDkBkDFZ0BGByhGtpp3O+0AQp+QLaZ1tSSCe
UEDAlVQb/bsYmF8fSwinotQZiMYlwXHazDfBWaLC4ujkzkPWz7E36QHMkIys
zT3mwo0a5NXsYJHk8Kqq9QnOqdGUYseq9JdZzB9Yax+p1ARK7mzfXKjTN82e
nL7YzfCTR4T4fZ8ZId0bWrtWc+JmnTQJvvKsxkRe/V8uNy6dfdAQSUpLM6Ux
RL+9uoqP44HuMvOfLN+n1udDsAsda3xij3RiHGSecTi+t5FoejtemFqiZ+Kk
t6d2+lEVXwwQeM5Ey1jekKFhopR/sjfPHhB36Oh1YR+H8NRNY5qmSp49fvXU
fT1l5NpVvo2LhKta/f2gBHOKWKVuRAD6joB6tXevvKM005XRkbuCsNgQYdap
hrAOuzQkxu9bIoFnDLmq62xnXiVVnF3frOr5wsKREq5eMo8SuDL55g2NOnm/
wx5IEUazAuvNXbHPJVn9U0EMJRYxMNbLDH+TPEBbn1JiB9DyUNtwZ9fQFoWU
7+yyExU5pxePLfyQ7Y6R7yYpq7Qj7+ZMTXHkildErt8ZsEL1LRgx69S7H7M/
CfUvFKHEd+0dbjIpMgcOhXtQKpMD9aRcUrt0sHqwPN3sqMcDqnW0KbcGwuqa
SFw/DsQ9SU1N0C9wL1ip1e1uVlnbwL4q+QnoAFsJ8Mj71tDv6Waq0oEiRDF0
mCfz49J7AHN7GtuIEeUI5OY9vRD7Cm5X/yJcLVKvdC95qSQEwYagoWaOY1M1
kMI7KzeRfcf5cp2X8AVXyA5C/BGBZqfVSa60C+Tk55bFLKAtcJfgvHY/X+0J
7FmmgmyejP1sbiL4QC4o/dxpSP+b6F1Y1/Pur9t3X5/aHE2KXX//aHFOiEW6
m0bTFNA48INefbERXIE1CoWA5KGJrw7Pk6Ah2qZIr/2S/8/DGffyiOIeER2I
5P0e1pI5o9XK62Lf1hXVZn7YqVA/MUaXvygRxiSUeEBxsbpx+PMih0LCkP1K
nXnaYOyNVoXil0d3iIEQ4e5rU7UREn474c6AIpbaz7KYcHGXGKoqMTtXEYcz
R4/xvprkSR73pRqpKEK1LFfmvxvBg2ObpY/lSegil56JFMWPV1qdPGzQ52KQ
TM21WIoH9v6x5lLCk9HLWQYuDeNQtnl1nI/SlE0CTIg3+M6S5GplE8VHNcTK
ynmuUS2ZlixLKaPssbmlniZGg+zFr7ihr2bRIz8jqyBjSxsOmhiN1IuPGeO8
mCtCSS+Y4HRMqhao57K+A+nLegu8wZy8CQHlooHW6A2VymEdr18np+H9gTEz
WCeEO6Fr68kvettQRSX4/WUp+wV6TXbFvTg0rIHq09fAnUN4LGAv88p/VEmw
39TB1nHwrcXT0+lk5PlY3WRnGCZNiWd6t9Op9QPmB0mZvjGDK72DJ2p+W0uQ
bg3xBnmAP+GT0nW8L28ZhGTGE6oqlD+heEDODC/4iBdezJyIDtIk9NxQfHYU
QjFL1YIToU37U8XdFnJhrKdviumMVEJmWCMsf55b0ehWkuy2pa/vR6l7bQUj
F7rJ9+Qx745TFNSAkP8m6LfkCgqMGUhD11xkg97m3atYVk/w03hfVTEaTOrg
84+x6xk3baC7pg/1NMzV9oZhZ0TrM9pWMCkIuS7dndaC+J/U9hQQ8Aut8WKu
yv2CQBLcI7PLCL//XrmVhcPTGIjYfEPDYFldBuonrpt3eiTpozkKb26BTOuA
25j7n/o7EpdA1SgAX8T61EME6zwJe9414cQX3KP5mr8ASjNEmnKyCgjn0YiM
44yCXc9NDpa/dTpxZjoG5RAhFUXHAikeWPOrP5TufMHtH7ub1o2Sc6uDLWB6
bMOrK++UfAcYcDrsRns8JVnIePx716LKfRhypRat07Nm30eTc1JobghQ5snH
k7ZscFBz6S3cgHtVwfwArz6WilSazQaTa5mK+/ifqPY1cFyjfACHrClWPeF/
dXwGhXp9P7lmkyrRBliFhNJXDnQSejFD4j16M1h5+azc+9/pHUwyefbQTmcP
+beWK4t8K+qvuy8ys/C5751Sqys3p1JcxodRPf1jaztgUpkM75EvmyiOyXqn
d4aHejhY3KVDsz5evzHtu2yrgvRRPJbkOuyTF95Dl+u+YGo/xxk9CHOxNcMt
MU0HyvcjOdMknoepqmefQDjqP31R9YoSLXIxDIHWEAdhMSjckMUATaLV9o8a
sO00WfsNUv+6LhCKM6V++a16o0k/rX7xs1z3FJ3ikSpksXV8vV0daCSFevk1
LfynDoAqcFn5Ayd/kham34XEYTcLAvqG99GkdgyvtnTtLc7mapUzmmlGsyBW
6ij+G3ISXlu9fpgXgKgqWKgvkaAdMD+aXVwnCN3cUbC6fBKH8BZaxEdeQNgy
ZmU5/boj2Bg0GYLazIYmsp2ec6GgnvC321TpbEyMLr4yv2F97a73dhIlJtuf
Pn9P8r8lpKx6qXysDTzfFp4xQUhHkZPerQVqmSR7pQ3FT/mVPycyR2DNiqJZ
pwEz0XRH7hcw8+S4YGjyhKoS0HYT16Jw16pupruqsDsFHa4M/33AjKkhFYKi
T5Fnp2u1P/51TFIOnR4GnWRD9B9SIFQdCs697JC1AJQ14JrxVo33va1BvIhP
4foR3FfxPXDZ/e1tWa69Ls8kN4IcyeOAKnTDTy9DoijWkfEuxbduqxWOVwZX
XTkT7/FkSzN4pgU5vhHBF7bezhb9eGvM93D6Usb1Y1wQuKvdaMKVFlH+JiPb
x9EBea3WON+a9w9ZraJ5jAGXIOsNlh3C0EohWM2xziOeq1Oxuckqe2NIHwO5
YEnyxK2wIaDNjTLl+yz+hBZwGgwJXX0DfMAF6FdTra6xWwwvP5ij4vWvGFJn
B6KNDL1DbrC5V1i8VD3MfnH/p7U9bf2nkJJpVmNOeJtw7o1QI/1UvUz2AQ8n
eWyytyzaLbwkmqw8fNBccLLXhiz3VF6Aq0v5S9+baHl02ArSPTq2ZXk4UHav
TPfJ9bT1gDoB1v3m8/s7knKmpfs3cCtG38zo5tMAPJb8O/ej6KbFyX9R8rFa
XX+Rg3DhAZNAQfIKrZWVhE3MgoNG8uQIg0SnWlTJolRlp6bWDjHjU2v+44jw
fMdkmvgcFfBZJh3cXVD9QVuJ2uiAiGlm3gGIQkEMc9Vxn/6vyhyKWBO4E/+u
paa1bYJz/C2BfQwBu1/gPtgibBnRWXVECKwOinKpYirDA/xlloQayYuaFSMo
+Mly4LSa6VXopQZiOK6WgOkt8MEJA5o+uz8jihTRWeMncEDpQnaMHqQ9CWuf
YrleroEjNJkJ97EdEgxRWCFyjNQHuJmQaQ1rsGnOsMqYI6htSKX0/83Va4J0
sT8wMpgmddlPib4AGS9bQUuDPqky70oF5bnnYnJeKiAnarKm22bNpx4tNDln
2LpTdQBfaK248fIa+0oj4mS36IEAMeAzXM4h5EM1uXA5l9c5ZtSjPyR2MO92
eLxYV4Z4fzb5xz7jujQDFK+GEKSbQ3NO7OB2eMxI+GGDzGbwS/8df4nMT5WR
MBOsx/+6GWLbfutaFFRl5COoO6JCKrwL0BUr8NMk/SuuySJmFjXxWLQHphx2
c7PSOHHYewy+0i6tnzgyGUUKLdHzwZ5ZbwxzpMNWO3/MRoaKcxU84g6NhLPL
cOe5qeDhMlZsbUzQplFxox4T4sUxPjjuir6DH/jz6dntJeiuULHaEABwv64E
Y0ZU/HCvdPILxKW6QOz5pGXSsx5lekluAp6p1zoRReP2C8SQ4qRu+2N9oX0z
7vEwr7ibX+R4sB3GcEddDiPEKW0PiemeJ/iBHIC/U/gcQyNy6qkEtQEFedBI
xApll9F5PjMINQjgUmdGo8WyTkxqx2tQMmVwkKUXnMWFSPf8fNIIbl3h93nr
6rYOYQ9esAH/rYEIcOxuXYlpWxmPrTgoHlzQJkgPipsV+hxqJBRQm8mzVpDl
i9f7JlaEtmVZd39azcNjL/IXK3EJJCgUDQ3FDrfc7YPdobB0iuRfkDcx4trb
ZAcmlyz6opp6BHrKUGEPqRPqhopC0504paTYuqRBJP/Ba/hLij/KTsKd0Akl
CJk8CZ4AOr5t4EDF3bUAT8sFxD/vFcv1YgbwRqVWCqnmi3rl6W2lFdDFDtTp
xfpNgx6RLFGsqnHmS1WJ0apu8T+Hvrgz+Iyz2WP+xQeFYiU6bO+4Dg1JNxmj
umDb/z1tdMrubveRjYs3q3vQvjMfYs10apsCJNZjgEwDPFT/YmQGVV2/N5jj
mWwJE1x4b+wryX3D8pT4f/ybFgVJqL3yD4SB7n6pmr/pN2drTHNRcZx9M9mL
DDhaJO7IbnWDn0dMCLaaVNciDJDsVVSCm65Zto//sLFsXZozFiDBKLJU4Zfe
PNgPl1vrorUidgc17v1uixxaqVjGrGNU/oNRC/fwm6WznXWjGUOV1W/0/k+n
vS5ly3n8s+7tgyzcTQb3A+raO64UGyaBUX4WjubInKuQPGSbCw6lztF/VmPd
mTVEqDp1PSkdKJSpp+8mqawmPJ+w4FIEpEupypKOjXkqBD2SL+EGC8QaA26c
CMrXKT6V2GB4+GuHUpHC6rbuyrsdb40prPG/gdq3WU42Od6bjhW7kiJuBbEf
J/L//8ACQGYmyzDM50KUaOM+q+NmcFPTscJDJiXswxsMfizbnI1vcE5M5Vck
AyQZn1x0TN4eX+IBLqBTcMUQ3GAU6XRm+7T5rr75p+A8RrZYap1Bv1JWhqpL
dfl2iZkAxPhQLu3glJ89kYmjqx490HR44ErPj7kOXrkaZdXh4QPAMKb5AeOX
ztWQEH08/+kTCDiZAxWDfMmKJIwBJ4GWpV0Q+EHbVykoprIXlCanVYYiux7f
HZsC2IntiIrM9olF1nT1jz417Y5/aLZfPXdxbSEgB2NwGqFklGX/NG1Xax+0
GbEjrvyslj+CLHTBDjOoeo5IdogJmixgKHxnZ+lhnbLr38ojwyqPOOOfPuTP
kx7sNF9n5VsdG/GzU43gonGHmVwMwUCW8XQHSWSKFquZVeQCRrmP7AjY8751
aeiXhFshfLaWTR29/qT2AQuQzcdr53zSj+6V3rVU9vWnUgE/FSUeXeHiz/9g
2KYCR7M2LN3R8oH5Jx1jxmTSn08aGajbZ4KzD9+DWbsnWX8tgpP9sWFFanqE
bW2I4McxePIHCBIpP/7upabmnk9xTZPaRFvF4d2JNISWkyH7AFGybRK6rU2F
FQBtayj/V5DfVENK1B584uo/xaLwwzXUrLIjFaUnpyFNH8V7izNYdiNaxGyG
g0DsJO9oLsEb3J53qB9Dl0mu6QYuNpV5KfjsvmaRRhwBr7hO/nX95dUEUGoK
4b32TqLmUHioBOmqojhUqEGcrM4/j0h4sLyRUHSy0sxSCAQudGll9OFm4Vss
7xLnI2i6OtPmqTFAUT3d3jJKmEVN4mAirOl7UfAi+WcVhLG8FNW5E/oTTJUB
hcjsmNtXa4b2MHFtK+07VcW4kowoXUqba93VIuY1B8671LYeIevSlxfBKxAY
PqekLVA8X+fQMTdZ1pqEMxi77yTCwMHAaqPGMzhmph01goHlQaOynU/io8Em
2aj0M/pR2Nq4EynN7LGRBX1DY2+yrjb+iHCcMynisVsQ4HwyETUr9PBzL3EV
gMuoo8Uo8ILI09/3+4X2zmehvIildiDS65aaXnrCv/xfZXH6O9NVhkun0fKX
FArnkAfKFfIHFP7EM+YDuj7qcJCxGOShEhCREVCPkWQCzfDrrwAyNCalxOAt
wgrjh89oI16YD4G04TFLMZlB7jzKzGvKe0P+2dCZ5fQBQ+j4mTdvvbWIYi1q
oznXqhjz57I3292JVwQDPEE6XvyIlLPF4S+DO/F+wSVWz2YGJgZwV1ohD/Uk
2bl4J2xtUouqreJeTo8SrpsKmAgpuGbNaNUzc/E51knDSKhsjVswsqHIhAhY
JCYvqGwcdOYbLg49xkwdvbq8KI1blUTnW9dwC1Zy8LsGb4MWRTp11IIL4zUm
HcqH1eQYluz4CwFYyQVvzrQN6/glGcLInQvmMrbklYv9qD5kGh49DZyMN6Zh
AfwZl0PaGGtPY/W7L5AOkJEJIBw4SJhqki/hRM+1mBeGaZQ1lsp6BU5paRH5
aHHialSAH5oppAeFbZWdR0EFw0IKFQljwWV2vLN3MH1yWLJkyoyP499hTiIO
xQ7eKNapkgTXEFsi7kSK+3mimAz0FrzF0Hd+3//lTd4P9pRrZGO+rYROj/Qu
le/jzXcEMgRBLAexEQn/1xWVStNtdUSn9dyPgEPbApgo/gKIuWzIAMyahKA3
H4B8f2LyXvQYi+MmM1mHKnPee5fG/yfJ0XkrTZkz5dvNhjP+CtBzn4QzpuT9
xM17U/Rz3ocNKXR/4sO4jsYWqQHPC1N2+5ZeUQNt7QNJfCfvWmMhG7Lz5KMR
WPWz2qmxeAyxHFy2EiMx3fb31H0LQ6EFfQX4o8/Uw273vl9eNdn0A7caH4hp
ATT2kx/tDJe8qrR3nLjzQvYq282WHcuO/O7CMq9TLe1b28HSwz0oRiJBLkNG
P4m92oLEo6tG+RvL9TUfJmOYSJ7/ytyRJD4K9sm6l89+HqnsbN9xbSZElOGb
rHHpDhtQhei6Kcmcuit+KKwYYLC2anuv/Gh9KXio1tfQrvBWXGIE7YeNEq2C
YyUnqPvi1VOF3ueJ3SqL+KvAvXX7TqlYdcl6x/bT3TAf4zbXMTvDw5nXKosv
+d7MEjmpEfr7UYxBctc/MEEPjDKtuoFvC/2taRCqYsmW801l8bcPM2rmCIRf
nMVELNRWAUbfEut5dVGzLvLptBvV65fUqjBzvW5MGUWM7nUX0BA2oG9aK1dD
2AlJkZfVgaHxk8iAek8NJkC7EqazEJbzLny3wk5U3tRMsqC/PrTKsKmKyQ8L
3+wXK+UUiUUvKl/Xk3ELyaweNurO9xrHjRHzr88qFgJb5nrHRihnaYTpP0ct
5IU/lm3LfA9Whou/raG+0/Zp10sLvniHrvr3dUXcIH/iW6VRnfQcpY+BgyWh
X65pkEMy+7WMUk4jK/CpfRSsVzlCR87zlZWNkNl7oooVrVcqR7EGXOOQ+MB7
SS1CSiuG1cZXMzss3To/VNb8PYbDEBMjE9upnCzCXASV+VJQudtqLZrScLlx
skM1wzNyWjAdBJVGNBgdlGHAboweE998ym0qbe6PXcZIwu6biIf9GcXtn2gK
ef+3XKvlrAOUN/YviYbVYlndv0Moq6KYFpm/Z3GY+4IoDmdo8dz23Iql1VQK
MjPz6jaUiHyGQhtRxHXM4u663kLVWBgc5PhDpQn+XC70cGbaXgYmitfV4XHP
8J8jbYqHtTrdILLbBGphqQXVXXIK2oHoNOGifjjU+2ghaxAfC6OZUbL5fKdv
DtpHch0k9Lvnt40LrpbeyKUqq4DS34+cIe0LwaVXHKHb1V0G1NRrDxB8eDJr
y3oWqOAfxYpc1aUpx4JDOJ8rczTzpMqqkxkngD4+BnaX0ZSDuNgxnZwcHB8/
ua0/412zP9z3XEJNaSn+e3xA5VWVN30heWrQ8IIcr1I5MMFLpdwvY6ptgtiL
hmNHk+CVzm865uvgqbcCx6lg4KiCQGTcyTjbPg+D/fNBB89sURJAK2YKFaFZ
aNzdXwqJfIuFf0ED5A64ywbiHEcSevxi0C+E6XYUuX+i78aJ/ZX7e7+3sco4
fZKd8aTJfQZc2dPXydJCgEfJ1H96rMr3NA3QpYV06NgKIM/8d26Tyzb5EHQy
HLOpIR+TjYrAVtYH4TjKr9SHAYuZ3AhPP1ZRHfDe1wKRxNnA0MmtRP1O5NIR
U8/JSaJPeC+bL9nfsL3VKw0uSOuSbbULwT5NG6akQEYnTug6faZquExft+7C
6GO5jm06gZQj+6MrLPL7Kkpvs8+KZdO4M7bT+NXjLRgmPhrYfYkSGs+HbNcl
fhdfjfaxORlC7WErlG7/XJpqKMOEPYMcVPgEMz1CEtAViQMPKZ3+iIxZwhOX
NGB2RlO4iJr9nnBOXIIzq386DEdZUix+UbEVJWZbLZah+QsJmbDo+xeXLUQw
d2fMBILystBOErLjAsbzvaChTzyFRkfokFKZnQkq1Kh/7vTnSHOznixuAIYA
/1vMmDMXa0KzrmPRxj1cqheuNiPMhBLeDp0jqLTQDOzO7TIKanmEkDl2EP1x
WvR7aNKn+c+htGnz9+xLova1N+xqGpFDSIoEzSwbl1ZzcwSTgXoyiQa5vHzI
jnG4+IJUFkHmD85PXKxK/qchfPB9SdDX8gm+bw3/4o2Y5iTpNuiZ38NxXxOB
/LNiu5wEWM+baTd46q6aNw1IDlpCjtl968UNfzVxF/4Fjh/ttfU/P0qP6uQX
gerMP70/iUPbLhDy/MrUArh92WIDc5py5PsU+U7VcZpbUnwMmBHaEbsU+YwV
9TpDDSp6sB486/oYdetq6dDXeTtiG0o1pwEsV67/k8tx1larmfn0PHdIfm82
RrE8gvR8jIpwD91E6m5vmf0FwZzpQx7SsQHrw1u8w4qmpohSNvcwCGl0XFrE
9ltISAMmFWqiMwTp3G7BqtTLucSyA0QAjnaM6co5V1TZxNOEkj7IGh+Ree3P
V0P2LukdiOmiSwAAPNTaOoezuC+WETK76AcVQzFtK2ssJcUCeWKAhiZaVpjs
EcSahkx0iz2MTNah+tlWbJRSOjzaQK9zgon/HEw4NdCLxfLXfCEG2ot/U3QC
kOhz6uBW7sCOTTJdLmNcVAwTyP2F+Rkpa2DNqtGuPn3UCibuxLsRawCFKmqV
aAtQaLkVDrfNrNKBXxR4AGe5YTnpgU93pc5uqVj3zSkdmqxPVcMCADeB6br7
oifRCzYJ0ttmj8/qokEh4c7GVQXav3Lno0tSP7CdiqGe1Y9nk+Q0McL7NePl
J+/jWH5mKK7LCVRz2cXmsxTEVW9s6M6MYzsW02eKnX5xdGDJ1degeyxSLO4u
QoaGdMp6E+1ZUnsBF/xc4m5diNPnDhieJwP9C8/BnePy2anW4Tc3fEx4A/Tf
ys7AC9+6gahymycDcUE8KKNT6Kdd/WuIiuYkiaBuripdhm816tpYsn8U/F5p
/ipeGcOZSziNutMKbg4c+aocv9gV3zjnpYJG305/1gFgRXqAa9W/UdiSo4Vy
zjIb8qMXh5RmqKen3IM37Dqr/j40tolCSYrqgP76t6YYRIuZJ4PzMMrAIbYm
YldEKrF9yK7ZLKuhwtxUz7dO4Fzin+q059C9wY+CHawOW4AnOZw/p6wpNe03
nJBsWXU+RCPpJ5NUx3iQ/6szuEazk0XQxuHRkHk7ssuF/LS9lCHyQnCW7+D/
KxNmXgY7FdyLNrpeNwErHFZSKNPOKdcLWRzsSuYcUb39zsLLX6gDn06HfGsu
GOk4rJx82wYjadXD5TkTVn/2btZUERbHKUVW9Eg0SrguLRgmLsudZFIDxEBs
BraT45MSQFZBO9kYfYNK4nXgjLRyhe/7pggP8O5i/JwwqE+iMnXTaZQFiUlF
xA8h/iL5baC1tXs3Clh6BSIcSbaOhEFsnw7Xr98AIw1vEXuGsxREe+MIcJU/
R0wqmdy74j/v93JkmCXFI6ZPSFWI6Qep6C6vkMOYZ/bTW8hIBlKurDXwoiMG
uXYQIbhyJGGzLQ5b/AMnzcSbbxqvig4nKR1ESFTcy8ugXyLRV3hE+TjjwQeN
kxOMjflAthAiLJJRPo/myQTZwzeX4/WrFl3q0HpONvZi7vPy5/nagRyyxH/n
Cc9KgYWntQvem4B08sSl9Hxmc+sNmPKQJQfH0LsHyCVm5d8qZuD+XKn5lVr7
69EawVT57BAXyfvqK07SVeL+0CROQCt76MnUecL2KUEXT3Sk+3NrDtOs3O9T
4Uhz9cUY78uOTuGa2hSgs3TxxfxdFrwhOguEfNToElGR5yDz39Ndh11SFPFI
6kB2zUm+d9eQvlLVxXlHm5wxkLsynp7o8MqB4eTEJ0G9KE8c2CmcmxS7yUEA
O9ILaD9sD4EG0IsuOTJW4+YiuHXQcb413wPZduKIwLXzLyZJZBGd2rKfyAzV
R5+Msm3ifK7kt/LLCnh7DUd4Xw+CjDkwVvzyBlbblNVWS3ejBPasy3kkRJJc
ClmOoMIDNeJOf0lRvCvzhKX+zSXRLO5uNtHsYasSxqBtSkeCRBtQP1EQ4OCA
uJ6qZzitqXN9T7GHP1/lxGl+D0EGLLkdIOykgdZjw/NAldJXBsQIBKpDZd0H
BbIvEURjnXi4VMmJ+6SmvfVaMRN+JeBmUpBH5iAe6kWbxInKj9WMVFDwwr1n
Mgpdckq4TH1i4XqRZl8oge/AbnZ7pjUpWb+O/993xtfPSRVqRQnhQSozWI/a
3c5z+pyJo2PJW+tJLC8mT8x0zS6yYMS9ZSlY3pN7D0mUlTKMxKhWJUngmtLj
JMr6jXU6mwBOHSysMeV6e0me1ISUbhzz9Y2lpS8/gZa43YsJk2OXF2429twI
A+NPZ6y6r9k4/9N98FpHxYr2FSuEzLNTjOYdAH+Lr4A9tNPP/czVG1bxy7Gp
trLFxE5ltxgACZyB5ggoqWNwOClMCaQeXDIVrlx0x9X8tDd+aMsHsDRmG1Vc
TCoOqI0RBnEzNPiUG/MLiVtUT3Yhq/wmNxfG7jsGBsmF7126EhHtUm8n52ap
1+9RloC+CJAK7ecsCTyg9FphATEb848bl2P39/uFeqHQK4DTtr9BOGvwV1Rs
8cMUdd2W50V4xD9pYs9nJ5fJYfcrabeqBzeLssO6G5Huebs6k+U0TVcl7+jr
GLWCiN5a+/q1bAAEVi1xzm3IwTAtfnq4zGrjGGv+Avn8hdm7UV1EKwIIquxj
XK+g6y0CNa0YW2cVSstg8+gBCIgrjrek47pYkHITAzsXBaiwFEVKevgU495a
bYvYku5t7KP45NE8oh/WD2lj/HI/IvJgqOxF47p53Kghh97fFaF+HYUBYVdP
8W8pzQxWvk2UapS3LAeFdQ9V7rJY+j1svQwoJXqNmXfBaBUScAuEKyUImVt3
01MtOVjV0NtWc0CPuyvVFQguolYlH51gA5F7vzQ11i67w8O6mCy6hdkppjjs
6K8U+RHS63SVKZOx807XPsfmsdSXq6X6IHP7OxvE7Yhj7Tk7JuhUniM1bWgL
7ETdvKoc9Sfth8t45CgY5NOqErW4U0KJp6sKyFo/LAsOidas7NKSGuM8glqv
Z2YsTcv9NFbtiEQJRg/LbYK8iuKJYA2bzMrKsNg0F9x/pDguXdGe1RjXoLFV
kk+HXA1Hx3Ghw6Qw9HtD7oRkA5FTGnyAdEQkJyDv1JIGJImjigHbGvOpw/xv
jZmmp2RJWPixcx+oJIi3MFDSu+hIO5w4mOoENzZaowLF8YpLqb4IktPPMTag
B6R+6KAJSISdCVlWB2K0pKFpPfPhgocBLcSTlz/FKwyoZAiyFekwwPokSmL7
kmKcLJBvn/Gbs44zwplfvCwBQvQB3INiB0ZIMe94rWMHnBCAXkYnExtE04b0
3ToKcv7qhSDaJsUhL00/dppd3v6nKMZbIbhSuKutCCj2S5aW9S51cHAMwyyq
CoMnWKrQB2lyu2KAJUzP2kx2upMiJHa8E/n+HS+ocx3mRjGRATRXm4NprVtI
T36SbDkvb5qvcXiAAvbAkpOhBwvTGTDRGKFFgBv1hGKquXdS6G41LXF8Vj/k
dRWcPSFNzjSKu5RaKMfX6w6HAkloLn3/vg5GgiexlmJlGqs0vpwyAWBGBKvB
r2tuckS+Z/2T7KnsM+m42ULNT15WPo5OGhvZGG96Os2QEf8B2SiL/zZYLVVq
HICcI5nGzmGhLN1jwwLpyFwjI/QNhLta1bLyMaf+EWFZEVqEf9sQv8dvWdnH
61Bjy/luX31mKVFc7cqUEmPQS1q3uzGVEs519l8Q8LQSzEyB+JwXRWlHPukR
7hjJZx4xMAXVrH+zJv896+OsM435hTUQlvuWEvBc7sd4xxYuHEZAYhpW38EM
ZUMHaSwhe/A0isnAPu4xNpL8Cg29x1G6ehUE5X9qyjVFgnbTWCZPDiwEqLUO
RSKBMC6EtmIS4nN3c1e1Q+Qu7XUxOfhcuJAXEMf5S/wpta8De9kcmGQvljGH
1G6NCFEmPGhWegFo1F47YpMcq3ie20Wz9wzMDPhhiEfkYxY8+NBJKh37EvM6
yDe63zuGvwVjqc9aLoK3HeVGUrVkNxJdbJajSnjF13fKurfLov3sx9wYVyxP
5on9+CcCP/fNG1J4mZkkoWUv3p6aivc2jij1VSssO7xWHEgn1a6sQ2+IBXEf
X+RGoxYsncJuuWak27iDANNulcxiZTeBwEY7aXvI+Onk+0IgQ5rhv9KTQkPb
4xXEYjj7MjUEfY+J4rpMdFqj00MjxxF280MQi8bVJ0m0NmSTWMEvLbkrQekS
3OD1afWE3xDWFpfSrRdg/dgy1RsarfQ2hXlkEYte7Z4UjdKZ/f06UoXpscoo
McZ4Fd+hxKjjfiS/foeIF40eDSgmkwxO+XYsC+U2L6MuvUw3bvHtSLx6SI25
MzC/71llg4p3WtxndpG1SaYz7o7NmA5unLX1X3rMEOlxLWwouakC9Znivd/3
uVHOzIFz4zQKcifR0YBFjXqCQMg9qA5OwBny7EK9wOoeeXZaM9KPU3+Jtku/
aEiDE07u2b4VFl322VyJyIvvacePAm5KgCLHlgo8jCXdsQMDWYdfQPtElGLA
C8cIDwrtdeU8Da1ewwK6NfYGdrDwi4X8bIFovRsfRTq/IxJoLw1Da2nijNnk
AzVq2tb3tVS2gzV5mPRir9KTm7mOeHzY3ZFADLRO5p8AXiAhHzLr7YXz583N
5s0YLtcc0wPKs9M2ddifGN5Pkj2OxjYkdopxWOxD2pOgV8lCMMqKXxXiSIdq
Cf6XtDWwtSWIzNpxIws+qDKbswEyHJxcQE5jQ68wDiCT5h2durzK8/ANk4Qk
Vfkjv7XVnbsW8ZmPWUX7+lc2mF7HOfmPumSy3A62RPPUvxFe/BfL/h18Vo6g
mMCdUXoLRz5Z30tQrfFQjvmZy8SldGNzy4iYWp50P8R9jYNPnuXX02i2L+l4
cTt6IcE1n5qYCbHgvJrJPVvrV085MzU25XxndMUcvUIfhjAlGJepf95PArXK
S0H8H+la/n0DzOr6Z5qYdEtjwFn3AHXLxy29wuadFZHv8KCI920Qk9lKwvzO
iy4RaDdyAAzz18ptsR1BwZb46ybEIxESzwdcPMqerMHDQOxM/Pi7Yg8biCga
XCT6Tye9FTJGA5zb6+xMePQVcGyZJMg1fJ0Zc5HguXeksITUhdZjUs27TURe
9xKL1p5ewyn2wZC9zJL9js2zjTitabMlKUdfTrOA3RBrhkqdddymRXmfdGDP
mdnMswT6mL8+nPnN92Zm6DZ2h8K5B28HlI5DaMA/97AoiFVX1HDdJDNlzOOx
67UstVEZJ4lZvarviqA/zo6qEoZihidKvWFxqQNaVN1opc0Tqxf3r9SeRg+d
m+q6be+BSnQlMDVwy7IiG3qnCMu+fQxBLK5kke2NuqZ73sAJK0vAbuIW5Jyx
ajZIYXlqHgw5AZRHHGpgHSDm6s2yDJTnYxF0r+orwzt3b8Bpm6qUZyhB5YpO
qSVWpBiqAct2kreaSE2ufkIC1K/wWS7gbDx3FbKW+F1hScRncuc0ZdhD4v9f
iE5VZ+ggoq+E9mjELTSo7gkRkaFnVQGF9EvdS8vS1h/mXqqVDnKi4hSSoONl
jfFrHYhPoter9dSPegCLLdKuJmnmQa7LOGetLIO8kUfB1xcOcFJcDknQ7Cty
dq4sV+qQfQ8S+BYoN+lnxBrHLivCo5qDGuYa+0UN/DHp7wsdTlQgy2ji8zKR
+PVlatOYhRsI/l4ANeV5+hE2SXLAj/scyUjTttaCBGSCOuDdJZJWws0qLAih
k1FkK4LkVN73n/xjVl4kF0uU80LOTOl3KfhGUJnoglaNumTvEBe/pMvncC1K
71/bgicQYwNQkIAxO1QtikZwhdjIXZRlcJcddEhse9qhMBg0wQmuS4o1DELP
ru7HH21azJx7jBsfm7J4EQ8bTK0VB+UvbEFpf+mNAYBnytQHDtwM6V4jo/nz
QQYmJGpkc2w7EEAl2Svqab7dUJ4YXpET2SkAXdCWZQzFKI0y9WGlJgTE5c29
dRna9CG/EgMoE5srZis4dmIHDfO6JwXJznebMAlDTEcEP9yqWYcFOiBf5UPe
qSZV6yhNkBN7OD8+X/id2NjOps20iQJHEm6D3Z0Prrt4GySD1NNgkVo549p3
nTtKsRV3u7rIoF82+KcHnc3dflYYqspb24DcX1v7AvvKlzRawiQIDN6E1O/h
gqZTk1Mh1e2iZXYyXlzuqplWFXZqFg1KfoK25IvI81NJLMu1LGxEzjCtcFCn
JUovE5smvtXu7U3DzCmQ3ypdhfLcdJ4D5uTjjHG5621pbjfrUWe+1ehgRRbw
eW5ii4qj78vOzXjmaZ93or/PDi2rTX8sDNz54VM46pchL/uvgXBaPLK1sI7J
VerssCv/O30SpiRGd6A46nSGRUAlF4x1VD4ATLF+YSHfcrdfs7crlY53X5l+
EzW7auyV+E+c5WjQHhhTGFXHxincShWoJsY7m8TZJ5RrMADxL4qSkAr9Ayuc
SbBdaGhIyfdmzxKwsPY7mTO+wQiz0mDV2X0nS/RO6zsphObjuKoHeSlt5cFK
NrkzWMX82PpsTGNNTsBhffQk4eSz/cSDIhsvKCbXLIsZ8XN58AEyARC/O8lU
VLq6uwsdO405Ayr5S8TzVBxYkyV80NWgYWT4LR5ygk87Jew9qotzLWIZaVYy
ePaaZmUuaN4v7HmhuszksCm/qchTWTpui0V/kEfD0GkcJKbEs5H0m2DVylJP
3ab3G0mDflsYO612YXO/ynEKxBKfp8+/6JaY2sk/IfSeO6qDl4UrYY0xg07n
9V6iWGzhH3AGGHtSZ0EncI4S+mhtNle236Qx0YnNHyqlB2i+/Opi6D9dCIRW
qaFuifqImKW79FAPAHxMY3RZVj3zEJYlOlE84O/DzRzutkD+WSA8ZFKK9vfq
dEJ++eMJqcd+Gdv9OIuQmojRJXN7eeU0apsnto5zHkOn8mcBIbsO3oBenTZ9
qKx1x2ZuUEm6uqNrQVV12NO9agpirbTov0d2wV44jc10bG8sX6dr0XviYiN/
kbYJbSwLjHxNTD2TspsMNPYntEN4hfGAKzqpSeDSqUPtvBDo+7Q87CB20P73
NgOaZ4KzvJFnA+NBID5hDUSfBFt2wHonm7vgaRJHkKKL21XweFpQ0UfmO4x2
84sqQ1/s030bmtL2AH5Cim4wmEHIruhCwFVOkYbYFpInIbUeztTB6tWn5I8m
7il4H1YHTo4PALctaV9SKwUkfKlgw0NJFnsif1aFU+VFbdrA1Nzbt1zM2aII
RpfgfWW7TwgSneexar6xw4a6DnwZ2HclxVTCm0u9qNK6VCau8hGHkmc7wJcp
z1L1GywwoLRd7i0KSVwAgVIBVyZcQMpCC41e1xTv2EpjJ8LwdEW/z5fmt/zV
lMS0eamA61ouDnPVzVv6SC6f7j63wLOCAVhFsNxRJYFgvirjufewfobOdW0N
FK7cEQzh6Nf9Me5RLTs/ErI8D+jo7Dq4KV4EiVPy44hHbyRBoWKyertFDlsP
HSuX8+uSTM4W8AGo5veK5uoGW7064UashiDBuepYV/7M6navNTEQKE06fMzq
1YoFez50mHj4eG4NxrHaEtScEaX3PoUn61A9Fq2zMXpD0Pao1F4mxeY2tqJm
2Bi/EH6PYj+8y8jtKve+fytzbDZ2p2id1T5a20agxtKec1bK30lhxCBvTiaH
U/KgGgbFfHIZZGJeeRgyHtYLh5J0uWkDOPwGevI74MwDmk003ib5jdqZMIt4
NSNUU1EOKn0Wfuy3sZ0vpky0d09AsdaSUryR+F/GMK25Hd9DTdUTgrybcKr6
e78t/4pz/0PUV0+bsLACkQn4iHfjz6WkFg0qSRqwe0bXyFFhsTlTqKZ873XK
ZLCRucWD4HsFLiokis+gb9/nvbD/IIMLwCcVQe7h0Zv4IS+P3b8mvRA8nT6X
Eget0PyueSX1LJKABLXBCT6MO51DdFGuAflmUYqXAuJ78RbzafK050CQxUt7
MK5OS2E9ZcgJZNpP+JkXRyhAl3tvNPi720+GRrEcJHouHXyuVJHaq5RRcyD7
deTTQzF5E6XToOfFgyVdm7tRMHJJ4Wf16ai6LyxdBX47kcQTcj4nB5wx0i+i
UcjtKA2RTuqn3jZUPb/Lqr+3FH81P2Q0gpCiWEk0xbEOqTwkSt+0B/pL3fXr
KXGTaDp+V664T0aK8EhRz5sfgzDNdzxUoSB46l2S5M203yi5k8PTsKSS6ugi
rfyuu4wrr0jOOu/pyvhtcIj8fhm0rSAIdeD8dPYVHvC/6hwz8XEo8MEyOKpg
+5DvkGz5V6ecMnqL/kwM/5fwtCInASuOo5Xz3/DpLcru6nBt4KzPc63FYobH
r6eNXEs4bJLC1gPCSaj/5dmD0ICHjRMk3c68Q9pxw9SJnWwN1BAxP8t8rdNt
CFrNnk1tpXDIFlPG48DKebSTi0L+DsYqD/KueZ9rhWvyVO4IMlPuCUURIYmf
+NyTuqKN/+zuKTMwQDBwdc/880VTVvFz3Oj4MPC6av7g6RxKX04S/uRceZeB
KdmxOWOZ9cZ9q5yHC5Y4LCifO/NM7WNz9ayd5Jq1D8HWS6gHuZhZObbPZsfo
w3hcKhDaNjNvB4JNKau7I7smeh3abKUU9R7TI9Q+0XLs1PUjtd4uAHUc2oAi
TZGD2AszybF/csbB6IXqy+LjZnBVtcr0FX/jE17BALAVfiWZuV/UxJxcuPa6
IE/hB0HeAlnhZp9kFzB9JL40gjCAtvu0ETqIKAWE+X/RJfbLUlPH6TJeFLyY
+cXXWu1nKNSMSsIlqfF+w21gdkYFJxqBgcvbaOE1yvxu8q2cLCC04mTVORtC
fh01+fgd4qv2vCYTlMhozxCNWOHwEZMkFGDCmWAYvSmMFnAKgUplVrBJTBTz
gf954MBp1d51j9nIsusVBFYbzcIG2X9uPZAQTHfDfWg2i31cxbGZ+v8T3Zm7
Dtp+4iyhK62UCwsQSDEgvcz4ofIIBFOoBoqAZS4PTPsbG7VZCKOb9Qrpwjul
hdEL57A9EFIwDInlJpFD0fZuS/6HxWZzrtoHpUbSVngD7TV7Ah0ucgz4SUkn
/ulFhWOow8QvakF8aJTCpJtd7+3LTc8PwQauQu0TpNDdBDrA4AW3inSL6Vy1
ZKX54BQaSKQl5I0D5325f3xSD+q93LwXDLU5DIWMxhGWRLHTNGArDWdySsj8
1icbF6OhC4mzjMhGeflvZR1s+7E6oDGdVYpE7BGrDrviS9HL+E77icC1s0Vj
GxNu3lI11eXI1t8VEcUdF8TNNI0HV+uhJFvwHL8nsbFLxGhYpNGX2lt3xatY
BIP+EmR8zOgEiO3+4MlGaXkgcryGgIIORLiZdRRZyD4Fky6hQIh1klGKJiCw
7fJtuamzdwtuTxc/Bu1eRwL/eV5eRPrnPrDIFYEOIe48jOLBE640MLlFSsqT
nnXrgf82R7DKERWykcOgb8CgWJgIa0bzCmigVspaHD6Vqu76nhVE4oAMQiio
oNBY/xIz9BnqG4EuutgHI2yZ6fIYosNM+nI7sacKpiL1yIdeRC2tlz2kS7pe
GyZSDG1IxHNzFF/v7xHbBhI45F+wjOGawIYnNvEvdmTKz4qP6m41C7Qut1kB
TyVqM6JBUF+HxBIkPKuR0FcAnjmEr4wn1BKr93xxbXOHDy4NVlaqWKrv0RUs
ZqfKVykn07DSAmQOUpN6hbl3tf5W7NxEJr0t2uD3TA4SJwKpmkXxz8G3ELqX
yZ2vddP+LzkubXnCDQwqO+s1wvyMqmKiOwA/TrIHt2VJ94jxDWojvwtdGZfT
EPvMFhRbWdBCZVUqFvnol6qeUNRAQTEfgcTu992X2lkDtMVzZD5LZRM3rY6g
AI1yHO1CzOEQ2KG/+a/iNq5dlcuIUaObPhUYHxuThabkD+x8pXS4liO/AAWb
lCsErFP5N6/cGIgHrjupqZ6WHLXFccry2RabM10HcraZ/Bb4hjpcV031fMND
gvbb/QbIMd4UEhxU00GeSINXvxYnGstjAaQSKLtLltzGfv425s1IQP1QEUCD
aIEyt4xDnvXGUPiIzbDWhvWis7BXJjL8s0z/ZxD+IHDrp/4RnYMMYCeJKir3
vW1Zgp85j4ZSDtiB4REqqvbxBgSsA4sN9aTcoRgY5ta8eLFCyOrYln6krmag
f2ArnT/S7t7XDFM5xK8XbvNoQE6Y+S6a6IKN2G91vU2LVgTC4J80gAsJWrXo
H9vpOg+DFVMCuRNedUWwzSld5fs6elqtg7uRP+hPWJVnqW43BUAFSyy4MQMg
Klj75OVak8ZQfp9KSeV/6jQz42hwz2rM92BZ5BexDwgOcPupplaYcxq+YwiB
GI1rI+s6iWQ/62AQ9wrgzhOufaG4P7CzKx1WWQL+7FkMUIQORyRQVzCKG2za
n257XPjgpuNPmQoeobDy7zxjOFlV6uwSVkLZsiopQtJqksh3sqTEd0J9OAtl
UFNcW9WWsBmETGUEFA+atOSprE6yLSjoUEL2xRyVncoNOY3uQyzTBnOz7Thf
/JMp3ZxosR4fPNAFaUX66e6jb/b4/cX1URG4t3kW/o9gwvMERJqkT11dj2/S
lV52/9+zW+57KmgvDfjWYELusmibNzLT9HCbVBHRcARwDr/VBkS+yxxt66Wy
hznn3OMqxMXiLgCZHQTLTKHlhEq6r3RFXymWk0k0NbcWnzgz+2f15gSX+iEA
JiQMaew+OL4aYURpgCXTylobAYH+6oCV7lTJy7EeRPqjaK3e5CjewKWEytS9
1k1cBb1+P+T0Z6aeBjNkKPE8A34sWLBdcJkOvlL5HPJSFaykTFSxzgy4rg9K
afRrJG9hdnG2m7PyYhFyd/o8llhAAY+8fv0HxkaS/2FbegRIyFdoy71sAwqi
yNAysBwP9hcVXquRKVZrDMLjVf7Nvsne1a8adzpWH4r6I8gh3jOpt8EzyqzA
sgvGNyNiL832hAJVcePW5jWyzdBV2hWcqcKVMCo9g75nNFOnWrktrmOPhx3H
mdzcD9ftjd6zz80CtleSctyifI3m7ET/fEyN9LSyn9I/xocNzxvjMI75Aa5+
slwuNlKI3rRouUXnwUFcUFvAs1Vr06Am+77aUYxXu3lY2onL2em4/sH+hEwD
cFSjlt3Ba5c9yY1tgYmKmHvz555F88gf+0fHLxaQD+8IXGa4YJKU0s8Jq4kL
BfQNABHQ0EFY1qzG1xjYM6u1qAxo6Ob9W0/wFOWWgY5Uv3/bT8v2FChfzJK1
vBIGRElZNOEUIO25URQc21hMFhSfB43uanVFQgh2yZ8ojwWh///ciTPDPuO+
P42NlyMCtSf7DYQYbVnLyEgVtSPDtSAz0sWVh1Teo29/+5Uli3Wme+8DPZKQ
91FaNknXW4s1gYRNa3V5LxHGtWz8RsRRTRS0BuDeEnRuzgxX4gFBsomH/Pcb
ssYsJypeZerdiUamcWtaaaYeiPN8JKQXRnFnNoJGHH1F+onSKZdIZx0/o7qY
GdkrqEiIe8jB7RSvK+VGZOreslkp7nI6RxsE+UUUnQlgKTZThQFtOoJF6F52
fsru0x1QZaqnselKIMb77NqJhoOGGDsr0usNOH6TcZAIuywm4XqLHjeQnSyH
Z36ECEJsP4f+MHB8jpxuITUxYzXrAlDqb2UBFZ5UlXo4wv8MtCdHl8XAAeeh
ARJhl5jTHBzB9NvIBn+mXx52okIylWBEoDfLgusOpuZtd98Ce28Pu2WlxT3m
r8G+16SWhAUH3FyxOO9A3tgrvC9Sl9Pmg7ZY4QdJQDBKFcarZD/LsyNyvMp5
PiatN2TDb5Zl1vJz5UUWlv2XrgWee8uMLYRBnvDoPZyY/cDYaP1f9Urodc5e
bW3FBnXIRPQT4gkz8zYFc0IbYk5Pk8NCt9xVoXebEzMGLxeAOmpmEsSTMcDb
0Pyu5I3e5TPkySijGOMKvQwjK9Ksmri+tsubBH+oT0zyzhiWWWbOqh/me+5i
ic7F2lgwVEi5U1+trYluv1Wa8b0t7pZ186LeubHHEFhUhPzaZT72tlpqdokz
GLGT8jFeqKlEGk8Rp6ejr3MED+BGgWUeTj2ITXqmZFhILrE0r7c2PiiupeyM
NonM3SOyjNFacEuXPkp3qPDuj3G4AXzGTtJ1iHZKMBKhOFWeHh3wto4K6Oaj
T5uPwg3T2clMCSIx9Uk4y3NHqfYgIFOJo+rkKR2av+OGbLD19q0uDGV0i6Ee
rrHCYZcQkx8CZDzrqmxRy1Ou1HxLRM1LsG1oqzXFDCCgojnF/OUQKIYpzIX3
VfQN4Rwolt5/CX3F/4CSRjQC4rkoWJ53drPMv9oQ1AWtTwXtLa8weWQu5TDv
fk4GSdw7SgkjvXZ1V/5mEY+ln89969jP7sGQVHZ49jRirOF0KC2izyBUt6KA
D+FUszanv6uLgPy4LyCMuBGjlUTyzHHzsVX6j1aoDCgLfuE5JfgL+ICyMTOK
7SSI3Ge5Jw/BXfuUQeVvai3tUCQdhBOFrsZ2Sqn5/FtjP6PExVxpqNCg9wnp
5gNiWRKQ4DG9Jc2joUCL+ZRtp3RLtmGKwXEarDL9Wq8DTpapqmvlGqFX2sLA
JBcxLTJxa+NvyFiyejny2b7pI4IMR2i9js3KZCnKVZtSqXHdYlQS44c18wDC
EDYNWTe3a2gxeaub5byMfMr/6FXqmFp2mvetj+UwJ9aBJ9zINCAIoBKZDq0l
v39rxP1dAfVOzn0Zk5O65U9b0EJV1zz2EbGwIZn6HSCIqjeDzo6EtHFAgf4m
usOY8rPl54Twzy9cp0B8lXZxT010Nd/ZWqG44B+J2fu+9LQK7pDid8Ezxpum
0H3X/oDVS0Oz9H1rzn6BQNitEjNx+eG45jl3PCmzJOajLAFKigp9P5RzJtq4
4H64rYPetLJeVwXJgholER/niWyYcyWqP5b2YBJWPiorkt3MuuPAp6nyVzza
UAb5+7TSZf5DCz8a5i+NPJ8JlzHhxLT2FjJCAMr5/Bg29mtUTwe3kla6fRrI
ITVYV0wLKvFtPEIRgLMouhqVRUkzSPCm7GVBXTeEF5WeB9sFELON+9VfVqcQ
oFhkUwJnwAbwZThbrhiGvb8U+FDxKPu5GGGLEOywmH9DXXK+Jbta9lh/2LoV
+39Jn5i7fGb4QyIT50mMjukLJZd4LtfATmCYBGYNHxBakk0PhoLV9VfpEy1f
ZSav3He9ZJfus2TrbKSypj1BbuuOxym8wdvJmush9OY1wdGTvMQHP3LNvNNk
/EjyYIbBHuaISFC3pcZ7Eipe4XTx8wSRPUhorxILxjDdJTl3bmCC4VeXgb+R
OYgfpcfFhSH+OVw00927KXmbWpRvi/VLVifHR1bYos4JjtTDHjDlFTBnBrTE
Z8uINGSncWliQEAAcSEhDXhDHw0tk+TFVyQ02B7SP6kBKj6Z+XTJchvT7Hp4
JKbd9/mJdHTdFJAkeeObyw5veGPbmduRKbidwIOyS+NJb1NGOay1D+FMsZT/
8cwL+q0fZdUQGvbejUvnBHK4Ja1mt7KxwxZ5Rx0mnD36vUx/d6psgjYqL4pe
/ZvsfvCXLxMrQFRk6TmJUH+W4qPOC4HiRsX8mD9fnChOEZewPrOWq38mgeja
ojW/Wvlkyzt33UsThSIzsCYDEAA31zTmLkSYzK5nIZUHeOG2FhyUwARZpR1t
xt4nD5CUSg3MpUN2gXn8m9cOZqn3uAcZWv/WuvcgcT5Y0XXqJ+t0mn7slYxV
OzdNlvBVE7F7ll3tBvYiri/S9JLRR3W+njpza9BBPWVMN6wbW+xoq6HWKkya
SS7Wzvqe8SoCcrZWUkiYInpfoGwEEAsv2y3DafYhDiSa6uvRb5aistuowk6T
QpDZYEF+NC924hm+w5eKrWg2kCM+3al2aPJ3s2ln/QMwNS3Gh9g+Io6o/Igj
DkX5X4R/pERa0Ah2xz7BzSDacQBLi/OFGFeMpDlL3TcoEGYkksmISZ1AJJaI
LSuzCWqeqZKKnKGw6ZGyCwW8pIRi0CKXVSau5aKdnHHNviEKP6qPv7A/UYEQ
htK0MPOZUiWrgEn362LAQV0SuoXbeMz2zyHsBvYlndplwEK20tyF0wikyc1d
7B1MeFL+sY6R2r7qz4KCcggcUxlEJRimDbxqnzM52qS+1SYHzy+5iJiBbRHe
6XMQdSFNxOfv/skelPdBHcnc6uuRmBT/noYGGZqHZwkGEmhl3XsIzOzh/MfE
58IERM5Lqo5v/9ibGiSQyKyduvpWiTO7+qMDaa3WDfkvDKRTrATvV92ymYL+
HL0zuyZEUt2VdIkkwgbbmekBxKs6iy0FkCp6fHg9TKnh+wGWJ1Xb5mFK+VSN
7Eq+mqDGy1bDS+991eGjEPzuDWxSYF+PELfFSedA2x8FNQUOUFSD+Gjlz2xf
WwHmxOuP/SUXt9TPBnN2AucqgbcX6hSOE5l3fS/rP2KG8LeGyeW89PDpzvP8
+X1IkR/yewikcyBK5NhP1Td43tyHPN7QqTYZixkIriemBCfeZuO2r1jsQ3YO
EHuZYlHd0kbxw5FfPgVL2N0kEeKSBYGUPpUwzGNzLZSluePYPusrLBGbtndo
dDgmLIdZf3whZmX1t5VihCmjGzWkwGtbDI/Y0a4FWtgQnnuTPgSKr/+1pd7J
H7UfDG1SGntKFI7J2xc1VHqVg6clzwt2kyYVK9w0W9pjD2NS8quiEoJW0mX7
NgZDpePEIwtR/IQGrIklwaGxk3k8BaksKaFPt0QNbKd0EN8bDpztVxR4ps8f
O4ZPPNxqczQg3gVGgVTG4MHUefJ8WL0RZBGPGr4iUSbcRjIFeZDbUWIbWE1i
QJ2OsadCcpukGMd1LhzhIsZC8P4xpcu9O+MNJbuJ/aZAggABuxf8YMGf4BLg
Z/S4fFC1aVnt6l8/ADzq6xN12i1i9cdXnQB3hEQOn6W4Vd9fO66TqvJKmu29
5m6wLAHJHgDPtFmpZJAPCTp/Godb0V8WwYfJLlHmjEF9+hyZ8QRoG8aAid5D
+OHXltNoLxeTFOfItUZRBeOIckOS3/kzH1yXTy4E1Jy5mPfdsjqSodqWfX30
X4YClRuC5XT5JqNylof6RIghC/7G15ev+PIyl50/En2QNyoWepE9tHnBL0K+
0rTJTSD4QYf3gIginy3iBq4s7pu0emHN4JVuMKH1m/in7pIxK9RlX2+NPV5z
ax84jsznpSEQTtGfDj3byKSMghredmlgAaFl+MwKd9YtPEV5GrcZJXmfN7uv
Ibb8Go2uC1kAXm+DcZz4HfeFj2J39F5Zb88OK8ToWHX2QfbYh03jn6TnMUIO
qgyFbL4h4EM2v0lLoXwuCtC/b2wgiR6FRvqnxZFSbCmWGg81a25V9bTnyecG
QSYnjERjs4jsiafHy5WAx038lQl42CQqEmhdAOeYBuFVjVicPG+XeagFgz81
zOMlwSYNutBBiMCDL5xwB/7HewlAXRSdPo8ec5fw8ROWaufsxqGvHfQ4lJQL
Q2PFAFUE6Pd/pTAlRQOaamugD3ga91LMdsIP7gp/G43gwFVtMkXc+PYCz0yL
nGYvx3ZdBMnKqs/pVBIBHyGK/U1gE89aYaMqJAZN77Gqd85Htx1gwez1VkTJ
Vy850ccURTlW8i/HjjiX/9J5W4MotBioNHDpHQUtvA63YOebGfkzMsbfuA9l
g7Cweab/sxG/d4RsUwsFYw8TG/hc4XPFH5BcfzOiWDHr/qPOuXLYSrwEZm0g
frmk6Z0BBiUgmZoxjGADpx91dBRF43dfObE3M8EdIdcujhu3RP2iJ6uZRz0t
NoQIA3Hy3bqgJjFZ59YO2vomeyfFulWxqhZVHYK8fR8KYL3dyMKPqxq/Zidj
MELLpfCZWuteBOqpDChBI/EnW4ZSqIZBUslIn8CjpP56+7U73TAmpONSGidt
qpP7BdB4QrZEQtTUM8ah4WxY0TwfLHe4/MGznj/E/npW/xzI51IlBPmclp1s
KoI5+3i5POwj4EKyo47HhzIGqQroxMaYGSw1sKAHxn7PE7i3bmNswsAt4DAU
nq6mY8vZhVnK36y0Gieh2H7X0zzxM+BP9OnIH/BspLkKqOmixaiTiAPfJtI3
gQJbqLsQCU/oIZoGrUgmsRiOTwQXUIHgMm0lG7aB2r+1GcC0baR+di90C6x2
OLVx3ELLYAIYsg1P3qks8/Mr06bxwYV3Q0ElA9+zalXwkoUdmmD3fvNCYuh8
+FaCFZJTzly2As/XV8qDG85sMgCl+1iNsMBcqz3evbZOe9PxUZb/0X3gJ0+9
HbqX0rzGiUPkUaa2SiclfM1o8U3jcWbwS8oCkLVKbqqpYQS7PZoMqlBJviFt
soVx8ehv6f1HY6uerCM+MDmRRebhiN55BCUKaMWbPdDDg12zyjArfcMKkbES
CNMQs29IuGKZVTmXy7p+cZkhUxPi/skimR1DMMbJAYCXQ+TWbVXlHIKiJ1IS
tHd4+kgT+dqqT+GuLqAUT3ZWVxmV9A1Ba6EvB2PtYtFg3KdBpkNcNCnnYq0K
tpZnDUB0pGjnu6rcovqtUPVhc+EzVZyEbP+Xc8OjBLlvm32OBn0cHklpP7wg
GXjRmeVPcwYpPrOaXkrtwhH4LWEWCwdXBa0diuLtO9eJiQ7JOE7Hxl5+ru3R
eW4dmFkNM3zDBPZeV03TDo2YX233VZH7g346b2HdDqyQoopz1WcCial6+igf
mgn8YiJxKfA0QBhGdDh0RUi1C4j1tOZBF7LLeHgCCPdmqRqk4rvBACpVmVFO
p3Q7vLvRx7xRzfFpcNAdPA2yNfXisFoJOEkjGUJVdk+ZYBjCD0mLkzRvaddT
YZR8yP1mNlEhaNEjcTXWODHDI674ROTo+SrjCXzzQPRJapBZQC92l3PzJsGi
ECPMMkORcQd6AeHiqMyavqOi4gmmBQ9IEZ9uCv3sypsLPAfq98Ld2ONkrZ4B
DVkhaN9OfclRb2JcSoijLnNzz0e8TkzXXfWg+iRaS8UB82ZNcg4aeg77H3i2
0lHIgZFaJMVX0vtbIkXwbLDncmQQqUJHf68FsNUw8boZyvrwyD+XN3AeM06/
Koz/0/ZtlNBrqQWOIx4yQRw5X6hkN9q6yQQ9fhnAvwcRGqR3J7fOvFFDTzFY
EjFS7aZrfmS0MLTdkupjpLYl1kFBFrnb7XCbsgk+iTPpWUN7kkUrr0R72k9H
tFhFCQEOUg28h+BT5/Eo6jZLJ39/u9fAwz3obcLv3pydmFrPYILvXzx4S9e2
si6YFtalBDgjTx20PiWWSPKA9YJK+PGGmMigE7y6GZCirbIP6A8guUVjW2MW
vfOr6wXXlVwn4GlkvzPeoAIDeGJN1UncRIkvFysLQhgtvKWO6HtV9mmSsafi
37/yJ6wZ6IxkJM2AlT+Ck1RJr3fRPGNvwRSLy/hMXX8HBySgmJ47XVi5RNyk
CVpho8VuayW4X5hBcKIIT196LZENWGReKSP3upCJfQxXYQXBG4t4+vnrXrZB
M6+4ldjTx2oA1tyJRUCOq4XZa6NEBpm7+Sd0jxXHU1PIEqhG0bUKT3zeV7Ua
f/z3gi5Uj5YQIpNeNvXai6N+FqUcSGJVrczGxu3+JOvBe/OYfCHSwUc9IMmG
t2/IT+K3zna+lJkQusCgluUKduVa5o9xtC08SAVB345HkGPsrgbdCQK3QU4R
tNrMFeVtQc/AHXDAWUtmGUQpV0pQfctYdkvFBaU76f0yP0biHDkrhN7ZnXmt
riY03sid3Zxns13+rDbADm3wongaQ0h7IdON94O+k5aqhbs4MOyqcAY92w10
toO/euSh3gmZD+spmsIpRpQYeG/JsYEfTd5LNiRZeM2Tlq06wUV92JkQMnMh
Wa/KPl8L4LxgN2OuMHWEIwb298OIIk38QB/dQCt8ws0oqAAqwZuQom7TohPO
2JLn0w7IgNnreo5OkYBv7EyULZT/hv1ArpXgO/mjhP5c83H+M78KNiVYjrUj
DQiZu1cdRLDL5R9p4lObA1ULQ7XKiGMlbS0jcIiqlzdq5+Kdmm3HZzWKdokI
upIhsL35gXgSKqZziGxnkw6WwxQsY9nOTTG/yE3umSpobSOZXYKUmL2A9+OT
kBEklCLhRjBdv8b1zPRVhxIKcUBIcc1nB1qwlph7ITs+wHuVmKQEJClU9afU
IP75GpCCiCybATkA+3XLezeoAwSjqRjJ3ULVPhQMgzUKq9l0f14vI8Jc1s7g
NIAGTbT5eu7d1FVXxQRwVhuuV0ASBwtnFLmTPNH29t2vQQq8WDBPfjv4Fr5j
qDuSl/b9IVsQlC7JkOLpdH7ZrWep2fnW7lKO0Ux9tYbyIJsc8JW4OyPMpZNo
2oaiyM3zbTiEuHymnEJ+Z1uV7p26rQ/BI9Du+a6bBg2noEvCtJnphHnp/822
tz1PUOXbRfaBP12/Qy7NEFvW53JEBWS/OcqcJx14eIlIRW5t+txIHPbE+OGb
STzS2PKi2ylkHFdKkMDnjfKQqSX/fmxCT9CqZz30As5YK41kj1PLjrMA//a7
9vlns3uMWPugZyUGYH8GHuDcPS4NQQz37ya+DAtAVZjTW+s7yUBho891LpBA
S8o7pDGwAsTLjTAtXupD2aTqRaX64b+v86CgseTN9KCrL4Eo9IKp47IX7hdP
d/TYPZ/5VqgLSkRb8HUgMiA7NM1uQLUhzapI12wUpqAjASzhyIt2qVOF96iu
Mb9vQHrg1zSUqnxGKtqF59ZXcGDUEmc+DUdWhQ2q65yH7bydIhpIBoNxOY7i
1r+L5LLg/ojAfsyVV/UKabF/FbkVA7mWHlfMdSn0bSJVunJo3XwWozFlWyxN
cJ99KZ7d9ZM2zJhCPjNoK+9FFBGJ9GR/f0Ra0FaY9sUbisL3lc68aCgX76sf
0vL+TbBlazqDbcObnt+/8m7dwyz4O044apEAb7ftwp0JcJFBwv9FU/tFm47C
NabtLKTKPZTnkbnhNq0mk2s1mwgu1I7jh1JnY64XD6ACYpdUBbjijRZaBIv+
wjNElokXSgh4c0G8PYLmaCwyBN2YQvVZTEG6UF2fn/b8QBDPcLEPxw8tVdLO
RWDqmDIOuqnlpQrtIMhDi7qy6Di22crs8X9eOiZunczR+moCDrv6JbbSCK5B
M4mg4t9zj5BqaWvD6kYMFg0rig77loffX83aIcLombm7lNq7qMOHn68MBgkk
/JgLIVrmIcw9OF7Dd638wXDNRxs/QxEViMZnCtZxBFDQ+EWolDTyWESl6SAm
qtuiXyIZp1+q/DvNTrwB+Hfhm1XVSIC6Eu4AEpLod2Lkvz6C3Jr2XWYYvbvQ
VS+sQc/LAuu6PRRvwR0HFBL/Cr5BBaZ0DC3cuIs3e8s/KNYnNO6Dm7EVdTDv
FJ9bmoCANPZ49tKld9uFHwaa2JCRt1LFy7seOibJjn1C3TBiaq3z79my/K+A
kUUTtzJdAonAbPT33vmCZ56+wA6Ie4NnTW70a6LK7nLm3u1MdIuU4LHi2bzi
UxpnXbeyYKxBrJRj9LsM9JkWrF2kDYyRamEp0jWDI7w37ea4iwxOkBtgQF0C
mwjY7p1kzaVwwdZIeDMe5M5jCR03o/vNBKWSNJ2BhO25Q/DMlEv/pKSknyqX
+xG3hhH7NQcFhfWSYr+oN6Yytap41PYr7tGo52cBYTw/+Fz1i70ehLbyL1Mp
2R37TxoYT5PHGYnHPSIHq6tqmjavNZsbhFOhvgTyOfcfEeREC9mhZ9RfOvNG
qt9GX5O55u26SbFsi4W4oEBJ6qP7c71sv9AhG2dVo79SLGB0yuzBmjGXEZM6
ZQBDXptn6vlBbBDpY/xw0QcDmmLRYjap/NW1KBR2fcrGFleW2CEeSj1JbSy7
5et7PnY7ImTz8Z3rioRLYFS74OM7Ih4mV93QNVLsg/Tubys8SEs0Gn3AzMn7
TcV56cc8xexVczxl3naW8R5/AblGCYwtfR5oGn9A4UJteRlWIUAkDRgBKJGm
kl59fk1lJu+iyoxOj2XTmnj2S2Jso9QHXjA9XLfvzTd9rj+vbSmOHwYQdzec
s2zjSVwK3SCpq0gKP/k3zZ16cSuyN4Bh5jNfSkIA4YThe77fMCoog+ZiTGEN
txdED5PG3+SDIg2EiamUr49PNMQbke3BsDEVTTO4EmUuP0nc3Xz7kkBw5xbm
6DSiyno3Rl06rNa0nJPzal/wEJ2+ds8pp4e6hcsFPOPZB4zD/WmXMN9bcIxo
ZTb7BEZF0Y3uMdAwrXc9ZAFS54nFoIgYoRMSEpIrqsPxpBuTe0GPMrX99Xzq
+qLjiEQI7OIYvnPVhEkhZo5G6+bnYZ8LeCgz6gq+qCmZT6x1l8I6ITukyEfL
Fo4fiU1V9Ru4JRMZeWOKF2OBF5UyjQcq+Mr03lyzgVAoueuEn+yzEXnYuE6D
i8ZP3dhpwbZEEdEBpagl0MOJiXWaPfsN7QyayyUT/fnShVWdPoTfmIHqTGph
VV+cjCC6PcXDbOtmC23F7t8LI3D/3klsdK061qoiDPXxA5aqx2/fGI4OKMjN
KCD94jH9GDA/kIfc5VrpBuYzX6SPxhZuZSEYjq6/0byhxbSFyVOw7OkKxOZl
1YgQC7HeiWAEiIe+hLZvD6QFVPucA5IYroZygWHD7PRfUeOyIjl0UJD1N6bo
044HKKQa54852GmszMrg1qYWS65uK/bH6fYvf9EzSnQEkU6QEzTbnrW1he/C
phOaQMesV1RAboW8LoVU8/J5wIM3iKD2lWn85I1sU66ApAtDjhTFZJiEdSh6
48VeyHy2mJoPqd/fTooG8osluzw+p0AaYlHSRFoAvMdep8p5lM85tMmkQSXC
Z7ls8/8onhj1wNXu0YSBMGSjKUiROZpfzhcRry4kbmsEfOaK1+ILYW1khztr
1Uwxf6d8EgpYv4q2TCW3H/ZOaML8SN/xKJnG+fm3ku+bnbSQdEl5xSPe0kR9
AoMQNpcNIv0TiL7ZcmpKS1baG8YqnV2RXQMqcVSVOVWbIZ2iXYAT3lfpE9Wm
Fjl2547tLrMcnVsx1bn2GyfLq70ypbNp9h6hhfOXfXyb0yonpIArWaPjrbqT
8EBJD+w5Y9BAgfb6dVj6DD+MPTWbwRgtdR8TRu4oEhC0pqI3SSsSUNjOULPI
/Kz3YW1xYtQLYlcQirS/xHbXZBxTuvc7pdTKrcyzx9b2b0SRhtI3KepdOxin
DG1IKDuYdGIju/3ttHh94lsZDKBICGUNrt87W+nipq/eD7fpb5QOMhf72NDI
Ixzds97+Vz6gaix73ul/dIsN01CkmaPl2vPLQGT81WozQuUKNPfPE7eeVB6C
2R+JFpFRmwZtwdmAql+GpWxeMngArV1jtVsvi2H7sSvWaYfyfjjaeLRQ/bxx
8C3bbwblx6JdFZjndcA9ny7IGtiZAOJZog4TBgXmANnzYoLKPNCuVf2uNVhy
meenNfdua7neyTn0u3GWiq2OxV7ZFk5lCouDlgcXO+GEidkPm+i4qTYBJY7J
1AkF9Ee9mv1fOLM2/xtSjeO3vnlKyyBUEZx6I5DQr60T5nT6k9HFVyVFJWpP
2ENnR6+8jK0TRrEzB+K2hyG+pTk4fFxYVs+jdoSB/sC9gDQfiB8Ze3pQo8bV
0PfGIsuzF68R/UBYthdY8dI0NYlnnHed8jf8F8cPsV3xkNNHEtClDHqdJKsp
aTUwMdl5oCZoz3oTkXK+y6GUyOZS7OkwkTOznUaE1IWUuuPTzJs/1/THFV/t
XABqKk+YmcHqL5lCtuzxDR7rgqxYLXFjQECi0xIBIER9Kd/4ViO/T/oNneYC
QcsKdqbNiRqoaxhYrCz53OEHAuWa/E/ZFgxb/p2hbG727RSeosC0bZK0HU9/
EgiiQFb4F1rJpd+SeHcMtNYMzYQp2YQGDPMQR7AOgJL0YpcK5bq/xr5s1jC3
UNQHjd6w1NkDufBaGhV1n4Epn5//L2tEUMbv7r62MhzsIHe06NCICqsZ6dWE
iGtDaS20dwElimcBYTUyUVLAwpZDBetMlWlrdAZ1zKc7Q3RNLqUbnCGUDZw6
mza7H1P/v0YtpCZPKx2L4fWYtViZn45Qp1gH+yjeLc71FI8UXI+eGZYhZzlb
/tneLW9Nb4okGjTTSCqnMmqcYbu2XUgXboZEW2gh1Cl6L5VbVMblqn15Jlm8
9G8ONH3vicKAfz8TCeyiF6cBBoOgmPK4RGI7g7GkffJ9I70M8wJG/IQSzFPW
6OqcKtqnQop3ORNRH1ahRU1+7HFX3E0nCoS2a2AI/kGhgUITRzwPQgAOJi77
iAK0fOuQethjCl7GLIoLO5rZzncHjOJqjzTvQztSe9jEQFD+0dgpzXnvnkzW
jpRt8lRNSuT0fMBYLuAKeEwPBAN1rwojzvo9ngpCdUzqQIsfhQnWBw1d8o5E
ARuA+CJEUTpYdHRfopAofRj4HCZluU7Bfq27IrvpdcaxAgI20cE7KW5l+Xzm
cYFVrtSpXbwQzSukJWWoFOk2FJRcdyi5BC1q4kqQEIeD/bLqSx8v/JYHikEX
rRW5dZKz4WOO1rdLoJE8QxtYDUh0qLoLSQAKKTStMW+hiNfIg0pplC2/tVb1
6H4MPbHDZDWA8mgw1XFyQX13Fjtm5UOFSrIRa1voM/nkB2EkkW2H1wiiKb5u
rGr7LSnWeMlKp8JKiO8c/uvysVvhpMW8Glj+r3MsPimdNYxeAGDKE68QluQC
o3FGm/i3rGnJkaV1K9wvGa27Ys4/IN/Jmf6egST+NTcsb1HkQQ+llmtLsifI
oqaCT572MGg4FmPR0urUU1jyDfDRW9tkbUHTXK8fSHSXZhEC+/yGflY1c8zJ
o+eTaDgg01JrGUMBzrumLQ2rOhYTJDeWadbEPH5MvBAlZ8n//Z2NWMLvRXlI
LyHgNR8fOuvXHBbykm+A8Xoou6TWHikF24+PyHcdDlZ9K3+Y/0iGE4sa55Q2
+xU0FKo/Xu2iHnryQ+c9RloptXbFMMrkgV4vEBcuCXE5KV2gd+2Ti1bdPKN1
iI5D5I3tXjdwXR8H8NC7Q9ooNldrZ4arUVWu9Leim+z9LoyfvltIluU7TQI4
/dQFxpLap+AcY6WamHt6h2IKcG+73xkZcVqJNtgdoKUQYWmOJ3FFiX+whLNV
8xojcbcCyXsNb2xiYBXUT8iIHIjGNfPXlXoywgAktkhALN+LQ8nZOJyz4LVQ
h9I20nFVFil6pGNpDKs6YoL3l7oE2P+DImMqYUxx/XRocETommP5t2dRvQr7
MmOi7ibBUDwypIehTdQdPH/SKHnTUofz9xsCUwbzB94bRz7ywFeAd/qvFM6X
HDf/0RjI4xJxYf6D/ElS3BAuE3ijfrAqVk4OWqA4B4G+WVxoFfSBkftKS4bU
khIzyQA1GVhsFz2JhSr6liX7VbFKSn8ki3/m9RZwrjrzbZsArUTbSKmZ/OgZ
OePCMDmtYPpNGuQMX4PDk0v2sk1sduYJ6BpqrTzzxmk6wj7lanF6WPLb6DPy
4yqSAXE+ubOipIkguMr/BjopcHgKCsnUqvXcSJnJxRUnWMM8n1IW40JNNhHg
hCd3LGmUXz0fwB7/8srblbiS7B5WpbdPGKSXJ7j5PimEulbNB19GuXK1tw33
qNdM/JeytrQm3pWsruDy4Ys0WmgAtFKPXNO+kDavJbhCbeq15LxRedpaIapx
8wW6uBmFwTJMrkywI/EbmqRQHbSe2UV2erJ5GA5zBjwXZadUAqIDbkDTG4TZ
qi0q/p0uqi/8m4tmYB8lIA5LRSTZ8BSOakHQkPKKDogTpdNqmfcrd8iJ9cPu
bSjztt3g8UbgY2SWl3fYiyAkn1eTwW0ILhT74PNe+qdX82n2UnZI4AfJoKyy
ej8T2pAYaTsPYOu66vz/VUKyAqPyHvRWjB5tj9RIvE91J8Nb/esSkFpGY9bS
OFLDeMWQR08TVqhwIGyeCRyc6w7EVsbBAYnNwgShen5rsSJPl8o0WHMk2x+5
j/jWjy9VgxdKqM4accdVw72z6M8wYSaHzSOIw/HS531aFFc1oaJ8mJ9GxrM2
uGcFWeVZLouacu/TxOmjrcgz0//FjsH2EGlxiwfdLe0ZA/uKWBnTA0vJvR1p
ZePPwTRC/md14oelaK09apLpzO98wL2/mpj/kclFJnQ0o6EnZa1D9E6EKvZO
4Y/RBDIcOHNlLyatRP+mSXE7EGg47jzgnhsMcvBplKW+fNMNig3kZ69WmHtn
V/ynRxE/GLQaHs0xe5ibtwzr70tgNNCaBK2scPXguMM0c6I6DT/7Gc6J3B/T
9XEEfTci7rHQrDXCDu2+5fy2za+ho7uvDm1gqTtrJzlXJo0FbYzr/pFDFlHl
nELuSWvoGZcpwVkXzcFT+hhx+neA0tdL638a5uImWbFakJnJJhOdI2dQLNCF
X5C4rF2hI1h29Bt7QcdRCa0PnlxNwUSgqlnd0ZyjQA+d9b2IN8FPVXUnbY1U
0HT6jDR3+2pP4x3Pvarw5yPZFi82Gb+0/S5SCBSWpeF+0HsWnq4ggrzlB7Zc
rfp+kPeVTpjtfZfckNUVkpCD0V3b7+SxnLTzFq7jrKY23Xz2z/ArxUe5m0PI
97XysHVqeA3ERR0t/ZJ5gjT1p/kIaBV17kQmKYDr+ka2bNUh+pSL7jDLVsT7
9LSfCT4B8t6J/LVNgzuFZVDAI0lK74f6TocSSO5mrbr/ha3cFPOb/di0c5kR
uU4zJj4XpbaHz27rt6Qk5RFPu2lv8YJlvYZ2nR1S1vGjNkFxIIstaegUPHCX
kMfBZXRAPxFsLJevgJdTdVPTrlCqlcQxpU5ZTxsvJSle0Z0gSEgp+K2uelQg
gBynk/N2MWkZaLWH41JBNnyCbtbpmfPyWMN3NZeLlJJhFpXfFPG/g5a8uEvd
tOidM53Dln0gahSv0OMX0gDeLluor16dJS8ujUZ25IOGZPbbEAaqqZFwO+4G
7AmJP7JFsPoEU3EdfPZouSaPlv1R7z5x8Sy5MQ7Xk7DrxlDjvpMarErBKUUt
L8+jSdOzvV6dxiwn3rOT7q1ACwySj49hL83E/v7UW4Bo2arcJnyR+F7DIbAc
0utPh2fQo3vX7I4viN5+dEPPvOTwzumkK/H1xsSDI67EB3iZV6lzv0MyvLgV
qhZ6SQYUZDwbP3/saQwxmlLdVXeSlih3UQuWppv2s7HXxHelDzm4wECVn60g
v5qVwUa3eTNjrXs9ruyx/x1Ib5D1muIYopWgWNMkvyYPAVYiph5Dd6Nr1BL3
e7+LMgVYX1xZjWWRsMYvndlCBGh8JBim9HIAasCohrE1EdMZIoKMPWX2E6R6
2fliFj8shskBmirXjXDE4gfExA0psYjO8K78qZr7tcxAzd0hFUeBAdznMLgX
MTyoQO6f3NDS6VJ3cY96juB6uXjacTsxzc8OEroKvLsZELxowsoxZzE+twBz
hnk+GrwPKAI9I28gZ9rNksyFGcRkGvXiPjq7vEzSZP1+ur56OPQ+rjmq4XxA
pQjhGRse9kE+dDTDfpk1IZbI+kQ6JQAP3U/wMFKXIbpiv4CQBrgP5MKrAYtf
pnrQh6kt6yyr3o9XBaa93V/Hdzihjvo6jHYWCaoJg3zjYgBjanBog/r1EI3W
dOcMztjRCPh4H8QYEk9CA63TVVqdpTlh3ZKOonsEmo6/sGo3A8yoYC9aUaoi
46UcZ44DChjNj3/YIlxwo+Tq/lXLjOU7uVwhJiRzy0+a5mWyscxorBEomvT0
Uu0rv+SJQBrUfALkSBXHftKZhS2TRrXryss7YGgFKrC53zqMB2EPyAkfSZCx
IZ5s10piRyWzpyoBdxgwd1Vq7v7+V8EktNamoPlnEFP5OAR1NyyzUxuNxArp
5IKkZv2OjwZwgZrGNWdqONSCS9Ey+KDH+hl49Nd+scnZQRDJOFmZYin7J+8v
td6NolFYzb0jCdBAUvOUjXNFJm3sdB8wDyk9DpjVdC6QFK/FlfSgV06oQbkq
2gPxGlpAj0OoC/5p3YXq/f3GRVPiMTg1utXeI+UU8ukTLEC+UQIStiCZztQ2
2lYjHOyG6EO4CWPfiWKufZk86ldNSdFSNRBER8NFvRnvVuzkAkN4FG/mpl7k
NVm8nLbUdu0jgn4GdizrjKHMWLh6chvXVjoESjzbla9bda2L6gCto3UjizTB
aohb43qvx+keyrdBaHiHFwHbbjBKpKQQvRO/vUuFhT//lbDr97fkBh2VRosM
awNCapVQ4AU+2nIBTgGUD3NAzBdIxspihYSOb6WMwKZ7JH4VFvCZ3EENms8i
lwYBjyaVFd5Xm7lI90EPrtBXoLarlSqXdK0e7B7sXkKebE5bfoBMRKu2IQ0F
lWASg24ct6bIi8qYPxUFPG7JgLhqCKvA96OnzGkCLBy7pqU7qENLmQxlWkJL
9tkvq6J/IQBPeywbVha7C4YCIiULqGl9VR3YaIRbXahTMb6Fo3piotK83avN
he4c5/6tSZoxxZkgxnlTNldYGLOXKdEXSPew+ST822rJWfA1n1tFSqkMjdKq
Bv0NSaiHjCGuD8KUK22Zux+vVOGPEUk0Xj6ajmiG44ovWQ9ATI0sNOCCHbV5
fwZ5Vh8ykHRsFAL4IQrIL7++gPBSm4DS6YZpDfKpSaYjAlLtHqgi3YSzPcQ8
jgwuKLuepjQzKz2TKPqmyuUkqz/UgVPNrHNlVg9YSmudSZAo4pmbXhOrVNXz
sip1AfYOmKwqmmmxrhEZQj045hf6sttLn/RfyV8dTOQk5VcZ+HScZ0Qjbnrw
g2mqhRyj9FnkZ/tAn9j2If6hygWipROZm7LoWstzulWKAjErWvMJqF9j4Ww2
i46fFXVBnucxXaRw5hZyUoSopV/XbUEM+2+dC/UnfyMTTHXoaIItpDvN5uj/
wyL77lt03q0sXqXPR9qtzO4wj/zTcJOHMt4f8ASBLknzYOklEGeHOm/l4g3d
a9xhSGk8OlRiS4EfGPxt3glWn/9pILyKAMDLXDuTQDZEX9mlxe5zVpm8KV6v
ZtBzsOzI5H1SlNgzgmNrGS17kRRCLV/Ta2WuJwvVChHZVSfGywi+qm7dBSWu
EmvLiqd6WfweNHticqcXChnrs6brb6KgtC+FfU1Kz2JV8TsCnGjjHNfza7yW
izpETOJYMZJ7BjHVG3PGaNCpwU/UAjwcbD8co0zxHZgk9ARuCm5mPYlfud6O
tx0ZkkDoc/CMMvcPJA0ILkO0JtJXZiOuUpzBlFKuu+oBVnFzXqubXqao0uxr
BZcniJiSNC5qg9kBz/9Ig3oTWDYCAuHT3KRjwSydFmdSzfQ12ml3Etge6fUT
3olKBeRleimrdPCF/KF8oM7Y0Kv1SVmFW8GkBmvrPRyryIvjTfh9M5RvCUgp
QNjddkOZiQMjRnINiZlZ4XDRyPwyeSGwH+CXi40PHWPwMCuyQcE6DP3K7nP8
6qOBCv5gEwyMa+RavIL7vc0nN4UjXsfg/Sbh4RZj2R1vlSc3E5/ss/wKVv5v
h6lfUvGpuU5NufK3pjpbWj/R3FkcmAOIq4+ZvavTj67Ikj3nFNRTFmfenH+/
2dHfFusLUssy+MOJnTr5L/9o0XEEKk0oemgMpmbMo0UYZx6597AHF+tgNg65
WD3Z4El5K4kH1r4OHP6DvBTVzaTCiB5J6TAzeRCmDXf7HzOAFETC9NOsq2sD
xi3Fm3aL5KwQVksY/dn691aRX3gqfP2DDAZJ7IMEEtGKGTZon03AL0rDSWJz
Aq6WvZxeRt7ar7NTE1RQXcehKEHTZ250Dx9dlODlxKK11tEMiaQpRxo9AIwq
oCAUaK6icJnbRqCnWYoNoVhAvR2MXheFanptN6hfjEgFE1MQ33JbBN/P1tQ7
pPERXrKf6gCwP/2JltKVIPjoL5KQr8huRxaBbh96xWK+Mghryyu1qfpx/1B5
66TWVAAXp0X62Jq8vftnQ5Lj5QLZeZQ97nN9TrSlutfLJYMGjMW3I06Y6kuG
Hp8TFEbHpzYowg3NCO4q9E3y876vH+HQFoKZehmCd/MM/EApfn2Lw3G520V9
s6r4Sfrffru6jacKduP7w4NUaoiWf1ERg6YQRvzZsbjOrQX3AUIcuJOH7rBD
Zpje1/O0+scIbV08FsXupaLhVyHHQWbKEQID2IfQDPAKs1jwM897rUj0fSq/
Cm/2pY0+Ci1ydHYbMUFrnvUJugvJXh747i6E5DaigndQs6Hwtt7LdlogZzIA
5wWEx76qJ3YhoGobwdrwfrffuvgI1PEyRVj5FVuppUJCf+K4cT1Ku8LQI+IK
jia/Z0nqFyo7yrE77+ofG0cYFVFmDDaHjas5/llQR2wfnZmR18l+2HGz/Svx
tCTgF/GjObUrtO2CwbCS9Cgk+VD7jSVuOaEXMT0NU0+9FOlBgEHAdrE3kn19
DmokthMAEmiiozx8+rRTJLz+uWF8hWTjdlws11gQQ3ziPaXS2vcwof/4Um/3
QAlx4AzKbGqDJ405GrzuxHIQmdzCGO1BRF7NjcEvl6TPcpZZ4bL6XlkfDN1G
wUFAy19rtTZ0Y31Hr1rpwvDmGFmA7jFj8bEqLJTv0WG1j5KvMwKyAZ71EGGs
zoN56FUwxuoMxUnYEOtYdbbFEFK4aLCi6+N8ZBUE2fRanGdkVKN9hbpifInX
6yLS/dAgdCexDY+VofxMs5A7A42iYxGXO2eAON4axx3yzy9Yw4c0DMLlrNay
3TAa5b4EEzeJBFmxX+x02AVtpuUp8jkADST29QxSjeryvxEpN9eFqC5OnaCj
Craj+tSto+Ui6MqYanjvq+62unQ+YDvqSskyZ3bw/GsQ8I4ri1Io0TNMBzM+
1wHZgQ1ROFi0Oy769vCE24QezlqyOWE/jsmalWAjkAHuwL5VDw5QLg1Ra2jp
oNHL4+iKoNBiIOf1YNyC2N4it0nw1YLd+pgSHlA01o11g6Swq4+b967l+cOQ
JlOJAhJ9XPjoifcEDHnQ8XDwmr6Zsrfj4IPbadYX3A+PMLV2kn9MxZpyXJaE
RhfJbDj5SBzBav35mIbjSgIKPl8ZjYuNm5f++e3j+bUgN8kUxx9BgxmjJKJe
s50FxIA+y90hqXYCw8MIYG2qyTNELdp9MrDSL24SKD/6OjqzjwhSFMSU6afl
vd2QsOCtBnU3o4y2u/k+ryO39TJeeBQDNy0yEk43jLH6IYTY9DhbE9hLyLK2
jZK6P7o6VBRz64W/GBIuJXs+Ep7TGLfBh9XIjjFWvjbP2topyXWTrZ7RJZcC
qEXGLzX0zgiKKjE0Uf1uww78lYYQJA6Rk4xAf3K58q1IxxR7oqGPPyF5bEav
f9CPuR33xhQioeBKsgC+OBKt3UtIF2IC2SKzHeI8mQHQjLMcSXaTYKB5Bmg6
aO1RxhnXPWmTISIJup4b5T99UHG76/fv7S5rJzu7vMYxb/Y3k0YznUM9KXoM
Dp8+7iMwSUqmUrIUXZE5sTmQoWd6nUfnGDE/tfqhgmivcoW8bcYRQoqfhq0i
NPSGZHAOS1wk3+S2MpN4TLdqAfXXx1L6HztIeXLvRRvTw/wcnQ5D1HKynqKs
x6MSrW5TLwEAmMmLxY1t6Got2KB60/8aHjOGFDiImr2NnQ9NRYwGawMaOzOf
t2Sx77dmTzCh8JBraThSexjLh8ErSEsF6+nK1dqHTjc4qm/74KPlbblFx2wf
HNgPDXPhsftYSzQQiHS83prGvy06lpJc+gCsFKOJ5Hoda0qgdpXzro8NWnwB
Wq1O2cMOaN7B4JSdMUtsiaIdbfcmTXXsXudq1lCKl66FwqDP3Tu3mM5EvQZY
6Th2s98caF3Mv0T1fqCoxgmeYWBJ/irLqaBscZLkjmytRALHoKfmp2C22Cfe
gUULiZCOxpfYKfffQUf3CaSKvdGdvF7m04180uJqOO85Q5hqj2ILMxTtk2Ma
NYlV2tiMLVly3JYcZfFguVr9i1xVc5Bu3aLeuwLxGTrnKRyqHQS5w/yErQ0T
rOTGOi9os4J5VBAmvUyendTG9stDzBm1vOj/qdSno72bct/1G9V5a6kqPiOw
WQQqxveOMsGCYGtpzX0TRPTopoSd3bX1XFAHodRjHZqCeEm97brvfz0DLmou
qK1c4aObAg+96OwZPlMelSCGPS8QaxiczLIOshLIIJ/IgFjJEfbP/csiHnNv
8kjrqqR7v36FqPad068L/PRiXwq77NAbWGzM9y7ciC7KerFlmtdGPJCI+RPU
OVAfz3qtZHhdkpSNrcfx+qiYGPNjoKm0cetAG3APcZwvINhXu1kwjPFg2H92
FEgdLXCyWmX0Kx7TRa+FWtlMvVp9YrBvo7QHJxgGLmTU8xbKnfDlPyJKMJ9m
VhHb3z/MNMcEG2rj7JgkkSeM1/3JbqRHGB/JZtK/FkwwzceOCf869W0jbkFn
HJsG2XFB6tztzr3ejN/chYViaETWRbf43jpWhawtEEGEHT8mNhc1tvanhcRD
bzW5vX7VNDlukUK1jShxIUxIY7+GDLb/AMjVcWQEJRGTrCOx4Fi0WyWuDzaP
7B1OnZ90xHAyY2S+zLYoTZ39OO0H9tx/2X8dbiGTIN0Ry3WRgB0zNhfN4uPZ
4z6SgaqX09LunyTM1nf+O0By7sXIKRRs3OozbiyclLms93P/QQu0jkGMeX2M
JvT6ZMIUy3IkDkJMK9NS0344fIu5ywdqZrHBI/wezKVNCQ/2kVR7ukzfRRgd
MbuUG3sc27wuwEHaKxZc/w7BczGLVHBRiImWCcUuQoKvspJ2FiYx9FCprTf8
S8Fpr7t/jLC4FKQZ/gjFEBUtdUXYFSIiTBuK9tCCaIneem2/PxaIafc5pSyF
7Nv/GKxOPC6MnJh6u/yov/OoFxHGRoN1Hf4W6FOuMLbF0FRxdZP8qy3m/lPX
xx/aP9ZYBCKT6ZiksGuT7TXjb+AD3eUvL9m8NSUBH7Zvwm/PqVoqzMoACc5e
UzSIrJbP4y52HuexK5KHEodRDi0wDwr9Q6YrndOAATyol+V1bG7P4xc3bf6u
iDfVjhG1452rjM861JN/gZcSN5r/Pc/SEsRlSHPTc0qwIkq09ujNgzMCG/f+
oqgBy2z2I0WlSobK9y8EzbiFC7Y/faBWX4nXpjvJdCo3WuVKgr/VRqSQc5sR
4ZwcT0Q4MmgRbPkAy9kKsQhWhQvD4soUUPTHV4I+XJcIiso2HZ1MpXg4TD6O
1AqjQP6UEemR2KfKFaAx5nxemSDwPL9d6872VXmEMVrh3js7/cUYSbBK0/Al
QCzre2dmi0mRoEm5kw/hQVr7LeVR8DgYo00yD6vktB20yiFzHiPuyZEwLQO/
ANbcnnQfkjLaPPRBwNfKc2banqYr9wD1OpJIGEmo2iUntSrMV9zlpAo7Kwo8
ilBzSY8wJSWCDaLMJT4Ty23or8PH1z9YcNk24GQwTgPBXGtRJHX4erawUNRA
87ElNouplmxw3nBXdtO8itej96nDjk43DsT8vj8EfeAKMhHvIVA4xzxvrcQ6
/LYaKffAq+4YxDNUc9OvYWz74e2zuKvCz9GFo0GAezW3GYfgP0SF4FMhTmqc
uN3q2QQijxQRu19/Jkhv8rnlJ77yM8bh2/otbTTAzjaa0oKiN492kExlK27u
jll3FWvtJfPOgew3291q1XWq4i1Btvw2imyNt1Cm6zeOL2F2kmQvGeqeUjCd
vnolA0m4bEhCUnyu+8IoOjXp/DVQRbnDqrqMYc4co+Xc+gGflab2koOdFKQN
w5idGMTo6uyxfOHFJef4Ww1wSLpJgjDg7kY/jNh84b31N5eD1hGVnnyouSMC
PhNZeSGDC9piaFSBbgBMCGkTNVOLbZb3Ugc9r8JNmjNv1QnEiMB7NafheUZ8
YxgxRloUjKtCPcWlu5fFqDXDMJjFPdyBqi9dHcFAR5LzZ/bMWUEgtJc+7grF
nkJFR0WWS6EljEwWCCkF5jSRulCE/fTSScOaGjxKZZAP2zCjhge8xTasfxUn
YzFejN2I+2u4bZivL95QViKDJF7HuwUuycOTO1D9tY7nyDEvy6ctBWHp54Ip
FKKWgUU4JRc60cpv/K4SI6eA30deqEKApztpNg5Pp75FBL6WzZkufhSFINWi
PW3RO8GvmRIer3cXVKx8dVSk/YAznKvGkpJtUp50N0uDeJBL5U1UiI88JLHJ
lI2mUpvTwwMhVeM55KxzybxCwUz9qRSTDQpEi8aJViB8ouxom/Q2ChDPnAPm
X08yR5Vq4FuTRH9LRIjYN7pGTVUsQVOVwhjz65MIbeAwGJObljtApjcjNgXP
5mz2DNPXsQtlqkt9ljBGvuHcFmj/FAUoDCamEcxiOCeKZpMCIH6f6XKUe3Mf
C7XbcChR7c0LK59IweoQYx792dHrSrPlGSOjN/qUxosQox7WlpoTDXbTOhsB
vrkUgS0VSe6jFU2FsS8Sfc3emapj7FQMStsyzuDzcbxrZDQeORqyKv4Ijc70
bcW1mN1ueoza3xr/gvAl767nI9xwn1j2mdlFVrZzDF5iZijkpV/rm0pcxMIM
cWlZAHi0qpRw0CK3I7WygogcrNlEoZiRgVTvhY0i49e49OFBn2N6ZGLQoP/2
j5rTtTo0OIcA+udpf+pUVQr/lcQB8o03QM4ahrEBZvxpG9DSpYpEFHqi8Ig1
/rYdCdQStdl03ce4Zxe0FFj5yzGSgnaxt8sttgs43lF5d2qFVQxbmogezmx1
U8bR7ipkGuBOS3L+BSRi7mbKaIHsIjVc0lbsXglEvKQosZk7NanaluUOqUgL
v56gK9WlULtLQ3DrDWcCuwFQWRaK9G8GcHvVJmmHTfL7QOfbQQkF52Tc5jdO
o7RIuIZyncS1xqomXayWoepX/A79bXZ7YH0Rx9V3iOXOYOTfYM9hz30TBc8N
j71mh+zZlVd3/E+vzpGo+a4GQHI8RBcwUmugch/tsBBsPq/PeO6I3/B1j61C
wtBsm45uV5EYGJ1Bp69TxwnivrR44nbovNNcpir6Uhy80p0KHa2IkFPxPV93
31W0mpb8V9YvZLDIqiXFW7+qlQag789mUjvoWCGfl1t7+Ctb0vrnv4CMPNbN
4gQfjvJk81gKVMdFg0WLWpJpDFGne6SV2ec9LNN2sNg8M3bWdmqXPm2LaTSR
FPD147SjyTM8xfCyf71inH9nUcNVqEKms3/ekNNFH9VwcXoQa3dNG8GPTcC/
Vkql1wIfw+tXVADjGV42Q1gIdpx4pZRQQO4ruhAwcs9SJmPrvgbpW1EpBEIz
89lK0lvu+lI1V36ehyjOHd3tMmgUq2NHhB8OQ75+yyKqQqUJKsH89Szsyk++
0O8udVqER1JFjPrGbRAQk1vICXK9OzPZOIwrl72lRFyhECCgLGQu+dXogSp4
ZIP+vWNCsjEknH0T+8utcLJpanBRWC/2EayXPW7Fe4JUfZeMmcMOmRKX4y5G
F4HwBbJOWG6r2k2wdjFkywgqn5gV6dEydMZ4Zmchlw2edEBYfGZvFx3ZKFVd
IVVK+k4u1dnBN97yrqz8psEnSSsEj/Hh1dQrhbyy2zoNYpl9mtDsCubtqu9d
HiHYD3e2Hc3JCayLHSTWYH38cexCCPICqD/uI3a/QeDVLiDk+Kj0pULiqHhn
u0QWgmi3LhiWLOI+ERpz46nlGOB+bqCG+IDtdTHd/UdFHcPPR4ZrkR/bVYoV
v52pTwrXArEFeABDjkToYO1JpEcDXQG2+FbdqXPzN7+HeJ9IuXU+sDQUmb8f
1rY1TwBTlZ8UYllRR0zsaMX+6yHYViLkjRoBtVOBP3vwxCnCm9ofJa4xc3B9
f16fiMOnezxOcD0o3QvBPvZOd89Ja33G7J8UDn3KS/P/1jvT/22o1TpZO9FF
hjSpwvRp4BcqRgprUcfqQ/iZe+jTXsepscVGjZUD8ZVIvoFZwdYwUYIpripf
XBjXE+e5fSZqLFxLCcJTb0NO36gOk8+Z6KiW41GQj7I5nclj+xKmk4lW8VRj
V8pNReXmo4wv/znOrPCtS6ac3E8UK2Ascvi8kj1FUK2Nn7MtSk8DrhLwUedA
KJLdNSkAOfZX40PFisV/gYvdL9XfPwBLntpxm1cfuoexSdZQxEfJPp8qAlJd
HzTFxQGAYm3cAMdS/02U464eOFWroEXW7FraDHF+9p6o5ScpcHk7Mz1keFDk
G94t6Xxy+1NkjMYFxzWwCeDPfuxu4L44Aknq4cRh0cM50dxwtwHmTYEJzkAq
1aZUxxoPiIo20ZPyrqn82YCgdqUDa408lFs0W1/Prg3WnCzcp8pa1ztoiA+y
6iez6O2cQvD/j8ZaomDEczx/VJjFovGgS6hkcD6hYOdcGQwGpSgk4FjXq4hN
k8xFj6+V+K94E0GLVTgI6Boztj6fZJ47Pn7CoPQrVxDqV0ayZaGA5pbfjDtF
pUkN/pGTmWQk7DTIJJUb+B5ZVgL7rxsmaeyu6B4nJqumB9pGKs8vXir0QdbC
o7C1WBUiDpiAmpQ71cZA5Kk6J09B3qfPq7nb2W8ruMlXvmI5xXjefnRzcgWO
tWlYb/DjPVs1jVU1fnpLPK7zeRrbHdMHU2zAv4od7CvaQJLGkozug7Cn0IZ7
OXbkERT3SdJEzgVFH+TGq3AVdEhR8i0Uh8+gT7XBDWCXHYBjQFCpKJVdjBTc
+Sux/+7rf/4MTgpqgTkom1PhXMuoRVBB5b8RQH7F95f8NpJ7Jyyr7/PB0BZG
LTB9cN55n9vH+ry37sVpE/PprfxOaSt1Dl9TfECvH9sU/iyxatWAgb0F/cbd
5MCaV7rn/h9HQkDf5/8B6XfG1CmLv7c7IqnpNtASXw66P5hWF1fXQuWWy9o7
Lk9NiTRk/7yVw9F9IUoRFlIfNPOXWv1+oGM4i59KN0ty7ON8fgNfn2stPoXG
qk9+lh+eeH5IGsv15r0qnMS1fThqqDrgptIOdb/H8iUPx9X8DnvU8l8UJF5T
oqxwLAY+/t9uGrXeAXEU16aBapLwbUEBcsj7GwAqVwLan0oDWTwTsISkhevp
J/m0hJBscevXZPLG1YhPHS3nbNXz7S+MB4zL00nerpvVKsPuisCkHHZWx3xv
sypcpEVMf5X0tyEOQAZL0Da9LgzAyXSQMoT9akMOoiN2RSqYVbHIhk45LHwG
+nm1/QdaAVPnyyfJzdosJu5xuq2yFl99m0rB5Kkl8LrxOaf2VxmurfHN8ddL
GSFM51zMidTSN5dvfp75DsZBbNLNK4wSIjaElIc7NK6FDABGH68XWny9vjiu
j029wDPFMYIgqUHf2XsttpWkPnv76TsIL1hyJaDLRxmhuule4fFVCuci4sLs
clslg3U6NAbqnI+YsOXi5FlBjgUZN3nRUGXvRQYJ1eaH6lFt/CiRgQqwmZTI
9UMfDVVcp8A3Yvt0TTR/SHl21ygJYWkm0FmDiOnDj4cNXhuMHwT2UrhdBPFb
tmhCDVYXENg5xtgc/JamVipFFXEEwMVYDdYgOU9VngYpAReY1N1imT0Hj7Ox
FPopECV6q43At/a2C49nPGGdcURTt0koibpGxHNtc/ZnD4fj/g1pMUm3HM/P
PvCSZ0G0d2bH00PGr4fHfPs1hwsihiv/A382zApJUe6zj64anzRB066qOPsQ
nWrwJKsZZ/Jak9742xEtOTD2eTER1bQ3CAsQkLWgZ35q4mdBNHhCkXQPZcvU
9We79deMXNbXjjNTO0FSTT5w3Cs9/Ketj0BNW8ORyGAlTSw/jLHk5taOt8fy
JTxk78vQdYKcV1mt7aq4b2MqoY47A+UodOGT+vExcHzMJtbet2dIH2wOgjvw
8K+zgLLzXqc7O4n783r5Q+KSK/Q1DrrtzHe38lE6X4EUWGlww91+IZmBrs20
PchCqu3axBBFnIkD3rAMrMtW9zcMQCHJ4+FpS1zODyFURN2YfdOLphBXZp9s
F30yzHIP+lTJ3o+BHRRslVeEimerTsWip5De5fpa5np6HdfAoSVPvyA5KNbB
ri371bCHStYXNpYCWpnvCu23XJENGw5u6Tn+p2sfR4Sg+Om+cSPkOqm/i6v1
Um5P/24INGWstsNG43nrZC+kuAFIOu1d0TWsSXf7FWg5bc/vyBo5Od9Op+lC
tFbDtrscvRrzf67uyZqG0ycVGEAxQ972l9F/lL/sFw3Qge4iEKnHdNm1t5pe
/Tad9Yj5P52IdbFYCdSFiBWNdemJ0m0J1iUE+e6NjYf1cw0nrNsW79poEw6c
1tVYo9M0af6oLwyAjU1eVtEVdaWDEFcDAnuBclnKbNOSFYNg0570gYvLE0Wy
UFJYLJ80gBVrRqOeW74Wud7rslGlbgq5VW2Twk6qGdZXUQOD5R7WexQ4O8gQ
x/c04IF7O/Xk2uxewp5POoIhwxKTXJyxmDzVUdPSYFfjU81EDOZzBLeRUy47
IXKsOVS3D5iZAopezPcQ2rGCEcfv0m4oYrgNJpuFB6Ua1Jt2k287ZQmhZkxh
vkYTLBuYd5vExz8X/25MSGUYiuPoOispvh5CB4CGVExz12zb/tMc6jJCyWg+
ApWHHPLZ77Ce8sjVdSFWA6vJ4F34nkMpHxsGLzxv60/u9+SK0Sbgys2/6355
u+dOYwT3Ar1AI6c13kuzZGpuPk9xrRWlpbJNs6s1PU1XYghCGhPTFj4IZyae
MWXtO3kvaxmItoFsLrNKaw6c4BmRl3+d02KAf/ztG7KA3GfFF4SIHAtmY1ul
9K/jsQxHVlGc3AJNoMVcQX8iff79tXf/LnajYhEi+BhxdsHXdTc05UVX4MYr
cOf48IYqzv4jQMxkdIdfLo4vcWNBjwh7QFozqnjAu5jRUOOt3RNPzJHoMjt5
+cfmibxN2ctILMr8kRypWZpLRIxnsIivHOLYpFHiIp2v5Yw2w5ZamezerpPq
vYrNRuwhth3BWOIWEEeY97uSYc1s8bBxXukruRiEJKmbQPYdmNwY2fsUt2m/
kWNT0+Jgvn6U75PddLXYWLk/ps0soAE6WldgHI9FcY7lHZWjlA0kxS+R/kaf
PRfFAHeFCDBu1ydaDJxmsxMuAVes5pUpClL5TBim9mW6Uv5rJOmn4PQN2JMW
GHnIFrOdMRPtt5PcPWD47wiZ20GEoJURWqjp/ns+G9t+qHdToRwHVpcKP1ud
GbWaxMVXLU8YjVRBaDWVpPynQDbVbcli1zBg8yoZ1kl3KZO6/7i/itdLNUJF
811w4rnjLf23aUZfZlzhj+L2hFWtyBrFYT2NcZibD36H4sb1HJyceTkOHfzX
WDri3mEqCO69wmEDpNP6jCW5OixW19NCFrD8sSwbtskW+mF+GHYNwZD8DRt/
lTla/pbHk0jX9VB58B2n/84YSEyu5ihEa5mD4pOfrpIMrgAhFPF12EEYjun6
x1DDuMuS3TATFwGiRS5VJpPcpP6QxEwGAiqkUc25mYfRYPqTsCVCWBLCKCRn
KK9iRlU5ttrhz3eEJezaR6RxOd1t1S8BNzJxCmc1GFSYPvCy+X/IU6fD3arh
ZonBlM0gTC/Bf7+dNdWWL3j+5SYwGV9Ztq4aw+qfzmXO/lx2KAYNs9Tvv5a8
HpZTzhIiH45Oa2RqN9tNk1dBYHBGr+SJJcjnac41IusePamPd+uMqO3nF6fs
Qhu4elorHFDgREaDRWnq99gm8XD2uSg5oc3X9Ibsap+thYHjFQoX/c63AS3z
Hn7tVEifQs3aJT1SiQGGwNMkBGrVfg3nCtbcXxb3SiOSTYplW2/qwFMIM0PY
/o9Lgqx/GVEVlgdq20pfbOshMvhA13zdWNZSOU4VE17oCSh3Xb/r7nj6TCRt
B4ueiZw/6srjYCk1D4Yq8QiT2ruyadEUlw/9FU4Zu/LFiqS6RcDvnuD3Waci
ZAtlHVJGdv38zX0jpmans1vT4Eua5+E+ch/JAUCR7Gh44pYS/NVhoyCR3e/F
RWL+hFGy1rJIpKSq4QAboCBlDWvL9JVfGHaWe1SInwwi9LbrpuJZ2WzIbHpC
TcH7RA1oIi8FMaYQOrPZQ0kFepbzDXdtykzPO5Sn+Wifr5AmLlBv0qOu333A
srM2VvTGDqBb/sb5qDIkU+B4DfMjDRPQZOkGJUz2Z6aLo2BJSz89NlZpkWlH
3Bmgtb+Y3BN5kfyoFkAMaxmuOiYLmUu6b21UdNt/U9+pfGyYzGL3/K80WQFB
1peuh/0prr3UnLVAW9YPWVL+uNjJ62Sf/xVtAl2Z7qG2IQUVwEZNgVyjkJFs
d/zkZ5dvIlyhnQofxN3yA2mU+rLTwruJMGJz1u4SXwTe+HeDfUbozlBdlIrx
xUFDOcSZoqwAh95ih4iRFasvU8voyC4ROh3A6deBN8TqDPfO65PcA7VoSQri
gwbREgn//3vGgW4rcOVgR/vkYJYdAQ5CH3XWAnDHb7EUN5N3yih/oHDlrpzX
EBDHr5nitvOkD7ZGlexXzu2CtFofAasRszTszDPSBHTMmkEROOgynwUFUvIs
ZMrISAUlm5S9V9iF9uhsRpJHUIzP5vEJAH9nGNDPMwUraqJAFss7atFVjXH0
upwvbcchgEwaHVemr4X/o6C4YZicX61uSafkazWeuHKXrTJaKkEVw8b+Y2cR
cPtgi84Y8VgGNE4wI3rpsIW9ybNmdo1elV2GznjLSQDb/IeGPclv8lmC5O+8
WJIVSyTSfvL4/CjqVtupEOENIMLnJ+Mfl5Gy7oFwaLT3wxRVCmwIBgrnmna1
6N3/fyg7yNKgZCBEsTmtpH2YCXZ7Bid1mAz+gaR5rkyuR/VBR1yiLatF3szr
oCf2fy9OpB19/XjmVrHMcbK5jETmZ6iI/KiE3eW6X2MDBWRjfP2RfF3NiHLG
EA1MnMAv6SUxBQysa6kRHl7uvBs/kNhYN4JE975ZO6Pz8POjPptfZ+yfZHQQ
2HBEZ6Dfles944kyCCHzIaty6Q+6xFwS+RlOb/XA3QmqF7XGlV6N6xbIO78p
9//CdKl7KaOunm85qPdRKInlP41sNRKrcm0fv0J7VEZlB0feJj0Ex0G3flPS
/vyGRDInaEwuFlQ91oU3X008VKhoxQSiZHKR2ih2PHBphg1Tu5lAbweUhxop
EQFCMWWO/aI0mGljaUy7/xCCElNVh1qg1AC8eUvaZirZwrBnwG/3YzK4sF02
MFChewB4Ver0GCNLC7w03aiimLlGK3kxdo9fAACY5MU7rLO6u8xgSAvgBrpm
vEFALoYwkXKG6Kr/hj59R1U+bhXx3LmLTC6pT2pxpGjM/aFvj52cABcZz5oz
IeR5gfLSnIB89zDC3lxhF0afZM8SAFJghLHT33I8osXm/G4MYiy7LWZPbwrW
ALORRreGm1LX3gmOc2wfPKiaBVVP3qsv9mZrl3/Z4/CyG9S+QtXS4/PLrIHe
YgjEJEptjoJCT9fNSuX8eQY31IhEEAdARuktOB05B+0q6HW7+P6lg+XB03nj
gj6f2uxPN8XhJnPvxlufpU4vWeA8KeIpIczxMl2mCoYABk9WGNJ2TDa1ftIT
209eY2/WMBNcrFoJLX+Hw2cuKEhFE7oduk2umALD7DHXXPXK35gjsKJJ5Vx6
BjnkkehTWxieu/iwBrqO3gXcKy/Q2Ro40xg1Oi10lDKwkGYDg4qs5YXzwEKM
CEeB11l36FWCslQQWO5s8SU+U+6/eOvzoEshmNl6SA2DzU7UvxGWj+iL6Ov5
ahpXgTHSx882LK8ezd8xspKkrXkYg1PsIs+G/81N+l/NL5jBsW6J6ocpPNgL
jFZ8zp9RbIVodsTjs50khyhHCU3D40Vet96CxjDDz+ofTMkINXrfHJo4z2Bu
oZ1mKaMHw4ZatYUwjPi7DvjOlipBPCUT+BFjzqzcy3ZepuO0v4zc+UTVG9PZ
WYpw0CPrmKc/ZSxjZkpMqMBoYhxGwz3oiYgPSuAB8O6dHQANfcmvopcM9TJd
U/oFNwJfivrG20PQ0x4Khzn/LFJDKsodLA2E5bjmvS2Xt7aLCcAC28z8TPib
5td4v78GkPUZ+ag/DEEWjN4w3tJ6qlOUFw4+74ajcWnYm6cDN8bQwmiGXw6V
NAO5KyOQ37cKaTpQLoUxj2jGIfyC92W8PvQIPMHj2C6Pl8r3x+EHDJnm5yOw
uBjk+nnsNTMlALhh0HJ3flPs/ODwRLzU3eHGNDxjI983PYgOC2lJ9iIPFzGh
ruuGlCB3c2ZUJ1GSnCJsLzMMW/x3pQ/W0NjzuGvhGU/B3dhGtG70YJgX4e23
otHwByPh10fk60q9mNOyfkmBUJp0RAETIQ/ssBXifWXh/tdgjRPjRWKs5Hhv
8qrHjvgiqYq/rd5S4dh+MQASGTgylyMU1YwZTxhxhF6ii7Juqp5PFgp1VLRn
VPdP8FrRar8CeHB+XMlZIByCiYC7Yf/3E6HybyKB3K4LDRKIsR9+RBsz9RYd
JrdXOgvDzlidd13gR4m+/1C+g8p8UeMwt+ifNxsFPLPxZpphBOtHsjBNt+uY
PI8SlIGPRQYbVQJM3Fbocf/Dpn9DPW8nnoOCxTxJmFpxBOUbnpp4oaBd0cb3
gnpIFFCghQuOeY7yphu9gK8Yi8RaU4FpCJABeeSkDdJivb7wOGOyzoVZNUGQ
DMX7nAwHoKjsEtP6gBgfyG3FjtB0YA6mSvhGH/WhssXxwa+qYjfIkANUaGnI
VzO0jjVNw3/HE67udDa8CF3Q5Rl1eB/rsBqhiWm4uhS5gvtRJ0bu88hdeIt8
omaTDZWOHhp3y8UiSgpw1K15Jg5dYLd8A91WQiPpGmOhMPmY4W3GDxtOnpaj
j7gXnJSCndQ9GYcE7bh+pL/wf7qrrqGJzQANe+IjBnHxHJHGi59HC/YBvGZ0
CHtJ2eLFq02TRhgwlDk549QdBNwvR9d6RtRT9C01Z3JmcYHP4ral568KPCyX
BPe9xK0P1SO4v5q6dsIt2X18g3C5F7AWffFz/m5KntvdPf4sVE96vKRtC/Vu
kn9N5OXmE/cx5d5lk9RWwf2W7vS/hliCukjefw8XZ18IIN9mDf2WWZ24nNza
kcCP4plRG4ZwHsQdu1K9BY6Z557O8hBFCnk6Xh9czK08aECyaQjuGzUTs6Lx
+YvLdZ00LNRGhO+lDj/fAs2oQd0Lz2O0QOpiIMR/3hU4lImWyNk9lfx0symg
eLDns5wtrC8uUYVXphkO71bEUtfjmVengi96tCPzlFZcZ2DpshNOnFKSKGGT
fEjJozyGflPO2q5+NU+JGxtWiDjIEqNhf3ZiwsNJAV+N3vE3FcMIqnG5Kpr+
jnEbnPys/ykn8pumTYktE8nQyEYUNjRrjd2VUuNEP3q81qsxwxSouz50YknY
8YduBwoIpaTnRo7Hjr4XDqE/I/BTUOl1syJfDMdouvRbEYea94D32SlRJwEs
dYjRJjSEaiLYSTsaz3LsuQsyooSfc6/FIn+j9k4u/XeTOq35hea0DiCNxR1k
/gWZyjuKfIGGbdWARMU6P8eoifjx2XXjG8JqHt0/KkYhYjMGvpUAtN5YhS6E
HTHE2Urx6KlHngAj0MAUOZD1gPNjPxa83ZOx68aLZ7O4F11pAQBJwL8q6qTb
KRD/71RWxXC6eww4MgqQcAbkPs69gkX6ewmslsZvImIR1n7Knvt+gNdH4s33
D7LlMOtmjFPIIc35Kz5Wr6wA581+ueZ6z2AGvIcNVrR0vpGO5tWopcofEdox
szA8ILoOzbyk4hm/41P7I3neHANvrwWvPZQ/o3y+e1OV+3110+IopggQxtb5
obl2jfZ38wWs7y+EfAJJY2kV+wZtpCFANt0pwCf6O264MsdqdmRkiSN6EexJ
N5Lz1nsIF2U31TBBYwJZUxnB37DtAGHRYZvt7Pi1Z54nUGmJWgc/MmVp8XTQ
LTBTmFG5uzY1Foz2AtNMVRTWOH8/4mFniBrOvDG0mK8hDNQiwJzX39sfDMKv
m+QY2LrgV2YdQpfr2qEptMPpdPebbb1UOO/ljiuRKkMZVcHx7LmIZ7+p8Q3O
I6ckCIW4SbQ30KBCZPDzy7cFHOdbFgKMjYhkcfq8JK30vbaWggHrYc5pIpn6
zLzYSSUR7GbsuGf+SYK6T+Qbg/yU1XRhpe6SEYtPuWixrF3tKxHIySsPsrPp
4a60olHKLvTGG/5Ukt/+1XDo8Ijz8YaXu1XlYnO3iYyVfuDqHGlWDXwDAhbF
esA0vrawlG2KYJpTuEmo83q9Dsjp72FsXadE8i1JtH3/wVP5MS2M/bAGmDYi
4du87DeiaHblsTRpinpcgnlLvnaUlcU0lx8WWwVdz3VGVvg6pWrxZO4dVssQ
URQ4jT1SrDCHEvmrRgXUwFjJ/eO8bIdMc/77jvRXAsZX6QAHTh1h75wu39Di
HFLpavzjEpxrPVhd3n3ufIvVnvpTIq0BodNFzWxMQAcUqrt3bJakRHtcCAQb
+lvMbdZOIzuQrZ4fZIxOv1cGUF8ZVh/AhwDtjzZr7mT+OqLYmxlUwSfqQOPs
E9qMHvj9W197iHCfYaPsWlH+E294ejtBfioUgHX71W/WbGy8iTK9MjizPHal
4rpjgnGpEYB3KtdCt3JesWASmMOgeqgN3cTlxGQyF20IyXz22mL4FOuxakjb
bOCN0qElkavhQXW+zNu+oz5nsA+sdP3NybvDb1r6pxzEGOUbBDPqCaxc8czA
SuT/bRSNiG0GZQWj42r7JOi1f/xWMw1BjqJWxRacIhlsYG79/t599M5T+N6z
GBVAs+8oFvBMldYrTAOV5RjAVnNHqKJVkMVWhJNQp6C2EhFPetYyJJb6729s
upv1gLOD+z7r9n7DT1Cj8M/q+sE1gyZ1iB0CVrWJCz3e8JXIoYs9INMWl2LH
KDXfBsuEqKc/IfAJp2hEzChcrwPTbYiDLnwE1uYE/HR/FzP4+a2LKcDUIb7v
H+En+Ox26oPR/UyH0Mhu7Rg8ftuWc6nR3GcH/HnoV877YbNglw8OpHanNJCd
aU9HOlQFNh9YubZ/UnUAzQYtjK2joVn9IwuQC6hGjSraRqx4uKtMrOQXRilg
bzZrE2xvzZufAeNz0Q44lCr/w9bsyymCaRRTVBPhpLWNBxkNFFlJWRubqYe9
RudCQ2zu948wEw5ptZd2LnO7gTUu27gZd1y9SKjZX9+dn7YJ6fpJtayMU6wX
ROzmyvM2iYKPhsLS//cN/E4nzdJaf6zqWoce0TkWjWzp1kVFdgHevecpafej
KogNtqh1ymQ+Z+uSRkLzPN0U2qJa4fDuGdJgLIlfq3Jld/S6IFH8XfcBgYFv
Efpxu2U09gkTRkr2Wg3q2sJgY5jwp91C79zrvubJfEOA4rpThWmtj/x19ROd
zqP05B3zK8qXsJv36DkwsaEsjLkYCYKvRQinsz6DEZlO1wHJOpsNm2flHJ/x
zFzRHy9ObdA14hLwzwgHyi81C/abJcOkFybJq0VrGxiqO47IjerSHjfISD2T
UQZxtO/Z8/8chog46Q66UgRtUgWcoGZtky0umA0nec/bBSWh7787fGNfjEqO
31KMZSnsozpqdeV2Z1X01SCveEm8BMVc/sR4bY1WRODJF5Th87hFnj+ZV4Ol
3dMcD0Kdbx+rYcWCqcPrVHMtoQXior7uVTqKoAM4b/8qEjouKULZrHP9wTY0
zso+IFQuZOug3tBfdStTyS7J00W7VeEn7BhJB0bKp1QcG9wDc5YYcZC1wbVg
yXqnJAtfDtdPFgKdR9Cc1fDFLgdog0/uQjUUz2Lhea/dfb4QGUMvNWhIuxLI
KV7gUMeVeOjFEPrSVbrEWONvsIQuf4ebFz2JFZelJ/L6Vn0OuNas6WsPihYD
Hu64SImKdSq+q2PLj9a1Om9bMnqaHdxX3ixM2XZuoZU88k6Fm1ELjH1FdExN
M383eYZs1dvoH9aLYMZquhJLJ4ytfb5DvZvtPLDDsZD3rdw7/vylcwiZ549L
1o2iAPD2Bs11AMnxkX60TVuuQ+59Y3XTLGb7+SFZzOKIOig0YEilD8UdsWXL
9NCdVbf6nl506sInXXAfguFlcWX52TXtmUibKX2oX3s83dXG5qewyVyamKb+
zKL26kJpZfX3MtfdbZOm3lDc/J5otq8uUr+KNreeoXlfK9nZHePsA42Rh5/A
Lqgr1BkPdYuBVmIbNXMr6apLE9v3KCDQNlNI3zXi82P1jJRl32G3nsNCZ3+e
NEMS3qH+lF09nPntR4xXJNk4+4w3vW/Tn+G6v8huIFu1KIzENDdpvr8Z8KxY
oUYwU5gSypdqxGCsdOC2woIm4B/NEhmA/voDh6tFbU2c1XQG7V1dUimOXrGQ
Kj/B3mqw3gpoOPLjAtDfh8am96zGFHnwfo2d5nRDT67ndHhgsbg7RQRS4iNB
vuj4fiZkwbsibUQ1wZric1LMdYJ2Tzcr5Na+y/pRyaFM7kMG9D2pLIyqarWx
rhgqEnbgb91NWGgtLzzI9lJLL8DWRlZdVWGP1YdZZR4buxFDbj3mYE4dbFT+
o+X37pZl1ybu+mV1a7uJg0i0xO48lDUdTdMA/pSDnecUMNOQIX8N6wjgWYdc
2P3Ovq+z5CDUi38mg5dQRwr2vkU7H8+z8HLaCh5CejnlW5IBdKvWoLMOCQ3L
VCZKN7HWPKzwKvAq0PSHeneNhTrq0eYeZj7qZp1HVTiVVqdswzQ/COcupNBZ
HIjWdl74a0zv3H1leDExdIG+vtBTUc+o/ZTFRNyZNMvNfuGjS8JeRf2y98v3
bPG9AAo7sA/UMVc+1xuqPItdy/woKvb+isXsCwHSYvNgbNMlepKtyO8xpaET
9ErcBlP7mPxTMlSMqylgcyi5c5OloR2s1PCHectScmd/4tWI8cFPfKGiHst6
C1EnCTPyBWAj82qy3f9yc9FXOh568X6CFFR47eqgOQCGn+ENWKFh82xVcHs1
ddvfiD8gFwIta5bjTwUifSyHKDv9tT+sBIv0mgQpsOvcJ1huGMp8Twcjqta4
n01BTrTRYoSnQrxaKk8dFynA5wcWWBLsx6dZZgjDlMGX9rM38orC0BgChFhY
AAI6I3ssRt6tXIDjVEveAutwwgGGu8XlZxYZpiRqA5YEg0KtDFq0SU4Ni4aJ
+BONFQoNPqpRnzDG2WCtd/mDrRut8K+F+Xq+g5Cd1QRgKqO1/LuJ49Fv3Hl3
Z6MmVXZlrM2rhOUtDznJhh9kCj5ccgMBbI6smrbu3yHAEmCnRVy6OFM0YzVM
5DdLrklAd2dLxNaxmxACObLF9j7qYdUU88yRvtPJ5BDHceexP64JUngXcYTJ
iKn7ZDFNFCvWGyZxNS/vO2EiU6p6Xg6J7Or8QRoDkcnIdpcHfhW4OeaDTvJv
LDYwyV7avDXLOR+lQJqw/IBwIvZXotmDi/voUKFc6GXG0h7gxsxND9oMRVxi
qw6jPI5uLOfvKyiHZ26hEq15upz0FplQRKCFSi6woMzIzL94nOjYyotI7jtS
JBvu36QreW0ENMTKRdrzSzubWggn3fh0KAQAKMHtnG47qXX+Num6WjnE3sXt
lIH7jd3PbUq0uyMbC8P2+VPiWl9qqwN9r4hK6JlMqPtf8bDtKnBiRJfvoq6B
FOnnv12WhfJKFSswJZO6cEkBwvfctiy7lJTFkzms4D2mc9yAdzOVzlFYiKLM
rZ5nvfC3OV//5/z0t54BWGrsFvhwmWa0WN3oULw7NwSKLRpGKeOLNAAnKziR
xOTQpVPy+q8PXV9wcZghQIRSfU7yaezrWa3uv5Lru+m0PKmJD6AiLGXzKlQO
FmmNzxhcU4J7oy647rdpiax/zRqivn3zsHGg+JvquE4C2CwkGxV+naoCV6ho
D8NIrRkn/5qjftueZ3pgFi26dW0AUHXoILCWLIASzSZUcE174Hex2sygTfB8
xgrbY8rRxAFvUsBxbRdwdc211E7x7m5RvQkn4iXe+JT0FUMNxKiINhpFG+pK
hj7xYLpG6vzH3sEUa4T0MBg+HB3eWJhlpYFVbvxogw0KZtX7JhdH90oiCbgM
6941DgEHXRt5Y6IcHilGOzmcCaqqhbntyBv4bZpCub9cQhJ+XtV6L3Uc148/
egZC0Zu0lblmd2gEHq4yECAYrcIvuh7tK3uL5KMX4EHo4jWoiXkuzxy2jJAz
N1WQnpLjWCrXZuaRxOp/yAJOb3CkHrH6G9ZSZ/9zGiBmPkrnXpI/9aYojvMj
YvhoI01w9xRXaX1wcJ94VQe8rL5ZwgzynA3RnqHg+ihvigIHpSfWB8K6VyJT
fj7MBJz9qSMZKG9yj6D2QKx0o+8TlxsZDdhpMsLucEk2BmP7JKpc0p4AFnAM
eYZcbwMPf8+O6AAQvHH2MNp6jVC2YsN/UGDrNDBrpdb2u3LYy8XMRQoKIZzO
LlLMaZz/bFNQNGlaz5vPLs2WYdjZoxH2eslIAEudS5fSeOc5MOgUbT/hncn0
aow26N9da6onuZK4LQWs/y/gPqWE6HUm66OE9DQCTUGtNqD2CeUaef50aa9K
PzFVrk2iciOOlSvxThlyArZv0h3JTtNwnyCeWOBFuZxgPLd916lwU4K5Krgh
D3RudCWFrw/f/0XnEc+B1TNUOgvluUPtfL5pRiKlOKjsfl060kNIVNX7Dijc
Anrxdq8U0njYM2Tt2qA5s/S6L/NyCnpPfasp1xyScf0LDKoAQt5Yup7GwM/p
srl2V60NAvQmTYsBCZ6TRBC0SxRqesqAjV/Dn+uDiOGagpw8MAH7SdfmIhnJ
NUYKz6yfgOo2Wzic9Zr8M5lfkxAswY2up6Tk3sKCA1fxbMfRjREFRN5xNJ+P
aCiXAv+EYQ0oL7cQ88uC1+vRsGoSqOmEtuVJcG99ukiOClJa4LRtqWs3ooNv
tBB0R9V9JUeSThjCAOXHaYJUJedKoAckJly1fPh6bVGf0wTFQgdxuTegLO1h
aKvRa9tBYhIv9Vaof/33cPOuSu+muOJQnGuxatwN9mrTLJBrCrvF8jyP26NT
Oyz+R5hH3z1ZbvZHU9UCu4PmbRhFgHc1WQ1x0pFywZibJZ8cyiJYQIJ8HfJX
7dzJt51ggarMKOgHLpBehlS5cgqX+67XKOtqDZ09wlhaPYIV5YHAEjnLg2Nz
a7K6MoWqBRLqx07lC0KFUdUw+Dc1hIXjXfQwGgrIHP8rhNtwoBONPuS2NIge
HgBy2+na5UDoEnap2/WWJ6OwknmpK1ED1w3XG86goRl58Ci6FU6kfh8F/1Ry
mLYskGufedA63ZDwSc4PtQpfAmNfDswOXGTJxsmIBTHUT1Nrbwba4CemTeBV
oHEq3czJfd/BSNVbXkCJULw0EUN41JWTVSr/KHhJR3kaKPDTcPiRGXp3tDRY
stydZiL0JJmbpGZ9fbYBu33mhFw3v9W86n1ON6EgMYg7mJ2N3zG0UD+9djdJ
bEynShBYjpkfwM7GtSXpD76Rrvx4fcLJ/m4R76jvhAANmVrz6t3QKlroKHlV
yjMTPIxMblInodhZMosNH9y2frdb0b1Nniwdq/SExw1EGvg4uCGoW12lUpUg
UyEz07+mDGlc9hZPh6H7FK80fh00FlhCLp9zX0gSsUvUGMFOW9skTSwCLBB4
ArKeT/Q/nb4w58+YPvEN3YWUynGyHZjCCj048am9pRBPUp4tlKfGmdfhRcVa
8lf67/H4i/e2DDQcZnOHlhbmmBP8ub+a2LWWHnOhkl7Puq6wjirWrRuvDQNk
ML64OTSmjpat0ZJLdPL3MiT9wP384nA2mHbLeiaLkM1mld36xouMvqOnQ7VH
7BmzwqU21XMbXbF6hD+QQviw7Mb98sCNeE+/MZhCAeFQSwd617F7H13MY5cd
XD3MeQOhtGVTSHAnwDhXd4IlzwxO487xz2buvWyCZ2sv3yI5eWXByGb1ZTGf
I/APYgMzRVt08ZjyV5HdrXYYFyOYJldqd6+/Pa/T6nvI/4elCHABwHLNATi8
VtcBYKOVsRAwp7vZQQ9yyKb5A8XYQFor/zf/h/YRmb6T1A+e4IM32evKlkGq
eWHAbGqRT4ZqlWxCXkYcEZyee97fjG+C9EJLM9+v3CzoLsaR21vzRXjcgQM6
Lw0PBUelbqFCIw4DKgWWsk/nWwsWtsJd6gIH2VERcE7a6ddGV8q6qcA1vOze
jrrCeDBk5hsvODbTvGR+10sUZoyr4DeIIALZ/nS8pKNKg8bujbbghvJabYn2
hvdThgCfOI4vFuMuJkxnzG+nIHQYc1kt2aJVpvQAXw7RWowiysgqwN81G63g
aB0ETd0Nx38GDVRrJptNLwqFjF8lD3dWN64lswix5AGbapwo7w8n9JOLTcmY
ck4aMV+JXKVSLYGnROUd313VieLsRC/Qy+q1YdV0x+WQPbm02yGSgVrTOtyg
Nng1oVcmDxRlBJbD9JPzSAZU2GIS7k24RG1YH+NdUkdUb5j8ju9hnWppvTuR
kUUrzK8M4p6+U1e0UgB9XnFZVHJ/Rt7WzxEafzkvb4t59aOZuU/9GCsdhNo3
+6xzMMtvSgXse6GQfdQ9pTI6XaY9+smzfJlV6N0/QXMWO8jN17/Fbg6Cf9qV
4mo0OieMyEjs7VpX9C3PYuhP541Ul2bGe8tQBbxcp33hQMZCh32p6EJ9HBff
yMMwJWtDw62S6gOeae4YNV3X1+zj/1CGeAejxJLdqHoPjfxtR1TspHniOthn
V3GKG5R00oUY9HAqANif57HDuBQqKih/A82FQubpFsQmAaZpf8k/VQSlyHES
lnTWB8PpS7jogk7AA94H30Dt9icsbWGP/cKfjBw1PsJLXR4yeU/S1c9zt3JL
wFMWoXu2E+tfScpBeun/TAsX4MA2+bfRO8AW3TeVuFMCN+ALDnY0fPn8Z9JF
Mhi3BYU42pzGc1mjgkYE2+iXIFSlnmndz+TBrRu3H0MBNJu24vRPx6wexIZF
hLcV/uwJdZ3DVLDNlFpgq+aKYf0rsdF8WpcAQrGxpnbQrprn3ARTKfWL8k1h
vDvoXO7qIIXT57A7dBCTEubv5UALIaEzsQeC0xkLDDhRnfXUKZAlVrLhoqtP
WoAuCv+nSEWtN0CGVpTtuFKyOewtSyrIPc3BKkhh4bNRX67rVmo8tTur8Pj0
bCTobY983Ke4/iqNqu4dj5VnrSxj2LtbWn5RGeeIHBOhDNLzbZS8kEaJm2Ky
UydLZ5gsXYMcI77WsA1FTMoyHOwjIW4OcghvdM4qhoP65ItpL7rU8CqjfbXS
6Bn2Zqa5juCKATgLGOH79tJrJtmGI6+EBAl5uIbE7gpW1/brRreExoQnwyUT
fzlopyfPidwpKapDU6PS0pGjhCIOWtiG5ViWC1ZG+eWTXwaC2eJlrpboBCcu
7pZJ6JeG/CT9Ln9au7AoXKNQwAZS3x8ro3wdICXiKzC6XzSCewlcFMZH4dLu
cP6fxXTlhNrcJdLmar2QJGFB5nc3M+dW4Mna4AE0jG3qg9TPqzSy5QCcN0XR
7BvYXv/ZZbK61zYgan527FByULG+7WmAcxX8+mA2IZIbmIyyiHbc9+TIqlib
KOno0QqD0YHoxJjLPM+vGBsxDFNkG7BeXebj0FkDQtJcJx64928EeLqQngXr
M4AMUymS0Bw53QcfRBy0ss0wxNlIgs2Enlv7bwUgcJyFfZJYGsbK3JtySeSv
CclViy0luYx+WeLXnjDXqe/ceSYbncHY/MGuq/g5kuNNzq/Vn5m2y34WRU8m
8ebWRQfqfySqxaFxe9pdG2QgQQM5HW3I/x4RXB2wHmepkEePtdNpmRn2e8+6
olWHI1hbmHyarIPxJXSAXCgUz+MsIuu1qRHxeKyZeWItQTgif33N8Fr/LAPD
kEViYKNgZn4CIKBfP33f/SjvifhPfKqPN7N9OpcK7CGP4kLVBNsgiJ/U9gai
Jn/a+9BgfVhGGboQ9WevmknBvKRT+nEnKYLF86YmwVMK9kPLFR4KxbMivRoQ
4xG0B/W/II0GrkNfpNGWNuUOriJ6uQyQRG0ZFYDwIpTvI88cFy4WsLFuxk3I
sqC+auhltCFwQM6kKPn0U7zMB70kkqdouUdczfCE1LRODCME28Ef2CN++IOq
s+CGYoLWyA8IkIIoZuvs7jNuS5wAvJgSXhjtqBlQvMVuW9+DbH/nN9YKOrGh
kwQGZXoRL6is2L3qVHfgREgjN9kPRbxuHz6RWUIeJ7NUlBqvH33mX6dRAEDn
zHWI/XJsHqjpkO7a4oOoGN5GXZuEWKBRg2oCnE1fqg2g2GLmfc2LlNwOz1Yo
g/lS223IYY5Qpa25JuDvnwjicC5C2nUkNc5kxdiFTEu6BkaLjwhun4FvrZKd
sHYLvPLjFGcApXjj7F4WRt7u/grzKIDC1KRrbqMc9ZlJQvCmcA8Ht89lQ3so
b3eir/Rju9bJ43tZSAYal1p6vAkw9HC38RsnrN2CooVdwTb3UgOggXxco7/D
DqC/JjxhInufBFXAtGCvhTX6DUOvYZ+dBUh+tEggfgWTRhK21FR8D+tfIOEr
FqmCY5hAuaPxXhKXKZERQk+vwNzKdZZjTheHpGxScznEQS9OF8w2fyYx+fYS
V28PWstlTmenQ4cH6gxjZbFsZBahcc9NkU+aGkElKOAHLhpcm2pSMe9U0QHO
xyJQ8u0XQH0t8hIPex1cPL/oNbesPfnm4+if7BGbLr1UT+GoEobIZOZvXv09
Z/amdgWIXCTy/yAX/7aip3kw7eORnSF40dndJCFNGVVnycDU3r4s1CRRgw9a
5LSQntzJgvDvEx/JPkyD6/wfJJtdZF9H2V40YiX1C+HJ3WKgIJzIeiNf2smX
J0XoVUaX8Lhyv8Pvuz5ZqpWyajOQPDctt85xWgK1E4MoHqEnT6iE9xqKees9
lMbYyQDkP6GfIL73hf50GyYCO9xuW5azHGizFL+uFJTt0Q6XMCg4wYZM+dGc
+3wGZBB3fNSqQ++67C2C5pRwoLJMLjjrk8IyquFThR92xFfhwxr+fPRWnTFY
I3KVYwD+1u+xho5shjoX8ATNiEtw8HZx124QM/UTSGAc28yNkdL4iemNtbu9
v33xLOIutrEg6GwePaxwSZmdNUeMO5UZNIY0j6gogSzRNrxXeJXNAmfcLhIz
DYCutdsIpVJ6BkxmywFqAGI6vSMTBda7lsRWSUMLcQXOEF8BhQOdDifVbt/G
IhE8QGnJqbeMWYThHUSTAMTxJ5KSaam6iVExOyHOAidfU8/Md7G8uaU1qbgu
CrbRMERz7lwO0TMzD/W9WtEXTiDrxGOYwV9j/9fCB5XyVp/g2C8vizeh7TJp
Cz90SvDZucDlvbxpcmaijIKdy7FaKx4ZABPTinpyfcNjV8r821GVoPuJW8wD
2LkD0wUQ5VvZ4UShQ+lkOQjhNaxMtvY43vfblGrKqbFTP8CYfVZ8zntsYHyk
8mRQqtBH38S3R6UtnyeOowKPelQjcXgm3U5qR4cnuDW7hI+fQ16KflsKikTM
a21mybVPIzmcMVItCHFhsNMA+88VcZ9xf0ID3d7eOWYo/YIG9opMjM51dGz2
6zewZlZ8UNGHFsH8S6jVnSv76XTONG6mhTsMu9CBPQxBAemqDTAKl2w/00Fc
cVc6iS0YTfuka9Zsj0xCPQA6b9giwwLhDRt0M7AybjJxyxrzquGK6qMhkLIM
kDhdi3tWPGmQq7unl8hjioC0FueStY7i04D676Pjmdk6IRpAhilAHQr9/ZNZ
cG10bnz1yHpu6iDpDjoOuP4ilAenzQjETbe/ZrMoU/48GCw+3vO8ybpww0XN
/3L6g0kAMVF7I6wra9aUWzeH9ul9yISjUn1ajVn2klq3vc15JiX4ErrqSyC7
jL5CaZL8oxeBXiwtq1yUNJLSH+offOivCGVLJWKy34ezH+vccncNSPMWnaHB
iNsxV1Z/BeEqaa9lLA7bRhCl/SEXatHVgaJjwIEmVtaPhrNAd5YfFcWqXYDg
lzamzL9WUOk8pYLjydlcKyn0a6f6nR4V4ex1Iz8BCbHywqxBfF/RdH/4SOut
Hv5ODy2UKnU8aPHRROejMR2gKC3hWtWszrY+kmflFJ6Ziq3UHO3dSDFHz2T6
eAgLGpR+smt++w5nrBMA0O3ls2s3Y19xvlKdsLkzks3kSdf5eq+sTLWS8HkI
Z9df1HfmNXeheNZ+lR2KkMv6WiPU1SRtaA5uOXDck+/tqXj5uWkEmaOd9nrl
P3McWi3Ou6uwxeFxCzvS6scGY3xhB6GA1keLVuzw0bKNO1LrnvWUwHQjGd6d
tCmiIIxCQh4IoyImJ8HS01Q+o03RLqMsxWpAw7k2J2xBhEBuluKaR85IIbQi
ettOMduVQO/3asvisUO/TGlXusO1d8o/GyY60lpIdThrjie9elNMCZuPn56I
2n0BIGme17Zj9PncZyXEzONlwobGF+o06L9TwxhO8u7QLP9Gi1wpBrTWCxkg
JY6l10mQUeTLWHtogTLyrRACGITodPwDjb0iTBrjvmt576VjPq01LTHs87YT
iCS87977MJ1RcyS1AODuMKO/pcnHk6PZF7/oIWrykpMwF7AFS8NiDK97Ag1t
gjKxxNMLRJAiZTfd1UpSd3jz76XfvGHaQ75n3mbTbsCvCFjHbDOhQRngB0r8
KqXBlYbzTcLb+E/anUKHcp49z6uLJ/v4TtnIvt9vmd/FuIuy4MLDy5V96COK
BQ5J+pudJiTkx1G2h9WHYWKSeeIcQxzpdu9yfefsagPhlvVsY6uUIT7bf5w+
NNJ0JgBMRJovCRsRpVJqzou0DO988HGoXW5heGVb0/gYfULGXvFslkoEGxUg
KChL9/5JZc0a00OAlPB2fY66ywjEqu+/9q8Uyo0LrTCYcZwRY3OWMuFwNwXJ
2fNhS0Ho6W7gUCUPoF/KwxpjczvMthxLCiw5Efs2l6PjnrM7lxCY3Ab8ZOaV
Sr/bd8Qs1RsIhQKN2rniFtfcdCB/vVu7UQJNMKaRQoPMvwbjJQF0td+JpE2O
pTdzyBLJyeCiLNQS1Zp1VcyzFIUvLCWTtH5IjZDYXnnDsl9JPnS1ypgrgRqr
5W4FpncV0n3nh+2m2ZDujNoJtoU+5KWWJc1bcGMBuYFBrzKuIpPVnXnOadtk
9NIOEvsPzVFniC3ge2BFEaj+yO323CG7q7wv44iMzFQxWuxH4ciprj7rLZlB
iA3Unk6hjB4EzcVJU809oVuzvC/hDxahKX9JmdOvR1lbEfb+Eq0=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+ErhCPKYj7L/sIHdU3rt7gGU4rckdNE2q4nN2ddnnCGmCMZNcACsgn4BFNWc1k3IlocaOQEY0C5LRDvzvN5bXNKjFfIhweYMPKTv3QF8FD+8ZkRtpYUeRnWXONlavE2tPJXcFAxs55wvgwXYmZT7CAhCGjIZeXMo1iQlDmZuzDXQSjwl8QvBY8yFlTonEyAyYm840CP0ETD6PWMGLriAG2LRcBCTOS08gbbVc1zK/zgB8+ujCcU9Y4MPVB382tTtKEjFneLEnlDKGfBS9wrUnK4Nxha3Cf1A3HeCv38MFhvxTkT+WPnH/pVKLorNQTOzmoONQ8J4U77yVityDpqqSmm1vz7W5VND+WYa3HkwNZcDA9jce8evqupTz1HzpbjJu2V1+HX6gafk1vHkya5Lq532dundaB4zpsaRIBWPAefQkAiGk3OfEzb12tD1KX2sfj05I0nQwejnIMtO4itqOiYxvjQA1rIAy7RSAowjuckEA89Ft8oqY9/RFkZz07xX6LGluS0IuTuDVa8nn6uPOTRojdDP6eMKX4FxRLy44LGZgdHjUrHqc0VVfmJGKp1XbX8ipvRtqdMR1REOx/501gtNLzIHxN5ot90WK9n/YDeQ7Hr6/7vThCyVHQbpq/da44yz6rsZbW3ffgAdbQtKtGEvkTKRHeTyNrFWKah87uA+mkHXtSlLbsd/67BvkYWd81Siv50/zkm3UkpgYEeN4EH/Su0LX4Dxv8h9bzbtp4Gt0GNLS6rHxS3Rmob7l4wyrZa0uHGopzHQIM1HuIJgoJSG"
`endif