// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WJLTCNFVz7QAi0rQG9IlErJlGAa2kNfeCl1bBNXNHdw0j1IJDachoSdrbBte
n+tzcgFONGzA3YpJpXkDdJZNxrv+QNtUjjWiFYqY0at8jwXubkB+82PfMnio
JBcAgUX1DiDz2mcXCw7eVDtEiD7rscFtWu4iOPVOWs0IxMFxYTI/SDqaYLaq
IRjPiSRTjeNICHuBd1eaQIzvKAtUPiWoqk6/mI5m6xT4Lo3ss2KXcYTl6T7j
UD8tjYCBEH20vXARzf2QnSLchhD5wSkWBS9h7Ta91gJwWPBND+Y/UQsWgAOs
t9UxLJCUTTOn3AAkEg0JgYs4u2gg2fKvCz3Zw7KTKQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HyvwqA/EWDqrYzmMIMH1puWJHvKIPwOzawJOCQLZLvTngnAJWzGfaAPeLNAt
2MsK9x+nE/45zaUIs2yrXsQkV42cYNAFmVsYJ5LJGxUTeHZDIIq/yyFE3O6u
w/r5py0WOeLb5X0WxlVqJ8KUNxB8lXAe50FrFPpD2eun+08HO4ZQ5AjTHnPd
NOBU1o99Fo3hfWT4+91cPPgPhfhwrHJYLMr0W78uKqID3/wZQ5pw3sHIP/th
Mx7f7lcXlTC74guWX4h8LMpugAB3SruwIJRnhtvDjYClW2oKDwXR2TF1Edow
ps2db8DGoCnq3BHeFoGzWPMVg9204mOwdQYXXem66w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QSh2MQ5vU5F24wd/rLjKzdPzrzmsB+Rz9Uws6j4lN2x3xOIcAzbhNg45CsPG
XhNPllPC2pIMhhGk6TM/G/81muNVA5E8QaXfbS2wMFfB9oGHJZVp7p4qD6MR
NpNz71BupGFxKyZbOxA8kb5GnwSyzygbdZH2i45rMvF+UmtkVTSLq9p0Aj2P
7geFWNObhXbUBNmqPWsTgZnIGf6PNXxsZFljYLjiZTlGrvRsxsFZFQpCVLtl
GuduQQ80onMVD71cdEFH+SJcb7c//5OZ3rRPKD2KSMqv+BUQaEkPWJvmsVP0
dUhlA8R8sez5BRE5SD+9gt3QXP0GAl9lAo3zaU4yTw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ymc0zRnEobiZ1hi5OxKZcTmrI2ZOulVyk2uEArLjsEkvj+wuqE7gdQEzyy+8
vqNHKZdAP01xkHyeqrM2Xr9dSuSOCoHz9JmF7/st1m1eFQm2zd7B3gxeGHuc
O4Um1Mtj4gYm9u6usYJw/BkTknymnj39Vlex7KxKhHloah3NmnAP+7OwckU+
qh4z5trDSqf+mE5HlOaahbowV3TYZUH3k4xwhg1n/4GHoA/XQKBL6SsSjVnN
c1+HTiD/g8bPf1VGNxpqxf7a2XAhXT3ml+yaj0UB3CpvR7sgPiLwSd9v0PMD
U+XgUQjlDWJAtuDfxT/HlvdgY6B64IXO7ilQp6dBvg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qfPouSZSrybIlhIqHoISTR9/vhm5cMHOhNBqO9g+y9QyoqMaeFa0scKzty9e
m7/Oy47Zf0+6qwoQ9UXVcnLu7gZuP5fZB0hciBAANCNPRkbfKjWPhkAHmH+x
cySWdiVIVYl7btSflhvSuXyk7EwbcyiNK8H3UGB6Om2G82KjTNM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Hkf3/l+PxUtNCzmIEMcKv2B5pP4VR9oe++mRVbIP2wmkaFjfGhNl91V37MIX
wJS+OO4BoYXJvn4oKReW0XH9/zRkdm5KDVLD7wQNEIwui7Db8bT0EVrwHwv6
vFoJ51p6YYebAqWD9FtwX/6awHPcWGNyVud+mjJfRbjfoGWr1CaVT6GcfE24
fGvm4oARRrnc8uz/rXcbAo3pNhuRpDs2ia3fZOltquKzGX+H0tq8MzwnLDgO
muScjAxs0KC5wilqupgVXiP1vxpgAtmaTHNf1XCBJd8Cg59IkPhCO4wYfWVS
Uly7T2d7Yt2yzKrywy7x4A7L5JaCXKc79ETif3eOlBXzuPdXKsvO6YIgD1GI
8usb8ATuXLYBgUIacNwbFvU+23Shmtp3om8N+IeGAQ6MRdG32cgB+DJfQ+7v
Lfo8wlLM8Tb8vYx22kC3K5kH6XTLoMOcw041PM4s7wipP/pKTfQwAcJ7wQVt
yWGZJ/qf+YlqLiXzYQpxgsJzbspzkeao


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QIJWFaYgzGaguAmZ1z7l4G9D5GqWhOlgBx5o9k5dzs4hZgI6lHtuyqvGlnhU
Mm+q9/l5Sg4uDAM3WhEJ4Tk45imrRLXaMr3Z4/gVzHjea25arvwsqPTR95lk
WfNipwONUTUmQf/Q1QE0glVK9BHaBwOB7+Ge/ybanE9Atrac8fI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r7dui3ADe7MjQKjPfu9xR0YRr17f9yekY8dcXjdzMphT0EYi4O9CTgjPHagP
OzLREPqB7MVHTNVSRTPo1r3kqJKhyjPRCtmQUaGRjtRUnNiJZIXnxgLg15Qm
BenL+FiwKVkHKUtY2+uGG7vOsIiKe1v7ZjGMtx1psATId74jkrg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1392)
`pragma protect data_block
XmkizTF/oVH8/zbEOqMmS5Le0p3WSsaCRg4ocb2iAuaPCNgBK5VHWV4dW0bL
8+smpWgDrb/ZWVgYQurWMfv0bGBf/ZgEu2ExAbJREXLLCvaqVzga0hNwElIW
gn3mFdnawR8di8LcVlbNTIcE34+vKmTtUCErAgpbUVh4gEkNPQ0F2OzXpMYo
iL6FqtsY5NB8LZRqxahQgpd+WEFwo3c7o7F4T3RErYrDIQiIaCRDNK7m2LTN
EtKSNRiuxSv5S8K7s0iNFOI2cz7CrzYTeCwB/CBxXExH7gyRw6jOKKl9FFgC
TOCrnWcCk5b72u5daVkUXfXFiSSShi2GOWILFX0yBbqx68ZFjBzfduzpO+k+
S7EbjwOfZXIACZy9nTiPWyttPWqWG/rxKEgFW9fIzzlwmEAh8j1JCZpkGQ5+
GZxfsAeI9ZVMASOHX9jtsjI5GdkpP0K9IFR+1aTk9Hecv7DeajbxpCA/jQgI
vm3RdcAEeMHz3lUC4vu/gkEWiwGsFzMeM6w08DFBx1+uzxZa+Q4ARrFJdDdH
SLDlVf5pL2dGqWOyMUzYbZ/kCLq6MchCNGgLbDvZfZu9NXgtKDJDSH2iXFtL
HW8CBFlwqeNJVMMRUiksP/iV8uLuqnoPBOce3vazl1ogJ5nNwDEmkqfNs8Te
BBLViazL7FS6BLek+tSAPwZuoNnH56xhmjSXObpC45XLuTji+BUHePE+xviD
xK+awqU+JuYNo4uy/rgNDS3emEizUSv2BuAIkMk7oPi5mICr9FQf1TUBFKQR
SaU32XlSGy36BNXXpQV+gqKcTClie9H153xoPYnBBZ3MgJkJ5oujB4dRUz/K
ZBYaW2rPxegZ7UYZC4ePOTRuZEv4/3LjMZoJhK61l9l/S7iEEAYjx8+TaRXw
8tfaTTSZXDm7mEFiN+CzJILeIYw0svtPTfqIbM8f/KTRIl2aaMkSGuAD2rlO
gWOsxsmHE8C3/xqTPH3+VeiX9JJRpER0wS5nREGNR7WqZv9QUTwQObtKPNMM
4L6bYf+dtx0vW2DE6FhP8evx819N1xPUWaAResdHivV7TXtTZZlDMvZn4lgY
CGNOkKwb+qk1Gq2Gp2EK01l0yelJ4Dc4OjcES1xTYfvw2L1iXBrv5fobTUXM
Sf1f/hJi+PcqoEJAwNv1mx7neLWkQ0nT86dQHhX6W5qjUfIm7F60+lWkaIIX
5AyVUHB+Ab6P1XoH04zNYcF6yFjPtnm0MFkFBc0mcX9m1R5pcKbN5ZXx8Ldw
401eBtDo7dH1Cij7s6Od2rXAYfwz3LQ/iXuW8/t80UiHYiGvK6vKWebfW5NJ
W+tK1VHbumEqB4UHq8T4teY3bV+ysY8BKHbxDPA0ROzxpyj/FaRK+VoUvXXo
lKGRGRmiMs9p++GTUtgsY9b6hCxCj0KCLPi3Ic+h7vnIvfvZJI612zaB9J9e
EGxYftpO3FCcVHOE84fy8UcKP1lwib4tWWeOCQJA+zFn3Ae3G2tR8FDmzEw1
IOO/pej2y4s9mTLb5uN6GghafYOH4XDQVDYiJ+q/i9fTwWbaBXLJ4pvePwEb
dr6GVN//1Mr4YK4AOORrLNKekFzXTKt0YGDs9F9woieGMDay59Ojt6C9u541
9zmW62VoXAXySYjgfGkiyens4ppdrx0h4q5trA0HKa7hGQWIz1vPS/ZDZiEQ
sp60MQB9SXGFzLKPIfT3eKaGMKED5zPgdEd8J2iVcpUNYIJCgPs7i9Ef2rM2
0Pt4+JVaFU1KzXvmfriP7TNflcJfFnIorAo4ecx/v7cEL+qPa3rzG8xBkzYf
geDzuH0yanzRGHnoO8rYv4kkcIj7oxvQVvBsx1RpNr4ZCeAfok6UiR31

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqeyltaEMPbIg+h0RRoODBS3wosh+stF4U72ri/aplFYZzVQiqtud8nHG5XsdqycdIjwodF4DBF7bBHPVpYfN2sCQRxd+ZNw3zVxUREVYxep29DlmEErmqUpsj1ClpX6AJPSW6r6PmZNvIqpod+sqP4QcDdBjAcVoKjt4UGDQ4imHeiSHA85rU0cNDp+np2QMepDDQzSXbtLnr3Qva4JC8IAFrL/D50izoXFY3oDpxE5eRHisGC07wUmb47LYJXEYWDrS6KqPavmMHRaSsQ+5BBUvoqswv2VI9pHGyNTIUkJ1f/P7jafuZ8+s9v3EUEt3Yx2AD2q1hHdfh5Kz3Olq62DCFHVL+ikKLSSM/QmFYe7kbyRDcCZi1Pw3nzWLr3mzz4gHYYemosSuBRE6hOgQK5CaIUF1qcNKILAEyGrTbMLTOKKfn0QmNkANDjmlgUzilv/yhAbzZCoI1IT2iupJfBOzJYgJHBppLFFeiT/oQcWv7QREVavfr2QwH4k9RG7aDX+gGVRNHKyV2ILxVYnhRG+NVuw6UyB7WUCpgEFRsPvk4nl7JjHqprfmBRUAfci9i3qPgG+LVIkaX4dVFpXXY3L3snNXyYAvxKMBQ/XZEnpKkKJvr7UUYT67wKeSAh8Vm/g8JXeU9oxaQG65gv8VmmlqQGKUMcHwMRJuntZ5MzOqnP8xVHsVEFO56kftep5WiXaJmTWrJiQRK+RJ9UDI3BevsZ2JEJhEYLpgbS+wO7RrvDDFK6YjwtlkakSg/hRQ8VsuRNTxGL6xWsQeg1NtxZn"
`endif