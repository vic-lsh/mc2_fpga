// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bR6HdCY6fsWrQe3pCKNSjRdWIvq8vJfnqu2T3STMSwCKTTUKFpz1u3GAhMhi
HoHNyM1agmcjshU+xY0mrscrCK74BmJ3yrwwBcmIDOv6fv5Jri3EaUVbM0ol
jlT5/KwS+aY+M6CbJpQE4DC4o4Mjvu3HgaU3BFCeSKZNTIpuJnerBBKQTIaT
KfvBYscpJLLDPqyYv/dX5tN68uV4EGhKy3rPSCPMzNoAMoME4qVjO1SOOeNR
uD2qy383wP/ABBN4Gxhgje3psibr7kR3iUznssujRSBnJYPEtRa2S9aJKR5o
eaSt7F9kQ364vsF7ozlIlPTjZ2AYLR6AJIX/ybr6dQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CNH7TNKWHq8QoCzZE11xPOrCxCRuilkycQMk8dzfhZv/d8k8RGsBJ8JtVYjA
yyzldXi+s6rEnstHzjRtQfLn4ZCK3dqB/jslmPIrIPgR9oppV0jzBPDPt/1l
6UTi74uXfoy50V/hI5guhBaQGzixmWspjelmPDYzPWH0AoG8a/Y24zRYjjcx
GOruTfw8EjFbxcGg6em/QVcvM9pTM2/MUmV9erUjzXaf8ed7BjJ5I+DMo19N
/3SO5iIFdMrL8nyIngU9fd2ZQUu77ioI5UKqYomi30pcN/3F8mM9PeoaREnE
mwEq6Y4Iv8KUk98pgVdue4MkEg7TzLCNB3PphRI1lA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UylpNW7d/aDRbqS+KlG08M5L6qYG0mdNxm1RCfh3KQ4ruywr2SfApinj0vuC
L4N5tK4B6H+wdrx0aRmd7bB0J+IwomP33He/GYbl0nL/5Kp9BHH33YsMpPl/
xrndxD1J0RYqp04xmy6w1IcqhMykflA1bsY9bwGkaRRBbHUc4E5qCb0YPT5T
GF+cPedoDrn4mKklWH46jFfT/FpsyRas0bAxIhojzQNpz/dMSnT8TY99Jl2w
zi/sowUMffCpkI70sXburPNos/Zd9T747nf1uY9nRMjSO8iD31xFedTn+HGF
HOcfQydLTi+1+ulDxz55hfssyPbrnYRTNNRqjYt3Gw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Hz40a10IQsxvp22A9TIkJq5tuaqSisxaTa162vt+3Lu+8WRtcgwqNMCYCKQ0
s951ueNctQOvRIH9TC+z/iwCHplRI+nBof8Rbjb7x+lMUvdcMOQDuUTHMraM
+eRcBL3QpGNNzYrjtJ9feedZR+4FjPCMFQnxNZMdX8HlBx5RX9Ot69WYQlX0
SYD8jJdDFbeHvm81b7gwxPdT8gntWWJBBAaBq2Q89ZSIo89DuNJrnlbPR+ir
tuLQ1qqsjmJpyDdJWCqDd6wpstaq3a1/Vad6R9keLQjb8sCVQirXV4wgIsqQ
ymThPiXwh3QHgNdC3oeuMpBPDiLyEsWgUJRVow1Sww==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OyDt94ECj5emYMB/veNOSakRlgF5wk3XbQ7bycBG0sfCaa2orxyjPXPqX9RK
kOt+fzd9VGCVG4DJ4fHj7ex26fkn6H4HTH1EMiRkhnkqhS8IZmYQiqBtcmGi
nFByc453vD9TOuTqM3b0K48c6RwgPC5A+a7h9iYtg0qKrRYKWXQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Sk/WG7vCvXlAUyrYUlw69aFGezeyAy0zwaSStr8coIjL6xZRq9vHUvR9Tq0r
+Uu6i6mj8OCFHvoGUitGOHAOZrbwSZKSZeRj6YE7sKFaYiP1vxJVZETRZQga
H+WNWgOw2a5Pn0i/OvlS2/r8N7ngJNy54psYdsryAPyNA2glqLYXDAYFVKwt
6mXjQ/14jfEuixiXXoGvjqcCLPx4oZIWGMg6jE2Dq4RcikuScX2Vbaa9+LXk
P5aTCPe06CNS8qjKfoyuF/mosIBDl6sSQsw2itPc+6dq1sCGG6B0oRT0SzsL
gKClew9DSGtMi+HdesxdFd8zfiEKsdv1Ks0z+9rZDaqptQw0WoM6ByjzlqK2
EpBcDIOcCgbSeEap5zmhKsN/CYmTn0+cm9HgIpqEFLK7m1Xk/qxQKfkV/r7j
gmkqZ0GMU0iEEETzQ813utMHbyrQ0G4jKZz5/jzX1HFxdBAEJzhBiSfGDRj8
A81b13J+tCU9p85PI37ayjGNQYfSM4qe


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NjvkQAeHVEOoaev8oKPWs69EsPCkd4/eRgONKIlI11TIM4soifnylPw4yKEt
KVZuNNwNvzm8VuOL07kQK89EHAIdnB/K5kMBC1QOvXDbW4QMc/DasPyLCMrm
albpfMn7QlwH9ormuZo5my/C30cvTCocYEmZ8Tp3ZHT4rBblOEY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oHQO0wNdzL0gTug5DZWU+3jAjCWd/8ns6t/ZBS9sHNZgCJ42ICkSp5ngB+ir
44weklK/xkuqU0hDfsKQcY0tdUhyPjF+pFwsdH3oCIYZDRQxTLg5uDiXc/Wk
sFJYh+/sV7GbrQBC8Bob7rWqCZ1o5yrFbDQVQ8S5O4Pnpul5gfA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 106288)
`pragma protect data_block
CG0maTuskMOs95ZQpyHqptpdSzNVO5K6D7AZ4JgxMhW0p6H6VryQ2zWZOYsl
RxcAY1qSIKD8VQodEb0ek3NnQRjw26WtZfmVJpu4wStSi8c7D2MV6FWvhasK
1x9W+5AscdwyaB/u3etHeVWfg5sOw9fPpa8L1wiQXDSXi9NX2EP6U/G7y+On
1BbO5MOyVUaEi75EJcuiRnP5mlKnbOOn2W4oAd5Puw4F//SDeD13PNAg1wd7
ZkBGpaT4YDnzyp3hZRTCbSB0GBNO4KcxUmDEPMmiE9NC5jpL4FWKhOAumC9R
tf1j5bvqLPqpZMJFTevLcicPi0WxxZBeu7mvz71J4xwJ1okbzhw0jHQB/5lp
USDH5sdEGotCSo/oX+pncoWzxbKSbac8mtD3jzZNZYbIWq/euj9jLCuXpCXh
Hz4jl5XiymOYIEqGEoUdbgO3Wxi9rvlPEAjST0yUQiHCxU0UxeoDmqnZ8zGh
aZJSZOA2hH/oC9BsYj5ZyRkYX569JoiAYAOWC73IfwWDxo+VRFkCdnHm6Jmj
vqcjK2+Bt2bEKTNsGjUTnUFA8L9mJUnUrUH643n+MHKzfBbDmKWGXBt7w+iy
iAYLX59dzPVIEan+VSCbhr+S+LpT34W770iJ5YWgx8XTAsAyDHOlwWPu6AWy
MRicg3XcSlkJkn3EhKZZblz8IINo/M0rgN6cM9YkK/keI+klCxbgmn+gipax
glDrq9L9X/kr3MZ2LYNT36/UtX0UQRwD54zH6IZ0G4EJon1FwVYBvGHpN3Ae
5rl0wY38AE02/BRivWocb6sOL13sA4HFJMVB/U20prv9/M5LRuBvjCzTSgK/
wpFKIwq/4VhLN4eRvaCtUxJGQR4tIkbeeAWFGbeGtRVp/8grdPZHom6tM+3b
v+uWVP8qsabt1gmCovq+6IEc6n3qIbmSyLs7lQUOq0VYf2xk2JWFATd0o4gt
uxq6PiYUTfW10d5tOoz22wjB9lPds/AWHH3oRtXmqisBSL0iBNuZDOezWPUI
xFQd/uEACNimYmI+FrGJrJmZeSavRGQwoD4nbA9rUSVDdp+AqIXR+DCWpyWR
AigmE84lmEu+Ig20J8nrLKDI50aJFw7i5vKhA60PH92jY+QnCYIFDIrEsoPH
9yxls16maOUa5Dg4xKIbuLv8fZb4U9EbpfSXQyEE7lTiS/SUhlUDU2eGpq0o
uhqBWsg+P7LrkRqwUm+1nqTKZ1wUj4qNzw/OifNRhi5umsBVC3dl6KuyXVod
uUJElFF4mwbC7HGCSa785nIxhz1rMq4bEv2EQZ6L0yTdEN1N/IsDp2OlifML
hfob3O8M7c8SocUefHx1e9DyrA2PTbzUXDXYTsHmMwBFuuCWIWPHPco/Kemf
pOmCYNz5LwLd8oHfzdNhnYk/XNDs+5xTcRbVZAjy1neWSuo2nneOayE01r7J
V9DhvVkUBnDWhG63Vjrtm9KKZSKvpNwt9PYEChbfiSvhUTv/Qwhk66QYyuzg
3U8FRuqsbAvAy/WqiW1iDlc3AYIQisubSSH1ENJsaBB6L62vGzM03xDc6JO+
jbA8mjhnzr0DewIzZqpHpY1zn4KZZkXPzaS6g3RkJRFd/r0QKGLL5kNidQcJ
Nejg0yYdsDze6/xzfttveX0fwLOX7i2XvJVW8PxtPP/CQClhNLIhDkNXpEbK
gsT73DJpqfFaiIzo19CrmYVzjCKs11c8wNdj9q0rsJangLqdJcy96jBzJs7/
1HoPg/bj5Wi9R54YTT8N5OBb7qbpfzxh4mw0uyK40HQdY8jr8wSUSdFP69rs
vocG+AdzlHqPVJwDz+4kbKuvdTF8TPZDKx1MOlLADtsOsV9kr4Vw4UDoT+zv
ctabqBbNiv6irLjAYs6Whi8Mb51m+UdyH7tU0rBJN74aIgw8sSAYCRxNBlWO
V3aamkDRVYQC/GZCtHhDk59Crl1n/bDZyC5tvL8IK65wx+iQcXnUMJv7js4X
BlieNdCWiR4NI3T9+RMqNP2tZUljO9fBrEUg0374AeJ5Zxpv9ND+TChcM4V2
IB4bU1kU3ZRi29JPqH2klbynUU0Ox2odI7Kt0HnZoHTWOuBC6Dbm4dK0QpwI
MBvcWh4uGK/fV8v7VFJcLGaEbYRfRcKmMy9eCadGbYY4jl/pUY4t0ei8Emeo
1rcc2WnKa3smVjYbMd7PzKRxiDuClQmtsX6aDEVblNS6gOO3L+MzYMas710r
7vxmRwnsY2yxYDT48dt/pUCwKrEJVRpa9KCiLh3wZhYqOkZfWJ4GZFaR6A3s
ipVdkPOqEqcLGk8+sbVO9jA9USqIzrUTODM+x9oqgvB2D1td1AExB9a8HN0z
UT2h0AxoBhbZWFuBlCbahAuoLEMGTD+AC8GgbD4HeOMD7srz+30aBlfPD676
KP2qwTA+Ajvna7ZNZE64Cvb9nzv1vgpQhg88FdvgihNzJFri0cHdanct4OYu
jx8PZPP7Z4GYlNhQT7QNKvfgLcPcuXJ9RpJlP5jpBUFK4IA48sQB5Pmaer/k
LSm1yaCXdpc6l6Do9LB5i3NKGApMPRMZu5ruhSzyZm9ABHWlQBK5skWY/aPf
zOJmgRkKKFYzZLuW7AFd4LyEDCpSxlPRSs89FFHkEepYPA+oE4tqqq/uJX2m
yQqXzMj9wErDqDo8Z0subvmunRKbYPHanREecMmJm/TqeGh0g330eJPMU0d3
QC4ZAvXoo+ChPKkgK3hZEC4mH7VPhxQPeriPiZIVqKVzAQkFNjHsg54hfIN/
2vCZuCbYN4lVeKRv2aiFak6MhqV9RejKpdnwVGWTuULd/Y62dz96rtGWfRFh
mqa2Akg+Q+wLUkySdz2Y8dw8gaLN+27JiBJ2KFS3A0m4TzElpUPHE+Kt2sN+
sWdl78JcOd42NqihX2ulyCNyv/u/D1QZm9IComXh4+64PgigjkE9rYiuecjM
F0wafAVskdN+/WP0xjVKMBv58hKS7tR03C3AYfspMMdYy6TeOixKXUD4wvA/
zgd0kQcYX8vw6uaEPUXiqI/Y09WWK1jXCijpmledb3uzLuYEpQUxYYWv1zZ/
oyDhiXsW2dFeFBp1M8ZjEBxxcAmlGHShaIaVEO+G2ONUaDNBVV87rIu3wOMf
SlUxjMG6v2dVd5i1zPOUET4jeLDSsNC8bS/AFuKQhq5Z2E+lpLJ6/pxbrbJA
ZQ70LzZYMv6BzVaLiuB3kRYqqcGm8iBdgtiuGNZjkmNvV+QxBZOGnd4kFfIp
ENe4gqnAJ48JRXrP6XWyKMQdn4u1mftCAd/0br6o0/t7MUQ/7NW8/fpi5k9N
KLHESmxIHD9EekIzs3e4SbOrg7D7UVRQfGqsikKQZDFXcT6fzeKWnmt3W6/+
Je+ocqcYeOGi9xCU06Tw/PAjBP9cj43IoPq+6U5C7hIJjqFdJwb9kEqhCXzy
6FFY5kmE/QiB1pMEMvqTQ7Y8SvqZ2rTDPK+r70wCMpLcH1kSGjN/szCmOX6k
8DR6S7JHR4MTnafowYRFYqiSvhpwKBEhEf7XpS7c+Y9pejHGnvcKFjC3PD0j
3jugC0uj0J38SHx6dcNLZfRRXxFPc6JK38v6MPq5hUJ/yVfNAauPKv7a6qNf
JfsMQvMXT44q2IqjBqte02CyKZpRtetS4H2M73s/6JPqC6JydlGpxKg9AxWU
Smzmra7mkqWIw4g7rqLCpKG9voVmCJ9K3errRwmjrLljrrCyjS9uogw7IklW
Z5/CS2NVBNrycKc+YaT67l2t5WcGlxi+PLfcGkGCm4Md/FltmyDG/YnZlIKR
IfSTPMORCUebjut2zwdXXamdPaKfg1/xtpKkFt9ObLZS8hB/CPNtu4slvedD
eA5LL7sh/3kRu9KF+h9uipqZFyPSJwictWTFJPrYHrXbnQ4MrljKJ9mu8rjS
IVARLDUywUZFhwFKgrC/RRRwuZDeGUCZ/bm2cYJqCbF0KEZuWz70HXP+/rda
HOYOPmefHvXWXMUGALFSbu5GLZnffDO3U4b1Aak2MJwpi282e3+gMwvaTFE6
9jyIZjgnkZSjjNbEL8aqy3dWYQ+/XEnfx4oR1zVl7FkSy+TJKENWvg7n4kPG
SYIN4jpZ+NIdYEjzI1nXuxm7JfKCmTF9LTkhphAzPh8SUyWCIaYVAPdyV8In
lsDO/ibTPMoNkEhgZYOYuPPL/q4yWqNeghJB8PvaxymKZShseylEVElykFEz
Ru7mtk6gGNW2qAthQzQ+3tTleRgL7FA8pqSBM5bC+xUJrkyRyLyybpd5zI1L
R/OZIezcuPxcOH4x+b1/gSAv5QHz79As+MiojqNVOU1JUsOW6mGHCFKJV33g
rz3+pOkeQ6ku0k4KaSrqJVkoAaIrXdC4UZAgYcQ1fWz1nGbJ61JwWrzS/Rps
tWWVMeaT55GxMxKQsbYfSzN9QBTRzIzuVFTdxbmfrt0HUHuBKxIHR7BG1mIl
pVaeP9l08EN4fVp4MsVqHLv/SsxwslgPAkPLo0wDKUL2LhqrYGnFN24CXD0j
n094Mfp7NRgfJ2EpNpe9oY8emXQze6+BnaPWUrYaTqc94fzlEjaAiFNUZMjs
SFIt14ET3xXyHn107PWgKtiTJBmY444v3HCd5LESS1Iqc0XjHIDAC3B8GV4A
hbUy9KcjeelBoI5bEAPAoVnjoynIJqyFWIpHPI6gSNRoCvpXNQiI1shKqTP/
qqbMRsvd7ZJ07X8xr1o3yv20+pTvpexwLevX1ogpxKiZRNL2UgpAhP/wPWsw
bcclFz6Ykc/tUX5xjW2Jwyd5yvz9zJrPLmZZC+8fcggYaQwwCNCnmBD2EOEr
MZ2gXMuGosh5GZhzJm/Vi935FzOzAhdNL5iaSwyKLV4ux2A1B10pY+LvAD8I
UmHp+Bk76k6X+8nbVuv4xTgAMSnHXgF6oCN+CXis3XuZQpNGxWcJhqJkxu7O
TosQGriGisjnVpI5mXcUuZx6FutFxYrUKTKL5Z1IyYJTuzpV8kTnhwJgpWgx
pt+8Qj9YTD9DxwuIY16BvkPkDrIrvwP85Su+x/AQLe4zD7LPbgydUFjJI6pj
lYmDZPZOsqYphKTihmiyXf9H4t696JcOmqs6hSiXoRraE5mbsfmondvCrPC0
hRAtADM/GL8+cEGji1mJV7mEfyE53ZNXIivwsfUBBBEgCNKLFupKzl+f70zC
M7OWL4zYYfQcxrhHQRYXA6duxHIgKxGq62xNaMPKMeVEimSz95ABKB5i8aWJ
EAZyvj3KHAJrKOsm3lBnLqxGenwPX/e5bIENK8HNhGZOWcsvjzlOcVAGEkwD
ZBXHk0KDU97OSg8Eh0XcM5ZQ7C7ODaLbkzdGCgVYqB9DVk8L5IkEo5mjJ7Gm
nssUD+wqGOX3XhT6XoWvYbpRUMEmdLEL63G/i/AgS5OVld+4IucsgxECChX+
nQrK+Lh0LCr5wMBp1mN4/4oPQ28P4pdjCaHrDmkGlri+0XXMBMEzNoaTL4gV
eQCTSrp8IKKSM+F9+JwB1dVz+ES4EOu4XMMrLisv39H3sFIjGijhyGxpWSuy
yoOt96CrXWlm9f2IrREuXUlZv0zC5kUVr68Qb5lb0Sv2B7NNHKx3eFO1HaQb
zH5Ex6RZ5dbCp00CZMn4KRe0PV6rJtNFvCqkxBpmVOHvO9vQMRuVu/oXESfa
MwZkT0y4IWj2n782nbgv/edY1Y8dfE4ceDEVQFCtbtZvOcSVRb8vzmEjpDyF
8oQGnDxiYJVl6ylv9SUDPCVvlR/EI6SPJmLm5FohiMATo4JEVgjSgTPserK0
ZDAbq75jwCudY44A5erNFXuNI1W9i4sJQSuFdftH5lj9wpS5XleCi7mu3AAo
Y+JB3aL0xeMccskBfRMpdF7RIkjATYaVRiK3R9wn+r279ySivZrg4kPVV+qE
knvYnFEkE3CIdP5zwaB7r+Cn1zNKIH973cUerQJGd5yppqaSHac9LG0ZQBL4
Jz/nvr7F/Z9LuW+6/UNqbl4KpBrVx0/Vh7cDsMvKMLNg5E4EWTa4/9+nEpFX
/dvqP07ucGV0G5Pv0Cii8X1oIMGKO6aTnaiLRQeJKhoo7puMSNmqETBbbWCH
w6mv38fMvZ2z0UTWkymrc9aVeibU6CFSLKi0WQYUbfzEUGPJLHdNOWHWXzuj
VYpeKOJVYvyLcBLwyomGnQEqL+M/jl0tflvA8P3RP3SMtgyqEIjTaDhx17TW
oBOFabpHgtm5tnb+xMFnBNZbkltHit6bAhX9UgGiFylJ9xSpIOjzqXnsBzCd
pshbY2KNJqhQIfa8Phs1KB9uNMwjKWjGoJ8BQfseh7FoAMyEK7wrKDhTrzuf
foamvbqOBqS5yanti3zFsZGk1TSDj5xtxjoA6aDv1+qMdkZ+wA4eP8q51ogz
N838YBgk6tzgOKOVSnvQJeB6oYtsPqCCCEgmwpAuDBMPSjXXT4bvA3glpdFG
Trac75xoUJJ2AWDM2HkQ/K7i3fV9uSnLr6gopBLUtR5pTXENaO38TOYB65oz
GaitoA16i2arPHvM/7XGv++58OCUJmy/v+Tz8NUA8gaP08hmaN7UGlAmP86w
+C56pILkp3efFaoffETPuLaHR62ttRo7Fc4bhaTd6LAwqQlAxcnvshNvVvQQ
nSLWVE+jWufVRMwoJJGReYfmRzbw5U8G1vDEu8guh/g0Tchbzl9vg2OkADy0
g58gtMcNAAigO/Ritr/5IKrlHA0AFQG0FPia5kbe1ehkdvgewhU2neMIm6kc
AA+doA6x6XJvKtR36V+BArW6ldyr/QmB04/aUBl2xFbnPoLlEvhisw6C8OHY
hw1rFDqpVa0NLqVlHZ7Kg4Ir1ETI8mRkkuJDVbde04wt1rara9sUgcPWur5I
3yOxdzr6Q4J9RiRX3wutewQfvEsHtfnaXpZ82lNzy0LUCJcfNu1DywPKvXlY
RI60ISIlSd2efrRB8sU6SaqWCapYRtpTNZlH8igLJofsDHM/jiGbSLFCWVnt
1xZ+NmPmOFqyvrTtaY+5y+HUeL02XdgD5nQy1eEtq5ML5wYrURkx2sOKV8R3
S/jcJqnCJqkAiP1JXT4IfEeA0LXRQXzPBqFsanJjxIvESdy71co6DsrmZg8l
JyJm9r1GcaHpiPOGyi9rJyq2UJ75y32IN1q2WqqKxRe/2xtfA8m4Xm3R4mMa
ey3shc3h++nQcPptaUV7k4+QMfBdHiWY2PwojE4V2Abezw8JJcR15ZG2offW
wpD1l/ac+O5p4fvQHbIkom1VGXEtSrswN1CiRwcKaZ8radNJBY863HrMzkxS
YEEr+M9J4RABi/FaMVEK85JYOUggnCSO7rGIKXMOU974tULOZcF6scTPbnam
vyo+SstNu7JmPvOgq2hzBJwvwGpNBjIRYWez6aZYhwTvxEzkQdrxd4xOr8MP
/atZVFaug/a0eeXl//4zR5fmWyCqCmoNHV7Jrol5JmAtDbCjiMqw+/DJnFZm
D+/36JEoDGQD4XHiF0qzq5Qt38LJHJICRi4wwB5GZLEeCNAEFRY5KnYghjVG
uao6kIy9S8KTtDvKuEn7zcHG1ciu7CiMlTPHfwYtdFPTrUAIYdCz9oVJdzu6
UieP87RCgfk6ecgbzeakdZcE6F8QaDX5C2fqcj79itWYktCEdrC3AumprQSQ
htY6AMPYzpiVceWi3lfhpteWXwgKlSNZrt86VF514wIn3f+N3e74eif0mLHn
5fy3xQyGQFDUQ4+A0zkPrU/jfH6ZhGAJN1sSKZrJ0iO0y5vbGtJ5GSGyx3E9
QJka4n/e+jKsvWRrfygHvJRnbsXJnYLe4SD10K9DUzTsW9mLW1z3Ls43MKyb
/A9Z3Kh13X47EVZEl4Eb3Wco2hMmNI3GKwpNOiR4PrfXIVhrWZ9nlPsIl0Ar
2SbYa/zsNLD0bVjhYJXYErzCL9k512dvROcg4Y/co9/CgZ+Imqk5qqCrwaRq
VWt3AGqrO8Rkt8GE+07hNbIjYiV++YIq6lf0CVaop55lJSaIYbbUM6Ty4ATI
SA4HDnNUWyeQfzqZn2/Dd4+GPsngunK/vBljGQB7827glxXvGw75+u/1oqFy
oZmXXoplkqGj+FOFXxpcqZ5W7PQIbTvnOH6zKPs8dcZBOrnvj/Ot5vCe1XS8
fNQ+NFBJzPWMV1uHRqcmEZ32bJKiyF2Go+eCmb+vfA5B3h3rKu0geCLyE+a2
Z3j4SRPKLSGdpT/Mpevusl+AMgTuDCo51jFSIqIQW2KemgaR2R+sIeC8Lq5s
s2qVJj9n6spy4DA/V3Pgn0EITCE9EpTmUIQT4E1KYhu8atICanElJrLUpt/M
qqCQqRHUQQ9/xwiopKXGkvhabTLFHyt7wpNxPZKwsxvOeP7l3UgID3ONdyiL
uM/Cq/gp5vorWsXebYh1EU154dWL0F0Uh2ck12YRv3TXrUq2azgoBxqG6r+S
/2ugIpi4/kKIeGvaRlt0xea0WH1vH326Xm/Kn2UD//bOQhLXDEC401afTWTn
cXUle4vn+Fzne4+4Kc7wWa+3jPFMYaUUKLIBYFD5J/J3C94S7WB7HqKYOLD0
rEI648206/2tpYzXa+vYN9dnJWzTv0yTwAwqMuvWgypW87Qu/A3sqyTP3OTf
Kx/nwsWCW9Nm9z5GyP6QV+M3VTXtkabQjgb6xZp6jnpmTDd39wONoBZ49By6
LRiSVhVOcNkLFVrMASkdaeq3UnwZ934Y6HGSjK2c5fA1nhA3Lab+Wox0MBuU
1QUnZV5+k9Jd+FXAuIlJ93C8975yYsHtew4J8bmwiVWtqCddXbKFRzRH9QN8
8IR8ulHW1twrqK/5cN16O3rbzLgjMqDa8jq7dkS1rz6KPhDafMSzPWAue3ut
XB7z6SOOSJjsPCxEOWrXL9NyzberBtW9H2cdyca99hM0paqc4QQxeJdbceOE
h1j1dg0wnWAVIh1tX4sEl+hiRG9T/poVcNZ+Pzb/Z23IKh1BeAlKhyKCQS47
LHopBFQtypOfZS5N0tBw21TGDM48UTIOMg60xQCnTekHMX9KZGtlUF4J4thG
HAAtPZqAm5uCUx8u/at2T5wZOtRjRQ4wATqgApBpphlhU7J3algt8v+WpxkK
wLQZ6KC+jtnbRE2Ly0WKX5WM109xzhXB6Uxe9uuDajlw1WUqQQpvQvKndoVk
eHdrSJV8o2AgKcnl9NhFHAAssZMpLTENAtj+5HwjFzAxzV0ZGsj64yEsfQPC
Q5DQGiaxiG8OFndydpzP1VUIFqhOP/XUOPvq3uaV34g3JT35+dzX5rzU3are
0+ng6aWoYDKOpf+hBmqRjh/xN5QPnA/Q6uq5GLuZPA0kblUsbJ1RuK21z8KS
vA1jQLmd1k3x60eFqiSIEwXTnbWVaxovOkVXolbmQ3PplcJGnvV82i/H0KrD
P6ufLqxJ5+zYxUS24PuSrU78lmbj5uatjmnvBfPxhKodp9gwMYBp5bau4eVe
z6jd3gexJyiw71krOn7pLbpbLrUu9P3V/3L9sn73B8NbWVBXzCqKoSjczhoO
gaeiMrLrLxaysFXLhkpHFZopekHGHWb90zbB5doLH6z0sVxn4xuoHape1+KU
LI8/e+7qBCpcS0yFO5tGK8ZxadfZ2qcrtTaZS3q6dITtvN3MdL9pZ3Ab3XF0
QWC+s1c42/HaqOP13G/hBF4CaL4pmGt6y+UuQcexycExJT0NGrW2ulUFzW69
iOhvXDyAhPfrfgqVyU/hT7hlXc+B/WEI6rvI+WIp+KwaxT/R7rx/7M5getiP
GjWWEgZDSV71vX5XD9tfn1/N9/Ftg/Zs1K8Hk8RdtTWWRsRLJHDxeF1ARog/
SrLuJFe8IZlwQFcSg7h98OvhJcm0kNfJyEQ21+RwyLJzPv/9gHObCJi/r9dP
D+nXlgL4+N7o93Mz3uf8HMNXQY5F9AIiphHhwLvogQyfEFNVeZLhf6jgrVVE
h3aVB+oCY9RvwzQ+MvDk/Vja/Eh1I+bI5bx6FI0DGZkve4hl1o5Tm+PbUSt+
muTQr852Sk7tTJPNrEYNuZKDhRu1AsnPmqHWfdg1mYZ0IsVXHt+OiMM/tIWp
8QskhzBxWKJkcIwwuQP5waLzb8TJchLlKiNFoJQ8NkFgH8U5UfBwbW1RKmNT
IjiAWFMHjsuA13qXS/udBOBq4cAQ746iEpgdAebjGpH7dunG2wD2eDpIe6Bl
9jzceg3itTKdcXC6AJtrtRdycJ5+6r0vZ83esnYayO3Pw+6d77Pc9CZYYldC
B/oNqJ1MGVZIp7bp+eUVpu3PHlaD56YXtuZw0aQ9xdDSblFEhkIwfc9UkBSs
yqFa/PUYYKwTM9myDR14SDvEvmRyJ8VqY3hImPs0CKqEq1GNiusLw3El7mgH
iFf6ChDsxXeM6VsKusVVBIiGwpCMxAqZbkAwv3Lo0cnEw7tZIhZyeIZB7DfU
JxisrB/5nzPdcPcivttDg7xiq1cS9jQ8cvsuH6iH64hAmDdfOrXGYAcx5G/D
/d/K4szvllkfZs/8/vaTA+ub+pskVfHBldTlQ40tn41cx//tVXNX9Yd/uE6s
lXnvvYSt98m3EcHCXu9MfPGCnVFIRGp7Gowf11yl2a8Z37y25sU2zxjoHu/R
41N2wEBUrJF+QFQ3/YCHUEDjaIfbFfmQV16xvsW/td71D76pNYmVVkqqcrJj
40tQyp3i7lUhVFsnkhQ+mrN7wI72DWLUxIDSe8lxrH3HKo9xD/hTX9DJtneS
PlVPOb84WL38QMIHl8fHF1qvQ1xYw0Itol8Em8ij8lQGw2EY8IVIKTkiodGm
gA4hV9kJSPnVzC5vOinA0kNmoeJWEXLbyx++TR/yotSryEbO2ny1jiHDxGjL
7bDYLAwjyF1To/0MTX0kBBKeFYjjaJDxwlyfbY1AJfAleGBahIoJansPXNEB
dp/Ao7GrliFryAJtAxNTOglo7BM4Kb7xCU41otr3IQhfV6/ikTNvtYD6l8iW
0PXMdcdmUWNOiUuHXH7Zjmw3G6glN93zSJh9V/yodOwY3ymuxLqfjyyIxWYb
MQ/Vf9msG/Cbsd7c3k6kd6iXlGazK5liAPzTz/RD/+0dP2B+Sv04aRLwg0te
pCaoXhmSRsD8esaTgZCHZA58RDuze7fvlYr6T1PvFowrRJ6x4f0tva6uXmfU
jcOrwZA4c9cICeyfw2yE+METWDbrigjWkuqE65TidJQ+3qie1SuAozLFdr+Q
onvBOeVfg7mFGMXgjaxNOcAJbD+wq2HyRW3avD2NOMhaZzjiinolB2kpEyZ6
bYjkieBh2TlwHA/erJLWTWIPuy1AAqXBOhiqpZGVsjnMp+IRbm2IjKL5EIjL
1ZXbJ8BIWVmouvW2UqWdb68rVhjjXzBXHCkGHLXXYrGrAIh+rYi8H5qchajP
Ela2wWmJYkGAK+oO4C2kT5Ib9vpKB/KQAaAPLbRr47WKKTiMwZyuEZRaylBx
xNOAAXJ/VNzY/n6QTtWrLrzZgcnSSJ1B7ZfRRxaBYYZE+0SyJFEAUM4QlZiI
HukDWO+BMg1UNgT9PXBeYqX5V6J/LvQiB9eOe29v210JKFtP/jTXnSbVHxxT
Xhz/51kXuuT/PW3na64vmbwkTpUDyPVxb7IinmJAUTze+A7Mm23bKA0chm7G
4B4MV2uK1giiNngeIXe4zq2mcgCmWlgzCXSyanlFiZFetpsgVmkSprMhnI2f
7BTsfkr8WfYa1xrWaMg/8OmDjIXAX/tPbJbJ0t77nS9gP/jsgFEPNSIUQP0l
pSoxizX5T6a1F5hLa9vK+4Wgwa4V8QlJTPjqwVuhNGVXfpKTE/4yMk06fcfw
D80cdc8dRqWJf+JBhSmtwxWjT7ORthFAcR02VwkP8IcXLNXMhOzK8pvbRfId
kLsfyZZnPXxRCh1xENUHZI7aN5kScAXX10tBez5ETNO3iaWyUNdiYWE5S7Qo
FMCuTSHxaKMm+++iXivbMIHaJizkUGRxTotko0fllP+FtP/JTpBsWcOOhkmH
Hu3FDlV39ibCAuha6qYvDI8/PB94aHEqOTwg7ytTwHBSqUKILJFaJY3V7hdp
Es3MT4rX/ugeLgP4i1pISYWkXIxh7jSdHDQ2da9pAQeJnU5he+b9nlhjGFau
VbwFzoGYY1McQcsyorqBZZdOS+hN0OozI6WvThvpxX8GxCQZbgLNwgBm12rn
rwWklbcz53Fh61iFgLIadELAG+8rB+vY1NUlrjrf2a+pcnWR33MVLn90ZW/3
bIBxO+i+jWRh3Pdne95nAJeemvyifidg74FAVJ+QuSa7D9xne93gxAWQumhC
tudK0d0FYb7pSWaa/G5/bevMnWfZ/SEfP5nyYQhzINdrsn/rpospiFHtgbgx
JlO5Q8zf/h0bhjWs+3eUC0Jmn7Ju34akZ7YcBGJ5yl+VQOrs1OJPbLo4k5Ny
gQ6pnJKnWQcj4/yDLs7yHeTt4p4PenDmMtp7JvccxjbypJM5y+ss+ABEayf6
BBoZ7zlegPy9Ywf80h3FagGuU5VUWDlQRzNMVocNbcmu2eP0e5Yatepf26B/
XZP5KJhKYvPPyZsj4SteZStwTv/oszw0e/hFIhONIw43/K6DiSwOiPqLRnOo
FoIxqZBc1EZ9+GIz85EYUCqTk33u0lpBMpM6518x9g3YumWpXJXNIxruaMi4
6uBu4RIc02ltEHOGMTjAUKIFlocXPQxVnzIsd9LxPjUE0wwnDM0GkVGpPjl3
XR1bn3wTPw/ST/YLDlYzqfqz78twOETLpP3aLby0SjiYHNM+KVOfTe42mASV
plvDUQkBvv6IZ03LU5T9Ko9Fy0WMIjwT6URRxds1dNUbgmDRzMCFZpL2C1tU
cOwlVTo6uH4cc3YwuA8DmsHJdTUjSo0QlniqmhmjK5Qkzij/iI/FJXWOF7pS
0mpZLxv9+zp7bA7a/+E16LjBVNrWVYChpbVu5xohjQ9um3SPFQXWOwAc800n
RZuBGgwrIKKVfraGpT6Rj2+wDSz7DR5w0UgI7DlEWiHM/qCRKdKzFhmr/zfP
0kL2tTSY37/h4Evv746iroFSzlIpBj2A9pQBah4qrnW02J6jGG/h3jYrw5Sp
13y7V0I/TxX2Rl9VwVWuXlhaYJjQ6usCTvsaHxEamlzxPUWVKskxjMMNzA7f
QYXs1qAEXsFM23Xq9E0vVQtF1YHRSLwE8ND4sOso0Yw0QXDUjL1+Yqel+/SW
ywBGSeCNNxAscYAsKMSFFV3i8KA1AZEMDRq2lT0jishjlE7ROcBUYgcOH9H5
em+ILWqzzZU7/7LZ+1iQBNlBI0O9shu9A688CbVudXxZmCRVFe5Py9vfymU8
/r2uOlZhG2G336vl1VZfx2Ja4y5cPlF8uy1Ai3VTLoNNmM+aISYfWLPnRVn+
CCdu7iyeYX10Qrej9HiAcPX7011SmxaRSSR/9sbKi9KnB+nnxmYN1CNJVEYX
DgKfwQjb172uSH/dboXv/3WlswLDnGrWaYDb/1HGUL5ylrpcwHeNZdqp4Um5
pYhFJGqeMlcO87SckoDtsU3lk4who2TMp5Tqx03WmHttmrJcIvFY+SdSKJOJ
nqZCtqyGG2o+tXFODRP02m71CZS77Cx9ircp1vkGr+GJOAAnY/hZvfU5u90M
035kGUEvE+n0/5Y0vkt6IBMQFW5E9pekXW2ovo66DORZPngsUzVnlBUqDbRF
48PnpPpNi7CbUPh5ZQbyHDFVhlwCTMCt1gvuuMRy+0xgNX9RgY7On5RCNiHs
9SoPSme9Jn6PtMRP0NInPmCgAKAiah/SrSrXdfW3k2YGk5ZxdrT8DqzKSukZ
IQv6ll7wWR85nnKGidF5Ysa5h2koY8vahjqHBXSKNiVnUWT4Rs20vQnEnvio
dTUXloNDovwTmukGClwN5Bi6ujWZQwGjriOiIpkIIAggq5DajRQQXaVFmQ5z
1jd+JGEMKVQBvlCvgH4h63yXwE13dxrP2k0vfIanpCTgGagpSPA1XGSKVfXb
wpR/kUW1ghWFhMsrWBbIx7n1SXrcaFkT9LPFHIPGznhuDy5gtV2rlu5GWjMM
V327B/OnYhuFnXIBa61aYYeSDx+anLOr1ZhNzpDr15lPiAkqOGjMePnS4S7Q
qdBX1KCM3wJqUaLMAXMFG4V/0lnwb0s1d/yrDxq8wSAt9vedExtff/iAuOkI
PQtbbCWotyfbc0JI494oBqLTaOOM508NLXBp9pMf404IV3WZ45riHRG7Amyj
X7vb6CpC64Z+eJkZc/kmpTQeHw2J5RE19dKyVG9y2h2NqWyvjwBhvZuth32+
ECekxiv9ROgZliHwopJCc/GoUrsiIlnmf2lgzc3eerXqeYMpidbeuqRMK9cy
ZgspKQBLC23sBjFDRND5xVSpJ4fz4L67Ch3tcegwHSzHOS9wbUH+1dezDjK6
ydVcQRh7noJRs21RCqX62b/72P7Pode/FjerDY85T/ONvou0RWqNjSnmVbLY
zLaqFhe0AtYw5cdSZRNYYDEkyIU19KI22WB+XQmKXMPgVo8GJf7Kb2qiwVvq
DEs1hEieL0FU58dhEU899GClk/SJ1FabfI+MeGM3HrwOJ/eX53ryzxxhHchX
RUbv/xrDvwdynpA4z0zGLwfpKRAAUtFeaKrt/FlbGC1jUMYlEH0/BE0QrNQL
ltQS+EuDqR8TKfgNdwdrQY+lUPoiOvy95NZd8cONfjPMfoIFLaqN3HcFM92j
q4frcFaSrepglRs0iwsEYqIyL4pCvNz+n+rXlEK9FeVLMYT0y5sUK6GFtZxd
dwa8sjIIt/tha9RfeXPa7SFPAnrSgGtBWRU0XS8ZkUxeHFGtieE/PYutG2ZL
/MKVQvwUEHtnUJmffdydtxdbE4pFjVzKiCOVk6QDf6zuHElT1idXTnLIaM3H
hx97oVLYptrKw6VSGd2jzaqJ0OZAKLddXjbFdEEgxd3Kc+47h6/gr8R4Riwb
tR63pF3aKKwENUT6tPZ19OVZoRBnjOMO8pkU8tqcMnHcExsP7Pn0uy4DUsMm
nrNniDzdi6SGW40GRBXGPoo/0bxlLpqkfe3/6eylxsFDeCvB/n1+rz9Jgc8R
wPbTHRjCKNOA43r7UHUJSbhTWTiA/63vWhUB/HeEDa8eVzrkBd1roGJk/Ab/
GexHmM77mxPPkCizdKi8D/0BI8094tTGjpf3smbFBsdUensrhZpUUGrY4/Ud
4T5XVUN88lhVJtPPdlFeputRfvz+L8yEaEz+HTn+zp2mT/iFrbSra+UW1hfA
yA3NmHwfsgvoeOr9109OxwHKLK1CRtm2AFaelNsiRKkZ1NkdpfQxTK1RlI+U
+1lj0vY9vEME4zSFARgZN9ZeYX+hv3NRHKAvGT72ZUNtrlEOpl+PnFEodfi1
iJ3XN3QhRiXyZ1A6G1TUA0uRTdHORNCEHk+nUB8oOqBP7+2X1qhhRLja2NUU
oHvITIpMVHE1MSgGz1/NTmSVCNoHP3Hp91E6Vt5h5sjEU3eJaPfM9CxW7SlH
/2uVEkngdKYiyj9/qy75NYgryHB1eceTV/hpPuAndJel8lwtuzFpanF2dYhY
2wAy5pJnXbjUwYyrreB5prs64KDD7E6qd4Xi443oFP9DYrd3OQqaoVQxt2Z1
2sO+IUpN0C0lOJ4GIBbeuw12wUNniDEbPEHWz0WZ77I5IqVNp+xwn9YwapK0
pQdbDV68gMC+PC2fEOlO00UPJKmMwJDySra/fJGzEH1XdEgo1Ahs+eEQWcYO
6Nj1wvsyTncsAgq0vpVXuHV2/O+Fo+i+nlaOVu4982gmrrnrgBodRA3cIUSp
uo7WquCKGGnXmuRiVmnCJ1PbEGr+Dp8OqvGHcHJJjoHllfUeZZLpp+QvKVuL
EoFofL1rUECFEQs4H7fIU64U/1dhq7L9RtyPD5lTeMLCtgYM6Laquik1eBR4
cqO6x+i2y4Xf7M4eTJ+BZdMCUK2koXkE1z46AtgVPXfX+FsBUn32U+UCnnXQ
h0bTVMfDZZHLceXpKlcjA9GxQrYQQ81HecBp7tYAvhHfDyqDFdN5XO47fP8N
1TvncGx+jCgslFMWdfrei5Xg8DPKNmyYNn55RWw2o1zArLeVHFcrNgTEYhmM
2+a7O7PGrwZDBxlbf0FBibd1xvXoKI3/Pwzfk/l/Zfm3X7YDaZZAl/GDCmsD
XeAW51UqnffU/5NTDWmVKpioyIkyTwA4sbFqrRjhtLmVoDIWc3Ti0iQMilZb
65LzjLdMLMS8USIfFZYvPsCrvntzSmL6OUfyhmJmlgGm417I54HReHTHukWT
n2dXHBiHTyjEFJGM1WfpwGBjEawoO1Mzo2yM0W/ykQS5vWwoGQy9dMhCU3VD
IxZTGqZS2gl+iHcCCWXyqUishb6UB7PVelX+UPXr8qPrnJQTw42Ic379u+Tb
y8cXdjaZ0mg0CIpf9/L0NDqld4G5ywtpuBZu0SioHV8SH/17MgiEWhLaBfw2
FfWe/L1Y5RK61pNWGiGBL+180+vzxgVYT8Xpkci14zWGstH/XFVsZcadBB8F
ajvS7JPU5UyKIrP8ZN5krXeb8SLhM2B319XpdjmTHirF/lAvhzEGRFYBsHM/
9wRGqAu4P5djcP+mdf9IUbhQVQglwlss4dUc+yALrCyUln9SOk7S+NSdLXmG
wUWlTatrTqK7WWUnl7YIRxkJbVA00ikLiuXyBf2VnCou4a2LPyFbha5/hGxU
19UGssSRz3Q57Ouu5JCbn6YhhhkugXL8/f7IHgbF44GeVrinkVSxfq8ZHEmi
1+6TLFiJSPc1XfbFK9FDoVw4Yfo1z6HiItJ3mQN0i1GNXpQkqp5Vzk9gjMRI
amgQ9raYp7qa7X1YlKxOyuOhyEy44A6mRZgdqjmiv9P6SO7yD6Sj2qNh7G89
Vz6CuTTWwBhiNWYeoHsvCi4DqMtks1vEwS5uIWj+/TkU+ngBFsHrVP6ddPJ+
R41pXRcWyghVmZYJ0H9rMUIxtpV7qmGDfL+m28q1IytFPKyhTj1ZCopcy6iR
bdO/O9QdFGY6usDd69nlBeLcl9h6rrzjVAk5eLb+/BuENKotOv/4rCa0m7IS
QMcDJpMqZb4M+M9g37qRbF4ULGGUZ+Rj1wuHbVCcdRiXqPWJgrXYHoK3ABNc
PcpIcZKBgNXIZLLyUVR3sJQyCFdrR3bDHessv7P+e0RGd3yxxQ8sJHWy4KWs
guyj63R7eNWIeGTFGEXZIaTC+tbbkt5CtUo14HcxpXJJQRt+CmQ1gyippQtn
0yT1eFOfpoB6Fa6vsXFQCKSwxZ7OujRHG7pQpunv8VsIBHkKqOZJcuduCnbc
VfzaalicHJT6aUGPwSe+LEPsoEHIl3/Tk6Hy1LrTBLWEE75lZOOm5AIHouTj
bhzfhIjQEJh3L4ktqWQG9GeHkP2CaivBvxa+x69B3Lell5kXXpgNy3uwW8LX
5RXUW/edO7vDfTy/94wYmOQCmdq3JKjAHkZveu3ITowh0iU9sm7LeXBAgdl7
Es01zugiitavXIo66clpHXoLJGIo4XS7SZNGwgWuunktIZgqhS/odlhTcy41
bXy7MWUl6HGEbT7oiwKbdXJKOBz8vVPzp+2c76IlklKgcKULf618Tw83XcgB
cfGyc4oss3EMlCU96JF4EZGT31bYzydTh83DjQ1IlipIUlWMxrvp7eHs3dwk
HgYfi/hsBkkoZ0CBiHOLK/lcSQZypfkZdh8pXSJWaYAC78mtW0XiU9npONxe
MXJoPQkgCCenc/zcDO/63gc5UaTVycntHqzz+ScTlyKc9dT4nZPlUUz/1xee
5Lp9kFbJR8R9FtzJeAltKtOnCICoHZVKYUlox/4VTHYCWIrvxQPu1eErPo7+
hR14UadvblRTou5UiAvaux4TZs3vfBu8ovC6Q7hVbD2uZAlBBjqNOaA0V49q
IGagSIIu0kRTGiS8T93XBMfzmYVyezHWfzn/YTiii/1DieYuDmbuIs8JA8F+
DxacMA1NSBvBI2oiOAU6XUivcv8Bf7KNlQBIBp0S8B99y8nDgs5FhszdoBlJ
3pnLpntm5QDuFahNrnkcRXFkfCcRF37kWwEQdkGw03GP59S2+MoT5tmICwE8
xDaNQ/mgR4orsysSv5/HTjsVZUQBP6O6bODx7IpYO03+QajsYKSAmF8iXZPN
C5u4Xc+ALNLn0GtxDqCC2L7S9DvDVXmbMGnZYymS5tpXXmZslah9lRyjMJfc
ccctrb3LRzK18fny3gWOuAERmJiohHmdEHGUJlZrzTmFMQcBNhHYwRZzeJvj
LAcWNUhkDQX1R7wbrRZAeJagCnVfmTGq3O4KJ5P7OxH8J5NdH6478AFogJ7g
UQDeHw85z4BSeCKStEFArXem/Y/tPsMIYBCVYSvuBT0lIr0UPv9lkakdZwhV
NHFmCf1tM29fFnJf9DQNn3AIO1zzvizJFOyNtXogjvXRMe3JadQ2fbIlapOA
odcvQN+OCU0YhRIEUvQEc3iSxtuw2eXdLNCsU9sN2e1lK2H/E+UssYCqZXAR
clibEjBcgjaZSaD7NhYMH/6JZ/GlAOZOj4Eu09C5+Fgtb1zufHvsyN/0UmbZ
XCONf9JCgy9RZVK8ehx+m3Xeeqr8xTxpqppGiaWhDZ9HLyUBkk5nUChGvvhz
F3H1Fk191R1KUFdWOt/Tq/vpKyVnPtSPMHtbgwAAmJMXlKLFPtMHSdSw8dKJ
Oqqj5DPxuTVNPhUpgGDwkwbrfGZsgJ4qD/Sjuxxb3ndwQBRpiXp81H6pTnbJ
Rj29lf2lzjy6HB3UGbC+8QCQxZX0UTm1/cOyYvBvyPcTI6L2kkslksFxOg/c
0ZyccPf4oelWJeF1AmeN81Jib9EqO88erfD/rWZ748ijqzGzwiwGI6ZXAQQr
Pj6IykLoGNpQDDNynIssig0prXwZIQEpnuEeKOBvdl6Cp/oO+u36O821DRUq
q5Cc0yM76pzlqqeWjcnHctkIiPsga72E2Y59PmDQG6oj19+G37ixC2EE73nu
lihRxZxSMaEnTsfnL0RwYn6rmd3Hw6pBAZ2ABb0K7mg+laDM5aPHuOFTlTYX
qJFa3sqKnRlaIYpbAP6+RuEhHhByy24A+OlLZXcXzS6sZyKrXBIaytaQhJsk
pPImeJ2iDDlgZX9aK4uxpX2kL20XHtIGhUyCQ6adXGi75gxSuU3vzXLaVLLv
8H28I0aQjmxXeLFfQpZitJeaqrvnjfzbGX8U3wF7fTeCAYnG0OgofhZV0cgf
4/EXPRI5mUfHtwILCKPfnTSusY/P4sQMH9zG9+sOUVE28AwAA6mxnwNpS9dG
0+b1Jpw5lrQ50KbxjdbxgeH5cwbqCRd8Nk+X4AEZexT4CSSbzz1YKWQUTfEF
RtPcMUfj4yGdPaqh+I2/4JVfxOXS9/fLSq2sJ7/tznSSTNjvS5FHrZ2xH8Sr
L6O4WjUJUtocov+iVvoRRv8uHvPh56YcoJivP2FH2bD471DGmRRDGVBlJOo/
9PO/bWEPPdHX/w+/ZWoW+utzbBKUm40toQBslYXT+zLbNU2hdzh127kTgvig
kMxPT0/37EUUDUS9v60DrsaLAOqQSwMR2P+15wMU7jaM68+IZz14OvKs4ojL
kO+jWleljkMm9NNvNr/gF+5Vzwk53BBlY+YIJ4Nuv/rcyH0E2Vek3Qu3RTwq
okRtZELATHRWwWztu7tyN+gt1C1JHBZ/bLqAh9aVSdCrt0ZDR47fp2vS4MDP
rBIFMFG8KbtJ+QzAMW2ycj4wwcusZtG/ZkSdLVDpOgpmRQmixyfM1uHEsocy
SnjIRy/grT3mB0/b3IwFFU7/rgF0an9MoZKvEECLI9m0nhT8hBE6zeLAQEoP
QiKKFu4I9O97+/8ExslP33NoYAtq+wkfZ75zGYVMbil6drf09UurnRnbMfmL
9Rt2wnD7m9FuQv5alXIvqp4Jti8XYK/1gpK2DY8qbtP9Bm1/+0furEfcB2ka
VHwd4gZI+zb8wLJGYpI2ERWaX0/g93X3Pr34HgtuMLm0hHgsTi/nhQPS1zfg
R723PVxmN6RoIXpTnvUJW5V018Q2VsKEYjU0llxMzYlHE/yMI6fU57QqWdC5
dVp3m9ZOIvefydkIaE2UGi3cb3Xk2my4OOCh3XbDA7184gqR5/oJccZgtsrF
n69jqsi35A28IL7F/RImu4amptzF6zitdzI1ODZIolCo3NJ1hSsXc/T9G14h
oY3L03WgLojXLbOk9peOePJwQO2dsTq32abwvc2K+UUu4A7gg6g0tdMHkfbk
obs/REWXEJWBSHeCun2+zdnolG/HgvFZQFRArUx1HyyufXiYJhrqoIswfiLt
U1PJyRb3EMO8VJcbpSe9YeWZFM+8qGD+uSNNYduKkpE2vHW/HAG+YaRr1NXa
Y4xSnxhyhL5rzMpqkFOJlqLFQ2P5lh50LMRjkEMUpz3D5bUsdfEkzhIEMQOf
VXQEHrFhpjjVY86Njz7HF0oAmtQe3GznmloUFM3mrL730ttWB9nAIC+BIcn6
Z024iQZXThT5JL9Qa2oecZLkfIZIJ9eAEdKSa0VgH/0l0qQfuiXC7g+3kR6C
hyE7ZuelempuErryWKr/zHp3TXL+YUAhgiP+Uat2pYCKe6CBZ+zoCBDFFgyD
1Ba0WsxhZjor8dLLmlxiQ97Q1vcW1SAZYYqQOnm9iNtcTD5lcq5/UMK26dH2
DRvKiZFrFvtT4lR9aCSSQUg0C46MPPYlDQ7Y41+Ts2TcKCSZP1rQYgeg8cnv
ZZBsNhVzqQx31g9n3JrcQvKpuseAb//8CxHTDDkaNDpOk9s+4Py9yLhvZ7VY
Uv8VYUru4oNYL0V/vb1zWxcneEPuypDmST08hF+lS36+rid6xDJjgR7z6Dis
+MAxqalNnRb+zzJV0BDhuUZn7vFbzM5LI+NTtkRbeVatqPCqVdIBQ8cd1mVc
Jwyg7KMSbr42F6c/ThLZF9J6UBceFjXHf/2jCRarCSyDayq1OTpotcDOgaH0
iysipwLaDw/rrRbKLtupXwY83ixfOpI5hEyIDAL2fPiKjE8we9XEczp2u6eB
3M1ovJWZEksN+7fatDaF0bg0cSWC2lcwXpecYDfYWwRYixk4w2JV32j1Q6Zs
/mAT/MDUo0u6SucrPilvWjt6eD39Fy2WDEfgeixltEtuysTi1OCyAkk0Ithw
5gfIfuNgewtxPoDJpz3l7RrC8rYn7LWu79Vmd66larJl/rs1sil9Z9VPOlqd
HIYAcLhpLBEAcxkvLDG9nkJ4o4YTb1rUF2mW8E1sVRR8xF0H7be3kMh05IzM
EE27mJLiu4vj4YBOxyhX5XBI3nH8rhNhusssXdC2dZ2wnijMCxJ8kecMVk7Y
vNhgKcUQQ9UmHsMHL9AqqVmwmuf1RHOnV45D8yduswx1EO4JxTQkP8/blciX
0HsqzKbbE2DYoGjYzCca+r4508q4xuWCnn+vKmw6Ohix/oIsQDRUgaSonCpw
TaYfPG8Oe12GTbU8kTGcognMep90KmgzRVk75rwAuRw5/gNPhGDUlv+kcgTE
pZNOjtXJsAn7o4VZv9U3ZUIZj/NS5huua3L1g0No+mDNa9orXGu/IUBKqkeR
gkQyW7JEL9t0/XmjWRdfUwOtEEB7PEOmPZCu4irtfuuuMP+TyoBaHHRfKbZS
23Mue7pJ5Ixzy4srtPosWsC4FkJWWheAGhiB4BFbu4AGlcdurNWZjUs/Gisi
mEbmeRcaD4hJvxKn9LvkhZLvQ/AKkeE/XefSeERse+KUb8sNNTqTHVid8ny8
qixbbzjwhD35/6P+cqMC9gs/9E2DsYGyfK6hd9+lpKE+uAwUm5c0KhabFETa
0eXM8k2/yvG9zGhiZcboNTUTZ3PR2jVixwUZ0e7uriVV4+urtv5YTu2Gvvpw
5CbccU0sPcKKrqs5jJiodWfIeFtMFiyhyqJDnovyHhKa+v6A+6I8pBHONQF8
Nn4YRp5CdH95NH0r0UDk29DRd6suiBN1xQ1qEafaKcOwMPPq944pUB5j847W
dVKa6v+Tp6WgWB3aT+YTmhK7aW0tDnWG4GnxRgq3SK+LyYrV3XPVtUofUrYH
TnBlgoLIwEiiSrVv9vc2WBoRhE/zYUNoMPosAki63YJUXJzxqhMIdlm75owq
RHPB6CuLh9ha91HA5pBU9HQ1XErs5Cvec1hgnXhfXA0xK8OzdCxdraytPSTC
4wE36Klb2i2DkYfZUdkZwWPVOHkF+5TX/cZarNyqy22nvGjqQROeNGus4Dqf
hOTZfGykojOM7lYgamTt6e4+6lAFOIphq+k2gDCqo0QR4zEZvnWsWiqPIy3I
vr09gJen1mFF96Tk3ilrfdll1Bt4FovaSWrDj5tlfVRyrPHYust/k1zVqD2U
8VyzgrpkuxkFyW51YHudBBUOrt2spM33tlgyI7Tu2W464t9K6PvVsxoye/cS
kfiE+t5qUZABS9gfF9PQSPcck83Nxb+yXTA6S5lAdypzmFX8++eMAFBhsWQL
WqwtDjnnmgP3UCirhf7qW7rPVKwdXLSPE87QfR95tigfrqOMYmMqBRXSPEB0
vP2ejx38F96gXnnSIWv5vAZ3A+Yaq+eOMObSbsP61OMY+vp7kDwqR8SqJYBW
WwvTqHjqQXpBkLjAZks8oodfzRsl7JQTOgf2bFQ4pHfi6Wz9V3/CxcThOvXA
AZCJDpqykMQ+vjoAEIyVs6PDY5+Eewhw3bDKzir9x9hwTdbEsCTWyyHEwvki
j2qT+NuRHos/wO5rFdK61PsHEEgsJZ5DW66/aL8zz15ksvr5Tu98fK+X4KQW
x2b+FxJyRQJfYZZ/WkQaanjLr7lLBEp96g2hWOH62hc4hgjbpNCE7baRb4pf
k7zPQZf897Le7cDIy6Z93UTdhEXum5hTD/JauhPxC+SfgxIgD5U4Pq7LbuhD
fZv3DjS0gBqNgy0hHR/M9xyzoBqriGAtpbZdUO5Z5CaxnKEPe6qlt9YuyzmW
OrprUvIIop5zEpqIx5Iy11aURwbquwKCeacd4DQnYK/4/UYs6qsyHiMLJygD
aFaXOrMek5ZT5Tyi15JafbL5LTSI7ljU026vwP6HvRbYxUJsmH4nUA3V5JPp
6ZEjDt25Xfp1tGUT7brMX4T7QaW1Cs2B1p3lLuYXtlnLiBmttN70HXOG8XSw
bW/0UIVW2PxXNliTOnVhKQnLhmO7paYVHFPWmDUKQJ/ZsTVALWNjTCzIVcoO
GQVSK+AuMRAyr6ACB745WyYzkLg5SS0Rn0Ig46oPvnJgtecFGZAJGhPj7Fry
oLtD/g9PL+oaiFHh5ps1XZ2033mNVktnnGA18T5PN35xggS8FoZ/56F/x/BU
/P9VUfCOwaJHvcIoKI2mEDxcch9i1G1aKYTb1kCr5sXEtcTtX70H6KyN8n1n
tioWRP5uPpFbYcumEBqZRFmK7vAMIXhG2A/YAQvGegiN30q6N05chyntTKdJ
O5f03/wr9AYRRtKhQYsyy5Ag46+hXgzVxMTCH4bqzsdabt5oNOK6HVAm0EJX
NjNJ4Dm4kg6oxp7ySDQHfWAhRm8TUxaWCy2MVzKFvsEiGgif1rsyd0DILytj
L7pNGHK3leQa9NAKEkvhqEOad4Q8lMHwwpRX6dGaLJXNLlLIWXTZCuURtmza
cOocMGD1qZX95dpypdMbH+IEo1MEOMi5rfBXvl3GGTZlpwCZnXtxmZkG9gjG
tyyCVA4K3uwmjPm8rPKidt9Dg/Q/Lhtm/N0c03Q9J0e/seLZoZIqCSnWEhrU
k3KDiiopRH/BKhewcvs3MC0lucbwYyaz2kOUFEh4J4IHvpJ/HV2BiDufqjm+
PTYz8tmtrorLXB7wYqbceKhTTp4TdCxEF2WYvz2k3MNU5CBSNBfVwReHvBko
wWIf6fXh+VMFoX32EfX7SYaglFQRYu90NP/3D4gUddZGjKDnGOd3TE7EF5tZ
YhL7hqqDgRwyNSMWy7z7AzAjLL+P6xRuFIrONyC/1I75ATmVsfAAePOmBv31
Kr6vOVtRK45HUoK84pM7ShL8iLVJZm8zfBASHaDpL1cgORFtHErWTPXkXFF3
pNLoqux11KWD5L1f7bP/QKJXXpWs+AYWhqJIAcbjlpXwVJD7jY5kgkwDvx5n
XTbAdK04qZzQSs19KjGohECLAkd3en83HLvt5CV2FcahRpcsbsGdH1goIvs1
BdshXh26GJ+FjQXYUF+fgT8eNinNqV5l4g/qFNKDojHIz7oqTRu4GCdDlju7
IYVJY29+orSWIVzp9fHOiephNvrTJOnloXKnU/Ve1TIoCaTg/BnjmOKRpspM
mGA/bagC8qdfgCLE9vUbRcvj8RjiN9mlSc4R0B1rNKRE97UHMoamH5nuUbTE
udxOF2Tf+RGlLRZHH1WZd4Nr9JBeKOxuUtrSYgDluxB+/RNwzD4+TG41B/1i
/ojpSvCeRjcGXWxEUVNWtpOP/TEql0wWicV01Q+bfIgT4KcIgcBovauc1juu
7Il3qpCOvvO9zVZ5lBi+QpYG2BxScsE1g5YYJ4qf3mC48fLweJoZ5875EZ58
qPO4bNsA8JDHAdm/o3kSWM/klYvMKWyztnm/a4oqyE/wYGtLGgwGUFwZVpxM
jPQLSdhy8ASmj+tyLDYvBpuRgCbfK+j1eAc/D0W+t8u+rIFBtKvgCdKPQU7a
NUmx4f/WPa8fgjAZN6Uk+6DCWWHNbI6N9AEkgvEvuUUhWR/HCVkNdAeyM5SD
vIH+PbIZNlu3RWICtscexdAh/Rh4IphaxQ6c74E2onQlqbl3+dyZsg9MG9fo
sVuVPXG0lQquHckrpUVYpL8VJkCDtdIHGyz1Sbq1h1cqzx9uFP3zPa2CrGUK
ASIRJYerF3ws1OmcpTo0oB8xhK7dY35dmtVVdJ1Ow/mvYkcpHBYLy5WRa74W
Y+3SyKtnAac9pUl1AQz4LJGTjpM972VVUF4A2zUYtVUPlYfZymZEleb/BADZ
pABy6eJ5ehUaiWLeF5d8lWJHuotfiMHs7S4dXPuk5icM1/VTe5K4KedIwBic
ZiSo3sc+eel3zHRD9Uz+Acr0T/vFtsBtzS5w75F8R9fdJr/eJYq3+jbmsfMc
I7m2h7kbPjPb58DG5IetPdApvGySzVgk2YAjARkld4zmOYcp7RjIoWKsSqM0
AKbObbMNXSjp0JV61UIlT3EvLQ5nD+wo9l+gPXXOLS5Mho2RhaJu2rZmaYtH
zSCdzyPwvHWDDmvYRmY1T/q3uf5/3tZPcKzqeJlWK4QOHziBi8ih2MnmUnKv
PlINtxQPZmvJjSPNRonrJer9ylxugPDB637oZ1Pla97bK/nqi4bw+b80vKTO
HJPw9zfCLU5XJYI9HJA8ff5IgSZrdUq3dfS2MEx8xxyaRKJwmVN7UofwHjeE
bcxMINZQVjdp9TlGEhE2vBGGtKLHdbHuMgRfIBF6F2n7Eh+yWh2lpJMcOwCR
sC2JOTERBFdNc5WK9QxBj8gb69ieHjBfbY+gTm7DfFA3r012J3aVc55Kx0zD
D3EkO4WyEm2Ks/Atri4J+Qn7bvbE9nZuq1HKhrXH6Sh/7U2Q70yAZN4+OQlr
hZCHC4aTd3VdpW/nELziDTVyfsOVc6IFZuzatIc1vAAN52LebN/6bc/nti6E
7BaOfB3LOXzlt4fF8PX2+6ibu26wTHB48j/7HB0Yz6+HvcscyR/837IXPmSf
eNijQU0Xok+RyiWpEjCEwkXph7PVFDDtuZcxRTO/NbJ465omPq59f48k54sb
SSj+Mwk+eLOhRh/k5/pzfl6idby7EyhPNK+vyartV/DFTwpH579pP7wuv6iL
/70GlR28In/BYKCh/jyMtMdjrtTKQFZAuC57wkvEPd/LNF0ADRuHq7wsFB3F
X4t3iDwMfx4xKML2Y1SSDAWmF+QZCDzUAuFYEo9wI7Zo+NYPjJ6G4TOYRR50
gLYVQ0Y9H6PsUFLXTiFj0DY/PTbVSMvXAqij2l+1n3qxOU6xppVtdF2LuaWo
cS6sL/Tjc+BkzrCcQhGC2KinFXE1YY5Vl8lm622kQ+X783bPNbnunWJEWB0A
K6D6WBJhoNKAaBUm0gjbdvrka5+5s+Z47V3O1ckX0yHZWhGiK1TJ1lSIlnzV
JL6o95E00Fg8kw6v9Or/phhXxkP6G1V0nDC8hVsGAFY5FYD8uhC/bkLAP7ep
Z5LgH3AfNeRyU3cBclA8z8ZoKOH+i+l235EIiJ3VqOKS8ntrM6zIO7wgHn+b
jSD018jsufxCdT5Dsx8y3a/EpUzmHRoyMwupZdPxDw9N1pHhASbtITegush8
L1f1nmA2nr89SQqlXe7n3+Ktnq9xZPNnQ4XfmVWmPUCd+HTl0kfgb98rqjL+
fN5I93+lGZZ8LhNk6sxNYEXcSnS8Kt9v5qbDaVFOKg8EJ2S82NhywOAtTVcE
VGSw2TynYliPOctpYicyUBntX4RgQ2W8P6BZpEx9/UUsPQF1bkDa754JVioU
Y1ZzpW9qTRvrNMVBPRxamu44BYVZd0JAEtXTrOoD9ppyNPOXz/b9jVhBr3iD
6DuxH3OuhB19jAawd5RCefmeSesgeUwhgGpH6rj/doB9apRXScQmRazAj8Il
q1WySzfQezrezxru3/U0/2korZw+mO0vbtEnxVzsNVmCwzpqv5nz8kCFBTJV
AaBPDFs/oL36DF+JMhHdSFPLSGX0zQLWY9zeg344bs3PUuDtzsY/r+z2D0Ph
dCZUs6z0PuMD+klFDr/4VN+nNzaSGTWYhxDeX4L2zHBNUIUjk32jtkfWzV/C
B+7mEVlqpiPP6F+dIC8dZVJwqIEYcfPn0btoA3u21oZ21j4f4+4uvGqWbhgh
BFcAUJE0qBJEwATsHHeLi7TKut6qp56jVZxr3RRaENizKg0EWDzwScdNr6jl
WRMCJMXqGgfZQQCC7ikMzOoMIW5RyG4HkwtT0CQxYltO2Ym510RERfS09S2n
jyqmXGuQssJQj32I5P9A3MwAhLt24f901DW9fHxA55VPIWSxOdKIjaiO7iXk
JltgmEv0P05jHfKbzvwJVVKKkTlAki+tchwewxeVZoALpkhOWqD9uTAOc8hG
iW+ixd5gtQbv1oCR3gxB9TcjeCodS2zXFyo6wXiZz1Q5YqXoKQ6dUQkDcMHL
Yb3oIlbfD+dyYFLBJcuGPOqoU/G7I2fjKh5+/C+Lfj4Dj5QJ/IE3JbYAffSX
RC8ZplXBjBZVCictaR+Ixmc7muCqtKMYy5H0EXJ/rMSZ4nk4g+vTvH1pQuWx
k3TSPH4EWh328nOVILXJPFmjhzz/GTTgfI93CXfO+pb3TNppQScc+xJ+cq04
sr63SeoVvqJNXZPTn/5lFHuGxPYD/GAz/omPYXwMDqhjOL/cVHvXZGVjEhpq
CCg2WCByQrBjBTCxvB/o5nnuGF/+Auy7CXVxk2BP3jSFo3uR+AHyvbHp5cVA
gGjuBenMUyeY+2j/11cFh9lKPs44x+ebVlssMpHdBQHdfhtgp9eWsuhs3X17
pjLMeq/As56W8saMj+ObV47I7lNAl71SKa4hasKW/qrdslw/RHnbkHcHKwvv
ZyhGtZJuAVZuBknZbfU9PR9Ap6joEnUtVavMau6GhU0a+6yltXAFnoPU4g0s
uGY3kzCLGOWhZDLgUa8ca10XcVKIYPRenBdOqFEcNAxWdPz7QX8qblyFve7P
++fhiioKTMY5soRlfPuf44Km8eo0so2mRvYM+CKj7aQfDpD/R0brHw0YXnHU
vkHV3lJdH9iloXiyc1dhMtEpTnVqT8RKXI4RGHU3lE/qVkbGQwq60e9VLe7H
I78zxlO4eHaWLxV2ZrlGJhVhQwrkU+VjixuKmV4a7Z76IomLmTpG8WbUqG5a
yOzAttk2QxL3iEmDxJUtI3FuwEV2O1omtPXvyWdRmbBDodfeKyb/PLkTBzvv
rFv+I0mhMz0eP+aKm8+qqhOd6HcYODyuqrLbANT7weiM4uSXREVgZC6lF1FM
IYBc+kmdq+XHDwsn9TsRS+QDaJLFQkoav5tp2eT9AwPXwbpVqBJO5tnDRwX6
w5rjX+mRRrQ/5ZadcOL2dm3AfBmWgmiIAWVrvumvaqK69kEQkBuQ+6y0kvqE
F+JE6fHGak8Xl9c/JiDH/VE6xI3KcQ7RJKZbLRIi1Cu61gj4xMCpdZYq6siL
zqMYUh2AnYMCnhcRrJ7/aOxv2AARerzDdtRo8+frmO5ZndeoqL77mEx3LUWo
Mn2EDjeMBT/hOIvsVDIw30tE0rwJpQa6VpZzZIH6EozCEh/iVDJntxFqTA1O
0toF6tk/WzLe8y7OFQtSXUhVfQYEuXifL8WaGdUrHLjew52GwNZW77WfajiK
i9x9nSooVGe6TbphDXVAr2e6M00CKXEKFa6J1S5Jdru+it0tVckm6RJvG5kC
lacVZn7aL9wytAn5luACMLNB3IMUp93GMA5InzDhei2cdpyCXkNY5u+rawfR
qTBI9wVGU8JtGW3QST2cNbTsCg2h1xL0Qzmh1GHnFCx9vj+fh3V31obQKKEq
ENqqn1ZuEZ+d4RtnqI9MxtWsV3WpIS61BBUwi4IQm7XaHS82ZIv0+7yHdl48
eGRMs4K5rftmGKsS6rolcVHdAs42UDPlKdanyzEi2Z5BKL8Zj3XMwe1ES4zO
0IJr21woqxiVqVl+QSgUYcjEk5atvIuZXTtHdOXcNaNNJ16u16I21kR2nXdH
OQT9Z4RFrZV+nfwAhvgmAKg3Lr7EyWyyq7nZuPitZVgY8K5VDiaJlT7omNi6
oTqCN1BVlI5jC9m2Z1CIawJSDovK1XnhX8BRwMqsvbrKf3N30vz4Feiopd3Y
Dpid8t8fMNIAyex/cdHEGwGvDAErTAXa3/A74yrSm+NJyn1ujEqgNhUTefbv
uyxwVRLpczQ/yr+WoZl09hfblbK18vHLU5Qk2Xwjz4maeyZDkC5ndPTRrkkj
7MgqkVcIE60jy0OrIsuMMDCp4yxvqQkQunWvrmeOmw/kr9o1jC5aVnPBrSR3
Bn8ATnGOA6xoH5hThtVSTERUu6HxgGcrpRp0UNcFDWQUig0na0BYG0LRDFzM
zD5Cmn5I+vinJzohhNYVqPv6X4pSwsCKBaz4qc+eKcqkc9W+3xlWpum+XXuR
qWkbLLV6lWkWJtnOikgLPsfQsdTGX7RxLcmBx5Agl3K8TuJYJmUf8lmeE4Sv
4VK6UHgq0V0VcQgLnE6IXIN9KINGIbf+Qy3oOd9/NqK6cuQAMlkVKUuHJa8+
BwOOUrHQWObrB18R34EHcJ9il/x3ciyzjZK9vAh5j+w7HE4zqlJTzepYGoWB
gFNeErI1+Sar3DhZZO/yj/x1kHrmuhi6WD7Nvu1sonGM22QATM9p/utt1O2f
SWxOJFA+u2nkQl5MTjUMSc/DJFySyONp1ZGtau1kHRNKO5z268tPZMEBAoRR
7s3e/GcYhyK1R8HtapyNxoYqJbozCEMSJIMrBu8MbzYQlRtQWL44tCPgfDxB
ACSBYMtbiIOaVxTDuuSEB6lyAi1gwAU2MIlxFNdy4QeKHLpEwE6jbPi4eWg5
lUqchNrQHz3PWEJYdhdh9tK3Z1f4SzquC/nJ29O/ll46nR/IUvwNd41j2lip
Twp3CdW2D5e5sSRwRDxIZOxDJIz/WZfJHHBOyUIGnyyIJ2ID1Qiui+ownXbw
nLJgzKw5JRiFWSB0oOdI9rfUHIbbJlS+vsLz71yd0Co98KUbrj4vgC18CFyN
pXbzTjYVRttjeR0CPOPX7715b6TQjCbR2lsaxxJvlZ4euImmcohBDVvETtqD
mBOoQn761wAyiqdlm2ZtN+qnFWnUL/6flCeTD0+DSBkYl/Wrd6PxxCKr5W10
wnKH//Qv6P/+/lq1EHMXITKNtWYyQZCX2cfQU6ngmEyXTRjm8fTM309iqBwH
c2lICcBSNRltIptSmtoiwvC3kEb4pP574Jpxk8ZEaJbNjK9LyK2pIez5MJRr
dY4uts4Ez6siX36I0c/fEO56R8NwtYDhfrNhE+hPU4E4eFrIG3f4bQ2sywJJ
lI9XNeTOTgTuJXv4h/jwSRfqDDGe9hbgBkCrxhS6VTmVJltKqyXyqjbLJ38M
EuCc6HZvcxT549TxL0VPtas7HbkRkL7FpqO1auIBUefK1A0MgUkD+cVf+NeX
EafwCXjlLkFy+5ND8Nuqtabu0fi6Z7bZNrzajlSYqTCBV9qK1OfUcDyT0Htk
VJxMGUSwGwf5k9KZvU+SG82I3JJZvzxZtmd7Fkv4UL9dIFSbMfmX3LKXLcU0
UVvE/GxlehG7+mb0iNuai8vwzFwy/tD71TXKmDcyhpAb0gPi41dJ++EXQJVL
L0OxyJRaMoQu0ZXoNogCKw4UgUNBZRfBLkoAZ8leRr4syRmXjNNC+mOw3bHG
SgmtBEiygb2olQwY4hDRhqnsYq53SABMWstqNOX26xfFdEGkdu9FqLKvwqUq
8ogKLp51MtEHq00NojZFWVfcUkOBD5iPzCSdHNHjyScdT40DY7SmU/Cvdbpn
u1s7LYZhOx0W4xv9o+fGMUnloHE4fVTdSimYiKt/H9yNT2QuY/BJJvlolAHk
asTmbj0UcovD6TkCSeWPS2OvCMOXc5KlizbUk0h1f68gZ6P6+Q0kQevqIem4
mFhoJljrqsaXwYxVd2yAkFlZHme2ibmptwQo7h4pNT/Y27ThMgnFnvHcuerT
DHFF6HLqiAFv2vP077Px9jHc+R8HDDp9EQiUJ48Kl9/9JI9tZZniXj9WREwT
roBTyuFeKLbk7rxqSlrfyiTtqJPZW+rv4olZtOEDh3uRhZAKvWP+uvFi2iaD
w9YStlBLJbMD4qj9hVx/aaChuzPpGqdjLLZK0g10GchkLHulGLgAGbK2rO/H
GeJlavVuKcAUm3PXoFhOEHuGAY/JuVJwq+8Zw21jfmohAmjGOkfS0ZJPZ7Jo
5pZ9HfEo3njRtaHzEcBklNxSQAZzu7thuTbwrnHLkUpS5Mrg0I2j5pGxqT0/
tMbcAoj5xkJ74cdj/5BbPfz6HvccSbOKPETG3DyQpXU5FkNFhcZEWxOuL9My
nB48Jrz77MgYi+BfoLHl+7qgRJYugBsgasGockch5OO+fzRLxYy3p1hOX7qM
T+4YqNgpBTxwpgGhgHMMABTYq47Vwc90O6e8eMQET3vmWghD/VHTLSGcuYlp
ikeyZxMB935yhginYxLoRnvphhcyXNCTEO/Jn8iNhXyca1cyowvcRWWGBp/x
cI25Vx/VZ6J1cTRWIQxwl+3Boizyo6FYjAjFt8PWJfq57r2+YUp6FzLIMSMz
02m5EBI00O2Egc6208Z9ke+yCQ4ND6zYhXU6sf0mF/dV0CNfvDWaQ5haET5O
SKqFSEVOJFKadJxaC/lORA4slXmABAgoaIaBnKKeVKtao+sIEXLfuhEmo6HE
gZINN0pMl0ZUFpZAj8lKhEGxeRoc3C2HikB6h44KAGcwIzNqrAQS0/jlfXh6
iU858bVI4jb0/KasPCiG/Th31Qg2Yzah4pOJ31NN+l5UaDfxcbIPKabnQ0Y6
ukQM99iLyUU+58EpQFd/nrqAgHdbN8LZf0wkVPM/pkbimZFF0+bpjC5dDbol
DJuvt3VoYmZLN8YCx8ZEIay/Ip14mv+Fpmp7WhqVDraj//k2vCBSgZitSMij
17n70fyi9B786PaZ5oqewwZEEI4wX952urnJV8I82WNL20g+icSlOJLRvSOh
EfETOfuqsB6dc83QDjflZO0IwODaDmoZMaI0XaJKTxH6eTqnBCnKD8IXjdFg
j7zh+MJirX8QGxGHMTHHlXsRQc8OGO8M2J0YCFwtCql0TkpFcm4oRNlDIFOM
D5G0UwaLg30xLNjopEaxKFLFs9B7jyisvqSGCIvQ1+s89Zka/b5+lEqQOFFP
De97ncxhZ4Wy2slmvG/9i20+ZpLaiGHxxg8c3B4O4e0qx+E2rcJtBpdMgyrv
ipTi41NGTHvY8zNCZUIIrrVdt9VEatIQzVkWkqi9JkrbsniCd2agwawedEoQ
bZCDNtDS4J4aRY0DtshsK6Ttoix+nPkisLNPToLCsm/bNdThjz9Wx3IwbQwD
ChqYr4q13J/PSJGVuT9RSQBgCi6suvaXNzNNUUzfFw4xZcwb1dhGUpmwFwdY
BxOtoRpW8+oiAj+pOQsNVf7jXr/fKgwbjKJnjpNMfX6wBrcy9TrUgNmFSeiA
AxlK7c2QKGRtGCn/qEj04U8CgugVaw0HYSZ8NanCqFTK/G0cGoTHsV7ZA+5M
6MmPBaNdXn56IJWumUW5eiZbQ85io9vqJGSRQeSqT8LsAOwaNrYkGNGurrzz
3SjByZ3lR3PPyUEl0RtG0s+p4Mpv3VQKYMK0QiIfkMX0zseML3/alCv2EA0y
li3BHZ9nMBLUK1ylJ+G4SRT2jlS9wIdg88R0GkZQgRQpTMtTRh1GDrXGFAmc
tC9Drkw8Rh5rryPdCv2fukZhNzK9W6thhHn74PvSTgd/YJvwnN3B37C/jWVn
fgJsXIN4OVN4RIEaSnc4NDRtX5ZKMbWKZkzHDDvS0z5iffFDJAmDD+bvmckc
DK7L/d/yl466bbsev7T3HsWKRaRV+5UY34Wo2XCzoThAZ39JhGER+AHrVtvk
uLJwPs8heANTZNPzAgP6tHI12GQbyRE5m4IaZL7O5UAUeP/5nE6JJr8u0KxC
CR/2bbdgZtfIVDGfzOM2HVmXousx0+L9S5LK2o/C5d/+WXrqnWBanAHm3p+g
301e7D8Qbk0/PV+YvRsQmXLp05ADJP3buHgfjvcWkLdHmAvIT1S914/W1dBn
OaRC65Dq/a2J3joFU2C5nTOzzGFjeGo5lMMhtpMZ2IlsyE2tPrB0ZKr6S34U
jeQeE0dxXWtl0MJ+6bo1d08GnawWOhOs7CcV4M7c1wNVpHvj4O7nB1DsWjhZ
nzKASdStkBQzt/k4IErpmiNLYO1IYtUXKkzYXwmtFHZY7leDmUbmFIteSo9q
o2R364o1SUABuK1i/hXiBugV8wBYtfHo3q+XeWkkcsevlxR6+aiQt6vHB3f7
Q3ASWeNyn+8PxdQwu99pkN+yRDnBWp/AltBHYw9uGWijdJ/MJDP4fM8cJG4z
YgAxc5vdNRifAy8xiJq+C0KtIM7YSsAVKY9YcJqmwlkiU8kBKYTtzjgkyJIE
teofk0ugf1Y3+l8yrOmCKFA6Zws7g5Iptt+oy45INolQ47vhHhRrvaMtPcLD
0W+X7yFYVIEzFZAiXacc68nOvjsrv35CnjildlW5BYtY58scv+eAx6r4eMSS
1bX6ny25O0L2+eSvxwRR+AEppRDa2oAt1qXXfEYZG8BDKpwfwjyGRjlHa0vh
z60qbV5WDEbB68QU+75Xv9Gn6kgcZ+R1q22cbObYLikiRq9OkTRfK9MmgCjO
NZ+9ejMtia2Mf/SkPGs0OBLxZymEZ2nUJ1jj8E2VIMc2He2pas7QmvUCUDXx
oDaUFFdfkKNYGBkwuLVbOVTv0HuSU8InrGJpWXYZKgyOPE1eWDTdV+iY57G+
32ecn4UDB2JYIMY7Ifw2JdX2RiZ3e4L8rifiRsotwzpe3O138NwrQFg2+zOS
hggelQ7ejWoHPopen4+HUw+Yml3vNcSbX4VRMkwQyN6E2McE81ZWoTterXgW
LvIwbOUrwv7u6snNt2JbpToYOw6sBn6oP9VjkkZGf+3pAeRhqvfJnRwHLkPR
xeRTqBDz4XZQX6TB7I14FLHmvxnVPYh1bAAiK2/ExEU1oHQkeDPKOc7EcQMm
3twjlTLQztp6C+G8ESBhiPy2IhmFH4PYIeXSCa7LFEZmY0HJDYitaZ24SIdf
kTLpz1VMxYY3K1AFgPO0vSfm8FrpV4D4VQ7gbjl5mAl6zZ3BOhbfFhlgb9sI
CA8k4ErrYWbqeaZfpZid54/H0PqWNGNHuh3R+rRpT+9503SxfLeBYJr+6NuK
QjNhDWyxnmZDB1F/vvjYCZ4a07ciY5y7Qm0x+/UMfMmj4p+Gc9xXa7/jbcA8
BrlyTBmnF3ary2kaXSBTZnM3utkGkIaUhwTnQVr9HxVajJTTfrespmEvOduY
4VkA/BswCu3pzC2qi6v9sytWS1Vs9HHOkSC9u+tqAou1Cnw2ucVsYNSF3iAC
H4FzBMbI3zNGweITyQL2wdrK4TuKgkLxQrOJOA+r0jCDdfn91i1VpP86mWa/
X9VcZ1gvsLcKWIH185p0/nnjZpXZ+j82ty2YF1yW7GarR5JfXFKO926C73QM
vjPpso2CmWdTnBwDjsp6tlKSRYjxEZb02Lr0/P53WnwLkCV+QuHFVH5Procd
ohnQ6Adzz50fYY6Dn7pjRzJyrnMTxE1uFoS1TDsIJl0d7/Fv5/iM5/ZGGwN+
246FqT6vnWwZ3HdBm6lIYHC6Bq1/Vt4JyHpoqZsZArCh5Z4o1YqJenagp0uu
v1DA51nN236fqGaJyXpeu9Q3TJ076SQbW+tiqB10FKZ+OE55jU1rjU1qVKTx
0zO8bToHiKcw4YoTEAPEUYqTStkEvkdESy3g0pb0aXHbE2XyllFbaZCB+9wP
TMTbGoxTFRRE1ZtsW6B6WlCoxbq6i0xiCr6nTvOZH8KRGENRpRuGTUlf7YgX
svLMzUhJJi6kFHa5+SPQAbfsIyaVzfD5PLKcQdLhoEDBbX1pR+wmyTvZ43Kw
PnQvbFQdbs3NHYDy38oR4WINQkSB0t/K4SDmCryhu/3RAU99OIQy8hihIUaj
Na3MEcgCXsNTCTf7F6BqthG/lKtMcJ+Wz4FDtoDq9Q7kv+RzFSKMzTJPI6ca
+Y1amw6xZnzHCmiyzjlKInlDgD1v7RXtr02FiwwQo1RvGQ/Nk9ZTZjFif0MR
X3rwOjTlwC0iHvIlodGPSla17+fzjmjyC5NUUZjY+eGnvcwpFOASEVtQnMwV
EwSRmER5b8RfUDXIRAR/zAYw6ZvSv9t9qR6LjYjaJ8T2iRCrAoMoZvm9UpSM
5VZFc/xhl6uBTM7UXl5nxmYFSUnF9xRWywglIrXLpfuistKKcWXyiHjKk1M1
5hIcbkVaL19dVkNaSvGX+yc5OKMAykmrZB491H/sK4lKZX5DtyOoZT6MTLF8
S5aDUmaiMkphuWDbosD1MHO6OeNgk/YDEImFCK067VbJOW2bOnU4pmbM+GFb
4vgImuhh6TDah61kOqC6eQVzGjvp7P71EclTdQPHyhOv8o3+7iiCDUZ1p2SY
3BFLUGR+8XBAYLIPTRiJrjnwJ39oS0jTa3+HrR0VNN3p2zkggJ3RjmHHYGfU
kqnFJ7Yw4G02rmuZTZK+1TNtksxMfv/V+kc1P3zC61Wj4WRp6Ekp1KEsxjIl
lwmO17FQFTdxSfTX0970D8HnA739ikmb+kBurQfNOy/V/azZOUmi2/SvCcYx
wLiX1EwzNhcLR0I2LTy83/+mXglmInH1x2m3rUi5+jK30cEoWm1vkT6pOGoF
k6QQW+PmfYiCZpVA9VrseGP2mnF2rZzttYzZZAkXp2EEhZcGLwpGfC54g7P9
BL5pt9p1xcnenZ6iHpmv2XlvuBXrWidNDJFRI2mcnwoJyzpd50gQe/nFok/D
uTVzEmCtvmpZ0V19DETcfT7Xhn7zdwF+KqbDiPwSKS4vPR4zydtyZsOE5uzM
G8itIxdusC8Lh7S8C0QeP68iKxBsrDhMLb41vti8KHzrV1JUo1Ns4Udxi3CB
vEiwDwGH/M7pWuyASrizkaXmA0w0lpoTuAnH+zbJbAZXEFnZcy/27NWp1WT+
+XmqscJ8jHpJQVjZnF/fcBqL9DpEpBO9cfqoE+y1E/KomZDE+FzNUKW6wqUa
dCHh25CBUD4rmP/JBNXLpch8gaISI9g0gJFpU9W0QkcccN4yQXkDK/9wJC9E
Y0ey56QBrJA84l6kJ7G4DtTVJtbYjbk1qAOWpvs9UItF5p6/nG4VC9USWPCl
qBAWMUQiVv9TPOAUgDXuzhJY3oJq3DNE4ZjR7yp/NA/D1j3MG0bS31EIq2AT
+JRShhW+4/ssLJhody2+pWzY4CeWrWX8rB6rcssZSNKj7zVM54zm1dXICH95
5xbSGjf9S7rQtIycT4O/1Sxx9W1SSGhQrezX8mUS8rHq/4+AeLaATl5iW8HU
75BTzFOxbTqH8N1UFJL4pNSdB4b+mPjK1oLVV8RyrJNhZk5w406UKpzV6WJf
WR7Zt4XKtnr2aOjYEJZCNdnKNZZ5R5AegkE592buwSxWr1ss7BkNxHyDyqnS
DkVxQZD++uqp0dGNFxWsGwg/mA67iirbcizJabWjgyeoMO9X7a1b30ZVbmiM
Vjkm7YDTjK5MM/mUK5gHT7p0zwGKE4Cglcsn3bA6yMR6Qae63MALLUNz0DhG
2TB563zzVYvJQDU462LaNABCIjAnKAvmvdnai5q/The+kwfEFVyMBDcGVVOB
Sy8PpbrJ5ZKdjz/hLDH/neKma6L4q/MdSk6y2hU5yp+URuxpax/FXRnkKDbD
/2FbQLBuYRbTaJEBDKGPbPG+airsL5mP5vfB82r2JMuvOOgK+P9BaM0J2sjd
W5JZO+hotzozVite0WYggiFmqzeTc9MFf1Vmin0MvtAvz7KSPK8AvlN+OW5Y
LIyDPPcHc1hncgZdJcc89rgs+CVSr3BUcauPgv1suBZpdZ6+j/QQ3ulPv7i3
bcF9H7pwYt9NoaBfmCsKiyG7Y4WWQIIaje4Ei+duAzMWPJ9/H+ANxYcb1swR
bUILWktYUFLJ5IG4j0D2jxAPgin6LHx6TKml3hIH5D/e7ysFH/CgvXP+F2v9
F6yxMfnsHE2iQomKwpfbuAGI+G868YhtMrzLrPHbj23eMf89lv8P6YTgu6G/
R92BaC3xBdK8xoU9FOUQ74FRijPci6LErFidnz8DeNlr1sTEgjUwZu9hRQc4
34L6nItIPw0A31kvuXifsC1WL1TvyyaYzmVHeCujPvPv88tfFYVd5zc6HCA7
qbzqRaUc5a6doEemAnCjUpOEOCWmXOKuUIgj9pDuEC7hPHmFxsOBE6+oPqPp
RUJ+wRQCfxtnf0jl8gy3lTMXOWFNHHsw87tUSCybyX528V/wEOB+zPJAK1V/
bjJggftHoK76ezLxfvVe7EsYvLsguHGgt/afGw/KXlFI4dvEuWVWisEyhq6L
FBtdJ9oBJ6oj6TifhyAXLcoErt4udLoLaFiTmlb3wSGeJr9sk9PD7NA7TNHk
Ssxuz2tMbyJflZxzfV5GNJNlr3wlpAPMmRikh5/QemN5Mv3uvFXVWO03FBZI
j/FxgKkQLf4141E6545metajSqtO1bc/nFmBYAAfdxk1587MT8VrqMQXh8PB
khSQWUpIJTDazl0AcDWIzQjnxKG3tPSAVhLqYmnzKlQ5IFpuAL8oV0R9cQzK
L0nTc7xl3SB2bHvPlDsiesyrea6Gtq8qOscHKZA37S+vhl5W5NamXsnfUImv
oK9t/L3iVH3xuqZbj4sWPRIHUGSu1uF35nPqChoHIJm8z1FbrsnotwAx1XfP
gfDM8YUlw2f1eDxo5CZNUhwRUwDF94CK5lrUFuHVmzTvKC0sf7ndn5S5LbPR
+3WVhDHoYy4us+eLWMa/QWDoVp436VvP6TL/S3A7jeVkJXQTuNeP/QNoqX9r
xoQgLDM9OAPVPryN3ozolc3LX30Wi6oTO38xJpQlPB3WzEg2NA2ZSW0SMSXX
XOWhuoXcZQJ+XCDOOaTmYM4Pzg+y6kSe3pSsCgQ9k9B2DTv15BiFmIC1ze5S
7TJeJOuYF/tHwjl5oWOX4ZX802JaUyZlexBM50OzQjNb/POn+WGVCE3C9rVn
a5yJR9s84EhW1U3hEwIVKZJY8YyVvJEqAHuUgWEsH7cIBtXfuAL36w0k1vlZ
gSVp5XjeP2layiE4TIfsDKgdYp9TukiaNZXIXlv/dPHVLYDPh7lUk8Dk93LX
9Rdxb498Yi2IxTHVqVy8b7yLrnqJkYTcECoMbI8M+y86vF+Xi00AexfTYvZw
9nb8IcWv52x3JVeVdZuu6d10ZyrGnNwB8TLAM5qYMw/HubgOtn67xGV/gMhE
PrjhnAKAFevItFUQ0GKq1jfzNqAEQOYbBvMJi4CWaGADiQvgCpXOHULJj4J6
bGHOkmn+CRQ33frMB/D9TO/lUMQAbKwSBStdlcapj59PK3hdy0y8fOpHyqVt
+PkxzLKi5P+mSrcmr6JXFNrysSk1kAfJg23NBhe9d0CgV+13KUah8BgqVkph
0g/pCwX+RydDOqTXVqvmyipJpi17Qsvc0GhHG8p2QN6A9eyjLcSGJUq9Rx6R
zt2A0hHZF8Mpq32oKbGQM8nEq8voDybY+9yx0wRVLU3iTNiIpbQqb0dCmb0J
M8BAT2fP5PXp3p8DE12ho042L1c7oqBig0zuwEJl1t0vjVQ7+0I/pt2Y8WC6
7pLkOmv0df8XSQmZ995U6MNcqnf1DTFlJKu1SVL+0uQsLBKNl+UJFAzaWnYf
ASw7rh0X45ybmDJVUNCxhdPoLBxx7sryuTdMibeL1HM1bDaklDGHzVAVf08d
L/zbRy8jnQ3aRKmKCbuMKdHhlZFMhkKO85LU80OOCs6Ta7DnLwctz0iV3PqX
mp7RJtIkBOq4Pe5edu9V3kzSK4vpAwMvwKewbodB9wSuxCOMoTGKqHEbuGWI
VBxpGAh3IfDkk/mfRFS0DPQwzvB7TgGAWlXbqATs7wFhl77C+dOOzUazpzyn
L+Sfs2ayiG48MoEGvhlj0+fFPsLB1raU1YgMQ9UDpV+qqgUhD6ZfedBSQ+dk
PRtb8g3K7iCA6iQb8A6QfGW2ANBNF0n7NyOVV62b6irjIjiSCiMiLN3XxlBg
mASJ8vsyfFOm0aKa4GVgJBcB5aCWrR6c/+JCymZdZWTrG8FhK4Mw0mSqBldG
UPNXcpy1h71jYgsIvvrCimcO5NxsIOrOlL7w3We52sliPXlodzruXxoI5XPO
IPrXJVboLjRFcBE7khPTZBeD2yhNEKDRE9L+Fp/mVmJNyIYNq50zyUwHk490
GL2VKw8m2IxyvRmHgZNZrhGebYr7RWcvELyvqnniF6B+3BwwdRhTbpjMbWUn
j7wzr+UwkSfhYRy8vcrdHtAlRpEJlcUNdBfPInTltdtyWlT+Y1EefC6cC8xz
h2cIp5K6jzKWSubr1L56ulg2tBjzyTOuDu0s09uUAZmtkOuh61tRGoszBe/W
xRMGo9BTaoo6RK3nnX2WhqwW6doaVUUnPcg41dND3kfs43LARgczzua6VQc6
3ORgp/tIqkYWZCK/e65dBrfr1jSmizVSAaOmVAirbCDkktWans+9t7RA72+/
q/kYn9sGbaGdDmYVmedPpPCbXWaEQ6AcoxjfBLHW6iSVtoyUDYaUO+cR066U
qVkQaLH6tnGr2bl5+5cNVcJxH7DM+CYzzmnzYmF/IEtrq7aLny55CbJr/tSI
U/dKqLXWTDLXB1AHEPk2VCkLlxfKhk1pm7OqDPJDsb4Xk6PaXm4EJ9HlH38+
LuNk9ZTL8ehvIIToi593avh+5tX86IN+MqZxQqeNYduZRUtvzMZRbEeCbcoB
UxOA4pYBDivfDN/Q4biYgwl5+G3dmLqhyLo8johuaCLJ0buGxw4uSWC1FVuY
kfVW5EOz1x/nG7MT91HTHSBu8CTFl3Xr79bhBNh1k2pF+xBQiTjwdpD++7vN
UeCkN1eQI2/fDawnTYxC0+L0MsQOYGueMy5oBnmM4iPtXFHOZdHpwHOGidtz
faGg5pnKkLNnsEgMGvZBFTtcuJpkHOoAkk9EFylRtcsG2Aj2E9O2BDBnIUri
GQI4FLjR7dNTLqE2GE2VvEDrR5bgelPqcsc5ySWdrLEq/5PZjycx5dZlDESp
1MuBy9ROc+PmGAZFbH9mAJIFNU8D7w9QaFY0ZzIj2Fsfjq2+aq3huPsKclQb
mK81saBJeV8L++4IGnWZTMN8GwiGn5Jveqf5/zpgCcQMwCyriiVxZYwBiFPj
sMr8lU+J12emH2PhlxIjT64tss1bFpPiT3CD/k/DV9uyRxoDkD3KBckN25/H
QgxdQYhnNL3N2ug7XN2XhcgQd+oTczoe24FBX3N9RFdh4DQWpaPxVDqhuYxS
u89i9Drfymbqn645nTLNrGFSuH28Cl8+Efqutzfvimxf9U/SZSEsm6YmdqDQ
PshV502YN3F9ICrqZa1vVaq1WQzkDvEktgFDAcpYWoEikAuWs4NZrb3QbSgX
m3lDBN5L4c9YMly5JmWxQQyKBbThDwoJxpncg5irjS5Dc5697PbMefAseYvg
mEjHyEqlDE2nwxrLKlKiuKueXQbP+wUs7bK2cjrNcnqhm5Yvpq/yCE2h1eaq
JGbIwiO7dK7ZJwpBWi5cLfgx7RQuqw0UUGiJmLwKA58f6jRG84k3qoJ+9ILB
S72EDw7CGW5GlWWOOZm/iqMP7Or9q6XvpbieLY+MPdzTsaS5NZ4yKD/RGwMC
8zTTkfDa3MtMpqH4IpWNgZaxoicfUYJjexfyO/fNC4HJ2c+P0hrhG26Ltuk7
LegtKa4E+kXoymOneiuUgbe2ukkisX0UbuOfgBGdr7A2oNODG0jM9xes9+u0
cwK3JQAuJxlGLPwS+co4p2JtPN4Rb1s5MCBQIR+Hw1LiMaXwP1xp2rmeWJBn
FH2e0fDVwNy6UfGpsiLEBgSCwNNiTdjx0QKJkFb5NMe7f99KJNiueuO99YUP
WSocv82Ji2qPgq8EQhAr7hyDcbBy3emdakLrBwPTPYuv6SQnZTkV3McWh9Hg
/jpkRs8SODxT6s7L6cb6XFXmlZ+brWAVZ6mkzuJYXA91slsl87nB/FZL1y5/
NBpYQB9U3r/V4lWP6bau37xwTRPljjSh09cmo0BpEFoA09KpkCc4q68isvKo
22wLjicXBPLGWaTbnRVE/ybb+eBz+P1PtCGObx9Q+Mc2SN9PoBiNClOEpnFG
8sH1M8fjZXpFgC6WSyOqnxYcBpJme8PT7hUboRyHLxfQw/hl+TXXYC6S+t+Q
C1eSj+TOGXYPbsqJf3IDfDQrGvNJ9gfYDpAByVR+kdNXKkjsM66XsJtzmBZQ
whCsfyEhpknjQrQW2y6lco3vqiZeNItKfhEnuDwe+qu8VNV62div/+2fhhOS
aC+Jc5Kb2az+hSB7WQdajRJh5fRfByhoeKTvLaF1dRG5z1XysZQax3A22LNO
w/34HDV3BaKzK1yKN3jqe4xJ8M0HPm5X2boIzGENavg/6OqEWRI7qEQ6BpsL
YmmtwwXWTPcMpZUaie9FwoZorJUKyGqmkp1wZJkE25tw75Tx+UGD3y04O5DL
PPo7KizedosnK6ZvbqqFy77Bmnfj+pxbvScmGAL/VfOsLD0CdHulVsukX2gV
VMJH+E4ZeJu324lUoBy6nCPC8tmkPld7QilkwcuGKI5F5Gn0s65wGGgr5qk9
qdU3J385jCNqCk56sQaG2abEY3QqVwoH4k1e0rlx1P5K9en/k9SH9x5HxulW
cLo1yk5rjPygtspAZa0J6ODwcMm0jL5GK+eusQGPg0Av4v46uBOhtXZ0XLtG
oOwwYiecBrwIKRlaaDSYd8XfHAdyG0elx1cCaohrNnfJzgTzc3iyTgv/L4WB
SF6e7Hfy/88D5KtKTXsNT/zyX085WB/FC0HJ1I45I6APuSWDeOTrxLH34HeR
+xHUn6B/xl1tGrawdkDGZjB49f5IY8bqej5Gf6YzPtN4EqfiGfN1KuAVEUv6
XakrB/Jz4OWRdQ7BBV5oj0gpCYVNmk3xJSR5DOxhNi7Hl3d6fWeoQQ1XlKGG
fJ67WHqxAwNc7rOcpRknmHPJ9s+b7KXr9NdI+yYzKPSP409cbeaUbSGBd0F+
bHhgu//piyUYJEnOAkZu9JNnjO+QU5C2H5O2UCp9qVXPFY24GW0U8Lai1bFX
xv1f+JI7KhArdJnf2AihhqDehiCDShT9JxgxNOQP7SOTsph60sUlKAUKczI9
N3sOq/LnW5vu/yTDlUWkb4pfJ0VLo/0kGNIzfqtF5WhfNk1x7Kn5c1Z11QCB
2FeiyLiDE3RQIBwpwryrqwLs0RJ59XaI+iEUjhIqGH+RP2PJBev15UYO8/1v
GG9Ie+9p1SsCMwGSfhBbpBmsTEF9lOEBR1QMt9PCwc7kkgzZ//FM6NfTneC9
Rur585iNU/oWOC7RaP+u0r2eXXU+1CBcy1oDNiPIlenf/4vnJGQg/XywDigU
zpW8Od/yJOIm7W8yjhPxz6j7Y+p6+KkCYagd9pzY2LV9zYojsKN9YHIHxbgg
2GX3E+iyvoDZ/8e0V6f+QB9NxmeCWFrtmuRI3vD6YqcpGM7xKRjsnbKBJ1Sx
4zleTNR1JEmExszHHjeWbPZGcAppf+AYmMRyh/+HVt6rfJalaTQNra9djl2w
5ep/ceR8l5UNjsKksSRoXNQ/iaAXbwkEs9IeTuDyaOTAgDIPeZHPIWJIJR/V
wTOK2t+tjlvjIq7NKPEGZzlsC7eCHYGmsWi6/JbsgKkvzJpygzu3tN2tbOwv
q0E7G1XQsbh76/Q05LekbhF1+KlNFRLIEcS/IPQGLqBvbLuRAV/F4OsbN5pj
YPFGI+otV7cSr1iRaDoaJ4cjEhlJa9q/soX4gABOvu4Vr6XbauQK10DsJ6go
LXQpFzTHzWAWycYmJNAzd662va+nTi+3R2UlWA9D5gmEoqwuKrErEDabnIsJ
H2Q/8QukX/pKtr0Lja+VFHHKzHXwW3qe+SjQmZKpqpkgwfh4XW13FHaeIlGL
ALqsx9rRs2kLAqZNttN1HXh1E0ebsr9a4uEX0/suSn+Er8rCm3ESRPZyRe+P
FsqzRXj/CNmTebGbmZhWhu8//oosUfIQsZqbPUGMBbysRFIkYk0vRSwe7vm7
V3/TcqRu5ib3W+sJj1653TGRrsAYKUuRmtH9JhcrsUSHfd8YDAFq8VTsSr7G
TuSr1CjETq5ieQlhHOycTWMyh39B/R7uEzC1SJiQDX2yUFtapyQcQEXrwDMX
mNgxsaGqKvVyhvhRp/vZg2NrpnuNgaXkxo22LjuectFiNpzc6E/vB2el+726
PkDvWQ+Kpd8oYEdXMSM448ckB46Am+YztXSArZ5uG3yguK8znQj/qasrEVsA
C0duWOiY+yWc+l/g6CA/dmT4b0mcguCHUtvS5GxUqEUbhgJVdn8sl/OAa88W
g0q/e0HHthihUpBd0wm3YGeWLDrGeaaCf/Fn2bPaSogbHLlzwn1Q9ekazwgb
8ghvZqt3ORsHGGgPbIkyqGBy10WTp75MuhweOv/zj3C7UJEdtdsWuTnbOV1M
PqG1NDdpE4a9ybaQ7ZzvIJyqumzhxOs0ZF1Caicwy9eKZ0Vqy8Gmx60E48eY
T8j9JNWa84x66Zl3TIrWsnIoVSDbJ1IsI7AHdlYDDcunKiEl3u9A7fdbiwDA
ol1NUzNrr9oKgvVzONMvz9Q87eHnV2SDk67/ZdLz3s0P/jSHvXM/HzQUdmhT
ykzSSuayFIHkTeEWAbyPKXfkBi3oSUGs4ZzXPFulYW+Vjjju9Xgqs68S6JiL
KhPb8NM3PI8BiPjZMcDGlBLuWDrYRX10VQm1vFMp7LjDLNDIjMAzyZ/4YQWB
4VGxXM05iRSW5nmaQX7uXwqFsbIzDeyYkTj866wA///ykLpQ5OU8x3SIENj1
qynMvOm6LkB+csBqpn+x/gYuBk20r3NpWGj8MBFCvseBkQNGBCtiv2X20tA3
bXPD/u28k2FPCyCD5en7+ZzXck6VG5BB3U4B4LOImILH5j4cD/pBM8F68W4r
LwGU33QmjmM3T+Za73C6n0bgXkiLpGg/qxlyM9D5QGXsr+8GfDwb6FE3fAJv
U5mvfZ3NCZ9dBs9wAi+uZyxniKjMnZ9lPcwWrkWjWc9Z4SQ3M+tlzbvbOjYg
thEPI266UBfqyDp1eRnTDVQxfF8Zm7X0UxDJ847EdrkedYPaO+cvGuIUpYvx
6/4fa/iCCaxuHm+JHROdcfO0SIExv7THTXHXAO2wZhH2C4SUc4SHS97Nzvey
0YecM7F0zIh362F4Iu7gXED9T0e3RmjWZ0wckQLSYCfAgfJz6psLcxfgSUh6
s9jqIfbMKTNsoFbSOmYVROVoAajboy53w3MWcRz57hZ/6eFBwzUjsBlgrRJY
gTPOEfCjMmVzvOCke39+qUalRAgEnGqfXQAYn68xPGc7eBu0TtirVuGchJPr
FH26WXCQS7sP0hKzlfylayjr3NzYBcmlejtU7Sx/2G0s0RoUM4thrrzd6p6S
1FrrKUtgO58L6Vd4yG3Kzebt7pK1ggW1KtbkAkYFw4uGUKeW7s+UdX1lZmEO
qts0IEJUxfH10hFNC01TMPj/CAAatiDXv8xuDDiA3KXkuiaHE2cj98qyQvvC
Kv+WZTlA/WdU8poDcGcVU9z5BIapX3Lia+SkGYpVWK92FeAFS68+OHHGJP2l
TUt0ePfRMqTNnEP/y9+OLRVPrwPL6ZQoOd5NGPcpSaM66giX6hJvmsy0UcTT
AsUBrGXDdWVIXDZisKjLUgG1GyEMkqK9ETFXARRYFbKAeuW9Ew0WvWWNCOni
gK6Bgvwo26WTzmbZaAuApAIphHdO+hLm9fkJG/75jW7DnlZxaw3JK1ZSWp9n
cn/Fn6OgFfBpi/wqHJlTTpGtLGE7bReMyPGgHsDo/wPqKQMdEenmrqk4Erca
i8XjKIdg5GnvSSv+yWqZnzeFssBP/kaJBE3bNxuRf7vobfqXzlGlDr9wnoYu
zPRMScL2us41vAex6ZzrtlcNryvoL3uTMPeQPuOxjPCKGLA7lg6UrgzF6Aj4
lvQg6lK5LieEf/OwYclEjGUdlnFZ67LalaPe+VsS6eg/0hZxBTHuoayZRuDE
50wKtX4sRek3SRBRwHTQxbckQLjHU8rCTEkvu4EF449vyD3dafw6bZWVMp6O
IjloLHPUCY4GXUfeo4czi8CSDb118/sjVydRmQza7l/MY7XQhQWP8upFul76
S5qNwRvKxJDO4adBwlvP04h07iUd9/6YEH3UZoTYwTITmvEE6e1MpU3JCGug
VArsldI+uS8eTvU+HPsEj7QskE1F3Pq9u3UtDqYRfX28tDJ1I3aGTEMghGV4
ih/lnq92CuEzdRbMLcD41Df+erHJ9Dv/1LBz8cjYR9emMlepnpaTm+jyfOyt
xySCnOlVirJHaohFQ9aPBphzQvL/fYVDXGoTG4IDw8b5QwntwUL4Y8/lXV4m
U0q0RkNFtM8/nnk/TEc111YhrWfXNjX2MYxUckCelB9t9FgI3ffJRwnOz9bd
xt1t/yMmfl1Vta/HLN0/iPhtP57aSXaRV+R6URGvnJkc+LGTdja/UZsF07fV
WCvqiFytJoV1xaJNGTVVFD7JrJKf6mVXngqVq91STl5anyrS3ByiUZ07XjSy
svHiMR00d6a1OepHw+JpbnRabmH+Y+H8glYQHmX8ppilGg/sEaOwrWNlc8/z
Sy5az+q5GixhV8XqVsWypfF9tK9X30Q1OIe6PnE9vW1/NVyXP5BEsmngFs9p
qWcJCx3owX0Kkr92pqvwQxuGB9mwlM7tb1FlfcDGiP1oSLlrGqr6R6Qgbdbk
sNjfmljJiGWbjcltu+KapURHOSP3MRqKWgYrfqGqcy7edlz08FstUe6bptu4
5u52dTLOKZZTI28lTjTWOTxmgHJZoi/Zd11Sba2tFAmyBM5pvlS/XlOBrdtp
OQa1ikoC0himVhaNIsRlVG0JDzZJzUJlUYmoxUca5iB7lELxMcTSCnQWXmgk
eZnzuuCCrr/xgQ3XL0M+2d1lLAfUzUhsM5IyqTQMPNsqz3/wxCpdCy1IxdR5
BBHV9GZYjufeB26W8TSnD0w6qrmbw92SWyuCvPXQlibg62pfS6iO9ZNsqumx
8f/sn2Sx6ITme8U/RR6CT6oW+XzD3a0oTNyD0L7Sb/gjru75E5TDY8oGKFqf
KXl0FLD1Yu6GeASPcZ5VqNhJy+WejC4k58uCNYCpcDBMvI0NlN96gpeNe/be
pRNyZXZQiPZO5tDo2P4whfjq9JL76BuUmW5hC4yGG8NsgCp2qlW8wxfa/ayn
hopBOB6pHtBDKF0hg0PM52uW+yUm04dAKLU/v40FFNoMx+WmaI/r4nZKI5K2
0r6cPfdkY5EMGnxLuV4VBLrkHWYBHnvqSEQWV9mg0N4fGots/71fSniY+UhY
z/LzcUSNDj0aFzrKmFIZ2fGvZk9qiSPziRvDNv32kY3OFdUb3Gt49dZzgrkM
o7SypGzmBbIlgkar11gWYANiFTYW7c83xa1+fd7epST33NCEjJHobsi4Fyif
hD5vMmF/RLevA0LMtXWjmeDM3eLei0LGwYWf7MVYNCcEZhCddp5UywqXHJs1
IwpJ6je86V0kQoDyA1u/kYwKk4liXE0+1Z49j3rMlcZqpWNxA2gaIbRUptOj
+D35t2O8DGeYX6og3un965c6h/JRvRjT4fiYAXGe3M8am7+Xk836ReAVFJyZ
EsoRsZKFUHDTs81Zo8T2r5S3Ie8lrn1tcrDyLXx2UL9oqZWhD2am7K+t3gFT
zMFqeKwbGfDUubw3o+JtCG3Pa20SbmVgs4mgRaMlt2o4/v5pfyz07CHEdQaw
OV+AZSUIFQ4MsSrc6nVFt9YRrORfy0A510KZmHEpRFwbwnDjHCON1Et3w3F9
U0sjqWSze2fMUuCW93a5c8mKk5kYpJ+1uT4ihK9z1nrWeOW9n0ZPlN9yeM3N
J06bvZeIhDvGzfNUHdYp2oYsN68jHZ6+ODXodQO5F3ouGYmR7Y60IgStLK/7
WrYIzsSnDSZ3rCMpjDh7Z8dape4Y7q8IOIltWwMyipT/GtC/o9Evne/fA1HP
1L8RukjO+hboF/TSN0qaOI5tiHbXl4PVXyHGwFPIR6gEbAr5la0OKwgGFdBB
0iyBTa53gdNqHiv69+ppCylKwNr8e2RaC9o6JsGT3BF7/Jy6cxIouvkWOMNC
59WGV8Bq+nVCTb47/4WoUUCrP8bHx+h5Ud/Ijo1cvQnht1wt5HkeBH7DNscK
yrKNjcENW0l5PbW8dxZYguiyNh0FbVJNS1dZ0AbK/i7dhbjLBVbtN+ZvSJsP
JInxCz4Vwu6Igit6fvzgCvzAIdSz+C+B27NvPbWNdJb+CscdMZDC+l6WVfJi
nzEGINHDu1FoesWK68tIEpb4KCpcG39fQNZTxWr8vYq7D8NB3DqvOtgNuTE6
RwPZ4cgMy00Bv+JHyfPjo4qZVNTNX7ViOCdg1En3BTdZuYDnchTTYQsT7A3u
iogAcJ1QoFzy7U0kSVZ5yGspkwFpfcpKdSYImEdW8NqDOvi1SnaFtj5BHFA3
AVfWqGmVYdlvq/TrdTIBPs9mb8LQqKcgNQyS08TU9iXSV67E5kqyxYcZvMHs
qQN8qriH7RKnwaFmmTLXy17VJtKgXsqAxqbd1W6u+4VHYSLmA5mZlloEDFac
kOM53deIAY/Aj7Rjp1cCapQ/aSsSrq8HyhYrjkbJaJ1m7BimDK+p23aMSMNe
fot+JTZv0cOfZCwcuzn831Z4u1VQCGHhyZxu5wDGCKHm/fqNvaF7QLOgLI56
fqPRwbqaqUhik1SJvUfPo69LVE53yF6sQTLo9h455Rh57jsJhhQfuBYWCyUb
KfzGjf2sb+E/F3UYYq2HPMHblS9Ja5V14DSfTh/glMq1LczGrVboFIFV3I9t
OWcjHziygxqeOIfcYkuLX6VbafSoYmMic7wjcLa4aq8NlXaKTm5e4Ce6DTKH
hEsGgW+lMYfYbqN8rBHeZe1fiUYcZCc+pdTqmXdGmhvZrMa1O0gej2wpmxpQ
YCAQPlTR2lGA05UmIiaWZsE2mPivGUX+zJnx6AwLZBG+l/nA6qkCBZQK29UQ
cgYE15u86mx0y9R1sKdxmmY6+len05G3eDF8hRTBkd7rcSekmVCms14RIg9M
9aMvMMulwcvNqX9MRC83y2v/DXXZG6mPbNtU/GSBGZYQDgSTFpHEacXOiX7w
ik4bx1yIxJUE1gjDi7TxvEUSlD59tZGY8EauHB2+oyKZ29xhlUnu45OTntj3
SlMmiH+3XtqsneTwZ4oDaJq4F/+VzBY5MsNaoivKd9Tx8dW0y6lqpI4x08Ja
sKzPyvtpjQdSf7MKQiOOxRxEWeGFWsSdAzoe4lN/mBQfp8tm00DgRT7L2I56
YoKmOcyNWssd+2nTAiaxberg1FKb5xhX8FUl9knQsfccgAEL0EHD7TKNEwmZ
vx6aqWeuxdoMJL7B49BEOwdVQ/ts2udSYZlcV6iKn3W7LglPWwxFg9tiicJM
05RKp/6JU7R+KzaU8aEQFYXbpqT5r4h3Z7ZTmO8LVdVBiK/mUmhUQ6R4ccLG
KjeORK8jDqIkufP5GFYXm+ekE6xey2LCm0qGgElSDAQ19cPX7uIWZfLmxy6c
ScmcKdDD6UpFyB/CMq27jkCuCACS6kgqCEA01HjVUO3cRhz0ENvvbif1f/eJ
igxH5C92Vk80ep5B720jnz8S5rsRlArzvsaOPlycrGpL/SjLvKTqrdSuH608
P8xTIxNQoVKaPepyDahfmD1U6BYFnkn0BnEBUL8/JHc6OoILLb0DzNpYowwB
BXiYmTVLM7/x0OkGYTKmecERi4MbWefj4d87CfdP8XuJr4edlYh1z4Q0WZf8
flAEngIvAPZYHoYKTxsqrxJ7OieMM7SQpeLbFefuphuwydWCJ+S7OK4AXg5/
wkQK4e8/UAoCyXUI0MiYVw4qHwd2fohqjZ4zJj3tkSUQ0ZNXN7QoLvjNVp1O
8FolWzN+97rLcvu9ukNl9T3AVLXNT+aaiL979YyytrTTPl7aMmq+ooUZ4Qe7
zoZnppKA7zOWz8eMRkGcodpk1lNyhBDV1H0K9ghHcmhAcGaxLRLjSZjhd+fs
4sBbGKAbo6Ixec5a6No5mYoaifbqMBi4uP6/nMFS36ewpCeSMXEDh00lwzjp
7kpGMiF75wZ0CXP7AyQtANGgqcKjM8s7OzIa/anGrlx7TZJYdPEkaB1c3EW9
gQUbtm3kXkReifN8N6PNkyFUW6NhO/lEcPUO4gQaHBnlov2QYqdVDgACV31D
P2a7AWs3KZwD+vCRj6HIScVkKjrV4lYpu3ijUTcbw0kFP/mMYwoR60LNFHy/
YgCw13VvtEIwnTqLhiTyPkZnleATd2mYdeyf9sV38uJu0oWqjw5Q5zicmXvc
Ofnb+pXs3+RYyF++EfptlCOyLWw/p7SPoy04dJXCQfwlFGizyjEdJ+lBK6RX
CbkZXBaR58pwwjebWwOUkFLrUdYqcqO1Kux+M77mmp/WbSyuMmClw9LKoAce
gN7tXk2FfYBj+aQYNU/aE8tDMrhCTKacLFuzYEfHv2Q7Kf516/OOWIxwEJBN
mtI1GerOgKw/jTtGr+KbCh9clbrlsMbO9uSkE5qEmCJWz9CpkWTfS0erMDzu
xrmzkytD9S7wfQLin2IFn850VVApcB0TSrZKGsyU7IzcKo2F3oWU5shDsZzv
HVmvedPikLKhR+E2UPiqQWHSpkNzLdMXoFtsygna9T1Eb1MsTK/zpEYu6vqE
NGO5PI+6bpCFYv++slfOgtCAUdYtuLJevXvGTi1tjGIuHBjimnGHdbGatA8y
5zFjSeZcXmB7UB3rhBDui/5ZkcyR0L5ygQm2lmVNvYZiyORXRcYTTlBm8u1X
qp6TT+wDld98EV2mDdVdNIf8Qr+8DFs/UwJKIXmcqtNuUY1V7nuL/htc1N2y
d4fM7WP+Nw89uANL14C5JcgzSiEcPNp76VXDsVCtSILgDMpQteY5wNODXqm/
5qabWzSOqNW1yvysvSpyLR9+bFcrSJmD0+OKxZUrFwOWSD54JcfDMyj7VB5t
aT4HJ+11cVN0ZevMW3hdF6zLo70Wps1W+o0kjk25JARoBRjkWKlFbtRUje74
WYJDnBoFnDZsDfDPhK+rxQrflqGXSv1goF+yA4BQBL3DsN1LsHqJ8PyNGZwA
eQST6PQ28lemaBBC0nKUCdiPwre7s8RC8uWQkr41HZpsVVoScBEG5AiZDC8Y
6oYUdQ1p7xYVYjS6OrqoWfytvj2QsaXxVj/up9/sTPXQ9nk5yhyxWBIfWwbo
dazsFmoPDs2Wz5Hh39jt4csCt+snQXzD7oj8Pu/Aera2B5EhNeAstAYO/jJz
W3FMDGyXCptlW+G+JdxydlqbZlY9lIReu7hyR24eGET7BXAio+LjRfbM738Z
xQkMRU1MCa0qcvXmIZmizD7fbNDGUNW+3d07E0IvFlpyQYaGiGuQOqgARrwW
BgAbzgZaf2ZyT8x4SU4E+dZ1o6nfFMUzvCSQULz+BvRPRl2TWqLBYxA2y9lg
LueVo3rpXESE+LRitsayNg4KpPbWQpi69mpd0kQk3sgDRuOUDwoG6iQOdSDv
oB0F5PwxaDlk3VX+OyxbaYPhlRF1kQBeMKTeXCYsxL4TZRdkflvUnWbBZ3IP
Sa2xVaqGGFODMFecN/N2Kl69YQe842/TSukZKzlXwHDJgqqQrsYclaw0iAaW
iNDb3c4GeKZozUOhNv8nOoUCpsXlbN613R/5BeFLvMk2cI0VO317ppEvtB6H
Me6IjP/AvuyESsMyTIUOMP3SBXTKWCkwqozYdcyYTDuNOhoxEe4UR/583WxT
dcdSUAsiEdC1e5Lrhs2LVgG0wg9fRkKGMlBUTxWh2zHiajXHwNDi/OCXPrEM
sUFk1nWglZC1J31M0pe6I60bsZ6GMZtu2oTViHxTsJmJPwafKXpuaDYv/t4Y
Mel6YYTJ/9eH8XamSaQtVU+su+O18EbzEV5vrW0tbeSaVakOr03d9/pFFBlO
KK/QbS1aROv+oTiTKjW8Y9qpZdSGxefJ55Yv5DxrhteHbID4F3nMX4liU48h
Lx4hNLSLxe5NqlsZG/6DLKFnD+fCI7JqYIxOpvahytMbvzH5jq5hyeOzEWUc
Fk5U5DvtAFUrr2KLnCWBLGEQNDR4Y/04oXG6T0H6vW4wOofQDLs5qg1E3A+m
jz9yHpSX4YnG5ggNwnh1t5+oTWXsl4gblQm/qD/VjyMM8sCK6xBaNDMsC03z
u+itsxae55QaoxSvzCTN4cEIr003OcMWcSUnnnz793wZ9sGCbVKdcH3NNXHc
GEQwt1KhOsA9znj5zFsswrBpQdA/rYdqrfe+gpAdxBTM+Y8XVUQRlV5DHoUl
WBjV9PGDQsoS83nepNzaNfYqMSs5fXBUMjiqPpjzZgxcCVDka4t9yyNod44f
1Yf9kQ9VHCMrGvrZtojquFvREtg5W3iHvc3T4ERU82c+60gmy5LSPtI6UHXZ
I4wqCaA5jx4ggFPZ//Dqdgd9ZWUaFyOWHh7J7mjOVy20SA3il5VKT7NDJfO0
nPqb3vEDGA37DlqsqfsrKFfPRVf5MAW2Ekda1J/20vt3wOqVoQNC0tcFowvl
A40Za9QLVeKqUolNUWiXUXisJCncuKesPDv0UH7y28jZ3kAecVineFaTCAGv
cd4iaxeSzBVK6yk56R/YwxmVCCLnsWUI9Fo/14fAQR4OXUbrjJxjRv6QzFTg
HNq+rVELzffofZwDo8lX0LyOuHSM6LpMzapKRJti1UknE0JC+rTkrnsjgz7a
fYuAZKMpJzwxY5hrtEvpLYJHESOn1B1nlhB8M1yuaESxfTy9K7hJPJqxZgk/
CagsiR4vijrOfyCAtIaQECntPw095PKFIZeL63myPwQsAS8F5su+y1ACXkyE
nDsCo/1MaX97kc9P0C5E1Jm4fW5XcwjUNJHrKLeb73JS8F3r0vhfTsgC2utT
aU3z4JHp16o7hLg5sfxdTq/5sUNWgJ0+1QdHIVRrYFZZb6Osg7q/fYaC+jDy
vuQQwi+nDG6BYNp7bYlF2Fg5i1Cj0S1hrs5OPef8syinkBD9IYj42nAk04dg
Ew1ujU3H59c472DDDo0CQLYE31xyvusNqGLIzfq2c2mS9SO3pWjyrVmdhuEj
hZDaUMrnXkHVyQTzBkfnXz45POsAKph0n0YiQ8TwvhVLVEP/ULdUPCd1Hnd0
EzhYwh0VTCW5X+HhCuUXbtKNw1hDisL4W6zXO+f0vLCByjagtms+DUJ/vZ/x
ukyAkpE0Ms7hStbuvfhF1mPoxtsh5PoWM06+G6hCUiXtp0gJvoQEfwKHmLe4
Zj6N58+TP3OrDKsUMb8RAur4WRX46belyOwbd4qL3kU2T4tXqw7kMm3/rBTN
HP5zhsc3oeH0KE829zdf1cydkDKUmli21yIBYfbk0qpENvexWNOetIE6AFEx
EzVkoRUeCjFbb5k9WrDKL8wS5hFlzJ0dORrLPpfpNVfXXJQqE0qtf3zsZEIH
GuIkD5zG3hYi8cuMgxqRSXy98dLMVngGOniBY3FDWw1lsr1kt1VekEOWLFLN
GfixTl5laFCmGceyhe9KgB/u+2dyyde0NYuTougOa2wkkiL/5Hsop/1/3q7w
F+GrJ2+h2USN48ElV8D7cHfAXC6QzeOiN+qf6aA5EOHpjN4Bim28NuOr0iN5
se8evHoSaic1b6Nc9bGuoeWm6Zu37OckrO2DLc4DN9NPxabqKIa0Nd85b+wI
Yl2zw6YBxvIQqw/KRYqF7pdQKREPfkSLMoz/yMDPJi2yim4poWtGVX3xWhBN
+NpoJWdv8Lbhe1JU96LUu1biswtHT8QfEM6Bs1LtmiS8qKLJXwnBRhkYT83g
Athya5yupujUPz124jm4wFgnMQ/vmhddTOVvpucGKSRjCkHOP1tv82Ble1fr
UIKKwqn8+83mNWFGuKq5juJ4qoNh2opN7zIH1eYAazwttpBjTax2XsW0u+Wn
Z+GwE0RGISODRy8KuiaXvsToZ5jSyxwzg6znks6+dWSNP3H8/GW/f8bo5y4f
cAc/NSvo2OMyNhJg/r/riZRWRQtcgNySM4y0408c/AWBjy3dG/z10YJAEjxm
uyXE5XTCGyIIM+FaD5/7Esp1Pk61SCl5tJBJoNG7wGKMl+CcHEzrQ/fAOMy4
yHguhgPuuXhLoLI/nxlgDiuP6TaSpkJf0MqpmXn2pPoVMU2InP8GFtQWZNbF
5REqnSzGKwsfmuE7+SQ7CN8D2LQxaP6WB3B2p6HkWnuqrkVirkMG8DBY7eSH
jCCbk4Mat/UhBF+3YqUv5LZ9YMtf0p5ZGjdjvuwQLMV0yPGHXT3/oOzWABAT
2YrUtAKv2Y5uFEAEFPYNdPjLCsHH6bPHLV2/1fx3AwOCb9NAOvfMw5LRNIdp
o1JkWuF/8ga3Va0/8D/L4XXY/N51csvufWRwPxB9vMpDj61107+8EA9E//lo
+gtTQqx/+/iAXBAT7GteM3a8sWbPB/Pwxh/Ir5lj4TVGHdAylBPDv8T9pf33
aeCsiekfjc4cYs+EmsR8GBblxbaLB2+5oM+Zu7XQm+a0kEcDYGmyVBkYafoZ
/plSzkpQ93Y773sYYAzSxRy6Thqudj1bINgkD9jMhvLXsoXkN/bNjjC2Parc
ftJWawUXyFCAqL8Dp/Dm9D/rTi7wkjQMlqlf1zkYFI3UrqRfTD+5h8M8gKxj
V8SpRQhLwwgE/Y4KlPCobxk5HF+jLtgdwpgYpKBwUtnupNRORBIXPgcUksTm
47jcREr9jzs0spdkSB0tKxJZ1ehdFtqk94KpS/QvPrEC7MWwcrE3DZL20Gb6
bk1k9VGIIP5080bE5nsNkbm62ztU2Br87OudzeTd3uvLD5+8WxMNGcSZluSv
cOr/pQnJW3ZX8z4/f1u3kwSOAdCHI015jMYIyMP0pXLKOOtJCbjqVCg32f45
N3GlukBn6Yzqifz/AeHIQCk7awvGQ+dhz9QEuMF7xywK9rmUp5unHSj8kNsS
zEWC+kP68FTPycRO39FThtBA7JtM5xOrUzSxKNee8pXrbPBOBNH3erAtqiFK
YD9ZJlbPAcdIhI9xn9NkICuE+70nRLdDXEAhoNCnqx6aAP8mj/YFftXnzYnz
HcaNoODTsirjqBR4YZ61Rl6Vd2Btemn2gMhUiKqKzkQCTiGRMnli9gIGVhKk
kSX/xTzFYtnmt37Iq1FTSHbgfVUep3ah0CX1F+3nVcFc89eRBHsHsdNw7cRI
yiCOq3ZLRREof/1fEJik5xTEhi64qE+oGcTlwNdCcYIpEz/nqXnEaNGEji3M
96bzPT6gFfTcRc2FvkLDLbWPjxs4i71mS5SQ7B2QvuP6wJOjRNLlad+gv/l2
iShxd6Rf+1MDWoHObG5/yML0HE/uC3aMZOEoRWzY3NNtoCRahyOtaMCp4lLk
QzceuhOEk0LzO3gA1oZKzw3cQdrw9m7w2pfXghvJGIZNBQwiSQdwCQZw/0Lx
S6LOopqN//2Hf6gFmPUZbn1GvIz20vZ8nFmtSKOzmxSHBDIvMAzptt1lye6y
Wg3s4k9pp20MfBce/QBI+BOdBITdMhzOWY3ELcGYz1cmZFN5d70xZw4sGXiJ
oCbvOsQPxd11z9btnOoJybzK90fFXQxAy1jGAvmJzeYSv1+mWvyLk2sfyj++
NmbkqKB5fPtVUUFOk4732xNxawri/NVPdLn0DFVzkQaEY9X6kh8B0QcObBQ+
ScJ6n5YZRisy+MHGmkGvyXYntZcat5vqFs2txy7cfDtRtrtJ7OyrmK+TObSg
9+N8WiN1l3wB/F6AXCCpElIU2zacmJEQjwHfWdhSzTdqXlaw7s+4YGgHzujB
G+Vv2i9P7Q9Np02VD+Msem1P453rg5kX9iTlIGDswtRvKsey+H+6YBtZMrDE
fzsidKCm7GfevBO0T0rvwizvCKp3laRTphbyCN5XJhxFD4fv+8XJeSWPTmbM
3ZJAjLXdZXXdWukGaSEl4nRAc2dI/eRIBgKlc7jsrrfq95ANa4O6HYdLexgx
4nr+AyNc+u6SqNLzbPbr7cENCSb2fzxwa6NVwR8g8R79rlXZIu7kgT9WgmVa
oBZratwCfn37UnKiWL7C0bKmd1r6jF3aMXiqsiwm6/sujDXXzrVxJUE0yhPs
czK7MTXAxPHjb0G97VEPk6h1FSLUz59jAcTLKEtXpzmtPeHDKad9RoOSWYMr
OCBaJVQ8TZ0JxXKIGrLi97DKEbDt5zBdrBhszv+26CLOD3YLLl7IvXk9GB+Q
j8aB+80tpCGKU2GRiSu6L85dBl7WnsNbw2a26lYfAbO0Y6Dbb7P3PfScW2Kn
HSP/+jFyMa9gTo0mJeVUbHhkuD3SJOZpmlDRV3lowPfN7mzU61yr5EdMZSbb
RnyWphF3FFHOhBWcjASZUeMvbbILs+Br09/cXqKMxrWM+i3VpTJNlG1igdYq
eFmaK1F91xn2YQ1CmNU9mNIR7k7g1aDprHfSs2DLLEOacX3piovHSWG8ORT7
zVn9EDoHGj1BmqBfgy3TBaU7HFsY0kSwtGt51fEgnmzAQ9TvBwqh+jK3sD2E
MpOf+/R5hdtHtCqrMoml8SMTUJRPBWIopyB99ROURbbn1txXdx2oGbJZKmrz
5V6VlaOmCMJsKPxNPg0T0NynfBTvL3GlcwsAv2xbDfJaLoi+rDYVRqLJrwnE
64qDRa96qUzXDzlrr3C45PbfhGSZ75zKlpU3EBfKiS3Fh8D9a5q7KdLBD/GP
neyxrVVjqBWR6I3dzfQQsKtkYQ67+NQz/KeRIBIE1bAcYOy8WnyB81Q8lRim
KMxYB/fn9P9ubxtAs+FU8kvCGw1woJyaTkqtBCWZ/4bpNFv0oZqEyONVERLl
ZduTZ5Hb6FmHlHYGzBVeGjY3qFYi3aqyAs3ZmxwzgIfcB9LPqj96ciBYu+ZD
ri/7RaXPGJGgtwabH9D/2DAaRGHLBgZRm2lRLTZVrVBWP9XSheBBvYvYt2us
9BOyMKME6wa5wTjfGbiBsS12h/TLJCE2kB8Z95KK68IV83NC0mKq6m0BIhhl
VaCEqHn9uDsqd/K/U4i9VUlIKbaIxlffEFvDajbJu62LEt1/XPaiLAo7/ozG
5j5+2ZziEFDxNltUfLXwYQ3vUXCCR+q6BrkDUECmNT4TRGUQktS2LoNsE5oy
aNqStk92h1lkSEGE7iZjA3z1JgUujGIhM8/xIXbbYibwi9jYjift68erA3FI
VysR09Cv5iHyvbf2TWcDuPhvdbTCRFU0+UJQCWydQE93ig1gd3Gvb+N2d5Du
QeddLrQ8VsYyHEta/vIfvf+N9ueEDQH8IDg9oloNjtHpqWiJkhB7wpPHsZbF
EHFRCZeMV7ueZ1mBexiK3EUbUtqUqb7FCf0/o60E5lPGQEvIfGv4Sd1i8xGs
8IIwMXqZ5A+FD/a5fMatVxqdr5L+x0nwrwVkumEpoRQ/f7Hj+ynLmH/4IbrW
XeZeazl+d79Jn0bu38xBtFsRDsxdthL6nFg9dixecOrE7D3nroVoO4Wn4Zng
j3XSAwgzpAdC0gDxU4J5sbR3VopwLmjBDg2eJVNLjLc1ZAO6s3jmw+MBDKaY
xpwHaiOblRXQhUIChkSFMaF4utBWGizDVJz1LbOY8DwNAidg47B/AjOTeqa4
BilOFa8kpHHgKNVHZCPp+Fnp50jfCG6TOxrOmLgQZOb4wVkC5CXYOgC0mq/T
WCAbA3ryItgyuHvgPXfht4EWy72e19VptRNZWO4bP6cDcmkxtkyv+yWPkgfS
6hNiEyH4I3eqTxv+5mrBFXoweRa+D0TsJc35pJ7UfSM099XoTWZoQZ/uu7Kf
XlrOCBdrBRlCrFf7IStkvq72B243BbO7NhaDeRuLIqhl+87vBFa93gh/1BVQ
s5O6lEA5RvWCvehSJlASdH4g3QRu1V3XwJZII3jztm9lgu7Nu5z+9KFvrebg
4Mxw2cjCKCrsWoKitHNiHpr+IhldnAsYJSmoN09Mfi4oIG4DKF2MdnpS/gGf
kSl/OvaGMu/1VArlgef0ZOrlOs6n7VosmcEXtxklHI4RpSp22oViIV3GO3P4
QLEG6qJoz2eZam4WkOapeFD7Pne7/QQCb+87KdRMu4w578BrtW4xn9OSSS30
C5s5cVki40E3EGQmsgl0nSEduPqH7kKlEOkIkywWtROnDBvbzEPs2uj7vvUF
Na48eLvRr8yRKJVFgfrokdFIhoXeGeI+AVFWkU0mdLdJMXeRh4X9Nd6ok5Im
EJX3blkNrhaLlrQZdZgoNCTdTR+qAj4wYKO3EOhsJv8OpAdogMHN3ulBw4ya
otIVcGv2AKZ0fWwvHg2v+uQ8261+5EjUa+wvRRY2zMUj4LXq/5q6ghBrfOjU
X34frjgjCiPKES3SMTiCmcxf7O8mQuSt3wOBxd6ZlSzdCpoDaqRMeWn+e78l
OvWyComKQwRyoqM49M1n66ziQc+WfEjWyOA2vdWX1crxHW1XbHq0Yc3EdqCB
g3sGo6ibP5x9sD46L39ytDybEqdyDFid+p5a2yVturtxWC8svq/ZDBDbT/kl
36TY9Uyw0a6gOavlSFC29F9FzG8rCwcPocbjeXcNnWXlZbNpWPP1sdnA2PsP
rW7XqwyrfX48U/pdQOEYK1qKjcTjDv9WGTAcT0Bj0c6ieQAQJnTEIIdVxcCW
LXN7fu5Z03ej7tmdW5wP01E7KyYnGmUIymVYdVe7ZTsBRzuxb2qOUN4Iopla
Is48PLuB0j38QdxmiGzY7iYM/lzmAyK4KVEGXl2T1SuaE5/e2tGzc0JRzkt2
OTteA3od4RxvEKSrm96HJIjv2LCyrmoub0lD8A3zPcaSLsXdT7/gl/lEl5jg
pIOW3FTKNhcyD1yNSGh7vmAPmkcoqg2GgD92jkeU4wAvDGYNgBDxjXhU+b5l
3rAWE6tXjaxm+evJOxJERmxzb0TutTjvXskj5Lol8IvBdNd0ivMDAx1Qt5pi
OF0SMCH2bDDoGvyYz8NWLFSBDbUjdDU3uavXKZEQe/WBm/4TZZRonrmgZWoz
XdwblGfDi42UDWMb1KQQ41b+TrSF6yic2nhv0lEqj7h62RucELQYbiGMixt2
/qbjSmcxXSVmpmJya5HvL7X6j92j0nA25fyCnz20KAbe4PvitcFq+ZA4+++r
nerk9nNVjJkXHAsoVR5gi+T5XzaxCVXw+DmUuTDRLk+sQt4WSN0bvOPbqtGk
7b7bX/DyuvUKS7uZUP0IOxvg6jlSWdBIjWoBmq4/rTikveaMaQaA4xkGQG1b
OQVxvj2nR3g0WT5WuwkUZah+5pRdgHC9G/nS348k07gXNzLqcwKwQZDx8pVw
L3BjlJu3sBuXxluvVOklWw8LUyj2iAsZdfrfDoYZAfF6m/is0A5GpCOX4jyk
DxJ84it9MKRDM29+lhRDDpuoJHDKocuyqORTdoFKw383XIZJDDjmGXEEKGQK
IoWMKfILbOrYM/tfRwtwufMRJdKdrf8sC5GlZk9RcXzLApKk2bGGpgiZ9zu8
fbeJP77Qvr4jfN6nDS/YI5xbvSr/5sJRl++jaYb4lWwv13ZildLxes0Karqv
sSuHhh/8MC26SFNVZdB6tYW2cM/5T4+cefccsJE1HkwSB5f17u0vGcszzYaz
p7VdoxoSoypzupDbMnfJ1nea6o5Q5ys4yQYQ6pnBIS6KWC2fAxdmcLeWlj8R
wdNBCgXYceiprmzF/Nkt6EddRSg/LE3ttulyXY5P3BHNtQjaFCEliAqMeBLf
k6MLWvajyC04oPXRFPGMe3bMgWZuxHqd7+2tMOJ4k7hIZdbCZHwljvFjR0cj
amTpFfCV9yTOcwxDRBT+fCW2vmNQtDNjwlXaluvCx00zw44Rpn3N/c81OIsD
k11DIB/E4uVC3rOkW880PxQ2qRCNh8ovq6DPHhCpd+UUHeHou9zslS/ZWTN5
eedTklZFK9843+Ohr9deX5JKTDm/D4PDkfGqmG1PwDDR+W7HP5KqP5oQqHI1
Er2607BXURP01708JGoKI02aoqnEvOiNfOwOefatxNDlY/P4C4h+S8hC4L1a
DSy/eitV9gLZmoQUic7EngHHD0UmqOND1tUQIyQA04olwzgISR69HO96xscL
rH9f8P5g7crULroht/GTV5bUXM3/ZPMQs/X683zAR3SvsHYKd+s4Y0vTa5/D
+Gbl0ovEBgDE7WxwQYS+pNsiCg3o4Z8zMAIfdZGbO3IzU+UnNMg6lV0XfUyD
0/i86o5UKUOYPGOqb7hvL6tfoOF67MC8NzwLJP/mGnKbc/ewGdYLLLIiDGsF
OSyXrAQI0B96m05lJGcUUkJdo/1Ymi3oltjDSnIBSd1kAxfbiTdzV9lJcDhl
9jeGI38Uz1Tn3gZwwZlBGXNnnHOQcht+TJvka4J/DMfBkFWcE2MUywPrABdR
Tirc8jLQHb1YEv41SGf51dNH4kZqRq2STFbexiGcjCt9Kkl64k//mCzKbIV+
FgP34NyuwawWvSQn7IXNlGbQsgTsGRiUFsoF5ohuFSv144QckNa90dW7Ujw7
ptlWTwvbseUw9uWolwLfZT/RA1hL9AgiYDLjW+8B+VLkH6XZc0atSha1drkG
yAHW/pYe/0ird7VXjVx9PI+6i2Zw4tdDSZUsBvnyJsQUbMzXciNkWg+V3cvi
tte65OdjyzDnAgGGkNlkmk6g1ry1lQPqsmCs+dhL9AM55qs6DYZe/fbWytxr
pYHKxTqp3rdvAaXM4aoSLiGV44AmDrU2bzTSWwD0wqzuNLIK+RXGZOj0qrAD
2Q3DvcqPfR/NUy1q/YqAkYECa9hEtuTmbyS4B86Di8rAxkaymg4uBAgrohCo
L0w6w9n7Y/OZh9PbfAp+VrGevhhVNlzy9QO1a3Q1o7lf3p1XDe8JPtHhpA/i
N/8uTQZDaqCysj6G1nowXShALlm0NClnq1oxYjH97OR847SiQtp5Z0GwmXLV
Ii6W1dZGrYS6D25Hl1+d1ewla2aGChSGE6SUfurpsYo/7xouIUqOeR0FXXl+
drwttjor8s+ojtPgF1yCXIedzN+vQYnaAXG2bxnCjYymAaY5X2mpSThRN3ER
2joGsgz468Hc/Ld+sTrGslY2fWoyi17Jcw4jYf6jdu4Xjbzb2Hwdm7sujzYZ
0L1eo4PmdiGX/g+FToYozM1VKMReQqzzE7YxkkS3vPJ3DZQjwYY1xqjdY4d/
g1MMN3QcpyW38wz+Q7wpGtAyEwlqSBJ1GDUdkwYR7/o2cwDep6WN1G30BI2G
02r25Xw+kzvqH+ndiNKeMCp5YeSPqgoxylrkJLHqC88CJHivo4f6j90C496l
hPZxJR8RUFbJQ878NvGqnjlX1Ztbv9ZvWYT+xInZysb89vVhhcLFpnmYNsVJ
/gkvZfqYUEnWHso2MMZX+dZDOSn+cjqYAYXhgy3pQh3BLuRgTsG15Xx1IKWJ
BMz8Tsb+xMEa5ElI7kobIP6WNQYVqiUv1bZwFOVgh8cyECv+o1VilT0UfUlA
xfSY9lAzHYX/uBsZXPtj9dTpA7ki3QRgNc4KUVEVjOVgNM1XLdAdZKpsyAek
6GRDzcANin5I7w1jy9s35OYd2tmnMFNSM3pWFXO+tnYHXQaNBjvPGwxvJM0l
fxbsXN0GGMnadMeDIBl7B7ruvKU0lgeWGrU4SEAMmdwVcVYlL6ykehshUI74
f/2op7dAChDx+r06fKTribPvOELFDssxxqJhcJ5qdB1AIdlgO4UqnVn5duGi
vBnkrphxVA1qcU8BceH9nMuZJqaDlVIsO2Oi3qtiVyNfNbPLeEn76oN/4SGq
+LsF30bmYVGsX/vLZCaSVNCmlyxhHi7HEAEFzqn0KujUA2OzB7q5kxDr3nWj
f1Ps0T/diZSNcEqqk4MD4dmJDDljm15rZZdZBtsBEIt0+MCObyMy+wOFg4fU
Vhtu/AhTtQLRywSGl/GqsQXEYvuAYq7NRHX/vfsyV2im7/Qu2GkRhnYXEwqw
xSCtfplq0t0S3bgXj2C8+O92W75YUIJc7SJPfNRYuehdO9oNzDl7nzpk78g/
vabnQDpVFifAiZFPZEAS6UICERr3Lf98pIKHZuSFoBpy4QFO0u9Y7a4nwLMD
XHw0V62mYnQp9Clq5BvwntdBRq1j7vnOkTO0SnGp3sW/XmCGai2qDnuHnZQf
TDS6B8bHN1Esl5Xj31/D/ZQ3C4dkh2ya/ZhrAizVegAsrmE4BJ4BEemEIwz+
ZkR3KIBJuFplODvh04QWbERmYSELeqWlMjdmRi1hyaZ7xyFF5+qpeXy/Y+x4
tet+oRn2RMFdkupmVXG9xlzxISOIuEvUn2VTAk/bd3DYgDju58t3m9Ef+Yyq
4AAjY3FUXLRba3kwzwsf6PldHuflhCXASQz7hbSE/CqxTFEtNynx3zDAI93U
y43CuhHr2Lw13RFdjuJbERKSbRsWNBioygEWxa7JKEF6d8X3YNq8kzvL79BM
tlKBMisFd5s2kheiC08/nioshbxXmhar47who8gfV64RlBdgLTxbTByCG7VK
ffS34JgxB7FH5ThT5gWCqIKxry++n57oION5yjI3cSKY+OFeMDn4/w/sZQxz
P+mPDRb3V3L43btiLuVtIHU/GQHRteg1dWTl2agrY/Ye9yreH1Q9HHI4QTJr
Qwzmloqx9lq1VW9OFmT+Wkt4MmIfirob8pAjjKL4t4Uho9+cBL9iO4BHDURk
1WjnxZV8f5Q2hgDW805oA3zPueB08sqaGUIxyYH3FIOFpANKPqFTzwKo4P9x
Xzvh3f6ifXzCIXAyTQfC63YLtfItWRYI6QaOEaxy/Y/yKXdKwgw8LVIGD+yf
rjd3pP83G9iURdClVo7IKyMaKBAMHDVuqMicItnEZnOiTms1sU/+UZLssg1j
pillinh3igSQnWG7pnecbEwr2paIiLX4LOEiKyxJ5U79eEvb/Tc437lwPfyO
/e/U44gKmaO5RGiyVMOPfg19M/RioL/sR1e1jxRcYVcHBbNNXHl5eYSQkdEn
X1Swpatv7vribVhI7FuJqlqGMncioQ/syNdzqA1+nENNwBONbgC8tqR6bMBQ
gU5cLXp0/ctj7yvJm/OPXAmgz6UtKRAeCyMHzuqtqZM8ApMdsaEkTztoOHHQ
pZ7zSjs7oHHUder8kM0iI3Nwj/zzN8o6nH5ja5HX0ps4iTORAW4ftj7W1ysk
vPxhFE4gYjc/VMtHcaq+3BNGPQZvot4RGbxR/4X6HtmjGX30ySdAUQS6Nm24
c4IhyUvC6UUV3i32jN+JNp5VtvQ/MGHUEifQK4WtMVtGRVtafx7DqSl/BP5B
1NWIpFy5Eg4mlGO92WooucGNi9Okrz3DHI3Y5RXijTCHCERd02J/5fmwdBw1
bWuXTMga9BcAK7Hs3RYNbgJGaqX8OJUNM4ZWqzSCChZe+1BRkoCpc8XdxzSe
NFdCmFLqKcTYUtWJtI2zls/nrp0qXBQ4sqFuu5fZTxUpusA+X2POkl1K8ebF
DsoZkjLwPiZ6/0t6OFLBh9GoEVDAleUBSC8n/5wM1EFib3KFwHJg2fsNX1P2
3AI2MaKmMhLMikTEDjWaMlqVrDThapXga6+ThMmA2vd3c+Pd4AbfjCD+h/NF
20Kr4CqperlmZ6t4ZGajVHZh32NHDaYjPKN5w14E/F/ZhqNSN96LOEwcWTBW
dw12eOfKm3G25UeA8Db52msHl344kiFmwi9YZjTqF9nsnhgg4dblhoB29izu
E+D3cTiOigCnXirpkw8lx2NvILUJcEGKzM7sP5GpLms6JRBc5YzcAr5ni3Xc
LxDPRbLYdjn9nJG6BdS3zWoJehZL9UzRcPHgZC4lLtMbL7SpuS2CaM/54rme
qmTicz0qZXv5g19uGtvfbhXVdFRlj28kL+9OrEnDr+f0G2OvTBWF+orBPFFh
ngahPIor5sRJxcNeF+F2QDzmOlGtrveYDo3+ngx4C4A4nfXXIPVOCub6o+6C
/+XXigOKwBg0M8J3M6trHD1ojz5gy/4Ns9fcwy/lPqQnV6GlaIPKUVmPWI90
oPyk/8JzDROTbr5TlqzIweMorOLn6MX83+OaKxTjoMGchJTShIpsTXXWqc0Y
BADrJdgx4zIxl/X65DooSAnIqLg9BDeRddYoDM43Bg7GrzIXSX6DmvQ+iueo
pDK3n1BRFTAPxsTkaZHUu4y/+CNinOccqEvsPWyiHf+GZ3UDpCA/h2i4YuEr
wSHw3qlV2om83I/fQPKFTwGrKED5qdmiX8Nw4Rnl/RTthBNj1sAaicMskd9k
AXmhffZ9NV674oeFiIJzTPPL/z5SgrfRFfvH2Bree0l4t9HuK8mF1doe6BSA
v8gTS0uczD7OLYYpvBUiobgEQNuJOWs5kWNHWRtZ24C5bfdA7k6aQBe0oHrw
P2qYBpN/994cmFJe531iGguBCykvEvkt9ycYnkWEDpSITwKblXJaN/o5sSo5
+FD+/919x9odBAdUnsKFV7G3cDkzyhJRsbu2QeqfCLqOXc8Ag+Mc7otmrH6v
Kn4cDeMsyqVcmNn4JTY70Td9A9w1H20CQv34T4QwTZ2To72n7rKVPwGW0yjN
O9JaH0ScMoxiezBVr55lI6FEhJhNuuGrNitDVAda1vjg3r72poXJDZgxNNj9
lebuCqzCMDELH/3JpqcJkph54vxZWn7pJP8NoNwJ5yqqASPp0naofXff4QX2
PUq/Z21vvlxz7FM/b25gdpnkW4PFNYzhulvlzFUUgXRRyLovO9hM2XVdv90D
YSapAe4BBNThGMYMTHtIFZo6Z074XV9jYvU2gUOOYDGY23ML8fNE/86iF/dE
kUDKy1bq4S6zTjjo/A0moEAC3hjinF9sBLd4B6gzTCbcsbE8154/jmshQWyN
JhLs27fR/L7285JnNPE28TkaS/6nz4Mq4CSfryJEKN03tU/3oLAoqPl5jb8D
JlxqGsG0pLlrj7kBBZBbikXAX1vmFmpl+cX03URVwudY+Kf2F+RuU+0+dX4c
0M5TivZ27Xqgu6NzDV6xps9xQpXYzB50/9uXkn6vUuKBvwDdJI9chF+0q6g5
tSe8q8vN9+xvQPb+mlcUfbhwgkV8t+/BnOXpt6MVbGAvCj7UMAuWpBgi6d0r
oIa3I7z2G+mMmQH6Y8txDmUYDEo670PeYeQxR4iiA1pZriwxBNkcrJWDGb6q
Lhn7taQwu7gAEBvCaEsOg9IjqtMiD6H+fxdvZMZ1Nzl6Slq5hmwgf7Y4kyGr
BT6iQJcfpo/JRXLmwQyJj6e94HIiIKfnXn2pK5l3e1mtY91lstOhHGUnQUJb
8DF5GDmB8GC7NYYvK0SAKKGinBPW/p6LzAQd/lYSsQH6CHic56gTjvduEUUn
qtaaBE1CeaVnSHmFYF7yT96P0VnlK4up+bfYpPpmhMszqzvccuM3fVKUNwAV
ASsWFJIsrqXir/Xbv8ikZkNrQCxWhjp7Q++6EhS2JmfWC2dktAyQr+ZNSyxq
o2VH8WQ4xwDQUYbnko/wG4zEy8AD0GbIidCqGDWHPH0srz2ugIs/qIJNOBl+
CwTWPb0nlv8PQYLe7dwXZITxkoMLBfvFH2aZ6CpjRiM/1NEtr85nALhh4egu
jDY/t6KdICBqijuCrNALjheLT4sWTTJZ4pvnoAt06s3ipa/Mu1Q5FCYZdQjh
qppid0z8N3jNXPenDgGx78KBx/iHEVRLHSsvdxbCZ/r3bzs72nGshSreLHs3
7R5cKOGxuZ1y8Uje/2H2g+1HjlsOstJgO8u6djq0mPbG4UM9RTofilOwjDfN
QRRRCwBQsnr7Udgfu36wcR65hdsRfdVPz8rqkawOWEDq1pi8OIJ6BrP/zBEU
GxJbZQsZw/vK/tLJxazfmD/5LK6SXCqBmg2LphKNatHCXP73fMr8XzJbVzij
qkj1kJma8us1omDDY9Ro/cDZ8nej2bciUkgNHhh9fSiYDEbpkw9Fcp50qd+O
zirwuVdfdaxMnd4/n510YcNZfpYMV+6eZ5Ku7xkJAtyKgx2f2XNyFnkfRnzZ
VOsrKG6KSt4jrsBgG72cnd/LBPt0ps5tr0CkRYjrZRy27MqoPcsU56IdoPCB
mFGIoBMz8N77d2ZuL/mYs3X7u1bFhmc3eM/43TGQYdNVx3s4FLskn/ve+2PL
pY6k+nJip4lCh+hG08lrFsHqb9m8r2iEnEz4EZel6LiKAoD3vbxPk8xMCP2S
68Ru2320LaHDdDl7feQz+6yHQIxsjaG+WvXoS1PrU1K86xlLsN8om6X0d9tV
R3OEAXFYzphUU1Nskp3VoI1E0awgOW68uSTamOdBINDf5qeOhMROA3gayF2X
fQVcnzlhuHvGkZQIe6PcfvwLAddQ9z+D8g8lVzCurHqa7E5k7AXlRnafgvY3
bivsBW8ZJBApZAoidiYf6SCCf80JItioUR0eNuD91xhL96WaXiArOBrda261
jK8KuVh23+s7+jnHD1hrVMWUOicyTQcV77pCnd0qysrKXFwFXRcetBq3JotI
Y5zeNS8DeGjF9lwGuOGmFcUkW/y+6RWKAOyEqqSOwlAl8FGj6vYSaJZrtaf5
RP5N+BVPSwuRMM+QDsCZrqUWa+cJ4w6iUpKUQcF2CrViNszaTsXkraxxZgd2
9zr2iOftZuamESVjTG9WJ1tFlNDY8TyN/9+62AFVRVsvR6EwwdgCWwrsMe0N
+UT7DqbQKYsenlgxjcsOlfayJhGaJIw9cHMonqGrykmPYq7Fmik6LZ9xCnFq
VTXHR7qh2ZeAbUsTvVqvDlVBiyRn83s5kXRbFkmHUdeTX3vrlDW3n8dRc1+F
n7UEz2+Ylq/j60Q3AhWCKCOGwdolK0byXaOgjtKPyJK8zLPt7iY9uvpw4m2z
4SrKo9LG1230rNhqSdn0MN9qWI22DrIwED+mZpIYPt1LiCZNz++yi+6dvhp9
D/mGynLGrErhn6hFVd8EWtWiGL5h4NBvTIa48/ddbHbh5s9h++BJrKnOG2Xs
kw/yGrs3x14BMMT8JArlIv7qA/8sm6TJRC+Z5O8K4OOYkti9lmMb6ROcNi/i
J/F7g+4V45eY5kZgoaYPuJh5DWfl2hoiFwXy06gXxySJjGSFOMo3JcndA31z
4ar9f199WluBSI+sHQ1QF4lpUiW5P6M6/xbe9icpKoBLG6iJe91d5RADfa7i
HC2HYECgV9GWwQLYnARnTAHKlXkJfnIZ2JQoyOhw1oH8ctef7beZIWBrFDdy
gOIojW9NZ++QQymDWdWBPDtCroAO7RrGonOKhhJIJm1P5n8Os69IeSG2mn3r
bVIiuiDqKbwh4/WjoWaGugFURwfC3OwrAt9FPWj9ITG7FJVw37kzg4gGVmDr
gb92W54lemPdNrvkTv5FaX9sy7FBWLYtivC8OGFWqdbTH1tjrc2arohbyNQV
Ka42a/dtmLqWwc+1GD/X/3YEp4G/Gn4CMNgEjcButbpiwfbonwC0vDRqwi2o
58j3GQClpdiO+roPDX8zVRWUpJZEzfqWg3z3RUowT1CynS7zRBzxu58gaH60
zukJ/hcTy2TRpuMNN4+2D3N/47HwFT3NFwnux5fFaGylTAcQvdORiH5sT8ak
LNgz5b1ylTtXtdx/yLBYOzHQOW4azL5czMXId4TGkIm4jGj4sAJqkuqgRnC4
efjHz9zEBaAPQv1fbTFYF7Th2qoCum9D3HzgAhMqTqIWGxSf8/bL97BcYNk9
E1UXyZkYMukqUROqkeFYEJxvI9uiWEhofUT82n9MruPPX6g5ED6T79OIDt9t
xmP7xi4O2F5OcSPIGU4Nop3PG24Uqir8R87tOp3JFkzj7uqkDSR4AxWG6R8e
ndPBOFL1355sfl6aI8sTnoTsS0clxubpYbAMSLkhsekTecm7tit02YmJ0H46
kOZlYKesLvmE0WF5YiDtNQJWORfuzOwMadEqupNBN979nr4QF/+n9l5EuQLO
alZ27MgrEzt3urboIMMincE2qZZ8uBQpJ/1C44761PQ3nr4qQZIQzd/Q09qg
esT0MdLJKZTK4sDczXlw1y1vQ080e1DgFvj7Qdf77i7/wfVYSdOo9ut12JDa
5fzsrlBqtd1wZGaghzb+q4c/ugTQGIgiuwO5fB1kX0s5RCxnykrPrXS8u/l9
W6nl06pZm/KJ3fdK5BWaV0136tGcVn1Foo35Rzlp9dBOJXjXvhOJpmMaI0r0
HijuNEwpTr65xgQDXFQi/BmLiKhe97TgkPTHuQCPuFYFQIlleed7/a+DyogF
RU0m2L83Z7/SiLUlwm+V8QkkihPyUjVk+6EwjjpG4aBZFmpeu00TrSXJsfzH
D8SuP+Xjs/i0qgPSK/T3ZtcT8ZBEGzNax4r8fwe5c9f5FLpaTDE34s8NxWSS
/vy1ADgu0kt7kJdwwkBJZSEsGpQ6Y4Vii7F/fPWB2k2Us3aC6vnA6nUER3tP
vUecSJueT7mlu3YhfQoKX0vmljbXmedJ+AsLGL0YzVZfxI/jqE7O7u4nu69N
5U5XgOSQtBgqti77phVuYhMArPgXwsWhNyNvS+UXcQOmvSVugqgSZzK8YrrX
iZxA4GHEXzC3xfK0JAgPMwVLeFWauECPSRR1vVnktIqEKyYEp6MqeQ+k90jd
sbDVcMicGmr9bZMrghUfIciCaejkgNYHPzaSjDJJjzMszd/JAo3Paz+XTMQJ
fQAnFCG8WkyzmUoSZzog2tNlZbhGXRp3M87UhRHcZkqdKxETXQDW6rO6gqCT
D5OA7HaLiYjDGkzRJzY2fqYB8G2jwjEy1pacz/azX2l7Y8pPJtBC0qiBTXkA
2J27zsSKLHBye/FEwXJtM2R0CgJHGbRTCeelosv8BOTykWdgqBw8L7WmnBWH
xJgLJVi0UAg49RabmouwgFNbv17JVaTqNx4FdarVn/9N5MYCS5Wl6PeAF+kM
b3Eh9OTnNYPTHpGKrpVcSb1bXED2HT8Lc4yilcC1opCjjYMCEKRKENbpVdYO
1aso1fgW3YyrdP9l6wfj7NL/CdtMd8ze9+wz/QHoP5yOi7dI6hfQGAw/2WpN
r0o8fD+SZGluz2LfTsuyGT1n4Rk/ZwBbFQ5MyNLTfUuPO9Ii8Fys6U24PwqQ
mu8JN3BzPdyJSnnkExv3Ks+JLiLAmprHv0ItCrFtrYKux5TS9mYDx/KKbCk6
Wkj7eSS7ZE1y4c4ni8IHWPcCMM0I/eTCxF9bc5uDpdresHjBb/6Eyo8ASh/I
P9ybbO89KIMnikAIHjv/lAxe46CL4O1GvkHT2KElPun/eFNHS2LoaayN1yn2
EQd3UUQBWVFty2lSO1zoY0GhrEAd0JZ5v8T+AxHBJsvi5KpwuvMq6JGvwePL
W2vx8hgXvN5wKZdSWX2NQpvT01wRDGRbH+CQW3mXCNBsVGmsN5nRDXP5YnG2
w+ULZNGN8ZwZfBLh09gZq90DWzmsg/Mlz2c/mTDajugg9JFpYzobeOgDkao/
vxKlyF9lF41EtGJw0u7ljS7ti+gYoCLUiOdlWTZlr1dgxWbomJ/mRz0G6pLw
EnGRo8CmLvL4t1Q4QLC5XGe5uazFXrT2y17nH6+tAWgMML/QuYlkUidiPiIs
/t9q3ayVsaSKZCvS6mixk634y4eZ5Csnt2KO7KNWzctszn0ThiHOg4HcEdI8
fNr/3sCDJ1W1yZhA111wZbMMznR58CpK5y2wTnurCXaHRJFhOWX/BAHAfXYY
HnGgXRNb4KRSHmVwmRAivs5ApLrI4yGhAKB62y1wbsHENUTFiVvPdoE3DelZ
druQI+WbWXziIiU9J+AigD9mzh5ZKDf4W54ymjznMUrPqclfCAfeYVaZqyRL
MsHn4WqQad3fPi2ktFd/9Mbc8LAglrCkHqlN0jHKCBS4e8iijaN6/t3dhhEb
Pfcj/7bMFBN4+socFjB8noJr1WyK60hiH9ag7ahxtFnIqvGoygqWx63Ez4qV
0sy89hUJgCb720a2E9nbCVAqt3xRzsD0mA6V19/tq9ZvwnuFkNOM1fSD2h5E
eicmQZmDNIadX27ypanOYsolEbegPbA4KuqHymmGcTv2OFQXXVZgYViimFYa
rcfKCSVUYrPkEO676VZAyS6viyoYPsGSCTcgQDvFUVn4PHNVgU++p/CsHIsa
LCHkJM7yuhYOAMk6XhFyOPKsGboideYaHgEB/dSEK3J0FXUIxGmLqvD9PeP8
do0yvsR4p1I5+kW4MawBpo/PaYVXwIkPtUet3eUOssQEfOSP+RMQUqtDiIgG
o2i+4deycwoWAWgoDfoDzaFCi7z3WxB8/cIhvgdy/bTvZOwCAqdL4LBJ1Ufp
9arVEXhcC4NzkhKHDHgLMkjxcP+U411ypfq7QlGD/rLE9mqGC6jIlbhVXUn5
aJM8Bw37Spm0FmT+HoJzT479/MoKKtTh5osJRwCbArSCjZmKl0ZejK/PsTBA
JTqTv/7Ys1BNZc4rXc2mq3bt35WRHD/0dnL04uov9dTa7S3LknBRJ2jEFYHk
qRvfObzjcKsr3//XeweRh4+0WvjDdnBWdc80OCjBb5Bqb2PZKv6oZum+i02r
rf/QmPcss6D3+SUzqLvoeScS+YGjyeE/SRexK0CHPlM+fcK3JRK8qgWbQXMO
oH7ymqp/iTaEPE1mbm3Qhb4QQGtOtthWQc0eU973yao+qEK0D5PpbJgWDsdp
aVeVyN/OWhAI4vxr49omxfPESLPDpu9nr7AWrXPiwenS/g9c0oPVnhWD7J3b
Sl9zMqww5vkPMjDHtDav9UcQJZDX486CKzZOhr7wmy/HaWcNTzBzlqcj6QZd
KtUA9Zg7iIzsdgwedZ+KBB5UaFe5Vv0O0LuLGaI7IrQpzUG5MbQ5jd3pL4hC
7yj8TjLWp/xRKMfYuzlefMJ4dUT3+5YURG4jQ76rUaLAIaaIIp/VcxxXTGDs
eVBAYZDFOVFZCmLs4HJI6wx6pLRwZ6Lo42HInHvt7lmvHkBXRQ32V3bt6faI
z2KyjdXDAFFEauO6i5EiurbniClPTyszLytFgiHEh1mUf3EXAOWuwAANCQL/
GiFGpx8q/P0LBYCFwcA2f6EUKnH49ItcBpt3J0E3edT/7i3JUZNClqcVwWQs
AhPvXCm6ldr4ou2H2qsR5BnjnStme+tzoZ/TSl0w8utK97Km/MmJ7HQ++p7L
Hoi+OWg46I7g/piEu9/rOXbfY/QqqoQQucGloXzrGbvTVoQWbeGcRVBr7WPQ
8a0UiibbyH9/JgiEIiY02F1AXY9/kR+IngZ4QDw9LpUx/ZsH9p4dKC7orpxs
2Y6i9i1MQrn6V9fJfOK4JVH1rNHudzYKhXoVI4DvnQKDhd0u9Tk5fH7IRGzK
N/gvX4EJKzyfpIR6PGzEq+8bpUEvbyb5oJh4r1jCpt6tOwwoPILtUqwgFKMe
Asn4Zl3pDar6U9dVVezzEhdOCzveNjT0ZWq3esIrnqvBAQYp7QOYTeazOj93
zRhyG6nR41w6FPMd6ELzZFAEWL0zFrsEoFp9kPKITq4tR+8Xe/wHltK4FTll
EfgEgqwBtkk5qGr/RDRpraxH1bYbxCxdofN5ory276RNCkepgJYd9ScjQhND
y8+b2tUHFwTThMV9zlFwcE+FProlbjIMu9UvH/uD7CH2jIpg7134gu69Km52
rDHzH44s1XVc7Vaw7kPFla5Oel0j7Be+3WVnSmsE8KwsRCpw+duShGFbQ7eE
nS+CruKZbIB0IKbG4ScOHcwrpIGeGJJQDakxWxe+6xDuoyHkPxu2qaFGg+7J
RRVOoRfn48kkofaqUM0LW0zc++8TkTkU5jSFKKx0Z5w1/3iHyK63IbzqCw27
XuXnapPVv8dKYuBFTmO91Sv8CvAyIZJ9c7lJEboYr5LfRTcVEiu5MAKfcr5A
z4oOLwczYbof0ifzwrmlf7HEEXB9xrITY5D9C5WsvyX3UEhD3pzyz9UG+gEQ
Std8CgvZ7ytNfc1hLZpnL0Dgu+248mBnPU/sU6a2yichmduMwyl6rQoFdYfu
mYZ0uRu+NtIMnYgqJo6kYIvO54CzVYvREofk10w5CuXu5cqh0+EtQzZI5FTo
YePuaAb+FKWaQ448sWeXGabueco3F3mS0O34h/uW9XPoHj3kPT5cFNJwJzi2
7JK7lwNuKLYYYHCI2fPakROzNTPmp+RsV+2gU7w6Ab7QCPYmbGFBHF43KsXK
myDhUv18YCpKXnF3ZPsvKfsn9/Bo3MW5ieOm01wxU3L+Y/5lNBRng35w1dTX
vvsMevSBSjDFvpb+TbDlr6guJ99zSxCKY/7dL6nt2xpF+R7GqtivQkMk6U4A
Lca6wpSTkwCrkB8k8snlyFUMOdoJY4ZaB4PR17Wf+R07dOUUfarghIduJn5q
u0sz1RIMFFUOh/vNOvD/aK355yl1CUqTSvel7BTaY4ZaE+nA3lUjpbFJcHYl
G8cCojDtvKJ78dg1AIAFuePlmeXKDB4Wa8cb4CRuY4dIOjKuwa03nthYLoMl
2U8Fd0dUUEzRASIQAWOjd0nr/Gw4+alGVtIugY6/pj9kvVlKib4Z+L4DQRdp
obshTv6eDZlqEb54kbl58C6cwn19vZfqarv41gLYFIeo9ulmhY+uhoiI0FlU
WxbKsuAxo+fGMmGg4+FtvkUM9PoWZSZ7wLNw0vT85nYkv6yNd7wAyjm/EofZ
t5M7m68UQvAl17Fb9/K6AbelvRoddqIEl2GhBup6EsZAfIUYi54HJhGR658R
jPfoj7Bxw9Yt+FvMtEsHIbRZhsRUPwzMcw/EhKM/yCOfu0HHkLNH16BTJi+d
GT1EHyzLjTNo5PZB1Mo4v+5WrQ8NOzXffJEToiODGPwl8cBvD/fV+TgOQmwc
H/TRjdgz5hb2/UzI/aG3MkylNQto++HV9DucXxoXgvd5/R/YjOOLq3Ml+x7t
JGMmUz28SxY3yLaeda8iC53VoVuvuBoD08cvVtJrB5MIGXR8IQVBUjNI7E5N
ng/YVvzdTDptp2zvxiQyeexbON1YdqCCWIyeVFS3ODmM2TngO9CFLwRXbY8l
sneQGf+VflZlO50jxfD56jABZfkXSkjgtxBdzYZi2twNjy9cqnla0uET8XLn
0G3McfPEXqQ5KZrA7QIaw11Kkiv7Qt4FKeliSTNRIs1K/QGthGf2VhqeBqFZ
goZKfNk5eI/+Ij2i1I/RNIe2pp7GreQhefmHbSGKSU8ErMHOMH+b99DaAhhn
IOsPwXVMvqkTJL1iAvzhXFK629JkCAIwAitJsWWyja4OJkeVPAESRZ4FXBmk
6gDNG1kU70Knyx+vRxLpJj/zxTENIiLPktqb2CDJuyIRhJjM7rfEeW+mTncF
K/Qsabf0hEuN/CFb29Fbiu0hXaNNVvGg5SbF1NWqfGa78YRJmSUbkkY4GAEU
1zoj2beE7XYBJW/s5sA1wYfyzFyS5mvyr9aL09n/f6aFXghnzJs7wVwkNHFk
iGywBklCYEIwzkHqpa1jWwVn/9A75fvQSjkYSuE7cpw1XNqTggnE1zD/1hGY
1IDxZqjMAZOqvzqH8CcyGXnfJb+K4fij29WWNYW3yeRjRLz42J8ferhDoPrz
lu3XuiVdBsa5qNmCW0vZYdTXY/3BzEt4mgzeSPtCEFv3pR88MFWizNOy8Ffz
WxeVM/JAttahd6bx4hie+Atgl//d57fEnXND14FS3vAdq25fkOvc8UPVRjMS
e31wp0yZhB7ZtQDQ0ePak0bfANNrruyyvf0sDVlGMqXCs6OrC52i5seY/Pwq
kEkSO/RUm0IcL6ZjzTIq26r88m3sVEgE9UJoAmpvYc4gMD0Gb+lY8AdeLICK
UFKXKzOMG9cd2O4rL7s3mtHsmUzdqL7P0DGgH6ooucD2+mfkSDVw1cTOk6zA
aVy97KWrJAgNSVE0gjVJSpE/4I6fSgeK2hY33XMjP8vIQJNwDQ4ubVbTl2pQ
CfqI7ex/7rZuVADDxWZHCvI0pX1YPPpUOIaVYSm95TXoMt8K6uI9FkvHErdL
Q2WobmmKqPDGvP4R6qaGtdLB14EKmQ/kDay7ejzjKOynywbfNDMZT8YGu1cZ
CJvFbIt+r3zRDEWPkCE8O+ct0yPtEm+P8Ji/+t1JQ4pc5M5SqosG1TAmu/Iy
ZDBDbUTF/31tAYROnIEg1VNK1Pvlkh0gt6gjYRuRWQa49hhuT+KERjGj1LDI
13I6ch18YxZD1Zv36mVanhJihuXlqEtQyess7whpl7yOVGzXAmPXnRPlYNPX
e4F1wmjytWWRJlW7mH+g5RIG0r2iUw3Q7kWOCYKRhA5dmWE/ZBagR4GA7oKU
V+slaSmrYIY1WMdIEWI/GNKyYSLOcQmTqoVYkvanZ03cfrY+s2ZF6M2S1U3c
Uu88Atb5WxwgFLxYVzJ47Fh2dS/SA8ATogyipAcKLSdzFbwjsJr0TwYlcFUp
/cms1HAa9RtxEfiTZAIBPK0XGTn5sfbObvNqcH1gxQCKI7rsz67cxvfSmujp
ipcWAzZg6zdFWV4qPE5Q8xXDTf9nsu32Fa1kv4t/0g5UJwUqS++WY02s4Ma/
PQ/PykMJnu4yi3ZSyZmRnu+70TOpP+U50dqOxipedTM0EdY5QGW8j776riGt
iV8jv1aXq6tmVDHVo/rpvGcE5JpH0i42vZpK5kOQbijstY+msxZ9ENEYj3/n
Z6IHRvkPyLTUno1U7WFvDeB4wRhn/8JNQhaCEvEa7Tj1GXBG0HYy/QxmXmd5
OpF7S+j+Bdt5Wlu4WaIocDPX98INwul1pPaiEEcgsiCME7OFi6/AY/vH4BH3
7VAj2hMWRCdRL8odjr9dzvevGwFOgGOucC+pFmc4RUN4Jjsl9eF28NJj7Tyx
XZq4Vva8vHxHN1UfyIcvBUKALwfj6BNo5o9IqE7ZB/QEK0APvaFnZRrWfZoI
3f30FcE+BcRR5p26Ux+OPIIs8hGwjS0/jBnHG0wesSuY3s8QaOsrHNxtF1DW
7yG4oNFHWFHRJtw/688IUcH4kYPlfdMjsHKHxgMxv9sF8RjmrxINW0AspdEu
6gLHuVv1bLRIEeFicvS9IyHc6o/yeZg7mtKULiT/Rf57k7Fon1YHN9QVRAlV
g2sA/rPIkmXq5iZ7zcKok0hNb4Mrt0gwfRmUv2btJ4hf1B9CzuVZ1Ee/ReFi
9MKe5afPxWJjO48qeXGYmFzWq8hNchiKmWqOYHR9ALaLeG180kdCyvaLIiaM
NaacbpCweD00RoIjB9pbOBef5/1CAa5aqMkc91+sTPCn2H1RlQ3uRZgzks0G
jicxBUp/cOng4fvfBD4ihffTutG0KuJODnrK2lCOriN+a/2Vm/My8ppyo6x5
DQviDoy8sf+owku4TdG2QxnvKdqZfwBcp8mfr2bXbkFiHgdQ0MsMZJpK0iBJ
SMYklRL4G4TUxp8VmLexibbcQCghHDQ74V9BiRzZFX5NHw1SbwusUIsQJYfE
9Z3R3Wk6286xndFOnOAvbDX/vaXEQ0wbKo/ThDI9AtnXBw+/+ZdijkNfV0DJ
V8LWbA430u2CQ9PqHGvx+lqJE6QQw/aha2DgfYDVk2dBINF98vJPG2myxDbk
rGBC5dEJ1AVyh+ZK6MNo2xS6R9t+F5rlmlRI+PugfjL7W7ZXvrjwvL85TVXu
KxC+iE4fC7JxaHSOY3W/DegnYoLxc1I9kReNyNWayhSwjhZjBItKsOE6sy3j
hMQHA4Q5FfLrXLr/lH6m9oHtMsrNgEBAdmSNCY4/tiiFIIB95rSGJmYoe7Rj
EtMIAW/Jae1IIG9qIp4r6wokEyiaM+DyHQWj8gprot+2Wd+C3wBVWNYdIT4p
Dd3Jlkoqspe0UThl2LUGf6dXhSE+Xp+GmHaUKcTkT3VW0QpdCjK2aX8U+c9x
JhucWpjdSj7E9nXRPXtRLBw4yjLOQwdkBjX8teClL3E9fbFI0yk2YpDwPZVd
Js4WqwYFAwl9vbIj91ONQEGh8NZ+8XrodqbNwu4T6h8oBiuyhP4phP2a4IZP
uKYwesaoU9doke9ailG3qPiYwtUTtUJxm5rhNTX6+CQiprPNhDhD08J1r/v7
1fNMQrdriNmFn23U7BoFuDqDfF7SFqE/QtiQcW9Qwo1VvPir42yFOe+X1H5B
cX/Hrz2tcLn7/OzQmBDmcgHf2tF2bKYVclY1lXc2kF4nskxp4mcdm7dbNwL2
KsfwDwDvOc3SoajwS0OM4NBtzmkqB7dAHVooXxkIQtguzDm11zxByzGOJQ4s
FQPzoaXZeiJUMFvx/xNdomkP98mpodm5d7opxsZs7pXg+sqoDklpemHhtMV3
YGjHBVmBSP3hez9b1W4OE5g0VSHP5OF0hAB74bKPYvQuBbivNthCP9owixOj
b841MCI/EteU39Gk/yrlqNbTpm1GyJSJg/dJSpZXrBOqPnYLHAdnhjTFatJv
nd8XTr3tm+zu2x5mVGbScCjPiIVeCV5/AG8ijw3cmc+OHPz30tLVhtL8q9M+
1MFgQkPofmxQ43s7ryF9mf8b35UAMuQxsqmVFby9b0R+eKSgwtnOFNZFdRXv
AiojZDjb24Eq/lE1f50kg3P/x2TXGwyQvHpA18wszlGYVUsgj5aaKvv3kiXi
7J99JvIw5oSTTCgXw7sp5mT09xbhGD3UM4i7M3N1o15QL8w6r1UAjtQg2xo+
yJfT1YL7JMN+R8VJbbXl3Id26M6xue8X74nu4/j2My9iHpGMJBRbpBaapAUS
4R4+Ch2Vr4IkqmuoWL5UiVM3LrdpYvBnkqI93/E8Erv2jw8bBMed/4aoqNOY
zCNV2JNF/1cOYWbHT11DiGAZAHPNpLqhk1O58r6ZkIDOTmNCtOVCf+LDruxg
5alzXKtUT0fFyvt9qBFcwGA7Z3NPvfhMaOBIIlZcFtkBHSp2L73xWMX1+/TM
vo9dhwjaubCwYdFsfgRrZhhyMjG8yi/HdlTm72WYSTA/Sn3ypEbBk8RfPcAp
6xTqp/1qRzmZDFHFqD7SJayepYoCKSFuOwmkAF/CpioCOdL3zsQ+mVpKOfCD
Ht5Dup7LjlTlLNcbjfTVWpq5RPoY9DJhxmM6kqqupekhpRwGnX6rkW70q9ro
fJrxCbWDIIoyENTLkpVfSuCg227wt6EMTDfnASAuRwI9DE5iDw5u+/GnsqTT
ogR4gozrtCC4L5g6PwSGmNWlLSA7JoZOgGv3ef/dLA66AhzAqaqOclqHQ0p/
MHr2FG3Ku5E2ZxLQ6CJ+otA7P4KHtd4IFY3F8E1vds9SzNO3cdtnDCOWwTe0
ZXsf6T6azfQ004If3NoUlzZZG36SWHYcc2csVoEkHx8EE7MpGFNCCYPHDha5
BhGjyBMg9Dut+RpYme/oxENF0VLU/tHuI1N0IEqpAmS/7TI6LWELoMuPLyKp
1/UoZp+T/Q3QPQzGjcQKmXS8M/eXiL9/Fz5W7NWVBCt+Zi/tyEObj+iDnu1i
4GHzdPKJLIuacWZg4BOxv8W6sxtuG+mnWjRFQKjtit1ALBT5TAjSSlW7+CjY
1SmTP0GZlzHUmDwnPhEfRLgvB7uy0G1tJUl5uAM6ySIaSC+pq7rvjH/bAbfF
RVHkys6sSLv6bkF/FC7PC0sVPk8gU5fra1uVx1pEo3GHqnlmHXwf0SXrK7rW
aGRBQG7KsZbHIKhZ5XuaBR7rfW4/i+TywJEbDcPogV5p5S2T/F2oXE7RBUx9
aayKK6nef3OQ6g9tuLGcyJA6EFtemkIQ21MvXijcwdlCCD8uvzhakV6//KXF
DrUAhRfT7wyW4VG7RFYfsxD6wFSDQ8HLpiEAoSa0E4oZMKtTLJJ0ZeYRzQdd
Nj1dJBi0jAidlayxFsTDz5TPoETYQ1Adshr+SFMUzPIBh1aa1ni+FYxs99aE
XOjHvbHDHPQyIPVizcj9aKOivOUo0cPbmRdSDG2N+WrvJ5VF7B3DKVn4hr++
L5jyq9Mi7gx0Ox+RfI43ndMzqikwXAG8yeFTFum+vKOOC/qO+g51n7Cp5AwZ
PGZmgBEJWtwkeJr+BL1vG1DkQTUf+q3p28XunQ1llzQBD7tVn3Fo3ks6QuI2
JuowhKF/LPy0ur2vwPOhx9M+lODbCSGsZPnKYxveTCgpDZ9sCMqxpi9leQbk
LXVoGp/fnqhSLGJ7NNhxPgzrBaf1FQtIZVAolD63TrQYDBwryb4BDkkXaGLF
rbGy+km3a+QVmC/aCwA2FotA9h2j8YivAt/kgiolVNOtRp8Bhso5Vkjmy9dD
ITtEVUyoh3jWVzNVSk0jhtvx4TmqJAEavBaeo4w3ukFZac6uwsTU6aKdaJCN
CKy1LOIyg5iZA8OaFGISWXsuhtL3A3oNrjk1hzP/cE6NJ7ZXsZhuWupfYCD3
IBEMRXit+9HOan2YfQ/W7XHpuAnwbJLhNUqBuwRT91zd74tNPU+E/42Ko0gZ
k8JscVRX/WZxvg8th0vcVnfXdWves2RIyWFjCQGII6CFPt738mNUknKlEsBf
Km9K3zX4oZQhiXFaOLINEuZBy0Wg95moaKuoZwxZf3G4L1W7JuQ+j8Pcbcbk
b72kd5hwqOg0TzmAZSbzFKcLx9yee4cPck1OZQz7lrVSn//vakDSVJNeI98O
QmVBXi2k9u0B91BFUmGrBYkrkyLmP70srwetHHYudJclt4YlEoS+PyzhoC/g
+J2AONU8g0B/YNMbwZB24dgeCToiAcY/sEIhl5ygsN6WjkBufYaFpYX3bXNn
UEd82bzOC/H3R69zgyMU0OG8z3qAg5hquYzk5XvKMpHpbKKlwF7SW285YtUL
g20YpYbGCceIR5SHK6fA/CGaa6WjntppopJZPtG7wenvhIrHgs5CAZgBKHJd
QhP1MwQfSNsjV6+AG1KqgT7GtKvJAOiP8vj4aMg3YgQOu71bV78Smw6528qX
eyPWI0fr7CmcodowbToL2ahpVWu/aap2lWi6h+Z2dhisahSPCm1a0y90As6N
QYOymdqm1VWvZ2JyxI+kHBIrkl5/jJBh4PdipvPUv473FQZS8rEsqzv3cJJ1
di8qP99TzlwcBWcmjlOYqPSd698hxe6jyIYojAlXc85aJxx3cF8eq265Py3c
vhURQ7rnDsAfy5nWGAGn6z6ovimKwZdDXvOuqJeapVhDqdO7j8k7AuV4Lh4R
+4c0RB9osxosi82AkYc18gDD8TUg4BHDSnkNZ7PZPg+nCDk09dubFdnlYgrm
cIXI2ONeqhprvTtqibadkH4gYfNhqF1d6goJfd1LSWRyc/2pOY+fS1kK6x1b
yuvxxhLfBrOR0Hxn4G/mjd07U888gpc8oLCdbLUjT8II3Qw11vY7qc9UCXC1
R+4NxMeq99uj1Nz1KMYODNECaMSXzBG8rlfaPY1CQBxSlyKnpCTTuAEJfBF6
WwChxsJs1Ej94/Fj/lRpR+7sDvn/IjoquNeR2qKSAXDMQ+4lNcNCwljfOq2j
mm0YtWFSo41mYlgmiQEPqa1R1KnrO+5XIjSqlL4aN6nNqMflOnXO2m+Jarl2
fkgtD7unEurdqpVU2cGt3htvzY0PhC9iMVUlXAgeMn66v7REaXZs2jlFcwFq
e87pwtc02LHwB64tdeJG6lQZle0idh1Pg9kILsqntK4aQSfKLNl14GUBciiQ
uCMrIgmhKJfTLoIqrx1Rrqnmqybn6ZWWxzcAO3vUjjcie1nNdtxoLy4DXr+b
5ZgRTOH7RtI3x36GO4Ogr0OfSNKzINDcTblWoRLtdXI7vqFCNvAGeHp+uU5N
/vYwdqUhSx+0mX3NtOHp45G2ILOPoIZQ0E811RJZY8EtCsxeSSzo9kcyzo48
rxA3LVx4PDCSY2yQsVvhmxyS54HQFPH7cPPlq30khsmdP/VWN4byeuIkakac
KFQAzpvelOKKs04XlOnmZsYuD0FgyAPdcTgQv4mkSR8hkYSw2lDgzbTyJGef
YvY0ChRSHcQvT1QGOOzT2fxosAne4vO4gk793fVHexthhBv7V1oWddtuzcpL
3n80ZWFJ+QLfSHcFYzUhjWqS6EmyY5L2bGO8JX61n2hGlJOnrWB0SLBFoo/F
MCiUVs2NuRx4ozGRmzjTY+/zD72nKNz+pg7utvRKxh39DEiV/+T2nSvn7tSy
POrew/5SWIVAQMTsbmhR6FiGGy2hWvGH7jGm7AvDzKpvo+/8Xi9KmU04MXg4
2EIePDtNfdgZO7it80CnhFSf69igCvkz3v0pd76x0levOhq581QdOdHz0AZZ
PiYySXIhjWP0Lpa3zqnsh+4Fw7XRggxw2464llNHVvCLQtX3Q+BYgpwZG6vj
Ct5ple5EUTB/wsU1Ljr/c5r1HqHt5+sKlnf45o7k52MJ6Kin+wPnAF04qM5L
wnORj31GLcPGHndnwOE1zsHL8B+ElqYLdZuAzJAwPi6xrYnOsZLjygDzxuvB
4FIy0UOXlyx/6/CJeSlYj0zsVyaI4i6YOc3zHSMllcoq99vsH01aDv/LBlLt
+oFL91/9LciPOXoNC67iX5ZORJOiegs8ix92J0l76wHvYuuC5O+FX6EOYkkN
bj3yiXQy674xQbTfiE9G+iIWksM9qH4Yf0CCopDTU9kv+Giy7nDkMLK5Durg
FcMWkX5zRfNCPJ3B9TIX4Ryai4V29fSPR21xYVbSCqszKSVprrKx8fPd1rMC
ukGvpubpJAu3WrTEiIdtOAOtOKrBU8ejPqAfVZwoQbCILJ6QWdseYqLA6y1M
+LWnAnzAQPjr+HDi80tO2Invvr6V2Cw4jjSbcuHACbIDt5xc1gZE1to5H3b+
U0j8wWzIQKztAYMp8SJsqCcBpNJoC7lbSVpdt2F/mlnMf5XvEqSAT1EnAZvg
QJwwlzWD0KKdi76IfzBQIz4b1FLeCnVV6/XIrtzsvLY7SCIULn6MN/+vtCef
MndOwR851j+bZkBnpjKFF+V/ILT0rKeoTImsKtPWtE2XMwp0C0yOLqXFOV2R
4edcpkyiOx1RMIlOWNAEgBTGPzHZqcjuVUPkJ7ZsdxT3zP0vvRJXmt1gB/Lj
nLV8Q3cPBujZHGVixZPqd6UGS8ujUx9jtHkDWx3xuYikdWcVaRgwMMQ59flN
kFqaRuxtWcRmGmtDtr9EPGorQXAO1IvntthQmdTLa6UfVfaX2g7PKi69BjZ5
QPkemPNfe5aMVjGBxFIBN527lQCBkq2jVdR70L/Gd1zt2WYk0Rk/khQ+3Q3k
KEu9JHqY95lOmZNATNlzoABOmuDFaH6YrodGNc/n/PipkHGisorXz2gsbuK7
VOY4942OlFy7IaMyIxhBvAJRwhit6nIDM2uhv4zdd1xM0y7XYXKr03rHjHZx
xqgbqNB4J4s/4oooQRcNB3wejYIL7RZ+TytzSCuDMckahX0f8op0ixVQ0w2k
szs1JXqbKsu2cTpePBwP2xGK4AhsqUah6tWBP5VbFG4fd/FwK+3vGxW5/F5X
pWzWpH4+o3964BZCoHUQgjC35p8n3Hb8vfhu/B222eX1T9Rbf5idUsA5YKgC
jV7BQ+l4nMsp/yZubls2EjVHT5RDXrG8G+MEd2wdq/cx8986wtomab/7Ml9f
TrVYyxwEQQ3OsxCurJbCHxYoELpMvigrYvOPX2A8yFvpJil0E0i0t+Z8eZK5
V+Q+/Abd3REGa5EztUq91W7jgesRenf+zYsETLvPgvDdnODRtjvY/5k7fWRg
vIRTruhVeWu7/ZSAdo4Ri3+qhMY5pO0ihGvj+FNk8l6ORqwvTQHhvJMeGnbM
jz5cJxbYqgft/zGl2WYrmjveuBAM3rXCuEWp11RbC2Emcc1f5ue3gaB8wHis
0rgv09YKU4Oj+38a67zqFuc0avNu2IkEFR6ML9haXzd0XvrOcLvEvR2MsaUr
2NzrRvfIwkaoyEeNLc6TRDIUATZfRoNjC9bSSMhFdKHpp+d5hgJNPWqOaCeH
IljABggDngU2n7xNk80LnY2gqH35febwA1kE8riEFLkFNt6d2m3ZtaYs9bgb
b78yCCqfTs1p73fj5h7JKTNDyN7Z4AKMMtx0wYnYBSlY1/8mEoczc6hdfIt1
gflYdBzWutAGxvfoLRkWoy/m/ltPHVXOTxvllBZ5H5xkPsNstJ7l+5H1sKy9
jKD8wVCurj8rsDUrtNW6Njkb2vSKyeKcpgsUbJ+QnofhbcdnlXr07bTYmbJa
rDhVU43Y72SEnq+gxIU4hcRw6B9K8WqwB1ZJwOrcXWdOa4Tx0IhnHnWmn+ub
T2eCKTUgJ280H00oeyDIMv+CKICtVCAZydzCYcY0+3v3mF445qvCP+O9VlFk
FD0H5FUqtOZXEM4L/YqlcrbfenXPCsnB+OvjHMZXDa+AFKDkVWhU2uuStsvi
mpt4+qnZJaUQ65P6i17FR1pIqGxEWB0HbKpzthXb1LNJ5kg/cgJtfz8Sdws5
07QWHfL+OMdoT0VENS2xdZgqPhSZ51UbNvh92XNSGhjUydVXTb/Ho3L6a+gl
81kfac3tMXt3WqKf+XJ115O8reUSZg2DmtG+SqKZkE64lf9QIsmQbcpLOGM3
vHs/nqBwsVweESTPeL1WNyWPWXiNWPaAwazTOjs6VipQy9+/GJ1Y6kEFMtP0
oQ8iLNTNgERo3ifVdurmCmWwOCsbEKW2lePMS+9MNNC7nD4MLQi6FGXtdWuj
kqLXtM45My6xeKP/CddNfCs08FgBSgWAunO+r67ycGxbt8+vkHsBe/h43CtJ
H/83PNYqo8dfrI9cRK3gJaEErgS6+auKoSyYm1tE5lGsDxzyXKGoAm/awlL3
Oo+1hDAWVbTU0UkrgBuZQEEi0x855nnJ5eJPNhSdHlYdnu1lLZb1UpJ8ppqu
bhYi3ABfaLMFTE2FsSlSRg1kFTR32334ivvvkUUfxNm6aUP9nrVCvdYNukfr
9s7XbSjHiDVp9glCrqKxsOjqAWd+U8xaRlYT3KAACWD6kOU3FVOut/3Mcj3x
V7DMm86Rvgdcn7f0H/43DRNTbd3sMtMarZVkebK6Sqwk+tnhlRjk9KsgDOT1
UqS/s8l/wFbPSVHY4YbAcchiFWxlHtHy4NWA3wE6P2r6QsEYcaY9qqQKJsOf
eY0NcpBwOKaGImLRoHT1RwzWgfT1kB0JwRZc8/WtMJzFqiM/MtkBWNrBwC31
0z4A6335hZWqpaA/hHoePNh2gzubEhzULwJTAn5Vle8Ygjamm4KLTlEd68Ea
ZdfhHfMBVfb2wKg/82RGPGO2ab2brnw5QXvvIGypHYNFlQaNOBL/sXSxBlb8
cbsJCg4JADjxgH09w4r33n0pvo8doELNaKF2x8D6X7oL7+GKWmNbkoHtmvkD
XfCd0bSHCefzbKpyG9O4h4xA5aErLpRBMUJVke8wwk8QEe8sEmGdiU2BqNch
w/uH7Sex2R7wlA8SRgmAzQo7mMo3FIzZeudMqvGIqMlSkK984zNGz9y7Q1Xw
4PO0RBmzFnKX0uYyVfQc+mrlznB3V2WrM0xSTpUw9CqgqeHMC48kiMBCt3Fl
YzhJR+eLQVx09L8du7BMP+RBMeej4hRFCPgXIp+DtNDV81YyLxytdEkXwW06
rIoRoVsaNl1eCtB5TXshSekGldweOhUelQvSMrOtGXo9axIpCSOu0ydgPExJ
HnA3d62WYBEvpUmqH/ZjZ9NfzLv+hUQWlz4+IhCZTN5G59aaPXZk12LB05rW
a+GkiFogA7ztyN4WYOpRnJtNrymcp+jZADm3NmAGDGnEONhDfEox77fBbt+w
kp9uzz2Q7G+FUtY1QaL8umf+HFpxQTKYKcUl6oKqS3wSw+j3+SXNbb9kEroW
u1YdhU4TL+QcGC17tNC11sbAMntwycTzj862bJdcw2WGyaSkzZ/OXyNs85/Q
RUsXrwYTucmxjd/eVYOvrc4utc9Gx0LtWQ6aOL6BJyWxFVNAAe++V5uScdlJ
+Mhf3Uxq1KI4bkSEYEpyafN1xRn/TAVN6/zE3QhAdS8TiGPtm7ZfA6mDI8ju
L+3zEtMOhUeycDJ8JQg0n7AO9rI3vNi0PuBljyodcKg7h+0r/RDQYpKIZ7sg
2oklDqMrLwvgy5XHnwPaI6X/yIGs1NdkDLG6Oq6UrOQ+faa7ktB1C/lY2pjq
qV/Vh8RxvbmGxhC0DMtiyQmFeEXYWU0O8KwYF6nEaadRvEopz/m65O93vh6x
T9DZHly1HiUciQn2LV/izVxrf7kS9Hf6GQIE/8SAY/CArlFuZwvBy7DdWZFl
O5DpIaxRGmsBr1K2zHRu9l2Mp7ut+juCTg4ny2ws1C81LsbEpKAvRSmOa3UE
hIHPYIlXjLRpkzADbSaANWp6VDMDR+CTZBE8xxJMSNHVzI1+C/05h+itweE2
xk82GHD5rkbTkGPCPLv3Do3uCKERGyx3bfgLt5LVrI+ohLgWLtC7lZwSqe6g
otOi/7tBMOqjMtAIbJiA+kBYGNtnIYzT7mdDaoZUh3XEYWTmHnyaugyQpMRV
yRb2bc4h/VkzI8QSu6PEd+klA0OLcBP7gfr6L8XBp5l+wVFVFBukVnz27eF8
6ttYrbB68l6EEc28umEjIakObtsflUOyF9grJCGICoNQKxYqL9z/MkGwa6nu
SJN5jpCICKV7C4HcL8/mXpzejWvrF2aCoF/j8AoqlJzdQFLtqlkDLxPDYcgE
saxMHEvKHNsaDdogmNlvJXq8xL1vabnDC1ddWkuW+yEU+QvF91uCiXt5BkyO
aYwTC4+Fh5yAbT8x79qaZTAzd7S6B0AiWR/XYqFHBcvQa58o5JrHvaRDbJ0O
11l6rdytMZD/iz/7rz/oWDNcCUeZCu8RmSPhkZql9o5Gu2Va1veu+b/KioiJ
2hkywy5ajEiv6uW6EJKU9bwHQwlWCBg2mi9n16SUT4TgmO883aqGApehfyY7
sxi27ET8PvEDSKjsK0cxvgxiNVQODdb5IYeG9FgkWLy/8NGAQQUwh+VYvsrS
GZPF5Nbu0VwdZq3rWx9eEAMO8XZYC7QbTZZxJ63qN3k2lop798iungYNQ5P6
P9e/ZcbS9TCUwz9lrknS+y85+57ntrquXCWaKO+mKXZf8fviMHhyd1RsQFo0
6BSOodqmv4yQ2dTIYTNQGWHxAKDHbUox8kUfxbO1Si5JM0F1ZDiEvdh0jyrN
seGkPrqENt9+BV7VTSWZOILtzBsSyNJokW0lpBqdTFQ1AM1brsv9i05FJiNH
U4I18n4ES1tNeFP/Ol1HjQQ/qjN3WkEChj9E+FuhSBGk8vY39bty/P3yO1Di
ZocO+JOIWswCmovQmVxnftSUrTQEaUBwr25DnEgjLhqV7gNneaOeRajEGwhe
e3+mAO6pK0DtubtqUqARWkktQtkaG4ELjVG04bbMsDbIgA59pBnoK/80DIJU
mfvpD7/9zvHStZ3WIKYRu9iqYI0IANOkYtigbq1O3PqDSCnoxTBMMqbpQ1yT
r+WjSYmYC38X0bLWic0YCvnhSUkkPDxcTLjTi/ZEdY7wk8JbSPl2M4dQIW7P
KTvWbw+Q7uCfj5XUW4M7hxeBbaxgxO9u1Fo75OoSVcrAjAxYvQ+tq5q8eX4s
Qb569+356ETBigYjii0q5uY0NoiYYuwQiP1V8tprQ+uL8z1VHdrRDiWuOare
XA+qPH2dxo4RsZ8s9cFTwlSat3pKe7lu3FgNl2D8/NUZcWBLldbI1k+gLi9F
k96ZbHjyyR76vzCWcdX1dgetPbYhdjtMuDNtsyiBmoUb7oVP9+k2EMVkn8qv
6e5sFoTx9BWFyEeYsWptI369TyZFvviYyIjp58/NZRqB3gzLnSKnzO7qNS61
MwgSx7LvlQvZEyAvXmWbMrYSXavQPH1K/ObXvzFcSXOVWZMb9UdJQMIRXGHS
Gbee33U2yWq7ry1QE2bioRM7fgpzq0lMXND9TMyb3y6mX0gE6mU0TRaf1ikI
rttyX+cdPXgmlD4+U/UkBi7zF4jvtbI3PUuA+nd0VraxNOYlH9e1KIJ+6hJG
N8xqcVJS4MQOwOmjX4mDfn6b01iSV+AbM6GFlKOiUfgMzn6OyezJfnBKGTrL
hgs62ShrGr4oJ34cmZtHN2YqwGw3tzsQRxFT0iCicK1fUoWgojoQXJJw21U0
snY+6Uf0mlTGrQ9P4Sh/dJEcsgLJ2bO+uZqbG3KfxcSpCnjoAGcmuIf8ywcg
AUBqp57V/TSOf+y38e3zqn4FVEh9brKUHK947VuWdxpuYDBcgcNE3EMbEAaI
vmdhsJeuwIkRFvap46zh/mSp+T3M1a3Rzzz8XnSvSj2y6x25RjJiVljCp3J/
+KV939SZpPFdZGgN7RDDq7iADPYU6dUvZp6v0ynUjhT9mV6HV8nYMwpW5I69
cMsSrx0tLGe/kIoBuhMxoEkfPCBbVbTCXOrMzuRks40y20LJa1n7N4r2n806
wnh/JjBtZHM/zXkaneEITk3h9S/+qlol0AZQ3G7JorFEyCz8B09u05HNXs1G
SBMfoekN4pM1J6FVBIA6W7BWyFv2y92wzns+Zyws1evKT/sQw0dg3btnt8W+
NIdKxEjWqlj5Rmd5RM1AbdUHC70fnOumx0SM+s338EnH1M3mMUA8gN3wTCQN
Ni+14wUBGlLbUHVrySXX5OvldQ/xQtRZiYZvmMtza2knc3PHD1wPt6UCmsRy
ZFwPjT1/CQ/fn6mQ/sk+gt99n/6MgDPpxw0GJZ26hXk3Ji7/Y+asYyAQNDgE
CvfDi1yO7vB54OY72Lws2LKw/OBsF6LEX1FsE5mng5V5O0l7REk0hIF7+FlO
ZjOMBx3H/szARKH1tirITYZq/KjfyB+lY2W42SO86FKy01hPDsjA5fzihtuI
sGXYH+pb/CrRmdu2qFG1Ik9aKPqPdDj+tUHexRSMwisfxe5Rax2k8uTPgzb3
S/fDRkVBfCqSr2DsO4vU/VQc3EPKKX3yBTW0kACljucLCs6nfdZgj7cEgqcL
BKkLOpoNjxnSUlJzYsbQooyvJxClhuspd00LQQssk0Qt9agRWhPpzFIC4j/o
yugeg1V7lQGnIwY+pdAVe6t0hEj2m7146o5UdrhmRQqemaQ/EeDxUDHpQcJd
LEJT6NSWzCDPpeTuMPg6Yhqz1A/0nTHdMf7nPoay+4mk53U7KYGP6Z+R+Sj+
OfO3Q75p9GPlmvlhZTv4OOJYoDPoMQZlrDln1Tf+VZrXf3a7h68RSjl8ar2S
xESAmBG2idLQsL7L4OljLcRDQfLKvzKGQn6TdJllwe5xUgDDcvVwUwpRcCYd
9jE6FQYx1LRG0ah8blJZvmM4TtZIyjeuItUx2SrYkEvbfZ0b3lBdoR8JLHEF
MrytL2dsPp+Xag6M6WV3wNVmi08YqNH3wTwLm3sipTb3QwdMPyRSHtEXKv7e
vqnIgb3kTGVxzJvZV7722KZA2MrKQXQX+jtIURiI2aNaYnK+YDxZXagDpipX
XBs7jaA/GqG0z+SALqF3rENb6PVG2snSRAEmr4TLZFXUnfZXJhCNNvhjpT/B
7PXLey/CNlh2n8iX3KKkraRlP1n43jxC3pfQCU+Jvy4FKa2o2oE8e6n+llzh
gXqsUi+Eon1rZ3NST88iwWvdNAttJZ55lHQIJn8Mt9lYkodmylm8HsRKO3KU
fI56HVi9imV51N+tdscl6HEkRHSR227h2W4o2yE7kHr+Ny3DyyMhXvtR1t2C
M1DrcDzEYBGmQ66ZbLu2b4y1h6Qm2oI4jIornbCSlxR2E6tK67z3CvVZi7CK
+l21b7BTYUXo3+IH99lGyH4Qwzu/QLlnZDQcQMvyXfGSldezXdhp+qF9DtvE
71j2uYPFRqFauWzsxEeiFN/i1KUVHkpvZw20rnujg1Fl6dXV7zHVEjAtEL0D
TOGRtWlLbAPvZDXLednUXQbmyLv+VwpTtPUdvTz3N9hGNWnEaB/RRZk1WR9S
eADDpQVSSuKBEzotNFV+pGNjNyycm2hFYzVwFe7gh+1iYRj3QXFPX+dElVeD
dQIiqUqcq3My7jN8yqeNM+r9U/eRrgrslMOu4ZyoJNjTLbCe7jJ/6pGjoVlq
QHt2PaQOpcNfd0Jnp9EvW4GIXmo9DyltYdutyhQFzgPlwYVRYSTCI+Yvu32z
MXZEmaxJesMW6B8uhMYIOvgHlwndiZwjTznHNXXoY0Of/qpX/+hlhHBJOqqA
YYQwA5JSlQhxfiBESxQKJdMc6Fjef4nxZAlVEzxwURw7gYnO/MW3p0ibh27p
SzpsycQ0mqfOFnZyDTD3gUs1I+URabm307M9oQPq8Law+XECcOXVrcF6VMe/
Xb6aZqHeM7Pbgjoq5159XlY6jZ4XQXlRXYF6+MNOjoqvkL83ZVQQMH0gxo7T
xd2aRVdJQ3wbycdfd19pr3o4sd1Hfuatu+uCLhXOvWkM49XpgM/b9ScH8H/R
RsYAPGJRaW+s7tuA04ZNFOYgoyVYySecPQ4oyZ+XqwKugl2seUDNPZ6qz1w1
QRwT+q80/cgqaVyCJlvFAa+csXELqCjFXkyKhVf7iVwM27N2ZsavQ+Tl6owj
Ax8t/hYUtgcVXmLHn2MJU3srjkFEEd8qQwKrJlKN6ySQvju3dzJQQO0YZq2a
R8s38beB/V3DueSU8fJsT6qcyQpNA6Y1PKAsU7rUGraOUSxlq4TWVIv8Sf+D
ifuYX3K2QBcagDDcqWum6kLhuszX65vjgNYZyEpT/cPnpRh9Go8jnzrxy+9p
4bK/EapBEKdTwwJfSrv1g1g4jJ2Kac75yev9lUaJqZF55mUO2eGUxBe/rq+R
ccghJPzi2sNtAkmkKDUL0PLn2zBJwEE9+kv+lI0iwa8bSBJKi95Ab32P1Fo8
RlgMCheDm9Q92l6YiPnJUmJ4RbWmezG7RJCPJttOxEGktQZ4cIVs1tlJYcXp
e1is544EmW/WN1tc8NCYB/8gc6AIQArrYwBinOtwgNxEPkzWvek8A8QRS60v
ExMchSpTJXOfKPsZeWg8LdhUT81QCm4o11kKw03dqx0QSv9SsVU8+FyIrIyW
HbuikQLGEDIqtpYN+SEw7ioKNaYFLEzZNFl1kuHJob4Wn//38xegpU6NYEfH
ZbhswTE6VlVPzKhOkOw/IzFWJ4f3hgkGpOk/R9ie3GHmvlSDgJWe7BZ1KN7E
45kOoDSIyZ/PZjSzBqVPrX54R5mOunJUfQMRXeZ5aCSCx5epE/TKWLUdqjpa
qs3PzVa7mYF/jwbxtqqnnqf9LBIcX7AvHZjTDIgzb/ZQzk/oHjQFOuoUEUgV
OVy6DW0yvQim6gQR9wp+xR1omq+TbjwaIKtpn9b/iz9ENTQ8u+MJWGTzEy/j
vIVxrj7A4RGe7o8teSI0XeMBduhBCdHwGTS4h7yBCo24cdsK1pydhji+oeKT
xZGx+8Cw/O5igYceqEvXoCpRT/ckGeN//epSxumHaz7aKHn/WdPjRAY6GX8i
tz+w58l/Mf3I5OBCJsBQYdxiQxbjB2uuOYkTe5dFnkOGnArblNJZNGR3CWxm
s8hU8gc/mbx0USWFArUD4lvlItus7g14qbnOc19+1jNXacr5NOcD4457zt9w
pAgIE/jJAgV1qSYJY0nnFZfxMaeh5zqryFyWs8dzTdZiuQroeJFt2EP2yrtE
98wxsUo9CE1f2Rlk9cG/Bz9UXwOBkA30mG2hf+IcccHFeT9CU1009VWIOwMb
kNi2ZIAyVdXcz6vzCPPNQmSaMt0OOFt8QC1vuj125+MStaHLJW0vBjeWVeYe
pVpnv6t8BHFvM99BMIVyhUHs9N5SzaW7em0GRZFarZOaLfiMmWqvlNRj1k44
hCdLM26gBnbrp9NdiJdtyvq+rWjnLwdk3a79lJxMUEHDUzLou+Wj44u40EcF
+JsIJzWc34uN28kS+LZ3eBSvWHPnC/8EDwfhcg9z/1sZ+1qPwLHGtVM/5Hgd
nnEGSak/Uk18G80NGJn0m8l82fIHc+fmeXNjSlOSg9TTYPNMJV3nh9DiNKpq
mxALbQwDhDQiaFHzfNlanVIt5PPHdqR9hPPeRs4bqyGmCARzSvCfV3BTbAUJ
LY3nOcVrNuRc9D7SA/5ZRRzF8kqo6VPCJRQc9wW2CgwHwJzt08BE9eWID5lU
YpTdgvq1oTgtiFm/ugQlkgv+kG6yru/Co61xK/fUEN9jrYruTxNwmgAwQE8V
9CfE6L5alpbU4OzsJDT3tIEDW+zTl1kvWTQlRi03tUN4P+4WEA3M0XbN9hpc
dhxVTIasdTKcpo7gIVLJlA+5lVjCwCecGkMZhBjna6kwx8PGBZyOB9tcjJTi
sUSZL4zyfDTqdJtUjlcP6QoAQe8j21ORVOxQ+Fb5WMZFaoxpTKLnH0YimV+U
A5FLlBFSTsFCF69AZ1zATCzC7Hjh6jzSSlcOzBdoYVJTd7MLArr/uB4ljIEC
F+rroAYOkmzuBO33qiTRcqdd2pZNSwLqxAKW0t4yT4v2Wp8bSOshUTd0dMWz
6rGbx7CElvCQAiY7Aw9Q1fhg54W8b27omCGs9QVD9nY9HXS09D0MQhnh6ysu
aq0u9T8OIqzCfCNw1Cky2gslchs03r2V52+iUsUprZOAFY3reYaYlZ6RSjdv
Ibhz+jh+UxQxiX2eIz6tpUXsiIdYxsuE2c1hcLXEXbm7dAgGqOci1TawkaUH
Ay+f9gQZ68zH7iNPteX1vVkCzRGaa0sMRky3tHcFchgjBpbC+Jb46j/LA04H
y0ASWUB45SaR7285vr4vLLkoJzSWyQB8kuOpHyQQu3/2TXpv2efe/WfuPL1y
fN5+LNH95AVPuHgjTWSJOcAZQa7zvBtirBYytnKVzPeHqmYNP2khZd0luh+H
tlNzzJwHyw0gCtu8L369hi5MXTDnzRg5ZUn5NtcIfUNeEQ+ZFA7KGLx77MVR
Iob6L938IPjABVFIrXJ5u5YEWerengIqFprk9tx4kC/xUktUjpHEr01sNNp1
sALMl4FifR01DQ8Vbk5qR5dZik/ocQGDwh4PC2Vwf/HX3FE8OQqRGOp8FiHv
d12ADgQmHxIhQP9i8EchcY/5CKXEUeK0eKNIlpj0l2qBsTBnbquWtdK3uZe1
BBvf7J78SAJy3zlWgQO21Z0oPRTRz/h7sQlmX8naRds3SLTUiIfDlPaFTsx4
M/5fkiplJsJpAWkAPBsys947dCRtCLsRqEEZDadMaHaDtySWZjzSlZ1fu2RC
jkvvFFl1FK+nqpskWdSk/8yAsHMw/C9LNffqCtAMSJ5ABVVuStnYahcdRKqF
p/Ft8lsjdzcPX9jnbTKHL1fKRUcAA0mV6c6XO4B3gKCoYLHd9nnCmC28z0VT
GDksvPc3CX5DnFitsnewSXcm+jFw1OWtxSjGJVFjgHAjIrwzg4xnYdEe78GG
DeUHjmoKTcSSttqIwN/r0Q1Lx/OXW4S17drjkPCfGXnpoLUhj51N54YdVDt7
Uls69uM6PbOoWO+zRUBkPxj5HKGpVoz8CE/3aKGl+p96UPIltHPtKpzBvUOv
EtA5y4XK1JEvnkNmZTVqFD9uD9F0VQ9nuLDL7GvA6vTjW66iSNxlPJ2J+EsW
lH8olClxd90EjjfxpKfl/HAX4jTMn8Vgayp8YfmKHmT0JaEDWe0/ss5MS+9m
Z/2XSmf1Bjl0L7c7Jmv3BrDJHNtxVIUmr5zcS0/nM50VJ56Bq1G5w+Zmxcgx
K6kpXj/PQvatytoEkIY+4jm2D9UV1yEYyBQAIs0MkWdYNJD9pWH+I+6eS+7d
pWgr9Mmzlya8AqieWyO4Boy7xhaeJAXrWffavFRTQhHHfA5XyggVINNOIKk+
CywF2JkLtjUFuBWPUE00yQJOrr53pTj1LP8DYkNSVWXf1239w1vAQhmY3/HE
eBJ0J3DE31QS7u5ktCfATbPNgq/01N/CmBkiRi4bdmzYtEW+0yAD1WdicF3M
SB9Y2C+BsFwVdOhPmEE0ChGzCpZFGB2Gj+K97whWuqLWyALCbGEErcYTul95
UhUd7xcgNEWzl8f65jdHPwDfl/NUjp4f8qj9hYp2BT+IAZMCVJl3SayNBYAU
EROQUV1OuaUqs8kcSv+KvC0iX+cv7CkJwiPPA9jm1h9DOiuYiV0dTKVk0rK8
1JwyY1fMwH0OHIXUo9Prh+lxjYmNBhtzECvWsEi8L/maa/8ETfRavxzzIzqT
bm3NLoWsAoy7fo4xmRROOTwOeXv5Yb5AlZvgcMoBDYH8156aOeHVWnqHjpuG
NPrXLut6UPjU3RspKF+dXc1eRkkN9EzBes7MZRk1rzugHT3LvRn7m5CancUs
WwRI9bZKMHW1nF/AyJJlUamTb9QjG9q4Ak0qCCECrJvl01UfsOF4sUvayZS+
8M3gaX2wAf493nrIyFKr0ttpERzg6J8G6kbtfGMPm/ZV6EgzOyDnufyzh6xK
LOWjxBdW7dVC/om3iUVFYCaFyF93PXrA5HsobtwK0+6hhoy7YdHAhI+qfOwX
4ltBjt1Rs3Te6wRMYZrFBZ3Ucj185g70iJ6yYeYDLK5gI7tRwErx3+gW8WcS
o0mGql7rsU9XWRbJ3uq2yfItPkNiWv/fbwcdVI7IC/i6ttdDLRMjk+ajsTZO
wQp6vQ8UxmVgi/CE/xxFbCkBAsdFI7z1aHSS/fYrpeasU7izZDcMhvF78o+4
qZg+5xTgaL03AE3VddYy5n9Atcd5NVC0HjaPIV0cdhtY0vV/FjCoXa4gVzxN
O+gEMfXTauyh5QtVjNV/NyzTxIfUVoV78fDsjaldi7VUe8bWQqqlFVY0rWzM
52j5gkMTXuNNxm+6ARnvn20Z4SrseCprTr7Eg7TNsLDqBx0PxNgUdLl7KiA9
YjQyR2/9JR+L2q7fUouzw94Gq+19fK8EX41zjxLIPZmLGz6huI79uEx1JRJ+
GvSmyKJVksqBPEc4YCN6u3S4XPd/QLQGdzliFN6nAzRMFx5vY3AKAP+8Y3HS
HnuIaSJaYs2C/JZS3ju163eG8r7LWoQ66vy7i9u1VYpTcTWrAByBOqHnp5fz
ftfQ2IPvmlfsKHLMxn+i6I4HXJVjdSFvUk9qg/WNX9v79TsUo7AaPfCkoxzS
oIk0xZV4BuL4gXA91urQDdBsbS8sO8ZDm2sUKVgvOs/E0S0/siTzRkQ6JCFb
3CION17jvNTLIs5cC+jhvV1/UTfuZSXeKbvbGQUTGoPEjcqKJSM/Whw1vfaP
lWL3u53jHlMy5xxbye2np8c6xFy/LSN7hpHPVtxWYu97PNvPq3kVv/pbNqGB
F2q7sXRC1GEsfM4cSY6Hvam1/BOi8w+0AmeNILQTYi6kVEjfY3Bk066jqKUz
lFNrlN4rK2W2SQPoEGtvbR8gpvvGu9z40iltU40ky9mwRDL+M4aPsy8LlFKa
xUpmL3qz6VnaAVCqpbIGyR2MLbUcYHn6t4yiGyD0ZNjrdmc6c5gNuhPGkfj0
t2syEnLMfjzl2KTcPUFY8ehPDtFmG1b0pTmgMcLYxBO0FjYzwfX/qYu4jy7N
hxhtq8TsEwyHOr8wg/CzAiplj3OAAP6zndD3xHHm/w8jLr3Edsmgwtmgie18
JqcyiVhiSaQzoh8xs/PoeF5F2M8m0HhZSvW7aQ99aTvdMJmQZ7wDo0+pzx4n
nY6bjESWahWKoDaI7N3xbuMvUn7W+GnGfOLmPI+jJSYJVchOn77nAZ1SwNjG
efTxEJg9I5KJCku931E+OMwu/cPC/gSA2AUdnGdEK8w0w60s3NvXeYiAWuMw
+XIyYFey0llw6bHdI/ahns4qVCnkS2JsY/8Bwswf3lpZjpIeWGT5gNRPis9W
fg9HBth96YpwYCz8u2QAaLwg/P7dbuXhZM9XDDxRvNoAbIIvmZESs6dLFqZA
MEnUfuGMbaZokuiSucLB/d1vTD+OFJxR+Bl1gkamjtyNGV9j2/fcihbYUD+9
tGqu2JG3QwYFTLO3URyb1i9HUD2wUxIOaUcAn383e8CXly0nCi0q9PkHoWCT
ION7X/Gql7AqQY8ygZH2u9cLsPOrvm3W+3tfRAPfK8wnKWejq7rZiYtcDtdW
eoiaIGfa5Hn5Y9arNyLRO56s7fzGdB3FRcqkIcCUHbrKqwO9QSheZNDjAt8S
jVMGgLowHNgItQrySxOhgjvE2UGBCMxVybqgH+tw04CXPjjKi8My6t9T+0Nw
0VFJSnXoywfkq9nofKGVNzmKRp4gpBUaEl+6fG6Ejoxyt+rtHBEFlo3iruGS
K2SVC+tXt8J6WRSoR0s5R+FVWXYGczdbe+JTErOyF7dg5rP8lTa+D7ASe6z7
CWvpnlNDgtluUoJyrkiACWyUic6IM1RdjT2lI5bAHwdJt3a+cax44Zb6qEIC
F0y9odeQxUNRePvkKECN2EOe+4US/esCnA+P/LUvTk9jle0L+cD+bNjYGRq0
hY+hyvel73N740OzJSXzsmRvREps06/QhoZThJnNurtpd3qT0aeR4z7vY4jd
uuz4GYw6racanI9jg28VKvTZyqEH+UxLNnnAP4lfrXboqBEGGoCgCPp+DKSt
KgRzzYhCh+VCR7mP/qQ5uIneZNYQwIBgGoxcbXKiADbfj20UPhcnWtpZ+rTO
cP+0dkJaJovc0e1BGPwQ8tDuVl/6yfsyhAP6zlM+zB6BtpsvwnyUQ480uFaQ
v5uVFeeMTYKB5cpV/z5y6qbzHHHV2z45QxOkSE65iTgDsg84hgADPJGLUqyb
oOxPLJzIrXepyS4YcM2u2+LG3zgHLUj5Tm14V+vUxdbvf1uJ3D6dk69hX8Nn
v5WkloU/IFg2N6kR7ewynF32sn6B/tvJtU9JKo0jsrvH/DIgQePeKzOIYNPz
JfSeMztyp4xXQqVCq7KUrIi+DqBpOSO4khTMewm1xLfAe4EkaA8Y9mABPDOP
1Fk5R4vO3LfYOrz3To/3ySe1yqUSP3iEconN8M4jL4tCtpd51tehhS1QLLP/
jRCR6TcB+viEQK5nRzgWYjTFpmLj71ROs66i9BfkjXzymZPGar/Eua4pGz5M
P7eLtWXlw6tOrA/9wcC5AuS+uq0Np+sbPDtEQ5VpHicbpNy3i6o/rZnrkVAs
3jppcH9uvLoE90PClyCyX30eyBrwo6q4jOyXIP3+8KYK1IGMjXwH2hXD918m
chhWFZopr+3iZQ7JNfusynVkr6gIEtoIVdBinXDUJDK4RCaRxAbASChRbAm1
sgjd0gFJ9v8oELeMrcLRcFiN3eBKJZJCeZI+I/b77Nq59JIJqkMLZtLgUW7f
iXLQLVVbnwsiAarls6/DZvewxkmtZSBDud9S5aeEegTvMXBd1h9WgE2ikNo1
ng9utIue9XWr0UCAR8sbaK2/NUg5ysFsMohnr7g8+PTSNnwpEpe2/F8QExcD
hcNCaqM+qNx8bpbnQUCsgaVZ4Kp1t4Desh05se5E+hUbWPhtAgxTCNPA6EUI
WbV6mIqY4uJeYSSvxIlCmRpWXrnao3M2e2NSHHxqlnX33W3hZ3qZSNy37Wcy
i1FqPpkLoxftDNjVuA7n9JHDLea2uPqHqbuHF04Ca6Q9Ak7oVgjtHAoUdXeQ
YPPfkUgAVgvmBdcYhagdR5tMxg8G2jjhHyXr2WI571FGJm5ixuv8ccW1mUic
YJ3Zlv+iLr7yhtH9U5drPVeGjOTLWuvDofIU6cYT+W4T2BYqzATTL4Q5nchq
60zFUyODdS4M0yVA4c8mocJLiK/42ka7+HAJLX/9S1ox8h0BIrm85Qj89XnH
Ca3CZEdOYvA81yb9Xxmt5BB5NxODTzkDg69Zh4BpWZvx79gf7Nv/bWwGA9Hh
Nt6TXbl33/UJN7c3bPORdwgRqdlu8EBAlyYVZIe86xm/MtbYdq/J8N7h3jxy
aVqYzxcucGBaafceqoc0RaCzkYhbggoc9yl3KQwkTMNcoytvL92WnkBxGiAJ
c7JODOvu7dAoG6X3bmlghw0o4yOKmC82yMF/YF0oYuA2CJp11kvWnTwxxJKM
SLknGraQeMSE448M4tEDUxDi2jv6yWvwhdfZuEJqaXFMao4/lTrKMs078z7X
6Zzazt0VRhirdqTuRR5RVdwQYWyOy0E03xv7oHuJPyOsnMp8v/ggq+Qj6Hb+
zZ3CaT7teeindnzhqS1fjry+MGPWZ/3+zsfR6QeOm/xSIPsBD2J6LZGgi0yv
5lWpQMvmB7TqE1LckmqeTIJ7Xj7o4j8wQc+Skq8BYkmvrm6YcEdqny3q3A9R
4gr1pGgFCKDLTVdCzGVVQ+9G+HWuuHmBjJ0o6+U5pZWqE1FDqvf2QEzy4pFs
Rwrq9vasnd6GJgTV2luf0g+GBFD7JPmHnWqH/A3B6yiWtyY3EV1GRSBu1D8P
RSE7HUHlZ3ycSZSz3h85vLA1JLP09KtYOFTYz38yFpVejapwgddxqCjkTmU0
ElJ9zoyrFCYvBl3lxm9M3nEVtM4udJxNeBRvfov9cpn0Ang6zL0SVuVAd3NP
fO34zSH6wgnYpiAORh1vvcLHGm/sZ5/NbAG+Of4O+/DDycXEfW5sXFJ325bD
7wWR4P0HQ+SiFMgag2Zv82eDC1SzUvIVGIAU5e3ns199HaITb1fQIpCWDjrU
GtjfYq9ZomjEYCe9IFdReyrnAk2/QEowX+jz4J5GABcAXZz7UjGsJ4c6GHsk
iUR5Uj0+RMrbYLEa8oWChvrSi+K2zFmjb5nTZIcaDc6XLSEV5ciT3iatVh+C
qQ6vf0C4YcM0cHiID/rxHfhz0KNBB9J8ZQFZsRiQT8T7/DrT9pQAM72MB7IB
Z2N7TqTVos9pLm1RF5VjftYW2baRFdechsMYdB7bq2EtQslrEmgrmuRMepJW
xzlCSs25BxVbBcpr4mo1Z8YOAm/RDw9x1QLq9rqS3fTMBc9Egt9QqdjfYGzM
cdONlGqj3qvpoF5TN+KYiM9lm10KN/LHJD5vcdN/bugmT12IscyZSF6Cnd8n
kPiH+rDcHU1hj7PbRDjhYHkJQJIJTdHXMCgIqbqKSP9d9W+kifE1+NvH273y
1wM5kRe6Py0euvoSkEDINHaqDU04NCHyt8/yyw6omBlmcLhFmO7SmmaS1Gv+
NtxNeUj13h8EUUc1QCUDfkQ/In2YeGYlzpElyDvYfto2n0z3CCIk1WDpyKJK
kzFynjhdb7hm3V4MHfcvhsjqPTC9gMYTM478LZjJxWXufG+5XztFy+6uaO3B
Eombqtk0Oj/WOTxpr4NzVD8jVJuSpt4lP44DT+9Du5TinHNkRpYWhwM0uBHD
7iwnwxlj8/HZMVGITVNeu3IoU4z9VtGp2XVtTo3+7znK4+ugrCMA5jKGyhg8
zh94IF3DHBiGGFbCPste9X4XsTqVEx/QJMgJ9C/PDCJJlY2DFc1infeahOSL
FF7l27TYCnb07lXtwhFkJCaxwzV3k0AgDeVx9lXxl+jt/1e828q3z6TmyIp2
Izz8RSREHEDPrysy6AkemuHBTB4LAUy8SZFprh5Hoo8x/Ortyqyoc01ctiDS
N1n+kN+8KnXXs8L0SAzJ/STkBdL3g2f6QNUnwChDD/nxNx/ilnKR2Q29IgoQ
Bdt4vBwl33n0k3jMFdLoy5Fv4821+LMEFjN2IE+v+klMfiVTiR5VqkRKn5O1
/AY2d4YQaLj7R9n8HyvzZAobS8h3V2E2TNGuWsF2x5UfHvkc+7xOhHP4mg2x
pf+z1JvIWTWc406pA7wEOX59mbP3pyErsDE8drUnFNGncWKKFB84z5w8amM3
BDFTTpMsyQDj2PcZHtt8zF/etOC7WhVKUjBwjuTdGrnHPv8nh8GgNLQfCC1k
2iPYdk9WOdBWQ8h6HHw97bPDwdNsw5J7XP+HMgKw2Ol5DrA0TLtwBbWyVIBE
ww/vbEBs50BM0OtcpZbT7jkiQEvkm7Onoob+v7uTeaWaLYQ2qxmZJvsdIcho
wLfx83fs5g9RCwbVMc82yEB9B/hcpBBXmReNQQM94hWdCTyOdsaqDbuNVEgC
CUANfcbiwzXKxk+wv102JJjjoPHieCZpaCuGwituHij7PzJDoqh8LNpfeHTV
m+XUy4l6UglUOJubCZETMLWIOeh4XoMlJcxtukqJ88ZEFdk/c+wo0N1MQ39J
YS7DdD3+FjH8/H8pub6KU3y+6Yf4VoQCwCfmzV6DizpoiiI+6zwBVWQJjuCN
9WCsOhZFGadtHiTsvCq19uQdMtB5lcXZDrrZSt7yqRlBTErqOL4tmBrIYiwA
7pxtDOnmxhL0pms78Iw2dwks7Yo+VNgOu2BR3iQNAODr/2P9q1bJ4B/fBu52
wrtv16o4MczN9Af39953B76C5Tvk7/HN13hvltcx3GB+hKN/CPy0e9xJ+863
C8Cc2eztAL9akKAveHQVehOZ9/JE140xVSDBW3selqjuWhWpiQBbYRggjsP+
qYFJQhTf3mxCPc/EzEsdVJOJ3Cf+VeTBiWZ91/PhzLbpQ4jUcBw3ao2XAtNp
bNaaMo6TN5y6v3mfdxGddn9GozAbhcb2lJA+aHw8Ro0ot231pabe3Vt32Us/
CQPsc7+xIHnnaRXgjzA4HHxjNHZqaE1mV7oWBRO7t+a4KNpoyQMjXdHlv05g
8hDu4+djvcXedyFP8mUUOejv/3vGSK76tD3EE833s/YsD1U0ls6D2WhxBsLD
tkgWmrdjbzpnFaAEkqgVhruFgDNc8BINd4FZPLLoerm72gBDRh8Neaywlv/D
oUdK0XrYeC5o7mFoMYjX+iN7oQra+xJ2dXJMg0YXSTX+hnmabf1+i8tvBMmG
PQopdHJ1CQdBnrspxPuPLDkYdvpjU9EC8YthHpupLajWvfAXO0riXMsK1Gvt
1k6c8ycJv1zUaFbnl21wb9H5YHR9/TXQrfad47Rhantr+rRbX0HupOtrhG8m
zdZliS/aHurKLXtgqDe3UhhJCMBKWOcbhtOmtsCz2KGmGodfVlgaWNSQZyh2
NKDVXkdaPcC8XV52z9uvZuDnObOLpwapbQzVwsxL/C4sf4deY+9bdhn/T6KA
lrQoGOQwCLw+IZDFA31NShrijTBJVZi0hnjeRSW3rA8gq8gObApfbuUG6A9q
IJLN8HTzxy8jPIovvDqk44CvxeQDi847ikXX6fTZ89JlUcKqlP6+cNiUhyBC
tLOsHkmzZPWGa274Ymfwb24SMpx9SPMGEN/5MeqrI/DERo6OXx/g2/hfoeqH
o7uP1SEGD2N/Ghi9re6A9dK74wEWRbrriMmY3XYLfBW6wQumaRDeukxskt0m
eZE9/FHGKNt5l28vuly41ZaTtEb8aSk4ZqQH0G3jGHY1MSvEBWhXg8Sw4bq8
N/7WFDb5HShw5WOqj2bscO1fNoqJVPPdNYJjzaT1Uk9zMdOrRW7eKg3c07cu
b9IFa2HTuVUdPA84bvRHkNvCoyrcYrLEc5q7+L56Ulu5/LcBDpkufimo9VEJ
eFTLDpJqEPmgqymiszyzcxYYlepImaVoIQ0hsguXg92eWd7BVF5gS1Yx6DlX
MV5LXiT1hODBDSucU0LmoTWn6rS10vAnfJOa6OCjBLqAqCaEgAD+gCDacZdq
+v99Oq/fYXy1kdXTVCol1pQpV5aRZ5wJtB2aqzgjRs0ClwBy1KjS8FNIyXce
4XFP3iTy6GicCGHPKliT2ARVQH1IKR0YHKceIgxFnrqpza3qBrjShP38JDSd
u6f5ozHf20S9mtXHrpFpk1/Zx5xkMWB1sUTDN/O51Qy08PeZlHMTJb1nqLm+
cgPstjz27QJ263V4y/YiC5VZlWBtPuAocBlL+TxdncL6VgDq9V165w+y5W3r
iH8CGDLKnhiVNWoLNH2RaOamNpPYGAvfqTt8ZDgLGdSkfIOP0VZRmKH4pBfL
AtziiCWg4Y+Au2ipS5ZFOyUcF18+pbZccUDuCovSE+E4LrAyHNlXHKB4/xCL
vyhwknMQitAMYa5uN6mvJ9megi7mdWuVBLhFR7rwkTmk3PEss2VPIadThIsq
d70YPfs7WpgoLXM7eGTMP5mM7LdYt7rVOV0GlSH2yoCPQVRZEUeOitS9XoM9
Dd2JxdsRsu/BW6JIBjpYDXEB7BXrki2wtSugv/Vdc13po3KCaFrsgjQcoiM7
yeAD4XC4nIv9enfw+7dzEvfM2gyxt3OcucwBCvCgEZxHWzvmsZqJD6gS4yA1
sjAajZ2BISqIRMx0YummzWFldgyb7pafTtknS27J9rm/1l5XSxEGAvOg0V/7
MBXNqM+1aqTU37XJE1b1a399xKgJF89K+z4jGq7dgNyKnYWHVpI6Lj/mqrTS
g2OIYNjEohUhHGsoMYEn5xyGd5DYHgkyXlqga0aF0Idl4zyuJREaEMK65jid
GkdmnldDA4n9kzXX4VyPvCU90UQtHkb1gigLcsKXeoLP8AtTEuhJNm13jDN/
Q5JKUkwYmcqStNUVFkqAlG1FnLEHqywDu+L2TmbVoLzbGn94qIgPUexEsbzb
lK+sqZIdBpKp2TUfdTibv0rxYSmuQqhAt9wmvYeLoTxyK7uE9xos1Uc2PJ94
xQdDKQyCQPJBgRwq7vEs+tRiAA5Lwl31lIl4hF88Nfjq8Lx4/9wGC3djfJWH
cWkLQbBQiURY//OxHkiNuoWI3CCxNLFGCIBE7HGmaTkShh0zmY7euSWON/SL
QDpdPpL7+wA7yAUOETR/+aIb9zqTq2FCdRPwOQUpUMyMuifXmlWAWub3tOLq
vWgJ9VbD/ikHyU/7YCBNj6UoEKEgyiApo/uOL5BjiHQyuULYqnQv7E+CV5B8
3HmHaS8H7J9GEmAj94aB4rxnj4+8KUP6Bcu2uEwYEblF12FNCCwcX47kdEt/
OF2QrDlGmInG4livsjff91auoRvRozL0+cdVhkmfGo9C+N2jShRKWYvPhos4
tBs0JT09VWqygvRPXvhPbU3CImSOefMAZgM88LuNEaemfk2nbrWaK8eGkfG6
Llu0GzZgMjPID+tE8L+5kI8EEC16az4GNFPBb5u0MKeJCsCEPtbIlQcemEts
0sR9VIwulQD7DdOuxcxj75erIz7l3MjARf1EWW/IMh8qnG+bkmD56ksTWcDI
UD7ZHU09zSUTwQxqKfWJgW1VK89KuvQQeBUFBHu5msUIPqLHOwMq5KVIH+9s
MXEKoPnjbsmICGI38stNkLDLRHYapk84MhoGMZp7e478ssUAgtue66V9G79/
YiI55vUVDL0DN86335lKZxJTEt8Wwes5OcEfiObMqWJU0yNN7ChVsfOoh9NQ
tV9EyCkgrfJJUN+25bueVjpFm7H06hzkVIHUqaVUh4/U1r6L7Rgxkmbr02qZ
hoAx6hBhyy8ZS09UuZ8Wes53iCo4vW1IQIJIhHI/d2h75gXEi3cU0Uglno0e
iKsSlXg8f4+iY5+2La98y6soS7zDu2S0V94EN2Tg1qKdIJhvs3m0aVKPB4wp
Zs7Zon56VtQVc/BKLrqZGNYpoXsKSeTahugZ/pySnlov9x0KTgZxYQiljGYX
ngBnR7lB+Fh/WToB9W1dXwjh7UQ3Z4XJvhvytm6Ge+04HLXP6Ha660DEKD5l
6Ad8x6ay6iuTLaE2LfWkxJJcWIY/95AAaIg8bjAbI5qNNItjLShVUw6kkMwT
OsOHbYfGkjfDiaE7SZmgmM8+66N8BNJjdYQb4kNht9pNRo0XrjAwUxX3/zd7
Gw/DwY3xA6FYhPDCostt59PKRi9IlpU8+PBK6Z1ptsN+fsPAgpt0P+d2Mtkm
Pq6y9iP2cXaz2933uipyNVQQgbGmVB0FRtV0fFjguGItm/KPebgOVoF9I4jb
kTpAtZdPIv35TyUKassvHxxIBGdxTVOLfOKENPJuvJSQs2wbzgN9dbnljvhp
YfdDG4wA9jCNxgEl5VimbFkJHUwjxDV8H4O8uM/BftH6aFuph+4bZ5sj9Eg6
j8ec6HNQTzMs4qBh4w9BvyV0h+1zAC1aOcSes/4YJzZuXpnAWPWsVmnLlnEo
xPzJ3nZHemiJSenND8g1YuTFnsyioHLFwgTaNEOciFFtNvvTzl07R4IQpUvm
YWe1EeoDAgu+30IT80JZRagm7PtrXMy5KsX4TEsF9UD2sT9ZtzjHvNnlGEgk
oPIB+20olWI+aBxoAh1fbmiCEq8EP3v+juFXzZyM+7iFhXLdDX00Wbzjkj5z
EbQTI1oECXNFNNMPa82vfEPUVxYI9yoO7HXN4fBI6vEjf6EMBiaNtJDrDF7Q
EAdr58Rfl0nG/cpmHX0NpFHrU3+oiNc8YWU6msoS7U87sHbMGqriGwTYR6Ie
zni3fyqBiIkHaxnYPrDwXWHxnh87NH3AlAf1eUQ4seWC3IrOdrkXXDLjkCVC
UD/z4Z+TLsIRRL6rpi1gztT3RcFS2/wWBOPcgE9XgJDsbOLSHjxwiWjgd5DR
i56QWUZu1KqmcJWl7eomvYAXUotaPF8epi/gAptZZp6lb2SVxyuHlsVP+IKP
+6fRNttBRh0yGk0x7o6ytB6vDc9DPZHvIHcza02dTJrRgc8KzWbJQ7lxWjAa
jW2lV8iNmOulb0gokWMiYymKWAcs2C4mSU9nz8p4OrycPC8//bJ9AX1PIzzR
tylTqb6n4pfdyWlBh2tjp7hCYFg1phKn4td9RZa/Gw3Q/SEREbfGTPa+FDcY
7NnYVVWBsbLLVzMVGSIMScgIrrnBYpaCTI+7SNQIRHTa2lxx9pETYLcODIO+
qzdGP1TVIfgfpyyYiipdziFOnIWkQ3LFTBraVh7VRJk2zV8bX2vs1o79uyoG
ohs/N4bs9QB4uwxhcZefmHVFxpVjcMyFFDsb1aN9W+ySK4F01U36ytA06lBM
VLSw8zvRBZ2Ev1Rtv/MYiiOxoyy4kZ797/e3IAXgh2iuIk1BZelZA1uF9b9x
mODjSrGZA3Sp9QM8CMAeA2edtpv3La0kBylEL7zfhSRc+qjBi9abqRhysJUS
QQzAvw3oxB8Le69aDCyQ8NNutXYMZTFt+t/oMEKBz+IVlKLtpu3ZG/LDdZRh
K8CYKEcGPZP/TcemiYQl4C/Ihfcj0mWZ1WweeXOC4VGAGhFmxRsjkbVxoKxX
LH14UBG6GB4nXX5IcNE/ZuIsmc8LVRVsdY6haM+XXNxEpHgfs3NTxf6tECj9
kGrU8FRQEa3SFe9A8Bidv0nJmyR8xqHlF118+7Jt48EXe2oD/IdBAuouaa2Q
4u3UrIhD4fvHJI3KNAuJ1uua96s6oEbSjP5vLt36l9JLcC54cjo/lk1Kz2c0
77YCCLfGTUzSofvkkh/uSp3FFw8FgDfECGWJK42TN6YvtGKESp2EEn06W/MJ
wUPEZb4bqE4Fs+q352dsG5Oo8evEfF2DjjVCEOfC47kqUhYV5ceGsrRGtaH3
61Nr5jJgDfERNH5ifwY8U9Lno/UmWIvfx3JUPlMqA8PaYIfsQ757RsShe5O5
yCVGooEY+w5tCKO7pZ0mIDZISBdETOnTE/QZ3rJU2uQe81C8ssazEOQxyV5k
KDhqrVEvS7CO4GWQEgki3yxRJsb+IblVOZkNb7NIbHAzlpL8RQJV3dbPOFNw
Ylku77kYYhvy4MgxiKR8LBjng2jD24SacxgZyucHzUNZxX9iQzjeEsDCrAdl
1P8q/4//RT9R8a9+hvE/Lt67GejLrvap4kdRymf7PR/7DL45LRrG5RmWdQ1T
W51FtFE9kTxyPCXHuD9WdOSBTEYg9caZjOfxkOQsmpfXLrUBEHmRAE5CxXfy
iakrnl9Kzor1bC+j702Q7ImkkTeaknzpis5JV4wigRZxiKAoQyZnRB1OIZti
eMPAk8VoMlaDPHyDxbWwd1+bYX1NktRhiAoMpWoe9rufYiZkKiErq/ErkxTw
j33bEX4EdlGtgROm5+Wxkc0lMTl7D2lFFQf58xPhSl05ODqrv3c+L2srHAeW
JM2fWxe28vOau+7xT3qsebD2Csp1tos4+cRzPd1FLF1K75vKltQbiclCtIuq
2VB/CQMQneepP/ISDOsd6bFn8vE7DlUVdRJYylZ4MHYlfCKnbkHwBvpsPCx9
LRDGlTkeT5IyrmOMuDX6x4TPLeiZ8Vsbp1G94RGZ1eEguZcnwfUezWhIL1M6
PdDw4f24IejJdfppkbOTASdy1cCchwnlUgZt+JodnAlzTGuMCCPHF1sQw9NF
Yh9ftO1GF8ZtvhJZYWqSFoQ9sv8wR0Wg1wZ9p4czY7S3aMli3EKWpJSdX7Vd
rBHSKHr9EJxzyhFxNdTZu6gSc1UNSzzkIZDG9kC2pYIWu6vmxAOYX//cLx6a
a2h1aK0NFy6BgE2volV3xIYfbVaL5MkEjLXAj32833JRnyqgNY4hkSte0XYr
tUQFEI56r32UgLYKWekaA4y/FS4PS7ydl7R/ZHikj8imNKMOqzG8ca/sNvfx
ET8coEx8gvzQetNrMs5d/+ZuYYL3xUtzETm4Jk5JAQwV7cgegdCwUrbVLq66
zjqImbMlHvPbibAJQaZeJxjOiouXdD+RZ1PwJfEbooIF8TY6cJMIXNfEjMnp
btvqIC7/PQGkVyF51jkR/wiDjY8Tqo/0sWcvb11pxQiaTfhgMYGeku+jc/nH
OhJKBSY55fxf60CLNIsPGxL1FWJB4n5FUmfKAj0tNiZQLlts/XsK7TRwIMiF
ws1t6lh00efaY2h4yXB4Zo5F6SLmHFDvXt4BEZW7JAGjseQapJ1oT4UYwPYA
kQ5F4B/u5WBXLW+j4v4T/JcrYwa6UI7XO4ZmvaGO6W+mpJbVg61PSGqIwVoJ
3jPSvJpZ0PvHv3zfLBCGfWtq7CpgtqEe+GLJyNmAZBXNURhxLgEhCyI8eiM6
y/1VgoO14X+G5YMC5xGZcQ8/otIxbcnSTqAY8k39YqcYCZgWMJLER6iWNfXj
R8DU+bvMYon45h8hkBZpPHxRG2ptA4kS4BXI1HfzWCs0dCHkarCd3uO37zE7
feFAAY8kb4r66cxFNxdx1aq+7OOHEZDVl8iGCtD3Gp8DP/hmHgHQ7Ro5zJwI
D+5v7CGnQRvi+GJ7idr2mxoYNjZMF7nfIvmWBY3VatXE6tAwYDAjz24aHyiY
ImcFkXqnHdHTagX8cS/e+0klEoSDCXKVmD55VeEV7EsqiahMwcVpzzPz90BC
sozaGfEFbMsO5umtToJNy+WCA7DAh93leHBQvXT6yy0VzKUbS/D2615NQcHI
HBI0grzH/pUt/1JLBQ7n2Hp2itbRaT71lApyAr37Lo75h660mMN+DgdiE29m
MpLEQPZts/lyWt7ayZNx9xT4dF3c6BslyHt0lMngOGqgeQdGuFQswJw7dqO5
lMwF5LfjwrTZKZPnRSdu6/RDjU1KjP+DqP2jabdf7mO48yO1vAiDSxGh4WcM
Zr5Wo/Br9HHxYGO3uGbSs3if0f+iYk87Jc1hH26rhuyaBKGg29Q3pMrIDB1l
bC9++AkYLAhprMecgwCYG3dQYPcKTi5/H8ipRQKKlsXI94SSqDHxnVkaQirQ
ikpr4AOjKGCIqx6MY2UtdvRiwppm0FnofVfVkijrUXdVMvkDY+Or/1URq9mW
bLa/6wyRR4Mmc/LrL1dBeGShYQiQloBdd5X2bXfnFTyX5tP5DOfJU5i90TPK
8Lae8DeFv0C6tUKmP+D81h6XHamLuQHMIR2TF2d1TzlOkVRcPBtjM+Un9484
Rh1RFpn2IdIM4Nfo4t1xKellgE/qJxvr4av1rQULimFHPwEkSMBBdBkbtYrl
yUZv9HXczOVJz1LAkVDjACnciQZOfYSnDqwj0A6y3zzWHGTjiX7ZzBnikbtW
oS8ugHACl1WyMfdnnAV6FwiwyFcQE8LU+xFPBEfMscdq/l/xwi5nExRu1oJ0
o3e62nZLpccu1VWO/HWwlmcDb9jJYP2dQQsgpeq+4Ciou2ZSG8bWGtnaithC
zA1doCAeIAykkNYJ2Sof4Z751hVNP6utcol9+xYD5n0zgtz/75ak88MfLK5o
/+Fuu2nypKnloU3qIKqMFYCFSVoMs4WQla7j3znuyRmWLqzqIAqK7KSfBG0a
Rp9lDGwvj+sGOeOb4fiTo9k6/oI0oyy4V4xl9qzAnt20GBozjEzQh9B2N169
EXrBHApXe+/hICpiq2dbj1qYVRIEaoVROWx4yNV8G4p+UXrRabNcUSyvXxsr
fIRMS7Zw3UEAMRAqJz3Nbzl/e0tVyUPvE0sR2n0OAAq35RKMNAxk66WVrl7A
SJN1YjFUVXuNTwLzBe14jP2KSRZYMLqAp/6PJ7yd4iSu+BtRDJf7jX0WHkOv
KLX1b9r/PKXtkjMrJPHc0hCuizbYRJO2OhCpwfQCsvmtVKOEIp91jdkkkHeR
HAoTAbT+V7wJfCuXxiBreJ/y9SwknIcSra0AmYZ0l0SmwMpfxP0hw6dJAlQg
rWhozj0j4JZn8Oet10di1/fUeiS2/LJmfQaHRiZQNdAU6WLWSGmuE5Ss4aSH
98bMpwYKmWMjX0q06BLvwozwil7rBhI0OcOqWudI/HLpk750At6IFpn8m1I0
l3+rFuZwZBJJ0zzVgZNr58QUhTlc1GlbNXKzos/jG+qgklvjYex8KDfnRkyw
iZCjbqp28J08oPzi+2RLHEt0qXlDCvfCLmaIFZAtL6y2rrauEYC/0jRX+ucM
hgSuFyII67Cprf+w/fbCcnV3VPnO3pLqQzyNQFIA66r6C0T/l7j5Yuzo8Hpt
9xyPDM6WQ6PoKt6YfxxXRME5ItpneJMmht1/g7dX9Rijq4fu6BVG+y54Sg1/
kBGaIah13Tp9aUyb5/UE6HdmAFTElU4CvY239EBm2odbsYDWOPEQaHXkvM83
jCRH8hi1/sLxEjadd8mRmj0xDMJGBYBKyzF8YdGajWGt0rhETY5ijbXAbcBc
X1vmUJFPTzboWuWXZRNCWQEJxZp6CPbUrXzMV0NOJfhDdA++kWtfR13fOHs1
K/yECxeNBOK7s/7EkB+EGlTh5PPcBU6pfbgacoH6TP8czuo+kJghzdkRfbxk
X5R6s21GZI7eLRHNEi4liXpoCi9ta1a5T4dH52aHZQHcbu/2g/DqXgmp0QXG
OndcnXen5Xt2t9uryI5E+JlhPmcf2dh16UiRqRFWRpXnZE3SAHYHKneklm6d
P+O9TSE9BcH3cryjYBpEvhZ38lgw8uKbRPm/WlkXeNFVFKxOI9Wa6elFA2fv
gM9xA+ktj+OKiXTbCsHqf3ZwkEjcitlKvqPrSp8ol9nafhKtnFXevED+7RL+
kmOMdyKbcOKlDcXRTJv1CtPnod9tUYeGPOkAlBfx1MpxfNmbw8cw6Mde5BzT
qHvRchhqKnmy4n4VOtfc2tbUywcrmaH3HJQd3LZWibatktXZTUS3HzslS+AQ
eIATEVx6ydFzay/F0+poPQtpt+FXdfSF8wQV8lSJOgnUjzlu5CBsoNfiz1l+
D1JWV2BKsMbPlJeZapokYaTNpKzKaZF8x3e6Eteg35WFy6e346mVGM0CiiWD
YuDdCA7A83xC8gApdL8th0nuHTRMPMzIksh+ebhEg9SXIoOqUVj2yx1QBUOi
lnIosJJbb6tZdufDB+MWZ7/QDvVMvTAWfxM7mmSTgsSyW434DzRWuCZedN9E
KSzNQa48ZqUPopJnhwyGre80dDguspYd4Z+Xs73xKYzWmlPblxczuCkNj43Q
UbdVjNMYKOHL+oGjNQ+uoFbdsnTWqZ06EnmudaJ/r/qXXFiswFur3eJsB4Q8
YjJSxhSTVG6heQGiTuBba5lXERXllJz49SbZ74YFPwEp/ZzPPBt8tlDIIaNE
jagmW+8FCVeYMDXK/94nNRMd1+1R/knXpEMmG0ad1wkQT3x7yoVth54EB7mP
6gfHpixQUtESlZTc0ifuLE5JIc+HPy2J7bcvMFyocq6POxXXDopi2Tt6mnkC
FDtejZyhXq3GCJCmnhZplLhtQ7WM7trxxX6ZLwnqFmv4GAEtyFU+/x76pzD8
chTCfbJxmP+j1L1tIoJeC3XsV6rEMgu99QDplIgSRVnQjGgXNNi1zg5flf59
nzjd4mGFEPgFpdEyNYZrcUksxk0UGOvvpKrUuvXFoYkNGk2dsYAE9Nu/qymZ
vxCAOqJqKGaG+gnvHy7H36r35YkIJ6fWkjEcx4APF8UwLVm9NhaL+IMmN/jX
I0FjNLhiA320VLjec5oazUnDU8ROdfASfBctnwVRaagr2mT3mN19Ypky5hYY
eLxQUeemo0MyBWQU01aUkRp9wBuekVYoXvAoyt6tAnCY1POkTWvlBdmDM9IB
QQKzGtUc0iPNeDskPXsqnK5yraFpBo07qzcRin8Up4cux88ym1drl+bELRWl
D90GJOCwEhtvqaFqrSu1BWIsuZoEv1XQgnlXy9tHAJfrnmwTV41BsDw52+/T
x2WPXVVBCoLlShH8LNniDqni/E4WWWDiXAX+BLJNJRjkMMfK6YVE6sPPaDpz
gR9O8h53G+QvMqPR7UOD2ftudPlyCmBU8rYnZS34SDV1YJBPISgAbb6fMoym
YQ/MCV4oNr4/BlhS8fkSx5yOi2GRtLMp4Vx7GiIpszM8OlXWMt2+/fLTgu87
J6CEGUbR5fvSWCplbWPhes3GnVNC5xkcyJN88/lj9Q9Wwutn7wk3NP1mu770
JAvSv94YHX52+UMVIUjQZGBI4uBaTZrO0oq8cOQ7I4DjNMFu0APAJNNetIVm
Q2Kvwg/ncv9QSarFkCT87kkdG8gCNctU8yJ8NgHXlX81lg7IIYZ0CizcsrpJ
T41j0lE8QMQXzfS53S9U/p0ray4TvgVAN4rOj9o8ToSn0W/0Li3YBSeHmCQS
d7HEvZhqCH7FpqdlU/Wp8zxO/GYVSVD4ws0TCk4TB4YAFuoEM8Fff4JsuH1Q
c8N6NZROFeGhEus/QjUJ9/RXFlp4XBEmfIxDwX/ajpe5ehYd87ZCFJ43U9My
PMQZz+JABDQbBibrwPmKB/RNDUvMNa6xrW3q3LdJH2qFufMQZ4kOxuHosMU8
ydcyTnwHEt6apxyA+WoHqbqhoAi4h6aJj8xbuxrBzTHDF5orKg9QN++Bv0sF
6+nU6tk9YCc7omDsa0UIuT5d6MvnmjFAIs6cgThKuTQ48NkvhZbENokYbqQb
NUmeQFXZ33iF0TXMBnzbKdQ6Aa3ZYHDvGKfBNynsqCOGLHDbhmaW71BBQkJ3
o5i7klpjTM4Z1mYNspwA/+KI1JgrDcRYtoEbVPXxha/Yrv2BsiGD15SfBwVf
RFIiX+mhKvAxEx5IfFNKDvxwywYoFtkcVL7BILSNkR5B4s2QniCj4dRpZLQ3
Q6rQ0NsUzQbUu963uQ9oEY4TagjYZteNWBoKOtUM11tVPodu7wP5fuIBDBhb
U9hHQycybRCzocDllEnjG5OkdrBnY65A7OYlMoJ12r/KnzbA/UtzjOwLNxM4
2reo7Vg1PJi5GxpNCMSYH63ueTVYJbDn+tH2F55sw1F7mVPISeM2+cMwGWbI
LbcEQ5DP8x7e9SQNB4PtUojmxx163BkZy9OB4xv8gF6zoQvfOWqlLld1kK1D
hpHtPJkKAZE2zZCYgZ8tXfjVjof04OOt9fk6CLmuZoXdvm7gu8YUu6bSQICk
0tIAVbHM31YnNjKYcSUpprSwzjb/yRj6SrJbqSneP4At7Rw2EqsJL7NBNkfL
+Sp2zZbEiesiQaI00MmDwodleVS4xqhVYTvu/kHJVqFCjhFTcqM0pn8hdso3
7Trhw8PNO5g1NNMGQs4eBRVpsuLKggdJt0w2u6vTuxm14JsXJd4mmIVX6H9c
0oWX8toe4HPsIkU3B35m8+Yla16cv4dbxKoaG+m33TteYOJDaUMgdq8g4GYm
vglJfPwjDAQVDQTFc1yEwibMm9ajLIT8149EEDmZAbvmjMny/SCjeDc0GOZ5
zrTBzA5TI9m21RbYwbC2GIwnZBv6vW5PlO5D/8dfFdahHWiPN9yqofSkfCwX
gL6H2zvYN+H8ihrOkRWJ9DSK1qHhPWg/BWHWYlQdPz4kVmlCcj0X87cjKUbp
dA6TpZXfG9Exk95VabjySrQjiEz1XVB89LzGIyNzinrXGN17copZJ6z1Xd5p
B1dQYVaPkRd44pTsj7ifMYuY0lQ5wiwISx+36sPhUuNdNGgUlhCW0xHOZWmC
mv5PQSeWc0wVSXYp2eW2rMY4Q6Tep/pgr58fpbhlXNqNOP0CctKgl5G+BxzF
xBcB/WoEOYSXdZ8BBVeXDkiXaIs7XvfiJxDNLVdrK86MmGNLXdef+a56qZg8
Dxp6DzX/tFlpob3tW2HucrFh3SM/JQKnTkSbbEDy7LNTT+NFGT9lFR7e2SaU
fynvYZi2mr2DLFh7nYsYVQxaT6izLJCVqHcPFIIvM2srMUhTk2oIuMPfCt11
wBdgPGfPhm96BA1GZ3940uYtF+Cf3BwTR82F2doNNA5VmRNhzDh7U0vxpok4
Lx0oLlJOadHAQuP0UhFnpcnzfWTzCfybVGwXeXnMZ25wXTpP8KtZSvojKgFq
ipIKWnB+ZGVWz6s2FCDE3C0j377P6OCeilPwtahuDoqBd5khZ+Y/WHtrGrty
ZiTJY2RKyzrHG9LpY3GGJsqhNSUz7jlHlNPELosWAx/yZQbtAwo9qKH9Piw2
XvM69BittdszA5Ry1J80he1j8ikSmNPz7/EOQGnsFl/9pUD5hhNZvzBjB8fq
5RRZ4i5UHPBS1WYgus8atCj02R2O2JhS6XGyw/xB+3TaRA6PLE4u4vJdYFxK
w8G+PZj/ccfeq/32k8xa7F7d8X/ybrPkWqBWXRz3nSGBTpcCA4et8MHEdCQd
z7SxTS+uQP9sRRsEdPkvH/YoFaa05J042r+Q0/ZsdlS55MGtjpivS74BByMe
HPmXSxtYiPXx4L+wEIly0Pv0aLYWkyBJ+MoOb+Mpdq+R4Vo/stPIjhueLhfL
RMXxcUU+S/aKZVH+3imVnyPiGIUyJPw+mgIPaEqjQR5bOJkkGkYCyCcEc+Mj
AYPh8J80dO2LFlpHsz7ameZQrF5kduCWX1HZ2BXzFPvDaDl5sutquDf0K5du
sNSLQmHZn50CqwD7jgDv/JoQ61EYQ0UfLvuGiTovSxMt24dQYZJNTp51ZT3N
0zihh7vl52PSancMhdxwHOZ0MlFb38Z636bjktRWO8qdhDk9qjPsdKu6L4B5
EJsgsLjDPXwHfKCceOYkyrUOJvdKAoYi378SwYo1xQexhqLa0Hfr4B6qIROK
JvHr4UWezVkSLZHvOQh999hCgeQ3AJX9+JFpCYAUpds8RAh85jNeXSaH2uQy
u2HAgfPJpi6nxS844jPm4QUoNvQKSvXrZf75jUX0344N7FQzGhgaCR/uBYyL
PsH6nz61sbYuKGktAWT6+Elxc+GAEnf+jC0xXpUYAXe5qj4Z5eRpnvW4jot0
r7hNMGC3k+JycK2yF06JGSMd7ymcO5Lgf7rkG1pdx7B1xg9U9vxe3Ngl97KE
bfyxcKBhHFJWNHYqiz512OnaYJE3YXsgudU0rS6qcAFf4JoQraa3b75PBSSJ
Qvay2zc5yZkvEVutcPSMbB4pU3qBxVpeqoW1C97gItdTl/HtQos7LPSWYtIC
nYEBeE5E0sp5DuHSNHAvEiK5SKvAGqe/pwkzhFBiPLVWgCo14peVn4hZAXpG
nKoZ4QVKbDkxdy0ElttNFowGtirgGfRfVfD7I38n39uNErrY8z/KFHNZTLmv
LUfeiNKCE8hvOF8j8mE7kIPZ10ZSvY6boECAG1r5dH9QmSyygKgP5kNG3n+j
CgPO7oGMIiEPWQ7gfpTSjUp3vqqBlEJ/swqAOVQk55+tVZAZ/jGtsjlZqtyo
UGqMfcUrkkzcg9Mrz3LTodz4H53MSLp7JKO+o6SMSHQC7cHpxbK47EEdRQ3K
zpvjPM8h3kAklfgU4xEBEcCCcR84Q0fl7Kj+TSUP2ZPAQFUd2vJouQh6OMPL
2SfdbOsB1UfeqyKA3ipZsRLrfzs4fVY2MiVpOSnkiB2zIb5XB5hJxzdt+VN5
ctieve8YpL7WGPyHom4I2R71ZoPPjaRvPnpRpcekHq9uni/kHpkUKBD/Vhia
CbIpg6hRoc4F/7iQh2l7GaD3vFxSmaWAigz7QdtoNT8p1E8rPt9gbOXuwEzT
AdtrOKpEjuun6bnoEqcxpDiCF4SNVXNNbkAKFnhmk+HrZqunwhJVVyljRxZG
mwttT4S7N1/OyRMv3voObXOrzwo2GVb1GpQ2Zp4onbxEqA7+76beCg45y6nR
vvsinj29uAuNaiNN7LoEuPjItmgQcCtVXN3OuhfiRT8oSu4OuQIRtWwfMjbn
L230cF5fRQiNzRBS1I4qqCOINHGmJken0NqHAYdRL3k4efKRykKlptapc0b2
iOB43T6qScUbxN7CaeNcb8+psD722q2246rYg+qyxICX5Dto+v/ECbZ+F3WS
P7rEUHCppcng7fFOS8mPJWhpXY0lgCJugPl9EywSkN2SiOoRaNjTQ2eKG9xe
+dC3DGENfJiZekeuV2P66AlP9Ls8LXkqQXDYqbdfRx1eE4B5e49NSoTO0MOI
in4lunsvEz83VE+wOKZnp2pifoMVzxpDIUpBgkWAxp+0S17X9yn6MOsP6wn3
YgDJp8Q5r8iEycJYgGxsr/BccpBV7PWZFnKFX/N7SRu/z8drS8Yeyldn3/0s
wqoRzn2kTW1L7dSdJfTvMJe28pFXEb1oJboqoXnumdQpv0WL23lORZLUvhjq
a32tnWHrn/fDiWP21SMFMkyF1vt6r7xhMdph/OUWrHiTiYV6p8hoRxiKdaLt
OZs0m6U9ScTYIP+9Vk8YPPO7jZtuwznveTzK3Fz8cHD8q+aUMg+2BPCgfhvO
M0tIfNTATLHwTUvwGE7FmWqkx3Q3szwndKwawERg+dOnlArzKEK/2CMOHhHL
zlSE0wOZc1HqgFmvbbdVoaSBYozyBWolh1BUzZy4+5L+sg6bAszGCF4G62lS
l1QVdFCpo04wz6LFfwaFwR0dQDtGp2C2QMPw+rT1/QCvtqLztpxcvQJI7aWH
acX3zguFnUCnTsEmpDhq0AuCCjLevXfHJ+6HgaV5fbwGmDoywFFnwpu8uEsx
7cuNX9S6CAXkyRK7R1zDte3W4at9atdr+ngtE2K7DWfMlAOKXPr5p6/AIME6
PrK9ej0xgaBsGdCKhB/MUzNDFyTx/YxY6Ix4glp27/89MGRpIHqGFhHpGDE5
v/OdpK5f3iqLlBtbKB+wfTf0pHS7kXiksZrhar2nE8t/YSP0b/qlE5w+91SY
lVBRm1AWrmOHUVrZ+YtrtcLedUMrZZe7eLFXaXOMxmDaAk/P5288K8s51tXj
Z/yutG+44ex++ROvaE+mnGhFMUxwCr+IGjaxfTDQS+NYlUKCKD4+7KmK6TcP
JyNMLMGh23zn/gJfhjh4Kw1Nor8MrrTtn8N6MYTR14o+Ts+TELX85z1lb92u
6oCsp0yErThYJ4a8OTTMJ4jGC3Ha80YsmbL/fZiHCIrxLcwxdAouZHpkNgJd
4duYUN0k8pGw0Su/s0hsSe7f2VaPU5iFp4upPfhR5TrfQ5ojDkf2GCoLhJPO
r5ZrsmJ7jNG+jZg8HuAWuhr8eFE/3j4xPt6AuTYt+i/a8mWzCSHYKKQRnD7U
44884P1okPb15RwwnMXk8kXJnXD8EQ34+sIqk0jGtpMnITa0BBysQYCMp9XI
EeDE203c2e+NQWQEmuSnDGbWDFagl5sNAum+Kv57QmrduWGIy1L29/JwAFab
UG89D8GVNBNMPIhOW3R+gJfcYMoxPxX7hc3TPVP9WUzxx1JWPABHn80XUdij
iPvvbok2yyASPsaNLfmQ6JYkq7/LXDF6zBl7h7juvBG/Iu8u6w3YCf3Rwg00
CtOi8g6Dx3ti3fYKeRyhQe0gpQAeNWIC0bfST884Nvp8LdWBuo6iXoOBkdI1
Y70Dps2wX2ShercgpbM/zrVhRPIFLSowPBPvVDYNUMchLBr8WpK/UtkfysYb
JLHaxAEbLs5gPh+a5qdbviQsloCy8UIAD/rnFkjYoVqn2SdtHlUACJwQWCOm
m4pg/VnN4pZeAAGBTbCUDshn2+jw4VVpT7GnL2MBNaR9nNfdBfy/+Q62dFEt
VFhNKNc7cbABXGqpTKLeU7bpcowNhG/BB2uniPDwSu6/zVPampXmzanAobsJ
V/UyS9Nm+BrxC5RpLPhUCmkSrBXM4WS/+0F3RyNoeKe2tqGU2c8oNzSUgCXl
rt7vTL7ExJLzUiadJ72DXnodFHdvJ4MZiwM9VqHN6GfBHW/hcTZXJ1T0Mae9
u+Zf8b1iaOjsDkjniEWsC6ifI/ZDTfL6uz92Nz8J8378P3i+FjzvET7aZoaV
iMivOSahtQvzYsrghmXG0AAulMe/x6gD/cnCSl3rHYwavqJYth0grQVTpheM
KF8Pap52KnNI+Uvig0YT25sLqQzBMDA9fWFN22DHNejG81CgESQqPBEey2po
Sd/+XEmtFR4ZlqOoq0EVOg/C898wP8GU1tFTdT+mmIv1sFj01my7XSPdlEG1
QZi/S8YjIreYmFqE1ZuERPApRg2vOwHuGC092YHnsN4XS4Nfkq9Yr1TtaWEl
q62bTNkObkzO+kdRROwFOFTmzsW5MibRmNYFFg4V3GnE4iTPvE2noh8ecxE6
kWTdrxAhd9vRoaEnJ1R1xOcVtZzPKBB8h0J1xJahg7o/iGoyVXZDhcTbzgMf
kY/e3MArvKnuGlFPs9oDN38H/oYcw5dUPQbTRf7TBxNXMQu4YfoODuKD63oK
U4C7WRgYGZfGCVNhTnymA/Dt+wuYT9N7MQvNutJw4KlvQoPJBGb1XyDj6nMd
g97nDn71Nxy/+5kNa5T5ibH3QZsbyrjfs15IQWC4jN1z37LdXFHVkamOSedB
lQsAlkaZxIf5G6v8PH8PuRJ2ihbu0mV0tWMd+5+2pYcBOLo97noIWG+ohz36
ekMeGu/w66TtzOXATNMg+WcSouMuEDGofhS432416MPQBTyaqzBqPaSKrjDU
Cik/7aiKtMNcXugvEuPI5lfcPjDD9uybAEaigU3uhOfPR/n0aaI5vt/hLfgG
EnOMysldQD/DhaIxTmbVCzlNK1WH8BMIwdv/Q6j1YN2pVG7bPeNaq+Z6vU9k
/J0E2gthCnNmfppWs5R9vPbzSUrEEc5l/lkXfU9Bg1y5zuFtdqcHtON0V86E
x78/BZQmYBr8KXvQ0TzXWN9f+yVeHHDYQ3x8rihs8eYxSqsqDewonyBVrSRB
9Fdrcngj/ZP49kaYSSRoXZaaJcdDFafNU76Z8v6Fb7/J49axANuxsi/rezKl
Q1BS3R4EvE4iOHjHzsCVZqYQfcP2XNr7VT0TbU4qTFtE/wHJiNOV+3jxXaTQ
SNJmJw+KQHfrrOle2Jb9oFN/2KGVg6eYfzbhCoXWxQ1e97ZrzzX5ohnKv0Hw
RkOwbeCcb+GyDyt9omJofgL/gKInQP2/ApweVoppoe7uj6ezSPM4muGlIeuL
C0PUKnyel3GFTVVR9FmL3qtcHTAf6OQ38dEiTG5rocBJhyQUrYybuXzFWjNF
yCE+EtTWJUSf/FbjIxnyXLoNR8hhD0p0kemcdNPQPcg0mCIKL1XKJMxERUxm
UNMnUqJVw2jqMK69I3JiaW4knxw0y7DMa9PF8drZ7I6ZWculsmjVYLA2pAap
DWGFNY1DQhiByO9j2/I596OyQ9hmDCGpTdXoQQvnAtGHBHjeOJ77t5j4C4ly
JGvDmMfFQY2Dc0wAelIb2NgQQWQG3D3Ep5o/IWq11BEShaTwQt0vYnaUkzGm
vZcr7DPY1oPbRY0l68M8syLyNmlSDTIo+BCl2cCza2JX46i0c0rAxokpatPc
+HCtIkveluDtwAR14HZAoy4Zp2xSbWDN4HhEhg3dttjds/hIJ8O77jl7Hn8u
xCYtrlMnRZU9QeHrjYKtw2I0XxI+9SW1XJsefcxetzkATwtauhUaqHxyU+uk
aD/ZpjvFf9Uekgc91cXSkp/Z6DaWzdsMYbM3cISKTU+tuF8ydWb+IerVTb0v
37POTZVnj7zWonuiSDYV8ovP2HrmqVccpJO3aTsXbiTvnfqsb5hVP3CWl+3/
rwPNcP0/KMoSWzLV8KvIttxD4cxmDju5JhWEPq1/J/pu5ag0gCnC2Df9Lk57
XNqg46NKXhj61gPuNqb/9TI2rUtpDPMD08nx/n68Of4KWppFZHACYy9nz3b0
fCULOHM103+l4wK8trOq6jEAIl7uXOUfCr0WwiIkQUNoWLxUS/hKbJE9PY0v
lSSdA8BFtgCQts5XF9DHENxuGv3UuoxgH5v2enqlEVhX2JYuDZhRxxQs2wwx
62TEK33QeSJoIXAW6X4WHvQ5BZSPJ/45Wk0IrQ1rKvTA40pqujudRzGgKQ1q
Qb/JBTXc+c5HuQAQzb07PcpTEsPc0gVn1ZJwB2LNKIX4BbEmuQDtRpAxuWgT
X5AYA4lOzUy1iTII1L3QOIK1LrGI+quiBgaIWHUBpYBRZEpMwGKdgMbgEA91
z2xHUxmVLweJkwZAlj1HalQqCb69INBL7BjLRHlVQDsbc8rvbc42VZpwPuze
Yy2a7zbnim/FMNnHTQkMiA4wvjGwhP8Z7liDRMB7vw70snSGyHjFV7XP7ZZB
80F+7xDFwJvw5IJtCLU+OVspiAspS5zK1T0ub3h3d0KvBxKkUfeR70EWE6Sk
0saSRC8RX005BLNADofdCLIJIIGoPLbsSIyMnhsqLCPpqxtXUmXu0ngtjHRr
qmA7imXPf/yUwaTdFr/xPHzLJDZw76+lzxdmQ/f149pz7PTv9Gw/UfugDv4I
HpDZYA8fAE9sVxndULovhqIIYQmm/voRLjbECuDTvIKI00dXtSWevD7QWH/A
tvdAmLqpcKGt5VXkmhR278FooQtoC5Bd/FIah0g3m/dy/LPow8ss3BBXTtB3
pQ5g9FW3bERhUdBsjbgq6w4dV0Ii6gnW3aVdLP/QkD1Hqf1dz1DRjXjuRWKK
AauiUP8IEjxHXSd35dG0811ueDgtJBM/hS1LRHcqWzSyI3B5fsPITCaOBtnb
GK2CF7dHdxaaTd9Xwxe+SjzXIep5HR7eccoMvgpOPjpUzmIF4OlpJtr2mexn
mN/4Vpj0TTsNqRHITS+pp9Tj1k49xhNg5k8lQrMHlIG4ebc2ZLgxBmZ+m6/t
v4x7TKLH/ifVQK756U1xN8V9fJIOcxNIKb2GOWkpitXJfQnpu3M/CbGwoO23
aLMIK1sWE0JUZAMEJrwMb/43Kq6hyML+9uUYyDOnaueKMmFFzX0uUxr8o43d
tT0mkBqi4he+jAUwmKhCRT+zbUM8+wSQffTef9jseGkVnn+Yv9ZbT/hehNjW
MtjdktpI2Z47Z1lUr2FbH2sY/xkapS39ljW9sT8XlKwTze2pBxrE6j/nlg0D
wwi9XkPBe/Sa36cNx8KigWrGK8F5XD6IqQLjePMH8ps+t4Ju6YjLbyK7zxh5
bX+OPLPNM+X47DS5qkj5SOQAJ26cGoR8oMeayZIvoDH1VpfjVFendPIxqVbc
ZaNKi/9/VuddtuZAN8Q6kWDNW69gsDt9tYmyP5xvQF7hp+S1loMRT4hgp3fJ
6MP2vyWr2BPZOyu/W2BThdPjTu6TM7tBwzOTzRiq6SQQsqmwlSpLa0uOSr2F
Itn87d5KR9lcWp3qoh6aDDiOYvdtq858RSpWhUpxyr29PdQLsQs7ZUZRb6ol
lGo9v/LL6C6f4vmgmX3pFa386jsHITVJc0lPr6OQ3O0kWa0IdvOjXsp3naYY
iJBXKyh/iZa4kHqebxFoidFvctzxTtba5ROGx8rN2c8qetCjSiclnPLWqzZn
oiFEr9Ag09lkBWuD02ZJDq3MOqitp/imYTRhe3UySyXQjB8LaPpALUmBvajY
uxdyQvWFV+VTd+IAr7Rpy2NmfQn6+zkeZxcI1Yx7MCEYHmcahPHwUEVItvF2
XnIMIDnktMkBIOjylWJeogwvQF4k5BU+WHqrX3HDH4eIrbx9MuZ69+psSykS
wzASQ+L/VmJWHaaaqy3sSYtmAqeTi1dn+b3yLvQTc1HuXEI7lm3hpftM5QWW
nCuMGRWQmUm8VBC416RXgx7NKQxExDXzRJ2W96j4Jss86ZDvD4Qee0Z9J1/e
J42Cv+FFUev1mGZs2DtqNGxZ/D1e6HzuazUJanxq8+eswB0VVRU/GgI8NX2d
MEEOpBly/+AD8CS61CGJVcPXEiHFvEL6R3UC4ifQDjeJxucIGd1lH9DG7TRN
fC7bIG8Yebfa77hiZhjovy6h8wpWQfvwRtm3mQIKzHMeovL2VhGBqcYJ0h1X
dRc4ZOMlBbDTuA01UrnNdgXXTcH+eJN8B4AnuLDBT+3OTnTMTde907qujX56
liS0iGfg/Ev5JvwpGbKvEih4ShEvDi4YvGriXSy0Uo06h2x8vj3h1fy8XqEy
sjZEhJi4UOJD3I24uSgMSOxkIA2sGoamXyW/TVVz8J0Qz7bn/mEXrKVJ2qhB
34j8HYjfwGGRnSYtafDl4UBH082UijEjhGyyUKL5Ik1fEIAk4vkLbxiZUgau
m96uFLrFcvv30e5UB3n9DQrQp+ae7aF8BEytpAGP7VTbu47qiZy1tok2xuVM
JBUUO6e5rmImgJ5xxxP8gy5KWFFpNNKwOSMV62cYV5bXGkvXHnDsw/DdUy5a
s4ZFSQN981P7zJeylRzCmOd3CBsQMX/SzQshfVgBiBfDLueRzV71XbChWHzu
OUjvO/TZTKw1WwiHMOWZld68GDz78ndQUbaZSdndcYyqYaUWQpbApcsaeuiN
RiF80sALpU8fJfYrPa/pwPYyLL2bLmtFFULMDwN/bo9dmnOtxuLxkBhV/zc2
loBTFR+0oyREB3r2/RelMZyebI2AyJMk9REJgF6hn7rlVz+2lLgBAXS41paW
coNmb7gXMMkIgREYzSCNKpNCWuT3k8EhHwJjrpjJ/166bptGkjT4W1pXNn1W
jhix3mKGRz9FYLuYr0DawLk4zz5sUlYNNRdh5TMHwgdqzSOzozGvHQ1VJ/9C
ev6YNICjVBuErTzcUMlUV5dNV06Xyk3VQfAzAZSBQIFGLwN2WNjR1XmnLy1X
e2hMTc8u/pZ6IEdjLTvRx0AkSs7vqJQ1bm+epP64wV6SCfHBhO2iDbgCzFbR
kIoAD9sjTYNvjRSjuTCOs5jd0ipGrSX+rD6TCDxR+/XLXseAaSBsJLQd/0tb
vO7KSa4BL0Mc2NN9N20Sj0JmluJYpd3574uEqwPr/H7E7zqPUclCBGae6u2h
kQz+mtRDlfaE1AnLirTwMdk3AzNdRiGhs1V4AQoELZEsdsEwDN1+tF4Fznng
7mU2Omar22pDgw/jlsIiSuutU8HdqiAS2QQvDk4JYpG5osyPf/42nVv4WiJ4
D9icMHK9nG3exFL65N4VKBNWxWNoA5tZv5NcoPqlBVYhgNWlrLRaRBe5Y/ai
lEeiRiVT/Mm7O7sRqh1mZwMkE6mb1OPyRuMmu9WOEO+/pPGGkqtE+F+AOyuw
kngIE3gqa1ChiW/8BuEhIc5I1FODOMq2zPThNbsP98cgeXNgowAAIlmwST12
hRaqcMdPHYKb4HGadWLJm3A6IYBlpup4/u9hfx5pFVI+jd0eaaOZmAdSSM+G
dPiGKOwY4kIvAsrUD72JKzfYnukRrfXqILdw9c1eoLQqps/VV/fqje64jQu6
eiMnDocIqGS8gVV3QawlU1azagNQ37VpnEyz6gHmDNtMQ6yE7PKA1mk/vXBh
bBpwjey/moSNqAhJXQf58/EGzvyhBi3sHX930+oUB5h8SkWplOjJJFKbk/aE
NzaKTlHqVXPjTdMXD9LJqLgVYeWX2hIUJoVtVJVJHV69Ms3XAc/yoeMzyfh6
1JZCw+7A0660OiCRUL7YL+dOZlrMQ3NasQXlNYre/mE/mqLlrmwP0+Gk6zGX
RdhVlyzGGObM1PH3xToREcb9l4UboEDkzpc10iPwuAW0UAXcmo8mHUaawlyr
Z7Weev8q6bRkZ9hHOuk0Bm5DXkjBuPpfkWJHVQh2v2Kr+9mp+hKYqBgZcYWw
qvqynl8Qj9ptk/Cenem0MHJWNyt+9DPBh7k0QoHOdOVz9nlYOYnnBnSrre2z
EfFmfGtMLBVx4LwU1/Mgq8J1akVcMrohO2kqtTyJDoH1zkjpOJbpG5wa1Fuy
40VAi0o9Gj2VlDy1PzzWdjGFZp+QDvkHqSXNo6F+z44oVPxg0RvqmAYtPChL
Q9uQ/ck7qTy/8q6a5hRWKJgv7PqZCv5vULFpno3kBKXkn7x0cSESjZSs4IH1
3kra12J/ktc0NDHMt/GMqrRMu8tRi7qSNJeumahxRtBA4DDOOxtyHa7uJ699
GAayeZfIfm482+1UMZI4o7P2owEHkDUyxqlGOFyahEtXhCPZ9hG2Y32SYxGp
shGW+uM8kyp7boRrqJWVujaXuJSlwXlzj5YZgPtqtKxGlzICBOluruYlfTmj
GfPXAMyBya6yHi9Q/68kC9ff2nPQ+K3jsgRNN1JvubgPrmKswa8cjuMNamU8
EHZp3Z2uFiwPSx9aSZ6QThlAyIqITX6zxRdvY9IkvX0qzmJ5Spca7SycbpEO
fHsa5twPZC4GzyuKwlhRg2EMpQoupRHP5IK4WpszTlVzXASOohxmckDWCo/s
yX8DuhLCZhLLMdyjb8ggZYxzhUu7nOiKmG9f4NXnvt1fwmqj7xRcIu6ssNk8
1sqCtonGsLVt6ci5+/hntykjk10tJyLnT0vONGe9CKBzCTRWWIExj6xqjXYp
92wP+WUEHWjmhm06OB3nOp2gGP0d8WRlWbdEJkuy/75PSwDi1esb6lodq1Ao
89dFOIlKZFj5qO1QPLe06xfIzLBAeo0UUvqywyGp5sEWifY7KRnUUL++sxik
WkQaOhsS3H27jUM8ZQZnwxp9g5fdyLI1gmgCDKYsl7qMTeZGbxayDfhV9j1m
WanIUN/qZ2/2gnvH4cR+iQEdyXgAP3JFwxlOWZqSIXC9j+ePgFlLDDGV32yq
X6hhuvphmylgCGUHpGOibfVa/VESTw+2WK64hOO8mMNNQ/6hb+pLu5Yb/QoL
x2C6nYEjs+sWMHiPUb8q3DJsOygYXRdrv9PAO0lZ+nlqK3M/Bqn8qt9xIW9k
SJz6QotI1FjAGAIIXDTCMlhRdao+1WSRIH5igQRpAO3ZDM4giSHlbZqxY5zG
8q/x0rw0pJ4usb8dlAPsJMuhNlzIdMfiywT81ad/CK5e+hfF7IWmByXL4X9n
FORWV8+4O1NFt4u7Q6VaGGrS986n4sPFynXabcNX9ZnsR9K/OgqyM1x6wk/I
digzkcECDBn0ObJ12+ubu40K63M8V+WVA3LrGkbkvvbTq2KQzOzeoxfe+iee
QyYu6FUxRxNKGKXzifksKnrDqxxOart3n7oGgkq2/dhcYZoz2CRowFvV2OTW
0J/HpUIzyubwz2/EejQCCX/1t883xKcZFZeLOk3CrhrtlToPWIBMNZd8/b5o
Z5airr2mhUmQjutzMg0BCnw3cE0hx4gmR7aIlbFKuanTIlbJZTea0SSB9Dq8
XSCUkl2YofIhBX+5L5wQN6G3WH7zMWtKKL0hA8aApmFYQiQD0/WHxEUdTc2M
4AoybVHnDSh6r7HaO0bgao17RkRtU+VEEqfsTiZZPsHkLyUQqAhdICokdL6R
HlyYaxdn3gfufNTFHW9gBc6IbUlyo/PJpZIQbf9d3OW1y4VWt0OMcpi25Zfe
hTZh2xh8iSDhm4GKF5LrL+J+pmlyCpNG841kmJBwGU0rWa12KQ6h0trOv4Of
eIhVzpGA8O8Nv3iOrL26uB8vn7RjqCORXV+NX5TEO9Cgdg1PQz8ktF5eAtL1
7pNyDvtph9rY1akJe8pHbPOG0vqokDKnkx35y/WCO94xqVXnvlUsE+yQIl4S
T3N4boNvB0TSCVS8NZQelFHCquFnk4f6Mp+YggUi+iXNI0zWJ86TIqmto/it
vjfN9gQyPomn1lENWpxJauSE16UJ4Nt9PPetuoxe4vKKl8Zu3/6m69t7/pr6
jyeTJ2o0QluGgTd0pzZ4oBcv4l9HZdA5TmHWptLV/Owf8ofJrK8afFr0aXzW
b832T5CJgg0ffyEUUA+/zukvLQ47n7l9tdIXwb6RONOkxG23pbYVomsE0HSK
Awe4QqVIxxjnrzg5V1K1cDPYmFvm3C+1AGZfiLlY7CgHhzUbCtgf5NVAiM8+
IQ4dRiIKJ0mjUhSw4OPLNtsB4hjXaO/G3gNhQiqzHpeYN5V7+JQaG8bC+VG9
WeY1ToY9xu62GTd3qlLvGNEKhwqA2BKGPcmmuGdugxxiJrEF0QHIlQ9Hpcop
sGv2GclyfpShb3qMNWo9oFCQ6UyBhvYxZoB3ZSoHzHSF0pL+7OwYqnDWoiYG
CdjrahIW0+qMjfxvd6z97pSnQdbcynEvoK/rrMIT0mp/c5jwioMkYZ5LL4jF
Ad7xhusc9LWsX8xQYi3jnylMBelT5lucIexhGnHa51CpTO7lMOieID8HIQ90
jKhFMd6bpMx3RCUEBNgMpNb1QtW5OPRnrBdVVJGCDtzo/2swHyplY3xdkQTe
OJy/XIhWfuw9m/8FWiFV3RLZxqekXqU1T66WIXctbABXqeg0ELz6s2TNl+HN
jfEv4+TCyMVS8nM3aeB5Qju10kVSC9WYhPvDHIKFHwa2L5yElFSn+4CNDNkY
r9IXCLfWBalQycME57lcRUqUleXvlRN1CriO743Rv7RuBTB1Vkt4RM4CxIlH
2CNZzVfIMWGryKpRzJ/nUAO99sCQb0eSFHCJDPWzdnIVxjY629+RsONQZroN
GujNMxZ4XHbspgWO2wLtuOB1Z4yCcawa6oaJGnE3bX4X/gqFmFyWbQ6qfdbo
LwxC/L1WfYf8MT6RJSTdI6xhswgO9VmwFevbXtHdS/I3niAWOHL4yztVo/za
3yJIbzoHHZjU4hUfWD5R82hu9tBbCUwhPJEA0H7nIMaQ3rJOgfsr/BrJgG6k
SNT72GnVgU2p3T2v9zYJABnBuxV9hcIXc7NTQGc3fZnG3Y/6jMhk8vyWrJ9x
+OlirvgUluDbX1cCHmf20J3Sc6a4WMmKaaXukNDPkN6mA/uHWUVBcY+3Kqkj
2bElk2qEbf3hGiD4xkfAjA8v+DDWKxIwbLopKaGuCjHrnlgYOywiKZtG3U4x
glIsEIPb8sknBg7JJ54SdHz3cq6sRxFblMxTZeDuMIVdgO89f8TGQHOi8u78
lTnHx/0+e6huFgaT8/eOiShxFwvT5woPlqYditk0HqD0Y8VwRv4A6lulkx1N
991ecJyunLc4GhutA25fggD3JH44aSwBZLD4MKHRTyCn2b0fLzxD6uG5CVBm
vg7udF2dy3neQ5hH4qAQh+puAR0AW6Yr4IvI/Byl3esWEUljDFdpWQbDgdmn
w0+QW3746jspZiLEFi1v54DgeCRhyqgnvvlJf+BQg05nEpe+EFJ0vx1PvDlm
k98GvAv+Hxcc+jseALhgN0wzZITFaKAkQhApv+JPoF3GWr4gjNEyvSwI86hT
F6VRpDT6ClHoGqNkoZHFHMvkrIyrmwFrlYYub7+HqUNkuAHg1lyj0m8BZh0+
NdiBGt6yLzM9L+yodNbPyRt7eEPeB8U3I1Mu9bWEWqAeLQWyylphQGAXgQ7K
yb7i+QMzrYbvGJVrQ+biac5Xoba7KoUDH2+97W5bHL48VKAPcan79oyH2KNv
4UteanxxDUOqXr3TYlTWr3N+ewW3GUYdLNFeB4rKpgDUBbEyMlq48+CGcrwG
4ZuVrz1oSY464u/BLTd3VIPPUzchkK7NuEyqUaFqKYp0gh04SvIhfDv05jvQ
Up1g9/7Y8N1J6MmkCxHf563sTgaJ267hI1sA9hv0h4rdaz4zaMVtKIc+Fo4o
1U0C21idVXvoHZR9aDUioLRgaYrhZ1lhGSUQiOQQsZ0MGFQ4uCwx10IEqo/s
lblT1tdfj60q7+kH6BQ919OeEJUIHQ0jPzuu3l7ynczcmPCNWCV/CPAyLg5a
0CVpPZ57XVHIAzAq/sn1kOEEc8vdJ6azPcIPZpXUpNDiR0DeEOcY6zRhXMMX
brJSnbZ6KbZM0FuRsCHCvsteHbhNhzFBt9Tm+uL4muRl69itCFQduIB2gP7Y
EmveINTfCalfO50u2W7CsznXFvdoJKGuBEtJas3PD6dnBB9XdcqWfgnCzfyj
P0sk6xRPX1dotIXsU5UQQfY6Zrhb25fKGRemU8FoNoqinlu9T0M49sppRSM7
udMFeMMg+89/mJAnVOlwVJC4IfjbvcNhmdgz3fAPFAYfoDtct1h3LQZ1bBIU
frYdq6gUqC3Ei4THxuuvtSXP72OkojzushL/ssFtX9Rv2WSHYUGjnt4ZSAQC
hrZ6WX2EL+SpIy4uklA0MYIW8OQSl1wdXJA6Qlm8+07I+UwC+NDMLdpUBEfJ
bkk5rTT/IvVew0aFdtLF7zZq/xicf2fba8OeyN2KY311dQt6qvaMHJgd0QWp
Wu2UpPi93zeyWRsLYTuWI88EcUBOF4kfalmixwc/sY07oFUKo4Wh0afow4Zv
lVq5lJl4bFZUiDMtMKYyQc0j3kv+c1VYN/04O5KTC40RWJQ6ewFf03ddFqhu
oNPwMXF+badsFYZOkuFa8tFifmvCJTuXI8AX1hGTb7l/yrOFQxpyyeRB0MAL
MgIKNPfxXJe4jNOKObBtvxuVB4W468YdJJZEIgx5Zmm9okq2KMqa7zQ1eGRk
aujHXn19ZwVRHk1UuoWBAsMTwRaTDQD5UlrR48yik/wZ+yuNTMESVHt1Q16o
vxNG3VO+FaExpkfZpjmTDwvwjp9rctML3JrhUPtDTnOPJxlRwPk3nKE1N8iF
KvWNm88F2yCfNbUx+BrLdTe8uHlRz/MOy4hsvte9KpnUDDHWKBuc5kZLPG2p
tcEwVieeHEvJGHhsnGWUpzqlelmA1MbmhFH+aNQPwJL40r/qvzxMSf4Sgvvd
TzwPCuvSkkzWvL6Btm5NRI92TsnVTcs4iCKG1frX+leuqPjs4nPhIPYzPpHo
aqGsRezAiV8qaAqv7tCIgGEpC9tDP0WU1k51AfE9vL4v+5eng9tsmoCC46Y8
jWOmGEd2fOhXLXOnGVUmKyOME1xWVOgGPESk5UMNfcDT1XJHvtz5pvyqhzLu
DdlG6M8+t9zSlpAg/8ryYCWJz4EOWQoFFAQfj/g4MWcnWSqlJkJa17z9Iqac
5ZZsGFwJFt2q3cV8OXQghRM9XjT661rYRol6dnXnYut8WuL//+Xg9penrX0r
a2yX1e8Gft4OHiwMLianBude8cVXIAXGf1/aO5VLLYJ0F1YjgtR1qr2fGnIZ
G22k+YD/oC3RTXUeIOzARl8TDDE3hv8O7dJgP72WoXIOu7cOmDr5t9Uli5EP
Vpaw6bOJy3DFtuZFCpFk+7aJvFfgATqpwpE2pAv5FBNE74ZrNZSxHNpBMZif
pwdBMYxxNTsaq79g1w1OYqtQ8xTsikVDoGc0xye7kyhQU7Z7W13+3M3co91G
4fLQ5sdbzP9q5OzYPJX4kG0R6f3BBEKubBUiH/ZklXuwumtKoGFg23sGmGL0
Fyy21WEEBpRqeOP4aiDvIrIaYicJ27VYP3FiQIgW5fNzj7cnj/LJbAmaa56H
462XN3Yjrwarbmainr6tdKbm2abPihxPjNA1wgGlD/eArgKukIBkxUhBvOt4
WIl42Rpvyr3VH9pD8bEuVo4+exiuw6CboBwBsblfbUZLnkscRmqXMeKSVUED
c8/AvhZx//322plLNlXX5Yg0EbbYTfa514DDjCwNSzrXCdtWwPZ/wb+UeYkH
vO+KW/P2enENE7N32m02BkxxoS6QuYY2Zs2QF2HwEkrjZN3Kqi+1CprvB91N
WKCKyBPxnZDGGno/X1SwqQ7ds3UarNrh5UyIBPMupGwAf311o+HGSqZha9ag
GpACGpHhQV0uKVsPvb+OyCr2GXda+55B1PiBlAZCYptGjGFyjZEPtXgJ+OwD
PXFRDDqpN1Ia2MBd0WNK8pXmwUSogYy3r9nJPZX3zqYESTkzqDoz/ONkPTCG
wdQxg4vtw3t1THCUS4MFRonBaga3vknRjnuMelnsJwcwKMpiSmqxhh2zzhI9
FGF+v5ywnSLw/hYkpezlbZn6xkl9tZD8USHqg235SzyTPmfOaQwptahB/3UT
nmFlcEhVa8L3Tdf0Xhhum/eVZwfLuBZ2eDADOUVjusq9uY4pH0tQdJdCxrkD
Y2C5FLcl0yZR4W30Bpu3t4dA0eEUvZjRsZuRTCNP7M1FweytQElC3eE+1E5g
y6RLWhPTkS5vUA5chlyzG1MW/k7DEWhi3ZTsKRF2mAoduYMlAtqxr9sGz22V
6pcwLLxhaSFQaSB6f9eb/mLzTHwcZdcTZiNdOVCXC/XmDCQVE9E3TPCLn+1g
ZDRQyu7ji4V/uUwRPnIkfWkPmQ4FBGFO4jGd3ttgZeV807AFLBvp91F/qU6D
YvZKzSnv0HT8TVE01bvyoHwHye0IAZAQwcOnIXZ4dTEhUzaq2vttaiE8Vddw
TyyaPzf8BfqB67oRJDHaEWim+tYyNdv7CYnqmzPJiFLjlZAarNr6DKAm80LJ
4k1oU0ZaWZrx0VWSimF2JjoM0dUJIrzi5z2Av2+rTbZ4nAWMkHjO7sp8ER+C
YUZuuoEPTW1cir1cp29jNm/U+vcye0OpEvDlxxFsBoTZ8gJ/ftcPBHeOhAVr
kA08XGdEMFQtR9hACogDk4mJRtMqg3dBiHUvgQVDKb0VpC8u1+refQeDVAmQ
Ab6LfaDFDXJ/ye+nWaA9zmthEVDhDtmGXIXJOircxs8DaS90V6flLvo6ocgC
QTAC0VzJna9+YnSHTsQa09pSS3wVMiShoYLmOCxtys1t2e3N63yqUCZx71E2
QssjaArBHdmKijh5Vk3NiCpT/fgll253L1hStqvU/LL4qQT8OCklVTuHKlFN
Oa5RYTuvvnkwNOP3HEaD8DvdT340I4TkQTaZK3lqhdt8lTarzQJIKgm4H8dL
x4aeSo5cOWwyOjQ+zT8pnbtlOnAzJJ4jtTXUigdC8l3LHNDS7VhIpKx9Gzuh
1gYwuDJVcFj6vQGcRGP4fc1/ptHPaXpRjGUAO5c1kP6WHpSUaBW+6uAzslmm
4pPCENFaWTJF3kzOIWZE5f8JtoQprqWNouC7X4vsNxbI0CotMnXJiOk9xVg0
aekNzn9JFwJ1EijSJrYHjT4QGefVR4wMDYw4puH798ugmsquw0fv95lsVlh0
5gMof7Vznuw0e/UmdK3fsIaREhwaKe18V6PZcbTbjTplsck78YDpK0fnVr8n
Bgv4ltkbia/duy3ccehp+Xi5Zxaj5mwTCOhzyff/yQOsr61OHeW93N5x/VMF
2pfYT5EAjzwUaBY08vPIcuy3/WsDkVGIH6Kyz7PY4SfR5tWplH0AURtDXuP4
p3rAT2z6dJ7l12sEiY7jlXnVda9jh2PbT+PNPEmhiBKAALiElyfh2p4/ht4A
YdFuNFALZWdmh4ySx26Ccb/mM54iVHf7Xl7cnYxyj1v/LnRF+jwU6GcMUQQ5
8q+qa5JmXlbagAOwf8fz1hfDfKSsO+e9igbha7cQ+zatcjNny8MOnmnZ0bdn
V9U20m4/1Cm8pwT6IDAFJVWKZOfItNYGXSOJw3Q+n5lVPyEuMMhf2IBVPIUC
j6ZkpiR/4dCkWmpw5B/3Gy/+iarb5WUCd0xD7JSWCnQOene0mJIFpl66xp2E
oa0U9G5gDXxls4vPXwTnDKmQGSh3RtWrRa+c/87Jxjv2PZGwysiY0VjQLooQ
zxyEU80g8hTLpLBLhZfJA+bfoDRGiRan+9+ekUZit7kuSPF7cLBS7qZkEjks
1/K1i0oq4ddeBL7x8f20znuViJq8mYeNyJU06rpfG1Tq1STrXGmDLYsHpc/u
LF91+M727HOHLtWj6OLPhkdMOE8OxCnEo4QsGzujk1QIuIscSdPm8M6Vnz0F
cR2orCYkHMsB7UhscyEy5m1/d/V26kS/MyGTWpnUU58q1Frg3MhKPmNyeB9A
LHy1uPrk/VfiEfTlTvapzoLPpvZJp6kTNFY85CYzxyK6/YpkJW5Mm4G7r2J5
tJVIrY4EegdGm4XUQee0oIccQER+fNoY8KQCf90gLTwmK7F225ZVgtro4fh1
YHsulL1raBAM98htPfP9t4aT4xA+kvlWpN492GhOPgHlCLoqDOcJFQ3WG/jo
Po92JG0DhAMWn1fBc5+pzesioZoJpBgctLwYSQ0Bj2uF8R5OvGdT6+y2pVHk
tzjv+9l6yPSEyHGknPDlHIVljUgIuGjKqHask+EJov9dmaBILqiqqjAoD5ej
UzKWyJz4LLGyyWJEHS1FCJnOClf2j1qfW6ZLk6p9jjib1XeIxCiVClrzmwGO
fMgtw9OtvO5qN7FnjjkHjioc9kW2hDYviJucrQ9+HmBd4GHIvRb6igB2qWQj
8pwms+CP8SEeHZILQIJ1VRfd57paOJe990NB+maBmRGPu+/9PYLKwH8nSOK2
B/+Fp/a7oF6espQbbKmxSrplx4ahtq8wouVFnzoInP0wiMkSwzg1bXBT+UVG
rHv5mFDabLjn40QVbS4Uakp7CcyvDLHXpg2hy0MlVXAXBaFi5pntBuaV+9AT
oaNgrn/Le725f8pjS8VX8jEV6H6kpMqlsrdBI/zxJxsG5HtWRgRyZJssNgK4
tY9IOttLNeyiVQ8SsMORlA/2yZiD+VCDK56pH9UNazuwJvKOhwGN21Biakb4
WWrO/DFuKB1RHU6x261vBL0pB0in6+MLEQ+iNxews96xPaHUjSEMHWzB/6pd
ZosbFCfnxi2i2Q0QQXxUwKq03j9V5U/H1FqxXNQGi0CiRugBdVdtxIe+BPlN
IQqNAQABzPWhM1z+P7Or7XjQ0llvWfplj+qr9WMUeylVPfjf2LecBcaVIbBH
TdHo75m6tKJjutR/34SMI0pmZGyQs/AzhZa0b4WDeLr+5wh3UrvMH37H/8Vp
2iJhGCTyfmBspJtIiKMKiRXMQmsQ1fizHD9uljPaqv2Gc2tAG45KzBVIB+LU
Xm5wlD6xvHSZHKjLsc5HY+HvA6F5HQl9vaa5l9lc5Eb9AjRaqLZ2LSKLEYEz
JYPQ5NDuwsOdBCDoTcyT0gbo0WxswIPgw4DMRHfK22ukpHb95GSM9qWrg0Fb
8qcwG4NRahwrk7KOfe5XGZ+E4a2y34CndY0uuO/lMFA0FmlM+6gUwWBskkBZ
WaN6216WN8fIUgd02qMI+zybSCBNqP+LQrCPZm/ZFlEycZGTG+mbO7PRk9gB
/DfgL2UJmK28HV0UVYrCHw7T+sWRugOhIH2Ruuz3upw5N1T4+80jxMRnOd87
lXkjyncn/+PATFdAYqghvcGWzfvVwxUb8X1ieoqs9bWovLOe8RiFMMzoxXJ3
Jo2xVl4a7Ttl95NS2onwbP9L1kvbTOJxQgE/2hQOjUlpKuTSWA/EqU0kDykx
BT08EJZ7shwQ5lz3v9TnlLhwNibtr+wW7FtASSZPhNiHY8HYk/MWQ748GNjz
wD7X0Ez+39OJfG5JNWkWPhZMRc7If74KU+wXS5RmQ1ZRQ43EQEfg+1xlxtlN
FCdpH1Lw/0FIUiaTtc9z/ZDStOP+54BsrK553UYrXgILWZ548/MxRhP+UUNv
F8j6cKmDW5RyGOLzUr3cfhSjlUGB9+X/k+yATV0B5wuFPSKMw/X0H8P5Sgui
xvqkwgUZVmGreRaxEnSJ176Ir2jd3BF/spTW1q6y359+gv2LyYJBSwM0DOZ7
ihq6dPtdDATQA61gj1y8KRTD1CdoyeBnjLZpIlQJSIBkBQ05GmmLv5+1ni/2
zsHTiFzAHVhgw9p8b3RYw85bUfgTupUvjxs3bVdWN79l/gQHKgDgbTx1ESOm
dBktXGBNVGmJDYsK4Rn/fd38e/js0rriOEqR8aFXPIwD36kPBgV6Gy3Bkr1S
mcvqZS1HYmhXTjpFOp27pOO5Ta5oOGcdaJ3WiIj0S5620bKOz0EYLwS0k6c/
Zhye0nbYwCwKHZ9P26xD//qgqS/FMOU5/479nilXcwoOGC1EVO7BlGt2lyFs
P+woqLlxXtg3+DubtWyKz5TI2DLcI3OMCBV+jMfBcm197O60ietaN3eKRuyy
QFtbozlDAPEAdgJrV5+UstA5PhESPAoff+5kJZJAbO5oPEC0pF2wXfeMlyC8
g+c8i8oHNFgGDu1REhxqsxy/XiUqgAhgqS5/8kklkquNVisxcBfv2CnUu6me
LhU8NmKBUdIhHhQS4wQEnGJQNALl3+SFLecvs1vNSG9I/Y/ht9Z5QKH0pfcb
w+DYvzm6UP1VsINmGxOer6+bKOBQkZmARSnf4TqAmiyLeDq5LpjEVpEL5V4D
D6u2KWiqwsTK/6YF4KiOGjQJygRjVZdlVtvrHtUq6gQTgJY/eVQ6rX4qkvaf
3vtVMiVay25cmIXMOI5IgYdxEQhHLzChoBh1Ymii5EoNr939qfD/O6qfFG97
lafXldKq44XV6dNXhToeJi8Zwapc+oHxBwlC1WQf0dDU8xwWPagPKtQp978a
es5OMEWFqGxZFBcb341qY9r4dj6lzf/2dGfAzwBh0mMZdEdcJFz/OCPbOFCj
9jNTk93uygUgSNgM3Q6IRd4b1A0FW4duVaifvJdT8Exc4ictplwXXzhdUZDf
Ozy9PaYZQlqO9LLny0O/JJ5maTEsK2UrWhg3EdPPFl6bI7rRVcCIXCCZrkFk
Jqc5auGFolufxtONQd9H9rhCd7YYYsojBDNZIuVcqr49VwDeGRUVbOW2YVhw
/mhLJ2aP8rkp1nnceq9MrI4rjGWTFHgbZSqSbfoX22yDPnUJLAjwwlVlUiZ2
ky9j4Kz105Yq+eGh2ungWlED7TUr8i/r13KCXNwVGFtSzo5JyZE5IlDlvtTw
Pm3jFI5w4BahzQYUrB9JtgawQ83YFg+0onz/fQfE4Sw1EO0/unz59oqAEpQT
sTe4ybe1T0OCFiijdYRmLnoSCRWuZkPMF+s7qc/pF7N7aSKn0s10td+V1FQi
l4oqpKpfkBYOYnM7IE0Adh76pGAQalJgXW+F7zmA7qUMcOVrxnSFQv5W8dHA
h1QXfKqkPD/Rs3eqBUZXccXHQ5zJq0LrJB1mG347kauuVBmiXF2wP2nvrrVF
ZZPIUrywMNzqcCWn6W4B0YkKQUxCKTaYen5tnvoA+Nr8ewlsvIs/kvzjazC4
f+NijsA0j+/yp/iqh7vy/lv9b6387iWTfIye1V5tJLx41zGLcPWvutuoEILZ
0GMxIVbskwUAj/E+XgQrWjyW6vy396dRDa4UrC8M+tpMMojUUFa+QLZr6gMg
MExVeRuTE3YGaIK1fslQ82pUBeLHXyJ3SMpFTwfvXDrEahXzIz3kk+4lNvO9
v+yB2jS+A/XfsOMvTF5cRnjNhRCsMjDMWAkXPIunjI/M0SflOat4Yq+4L7ff
cALYsNSqr1YbPyz7I9kOtslAMTCYdk9sy9d/WYq4nuzVAoHD1vkfSxSujGBu
KD8dIb/OC4d7FRBgCXfPl+OByGQaCrlfaRNyaUJDeDzqMXxU/aw3PsdVqZUR
nPxDaAqb9Cjn7Ur3DyrRbRHzgyRmQB/mgy4TRSVDpA5mSPGYlJuRBmVrFtX/
9DpdjlX1shgP5y3rFEkcZCuxXJbR/oENr6m0Hp/Vo1LjySN88yjduTknsVmH
6vJrLK9GNjqF3bR6LwCsfPy9+bNXXABabPpq0VMoXmwl4r1KysdzN6bcNwfz
MJ55ywCB6ek0i6+ISnA/CM2Tqb3QWVaYEwKHr7Lf/Y0U/mcQqUkqsaq3tt70
IwbNNiO2VlgAWGkhqvz/4UsO8gEEZ8xB0XHdoOpfv9Qo99A3ofopx7zNCU5r
UL3GF672+KhntFG5B/XhXxgXoybohmNf9qfXPiWuQ99ZY3rqTp1DJN2o6jhm
yFxCG36ifMz6EebhJ8duQ7CJZ5YCj9xrM37P9eYDRQXuqkf6wyjnjsPFDSSX
M4GGIU99i+qmK+Eq6sDH5UPhHVbgJNjpm5R9yNK24a16UsrXI17qR8tlbic1
SOFkH0X9SilPIQoOGWxY397oTXBdS/+3dgkMO0jgLNCMNEoZJrMJepcKcWq7
NSgsOhpX7nb+Ru6bRohSPp+VYtOiG4spqoszJ3m1/XbRF9medGwD+CAYRmcK
8dj506tAmboR6QRg1RJiHMS7h/wDZv5D3F7t3khKJZQ8Yg6Ra60loSRvWzSu
v54+xjyybgBkb0dGFosCUgvqP395Ec1VaFvHEAP2wmAJ95HQSeuYc1PbgtEo
wH4bhpkiJLi9Aqvv4AaXlCK5Be0VXPBBEwjTkJFwV/Q93a91iUe5BsK3lxdN
xqu8iS25A2br4gASEFyluSUB931fc/W6+Y8cGBRcVCV8EPCiSaSNDa5d/6hd
IZT1e2B8laChY06Lj+p0QmHFXm6ThL9mXCT0SpxEpI7QqH6BAwPoIzWaA7Zq
g9Vd44sStE0PLfplWJZQSuWO9dtTx1WmM7OmyDdDXdJKbrsgxJfHmfd3+1Wt
90RXdSj6eLkQsIX582ZMD4f5NcI5gH2lI03hHab/1kSmvDbLGu0o21somblP
JeX9bE0AsCnJnAinCGLP9He269irgcLCfTULigGpCSTDSv8ahq3ulOguBy98
a7BHwcQt5Nm1MR7OzqRtCvjhLlIX1PnXLGzxIC+hrLuRiUisXxWqahnPdpQY
VodhoMEz+UhsP9k7BTcFN3lzf5CUQWE+mRWb05tzcckP6OzbL4oKH+TY8Fq/
GCt21heQMM0hsjzE7cX0nnYvfMVmas8izSvfUi2HYvZFaPgv4N4erm4Unfkj
YKtRIamSmQSxGjlh4+52CnDnt1czo6FvCMJX5WVrhiMNgSW2bYpUPkeha2fX
lKC1XNKAjvEzuFMcIN/8E6GHX7VGDQiUr2CaPcpJtEIUpaMYg1PKO5fIUf3C
aGEmMQ3nDYjGE9fFqvSqkjaAHhh50hWTKGDvS3wtRborWux56SSF4xZ7QN3y
A8ZGsomkv/0ZLN3IzQ+Bs14FNuEiiJiEP8A6SvklqulcyBB0vk0OHuEi4q+b
FbHrIaOYY5fW/19r3j92uJ0aQ+fR77O/DsWTL3q5qOxNTIctufZS3LBKcMv2
TOvMDCo2zQFQ8FX20fOMtTfdKfLn4tc1ePRD+HnpFrcdk0nleOIrObXY4dti
Av88MiDFr8YlswC5Dma3nxmVVZdvz/RhzpW98uC6gRUQ3EMvbopcHd8QCklf
M27MfrMLioXQRVpiv2XaNk4YaYY5OPgoekLG60+h+B5TRHuk78dsMb2hSFMc
wFvXKvXVOfkQiGUXQ2UEhz17tF1R3MFrwsI+iQbFdwFMikfqIVVLfU9yx/o7
VSu7NGu4dsJ4TxsMrBfoRFP8jEkbVJ0m6Dwgk8EuGUTUxxo0X4SfRRlJSz9x
um0xRYzZmyEyY7L4Qqyuf1kKq9SAOvNX8RdU36lY2mr8vOrxyZZ2fkdYzdKh
3d1Y/vsJBinFHJB7mYGHBAjqZs1RWcUEVzJl1KrEkAvzOqQPGH9EYgUJQun1
Bhrlm5H9H5e1dB+ePtQ5LCi7ZbheIxjm2vfHhkQ2+Mt6+D6n6sbVft1Mh6co
CihAzNEvcqfUCID1zVwqzxS9OEG8FW+/rrNmbFGYx6t6bw8wEzahNDRR8SYm
nPyM4Xj6Et+x2ZMjiPP1TQ7r0Fv5vSlO0VeWQRvroetRJesyzTxTs6b7IJ8J
H37zr8VICsnHZjSZU9o9BmrwplL9JXLTTDCWah9ogvOID5nD2n3Ejn/57SFH
m710+6S0rA+PrzdiZmN2jH/3CM0ET23JgGzD00QYV/JNZNM9UilOY54+iid/
kWE6uh7jYq8A7ljBnk4rMn5uImWeMaJzscvZu0V7Hj4uhhqVteHp7S1ueG1r
IOdQJHrb3+zNcfQtCNrsFVJPyP0shHofBsGPI+D+igt3FegNqRJZDG/1n2I1
BO94W1bk8e15b7gaxOyJrO/sQljTqgaCA4W4dwqaYPWfWTRjPFrpIMs8/CK/
XWqDsiYcrrjkNdmWQJIb3ZWGtC3JBO8gsuZMIIcf/aKgPTpyYIOHhoaZkXTt
tJS87z7jpupMGQSrwttr5K0vSAN2ZQ1m9Mgcy+zc7mnQKYkRMvHN7TjueERH
/5MsNMxY/ioU+gj3FXUDEOjvRsX95QSR+NgGimRUSd0sXjINVEsqo1wWMJku
5F/1KHAyx6VjsXqO7dzhFzVmqayl8NpdOOysQ61o0Ma/sK5UrqlJAYnnACFo
tmchgAmVurEcUw0RbByQpW+mTij3NvKgcRtPHgX+XgZupRJ790x4kFbdaQ75
WbhA1kt7WuXEXDLBHGRmeX1TyLMBlwRTGW3T2N02RfstmFXrWq0hOnr509ZF
ofHUojOANn97HugF4BsI7VHF4EHAUfOTtEvhLYUpAk4oMSeUm4aE16P37UtK
MRD2fsn7Qk6jIY8U+SDc2eCUkELQp3pUf4ojNcmOuR/Y1UMhPHmR//mq27bv
eApUOg6se0Bd+tNwH7kOex3PlQJUg2f3L1AhF2EX2eYwUCfPExFgFBI58hjQ
SNe4reUdK+/ls6mHxvb3F6g8jFmBvrBs+xiq7iEIIkwdHbsErq1J9Kru1ZYK
Ov3ILPJxM4GMP/gYa06eB7MvQ0OQ1Di9tUx65rJosbeEd8AwXGquROgr3P5F
1ZXHpx6krgZgV0yhhOpp7v8j6zs6ORO0Ot7ZxXRWTtSwodWegBSV3CcxuYme
8QF6iNoqaWXhf/BHu1ULP3vVo8CbI/V4Ex8rwosi2Baf5uoQQgdTcqCiZip+
7TI95goZy8HWlp4J9XzMkZ3NcvsqNJrz7IvZ5NXPe+yXkAv6Ua2/znnVTdNY
+lw6+G9r1tm+IxVo2rAxAtGqn613K4uz4RxiAamqIeaCf0AJTvxTSXbJwWkE
dYLDENJniw5lylT9novs+7unx8uyKwdq/sPsOF9fDT2qUFULZIl+FrMjc69Y
pcWOFXdvOF2MrauwuQ8QtpXNHNs6jNokiecT7JbM0Lof8tDlgc+ztYifZZn6
gebPZApRaIqMwVK2HiTM+47FK82IhT1bprsbq6CA/trbrv9CGkQ4WsEQKieM
jt3RgLORs2WEeB/Ta2ljgua+bro+SmggERndMI/xlF3yARgwfmzWzxUw8Srx
Jf3odgpFDsC67vyqv99+alO1rPLCnf788p0WbyLBtxtC9n+9uBO7SjUme4h1
iLqnyuBBc4vZbyYRPnn3m/9xHNKNJ1zFbCSuc2GNehHrjOdL0IOK++rIMoFA
XWDyM8flBT7tqeazpIe1o9Ecb4v8Pi5j0XhpYZzi66LxP9W2vk5p1TA3mpIz
WPnUQKSdFPGobTVqzCIxWwMrAwL/A07KX/wIChr28Nj/RPw/zj6FrRn8YtA5
riz8l3jNnex9rHStfwJrJPtaRmfTmYxbWb1cZAg7ySIqYk4Wvuy3/U+ZfvmR
UuoQc/TQ+PjaGLHUrm5vXuFXgVpygjz2cxxuEbMjOjn/sVBr1OnYsRkWWMZr
B4jr9NbIJRMJa2xZnUbeKTdY7tX3rsgcNcNj+Xw0LyNNUMrwX4+n0dr3uVhj
Bdbsxww6pOsnBKBJjVkXgXyI//+7R8joYjgeZpTb6b9sAw9BGv3CN+VLG7eQ
4UjTkGPdJzEI907cxng8gj5bts8AEO1z25xAB/EYGIQE2xC2Di63OkyV4wx4
BG1Su3Sk7OvGKJDG3lVkVOdJ+wrXv0VWAgfso64cRE4zAyaDO5gFFTpA4ioV
QGBemKgtSQhDsKk1/h5ShhRbB3UU2ddJrONG4bCiN/pmnIjI2za3S7RiucXc
tc/8y4Ily0YJ7pVur3TU34vpT3ARHdY+2LcsmFd0ddVuPbihfD5G/OHrAg6b
fVwmvV/YX4ACKDUo+6ITiru3c0kd4X7wtyt9QT/A5Lf169QhVddHNTLgITj6
dUdRLNAUwj+ZB7KE2Vbz4B3FhyI80MXOa6HpSgLOQBRz77728inHIfugop7b
kSA+hmEtxBcOA5JQfMrdJy1uOwlwMJHghExCN4lMLid0FshYpbncerOln/EE
ORDZkbQFOiQcUFehbejhcIl8fneLJ8nka3vsM3hagptf6RwSXy3e3274VU5M
aaCjxRlaYIW7Astm6Xcv2nLWOuZOfYCSmwVFusN+Y80EFlOslEJox4End6AG
xPtE3LB/QkvITD6GtfJAFvBbKCAFipvaxjRZePBNLJ+uIjH1FI3Aays7RTCt
ONKZ/T8Mh0y3F2XDP+ZPXbnHReeGY03NYL0c/DkqruIVb0qjTUUKdRtFh7ez
Cln9zlCZARmFNClijx8cbVNZmePKSPupYZUGQzKVPXna3slTM307tTwwIvOn
HdiWkqBmS2pgkb6BwCU3qX5TGD1eM0BiRXJ8539pIfc0k98POpXngnousEqW
dLWO2acwsdRFVhFq4V2qn5dGTaPKkpLlnG2h1qfKjiZbFll0lKucsZHBJz4x
23VhUm8wHj7El1iaMCBtmjKRoGoRTHTm8t1lkBqbto1pp7CJpgOY6jUdex/X
vLR+0D72OArBPp9hHNUe2T+fJD/NFfjfNiwoGr+Ytoc0ehB7tn/YuuAhgIxc
UA8+/i6VPMmUdgNV5fFVuOBXhePURFhCk2tNIJOjyyT5obj1f7Hyo3l6f58l
Ju5tVF6CF+itGEZIo+lqCBY7HPV7D8JrHInzDhgLqyBQHv/7b1KfL6iDnXCY
JhEXMdSVrPbBym83Pjg/xA0x+sjTr57wCsr6vam4q21Zac7K6yN4tK3ajMQF
iy5TRK//99knLDiX86r4EVVlvxNTNhYoYTMcvQ85tBl2vyYmJwrU5JMULN3S
ryqugYN9QDicYet+jqK3IdmMqdFZIaD7ebm88sjpPIrBVMHTvRwVVtnb1VNN
VNTWVO9qFPpEUy2d3M3ScrCS+/QeIMsWVbQCv40Yfev/Uc9AUEweugk2+q7V
Gnzgi3LGm+xqWTxH6IUZH9Lple0QrXUGSd4q0VDbCITgEHMuHawAZ1i06hSx
9MRWQrIW3CFI5MyiYuiLZVK/7MBl2/lxLCrhNQQAfpBpmRyl37+GSW1NXsTF
ZZayk/pDm7h9UDN9tr7Uhyqi+R+IlU9Gyni2p8sVHY67zjudxDZd8vlARkqi
etPNe9Vs2hL/k3VXJiKaEwIunPlG3HnU3bc/HpM6fP8UG2zNktfYTvt+6dTA
bz8pNMf9b8nQPsbfQos37wYmNQQA+e9esFXtkdkgrcmrKHrOlNVKaeuaAE2/
DwLOG5JkN3PyYbb9xIh+5vhDEBIuQK+7R2QwlFRMfsXNbZbU7JpgJ1vUNMwb
+e1o2LTKLpB+hB/M+q/0htdDHSmpXFCIiN6XXkyx498IkEh5Y5hnYsA8EZrG
00GlrrE5or78FlhxiTskCDmxa6VJKAMCSFPaUwSS3eG6+mn32PTlM2FBAYGm
VFC0H5QlgAzl635O6R563unwAJXm/UK6MhoMNdF08/5XgmscWAZ+mlQpEDk6
aPJDANjwL4MvwfpJfvuxHJgPY070shBOwcW2HiCxksWcyR69jPnWjf9/rLOL
2Zt0+tV54wrl50le8zv9tVytVHz2/0VGxaCMvxgj+ntDo//UwcExpEMuQXgk
mEIJxZ5mq16ctxIUn/Pv1dOsEcsAtHAsev/UgFMRilSr9hoK/vldXF8I0vt9
hO6zCy04uKRpzW9DdnHlFuuOWxcQ2sIKoPpVTGP/QRyDXwEZtG1H6MgW/Pz4
SAJJGgacrJUbYlFaIm3cvQVIlEGzXle0U5njlNenJ2UYVMar49qsSoGqGWWJ
PbBVYp0bQw+/n7tcNCFJkzOGmkGbUx8dqI+LUmtY5vu03AAcBMLehjG0JEEC
Y3P/NIpF10DZU/wQiYhb450s0+c19Gw2vSL/2Df7krQYYzJHRMFtApWVb9kH
0vTz1S96N+d7JIdJp8V1jR+1p5tzKFGDp4IZJF0DzoYHopY3pIgjnB6M5NAa
cLVTEGqqAsK13PB7kUdu2rn4X9DxUu83E3DrhNwkrE188StxpPN7Qs28RL1J
3AavucPzHwW+30C7A74I6VccJsAkdjaG1UWgiWvKdMTp+tytiyvKNk+0ffHt
hILQnpGHAE4+q6OwYDDGpL7N65+NpHLp3BHtXV9lSH8qChWgNuJxPDmuGmKi
PYAzTje8R9vZg/CM1J38B7Nr1bSkHEKH+8B+GMzIcq+1OeB1ttFLMBb0mOTq
RiB363RlfBQo1oTHJeS/UcykmveB3DTXqAn5YhwgR0BzMrPN2Uaf7QHa0Esi
B7MStBoCO45T7AuCwmAkNla6ThPdKdeO0PE5fcqJblTwx20vIWezgfLy5fcX
TGLgbHP+w18hy1HAccOITefMRczS1IuIwGYC0p0CUVNSyQLd+VeVEBSGKhR6
osLbOnH8NaLscg3dwp0Fc255fTKTXKCb5UcCsPYwlkj/fKMPfFsi/zMzNh8Q
4Zsw1b1NLGhU2Ele+InnEFbQt/5h7E2lQtEZ2DnoN6uigKqNNK7UF1q6St1d
zQEKCueC2Ov97vW5vqXwtG/C3Xz7saWwqP8I7IOhojlOUjwQAbj6kB+pepSC
FK5F3ZjoOJlMgjEt8S5sncv51iHkpALYL1lRdJtFyVTqkid/DRphnzfismfc
WGwxuZ5U1HVw7SpcJNj5i8TZsdgo+fZ54w1vF7HY8lJZl80NQ9oeMWLOhNA7
nL6/1X+0g0Izr0slBNTMEUqMfn8SaDbC/pnIt2XCg55CETdV1Bn2gCigtfna
Q+00wmsp2jKDTIYKYHNQMWi38bRi6c9MyUr/yPvT8tuLZpiIpAt9QI82/Hwx
N4Pij6RAYiGVitmZuN7R5TEZz8thsM34/Ygo/nKZrAvDVeOEfkIa+YPlVu3k
RuKsB6/UfhBaOZNfbcRTfhp5hfC2oAJQ4M7PZT6DMsCKtrQPyKLhLnnUr/0D
pNs9o/1eIU1j2aARLVhw25xMANKHedVLgFlUpW4JP4YBlBeWWfdk/Mh0NT6R
9x1yEUC+htC1ZsAhRWi5l0q/3ciVGg3+TASeJWrI6ioeaHO/y/gtUltgwqTX
1LlrE0s+6OEXbYQSREKuhyjAtfy6ASeT8djfSAe8DO5f1ETZMeFXleh53tFM
utEOslhoBqgK4PUYlji3z5ySJtKWhxTQOVE1WgzYJpskIkrSrL/a5MXv71C9
dC5EkzMzluehaBhVLwrlOiZYNN8O/TfnuM9MXzM6GntEfcF2osU4am0z+In0
5aCkxUjRWgvZKyeMt0teUQHidM0Z+xZRyW0o1S8ZW3+9lLiTxDxg3J2e75NE
WL/G+8jR99LpEV7cWg1c0cOKneYcvendZkvE33p2vpos+oP7gbZ273QZNHV9
HjODUlJyXg0+lqLdS61YJR3RdruiAWPMCLYgaVrF6lBmbxkER5lcxwOqJdrG
siyoXRtrp61dlEIt5IXsnbfRkSXlWl6UkHThYWI7cYMi+jm0VZru2GFa0Z8J
o7nMaueqb1U7cqbo82nwaD+q1U/g3WEtoHVksEkLYkmFmRJ/Mc95BBZv/Iwr
wd0yiNUy6NoRvVW5A6fhJPtMM8JxCG9aPOVmFlSwGlBhn8CySu7RJgaI+Ehp
LSsyf8nr4imOrS7GgZZVTcXgaj/uc/eMRd0bulvGKAETov/ZPf3oxb1u7l3R
3VY4OXgwARapiSJ8LtEIVqxaCiSvISlWc6FPfEyQcJRQxuoxfIF6rGcMyihV
OXuQNsWbnECWEXYxCaxgebjPQIruxBpbrEy0O6sfLgAVZgaqQMOdqCNG8tCx
JhLnOA/1e+TWOIWH75WnvuvKgHaSCnQXSeF+OyW/BCvSiCW+omzjKzVccUMP
5Jb7YsVEMqY+Q14C/jxx6VypWVjbDv8elOSRtN+YpoPLQHSTBIoC96pZ8ibp
28QTAsCnjdfW4PGzuLLf0TdUVDv/ccH742DL6W0/p6ckf/9wPeUw/jv6VWw5
TsE8lRH+jWf6/j0nDGSihvY2jEzOhY4ZlRY67SD9W3XFHuMfL1/rz7WZwagM
mLAtgtM4Rx+mBrrrV04QD6yik7aTVtQizVSB1p9tkBMOvLEb1K0uXvWBfVxc
N4hmAjwukR5NgQyBtBSsjutwidxqvRawnLJvrBPQH4hZvbiFdHuTAmaq+q+/
c0Mr9dt46+4hb5jw8GV85hbNnCPFiW8JwfYGUddaPT+OL0Oewgn3bhc+D5br
aVBp0pHB+K16AYH6UPkFktICVjbsDs6LyykpAhqXl/IMvlNes3ovsXZ6Uw6e
9IEbqdfVe9AeNFL+MlqQbHeiID/ThGeBKVQCRFE3ykk+Y+Kc6QumcXXI1/hf
uSi6X1NZQBLMzU6ovrRF8sn5YZVzc7QSbTQYhlRDSNopHjibGPsL2KenQdNS
OJU1r8y7eLDxG/57Dh69lN2D6CDNbkRmVWUbiGN1SM4TTPP0tJQx2acaTYnP
6GJjzKdJ1oNNv3fludPJZRnneM+Tuht4rOsWeLp10UwbIhlHwtsoOj+Bl3gq
8MlQn8GXrVDhhJsVYfXtfXC6nEUZGcE4G63/ALAbIDUMmpr/F2OpojLCMvdT
Ue6j/sCB21X1mgWJQPwDL4wZ+7dSFPY2VAKQtFVVPgKl2as4pZx8em8v1/H0
ySdno6MFVUP/z9ljYwRXi/p+HznkIoocVufBOFeatixVeXJ+ZJfGaPeBneHu
DAf1aBK5TBNf6OaopQ4npeyRybpT2/haQJD4RFxcXofmxsPZbCuYUiC1mEgW
MtcVlb6iHESvfiCxikyc1Wd4PhTT/XnLmUDG+VyAieqNVr3FgEvCUY3PGk9o
nsPDb1Gm1KIj9OooAKv20F2eeQo3fmLrobqoc20W7g7tu2ZAxvoVOvYjuQ1R
w+sEdUel0bek07tCdOhCb9e2bdmRmF/eSSXzvHYJnhE3+2REpgsj1yHjlWy8
bsPZw421Z+HLF9n6kmxPmfW6ULugI7owdWtebRUXSiOlU1yAdAbllre88Yfp
OxGnPmnT0FBm9GTZu36cYtYf8lD9Uezs26+wcmvafNOK8eNDxPTdhm9wkcUX
Esd7jV1XcjfEHJ+YgEyVYgE0D0zo5TtqYqAMwEpyVAoaqxoURA/x8hiWciwl
P+pZMKpxHnlcR5Nh96GIPpF04V/PPn/28R6ILt2fesmi7swJZErFUEV1rWq9
ZWqtbGLo56x3Lbd+4TpoyZnDz7kMwyjB6AQ+C5+Pns4UkNyS93Ey4A6CcBEX
dkzlcac5J0Lv60ew6qcruwNGu3RBmBrYQQ97ehwU4VWwxKjf+l8wGyIYlHDY
tRbgniij4aXrZdvm/HTNuRRvqQCVx0xvyGmllotpOwniCevH2myN6owN9zgU
gyhTfHbFEQw2lc1iNoRfT6cs0dp/jtBFpxFxMAQTChwk2pwf1tXoOf1xNg5E
nHyFFN50kySYi7MalyzQZnCWR8DwDnEg2prgtbmMdpHT2JqwNtSgMigpvwh3
sIizgLGsoieYOlFCFSxQsBulQOK7o32mUKMJ18CSwa+gSCeJbbgu+ma/os6o
A+QBi/O/MpvyeQvKGiLMIpg0p0wh9drOke9Fcd4lkw6sgkpjX7sIibKS3Zm7
2DMsLeX/X03F96psR1FABc/pVZwWZAYLJz5Fpql1Z7OMQkYCVA/R3NAK4xUk
yXK3ovrYjOn9cHkxVMYq829yiiK0AL55+3Agf8QmAZZdrIR0ynhGXzB4mzuy
ivApUbVidCNmHr24XFN2l8oXT9IiEa/STFTqJ/L5IIbBnPTfPbh19JD37FjX
HgKtA7JdWlwP2TLYJNNxZK3/iV0Iu7B6id1lMMaYbLY836e1cY7ujHVdf9lL
wuV8Dk55OcIpDqNB9a0afBovlj32xaBhmRytakvQdszcYiDg7DoKxbjjEPCt
Jt8npthoyVOnnoKegTXWI86OAW5EnJzCHb4q250DOiB5PJ7n4Eb1iEMWk3Yw
85VtQmhN4JMAdDgKAwPmKmB4C3L5rX4BHpGHPIIoHxpl4cWSqUTlyKF9ueOf
w/7CjNb96FxY7s3YAm4BYDSfRnXJ3j4jiCH2hkPigWMufkCBcdwyACSz2ET1
F9y4GJQvBIU8Is68sQWDw6FypQ7uswyUhfSspadhGMTKt4rbvA3NY90vregb
y3fKnW5DutdQBbSjU32cAtpMX3h0MqC/UBb+qVHV3ZnVx13e1eA5etF844xR
ZUSKEhNC3aZ3J9dZeZGODYp1URIIzM2fpl2CG8WYIRNeaxEUfRd7rTmHIlxS
fuoIxP3tEJerr6K5YZZYQn9gtcgulG2wgckoEmxAf+K6O+k26/MEswjw6trk
Rc2Nn5VlLAG6R+KqaGvyhRcLyl91ZcIvoJFtH6LLlTvxk3A7Bcrmwx8cOJjh
uMHXNBzgs63sRe0wS5XKbCnvWcK0HroX5LttO9x2Py5iBDI0sZNuoY1NBAju
/PHFSRYWKVvDAZY+yjHfphOo3Qaw6X9gIX85dfjFN4UP3IDTqqSDlkfk1ZqC
gGXDsbDXUx5zh4Jk+1ZJTWshaNjexZmca6/5XGGNOarEeG4l4MVEDEVTzndM
/My3viKEyDztVqp/Ba/NkeO4Lgf4+8nbAjHQ5M66PM5eDal4q+POaFbxVpTz
/utHcPgmCgKIqC91gOPtAGI5I52ztK/ipcTEfGC5zatflY/LuVsbpPS+DX8c
ncbv9OoiIJLrrb113CgAjEJUn1EIMABrzIdt2yKF0Q34RH7X1eN5UqMU+P05
p4nCFJNgVsRP7L1qo3R+Z8TAsR+Ocr+pVRHRVI2f0VKKdxk4Y53xODZHB373
V5gfpmkT81F5vbVHA43xlc8sxQghlJnRYX9PJMQsJHe9rSUitpSUpv8b5SSF
Lb3t1Xx5s7O1qA40BGaAuUSG/BeRYXclCjAMWEIK8CzlheT4rG1gpspRx2LR
BQa6F+UfDAJq3GvHyRaeSrTmmD9l3u+638NmnazY2Jm76ypf2hKuduNTNwj9
xDDfM1AwQLK7tA8i81J50rsomcOf5qcJx+PkolVP0LR2PvgJjy+/9KXI7c8I
cyTRxN5/wMhAJBICFkh7w3OJ4kSn/R8bPHFGrY5DvwSwdWKZymzLfNXGbTti
Tjgs8aWY7sYQHmWUyGBETtjXaccIOT40KSdjj1YvCfeSyD72wpL2r01Vni9/
2ryb0TMnHn0jg9zFj5CVbRrjV65OAxoutA+v4qIJOqfyE5pHLIynKeXDcUw5
FVcjiRRIx03uKvbz41C5BvwirmvWl7cGg83hvLKmX0GgnUsC2ocel31OiXJH
etSu0hpTiaAD9BCPWbjmXyLcyED60mHOfnnz6DfBQ6mmoc8oFMaO+tFJllEC
EnBsFBCIhxZy6pRqy1SXJFegbISuqQbs7nKdwvO+aGzsz3NFRcs8TqpOx2ss
5hMrNZJ17RWqOQWKbNxCgDA9cAc7uLXPk4+teGHzzfULE+bGt9+PySwi/QoN
QwSmmmbTKMh+H86V8KxsHLKotwpHlbJTYs3GB8On4SPdOYb4vIl+2fIwkgKg
RH6Ax1k0E3luV7NVjvO7QZLjfF4KXCiqMwLAgyDv5VxJpyVYQnXwVvC+pw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Eqcy8tpFXKDnX54LqDwOTpEaeQag4lpXP/UEo4AkqljhqNqy8zuI3Kevxnw+6dBlQmXb21Mfzew/1Mq93CpEBnI3xLd5SNp1Q6pdoHwit7j0dmpFzZS3DA5PjXzJjfWteb7OYlQ1jKJAcL1fgfLYZx3Mv/1C0wev+1NemoIb80E+DkGLalv1j1c2GYHNj+jFu/EqzS4vapdObENki63qbhib05c6RHYGBX5MUVDr4Ofyugs2wivWoCdmWiLS4jW9P/XYk6Ly2gQK5L/kuLT09uXVL6aE/PQfRzF9G5lxKSHW0v16PFZI7jBbk/7M5g4RpMMJQF833ds7Tr/wZ0MDlaBhAC+Tg1x95NrfzxoGJxRZE8dqoXf0inm8B5/OQJ1X8GG2zr5nvGRAkOGshCpIK+jJw+kzmcBLS3N4TFNNXfXqQIcIQLt7Msh/k3I3gmdS4Fox0kcWctksTpxBQbhU93l/G20jNhlOuP8iVPbDtHTNalW6LdE1vtNY2lQ88mC397jxskL16Dy6jzV5hNYk6x2D+KUavawf8vHCciv4m3F1uHG9Z8pAw1CY4II4bM1vY5b8Cyzq0QMH3SDetgTJVHiS2qTBfzITumZ/AVqq0SfYIbFSWViWYz11tmVNvth7I27ZHgzRCRYte3QIboIrX9vhSRLwihJSd5lIaPMAE954SvG1LWt6z7rIh6zKnhJyDnPOjcSmdehh64BZcxopN3JobQmWNNg/wzpK+yOtzlCKn1YRD622N8BVE9aVJ8ZdIuUTHTlP0p0jd4VQoKbK2U8"
`endif