// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AHuvo6VvehUucBA8clUyAYyvU8sLHYwksqwZUdsQEIVqlDJQ/dlHjBe4wFJ3
pyTPmqQLTu5imEUQd/gUsUEzX9Gj/6pZNOx3zKgQM6dMAHvWByl5TZurMZ9X
NIxOc1TD8sXJPi1R8xN4d/G2zI9g8JvsNUdVu+SAb8LNTlKHy9yDPly7pjen
CoYCyb1oO3wDmmjcQJ/eaMriVfKa3noOIEpKtWtLg1VL6KlqdQDzdItxPu2H
++7iAuMNmca5ZAFghUTYKPpa5cAjVv+alEu2RaytrzS3z7LwH/a8Oxe1mSl0
hqek8C535czwebc+0R/7Nouudd5XRG79oMdr9MbysQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TQw0EWv8ahY+pXbjFuTlbkrRseYRWv3UuQEC7N6KM6XpDZwJ9QtzTHLNaIY9
l8m2KFKnqmDI1fvLmRwNUgYnGBx/emprfKX8fvJkW/RVcMnQXiiWqiob2LpS
+4H0qTIEPe/4m4verFsYhftaEkM1FObnBsBXOOMqvK9cO+yJAyiNf96AzNEz
ZT6MW7h3CHHGgAw80ABNpCKVq1P19McIcCYu8morOnGhvx6eWsC+WHVKXkCQ
B6woaRWKIkupjRMHhusMbmS598fRpg9OIP0XWJMnmGYPJfcr26pQlJvfMpvG
id4beQEdwtP+rjMHBLzsLa3aaR7wNWKv7nbVhEIcYQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lM1l0O1Vn7K006HwhdMCztSYAuw29mpvxaiBtTAyCGAs3VIsmx6ao2+OOdYz
7GWkltb+rEHCbdpGzt2D1ncIQu/gWDa/nAgo81RABM5KCDkSPAIWEht/K+0D
gfXfcR6Hxfccl9by/IG7/Enm2O7jBrcC+8eEA7X37L/CnRekDl/7p+uhOpUd
+FqdqIdSODVXkZq2obNbCh/hRuMMltvjTeIFDIOUr67kXlzEDjHDnEBMdxlO
JIhXiGwgxxM9GwfWklXa3FNREN/UPoVf2PdxygHlXed5GZYL+znkSMdZ+d1w
syfbYZOSvxij87NIZPZor6JIw32coYuzIyUNQ9QODg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FcNLhlAXQnKgjkacZeN6awIPdB32Cc/aLdIuvAU6VNdsebu0U0z3Vzfvlbuy
YjDWP4baUIPhOjfc3r96bj9BvKXoXibBCiBAxzYuDA1gHTiSOgKik8mWYtcl
YKvaxu8286uqUmolVS1WJE5pteN7DggX6ETzVuhs4lRbJFLwHUrKRyvlr/OA
6Wtq8KDDeAMac4Ww90dmpoSKPvr5g/gnbJxH/oXk0oYjVTbcSluVEsmC2KNV
QS4/Nstt/6EMu8H89e0lbssnfppIVj05OVGOuDfSUghMph1yCVjis6nAfcuf
c4M39D9e/KePZlKR+Mvrhx6mQLVZgzXy/86wqdGXKw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kcTECizF3D/s4iGcyGqd+fPW1vJvGH79OYZxNEUkB4DWFZ5aFDWjdVdf/UZY
sNMuoXE5QVIY10CCZcERZMTVpdw67VFGFb6ApMRbKOksXLQxywlROtUBVW1c
4WyW8E1MjcdIYznAZoamKdX9Ly+VBaTU6sZdiWc/zyQfBc8Q+hA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
EnoaAd0ojCwP1cpZ+yx3QSKd5sYsqNBH/T8v70lnQxlddC3/YHMxr+mKXYAb
5usNiUzvzC3srbKqW/nAJvCFhSjiTB8oKV5UsOwvtEsRuP1o4DgUjd9LdiiE
ko2GaojlL5+fa3IM8ldwt9taxHNfT7sNmu/Lz1jbV9Fy9xXKyvOo7dS0dHqy
32Q3XVhpMTfe8+4wAyZAI0l2p+XofQ6M1KEOnKGZR5qyRofspqedmn3gpYUi
lhvwRi6VpdweYqJ5HDEnDffHOdMD6S2Tmn91GU5AwhSDVkug6mDWS73jB3I9
SeB/xXPtl6U9NoVU9BJP7/yrZEocBM849FueY7TWjQl3uaeQQETaXoKKovkk
7xIXlwTiy6v9GPiG7mKUG1yyGEHOQgKO49bAxUIiWY+Jo4u70tpDaK/Wsmqc
VU8TL7THykWxJpfuPQVsg7VmvV66odyfNJu5h+0bZasTrfgNF9GTax2liPIm
so4nL/OBevpyV/i/P87/+tdM10N4jwBw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tBH18Uib4lRygRg2izHaxrNT2m11eNYVyQDuGzbwkw6S4Dh9uVgzlBfKhQuB
bPkt10KlkDXsoaODaYp0WNW8/U0ZTYU4o3EqAkk+U3ZgaF0Dxxr+OmmPcDPw
oTzH19vr7usjXmwArCeHglnQvuhiVpmmUKm2+3WZN0b25iYcCA4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L/1TZC4/uc0b2Gk9yRiDvjlaSikSXe39D8xHtMHN9gNK6ldnSXxfQUjceQdU
cMFIZtaXdQgRycQMyOom6oN4dzd7/0W65uDRJx0cJRtRQ26JiFVtBuf8xH/M
fYFNawW2OEvUkdT7+N9HJZCmln687TxOlIazhWnwY8oFHrx3JeE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 17520)
`pragma protect data_block
Z0tPKGdfiGoNsRO6I2/fpPprD4q5C/5VRlbqMwVhWUw3xLL7T1ABKHdHLA4P
NJTkikr/uAoJBN4YVE2wnGglBf0hp2Lr2jfQiFn+d6pA2sf9QxoWk1A95Ow+
QA7rsV7DQM4qEeRrrR1UAH0nTHi5UlK4f+MfdXtrx91ZSXnPnYZYOPaJW7MA
Ocl7DI67X1Eybfd/DrdsRHKeb1P+pW+f0J3WL3VXW6KUYcwavtTbef99U6V9
SV7I+JL3attOzPRWqYWTbO1vdXdUr9AyiASuQB2+KL/6XRDkNH8jhgwx7Nb4
vQHdLCwO1/4N+ykepjPdOaCHDeP8AbLva8SFxuSRmATUmkFtFJw1lKUzmuRh
9Rxf+twPTMtwVKLCwjARFHhYkStnOw0ngbtw5QX5jvnW55GSmRlmh1dE/dXx
EcOOqmXN6YG1VNPmg6OgZTpA9PflSrXJ7O3N7qloD9aAkGi2dORVxCAVOAnf
DHbtn2RGD4gNPFGxqD3n8JTZBChQLBb3TRVi5ZPMFmO/+bf869PBqUiAWYc8
ROJy5HZOZwEcyn+T+rr7w/6dykQ7SryPPb26LkT/nYFCnWvBKoHJghqJhh1M
sIgwDMHKtSrHjZMKQEBtW8DqxYWdyoryWFUlCn2E4yw2OfQo1CKGPMxyQIXL
NnQiWS/BR+/LN8DT46Y3iAJ6y15oRNliiblOIYJkRNxJvgwRbNr1Lu1sKN+C
T3G8T6b35/IZgZUkso1OD2BGv6O7nUN2x7ukvAOHVAkBjs68C95sqtOwzNpR
V4ODtzleNQYBRTeQEynR/uR0iPI7dHTZpTt1cv2rwX0FsktYn0OIZvbEZyjv
rU44dKJG8m3Z6y2DYbkDvJJbOU450db7Cq7Bpqv6+EqPWYM9CUlvRmxEjPqG
egkMrtd8w7HFpVEhTiQ3P5NV0dxoF4IpuvOQGcgJGxo/kqm8GTVYAZb577of
g/Qr+tvzoclYIOPg2MuDcLUnkZ/nv1MbQeZpkr6vupE7+Cy83998+tBD9l7/
5Up9QWQnCkcfH075R9NkHMWdW/DM01zNZXVV63pFTPdRNDCHLlQXrwladWLC
pm4C5DcOJ6zdAGf3qcg7r8ospdk8S73VZ5R9/2vNJSLC+T7oKqpHDvnPjPhp
geWb6F9A5/zKtwUoXUQcVxuDmkZEcJ3ISDWRGnSzyOiWIULY6B5OjdxmsCLP
BZ3112qge6HBRfD74ss8pMEbHQ/DfSu/jYjg1KW8l9l5fTSMauCI56RebAkv
a3v78SL5gK0qUKB6tWrXPX8rKzuJT5DEOwdToyF8rhFu6uNyrWOGnjgeE1te
EQT6Mvi/GukBaezLIidTMDygNvc7mFnnhYx6+m6aVuY1Shd0NRyR3KsQP569
5sdrbF6KS8CPTvDIet4g0rR7SUrYGk9BjBPN2gyWqZpPfjIweIpwKtKDOMvG
gnVqXpMgJ+rpb/fp9RvqdmRUjwFskCHICWcUSFJUvcUZTJviEocsAeyUptjF
+YG5E0chGaUtCpSM3RMvr6hK2e3BwO+6HKs5cb//lYmr4kzJBjgE/+hj6aHy
+iQmzH6ShhjYSIfg5hxNmtjAGcTxwfk7Fi6z4Q/BzJ5dp5OpererwnXuu1bd
vaMA/H8DJsGT1FIrIz+k5EUKJq9wfcmDSjQGzFwAdeD9A0QLCC2DiloKfDao
G6EmeymNKu1tASDVBTdzKBqORrc3GWkBlBxoTxxWtcKzoTSbZpfD6or2WGti
0Cin9ZTOyF5vEcx70VCbSC50fRZI4l+GitZ3a5rkW1euY8ZQ1DTLglEkIt65
42E0wS+sl0urzTyM1DVXLIIK7S0xX1Pz/dGBdjPVydO3cBwqIDuD5hUcj3k0
xNL6tkgVMTeHo+wKKMO786y5BHOLUlqudf74dNu4X5Eci0eTeUJItXRof5yU
nJOhAc3bQ+L+f3QmMk0TXfLhjSiK7y+5+aqImTbjfshuOLOobc11CFUEI8KL
1ApqFKoiciABYcA27d30O7I5oKyGDaEi+9q3qfmkZjI7DdeLldT3Q2hx7EYp
xKnCu77nPTYqX2VifiGcD0dmPyiirinlUTwKujkBlsDYTHd7JRZ+IeBXkj/O
A0yKz7Rw8FDJPTPOxN+LW+S0SVJwJM+BzJCoMdIWyJtHNPGx8HQOoSgl5Ty0
QNSBFFiMgirTPdk9BvIO3pHYSDMn32Kv7O3XzBNzVXtsK9O34WpIVY43Vvne
uUUjBXwDuAT8E/QXcaASkO4ZB8K7DWDQANPKBsaiJ+RGpwO92KTylFMJX/pY
5Rnj1qUJwV4JRbAWAGiVxpC3fTNWPdCRKVLXKoJwblQb27fNEaHJnBGd+GrQ
octaaW4S7ea9oqOP8vVArLJVVOFwHboY73Ofyzl+synyD135RLa1UkYYisT8
w03HcIrJHkKBnf3L8vqO0/Ze9qKd8fKGCuzQUzn257FeBUhI1xsPkX8vMfXJ
cLtrA1jNMrhw8KhAah7jq48CXesJ/3Ug7PE6HGu1smIdPRL7CQOfZj8oTuUO
Q+piZnXHEMWBUU5YQ252RkiL7fZBK2d5TJZBTlDbvwcfsqQKrMGDooB4+TR4
oUEcWhHUwiVhISB0H5QUOJFIheIkNr36VcDf7jS2sNfK0Prh7zQCSR4uv8sN
lMTTtL2CXEFaQysegcRTlByVHBhgNI06EAn+TT5tILoVEg22RNJTF9/S0Rdu
Q6iMCEjmsRKcoPBIQ6fWspV1B24/THlzpdk7UjBoKF/Bti5sZvVMLahTfM+2
7M22gAj6uGgPwVhbtqkpyTV3S3trXadvO0RCTCYPrEKjeggVL0z9EeoN+FPv
bZowoiZUOCgYQdMo11GxGbuGO+U14QUt0F6STtnlVV1HQUIdG9eSFBPkDMhD
c/wO8UEmAdoScd5/tS1o7KAoJszigDv7PDqOrrSOZZdFTvmUWPaV+BIIvL8u
N0H7x4HXoAI27J18PKDT6+Aw6Bj8d+rAQI36CHdZraViDyqDKXPWVCZk6ElU
AVxBhRP8gM1VEPRWrWW92XnO9Ow3/BkEOtZtcz+EAZ1XDqPA2tr6/W1rbghb
AaaRkNRvLsHsm6hqHZyAfBI/oW/Xo23VXsuEoLpPI7JYoxVlKy7ACjLyMuHh
8p/xyJ5rUshtZO+Q4mM0GUtroVNZnh5XZYasyjNUfS9e1QVRByIYjJ9VkIsK
w/Td7CZ7D2e2Ho+sxRer73a0D0kTPGoimTOgywYUsUGuAAV+IGTqZ0WucBLr
iGqYl6nKJH9CCqMJvgrLpfVndvHTbk8r3jat/Hr/cELuYYTBnhiG76PStm82
ZZKr9tcEMf3Qo6iz/bsWfmKLMUIzerBwf63qWy+wi9YBgtOqzxK4/WdeMQqI
GPU9TZ/p8P/eXCtHsX42e8FSGqs8kwBrzzE/VPTMBXikfKTZ2DaF0SpQHqOH
61POhttsTOLCABTQ8u29P/uMe1KID5ge2nHSaMpeYcOiH6m1KennWAk5p4nm
H8KNbFj2zSpEarl2PW47RGLdlng4LXqneCnZhMLcIREpkiHRywluQTjlXDWv
mjgGWPDpT9euznggmQj7RhgxXnAg+uFqe5PS8KCt1qAPZqWiwLHDI9gnzZKu
1eBUMtADagLWTiWi6zDPACwhHVkxbYYmEinClHr1KEubWbGztxTLlZw97LGS
15Y8t7IJBARsjaPxT/N23RRiP1kStxcWQEBqbJhuThhu9T5uxoZnoREFkc2e
czpeUFZi4rPRUksFeLfEVyYmoph28bXtL5F8anJSbaBFNQyI4YUqL2KSXzB0
RtcWaUCUjvCYO52GcGzlAOWzCvDpwRveI3R6cU61bhH3KIr+sh0nfGleIO0c
eZdVrfwJpPkXQnmPAwA84SUo8z990XbCkJN4yuKSPgTCCzIcLPtBuPr/kq2+
tvmdKDnr4mDKtJrrghSx0BYVcCIZmdOoTa14Z7Lbtdqd6XeKOKKQc3gSvzu+
is47RRz+WIlycH5KQbk0y81OZ4teuUeTsaEuN1BA7tc4fKZs6KjxDLOGXYOH
WvgO81Gkzgx/uw+B+DOPOsAunuA3KMdD4XBVyQD2wSwbPRYy58OExRP0Jtsq
agrOEQ4Hf3Rw30IY76gzQTCAbebek08A9czJ+jmfWuCzrFf/8Cyi4vCeHMaT
tpUlZ0ixyF90FEi1IoUxwlNBmvSKe/mRwWPx1QSJkv+VrZuiLfkENlApq+rW
bMx7Cdsaos6OInXo3dru3GWc1xkhnXaHLNJd29vf58GIy689w2sSDTf0xsQd
dJ4x5rc5O4oia5d+6YEsQD65qMRKPOGM5spBfHUqb8pN50SrGx072FRJIbEE
/2qruMhdT37q/y7QZ73Tt2CY9Qip+rrSCN2xPI/k3gyGcCFt/khknP/BsdQu
5FUKok1t35AZUO5dZwAjn8LLE5f6qVnRkTYQ9sDrZF1IMLw/FILhFB+UnSWf
8RFmkDW9SM5PscDxR/o//CENNuEc+iL/9qh037g1+lMasgf+52p2sYdGizde
BZkWslCRhh7J0dWAytCEJJFHtQ1pPLwa1C/zThtw5XyodGGH3MFufSYHsLVg
E1FQxq+97ko+oWZGSXZUZebyhr2pKFcbdb7Pm41pDg+FdVldOwwDLkBOOR1K
bt7imRgLDQN6ImHgwDBrpPXm2/bWrdm3EzTnZwV42+7XkLN3jWi3kJzHANpH
o6AzcSLqN/FAQrX3cKAFo61SloO6dpb2oCCzwYF2mwRQE64CipZe4klG2jrV
8VlmgeP6fOvu7kB2C1V1tdrqp7ve43LNDlSHRwWTpVaAsin9hm++FPWRL+yF
ruRd+gstjFyWHLIfvSXrIP4Eberalhuovdp54wTcbQYy5G0aeS9Y3+YZCm7H
mJLCmQdbwH88apRBT2m7Rc+g0C498SsRagA7wPUEsYSd882WZTNPIfVeC6R1
RgIvQzDH+8jnT3IOjlupLiSw5JGlFKvKlZSzlILorRi/4DVYsLc8fZK3h6Rb
OJminxn/ELKKp6UH8yDMVvnPXibKUzAB6TxNhQtR3Uq+0wKKzuWTAiRpciaV
KDXpZaVuK29aXzT4oTJi7F1XxEq1EpQ6ibMDc1Blgyo14Gh1yoNr2JbrHV8u
XWNM5nHI2AoteJvkemZ1WoLGz4DjAz28roaTEkaC/chMlD57cnviTE6c6G8h
GnC1bzoCOW/MJlpw8AMPgnml1U+l6esLTylrvpoimlZAOF8Ngf/YWBuDnPhf
XX5jdy+FXoVdL/1B0d6I/hcNaiU/72vrMnXrEq73BbBJM64oTwfxOjpsn5Kv
/rU8v1ItNOS4V63yE73nA5OOI5kce31qEukSTyn5pHwq0oMSuHPRgStOPNhc
CtI7dT0QlY2uB1XO76YKTPsGiEHErrXZ2TLZ9na4lJmLwtvaL0sZYwjen1BM
9sJ4zR6gb8aJOp+BOePmwuUzyPUrmNCXak9yI3nquSRTidgSP8FR6ImC3c8D
7Kkg1EYBvT/qXRsFOyCxADRD0WBKWyYP7dIgKnQF3B6TG6MR81ykbzWhuhwo
3EhFyRZuHE08EITk2l+02uU8IsNFhbBfw8Ndn5rGTIaJLR8pQKXC70Ye6xa/
/m7i5RDh2dqQT615rynmioPIDCvqW+DIPV5SOIeGhj9xXNpiPMOLEEHllLN4
24gUDU8cGYvpV+QXySQqkjRdSud0L9IOIDqz2WHcAeTlsLDdRln9Z9gBtYZ4
vQWF2vE9Iu/HCrqb41RuAk4zII/z+xkAYbsvKojDmU9e2JGKtx2hgS+RI/2A
yQKhnLhSz4QIKfWiB0LXj+A3yJpPiC3B5JTIge0mhp23rPeVVs2yWzi/8tT+
+D1mQp7lQs6S6vBr99DRsk5Z0f90RZwz7ZzM2KTkXZZF+kpchQPmCom2IhDN
zUQsqbwmXNf8XM/1lxV/8KFmOzlJhCJ32I3AL8TADhD1pKf+Wowta6SqyYH8
HpEQO2zuH8D7qCLdMZnHiCrLbJ2Vlmwh/Q6lH7h1N3+NXpasWnB/SJtqhfSW
xGoc5Lg7lWaqbum4Mi7wB9RAAUE0e7nkEAD7mAXDqlnF37JlRX4ZGON8zpLA
f/ojwprWOTRGxfaa7HFPZ/TsS96c/qAy3sKDN+hVN/3NR8/KDbYwhDuhwhbi
deeYZZZm0ogEHgq6+VtCqCX1JYYRhmf7xX6DIBPFRwlpbXcpZwuxKCRz+f19
073PCgQ+AoUU/j/Bn1rXj7dRICvtM5wjfwBMcEflaz9P/s16tYwmFbZeg3U3
22cNfaEkGM0sKW2uP1juxZZezEKUCFvqTm045+TCYF3Bxezg+guuzfaGyMNv
RbpssLDLzc+tQbubsQj4uhDmJPRUXgtpz/tRG/f8vn4kTbrEkdAaEvocJxE4
I6Bq1k5x8dwcSQLiIHqdluRFWniBZ77OSjGcEjeNeIc9YHf5R4y+YpERWJgm
r3xKjW7sHHIZuAU3+AZifAR7CcMxlUXW0004Suzv7d+QX1Wo5j48dDUqW6WE
EduhlITAQXjanqB6Glw2nux1KMQOFiWGhK90CqecjehhpK89+zdO8WqwzTck
kTE+z6F5QMMgchvqFrcaGmUW8Xjuq+nw48y674yBmtu0Tk/nMuBZtaHGIjCI
fc3DnVdKNjaBg+TTu7gxcM4he2AsQx7HnJpkMyo1deLcg4BkCj8w9tLokBC+
1xd20vkAi3/2EZ05790stCIbC3BeFiCt886sEVj+1rdBs7x629S11Zi23zgf
Dfzx7wsH2WS8MjlGykq5XaUCmwUBnfZsAZMsp8UgBh4tWWjoZhYJzD1zyVa5
/xkye4yoxb4wQpi/4CIggyZKFv39Knd8nyVPVHEcBGdgSmCx7rjvSau9MlTv
+0uXb7IGuSMBM4QwhjIvGLvBtYZGzxbyQGOTBqHE6PNwf3taK+SakxrIWOkh
TkXTt4qyzkiBdY9a28+pQ2FaKQQuRt/DQtVLIafJuTM4GLWQUV2yaAser+0T
dd40OpOsYGZqJ0P5wlV1TqSdggJBsBT/M/6aHVv/B0xqN/zKSWyIOB88/zg8
IwLuE1S1grQjLsQ1nwejhGzn/UAT+msaZAMyYvyZDSnHCLmu5iAKU7XjTag1
eRGx1S6NrlB4LJJ11BVSu/qt/sGC733/soaUojVhL8kpNBVvsnN/OAPle57I
qi6rX1wUpi96YOlSDcwUkg6qkmSQUtZXmhbV5ifgH+ovkx/TGobmv/auarB5
4PZAoiXz/2WQ/jpNgK8hJdF3AuzHHlFEuDe1pl5PX+CACxz/UFFN3aBW/JjW
EQzwrLJO6WkSX+Qc6D20GzdFgncZs5aJWjup9KaCeKje0LJJfs7h6xSd4G7H
Fi2eZAQpWWSnuDhh/TW7kfg+k9dJ/pnTPgC9X7c2gw/CpXIrH2/m+aF93+/+
aLUAIAVtdqSyvVMOAynwXljelkENNOAgdSpSegIdUrDbGqp0G1hY7o16bXZf
VN/iuost8ZFQXeezvSfs4CKDYHIvux+8XjNflbZg8/VwQznT7hqOPdLn5/sX
hEjENRt6okdlAxYFrjqZOjjzpiywGKvyak/EMCxC9UTWwPKiU0ZPABOkmoQN
QF/3URgIAniuBQXuDhc7ScsVQJadhc9CIdxt/LxmiBp4wecBsm++B2qBHODv
W+/bRDilrod0ueE3KXFbN+RS2nT5U7h7szmTyHMzjstn59+sReRTM3e8rHw5
4W2xKsYAwh7jLZYwC0zfck8z9RrWEPOHnHi5ZVB95+Sm/hWGcSyDB6kt8GGU
xTgNXM0eddHAApQb4ZAsuhQkSzrNMbADoGCv8Ruk2d+BmbQishix66UwkZQr
26Ba/PaUJBy/pq5y3p4mm8VIpJUYGDhJTSrs34aqQ6Rm84in51B5pFgyi1gc
K7lMuI6UUcdOiM8gLsU4UfjJgckDA8wIEU4uiPI7ZuQUCyXUoSmygEOZoGTg
JZxm1nYdVfG5j5iukm6Enh7zWlKi58iECDSFikPXsNVdhk0sVpfLWUmnY1yE
9Q3TEbOf+RMk1iIjOOSWcBmSx/RdvA5xC++UOYomOmAA+5PBKOuWxzOnzpVI
vNSlDfqz/8v8254enR29+aeuUzXsNw1F335zBiqDqWP0rxfCvTZCXV7f3qqL
XC0kAvzLyOk0YFNXYlVsKNcgUnv+EM4SqtWQOHUyXTTuC8jHySSrTqX79VqL
ytCIYUQZrLs7SR81oyjgPTTpvBxBhVJmuQAtv+z8rnKAiMXDWRqsfvQydrfd
XaGmUFst3+ZHVU0CT+MHw5Bkh37rOETldr/kg4zGhUOIIcR8f+hLgF7nYtC4
T5Ufiux3Aa/07CqiD779QArN/MC8i8G/B+Ll5WSJ3GX5Tzf1a6/Jgvo5pB80
6Hs4tsFLQEXkkgNR3NKRG28cmsPze7mHJnnFlnhRTqJVsg8xM5prud4otJut
NqIhl02s5wKGHWNo5NfWvxVYDpfVMbqTfbzv/EwUs94zkz56h8X+VVrvdsDk
+BmF68IniUcbuK29ZP2u/peWS0lPZXwqC8eRLSEt9+fJIM/o84SehDu0jJY4
lqv71rQQAA1f0emAgF0xc0NZOdipOD+FvbTUfkH8j+K6+KwAoZxHd0kNzvhn
LwVOjH8clliPppFcuEyM5DXoL5zpLUb0zc0rIpOJs0aJIgOSGs2CN94xROk1
guqjFQJ8UjnlkXXvdWnbZfMAbHpsgQcOcB4m81pk84T6xLe1/83gd26VD4IG
/gC6/DS1C0AZgCxkD2rfC1eJj7FemAyCLfU+wzwsvcp4TYSBVjUrX4ZzPt6p
BX3ygQ71zIH06lXhMRk/ibs+VBgD5lRIaiiWdirXqUqbdmLF9cku05rnusn6
he8fQT5adzGmk1CAdA6yP/8Scpke0rZfgmcAOKc61ZCEBAsymhiLPFbAmuaA
z1wzGlJilcWvlupH+3b5yVbDVtWcLcz0r0atsnAbjJBd3HTF1v9AiEefQ28R
qxB1wC5ACIEHSmXTMRv9pj9u920ltzsLW7yAtuOjFYtq86Vjl0iLnQKofiOz
e8IHtI8TBCaKVczs4+zNu8vC2j2aLeTBJvTopwjDAZMoSLHYQxUeQBFySN8A
N1/UpLxOyn2uw67+Tpk9mLsnRzd74fEJWW2yAGwdN1rcNQ3RXSPXhi2ti7dl
+32kmZEP2xOhL/+Hq8NFa1QeKe66pCQuSISYpbi60dTRGtxW3Y9KgNufSCVW
6CbrRUYPb5WwDb//b1BvyijM3Jd5xTg6V9rUW0UCeLiqDXozBGWxnn9Hknil
RkHNtXP+YGUNWST/fNoEg8IR0HbHxg45nTMSlK/CyWzUxWkzKhmyaavsVR1z
go5N8IeURuYrZ6ARpsS6Y02c23ZpkgngwC91I4fCBvR9EgQ6VajfHSQcwrZW
3SVBHmVgyK/CXxqub77zcKNiwJRUVzU++NKIm02GIkpKlgoM+YWyATS9iuMy
m/DlJevP0Sti/k9xJ9HN+apaNIaPFZ+Zq9PFqDCgApiOGCgCQlTbT6RODoQ5
3W+1mdP4y0EUa8xuQzn0Itmo5Oosgaii3A87FnBgwMLfjF8vSHqIV8a0kd2Q
Fzz/ppXs3StnQCWVA7azXhfZhgtW/O+SgJQsfPsVzpT1r7Uf8KUNkeVhFMtS
VvG46T0R/0Nvog8D4UElayROiQfJiAuaxpUtoYuHPCM0AJimIc3dksZTBG+9
yaguHerzfxPxbRjnzkcm43LK5AFL4Fg/2W+LmoAzPQmz6tXs2f/R/93vmsIO
QjyAWP3K6xzMyztqzbnvH6NyWVD0sLAT8kemi/Wdyc0QLvJfcZURT6D5RILn
OrUdJYq4ItLNcSHDao7VxMC1e42jSgNpwt4HWOItFaLu4M+2SJc1ZjKz09W3
pPK+4ZOnqkpfkoQpUZcAAjxB0HayhZU03+t9wc/Au1qvNwhU++P553LEjiMs
DOVzY/mTFVEdo2X8winagwcu7+pnrJW9IlaLXr1patkYUlo/YFQGiF8lospP
JuIChVCyqsVWGdPR7N++Ew+5SfeHyNmi/FLFIrl3oGSJxr8tD1zZAvEk/SJ2
7Oh7OxQh0TRZBsDdKoP5GWQ+rSA7Vl0/iJGNAT8qb6tJE6IWHv1duZWoXxUX
guHQi9/3HzCbR0JDg/gBEG8iOponXJZfmgUDmSAVw4ymciRME48we2w/IC2L
j/VDKFGXdjCzYiuyCGMjBQWJiRhU+qYSF92hl0qBwiz89nTmk26a76Vs8i2k
UG0OeTIv/fgmI25BJv+nrl5Yw9zIDccbRInpb7HijnoQE5HipvKhNpEeOP+w
8XbKbA2VY+H5rQ5p7jK6gflOv6vbdCmO4+eRXTH8KMR7dWlTO9fY+JQGVsFJ
G1P9Tqk6bHJiDHbxp3dgbNH7z/ek7Yom5FPakXsBbufYB1xq4vMTmGrVC+6N
EzrKNhlhMoa11cRF4AKWmUgopR6wGJNPBYv5XXk2sd1okzAvXyG35iIyVaWc
zf8P1YM2Z8x+Ya+aESd2HV8xhuZZp4XcM0cUjqZxIxIariClbY8PGwIVJC9u
ZTmXeah7HHRRLcwkhCuLkE5KQfjJHJ9ur/absv+eyuTrzvxLhVFM1R8cCGRx
eXTrWDSt1P7OG1TTNlKtWvlEs9kzdNrCwDnRaMCNw2aVavy1PzjG/MYCAERv
NSMs7PDB94Dy8UP6C1H5Wdp/Yr2h+NNcqEjHphRLyCViyWVxt0k4107vjwq+
WtSGjM+TQOEXVi5AfpGj1MOftERHk6QnJ2fVSUtjx27LWViybMu0exB33kTk
N3uMXOxw8IYe2AKZl3D4YJvLyxJ9gATR765pBOr1RjXLwQ30ds8USmOAU5JN
CDnCQfq8cgrUfUky/eP3LrkhfXF0EP6Ra38JTcvYIpYNsBxrg7KX5Nqrp3eo
OikvSa/LvVihijUi5/I1w5K1I8KxJJVNWzmQGoGdQKuN9zDhp2rKQ86G2Ey8
V7h204J9s4F1SGXrY9m4e3utwkQ/UVE3YaIhieTNKrvyuILI0LxFHwlJkpTu
KBiZs84u3xIMyYsYq6ntIQBd8ZIljdjAKG2lFKF3m4sQgvVdZRF5UE6PzTnQ
zwFM2SfoEl/v9I+xCgosoavS3QzG2nqT61xXC2v2RMU1Yd+orzVtdhCCGoUc
qJeVMyxzUk9m8Fj47GYzUvtMqxuNmCMVOO73GnN8i5I2UcMizRszGlmuY39P
Q4c2iQyCar/2mxq2++D/L1xLTtuwMx7T1HXGim41nyNCOr5tRUEaW/3Mdem5
DANqUxnJSfrqzFgoGv7iznOzEh/nOXdn4326VyfJzdiIf71xAz1IP7zrEtl+
CGhEahOemQ4lRfi+fyoHcJuPheq0sXCElLx8IDIMuEIqueZ31XIDa7u8xPo7
DM/Y2QRdPqePmLcDWwN/y2ucmzDlYWHHvtE9JhzWmG9I5CYUw5LLCYZzuHKb
tMIbcSWh5hY5IsvQMnBlFmdMbasIpmd26vvFcmZIv9AvKhWTxkCzIhv81BHA
c84wZJ8s5DiwCmn3KVLkVAmRp9fVR6srNc5GB/oV75dnOtlGL2Awm+i0Ugn0
2k5gjh7SYQ62BtT/vS1giwnWaxmTkJREzyTM9Ii1I2mOIeWMJIWURrtaL6kz
DO/MaiDEffwRp85QEycwPpxtinU8kr+tPmPbM4EG0ekwMKXCD1F7aFk87KLf
cAYnkB3XKXgd1/1f9fuxYQaDPJttZ2wpqKkVRqFTr4SZRKX632fuuE/sepcp
ubnSasEBAlUTa45XBvyqo5pAlEnrSDfGUbV9HEF+EcxfOZmpbfe2l2V5N3JI
Db4g6ryhVP6py3e2nqUQ6ln4k0yC/tJpZE5Kt9+xraPC6Ypr4V1YLOKlRici
vyEpuooU8iyR/f4k2SeCFLf96fxlCKnJfE7Sl+X1iUFhcITR4VUWS7sKdp+S
nCswmy5SgTlOw1kAYf7gxra9w8wlJp9hF+yXrsunjxAy5/PHRZLhceRr6Xw7
qBVN3vN2eHKGW7xyk8r+Cv5apsjSZxYXNU5xcxHCdk/A+ov4Xdkmm7R6UZ+O
Micdy6oWe/Yq7MLiFfeW4LedkQgER2Og6Cm24D0N2RYu8XnJeE1S769+INRE
w7/J1EiSZHFcIVIsN0Oc2l9DBk+8yMzx0upe/Nw+FoOVuFNzCGZ+bEdqxDh2
3h9yPoRTBQmam98xIOJi1TcKdHCBcfZKkU3+csLJOMSz/vyPLERMAZVsx54H
1L9+hl9t7MPc5Y/C9T/lSHnHvRfMnxPTNL97x4A1hTSkRkVlaaEZnn+xXGgv
UIWfKDPdkiAz3WgEC1cdBJv5ySW9nFd6XOptzw5HZAjZ7LALtk45pqFrak9N
+gOzBmC9PbEiJEB8QjL3exZ5anAnHqarcVAVLlE2MWuu3BdY/h3oeogjT5/o
ISqBDta//PGNcql1wMOGPiajVWK7H/JQAk27YnJrdpNxIgJzVlEY/4Pb4OTZ
GyGxgzT0I/oJsIm1KK6zJAObFY0QIjQ3epi+JvSPLzv7v9iEWJ4lVXzGCN3x
HrBlEmznh9iGw862gMVnMJuygpUHZfVROPpThF+w/+ZccffbChkXcVq05f03
zZZFm3jBI5foJhDEPNYH3L3DcGk3Y8vXaVmZEdxyvks9dkVKIKni6ZrwhhjW
xiajCnVI/njeaLtVC0kOHey3POUttCIeDxOwa3l/4UlMBOmclL52CJVJrDZ9
BaCDy5ngoKg3mo9HNV/j/f6yLPoFp59RaxRGIFQFgeMk7dJ0fM/tQnPiy4YS
vl6ggwi3ilKUcBUnD4uSfeyBW6o75pTh/WyLdy1ZyefaVLG8CQ6e9ZfTAy78
Jha//3B2m6+eQFq8VUo/8Eq7qMBNDMn+l9XFh0akVcLzWI0xEjp59+94Ee+O
psHkuxBIabkAifhkGdV3o/RNtVYdDJ1peXAYRwH71LQWsEzOdOz8Qitc5rLS
A82rpkt6FVD0GfjTYeRzSlmCk0MLPTjV1pCbuM0qXrEA1oEFQI0hMces75us
EfQViOktO5P44Nc556FHOjAF4zSPb1Flm3tBsCVm1D5u5zqmN3jlbIf2pszq
fhiIfop9dFXdu6PY6yRxLwvmZME2SrrX9JXzJu1ENp+e7mo49vh8namVV04U
SzfnJK33iu+ERdJdJYZYVZkX/5u66Q1ewNQURqHj7S4qkO4cjwn343nvtkbT
m1ct3Tc9m4ruMparXn5wL1m5dvyU3wbe5a1Z/aHClY076FiAEQog9HrEIJmw
oTh5lsrUeIVnu2BTTH4UFyb7rLnylag+KLBojBBIoORT8nM6xanVDa98C8Y6
dCRdNufsiIgOoianXACtG3l/c5P9H8K6OmmtIbbQPIXBJ1TA7RTVJuOsIKqh
q61VeLUQPj+XiI5tYsyLz7rzDA+q8svSC17mtPXyN1I0GQxVKdoCxMW2geDl
IWePV8A7jKMmraMO/MfOn0qFzq/ZaOh8sfOQ2LQ6XQ0UsrAg9UdzRZAP7a5I
77c9A+89ywvb3D1bPqky4AO8is560K2OJ/LrIXEeJNz0ND2rJmhaXzDdT1Z3
kcz/838nymqeqOh765hYbt9ENrfIHl3ANCTD9iz29KmrWXYlBqfZtJodBQm+
tS+Q7cTw2rtN9P92O60pab6CbFUxSc4GTA8HQR+Q2JrOBrA4zWbWcRaDCIZq
aHApu5gCh17w5QJszH6WS/uZmpeMmjhWyYBNY3W0txPAUTUmleMJvjgqm+IY
MdC8+YisAnruUTVhSRyQu3M2e4shzzcmtLgTZPdyuvWRK+ka6VsYZv8G/mD2
ANXK+AHldPo0VObdz0gxSTu4tNLfjxpMswJ7Eop41Alk/4tz19/eY/89sEnT
9m7PGp7WIQVDKvVKGUIOaF1wIbrUnOAq18q5WCvHbcNIVgQwuJbwkB3Sm19U
Z2mpZO2HsOtKjw9IrmLWgnUjIAjnzJMCmt3RD2B3aNtnyUM+1QoxbzQkLSrB
GiBbSvcjQ8YDaQTOujaXeR7SJHHr87CRSvhnmqYOJQXS3L95rYt3mJvd0x4Z
aESFrug8iS0QqoSm0vRj4y5ttPGP9H+a6x6vIDlGOk2BLTGByZUJrvyHMwju
3b+FIrhIuPxChGZA81Gc2YvcMeoyayo6uIQMdQL0HwnoVWUFnMdtMrk3jRMm
i/Q4NtPGq7UyLS9BrjynxBq099EgjVz8PLQB7cB8w2EVlywzzGvm73NJE2Dg
52T7UgP9/ozDuztU1AEcXUezc2m09lIcjnBrtk7kfTT+oj3XTgxYGpOQPwgH
5M46PMdwNyZOqNsVtOh6URlS3nuuUZa3jae3E4jGGZtOre/I8reSxCFULOXz
4aoMZUr4U3Ee9psTjtNyHUVKpou5DddZRwvyr4P1nL5QbBb1cMaevmP1FtJx
1wxtIVfOT15+z57jSgukzCVJuckVOIcEtYHBwuP9KNWFh5YGYOKLRtNf7j7x
5/yrDzcb+7YAuaMRzDc4yCny64LAeRu6INuBfiXsQC6Rysj3zr8maiLLt9dW
a8ZqBYApjbHpYI2USiwoeEhWyrKyvbBOY0A1tTX2y3EthZse2iH63LjZdqF5
UfrDEeRpHeyRrL+l0VcQjuTt63nmKDB2CcyACyIeDJybXMKm3duOZeK+uIZe
cxj1LN3oFRhJdGRTOwQv0js50OZdxDE+nrYffSCBb4mbI9WOU9FHXa8q2Lnc
2PTKPV84rpIxZ+YvqO0EHLnFcZG8NgqL4mJZl/k9Yh7EY+1N1eeIImJsqvKa
rXy5zMvTse4TFI/SzzpAjFg6lRg/MOMxfV3HKoLRVzt+b5BMA2DKMRl2H2cO
H86XUfBV4W9XMYMREgf7KkeSQ6aW5QCJVMY3ghaYfOR0YGKXfa3yHc7MKg/m
i4TxWcVj3HGJp0lTz35ytDARudnPNtlZvU4FpLMRb7khT91No42Xr1N7WPZN
s7ZSxOvfoBcis/b14eg6wEfSe2xu6vygO+STglhLqLOW4sAgnEibQgQ8qWjC
MScNh+yCDM7/D+E4TX5NXDm5OS6qcldeVlbOpvvdnU9YDCjjkwpfck7V/cHs
uFerR1o8hKIhhvBPFW2ZXHc0P49euypOxXaYtOSwplrb5KzVnNsj5qsbEH1p
Q3x+IcdH68+f+NODVJBJbTbqW7V0PvomdiejVdyMUvlBoHDabeI0mbC9tWLp
z1AhGnptKsa7PmrwPuJiIEpE/7GLuuhLzikO0theoE+nxYM/Fkb2mZmo6rS2
EibpBRyzl71FxY+e47at1T+EY3SvzcdHK8I6aS+yEZEYFntcedHpoVnlq4Fp
JoTaODW2Wa56dcjBmR8FJePEgaChWClN0cejRbFQ4wGshQpPxaF+26rvh9FK
HpysieGsJfS8TlGV6IQQYIdlzbbe1dw26U57CimoQbL5sRQ/VycjPk8tQspo
RIMQRQInNeS2GkxEPD6M2PV0G9jWqsBMdIEdd+wa96rWqwZg4oArPJSc7pYc
XtT8B6kOvTBUz7aedRPJKgkSR3eoSE26ey/9+bhTzgRnb5S1OIk1hb5TP+ay
09uEMN/uj9Vx00HhrNP4rYuJp9ZTlVmu1NGFg/7I5lICqNAdtZE9km1bm/6C
lL9NRTwL61iqql8EqP70MXpgy3Um7EPzzQ347ioJxSaply2RoMERI3JNpn3Y
WkNneNQF9A+XmYcWZNTqnATdpTws4awjg3831dXWnyJXy1KcPtslq18/PkfI
4bWG2D+4MYbOQ+UupKTgQuB4/XgMDOqs/tcYAf6WYIDFRJ8EM9aXbNRIV9fz
jZOTzu9NBkxzcBI78B7biit/CP+SydCF3ndPaU7/hkuc8N3h9fW8bIc6Z1Oh
7U2ApLOwLfwYk2gJZtyYibv1CzyfqKM8Ft/rN5qBUjMqQ3wjhgNposi80/IE
m2TV7vpxsB6uGbiSHLD188YrmCXq3SKNws03YErxJFyTDsIKZcn5R5X9ZEAy
+DRP9ZOZVp8RJeV7qZTScW0pLE7r8veKnxrfSrPN8Pour5+byhKQSlSXMbYP
wiE0UmKGj3+9s0Szr+yubKRXwo3zZWtzYnXhUgfzCApCMh0INugIcY/kvqta
DATcrZiaNnRzUq4iqXCzS7ZtiuzusAtqX8C5gF+RRpLUMOFIGbNCKSOWX+je
C1Tmnm3qVn6/h06CtjIKj0dKwH+pZorbkQAA5uXG7P8NoEKnTppKIxj+oxof
cVCz+xbbzVfK6/KSy0C2RvaDfYYNDWfl6NxbkBs5Ud4kkp6Cxjk7d8dnkKNV
xIUW2WQrDnC1gFpyBCdQVIESJNBy8jjP99lLAqxIEKh0zXIKSbI6iux+sAgG
8L1Ai52433xLEug1LbHcbadxKDbq1FfHEgrVjjXCkrTCG+1ppewokncuMNXG
crW1f/utSzhIyHXMT1ps/H3HOTiPSA6x6dB3HNB6+wmBQ6eQXf8MXKoHiLIh
sKKGSRJlCaJhsReEYrnQFoyz/cfvrbOrjqlK7dUElIC7RSQ/zGIGedZR7x6Y
1AcGJ37SzrQtduK6BDN6ouorgSPViiu1xlWizEzRxmE1aTeupGC5OLW2jhcv
JAjzsCWW54Hys2nicH1OsMtEkGVMn9YPic8nI+9IYUbr1rcFOwBfbOfr+9qY
n61RpCNLAJEE4NfdCaM8u9w9cgCKcA1qAUVUg+tPRDWxLI2qlQXc62Ff9VgA
q/jyIwlSKBFSVjj7J4rdQpB9jH8ulserFj5frQAZqg+NtVraONMWjvx/pHrX
gzGnIkWKBuSxQmaZlv7fSpcX+v93G6vKNiED0Qrl35SvWy6rXtfJ+HQMdRV4
rbn8a4YVusGaWJ7MnGMtWBEZd8alZb3Pl6SnHrTAbwoacWNE2WeGW27qkaI7
eVM39auCpbeXuFckRwdV5AIwOo/gfrYb/5B2EhmTV1Z4DVzkrrlrNV5fbRPy
Yj3Hdbx7be7Ptc/8BYkrGT+v8xeriRXxaDJUVtD18vvx5+moptI1viADaElB
qfHs2gTBvdxBCPWgJ3de3p+7mt0aQJjTodHoUV2gfz98mfbJgDn+/UNUvE4U
Iuz0yofFag4jTjNhcz2DpvQaTBiFQkgg3UJpOZaw1JCWpeBJO4Rn5bcbEOtQ
sZYigAec1gJUfAT/XvhFi0d/scKl2Iwwz8kiDlMTN9YWZlOKc7qTCWtVWzBc
7CClR/mnXOhzQAdoTQJ8N9kRViO6mCQjg5JXM2RkANGA1XWSH44FA+a+q9og
R83Dzkqp5iSt4ResFskjbxVsCu/LtHYHhh7K6PB0vhSZZ8JXLbiSE+/+ky1B
RAl/hTEs6ilZjcCfMvAuCDrQdvhT4dMMOPJBIarZ325520fmhAvczzf3QYNI
D68nXCx9i0KryPH9ClPw/dner/Cmi6yuJZY3L9nfRYCvz/WpWqsVuB4ydCLD
v4DgwEF+IPmLAFyVHvqkyq1vMb0/g9CfrquTXVIpltGbuwuZBncEIwy6Dlqh
IHKbHnjg7L4g1/jB9kAgmp3KRBRrVbpR3OKkcacadFBttKNOYUQrORFAO2YK
yIPpP3ZRvhrn9hUqQOpXgo13M9l5iQg1qFc8THnm35EgkcYeAuDwnZ8BBVQB
hIUWiAcvAlbvi70iozS94u9M+7CkxdDF9aBwPVN5NvUvziTFXdBRbCFJF+Ow
0wHBo2IPOhzcqEJyFZDeOcEeXPsn5ttbDht+W1FQeSC2qj77Tgn8YeKFTeIt
AXloCiBELJUBXhsY0hp3vg6tNGv9d3HN02EFRd3hE2Fy1q9CrC+uKHFF/UuN
p6Elwr6Nb4iBBnoHVBGWMM7po4FsuXF4XsCqIS+z83ILXUEHtHVezUGcInfJ
s2NSSpbVsuPoqerizkxQsEwUPfEJY1fldfSns2QDtuKowkL94AD3TTA8hl94
EzogwyGSy+NUCLNt9P9EO8wDLw/2KzUyjKrfq5CbO4I/XgrpBPv11xj7x/cL
Ccj02it7oUIEqJyp6BtujPjl9oR6zjWDOdcdGcHKeqCg9JRUGFTLGZXGm4ge
ZAwTHhQyGM5W+1iG+JsjOWgGYoTL9qsUh1uVSzO0nduNrs79Wnr4WNpWq+6Q
tpAGT8ehptU0a+3e9vHJqTGs/hdo1yLF99osY+eQCk6o70Zndvsx/f6Gs8Nq
GjeYgnt32uH303Dol05Le0pdQ3PmGzeXYDKPGWY7zdRvrVP53oU8bNev3hU2
JaC5bicl1LNxRR7l+IRoMhwKh08P1ys3Wn7rDvw2A3FuQqf7FbZ4u4/JRIXD
TV42GoBDMaF/xOECc/FYNO3iM/tuIrtUv4PcTRWEyJcz2trwujkGLMu9Nl8K
IHD4b65hCaya1MXOulPoIoheceMCIyZAHTdEBV/IfE69OYV3FmF3riWNbsiG
gA9ifl654MP1fS5kFG012OJoyuRwH1BtYkhn14QNDUWh0AtqhJJTKwDbWqXQ
BoaN7/5SuStrSIW7V9m72J2eVhPBToW8R8aJ5yfSnfUFdeztxGTQDm2K/jj4
hvzTAHz2mWnmEWDTpgvPTwZm0SJA8pEx7ZCH8KAR6VocJRsfxjOdUZzQ7NF1
1fj1rgEghO7pMyBHe0gnBLN8GFP6dDhg/gb5skpwOpyuzEfijfsEnkRonweY
4cQZTlQ+n6tcEO2lN1OEDmjcK4tYp9dp47kdqVwF0QTrgl4WBy1muUJzL+FF
Dzj9rp/Ot9S+GkZXxZSU2fuV+ANj8lomHFnKtlh+C76fF3Gt3SrJaWhgCB8p
fx2MlKod6prX/v7Ub0Zd64VEknpTLUKkRI/Fz0JYRfn6/3bdn5ChNonB8VHI
BkhiYRpG2K/pR8oC/v7XH1b0aQzqcxrK8ffaw0U4nVJOoxJN5ChEVWVRJIui
yWYofNoFbUb1cwO+7uCSuz1aKYkw7SXU3kICFF6BPQngG37qDWz6macYkD0C
U6+fhthR0aAI5aW9xHK611w5TTO+NoH3dpxT6D6loyCUwDFkkceb+tEMAqqu
UEepVGnanN5H4/OORV6cNkBUmhM29+kacvUR4JlYDzUV8IHxHbUJGNfj8o85
f7A3jckJ5x9UDAGxrTSqD2YYiuGpmc2wyouPb6637f4rI576LNS27mbvSdlA
Z0fOMdKr2UGrOeIHsXvoOpruCueMFbVSORNC5P0OA1XQLovozkpYIq7W3JjP
Yr0OnOY5heYcE6ZhVtCpiv0YeLIMRQDnsm9/yXnzHldE2ys6Zuk2CoJfvMHb
lvLhq9dYvshtK9gFEJbOzxHi6KfsyW7wArxqFxJHEFfktfNTzRJtafFGxInT
hlwVbT7ZxF4vmH3FWyJKSN9xZToIJkPhYXE+hkUy/0H2QTntdRIQLRfG1L/D
0SyTK5mgd+ffQpfQb7+F7FvSW3ysaD/li7niQt518KzWRyJJstUOqYD+XCdX
V57af6JqtKCh+yK0WuT6/jPcFGRkf7VHLyUqyXTCY82ZjKKDQq4h0EB6cBrD
hbjJ7Ic9nIIJze+yapuNQDIcSYb0NcQVo+1Mwm9mEL6RZBz0ZGPZWQDnWQLJ
VVIkFz4DtSDKtE/P/8Tx4Pm/7VUWh8xQAMv2A+3QxgDM2hJQcot16vH5OyEk
vUrVqBLDQg+TRseY2NSJKbdCiw3ztOkJzsxRw/75jb+U5y5QC/QXzUPkhLef
FHLtvAqnnZ9SfDR2ZNtmMeeeZT4ueoryvNLVM06Zu2NmD1dor1NoqNNpyom+
szfrwRmZfoweK73FvKbVipWi4ZsLN+oOGzzMTCzsEKhZaMppojbdB07bUlwA
Q6gFgQcybdq1UposQbK5RHyzkNSwAThPSij4sD7gbdnj/ewuH34LFbToTJCI
U0Ge/F/c7IZwxDLNTx/K5Qxto2SknPDpjgHSBgpf1E0dYcq+1HIH+8oo715A
D2mSSckeTOQe/KTyBxtSZWqJvHJ3Th0XgLKtrZMRrS9vzAKvcpq39X9iQpfs
W0632JuwOAzWzUWSYgGLrD6b0cgZaYh+kr7dsqi2k8WBkgtPl+UcCSmpkv6/
gFbK+9TTGTA5SNAKA8gR2d7vUNEU7X+MJFEK+6foBKOh6LDM0t2MtFrQWmg0
XiJy3YD/7BxYOHD/VbfwsNfDozjWNxMJgaK5X4+vBkNltUEcKrd7Azv3wy24
25XUka8Jp0KKOEI2Qid2xFPhlqjr47PQeNRdqj9AMhEA043pQPZQhIZ06+vH
IFe/uOE/NqjT7XUYmpuhgRDuaRM9rtZPUqze+0SgZnYPdmqg8JmhYxdKnUzR
pnI84ZH3L61bqQKKkJ9HeSxDK8p4X+xSg7G4Mm1vO8sIi4ebT0j7qVkLYay0
CYxpQN4IrnItIM4jdJtB1GIMdyEd+iJmFcMZD49ZHxsHsjmiK+b2fs1kLv4W
icF3go/6HGse8accBHPXedDBmac9hK1cYy6sKjZN639bz+rF9hQ8IEHxC0dQ
+RvdoLE7omglsvgpSrPi8IMQCm14ed/1alrfglhXg/AVznH4Dg9gsYuxpaIf
8Ch3XbtXWFehaxVQQOCvPqq/sFaJ1dQ7SbhKR22p0NlEL4tSMrS9Q+EgM3T6
Ym4DseMGGnroUNp4zBDzo3Ks/a0jVOjmAHl/AP0hbrCNLsD0acLMZfYPlgZm
xiqkfSBzE/TuKEp+Ts+YAzu9rvRr2PUHdBF2/9Y137Jbo+WiFVBDQa6vrlQX
kuFAwDTQZWIyybcLIs+2fqT+e4i9xke2+XbmEth55soIdbaxHggX5VFWd81V
RDUeIWr1NurLKTaAABdiKdZBCQ3sBHHTSkpT4j32iPWkKInRkWgH+cVukzkt
kAxlBtqAQDpVcc/0MeVV5W+DYrHj4MYkPg7O6r+7T1sGUHeWn3AFSJMjFveD
fW/sEIrsRRaZPJ1Zd5zr5BeSzykQ2WuLQxZ0GWnA0Mn4B98Sc/mC9iGHKTGQ
HpID0Ajmtag4u/cha0BD07X/JGewY/3zzebSH7PO8CVf+IQ4Qq3UZ5iaOfAX
VA7ShvxTmLYta6ufzsV0ke+k6wPIT05AcW1mBXTpcJqZxoQ3cRU2IXksanVF
TwUJz0OrivGnpGBawbVJY6SoogVBDxZJNh6MXLQ88RIwSZPlh/PAZtkgM85u
VbsBtCGcvBbtivFx08DBepD0TcMLVyVprN0nuVfTP1cttiDcvXaPjJrwbv+A
9zUk86xnPVZ40rp95LyjE+Yeg/Dca6Xec+XASWTfWXd+aKic2whrRTtG9sCs
ZuQhI9HdgYrx4Cf1ZHUcofamcU1vWRDfJwZo7Blblhj5qyfc47SnzgCQVZ1M
aEYzXe1mifSfZZdbhHZZ+zk0UfA0Hoh1u4dY16OElcDlISRg7IhPh88tmeOc
2q9ykozRBGkvOSdSRYNpwAnw7EswJDIK2wxePfNcoNtkveMa9nRmWpPFkz10
0K9N0/7lZ9DOba2Qrw6JFaCcTym/VTiOc9GInWSJdz42ELbFC1/QzU/sKkf+
ebC6k8KvGK427vSqnPTEx206HVFXT4/oOYHDSsnJ0Aq6BkUMPdfXshFUIAQg
20iCrHfIdEK117UJ9CPiZB8ZVpUo71AMr6qD0/9ErccOTvJ8hNyKpF9bg3Ea
KRC9ga7BR62/KZR/COGEGR+mz8/1+vqLi8dZ4lvABC1CLrPrF29rXPGAnF4Y
XVygALmSTn0FYSYE2/TOTeWuyLKS2C6y9ZNQEr+6p4acfaUwoewECWXVUZIh
qUnC6XPEKF0X9KoQcetdYOsuIhmP4I6IzGRj2D6GGijaj+Fcn4uhaz35y1BG
TvdNZqf6jD5kSM0tKUudVJPdoZg+lfXxN79S2xujxVOm5UPlrCokYP3v2Lq9
AWFsTL3Cw/khh60TbeNHnA2GIOj0j/ehdT0FxGgofxyBlSPOHIWekJgJkgyo
e0RPCtCpo6I2TkYY0yADDpmNqNGwbm2zwk5XEG6y7CHIfBcSvDrwhho1KkbV
nd65yFo/dMVo8xg2X8BClFpnaoDKuhpsWucVCsbLEwhgOpOZh5BLgCCGpDZ9
r9CWhbL9m6egWeJNUsA9QVSBvVzLp5Ofn6sc+zZkK6JPnICnt9YkZwLvl54p
D+Gp+FyBeNjjhxDeAnXJFSOeTL3igXDlqrnmZodT9XGwUXcxxQLOHURuFcng
75k0c3H9JPCEkY5MchfzTSU0sxWDp+I0Xvi3tyHaeCVTLRQirqyMIWJ8Ou40
P0PQw44zrFG3wVOu3xMc67TmNERwjxo6EhWuHwzIGFGo4zaRBna79V19LnNq
3PyG/Mjz8KsoRtJoexsWUZbDoi9z2OBoUc0dhLg6KludF37wnoUg0lkHT0Z1
uo28RHYmpQE30uBe9qqCE6xr2ZXWOv6kYHq/NuFvJTvu7Z7p2Py2VbddvU4H
7iASIVUzMJo+JPYbrHZDfN1hjd6mS0NU0KAIvXmwqq54NynTFSTatNZ6vPd/
v9WzmwyjaqAuxwjFHbIlNDSzFBdPO9JeVRHMrirWW6ZV7nI7JQ0UR1QnTfMq
gE7LCPIjqix9HDGsNsZf8YfHP0iybsz2DDiGYxADoXU7ZpjOXco7B3C9wgup
ge4hmQamhVuTqUh7lOwPM5tp7wrgd/KztzdcArklUAOhWtA16fz1E6HaLjRx
vk9PMl3nw2qNx/HMVqLgd/N3wKa559EIOSgziGgpjH0pR2acZ2chfAM+pxe2
TaJjT0wldApxOmX+THXRyyfAby68lHsT4ALByDs9BPh2wrIoZIPou1Tprc37
Gq5Dj1S1SI5P5OmwBk/UlRJQbNqbeTGtUyyjY3cPKqRTHtBKFQQ5IroBNszI
EjkrI9COafr1FKjMjj/8mX+G3PQV4CC827gUQLnQosTT0qK6kx+tvZKh3GYN
87cdWxV90mUUQALZu8d2c+JAi7I00rTVz3/LcFsSeQ0odHuzJ9mczBpPbMiC
IZmH51D1209SSDD3+1VT28oluQcrkZoTfeHfOc8G2Cc0IZsrEZ9MCoRrPwSN
noIYX0AdeujPytKkcyYhk1LBu0JZupETiKBSxdJqdbMEUViRxzgmigkKGtO2
NoudmItIkGJZgS+UuhlcoW+a6ItWaB9WrdnO8UljXsq7hC6wWyrZntPYmdTa
TrVSROszLjTBCIymAnRzbITTDIY4vo7HlKwG1t4KAMvXBlpntXcAHXUmYHy8
fYOMeD3MWHG/ioSArsjueLqD8CPTVUuVk06H83vMEHaeUVIyeP9hl/YGa+ko
xuDqR/17iAU6XfRwIGVoMhSEGWspJEir3wn/BFOI/V9pJTenR7tqCMfEYWiX
T9hQTHNS3rhAc2fYopRTW8bAkOifzdVAPttD4PHn40XYNBBrQO95JqdZnljq
x7hkASWCAi5Boi9Dub4Xh/D38GNxb2dJttsG1d4wn3w+29QzyrM/io0w6nOd
+uQH7kE/zJPdg8Ykc6q03ljeFFfC7fEdc/JDhez5DcvbJBxqH0tEnMi5jhB6
OmG7/fUfRGq+9gofq1Ys

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EoFUsywSfEfrxkXpAXyWRgKGGLrcksMAP2CtI2MwTcTRk4hkLiPhrA+uVpbBIeKBFEVSDkPkH/Og7K4OchcWpBeNwcrnyA+FJp1S2vmrtGJbpXgrl3TxM/zWvrD+m0QxeA8pn67VWspB5h88zF8nyrFg0W11wwGOo1e+QfUvRZXhMVucA5PrLp1GnNk55WiiPmdR7r5+agVh6QdcOxMNqKhXkoYL6EG2IATXybxQr8cRx6TJqMDfU6UUP5vyWFBBcK10vG9HTY8k+bJGEUZwkzstafWKxUaL7UFqUd2n6g/wpqtuEquGzpZpR2cmVV00enZz03OGg5DlxjFYfXBev9pa9Ah7jrUT0NjHWaQumUFNw7zhRHiAzaPWiFasjYZv33i4maiyexIVqXnyFaLxxGr1q+icm7N2dPV43qdcwU5GwOMGsEJI6unQpceO+BDJ1cSB8UW9gw2ZfX5HpTs7F+Q96Z0zAJkg9hE7ZauyhyLqnH2aAK0kC8+VvS4euhbwkudE47YN2DpxL+4LBjaIvdP3UoQyfyyB6aKvwwMFoPTp9rIdJOFH9ZbKw37NBumtLG1e1eqjN/mtGaAJk+fzzQbCZEXhaixBkM7ODUEISSUMz0cjXj+/0JnP7W1i3QRfUFq0NK1AEc4xtjSP6xJfugp37mBG8LFvB8qGz3yrUhpC2zuMIimz0oJyU6hd9fMoukyGx6GxosZKTRopYcJGaPMtV11IU6OPvfZzrLwSNJXERFfPmtaN7o34XiAlb09Q0LkEC4lp56H6eWzpxQ2W0qE"
`endif