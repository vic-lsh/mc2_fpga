// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SxO9FLwjXcxm+G+jmn4C93iQwgf7dV5x+pDXl1twhDX/vHOPLz4byHqojc9I
0gg7sG6AhEBVe01QZb8B/jSYFT/6l60dtFxzeadQIFOAfx3f7y4l54P3EQWb
8IIE/fX0tbbxPR40dpeP6IQvhwLRumdPtei3IAd2n6crv8W0E08LlSz0HXhF
n/iqQCVAvTV/AConL40gbbG/gf+xWxqVsaxx8mJ9urBHZfvL0o0amK0x48No
epqc2oEgrBkCjUNS7UHEojaWdRMaeddpBHwH9qYph5GpuTLfZPdMKa4XmUoY
yIbB8Y4s0Ut2GguEMbANdyqaTfD6d3hEO7ExjFNm1g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Vp1ozUBQVL3ka6jXy5B+H1/3MqYfwICnOo81qR0ypMJNURjwjdRthMmS+oOh
NndidULQ2Vipl2dtdBFv877FfLASORSI5S+JBM4e6P7OFJ5CRIDVw7sbQUqd
SQxCqyg/mRYv46t1vi5u9alPPoDpVbs1cMxGPvKHXf0PJsJAKbjF5OLEYCDu
C/lBhH0sXtREH2fJXNMtZxJo5/SXYVH2tOETcuIINNl92e+mI2QsJaVonad0
01WKPb6YDG5T5LZ4c5ctDez0nKn+TQQrxvVu5PooMrGiCchrIg8TkRZ3htJU
2sAjRsJlzHxLOUlUtv2bl9x+deDbhYGc9cp80+LZxQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JGDGmCve6O0oGSzKEmVSRC3SPuALeeUqLDRvyXf65CGuxEPVRmdc0s5f3DUp
mQE/GzGPSeJ+7zL1rXOR2y/xK9KtDJ/X3S0b18xIVZ9YYVpR1daRMVgXSP4W
WnDT+MVpsqOJv5jGodx1GKg64DYT0qT2Fgj/eG/ue5FiXsBLQlhUYWZMe5B2
yLH6feluXh1DuPL/EBE4Ah9lC7srw1TBIgWJ2T/5VPjJGVfUMhI3xozCH4OD
Hf64ZSb88bDY9i5Ct3QUJ7MaXZjoK3F3MjX31EQW2mvftojFdXz77Csduusu
HYM2WC42NutcuSZAB0WFdbYWDYlNof3ZMabMlMY8cg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Xyb9LlZwA5Z7vx5OJo/5/uToxQXc+4k0kCMwCR6itazn8C12pakFIRKHhLdi
QRCnxIhym5TRhPbAAyMAYqPtCDTRgjwuPgavaQdoooYFGfax412IYvgS9TTE
1HUIGgs3413ZVncFa3yTMlNlILBxmZ1YbeaH8FPqjZo7MFxAIsFkg6cU9+pq
NUm/OOx/JnML8RKVVdSfr6G0VgKDiS5k8VWzMut9dFONYDbmrL7gO+k7a6x0
qAqB1YhcwhbYRzOslBZ9Xj9ZJaD0444VktT1q6JKP6Id7z93m+E/B1T34twT
oAY0IF+qRs4MlJNtQP/oEQsYfXc/vKPDNff7fzb4jg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
i0a8/dtlPUC1gQZzsQ1cwc2QIF/pwx6k+E3kmO4zeiYNpC5HuhWd+rVCiYXO
mzOZfvSAYg+HwER6KBSkII6zWuCiwVhe20Ua8c298cYe1SE1HMUAB2cPg6Wi
7n0bIK2UJh2N/SPDttAlhVn2BtQTxVHlqn4W5FwVYm/jj4hsil4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ajQO3+0u1X31iU0rXmnp13Knr12G2xIoUEkj6VtHrp9HlipijwuZFKEaRc9G
cACB29/Pwh6YmOKvAH13TKQnaQwX8zXtJ1bNRgHNWnGZ8zW6/mwC1luYq0XE
+oBhZhf+B10WtDwHLpvGs+mXMDSw1uZ0YVRIW1N0yRz262trnFU8moC9RK/F
bZuQTZe02r/PHZKMoYN4zsuAJoKzMuaFk5005bMPCH3PYSJhhfBjyNoN+XUN
h02M52zigKc/RxCaEvrVakrvyKUlqUqX/GcZ0WZ64xKLnQrXk7w5TyALWplc
0Njfg3OL00rIwLUFeynz9EgLPuMNgTJiS7etOkIgaYzcLIX7K3BGfeLebIaW
YC7UL6sIIVMc2L1RI0nVudce/chILXUpEv/RsgfPFH5hIMgydDTZwWchWdk6
Si9FSivWVzl2y9ERTSY6uDIgjrGDqCTXfcEtoJThPq7U8DmsT5FstzdviUyk
igRao3cpNpl0Jf6Zerxt7CnpN01rFNaZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bIPrUtkplgJsfe6U6LR07BgxaHcs1Daf4qCKbRSNKUUdxkXdtGO6GUbJCnSu
cvF1CGOfK24wi73udLGTn8LtG2fD3Rr/bCmi/E6LECsospdeMnUxuwH5D6Xy
qMv69pyhKKbXakCbyQsykirLZESw5Iw4VD+ry0sWUDZDEDvJ59o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Wz59fn/8mg2JWi1FXwtLIhVbHnFcm9It5n/0wMy/uWYoPGjIHkU6G6yJdX2P
NSZq5s/ahbgX/Jr+tumlXuByLSGrT5cfCe+Da6Txjgv/0b1l2IzMnxVqutKE
fBIb1rWeeuK06DGg1p1rg91iLtFDX4X7Caiit+4JnJeU2Y0+ajY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 49520)
`pragma protect data_block
YTs/ETqM+m/nfAusBklPnMs8fOaISCtEDic9mVb5nDPfZtnEKXKpr9aO3kBG
Zh+beBMffIJMC3TUucsinwsaMs4xirR99dDSUQcFFOWY0NvNO4dJg4vlO4QQ
UOEmhIaEJrIWgrU3NMm8vdXjeXP7u3ut0Y+GDXIB06xpFHaWq1S1XTIJTpkg
vTburWmGYvR22b6RX+kTkjX+1pr+ljlnRc4xVBeWYUj75ywcK0ZcjuNUrcyV
BaJkaMFY80Rgq5IN9JuzG4Q4zA2/+xIxZk/FMikzH2YDR687ae0JS060udoW
3PlA9xP+tTSVNdfJbcCKA8pcfPVD3iTYQwpUTAx/O1l1I7ucVjigf4nFLkXr
6EHMzRDlb32j/NRSZ0eBUjL30/2Cb6BdF9fRYFZl2ugrM5F0BvfRXWxG8IoY
gBACzHkEtSWu/e1Qak88eWFd1Ws3J8rh3SrjzItBkKoRvnZXPMqKG0BzN51f
UoSFSg0DH/SIw74TX7XpbtP0ZJnek5rbAD/4NXfQp9kPRiKb5sPZmwFPRqmE
56BhnleRYpcOe1ASxTtNTjtElAw+cRXrDqQnsua9tRRaijQTEPnE7c1tYeuH
1nyrFUb8HLBd6x7YiXtrO9DusZHo88KNSvwXbBmpH5MYNsQLIXRTP2hEos22
1T6GGAoyAIXOtWm+UhtG+3qcYGZcGGOCcCYHAxb29BbKQLHhO1GehcHfCorq
/ksHhkLvAeX+mDq/qntCPhEzdjuzUITGh3XnWCtTu7Q1UXTrYHNqfSf2ovQF
/mh85eGqezwqos9oXzy9vTY01zNS8lDoJ+Kvbl8Z6UppD2+0ytxQfecC4Fma
PAxPPhnvN3GJ1QtWT/NLF3H5vg1mUoCgaELC/kWQykFB04R8fNXfZ0kkGPqv
/+EQTzqno+4tNd1dvtpvHIU8/02qLCNR+FQricGJD+lVre7/lP1rrcKLc8ck
3eMTu/T3xFi8kcuGhHR5ehH9/AT063az+T5rgY57wELKyh41bB1c5CtmYlVu
nTDE/g7dfW9eskj7a0/TqZyZAtuzrElgAXE+1XVSWRZGsSxYjMBLAWUTeah6
7El6ILeXMv6YwquFEiiZpcEjYdMnTE+nPKmmGd9vCC078gJG6L63E0zS5Go7
I3senJQObH6xCYKsWqUqyaXcNzjHA1OmumVn+f1s6BluBkLWEFM9wD3bfDAW
KBGXGHbGRod1BqrbrGMCGcgJTdJH/EyUhRaCMO92G0Ku3H1ZWK9+W6uB2iGd
0vsAPBZBKlTTJ2Y4e+cSd/lBKX/JMDv5CjORyfiDOzY7xWmUO3Nzfqtd4Bp9
XcXbwu/p7sH6eziJyVY8oUyevtYkAz+OaJQcAr9hAAHjFoLEzVpppU35NC5G
LGcDnhrAIvFyOvI1zgaQFQNRBaxViWe3ZSQH9OBWNTlXbytLluK79pOIHsu3
9+wGG8UQoHfP8AMTRCEzDtibbyGlnH/Tc60BW3YSFw+xJ5GrH4qSSphIChv9
+krzrmcq6VKWaJWz4S43loCrGghvHNypCYaFTpMFJSN8tz/8KL2ucLU+SaZF
Te6xQCCEkiOP0Ouk4ieffMn0jMLwJe8f2zbsru+6YMltcce+9bj7P758kc4W
rrv83RepCl31n4nwhGJqrvoEqBFxZ1GZQN16RdngA0+eV6uRbRN8z0GwgBiv
hD5JJRIx2YdDlb/s6WuwS6aFkMIWbPaLzXHtL0lXAhGEfsEMK6DHPc6dIbfx
E5+ASOciZhmgJi+w9nEN3QX4VjDeusADZWVbSS0n9gMDd/z6jDBoVJB9fAe1
SiCJlH/98y/+TJLSuyaFiowdUDlEy1JvafiboE6CCtGeidox/m0g2w7Z5BLf
PYp8IXuErv5lmHQ7YWNqfRUwrs/+oP98PJC7wyjYYsDu9fKdBYzbx/SEYGV3
1aIgQa+sWaFeVwTuDH7pb6tNTZTlVnSk9uetFkIS1Vyydo5FPoxgtm4G5Lcy
3mmmOC9icXeXhH/y0dbU3JCtJEBO2J9Ley+ymjwyeekCpk+xrHqPNSxbwvEb
wiGG4LIRWIkGjvSvIO5haYrzr0DhwmAu0dhqCvFHLran9FUHiC3c7FDhieXk
fdE5Q92bqyt7/Nn418a8ZdI6nxLJvTg82LFu6OkNs2uKmelvcGRi9RGXvr1Z
5FEL78jba2oXy950oo7bFZPO6ay7hEVvmfpfr1oE2XTUa9hyTpObPibPcrUq
TPcD3RfPWILUebcpMNUp8ZIb6hTRYN38uqw5RVsM21+UTlDDH8y/qP77Jqx0
ydhZBMkqDU/Xdc9iuOKc8gIf8hiXp38zBBU0xuuFw4A36fXz6T/QRGu5bKtq
glWxoQxH/npeS7kB0nJx8J5r27ewaW42HnHH1rPPtulaANsmcWgaxOnDE4js
es+Czkh6Iyq0uDcCFSMmUYnz0G1Gsu3TTO0zdLZbp8tp03aBbp2SXIywVaMh
QdrOv0dfqrNQZfPFTWtwVD155aigaVm1V8jE4cvTy8Nw2i63Hg84tGNJzYol
cT9d1NPz9dEpNtoe265jyrp3ZfODSh/uQakKIhhdPPNYh1x/HmvCF6VWalXi
o/1HiGntfC7WlCjZ5UZ7jPitzhuAu9/smiWYiU0a1deTqp6ycFoWYzK7n3Hx
ST04ECr2xfY4Tn4NyN3jG2GjNUk3UWDNWcI7LeioTKVdD0D0iq9mKSmDZf7i
LZbk83lmVMF0tUI8Fx/hOp/8oOaKDikpGDJKTtMyOuS/WQ0zd6TsB0bWcNYW
PgF6HB14D81YCOLoL1iXK/Tt0JOEFUselJwyCG/6KtGbVJ2ZKwjgI46MIKbA
EodRwYOQtUrQzkhSY4gyDEzL6W3V4YiPIIZ3+maOgM0NDIKI+rHeMc/zeREe
MrPUX+d8ynMv0kUP7DD7rqsqH9VEpNh74eEkzarshf0hX00sMFgkRPYFIj4L
GZT3FcC5/yMReu6G9Wwf7tyfCqRiW7CLQCgpySWgTG5St9JZ0E4LxJmU9ihY
vXAX5T7/jacTLFrY98CP0PC42eYrd1dgjw2cg2IYXkuC3mIYsQA0oPPAg01B
fp24J0P6FFqm2jDkIAZJLHDYBxkEjZ/cHQBt8BQnuBpoCcV8qzlghpf4tYdl
5UVVDpFgSwGp6mvj/mbg4AanSNbXr2z4K1FyaU+K/8GpNjY5xMtzxPBFYvRK
CgjI+Nq4J31ezzcYbactHicxOA2vf2JioU+aRu2Ssl1LwG06PZsgmbXlhkW3
6nFnhcZkA3JiL4960FZpHyqH8bny524GJaB/th8166FekGiUTFq6w4gMbu1N
1JUGb0Q64Fl5toLS/TioW2ghT/sI7BWFbz4wie1oAVcqVoEBaEPa2Vu5T5fr
EThb92bXxkzObi8d4LEG79ZBADRYHacMY0f4z5yooRDasrj+86zwcPhDGCTQ
0NLJjyWM9jKOy8qLMNpvHLll9tSB2weRA4XWbeZyuIAbylpELS/Q8qEZE1rw
riO/Avs6XGWKmA2layfQ6/ot9xM6cIThshLSsrAOOS65VG1RZx5YguT99s2J
/+p8jSECqlSEYzyAjoOxsmOWR8JHhdAzr8LjZ7ZICovJRb10c3DOndDK7D0N
BhNA8nR7nRwZbDxxEwcYuO1KVXKy+2+ZpQ2unx77eAukOthNRbe274Egrnmv
ebsPrDpDxdJzVoYyQsNDjvca2MJQBRe8RscfW0XYbt8lC0ez6GjRbBxM1hQz
XxVDT7Gz5H/mUhHWD025Wfs0LAxMx+dM7ikzDXT2zqOvUSxOSitA7YA+i8g1
YCq5l/LlB79nwjOVUKxu8WbFw5tbQ4YBHtuKS8PUeQEEG6PFoNmi9METa6QP
TAuT4N5QRVT57OZ4ry3gRpj1xnbYbYPVOLKXa1zc3vQpIKSna5D6mqs1Gumz
L72uF8I3O4KmYdBmEtYznLB/UkfD8fkHRD1ARZa4YSDnKi0g/aN9p+IK1fFe
an3BF9UtNmph5zOwRY8aibsztR5iaXAcSmgIy4dUhY8M8C25+Rw+U3iGp+hc
kAmii+EQf8qBF00eMq9laZuL54fZtkWrnUmWZdxgaxjmpwcjnWWQMBMLdn6M
lIdiO+4WaC/xD06TgwM0CMaeBGU8eNGWpITNRyvbQ7wxydWmdJE1GAqNCeUT
XagkiIpsr/nMsdo1Rox8BJfRAO5NBSkIVZ2L+JwG5ewQ37xYmklbtE0MCzg3
81btD81wpq57JViH6j5RH8uuVrGnmsVsYIEIj8q3msDL2jnYMGBSPkvyT+nC
fiYnZPlv+ptdJL4nWzerR7SyiOny/ht8/MXPgS5XTJJEeL05qITsjb7K5WlL
jnHlcmaAO5/0b7N3gOa4YA0JPNy+9CuY+ahsAFalixfK8wicf2/jQ/zK/xjM
6sxQPsM6dvM9+SvPnP/bqb6FmNZ3WC9P4XQabMgu3lawiJenuvVTubbd1qwl
2Vep5a2/iVBAPUp5hLy1Qg50o6R++gXzgWnUab9KsO+rvMFG78PgGQ+tJqXj
8zyio+7FIu6lFg7u7lAFg4CQYwrZmwh2hTArkugbzqNqM/+QBKGgGx4hIkB9
6KCh73PexnOF1JhagHiQ5BL6vLGcxnTBrDrICY26Vio99PGeB1s4yTB0bjac
sWlwmDl7WcwpYcBsk76wRsNZta/tH2COXhAt3wLrWIQyEetJQQzJ9NRK3qWc
LvbQo4SvPFp3v3sz9aaHssq8U2UmXuf4u6QjsJRA/+xTZi//7p2ZaIRtsboQ
c+NNzCzwmMteOz3AWyhrwgZPSoc3kVng8pAOfp4B4GGBd+nyExd6zr/0eHPe
U+1uAKHnch5apJji6ow0/Uq8AAHQ+85RjxZbezJVPnoMwf6kFxKMTui4iBm4
EVco/es8La6CGi8SMc4Vt7oxyKQOOOKe5Bb5hLoi3JWI/YShPF3+BNWHDtTs
OlPM1VSIw5kzPporstYZkwTQXXg2QgjR7V1ZiYqzgdqnvzEN2LwfjVfoHmT6
obJ+5MUKwSdOIlK/c0ZSOVoERlu+TXWTnl6k9urOjGTF2pNGXVTa2lZNFFvH
xrYwxeIJgZmPPS82dQ0CC+va98E+NuADSO8cFlW+P1PsETxnRYYSP7l811iu
P8g2AOc1RgRHrZI5KXtvHxuPJnOPQSV9uiZWso28mIwdi45CKyroDnLUXb/m
9Nv4xHAEdLf/s1mzpYq8GJHkE3J1QBoigieJ6mFy8dZjEjYc+D6LNohPmHPp
OcVc53xDND4HIrjISoFWYcjF0tEIM5OahvUKrfC6MDpaoq3LiXMyQwhzG2vD
x+T6r6X7tkeTR4sqZMLrociSNg5UGASWByy+t6lZHr/T7rguUOOKVcW74YeP
OFtrV0xdfVUa3h6bXnL0OCnGjRPYJYM6uTYzAzCZoYrcbdlKanpbRC/udT8O
7yJWFhPzqEYn72dz6AlkW1SxUq4EAuTSkxXMwVuYaKuKJn+NWNLwZ5kM/nH2
Bqbue+XAamqH9FB/jfE+87AVFjMsqmBap9C8E7r8OQ0nqogk39L3C1MFkA37
GpWsRWuD641I2n8KmbbVDaKB+u4q52KAzgjpmZgw2SxXVLruioyLTb4M0xCV
UCV2FiaO6qh/FGQ1cGXxnEEhmdPoOLO7TxLXo18dCNY8k9P1mVKUgRIbqFmQ
iHUOvh/+e4/2jp19oInj47MvnJbIaXcmT64g8v3cdziajkCM4L/JdXmIrLd+
mruvi41FjNUJJ1PucYjsBaoQXygfOCXJElQjZxUjA9Y/EkC3T1ID3mx/M5oP
RwVrU5hjHwCLCk3Sel0GX5JvfIInVQpTJS6gB3v1NKg+u1TJLAv4hT6CP3r4
DAXP5wvszJ+kPfNskuX2r0ag4aTi10FUl9Rg4Aor4z1bh531YmIqaYq3TRsU
oGJpVCOsqfWSs/LD0e/KGkwoHHdcsTSfzIMW0hOktCtTbCgDayV1NFGlpp4+
5WQ5HXapGtConDbUn1XxvErGX8rL8oUMsOD2UzHttO6tB9AKn0RYx/uiiLrd
G2jlwUlNAYS5+F5ODCUrfBRyTeNce04O+42kuTqc4aRDQMUFMYI4P5reFjV2
kP20TKZQY/tPk2MS/OJUK6hYpeiU6mqqYAlzMLSGBQUNDUqVp5ZLeyH9iThw
f1CwfgB1tBy2qGhdYM4X5Rfnw+JlvLR1UenaAgq0RH3BMWldYY6GhuuarEB1
tkAghnpkvMN6B1o0BgfNNOJFtENuWtq1BJP9tEvDxWRGQJ1zwWYPJ+RR7rAL
uljrFam9jf45w3wi25UxvWhoBcxH153nQH4WduU1vGb44y9IiBpSRnIPMXqL
cOqkbEOs+QqmaL/MJJDyFWnj9l/RNrRolVoa7apy0tQQ4sjmzjhzaviNrfmD
njRLHgJb0L0pL8LxFygnJcH68BzVQcZcW8qWMB3mgXLhtjIROYJKmHY/WFH0
KtUAADTQnQwAbhM3Wrs5/urMX6ATqvt3oBIzPVXa959J0MtpXwu8oW3IpePT
bB+Xovry+PtZ7VyKhPOl+S3W7JcHVs6QssUrYAKVGGKmDDa2rb0B5Num3Nfr
TyJmd7hMVUmzo3JOSZCWyc8qO6AWctrwjC/cCwmmF//y2fAAN+yr0vHL8Heq
D1+cj48EXS4aHbVHg1WKHCexvfKIQ5jQHiuOqbft4VBKau6pD9i6MRXj/4IE
DAd6pYepHLavvvs3NejXJg8QKK16WR2ZOj8n0gV+zIxbr+RZM8mplSaWHfC9
6nbeoHtc9njS9+Qd0dlfwo4VY6yzp4bWKfP/mbD2fJqql/9OqQtbUm5OBwlP
FAbDeyGgcaapAEvklkp5w4XSOBVdKVDPQw+D2TNqBmPTZ+7jItMAdlJ7Wrwk
jTVPGs9MOwO1B4zYcfr3GoWF7NvT6q0bWaLHGtebaOYfLZd+6PEtB3m1QBrk
XJvLvSOmabMVjR2NReVY6DDjnSpE+/a91TNf3g0Hw6GimwL/nKFQyBnucLe9
pA9xEuw/RVA0L9BdI2EYHWlzIRMnFpTVXvSemVJTbTfQKB5tIC1tkhjc9a9p
fpEBt2MOwSR5xwPZS5DnNcfYMpznXs5qf5Wo5JwJ4Xu/6cTSxqXAmx4aIjgN
DWNROu60iypBI54OFBrZhqALW6JsDkM2MFuxPUTkvut6MrP+4ARnsKrGQDu7
CiEBQaXAx8dIr4nr7xbSCQcozKRj7AvDB4xBkZBA/sVp0mwz/oeeG5wBP1nz
gyA2xnB4nK+MDf9NCy0nakNbOGvZ/T7ofy3JNx2vXdgLjJ603wyE1MuP5I+C
f5KjIZkSVsfM/ooDZxZqLpW+7RAHOdKQb/PhShKcj7/NRE/DXbNChQqI2peE
gj920XbPe2Ty4k1ZdMYKuulehmDr/xwG4ghErL6vCBabryrCL263NqpE1ffd
MBbu430w8VP4Jy5JTEcC2/ihDcw6P1vOsX02EVHMPXuoS/+cYr8ORUVT8R/A
BH12g0P35Sy5OinYxrvwAKrhQdHen7sQguWW/le7uuwBxs3L6IMEdS49IdB6
c2dxvj8vkG9DG2ym+AHg+qyJtB43FEcztnZOJ28Ah4Hv2kBWVZQj13HrjvRx
/ZiRKJFKTsVecpRiF7PJazYrgKNdo8AhtXJZ5kCW5S/RF5h60ZGhe1dGk57p
Mo/nrkD6lbJiRZgErQS8Xurhr3/pCRPFH8yZ2c0HlELuAN7ft9VRDzJtBR+q
+w+fivb2WqUylFE2/9ecyJtnC8DItoiJrKfuaWXtoxNZFBp7g8HEVd1lkjF9
v5vC2qi6fbWHo3fQS5FY9es0EEVQmMDtCHC0g2T9T+B0F5TmnScyQPM3WBQH
+Dq3shO3dJ72E1PDN09ciEnoplb3BlaPu/+bwezSKFbh6MMTiy18Hy0xeWyO
22cBjGBWevAcGC5VjA5VUoOcOUSEhnwGm/X9WbU01oM5JS9m2Ac01UhFQAat
+hWY8I/J3wRf7VF/8LpflVFww01mPtAgyFC+20vnZSg9J3eqTIk41nrXHFHE
Ft92HtiSG6/5n7O87IXCQCprspWmRxZPS8rULUlgoZasUQFgDUiZelreTKQO
RirzFlleQZN9DIZqilvDVsR+Qow/Ke8HSq8KMVF73aMqrWbXRLi+85wq5tNU
MTYgxaQH3Kuj2WjiRVGNypV4dcT6OxH/SIbI/2+mzicW4KLTLVfPpklPBCG+
040eGD3hxbGmBSc1q65iWJulNXs5esft9XwQWa1bh+xmnRdR8CGgYUhdUqW9
n3Jg5Dnsoc5x4acAA0KRbXuF5Ah4uGVvLl8GYCv3RGEc8fBbU1/qhJZcQ9r5
eRvLByyLvWpNpz2Ij8Yw89zIT0QKik27SonkJaoTWvplEQ56ehzsHD0kQRhY
BJJAl+AmhS0kYdrSc/7Wf89Da79bxNLRcWmV0EUBMjIzrTCdXdCVGOUcDZ2q
ku4rsdYwB8KxS1tql2vnDpL4NXP53+oObNqP9FPaaLw6nGYmfcARluqUbai7
Tw/lZNlVuUKFtWs19vGH1azjOLGPCa5OSJKirQabeD6C672B1LdkeC1aGp+6
nuihh55t3F/eK272JKbUHdwlSlb14DUNkv7vGDTcCiPg22akz3gXJiQyuGfl
Stv607VrRoPQbqd/e+JHl48aSQf1icv38Gud2vdglYLhHUOScadXC8mjXugy
q9ka/AGJG/N7ca69ix0l98ed5mXSLaDc1WJWdlWXp2LMdBImAJK9XhqRq1Kx
GBSS2QuHFaFiZd/vSvFNc8hKphSa1KKM6bDlTUiC4rElS91SOQcQ88JBWVbs
ORoWbEticnt5UpxAj7EVp/oRLmvA84O2lV1Vz6SHq3Q3ndm+i6yKGiIEldJl
4S0/qb7doKzW5z+Jwx8crXZZY0B8//o2EU090AMyftawyTKSHlNSFz702e0W
3kih40w3CCrNr0ozx2yYXXHZufGiZGK7etnEaUKHruKAvjNxqN7Dl2tSrCIe
KUA6t1NpgmB2daVQOwBsmujoVswLbUUdQYMDzrXLPUMulTTOLdLqj91WUF2z
JE76uzL4aZLZKLDSvx9BV1sSXkFGb9vIG2qyRrUFfbC76FgUKTDdBWD+0QYS
iPAsW4My8tXRbMI2kd00mKjiNUxFwQwLO0dcsZFa07DxmA2wp094biVPL3bC
fHHi/BkohWr2bHdokI33ES+lsNaYHzIkDUFt7emK8F0o2iO0Li4Dq6VAoiTy
Lnp7+/pPypnTmpiJGkj9ve2oN2eTl69Uqp3tsd38XxIMaueYos78+eGzGMjv
LvR8wp+/oGIG110GZts16mZJ7Q8DYW98kD4XSpTOYOx1bTDnIG1Prk+N74qM
w/v1FDscfgRBlrtSEJ65jvnOU4+2+C4pAj6hKxyIBvnyjKxsog2RG2ULXjyI
qI8BTOyTAG0uvDczwG3RBYG9phvY3C+gIrxQpuMvPvuzK7WlpOMHycadz5gL
yUFUnoCuqzbFNO4Kx+2Eu3lNGalzkAEbOqxDdKgr1ZcJpG+xTXG4RdS5RPRA
8z201nMfpUQFJhxDSBT8i4iFaM1Pf9uDyaaKlsmwMPJ3zuqGD9xtmBx+IiFW
G1FRJ8WZ2QYl3eTCswUU3jq9nf6J+w5HlGaCO4bAYqV4d8oawD8dsgOt06K0
jTjBacqoIva3LSUMQsAnEGxD/u3/HtOgYQhhcwn9IoWSpqxzpifqvu7q9OT/
AXG230BvPxoptyND/BeI/C56MHMJGrsbUUsaJIMKWGr0qkMthgGjCGpQQbQo
k1cx0KNAYzXYi1MLFLXKdQgwGGl2UukkstTn3yCeyKwgO1Wp1cW3GcNn7t6e
agsT0jBhN2Il8WT1J+5zVGHZjfg9Mcdta569PfGjHnYq0L0CWGr9YPTxiVQ2
MstoG7TllUL/23audAMhwrrJirCWPQnp/1s0hkcgUdR61L0VUcyQvjQz+X3l
g/YVQTeeNcxB7rqlymvdyqA+ifeHegJpZg0g3RgxjxKx8wPYh7McR3xfyFas
q0QAYeUa8z9i2YYd+i6UsPTMGi7LptVB4UE+Pr1lNVQ8GJgwssyu80D3AhVh
LHGdzodsc2T4IScSIEOd8lW5laXXvqqgU2kRGRkN2JUk9iC/JUttx8dnFeDH
D4Az+auA11fRNE+h5qapJK4uRGrwLJSb8tPzgMBJ+8VJKbqunWkgHSkqCRJ4
5IVsvjNxr2+bat7wR0+KExRdtFfktyvqq3lQv0kVOkhUfrlpBTToBRCsU6sU
XjO7Ret4nmq+kGxEYjTWrbVPaDsi/aGGC3mBXdW7+XlZAQk8i8CYdN3wZskG
0JPBVUH5FiObu+JjIj7gJsY0t33eirLbD1Qgq/+RPRqFEXIIB+ttxi57Qhgs
8w0xnPbueIOs1KQjlvokTunQIrBE32uwc4wehoYb1lwLW1+8bI4TUY2/hqXn
BG81FLyptu6+NosJFbVDzou/bHiKq6twuKdz+QG1sH8y5dJuqfyyjhjWEG/0
9FdhbMCJocL6U6X8soDZVJMrPHVx3GPbBn0NWHnbqPB4MsEq/95gUdLEugdg
iVXTDKlnvyC0jlGfT4HYmogPAAPkMRhOc2xDqj9vTb2Li5y1u61TWQ4QG9/c
cn7PRKG0/jry0xdEqEKfQIk0y43xDWbfg2JE9JzZmCgr7XoAQx4xIxRowhnk
xKJpbpNbH9OyfkpFbEYI1Q5kOuwvdHUIRGGVNHzU/fRYn1/qunL3J27bbEqX
drwf92BeLyBhP8k7DvdrcnnFAJ1HsyqGGOi76mpcGp65Ov3QJ16KcMqn6d43
xML94+gANMssx4tAwNUZLYDqleVBeGoEW+CrILHCHn/av8Cjy6QcYeGGUfav
Oj2Si12DrMKEOklyW/N/etrq+CO1/V+8eO8gf5SjBMBzDHFKn1etggr8Avwz
TaIZ4wZESvSRbIoK2FzmhqR2cWeOLpGfSkg15STF7JbNVtfkeWxHOmRF3HWZ
O7cFbG4iQGeHsCHhIhrEI9fDJfkYdyQelzd4BTJ+mEQCGSMD7reNbKFABOCG
mHgcc63R/I889doz2AFDHOILQqUbdO26582hvB/2ONujjVe5uAvFuAkkVlSz
g0Y3jmProx4eQOAVi142Ye85lpG0a+d6BbPrJzPbqc2IfBKQgHKLzT1cR2CK
DYpZoJFSrN7nHLGnFArq9pvy6eUp35P5KUU449rz4Pip40M7JcjqQgeQ4uyV
SyORlcRIS4yly108M1JfzA1NpfsyU26jTn2C9fSzYc/X7tr2K1O6vpT7XlJI
9YgRAO+ZKZjCpubkGtcZUqX2vhqqx+WluNOW96dsxPC0T5q4kiSdKKC2Fyo/
1Py7Wq+tz29QqoYPR+8J4OhuN1/zQCYeoFIzGKkzeGtk0r4a+y6fchTEqVUA
uApA7iloX0knka9gFkp39pDpuNr2rZljIbN0byqTXo5u+f3ay7AuHyfWzhzq
+0prHWQTAphi2g//fR3YPJEydR9j9FIDoGqWmyVD416nISymaT2A6TSC8Nac
lDrNRnhnyhTWAQJLKjbdJmMcwWXFa11yfRXIU5FY988hwUa+U7k+74w/z6Q0
QCWrWTShmtEe4s+z4MJd/3kK/YYlxUroRXEKI+PG6fOROGBXNa49MUM772fq
qoDn464CszbvKkX12EaSPbss6RMfq9E75giaPLKZgY/w7KizqQp4lKxENZ9/
eQpmO1572QhRqeEbVubjtBBg28yNtiMCMUDsx35gAgErL2u7aleGN/rW4bSl
xTq2pPdLlz4O5I53jSqgLol3YrXj22jZAIgowaum9xoon8rvlPhjDta5J5rA
CXTXb++j7SlZOjn4YudGzC8keO+lqGbyVXKESCjnqwYV+6qOi+oov+5h09hl
vOf8w7Q5hbBHC03v5ugvjHWsrr6OuMw6IjjSC8YzDSisi+ItmNORDFbbs/Ff
1dJ5OpjnDV7aq27zhFzhgLWIKJrv6XxsWbGoHzhgcfwZfWQbAjDluk6xF/Le
Fp7R2aUPIha+Y+AomtU3eN85StvzlYAbb4WbQJProuqwFad2rttNOEsSkqFF
ckDWY4Ot+/3ByUIsFMcUgslNtWjr9oRFLJvzawc9Y2qbGhzfOnEpAoLlbCJS
mBTzl3+uHhJudYVDgBO1vm0nxCpWItypXjE5VaapZZl9EKFoXdzs+egyV+AD
xD+pdb/rFWJRt0dnY36kYXZwR8aFUJorPknytBlb2lFwEvbBULfxAyykji+Y
Z7C8YZMaqDQ+E1W/+U3Co1aUnDyj+xp0BuApNnoem0SOMpPX8ML88D8GT7nG
TV6QglYKxW1tLHbcPkKQ3fUHFrLwWvgu1PppAltjq/dGAPF7HRmS+e3vTvFy
YYT5ihe8YkNxHDMytTu0dO+tOCSKzK40GDvJ8KHmyQrPAAwPLdEK8MrfsjR7
gWlpRpggJT7/HefBY2235KVluADonTm/HT/q2a6+mj7K6Tyf+ln7lXcf2h8x
tnfDaAVI55j0tRm2cwMtqsC+hT/s73fLMElPTE2VRGjELJUcsXsV9RKL8WIL
+CfxY3A3hs/7x47eJcTYqDFTry9FGxtMSdSiQNcakA37A5Vdou0Kly8p2CYq
TjdiWD6YXWttBgnac8muUhd2RrcSZFz+TKZevzYaLMe+JFswQWeYrUaa1ftw
jojS1AMIO3mclmqsPPfmuANPle5ah3rUsQxT9d7XOViHIlTGz7XTViCK35fg
+SnbjwA4+9AmokTnisywAvrIK0gcgOd+8l1Gpe/ec918m1yvoQaPsBKR/254
qghAF/oRo/8gIqbFpGhmycgi/kUmWVQPpexRpyt4s+Nxg5Jw3Wry3TjfdEP1
5jgQjhz0iUbAowwYkHGa/rOzi32y4pBYCcA4B2aFviWAJOfrQRgJ/H8Y/tmQ
JLz45Ube54kABshonYNnBq7AIk9QaUqRfzL2N2I8GG4cNtUv4jT6QaNoWStx
Mv/wK2SLV8afnltcsgkn2Ha26Ngn0Gb5YGecNU9chJ3CCb6VK9gDP/8a9dm9
d7zhCgGWoMNTim9ag30WasLOhE7T9dvxw8nyIKKlAyBNdbST2pSC5Gs6L+VD
TUynMf3J92ZxjRZl2UuAQd5Eimmiq/1h16RrzBNHW5JFRsJMU5t4JthCkemM
mdXj9YmzXuNsxbknIXdKouMR8E5pRCr1xLTfjS2sD0WAodxy2ksvjpORO9r0
II8GuYVKPpO+3xJkysgDAUFecfdgMIBUg4/dyJ2sxX8ImjITQrK9kQSvJrCF
lCZbIRRLbbrstxgOcZEIxfrqAWY4qlaG53V8dky5MaiiDq/+zmPsVziDI3Lf
8RZ1QpRs4jVIEuK0U+fqBU5oQshB7vompXKEES60fatenHSNwS5Et/zFtZ+G
74hir4Q2/UNli4cJnjXg2qWKWIVctla1Yr/Ww0jxE4X8lzIzcFINTXHuvd1g
TYCfG9OoIs9CX8BfQFtB6xwXcJkJyiXGH2BM4cs/JGTQPFKfdSYQjkT5aANo
0zo8TlasgBtEyLCeVs+weS4dk0Z6U4Gs9o2bRcmPvQDTJbGkhq83zdYckOLj
//6JABsMMyYUSKS7ibqSHwWLsbJUYee9sq/1yjH3IVa4FzCpD2tMF47gPAmU
Rpfw0enYDjbgJP7gMgAX4Kpm2fuLrO7Xo6iF350bnnyzZFW4jfqp90Prqj/S
1DpyQSrPsGBjFXzOasKNLmqhh4mUvfsgQ43jlmWx5DB8SfbAAWdkJRVa4RDp
OrcZptwvu/sXXZQercaOviDKlQCpq+fMsfG47gewQ0gvUxugjUtoRtf44Gjl
GdKmnX59GccdFsGrddCEtQuzphKhQMNB6mIx5PYTcvZgrE6lE5kJ6HzBVtst
2kWLnPevIjRxrEtnVjMvR2r+CCcsRlY2/VCsoxyxoFhVx/P/oodZPwD4nA2Q
C82GDiTNztZjcPQPWSFVBbICKFyYIhohNVso1VJgDGBQYF925VTTr1kh3tRF
0zWrBJTPIvq4k3CLoZNyHYgKv4eL2dOwsGC4dANQaI8a6maLHLJBPFUHCXYC
FWH9LHiyYBMg+wCn0T68jEMRK4RlVLA+6ZkE9y0c5oEpP/704pDGAX88H/EO
1N/4fzpV/nxpKqJKQeg+OIlN6zaezpoTPEO6bei1FU0+vSGnWkQEGNcGX4EP
sdMBmX473awtx33XpJYHj55MYUdXUEC3jK34KI+FwfVmsgIQnQKK6/FJ0NYz
h1q58FD//1mjwmEA+aoqnVz+9e5w9kVqtcXigkRkEzrZf2q2GG4cqWWbvrKc
oBF3X8qcrEfIcXsdFCINXlxkE8kFtyETKxx6gh563kd5BD+PXRHMTKg/ZZxH
yVYSi+JXbJ5e6YzrcT46QB22lu72p+zaTaax+TOjcOXHIN5yvEM5LoscyHG2
L/69pO/uApuDvD8OiSd4GxZ/NWQRbsdKGOfGZw0aGqKWU1lJ4XCPie9Pyq8z
DGrN9w1HUfHNZDTOfklQou9HaN/DRcTgL7ojNF6EbgUrZ0XKCZGJw4KRIXuN
7QtpblhLFyD/960oaMqXnl7CFyOdgkS8bdhzqXLsIskBrkmd/fIN7lbjeEOc
2YHr/xhfoUqfxaJIYvCuDREczhwWHd3Ah9Zk9DKrhhwLTyj4LP7SVq7ZhYSC
HebEGUwr7XhDZX0LV8GsXvwYF9MdWQmrSrfqBfopda4kUjq33JSfRs3D8W5x
JLclxAw3afQpHJlcMOH/j1AbIkF8dzv8pCcl9kE2Wttuwug3lntHNAdbWOni
A5XgDKMv2hJJwYUPV/215jqQIsaYsBtJ6btubWCBXSrEvIMNv0HFgdqTPlBo
/RJV+Pvk9PYNmfZ84JgPF2siFsW4z3m/huyERgcmfDcpoA2Q7t4ap0QBHzF3
p3Fs2z6VON4bdcefkRp7mFde8Jgu++2g6qXlgF07RJ+LBlIpORrxQEjOeN1W
+VbmR+3Gh5Ig2G4X6DRxiOMYS7UBR7b0XhgcBKVs4zRuQAtPl7l5o2vGwEdH
VBCw3hqDfQUiOWAjxVta+dgQ8dQr+Kdqd3iUl6Hk0g5mqj6Q0A0TdcLmEaTA
9xKIGbYxAaulk3drxTYQv4d3TGqhc3zDWTywjFG5b35XyxBCiVsQc54QKkte
ujzOjXS7t8cH1aGASsfWvwCanwwTkIL95nmvGipxlAnaQrUdWS2041q2QB3J
qksQBNGWXW2Nnhc/cViTpJQsw/bw0VKbSQidHmEF7RvsxVVPsW37U5JJDBOZ
1gHmppiHTwev0TUS8fN2a6tgFBywz344ymhpktyAS4HqLPQZWhXEUqLtEgyt
QqsAJ0pHeOx8TRIpbqo2X8D/hEUEFWtakoeb3jkCoeSVELAIFYZVx5nVazio
fVIc+v9eozxsiDJp0ZNPGUeSHvJ2XCYOIsKD5aca6HM4gVOc3XFcA93UaTYe
CFtSdbqbhxkHNyVcp5LoQ9AZZvPOOBh8xxA9P/z0eIarmMdjrp7khxpprbMo
G1Lq4Yyq4peRvt2SoZElXn2EaHSUf97O0+F8hKXFePrJiQkkUBW1PnEqsxqh
YXYkW66Gxt7LQLC9ErlhBtrYMKNP39xgvwDhK8Z+n8czULejo68AG16cbuNb
mutiFd1LkNzpjjoEjeo38yxyNzBT/mn/ZMFj0Lazr/kUZUQjJg/Qsn7TQLyr
qRMgcla4lpaB62PLDivGPFnxn/s1X9D6V1lvOHYDIz0WdkOLVar2YfSVTWuS
xG/TR+QGEepTe7azZnomJ2LHmlKZJCEiqeq2a42Vr8cvkVjOEjlzQcF67fgn
zuqRAlHbZDv1CVSBoBG0Mbt+rq3mWhyB+5Cxw6RUSGPzf5CDSUjvLWbGDyOf
jFJEzzl2bhkwlq5FgQJvDXfMoA0YwOCIt5ik5m93/dKgL0jcsMrTaPiidEdM
7JNb2xbMgwZknyKlssPFY1KHmmzRwbjyUIYq+SPkz0UPLPTZEZ3uCtbBHX4X
76S0POEKS8pjTHkElX2BaMSAUJFvNukA+v5PRwgDuV+wRac6SYAo2I/WO+8H
u+64DvVG32+dRxNaFeQIhzU1R5LVn830QLxQAMzqAGZ4Mpc16gwBNgzOJ63D
w9wrtTROctDdq802Vn+dYLzcTtHa44sV2SVuB4mR/d9TkSWsYk1Z7ueMvWZ6
TxpNoXXv72HdmlzuS2G8WT+4A90cFJH72PVziCVyUeFP33354A743/0OjU1M
77UfhBGIMZAajt+ljaFM2XKv9Vu9eioKaaHjkKdAfFNhM3ndteyBc4kpxtvi
QYdNVhMTKeoiLOxKZWMJ0OiTQ3jbckSXUakM5wMWJwLr10OSgg3hw45Bwign
amZGTh+zysu6Jq6ZCrdow7d9YkBQkQJwYmjaPuKF2Sc7YiqTIPmL9/NREJ5P
YoHEYx6urgl0xL52WVQ9wpMhuBnCNAOlLseGmEeMi/dhAb6zSlaZjsB6JPO6
nfXTEMFTErF5XJ/m4UyoWi7IyKq1ygZfhsdqxkv75iNqjguhFOccEHbIBck2
yHuiRv5CxxKFo2dJhmlpGmhpgb+ooz+kZQm1O4jfTzx7bUT6q2tRx0ZPblya
nBmmxaLiEoDqbN/nQBPPX8R68uxL60+MNMdcmnD8tc4wgIrrMYTjuPRXrR+7
2JOUak4oaN/aPekgHL1t4O3tgNGtPD8yRBR8ajHHrhb7Rqa4dLVx+wTq9CFi
N49qH5MwN2NuQMb/on08XKD6TBFfCr1+1cWnMZLcDbTd7L85fbhwD6hLYYo3
zs8Z5WcX1Gc32JTW1+SZvRA9bvopM0jmedJHB944FRGNBHfwfYvAJ59oRufM
YOZl3ExW1Mv149xXZXhQq+YfUZ6rEbSusKphoNBFvgqjcFzSj3bjUq7yX99h
KBby1E5mGMt3szCBGk0Vxy1M6VDiesVfqgMyuvnTT2wLuF/MXvcxS4ZEj/kK
j9G8sFxkVeMmhk1hHOLoayxKjvXndtoY8+a50+zB8R1o2tHm8fSEi03p7RiO
6WouJ1EeHJqru1k4O2UAjCpYj7SWiDEaZZ778Js543O9IHiObuwThQGTCDz9
Dd6vDD+P5g+VMRxTzJJAQ2938sovaQRTwWYZaNZBDw83hZJbWRvBxN/ixsbx
awbO8OYE43zsL5VbWL7oEGOHsmwvFwqjJ+hQamd99BbTMvyHLd8GOdRjJT2d
k+AmLVi2DwUc5Gr+2vERoS3kUWLWw1uhYqEb3hlT/nUVfr3T/A4gWM5wiTcW
lWnB3LznSEDqMhC0p6XEykJPWe8+NQfOD4eKZpZ+NuLPojYNBRP521ywDQTj
+l9b07FvYfdCkENgP0Hp8CisfxrQ+27IvMahpJeqDjAJdcErRp2uz/sJUWlT
8CkDTqeUwnJ7JAPsnIYh+79dp448Ikll6m0kpyTcHKty/694fcIKGrG86Ri5
t6lhpw4EY+Ky+fn/5bBObKGXTgAyMJ2fYZA6qtrBrbWw5AsLGRbcwWkyV3fg
kUc20/rpqIg2y7JyCIpK6GZnhoAEZRaTvJSm2x7yNLYtgXyfyefj58XKBZFO
DV63B4wqlc7ZDVotvnLhlZ2scBkmi24ryS9Rnam+QDyNI/e9ZgIxIZkrq9GM
GDSSEJ+Sz5SC+9zORlBzMzHkGxvkmvWVhdmDH/CDxBgyXumjpkpA/4wEuIir
8VDp5I1Ivkv9gcM1t8HmupbCL1EOMeYDY156aSapZmCCT0+PGh8isQRkITvm
tzvO+VywZOwvwII3PRnb4KYgdc57fVGZgGSRlahvmlpgLslGuiXp06gm5BTy
rrAZn3CtLgrZN1+bKONlW4EbejXrs0hNRLDmSLodX/D41AmDHexYpMm6LnX6
gapAyliSiPNCJHgn1b6CJ1CQJ5skII8pUgLI/TSZuZKBgpMiFzR1SZKaDTDQ
B3S4AKv3AFcUayY7o7gevdWQ2bLHuhSbdLg3ymDJ91i4+qcb/65ykDksJOdb
zxUwMYkNUhMCGFgcu17jqUhubxF0uoC0QGof/L/+/FGs4SJJLquNdwy8r2Du
XSIgBQqv4KvWRQ8T4FPnPuC70rBNGDo7PIEKKwKxEzbftsiArPX7lM189hHd
EYRm4jLY/FgirhbHJIJDeM8/oe5ZlkruaUC8ihVrKLmtKMbnLfnnfWP2f7Jj
8xI0Zk0oSbaoGMrAGvgHuTxODTGQBs9R/Mnzsc0imqr/XTb8+0wgzjE2pbpx
1TX4oE/PYGQm5jSKHYUZ0dBdlks3r1veXpLl8gIXIfoDXbxLtxHtSCb4dGzd
ozVdeeLSZHQt1wAUqagq4Xhd+91dpoSvg/OhRn52OZ+se49Ly3Si8xIix59A
lECWdH0sjTFXzbwOFQvt0/IM0KuKfQdvNV9Fzk7vwt/TZk2wZDE2n0YNX9fg
HPYqQNYxB/JaYYqls/4ElJqOm06gcuVkAA5ZkPybIEo6Ss6b9d/9EOW4vWlN
GxGdLLWr9qb0W2GpZ+ESdsE+6hulZM/HktsTb1VvIYqqnc9kBEdYLgLDIDoQ
QJElTz5r0IHeRZc135HpNkmUkKoubIYJtCONV5ibc9fHNGGbn8iD0hTAp8WM
xmFOoZbgvhCpRPiSxnLjKFJ6qUCnDsYkwJGjYi2SjlhreXbqYMSM9saMMG9o
EyB6NsYHQCAzamkANaLDrXBtW/xglhl8tS0jQ0cI1bvdoVRwo+Q+Oh4TcKMZ
muTa52OIyvEpMSf6jsmW152mx1wmbTRwNiEU7RqaBi+7Y7LZljht/AGUxnzY
9ceQ1l1dZvJRQSbsCeMOZb3TaIonqjhuzKuDPSjJwAYwFyZ6FP6/dtbr0sDz
XhInVl8aWVYalWdgsmTQLlR0Ai6HyCdmuZFvH8cDbyWON+BGITbgbzKnB+HW
JLJQ0B4ZOTirVC0xUdoN5artMRbjuaNLA7wQukA+DwQZ1SDI1sJqYPydL7Dl
pj9JglZKlUgJjoDx7d/A2HXBeD6/AFAeq1mD2DbvjI35tLReG89XBZr75+BQ
uFdNO315d65jmmZd5BFN0DFFtJAlBDGGfCpI9LFQzBiiFvKlzvqun/yzMVPM
VkXLjYL1Y3+DE9NYUYsHmenSN3LLIuYl8S9pN7MmwCKCs5dsT65kqXpyM9qd
dh0jJ91lUSHiLei8IoMaXvHocDlw7+QAA71mlohHsdHyvqs+rxkq96Mxcqo5
8DHmYYxlK4wouiZdt5/ptyWOVGaqlsOJ1SrqrnpyB/hDrD/sOc1iuksxqciX
PRjCXZsl4xoRjP3R/kNzOeUnmkFUwEiRFOPu7XGdmrXsn1Flv1arTYw8pYxb
LdJ5gr9QoqJM4isL4vlVPMpJiQ3GZ/y3GpTin2q8/gb43Qeo0WRnQ5zvDeCa
/z+ooxiVkf4vuohTMaUxXidxno7mMrep7DlJ3wPc94DhFfzTeg4WHmjCtXSU
CCkYVVdEqTfEF210nmJKJi/BzN1u72M+77KZ4dghsERXakCpYktRNGAJsNG8
OqyOwcRkfwsRE7coMDstU0YHdpiwCZ/crC8Oxq14LL6freRDjUenW3DoVa5G
ZPTICsUNwXg3e1lMIvaBf6dRvzyes53ptKKO4z3u/m3QYkSLz7CEG8o3RoNS
+1EW/hqWOadWEOLPE45PcTc3Ce0fe3fsZHHF6rp2nnWwFinVnpN/AypFuQqP
XQmefM9tvNUFwPazJJtkzKgU+9nDDKwhK0AkvD3d7m+mTTkhsDNUVvtyfPy4
iw/795lj2oGf+a9ExeyJG5/aTBBt7KL14aek5BojnPomCNmJorhLZVFt+Ilk
otC1P9+QoCXodwsS2dwgfwxzfdJYQN1JnxqxF7vKxr7rn5aBgrRr/qLxnDwx
mg75lII8IlU3h+y1XK79KDkQieltVqXWWBckPf3e7M1JgyvGxDRzZ4lJLMYv
uU68th624emuWYopoliBbrK1GWnOaj7P+rVKixctQKn0vtr9udnjdp3k1Cjn
I8P0OiPfyayXPyWaSb5oyRqKCOXcL836dvdgWx/dLQFRvXJ1YCoXiypT18Lw
YeAy7mwLw1Xtjl98fhzjMLOUR2rI80PLefexRq8bDH/U5zK/xInE7LS+xq5d
h+JlsCHT0KcpH7Or2w2ToYFh9R7bevToXLI1UsKRX3QUc+5ue0cEYfsP6Y0B
r8UZXP93r5UI8AbyS8ZwCvWMcMKHGBkU3PL20ltrzPxQzgX3d7AWmmrRDXFw
D6QySbazMTuT8+ZnDKS1jgJoteI4PpqjVL9fwHR4nwSpWSYe+MzJGqI0bswc
1fRS2N1mAp4J0aQAnI5BcJ6GlMVvsmXMQ2VQmE++JYmA4lIccBrkyKm9To2X
Fo3CFdEaw+Mxc1CQtUkDnj11GihTaABVLkodoqA9k7b/4vwykug8uGsK682j
qnKIA0Cyfuc03+em10gKDgbN579oTLUleZLGyu7Wu+ifzts0o5s8WRx3A7BT
uigDz6LNfMblDZZkqeEQ3qqKFNVa0x0YemE5VXW68+0zGWG7d+aFFEO5/PHc
IDz8IoVbSCvNPfrPlE9Fu72gLjLr9kECV+4KPX+G7JZSYUb7n+gW6V3BVAAq
r5e0Bn6Hhn9fjSFnTwn+wVzx32ZDmI6mQC6xYu7yKC5CpfHpcbiaLtpVQ2Wx
Qi+c2SZxXhNHRxndEQtoPBSR+9A4g8QQVsc2j7dVs5IgRwfcorfMh7fyhctJ
o0LvtciY7G1JeLGCAtWEDgKgMsz6bH5tb1YPq9TTUCEmfjXwONWi1OgBclha
JWMIt/e3Tx+6t8Kn7ViWPtOh5VnFFjuOt7GUcv2irK4buASmcpsjb+zRbTit
FFaGARuWrIVP8Z2VLh4wuN0sSDYPs0eelVIGUJ118CueY9v16/EBBGaXLpzY
dZT4dxXDvHPlDE1TPPJnnGjB+XyAhELM7gtOvu+EUnzAf2r/ksbz583ZGYyR
5iTIE4nmNsa09kmGlQYU/sTiotM5k+IzctK7nk9FcpkFvMqlKDn8buKv+Xs/
sqj/j4xLz4mj10DuCBF70polzf1RGHW5D8DieKZOruWg3eYWS/9FRHLg6W64
UFlys/cDVmNt20MCwcTdRXgtYTKg7rtl4k8ZggArOCOs7gmnPSURFBWbcDji
BcDiaWu04F+cqFOJxqFH4uC++BuFylyvfMyvsNIpCmugFxlUEKsTG58u/2Jn
WzfhtGXwzfjlKjHwO3J6U2SVX5v+lgXJtbZzSgoaKUoZZt0QiwBJsOUpUbYX
pAEtVUxuVrK3I+X/k786DyNfGuBA3f6fg5m6ulVEwFxgCA/7ozmhW73QCyqW
JyrVR4BnI8W2UkjazWIqJzLcBZjm2XYBxtB4eNIl327jrfo9yhGJrlODwbw5
hazJZVPFTCCcATpHrLtVWGzx/z31CUApIoR4DfYke8smmlwVtDlQCX0xV4l9
Lnf6k6OUxo0O3a/v4TzYzhwh3My71raHcACZqzwyF4GfT7FphyVVqI+JjHhW
xrdQW53dq/D2Io6h2kKkBCWBdYgbUcBj0SmOnS5BAF66L2I208Ds5WBT/jO6
QdCTga9YpzPhPuP6ZuHtSuFkwp5SuDksjCyWIgVgfMjJL2n396KwNvZ71AoT
REwQtQxKHjbxMj4xN2scx/DFuqCua6pIGeaxA5Ux6OLe1TAdSg6c9BS+Yvwv
QOhVUz+/Zz2zqzqtjSJnWp8bKRiljg5SjlQx9c6qXrn4A4y/yq2HfNHx4hP5
SBQh1egM7+adhPMY2NqwlxkdoMN8QJAe0YSZkza4h22E+pmNHIOAlIJsqSzM
0/ON1Nl4k6Hool3DcWdCQRR0pTfu4W+WvO1RRkeC61DYIkzQyj4Gis9iXzp3
YmMYXlDU507DBxXdFkLqBHJcJWNjnZqmEylRs8ujaM9rTLRpY6Z9FVk8CVDK
SeOZMlZMot5IG8pGtqIF8xnMKeXePu32G3OvnjFN90dAYpzl31sLND4cu4Me
L9zDuRLyNyaHGjbJy6noBm2pSVmNlRCrOqchR1QdSLNl83stozmvLg1KUDYV
tv8PmISPF174QeJ1Cp1uI7rvnDhr+s06mcP+sdHi+a84voijuospDdJOFvM0
We2xEO5PZG5+AjfqqR8VE3sZJ4UEXEp2OoI8YMOJQgQws6OZvbzFdG12fLm6
+yH4/E4IoizgZ2HWcdLPxbCU90PDVNVFp8ybhchMGsj7JjYk9Ct9EHI5ahEH
ZBjN5mE4Ya16bkIDA/FTcpvxThp1096g79NuGAcOAfc7LOTxWv8/4Ywa2f7Z
e+JRPKl2AqdUy+nj+4gffu4kc9FlzNazD4Y5SnqJmsZvhNKW5CF216lC8LVh
FYXeukLXXrCYkfCoeTq2PFwKSCWAijNoYYoxBoLOYlSdwmN6yTdr88BWrvej
9TzNel40p10p2skMjSYmjCL/E7UDnINlIyxkB8ZDKooh3UlSLlCeVN/EMjJ7
AhYm3jinoTcs5ifczhi+23DaV+P+2X5nnJZ1/aW/72XhyWSW1auIWqEGLWTd
BJklXZCpmnhOUD+Vylz6BfHPUAmuRotUw2JZe1a8fzCvKNkAWape/5f0qJ2I
S/62U5OCbHK/xWVjwHTUSggQRcnRPCdXV6/NT3vC8jU5zNBcQBb/JTb3WeRK
T41y1s4VEPeZJBSo48yE6Ut95WaQnENUWxGVUpIV3Jff3SMRrHyukQ7QwegK
XDeJ4D6cbg7IDh3ZUJMDmDI0iKhHUA6t8s79IWNz30sFbY8M5K8Xi2kcwqZd
u1FZ8nmz2CCDzW3uoAqWhne76Db3rUD052tIlMhcP4IoPprRnkV/o81gkduj
GuJSm/Z+KHLagGQ07TtRiEe8WA9hQQV3efJUjCd4INvquUIadcvcsOueFgBc
QnywN2jJ6FIAMdyySRZHMHG/rkKoquD32xD8aeztMsVT6Xt6KZBeGLg5QsUs
ZE5cuU/xjXza6b1CifQ8qPnaPAQ1+MH8BMEjudCmU6hSUdL6u02efsBfKGEN
cROxtVHkT0YBlcXd8Sub9N/H0/MLLbZ3ALU7cEwdYzpQJ77A9qUQiqKvOYe/
sxmh/xhXeN+du0xsjzqqzCdqdvUrhobZfuHCsWShTIRkGUnNAwPUX50cgpBb
XsSXWAunrbIPfqUbqMWdJ5AcKjkfGeJU4lA0yEkTA5V327aojCWcSJEwXpBG
eojl3q74U3jBqDxyY38OzlPhlVs12iCo4BMyVEksxnXb2ToaLYYG40fZAwsp
DDXQDTxh2VeHoTS52K7PdvVyeW1YXtIrhOyYWJoJWaNaY3w9311ZVynb6eeI
h9xZm/WmatDhlKi15U4uJ/Icln9MrQoh/HcDI2VTp7A0euvBlIfvWFCZQqM6
ckfQWszqve4leet5ZQ4rttVnyYAUdwEFuoZBAiuXGJk3nZx7OzXepjtBJs9I
opCnv/LDVx6rIpJ1c+wljV2sCPTlKb0e+RH1nU+gYUxu31A5LaGmO0kH1pZh
Syc37sY1HESlwBDH3m2YFEKUhQmxgTopsVzVmmdHB8+vd61bz3jXW7VRJLER
82JQPZ/6RmAWSj812ARG0PMzIuqf1qHTSUWvJgvw3M8IemGSdGzkjLZampYT
neabaRKWjjE3AXUJUwGcyuZu3nOREWxgaWOlg8vUMx4mPlwkMJqry9Z6OS7m
J4FDCsV3fevRxhrMuOvWl//wmC9nrSz1Xb9tkD1WaToaQESZjcqAP16PFKmS
zYiYilnDLab7Eg5d7M1hgNok/1zmj+n2vCMMIWQZrq8lJMshnr6M3zykCA8B
oMsXZ5Sp65xXp6Sr5wt7wzcwNVfS/opVWbrG8SUFTHANs5zPo7VWogg901Ti
m9ZYqdFBZYPMGJ8MgcBAYx0Duk0u5oVk1uBx7E37ClB9Z5rT4yd4hclf3vA7
KcIxdePhwuHJBEy8Snm4FL2plH6za7Yo64UopZ6NH6t9JS+hOpAUbmjt9fxd
S4eOdufdWnJLSe+caqWcgNV8BBM+KeHdNpYZME0kcO9PlbmSp6AevKk/LPzm
yy3B8kpVDAk8sUymcSqucMNKRkbyueGhYUHS2Hln7rBjF03s2VkVmS036Kl6
CrNxtyTDW6Kyg+Iom7NUlE7qcHmHRRcNAckW6b8wBBcRqMCxB0M41j7Vp1Mo
lznfovw0nCs7qk/LEZwBiYoTthNeR1vK5terwVVXnFP7nKHArqS5nyxxM6tz
dgLrilqlgj3o8SHUGqDtKiiu7H+QW1DKyeg21nSE9NpeormZmbFuxy62V5rP
/ZaUFuFfEj0ZJCuBLdsy8e0rASa3tgf9cffUl2E15884BMuURMzNDySPLwGL
55RQ8hR7/UOhcRJDtgYL65lOlzmDx45XJU0DFNDkrriP+VtW+lOb7C7U2Rfh
vatUoOWzjUr8bHa6NcDkp0/A9Dga46QclAHT1P9X1/x9dUVra3y7Hs9ftO1b
RFzKoJy3snwRgWR6ywuTVOqUF1JOpJQg6QgBVh/isLLYgcBESOlMiLkLpJBM
lsYlUHu3N8ir4L3modOpJUIK1BYoKR1qKSLO8iNdF15Fw/vXjdxMblbqsHOj
ejSyVJZ6QGL8oM2FYlXHtBeo91dIoHx0boHG/IzaGIWlweg/cQ4p5/0H1U1k
ErkVtcMsU/VIOiD9xlW/iqmjUt/clc3PHMuWY9CAAv256s7HJgC3FMkF8jDf
BAVEkVtYSyLFhE+BWyo8DidFhLMMmswmrhpTJHmwHQeTYYTjIaBWanI14g++
L9OyBsPDqQXHum4YlVBFDp8wmZ6AVAtKmB6L+yV52LovUFiw8ILBCGWU0UNn
/MznAOqOIqAc933aMh/UoH0mDuHIGtawO2YzKPMnAFXz5nZ5tJpKKKWhW5St
ae16/oKkw6wfcp08KvDsKidbiGEgFERE8sfrnDcMtRzOsPTEMnsUPDgokyys
e9ETW864YOgb8chdiTIjZOwOU2TrQbfm+o+68ZEWygEPhGr4UX1ZmAQ0AtTv
v5pofEiy7CUjzAgGfpDh6b9UFVoPYoFHTeZMginNKpz5Yl7lqlmd+TAELOlu
b8daNUqDYJZCB0b+9RjBFI5N8+gwnS8VYKeiU4zb3nUAapxvBYab5KsO/n6z
6sn8IkKhrK6CT+nrEIDhVTFyn2K5ZskngUvRiV2UErfI5xkKV2w14DnK5LHV
xuClv/OYpS6VFYSIBk3tCFQZ2q0FezWF7LGNBgpWCfGfHkkQn1HZzEgi3S+V
Bdyh6cmG1vZNUccKIXdY+a4s2W+S9XMMJrE/Ct2OqSCzIW8RvnA3oNAtlsrq
LrAmlrM5LAKgaOJD5JFg0g1FhRkO5k6eoYN9slKCm1vvzdNgYf0AHoEc4wx7
bcIjsmU415NYKHAJK7rdQb5ubfIIli7Cd8zgLybNrXA3LoJoDatBdMtPuXwv
1D0e0UVL/1buKMge3JmNLegW19wlspIy+1TFpnmacqWJS2Dh4m3B0LqEfrFw
dv/Mo5frVV3ziyg9ZAJjZgMQ2IhXRTFt/G9zXg8dpDdIm3R+CB5oDh3ZJCVR
jgrEpRixZ8SQgOVqTBoPTyDGS/9yDBWDnNjc7odJ87kCZhbB6DO8CIgoGWGG
F3qtNjW6hi2YkX9ZI2bqy+KXixl2dbmEeCEvllK8LE+8ZUM2dQIjUU7Chr/x
xUT+MMuL0zoorANBKMEIhe5uYq7kOjrkfCTzg74xblk4ngoUSgcb+r3rmapE
iOvUXWiB3TTwZ3HrL0A2gwxymv3neOQuMC4HAbt4O1VgobIEfHfitVBO2tex
Tl6kJEfb/+v7F0T1FjIwoqzMMBxFZhnnkbC4keBp+qwRng/cD5oMuQsnUfwl
ZxJ5Ior/S5a8uFo4nKorERvJdVecVxWkdi5dl5+y5zljuUcK9FpaqNoyhjl3
Fes5bQ7l4zxXmEBniw7Kk9fTQzSkyp+09EUN1PslEgOWyD+eAZKlfNDPUI2O
aGAiapcqqt54GoXogopQJQcShi0o55eSaFAw5cfNvKaFdTLeemPfpeUxUfa8
ZkyFKzvTVPZRAxU+oPfrk42yftyCor4iBWi0NJHwOrmvSZtNRWVamF4yTSNM
fJKhXH23ahI89Lj3ZwkWRHWn+IhKAfrz0SB0Usu8CJbPA4PiPGKOqAdsNM4C
rPfkEXhXFLalA0P6MDSezcTnw8cy3qTc3C2+mNZYEUpFx2bJykO27ZTwc8Sy
qK9RaaFKYFbpszPpLUz/OKXPifSjAnnPZN4EzrN++QarXOAS6trGhUf5sRJ8
ZHw47AZ+2B+Odz8+2BadHuzo7Dh7DasWy8xUPr6tSlLsyFdG6Wk7hwrgU6tT
ERGQFlRk9ed+DBMgCYbrwoNwIwi0zHooEq8JkRIJMqTtdkCwLw/CXSiCo/3K
e91UOS65AzJAjNecrpv0CV9ZcUIzAW/yEdyYKPRf/NE0DCPTwe96+f2F6/CD
AOgjvL6XCKuWV+CiLvEo5UjM59NF8URXWN5sc3SU1M9As2PZIMu0rnD5oVrK
h+734z3J0VispwAvf+L4jGbTvhs/zzM9JQ05NnJ5djPxTK+rpwF6MMauhkY+
n6tHciEnmRT/TrSzpx/H445N9Gqhy9DCtUrccaFn62QU+6FlTCvqeLyXRh6c
R6GgYyy8YdxQVlBO+zJa+//1dXd9sAdAn/WJBwhzJiFRmWLxOqDpwBbOhso4
mgJR0ynG7x/F9iCvAvGCvYtCDXM6vTB4CgZncP9oNCewhoz9dkA9QtZwU4rB
sQYYnl7kViiW8sEpvTEbCZWz0L/X0IrqiBAI8sRx6ltU8sUYr0sqeuMwbyxz
8JVtybhxqGGYAHkkre/AfaGCY5AVvC7V2G9aiE7xMQK5pj0dATDPeaDz+Ub/
V74qsQMGH0eDLJ0lw1kPz0FPs+Pc92SMk3UUXguiIFlAa6LrTTG33qy/40Ag
zdfxZirZstbrfSE/EF6UoUekDguGYNrauxuI9WY4NEw3kqW7aKMBcdIBwzk0
uSwyuFBkUXzelqUnDwT8VFno4OURAciANG5YL2iyhZ8D6dAmxp8/0UnHuDxm
S2IYTRWqWVM/MpA3JvEhZDICgrJtQ76576tuV8z7aj7e/4fVJOq1+A40BPnA
539fZ4XlcTYax7hIwFJk9etWTnHB49LP9LKm6MgL3yXaJntMnebkYJRpb9In
kL6888huOXPU3/gcOec5CmzVhjwzUJUcczYDZ6H0eZXDSWjz2sLgxGaPEHGy
BTsbM8fRcwA8fxQ1HertMCSz9sSgyMFc1hOpq8kioFVqLsOzhCmU8KDaEFgM
vBmB1uEvnpSXBBBsjgo2uwyFtdOdyF6cyQGz7UgWlTS0i+fjVYFPxcUDE2y3
TZSaoIA3/VOUqkBUUyY2eIWq0MjbDm/MYhK26Fr4frYwBdJARJozkdFeCyBO
9yg/88JsDz2xX1GHmT/MWqr6x2WmQVLo5+YSeHV2TBEUj3KN7B1uRDaUSkze
dqifmCFVCiRphFHEQBIcZb9GlvBP2KQzBO5EtllRJvu35HYedu7Q+XvxH9uQ
/TvU9BPbaGlAxnBJiqatJtcMV/AGe7IS7mXxihju/vLvT6olklv7l7tLTs7k
t0HjcIgwSlu13htvccoFH0MCa1C2uLR36Fa8r2vDDeT2l3IQ58+dUt2vlb4L
VVaP5hDEnWgE0owjLh5TMbQWH39rF4cr7JWbZGUloD6O+0MYKd19S4l7K8ow
UgjuYNKBFxbK/jp/2xWL+CEspVsGVMzRSaxslp1PSSwhcei2yNzIhc9wCmor
287LxzFpHSiEIaNYYRDLpLYMZ+rWScOY35hWUETaYglqzqT/chmZoI5KM8O0
vVSbvUmJpL5te3sb1OoXC2D+cKoi5/15zToHlfkC/GAONh8XDCMwPdtwq84z
gJT++1mWCqhIGRTVWp9779L2qrI7oP6I55GVAss7yX4Dsi/FC8z34bTiKwCQ
c99P4rC6zLZarxrsMGYvOrU+b2fdrMi83wNjFNJUtwRueSgzDUg2lm0xOah/
yJxuWNIQiP4zghkfQpETzKFhO26D2P0W6e+ZIYVWlqCY3uI5x7g9MjxmtqAV
ez24YljqGka2XQ+7ocqJabR2E7t2JPVKEZ+h2KcHzI2v0+ylHZHv8YHShl2S
PKxzFjdUkIVF1YenXe8zxOzWr+WJ1cZngdOzOupFB7AMkEpUefOvFmAH/CyU
BXZ/ILwSpWkOuChaf95k5wPcSj3Y50BSYXusZTaB6XR/Bei+dvTWZSNf/NT4
3cu/aIfTpv3lA7pwRnvz47LaluXzKftajWFIU61GE4Gml3Njnuxp5wuTgRN2
b6eu7rFDC5sxDBM5HeXaqEy27160inAr/nnxNaSGLGBL7E5rvNrOxU3BMXgQ
n+LEhFW6WzOWFKvMs/tSevOs0um2WW+LFLYP+pkD4Q/w43QlxZazUYUYjfhN
+9RGVWVr0ZnLX9dGtDOJ190xJOiYQDTu2mLcJOjrDFMmhpp8D5nqNBDCocCl
USh5OF+i2vbJ99f6zuq7gFdeNPZKvpiUZ8ltHqi6oPoVk3MW1jmq0r2daqcD
pzkgztGoa0SuJS1MQfPg3XH3Ccvbmc92MihwdIfJFraAAVOTrkeJ20ArXjSY
5TEUWsc3VKxf/AgIJ11tyGazNSJ8uZJaM76WqCfZFST5cAPac1HoEBYN5t7L
4GNjQXSngaIqWOkHdT5YolSgiRh0WBbrSPuvySQYl6A9w3O2CLek7CU14j4M
HdzEbN31Adqq6adNMX9pqBWNelrwHZayvb6piBFSDsNkOXlVNMgeO1gOO51q
6YXF2z0LZeo2pzTKeG/bjo8RUjOaG39KmQ8DkkeNzwbNmExYomjyygBcLL3k
N9EtvvYpi3R6wBGXleXwMUuB9i+aidCdyZiCFw1oP6uetL8mxz/GDYN3iESo
3YX18ZcTeUfMXBGmJQVDZSp2mvNT0n3xuHJaM8TlBJCZO0UI5tIzls/1hzaF
mF09M7AfLK++x0HOCjLKF9y2L/HzsH9wlCQWybpaP7AUnVh7mXgqqi0uRRTP
jXKqFzvWIWtOkAdPuPJUmqE8i4G2tbIsT9A6T2muFw5fP/SPKV+W+FI73qqN
k3PUJNIPPs8zcvbzgP8AvK4nQsxUsuu86o7UCA7TktQ1lw/o18s/USFUnJmz
wH4r4dClHx3YaZDu/P/kgLOhl9LTjYZArlSlbEmoVpe+zTvlkzyfiCQix7EL
HOY7xRegHJttr89q6owdh9poouwWizX7XZp/LKJJxTgOJbHg8J4DeE9pH3LN
7qvVEtus3tve2asTEYbDt8KnesrRE/hcS9sh8N7Q5L2K/gZuV9NlNpkg/GhJ
T5S1bZyqKOl8FS/Ig49duoEugx4h9hgZ8JaGTKt1VmySPlti1GsmSWVk7w3G
K9q2V8S3I1OOcnFdH9wi6p09Pf4YctH0TbYZ6jWCCzdKNRblqsl7FkPYuz0w
TxU0dvSAPAGQEgPxu9TzuqfaaIHkxekZOInRjmGPSsrkl5+TOMGulf54mFsO
KhPJyeGDZiYI9cCRazoqUPao8ZWzhNeJfX9BeRjk2KT9p43hrdH1BWFz4Y4h
B8+aFucxmVkxWv0BoWmQcL+6fOoCEZzuKKevX5u9F8jToW1QZuqbhvUxytsZ
02sttxSa3789f47B5ycq/WPPFM1Ne5sPwwQy2WaVKKDkP4hwbDysjTRx76Uh
4EHgIqSOQm7cTbzwD1t+FBGDZot3Vy0Hz5bLFO4xrN0Jz7KDvLj006YuRoRr
uH1VqVlDio7F2X1kuh9VZSRZhMN3oINjhtRBLYZQGLO19ve5MWEjo8tHVrao
81Jn1XU7cDUh+Ndbsa89S7c763ybp30YqFq/kpgQm/rALujMkDQZomhZ/K6g
5FleT8iSxj01p+XN3r9ns668cCI7f//j84b/enQfMR+PhgHuK8cevL4oHVm2
Kaf46YgdnTy7QxZeSBGIleQAg6YXaXxpeEXD78VBtPd3GCFMVkhyRiNKKcVu
zYDQP7//ur25tFLjLU0ujq85TWEfDA4rfWAG1OwxoXFMuS73BRrxHZIULY8K
pNvcbB4jvzhu20N+rSekVBbfWIO77QOPD5X83uYEII+cplAj5LO/SvVcqDZq
G2Xmm2XN2DK57S02mqWLczHYfpzl4Rfv4p9Eo0hxfKoETUd7gpE+n+H2ZSxG
8HGkGE5iIgUFRDy/ZmTcsS2lXK6oYUKCRFwTZ2rblbmFwcKD5Sh9IdnwE/+a
UIdhec3N347MHcnoXCdFE6Urp9XQR69dSGzoBxP3vTvsxMCvQi1No25wBDeu
LkCpRp508fdkX8KvyiCxEqFfK9PMogHKg/c8W8xyZrlkT1RKoNmvR8zC++yY
4mFx40GxguezVAq4ug9qWeCnBRB4o+p291DC0O4TrKkOLrnF0UHMW06YBpiA
5Pr9ZxyuFCa9Fmc2XHK5a4aoxxE20JyEnPWHqhWMfHDWv8MvYmmOy56JUOca
tAoVkehjfBA400QXhFQmpZDm/HWEbjApUXtx7tLH0ahsgYZKAFWpVoAS+ggS
H7HX+p6f6JNJ7Tf59K79Dl65Bd/vpuz8QJpZW29wIj4JdF9CQ3ouJrhyFzd/
xw+KXogr5pM6ccy/6zZ3V/EjtHBGeJecDZbAgJ1pb70wKqWoXV6uxhSxrWr7
SoXyvJlxoxUZpOVdRUZr02bRVjEsSEIOotubK6FLGejOL8c+iFTvQ9PFgCrz
DIhYIOq4tpTKpgHGqvMgqpJCmlHKBlSR27cTHm8/MiktPlfcahSfZuod9uD/
hB2n2TfzUj3xtQqBKekJ2Uj9ORnH9pRjxN5pTLilu4UZBST4CmNZm7YRLF1c
bnaxfVhTLnwwGQ6PFcE7ldo8YVxqsv9YSdf/h64ue/pmIKTRw6grjH745sw/
pkNUhgt4SAD2nCKeDQFRdNpScRtbNY/X9rt4ei1q0w0U2wOWn2xkUfaviePn
eOVArTUSzPsHWwazf33S2IDM6s1CluybEty3Gij+2YYnxBH6xMe+8/ElkjCO
mFipzbHCm/8Tb9/aeu+gdKTpnVoOrJj+G+YozGZgkxAw2e2iKrr0eSksBC65
AMEf5CWktaPxZK+mbQqnNQou1huY0BjZZGOf5dqxBykkqDrTqId6GQyMCuMP
VK16lBody/RmgbbTM1l67NunzAUy6cZZ6XuqLuruyIl44TSaYCZqtTStwNkX
XymHUCu55ObO4wDBPVRh33Q+IxsCmJXFbuMrWvSrv8/+ZsTzRdOBfE+vbuMR
L4yMr9XXSlcubBSBMdD+TzF3NdFgW80Q8bBcWv41dIviYYOlSzlAAVToH44U
fQSfSoSIL+FxttGgSiRS4mtZd5nDCf4QgJX5NVETN5lNlXQoUDy8UM8RWgNA
OlQIlLyDHsi0UIqrPz+TG5cJcF8sESokj5ge8LmE4COoJiXMDA3gy+HEG98U
lUdBAPzUo5UkSTCWgO92wG0KMWiYfHk67rIxhKPOtMeMLEAMSWlBJ4vPs35x
QgIm+hZ3cbdzKMAB/3Ky9dQL6z+cdqj8HtbKA9g/MVcKPMv6tjfpMV88T/3Y
mZkX7u+HL52vWlHIcu8MCSMx/dYsILrqwcXuo6kP+iQBV84fdNnBJwpuEri5
487nyapGcxjWKgDfqMWBIC4xSEEnuCvKpcD3NL0wjtwrTFcYDmiShJBYJ1VP
iHwWx6DmpUIyEVi8GC58CvB3bSuQ3VgbexvNPmAV8R0cMLBjwSFFuUdtyvTx
F5PAWY0eY446g+TQmlEWjX/NKJmgsTLgbtHX8oRBEwyV620/8b7xonU5BtJp
hrbTxhJau5g7CB1HNGxU/xwUlmtRSF5Z7dK3FrnOFIRT3t3iLbmS1vBGYcvU
gICi6sNQIG4K6l/4EskyDYXB9/EXHjBu/F7MMz4hUd6ZopJ3jxzV92rJrVbo
uRIdkNY02cRZO4Vsk6CJ8RcwKo+ZGcV89ZXqvzhO6vStDNyn2/+QYRzEFNOz
5keTANl1ksTcllBSb6mXd/GmXEK+NxdDSBEmcuwqYCvu2fTWYn++r+RTomN8
MGuuPe2CBjNqoXfubD15cGjumjndmqkEVL0ujU1SYaqdAnIFkvJw7GjO1MDK
ELH/OT1TGOtrZd+t+6OOdaHf7p+6QxjZVxGwr00vgTg93hE2U8kh226Ej3re
WB7E48EcfVDtXOuDUYyDQAJ+inMYXwVHuoJD6Lrccpc4k88WUL4BKB6f+mAB
5HQsuNJc/H6OdTowR2pz86hdcY/sqzUyzTp4E7yQQfjnuMQhXCofytXND3Mi
zJ/Xuro6rYpDL+GEXWtpipk7LyJORIS81moHx2fbEWPIKPZobZ9Z5K72A2Im
FZVoC4v9zzKjYq/ho3ogPViUPA/cHp2rHhSZfB+PjmsQOKCJehqAiAhYALul
ezqBitWYjhjyxpGX0UYxEtiQbCreimzb9v68+Crc07Vxev7QShS4PZbCVkQD
mnZ+UnB7K8ojcMlfEADv0UVR5ulOYJHya5oAPA9UezjqMaXhKy+WnDfxcrEs
uZkv6IDXzOdoqrlAon0G5xfHIZdHXyXwhQnRCvTNO2Q8x+/Gjb1CHmeSiMVk
+wVhJUHfw799QPml9s7qXZ+ss/P60hLi/dtiPQ4Dk+JXhpQHDXlJS67v+pFO
1H6n47dapjH4OocxtdMY3noWsUhy/K2g3rMAo317OGWm4LpnvsEQAyiaBYqf
+WHXDm8U/BNBwBTX2OJ2rK6Wk8kmDZ54paayL/fEFCmCM0EvnFB4P0T/pP9b
UAb+sDj2k9Z0/EaK/Goz5o0yLOes0q32HvXeMOPAwXeFDz9PSub0TwleZYbj
xLoWNfgC6asaBKayLlAIi1i0vnjec4f0ddRBEMNBP4Ov3W7iLoUsAgpe3Vf2
YnTzdb+J7tlJ2BqFikyGG1eyLn0pKJg0j6w5hr4Av5i0BTjmEakS0CfjtfU5
cDDYsK+eG1KvLHpcVY6PxhcdfCIGEKzvqu6Dm0K989osCsDpnqP5Wa0de83e
OEaYLhn+ghQA3esuf/FVzzPqdp/bO9bF39qCVpx2CLQ+LdLRHd+Txen12CbW
Lk4/2KBazHZYWXF6sXSBj3OMYyAQ6BFNBgbX4VseuOAr74Vad87W0/GVmpTB
Q8sxsnJ6StvRgX/lxyn8RgfTI58cGGYTWuYWIppjuLBwDWKAFYdz5Y/LikGz
1jV9mWJAoP0w+vKE0vyY6VZfWgFpxfXTkeVPhq8PgN3yDgF3Wm2x3J8vYbSQ
OJnkacp4YuaDKUxBJkdEYprGKIoqp/4R7A4bqBgAQIXDx16tUewXC6CHi2Vr
9bujQEtUvzcLw4pKqdyKBg/9sn/BrkGFOlMbutTy/i+wAUUovUfHHF3KCv7N
4n+V4A+kMec8IIbzi62VGLnennMtwE6KxvblAUspdyjg4MJSBrgT9FsR0bBO
9gWPR89K0bU3Tffch055kNpx43XW2KjySNw0HyqLp0jR7sooHXNXLRiusE+z
Wt1NW1UvYphnqgpmWmBWBmkTU4vyJTWrSvR+RvRLhyYvlWIXTo1iwV0Dpphq
NUMQGjUC+f3E7khq49vssZb1Sy5IW9XDHlbRVH3e5SxhUs+ZVPgzd291qxyf
/qz4Uj5MvgKDlIdEpTjgRmeALq3909vR7EUj9CUlHhJaSJJUI14BX+N+OfRw
+hr4fURw3SoyWoxx7flKu4x5gyqX4Hc8PKgoRAWwiXM8DpRsTG8WKKpULMcJ
cthdKEmztnwL8UkBb7XuagDpYovqzU2idV1KVHYHZP7587aGcbeLNLPFC6Yh
xui1z6NuABJInh33Q/nhwFKZUWw+e87pQNvVRCWZYtwy2Cnna1fdC8a01qdL
FqUkSM+MsVk9cUmg4weppre8XuLAxMw7IVkFzShg/yNlBGDYs+sge5jYAM/2
mueIJi+g0jic//BgZLbBhIWjL9u5JQGXtZMQEJ3A98zVBQuoj7/r+PhSCUKR
3zW05kqNNCIDxBBdBHdmbtkLIbjDEoybM/OEOOAkub4vwuV7AkbW0OsVORZL
EkbmOr+kZH3ijq+J8WakObFyBSqJW/lyqo1zN20cWfJfuth5Nsw3o7vFlQmE
msOrw4vhXK0XBln6cYbOyHPGHzlRoYQvXA46w3ObN8cSZAURDHmMu7Oex0rL
rCgtYWOkYYcv4QPG6flUDdD1pJgkGsOIpFwWuistMCw1eXfTiUS34xZEFfpJ
rTykfSw6IqqXSwcBSJJO29xrQlUZQgUnpIGOll0tbK8Wl2Mm3zaWFHuA0XjW
roffr7UIjGqZ9R9h7R60iofqL7N4RuTj2hkfbBAxDB9PgLoUrtLoXJv5E7i0
KLRAJb2QUPVvBn6IErc2RmdtLIhobnF5mYvwMZ4UVscpSEoWmPftxsca6uXe
fpQq6+MCHnu3Q7VTPhlavZcGRnEg641xBgYp71XCiu5CwiiLYvoa4ruh7XB8
gYxKf7WUrxkSNGaVIfad1eLrQtXpPrDMJM14CU3kVD+yCfbLPf24aeAWvOc+
VxvVE+IxsukXLR4JAd2vt/aWSweg5SkIcEsb2Purrzo3aNofF0fUXcNsRIK9
fVBRhwEx7qgLsajqNYZh9XlE1rBFd91W/iuh1i4g8tZKsewitZBSLWmw7f3R
EMH/H6eJdtuSlUSrM1i0g2J3dLFptXUc2SLCUxqsgnQ+ED3sES3GKLAR2c1o
t2yl9dTwUDPJUPjN3U89e1+Mw1nZ9QYlb0i6F40tMkJDscFJ9mom2IGyHXz0
l0giOlyLZJu98/tha9CPo9xAJhed63DO9BfQJt/yCuru76HcSoGM2v65qOcp
HDtIcetb0fvIXbSbhldwn3bhh+KNVDhr5wI4sTdG4WQW144Ux6sDnykE7MHo
FHbzFWtUPFsCyJB/DrXLAtNr5pp9xEhouvteqd9q2rI9fHJU7lKwy56eYU43
jGYIzNdpRG7crIZ90R9t7JnG9mLjB4qrwvTy0ag0gMk/Tqpg+qRx9jKKSNH2
+c0L4tooAc3pdVwXtXKjlzt75THk5czYtep7jRLjurXjabTDxhjVKrX60cjG
w0EsC97djPRvHM4UgOQVtzRINez4V+GZ3eL2MPi1UgEfC0xrChMiKat70AWQ
O+qj+0FU22vzQ0Vu9ZcOSr654yrg4ALUMaCFCMzYAnYwZo+CICV912KS16aU
2CM6FcYlmoSGdE9dOghCcduQePYUinSZMqSTSVxC1C6SNmxreCayQ5sLB50U
p6Jmcw+Ipq+jlyZA69gg/A4680+x7nnblh1f46E10E3BHsbmNFBDoixDHU7r
2k6MTTa2C7CpPYxqPo7D+ZlKXgxaT/Y0gSLbyly8jp4HMnenNyBrIL74o+bI
X7+QBRHQT17KAW6DeBdCvUNkzitVFKNb0G9p6x3oLrpk6crNtca6xBLBvK9m
Z7f0/3Rg88qY1NqFjPl2VRU3U9l/fZbqHuK1Bakm7/0V+OoPgla5oM9aYOXf
VDV1MSkkpgT9JCAT47CjikXwV7nfSRrvty6ser4jTtbALey0aTN7JSVqueAQ
V0GcvAzkrwYwdyth70KWTa6Q+cE8/hA7vji9qHlAY3hMW5eJdzEWGwVCID3f
8JQiFU/Yd6/cJpSxmONOh97Lt0ynYCYbaDOQ1oYvaLt3FOiPSsHaSQlmAQcn
HB2PtWH6ZH9E3QVYa0g+U5xF1+sSw3rb++icE+J+ceeuhbFTNVSP1tsrdkSu
UFjgNgiyhSOFalTnKbA+YD0laydW40Qpax6hiSCYzau5pZpagsLwqLAB9ukE
G0edxAy6eBVWg/FNnoXQel9neQi+M02mJCDAMGxKbIift76eHXHso/U4yo6m
dkNVxmDj0vlqXRRB8sMob1NfhO0HNx40B1rJWy245supDBPxUY2Mwps4LDEH
P87/TxoulK3nEONjJAcKNHyaRR8asmaUq3YL8VnTCPXFVIttRbXGgotTGSHb
HrO/D97BaEzH13NC6eLREjIZIDmKWr8VVLD04wdfBjratLGOUcwQTEvahiDB
zyuc6dqA7iaWvePhaQ3msC1oaVDeIAnBIyQgbHZb7mrmlw4TJ6ajGv6fXQoZ
OLQQQFR/P+vL5e/MnkUmPSd597Y9uQRUfJctLkiuUkQmjfpvjAFrIp+GyBaO
p1lnqOGX1SUNibKCxCtBaDzL6vIEW+YIuZhAeQFRxA8dUy31Ebw2FtBkxD/9
ekwlwc+XscTwsa74RWvtMZxPeTKxJ30eqbNVvIR3opx2qTyFRy7xsgN1qs5m
E8a19UNPV+2yn2jTeVbIncNQd68LgAeH+QUwZjvvk440Lm6hL1zf/bAy61ol
rEzhx0YrVvGRjH11ucqNf1r7H99ZcOnCzcONyq4FZEg/MxaRjJUUfiDii05Q
+e9EdfjjagWE7DtGAEysHQxVWwXqiWycl2kAs8MopGyym/Di4gAmbSie6F5f
NqfCDKmcV5QjVTGeitjYnkN/C12EldNLgeBfaRZ4BHVbE7TqIODCzOQkjHXH
2gprnLVCxX5rij6gGDSSvr/U7ilrrF5YVTYd200AesOAZ4Mxlj7zTmD5wAoD
aXF6s7hrcLLOX06Z70FtDEhQ1LrKA9Cy1SPjZIL9kpvRm2ZGdhbvhUwOXTXN
3ipaYjMP+ItDM2OWFVLFN4lWGjtHSXK3TDATu2g2jmH/27Po2Wgqs34edk3g
L5iTqZejuvF9viJSx715EjYbQrxobIkHCGccliqBdQHcpoTpXVQqeI68k6ys
33UggdEqqekpZ81/gVJq9nRHjqTxnmC8t26yv9HI2vZj6vZbIuoxmjxxjLDT
YFTJnKaIQvckEr2VFmUmub0hLLLHth1VHIO7sJDjQzgjSBwO+bQDJUzFOp0s
+1a7Kpb/KAzAjVo1/0ztE+LmtalME0gWFNaA5utr9aQe7BB3AkNUILLDHgP2
XmO/dS5uOBTtMlCLWpR2ixKWgBJWB920VxaEKJM4m+VAev+HI0qK5aReRYnE
8+ScoPhZdxbcC7Ca/EHTKdjjvnu9WBBwvYp3tg7Us+l6Hh+AA9sttlEUuh0I
j0bcamDLIUxGx4nFY9S4BGIIvP67rgdY0VXf/InM3FwJO5Fw2WmMNdplayxg
4dUdoeU28FeZekq8ztzuxjLzwUunDgMp8reHJwQGglsnjGdtBpgkL250pM3G
bB30Vbc4PJz8sAy5VmE1r/b7nJpE7Oy87VbAubwmV02i3+HtoE1EhReoaDUl
lnUXR7BA4pH7s3Nr4fPLoTSw9bmfaO/3Y7cKax/jDHe7ckf+5OGHaCHz7pBv
IA8W1VSMFOEuuM5Cu2XZFEqnCotKuXcOZTFWxIZUi1uPCGE28vFiep7pJsu3
OC2YUY6Mz/2U/yTTg/8kCeb8UF5QwCCrF7OHUAAG/E9TgumltNTsaHmZbtiZ
NfMZCMR7Q8Qo3VSMba0ThwrrcU3iw9NP3dE77ZYzgblexTRjOYiT2uVFks8F
dET++Lq2QeI2VzsoPpHERRBzQQ9IFX1rSoOv7H6bCXYuYsn0AWFpnAd0vJ6q
o6Mu/GmMAE1ZGOKBsrI8Z1mnL2plU1YC4nv7T7/bo1P5HvJd3jOxnodpxjrl
eRvRZo4cKcs57wQgvS4RZLC68TqM9NVxvRt1z1k4MKaPiSZJSjFfU2YOlSa9
hEVfm3/9xhB0xBW6NFLSshonnT5RPCSDeYcEnZtaDwdFahbRTRqb+dWcuDGi
4GvflzYp1nFmXbd96QKjp8hY0L0tsehDFoNo1IMF88DA8mkDzW2YH4zmL/hk
PkJnk7FQru0EZSf8O2fvn1gRwczbJvgmDX39WIrucQqymFqTFg6ghU0NAY8u
LvQqcUaztOpCpfPSfZgAidZJi6SZLSzKDC3UmFhI44U+aPQf2jEqvx4VKm4X
aCQR4Eu55zsepdg0SnIHHlKVzMZeKg574ZVNywXqzJ5DRq3SCXuNcybRDnyY
1mZxB6Yogvrk28bw+yQ5rPoX3q9eOx2gGCUvPQ1FuxjEUuqGzY81cIuhdeuv
SWWXnlioTcq59VLPa5AFup2hl65gp1G1l24qjS43pbGUTYSpR422URYXrfpo
pzJDQC8lsiNemWB3y8ReN3dK7PC5KxhbbOupa5lCX045LOSS8gtAOM92FQAW
36STeJG7MrO0w8z+X1+WLxzSi27bYeMFk/DRCDF3tZsIgn076sgQ7tpoc8JW
jjvg9j2IN821zCQfm2VYfpQEjELEGTzmFmCRM1sP1lmfn80qxtQ7SEbuXpgS
D6NCyizYw+FCEk7CjqbJvx3OTg9owr6QNcUgrOMf7E8bc7rbHWU25779kAjt
I/DEKZK6RBNZS7mDvQe5LwCt/Lo9K7Zyr8p9ifkZDfEeJEdiqUx3XfK3qlge
IerQwL/GynLqey090CjcUUFCJTPl7LsCifvgSzAGMB4HzYzoo9/xmjEJ+dWt
YxCcdREtJL05A+Z27vBJgWZ0BskhyPvCCWsoF17YSQtLFblvJoTgfI6rRsM2
3iZfK3fl2hU0U6f7UDYUaw6RBMnBYfC/EAgtGM1QdzVgXGxuzrv+kallO0+f
zO6Z0935BoR3clHlfgdn/q9aU0QblRaBPLyU0wY+tv4eigzfCoQUXCk+GavX
zo0ud5sKQg7pQGcsi+kUNZbcfE1yF4jhMnfLwJbitisIAJh18IgbFFtfINGY
x6/8yJySlY37ONE880V0JGmuT9j/G8WtfSd5pTvMpDvcPRgMdPCeDsL0NSBH
2t8n7cA9SR5Q7ko0NnBNkwQJiJQhA5LQviE2ttLzG5TY8+cC/wUNe28IPbEo
ijpCDVXT+yhtFQTXYm59aMXKwYoxAI9dWMO+cZcR43DS63ZIt8AiD3iYA8fr
Y4VeUBXgRLi25FCK/AK+OPUH7ErQTxo1k27DYDR+3iT4oNoPBp5iNfwiIZ5p
jK1EVMMZmr5zbzuQg50hShyNIwF+Ri26R3wY3bPKS17iHEY2RNQx//4gPKQB
u4zSfFqA7u0ud9bQBpegW2wPBLtU9vaqPuWHeikX2hT5AMisSkdyqpiy/WHR
t8ezL7pBTstLtdXRfU64rrr73zmVnVMzd6+mJNNsp0sbwR9q/Ob+r/esH01c
Du+fQ96GmdayOjWSsDSxsCQbn5HgP0vAbVdKd49B0Jfvmpx+pjlyc3rrvpkr
VRK0LCq4KDu8RJEvYLRCBvNePEe6ip9G0FEXsBjuOrjqdSN4UZMtdOw4SqV6
imDqCOZhHrD3IPz6HjzfKS0QU2qVSNIWhz+GLYIlt4OjpY9aAgW8+M1Cqb4L
hqYSQY+zCFuetfVENwuahAa8vt9Y4PjXWQmvhfCdYoraSR94e20rdAIJ+K6z
jdoVBk2FZ91OhjrTGuWMr7W2CwaYAgvLBjC6wEfK2xdXx5InW5R5M+ixUmYM
LyNUwFMTvJa4B1oWc/kwZCO3s7HEzH/DJilTUsYqrV0Vy/RwTdNTxJLBOsa3
rMCsxxNEWB7+nm1o08Nsh19CSKH7DgaXc1bzF6hJIxFzfASxHy7hfkkhps5q
/Ol1OeqBBPATezZ34kbZupVS9f++h/Qs7Ds63Rp+BetbYcVBbKFsvJLhckDA
mzYQrc1UrSKXxgKuDzv+3iX0EuTbmjoIq+s3/dE6gxhY7IaiXEvSUppDZ8iO
/eI2mkTboVMdwpi7CentI9YlEeRXxAhYpZqrYSWBlK/0qOyJLSAuPeImgYdA
EOhr1XCJ5u/8+ZvBC44Kzlskv2Z7xLfYhcbuG9yhDFK+oYW8SgJrF1Sqq9Fe
TmeqQpx00Op+MehX/3ghuY+DfLEpTbZKSFo55qCOj5KCmM99ZY5J8kEnQM0O
lnHf7kMSRcXGi1rwyfwjsh780kjGdsqjLnf3POsJJP3HlASaqQYuTswypgoK
E/MiT7LDHDjKhp6xN1N2VW8YwYDpP32Vt2wFDi2JdoZiGAJ2r6q7D+q57JhT
wA+8hkEu3VjPJn/Oj9sWNo1vN+DObUww5jZKcwfR47kyclhK+GRLMFu9KQc6
ryoZHKumjZsKPZzaK63V9s4QnrrOtNdXWaXQXGh1The230F42Z7tHFBiee/m
1BFFTl5EZS35fPJrwnUsSeEurnZKl1de+6JdY5RMfYhNWUxLiUGXl7rxrzky
QCAyr3m4qOmJ/zDkiAWp0fFu/grAvKEnJhQVW+Tj+RsVPQRDXAb/9ePVU9Oz
Gba6nb2ZSJzUEm8BChS+TSBy9xCKfqstywCi767C1ae5kz+3dI6asmtmNSt4
REPRR6N2IBGyEYoQwET42nIQyoKREsxcQYdg9QtHJJW9TuupujwC3AoHklxS
psEduYlBuFFH+XoEUDKox1JpBmXk2BbSOyPlOIHB4WIlN7mbBc/fMzn96Jt2
mARWxkbw98F0i8E7SyYsDzpb0fywq5sFTbfZX3zvvm7StuojeAnD53SZNl8t
L6Fc+2EtDTBmCvCUgHAYrwjmTMDM/ez7UmhQmb6QzMP5mei3mXMov1qb6NaM
p10Kx99BECll2xn5IgmFF5m6NV6EfReetwOOUx+NTxsQCDNdyqMiN10hYvqM
ts3VGajjokbGo7hRfFNkUn4BnrGKr2AdB6A1NYh5XQR85KRN00fLoaqdoaEY
rDw/b4wpjmIlzf2iLRCXnI5uNeVva2a+Orx9QvPQgwsxWTjHL+PK9kuSmQ+8
XbTardOgw8xNyMQfFXycN0WwapCz21mKsstyW0L7tZcDQqBi2T8l0IaiV0Ic
Nou0P7/SSydmnfzVleyH0WbkbvyV/V0IzYr853DBQA30oRz+Ba9PpihNUtnK
YlOEZT7baSWm/wr3aeCaGw3In356smuovwie0hQ4KarOA7nlUKAc76XDGULo
/yN8TrIiZy+EBZMSn6ZsN/i8gtp9JTPST5qIA/CF1aJOVfvg2DEw0jh9/SHT
2DYNMkNhH+ECRNT5xodo6yxV8ZzchKukNfj3accrv8kYLqMAaWTsi7UjyZZn
zZXtAUGgVB6wJrgR0T3zjI1Y7NMQadllq6SlTHh4JocVUk/jpuUejzpIUMKV
4Eq2XL/FSJMIGBeVEA9S7eWPAVHCtmtH4gtam5deekKN4BNNzvcWCCX3SCch
UQuBVBb7icY6nNb7EXRmQcuhpdL54mobgNX/s1eUZdz52IDfRCmvttrH/fVB
EFcUxLyKl9SxkLfwAapWccubRXgClCnatAY/s+7klIsc+vNXTWtbAt+GJX4s
QfcU2ga4DRKeduOuj+vm2lJ7UgDzsqtUQhXw2G6P254cZKZOUUeprOzdDNB1
ib9ictHR2ysy84EzZgMUpgR6+gIOYpSQNceAbzG1nMS7VXKouByRlntTeOq0
DRZFmQk5WvKIfi/SPbv89XbCJdKj/BPe6K6iKam61/d4lTvBLnBprbyoJu56
2GpN9EZj2SG4CvBWSLlg85qC5nmMhRPyehjdGwuGyuyjJGVnq+tavKTVVaWH
nU3cmkDBkUM8Z94OKQss5KGnF2IOGhZTnYlNj8/5IyfHF7fF+NreozKriAgj
2AOM0f9ZlDkK5Q18AsOPU/sS85e5mDLJpPyJyNqtjag0xi9BwKyUrozzxcEQ
Hn4P2RllyWWEn+CTxHPBbrx5mTYe9N0SNtH9Jepp6aYS0VGgTh1INKG7mlVr
3vbdRWD715+q6ga18RpcF3LeHWSuGMrmgGXBGxtoldl3977dWeSZ2AqoRlOo
bgtBm2JMxrAg2QqKhRZu8q0VtkSxb3cg7NCmln4GqpJYqk9pJvi7WFFejKZN
f2romvq94ODgs+AlBLFHG/N7OcwhLnKXa3XKownJOWJGFFU2kNHDrJIeHIyv
BOYUpLtu0Hu+jANtJur2//hyrhYOwMdRs6f2jFm0lNjLD/2GVE1gqdZb/N03
4SOAHK7tBIp/VGVRU6gAM8yWEK+mXTePbbub8X9IcT8AUfdxWczbneeGjdwF
wPGKUDx/0DDGeoUrTr2B6CS0SK3CMYw++LVmVAJHrOokmbL7OK1nvqugj7ON
j7CZIjwgzzr7o9pequ02spPlFLYZ9q35+42siU810M6wHCqq4P+kXtYEU+Qp
g/UPjxV92RLsBrVnxWRhDmmKzjCsavO6YEQxXagNnBdYJhmVaV6IOdCLm96S
WGTbY4LZhk4gNuDu1hAKzYDanOZZZdJCWjL8gGO5I8Kg7K9tfBYz7j4nSN41
0MKk1vkHnkhXlXVefzw/mdOvBcuoLG4SBbIsLElPSMQkNJi0drrq2HDHbVY9
ac1XCon7z1G+7vbHk0WRXwI/iBmPTrk54/WJD+9CzzcdBYZElvYCrkixVLgX
Z4EIPLfB1YgjfTJGLuFeO061jaNcoq3lWeVzfYs9tHo6mTJJfhe3Kd7rrqLh
aHbATL0zfjaTG/HfxJjAwLpSzOwiBH4czeqW0UqUPCDJEJ67DMu91YB0kWdh
dhEE1sSAmpbO8yv1gLTiXPbEpqRc9xFhYhqsWSJmjYymzckr0q/E7HXTYzaN
d+8IwdLhNORoH8oSKSrphcz+or5DkCwDytfFvCbOlXoNka6edB95KrNiJaDl
B7549jURrObVqHua5VD6nrfgLlWW7Gp9c356OLttU6fSTXAhuXmWioIDrVkg
qyit6HeEPDfGt47z+tWuh7u2LS4t3/UAdSwVLuzqhLnycx6WtEFfMO8Dm0s5
Xnmw3KuTY9UkB6ScHdqeI5C1oLEKR0zMRbXU/YI9lMs4T1QAVdcxX64dN6bp
JBkbQ4AlGQ++WdnH15wkC2DWmm46ZwyBsu7Xkgy4hSpZpD7m4E+nA2zGDCVg
FuN77iEDTl/AQY1m+lKQiOX7uUIWeDve7W+Fcy5YsXeefHZfm04y+4RRwB7Z
0xwafRCvuRSvZNPuQ2lDCNr/nbTBw4Zu0UrhitCDehidWr+pIpgGhXDxhIOE
Ue8+cb8iJvzk3DjmzBSRf9uixmlY1FcQ5oZYW2WUDeXUnYmUAeg2/+YMGka7
OzVJoNHmEnbpzDhv5W1sBxCdaP6lt6ww4PwgkhPVAb6DfUXmICwfca5HC+yv
y0RqAfGiBoJ/1CPqlPywxBGI8Ne+upcpK07zqyDdol50CvR9nhet+wkdtY3g
i/e1lN3lwNqgwXOpHaSX5XKGojpXwD6RzblsMT9PFQzoPvyWBntvUJCaBkAw
WU08CgJUCTgXJ6BRHNZ3U6/y8FwMNTldd0h0eIqx3VH53zKPbLeD1rzI49wx
iN38z3x66KLtXaRHqCzY1kOvyvfftel6RZTvFwym/GqQwBfcEFNzxgggxHgS
20Jkq6mwEwAio2+8I9pbhnPs+xoDUAiOAvbV8I135aU5ZIFwvbzIDX2sskou
fLFvy+rdEE8EnbozugpOxck4JX+4arv36YPFEXS4+YRpVLbekEj+/pwzWI51
mDH6zuS/aeaHEre81iP/q0KG6gBtRzY7rGujKinUsvTawdC0AAz38aZW1NBE
Ig05rY17GtkKfql5ReuKKUYIwe29WooeVSkJihq9cuFO4WPlvqUg2y30P2O8
CAEUVTA+QV4+/tS9xbvvdFILGyIQspkdC6SIK9WCNgr7OsMYk4pzjBK5bmy+
CAyOEKmfyZoWcX4kCefzx9s04JbkehNHjjO5q0C175d8UL3lBRAN4jXuUQqa
u6SdD0+6o6vdplHZtNrZLRIWb+svf67luC8h7QXVDyHBzgW6fkWDoJDU0GbK
D78Q3EcPLbIjfJx7ujSxpCkHopnnSBc4KA4tikF9yz33jTVgw82ZyJxjTxdZ
uVC2nE7XCld//b8gywAhSJwTolx3b/tmXT3U2+nfSnlmOxUct5Jrai87I3bG
eR5+Hc5M1WUMWswS0d0zcok3EOEbaxZu9MZcgrKIhsMSvvydL05oc/SL+Qks
Q9sTcWYtVVnR6eckId1d66i6UOl5HlPpFxPbXmrmsUvFdtz1tckZqWN22Ubf
Eu7qMFH9g3JJsCgAQnipeFdUuZgf++FFCIC9bMr1J88/EZ2mC5kDaVRqPnJn
lvn6SXRzVs5WpePPq5iQRMRC/GVZGN3+CeWIb+46+T6JKTmAz2f6OJr5vvy2
HkOiCDnUAsKbd8lNX1SZK4AHEXYxBP+MiIO5UrePCCDMHgexbapYVJWm77+5
tHFtinGYvap4gNSjDdKzYzHThAgOHq05OfXddBpKhHZzf8sOFoIbUSZ0jeDn
7SHh2Sv9qOFPC0R7rO6C6vpLKhjRIrOyRDusxJotpyMpd+doOANaM68FoGBx
czgvhh17YitjMILsVYAhGndc/RbDMOos2IRmCp14CHGCHb1W8OqQaOsTinlD
7gfXUJSwEh404CscCVWgGVdVP1fXvEN5yaJUmDsByvr7JFcV1+kjSFhx9r/e
+yzCjGFFzXieY6tI15z/8KHnQbZw3PM/VuqfCT1/RQKoA/V9Vh61XHKc/4DL
mljOmtwLrIP+b6F5zQ5hEP4joEDZUiWdpvzSxpbs4fTEb7ohoS7urC7USjQx
D0RZ07tiRBYd09uKQf18rfw/MWida/XM/sIEnOIzmszDAUF4CiR8gQEycemV
Yk15jSxiN/yTBj5xy66mQhfMHtm5hPO17SZQRE/B5NDOjQc8NlQhuLjPPH48
DMiOn4E83nOf7aPKQTeuJneY2HvCS5SnYR6zfNm7LqPh0iLPBmZwtN8X2haT
PxCa2KH09Vbglv+8fuoOZwJnKlYhiIbyjlmOBIUfkWK/Fv9oPcn9cbRr4J5V
5V456QCZ1SINl5MdlqRMxhFqET/nHm51zJ42Z//kAi+nCeJKZAm3zyGSS8gc
4W6ZBLEAxPhOgLq5sKwYM0A+BeRIQyp7q6wyiMT216LkgziB7MiTKellYi3a
XYgc7Xb9/v8cBfxK0JbrMXNYbxQs8UvXYa300LsyOXyEDQIfQ+AKKbf35//K
pe4gJKrtrj0mEVZjeBSjHte0a1OTL2Z8MGJyhX38v1Moizq341iodPgNCC90
OwfPgK7+n8XCRol4qQwmwKqANNyDzsqTJcXtitkYkr3/yn1wvMzaiPr3ir/6
CHeK+uRYUzUNLm2HZTvLEbDP8TLHI7wHvIF0QMQaZq50gNmBvWJi8zMH6BFH
rLJggJNYmb/+kLuUpc8G+QtJw0Gl9fYjt8s4UnYcKdDhq2XEJ3jhOk105PBD
+4+j2zDgFBUSl2PIkBjjLRHlMZSwdBoCm+PL3PsRCP6bc0/oFDLJHm7x0YDT
B51AQtGz8jv+lUyDTOMGmZfw9pMLV7HbpaO1zLozaxw1noqTxKG4q7m4BWck
DjR4r6RGmWfW0G+mof4MzjIsBDTIjnDP/26hHwkZEE1PvVmP7HB3irIU54fG
YbG1TCG+tmr1tlB7iV6FoPb+zhg1uTiTj6MYq64Gm565odoJf59O7an6w8Et
Wkduf3tGfUqvIpNlG9fazxHnGnHbSCWO+q0CJ0JyL5GK64TKfLHc7pLutds/
VHua9BGqx80S9b5SX0/kngu0sVeEZIt2wPmorcTn1SjIarN0DNig/siKn7KK
GD8UMnOz6ff1N+ZICeWf56D9yidkb6ZhtX3PIyvWPP76FjGUt3BvJiztatY3
tgkFzZe/TzGpKMzTcKLhhL4DYajtX/mbORa5dGglS6q6pXSR6kKZdro3cLva
WQkdVaAo9r7JhyfTKhQS2fg3S1zlObRMSL4Cpm/yuoyHRs6oa9m7RdWHAS1b
z9G0MpwuyF5y3Gble9RMmieKyRP5n06HSgeWoe1BU0CjWv4YB3SlxAJgtZB/
B3SYq6I0RjhHAKZIA8qxOKIaAYcRkzXQd5iBgkq37isDhX5/M8zVxYmxNpRb
s0d+iLtD+wHDmEXMSUuCX8KJE5E95IQL4oP8IpKP3qf684R8UehM5FGkudZB
k0kSwB2J+USh4hIYSSEueDlHkuqZVx7QDmDhTekhGUTpRiScy6g1MtL5CT7m
7ZKsdEM8PghkuqRWno7ju3vIEdUXxfSJql0PaA4PGAL1tDjRh7W7WKE2oDvN
XLfsgXrA1Amj5rJDeA6KoZPR+SJHwSiJk8Px9bngeLYx+R7a8huVPMke1vBt
e0OShqyGLhDFPbjUpYRKkiY734w2+CAN9osEMJnXY57CbpHOPwj8O/XqWqFQ
Keg6tdOXh4oR5nMSqbVqYgiu2GMyZg7B2ARxu2eYOkA5Vd6Ua19RtbBPbEgV
hi7W5MsOArM4TIYbPK1PEd70dNxV/eC1Ey5exfE2NLN0XpBcO4HG83JvjuxO
8XD0+ARfM6ZuvqS8yIq8z02Ud1QW/wX3LoleIl/VcRwxzQ+IPBOHxYKASJas
2UZw++G05AGjEtu6gLzGA+w1wcPpIgOyhbZWQkGHWWWvU7b8jlfpE6BWZ1rb
0eaFPipr88eCfqLiqXSH5j9pi5F6Y6M6LvbVlf3ylFrS+iSe/MvecT6gnZgA
hssBbKS0ZOaor4Nv/ao0AnDLgPzDD7OT5O/78nVGyix+8do4kCXtoF47cTnT
1tqaWi+svPwROutMydt+cevWWCMxVZWSGV+9KhDZTFpkuzoCiZtcWjFViXfl
54604r0uyPrGBP59hwA87ie0OXSaC9JbeQiDjg3bOfQXjQMwnqESxhddfYTx
ecGEm8fhh34QOBcqjPYiagIHybOOw6o3Wf9ycUJTfl+QAUMdUmyoFLkaaFTz
xxNkQBdCEHqj337Mh4NSrPt8UgnT1xDV2NrKNUiroE3wYzHiiuuB9kbSudTb
ggQn817TveyCwK7GxwGzIKzO/o/MpCig8wW9RDzbXe6OUWgaXX79ODh1q4No
nDb/wc8O7034wTqr2G5Vc+kTamacorUJlakJeWzPkIXihF/tHGSuNs3GOOfH
wVH7suE3GgmhNE5MMNh93/bIZXcY01LsURoNuzAqfT+B1XC8PS3qMuYERPqO
aHyXzzsw607IS4ttnA0/l1+M33nvoeVl4omDDZow4gAgAyH6uHYZ0XRwG4aI
kCCWXN9mIoew3UJOY7g8+TApEosG2puO7KZhWv1nUIy4hDZWedyyTlzcN65P
eww/DwktEobzmbwaSV3qWLYLrBN6mMa6ScZokXjXckHqIB+6irCANY90Jsxz
K1FG1Vih+jo911dL3RicBUsGL591FRlp5YJGPi5u2Ojj6/Et8PFCz1+CEWfI
aiBQT0gPRDyUym6W0eekm/CtULEuPgFWnuYQM11SrGyjMa+dFwwihaiWpTJ5
ndbXwnLT9i4EQNjPqk0TC0/Q+tJNKEVoajlpooVoHk/rvvgKyQVzkhXc9tJT
M9yqIELmzfE9CqYbnfGRqXUx+vwOCV+y8VmquBXAwAc0MaBbRQCcahReMHMn
Lnib8H+0PHFAiUOeU6huD4tXvc2/XaakVfIW6eIDVVJy/nG1ZpsI6YKc1zmU
cDEVmp2ywZrdznaln6fUxO9nqPvTZaHZEG9U5jS6FSKMiomuLRSV8c2SuT9Z
C1It8iVKhMWmWNNMatk/CSCmYCt8b0vWG3wV5ND0Ii4uZHG4p9OpqENczmCd
E4kUYOjjoxsezP4UA60gCA1ts/6iIKCf9QeKMEQneXWryWnRRVXvfOZ0WNIX
uLUNiEiD/rIM8Zv0zpu9s9hEUXRqzqsd6YuXCbnBogR887FcAOUH9Nc/foUg
9RgvCFwiHQFKLkrPAphZ048pi7luXkHako3L631BAZpzLGJ+xf6SQuMN8DY7
ew8tJRmlznwt2u/+EMm010S310ehJIZvUr7gHrJyQUySIkRQWW4pj+buQ8EO
1M+DM3VdQeYSES3YGKZacNnxuBXzjFVcvHwSskh90cKTgv8KYt5GuwSL4DQb
1x7BtlzpX8l0x6KL7ccWM919n4AIRYhm0Bj+oJ4/niORIkJMK9KddyDsoxh1
2hWw3ZmrNoWsPMv6RlIr+wdsDXbHVLN9AXV3R/7LoWw+4nPvojYlU6JhkwOc
XQvhQExRg6+moZLgTZ2ly/Jka3xsXZ0EKk/S0JiK+PrHQXhLVGhQ/oRGitS8
ApmTH8yiS2uLv3mQZssFGhOcmLob/auPo6n5DktnBN3v3IFAFQKJCFeGbVTP
fSOQKWF3wWCdHdJ0RiCXTZvI6gsI2sDvS+M1G9PpA01K8dQjBO6JvuHoeqb7
kKa25XxmdsFwzYi8yR4FTWxuS1CY7U+OA34dJBnMO9TBi4OXK0D0y85vIvwU
4q6iw9Av4YlzHnx6ODOTxQeYbQXzqtazJxjxqQQUcBkg9eH7NpdRfCRmYCXl
D9ayYBrfeGNuYOkEzvf2m0dkey+k4fuJi69z84ANM3B6hNq5X5Mo1QpKuZPC
xYNVP8ILmlI7j49kAttAhQbbayITBnmYTBaizsRYiJzagBevzISA3wIYiTX+
DYHKNwJ3W+xk8lxrv82onzKxM749ZCwrlDMsf2Baff5pZ650gE9kaMz0jS3C
Knfg8ZdoTKAXp51GHIYLuchPtaX8Q6oRpXHoxr0j2/CBNeojyZEkwaqGKOjK
iUnLDArPnBYJPPAQH4o+/x/E/eOuk7nsMT0fTTjxRkBz+Tbe9RpkWWwa32UJ
df5vUVI1xI/fggzrpYUxNblANgXsycTAoBREwCV3C77v8njnVtkQ3BS03vS/
/cf843+VvQoFBIbRZ0Ulh09q3F7/kXCvMBI2jiFPkhGG4HkT/xbKN801YB4v
HHKg57DU8t3uGYvetORwQAR5atQcIDbfNU6Q4So3VXV/fKNe13d4VzpDm70F
nM7NWYmMBBTb49lBX2e5qjuM5Cd1QFBiZK62cNsMUmtZPseAFDbLrjn0DTm5
lbV+Yo/9A2bcj4sRZNtnpTwotfteP8SM3b+it1LzBInG/hPuWvJ21ZeWfpZY
vTXXy0WiRONRrPWFtgdjJhfL/CFava8oNKXFBHuEJ0REtL4TAC7NsSDiigVf
edlKFtUZo3ToQr9Nci9fm8SDPVBuuKmrMeOXn0fvsaiFHo1muqMlJybq9tVm
xqed27upV8yg29mLA7YO+8QNVmCajduRzu1qBrK0VMu7ycoAQotQLN5xj8EJ
mwMUpx+LT8zs0mnNvNZQj9sQRB25WQzC2+PedvgMz1YoVd+duvoNMFlsMyVV
NXlH7WN83nd3LYlmDrMfG4ZnxtqvNUg6djjnq7vjwfttUL8HDQsEMt05mCAe
NLUpvwLhFEgBZ40UH7MBxxoKhd+Uk8pL6qhiE4WM+AXxaUxJo/yKT9G0j50o
6vVnK5DAQb4krA2WkB1C0mFXgAPr95dPFXqS/psZWVgdjG7zhiTDPOl3q62j
44A1vSEkm4faUHUsweyeYQUPjtxKQp+z9VBqugw8xZV0L+V1v2Z8TeY4LDiK
/f8v88Yuh0/Zj9omsICAuV/sOVrH7c5hApyUgFOpmilRMOlcwtSQ6r9nbluC
xbFKAqV7SYrpH4nGfC0vBQl74N9Ukxu8M7tPqN1bM4sIFGOVOA8Iju3H3tN2
QbviS0W2WwhNLt+LdKQgtOwtshHJ7PL6+BzpkUP7Hd7r7aiolfiTvG4WB54Y
uY9TLmEsVNxZFl78K9NFOxenMRgBTyGV2bU6qQIbzzj2fmedRyCrVjdPZXDI
Ijr/H2qZbnu6upn5i0UZShXCysyJ8mlHfnJj7LHcR/pxr6XCta8nLZB9LD0h
Q+Wjkxn0FyrB3vNXZA6kYpPmSAIxxWS+Zg1hlISTYAzogH3E5Cg869MNPmWE
NaOGstT31dJGDlxgOe2qGOLeMIYXNkKfnE1T4d3XVEFI5OS4vKhb+TjyQelV
nYHVrAN3Z1p+zOVKQMLHyoTJIzSR2gby2ETZ5qT+PSHM0AXhUMXq/alh05rP
LqCM9Lq/eFQuh03zl7/6HSgoZDenhUpxaQH6JIubp+sMYEUVpqV9Iu4epM5W
TW1Gf77+VMEziruXeG1KkIgc0Slqp2w694nbGj6sYx6/ZOuoVgH776J69sJJ
LIAu1FK94oGP+KcYH59tRGmFiMOCF3TV5MhZ/WxoGSzc2HdQ5w/G+fyQg694
xrbOlsuA3i+esX8qbhcOwUT0I9ZB5c3vF5abHDc1nffepRobMUKHkKjIxAtP
67kcZXov2JPDe+Vqx7tfBzegu3+4AFzyxJSQFxiZJTZJfCPAnT0wb40ZokDD
a9azYoqitBD5gu7dfZmO2wvHyZdgXtvNYADUFIFLvDxqTizXeJ1iDj65X81v
woUBbA3SnUCHF5TkAX08PwJQyBAXDI3RNebyHvMgpWe8Oqh4oQGLtxRUjKH+
BSctML/jNlzr0SV6gQIEexynitLaT6IfKE/ldJHCiYh2NWR8aqS5iegjqHeo
zHGnTOq8t54bpJM9NTTLLf9DJU7uA7qpSYnLeKR8jk7U8QJZfG4O1tweqgCM
KJqfLhGaTHShps+/s69DGeYceEG5EaISWbB7vq4pEnJqNXG5+QsIbk4XzoEV
yN/BQ1ldUCKDB5KnxkXX7iqMeT6XNcW9IqQvaNU6ccqJYQyCV4oitXFLsmUr
SL1CuNY9q0SjVqo+rVfSkOe8v6y1kunOcw5Zu0qcuGIcPQ5Qz5UAhoJKKHzX
dE1oLk8itGIbaTrGCOScte83ophgBSZloOWs0rI71ZUehjH9GShba4o9dX98
J3a2jzi3zm5xT3P6U+c7HCHq/kGU5crIyz+V9EBtT+oG9q5lHOnNRBWdJMtw
67ia1IJRpcYCcDd5hBkj9x7b/BXZfmFO+RmJ3HCAn97nqKsIZTGRCochQJEU
LX4+Mj/A/jZsSKERKM2apDI1qnc3Sq72WEdcFDNjDI1kYR4+jpHX4fBQVhd/
Vlx87S3nVOVb2iRmzCVHvY/sL4xZrxj8uaZG4GhtdwAEYVBVYhC7Q+d21r+Y
WId89frHXOfFvmyUns1oPosLf8b88K1tliWOdGWn5jGOpQ9h8r2/9UvJ22Wl
vF7/wouRlnTpfX4Q7NCE3Uo844wIeWh3Su0D1kwwQvFLBN4cr0wvySI0Z7Hj
Vfx2rWTt55w3Rko9HEXeUjLKRkCR7upI9pOsGPDBz252QKCC98e/2Qfg7f8y
pLxR4+IS6agH1SSwgROk1TE9HN6krVo4QH6u83ds5OD6fOQvMnmkef4f2/iG
JwVHR09Re/ZJ49awKf02rvGaPOgfXbI/mMCTrNqGADML3Rjd+nt8QRuW19/S
Hcyy7qwsCra5KR8E9zkQaVFBGxxtAyBo8BmT4yni2a9XW1OCPutMiuIL5N6y
aIJGMtqQN5a9jarYxdZdZNK4Yy/+UXFBhy11R/PCIZLnKzgeQ6r8oEfxgZJn
27wqQRPzr2rw4gjEbKKaTKWnfeAggK/YN3q6gbeKoqTxLSTNROUztfSIeCo4
PGHcYTuAhuRCD95V2mZsNXxxdgyoZPQ9N15tz226V7ONhXEAY6qDjDyIeSrs
XF99FTu7FG7y0CcJo9LWiA1kJZZaRfRHxk4urTff0a9ByYe3afoWl3MwLsAQ
kDqDscc2tapbd9HP0hDVyvLKEg8aHW9hyChzNJm/W65otZiCwvN1uxZ46yYl
Y2LflTBRVbDZJSrXzDNhEi1VApEnP2cwFqPwyzn83xLJN+ZNh8BiO2pP9OyY
ugeiScVwus5IC1QLIXhvYrZ9Xxj2BPFCFLZWnvArAo8cAoAcG0xCG4rRl0xv
QUjV94c6aUG2u9LLGk8IeNv095Yq2DxW14B06zrlbAd84EOvwtJqVb+60AMa
pS46DXuXDj5sxZLEqcC23Q708quBeAtYJ3fi0tsYQ6lzU6Ro1dteZNF12K1P
cGKc70GZZgz0F9bLgmxMehcZDOYpsWo2DyMS+IkxXEN2eIjMJ3JVG6DF74SR
gBGIym2rVrrxmTfU17A1vi4B6emHeQOzuLAN8sVWhaagARI8CAXs6s9XeUyG
zi98TUu+lqC20QEQ0kLblTuxdz5n3g7C0zMX98hkf8OF/S1MquC0bsrc6FJp
VU3ubGT+T9T6nbY0hgliWWjCVYIBSy6TgWvwYecXr7eyksxvnBO6bpsJa6ZH
CtZzpuQ631VwCh0HDD93nECBobYM56A3WSMpD0ZLvG+BVBbpSTYg1S0gYwOK
Kk6eXzu3q1xlhOhSADYNCliG9T6oaSGhgXy8Qf/0/5us6Jj4x1+CVzO4QK0I
yyxFNFiTcsM7euP6Ouzc3a5+ki6szHIn7yPaQjPheICR6VkbxwrRFOL5Esyx
KUqNhb9rNIr+dBD7pqXQqzC7mGX0ABPQ++5eNdOVCvZGTLshGsBD5KmuVf8T
BdGeHxQvNYCUL1SKlCQMTOKQC+NNOP66aIftm+SgV5H4dCt9R5HUHLXV5G6q
ziCbKFqdju2ZnPoty3/FCN21+DSEc/1jtdL0aHCoKxOmAUxG8Hzb4+7s01l/
EtiKl1ELzYCqFw8dbWIhK6zz8EAtXqfUkl36j1XijiigMh+tYnbnQqYAf39X
ZHxl82p8e82ATV9VSj1+Vy+d9Vkso57ETCM3xNLUvhqReIOURXmstMrHGCLj
mdjxC4kvRvNU3OvtyW7E68ZP1zTpjyXIVH2md9QmYG8oOJmV1Pe5gMv8xk4q
pijd3f3Vkik05bKUglvIR5vy+HKuVVTBmxWt0bZTjWa5oxk+/VLmwjyCudvn
ZNEm4KbkwzWyWq9uMQdr17l18kzSAHRrQG2Onbq0Ho1r5JmBJXc6MwC8ShhJ
Pgu9yEMMPETvSUy8XQSWHizODLw0TYD+drF6dxBHZHeggpm+QYT/t/paFaDC
WL82ferS2+9d4ntcDx2/yc/7ySh/7TPmNL6k0eO7qoagauXgQIut8ov93FR5
jyQlLup73kN+Nucek6ZM88bZIMpVtEqOZuBUtZIineA67hefrXnmJ+klOWjL
xtxuNpZZ5VkKU0UKHiQkDtms2CCAm/YavMwmkCFOFwWz8FQBgqWuXoY1Tf2G
OUl+Mbsa04hUUanNxnk1iQUnQzMW7lc09IsIxEfgB4kHeiXbcoBaioLvsQTl
gj1C49RD0JKZMm/ri9KFcPLh6vFvCqUn7YC44t5bGkeAPRSSfKuXje3dJVdU
IldPxeNOmDx4TLl50Z+JEv9AlVVwlcEM+P7mJwd/walpObMdhKX7sxia+sdO
DNYAUbu+v44pVzO6bmqA90J+WGnbw0seQAr+4Hi655OOW5KH4HDLaj25XcSp
sEQZgbnLdCfazKBuk+hOjuKykK3+I7vFnMeTzKEd5GZSToiREoN1tq0cnTWL
nK5YaNrct/V0w/nVtOTOzGqcMGM38VfQxks7dZJv8REwb7y/rTTVSpCs40Id
H0XT0WLVI4G6jaxt0ZrX+724Oe/EPpXfAhLPdFS/SuVd9mEBl8dxjwlVYA0a
enrPRM00Hj9nwTmY5oqXy0/Q09ycgz2vNteM2Qt5dyzc7ZQqVh79l1o7626t
YlcjUTQhKx0RVo/tNSbp2ul16KQV+bJ0BlkzfpfflkRYdtCRNxMjr81CP7Iy
ouL8QtRk7L9zA6v8nFJbbXLCp8By1HFjEcltvCj3Yj3xZXXTObpsvIFtXlcl
figc2UJp68zqNNP/h1YEnPphmCP0eBd0Ognf5Pkdcij05WZUxHLmICdFHmhv
yrZvzzkXH4evmK5MFD3pAOFqKwFY2oWfEUCvZ5l+r6gFhTjt1LatGRtSyVcW
v3ECnes3/GCR9l8OzgtQCKqns951P+mmuW08d+Kj4xlRQWaJIdJQ8mKRFonh
luNsjeDPmR2A+dk8dpDYP4D9fN2RMJ3XF2KqWD0j21lnGuJnFTHqBf+6PJfG
kgpldtdnU1DljSUG6yzdzufcDT6Dwzm+xx747EoG6ij+gTslqZR7LONg6hHc
27X/Nw2LXhMad57faDxF6ZcPpYPVv158vxIkHqfg5hrxzUFU7k+YSEqJh8rI
XGwtwRhVeNUPdSYnlQgozxggtVOl8mlRaaP0FAYKEsQD1MI4bZ9cFoNr8TM3
ZfVHhbJaFegyqniX+NLz0024RjREHCbXcyVZuHxBWYrh7DcIfhZ3qASFkQXN
z3bhOCOZ5cC4GrlI0Pn8PQGLevJdrin3983aCf8ELVD8tjeRDj8plW/SDDzo
fom+j4rXG13IYXJRpdLITINQ7pyqyJt0NcuI/jFWW6dWbc/denwo9bCtYV0T
lfVZhA9ygLA2BtQP1wo3UEH6qxCV9F+DCGiJrvWVUISBfn6Q9G40+1T+EIC2
Py4RM+1hbz07e/6xmQOxJnKsWWKimbSjjlxS4zkj0Fv/lKTR+DWcrDsBPIgp
XrDcEoTtE0wpQguu6wLiutkeXUh1rMNwe02VbRDCDujmI84Nll9eHSqVN8XL
la2CWvtRss2U4O71bTJ+d8Niy5qzu+IvUaq9hs6Bnnxc+r6fTuBvbDEBQcA4
7fyAHCKFOjaT+Ng3tzltd2WolUvp2forh500Q0mhoSyj15tUa/vxJQAxJym7
R8OsSa/HHuYtK9HzN/gWa8iJNkXRnjG9FYQxGZk71lLhrD3tmeKR/vVagAfN
9ulX5gazmqRmrBxACylxK5c/cbvbu9eePdQtROxWl3AOT5PSX2uXOWKK/gzW
5Bzv+Zq4oAhBrenYVSL25sT1al2X7rcADMejgZio8nQbWUrSZ0Njn5N9d6U0
rmA1lLXb3VORLp5ClBJErzqQ2FulcTfiIPtYaBc9057JG6lAw29PuPRIzTyF
WSzVpg0aSSuu9Hr2bTPtdllzED1WswyfSxl5DYFV0IoT59g2glNw16OR8zgC
1RaB/gFxDVkEOadm0cNtZOah7/BDdop1lLp18jfv7ccaRXnpM2TMB6oHaIIn
eFXrJ7R9lcEvEvtOhMLrl3N0jSpRR2tQwvSXxoJSJm+wf+DrqtS+C2UgrP35
5I+iOb23rsEeJuEW8PMlyuBV/LsvNqAgtaLGQynl3q0zIax/6hR1lFnvugfZ
kKNw11LtDtH7triGA2PbCfF3lk30Ap7rY37+gklCCoCfiHEaz7Zj5ZaUmidf
hZjKiKoTiCXb9+/6EhrT97LIxizhSyPwKvaWwbntXxoXEEMl/zvmWg4/zQCW
EFF5+u+xfKaLz/paF7SFpYt4KXaSfiODyvI7zGm0rUowvgBV24MeMnrj4yLQ
1JaZq8OBEVoDVzG9xilQpgFPbcZoFSrfi9fYxXFhmyrG4P9fa0pZOQvA2qtx
hDDoGjI2PVDkh8yXAKEFrhIKpbQMOBtyU9cIffOvStZbPFKGgKnjapypIo9h
R6JAWsFJFrQkFpCH+wUu2ZMOB3pfjFRhWHAbRDUXtVm69/ubkeYwUEwi2Zbr
/MRAkqXUisq1pk/Zd6xE+3wyN+uhw0G6DUKeVLUEP6S2xOzYkdz0Zm2XzfVy
1DR2/qbKnruV6sxKy8F5DbVaosFy6pqkS8o7c/MjesoMbl7tidgbL46cWF1b
mAKbj4fTSyW3F8uxRVksFDKFL/lDtdycMQoItHqqxSPcoXi07U5/jCltnYez
1xr6E926KIoxZSNPiXrwC8DkVNmXjg+5/Rkf75b9tFPgVcfRZvcMCgPp3Xjs
2RcmuGq2DB8CEHJUMveS/SDp9kB7p5NSXPSFwQjFEwBFybcQLGW2EIQFzGig
QWJW9cjBHr53ahFL68jJF2kDmw2uCUX9sJ59QDTlSxCjIydvX7ZvvV7ChgAW
O7TQGqBBl+k0+iliwUlU4cNKlreNbBsVIrHANQR6pP+tXOsgzRlOAzBCrECr
sR55pmVWgBkRgKe11cGp1tI3XrXh1GjO4QS0wxn4iL7Ujf3goh9+c8f16tsS
7I+b0WoULWhbKehbHR9aTCDg5/lMyitZpJr3k1+TnItWJwaYRC1XHi9ivR7P
+AVVtv+r1EQyqnokuHhh3R8vT815d5kubNwOApzNX5KVB1IzV4YC5TtLvwnw
8DfxlRDAbU/wSJGkqkdMEm7gLsZqm3kIX7r9ZJIpu6A7m3dIFZ4bq0QelQr/
wzI9fs36V4wtsZf9YAp3v6fWqgqgig8/LUMZiRCTrQR64fQsXCfIia1C3GZ9
8WpTUnIoHiwFEOuJKaj3bIfCNEuNnIcUR3qRpC1Qi2YRMpf6QL7BCoXhNojd
C+l6z+b1DiJ0ZX1SZ33PJk4x/DohiJw7AMgpDuMqGkGvljXHeaeciSkeskIr
HrCnO7JkATpEp9ePdVFPrr5uLUFix7VYm49Rw4m0VuD5DUhV3KEk1FnO59bW
RIAsEEHGbu2uN9kXkPJQg+GRuUcvZNJI5/5ouBO5El0X9D42Z7j+XKcYFj4Q
FlDeuucqMIvfm0+jiGl1m8TWdgbdhD3bnKXG4rQb1HAMSy22P9kBaqzfwKPt
w8L/vnL0X/jE/CtmdTvV/Lbxw/ZgtUiNtwz089dM9sWLysLW0jIS07FxkRaJ
kQhFrKVK9ewfESff8ozDG8tvfYH+L+XLn2CT4WTq29kqchtmrABO7wK0spog
FfNsHZEfPjexZ+/PBhveBmeDQ1vWfA5TqxqRxZCiCyAo+7g6MkD0skUghgXr
KMtwBhs99bP+osJ2rMFcr4jAcUroy3sPI4XDicwznJNySZ4qMpVpjJZRvHrI
wwQKH0c746vlB9LzKJJtgzbqHh/Wisr7pszpPZ/41DYPF7TOUIkuhoptO4YE
2uV7hosI7dgeaGGFSPbelHQkbt+hkHVeKQt7T+WNK3pwcytHc5QkErXNR3BZ
pnRJuK+ZD2NdbMq1fHd2LUqZx5QYWqYqhxxO2wgEuYFXeDnGaaXdToXBPfzg
pYkFeSO44PcSaj89Hd0aRZY9L1ju2TdzhFDWmSK8hY/LoZ96lkVDXUbaB0GW
coGbmQMo6Ygxu50Sr0nZ9kMBAHdtVsdysiXFlXJRrMWL63j2OGzmJFHMaBcB
EtpIYwjihhpAilNp1someFFarityuePBxa+Uz0xj3U0hMG7WCu1OZSV+qCqY
nZzjcjbJNMO4jfF2XTIvpPacFcd+V1EdiD0475Fdciy3AfiJIDaHxzU3Whrx
9ez+kwHnKgwXRa1XeWBgkSwHB85PDe3RwbfNUa6GyUz+3PWjwqddx6S1Ib01
wtgPTBHyWjMUvz/oSiCWZQIQH7LngZ7Gs1JxwMFui2BsyD4b90MqgKl+odFs
h8+ruFp+62dgMgeDGoCeRGFmYaYqdMe/SlMbk150kK8KuTS8IIxeFldlE1ey
b3oijK0PLxPg2biPqDN/S8OLnh7K6CjQzrVOpHcP3cdxemIdaAcqv29s+57f
VacTvPWxCcmLyYvgGG4svoDxagOjs3mTlOMramrKDEC54TfEZHiiZFsxSKU/
GNdyzfTpDKsKMDz5Ra9kfUCiaftZ47IvYi+fEry2eUBkEHj4TvoPrPwynqUp
kG0rgrbxeYUpBBamyfSFT2RJ37oHqph0egj2rBG4tIk8FEgW0c9xEvzrTgQN
TGGjW46tIhbspM7iYUQckoVjLvvrxZgjw4yDa17+JH/GqdYZ9YRBcx/Pubio
dh6Cvlb/d1nLurKgQgoXJlK7ktJmzobHOTbTk7/wMTRLqqEGvRRNgF6l/+66
Tyn6OisnOnDZ3uLpHDDxZc1B7nXV6d/1LGCLYEDSWSbrLGsALlW0ZcrhUgSY
nQ0Np2UAUuHJNadf/Xeg4yxtRoJftHdeYfB5kuD3rrxh+NofXSzOlKGL/RUx
g9H4+GrEE6R+V6ypVAQz624Tc2xviTGlmGUibJeIHxh436q48uQA7Lm4np9o
RCug7/6bDtEvl0HgEOV/zub7thy5WyC1GJ6kiOZ9X1q1tCkLhhYrYnz5+M5v
RLiAs2PI3bSvN5L9uNK+6byE7SMPaaFnPdTgRZnwT2Mpfbp4X8KiJUrwzdBg
jD9DyH7820gZMIm3Bsqe50VCx54n+c4XLdvMpqeThIfSw9TVldz0QQ7uABto
eT6njgRjL+WjMtfu+gvHU6Sv8RIdyi8AtE7ay+wd6fnFp0mkQYZiFxVyDdPy
Uvv5BEiqIjDCGHjr/MblUSik2VPgJ2g4WaDNfI9Qca+VYAjlgxaosWZsWDhf
lvXQSauLfUibYt7ue0pRkVUyom5e+V4qvok5u28/nJIi/9d7JlbUlFNb3MBt
sXohX2AfqTefh2o+8qfn1u1b0Tn/vg4if/dlE20fDfdKhPI3KkCjyhryB/9O
4amuDS0FuYA8Vv3cJ/KScjaXdyzSXuQWENBpW9S+8epbwmD8RdKbXqNm3OD4
sdkGZOz4+TLqRXvKWmp8fa+5+hZSbKQwf4pxbskSBam4r0tovC6piQNrT9Z0
aMlMbFwNKeBOEn5qdmWI0oQqbtOYP0y5N9SGvCJE8jHzMAvAj0AU+RN6jcIf
ZmVak7qkWUaQnLpJd+AqU0mJpvedgdICthfdw/6bAKpYBF/91WM50X+cTcHs
7JOTjeuIdYG/CtHEakn5UEFNM9NW2/w+51moHoJwMZ5AozbkdOZUAB3x2gQK
vjtWj7hDgDsKkBtZ2ccdaa+8YZzSmDPExxE0yvvzW3WT+ca2LgkRE6c4eI2y
rEsOQP9BnNksIWQ+M3uvceLYYkwL7KjW7GmvLur2ZMvLDOtk+KHlumCIGvj4
RwlnZIWjRWZx5aB/hiQn2OIkLGYH8VbhZc9iRbQs2Y4EJD4E02BkouRCmkoM
yqQ/BOSULETg5JmELuYDSCSEHtelTfQ+o2PCEFbAU2chr0buT5nfg4IMCn6l
I/SsoDcSrfiAE4g8QGUPjbuKTuAzozMcovDNiizP5cFHfD6o0UQcqPjioMFi
K0wF9Rf73er1z7oSEPpRE4278/TT325wVpa7H2evg288UzFW5XMCTXrHgOHz
kxJmaJTL8t3jvwpvFmDq3bN1tnCWhf/8UR24wtOfCCGTh9NgK7y4uYHaiZGB
IbgGk+I1AV0KL9WBY/ObIei61i+mxZZDKRxvTRWfvpdocHCQjTWkIcG0MjEj
6N6FvValvzX75QKuWiQNa59uzkv9zODSHtagqF5EWmsksbnD5fi6NmoqdIrZ
R+LaobmULkKxvofMN7LaYCDkFBPby2mBmnDwcKtNfcqfyVDW2iZd2MUOikke
mQh5cS85d//LmFGZjN4stqyCw989BGTAP45KGFb0bwHCEBA6TFWS9+Gq/fk7
eWAq2dxPiFXzUBxEj8tWgDqkYL5EL0NHCHu5XGHfuab7vAzpffnsa9BJ7LsH
veiAYzz2aUP738kg/GdY/I5MBNHRVk9Toc/OHHs5oOH8CrLuUfvMqEV5Si7t
ZFXA8gdGKrbuJUkNludxZbNu/ladWFEd0SrMGQeN0hq3mF1CwEGaCJC/nQBt
TVSfc9rIRJOz41GOy2SmBkfm5J6sNJG6RbwvyfjOxPC4SG4dxn1OMUIUyZlV
inXlR2fM8SCwe9uccKun7f0omt0b4dSC1bCCJqQoQPx7F0Ew9TsM+T3C1UqF
UweJcABVfLllwZhIgjV5z31yJwotMHphLVrknA+9ZAgejZi/RQZQUwgQVJZr
tH/5w49ttdKEVnbUV9HB5gDKGJ/NiMgy/PF73FvhILfibroqzG0RQrjmrFxc
7UigfUMtuOe3amhrjUHPacrfNRmRn6NHZunRnQ+I60fh8vmrheGmWUrjW9vH
EdQuhjKJ0O6WMLKfCa0BMR9UlCuteK1Xnf67+NuEhF7nf02xoJI7b/cKFjPN
f/PTosay8UfNIb3bajgoOKdPAye2ElP4l4y/L/kEHrsKDgtPDcFiChF2Q3oE
eH+Jbzv/VZAivqHr+ZEharvCgQnJJ2TV6sltrecSu36/jjBlxSCGHNQpeXcz
j4eMkdvyhN+HG5k+PL+Z+LexCuIcP/Pl5OJBdnEM/C58I1vJUSMCw/ELsqgb
TPOAAwiVavXRKh/jeg+lzcZxQZXntjzIxulctRoaFvi8k/hPKZSIj6+ZY0Ag
ded9N+RpigJLrow2wCDR+CHnsa2Kw93lMNVNyPkMcL9XfhRzTflmcGhuIKgZ
9UqhZH0UtJ5UlA0MxyPydvRH1oQ2R/7JKeTsfIs6bTBKQV+yJlYgajoHbNYx
yATF27oPLuEoASbfL8X8Ks89qPEGshEUVFCKQZfk1XQ1CjT/rTDsL+JqclKk
nZI8Ga9OBI10W0aC9pMMjkeO2SELIA+ZEy5up+hjNsXShwBr/fbpQwxkQazg
nPhH5nlygX/UWdrOaOwVDbfGAgGND6X+H+5Emnzpr6u0lM6a0c13HiPLv7ME
jG3LETDAKb88PacKQfhGEFJWWA5fWBbBQRzW60DZ8edi1jV3N7dmtyVp1Go2
/hNDoTsUrgqohrWdx5MHSX/yJ12DXnAkg6co+IL75/WNxOoP1DHyzjenOpIn
ZRk6rE0Pg5zUZIrhS+lYhGKrWcAz8bvfVmge7bA9jcCBfT69t3G3W0nmsy2H
2xq6kipZoesqi/HS3ZFt97wm16V0EimE45ZsEASBxXgyBri62aOKWDv8SsQ7
FuM04p/mZ5+Vk7q7R8r0f+hOHF38njnqDcW34Y9rgLzzl/YbYcZzAohFqPkj
Laq1+hh92RaZsUuhRVfc6lk8MmmYQcP83juksvht+IR3jiW8YvWXa106JAK2
DHE/i+H+zVhUJhXy3I6TtadI36j6yasW+VvmOkwsOGHopsow92cq2AVd7dl1
SalqSLRriKERfe2LLWzgPa82F8iWtal7M1vPJOSH0use0ji18JZgEzuAsk4L
eWN1SJhx9To+TRy4U0czTpgcM+EgCFs0t6wqrpJhJVKGCq0vNp27KgtAg1pI
6awUecRzzKVGOLdyKchUa/jeYcSutSih+PR2iKDnP07Mp5U/lLrgLdGTTKyC
DwIo546y9fHQGGNmHRiTwP63cjyFhMhSU8wutETDUHEWbDS6Acefh50XYfFh
gxItvNC0JdycL7zynqhdx27/r4mjJgl/yp0puHuMSwRgWipZeO3qqk6Q1ThJ
jC8Kl2wfGGkZ2mgYaSMcJcQQ3IF3lj6nRM/2qY87YNxfqal9JtTzV7VYsGvr
l/ZT/Afq5KeFwd/F3pzEhQ/1MtGJhNueT2gBOoecerrQ/WupQhr7sAJrAVDt
cy1iQqoBHD5pjn9YIZbACY61oVbqy8JouhElgd54PwAImT+VQKXhQgPwK4gd
mVMoT/6dtF0u7iX3CXf8vasKTkxtwaSzUgsR7/0FPjVcSIciUltNXQeFku8l
zAfcOVXEm+u0LLze19SwwqiM4gxeEEKAbiip+ll5yBj7tQXum1AZ46biewcC
5B7honRXZxWEA28gYKcVFgUywKrSmU3+br8QBn94qGWEEXa6ZaJL3PCpPr48
mnSTmnWR2rQ0QCDFXIn/wLBDbmgQcHBQ3lfSNnYIZbR+AbvqO+CJ7xac3RwS
FqtB1Yfnw5MvylvzlsKJOTQldFSXLz/K8rwj6gXMUCfqD38NJRkpDxlDglla
bw6pvCRrtga3+chQ6FaPJmg3yu4gdx3t4oMaeH2h7oAONUwGI94Viv8KuTWz
vTOb2GgWkZvIQjNM8n0/th/RfWF4D9VRGtmLokoDWPJWb2Sm9jKZguBpCFyx
NUoWe8fjlyU2spNWqNQ1BNZgF+LuYbdfdJUBHV5i4uoU1LrptYR5g1qb3DjG
CtIN0OaJmYmgD30CyZ3aw8GiWMA8TAbvG72Dmc6nr8FPiGGCfX5xF/dIdTKj
2MO9E0HRIoPq90NtCVp7em0Qp6kTgArnBAFX3A+4qv4p8NRCRKP3QcklrWOJ
0HVknDQQ+bgN5mEzZ1bdaPhxdjxSI1EyZez95hCouhoKl2koX8g/o/JRYxH+
ThBYqroGH6VQcFcayQDwQ6Ufw0MoevfKosoNSJsXXBrR2r5Namz7/ARLipwi
TX5uw+yhB67b7j1xf3azvA6ZqrVxm3ThmSzgyd0AXZCSasmiEWxUAApu5fT6
NA0sWqiflSjzv/t1EXveMO3SgEwBcqaOvlBlOX3kJEkg2wKhrvZawTMTvKg5
K1P49GL6cq2BESTO1mB1BV+wuxsO7F/TXvv6eMGojeNckhFHZOgJcDkRQXKK
qf0ObW4uOsIErDQmA58s7UfaNAjZvVsxy5QcbM/PJ4iwzHesoBQvG5deB4Kp
GQeeZ+PhOqNFdCLuSCsWW0OWXM1ujOUeMiABlqTNNVifH+qicr4uqyf/Zr9E
6q4R2ahtnIZgALDnxWLq9ZWazEIquUGqj3ElOXhNU5nV10UltcE+IdPm9+dd
YTWKrcM11c9SJnaCVhv7Zd43hDl9EkwYmZzAT/DqIPPH5BmXFfIKxWjEWrma
DgAYtKQ7iokiDJEUo9Up42rEkLBaEGppvHwD9ckuQIInCb6m0hs3RAwHFv7w
aU5KyaNN8NBX0/WbsU3Nv/LPRFOcA8IynEgfSnrb6Gv9xdML6HmfYHrfEZqi
m2+TjL8ZTeynTjazp80E7G7h05nGS38ydodZy/JOJ3iczxZyLW7b5jkLrD0p
y3L9lqYeAY2eKRjubb5kqe9FEBqSrHCZ9Bv0VJo2RoWsXFiCAmTVkkI3m5UT
/Q7qXqJUCSpKhHBUmFpFNEXuHMLu6RGpA0crLNC+SUmkoHfXcJXP32McOh+K
5YNU+5Vi8mpSTU1hzChRYlTsDqu6Kl7BTkQuYR4gaZ/hIhG3hUXCBALXwCgW
EuwkFqf3Jke66IfC+GQTdPhn9uALWzCWk7qzLVD26tQvd2Zq2hUiON1Pz2Uc
g/lT/JdCDTEflBCdF3/DjDzq4Rc+5zJMzvJFyzQgJssRcm1T2PZirW03bxt9
zD/66DVvi6b+1mBQOfDAxBTkkt/m9Cpe/9rA5D7K25Rg8vnay6ZI3Vrv/In+
/1B5QNxlA+SQLlndSBWjC94QxmZOoPO0NwTZD3aPPvMwhPfS3/TQYE0tsf8e
Jal7sJr5TARsrgP1IYqUSMEp55aKE0q0I7iVLlBnkXzeG8psoP2L532hzBAx
UoXrLnZzNEPq+OxmKzTvsMeX+j3evH2edvj1oFxnza5DphmPc36ERMpO1srW
V12ThHbAvJyHU4aA93rwGr89miuU0kdenNcXuNfYykELJhvw4fA1/sh75uD+
sduiqqLetajGgTd2yvr6xeHAiWd8Rsthy62acjSOm+4LnZg3SYcGYNhCTqr5
oFEZwuaiPN9uvxzuuMT3FsnY8Wb8rh5jfDmKBA1VUqyasuHoYCpNfyv94f3d
x3DKHzN3sryBrBQGOXCkNDTB92CgaSktLzEH0eNWPUcpeqsdO0GqFCnUSeOo
WDDJ/rqaPxzGaH9/9O9z6pc+yOObcTA09VP4aVJPkeMMdnyNHcY7K2KtofG4
zJsWwLtR9BgK2cRCvefClSSdpUQjaVjM+WqxYXtA60hOQ8KQtAGnPjG6GaqK
fj8mRMGbc6WmrnBXWZh8r0YVZ1LUIgkUPZV3O0A33MYcoS8bSjZEmjQazXO7
Y6enJGiCjMoplAmMDLsrEZ46RHjdVMfmCPbBqbRqWbMwbRvcuuDr2+CYbG2c
BpMv9j6zKIRCBJji6u5qb1SK//vz6Bz5G8BOWl8hp73Mb1M8jkf3o47Dp5Rs
OaAXJz+NjGoQz5hy7+f1/ViUhHc42EHcbOe0APGBfEr2VersYJw3Ed8xUdqN
nXAXPPg75p6jdQw58mjb1eVGdMALgiwY4uNBah9+oPBmAoBZkAJiImtLE0uk
DX76qJwn5laSwM5YWm0vMlHHgOWBI2m9mcnbXwLq3m6FkYlSXWN5t7RE/+jy
UdTcbpswGywdV+GPJS0zx622ou2elwurQffaXA4z8cU61jRbwxH/DuBI4wqT
2oIMDJy5YM7OEV3+8yQQYDG1IGz5dMnV2WRaF/IX9lR6aT0XtMO0PUnuw04s
8a8Ilr5epM20ANuBjdcJsckxPJKvEfveAdTnZYgKp+GSGX1TFi4KLnnbfiyc
+tMcmOgbLjZHpPkIwPiTKbuK66FyQHiDJg8MPwvDBJjqnaAguDhjferePofi
O14TaOgXMDMGYVtJSx7xuNnqPGvhdpC0lUsW19C85i2x8aACmhSxfG6E0PsM
DhHQb2JRBhwJJFmf60wRRsQ4JD+m0vfzf7MMpinwb8+M/6dm6CjoBnQ/rYAx
DsVYnn/cHjSr8MW5JmjnJPafsdquCJdsbbcScWkdfk3CaUVRVeeCCs9m8VmW
fbbasnQyJsIm8SQHqoQ4Alf4vLa6zdSUvmkTdd5uRVNeRt1IvQeenWPDch4l
vbVp+hNNCl7c6wJzAVkyq1tzweH62Hl3opeLSx15bPZ89yKioLtKk+8mHDG4
joENHXN2wHQFdVA3upOtfjooXAAMNVowY8yCOFlzQ4Do9vviBDofLV0RcVUe
CbCtE4HOOb5vnZsrdm9SZIZuPu5zs3tw9vbSNMfp7db3uj8iqLVG4rnVty3r
uqGWhjAKLh4j9uQTTVIw7e10yianV16KCK1AGIKsgCjAd24sjVZsCiJ9ZILH
+q3Z8ptsAeVCgubEdVxroIyCVO1ci4GNIjW7Vozkr+HVgmKG43oxj4cd8d+O
E9r4hLqx69DLo+JVN+S1SV8whrVkVH9D0y/SYt7gFh1TFp+QBukcozZ8ibLF
bVoAI52T6TeYf/+FS1EbkQmKasog/97RB/Xf3mn7nhhIp3txoOEG5vAG84OP
uf6s8pm/pjeZOY0aQtXcDi2Fwh9kEi1SE6W+VAmTO2hckYYtmZE+LwYLcgE5
8TEDYZ1NXl0h+lCAw9eEpCqFGxGz+jST8QleiSshR6es8gq8j1XZQXBcnZX6
ESHhVj8I05MBUf6stGVVHSUwxD3rseruqQQ3GcQ++RIt+Nb3xPM1vZ0NxOb/
zZy1AhnBdFYqQ81OTFJk9oA9shRAC2LDRh+aG/GO6On11/d3dCQYZi0Y7OII
uMLyJ1V88ihwuH7Klyg00bgv0dIgU55MpDPdAUcdEI1DzNIIKD3KcZbBonOp
QinrrSMvxxOtRbdrZj0QG/CSo2wZ/pAykdDz/qAUTZoqp0KxJ0+4OlD2zUW7
ZqSmoUenfl/WdyanhpkAFPgp40CvgCjywu5w06m3IraEYzVKDPF1iSyeoFTW
MyFsDbpDiwsR6XajPoapsgnaQ+w3Y5AkLUjQGyANOaEUZb1nUtN89dnpJ7ob
YF05fDTqYO+F7O39Bw5KYy3srFCiwAWRGiIl1Xx+9oOs9b4isfLPZbfFk2rO
yKQ3LjD/hofpfvmkjl2FfG0PqEu/7gib4SvkM56sslPacotE+sUDmuUw2eHl
UU7XGEe/JXLysUgnGZfHVEn3ISBDluQbllKyz0Xty2WvW3TFtRCUENgHUl+p
1iQmSker9sr9mOBVp1xDphvkhOnJjRAOLMg/7eKd3v7ierXIlaVbuHUBqqwW
sFkxTjf2PZUS5zSzShYdOaMyYd87nrUEsrfpFfIYdpocMNtBAdfSrfAD3h+2
5akZsWZp01jAt/W9EpqBIZI74J3gAArZA727AGeDNw0i1WOtVvCK0IdB0J/9
OM9yKsoY6MZ8K5REobGugguUhMpdQ8HZUCQqsQvq0IwQ+d3qU4w3PhCWEc0V
u1hhdvTvkrASN/pSUZdvrKPbg3ENHznz3Pd5sCG416bo0uM2iNNZUiiDe0sO
kcfBfJCqYq2vFJZ31FNAg1a4dLgGfqGbwWF0IHM5BIw/N0lXHKZcZp2Z0HvE
4d+rgMoGaPuNvxACaDwHT2hiDQginvJWvlF8mZzv5Q48so/DsNelx6r4nn1p
q0lG2VPjdNJ+QIZz7KHQxdNkO3w/0Gl5B40UOsCB9PuvfewYrMHNNPSMYzyj
RgJB/Wdg/H6Q8S9FYZu7DPTbQSw56aonbaE3/EWORrbbiyVcw883zyoFgy/b
kSGONR+rsYr+mPK/CswXA1X22P6RRfg5T1XbI36nbv0DLGWFtj4fsIZ4TyDM
cOY0fHjeC0WsNqfdpglKb8/CuSFDRzC6b23jh31ZP7PSt0CZ2CWiXtnaJ3Pg
p0eJLLVLu8RTl2TG6DpUQxeHCvAdtyif3KHRavtQBDv2jaT5wYeFrpuahrWC
oQ2EnbebTRzxdQxLwaQPYnC4GC1B5P7MxoTvV+RBjo3SDm/8JJfsuw9Kh1Ua
gnLlpRUgXc9truKZjRnlpTOjahtTp1JYfArDUmPuUEBrqn33I1pWNezoNKCZ
YSCPI0pqxeuXdt1Fv60qxVyTPMV6M1yDnpZ1Cu9xsPbeAshUnlSsq42df2ca
b/NBtfNToBGag7Jk7NR1VNC1oNIJe/hVqj7MZM5o2yPfT/2nqoLCBLruSmZl
3jcA3mO7ybNgKtu7t758U+NdpvJRvFPFeSf4rFJjgPwSqV+1DafWB4pQwGGN
fPhBm4/INUOTjtMEqK3jKuWJP68iOnG83vzLKus2jFNUUYo0UVc4GR1eBKqS
gABIA6Mal3lM7jCg2gzFendaBmfcQnFI6FN7N9qDEueEy9o7SB4r81H3wiSH
71vqOzlMdNI/d8VamKNZmvhSvYutQiDFB3Q9Oo0QgwhOUomZIOsn/tajr6Ip
ldUze1bIUcjcvSEyEMuX/WSQAtc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpeg6T8TGqvSw+z96s5n28/+lazrR3cjaBu/oWEczCwaECvC7xHV4NN4BCf3iTpG7DVpF9XQz3pDW8FdlJ2tFBvMMDVzXI0GXHUbdr6knlwE4bJg02dye8uRinafYVWy5D1Po9Db7hIZL+cDPpzdJ79QrV2tQ1SsFpagrkFE1OOLcAXy14IrLIRvcB47N0e+07U+8HJ4tozs9SCsGDaFOreUTOCxiJ/21nnfKfCKLUXUpQ8PsLZ1NlhqpDkyI3sX2psoxKqPb9wdfao9oV58ztKi6zj4TAzCZIwitM6A45MTrUu98pW+KyZA6f5g+Q3PIAmmmtYVwbq0EMA1jzmdxwDMa3d2OjcmPhJAKmF0YyJiy2Rj8dGGprWB7qRYuXOfB9Rc1BqJT0xLEWakVtafaMDEYHyR1Fo7+bIaKlN4+P9usxP7d9TsjkghPRjgn0PiIOCAC6KKcYo2ZT93RCHmuxX4MoW9dRJp/skrH1XRZKxxbcjbA7/EHOrWGAt2q7DCgpXlIk4Sc0Nt23yqFzexS68xpFL3Bimh+ohsnBv9OIiPeWa0dtUBnWBOCWrB0Xk3ZkipFcKbTu/qrbFlDhEfDqFBqL7rL8xtnWvZOqS5B825Kr5Pe+sa/BTkDrfhsx6sgAzsASbK3qpBckSGZs3QTqGkUfPmG1Ep3DuTLAALT2dtvzcKxrkc0BN5rPnFA7NZzn+uwnT5i7RXuxXyYDt3bJ9PR24ozO+UQ+7XdgAceSHLQiqvBdwIUgLRP90EWuD37J2Ld3njoNGt+JhdF+ZT7/EuH"
`endif