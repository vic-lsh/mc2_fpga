// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iXsNNxaTDRKrH3cLasHiZH+0BvNDsliQYt3FE2C1aESGt7Uxk1M+2z6NLPjv
VQRuIqCDTzVTM4pvncgLV1adIVP85DM4UcrwUo/YY0ElShOK5LLMZ0Gsqc5z
VMSP3R2e2frbXlAA7QkoaDv2eYg1weeXAehyVsFke1dEXg6hd0csIhlFyr7n
Q7Krri5ZZTVVwu4vSlbjvg5K+lPxDEJ1cGnj2e/bRMIJ55rEtLX/AR/YTlIC
UysB5U62Q7MRsCpLE/xerm7p0MMElbh3HZF9Gg/t0daFFK3s+Y+w+u9Sen+5
NLFJEuZunTaTWhGzYM5kZJxGS+iu+uKiHdTNyEh2Hg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b2E8Zi5fYQG+JgjSm33eGcOpgHukPrDVvLpBppHqY3rGtuMD+hk1LAQEf994
sW+doDiP/zwplZj+q5Cru2FGUSNOMm1rC78okncQDZfCI5YSVTgv6lFZ8ik4
LqSv9X+J62wgSsryZXr5SEau0rusMBVICUePV6PglKBNeeXfglIsDQ3CUKe2
Z1eABvfFuZ23UGURkpEzxXMnyw8rQMVO2c95Hfmbn0gk9JZs6pIfU5bGDsa3
q5Fi7KmDzU/o0DTTvImpYoAOYN+3HnHcQMRtIrIIyzHBC2Q3M0Q7DaB8hp4S
QnTTiR86l0PmbIWfsB+f4kd8k2p8jmKmm/NsaH9S7A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rydanxyPeRfZTfJCe5zBI1BylUAMd3PHywRJknA9svIA3OH9NLQBSZEXxpx7
UqJr36ww2iD9HHR02nyVz0zK2oTk15QIEAylsIHP07hv9Wtl/jd1TBkrzPjf
PLFIYEKV8rs3fKcA28wIkhsOWeHIPWi1dX1zmx22SFp5XOuI7zHAc2e7loiW
xg6+bd3g64f3Pgb4Ib5Bfg2kM6bRfS3Djk4sZYeksfebagusCySl+D9V68Pe
tAn0CbmKx8vDldaV9U+UR4rDYSunttmfnQ0jxqRLOUNBuJkuu/Ygcm0hl8WL
rtX5a3nQWiFbLJNfW26ukV/lqLZ5jUDNgZclugZbEA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UAZFEb9oPXRBgVI3/dXYyTVgnfzxYPE+b6AuUMGQL1g2BzfUL/FMr9nJw6Wf
1GsWdJ7VBFRjOFREWP/4+lHgwngjyUVolF2cbfu9js0R6HTmvCR0byhOGWZa
JOHJW+ozrPSAqy87fLvJjjZnrbVa8EsIRnJZ7t6cjKfGDNmy2axYRIwWI/uS
YBg1upBlrxXG9lNpposSfo4ZPOOTm3+Jw6Y4rDHUYHtz9dLf2520/cFnmQYF
oXhgM8srOSNEYbw2lGYNbnzO4UC+P1fZ0NvXavIvYkgRaDweoJmeuci+Cgdl
PKzu6vUe9+IvdH6fWTunFXD9OmVMpQLp4AT4V1UMHg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gzmTuAVmFULYQ0PSjLN4qVT7cammwRbE71E57xkVU+aAtc8TVCwhYzwIs+uU
KZasEkgE5D3jsytWlVSq+NaYFoze2UduWb9KPUS3itkdq8vY33h5ru+nvqx6
PCT8C77iTXdiak10aCXEvjFGc1eoGLP7UHXpxoq5fMliQgX06HY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
l/ZuhEyKt4tj9EZvbEDQPdtJQIABg/qeZ+xsxOb0nRYOtSiGsc5jioPj4V4W
1ksP4ldGP/3SbP1GTE045d+paJdjafpwmHfVmyNHMj70ZRO3LiaQinsFOFk9
QeEN4EIFnFjqqtTfhmfl+BhLsgV2xjTrZ6B05P1y+78gK45gy4/OGr0sKUk6
tQzSKPkNbdRLVEebZ1VOonsnvZyoiU8cgljjJltEG8SxcKpylpZcZB/RgfQz
T77EtPE0fZkL+loYs+bwzDem78Vip042liaC+4+fWVUq2ESbZVyCYiZWAODF
M4UscNxJbJ+mkr7ioPv84eX5ayy/v44D/pp4f2koy8e8qRdXjGg7H6mznYzW
iajag7UpqlRQvWsqnHzVqpdSVvvfF46tc2rVo8pbWXTMuXg5J4rBJUlkSkep
Zax8/RhxooRBsqas5RUX7NMAdXQ1MANkaVkF9NKajDHTNbFcR/DjEAyAByZE
m0MbUHFgD255qSu8CRjG/5KcpdnBgxSa


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DgIHCqTiXE4drXOZWvycVCEtT38TY2qpyMb+PJZ7OCvlVaPD41mjb+9FROeS
UevXctBI+XHaUd2U3Qv5XzMHAn6EYOkr9ZzjaDrd+15Uuxk8MrNfLwLeXf++
jxg36CEcuE1rqPfy/iyGe14lrqbVmOeCashfPwDPtT/wD+X6+3c=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NOn0GINmq9hzbIVcC8VeYEV9Kxcjdfhhm7ih0gThmp3s/rEtf9Teo1ypqTzm
UWxxpB9JxwZyYFlMfhOnTdzahDheyTNpR1ClQsS7Ns+h3SRu+DsN5wFf5tnA
G+gfha8+agt6Nj9fF6dTuIsKgt+wFJT9ADHleX4mKiahO5O/ysc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13248)
`pragma protect data_block
BEwuQxAiOYhC4lDjLj5ARjEwJtIOAFPmxb+jfRTh7fHYJpD4YX0XczvlLTy5
ZjMXkiYXlz1ZEBW+8rKFlLNB0hjVwtWMDcCpgLMhN+6mL7D7iUZReW4jXhGs
yZ920PGKdX+zMjE3Au9WbHR8nRMsEQ+2+Zt5YqBQsJsa5jV6Bhr9AWSkyeI0
PId0cntBWLfJ8llEhnsQV+2ldRhwcS4hQUmlm5Za/ikTwSNiQ5xXwoJyF7E+
/GK4nLMEPjVMan4X5NCMhzlaJsD3poS8DDxCx2meKkTyC6XtCmC6/IYur1Iz
mux3rST4NTxH1AwAQGeI+TUERgWpajTMayExnZMcq9+yZX4TgLSBkZgEd754
xqALWHENIr9Asa19G/LHz3iN1P8npqA5r6GBobGCnHGIGBcIGQuFm1e8fI5i
Z1gpZZHU+hfB8H89LPgvMENIM3C9r97fdPqrzoC6QT0z5KGhJo9dK3ONKrMF
pMJ5if6hPVudduKlYH7Eu93xVwoyjsvaaU0gFrVRfHUekL4SQ0jMnXYjVjfX
V+4hOO6l7hnVNuTACS1l5dO0fSeUGuGcGZ3Fd7wIGQseILNVS9q7GcRw6u1p
RIBWpl2aqg1mbm29VlIwSIiJaRXhX/hRDHio5MqSn+sBBJYLW59VMQ928D0/
cjRYEDzdg/agCwGwgKYCm3ytNX6SKnUh0ikkewZ2cfJlUJww+CqtzBd+EGsZ
MMeZtt2/P6TbHcA4LoOUEXD8tgMjmtGdnB7lbqF1K8YaQZaBC/b6KR4WMGr0
4Jo+WjyZeIiyM01QllvFSPhxMnxKxSnhPsDBmujW0tm/A2qOgG6hMCD/yt98
yfbhZ2bLvCm26J4wfMA2b9YBI5baJJeOyg0Y4yD99mgL1lnjaNzTK17W6M9E
rtbyzZ0dQ8U178AdtnOvO+a6VA5iRD8ulMfIyt+9eJTuA1r6l4NzvmD+FnCR
anJRlAgxG+YJMqRDQHMmD+o3/bdkkg/RkTvNVTU6491YkoROUxEs/2LWE1YV
fLaJ5FOBc70sfyGUB5Am/wKY4Ixlc4GufaElM5JESLQv9V2MvCFZiNPoxrXH
AnihKeAyrcmJE6yipagifworgD6Pblv3l/26TXi+QRXVfjOC1zYIS6dSk4s9
SwdPWe1Xl+AgG0XtyavVz3mwjEmZdBUn7rVCyPv2X9ev8xi4cNo59hC1D6Uw
aGyeIybaXT5EMzba8IZTwCgvrJg5ybmfSE14t2s5oVPpkpLTNpKhcj00H8Js
vueATbtiIIQgGV1pwwRW/sppIdXdz9doASt2CoMnDZf/ml0nu1dDBbg9u2hA
q3aFOHaMKdxYsrfCnblSWtwhkQD1LarAsbq4sHLr34AnmLyAE4ZCR2qP6p+M
oLKySU50byAke2m1sCfc5kmWs1exWMjmb+uQxwE+gW4U77pmrsCxaebaG/VZ
CSpP5eWhrr2xIsVGuNmLDRFFIig9LCaJiD8T3dx46JVqKC6l1ZTzK18s87hK
LUiKGpwvjXIN2tMKsUnNOEf5w8JWLteelbIgPZ2gZ3RlZT8emHiIxF7LmnNK
fudu3KUWRNmksf8aLv392UmbGRQalhopIiRZle3AB5/Q9PR84+KQdiGRDQSm
58rdhHUUKiBs2WMsoRkJRZfKD5yD18L6XpVJ9SKhf8QIfBC08Z6m2o/orlvO
hKl0DxLIScqPyOYS7ZF+77ol20Wv4dCHbr6t+3ZqfsiB6v+ffFtInqMt/Pjc
H1girHCwPE0l7uqORp6m3ygo86f2Q1mqCpWafQBorClEuFm0RljIlrYSj8nb
f1tZ5fjegUQZbNCx6pgbSIOXEuCHUTROt7ZLdLeuUpQMUzR4mJl0LytZKQMd
EUDVUTjEGYyYqgCOG/gUNbe7OQy4BC77dJChJ/Jsum3imHZSksFXILiYZuJj
kERvQsZUZIpy1MrMJ8xNtrnDClknBPrqwNP9W342+BvNBrQG0pSZgriJpnHG
PrDkYpa1O9yBYbKYm/94+ynf0Cv4PVHD4AlLc9pqEto6Y7APJ/gisXkOFL1U
Cna1BuI1mDzkX3clOrjBiVmfq7h/+2aDMZjCuO+TClx9WDLjWw56Y6jWnYpH
HbriyxUH20SORUCGEME95mIj5RX+xgr8UfoW17t8Dd3608Dw2Pbdg0hZUJal
+hQlM4aW3PaCIb80Cc5wZ9+QRGcgra0L8HR9ZJXbVxmtpM8xAE0gQRkDwnE6
HIq6bgHZZ6JiOYol2eeZBKFUH4/eueoEqZH1+g7lOBorXshJNRh1qlygxpg+
pUCAD8OsQHFbi0pfWx4tnDys4RlQGILAOypbL9lfJZCZdlJ/r92/reLI9bM9
t80gdb13OvMY1qfFAFxAb53lxFbuJ2K0mouz3MyobOSOAP1mnovCXz2TwR54
KL0X5kdlznGFdvq2ZGIK9blfvX1anfixbp++83/SpxR1x14JQ11bRXUFU3eD
mRezINLqCJ+ROhgUkN0PV32tqjNhBD9sDBYuy18Gt9TZ0IaqF75n6LSa/bzM
3JgF37uug7GeZSt91MLnFacq3lX3RDxAy7LMu3X4q6cCJcTsG1+v3iKjWd+n
1SorzL4rGg4BNMk9AhfeZL6LTWsh+qq/gbPlMpbzAQZ9PLRw6x7jAEF16Wow
RTLCTJOKrGTB9DVpxlMxEJddM+BlA42jOz+u5Hcy4DK7USl5WfVOLq4l4zI8
unicI6QPrTMiEXMdUiH0C868Qqd0rlVYev+0MCgv8/k7nihaOQzcL1wIIfiB
Bv5LxY14/FCvY+O3OUWlcQl4DL2GWpAbakq8/2K3CyzR6E3UPBxku2V2JfT0
ttpWuMV0DieHY9m+5+cmMaQjPRi26qD5tqb209R7Ul6G3C123lyWr/m/dv8P
CA9f4zlzcs3q/eA2KIxDIEgiStE+U30RW8q54wFVFU8mqk4Y06+sJn1WAMpR
maTn3RKheFuuCyZln6wTpZQ7r8d2hdPYXE3qwF+aizNGVpD6VK7EGmL6uosu
UoFNAx5I6422c4bkRldXQqWCAt/n25f5Up4uQKEA/Lj5vhc6mg3ob+TOl48q
YBq3gCuIEoM5eA1j/xhsMOJMTYvTOg0Rx50+jFROp3fVAlT5/N9XQek4SjFF
kt3kYLzC1cTcdk1f8QpXT3g5diDT+X/4QS0Wl5P642WCNf/DadHOpldYg5Ja
DkTvBRtCqIFbus1rxwj3OfUOM+cjt0H68sm8rOElsX/H5zfvaI1A0G4nrAvN
NgQJ+sY6uPDGuPv8EWtgX7MRk3Lnul5MDKm/9lhbuYbujt5x6+/VyukUKYzW
MoYGeXzD53+6kDzPzdxcnBqcBi3PkU8cBwu2AhThf6eNOjPAyK6LNwsI1DF6
QqePl4L61D7rOuRyAlyxi8n0CVh/HN7Pv3lYkRy3mrCEqwY/2X1EWlS9bRo1
9sTNxjNa8u0mgNFnQH1el8LSHqKea+LwxSGg9BZ0Kklrc3MD1AhO7naNy/iu
QCh//uGIlEJgwAgNlhsoTN3NvaJoBqs8sITQiTRJ/gFrsYSOmdwV3roD/s+H
BCxcoLisbehNL5gt097YJwzOyfMHHWACLVp6yvqEIDMdcDs/YCKUtxt8UL/W
MphHiM1pg3mrA/VmH0DZSTaiYTT/xExBZZdnyzAQyZ2bcQoLFkNvr1yKOhXa
mOoyfI+i4oW+FxfrtT9xdyHle8X3eELpC412IOneMayB1uL5sKRjOJ9huFir
IJZdQX0suvGW11hVAWUmidMLp+IDRHdMN48FIbQsl7z03a9rXkNlDqewOdtq
vSAMNXrygMwEcFS+N6VTkxtuAhVB+ezMM65RfSjfU/zfzZOe+ZUtmiR9UH3A
Kr+CaQTMwrj446b5kRiK2kSWHhLBNacu7ntwq1dmoKf27VNrxZcIy/xI8Tkc
KMk82HRUYJcws+StpZZId9EcB3waCXDyNtuOo4voOLYJX9KqIGakY29Kpbhd
TGkxCXD4MThhOz1JP9ftz7a7pPEoYjaZEOfWvcf1t2B7Xai/FDWKTYGYoieL
AQfcTJ5JI2fugqHIQxfxrhR5X0A6c7/PfukmJJ13F9tDn67XKJyKXFCjgVUi
L03B268a4FP+HimrcEg9Zi3fLrGjcN+e7+XOrthrp1Aie78DhG4L3GfUVdom
Qg6xxZ7aJiFdj5oP8LWFVTzrhNGhvwZ6pz3/mXZYLkRJGmp81xoARTM4Jwkr
COwTEGPgGTzupoeHwhr7tjVlF+O0+75/ETFC6CgZ7XQsbcvSVqBD2tga9Oa+
2yZmC/OsrY4G5fQvmWlBt7Yf1Vo+PJ1zvpA+c11xX15T4ps0TTLKHohYhXQr
n1zx9LnpObnpgPJxEVIvYKoslsKfxZH92VsI1pqeNOsgr7cQAgVgQx1OvK+U
W62phOgdmIwCU0qfCBhOp9ZkBySom4sas9Et1Yrgrw/kehUujF0R6hlTw5+j
VcPeLNkAJT4G6mm9H+ZOESTU7uTpTXqdZt442OjybteLcX/7CSlns+HpxJ5q
/JvYFJ/Pq7hqWIkF22ysjixog6GWNADP7sPQq25KofXOm8viUiZYL5JguICD
ZVnhchwyzhdAda0t+3qwKwiYII/6s//v9FsT0jDQXzWCupgYSfPk3JH6c8iX
cKgMtNgew2LNZiFLcBs1Gma5a/19EQFy1Ijn0K23x3ug7mdAnVNtNNMnCj58
/vTpgjoky7Hps0AbjPSMvkOrWMWiE3IWct9KPaxaKzRuKM2dbqGmCsl34DVA
OO1qC2n+tNbSKdK3xA9IKj6sBGVd2qVbBewPUnjsoP/nYyLZkrxS9v4Gn8cK
BUr/KgnjSmQVQ/K25qfIglMSVTcGo0cA1yyJFoOGkmEv7PJdNBwf0TQPSwDG
TaH8smLlX7sRfyA+nwvOCdu4tjcXy53z4XrLu8BP9Y3FSkIaud3RtlfIPDPu
luciAx8hHklNKy9bmRoV29/D2nq1xHjP2JNtL12RnQ87gU7Zaqe2EbenZfUC
a7qo030wNB9EWHJaMEUlL9h3xRFfwQYAM5SimH1TxqBJZv2LwUhjWbSBhbgC
G2o2d66BI/yir6Fem4GtUlMGrgMGoX7HwcEBAIhe1X/xUVXWykcsaUcyDJoN
RHLKaH9svE62Tt0dIeJkddpTwnfXBi7tT7QoNnuWGTCAHzClTazFswd8v3RA
njekhX6kW+pKRcQPEPPHm0ke/bcea7u9kDWohxxN2zIqUVvmbrmnUd1d+mnJ
frjNgUkqnAsgKSQkLtolJrgl127OATzxmVRvwccuK25m+BWBk9InDuMYVb7q
wHouBIixKPjomDOahtrcclT+fprp0GYewdTfvMizlJLwEQLJHn3s7VwITCag
+Ok5QqiH+4sqR+cHDtd/8Rp4NqgmXLr27WVjMnlcy3s6jCm/9ZpNzp7LSyJ8
40kekE5IXHonUuEdrqkzTkhadUxAjEhNyoKgPKwB168UMDGCOAJk5IrIK/fG
EFT6qepneUH3GWPODN7WtCYxP942QeORq2JvUI/e3McLlId9Czdz0ENRF7l7
++zFqOSLVwMalqP46Y2l8LtD7Y8/887M4DxoihongyaY+Hc/wTU/gewkATWp
uZMYUboUXhqYclYxwW6A0be1N7GdopXoPCtyicLfjyYKZpmD5LTOySY+0AgH
nDvqT8LWBEhJL3ZPACzpeLdZwPqHW0tqYtiwq/RW98BwlndBLBbf+6wp485v
D275jO/Fy9ywXvCoHDJ+KgWIitRj/DHtd9JLa8ZAFfEEFS+Xq/29b+wWBGSr
LU8Bydwg+bgfKi8EkZsCwcdc6yt8HYJtsHAZ1cNuFaWfZ37Qs8wPe7lv/mYe
s+KUMAxjvaF+SjKq68gJOTW4WkWSmuWg3cGP4vS/UD8ede+lpXsAKnB1bv1h
jGFfaiZl2uN3p0w38wQAabdwnBGSrboqgJQ9uwX0b4F9f1VyDMhPKqGsdV2p
MNHkD+3F6dYMzlwX4a7qkZpYf2QQ9FJnjvqkTdAvsoXb/qo2XA4ppJ9tk98q
BeG3COAyXcx1ZD599iq3sSuKFcvUTeIBBQ1heWFadOe0Sjrez6JyW3g7xRQy
5+KnPJ6khIcyAx/f27D0YLOT9zRPcCX2e8gJrMIbPrLGuh00EiG30fyzN3pD
KPTe3LNNzkMgd6LUIuuFNuj/x6An2ABG4z+5CYOUJF7a6eTUZIjR3CJwtLCE
zpD+x75jxT7IBd8eIUWzSJL/xInEnv3pjn5jJl1YCSTC0SlNuS31uSm9U9Yq
m1cShQs0n50tzqDbHkz4+soyFA1sthCJYCfU77ON5ycfF8Ct3jnxZoBd4TJp
AED8hWPjXXP72dg4D+cFL0EqQWf0D07S0yNBbnIt26JroB6K8U6rT8mcED/R
omfVZM++fzgYO1S5bA8A1eJIXU2elmzoEk3qYeLDjdPIWMBT2U4t/JlXukiX
a7pPKpF7XCSENffkhhNX6I0x6hVpRDXPgJAT6kJKExuNFQ+bwy0yZo5+SFOm
DMQiJe74vwWj5pPE+bSus9mi+NKfUhq43Wbbddr/alOu+zEBpenX3ZvVaa3n
dT0cyvhwUkQ8KD22PXaN5GbDry8+Fouc4/YlZERNVmD2i6j4XE4XNULdp+Wm
fq/Io0LnasF2BuBthqAnD/3r0MoGKhXyLmu4exhIfrhTDWeYNGzhj0PXTeDn
bCmRSHNAKVpb1nKsLZ2z9bc3SLaw11MohWEVNw5/3mv6VH6+A/p/rf5NMGPh
WlPnIxw58Wac2Vqx2myYxCZUE/UilTABCtYzDdPk8Yqdxp46YN909doiNm9W
yKXdvPztWwrjrbYRr3MJeEq9srGd3zbxdZM2gbUePvXdB4tVsN+0PXvOVJFF
oPzftrdmJruo3SQJT+tCl+VTeWq1O7PTxJaAob8WpbCm68cuXp5PEqgfaBNN
fHpl3/2y7qZ7OVYZMcypO2YWLWC8bhnLIpunWvr+MUX79Vge7o6Y7dbMMGbg
707h+FHbIVunZKlfAz9nFxU2rjYO6mJOuZDU7cRLmKOs1+p5wI8LQZKwA/HR
lglS2oIdII5FF8KT5XKIwJ5kXau1am12EN7KHozJE0338l60frUxY4BTePM3
7dsbnaGSCA90JC9TFXxIPkCf754L9ix2Qe+Xzz8vC2lHgUe0JiSXW4VM+CFa
dlbbco1ZF27XzJ8KQE0kJyx7SiXZF7aizHO98B8o56GMZE5AQsxBMDBkzNh6
Vk8+lpHsR73HhtP/Evo4aYDAVaGy0NiV+O+Bq5CkqwuvCePUXlkL1JNEzcJ1
BvMe7FCYVU4kEVstF7vHMVEOm79Vl/0wVhYuk0ts0I7H0sMYmUfY/c1cCBKt
9hAosRIkGTSLK+YJiqrI4RiKE8a3kNMJdZVfPLvP8QS8uV5CXJ/JLnG9Ga4R
tWtae5hgB/DpFc60TH1Wt60TBuB7xEkThWfcQBCQrWS1uAnm6hfgMVSVqTZs
9zmlKtbMEeOpXpgCGbsQ5ccvftfHU+S98SYpPyFARwXw73aNDJntt/lgu2Mf
X4ezPmHa82HIWPT/j1K0mlvzdECStFxOqLocyiJNTbPBlTEiO7YqRzSxwjdF
ozAI4r9IT+qnQFT7WgS8OpIsnx1PPChmDYDH2KAhtwyl147uvLpyRzfFONs8
5PKJB1SIXn9Mhfi11rp4V303SQsehz/zmVBaLrzUi/iTyC19995ltlfZuKaB
xJWpzQg/xzylALHdlPqUezRinomou/Ux3d+4hhMdSBl+ViB4FFTrtqIu54iu
N+ewopvRCHr4GK41k5pfjhVvVclgsaANTFCR9uW9L/ezEgzNMxtYqDf+ZHHW
TotXaJ94iMYtT8Kj6MWgR7exF5uzcAoWYHBSNThWW5z5qhG8M6sFeqgQvVP7
v0UvSv3xDoX3N1AhbneghPmpQLwRMRYdOe380T+pSXlEjdNaerPZrWx7D11O
87ZbFj1YlRq1P+zyon0mzU/n1fZk5bPhxPolvxipuSBsRNTErUnGaAMYQbMW
HR21vQ/sSHG3pHh/HQEU3QigDy0MIggSz8OGkZH/wwNLo1uDYgw+wkJvhCgt
3r7ycmX1hsd1AHUSo2tgo/ItV2tDQ+uPGbETD0cKOD13cmhSX7xws8hPRDHM
y6Znwu965IlnLxXMYH0qdutUrXQRcGS6oSM1ze7wFI4OoErac1RDdCRjnViV
PsRn5r0sMpsjkdVHIABO1A9YufMgCmskpvEpfRwgOM85ljXmMRyg7rCUTOrw
+oePXwmBi+sT9afdSoHZXYcyP6O0FkVj0DuIydYPViu4wNoN74kDr98Y7Vwh
1YL9Y+pIjRLTnVlYwDYVHA8G6TZA5/lhnn3tTXZhGixzT56+Vkqc7FzWC9sK
kRqMhGp9BspxUQTYmJsVSExCkveDevv3V7ppHaH562Nzlq3wxAfpSGu3fyul
6tHANVokGqZZ4QBHC1g43FNpODeZ6/1MPnLPKdrBt5zgpkxN6PFpOrJWCrtm
XN+3aHKjQrv/Q+88TYIFmSGO1SBwKxgI677s06Gs36p2ezKbqfy0VVzc6YJy
V8/bA/D29LdA0nPdgw3sakIWf1ocpnLEHaIvf4kEmRJYTo7O02VHN+NDImCE
qgevbAsStGliaNCMO6Ot7R2aZpov8JW3Qks2Blz9uukuV6jb0wUedNNPNunx
wiOkMc69Fuzqm5t0tU6WF0MgBW6+cyaH3v6S3jU27FI+3Ao6rWFkAZjON3tt
+YRC4nlPvnVlqt3WRzJAZnbkcB1emdXlNUM3luFowV0FxCU0B5YB+LPPuFGb
enwEiHPtYcGrVnvaDNKLleTeFKJ8BNnD2sRU478wO5CY+RVa2NlTmeQN5mhj
YikOrh8+c8fbQVetykH3NHaHLXdhYAZQ2kIvZA5V60NEOvoBHvALTFZCzc0X
+t014hGT0WpFNNK16VPgMY1Jv9YlkjM5hRY6yYrdBH9/Yyd6r0I2UUqT+Zvg
pg2I+14SIZzYxVUmKTStlNWSBNTFK2ZL0cuCOfkGp4BGcwKZ8dvxdVmLoBJN
2Ri4kErCNb4cgRW7d18NtgjwFA6WVgkAORXhS7T+idD5RemoIENJ4tUFEtsg
SPWvv5g+lCM7AgCaCkasTBuGOjjCpgJoeWduUtkfBd56nmSG/ZkvYJAAzUnc
1I6oSaNJb1zRq6ByPUOl1RN2ms+sF8g3v0f/RqKjvYH3+2qgubi/tY/I6QKM
NCfI2fGtxhtVTadldwPmKkSVXIlvFrUcsDBMV/w+YzIDwZ1NrQRFHCIMkj+E
xeQ8sIWUI+BLiYi4XfBkLRv1uvYVHc5yE3pdS9xywO1drviHEt4miWyhSCeK
xxlYtzBFSyPebknjDKZZ9NA4YifipHlYuazp5U7uPZ2FzwjAHw3HUrQxKyB7
ng2X1YlTYn4UBT+Z7HpiF9ky1PgyuU7LpEmP7412QQXSAWiV2ERlZSjzV3D7
fYr3kMWEj3/MzraEg0vcm1SoDC0PI4AsvztwZxn6VbvrHYIiyDFiFibp4c4E
OOrgvz1t/CDkve4SRFHrx44Fo5W350pivWgHrOYy8/41r8urfYd2E4bzDqKx
RAS/vNDwDPVcbTQXSGUl9/lJ6s/n642SEgXbx5tUkF3g0i3wrCTKSmJ9aqDK
E22gOClabtYvvZphuMWRygaGWULoouWQ+vOKVLlGm/ztqJGWxuNp0PQ4W5oQ
9hQ1QIRbDo8ygNJX+1OkJlUJ4cYWsbswFKDsInGxfqrBP33eyKg7OGO/PNXZ
Xye/2JkeJWal8BgqB+G4oBczAB2GdvYjbTfw1AR6uagj3H3YdRuZnk7ip6D1
CYzb3bYSabAtkREIqjX2ZLwHB+yslnEDbohxTF0mNLj6g2Ri66t80HFnJQEd
SIGjQY5HTD7Znz6P/wr1hoS74LuWevgecjN9wL4pLoxyyO1xqQ8eVIJlJQU/
FU1eei+qVrF/gqz+OhPnYkNSEmC2iol+OlORw5YOnNKgCza3sa7N+2uWUEei
Mq1xPmMUIS4fB6V2yrSOVv3iiYB+xP2zkjrfmd+DBC1NAQLv5bG+3gnQipvT
GJ2YvMqBXFF+AnIFB+1mGt74x+w3UAx7H3Ij3P66kZpQG36VLJk5s/abGc1S
zlwZ/zVq548dsmkMcD1j2vI3z4aP7yKHMEpVrKAzmde0PLT+kYJ3oH72k9h8
2+9D+/C2zmDbBqxqDnVEDbdbvbDE1WEDlaAkFYcSTnAfuU9JNrHUhL2TY+MX
uRbi2lKxRfuw2BoWLZAAjVNlNDjfZtRALE4mlRQUNCxJwi0yHnikveWLqDkf
nAoaXVO3K+cCE/bbGW5ZKQ4aLpgDLYzAwzt5aL7qn82K+Dougjn1NS/bisa6
YLbbjDoFl/XJ0RE+Dhu+io6Apo3ItK0aQDn0XAmhgdxCXrKmT8Cd3nMZrutq
OMMTIqLWdnoIEhlCRol2s/k+ET6YumkVRYKYatDr1bJOpzr2dGwmDW8jQAU+
5Hg19tVqZtdoL6R4JSahaNInQqaFGAkkoZxStJZP1gZa8rLeDfSWJsjhR7YT
5BCrwQvvYLr+RolZwIuKcXksrkTah8wB3LAnxVm8gWC4FHdgwXm2XpLbWxcx
e5lPbC6TYJ+8bsSDhx8buUTiwQgaWGBmJSwM+l2tt6iRKaCDGe/MIQCNm4bt
s9eYx6l7A/dN32pSReN+kXZbrfs8pYXeCQhRBRlX6dFkn9QaK6WGEBX1S+o/
+PaGJCoj3Lb9khaHGHIM/wqVM0tDSD1FKCaVX7MCxIozWtU1S6IU7RZf6vZv
jnVyMcYue+qqJitKn1UHAOo8SI3fnXBvvNAaVJfivmloAXx5QFko2yTzm4Gq
ObnW+f06KzOXnCXW3rR7Q623nBjWXaIXx2WaPFsHwgnZfuwWnXm6zetGo6Nt
Wuq9PWtDE4He3blY0dV+22pnyrXShxRsKX/o7XL+SGRZZQOqs8p/8RHsTDzY
qEHwzKBjh1dUSOg0JH+P0dWvr9pr9RAXyr2RdvM2aTMatyXaoy/9f+qY30JR
ipzO7fG3HgbkFR1ESjMpXseY/WeLUp+GP8Ni2VTXYY9VlkrrXMKtck5wvGWj
lx4KGOy9F3z8I0TtHkIKz0fkjlAaB16A5eilyNx8+LkiO9s2BTsO+fAixRLI
CKcU5r45HO0T8rSXZ29jKkGqxO7sr2UYoulZUPAAw1CZq5smn4DFFN61dJ2U
hCxXnFUhk1c6FkWHu+tPMnG4D7zyhdri76lpY3BRtcyRDaT4LxR1cCNRwGSL
lECcYwj89La8MWf/uEqhf2P+YAhYbu/RUZzB+DbX67BnXeC2JYBENElSXr9t
+/Apc1LyI+cXAhno4yV96orfzVEQkoDsNWFF91za3obm9ABBJKKJDFedIyHn
SRRCUt82DfszD3w7wJKMp6RlyrhiTh5RJPKzwhrw6hiyEIYxdecAWmFD3vtt
zD2HfbCETMrZMFYLvT1al4DGaOuv8YcSy5srvYdy7FJiemd9az9ZgWO2gZPY
zBp4EzJCySWtWjKah79qQfA+EcUBGVJF0YGa97Pb2wkSf34yCQy+zGXkTPI8
Mv5LW0DIP9/FQYeRVr33rK2QpJlaANulFLFBZUbWEv1LjL4s227FXRClfDNH
ECYURP5mWKMEgkRgxGtlpFO/JFDlb/RwZwHlGG0VALg6fS44GM75aIdvgqjJ
tfJv+xMfdPc2cSHQ/7BERb4QUVz5OsC2GtDMCrWXEB6EIrF2WwqA2IoNi1hJ
n1TfJt593LXAhI7TrHslDyhWbPXqKtaZpVd7dwHPGXif9udW9cfe0f3Mm3f4
uQxikIrFwgfTiXT27mI2tZ9lFDdOz+eGXTA+JkXTroI/v+FPfx4ZUhHzAS+G
tPltE9+9V3osL8C3lu15lFMwxEZTHdb9ERcYbN2lpwRMEXERtkzl++dGLcdY
XEzv8KIrMeYcXSAsvrVk3fpbYBPBakZTdeE/5kkq9zszO+X496+9sg2ROMLJ
Yp95ApdVTtwAKX65inRUTKvqBQddQTAuVAP+xZnLrKbmdL8ZtN0xdiH4RHD5
JrqMOdpe3fdWQ+qxFx9iidEwx3VmXXa30hQmiLmMoNZsTzbDasajOaq01BTC
BTFiQ6ifEkCMbXi0tAOFAbKAqtBafddUzLFIuJTAm5u75ZQ7nlopeNsgd4oW
nZY2o5/nNxp9/r10c1R0Xa7Yttygj3ZDR+RQ1ELZujS8Im3+RPB5XPN0j6Hv
7KC6mHC1GNG50YiF1B63UMY1oKEzkkBKR4roe6BWcLYpGoUUe0LDbP4mRXEd
s/nmyVC0v0mR39eu2xnqSMFt6VN7ypZGNz5/bn5kCi4BF2PpoSaMEwBzeVPk
BOjKXYWsO2M9439yeJtLMsYcbD9m4c7ISnMJ8HOq/kiQ6OzCyPIPcQqYnh0E
o1OjHwHp4Zk/RN+CxeYgd6qF3MwzdoVq1wCfpAyw0eUNEF7Tan1Hq5O3GIDB
FAVNhMzoJFWs3XAnRD8SH3uwCCbMof1BgJ/bnf1hQnQR2rx49d2kOYOOV4sl
VIAmMxCg9JA/LhnP50bG7YUmYPhY9HVXmI001Vx98efXmwcFIbhlXxgq1aoX
HAfFKk0pPqcRvinKxqQOpLE2y3CNe0HLTflpb2TG4WFWL6NCpcIRmkiRpGVd
dlf86yL+MrdQxAvexo2WNskcslEYarnn3uCrO0J7sNFT+QxSWtR7hjFulDfM
uICrNgT+2INrw1olfZH5LYo4J3lBtAqToF8UMDfdbl+cZ1CNiQuC2XnVvdQ0
MxMMugKJLixMcCnB6OhZbIzM4agyNLgUN9G78RkdRJmebkynPweOfZ/S00br
2dcceaxFTjM120pg2fSpxPAANhL31LQIZTzCssOBCEA8Wwhfb6Dd7C26B8f9
m8sZYFu8UNoxjUI6yx3oGm/UwrssnnvHbUNscSy2cNb2XsMHuvqW/YOFML/q
98jn5KJz3HX+FY1fyAsvxH4Wr5zUrIL87y/iJUE2SwIK/JFFijDhw2LhQM6/
yyNBP7xKxgLCTvsejbUXjgeP3KsFIowsKp8eQlvkVUS0B0VXBkFFqTahXxCi
i8R5LdMMsGEpCL4iw8iEbGGAJBx7EeVivLLDJues1DqKp4Xlyx6y974sYnof
2ZKYuJUI1QJs7PqwNjnjKGanEGsN5LxelzjjcRxHHopfIeNHoD/166HdOPtu
W0FlhegEATxKVYYbpbOiR5dI+2hJmZwbDFv92ry0Tt3ne6QRAsPAgyha5MxK
UAn/9UwGbh44pKFF+lhaSiMyQzLoeukuAGiYl8oCwYBiT35OQ7HFWZpJGItj
1WZx6FiUKAV+nEEKyedBe4Ef1oOSkZz5cjoIbg5+zjEk71oZgXUSSv57YT+U
NcIE4XBZnBZCqQTPxXmGxWmO0MNkXyIBxtuSNgPZZ8ObsDVBO9z5BOgG06wh
ns3OJ03vqndvTpkYiPYCISXlCitEOUPkPDy38SG1ivhgK2SoKPbzqO9WTJA4
3w99DPUib14fcKpatWMZZHMCASihqLajflO/b35pYmsr7jnGtuaFHWhEkOVv
K6uzTPhATTCjqIGu6Mvm+nHskhDPbaZJOKJykKQDdprZw7peuPdWpu2zldEY
Fr5TzQVoxl4hxi7bDt2bLlTpPHBC91I24Uh5t5qWsJYRGQkDBxuDZvwTUPML
/OTqkaYII8Iw2zeZSdYGcyAgc05eD6F1sk5M3UQtJkYFVUdzbqWlOe7VRc7I
ZgTNMXQBVc8LJx/kjbcM3D6HbYRHPqblb+UIF6ldrEJbNXPqhBnQT0Zz707l
RHft8WzpiyObasw4kZZndjsYvb6Jve1dkR6ZCmu7KOM3dngUDkVGhvZlgicN
e7K3SrKUKpNSbhyV/V/ZEJt/sjc7wqnnwvu2xe6KUa5TKiJ39UtN+UchNSFD
AVPxDASiezWhhX5l55Z91l/YkvfJH+L8QCrIovBcYbZJZTx1IQJboeanJPNd
KshWPgCUrnS/fe3/5VBesAiUk5kwi+ZdxuEKsO+pRZNOVyCU/I/9HbtfuW1L
aSKyqKLN94b9V5UUj0vbuFLiU9cZRv3fj6t4zwYpoISCGvQh7Gsz9W4uL/1Y
DiVi3P2BIZPRRiPgQvI8hluZhfP3uTZw98Cu5uqz6ZlXW+tIi9GsAVh2vISh
7WsYCzfBgoqrVx+jWBlql2GOkhRxAMdsDbvRIZjvslN+6/czxHDcgIZe8cZn
GEHOOFRF+6o8ynqIAdNgOllVErQxIHMd/GVYGNgBcqECk5RyHqpz1myhqNM1
EfXECK3BSLTwZduISYx/1/PHqaO0TuU6hu1hbXY0BOQSWKbaeGN5ob0V4DYs
M/x9mW6ejSDNIv13CLgTZupQsVKd0VqgmAqSmCpskr5S6pxah6za6HAlldlz
EAv6gCI6pNc8OE4lHAZJGZixxaB9HQdXDpYAj907PMpbDYLaWra3BtQVR0By
6/qjA4LCskY401gobTOhBRyzmgiuFLeiMV0NBEPRhjdyXQnDIKLOSPpQbG1N
F2397+xpisOavM9Z3l12/Olvu3kFevCWgDXjsVekNDnt9b8rjupuZWjXrMiz
ATjNa7MNFIT0f8Tur4JNp/mzd5yHyo547mc25QLLtprd1wRQ+YV+GNvsopJu
oXtJXGP4iupVPFUyVdD0KasCXgXlkcPUN1arMxXyY1caVNmCfNFaDsquueIJ
fBaiL8JavsfODUwX1Wz1XIdGxthUlgy69g2JIDreMZK43EuaxRpLCQU73tB7
3ZxIomiXGVKZPPCh7EJKkAyk5YB5u8AC83O84be5K0Dp+9lIopyI8Rl/EM9T
a9S6qXgV2jfruWL433A/1IFDUBIvxvhQkFmJcPeWy3Hpi+Jbs9t2tBP0OuUk
7IxI1LokMv97FKPBErL0YmzF6Rzold+zDFdjU1KAXRcIFqNPvKzCRy1hhhZX
sgSkWL0aPw/Rb3mpfvZfVKSEm3+CrzxjGbhofNwZxtDOeBjn6Ld8hBkGoSli
SuXOEYhrmb38RvbsCPe3fJDbPet0tvOPCZzNuHLkS4MRpRLppQDVCL8R5Ffu
KokNOdFhdxoBROUoCs3JYT4Q6L8zuSrsTxCu+GmR4GMFrq7OoJ4OpQHFHqPJ
hMqCmMRrDZOsDz1XDX5OXeUVHOyehl2xYQvjUfMfsK0KH76LsYS+xEr8g+3j
ge8hsNLX5fjp4Dkz0ITUGvGTVUEejH1OIxWXB0kNTKaU2Fj7b6AZPwZfRT7X
EpWQb6xyY+vtXI/lOkIDErHGtbbZpk3DTxsSQ8FseZAEjWWAzPNAkyDup+Vm
4Lm8pdiSv24lD/8VFuId7/Gp+W9C6KG/GSh64q8m12nrXlGoHZPYArY22u9q
nIk3inWZGvUDlI8CF4ox7qPx1+00vey0KsAlwcrYZZCJk0ObNMxxnFoPb/wj
UJoa9N11i6EqrQjb3Kkmz3zLte8hzrorCCiGtRfG9AO1EraFAZEeWF194PAv
f9F17YCFzOJPixxFOMK4YUB8eFXYPfS5MbfAx8YlR8ZKtmvWz4bZ30nEFIBX
H8GjNaObPqx1IlIIer8rNkYyo1dzT50KushLzyl9m7OZ5Xfcfl+0Mkq4IFxE
9R6m0TafCjpav8Vt0fr4SLee8syKHjgkosMNLuK11CltPX1SfJWcTVNPQYvw
cpYAm3yFQnm7wkoTobdSiOOb43lHuhe373/Hgwq5X+yIrmdFu/PDGa6Gs2WS
psmNka5i/Ppe1qhqCiJXNZK8jVhuPFWP0JV6Q/bXOgrsBlx3vebxEgpO1QK5
jSQpE3f4EXWc+gq/Jt9rYZ1onsPIKvjwoqwGLALpoe780DfOSa5sY9ejft70
a/pmL+KzMNAcxmceIaPRW+XwRn+v2poXA9cwoq/wF/RJTLpRYi+6LfODv9DB
3zceFjJEIZ5EBHWv9vsodrPmXg38h7TzBHiptTDoh/0UVzxSqCv+7d20kogF
tdxUnqGUidddO9aWq83qi01/eqRnAUvR/MEffDqyapz6Xg6kfOdQA0jl0d11
b69uL9sROLLsVZkjTzXj5g0pfQdz3UMTSqL60Z50Ei02olx0zoBoXuY4ay4u
Gr96yg6EFVp6EsG5PY2dTTlfW/ZQuHAWbEPoeH4c13o/tg6wy1+qFkPsXIpk
r7LsH3GP/06AOpp/rNthAwcXOC2PnVoolhqDD37c8YxKDwWIMoVtAUDWBBgL
argMoKa65lKyfVlYXc6ufGfH0iJRs6yM9aM9eamiUmqBR5m1VZ9Q6lDnSHRW
aMcxrnErv+ofCiJolSEuWnp/XMgVejq/lRzLvKDMW3Z3aJFXrdf/UrcenXEK
JlFrYlITD4W5CmJNtOdcUILBtYPOJf3NZaGiZiMgkmJeBine/wvwcwPtRRts
9wD2LjH3IMZmcEtluB5oLj7oxPxBcRrR0Qoh7Pmy/jdtp4O3mE0qk7z1GpCo
JvmQzBozk/jEp05kNsXz8PAH7UjE0zkdciK2C9iK5Oj7nGDc1Dck4ljEimRT
TvLrg7U/W22zbrRQ90FxPhIzZPJIxUPwns/JWtZ2NGnhlh8ZXsqUrYddYMR5
0too0JfIGdZk26HwSc3MudHBQFKQnSBCTC8LtFNMe4AKhHTVD6TiHpRklmkj
ajE+c5fFifJEkIF9U815GqnWLVP0WVaktU31Hdu5scbP66ZuCorkVJMVfBCi
CG/BTmIfcPgrkeRWHq8/umqd5uGsBa1ajrB/MCIpHZNW3GNrdP0DlJKqE5Kc
t2vWjnfe+LzC4LeQ2lxVVVn531N9jpm80kAQw2+MYa/zFocc07MrVwTzoeQI
Mo8YuTYYAA0MjLYteQ6AqHjqJSQXMqrA+DuGHShYaBgxxwoNTqSoWR294M0h
imG9rMZyVsL37pdxFMbNRQqwKiZdpoEp3XPmeDgnefLj7N71wcSjZv7vwZs9
DlAKYjrbAhEKEb1aXkXPXqpMRFHkFDBPPgOHgZyrOetZn33VZ5PO619sTXje
y/YyMNxZ6xzkQU5AL2G+gmwvk3ECIIM/xnztgfikYkXYj8j/J1caZ3OnhBs8
JDofyqLZT1RWe8cVcM9hISEuFMNq8JUOzz8Cko9LrrTeASEMeBw4QQ+XX/JZ
rawMCwaBA2AL3bHUySuOaYTvPuMUCSQoFAG7c00C111VMYpaWfeo1pFmra3f
c4YKxGjza+JTjgbaoT4+W8QaWkoBM4FzpERTdtccBFKU2jtH8Mj0sJ9S1i6W
rzG9vA1f+ZhyWFnnvgEI1yQbZyvPzhI1r8fpU3wmFPDfDbAY7I7vsImbG1v6
eXmigarPJxaXKUYifq6+VeCse7lPlsbsBfp2JvsgOx2A7Nn4oK9/NOiE+WuB
eGFMkLHc4KqhsM8w4EtA19gTr7Ku4RKru9scEYBlX3MAbm4HjhBTK7TPngvT
M2/3ZTJYt+H/H32pN2/eQnjQCcsKFJTgkmRMy+JBXyC/L9+sZgUOFha+9m0G
Yat0wesM/XbIzBtpyn3WB32ixwcAChtnRzYj1MpXkmQ1+aREB28GfGZiJ/qf
mXFmjdomjjHZGej5fl906HG1q0QB961+IFaAAn0tZvfoNzk5D/h+r4F6Gd3F
K02IgBn3UlUu1WrDuL18AGXpQWpdRochgjRnJ/w77EBarmNVq4UkGKD2nUH/
kbL6pTII6P2L7dKGO79wkVbGEt9lGQ59LKyoh3I38SnXPDwVfspWcXYdKNG9
eKxwnW1yFG1b1sfhDT1XQbD8

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "9RW93T28GeolckbYRvHffOsKFRFmORm+azyCUYhudrVC3P73ufaBfyRVMCXUVPfCA/gVx4qupGWo2/MTXHrbiqujt9kp6+gvryDIvlW8esKlSeDbKqIxzhLY+DL5yFAjg+mCmTKnMSoiZ9J0N0zgOO806IAkac+OYN9FbEIEFuaO+G41krhhxrcYAZ7qVX+m993ig0jH+TdTkf+bgk6VV++svRquWf4VNDUj099hz6ANJ4xL4kpKLH40ZB/PPAjpl9Lemxz4Rtfng6Ub67Vdg8+rqy3TbUa02cbrTJFKc45+VFELtiB6QYj7oNH458TiNRkITYR6Q3uzT6YhJ2tumIpF7Jc+aUilmD/s1y7neMyzEx/zdYYv6Cer00jKL+1CtvWQsBz4pDlAOds/IoePNd5wZ+cLHxeFJhbYyt67jVZ8tpbw9aDG5rNz0teALCTQF/P1YPDLnuN2kVorDa1LKBewgt6YRfnNgWUoo3D7AvjqoeRZMPEzuOQKnOoMm9gseBNEYgc7mtD1gC+C2haguz3Me1EufM+Czm7dXESt/JhCzowqHwRgWtIlwFAwNozOm07K2oufVqG5l+6Y5WHuqbs7pM0CkZADFOrkqu+dKqM8zkCpMdsm1Xv7pT794ToQ8wPtDEN6eHWZXiehiP2kzQJOz713RnBNowCY9WVJGFAXPuTA+3H/Ipqi+BPX57QgL111aZGUzDeOc2WM//d5lBcv7/XNolGJc6Z315AzLoMaeFAljF31H/Ozg2nnw4Ac6DijntOD1f5YyqyNaYTwJYkra80eKMBXDmbxWyCaQItYsf3NDi5eekqvd+87JBm2NDUliWxisovmRyUw3KIKc1J2EnfQNWzxZoK/QMbh+cxYd6vwfbzsLZtOGYJv2zmKbnC3HnSeKJ82dhzvgsQ/DHgRRZWcjbdmdGGxPH5l65GndJcOFEQmPfTAwNyA9vAMnglTlLm0NFHGqS9NwYV123o8SUAIN/Q6lCdzKhc796+vFQ13Po/Uhg2jKWtAzdT5"
`endif