// (C) 2001-2024 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


module intel_rtile_cxl_ast # (
//CXL sim time reduction
parameter qhip_rtile_pipe_mode = 0,
//CXL sim time reduction
parameter qhip_csb2wire_en_hwtcl                                                                                                                                                 = 0,
parameter qhip_mmio_enable_hwtcl                                                                                                                                                 = 0,
parameter opt_tx_big_buffer_hwtcl                                                                                                                                                = 0,
parameter opt_csb_pll_en_hwtcl                                                                                                                                                   = 0,
parameter opt_d2h_req23_en_hwtcl                                                                                                                                                 = 0,
parameter opt_cache_formatb_en_hwtcl                                                                                                                                             = 1,
parameter opt_chemem_flow_err_det_en_hwtcl                                                                                                                                       = 0,
parameter hssi_aibnd_rx_0_aib_ber_margining_ctrl                                                                                                                                 = "aib_ber_margining_setting0",
parameter hssi_aibnd_rx_0_aib_datasel_gr0                                                                                                                                        = "aib_datasel0_setting0",
parameter hssi_aibnd_rx_0_aib_datasel_gr1                                                                                                                                        = "aib_datasel1_setting1",
parameter hssi_aibnd_rx_0_aib_datasel_gr2                                                                                                                                        = "aib_datasel2_setting1",
parameter hssi_aibnd_rx_0_aib_dllstr_align_clkdiv                                                                                                                                = "aib_dllstr_align_clkdiv_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_dly_pst                                                                                                                               = "aib_dllstr_align_dly_pst_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_dy_ctl_static                                                                                                                         = "aib_dllstr_align_dy_ctl_static_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_dy_ctlsel                                                                                                                             = "aib_dllstr_align_dy_ctlsel_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_entest                                                                                                                                = "aib_dllstr_align_test_disable",
parameter hssi_aibnd_rx_0_aib_dllstr_align_halfcode                                                                                                                              = "aib_dllstr_align_halfcode_enable",
parameter hssi_aibnd_rx_0_aib_dllstr_align_selflock                                                                                                                              = "aib_dllstr_align_selflock_enable",
parameter hssi_aibnd_rx_0_aib_dllstr_align_st_core_dn_prgmnvrt                                                                                                                   = "aib_dllstr_align_st_core_dn_prgmnvrt_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_st_core_up_prgmnvrt                                                                                                                   = "aib_dllstr_align_st_core_up_prgmnvrt_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_st_core_updnen                                                                                                                        = "aib_dllstr_align_st_core_updnen_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_st_dftmuxsel                                                                                                                          = "aib_dllstr_align_st_dftmuxsel_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_st_en                                                                                                                                 = "aib_dllstr_align_st_en_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_st_hps_ctrl_en                                                                                                                        = "aib_dllstr_align_hps_ctrl_en_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_st_lockreq_muxsel                                                                                                                     = "aib_dllstr_align_st_lockreq_muxsel_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_st_new_dll                                                                                                                            = "aib_dllstr_align_new_dll_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_st_rst                                                                                                                                = "aib_dllstr_align_st_rst_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_st_rst_prgmnvrt                                                                                                                       = "aib_dllstr_align_st_rst_prgmnvrt_setting0",
parameter hssi_aibnd_rx_0_aib_dllstr_align_test_clk_pll_en_n                                                                                                                     = "aib_dllstr_align_test_clk_pll_en_n_disable",
parameter hssi_aibnd_rx_0_aib_inctrl_gr0                                                                                                                                         = "aib_inctrl0_setting0",
parameter hssi_aibnd_rx_0_aib_inctrl_gr1                                                                                                                                         = "aib_inctrl1_setting0",
parameter hssi_aibnd_rx_0_aib_inctrl_gr2                                                                                                                                         = "aib_inctrl2_setting0",
parameter hssi_aibnd_rx_0_aib_inctrl_gr3                                                                                                                                         = "aib_inctrl3_setting0",
parameter hssi_aibnd_rx_0_aib_outctrl_gr0                                                                                                                                        = "aib_outen0_setting0",
parameter hssi_aibnd_rx_0_aib_outctrl_gr1                                                                                                                                        = "aib_outen1_setting0",
parameter hssi_aibnd_rx_0_aib_outctrl_gr2                                                                                                                                        = "aib_outen2_setting0",
parameter hssi_aibnd_rx_0_aib_outndrv_r12                                                                                                                                        = "aib_ndrv12_setting1",
parameter hssi_aibnd_rx_0_aib_outndrv_r34                                                                                                                                        = "aib_ndrv34_setting1",
parameter hssi_aibnd_rx_0_aib_outndrv_r56                                                                                                                                        = "aib_ndrv56_setting1",
parameter hssi_aibnd_rx_0_aib_outndrv_r78                                                                                                                                        = "aib_ndrv78_setting1",
parameter hssi_aibnd_rx_0_aib_outpdrv_r12                                                                                                                                        = "aib_pdrv12_setting1",
parameter hssi_aibnd_rx_0_aib_outpdrv_r34                                                                                                                                        = "aib_pdrv34_setting1",
parameter hssi_aibnd_rx_0_aib_outpdrv_r56                                                                                                                                        = "aib_pdrv56_setting1",
parameter hssi_aibnd_rx_0_aib_outpdrv_r78                                                                                                                                        = "aib_pdrv78_setting1",
parameter hssi_aibnd_rx_0_aib_red_shift_en                                                                                                                                       = "aib_red_shift_disable",
parameter hssi_aibnd_rx_0_dft_hssitestip_dll_dcc_en                                                                                                                              = "disable_dft",
parameter hssi_aibnd_rx_0_op_mode                                                                                                                                                = "pwr_down",
parameter hssi_aibnd_rx_0_powerdown_mode                                                                                                                                         = "true",
parameter hssi_aibnd_rx_0_powermode_ac                                                                                                                                           = "rxdatapath_low_speed_pwr",
parameter hssi_aibnd_rx_0_powermode_dc                                                                                                                                           = "rxdatapath_powerdown",
parameter hssi_aibnd_rx_0_powermode_freq_hz_aib_hssi_rx_transfer_clk                                                                                                             = 0,
parameter hssi_aibnd_rx_0_redundancy_en                                                                                                                                          = "disable",
parameter hssi_aibnd_rx_0_sup_mode                                                                                                                                               = "user_mode",
parameter hssi_ctr_silicon_rev                                                                                                                                                   = "10nm6arnra",
parameter hssi_aibnd_tx_0_aib_datasel_gr0                                                                                                                                        = "aib_datasel0_setting0",
parameter hssi_aibnd_tx_0_aib_datasel_gr1                                                                                                                                        = "aib_datasel1_setting0",
parameter hssi_aibnd_tx_0_aib_datasel_gr2                                                                                                                                        = "aib_datasel2_setting1",
parameter hssi_aibnd_tx_0_aib_datasel_gr3                                                                                                                                        = "aib_datasel3_setting1",
parameter hssi_aibnd_tx_0_aib_ddrctrl_gr0                                                                                                                                        = "aib_ddr0_setting1",
parameter hssi_aibnd_tx_0_aib_hssi_tx_transfer_clk_hz                                                                                                                            = 0,
parameter hssi_aibnd_tx_0_aib_iinasyncen                                                                                                                                         = "aib_inasyncen_setting0",
parameter hssi_aibnd_tx_0_aib_iinclken                                                                                                                                           = "aib_inclken_setting0",
parameter hssi_aibnd_tx_0_aib_outctrl_gr0                                                                                                                                        = "aib_outen0_setting0",
parameter hssi_aibnd_tx_0_aib_outctrl_gr1                                                                                                                                        = "aib_outen1_setting0",
parameter hssi_aibnd_tx_0_aib_outctrl_gr2                                                                                                                                        = "aib_outen2_setting0",
parameter hssi_aibnd_tx_0_aib_outctrl_gr3                                                                                                                                        = "aib_outen3_setting0",
parameter hssi_aibnd_tx_0_aib_outndrv_r34                                                                                                                                        = "aib_ndrv34_setting1",
parameter hssi_aibnd_tx_0_aib_outndrv_r56                                                                                                                                        = "aib_ndrv56_setting1",
parameter hssi_aibnd_tx_0_aib_outpdrv_r34                                                                                                                                        = "aib_pdrv34_setting1",
parameter hssi_aibnd_tx_0_aib_outpdrv_r56                                                                                                                                        = "aib_pdrv56_setting1",
parameter hssi_aibnd_tx_0_aib_red_dirclkn_shiften                                                                                                                                = "aib_red_dirclkn_shift_disable",
parameter hssi_aibnd_tx_0_aib_red_dirclkp_shiften                                                                                                                                = "aib_red_dirclkp_shift_disable",
parameter hssi_aibnd_tx_0_aib_red_drx_shiften                                                                                                                                    = "aib_red_drx_shift_disable",
parameter hssi_aibnd_tx_0_aib_red_dtx_shiften                                                                                                                                    = "aib_red_dtx_shift_disable",
parameter hssi_aibnd_tx_0_aib_red_pout_shiften                                                                                                                                   = "aib_red_pout_shift_disable",
parameter hssi_aibnd_tx_0_aib_red_rx_shiften                                                                                                                                     = "aib_red_rx_shift_disable",
parameter hssi_aibnd_tx_0_aib_red_tx_shiften                                                                                                                                     = "aib_red_tx_shift_disable",
parameter hssi_aibnd_tx_0_aib_red_txferclkout_shiften                                                                                                                            = "aib_red_txferclkout_shift_disable",
parameter hssi_aibnd_tx_0_aib_red_txferclkoutn_shiften                                                                                                                           = "aib_red_txferclkoutn_shift_disable",
parameter hssi_aibnd_tx_0_aib_tx_clkdiv                                                                                                                                          = "aib_tx_clkdiv_setting1",
parameter hssi_aibnd_tx_0_aib_tx_dcc_byp                                                                                                                                         = "aib_tx_dcc_byp_disable",
parameter hssi_aibnd_tx_0_aib_tx_dcc_byp_iocsr_unused                                                                                                                            = "aib_tx_dcc_byp_disable_iocsr_unused",
parameter hssi_aibnd_tx_0_aib_tx_dcc_cont_cal                                                                                                                                    = "aib_tx_dcc_cal_cont",
parameter hssi_aibnd_tx_0_aib_tx_dcc_cont_cal_iocsr_unused                                                                                                                       = "aib_tx_dcc_cal_single_iocsr_unused",
parameter hssi_aibnd_tx_0_aib_tx_dcc_dft                                                                                                                                         = "aib_tx_dcc_dft_disable",
parameter hssi_aibnd_tx_0_aib_tx_dcc_dft_sel                                                                                                                                     = "aib_tx_dcc_dft_mode0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_dll_dft_sel                                                                                                                                 = "aib_tx_dcc_dll_dft_sel_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_dll_entest                                                                                                                                  = "aib_tx_dcc_dll_test_disable",
parameter hssi_aibnd_tx_0_aib_tx_dcc_dy_ctl_static                                                                                                                               = "aib_tx_dcc_dy_ctl_static_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_dy_ctlsel                                                                                                                                   = "aib_tx_dcc_dy_ctlsel_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_en                                                                                                                                          = "aib_tx_dcc_enable",
parameter hssi_aibnd_tx_0_aib_tx_dcc_en_iocsr_unused                                                                                                                             = "aib_tx_dcc_disable_iocsr_unused",
parameter hssi_aibnd_tx_0_aib_tx_dcc_manual_dn                                                                                                                                   = "aib_tx_dcc_manual_dn0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_manual_up                                                                                                                                   = "aib_tx_dcc_manual_up0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_rst_prgmnvrt                                                                                                                                = "aib_tx_dcc_st_rst_prgmnvrt_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_st_core_dn_prgmnvrt                                                                                                                         = "aib_tx_dcc_st_core_dn_prgmnvrt_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_st_core_up_prgmnvrt                                                                                                                         = "aib_tx_dcc_st_core_up_prgmnvrt_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_st_core_updnen                                                                                                                              = "aib_tx_dcc_st_core_updnen_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_st_dftmuxsel                                                                                                                                = "aib_tx_dcc_st_dftmuxsel_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_st_dly_pst                                                                                                                                  = "aib_tx_dcc_st_dly_pst_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_st_en                                                                                                                                       = "aib_tx_dcc_st_en_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_st_hps_ctrl_en                                                                                                                              = "aib_tx_dcc_hps_ctrl_en_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_st_lockreq_muxsel                                                                                                                           = "aib_tx_dcc_st_lockreq_muxsel_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_st_new_dll                                                                                                                                  = "aib_tx_dcc_new_dll_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_st_rst                                                                                                                                      = "aib_tx_dcc_st_rst_setting0",
parameter hssi_aibnd_tx_0_aib_tx_dcc_test_clk_pll_en_n                                                                                                                           = "aib_tx_dcc_test_clk_pll_en_n_disable",
parameter hssi_aibnd_tx_0_aib_tx_halfcode                                                                                                                                        = "aib_tx_halfcode_enable",
parameter hssi_aibnd_tx_0_aib_tx_selflock                                                                                                                                        = "aib_tx_selflock_enable",
parameter hssi_aibnd_tx_0_dfd_dll_dcc_en                                                                                                                                         = "disable_dfd",
parameter hssi_aibnd_tx_0_dft_hssitestip_dll_dcc_en                                                                                                                              = "disable_dft",
parameter hssi_aibnd_tx_0_op_mode                                                                                                                                                = "tx_dcc_enable",
parameter hssi_aibnd_tx_0_powerdown_mode                                                                                                                                         = "true",
parameter hssi_aibnd_tx_0_powermode_ac                                                                                                                                           = "txdatapath_low_speed_pwr",
parameter hssi_aibnd_tx_0_powermode_dc                                                                                                                                           = "txdatapath_powerdown",
parameter hssi_aibnd_tx_0_powermode_freq_hz_aib_hssi_tx_transfer_clk                                                                                                             = 0,
parameter hssi_aibnd_tx_0_redundancy_en                                                                                                                                          = "disable",
parameter hssi_aibnd_tx_0_sup_mode                                                                                                                                               = "user_mode",
parameter hssi_pldadapt_tx_0_aib_clk1_sel                                                                                                                                        = "aib_clk1_pld_pcs_tx_clk_out",
parameter hssi_pldadapt_tx_0_aib_clk2_sel                                                                                                                                        = "aib_clk2_pld_pcs_tx_clk_out",
parameter hssi_pldadapt_tx_0_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                                                               = 0,
parameter hssi_pldadapt_tx_0_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz                                                                                                             = 0,
parameter hssi_pldadapt_tx_0_hdpldadapt_aib_fabric_tx_sr_clk_in_hz                                                                                                               = 0,
parameter hssi_pldadapt_tx_0_bonding_dft_en                                                                                                                                      = "dft_dis",
parameter hssi_pldadapt_tx_0_bonding_dft_val                                                                                                                                     = "dft_0",
parameter hssi_pldadapt_tx_0_chnl_bonding                                                                                                                                        = "disable",
parameter hssi_pldadapt_tx_0_comp_cnt                                                                                                                                            = 0,
parameter hssi_pldadapt_tx_0_compin_sel                                                                                                                                          = "compin_master",
parameter hssi_pldadapt_tx_0_hdpldadapt_csr_clk_hz                                                                                                                               = 0,
parameter hssi_pldadapt_tx_0_ctrl_plane_bonding                                                                                                                                  = "individual",
parameter hssi_pldadapt_tx_0_ds_bypass_pipeln                                                                                                                                    = "ds_bypass_pipeln_dis",
parameter hssi_pldadapt_tx_0_ds_last_chnl                                                                                                                                        = "ds_not_last_chnl",
parameter hssi_pldadapt_tx_0_ds_master                                                                                                                                           = "ds_master_en",
parameter hssi_pldadapt_tx_0_duplex_mode                                                                                                                                         = "disable",
parameter hssi_pldadapt_tx_0_dv_bond                                                                                                                                             = "dv_bond_dis",
parameter hssi_pldadapt_tx_0_dv_gen                                                                                                                                              = "dv_gen_dis",
parameter hssi_pldadapt_tx_0_fifo_double_write                                                                                                                                   = "fifo_double_write_dis",
parameter hssi_pldadapt_tx_0_fifo_mode                                                                                                                                           = "phase_comp",
parameter hssi_pldadapt_tx_0_fifo_rd_clk_frm_gen_scg_en                                                                                                                          = "disable",
parameter hssi_pldadapt_tx_0_fifo_rd_clk_scg_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_tx_0_fifo_rd_clk_sel                                                                                                                                     = "fifo_rd_pma_aib_tx_clk",
parameter hssi_pldadapt_tx_0_fifo_stop_rd                                                                                                                                        = "n_rd_empty",
parameter hssi_pldadapt_tx_0_fifo_stop_wr                                                                                                                                        = "n_wr_full",
parameter hssi_pldadapt_tx_0_fifo_width                                                                                                                                          = "fifo_single_width",
parameter hssi_pldadapt_tx_0_fifo_wr_clk_scg_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_tx_0_fpll_shared_direct_async_in_sel                                                                                                                     = "fpll_shared_direct_async_in_rowclk",
parameter hssi_pldadapt_tx_0_frmgen_burst                                                                                                                                        = "frmgen_burst_dis",
parameter hssi_pldadapt_tx_0_frmgen_bypass                                                                                                                                       = "frmgen_bypass_dis",
parameter hssi_pldadapt_tx_0_frmgen_mfrm_length                                                                                                                                  = 2048,
parameter hssi_pldadapt_tx_0_frmgen_pipeln                                                                                                                                       = "frmgen_pipeln_dis",
parameter hssi_pldadapt_tx_0_frmgen_pyld_ins                                                                                                                                     = "frmgen_pyld_ins_dis",
parameter hssi_pldadapt_tx_0_frmgen_wordslip                                                                                                                                     = "frmgen_wordslip_dis",
parameter hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit0_rst_val                                                                                                                         = "reset_to_zero_hfsrin0",
parameter hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit1_rst_val                                                                                                                         = "reset_to_zero_hfsrin1",
parameter hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit2_rst_val                                                                                                                         = "reset_to_zero_hfsrin2",
parameter hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit3_rst_val                                                                                                                         = "reset_to_zero_hfsrin3",
parameter hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit0_rst_val                                                                                                                        = "reset_to_zero_hfsrout0",
parameter hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit1_rst_val                                                                                                                        = "reset_to_zero_hfsrout1",
parameter hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit2_rst_val                                                                                                                        = "reset_to_zero_hfsrout2",
parameter hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit3_rst_val                                                                                                                        = "reset_to_zero_hfsrout3",
parameter hssi_pldadapt_tx_0_fsr_mask_tx_pll_rst_val                                                                                                                             = "reset_to_zero_maskpll",
parameter hssi_pldadapt_tx_0_fsr_pld_txelecidle_rst_val                                                                                                                          = "reset_to_zero_txelec",
parameter hssi_pldadapt_tx_0_gb_tx_idwidth                                                                                                                                       = "idwidth_66",
parameter hssi_pldadapt_tx_0_gb_tx_odwidth                                                                                                                                       = "odwidth_32",
parameter hssi_pldadapt_tx_0_hip_mode                                                                                                                                            = "disable_hip",
parameter hssi_pldadapt_tx_0_hip_osc_clk_scg_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_tx_0_hrdrst_dcd_cal_done_bypass                                                                                                                          = "disable",
parameter hssi_pldadapt_tx_0_hrdrst_rst_sm_dis                                                                                                                                   = "enable_tx_rst_sm",
parameter hssi_pldadapt_tx_0_hrdrst_rx_osc_clk_scg_en                                                                                                                            = "disable",
parameter hssi_pldadapt_tx_0_hrdrst_user_ctl_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_tx_0_indv                                                                                                                                                = "indv_en",
parameter hssi_pldadapt_tx_0_is_paired_with                                                                                                                                      = "other",
parameter hssi_pldadapt_tx_0_loopback_mode                                                                                                                                       = "disable",
parameter hssi_pldadapt_tx_0_low_latency_en                                                                                                                                      = "disable",
parameter hssi_pldadapt_tx_0_osc_clk_scg_en                                                                                                                                      = "disable",
parameter hssi_pldadapt_tx_0_phcomp_rd_del                                                                                                                                       = "phcomp_rd_del2",
parameter hssi_pldadapt_tx_0_pipe_mode                                                                                                                                           = "disable_pipe",
parameter hssi_pldadapt_tx_0_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                                                                  = 0,
parameter hssi_pldadapt_tx_0_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                                                                  = 0,
parameter hssi_pldadapt_tx_0_pld_clk1_delay_en                                                                                                                                   = "disable",
parameter hssi_pldadapt_tx_0_pld_clk1_delay_sel                                                                                                                                  = "delay_path0",
parameter hssi_pldadapt_tx_0_pld_clk1_inv_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_tx_0_pld_clk1_sel                                                                                                                                        = "pld_clk1_rowclk",
parameter hssi_pldadapt_tx_0_pld_clk2_sel                                                                                                                                        = "pld_clk2_rowclk",
parameter hssi_pldadapt_tx_0_hdpldadapt_pld_sclk1_rowclk_hz                                                                                                                      = 0,
parameter hssi_pldadapt_tx_0_hdpldadapt_pld_sclk2_rowclk_hz                                                                                                                      = 0,
parameter hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk1_dcm_hz                                                                                                                       = 0,
parameter hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk1_rowclk_hz                                                                                                                    = 0,
parameter hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk2_dcm_hz                                                                                                                       = 0,
parameter hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk2_rowclk_hz                                                                                                                    = 0,
parameter hssi_pldadapt_tx_0_pma_aib_tx_clk_expected_setting                                                                                                                     = "not_used",
parameter hssi_pldadapt_tx_0_powerdown_mode                                                                                                                                      = "powerdown",
parameter hssi_pldadapt_tx_0_powermode_dc                                                                                                                                        = "powerdown",
parameter hssi_pldadapt_tx_0_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                                                           = 0,
parameter hssi_pldadapt_tx_0_powermode_freq_hz_pld_tx_clk1_dcm                                                                                                                   = 0,
parameter hssi_pldadapt_tx_0_sh_err                                                                                                                                              = "sh_err_dis",
parameter hssi_pldadapt_tx_0_hdpldadapt_speed_grade                                                                                                                              = "dash_1",
parameter hssi_pldadapt_tx_0_hdpldadapt_sr_sr_testbus_sel                                                                                                                        = "ssr_testbus",
parameter hssi_pldadapt_tx_0_stretch_num_stages                                                                                                                                  = "zero_stage",
parameter hssi_pldadapt_tx_0_sup_mode                                                                                                                                            = "user_mode",
parameter hssi_pldadapt_tx_0_tx_datapath_tb_sel                                                                                                                                  = "cp_bond",
parameter hssi_pldadapt_tx_0_tx_fastbond_rden                                                                                                                                    = "rden_ds_del_us_del",
parameter hssi_pldadapt_tx_0_tx_fastbond_wren                                                                                                                                    = "wren_ds_del_us_del",
parameter hssi_pldadapt_tx_0_tx_fifo_power_mode                                                                                                                                  = "full_width_full_depth",
parameter hssi_pldadapt_tx_0_tx_fifo_read_latency_adjust                                                                                                                         = "disable",
parameter hssi_pldadapt_tx_0_tx_fifo_write_latency_adjust                                                                                                                        = "disable",
parameter hssi_pldadapt_tx_0_tx_hip_aib_ssr_in_polling_bypass                                                                                                                    = "disable",
parameter hssi_pldadapt_tx_0_tx_osc_clock_setting                                                                                                                                = "osc_clk_div_by1",
parameter hssi_pldadapt_tx_0_tx_pld_10g_tx_bitslip_polling_bypass                                                                                                                = "disable",
parameter hssi_pldadapt_tx_0_tx_pld_8g_tx_boundary_sel_polling_bypass                                                                                                            = "disable",
parameter hssi_pldadapt_tx_0_tx_pld_pma_fpll_cnt_sel_polling_bypass                                                                                                              = "disable",
parameter hssi_pldadapt_tx_0_tx_pld_pma_fpll_num_phase_shifts_polling_bypass                                                                                                     = "disable",
parameter hssi_pldadapt_tx_0_tx_usertest_sel                                                                                                                                     = "enable",
parameter hssi_pldadapt_tx_0_txfifo_empty                                                                                                                                        = "empty_default",
parameter hssi_pldadapt_tx_0_txfifo_full                                                                                                                                         = "full_pc_sw",
parameter hssi_pldadapt_tx_0_txfifo_mode                                                                                                                                         = "txphase_comp",
parameter hssi_pldadapt_tx_0_txfifo_pempty                                                                                                                                       = 2,
parameter hssi_pldadapt_tx_0_txfifo_pfull                                                                                                                                        = 24,
parameter hssi_pldadapt_tx_0_us_bypass_pipeln                                                                                                                                    = "us_bypass_pipeln_dis",
parameter hssi_pldadapt_tx_0_us_last_chnl                                                                                                                                        = "us_not_last_chnl",
parameter hssi_pldadapt_tx_0_us_master                                                                                                                                           = "us_master_en",
parameter hssi_pldadapt_tx_0_word_align_enable                                                                                                                                   = "disable",
parameter hssi_pldadapt_tx_0_word_mark                                                                                                                                           = "wm_en",
parameter hssi_pldadapt_tx_0_reconfig_settings                                                                                                                                   = "{}",
parameter hssi_pldadapt_rx_0_aib_clk1_sel                                                                                                                                        = "aib_clk1_rx_transfer_clk",
parameter hssi_pldadapt_rx_0_aib_clk2_sel                                                                                                                                        = "aib_clk2_rx_transfer_clk",
parameter hssi_pldadapt_rx_0_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                                                               = 0,
parameter hssi_pldadapt_rx_0_hdpldadapt_aib_fabric_rx_sr_clk_in_hz                                                                                                               = 0,
parameter hssi_pldadapt_rx_0_hdpldadapt_aib_fabric_rx_transfer_clk_hz                                                                                                            = 0,
parameter hssi_pldadapt_rx_0_asn_bypass_pma_pcie_sw_done                                                                                                                         = "disable",
parameter hssi_pldadapt_rx_0_asn_en                                                                                                                                              = "disable",
parameter hssi_pldadapt_rx_0_asn_wait_for_dll_reset_cnt                                                                                                                          = 0,
parameter hssi_pldadapt_rx_0_asn_wait_for_fifo_flush_cnt                                                                                                                         = 0,
parameter hssi_pldadapt_rx_0_asn_wait_for_pma_pcie_sw_done_cnt                                                                                                                   = 0,
parameter hssi_pldadapt_rx_0_bonding_dft_en                                                                                                                                      = "dft_dis",
parameter hssi_pldadapt_rx_0_bonding_dft_val                                                                                                                                     = "dft_0",
parameter hssi_pldadapt_rx_0_chnl_bonding                                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_0_clock_del_measure_enable                                                                                                                            = "disable",
parameter hssi_pldadapt_rx_0_comp_cnt                                                                                                                                            = 0,
parameter hssi_pldadapt_rx_0_compin_sel                                                                                                                                          = "compin_master",
parameter hssi_pldadapt_rx_0_hdpldadapt_csr_clk_hz                                                                                                                               = 0,
parameter hssi_pldadapt_rx_0_ctrl_plane_bonding                                                                                                                                  = "individual",
parameter hssi_pldadapt_rx_0_ds_bypass_pipeln                                                                                                                                    = "ds_bypass_pipeln_dis",
parameter hssi_pldadapt_rx_0_ds_last_chnl                                                                                                                                        = "ds_not_last_chnl",
parameter hssi_pldadapt_rx_0_ds_master                                                                                                                                           = "ds_master_en",
parameter hssi_pldadapt_rx_0_duplex_mode                                                                                                                                         = "disable",
parameter hssi_pldadapt_rx_0_dv_mode                                                                                                                                             = "dv_mode_dis",
parameter hssi_pldadapt_rx_0_fifo_double_read                                                                                                                                    = "fifo_double_read_dis",
parameter hssi_pldadapt_rx_0_fifo_mode                                                                                                                                           = "phase_comp",
parameter hssi_pldadapt_rx_0_fifo_rd_clk_ins_sm_scg_en                                                                                                                           = "disable",
parameter hssi_pldadapt_rx_0_fifo_rd_clk_scg_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_rx_0_fifo_rd_clk_sel                                                                                                                                     = "fifo_rd_clk_rx_transfer_clk",
parameter hssi_pldadapt_rx_0_fifo_stop_rd                                                                                                                                        = "n_rd_empty",
parameter hssi_pldadapt_rx_0_fifo_stop_wr                                                                                                                                        = "n_wr_full",
parameter hssi_pldadapt_rx_0_fifo_width                                                                                                                                          = "fifo_single_width",
parameter hssi_pldadapt_rx_0_fifo_wr_clk_del_sm_scg_en                                                                                                                           = "disable",
parameter hssi_pldadapt_rx_0_fifo_wr_clk_scg_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_rx_0_fifo_wr_clk_sel                                                                                                                                     = "fifo_wr_clk_rx_transfer_clk",
parameter hssi_pldadapt_rx_0_free_run_div_clk                                                                                                                                    = "out_of_reset_sync",
parameter hssi_pldadapt_rx_0_fsr_pld_10g_rx_crc32_err_rst_val                                                                                                                    = "reset_to_zero_crc32",
parameter hssi_pldadapt_rx_0_fsr_pld_8g_sigdet_out_rst_val                                                                                                                       = "reset_to_zero_sigdet",
parameter hssi_pldadapt_rx_0_fsr_pld_ltd_b_rst_val                                                                                                                               = "reset_to_zero_ltdb",
parameter hssi_pldadapt_rx_0_fsr_pld_ltr_rst_val                                                                                                                                 = "reset_to_zero_ltr",
parameter hssi_pldadapt_rx_0_fsr_pld_rx_fifo_align_clr_rst_val                                                                                                                   = "reset_to_zero_alignclr",
parameter hssi_pldadapt_rx_0_gb_rx_idwidth                                                                                                                                       = "idwidth_32",
parameter hssi_pldadapt_rx_0_gb_rx_odwidth                                                                                                                                       = "odwidth_66",
parameter hssi_pldadapt_rx_0_hip_mode                                                                                                                                            = "disable_hip",
parameter hssi_pldadapt_rx_0_hrdrst_align_bypass                                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_0_hrdrst_dll_lock_bypass                                                                                                                              = "disable",
parameter hssi_pldadapt_rx_0_hrdrst_rst_sm_dis                                                                                                                                   = "enable_rx_rst_sm",
parameter hssi_pldadapt_rx_0_hrdrst_rx_osc_clk_scg_en                                                                                                                            = "disable",
parameter hssi_pldadapt_rx_0_hrdrst_user_ctl_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_rx_0_indv                                                                                                                                                = "indv_en",
parameter hssi_pldadapt_rx_0_internal_clk1_sel1                                                                                                                                  = "pma_clks_or_txfiford_post_ct_mux_clk1_mux1",
parameter hssi_pldadapt_rx_0_internal_clk1_sel2                                                                                                                                  = "pma_clks_clk1_mux2",
parameter hssi_pldadapt_rx_0_internal_clk2_sel1                                                                                                                                  = "pma_clks_or_rxfifowr_post_ct_mux_clk2_mux1",
parameter hssi_pldadapt_rx_0_internal_clk2_sel2                                                                                                                                  = "pma_clks_clk2_mux2",
parameter hssi_pldadapt_rx_0_is_paired_with                                                                                                                                      = "other",
parameter hssi_pldadapt_rx_0_loopback_mode                                                                                                                                       = "disable",
parameter hssi_pldadapt_rx_0_low_latency_en                                                                                                                                      = "disable",
parameter hssi_pldadapt_rx_0_lpbk_mode                                                                                                                                           = "disable",
parameter hssi_pldadapt_rx_0_osc_clk_scg_en                                                                                                                                      = "disable",
parameter hssi_pldadapt_rx_0_phcomp_rd_del                                                                                                                                       = "phcomp_rd_del2",
parameter hssi_pldadapt_rx_0_pipe_enable                                                                                                                                         = "disable",
parameter hssi_pldadapt_rx_0_pipe_mode                                                                                                                                           = "disable_pipe",
parameter hssi_pldadapt_rx_0_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                                                                  = 0,
parameter hssi_pldadapt_rx_0_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                                                                  = 0,
parameter hssi_pldadapt_rx_0_pld_clk1_delay_en                                                                                                                                   = "disable",
parameter hssi_pldadapt_rx_0_pld_clk1_delay_sel                                                                                                                                  = "delay_path0",
parameter hssi_pldadapt_rx_0_pld_clk1_inv_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_rx_0_pld_clk1_sel                                                                                                                                        = "pld_clk1_rowclk",
parameter hssi_pldadapt_rx_0_hdpldadapt_pld_rx_clk1_dcm_hz                                                                                                                       = 0,
parameter hssi_pldadapt_rx_0_hdpldadapt_pld_rx_clk1_rowclk_hz                                                                                                                    = 0,
parameter hssi_pldadapt_rx_0_hdpldadapt_pld_sclk1_rowclk_hz                                                                                                                      = 0,
parameter hssi_pldadapt_rx_0_hdpldadapt_pld_sclk2_rowclk_hz                                                                                                                      = 0,
parameter hssi_pldadapt_rx_0_pma_hclk_scg_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_rx_0_powerdown_mode                                                                                                                                      = "powerdown",
parameter hssi_pldadapt_rx_0_powermode_dc                                                                                                                                        = "powerdown",
parameter hssi_pldadapt_rx_0_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                                                           = 0,
parameter hssi_pldadapt_rx_0_powermode_freq_hz_pld_rx_clk1_dcm                                                                                                                   = 0,
parameter hssi_pldadapt_rx_0_rx_datapath_tb_sel                                                                                                                                  = "cp_bond",
parameter hssi_pldadapt_rx_0_rx_fastbond_rden                                                                                                                                    = "rden_ds_del_us_del",
parameter hssi_pldadapt_rx_0_rx_fastbond_wren                                                                                                                                    = "wren_ds_del_us_del",
parameter hssi_pldadapt_rx_0_rx_fifo_power_mode                                                                                                                                  = "full_width_full_depth",
parameter hssi_pldadapt_rx_0_rx_fifo_read_latency_adjust                                                                                                                         = "disable",
parameter hssi_pldadapt_rx_0_rx_fifo_write_ctrl                                                                                                                                  = "blklock_stops",
parameter hssi_pldadapt_rx_0_rx_fifo_write_latency_adjust                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_0_rx_osc_clock_setting                                                                                                                                = "osc_clk_div_by1",
parameter hssi_pldadapt_rx_0_rx_pld_8g_eidleinfersel_polling_bypass                                                                                                              = "disable",
parameter hssi_pldadapt_rx_0_rx_pld_pma_eye_monitor_polling_bypass                                                                                                               = "disable",
parameter hssi_pldadapt_rx_0_rx_pld_pma_pcie_switch_polling_bypass                                                                                                               = "disable",
parameter hssi_pldadapt_rx_0_rx_pld_pma_reser_out_polling_bypass                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_0_rx_prbs_flags_sr_enable                                                                                                                             = "disable",
parameter hssi_pldadapt_rx_0_rx_true_b2b                                                                                                                                         = "b2b",
parameter hssi_pldadapt_rx_0_rx_usertest_sel                                                                                                                                     = "enable",
parameter hssi_pldadapt_rx_0_rxfifo_empty                                                                                                                                        = "empty_sw",
parameter hssi_pldadapt_rx_0_rxfifo_full                                                                                                                                         = "full_pc_sw",
parameter hssi_pldadapt_rx_0_rxfifo_mode                                                                                                                                         = "rxphase_comp",
parameter hssi_pldadapt_rx_0_rxfifo_pempty                                                                                                                                       = 2,
parameter hssi_pldadapt_rx_0_rxfifo_pfull                                                                                                                                        = 48,
parameter hssi_pldadapt_rx_0_rxfiford_post_ct_sel                                                                                                                                = "rxfiford_sclk_post_ct",
parameter hssi_pldadapt_rx_0_rxfifowr_post_ct_sel                                                                                                                                = "rxfifowr_sclk_post_ct",
parameter hssi_pldadapt_rx_0_sclk_sel                                                                                                                                            = "sclk1_rowclk",
parameter hssi_pldadapt_rx_0_hdpldadapt_speed_grade                                                                                                                              = "dash_1",
parameter hssi_pldadapt_rx_0_hdpldadapt_sr_sr_testbus_sel                                                                                                                        = "ssr_testbus",
parameter hssi_pldadapt_rx_0_stretch_num_stages                                                                                                                                  = "zero_stage",
parameter hssi_pldadapt_rx_0_sup_mode                                                                                                                                            = "user_mode",
parameter hssi_pldadapt_rx_0_txfiford_post_ct_sel                                                                                                                                = "txfiford_sclk_post_ct",
parameter hssi_pldadapt_rx_0_txfifowr_post_ct_sel                                                                                                                                = "txfifowr_sclk_post_ct",
parameter hssi_pldadapt_rx_0_us_bypass_pipeln                                                                                                                                    = "us_bypass_pipeln_dis",
parameter hssi_pldadapt_rx_0_us_last_chnl                                                                                                                                        = "us_not_last_chnl",
parameter hssi_pldadapt_rx_0_us_master                                                                                                                                           = "us_master_en",
parameter hssi_pldadapt_rx_0_word_align                                                                                                                                          = "wa_en",
parameter hssi_pldadapt_rx_0_word_align_enable                                                                                                                                   = "disable",
parameter hssi_pldadapt_rx_0_reconfig_settings                                                                                                                                   = "{}",
parameter hssi_avmm1_if_0_pcs_arbiter_ctrl                                                                                                                                       = "avmm1_arbiter_uc_sel",
parameter hssi_avmm1_if_0_hssiadapt_avmm_clk_dcg_en                                                                                                                              = "disable",
parameter hssi_avmm1_if_0_hssiadapt_avmm_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm1_if_0_pldadapt_avmm_clk_scg_en                                                                                                                               = "disable",
parameter hssi_avmm1_if_0_pcs_cal_done                                                                                                                                           = "avmm1_cal_done_assert",
parameter hssi_avmm1_if_0_pcs_cal_reserved                                                                                                                                       = 0,
parameter hssi_avmm1_if_0_pcs_calibration_feature_en                                                                                                                             = "avmm1_pcs_calibration_dis",
parameter hssi_avmm1_if_0_pldadapt_gate_dis                                                                                                                                      = "disable",
parameter hssi_avmm1_if_0_pcs_hip_cal_en                                                                                                                                         = "disable",
parameter hssi_avmm1_if_0_hssiadapt_nfhssi_calibratio_feature_en                                                                                                                 = "disable",
parameter hssi_avmm1_if_0_pldadapt_nfhssi_calibratio_feature_en                                                                                                                  = "disable",
parameter hssi_avmm1_if_0_hssiadapt_osc_clk_scg_en                                                                                                                               = "disable",
parameter hssi_avmm1_if_0_pldadapt_osc_clk_scg_en                                                                                                                                = "disable",
parameter hssi_avmm1_if_0_hssiadapt_read_blocking_enable                                                                                                                         = "enable",
parameter hssi_avmm1_if_0_pldadapt_read_blocking_enable                                                                                                                          = "enable",
parameter hssi_avmm1_if_0_hssiadapt_uc_blocking_enable                                                                                                                           = "enable",
parameter hssi_avmm1_if_0_pldadapt_uc_blocking_enable                                                                                                                            = "enable",
parameter hssi_avmm1_if_0_hssiadapt_write_resp_en                                                                                                                                = "disable",
parameter hssi_avmm1_if_0_hssiadapt_avmm_osc_clock_setting                                                                                                                       = "osc_clk_div_by1",
parameter hssi_avmm1_if_0_pldadapt_avmm_osc_clock_setting                                                                                                                        = "osc_clk_div_by1",
parameter hssi_avmm1_if_0_hssiadapt_avmm_testbus_sel                                                                                                                             = "avmm1_transfer_testbus",
parameter hssi_avmm1_if_0_pldadapt_avmm_testbus_sel                                                                                                                              = "avmm1_transfer_testbus",
parameter hssi_avmm1_if_0_func_mode                                                                                                                                              = "c3adpt_pmadir",
parameter hssi_avmm1_if_0_hssiadapt_sr_hip_mode                                                                                                                                  = "disable_hip",
parameter hssi_avmm1_if_0_hssiadapt_hip_mode                                                                                                                                     = "disable_hip",
parameter hssi_avmm1_if_0_pldadapt_hip_mode                                                                                                                                      = "disable_hip",
parameter hssi_avmm1_if_0_hssiadapt_sr_powerdown_mode                                                                                                                            = "powerup",
parameter hssi_avmm1_if_0_hssiadapt_sr_sr_free_run_div_clk                                                                                                                       = "out_of_reset_sync",
parameter hssi_avmm1_if_0_hssiadapt_sr_sr_hip_en                                                                                                                                 = "disable",
parameter hssi_avmm1_if_0_hssiadapt_sr_sr_osc_clk_div_sel                                                                                                                        = "non_div",
parameter hssi_avmm1_if_0_hssiadapt_sr_sr_osc_clk_scg_en                                                                                                                         = "disable",
parameter hssi_avmm1_if_0_hssiadapt_sr_sr_parity_en                                                                                                                              = "disable",
parameter hssi_avmm1_if_0_hssiadapt_sr_sr_reserved_in_en                                                                                                                         = "enable",
parameter hssi_avmm1_if_0_hssiadapt_sr_sr_reserved_out_en                                                                                                                        = "enable",
parameter hssi_avmm1_if_0_hssiadapt_sr_sup_mode                                                                                                                                  = "user_mode",
parameter hssi_avmm1_if_0_topology                                                                                                                                               = "disabled_block",
parameter hssi_avmm1_if_0_calibration_type                                                                                                                                       = "one_time",
parameter hssi_avmm2_if_0_pcs_arbiter_ctrl                                                                                                                                       = "avmm2_arbiter_uc_sel",
parameter hssi_avmm2_if_0_hssiadapt_avmm_clk_dcg_en                                                                                                                              = "disable",
parameter hssi_avmm2_if_0_hssiadapt_avmm_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm2_if_0_pldadapt_avmm_clk_scg_en                                                                                                                               = "disable",
parameter hssi_avmm2_if_0_pcs_cal_done                                                                                                                                           = "avmm2_cal_done_assert",
parameter hssi_avmm2_if_0_pcs_cal_reserved                                                                                                                                       = 0,
parameter hssi_avmm2_if_0_pcs_calibration_feature_en                                                                                                                             = "avmm2_pcs_calibration_dis",
parameter hssi_avmm2_if_0_pldadapt_gate_dis                                                                                                                                      = "disable",
parameter hssi_avmm2_if_0_pcs_hip_cal_en                                                                                                                                         = "disable",
parameter hssi_avmm2_if_0_hssiadapt_osc_clk_scg_en                                                                                                                               = "disable",
parameter hssi_avmm2_if_0_pldadapt_osc_clk_scg_en                                                                                                                                = "disable",
parameter hssi_avmm2_if_0_hssiadapt_avmm_osc_clock_setting                                                                                                                       = "osc_clk_div_by1",
parameter hssi_avmm2_if_0_pldadapt_avmm_osc_clock_setting                                                                                                                        = "osc_clk_div_by1",
parameter hssi_avmm2_if_0_hssiadapt_avmm_testbus_sel                                                                                                                             = "avmm1_transfer_testbus",
parameter hssi_avmm2_if_0_pldadapt_avmm_testbus_sel                                                                                                                              = "avmm1_transfer_testbus",
parameter hssi_avmm2_if_0_func_mode                                                                                                                                              = "c3adpt_pmadir",
parameter hssi_avmm2_if_0_hssiadapt_hip_mode                                                                                                                                     = "disable_hip",
parameter hssi_avmm2_if_0_pldadapt_hip_mode                                                                                                                                      = "disable_hip",
parameter hssi_avmm2_if_0_topology                                                                                                                                               = "disabled_block",
parameter hssi_avmm2_if_0_calibration_type                                                                                                                                       = "one_time",
parameter hssi_aibnd_rx_13_aib_ber_margining_ctrl                                                                                                                                = "aib_ber_margining_setting0",
parameter hssi_aibnd_rx_13_aib_datasel_gr0                                                                                                                                       = "aib_datasel0_setting0",
parameter hssi_aibnd_rx_13_aib_datasel_gr1                                                                                                                                       = "aib_datasel1_setting1",
parameter hssi_aibnd_rx_13_aib_datasel_gr2                                                                                                                                       = "aib_datasel2_setting1",
parameter hssi_aibnd_rx_13_aib_dllstr_align_clkdiv                                                                                                                               = "aib_dllstr_align_clkdiv_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_dly_pst                                                                                                                              = "aib_dllstr_align_dly_pst_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_dy_ctl_static                                                                                                                        = "aib_dllstr_align_dy_ctl_static_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_dy_ctlsel                                                                                                                            = "aib_dllstr_align_dy_ctlsel_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_entest                                                                                                                               = "aib_dllstr_align_test_disable",
parameter hssi_aibnd_rx_13_aib_dllstr_align_halfcode                                                                                                                             = "aib_dllstr_align_halfcode_enable",
parameter hssi_aibnd_rx_13_aib_dllstr_align_selflock                                                                                                                             = "aib_dllstr_align_selflock_enable",
parameter hssi_aibnd_rx_13_aib_dllstr_align_st_core_dn_prgmnvrt                                                                                                                  = "aib_dllstr_align_st_core_dn_prgmnvrt_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_st_core_up_prgmnvrt                                                                                                                  = "aib_dllstr_align_st_core_up_prgmnvrt_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_st_core_updnen                                                                                                                       = "aib_dllstr_align_st_core_updnen_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_st_dftmuxsel                                                                                                                         = "aib_dllstr_align_st_dftmuxsel_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_st_en                                                                                                                                = "aib_dllstr_align_st_en_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_st_hps_ctrl_en                                                                                                                       = "aib_dllstr_align_hps_ctrl_en_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_st_lockreq_muxsel                                                                                                                    = "aib_dllstr_align_st_lockreq_muxsel_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_st_new_dll                                                                                                                           = "aib_dllstr_align_new_dll_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_st_rst                                                                                                                               = "aib_dllstr_align_st_rst_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_st_rst_prgmnvrt                                                                                                                      = "aib_dllstr_align_st_rst_prgmnvrt_setting0",
parameter hssi_aibnd_rx_13_aib_dllstr_align_test_clk_pll_en_n                                                                                                                    = "aib_dllstr_align_test_clk_pll_en_n_disable",
parameter hssi_aibnd_rx_13_aib_inctrl_gr0                                                                                                                                        = "aib_inctrl0_setting0",
parameter hssi_aibnd_rx_13_aib_inctrl_gr1                                                                                                                                        = "aib_inctrl1_setting0",
parameter hssi_aibnd_rx_13_aib_inctrl_gr2                                                                                                                                        = "aib_inctrl2_setting0",
parameter hssi_aibnd_rx_13_aib_inctrl_gr3                                                                                                                                        = "aib_inctrl3_setting0",
parameter hssi_aibnd_rx_13_aib_outctrl_gr0                                                                                                                                       = "aib_outen0_setting0",
parameter hssi_aibnd_rx_13_aib_outctrl_gr1                                                                                                                                       = "aib_outen1_setting0",
parameter hssi_aibnd_rx_13_aib_outctrl_gr2                                                                                                                                       = "aib_outen2_setting0",
parameter hssi_aibnd_rx_13_aib_outndrv_r12                                                                                                                                       = "aib_ndrv12_setting1",
parameter hssi_aibnd_rx_13_aib_outndrv_r34                                                                                                                                       = "aib_ndrv34_setting1",
parameter hssi_aibnd_rx_13_aib_outndrv_r56                                                                                                                                       = "aib_ndrv56_setting1",
parameter hssi_aibnd_rx_13_aib_outndrv_r78                                                                                                                                       = "aib_ndrv78_setting1",
parameter hssi_aibnd_rx_13_aib_outpdrv_r12                                                                                                                                       = "aib_pdrv12_setting1",
parameter hssi_aibnd_rx_13_aib_outpdrv_r34                                                                                                                                       = "aib_pdrv34_setting1",
parameter hssi_aibnd_rx_13_aib_outpdrv_r56                                                                                                                                       = "aib_pdrv56_setting1",
parameter hssi_aibnd_rx_13_aib_outpdrv_r78                                                                                                                                       = "aib_pdrv78_setting1",
parameter hssi_aibnd_rx_13_aib_red_shift_en                                                                                                                                      = "aib_red_shift_disable",
parameter hssi_aibnd_rx_13_dft_hssitestip_dll_dcc_en                                                                                                                             = "disable_dft",
parameter hssi_aibnd_rx_13_op_mode                                                                                                                                               = "pwr_down",
parameter hssi_aibnd_rx_13_powerdown_mode                                                                                                                                        = "true",
parameter hssi_aibnd_rx_13_powermode_ac                                                                                                                                          = "rxdatapath_low_speed_pwr",
parameter hssi_aibnd_rx_13_powermode_dc                                                                                                                                          = "rxdatapath_powerdown",
parameter hssi_aibnd_rx_13_powermode_freq_hz_aib_hssi_rx_transfer_clk                                                                                                            = 0,
parameter hssi_aibnd_rx_13_redundancy_en                                                                                                                                         = "disable",
parameter hssi_aibnd_rx_13_sup_mode                                                                                                                                              = "user_mode",
parameter hssi_aibnd_tx_13_aib_datasel_gr0                                                                                                                                       = "aib_datasel0_setting0",
parameter hssi_aibnd_tx_13_aib_datasel_gr1                                                                                                                                       = "aib_datasel1_setting0",
parameter hssi_aibnd_tx_13_aib_datasel_gr2                                                                                                                                       = "aib_datasel2_setting1",
parameter hssi_aibnd_tx_13_aib_datasel_gr3                                                                                                                                       = "aib_datasel3_setting1",
parameter hssi_aibnd_tx_13_aib_ddrctrl_gr0                                                                                                                                       = "aib_ddr0_setting1",
parameter hssi_aibnd_tx_13_aib_hssi_tx_transfer_clk_hz                                                                                                                           = 0,
parameter hssi_aibnd_tx_13_aib_iinasyncen                                                                                                                                        = "aib_inasyncen_setting0",
parameter hssi_aibnd_tx_13_aib_iinclken                                                                                                                                          = "aib_inclken_setting0",
parameter hssi_aibnd_tx_13_aib_outctrl_gr0                                                                                                                                       = "aib_outen0_setting0",
parameter hssi_aibnd_tx_13_aib_outctrl_gr1                                                                                                                                       = "aib_outen1_setting0",
parameter hssi_aibnd_tx_13_aib_outctrl_gr2                                                                                                                                       = "aib_outen2_setting0",
parameter hssi_aibnd_tx_13_aib_outctrl_gr3                                                                                                                                       = "aib_outen3_setting0",
parameter hssi_aibnd_tx_13_aib_outndrv_r34                                                                                                                                       = "aib_ndrv34_setting1",
parameter hssi_aibnd_tx_13_aib_outndrv_r56                                                                                                                                       = "aib_ndrv56_setting1",
parameter hssi_aibnd_tx_13_aib_outpdrv_r34                                                                                                                                       = "aib_pdrv34_setting1",
parameter hssi_aibnd_tx_13_aib_outpdrv_r56                                                                                                                                       = "aib_pdrv56_setting1",
parameter hssi_aibnd_tx_13_aib_red_dirclkn_shiften                                                                                                                               = "aib_red_dirclkn_shift_disable",
parameter hssi_aibnd_tx_13_aib_red_dirclkp_shiften                                                                                                                               = "aib_red_dirclkp_shift_disable",
parameter hssi_aibnd_tx_13_aib_red_drx_shiften                                                                                                                                   = "aib_red_drx_shift_disable",
parameter hssi_aibnd_tx_13_aib_red_dtx_shiften                                                                                                                                   = "aib_red_dtx_shift_disable",
parameter hssi_aibnd_tx_13_aib_red_pout_shiften                                                                                                                                  = "aib_red_pout_shift_disable",
parameter hssi_aibnd_tx_13_aib_red_rx_shiften                                                                                                                                    = "aib_red_rx_shift_disable",
parameter hssi_aibnd_tx_13_aib_red_tx_shiften                                                                                                                                    = "aib_red_tx_shift_disable",
parameter hssi_aibnd_tx_13_aib_red_txferclkout_shiften                                                                                                                           = "aib_red_txferclkout_shift_disable",
parameter hssi_aibnd_tx_13_aib_red_txferclkoutn_shiften                                                                                                                          = "aib_red_txferclkoutn_shift_disable",
parameter hssi_aibnd_tx_13_aib_tx_clkdiv                                                                                                                                         = "aib_tx_clkdiv_setting1",
parameter hssi_aibnd_tx_13_aib_tx_dcc_byp                                                                                                                                        = "aib_tx_dcc_byp_disable",
parameter hssi_aibnd_tx_13_aib_tx_dcc_byp_iocsr_unused                                                                                                                           = "aib_tx_dcc_byp_disable_iocsr_unused",
parameter hssi_aibnd_tx_13_aib_tx_dcc_cont_cal                                                                                                                                   = "aib_tx_dcc_cal_cont",
parameter hssi_aibnd_tx_13_aib_tx_dcc_cont_cal_iocsr_unused                                                                                                                      = "aib_tx_dcc_cal_single_iocsr_unused",
parameter hssi_aibnd_tx_13_aib_tx_dcc_dft                                                                                                                                        = "aib_tx_dcc_dft_disable",
parameter hssi_aibnd_tx_13_aib_tx_dcc_dft_sel                                                                                                                                    = "aib_tx_dcc_dft_mode0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_dll_dft_sel                                                                                                                                = "aib_tx_dcc_dll_dft_sel_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_dll_entest                                                                                                                                 = "aib_tx_dcc_dll_test_disable",
parameter hssi_aibnd_tx_13_aib_tx_dcc_dy_ctl_static                                                                                                                              = "aib_tx_dcc_dy_ctl_static_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_dy_ctlsel                                                                                                                                  = "aib_tx_dcc_dy_ctlsel_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_en                                                                                                                                         = "aib_tx_dcc_enable",
parameter hssi_aibnd_tx_13_aib_tx_dcc_en_iocsr_unused                                                                                                                            = "aib_tx_dcc_disable_iocsr_unused",
parameter hssi_aibnd_tx_13_aib_tx_dcc_manual_dn                                                                                                                                  = "aib_tx_dcc_manual_dn0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_manual_up                                                                                                                                  = "aib_tx_dcc_manual_up0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_rst_prgmnvrt                                                                                                                               = "aib_tx_dcc_st_rst_prgmnvrt_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_st_core_dn_prgmnvrt                                                                                                                        = "aib_tx_dcc_st_core_dn_prgmnvrt_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_st_core_up_prgmnvrt                                                                                                                        = "aib_tx_dcc_st_core_up_prgmnvrt_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_st_core_updnen                                                                                                                             = "aib_tx_dcc_st_core_updnen_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_st_dftmuxsel                                                                                                                               = "aib_tx_dcc_st_dftmuxsel_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_st_dly_pst                                                                                                                                 = "aib_tx_dcc_st_dly_pst_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_st_en                                                                                                                                      = "aib_tx_dcc_st_en_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_st_hps_ctrl_en                                                                                                                             = "aib_tx_dcc_hps_ctrl_en_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_st_lockreq_muxsel                                                                                                                          = "aib_tx_dcc_st_lockreq_muxsel_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_st_new_dll                                                                                                                                 = "aib_tx_dcc_new_dll_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_st_rst                                                                                                                                     = "aib_tx_dcc_st_rst_setting0",
parameter hssi_aibnd_tx_13_aib_tx_dcc_test_clk_pll_en_n                                                                                                                          = "aib_tx_dcc_test_clk_pll_en_n_disable",
parameter hssi_aibnd_tx_13_aib_tx_halfcode                                                                                                                                       = "aib_tx_halfcode_enable",
parameter hssi_aibnd_tx_13_aib_tx_selflock                                                                                                                                       = "aib_tx_selflock_enable",
parameter hssi_aibnd_tx_13_dfd_dll_dcc_en                                                                                                                                        = "disable_dfd",
parameter hssi_aibnd_tx_13_dft_hssitestip_dll_dcc_en                                                                                                                             = "disable_dft",
parameter hssi_aibnd_tx_13_op_mode                                                                                                                                               = "tx_dcc_enable",
parameter hssi_aibnd_tx_13_powerdown_mode                                                                                                                                        = "true",
parameter hssi_aibnd_tx_13_powermode_ac                                                                                                                                          = "txdatapath_low_speed_pwr",
parameter hssi_aibnd_tx_13_powermode_dc                                                                                                                                          = "txdatapath_powerdown",
parameter hssi_aibnd_tx_13_powermode_freq_hz_aib_hssi_tx_transfer_clk                                                                                                            = 0,
parameter hssi_aibnd_tx_13_redundancy_en                                                                                                                                         = "disable",
parameter hssi_aibnd_tx_13_sup_mode                                                                                                                                              = "user_mode",
parameter hssi_pldadapt_tx_13_aib_clk1_sel                                                                                                                                       = "aib_clk1_pld_pcs_tx_clk_out",
parameter hssi_pldadapt_tx_13_aib_clk2_sel                                                                                                                                       = "aib_clk2_pld_pcs_tx_clk_out",
parameter hssi_pldadapt_tx_13_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                                                              = 0,
parameter hssi_pldadapt_tx_13_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz                                                                                                            = 0,
parameter hssi_pldadapt_tx_13_hdpldadapt_aib_fabric_tx_sr_clk_in_hz                                                                                                              = 0,
parameter hssi_pldadapt_tx_13_bonding_dft_en                                                                                                                                     = "dft_dis",
parameter hssi_pldadapt_tx_13_bonding_dft_val                                                                                                                                    = "dft_0",
parameter hssi_pldadapt_tx_13_chnl_bonding                                                                                                                                       = "disable",
parameter hssi_pldadapt_tx_13_comp_cnt                                                                                                                                           = 0,
parameter hssi_pldadapt_tx_13_compin_sel                                                                                                                                         = "compin_master",
parameter hssi_pldadapt_tx_13_hdpldadapt_csr_clk_hz                                                                                                                              = 0,
parameter hssi_pldadapt_tx_13_ctrl_plane_bonding                                                                                                                                 = "individual",
parameter hssi_pldadapt_tx_13_ds_bypass_pipeln                                                                                                                                   = "ds_bypass_pipeln_dis",
parameter hssi_pldadapt_tx_13_ds_last_chnl                                                                                                                                       = "ds_not_last_chnl",
parameter hssi_pldadapt_tx_13_ds_master                                                                                                                                          = "ds_master_en",
parameter hssi_pldadapt_tx_13_duplex_mode                                                                                                                                        = "disable",
parameter hssi_pldadapt_tx_13_dv_bond                                                                                                                                            = "dv_bond_dis",
parameter hssi_pldadapt_tx_13_dv_gen                                                                                                                                             = "dv_gen_dis",
parameter hssi_pldadapt_tx_13_fifo_double_write                                                                                                                                  = "fifo_double_write_dis",
parameter hssi_pldadapt_tx_13_fifo_mode                                                                                                                                          = "phase_comp",
parameter hssi_pldadapt_tx_13_fifo_rd_clk_frm_gen_scg_en                                                                                                                         = "disable",
parameter hssi_pldadapt_tx_13_fifo_rd_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_13_fifo_rd_clk_sel                                                                                                                                    = "fifo_rd_pma_aib_tx_clk",
parameter hssi_pldadapt_tx_13_fifo_stop_rd                                                                                                                                       = "n_rd_empty",
parameter hssi_pldadapt_tx_13_fifo_stop_wr                                                                                                                                       = "n_wr_full",
parameter hssi_pldadapt_tx_13_fifo_width                                                                                                                                         = "fifo_single_width",
parameter hssi_pldadapt_tx_13_fifo_wr_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_13_fpll_shared_direct_async_in_sel                                                                                                                    = "fpll_shared_direct_async_in_rowclk",
parameter hssi_pldadapt_tx_13_frmgen_burst                                                                                                                                       = "frmgen_burst_dis",
parameter hssi_pldadapt_tx_13_frmgen_bypass                                                                                                                                      = "frmgen_bypass_dis",
parameter hssi_pldadapt_tx_13_frmgen_mfrm_length                                                                                                                                 = 2048,
parameter hssi_pldadapt_tx_13_frmgen_pipeln                                                                                                                                      = "frmgen_pipeln_dis",
parameter hssi_pldadapt_tx_13_frmgen_pyld_ins                                                                                                                                    = "frmgen_pyld_ins_dis",
parameter hssi_pldadapt_tx_13_frmgen_wordslip                                                                                                                                    = "frmgen_wordslip_dis",
parameter hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit0_rst_val                                                                                                                        = "reset_to_zero_hfsrin0",
parameter hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit1_rst_val                                                                                                                        = "reset_to_zero_hfsrin1",
parameter hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit2_rst_val                                                                                                                        = "reset_to_zero_hfsrin2",
parameter hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit3_rst_val                                                                                                                        = "reset_to_zero_hfsrin3",
parameter hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit0_rst_val                                                                                                                       = "reset_to_zero_hfsrout0",
parameter hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit1_rst_val                                                                                                                       = "reset_to_zero_hfsrout1",
parameter hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit2_rst_val                                                                                                                       = "reset_to_zero_hfsrout2",
parameter hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit3_rst_val                                                                                                                       = "reset_to_zero_hfsrout3",
parameter hssi_pldadapt_tx_13_fsr_mask_tx_pll_rst_val                                                                                                                            = "reset_to_zero_maskpll",
parameter hssi_pldadapt_tx_13_fsr_pld_txelecidle_rst_val                                                                                                                         = "reset_to_zero_txelec",
parameter hssi_pldadapt_tx_13_gb_tx_idwidth                                                                                                                                      = "idwidth_66",
parameter hssi_pldadapt_tx_13_gb_tx_odwidth                                                                                                                                      = "odwidth_32",
parameter hssi_pldadapt_tx_13_hip_mode                                                                                                                                           = "disable_hip",
parameter hssi_pldadapt_tx_13_hip_osc_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_13_hrdrst_dcd_cal_done_bypass                                                                                                                         = "disable",
parameter hssi_pldadapt_tx_13_hrdrst_rst_sm_dis                                                                                                                                  = "enable_tx_rst_sm",
parameter hssi_pldadapt_tx_13_hrdrst_rx_osc_clk_scg_en                                                                                                                           = "disable",
parameter hssi_pldadapt_tx_13_hrdrst_user_ctl_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_13_indv                                                                                                                                               = "indv_en",
parameter hssi_pldadapt_tx_13_is_paired_with                                                                                                                                     = "other",
parameter hssi_pldadapt_tx_13_loopback_mode                                                                                                                                      = "disable",
parameter hssi_pldadapt_tx_13_low_latency_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_tx_13_osc_clk_scg_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_tx_13_phcomp_rd_del                                                                                                                                      = "phcomp_rd_del2",
parameter hssi_pldadapt_tx_13_pipe_mode                                                                                                                                          = "disable_pipe",
parameter hssi_pldadapt_tx_13_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_tx_13_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_tx_13_pld_clk1_delay_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_tx_13_pld_clk1_delay_sel                                                                                                                                 = "delay_path0",
parameter hssi_pldadapt_tx_13_pld_clk1_inv_en                                                                                                                                    = "disable",
parameter hssi_pldadapt_tx_13_pld_clk1_sel                                                                                                                                       = "pld_clk1_rowclk",
parameter hssi_pldadapt_tx_13_pld_clk2_sel                                                                                                                                       = "pld_clk2_rowclk",
parameter hssi_pldadapt_tx_13_hdpldadapt_pld_sclk1_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_tx_13_hdpldadapt_pld_sclk2_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk1_dcm_hz                                                                                                                      = 0,
parameter hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk1_rowclk_hz                                                                                                                   = 0,
parameter hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk2_dcm_hz                                                                                                                      = 0,
parameter hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk2_rowclk_hz                                                                                                                   = 0,
parameter hssi_pldadapt_tx_13_pma_aib_tx_clk_expected_setting                                                                                                                    = "not_used",
parameter hssi_pldadapt_tx_13_powerdown_mode                                                                                                                                     = "powerdown",
parameter hssi_pldadapt_tx_13_powermode_dc                                                                                                                                       = "powerdown",
parameter hssi_pldadapt_tx_13_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                                                          = 0,
parameter hssi_pldadapt_tx_13_powermode_freq_hz_pld_tx_clk1_dcm                                                                                                                  = 0,
parameter hssi_pldadapt_tx_13_sh_err                                                                                                                                             = "sh_err_dis",
parameter hssi_pldadapt_tx_13_hdpldadapt_speed_grade                                                                                                                             = "dash_1",
parameter hssi_pldadapt_tx_13_hdpldadapt_sr_sr_testbus_sel                                                                                                                       = "ssr_testbus",
parameter hssi_pldadapt_tx_13_stretch_num_stages                                                                                                                                 = "zero_stage",
parameter hssi_pldadapt_tx_13_sup_mode                                                                                                                                           = "user_mode",
parameter hssi_pldadapt_tx_13_tx_datapath_tb_sel                                                                                                                                 = "cp_bond",
parameter hssi_pldadapt_tx_13_tx_fastbond_rden                                                                                                                                   = "rden_ds_del_us_del",
parameter hssi_pldadapt_tx_13_tx_fastbond_wren                                                                                                                                   = "wren_ds_del_us_del",
parameter hssi_pldadapt_tx_13_tx_fifo_power_mode                                                                                                                                 = "full_width_full_depth",
parameter hssi_pldadapt_tx_13_tx_fifo_read_latency_adjust                                                                                                                        = "disable",
parameter hssi_pldadapt_tx_13_tx_fifo_write_latency_adjust                                                                                                                       = "disable",
parameter hssi_pldadapt_tx_13_tx_hip_aib_ssr_in_polling_bypass                                                                                                                   = "disable",
parameter hssi_pldadapt_tx_13_tx_osc_clock_setting                                                                                                                               = "osc_clk_div_by1",
parameter hssi_pldadapt_tx_13_tx_pld_10g_tx_bitslip_polling_bypass                                                                                                               = "disable",
parameter hssi_pldadapt_tx_13_tx_pld_8g_tx_boundary_sel_polling_bypass                                                                                                           = "disable",
parameter hssi_pldadapt_tx_13_tx_pld_pma_fpll_cnt_sel_polling_bypass                                                                                                             = "disable",
parameter hssi_pldadapt_tx_13_tx_pld_pma_fpll_num_phase_shifts_polling_bypass                                                                                                    = "disable",
parameter hssi_pldadapt_tx_13_tx_usertest_sel                                                                                                                                    = "enable",
parameter hssi_pldadapt_tx_13_txfifo_empty                                                                                                                                       = "empty_default",
parameter hssi_pldadapt_tx_13_txfifo_full                                                                                                                                        = "full_pc_sw",
parameter hssi_pldadapt_tx_13_txfifo_mode                                                                                                                                        = "txphase_comp",
parameter hssi_pldadapt_tx_13_txfifo_pempty                                                                                                                                      = 2,
parameter hssi_pldadapt_tx_13_txfifo_pfull                                                                                                                                       = 24,
parameter hssi_pldadapt_tx_13_us_bypass_pipeln                                                                                                                                   = "us_bypass_pipeln_dis",
parameter hssi_pldadapt_tx_13_us_last_chnl                                                                                                                                       = "us_not_last_chnl",
parameter hssi_pldadapt_tx_13_us_master                                                                                                                                          = "us_master_en",
parameter hssi_pldadapt_tx_13_word_align_enable                                                                                                                                  = "disable",
parameter hssi_pldadapt_tx_13_word_mark                                                                                                                                          = "wm_en",
parameter hssi_pldadapt_tx_13_reconfig_settings                                                                                                                                  = "{}",
parameter hssi_pldadapt_rx_13_aib_clk1_sel                                                                                                                                       = "aib_clk1_rx_transfer_clk",
parameter hssi_pldadapt_rx_13_aib_clk2_sel                                                                                                                                       = "aib_clk2_rx_transfer_clk",
parameter hssi_pldadapt_rx_13_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                                                              = 0,
parameter hssi_pldadapt_rx_13_hdpldadapt_aib_fabric_rx_sr_clk_in_hz                                                                                                              = 0,
parameter hssi_pldadapt_rx_13_hdpldadapt_aib_fabric_rx_transfer_clk_hz                                                                                                           = 0,
parameter hssi_pldadapt_rx_13_asn_bypass_pma_pcie_sw_done                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_13_asn_en                                                                                                                                             = "disable",
parameter hssi_pldadapt_rx_13_asn_wait_for_dll_reset_cnt                                                                                                                         = 0,
parameter hssi_pldadapt_rx_13_asn_wait_for_fifo_flush_cnt                                                                                                                        = 0,
parameter hssi_pldadapt_rx_13_asn_wait_for_pma_pcie_sw_done_cnt                                                                                                                  = 0,
parameter hssi_pldadapt_rx_13_bonding_dft_en                                                                                                                                     = "dft_dis",
parameter hssi_pldadapt_rx_13_bonding_dft_val                                                                                                                                    = "dft_0",
parameter hssi_pldadapt_rx_13_chnl_bonding                                                                                                                                       = "disable",
parameter hssi_pldadapt_rx_13_clock_del_measure_enable                                                                                                                           = "disable",
parameter hssi_pldadapt_rx_13_comp_cnt                                                                                                                                           = 0,
parameter hssi_pldadapt_rx_13_compin_sel                                                                                                                                         = "compin_master",
parameter hssi_pldadapt_rx_13_hdpldadapt_csr_clk_hz                                                                                                                              = 0,
parameter hssi_pldadapt_rx_13_ctrl_plane_bonding                                                                                                                                 = "individual",
parameter hssi_pldadapt_rx_13_ds_bypass_pipeln                                                                                                                                   = "ds_bypass_pipeln_dis",
parameter hssi_pldadapt_rx_13_ds_last_chnl                                                                                                                                       = "ds_not_last_chnl",
parameter hssi_pldadapt_rx_13_ds_master                                                                                                                                          = "ds_master_en",
parameter hssi_pldadapt_rx_13_duplex_mode                                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_13_dv_mode                                                                                                                                            = "dv_mode_dis",
parameter hssi_pldadapt_rx_13_fifo_double_read                                                                                                                                   = "fifo_double_read_dis",
parameter hssi_pldadapt_rx_13_fifo_mode                                                                                                                                          = "phase_comp",
parameter hssi_pldadapt_rx_13_fifo_rd_clk_ins_sm_scg_en                                                                                                                          = "disable",
parameter hssi_pldadapt_rx_13_fifo_rd_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_13_fifo_rd_clk_sel                                                                                                                                    = "fifo_rd_clk_rx_transfer_clk",
parameter hssi_pldadapt_rx_13_fifo_stop_rd                                                                                                                                       = "n_rd_empty",
parameter hssi_pldadapt_rx_13_fifo_stop_wr                                                                                                                                       = "n_wr_full",
parameter hssi_pldadapt_rx_13_fifo_width                                                                                                                                         = "fifo_single_width",
parameter hssi_pldadapt_rx_13_fifo_wr_clk_del_sm_scg_en                                                                                                                          = "disable",
parameter hssi_pldadapt_rx_13_fifo_wr_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_13_fifo_wr_clk_sel                                                                                                                                    = "fifo_wr_clk_rx_transfer_clk",
parameter hssi_pldadapt_rx_13_free_run_div_clk                                                                                                                                   = "out_of_reset_sync",
parameter hssi_pldadapt_rx_13_fsr_pld_10g_rx_crc32_err_rst_val                                                                                                                   = "reset_to_zero_crc32",
parameter hssi_pldadapt_rx_13_fsr_pld_8g_sigdet_out_rst_val                                                                                                                      = "reset_to_zero_sigdet",
parameter hssi_pldadapt_rx_13_fsr_pld_ltd_b_rst_val                                                                                                                              = "reset_to_zero_ltdb",
parameter hssi_pldadapt_rx_13_fsr_pld_ltr_rst_val                                                                                                                                = "reset_to_zero_ltr",
parameter hssi_pldadapt_rx_13_fsr_pld_rx_fifo_align_clr_rst_val                                                                                                                  = "reset_to_zero_alignclr",
parameter hssi_pldadapt_rx_13_gb_rx_idwidth                                                                                                                                      = "idwidth_32",
parameter hssi_pldadapt_rx_13_gb_rx_odwidth                                                                                                                                      = "odwidth_66",
parameter hssi_pldadapt_rx_13_hip_mode                                                                                                                                           = "disable_hip",
parameter hssi_pldadapt_rx_13_hrdrst_align_bypass                                                                                                                                = "disable",
parameter hssi_pldadapt_rx_13_hrdrst_dll_lock_bypass                                                                                                                             = "disable",
parameter hssi_pldadapt_rx_13_hrdrst_rst_sm_dis                                                                                                                                  = "enable_rx_rst_sm",
parameter hssi_pldadapt_rx_13_hrdrst_rx_osc_clk_scg_en                                                                                                                           = "disable",
parameter hssi_pldadapt_rx_13_hrdrst_user_ctl_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_13_indv                                                                                                                                               = "indv_en",
parameter hssi_pldadapt_rx_13_internal_clk1_sel1                                                                                                                                 = "pma_clks_or_txfiford_post_ct_mux_clk1_mux1",
parameter hssi_pldadapt_rx_13_internal_clk1_sel2                                                                                                                                 = "pma_clks_clk1_mux2",
parameter hssi_pldadapt_rx_13_internal_clk2_sel1                                                                                                                                 = "pma_clks_or_rxfifowr_post_ct_mux_clk2_mux1",
parameter hssi_pldadapt_rx_13_internal_clk2_sel2                                                                                                                                 = "pma_clks_clk2_mux2",
parameter hssi_pldadapt_rx_13_is_paired_with                                                                                                                                     = "other",
parameter hssi_pldadapt_rx_13_loopback_mode                                                                                                                                      = "disable",
parameter hssi_pldadapt_rx_13_low_latency_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_rx_13_lpbk_mode                                                                                                                                          = "disable",
parameter hssi_pldadapt_rx_13_osc_clk_scg_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_rx_13_phcomp_rd_del                                                                                                                                      = "phcomp_rd_del2",
parameter hssi_pldadapt_rx_13_pipe_enable                                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_13_pipe_mode                                                                                                                                          = "disable_pipe",
parameter hssi_pldadapt_rx_13_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_rx_13_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_rx_13_pld_clk1_delay_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_rx_13_pld_clk1_delay_sel                                                                                                                                 = "delay_path0",
parameter hssi_pldadapt_rx_13_pld_clk1_inv_en                                                                                                                                    = "disable",
parameter hssi_pldadapt_rx_13_pld_clk1_sel                                                                                                                                       = "pld_clk1_rowclk",
parameter hssi_pldadapt_rx_13_hdpldadapt_pld_rx_clk1_dcm_hz                                                                                                                      = 0,
parameter hssi_pldadapt_rx_13_hdpldadapt_pld_rx_clk1_rowclk_hz                                                                                                                   = 0,
parameter hssi_pldadapt_rx_13_hdpldadapt_pld_sclk1_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_rx_13_hdpldadapt_pld_sclk2_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_rx_13_pma_hclk_scg_en                                                                                                                                    = "disable",
parameter hssi_pldadapt_rx_13_powerdown_mode                                                                                                                                     = "powerdown",
parameter hssi_pldadapt_rx_13_powermode_dc                                                                                                                                       = "powerdown",
parameter hssi_pldadapt_rx_13_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                                                          = 0,
parameter hssi_pldadapt_rx_13_powermode_freq_hz_pld_rx_clk1_dcm                                                                                                                  = 0,
parameter hssi_pldadapt_rx_13_rx_datapath_tb_sel                                                                                                                                 = "cp_bond",
parameter hssi_pldadapt_rx_13_rx_fastbond_rden                                                                                                                                   = "rden_ds_del_us_del",
parameter hssi_pldadapt_rx_13_rx_fastbond_wren                                                                                                                                   = "wren_ds_del_us_del",
parameter hssi_pldadapt_rx_13_rx_fifo_power_mode                                                                                                                                 = "full_width_full_depth",
parameter hssi_pldadapt_rx_13_rx_fifo_read_latency_adjust                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_13_rx_fifo_write_ctrl                                                                                                                                 = "blklock_stops",
parameter hssi_pldadapt_rx_13_rx_fifo_write_latency_adjust                                                                                                                       = "disable",
parameter hssi_pldadapt_rx_13_rx_osc_clock_setting                                                                                                                               = "osc_clk_div_by1",
parameter hssi_pldadapt_rx_13_rx_pld_8g_eidleinfersel_polling_bypass                                                                                                             = "disable",
parameter hssi_pldadapt_rx_13_rx_pld_pma_eye_monitor_polling_bypass                                                                                                              = "disable",
parameter hssi_pldadapt_rx_13_rx_pld_pma_pcie_switch_polling_bypass                                                                                                              = "disable",
parameter hssi_pldadapt_rx_13_rx_pld_pma_reser_out_polling_bypass                                                                                                                = "disable",
parameter hssi_pldadapt_rx_13_rx_prbs_flags_sr_enable                                                                                                                            = "disable",
parameter hssi_pldadapt_rx_13_rx_true_b2b                                                                                                                                        = "b2b",
parameter hssi_pldadapt_rx_13_rx_usertest_sel                                                                                                                                    = "enable",
parameter hssi_pldadapt_rx_13_rxfifo_empty                                                                                                                                       = "empty_sw",
parameter hssi_pldadapt_rx_13_rxfifo_full                                                                                                                                        = "full_pc_sw",
parameter hssi_pldadapt_rx_13_rxfifo_mode                                                                                                                                        = "rxphase_comp",
parameter hssi_pldadapt_rx_13_rxfifo_pempty                                                                                                                                      = 2,
parameter hssi_pldadapt_rx_13_rxfifo_pfull                                                                                                                                       = 48,
parameter hssi_pldadapt_rx_13_rxfiford_post_ct_sel                                                                                                                               = "rxfiford_sclk_post_ct",
parameter hssi_pldadapt_rx_13_rxfifowr_post_ct_sel                                                                                                                               = "rxfifowr_sclk_post_ct",
parameter hssi_pldadapt_rx_13_sclk_sel                                                                                                                                           = "sclk1_rowclk",
parameter hssi_pldadapt_rx_13_hdpldadapt_speed_grade                                                                                                                             = "dash_1",
parameter hssi_pldadapt_rx_13_hdpldadapt_sr_sr_testbus_sel                                                                                                                       = "ssr_testbus",
parameter hssi_pldadapt_rx_13_stretch_num_stages                                                                                                                                 = "zero_stage",
parameter hssi_pldadapt_rx_13_sup_mode                                                                                                                                           = "user_mode",
parameter hssi_pldadapt_rx_13_txfiford_post_ct_sel                                                                                                                               = "txfiford_sclk_post_ct",
parameter hssi_pldadapt_rx_13_txfifowr_post_ct_sel                                                                                                                               = "txfifowr_sclk_post_ct",
parameter hssi_pldadapt_rx_13_us_bypass_pipeln                                                                                                                                   = "us_bypass_pipeln_dis",
parameter hssi_pldadapt_rx_13_us_last_chnl                                                                                                                                       = "us_not_last_chnl",
parameter hssi_pldadapt_rx_13_us_master                                                                                                                                          = "us_master_en",
parameter hssi_pldadapt_rx_13_word_align                                                                                                                                         = "wa_en",
parameter hssi_pldadapt_rx_13_word_align_enable                                                                                                                                  = "disable",
parameter hssi_pldadapt_rx_13_reconfig_settings                                                                                                                                  = "{}",
parameter hssi_avmm1_if_13_pcs_arbiter_ctrl                                                                                                                                      = "avmm1_arbiter_uc_sel",
parameter hssi_avmm1_if_13_hssiadapt_avmm_clk_dcg_en                                                                                                                             = "disable",
parameter hssi_avmm1_if_13_hssiadapt_avmm_clk_scg_en                                                                                                                             = "disable",
parameter hssi_avmm1_if_13_pldadapt_avmm_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm1_if_13_pcs_cal_done                                                                                                                                          = "avmm1_cal_done_assert",
parameter hssi_avmm1_if_13_pcs_cal_reserved                                                                                                                                      = 0,
parameter hssi_avmm1_if_13_pcs_calibration_feature_en                                                                                                                            = "avmm1_pcs_calibration_dis",
parameter hssi_avmm1_if_13_pldadapt_gate_dis                                                                                                                                     = "disable",
parameter hssi_avmm1_if_13_pcs_hip_cal_en                                                                                                                                        = "disable",
parameter hssi_avmm1_if_13_hssiadapt_nfhssi_calibratio_feature_en                                                                                                                = "disable",
parameter hssi_avmm1_if_13_pldadapt_nfhssi_calibratio_feature_en                                                                                                                 = "disable",
parameter hssi_avmm1_if_13_hssiadapt_osc_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm1_if_13_pldadapt_osc_clk_scg_en                                                                                                                               = "disable",
parameter hssi_avmm1_if_13_hssiadapt_read_blocking_enable                                                                                                                        = "enable",
parameter hssi_avmm1_if_13_pldadapt_read_blocking_enable                                                                                                                         = "enable",
parameter hssi_avmm1_if_13_hssiadapt_uc_blocking_enable                                                                                                                          = "enable",
parameter hssi_avmm1_if_13_pldadapt_uc_blocking_enable                                                                                                                           = "enable",
parameter hssi_avmm1_if_13_hssiadapt_write_resp_en                                                                                                                               = "disable",
parameter hssi_avmm1_if_13_hssiadapt_avmm_osc_clock_setting                                                                                                                      = "osc_clk_div_by1",
parameter hssi_avmm1_if_13_pldadapt_avmm_osc_clock_setting                                                                                                                       = "osc_clk_div_by1",
parameter hssi_avmm1_if_13_hssiadapt_avmm_testbus_sel                                                                                                                            = "avmm1_transfer_testbus",
parameter hssi_avmm1_if_13_pldadapt_avmm_testbus_sel                                                                                                                             = "avmm1_transfer_testbus",
parameter hssi_avmm1_if_13_func_mode                                                                                                                                             = "c3adpt_pmadir",
parameter hssi_avmm1_if_13_hssiadapt_sr_hip_mode                                                                                                                                 = "disable_hip",
parameter hssi_avmm1_if_13_hssiadapt_hip_mode                                                                                                                                    = "disable_hip",
parameter hssi_avmm1_if_13_pldadapt_hip_mode                                                                                                                                     = "disable_hip",
parameter hssi_avmm1_if_13_hssiadapt_sr_powerdown_mode                                                                                                                           = "powerup",
parameter hssi_avmm1_if_13_hssiadapt_sr_sr_free_run_div_clk                                                                                                                      = "out_of_reset_sync",
parameter hssi_avmm1_if_13_hssiadapt_sr_sr_hip_en                                                                                                                                = "disable",
parameter hssi_avmm1_if_13_hssiadapt_sr_sr_osc_clk_div_sel                                                                                                                       = "non_div",
parameter hssi_avmm1_if_13_hssiadapt_sr_sr_osc_clk_scg_en                                                                                                                        = "disable",
parameter hssi_avmm1_if_13_hssiadapt_sr_sr_parity_en                                                                                                                             = "disable",
parameter hssi_avmm1_if_13_hssiadapt_sr_sr_reserved_in_en                                                                                                                        = "enable",
parameter hssi_avmm1_if_13_hssiadapt_sr_sr_reserved_out_en                                                                                                                       = "enable",
parameter hssi_avmm1_if_13_hssiadapt_sr_sup_mode                                                                                                                                 = "user_mode",
parameter hssi_avmm1_if_13_topology                                                                                                                                              = "disabled_block",
parameter hssi_avmm1_if_13_calibration_type                                                                                                                                      = "one_time",
parameter hssi_avmm2_if_13_pcs_arbiter_ctrl                                                                                                                                      = "avmm2_arbiter_uc_sel",
parameter hssi_avmm2_if_13_hssiadapt_avmm_clk_dcg_en                                                                                                                             = "disable",
parameter hssi_avmm2_if_13_hssiadapt_avmm_clk_scg_en                                                                                                                             = "disable",
parameter hssi_avmm2_if_13_pldadapt_avmm_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm2_if_13_pcs_cal_done                                                                                                                                          = "avmm2_cal_done_assert",
parameter hssi_avmm2_if_13_pcs_cal_reserved                                                                                                                                      = 0,
parameter hssi_avmm2_if_13_pcs_calibration_feature_en                                                                                                                            = "avmm2_pcs_calibration_dis",
parameter hssi_avmm2_if_13_pldadapt_gate_dis                                                                                                                                     = "disable",
parameter hssi_avmm2_if_13_pcs_hip_cal_en                                                                                                                                        = "disable",
parameter hssi_avmm2_if_13_hssiadapt_osc_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm2_if_13_pldadapt_osc_clk_scg_en                                                                                                                               = "disable",
parameter hssi_avmm2_if_13_hssiadapt_avmm_osc_clock_setting                                                                                                                      = "osc_clk_div_by1",
parameter hssi_avmm2_if_13_pldadapt_avmm_osc_clock_setting                                                                                                                       = "osc_clk_div_by1",
parameter hssi_avmm2_if_13_hssiadapt_avmm_testbus_sel                                                                                                                            = "avmm1_transfer_testbus",
parameter hssi_avmm2_if_13_pldadapt_avmm_testbus_sel                                                                                                                             = "avmm1_transfer_testbus",
parameter hssi_avmm2_if_13_func_mode                                                                                                                                             = "c3adpt_pmadir",
parameter hssi_avmm2_if_13_hssiadapt_hip_mode                                                                                                                                    = "disable_hip",
parameter hssi_avmm2_if_13_pldadapt_hip_mode                                                                                                                                     = "disable_hip",
parameter hssi_avmm2_if_13_topology                                                                                                                                              = "disabled_block",
parameter hssi_avmm2_if_13_calibration_type                                                                                                                                      = "one_time",
parameter hssi_aibnd_rx_15_aib_ber_margining_ctrl                                                                                                                                = "aib_ber_margining_setting0",
parameter hssi_aibnd_rx_15_aib_datasel_gr0                                                                                                                                       = "aib_datasel0_setting0",
parameter hssi_aibnd_rx_15_aib_datasel_gr1                                                                                                                                       = "aib_datasel1_setting1",
parameter hssi_aibnd_rx_15_aib_datasel_gr2                                                                                                                                       = "aib_datasel2_setting1",
parameter hssi_aibnd_rx_15_aib_dllstr_align_clkdiv                                                                                                                               = "aib_dllstr_align_clkdiv_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_dly_pst                                                                                                                              = "aib_dllstr_align_dly_pst_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_dy_ctl_static                                                                                                                        = "aib_dllstr_align_dy_ctl_static_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_dy_ctlsel                                                                                                                            = "aib_dllstr_align_dy_ctlsel_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_entest                                                                                                                               = "aib_dllstr_align_test_disable",
parameter hssi_aibnd_rx_15_aib_dllstr_align_halfcode                                                                                                                             = "aib_dllstr_align_halfcode_enable",
parameter hssi_aibnd_rx_15_aib_dllstr_align_selflock                                                                                                                             = "aib_dllstr_align_selflock_enable",
parameter hssi_aibnd_rx_15_aib_dllstr_align_st_core_dn_prgmnvrt                                                                                                                  = "aib_dllstr_align_st_core_dn_prgmnvrt_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_st_core_up_prgmnvrt                                                                                                                  = "aib_dllstr_align_st_core_up_prgmnvrt_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_st_core_updnen                                                                                                                       = "aib_dllstr_align_st_core_updnen_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_st_dftmuxsel                                                                                                                         = "aib_dllstr_align_st_dftmuxsel_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_st_en                                                                                                                                = "aib_dllstr_align_st_en_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_st_hps_ctrl_en                                                                                                                       = "aib_dllstr_align_hps_ctrl_en_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_st_lockreq_muxsel                                                                                                                    = "aib_dllstr_align_st_lockreq_muxsel_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_st_new_dll                                                                                                                           = "aib_dllstr_align_new_dll_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_st_rst                                                                                                                               = "aib_dllstr_align_st_rst_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_st_rst_prgmnvrt                                                                                                                      = "aib_dllstr_align_st_rst_prgmnvrt_setting0",
parameter hssi_aibnd_rx_15_aib_dllstr_align_test_clk_pll_en_n                                                                                                                    = "aib_dllstr_align_test_clk_pll_en_n_disable",
parameter hssi_aibnd_rx_15_aib_inctrl_gr0                                                                                                                                        = "aib_inctrl0_setting0",
parameter hssi_aibnd_rx_15_aib_inctrl_gr1                                                                                                                                        = "aib_inctrl1_setting0",
parameter hssi_aibnd_rx_15_aib_inctrl_gr2                                                                                                                                        = "aib_inctrl2_setting0",
parameter hssi_aibnd_rx_15_aib_inctrl_gr3                                                                                                                                        = "aib_inctrl3_setting0",
parameter hssi_aibnd_rx_15_aib_outctrl_gr0                                                                                                                                       = "aib_outen0_setting0",
parameter hssi_aibnd_rx_15_aib_outctrl_gr1                                                                                                                                       = "aib_outen1_setting0",
parameter hssi_aibnd_rx_15_aib_outctrl_gr2                                                                                                                                       = "aib_outen2_setting0",
parameter hssi_aibnd_rx_15_aib_outndrv_r12                                                                                                                                       = "aib_ndrv12_setting1",
parameter hssi_aibnd_rx_15_aib_outndrv_r34                                                                                                                                       = "aib_ndrv34_setting1",
parameter hssi_aibnd_rx_15_aib_outndrv_r56                                                                                                                                       = "aib_ndrv56_setting1",
parameter hssi_aibnd_rx_15_aib_outndrv_r78                                                                                                                                       = "aib_ndrv78_setting1",
parameter hssi_aibnd_rx_15_aib_outpdrv_r12                                                                                                                                       = "aib_pdrv12_setting1",
parameter hssi_aibnd_rx_15_aib_outpdrv_r34                                                                                                                                       = "aib_pdrv34_setting1",
parameter hssi_aibnd_rx_15_aib_outpdrv_r56                                                                                                                                       = "aib_pdrv56_setting1",
parameter hssi_aibnd_rx_15_aib_outpdrv_r78                                                                                                                                       = "aib_pdrv78_setting1",
parameter hssi_aibnd_rx_15_aib_red_shift_en                                                                                                                                      = "aib_red_shift_disable",
parameter hssi_aibnd_rx_15_dft_hssitestip_dll_dcc_en                                                                                                                             = "disable_dft",
parameter hssi_aibnd_rx_15_op_mode                                                                                                                                               = "pwr_down",
parameter hssi_aibnd_rx_15_powerdown_mode                                                                                                                                        = "true",
parameter hssi_aibnd_rx_15_powermode_ac                                                                                                                                          = "rxdatapath_low_speed_pwr",
parameter hssi_aibnd_rx_15_powermode_dc                                                                                                                                          = "rxdatapath_powerdown",
parameter hssi_aibnd_rx_15_powermode_freq_hz_aib_hssi_rx_transfer_clk                                                                                                            = 0,
parameter hssi_aibnd_rx_15_redundancy_en                                                                                                                                         = "disable",
parameter hssi_aibnd_rx_15_sup_mode                                                                                                                                              = "user_mode",
parameter hssi_aibnd_tx_15_aib_datasel_gr0                                                                                                                                       = "aib_datasel0_setting0",
parameter hssi_aibnd_tx_15_aib_datasel_gr1                                                                                                                                       = "aib_datasel1_setting0",
parameter hssi_aibnd_tx_15_aib_datasel_gr2                                                                                                                                       = "aib_datasel2_setting1",
parameter hssi_aibnd_tx_15_aib_datasel_gr3                                                                                                                                       = "aib_datasel3_setting1",
parameter hssi_aibnd_tx_15_aib_ddrctrl_gr0                                                                                                                                       = "aib_ddr0_setting1",
parameter hssi_aibnd_tx_15_aib_hssi_tx_transfer_clk_hz                                                                                                                           = 0,
parameter hssi_aibnd_tx_15_aib_iinasyncen                                                                                                                                        = "aib_inasyncen_setting0",
parameter hssi_aibnd_tx_15_aib_iinclken                                                                                                                                          = "aib_inclken_setting0",
parameter hssi_aibnd_tx_15_aib_outctrl_gr0                                                                                                                                       = "aib_outen0_setting0",
parameter hssi_aibnd_tx_15_aib_outctrl_gr1                                                                                                                                       = "aib_outen1_setting0",
parameter hssi_aibnd_tx_15_aib_outctrl_gr2                                                                                                                                       = "aib_outen2_setting0",
parameter hssi_aibnd_tx_15_aib_outctrl_gr3                                                                                                                                       = "aib_outen3_setting0",
parameter hssi_aibnd_tx_15_aib_outndrv_r34                                                                                                                                       = "aib_ndrv34_setting1",
parameter hssi_aibnd_tx_15_aib_outndrv_r56                                                                                                                                       = "aib_ndrv56_setting1",
parameter hssi_aibnd_tx_15_aib_outpdrv_r34                                                                                                                                       = "aib_pdrv34_setting1",
parameter hssi_aibnd_tx_15_aib_outpdrv_r56                                                                                                                                       = "aib_pdrv56_setting1",
parameter hssi_aibnd_tx_15_aib_red_dirclkn_shiften                                                                                                                               = "aib_red_dirclkn_shift_disable",
parameter hssi_aibnd_tx_15_aib_red_dirclkp_shiften                                                                                                                               = "aib_red_dirclkp_shift_disable",
parameter hssi_aibnd_tx_15_aib_red_drx_shiften                                                                                                                                   = "aib_red_drx_shift_disable",
parameter hssi_aibnd_tx_15_aib_red_dtx_shiften                                                                                                                                   = "aib_red_dtx_shift_disable",
parameter hssi_aibnd_tx_15_aib_red_pout_shiften                                                                                                                                  = "aib_red_pout_shift_disable",
parameter hssi_aibnd_tx_15_aib_red_rx_shiften                                                                                                                                    = "aib_red_rx_shift_disable",
parameter hssi_aibnd_tx_15_aib_red_tx_shiften                                                                                                                                    = "aib_red_tx_shift_disable",
parameter hssi_aibnd_tx_15_aib_red_txferclkout_shiften                                                                                                                           = "aib_red_txferclkout_shift_disable",
parameter hssi_aibnd_tx_15_aib_red_txferclkoutn_shiften                                                                                                                          = "aib_red_txferclkoutn_shift_disable",
parameter hssi_aibnd_tx_15_aib_tx_clkdiv                                                                                                                                         = "aib_tx_clkdiv_setting1",
parameter hssi_aibnd_tx_15_aib_tx_dcc_byp                                                                                                                                        = "aib_tx_dcc_byp_disable",
parameter hssi_aibnd_tx_15_aib_tx_dcc_byp_iocsr_unused                                                                                                                           = "aib_tx_dcc_byp_disable_iocsr_unused",
parameter hssi_aibnd_tx_15_aib_tx_dcc_cont_cal                                                                                                                                   = "aib_tx_dcc_cal_cont",
parameter hssi_aibnd_tx_15_aib_tx_dcc_cont_cal_iocsr_unused                                                                                                                      = "aib_tx_dcc_cal_single_iocsr_unused",
parameter hssi_aibnd_tx_15_aib_tx_dcc_dft                                                                                                                                        = "aib_tx_dcc_dft_disable",
parameter hssi_aibnd_tx_15_aib_tx_dcc_dft_sel                                                                                                                                    = "aib_tx_dcc_dft_mode0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_dll_dft_sel                                                                                                                                = "aib_tx_dcc_dll_dft_sel_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_dll_entest                                                                                                                                 = "aib_tx_dcc_dll_test_disable",
parameter hssi_aibnd_tx_15_aib_tx_dcc_dy_ctl_static                                                                                                                              = "aib_tx_dcc_dy_ctl_static_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_dy_ctlsel                                                                                                                                  = "aib_tx_dcc_dy_ctlsel_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_en                                                                                                                                         = "aib_tx_dcc_enable",
parameter hssi_aibnd_tx_15_aib_tx_dcc_en_iocsr_unused                                                                                                                            = "aib_tx_dcc_disable_iocsr_unused",
parameter hssi_aibnd_tx_15_aib_tx_dcc_manual_dn                                                                                                                                  = "aib_tx_dcc_manual_dn0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_manual_up                                                                                                                                  = "aib_tx_dcc_manual_up0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_rst_prgmnvrt                                                                                                                               = "aib_tx_dcc_st_rst_prgmnvrt_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_st_core_dn_prgmnvrt                                                                                                                        = "aib_tx_dcc_st_core_dn_prgmnvrt_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_st_core_up_prgmnvrt                                                                                                                        = "aib_tx_dcc_st_core_up_prgmnvrt_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_st_core_updnen                                                                                                                             = "aib_tx_dcc_st_core_updnen_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_st_dftmuxsel                                                                                                                               = "aib_tx_dcc_st_dftmuxsel_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_st_dly_pst                                                                                                                                 = "aib_tx_dcc_st_dly_pst_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_st_en                                                                                                                                      = "aib_tx_dcc_st_en_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_st_hps_ctrl_en                                                                                                                             = "aib_tx_dcc_hps_ctrl_en_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_st_lockreq_muxsel                                                                                                                          = "aib_tx_dcc_st_lockreq_muxsel_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_st_new_dll                                                                                                                                 = "aib_tx_dcc_new_dll_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_st_rst                                                                                                                                     = "aib_tx_dcc_st_rst_setting0",
parameter hssi_aibnd_tx_15_aib_tx_dcc_test_clk_pll_en_n                                                                                                                          = "aib_tx_dcc_test_clk_pll_en_n_disable",
parameter hssi_aibnd_tx_15_aib_tx_halfcode                                                                                                                                       = "aib_tx_halfcode_enable",
parameter hssi_aibnd_tx_15_aib_tx_selflock                                                                                                                                       = "aib_tx_selflock_enable",
parameter hssi_aibnd_tx_15_dfd_dll_dcc_en                                                                                                                                        = "disable_dfd",
parameter hssi_aibnd_tx_15_dft_hssitestip_dll_dcc_en                                                                                                                             = "disable_dft",
parameter hssi_aibnd_tx_15_op_mode                                                                                                                                               = "tx_dcc_enable",
parameter hssi_aibnd_tx_15_powerdown_mode                                                                                                                                        = "true",
parameter hssi_aibnd_tx_15_powermode_ac                                                                                                                                          = "txdatapath_low_speed_pwr",
parameter hssi_aibnd_tx_15_powermode_dc                                                                                                                                          = "txdatapath_powerdown",
parameter hssi_aibnd_tx_15_powermode_freq_hz_aib_hssi_tx_transfer_clk                                                                                                            = 0,
parameter hssi_aibnd_tx_15_redundancy_en                                                                                                                                         = "disable",
parameter hssi_aibnd_tx_15_sup_mode                                                                                                                                              = "user_mode",
parameter hssi_pldadapt_tx_15_aib_clk1_sel                                                                                                                                       = "aib_clk1_pld_pcs_tx_clk_out",
parameter hssi_pldadapt_tx_15_aib_clk2_sel                                                                                                                                       = "aib_clk2_pld_pcs_tx_clk_out",
parameter hssi_pldadapt_tx_15_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                                                              = 0,
parameter hssi_pldadapt_tx_15_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz                                                                                                            = 0,
parameter hssi_pldadapt_tx_15_hdpldadapt_aib_fabric_tx_sr_clk_in_hz                                                                                                              = 0,
parameter hssi_pldadapt_tx_15_bonding_dft_en                                                                                                                                     = "dft_dis",
parameter hssi_pldadapt_tx_15_bonding_dft_val                                                                                                                                    = "dft_0",
parameter hssi_pldadapt_tx_15_chnl_bonding                                                                                                                                       = "disable",
parameter hssi_pldadapt_tx_15_comp_cnt                                                                                                                                           = 0,
parameter hssi_pldadapt_tx_15_compin_sel                                                                                                                                         = "compin_master",
parameter hssi_pldadapt_tx_15_hdpldadapt_csr_clk_hz                                                                                                                              = 0,
parameter hssi_pldadapt_tx_15_ctrl_plane_bonding                                                                                                                                 = "individual",
parameter hssi_pldadapt_tx_15_ds_bypass_pipeln                                                                                                                                   = "ds_bypass_pipeln_dis",
parameter hssi_pldadapt_tx_15_ds_last_chnl                                                                                                                                       = "ds_not_last_chnl",
parameter hssi_pldadapt_tx_15_ds_master                                                                                                                                          = "ds_master_en",
parameter hssi_pldadapt_tx_15_duplex_mode                                                                                                                                        = "disable",
parameter hssi_pldadapt_tx_15_dv_bond                                                                                                                                            = "dv_bond_dis",
parameter hssi_pldadapt_tx_15_dv_gen                                                                                                                                             = "dv_gen_dis",
parameter hssi_pldadapt_tx_15_fifo_double_write                                                                                                                                  = "fifo_double_write_dis",
parameter hssi_pldadapt_tx_15_fifo_mode                                                                                                                                          = "phase_comp",
parameter hssi_pldadapt_tx_15_fifo_rd_clk_frm_gen_scg_en                                                                                                                         = "disable",
parameter hssi_pldadapt_tx_15_fifo_rd_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_15_fifo_rd_clk_sel                                                                                                                                    = "fifo_rd_pma_aib_tx_clk",
parameter hssi_pldadapt_tx_15_fifo_stop_rd                                                                                                                                       = "n_rd_empty",
parameter hssi_pldadapt_tx_15_fifo_stop_wr                                                                                                                                       = "n_wr_full",
parameter hssi_pldadapt_tx_15_fifo_width                                                                                                                                         = "fifo_single_width",
parameter hssi_pldadapt_tx_15_fifo_wr_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_15_fpll_shared_direct_async_in_sel                                                                                                                    = "fpll_shared_direct_async_in_rowclk",
parameter hssi_pldadapt_tx_15_frmgen_burst                                                                                                                                       = "frmgen_burst_dis",
parameter hssi_pldadapt_tx_15_frmgen_bypass                                                                                                                                      = "frmgen_bypass_dis",
parameter hssi_pldadapt_tx_15_frmgen_mfrm_length                                                                                                                                 = 2048,
parameter hssi_pldadapt_tx_15_frmgen_pipeln                                                                                                                                      = "frmgen_pipeln_dis",
parameter hssi_pldadapt_tx_15_frmgen_pyld_ins                                                                                                                                    = "frmgen_pyld_ins_dis",
parameter hssi_pldadapt_tx_15_frmgen_wordslip                                                                                                                                    = "frmgen_wordslip_dis",
parameter hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit0_rst_val                                                                                                                        = "reset_to_zero_hfsrin0",
parameter hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit1_rst_val                                                                                                                        = "reset_to_zero_hfsrin1",
parameter hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit2_rst_val                                                                                                                        = "reset_to_zero_hfsrin2",
parameter hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit3_rst_val                                                                                                                        = "reset_to_zero_hfsrin3",
parameter hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit0_rst_val                                                                                                                       = "reset_to_zero_hfsrout0",
parameter hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit1_rst_val                                                                                                                       = "reset_to_zero_hfsrout1",
parameter hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit2_rst_val                                                                                                                       = "reset_to_zero_hfsrout2",
parameter hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit3_rst_val                                                                                                                       = "reset_to_zero_hfsrout3",
parameter hssi_pldadapt_tx_15_fsr_mask_tx_pll_rst_val                                                                                                                            = "reset_to_zero_maskpll",
parameter hssi_pldadapt_tx_15_fsr_pld_txelecidle_rst_val                                                                                                                         = "reset_to_zero_txelec",
parameter hssi_pldadapt_tx_15_gb_tx_idwidth                                                                                                                                      = "idwidth_66",
parameter hssi_pldadapt_tx_15_gb_tx_odwidth                                                                                                                                      = "odwidth_32",
parameter hssi_pldadapt_tx_15_hip_mode                                                                                                                                           = "disable_hip",
parameter hssi_pldadapt_tx_15_hip_osc_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_15_hrdrst_dcd_cal_done_bypass                                                                                                                         = "disable",
parameter hssi_pldadapt_tx_15_hrdrst_rst_sm_dis                                                                                                                                  = "enable_tx_rst_sm",
parameter hssi_pldadapt_tx_15_hrdrst_rx_osc_clk_scg_en                                                                                                                           = "disable",
parameter hssi_pldadapt_tx_15_hrdrst_user_ctl_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_15_indv                                                                                                                                               = "indv_en",
parameter hssi_pldadapt_tx_15_is_paired_with                                                                                                                                     = "other",
parameter hssi_pldadapt_tx_15_loopback_mode                                                                                                                                      = "disable",
parameter hssi_pldadapt_tx_15_low_latency_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_tx_15_osc_clk_scg_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_tx_15_phcomp_rd_del                                                                                                                                      = "phcomp_rd_del2",
parameter hssi_pldadapt_tx_15_pipe_mode                                                                                                                                          = "disable_pipe",
parameter hssi_pldadapt_tx_15_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_tx_15_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_tx_15_pld_clk1_delay_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_tx_15_pld_clk1_delay_sel                                                                                                                                 = "delay_path0",
parameter hssi_pldadapt_tx_15_pld_clk1_inv_en                                                                                                                                    = "disable",
parameter hssi_pldadapt_tx_15_pld_clk1_sel                                                                                                                                       = "pld_clk1_rowclk",
parameter hssi_pldadapt_tx_15_pld_clk2_sel                                                                                                                                       = "pld_clk2_rowclk",
parameter hssi_pldadapt_tx_15_hdpldadapt_pld_sclk1_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_tx_15_hdpldadapt_pld_sclk2_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk1_dcm_hz                                                                                                                      = 0,
parameter hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk1_rowclk_hz                                                                                                                   = 0,
parameter hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk2_dcm_hz                                                                                                                      = 0,
parameter hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk2_rowclk_hz                                                                                                                   = 0,
parameter hssi_pldadapt_tx_15_pma_aib_tx_clk_expected_setting                                                                                                                    = "not_used",
parameter hssi_pldadapt_tx_15_powerdown_mode                                                                                                                                     = "powerdown",
parameter hssi_pldadapt_tx_15_powermode_dc                                                                                                                                       = "powerdown",
parameter hssi_pldadapt_tx_15_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                                                          = 0,
parameter hssi_pldadapt_tx_15_powermode_freq_hz_pld_tx_clk1_dcm                                                                                                                  = 0,
parameter hssi_pldadapt_tx_15_sh_err                                                                                                                                             = "sh_err_dis",
parameter hssi_pldadapt_tx_15_hdpldadapt_speed_grade                                                                                                                             = "dash_1",
parameter hssi_pldadapt_tx_15_hdpldadapt_sr_sr_testbus_sel                                                                                                                       = "ssr_testbus",
parameter hssi_pldadapt_tx_15_stretch_num_stages                                                                                                                                 = "zero_stage",
parameter hssi_pldadapt_tx_15_sup_mode                                                                                                                                           = "user_mode",
parameter hssi_pldadapt_tx_15_tx_datapath_tb_sel                                                                                                                                 = "cp_bond",
parameter hssi_pldadapt_tx_15_tx_fastbond_rden                                                                                                                                   = "rden_ds_del_us_del",
parameter hssi_pldadapt_tx_15_tx_fastbond_wren                                                                                                                                   = "wren_ds_del_us_del",
parameter hssi_pldadapt_tx_15_tx_fifo_power_mode                                                                                                                                 = "full_width_full_depth",
parameter hssi_pldadapt_tx_15_tx_fifo_read_latency_adjust                                                                                                                        = "disable",
parameter hssi_pldadapt_tx_15_tx_fifo_write_latency_adjust                                                                                                                       = "disable",
parameter hssi_pldadapt_tx_15_tx_hip_aib_ssr_in_polling_bypass                                                                                                                   = "disable",
parameter hssi_pldadapt_tx_15_tx_osc_clock_setting                                                                                                                               = "osc_clk_div_by1",
parameter hssi_pldadapt_tx_15_tx_pld_10g_tx_bitslip_polling_bypass                                                                                                               = "disable",
parameter hssi_pldadapt_tx_15_tx_pld_8g_tx_boundary_sel_polling_bypass                                                                                                           = "disable",
parameter hssi_pldadapt_tx_15_tx_pld_pma_fpll_cnt_sel_polling_bypass                                                                                                             = "disable",
parameter hssi_pldadapt_tx_15_tx_pld_pma_fpll_num_phase_shifts_polling_bypass                                                                                                    = "disable",
parameter hssi_pldadapt_tx_15_tx_usertest_sel                                                                                                                                    = "enable",
parameter hssi_pldadapt_tx_15_txfifo_empty                                                                                                                                       = "empty_default",
parameter hssi_pldadapt_tx_15_txfifo_full                                                                                                                                        = "full_pc_sw",
parameter hssi_pldadapt_tx_15_txfifo_mode                                                                                                                                        = "txphase_comp",
parameter hssi_pldadapt_tx_15_txfifo_pempty                                                                                                                                      = 2,
parameter hssi_pldadapt_tx_15_txfifo_pfull                                                                                                                                       = 24,
parameter hssi_pldadapt_tx_15_us_bypass_pipeln                                                                                                                                   = "us_bypass_pipeln_dis",
parameter hssi_pldadapt_tx_15_us_last_chnl                                                                                                                                       = "us_not_last_chnl",
parameter hssi_pldadapt_tx_15_us_master                                                                                                                                          = "us_master_en",
parameter hssi_pldadapt_tx_15_word_align_enable                                                                                                                                  = "disable",
parameter hssi_pldadapt_tx_15_word_mark                                                                                                                                          = "wm_en",
parameter hssi_pldadapt_tx_15_reconfig_settings                                                                                                                                  = "{}",
parameter hssi_pldadapt_rx_15_aib_clk1_sel                                                                                                                                       = "aib_clk1_rx_transfer_clk",
parameter hssi_pldadapt_rx_15_aib_clk2_sel                                                                                                                                       = "aib_clk2_rx_transfer_clk",
parameter hssi_pldadapt_rx_15_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                                                              = 0,
parameter hssi_pldadapt_rx_15_hdpldadapt_aib_fabric_rx_sr_clk_in_hz                                                                                                              = 0,
parameter hssi_pldadapt_rx_15_hdpldadapt_aib_fabric_rx_transfer_clk_hz                                                                                                           = 0,
parameter hssi_pldadapt_rx_15_asn_bypass_pma_pcie_sw_done                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_15_asn_en                                                                                                                                             = "disable",
parameter hssi_pldadapt_rx_15_asn_wait_for_dll_reset_cnt                                                                                                                         = 0,
parameter hssi_pldadapt_rx_15_asn_wait_for_fifo_flush_cnt                                                                                                                        = 0,
parameter hssi_pldadapt_rx_15_asn_wait_for_pma_pcie_sw_done_cnt                                                                                                                  = 0,
parameter hssi_pldadapt_rx_15_bonding_dft_en                                                                                                                                     = "dft_dis",
parameter hssi_pldadapt_rx_15_bonding_dft_val                                                                                                                                    = "dft_0",
parameter hssi_pldadapt_rx_15_chnl_bonding                                                                                                                                       = "disable",
parameter hssi_pldadapt_rx_15_clock_del_measure_enable                                                                                                                           = "disable",
parameter hssi_pldadapt_rx_15_comp_cnt                                                                                                                                           = 0,
parameter hssi_pldadapt_rx_15_compin_sel                                                                                                                                         = "compin_master",
parameter hssi_pldadapt_rx_15_hdpldadapt_csr_clk_hz                                                                                                                              = 0,
parameter hssi_pldadapt_rx_15_ctrl_plane_bonding                                                                                                                                 = "individual",
parameter hssi_pldadapt_rx_15_ds_bypass_pipeln                                                                                                                                   = "ds_bypass_pipeln_dis",
parameter hssi_pldadapt_rx_15_ds_last_chnl                                                                                                                                       = "ds_not_last_chnl",
parameter hssi_pldadapt_rx_15_ds_master                                                                                                                                          = "ds_master_en",
parameter hssi_pldadapt_rx_15_duplex_mode                                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_15_dv_mode                                                                                                                                            = "dv_mode_dis",
parameter hssi_pldadapt_rx_15_fifo_double_read                                                                                                                                   = "fifo_double_read_dis",
parameter hssi_pldadapt_rx_15_fifo_mode                                                                                                                                          = "phase_comp",
parameter hssi_pldadapt_rx_15_fifo_rd_clk_ins_sm_scg_en                                                                                                                          = "disable",
parameter hssi_pldadapt_rx_15_fifo_rd_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_15_fifo_rd_clk_sel                                                                                                                                    = "fifo_rd_clk_rx_transfer_clk",
parameter hssi_pldadapt_rx_15_fifo_stop_rd                                                                                                                                       = "n_rd_empty",
parameter hssi_pldadapt_rx_15_fifo_stop_wr                                                                                                                                       = "n_wr_full",
parameter hssi_pldadapt_rx_15_fifo_width                                                                                                                                         = "fifo_single_width",
parameter hssi_pldadapt_rx_15_fifo_wr_clk_del_sm_scg_en                                                                                                                          = "disable",
parameter hssi_pldadapt_rx_15_fifo_wr_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_15_fifo_wr_clk_sel                                                                                                                                    = "fifo_wr_clk_rx_transfer_clk",
parameter hssi_pldadapt_rx_15_free_run_div_clk                                                                                                                                   = "out_of_reset_sync",
parameter hssi_pldadapt_rx_15_fsr_pld_10g_rx_crc32_err_rst_val                                                                                                                   = "reset_to_zero_crc32",
parameter hssi_pldadapt_rx_15_fsr_pld_8g_sigdet_out_rst_val                                                                                                                      = "reset_to_zero_sigdet",
parameter hssi_pldadapt_rx_15_fsr_pld_ltd_b_rst_val                                                                                                                              = "reset_to_zero_ltdb",
parameter hssi_pldadapt_rx_15_fsr_pld_ltr_rst_val                                                                                                                                = "reset_to_zero_ltr",
parameter hssi_pldadapt_rx_15_fsr_pld_rx_fifo_align_clr_rst_val                                                                                                                  = "reset_to_zero_alignclr",
parameter hssi_pldadapt_rx_15_gb_rx_idwidth                                                                                                                                      = "idwidth_32",
parameter hssi_pldadapt_rx_15_gb_rx_odwidth                                                                                                                                      = "odwidth_66",
parameter hssi_pldadapt_rx_15_hip_mode                                                                                                                                           = "disable_hip",
parameter hssi_pldadapt_rx_15_hrdrst_align_bypass                                                                                                                                = "disable",
parameter hssi_pldadapt_rx_15_hrdrst_dll_lock_bypass                                                                                                                             = "disable",
parameter hssi_pldadapt_rx_15_hrdrst_rst_sm_dis                                                                                                                                  = "enable_rx_rst_sm",
parameter hssi_pldadapt_rx_15_hrdrst_rx_osc_clk_scg_en                                                                                                                           = "disable",
parameter hssi_pldadapt_rx_15_hrdrst_user_ctl_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_15_indv                                                                                                                                               = "indv_en",
parameter hssi_pldadapt_rx_15_internal_clk1_sel1                                                                                                                                 = "pma_clks_or_txfiford_post_ct_mux_clk1_mux1",
parameter hssi_pldadapt_rx_15_internal_clk1_sel2                                                                                                                                 = "pma_clks_clk1_mux2",
parameter hssi_pldadapt_rx_15_internal_clk2_sel1                                                                                                                                 = "pma_clks_or_rxfifowr_post_ct_mux_clk2_mux1",
parameter hssi_pldadapt_rx_15_internal_clk2_sel2                                                                                                                                 = "pma_clks_clk2_mux2",
parameter hssi_pldadapt_rx_15_is_paired_with                                                                                                                                     = "other",
parameter hssi_pldadapt_rx_15_loopback_mode                                                                                                                                      = "disable",
parameter hssi_pldadapt_rx_15_low_latency_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_rx_15_lpbk_mode                                                                                                                                          = "disable",
parameter hssi_pldadapt_rx_15_osc_clk_scg_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_rx_15_phcomp_rd_del                                                                                                                                      = "phcomp_rd_del2",
parameter hssi_pldadapt_rx_15_pipe_enable                                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_15_pipe_mode                                                                                                                                          = "disable_pipe",
parameter hssi_pldadapt_rx_15_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_rx_15_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_rx_15_pld_clk1_delay_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_rx_15_pld_clk1_delay_sel                                                                                                                                 = "delay_path0",
parameter hssi_pldadapt_rx_15_pld_clk1_inv_en                                                                                                                                    = "disable",
parameter hssi_pldadapt_rx_15_pld_clk1_sel                                                                                                                                       = "pld_clk1_rowclk",
parameter hssi_pldadapt_rx_15_hdpldadapt_pld_rx_clk1_dcm_hz                                                                                                                      = 0,
parameter hssi_pldadapt_rx_15_hdpldadapt_pld_rx_clk1_rowclk_hz                                                                                                                   = 0,
parameter hssi_pldadapt_rx_15_hdpldadapt_pld_sclk1_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_rx_15_hdpldadapt_pld_sclk2_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_rx_15_pma_hclk_scg_en                                                                                                                                    = "disable",
parameter hssi_pldadapt_rx_15_powerdown_mode                                                                                                                                     = "powerdown",
parameter hssi_pldadapt_rx_15_powermode_dc                                                                                                                                       = "powerdown",
parameter hssi_pldadapt_rx_15_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                                                          = 0,
parameter hssi_pldadapt_rx_15_powermode_freq_hz_pld_rx_clk1_dcm                                                                                                                  = 0,
parameter hssi_pldadapt_rx_15_rx_datapath_tb_sel                                                                                                                                 = "cp_bond",
parameter hssi_pldadapt_rx_15_rx_fastbond_rden                                                                                                                                   = "rden_ds_del_us_del",
parameter hssi_pldadapt_rx_15_rx_fastbond_wren                                                                                                                                   = "wren_ds_del_us_del",
parameter hssi_pldadapt_rx_15_rx_fifo_power_mode                                                                                                                                 = "full_width_full_depth",
parameter hssi_pldadapt_rx_15_rx_fifo_read_latency_adjust                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_15_rx_fifo_write_ctrl                                                                                                                                 = "blklock_stops",
parameter hssi_pldadapt_rx_15_rx_fifo_write_latency_adjust                                                                                                                       = "disable",
parameter hssi_pldadapt_rx_15_rx_osc_clock_setting                                                                                                                               = "osc_clk_div_by1",
parameter hssi_pldadapt_rx_15_rx_pld_8g_eidleinfersel_polling_bypass                                                                                                             = "disable",
parameter hssi_pldadapt_rx_15_rx_pld_pma_eye_monitor_polling_bypass                                                                                                              = "disable",
parameter hssi_pldadapt_rx_15_rx_pld_pma_pcie_switch_polling_bypass                                                                                                              = "disable",
parameter hssi_pldadapt_rx_15_rx_pld_pma_reser_out_polling_bypass                                                                                                                = "disable",
parameter hssi_pldadapt_rx_15_rx_prbs_flags_sr_enable                                                                                                                            = "disable",
parameter hssi_pldadapt_rx_15_rx_true_b2b                                                                                                                                        = "b2b",
parameter hssi_pldadapt_rx_15_rx_usertest_sel                                                                                                                                    = "enable",
parameter hssi_pldadapt_rx_15_rxfifo_empty                                                                                                                                       = "empty_sw",
parameter hssi_pldadapt_rx_15_rxfifo_full                                                                                                                                        = "full_pc_sw",
parameter hssi_pldadapt_rx_15_rxfifo_mode                                                                                                                                        = "rxphase_comp",
parameter hssi_pldadapt_rx_15_rxfifo_pempty                                                                                                                                      = 2,
parameter hssi_pldadapt_rx_15_rxfifo_pfull                                                                                                                                       = 48,
parameter hssi_pldadapt_rx_15_rxfiford_post_ct_sel                                                                                                                               = "rxfiford_sclk_post_ct",
parameter hssi_pldadapt_rx_15_rxfifowr_post_ct_sel                                                                                                                               = "rxfifowr_sclk_post_ct",
parameter hssi_pldadapt_rx_15_sclk_sel                                                                                                                                           = "sclk1_rowclk",
parameter hssi_pldadapt_rx_15_hdpldadapt_speed_grade                                                                                                                             = "dash_1",
parameter hssi_pldadapt_rx_15_hdpldadapt_sr_sr_testbus_sel                                                                                                                       = "ssr_testbus",
parameter hssi_pldadapt_rx_15_stretch_num_stages                                                                                                                                 = "zero_stage",
parameter hssi_pldadapt_rx_15_sup_mode                                                                                                                                           = "user_mode",
parameter hssi_pldadapt_rx_15_txfiford_post_ct_sel                                                                                                                               = "txfiford_sclk_post_ct",
parameter hssi_pldadapt_rx_15_txfifowr_post_ct_sel                                                                                                                               = "txfifowr_sclk_post_ct",
parameter hssi_pldadapt_rx_15_us_bypass_pipeln                                                                                                                                   = "us_bypass_pipeln_dis",
parameter hssi_pldadapt_rx_15_us_last_chnl                                                                                                                                       = "us_not_last_chnl",
parameter hssi_pldadapt_rx_15_us_master                                                                                                                                          = "us_master_en",
parameter hssi_pldadapt_rx_15_word_align                                                                                                                                         = "wa_en",
parameter hssi_pldadapt_rx_15_word_align_enable                                                                                                                                  = "disable",
parameter hssi_pldadapt_rx_15_reconfig_settings                                                                                                                                  = "{}",
parameter hssi_avmm1_if_15_pcs_arbiter_ctrl                                                                                                                                      = "avmm1_arbiter_uc_sel",
parameter hssi_avmm1_if_15_hssiadapt_avmm_clk_dcg_en                                                                                                                             = "disable",
parameter hssi_avmm1_if_15_hssiadapt_avmm_clk_scg_en                                                                                                                             = "disable",
parameter hssi_avmm1_if_15_pldadapt_avmm_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm1_if_15_pcs_cal_done                                                                                                                                          = "avmm1_cal_done_assert",
parameter hssi_avmm1_if_15_pcs_cal_reserved                                                                                                                                      = 0,
parameter hssi_avmm1_if_15_pcs_calibration_feature_en                                                                                                                            = "avmm1_pcs_calibration_dis",
parameter hssi_avmm1_if_15_pldadapt_gate_dis                                                                                                                                     = "disable",
parameter hssi_avmm1_if_15_pcs_hip_cal_en                                                                                                                                        = "disable",
parameter hssi_avmm1_if_15_hssiadapt_nfhssi_calibratio_feature_en                                                                                                                = "disable",
parameter hssi_avmm1_if_15_pldadapt_nfhssi_calibratio_feature_en                                                                                                                 = "disable",
parameter hssi_avmm1_if_15_hssiadapt_osc_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm1_if_15_pldadapt_osc_clk_scg_en                                                                                                                               = "disable",
parameter hssi_avmm1_if_15_hssiadapt_read_blocking_enable                                                                                                                        = "enable",
parameter hssi_avmm1_if_15_pldadapt_read_blocking_enable                                                                                                                         = "enable",
parameter hssi_avmm1_if_15_hssiadapt_uc_blocking_enable                                                                                                                          = "enable",
parameter hssi_avmm1_if_15_pldadapt_uc_blocking_enable                                                                                                                           = "enable",
parameter hssi_avmm1_if_15_hssiadapt_write_resp_en                                                                                                                               = "disable",
parameter hssi_avmm1_if_15_hssiadapt_avmm_osc_clock_setting                                                                                                                      = "osc_clk_div_by1",
parameter hssi_avmm1_if_15_pldadapt_avmm_osc_clock_setting                                                                                                                       = "osc_clk_div_by1",
parameter hssi_avmm1_if_15_hssiadapt_avmm_testbus_sel                                                                                                                            = "avmm1_transfer_testbus",
parameter hssi_avmm1_if_15_pldadapt_avmm_testbus_sel                                                                                                                             = "avmm1_transfer_testbus",
parameter hssi_avmm1_if_15_func_mode                                                                                                                                             = "c3adpt_pmadir",
parameter hssi_avmm1_if_15_hssiadapt_sr_hip_mode                                                                                                                                 = "disable_hip",
parameter hssi_avmm1_if_15_hssiadapt_hip_mode                                                                                                                                    = "disable_hip",
parameter hssi_avmm1_if_15_pldadapt_hip_mode                                                                                                                                     = "disable_hip",
parameter hssi_avmm1_if_15_hssiadapt_sr_powerdown_mode                                                                                                                           = "powerup",
parameter hssi_avmm1_if_15_hssiadapt_sr_sr_free_run_div_clk                                                                                                                      = "out_of_reset_sync",
parameter hssi_avmm1_if_15_hssiadapt_sr_sr_hip_en                                                                                                                                = "disable",
parameter hssi_avmm1_if_15_hssiadapt_sr_sr_osc_clk_div_sel                                                                                                                       = "non_div",
parameter hssi_avmm1_if_15_hssiadapt_sr_sr_osc_clk_scg_en                                                                                                                        = "disable",
parameter hssi_avmm1_if_15_hssiadapt_sr_sr_parity_en                                                                                                                             = "disable",
parameter hssi_avmm1_if_15_hssiadapt_sr_sr_reserved_in_en                                                                                                                        = "enable",
parameter hssi_avmm1_if_15_hssiadapt_sr_sr_reserved_out_en                                                                                                                       = "enable",
parameter hssi_avmm1_if_15_hssiadapt_sr_sup_mode                                                                                                                                 = "user_mode",
parameter hssi_avmm1_if_15_topology                                                                                                                                              = "disabled_block",
parameter hssi_avmm1_if_15_calibration_type                                                                                                                                      = "one_time",
parameter hssi_avmm2_if_15_pcs_arbiter_ctrl                                                                                                                                      = "avmm2_arbiter_uc_sel",
parameter hssi_avmm2_if_15_hssiadapt_avmm_clk_dcg_en                                                                                                                             = "disable",
parameter hssi_avmm2_if_15_hssiadapt_avmm_clk_scg_en                                                                                                                             = "disable",
parameter hssi_avmm2_if_15_pldadapt_avmm_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm2_if_15_pcs_cal_done                                                                                                                                          = "avmm2_cal_done_assert",
parameter hssi_avmm2_if_15_pcs_cal_reserved                                                                                                                                      = 0,
parameter hssi_avmm2_if_15_pcs_calibration_feature_en                                                                                                                            = "avmm2_pcs_calibration_dis",
parameter hssi_avmm2_if_15_pldadapt_gate_dis                                                                                                                                     = "disable",
parameter hssi_avmm2_if_15_pcs_hip_cal_en                                                                                                                                        = "disable",
parameter hssi_avmm2_if_15_hssiadapt_osc_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm2_if_15_pldadapt_osc_clk_scg_en                                                                                                                               = "disable",
parameter hssi_avmm2_if_15_hssiadapt_avmm_osc_clock_setting                                                                                                                      = "osc_clk_div_by1",
parameter hssi_avmm2_if_15_pldadapt_avmm_osc_clock_setting                                                                                                                       = "osc_clk_div_by1",
parameter hssi_avmm2_if_15_hssiadapt_avmm_testbus_sel                                                                                                                            = "avmm1_transfer_testbus",
parameter hssi_avmm2_if_15_pldadapt_avmm_testbus_sel                                                                                                                             = "avmm1_transfer_testbus",
parameter hssi_avmm2_if_15_func_mode                                                                                                                                             = "c3adpt_pmadir",
parameter hssi_avmm2_if_15_hssiadapt_hip_mode                                                                                                                                    = "disable_hip",
parameter hssi_avmm2_if_15_pldadapt_hip_mode                                                                                                                                     = "disable_hip",
parameter hssi_avmm2_if_15_topology                                                                                                                                              = "disabled_block",
parameter hssi_avmm2_if_15_calibration_type                                                                                                                                      = "one_time",
parameter hssi_aibnd_rx_23_aib_ber_margining_ctrl                                                                                                                                = "aib_ber_margining_setting0",
parameter hssi_aibnd_rx_23_aib_datasel_gr0                                                                                                                                       = "aib_datasel0_setting0",
parameter hssi_aibnd_rx_23_aib_datasel_gr1                                                                                                                                       = "aib_datasel1_setting1",
parameter hssi_aibnd_rx_23_aib_datasel_gr2                                                                                                                                       = "aib_datasel2_setting1",
parameter hssi_aibnd_rx_23_aib_dllstr_align_clkdiv                                                                                                                               = "aib_dllstr_align_clkdiv_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_dly_pst                                                                                                                              = "aib_dllstr_align_dly_pst_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_dy_ctl_static                                                                                                                        = "aib_dllstr_align_dy_ctl_static_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_dy_ctlsel                                                                                                                            = "aib_dllstr_align_dy_ctlsel_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_entest                                                                                                                               = "aib_dllstr_align_test_disable",
parameter hssi_aibnd_rx_23_aib_dllstr_align_halfcode                                                                                                                             = "aib_dllstr_align_halfcode_enable",
parameter hssi_aibnd_rx_23_aib_dllstr_align_selflock                                                                                                                             = "aib_dllstr_align_selflock_enable",
parameter hssi_aibnd_rx_23_aib_dllstr_align_st_core_dn_prgmnvrt                                                                                                                  = "aib_dllstr_align_st_core_dn_prgmnvrt_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_st_core_up_prgmnvrt                                                                                                                  = "aib_dllstr_align_st_core_up_prgmnvrt_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_st_core_updnen                                                                                                                       = "aib_dllstr_align_st_core_updnen_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_st_dftmuxsel                                                                                                                         = "aib_dllstr_align_st_dftmuxsel_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_st_en                                                                                                                                = "aib_dllstr_align_st_en_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_st_hps_ctrl_en                                                                                                                       = "aib_dllstr_align_hps_ctrl_en_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_st_lockreq_muxsel                                                                                                                    = "aib_dllstr_align_st_lockreq_muxsel_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_st_new_dll                                                                                                                           = "aib_dllstr_align_new_dll_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_st_rst                                                                                                                               = "aib_dllstr_align_st_rst_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_st_rst_prgmnvrt                                                                                                                      = "aib_dllstr_align_st_rst_prgmnvrt_setting0",
parameter hssi_aibnd_rx_23_aib_dllstr_align_test_clk_pll_en_n                                                                                                                    = "aib_dllstr_align_test_clk_pll_en_n_disable",
parameter hssi_aibnd_rx_23_aib_inctrl_gr0                                                                                                                                        = "aib_inctrl0_setting0",
parameter hssi_aibnd_rx_23_aib_inctrl_gr1                                                                                                                                        = "aib_inctrl1_setting0",
parameter hssi_aibnd_rx_23_aib_inctrl_gr2                                                                                                                                        = "aib_inctrl2_setting0",
parameter hssi_aibnd_rx_23_aib_inctrl_gr3                                                                                                                                        = "aib_inctrl3_setting0",
parameter hssi_aibnd_rx_23_aib_outctrl_gr0                                                                                                                                       = "aib_outen0_setting0",
parameter hssi_aibnd_rx_23_aib_outctrl_gr1                                                                                                                                       = "aib_outen1_setting0",
parameter hssi_aibnd_rx_23_aib_outctrl_gr2                                                                                                                                       = "aib_outen2_setting0",
parameter hssi_aibnd_rx_23_aib_outndrv_r12                                                                                                                                       = "aib_ndrv12_setting1",
parameter hssi_aibnd_rx_23_aib_outndrv_r34                                                                                                                                       = "aib_ndrv34_setting1",
parameter hssi_aibnd_rx_23_aib_outndrv_r56                                                                                                                                       = "aib_ndrv56_setting1",
parameter hssi_aibnd_rx_23_aib_outndrv_r78                                                                                                                                       = "aib_ndrv78_setting1",
parameter hssi_aibnd_rx_23_aib_outpdrv_r12                                                                                                                                       = "aib_pdrv12_setting1",
parameter hssi_aibnd_rx_23_aib_outpdrv_r34                                                                                                                                       = "aib_pdrv34_setting1",
parameter hssi_aibnd_rx_23_aib_outpdrv_r56                                                                                                                                       = "aib_pdrv56_setting1",
parameter hssi_aibnd_rx_23_aib_outpdrv_r78                                                                                                                                       = "aib_pdrv78_setting1",
parameter hssi_aibnd_rx_23_aib_red_shift_en                                                                                                                                      = "aib_red_shift_disable",
parameter hssi_aibnd_rx_23_dft_hssitestip_dll_dcc_en                                                                                                                             = "disable_dft",
parameter hssi_aibnd_rx_23_op_mode                                                                                                                                               = "pwr_down",
parameter hssi_aibnd_rx_23_powerdown_mode                                                                                                                                        = "true",
parameter hssi_aibnd_rx_23_powermode_ac                                                                                                                                          = "rxdatapath_low_speed_pwr",
parameter hssi_aibnd_rx_23_powermode_dc                                                                                                                                          = "rxdatapath_powerdown",
parameter hssi_aibnd_rx_23_powermode_freq_hz_aib_hssi_rx_transfer_clk                                                                                                            = 0,
parameter hssi_aibnd_rx_23_redundancy_en                                                                                                                                         = "disable",
parameter hssi_aibnd_rx_23_sup_mode                                                                                                                                              = "user_mode",
parameter hssi_aibnd_tx_23_aib_datasel_gr0                                                                                                                                       = "aib_datasel0_setting0",
parameter hssi_aibnd_tx_23_aib_datasel_gr1                                                                                                                                       = "aib_datasel1_setting0",
parameter hssi_aibnd_tx_23_aib_datasel_gr2                                                                                                                                       = "aib_datasel2_setting1",
parameter hssi_aibnd_tx_23_aib_datasel_gr3                                                                                                                                       = "aib_datasel3_setting1",
parameter hssi_aibnd_tx_23_aib_ddrctrl_gr0                                                                                                                                       = "aib_ddr0_setting1",
parameter hssi_aibnd_tx_23_aib_hssi_tx_transfer_clk_hz                                                                                                                           = 0,
parameter hssi_aibnd_tx_23_aib_iinasyncen                                                                                                                                        = "aib_inasyncen_setting0",
parameter hssi_aibnd_tx_23_aib_iinclken                                                                                                                                          = "aib_inclken_setting0",
parameter hssi_aibnd_tx_23_aib_outctrl_gr0                                                                                                                                       = "aib_outen0_setting0",
parameter hssi_aibnd_tx_23_aib_outctrl_gr1                                                                                                                                       = "aib_outen1_setting0",
parameter hssi_aibnd_tx_23_aib_outctrl_gr2                                                                                                                                       = "aib_outen2_setting0",
parameter hssi_aibnd_tx_23_aib_outctrl_gr3                                                                                                                                       = "aib_outen3_setting0",
parameter hssi_aibnd_tx_23_aib_outndrv_r34                                                                                                                                       = "aib_ndrv34_setting1",
parameter hssi_aibnd_tx_23_aib_outndrv_r56                                                                                                                                       = "aib_ndrv56_setting1",
parameter hssi_aibnd_tx_23_aib_outpdrv_r34                                                                                                                                       = "aib_pdrv34_setting1",
parameter hssi_aibnd_tx_23_aib_outpdrv_r56                                                                                                                                       = "aib_pdrv56_setting1",
parameter hssi_aibnd_tx_23_aib_red_dirclkn_shiften                                                                                                                               = "aib_red_dirclkn_shift_disable",
parameter hssi_aibnd_tx_23_aib_red_dirclkp_shiften                                                                                                                               = "aib_red_dirclkp_shift_disable",
parameter hssi_aibnd_tx_23_aib_red_drx_shiften                                                                                                                                   = "aib_red_drx_shift_disable",
parameter hssi_aibnd_tx_23_aib_red_dtx_shiften                                                                                                                                   = "aib_red_dtx_shift_disable",
parameter hssi_aibnd_tx_23_aib_red_pout_shiften                                                                                                                                  = "aib_red_pout_shift_disable",
parameter hssi_aibnd_tx_23_aib_red_rx_shiften                                                                                                                                    = "aib_red_rx_shift_disable",
parameter hssi_aibnd_tx_23_aib_red_tx_shiften                                                                                                                                    = "aib_red_tx_shift_disable",
parameter hssi_aibnd_tx_23_aib_red_txferclkout_shiften                                                                                                                           = "aib_red_txferclkout_shift_disable",
parameter hssi_aibnd_tx_23_aib_red_txferclkoutn_shiften                                                                                                                          = "aib_red_txferclkoutn_shift_disable",
parameter hssi_aibnd_tx_23_aib_tx_clkdiv                                                                                                                                         = "aib_tx_clkdiv_setting1",
parameter hssi_aibnd_tx_23_aib_tx_dcc_byp                                                                                                                                        = "aib_tx_dcc_byp_disable",
parameter hssi_aibnd_tx_23_aib_tx_dcc_byp_iocsr_unused                                                                                                                           = "aib_tx_dcc_byp_disable_iocsr_unused",
parameter hssi_aibnd_tx_23_aib_tx_dcc_cont_cal                                                                                                                                   = "aib_tx_dcc_cal_cont",
parameter hssi_aibnd_tx_23_aib_tx_dcc_cont_cal_iocsr_unused                                                                                                                      = "aib_tx_dcc_cal_single_iocsr_unused",
parameter hssi_aibnd_tx_23_aib_tx_dcc_dft                                                                                                                                        = "aib_tx_dcc_dft_disable",
parameter hssi_aibnd_tx_23_aib_tx_dcc_dft_sel                                                                                                                                    = "aib_tx_dcc_dft_mode0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_dll_dft_sel                                                                                                                                = "aib_tx_dcc_dll_dft_sel_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_dll_entest                                                                                                                                 = "aib_tx_dcc_dll_test_disable",
parameter hssi_aibnd_tx_23_aib_tx_dcc_dy_ctl_static                                                                                                                              = "aib_tx_dcc_dy_ctl_static_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_dy_ctlsel                                                                                                                                  = "aib_tx_dcc_dy_ctlsel_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_en                                                                                                                                         = "aib_tx_dcc_enable",
parameter hssi_aibnd_tx_23_aib_tx_dcc_en_iocsr_unused                                                                                                                            = "aib_tx_dcc_disable_iocsr_unused",
parameter hssi_aibnd_tx_23_aib_tx_dcc_manual_dn                                                                                                                                  = "aib_tx_dcc_manual_dn0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_manual_up                                                                                                                                  = "aib_tx_dcc_manual_up0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_rst_prgmnvrt                                                                                                                               = "aib_tx_dcc_st_rst_prgmnvrt_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_st_core_dn_prgmnvrt                                                                                                                        = "aib_tx_dcc_st_core_dn_prgmnvrt_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_st_core_up_prgmnvrt                                                                                                                        = "aib_tx_dcc_st_core_up_prgmnvrt_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_st_core_updnen                                                                                                                             = "aib_tx_dcc_st_core_updnen_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_st_dftmuxsel                                                                                                                               = "aib_tx_dcc_st_dftmuxsel_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_st_dly_pst                                                                                                                                 = "aib_tx_dcc_st_dly_pst_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_st_en                                                                                                                                      = "aib_tx_dcc_st_en_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_st_hps_ctrl_en                                                                                                                             = "aib_tx_dcc_hps_ctrl_en_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_st_lockreq_muxsel                                                                                                                          = "aib_tx_dcc_st_lockreq_muxsel_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_st_new_dll                                                                                                                                 = "aib_tx_dcc_new_dll_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_st_rst                                                                                                                                     = "aib_tx_dcc_st_rst_setting0",
parameter hssi_aibnd_tx_23_aib_tx_dcc_test_clk_pll_en_n                                                                                                                          = "aib_tx_dcc_test_clk_pll_en_n_disable",
parameter hssi_aibnd_tx_23_aib_tx_halfcode                                                                                                                                       = "aib_tx_halfcode_enable",
parameter hssi_aibnd_tx_23_aib_tx_selflock                                                                                                                                       = "aib_tx_selflock_enable",
parameter hssi_aibnd_tx_23_dfd_dll_dcc_en                                                                                                                                        = "disable_dfd",
parameter hssi_aibnd_tx_23_dft_hssitestip_dll_dcc_en                                                                                                                             = "disable_dft",
parameter hssi_aibnd_tx_23_op_mode                                                                                                                                               = "tx_dcc_enable",
parameter hssi_aibnd_tx_23_powerdown_mode                                                                                                                                        = "true",
parameter hssi_aibnd_tx_23_powermode_ac                                                                                                                                          = "txdatapath_low_speed_pwr",
parameter hssi_aibnd_tx_23_powermode_dc                                                                                                                                          = "txdatapath_powerdown",
parameter hssi_aibnd_tx_23_powermode_freq_hz_aib_hssi_tx_transfer_clk                                                                                                            = 0,
parameter hssi_aibnd_tx_23_redundancy_en                                                                                                                                         = "disable",
parameter hssi_aibnd_tx_23_sup_mode                                                                                                                                              = "user_mode",
parameter hssi_pldadapt_tx_23_aib_clk1_sel                                                                                                                                       = "aib_clk1_pld_pcs_tx_clk_out",
parameter hssi_pldadapt_tx_23_aib_clk2_sel                                                                                                                                       = "aib_clk2_pld_pcs_tx_clk_out",
parameter hssi_pldadapt_tx_23_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                                                              = 0,
parameter hssi_pldadapt_tx_23_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz                                                                                                            = 0,
parameter hssi_pldadapt_tx_23_hdpldadapt_aib_fabric_tx_sr_clk_in_hz                                                                                                              = 0,
parameter hssi_pldadapt_tx_23_bonding_dft_en                                                                                                                                     = "dft_dis",
parameter hssi_pldadapt_tx_23_bonding_dft_val                                                                                                                                    = "dft_0",
parameter hssi_pldadapt_tx_23_chnl_bonding                                                                                                                                       = "disable",
parameter hssi_pldadapt_tx_23_comp_cnt                                                                                                                                           = 0,
parameter hssi_pldadapt_tx_23_compin_sel                                                                                                                                         = "compin_master",
parameter hssi_pldadapt_tx_23_hdpldadapt_csr_clk_hz                                                                                                                              = 0,
parameter hssi_pldadapt_tx_23_ctrl_plane_bonding                                                                                                                                 = "individual",
parameter hssi_pldadapt_tx_23_ds_bypass_pipeln                                                                                                                                   = "ds_bypass_pipeln_dis",
parameter hssi_pldadapt_tx_23_ds_last_chnl                                                                                                                                       = "ds_not_last_chnl",
parameter hssi_pldadapt_tx_23_ds_master                                                                                                                                          = "ds_master_en",
parameter hssi_pldadapt_tx_23_duplex_mode                                                                                                                                        = "disable",
parameter hssi_pldadapt_tx_23_dv_bond                                                                                                                                            = "dv_bond_dis",
parameter hssi_pldadapt_tx_23_dv_gen                                                                                                                                             = "dv_gen_dis",
parameter hssi_pldadapt_tx_23_fifo_double_write                                                                                                                                  = "fifo_double_write_dis",
parameter hssi_pldadapt_tx_23_fifo_mode                                                                                                                                          = "phase_comp",
parameter hssi_pldadapt_tx_23_fifo_rd_clk_frm_gen_scg_en                                                                                                                         = "disable",
parameter hssi_pldadapt_tx_23_fifo_rd_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_23_fifo_rd_clk_sel                                                                                                                                    = "fifo_rd_pma_aib_tx_clk",
parameter hssi_pldadapt_tx_23_fifo_stop_rd                                                                                                                                       = "n_rd_empty",
parameter hssi_pldadapt_tx_23_fifo_stop_wr                                                                                                                                       = "n_wr_full",
parameter hssi_pldadapt_tx_23_fifo_width                                                                                                                                         = "fifo_single_width",
parameter hssi_pldadapt_tx_23_fifo_wr_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_23_fpll_shared_direct_async_in_sel                                                                                                                    = "fpll_shared_direct_async_in_rowclk",
parameter hssi_pldadapt_tx_23_frmgen_burst                                                                                                                                       = "frmgen_burst_dis",
parameter hssi_pldadapt_tx_23_frmgen_bypass                                                                                                                                      = "frmgen_bypass_dis",
parameter hssi_pldadapt_tx_23_frmgen_mfrm_length                                                                                                                                 = 2048,
parameter hssi_pldadapt_tx_23_frmgen_pipeln                                                                                                                                      = "frmgen_pipeln_dis",
parameter hssi_pldadapt_tx_23_frmgen_pyld_ins                                                                                                                                    = "frmgen_pyld_ins_dis",
parameter hssi_pldadapt_tx_23_frmgen_wordslip                                                                                                                                    = "frmgen_wordslip_dis",
parameter hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit0_rst_val                                                                                                                        = "reset_to_zero_hfsrin0",
parameter hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit1_rst_val                                                                                                                        = "reset_to_zero_hfsrin1",
parameter hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit2_rst_val                                                                                                                        = "reset_to_zero_hfsrin2",
parameter hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit3_rst_val                                                                                                                        = "reset_to_zero_hfsrin3",
parameter hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit0_rst_val                                                                                                                       = "reset_to_zero_hfsrout0",
parameter hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit1_rst_val                                                                                                                       = "reset_to_zero_hfsrout1",
parameter hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit2_rst_val                                                                                                                       = "reset_to_zero_hfsrout2",
parameter hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit3_rst_val                                                                                                                       = "reset_to_zero_hfsrout3",
parameter hssi_pldadapt_tx_23_fsr_mask_tx_pll_rst_val                                                                                                                            = "reset_to_zero_maskpll",
parameter hssi_pldadapt_tx_23_fsr_pld_txelecidle_rst_val                                                                                                                         = "reset_to_zero_txelec",
parameter hssi_pldadapt_tx_23_gb_tx_idwidth                                                                                                                                      = "idwidth_66",
parameter hssi_pldadapt_tx_23_gb_tx_odwidth                                                                                                                                      = "odwidth_32",
parameter hssi_pldadapt_tx_23_hip_mode                                                                                                                                           = "disable_hip",
parameter hssi_pldadapt_tx_23_hip_osc_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_23_hrdrst_dcd_cal_done_bypass                                                                                                                         = "disable",
parameter hssi_pldadapt_tx_23_hrdrst_rst_sm_dis                                                                                                                                  = "enable_tx_rst_sm",
parameter hssi_pldadapt_tx_23_hrdrst_rx_osc_clk_scg_en                                                                                                                           = "disable",
parameter hssi_pldadapt_tx_23_hrdrst_user_ctl_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_tx_23_indv                                                                                                                                               = "indv_en",
parameter hssi_pldadapt_tx_23_is_paired_with                                                                                                                                     = "other",
parameter hssi_pldadapt_tx_23_loopback_mode                                                                                                                                      = "disable",
parameter hssi_pldadapt_tx_23_low_latency_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_tx_23_osc_clk_scg_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_tx_23_phcomp_rd_del                                                                                                                                      = "phcomp_rd_del2",
parameter hssi_pldadapt_tx_23_pipe_mode                                                                                                                                          = "disable_pipe",
parameter hssi_pldadapt_tx_23_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_tx_23_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_tx_23_pld_clk1_delay_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_tx_23_pld_clk1_delay_sel                                                                                                                                 = "delay_path0",
parameter hssi_pldadapt_tx_23_pld_clk1_inv_en                                                                                                                                    = "disable",
parameter hssi_pldadapt_tx_23_pld_clk1_sel                                                                                                                                       = "pld_clk1_rowclk",
parameter hssi_pldadapt_tx_23_pld_clk2_sel                                                                                                                                       = "pld_clk2_rowclk",
parameter hssi_pldadapt_tx_23_hdpldadapt_pld_sclk1_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_tx_23_hdpldadapt_pld_sclk2_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk1_dcm_hz                                                                                                                      = 0,
parameter hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk1_rowclk_hz                                                                                                                   = 0,
parameter hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk2_dcm_hz                                                                                                                      = 0,
parameter hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk2_rowclk_hz                                                                                                                   = 0,
parameter hssi_pldadapt_tx_23_pma_aib_tx_clk_expected_setting                                                                                                                    = "not_used",
parameter hssi_pldadapt_tx_23_powerdown_mode                                                                                                                                     = "powerdown",
parameter hssi_pldadapt_tx_23_powermode_dc                                                                                                                                       = "powerdown",
parameter hssi_pldadapt_tx_23_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                                                          = 0,
parameter hssi_pldadapt_tx_23_powermode_freq_hz_pld_tx_clk1_dcm                                                                                                                  = 0,
parameter hssi_pldadapt_tx_23_sh_err                                                                                                                                             = "sh_err_dis",
parameter hssi_pldadapt_tx_23_hdpldadapt_speed_grade                                                                                                                             = "dash_1",
parameter hssi_pldadapt_tx_23_hdpldadapt_sr_sr_testbus_sel                                                                                                                       = "ssr_testbus",
parameter hssi_pldadapt_tx_23_stretch_num_stages                                                                                                                                 = "zero_stage",
parameter hssi_pldadapt_tx_23_sup_mode                                                                                                                                           = "user_mode",
parameter hssi_pldadapt_tx_23_tx_datapath_tb_sel                                                                                                                                 = "cp_bond",
parameter hssi_pldadapt_tx_23_tx_fastbond_rden                                                                                                                                   = "rden_ds_del_us_del",
parameter hssi_pldadapt_tx_23_tx_fastbond_wren                                                                                                                                   = "wren_ds_del_us_del",
parameter hssi_pldadapt_tx_23_tx_fifo_power_mode                                                                                                                                 = "full_width_full_depth",
parameter hssi_pldadapt_tx_23_tx_fifo_read_latency_adjust                                                                                                                        = "disable",
parameter hssi_pldadapt_tx_23_tx_fifo_write_latency_adjust                                                                                                                       = "disable",
parameter hssi_pldadapt_tx_23_tx_hip_aib_ssr_in_polling_bypass                                                                                                                   = "disable",
parameter hssi_pldadapt_tx_23_tx_osc_clock_setting                                                                                                                               = "osc_clk_div_by1",
parameter hssi_pldadapt_tx_23_tx_pld_10g_tx_bitslip_polling_bypass                                                                                                               = "disable",
parameter hssi_pldadapt_tx_23_tx_pld_8g_tx_boundary_sel_polling_bypass                                                                                                           = "disable",
parameter hssi_pldadapt_tx_23_tx_pld_pma_fpll_cnt_sel_polling_bypass                                                                                                             = "disable",
parameter hssi_pldadapt_tx_23_tx_pld_pma_fpll_num_phase_shifts_polling_bypass                                                                                                    = "disable",
parameter hssi_pldadapt_tx_23_tx_usertest_sel                                                                                                                                    = "enable",
parameter hssi_pldadapt_tx_23_txfifo_empty                                                                                                                                       = "empty_default",
parameter hssi_pldadapt_tx_23_txfifo_full                                                                                                                                        = "full_pc_sw",
parameter hssi_pldadapt_tx_23_txfifo_mode                                                                                                                                        = "txphase_comp",
parameter hssi_pldadapt_tx_23_txfifo_pempty                                                                                                                                      = 2,
parameter hssi_pldadapt_tx_23_txfifo_pfull                                                                                                                                       = 24,
parameter hssi_pldadapt_tx_23_us_bypass_pipeln                                                                                                                                   = "us_bypass_pipeln_dis",
parameter hssi_pldadapt_tx_23_us_last_chnl                                                                                                                                       = "us_not_last_chnl",
parameter hssi_pldadapt_tx_23_us_master                                                                                                                                          = "us_master_en",
parameter hssi_pldadapt_tx_23_word_align_enable                                                                                                                                  = "disable",
parameter hssi_pldadapt_tx_23_word_mark                                                                                                                                          = "wm_en",
parameter hssi_pldadapt_tx_23_reconfig_settings                                                                                                                                  = "{}",
parameter hssi_pldadapt_rx_23_aib_clk1_sel                                                                                                                                       = "aib_clk1_rx_transfer_clk",
parameter hssi_pldadapt_rx_23_aib_clk2_sel                                                                                                                                       = "aib_clk2_rx_transfer_clk",
parameter hssi_pldadapt_rx_23_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                                                              = 0,
parameter hssi_pldadapt_rx_23_hdpldadapt_aib_fabric_rx_sr_clk_in_hz                                                                                                              = 0,
parameter hssi_pldadapt_rx_23_hdpldadapt_aib_fabric_rx_transfer_clk_hz                                                                                                           = 0,
parameter hssi_pldadapt_rx_23_asn_bypass_pma_pcie_sw_done                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_23_asn_en                                                                                                                                             = "disable",
parameter hssi_pldadapt_rx_23_asn_wait_for_dll_reset_cnt                                                                                                                         = 0,
parameter hssi_pldadapt_rx_23_asn_wait_for_fifo_flush_cnt                                                                                                                        = 0,
parameter hssi_pldadapt_rx_23_asn_wait_for_pma_pcie_sw_done_cnt                                                                                                                  = 0,
parameter hssi_pldadapt_rx_23_bonding_dft_en                                                                                                                                     = "dft_dis",
parameter hssi_pldadapt_rx_23_bonding_dft_val                                                                                                                                    = "dft_0",
parameter hssi_pldadapt_rx_23_chnl_bonding                                                                                                                                       = "disable",
parameter hssi_pldadapt_rx_23_clock_del_measure_enable                                                                                                                           = "disable",
parameter hssi_pldadapt_rx_23_comp_cnt                                                                                                                                           = 0,
parameter hssi_pldadapt_rx_23_compin_sel                                                                                                                                         = "compin_master",
parameter hssi_pldadapt_rx_23_hdpldadapt_csr_clk_hz                                                                                                                              = 0,
parameter hssi_pldadapt_rx_23_ctrl_plane_bonding                                                                                                                                 = "individual",
parameter hssi_pldadapt_rx_23_ds_bypass_pipeln                                                                                                                                   = "ds_bypass_pipeln_dis",
parameter hssi_pldadapt_rx_23_ds_last_chnl                                                                                                                                       = "ds_not_last_chnl",
parameter hssi_pldadapt_rx_23_ds_master                                                                                                                                          = "ds_master_en",
parameter hssi_pldadapt_rx_23_duplex_mode                                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_23_dv_mode                                                                                                                                            = "dv_mode_dis",
parameter hssi_pldadapt_rx_23_fifo_double_read                                                                                                                                   = "fifo_double_read_dis",
parameter hssi_pldadapt_rx_23_fifo_mode                                                                                                                                          = "phase_comp",
parameter hssi_pldadapt_rx_23_fifo_rd_clk_ins_sm_scg_en                                                                                                                          = "disable",
parameter hssi_pldadapt_rx_23_fifo_rd_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_23_fifo_rd_clk_sel                                                                                                                                    = "fifo_rd_clk_rx_transfer_clk",
parameter hssi_pldadapt_rx_23_fifo_stop_rd                                                                                                                                       = "n_rd_empty",
parameter hssi_pldadapt_rx_23_fifo_stop_wr                                                                                                                                       = "n_wr_full",
parameter hssi_pldadapt_rx_23_fifo_width                                                                                                                                         = "fifo_single_width",
parameter hssi_pldadapt_rx_23_fifo_wr_clk_del_sm_scg_en                                                                                                                          = "disable",
parameter hssi_pldadapt_rx_23_fifo_wr_clk_scg_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_23_fifo_wr_clk_sel                                                                                                                                    = "fifo_wr_clk_rx_transfer_clk",
parameter hssi_pldadapt_rx_23_free_run_div_clk                                                                                                                                   = "out_of_reset_sync",
parameter hssi_pldadapt_rx_23_fsr_pld_10g_rx_crc32_err_rst_val                                                                                                                   = "reset_to_zero_crc32",
parameter hssi_pldadapt_rx_23_fsr_pld_8g_sigdet_out_rst_val                                                                                                                      = "reset_to_zero_sigdet",
parameter hssi_pldadapt_rx_23_fsr_pld_ltd_b_rst_val                                                                                                                              = "reset_to_zero_ltdb",
parameter hssi_pldadapt_rx_23_fsr_pld_ltr_rst_val                                                                                                                                = "reset_to_zero_ltr",
parameter hssi_pldadapt_rx_23_fsr_pld_rx_fifo_align_clr_rst_val                                                                                                                  = "reset_to_zero_alignclr",
parameter hssi_pldadapt_rx_23_gb_rx_idwidth                                                                                                                                      = "idwidth_32",
parameter hssi_pldadapt_rx_23_gb_rx_odwidth                                                                                                                                      = "odwidth_66",
parameter hssi_pldadapt_rx_23_hip_mode                                                                                                                                           = "disable_hip",
parameter hssi_pldadapt_rx_23_hrdrst_align_bypass                                                                                                                                = "disable",
parameter hssi_pldadapt_rx_23_hrdrst_dll_lock_bypass                                                                                                                             = "disable",
parameter hssi_pldadapt_rx_23_hrdrst_rst_sm_dis                                                                                                                                  = "enable_rx_rst_sm",
parameter hssi_pldadapt_rx_23_hrdrst_rx_osc_clk_scg_en                                                                                                                           = "disable",
parameter hssi_pldadapt_rx_23_hrdrst_user_ctl_en                                                                                                                                 = "disable",
parameter hssi_pldadapt_rx_23_indv                                                                                                                                               = "indv_en",
parameter hssi_pldadapt_rx_23_internal_clk1_sel1                                                                                                                                 = "pma_clks_or_txfiford_post_ct_mux_clk1_mux1",
parameter hssi_pldadapt_rx_23_internal_clk1_sel2                                                                                                                                 = "pma_clks_clk1_mux2",
parameter hssi_pldadapt_rx_23_internal_clk2_sel1                                                                                                                                 = "pma_clks_or_rxfifowr_post_ct_mux_clk2_mux1",
parameter hssi_pldadapt_rx_23_internal_clk2_sel2                                                                                                                                 = "pma_clks_clk2_mux2",
parameter hssi_pldadapt_rx_23_is_paired_with                                                                                                                                     = "other",
parameter hssi_pldadapt_rx_23_loopback_mode                                                                                                                                      = "disable",
parameter hssi_pldadapt_rx_23_low_latency_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_rx_23_lpbk_mode                                                                                                                                          = "disable",
parameter hssi_pldadapt_rx_23_osc_clk_scg_en                                                                                                                                     = "disable",
parameter hssi_pldadapt_rx_23_phcomp_rd_del                                                                                                                                      = "phcomp_rd_del2",
parameter hssi_pldadapt_rx_23_pipe_enable                                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_23_pipe_mode                                                                                                                                          = "disable_pipe",
parameter hssi_pldadapt_rx_23_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_rx_23_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                                                                 = 0,
parameter hssi_pldadapt_rx_23_pld_clk1_delay_en                                                                                                                                  = "disable",
parameter hssi_pldadapt_rx_23_pld_clk1_delay_sel                                                                                                                                 = "delay_path0",
parameter hssi_pldadapt_rx_23_pld_clk1_inv_en                                                                                                                                    = "disable",
parameter hssi_pldadapt_rx_23_pld_clk1_sel                                                                                                                                       = "pld_clk1_rowclk",
parameter hssi_pldadapt_rx_23_hdpldadapt_pld_rx_clk1_dcm_hz                                                                                                                      = 0,
parameter hssi_pldadapt_rx_23_hdpldadapt_pld_rx_clk1_rowclk_hz                                                                                                                   = 0,
parameter hssi_pldadapt_rx_23_hdpldadapt_pld_sclk1_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_rx_23_hdpldadapt_pld_sclk2_rowclk_hz                                                                                                                     = 0,
parameter hssi_pldadapt_rx_23_pma_hclk_scg_en                                                                                                                                    = "disable",
parameter hssi_pldadapt_rx_23_powerdown_mode                                                                                                                                     = "powerdown",
parameter hssi_pldadapt_rx_23_powermode_dc                                                                                                                                       = "powerdown",
parameter hssi_pldadapt_rx_23_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                                                          = 0,
parameter hssi_pldadapt_rx_23_powermode_freq_hz_pld_rx_clk1_dcm                                                                                                                  = 0,
parameter hssi_pldadapt_rx_23_rx_datapath_tb_sel                                                                                                                                 = "cp_bond",
parameter hssi_pldadapt_rx_23_rx_fastbond_rden                                                                                                                                   = "rden_ds_del_us_del",
parameter hssi_pldadapt_rx_23_rx_fastbond_wren                                                                                                                                   = "wren_ds_del_us_del",
parameter hssi_pldadapt_rx_23_rx_fifo_power_mode                                                                                                                                 = "full_width_full_depth",
parameter hssi_pldadapt_rx_23_rx_fifo_read_latency_adjust                                                                                                                        = "disable",
parameter hssi_pldadapt_rx_23_rx_fifo_write_ctrl                                                                                                                                 = "blklock_stops",
parameter hssi_pldadapt_rx_23_rx_fifo_write_latency_adjust                                                                                                                       = "disable",
parameter hssi_pldadapt_rx_23_rx_osc_clock_setting                                                                                                                               = "osc_clk_div_by1",
parameter hssi_pldadapt_rx_23_rx_pld_8g_eidleinfersel_polling_bypass                                                                                                             = "disable",
parameter hssi_pldadapt_rx_23_rx_pld_pma_eye_monitor_polling_bypass                                                                                                              = "disable",
parameter hssi_pldadapt_rx_23_rx_pld_pma_pcie_switch_polling_bypass                                                                                                              = "disable",
parameter hssi_pldadapt_rx_23_rx_pld_pma_reser_out_polling_bypass                                                                                                                = "disable",
parameter hssi_pldadapt_rx_23_rx_prbs_flags_sr_enable                                                                                                                            = "disable",
parameter hssi_pldadapt_rx_23_rx_true_b2b                                                                                                                                        = "b2b",
parameter hssi_pldadapt_rx_23_rx_usertest_sel                                                                                                                                    = "enable",
parameter hssi_pldadapt_rx_23_rxfifo_empty                                                                                                                                       = "empty_sw",
parameter hssi_pldadapt_rx_23_rxfifo_full                                                                                                                                        = "full_pc_sw",
parameter hssi_pldadapt_rx_23_rxfifo_mode                                                                                                                                        = "rxphase_comp",
parameter hssi_pldadapt_rx_23_rxfifo_pempty                                                                                                                                      = 2,
parameter hssi_pldadapt_rx_23_rxfifo_pfull                                                                                                                                       = 48,
parameter hssi_pldadapt_rx_23_rxfiford_post_ct_sel                                                                                                                               = "rxfiford_sclk_post_ct",
parameter hssi_pldadapt_rx_23_rxfifowr_post_ct_sel                                                                                                                               = "rxfifowr_sclk_post_ct",
parameter hssi_pldadapt_rx_23_sclk_sel                                                                                                                                           = "sclk1_rowclk",
parameter hssi_pldadapt_rx_23_hdpldadapt_speed_grade                                                                                                                             = "dash_1",
parameter hssi_pldadapt_rx_23_hdpldadapt_sr_sr_testbus_sel                                                                                                                       = "ssr_testbus",
parameter hssi_pldadapt_rx_23_stretch_num_stages                                                                                                                                 = "zero_stage",
parameter hssi_pldadapt_rx_23_sup_mode                                                                                                                                           = "user_mode",
parameter hssi_pldadapt_rx_23_txfiford_post_ct_sel                                                                                                                               = "txfiford_sclk_post_ct",
parameter hssi_pldadapt_rx_23_txfifowr_post_ct_sel                                                                                                                               = "txfifowr_sclk_post_ct",
parameter hssi_pldadapt_rx_23_us_bypass_pipeln                                                                                                                                   = "us_bypass_pipeln_dis",
parameter hssi_pldadapt_rx_23_us_last_chnl                                                                                                                                       = "us_not_last_chnl",
parameter hssi_pldadapt_rx_23_us_master                                                                                                                                          = "us_master_en",
parameter hssi_pldadapt_rx_23_word_align                                                                                                                                         = "wa_en",
parameter hssi_pldadapt_rx_23_word_align_enable                                                                                                                                  = "disable",
parameter hssi_pldadapt_rx_23_reconfig_settings                                                                                                                                  = "{}",
parameter hssi_avmm1_if_23_pcs_arbiter_ctrl                                                                                                                                      = "avmm1_arbiter_uc_sel",
parameter hssi_avmm1_if_23_hssiadapt_avmm_clk_dcg_en                                                                                                                             = "disable",
parameter hssi_avmm1_if_23_hssiadapt_avmm_clk_scg_en                                                                                                                             = "disable",
parameter hssi_avmm1_if_23_pldadapt_avmm_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm1_if_23_pcs_cal_done                                                                                                                                          = "avmm1_cal_done_assert",
parameter hssi_avmm1_if_23_pcs_cal_reserved                                                                                                                                      = 0,
parameter hssi_avmm1_if_23_pcs_calibration_feature_en                                                                                                                            = "avmm1_pcs_calibration_dis",
parameter hssi_avmm1_if_23_pldadapt_gate_dis                                                                                                                                     = "disable",
parameter hssi_avmm1_if_23_pcs_hip_cal_en                                                                                                                                        = "disable",
parameter hssi_avmm1_if_23_hssiadapt_nfhssi_calibratio_feature_en                                                                                                                = "disable",
parameter hssi_avmm1_if_23_pldadapt_nfhssi_calibratio_feature_en                                                                                                                 = "disable",
parameter hssi_avmm1_if_23_hssiadapt_osc_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm1_if_23_pldadapt_osc_clk_scg_en                                                                                                                               = "disable",
parameter hssi_avmm1_if_23_hssiadapt_read_blocking_enable                                                                                                                        = "enable",
parameter hssi_avmm1_if_23_pldadapt_read_blocking_enable                                                                                                                         = "enable",
parameter hssi_avmm1_if_23_hssiadapt_uc_blocking_enable                                                                                                                          = "enable",
parameter hssi_avmm1_if_23_pldadapt_uc_blocking_enable                                                                                                                           = "enable",
parameter hssi_avmm1_if_23_hssiadapt_write_resp_en                                                                                                                               = "disable",
parameter hssi_avmm1_if_23_hssiadapt_avmm_osc_clock_setting                                                                                                                      = "osc_clk_div_by1",
parameter hssi_avmm1_if_23_pldadapt_avmm_osc_clock_setting                                                                                                                       = "osc_clk_div_by1",
parameter hssi_avmm1_if_23_hssiadapt_avmm_testbus_sel                                                                                                                            = "avmm1_transfer_testbus",
parameter hssi_avmm1_if_23_pldadapt_avmm_testbus_sel                                                                                                                             = "avmm1_transfer_testbus",
parameter hssi_avmm1_if_23_func_mode                                                                                                                                             = "c3adpt_pmadir",
parameter hssi_avmm1_if_23_hssiadapt_sr_hip_mode                                                                                                                                 = "disable_hip",
parameter hssi_avmm1_if_23_hssiadapt_hip_mode                                                                                                                                    = "disable_hip",
parameter hssi_avmm1_if_23_pldadapt_hip_mode                                                                                                                                     = "disable_hip",
parameter hssi_avmm1_if_23_hssiadapt_sr_powerdown_mode                                                                                                                           = "powerup",
parameter hssi_avmm1_if_23_hssiadapt_sr_sr_free_run_div_clk                                                                                                                      = "out_of_reset_sync",
parameter hssi_avmm1_if_23_hssiadapt_sr_sr_hip_en                                                                                                                                = "disable",
parameter hssi_avmm1_if_23_hssiadapt_sr_sr_osc_clk_div_sel                                                                                                                       = "non_div",
parameter hssi_avmm1_if_23_hssiadapt_sr_sr_osc_clk_scg_en                                                                                                                        = "disable",
parameter hssi_avmm1_if_23_hssiadapt_sr_sr_parity_en                                                                                                                             = "disable",
parameter hssi_avmm1_if_23_hssiadapt_sr_sr_reserved_in_en                                                                                                                        = "enable",
parameter hssi_avmm1_if_23_hssiadapt_sr_sr_reserved_out_en                                                                                                                       = "enable",
parameter hssi_avmm1_if_23_hssiadapt_sr_sup_mode                                                                                                                                 = "user_mode",
parameter hssi_avmm1_if_23_topology                                                                                                                                              = "disabled_block",
parameter hssi_avmm1_if_23_calibration_type                                                                                                                                      = "one_time",
parameter hssi_avmm2_if_23_pcs_arbiter_ctrl                                                                                                                                      = "avmm2_arbiter_uc_sel",
parameter hssi_avmm2_if_23_hssiadapt_avmm_clk_dcg_en                                                                                                                             = "disable",
parameter hssi_avmm2_if_23_hssiadapt_avmm_clk_scg_en                                                                                                                             = "disable",
parameter hssi_avmm2_if_23_pldadapt_avmm_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm2_if_23_pcs_cal_done                                                                                                                                          = "avmm2_cal_done_assert",
parameter hssi_avmm2_if_23_pcs_cal_reserved                                                                                                                                      = 0,
parameter hssi_avmm2_if_23_pcs_calibration_feature_en                                                                                                                            = "avmm2_pcs_calibration_dis",
parameter hssi_avmm2_if_23_pldadapt_gate_dis                                                                                                                                     = "disable",
parameter hssi_avmm2_if_23_pcs_hip_cal_en                                                                                                                                        = "disable",
parameter hssi_avmm2_if_23_hssiadapt_osc_clk_scg_en                                                                                                                              = "disable",
parameter hssi_avmm2_if_23_pldadapt_osc_clk_scg_en                                                                                                                               = "disable",
parameter hssi_avmm2_if_23_hssiadapt_avmm_osc_clock_setting                                                                                                                      = "osc_clk_div_by1",
parameter hssi_avmm2_if_23_pldadapt_avmm_osc_clock_setting                                                                                                                       = "osc_clk_div_by1",
parameter hssi_avmm2_if_23_hssiadapt_avmm_testbus_sel                                                                                                                            = "avmm1_transfer_testbus",
parameter hssi_avmm2_if_23_pldadapt_avmm_testbus_sel                                                                                                                             = "avmm1_transfer_testbus",
parameter hssi_avmm2_if_23_func_mode                                                                                                                                             = "c3adpt_pmadir",
parameter hssi_avmm2_if_23_hssiadapt_hip_mode                                                                                                                                    = "disable_hip",
parameter hssi_avmm2_if_23_pldadapt_hip_mode                                                                                                                                     = "disable_hip",
parameter hssi_avmm2_if_23_topology                                                                                                                                              = "disabled_block",
parameter hssi_avmm2_if_23_calibration_type                                                                                                                                      = "one_time",
parameter hssi_ctr_active_lane_octet0                                                                                                                                            = "octet0_lane_8on",
parameter hssi_ctr_active_lane_octet1                                                                                                                                            = "octet1_lane_8on",
parameter hssi_ctr_htol                                                                                                                                                          = "disable",
parameter hssi_ctr_independent_pcie_x8x8                                                                                                                                         = "disable",
parameter hssi_ctr_iopads_powerdown_mode                                                                                                                                         = "true",
parameter hssi_ctr_is_cvp_enable                                                                                                                                                 = "false",
parameter hssi_ctr_pcie_capable                                                                                                                                                  = "gen5_capable",
parameter hssi_ctr_pcie_p0_config                                                                                                                                                = "p0_rp",
parameter hssi_ctr_pcie_p1_config                                                                                                                                                = "p1_rp",
parameter hssi_ctr_pcie_p2_config                                                                                                                                                = "p2_rp",
parameter hssi_ctr_pcie_p3_config                                                                                                                                                = "p3_rp",
parameter hssi_ctr_pcie_pld_data_width                                                                                                                                           = "wide",
parameter hssi_ctr_pcie_virt_aspm                                                                                                                                                = "no_aspm",
parameter hssi_ctr_pipe_direct_octet0                                                                                                                                            = "octet0_eight_x1",
parameter hssi_ctr_pipe_direct_octet1                                                                                                                                            = "octet1_eight_x1",
parameter hssi_ctr_pld_txrx_clk_hz                                                                                                                                               = "pld_1000mhz",
parameter hssi_ctr_powerdown_mode                                                                                                                                                = "true",
parameter hssi_ctr_sup_mode                                                                                                                                                      = "user_mode",
parameter hssi_ctr_topology                                                                                                                                                      = "pcie_x16",
parameter hssi_ctr_u_aib_top_powerdown_mode                                                                                                                                      = "true",
parameter hssi_ctr_u_aib_top_sup_mode                                                                                                                                            = "user_mode",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                      = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                   = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                   = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                  = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                  = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                 = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                       = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                     = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                      = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                  = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp0                                                                                                  = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp1                                                                                                  = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp2                                                                                                  = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp3                                                                                                  = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_reset_n                                                                                                        = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                              = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                              = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                              = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                              = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                              = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                  = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                      = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                   = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                   = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                  = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                  = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                 = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                       = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                     = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                      = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                  = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp0                                                                                                  = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp1                                                                                                  = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp2                                                                                                  = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp3                                                                                                  = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_reset_n                                                                                                        = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                              = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                              = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                              = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                              = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                              = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                  = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                     = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                  = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                  = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                 = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                 = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                      = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                    = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                     = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                 = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                      = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                 = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                 = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp0                                                                                                 = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp1                                                                                                 = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp2                                                                                                 = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp3                                                                                                 = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_reset_n                                                                                                       = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                             = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                             = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                             = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                             = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                             = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                 = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                      = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                      = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                   = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                   = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                  = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                  = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                 = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                       = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                     = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                      = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                  = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp0                                                                                                  = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp1                                                                                                  = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp2                                                                                                  = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp3                                                                                                  = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_reset_n                                                                                                        = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                              = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                              = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                              = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                              = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                              = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                  = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                      = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                   = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                   = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                  = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                  = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                 = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                       = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                     = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                      = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                  = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp0                                                                                                  = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp1                                                                                                  = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp2                                                                                                  = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp3                                                                                                  = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_reset_n                                                                                                        = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                              = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                              = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                              = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                              = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                              = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                  = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                      = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                   = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                   = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                  = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                  = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                 = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                       = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                     = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                      = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                  = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp0                                                                                                  = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp1                                                                                                  = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp2                                                                                                  = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp3                                                                                                  = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_reset_n                                                                                                        = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                              = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                              = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                              = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                              = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                              = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                  = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                      = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                   = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                   = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                  = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                  = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                 = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                       = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                     = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                      = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                  = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp0                                                                                                  = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp1                                                                                                  = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp2                                                                                                  = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp3                                                                                                  = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_reset_n                                                                                                        = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                              = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                              = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                              = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                              = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                              = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                  = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                      = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                   = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                   = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                  = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                  = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                 = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                       = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                     = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                      = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                  = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp0                                                                                                  = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp1                                                                                                  = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp2                                                                                                  = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp3                                                                                                  = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_reset_n                                                                                                        = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                              = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                              = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                              = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                              = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                              = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                  = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                      = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                   = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                   = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                  = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                  = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                 = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                       = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                     = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                      = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                  = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp0                                                                                                  = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp1                                                                                                  = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp2                                                                                                  = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp3                                                                                                  = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_reset_n                                                                                                        = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                              = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                              = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                              = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                              = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                              = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                  = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                      = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                   = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                   = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                  = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                  = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                 = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                       = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                     = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                      = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                  = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp0                                                                                                  = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp1                                                                                                  = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp2                                                                                                  = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp3                                                                                                  = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_reset_n                                                                                                        = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                              = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                              = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                              = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                              = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                              = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                  = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                                                      = "avmm1_transfer_testbus",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                                                   = "feedthru_clk0_clk1",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                                                   = "feedthru_clk0_clk2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                                                                  = "pcs_chnl_tb",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                                                                  = "direct_tr_tb_bit0_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                                                                 = "phy_rx_word_clk",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                                                       = "sel_i_chnl_ssr",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                                                     = "direct_tr_usertest3_sel",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                                                      = "non_div",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                                                                  = "disable",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                                                       = "phcomp_rd_del2",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                                                                  = "zero_stage",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                                                                  = "cp_bond",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp0                                                                                                  = "tx_fifo_wrptr_wrdata_0to27_prbs",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp1                                                                                                  = "tx_fifo_rdptr_rddata_0to27_premap",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp2                                                                                                  = "rx_fifo_rdptr_rddata_0to27_postloopback",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp3                                                                                                  = "rx_fifo_wrpt_wrdata_0to27",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_reset_n                                                                                                        = "dfd_register_reset_asserted",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp0                                                                                              = "tx_fifo_wa_lock",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp1                                                                                              = "tx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp2                                                                                              = "rx_fifo_rd_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp3                                                                                              = "rx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger1_sel_grp0                                                                                              = "tx_fifo_wr_en",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                                                                  = "disable_dfd",
parameter hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                                                       = "disable_dft",

parameter hssi_ctr_true_independent_support_mode = "disable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_disable_phy_timer = "enable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_enable_phy_status = "enable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_octet_cfg_en = "disable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pin_perst0_is_fullrst = "disable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pin_perst1_is_fullrst = "disable",

parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_async_direct_rx_sel                                                                                                     = 254,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_byp_mode                                                                                                                = "hrc_mode",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_ctrl_0_control                                                                                                   = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_ctrl_1_control                                                                                                   = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_ctrl_2_control                                                                                                   = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_irq_msk                                                                                                          = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_pldpll_disable                                                                                                      = "enable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_second_pipepll_en                                                                                                   = "disable_2nd",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_sel_reset_assert                                                                                                    = "pll_lock_assert",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_sel_reset_deassert                                                                                                  = "pll_lock_deassert",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cold_reset_time                                                                                                         = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_core_rst_width                                                                                                          = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cpll_post_rls_quiet_time                                                                                                = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cpll_post_rst_quiet_time                                                                                                = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_adpt_0to7                                                                                                       = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_adpt_16to23                                                                                                     = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_adpt_8to15                                                                                                      = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_hrc                                                                                                             = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_pattern_cntr_data_sel                                                                                               = "user_data",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_reset_n                                                                                                             = "reset_en",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dis_chkplllock_b4_corerst                                                                                               = "disable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dis_phystatchk_b4_partialrst                                                                                            = "disable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_error_irq_msk                                                                                                           = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp0_sel                                                                                                        = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp1_sel                                                                                                        = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp2_sel                                                                                                        = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp3_sel                                                                                                        = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_lane_rls_quiet_time                                                                                                     = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_lane_stagger_disable                                                                                                    = "enable_lane_reset_staggering",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_lane_stagger_interval                                                                                                   = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_linkreq_fullrst                                                                                                         = "disable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_linkreq_partialrst                                                                                                      = "disable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_perst_hi_filt_time                                                                                                      = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_perst_lo_filt_time                                                                                                      = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_phy_lane_rst_width                                                                                                      = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_phy_post_lane_rst_quiet_time                                                                                            = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pin_perst_is_full_rst                                                                                                   = "full_reset",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pipepll_error_timeout                                                                                                   = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pldpll_error_timeout                                                                                                    = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pldpll_rsten_warm                                                                                                       = "disable",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_post_core_rst_quiet_time                                                                                                = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_sideband_clksel                                                                                                         = "sideband_div8clk",
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_warm_rst_timeout                                                                                                        = 0,
parameter hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_warm_rst_timeout_prescaler                                                                                              = 0,
parameter hssi_ctr_u_ctrl_powerdown_mode                                                                                                                                         = "true",

parameter hssi_ctr_u_ctrl_toolkit_debug_mode = "toolkit_debug_mode_disable",

parameter hssi_ctr_u_ial_top_cxl_op_mode                                                                                                                                         = "io_only",
parameter hssi_ctr_u_ial_top_r_credit_return_scheme                                                                                                                              = "rel_cnt",
parameter hssi_ctr_u_ial_top_r_cxlio_dphy_send_lidl_en_dis                                                                                                                       = "r_cxlio_dphy_send_lidl_en_dis_false",
parameter hssi_ctr_u_ial_top_r_flp_phy_rcvd_ts2_all_lanes_dis                                                                                                                    = "r_flp_phy_rcvd_ts2_all_lanes_dis_false",
parameter hssi_ctr_u_ial_top_r_s2m_drs_bypass_disrepflithdr                                                                                                                      = "r_s2m_drs_bypass_disrepflithdr_false",
parameter hssi_ctr_u_ial_top_r_wptr_delay                                                                                                                                        = "one_cycle",
parameter hssi_ctr_u_ial_top_rnr_ialup_flp_inst_flxbusptctl_driftbuf_en                                                                                                          = "flxbusptctl_driftbuf_en_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_flp_inst_hybrid_x4_width                                                                                                                  = "disable_x4",
parameter hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl2_ialinvratelnkdn                                                                                                          = "iapctl2_ialinvratelnkdn_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl2_vid                                                                                                                      = 32902,
parameter hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl_comclk                                                                                                                    = "iapctl_comclk_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl_force_ial                                                                                                                 = "iapctl_force_ial_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_flp_inst_sosctl_srisen                                                                                                                    = "sosctl_srisen_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_cxl_ldid_en                                                                                                                      = "ldid_enable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_ialpmmctl_vid                                                                                                                    = 32902,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_ialpmmctl_vmeb15                                                                                                                 = 72,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rcrbbar_en                                                                                                                       = "rcrbbar_en_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cfg_avmm_csr_k_partial_bypass_configload                                                                         = "cfg_avmm_csr_k_partial_bypass_configload_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_chemem_ctrl_k_perframe_addr_steer_opt                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_chemem_ctrl_k_perframe_cqid_steer_opt                                                                            = "chemem_ctrl_k_perframe_cqid_steer_opt_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_chemem_ctrl_k_perframe_slice_en                                                                                  = "chemem_ctrl_k_perframe_slice_en_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_clk_csr_k_clkreq_hysterisis                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_clk_csr_k_clock_control                                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_clk_csr_k_osc_clk_dis                                                                                            = "clk_csr_k_osc_clk_dis_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_2_k_compressed                                                                                          = "cvp_ctrl_2_k_compressed_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_2_k_devbrd_type                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_2_k_encryped                                                                                            = "cvp_ctrl_2_k_encryped_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_3_k_jtag_id_3                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_4_k_jtag_id_2                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_5_k_jtag_id_1                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_6_k_jtag_id_0                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_7_k_cvp_irq_en                                                                                          = "cvp_ctrl_7_k_cvp_irq_en_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_7_k_cvp_write_mask_ctl                                                                                  = "cvp_ctrl_7_k_cvp_write_mask_ctl_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_7_k_gpio_irq                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_h2d_arb_ctrl_k_h2drsp_throttle_en                                                                                = "h2d_arb_ctrl_k_h2drsp_throttle_en_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_ica_ctrl_k_ica_dbg_stepthrumode                                                                                  = "ica_ctrl_k_ica_dbg_stepthrumode_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_opcode_lock_k_opcode_lock                                                                                        = "opcode_lock_k_opcode_lock_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_aer_cntrl_reg_aer_ecrc_chk_capable                                                                           = "pf0_aer_cntrl_reg_aer_ecrc_chk_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_aer_cntrl_reg_aer_ecrc_gen_capable                                                                           = "pf0_aer_cntrl_reg_aer_ecrc_gen_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_global_inval_suppport                                                                                = "pf0_ats_reg_global_inval_suppport_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_inval_queue_dep                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_page_aglign_req                                                                                      = "pf0_ats_reg_page_aglign_req_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_ro_support                                                                                           = "pf0_ats_reg_ro_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg2_cpl_to_dis_support                                                                                = "pf0_devcapreg2_cpl_to_dis_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg2_ee_tlp_prefix_support                                                                             = "pf0_devcapreg2_ee_tlp_prefix_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg2_tph_cpl_support                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_ep_l0_acc_lat                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_ep_l1_acc_lat                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_flr_cap                                                                                            = "pf0_devcapreg_flr_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_rb_err_rptr                                                                                        = "pf0_devcapreg_rb_err_rptr_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devvendid_deviceid                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devvendid_vendorid                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_high_memory_range1_size_high                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_desired_interleave_range1                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_media_type_range1                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_active_range1                                                          = "pf0_dvsec_flex_bus_range1_size_low_memory_active_range1_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_class_range1                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_info_valid_range1                                                      = "pf0_dvsec_flex_bus_range1_size_low_memory_info_valid_range1_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_range1_size_low                                                        = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_high_memory_range2_size_high                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_desired_interleave_range2                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_media_type_range2                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_active_range2                                                          = "pf0_dvsec_flex_bus_range2_size_low_memory_active_range2_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_class_range2                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_info_valid_range2                                                      = "pf0_dvsec_flex_bus_range2_size_low_memory_info_valid_range2_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_range2_size_low                                                        = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_dvsecid                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_hdm_count                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_mem_hwinit_mode                                                                              = "pf0_dvsec_head2_cap_mem_hwinit_mode_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_viral_capable                                                                                = "pf0_dvsec_head2_cap_viral_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msi_cap_reg_extnd_msg_data_capable                                                                           = "pf0_msi_cap_reg_extnd_msg_data_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msi_cap_reg_mul_msg_cap                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msi_cap_reg_per_vector_msk_cap                                                                               = "pf0_msi_cap_reg_per_vector_msk_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_cap_reg_table_sz                                                                                        = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_pba_ptr_pba_bir                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_pba_ptr_pba_offset                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_table_ptr_table_bir                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_table_ptr_table_offset                                                                                  = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_pasid_reg_exec_permi_supp                                                                                    = "pf0_pasid_reg_exec_permi_supp_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_pasid_reg_pasid_max_width                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_pasid_reg_privil_mode_supp                                                                                   = "pf0_pasid_reg_privil_mode_supp_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ptm_cap_reg_local_clock_granularity                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ptm_cap_reg_ptm_rqstr_capable                                                                                = "pf0_ptm_cap_reg_ptm_rqstr_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_reset_entry_bypass_reset_entry_bypass_idle_check                                                             = "pf0_reset_entry_bypass_reset_entry_bypass_idle_check_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_revclasscode_class_codes                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_revclasscode_rid                                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_siov_dvsec_flags_h                                                                                           = "pf0_siov_dvsec_flags_h_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_siov_dvsec_funtion_dependency_link                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_siov_reg3_ims_support                                                                                        = "pf0_siov_reg3_ims_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_sriov_cap_vf_mig_cap                                                                                         = "pf0_sriov_cap_vf_mig_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_sriov_cap_vf_mig_int                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_subsystemid_subsystemid                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_subsystemid_subsystemvendorid                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_dev_spec_mode_supd                                                                           = "pf0_tph_req_cap_reg_dev_spec_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_etph_req_supd                                                                                = "pf0_tph_req_cap_reg_etph_req_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_int_vct_mode_supd                                                                            = "pf0_tph_req_cap_reg_int_vct_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_st_table_loc                                                                                 = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_tph_st_tab_size                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_0_vf_ats_globalinv_support_0                                                                       = "pf0_vf_atscap_0_vf_ats_globalinv_support_0_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_0_vf_ats_invqueue_depth_0                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_0_vf_ats_pagealignedreq_0                                                                          = "pf0_vf_atscap_0_vf_ats_pagealignedreq_0_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_1_vf_ats_globalinv_support_1                                                                       = "pf0_vf_atscap_1_vf_ats_globalinv_support_1_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_1_vf_ats_invqueue_depth_1                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_1_vf_ats_pagealignedreq_1                                                                          = "pf0_vf_atscap_1_vf_ats_pagealignedreq_1_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_2_vf_ats_globalinv_support_2                                                                       = "pf0_vf_atscap_2_vf_ats_globalinv_support_2_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_2_vf_ats_invqueue_depth_2                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_2_vf_ats_pagealignedreq_2                                                                          = "pf0_vf_atscap_2_vf_ats_pagealignedreq_2_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_3_vf_ats_globalinv_support_3                                                                       = "pf0_vf_atscap_3_vf_ats_globalinv_support_3_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_3_vf_ats_invqueue_depth_3                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_3_vf_ats_pagealignedreq_3                                                                          = "pf0_vf_atscap_3_vf_ats_pagealignedreq_3_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_4_vf_ats_globalinv_support_4                                                                       = "pf0_vf_atscap_4_vf_ats_globalinv_support_4_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_4_vf_ats_invqueue_depth_4                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_4_vf_ats_pagealignedreq_4                                                                          = "pf0_vf_atscap_4_vf_ats_pagealignedreq_4_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_5_vf_ats_globalinv_support_5                                                                       = "pf0_vf_atscap_5_vf_ats_globalinv_support_5_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_5_vf_ats_invqueue_depth_5                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_5_vf_ats_pagealignedreq_5                                                                          = "pf0_vf_atscap_5_vf_ats_pagealignedreq_5_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_6_vf_ats_globalinv_support_6                                                                       = "pf0_vf_atscap_6_vf_ats_globalinv_support_6_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_6_vf_ats_invqueue_depth_6                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_6_vf_ats_pagealignedreq_6                                                                          = "pf0_vf_atscap_6_vf_ats_pagealignedreq_6_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_7_vf_ats_globalinv_support_7                                                                       = "pf0_vf_atscap_7_vf_ats_globalinv_support_7_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_7_vf_ats_invqueue_depth_7                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_7_vf_ats_pagealignedreq_7                                                                          = "pf0_vf_atscap_7_vf_ats_pagealignedreq_7_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_device_id_vf_device_id                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_0_vf_msix_pba_bir_0                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_0_vf_msix_pba_offset_0                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_1_vf_msix_pba_bir_1                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_1_vf_msix_pba_offset_1                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_2_vf_msix_pba_bir_2                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_2_vf_msix_pba_offset_2                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_3_vf_msix_pba_bir_3                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_3_vf_msix_pba_offset_3                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_4_vf_msix_pba_bir_4                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_4_vf_msix_pba_offset_4                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_5_vf_msix_pba_bir_5                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_5_vf_msix_pba_offset_5                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_6_vf_msix_pba_bir_6                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_6_vf_msix_pba_offset_6                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_7_vf_msix_pba_bir_7                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_7_vf_msix_pba_offset_7                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_0_vf_msix_table_bir_0                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_0_vf_msix_table_offset_0                                                                       = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_1_vf_msix_table_bir_1                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_1_vf_msix_table_offset_1                                                                       = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_2_vf_msix_table_bir_2                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_2_vf_msix_table_offset_2                                                                       = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_3_vf_msix_table_bir_3                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_3_vf_msix_table_offset_3                                                                       = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_4_vf_msix_table_bir_4                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_4_vf_msix_table_offset_4                                                                       = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_5_vf_msix_table_bir_5                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_5_vf_msix_table_offset_5                                                                       = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_6_vf_msix_table_bir_6                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_6_vf_msix_table_offset_6                                                                       = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_7_vf_msix_table_bir_7                                                                          = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_7_vf_msix_table_offset_7                                                                       = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_offset_stride_first_vf_off                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_0_vf_msix_tablesz_0                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_1_vf_msix_tablesz_1                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_2_vf_msix_tablesz_2                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_3_vf_msix_tablesz_3                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_4_vf_msix_tablesz_4                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_5_vf_msix_tablesz_5                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_6_vf_msix_tablesz_6                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_7_vf_msix_tablesz_7                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_0_vf_revision_id_0                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_0_vf_subysystem_id_0                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_1_vf_revision_id_1                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_1_vf_subysystem_id_1                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_2_vf_revision_id_2                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_2_vf_subysystem_id_2                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_3_vf_revision_id_3                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_3_vf_subysystem_id_3                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_4_vf_revision_id_4                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_4_vf_subysystem_id_4                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_5_vf_revision_id_5                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_5_vf_subysystem_id_5                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_6_vf_revision_id_6                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_6_vf_subysystem_id_6                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_7_vf_revision_id_7                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_7_vf_subysystem_id_7                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_devspecific_mode_0                                                                        = "pf0_vf_tphcap_0_vf_tph_devspecific_mode_0_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_exttphreq_0                                                                               = "pf0_vf_tphcap_0_vf_tph_exttphreq_0_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_intvec_mode_0                                                                             = "pf0_vf_tphcap_0_vf_tph_intvec_mode_0_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_sttable_loc_0                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_sttable_size_0                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_devspecific_mode_1                                                                        = "pf0_vf_tphcap_1_vf_tph_devspecific_mode_1_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_exttphreq_1                                                                               = "pf0_vf_tphcap_1_vf_tph_exttphreq_1_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_intvec_mode_1                                                                             = "pf0_vf_tphcap_1_vf_tph_intvec_mode_1_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_sttable_loc_1                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_sttable_size_1                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_devspecific_mode_2                                                                        = "pf0_vf_tphcap_2_vf_tph_devspecific_mode_2_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_exttphreq_2                                                                               = "pf0_vf_tphcap_2_vf_tph_exttphreq_2_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_intvec_mode_2                                                                             = "pf0_vf_tphcap_2_vf_tph_intvec_mode_2_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_sttable_loc_2                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_sttable_size_2                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_devspecific_mode_3                                                                        = "pf0_vf_tphcap_3_vf_tph_devspecific_mode_3_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_exttphreq_3                                                                               = "pf0_vf_tphcap_3_vf_tph_exttphreq_3_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_intvec_mode_3                                                                             = "pf0_vf_tphcap_3_vf_tph_intvec_mode_3_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_sttable_loc_3                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_sttable_size_3                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_devspecific_mode_4                                                                        = "pf0_vf_tphcap_4_vf_tph_devspecific_mode_4_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_exttphreq_4                                                                               = "pf0_vf_tphcap_4_vf_tph_exttphreq_4_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_intvec_mode_4                                                                             = "pf0_vf_tphcap_4_vf_tph_intvec_mode_4_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_sttable_loc_4                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_sttable_size_4                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_devspecific_mode_5                                                                        = "pf0_vf_tphcap_5_vf_tph_devspecific_mode_5_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_exttphreq_5                                                                               = "pf0_vf_tphcap_5_vf_tph_exttphreq_5_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_intvec_mode_5                                                                             = "pf0_vf_tphcap_5_vf_tph_intvec_mode_5_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_sttable_loc_5                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_sttable_size_5                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_devspecific_mode_6                                                                        = "pf0_vf_tphcap_6_vf_tph_devspecific_mode_6_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_exttphreq_6                                                                               = "pf0_vf_tphcap_6_vf_tph_exttphreq_6_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_intvec_mode_6                                                                             = "pf0_vf_tphcap_6_vf_tph_intvec_mode_6_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_sttable_loc_6                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_sttable_size_6                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_devspecific_mode_7                                                                        = "pf0_vf_tphcap_7_vf_tph_devspecific_mode_7_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_exttphreq_7                                                                               = "pf0_vf_tphcap_7_vf_tph_exttphreq_7_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_intvec_mode_7                                                                             = "pf0_vf_tphcap_7_vf_tph_intvec_mode_7_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_sttable_loc_7                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_sttable_size_7                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_global_inval_suppport                                                                                = "pf1_ats_reg_global_inval_suppport_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_inval_queue_dep                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_page_aglign_req                                                                                      = "pf1_ats_reg_page_aglign_req_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_ro_support                                                                                           = "pf1_ats_reg_ro_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_devcapreg2_tph_cpl_support                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_devvendid_deviceid                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msi_cap_reg_extnd_msg_data_capable                                                                           = "pf1_msi_cap_reg_extnd_msg_data_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msi_cap_reg_mul_msg_cap                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msi_cap_reg_per_vector_msk_cap                                                                               = "pf1_msi_cap_reg_per_vector_msk_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_cap_reg_function_mask                                                                                   = "pf1_msix_cap_reg_function_mask_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_cap_reg_table_sz                                                                                        = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_pba_ptr_pba_bir                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_pba_ptr_pba_offset                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_table_ptr_table_bir                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_table_ptr_table_offset                                                                                  = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_revclasscode_class_codes                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_revclasscode_rid                                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_siov_dvsec_flags_h                                                                                           = "pf1_siov_dvsec_flags_h_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_siov_dvsec_funtion_dependency_link                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_siov_reg3_ims_support                                                                                        = "pf1_siov_reg3_ims_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_sriov_cap_vf_mig_cap                                                                                         = "pf1_sriov_cap_vf_mig_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_sriov_cap_vf_mig_int                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_dev_spec_mode_supd                                                                           = "pf1_tph_req_cap_reg_dev_spec_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_etph_req_supd                                                                                = "pf1_tph_req_cap_reg_etph_req_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_int_vct_mode_supd                                                                            = "pf1_tph_req_cap_reg_int_vct_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_st_table_loc                                                                                 = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_tph_st_tab_size                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_vf_device_id_vf_device_id                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_vf_offset_stride_first_vf_off                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_global_inval_suppport                                                                                = "pf2_ats_reg_global_inval_suppport_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_inval_queue_dep                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_page_aglign_req                                                                                      = "pf2_ats_reg_page_aglign_req_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_ro_support                                                                                           = "pf2_ats_reg_ro_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_devcapreg2_tph_cpl_support                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_devvendid_deviceid                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msi_cap_reg_extnd_msg_data_capable                                                                           = "pf2_msi_cap_reg_extnd_msg_data_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msi_cap_reg_mul_msg_cap                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msi_cap_reg_per_vector_msk_cap                                                                               = "pf2_msi_cap_reg_per_vector_msk_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_cap_reg_function_mask                                                                                   = "pf2_msix_cap_reg_function_mask_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_cap_reg_table_sz                                                                                        = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_pba_ptr_pba_bir                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_pba_ptr_pba_offset                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_table_ptr_table_bir                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_table_ptr_table_offset                                                                                  = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_revclasscode_class_codes                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_revclasscode_rid                                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_siov_dvsec_flags_h                                                                                           = "pf2_siov_dvsec_flags_h_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_siov_dvsec_funtion_dependency_link                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_siov_reg3_ims_support                                                                                        = "pf2_siov_reg3_ims_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_sriov_cap_vf_mig_cap                                                                                         = "pf2_sriov_cap_vf_mig_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_sriov_cap_vf_mig_int                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_dev_spec_mode_supd                                                                           = "pf2_tph_req_cap_reg_dev_spec_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_etph_req_supd                                                                                = "pf2_tph_req_cap_reg_etph_req_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_int_vct_mode_supd                                                                            = "pf2_tph_req_cap_reg_int_vct_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_st_table_loc                                                                                 = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_tph_st_tab_size                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_vf_device_id_vf_device_id                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_vf_offset_stride_first_vf_off                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_global_inval_suppport                                                                                = "pf3_ats_reg_global_inval_suppport_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_inval_queue_dep                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_page_aglign_req                                                                                      = "pf3_ats_reg_page_aglign_req_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_ro_support                                                                                           = "pf3_ats_reg_ro_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_devcapreg2_tph_cpl_support                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_devvendid_deviceid                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msi_cap_reg_extnd_msg_data_capable                                                                           = "pf3_msi_cap_reg_extnd_msg_data_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msi_cap_reg_mul_msg_cap                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msi_cap_reg_per_vector_msk_cap                                                                               = "pf3_msi_cap_reg_per_vector_msk_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_cap_reg_function_mask                                                                                   = "pf3_msix_cap_reg_function_mask_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_cap_reg_table_sz                                                                                        = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_pba_ptr_pba_bir                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_pba_ptr_pba_offset                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_table_ptr_table_bir                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_table_ptr_table_offset                                                                                  = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_revclasscode_class_codes                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_revclasscode_rid                                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_siov_dvsec_flags_h                                                                                           = "pf3_siov_dvsec_flags_h_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_siov_dvsec_funtion_dependency_link                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_siov_reg3_ims_support                                                                                        = "pf3_siov_reg3_ims_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_sriov_cap_vf_mig_cap                                                                                         = "pf3_sriov_cap_vf_mig_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_sriov_cap_vf_mig_int                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_dev_spec_mode_supd                                                                           = "pf3_tph_req_cap_reg_dev_spec_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_etph_req_supd                                                                                = "pf3_tph_req_cap_reg_etph_req_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_int_vct_mode_supd                                                                            = "pf3_tph_req_cap_reg_int_vct_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_st_table_loc                                                                                 = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_tph_st_tab_size                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_vf_device_id_vf_device_id                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_vf_offset_stride_first_vf_off                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_global_inval_suppport                                                                                = "pf4_ats_reg_global_inval_suppport_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_inval_queue_dep                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_page_aglign_req                                                                                      = "pf4_ats_reg_page_aglign_req_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_ro_support                                                                                           = "pf4_ats_reg_ro_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_devcapreg2_tph_cpl_support                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_devvendid_deviceid                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msi_cap_reg_extnd_msg_data_capable                                                                           = "pf4_msi_cap_reg_extnd_msg_data_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msi_cap_reg_mul_msg_cap                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msi_cap_reg_per_vector_msk_cap                                                                               = "pf4_msi_cap_reg_per_vector_msk_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_cap_reg_function_mask                                                                                   = "pf4_msix_cap_reg_function_mask_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_cap_reg_table_sz                                                                                        = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_pba_ptr_pba_bir                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_pba_ptr_pba_offset                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_table_ptr_table_bir                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_table_ptr_table_offset                                                                                  = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_revclasscode_class_codes                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_revclasscode_rid                                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_siov_dvsec_flags_h                                                                                           = "pf4_siov_dvsec_flags_h_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_siov_dvsec_funtion_dependency_link                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_siov_reg3_ims_support                                                                                        = "pf4_siov_reg3_ims_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_sriov_cap_vf_mig_cap                                                                                         = "pf4_sriov_cap_vf_mig_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_sriov_cap_vf_mig_int                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_dev_spec_mode_supd                                                                           = "pf4_tph_req_cap_reg_dev_spec_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_etph_req_supd                                                                                = "pf4_tph_req_cap_reg_etph_req_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_int_vct_mode_supd                                                                            = "pf4_tph_req_cap_reg_int_vct_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_st_table_loc                                                                                 = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_tph_st_tab_size                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_vf_device_id_vf_device_id                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_vf_offset_stride_first_vf_off                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_global_inval_suppport                                                                                = "pf5_ats_reg_global_inval_suppport_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_inval_queue_dep                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_page_aglign_req                                                                                      = "pf5_ats_reg_page_aglign_req_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_ro_support                                                                                           = "pf5_ats_reg_ro_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_devcapreg2_tph_cpl_support                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_devvendid_deviceid                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msi_cap_reg_extnd_msg_data_capable                                                                           = "pf5_msi_cap_reg_extnd_msg_data_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msi_cap_reg_mul_msg_cap                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msi_cap_reg_per_vector_msk_cap                                                                               = "pf5_msi_cap_reg_per_vector_msk_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_cap_reg_function_mask                                                                                   = "pf5_msix_cap_reg_function_mask_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_cap_reg_table_sz                                                                                        = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_pba_ptr_pba_bir                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_pba_ptr_pba_offset                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_table_ptr_table_bir                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_table_ptr_table_offset                                                                                  = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_revclasscode_class_codes                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_revclasscode_rid                                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_siov_dvsec_flags_h                                                                                           = "pf5_siov_dvsec_flags_h_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_siov_dvsec_funtion_dependency_link                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_siov_reg3_ims_support                                                                                        = "pf5_siov_reg3_ims_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_sriov_cap_vf_mig_cap                                                                                         = "pf5_sriov_cap_vf_mig_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_sriov_cap_vf_mig_int                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_dev_spec_mode_supd                                                                           = "pf5_tph_req_cap_reg_dev_spec_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_etph_req_supd                                                                                = "pf5_tph_req_cap_reg_etph_req_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_int_vct_mode_supd                                                                            = "pf5_tph_req_cap_reg_int_vct_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_st_table_loc                                                                                 = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_tph_st_tab_size                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_vf_device_id_vf_device_id                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_vf_offset_stride_first_vf_off                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_global_inval_suppport                                                                                = "pf6_ats_reg_global_inval_suppport_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_inval_queue_dep                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_page_aglign_req                                                                                      = "pf6_ats_reg_page_aglign_req_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_ro_support                                                                                           = "pf6_ats_reg_ro_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_devcapreg2_tph_cpl_support                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_devvendid_deviceid                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msi_cap_reg_extnd_msg_data_capable                                                                           = "pf6_msi_cap_reg_extnd_msg_data_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msi_cap_reg_mul_msg_cap                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msi_cap_reg_per_vector_msk_cap                                                                               = "pf6_msi_cap_reg_per_vector_msk_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_cap_reg_function_mask                                                                                   = "pf6_msix_cap_reg_function_mask_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_cap_reg_table_sz                                                                                        = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_pba_ptr_pba_bir                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_pba_ptr_pba_offset                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_table_ptr_table_bir                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_table_ptr_table_offset                                                                                  = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_revclasscode_class_codes                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_revclasscode_rid                                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_siov_dvsec_flags_h                                                                                           = "pf6_siov_dvsec_flags_h_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_siov_dvsec_funtion_dependency_link                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_siov_reg3_ims_support                                                                                        = "pf6_siov_reg3_ims_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_sriov_cap_vf_mig_cap                                                                                         = "pf6_sriov_cap_vf_mig_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_sriov_cap_vf_mig_int                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_dev_spec_mode_supd                                                                           = "pf6_tph_req_cap_reg_dev_spec_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_etph_req_supd                                                                                = "pf6_tph_req_cap_reg_etph_req_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_int_vct_mode_supd                                                                            = "pf6_tph_req_cap_reg_int_vct_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_st_table_loc                                                                                 = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_tph_st_tab_size                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_vf_device_id_vf_device_id                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_vf_offset_stride_first_vf_off                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_global_inval_suppport                                                                                = "pf7_ats_reg_global_inval_suppport_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_inval_queue_dep                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_page_aglign_req                                                                                      = "pf7_ats_reg_page_aglign_req_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_ro_support                                                                                           = "pf7_ats_reg_ro_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_devcapreg2_tph_cpl_support                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_devvendid_deviceid                                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msi_cap_reg_extnd_msg_data_capable                                                                           = "pf7_msi_cap_reg_extnd_msg_data_capable_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msi_cap_reg_mul_msg_cap                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msi_cap_reg_per_vector_msk_cap                                                                               = "pf7_msi_cap_reg_per_vector_msk_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_cap_reg_function_mask                                                                                   = "pf7_msix_cap_reg_function_mask_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_cap_reg_table_sz                                                                                        = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_pba_ptr_pba_bir                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_pba_ptr_pba_offset                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_table_ptr_table_bir                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_table_ptr_table_offset                                                                                  = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_revclasscode_class_codes                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_revclasscode_rid                                                                                             = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_siov_dvsec_flags_h                                                                                           = "pf7_siov_dvsec_flags_h_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_siov_dvsec_funtion_dependency_link                                                                           = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_siov_reg3_ims_support                                                                                        = "pf7_siov_reg3_ims_support_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_sriov_cap_vf_mig_cap                                                                                         = "pf7_sriov_cap_vf_mig_cap_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_sriov_cap_vf_mig_int                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_dev_spec_mode_supd                                                                           = "pf7_tph_req_cap_reg_dev_spec_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_etph_req_supd                                                                                = "pf7_tph_req_cap_reg_etph_req_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_int_vct_mode_supd                                                                            = "pf7_tph_req_cap_reg_int_vct_mode_supd_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_st_table_loc                                                                                 = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_tph_st_tab_size                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_vf_device_id_vf_device_id                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_vf_offset_stride_first_vf_off                                                                                = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pld_sbep_portid_k_pld_sbep_id                                                                                    = 128,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_powerdown_mode                                                                                                   = "true",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_r_spare_ctl2_k_r_spare_ctl2                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_reset_csr_k_pld_crs_en                                                                                           = "reset_csr_k_pld_crs_en_false",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_sup_mode                                                                                                         = "user_mode",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_addr_a2a3_data_pack                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_acs_next_ptr                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_aer_next_ptr                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_ats_next_ptr                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_cxl_next_ptr                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_ltr_next_ptr                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_msi_next_ptr                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_msix_next_ptr                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pasid_next_ptr                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pcie_next_ptr                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pm_next_ptr                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pri_next_ptr                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_ptm_next_ptr                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_siov_next_ptr                                                                                    = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_sriov_next_ptr                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_tph_next_ptr                                                                                     = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_vc_next_ptr                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cvp_bar_num                                                                                              = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cvp_mode                                                                                                 = "cvp_disabled",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_functional_mode                                                                                          = "normal",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_maxpayload_size                                                                                          = "max_payload_1024",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_num_of_pf                                                                                                = "num_1",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_acs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_aer_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_ats_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar1_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar1_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar1_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar3_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar3_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar3_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar5_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar5_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar5_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_cxl_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_expansion_rom_enable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_expansion_rom_mask                                                                                   = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_ltr_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_msi_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_msix_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_num_of_vf                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_pasid_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_prs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_ptm_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_siov_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_sriov_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_tph_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vc_cap_enable                                                                                        = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_acs_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_ats_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar1_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar1_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar1_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar3_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar3_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar3_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar5_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar5_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar5_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_msix_cap_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_tph_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_acs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_aer_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_ats_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar1_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar1_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar1_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar3_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar3_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar3_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar5_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar5_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar5_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_msi_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_msix_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_num_of_vf                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_pasid_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_prs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_siov_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_sriov_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_tph_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_acs_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_ats_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar1_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar1_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar1_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar3_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar3_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar3_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar5_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar5_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar5_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_msix_cap_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_tph_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_acs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_aer_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_ats_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar1_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar1_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar1_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar3_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar3_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar3_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar5_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar5_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar5_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_msi_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_msix_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_num_of_vf                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_pasid_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_prs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_siov_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_sriov_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_tph_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_acs_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_ats_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar1_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar1_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar1_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar3_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar3_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar3_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar5_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar5_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar5_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_msix_cap_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_tph_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_acs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_aer_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_ats_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar1_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar1_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar1_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar3_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar3_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar3_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar5_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar5_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar5_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_msi_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_msix_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_num_of_vf                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_pasid_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_prs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_siov_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_sriov_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_tph_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_acs_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_ats_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar1_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar1_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar1_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar3_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar3_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar3_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar5_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar5_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar5_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_msix_cap_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_tph_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_acs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_aer_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_ats_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar1_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar1_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar1_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar3_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar3_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar3_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar5_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar5_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar5_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_msi_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_msix_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_num_of_vf                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_pasid_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_prs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_siov_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_sriov_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_tph_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_acs_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_ats_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar1_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar1_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar1_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar3_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar3_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar3_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar5_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar5_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar5_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_msix_cap_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_tph_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_acs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_aer_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_ats_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar1_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar1_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar1_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar3_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar3_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar3_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar5_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar5_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar5_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_msi_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_msix_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_num_of_vf                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_pasid_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_prs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_siov_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_sriov_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_tph_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_acs_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_ats_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar1_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar1_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar1_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar3_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar3_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar3_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar5_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar5_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar5_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_msix_cap_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_tph_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_acs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_aer_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_ats_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar1_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar1_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar1_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar3_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar3_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar3_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar5_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar5_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar5_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_msi_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_msix_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_num_of_vf                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_pasid_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_prs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_siov_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_sriov_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_tph_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_acs_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_ats_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar1_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar1_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar1_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar3_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar3_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar3_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar5_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar5_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar5_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_msix_cap_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_tph_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_acs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_aer_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_ats_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar1_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar1_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar1_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar3_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar3_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar3_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_64b_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar5_enable                                                                                          = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar5_mask                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar5_prefetchable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_msi_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_msix_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_num_of_vf                                                                                            = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_pasid_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_prs_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_siov_cap_enable                                                                                      = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_sriov_cap_enable                                                                                     = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_tph_cap_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_acs_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_ats_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar1_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar1_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar1_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar3_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar3_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar3_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_64b_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar5_enable                                                                                       = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar5_mask                                                                                         = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar5_prefetchable                                                                                 = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_msix_cap_enable                                                                                   = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_tph_cap_enable                                                                                    = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pri_out_pagereq_capacity                                                                                 = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_ptile_header_fmt                                                                                         = "disable",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_supported_page_size                                                                                      = 0,
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_tag_support                                                                                              = "tag_5bit",
parameter hssi_ctr_u_ial_top_rnr_ialup_icm_inst_target_link_speed                                                                                                                = "gen5",
parameter hssi_ctr_u_ial_top_sup_mode                                                                                                                                            = "user_mode",
parameter hssi_ctr_u_pcie_top_powerdown_mode                                                                                                                                     = "false",
parameter hssi_ctr_u_pcie_top_ptm_enable                                                                                                                                         = "disabled",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_avmm_ctrl_k_rstrdy_resp_en_attr                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_avmm_ctrl_k_security_bypass_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p0_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p1_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p2_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p3_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_dfd_en_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_dfd_patcntr_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar0_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar1_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar2_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar3_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane0_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane1_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane2_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane3_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl3_k_trig0_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl3_k_trig1_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q0_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q1_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q2_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q3_sel_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_aib_sel_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_error_mask_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_sts_cor_en_attr                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_sts_uc_en_attr                                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_nparity_ecc_attr                                                                              = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_par_sts_uc_en_attr                                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_hw_mode_override_en                                                                                      = "disable",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf0_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf1_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf2_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf3_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf4_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf5_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf6_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf7_attr = "false",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_0_k_cii_addr_size0_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_0_k_cii_pf_en0_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_0_k_cii_start_addr0_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_1_k_cii_addr_size1_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_1_k_cii_pf_en1_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_1_k_cii_start_addr1_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_2_k_cii_addr_size2_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_2_k_cii_pf_en2_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_2_k_cii_start_addr2_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_3_k_cii_addr_size3_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_3_k_cii_pf_en3_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_3_k_cii_start_addr3_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_4_k_cii_addr_size4_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_4_k_cii_pf_en4_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_4_k_cii_start_addr4_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_5_k_cii_addr_size5_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_5_k_cii_pf_en5_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_5_k_cii_start_addr5_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_6_k_cii_addr_size6_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_6_k_cii_pf_en6_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_6_k_cii_start_addr6_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_7_k_cii_addr_size7_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_7_k_cii_pf_en7_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_7_k_cii_start_addr7_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_fixedcred_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_mcred_attr                                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_reloadcred_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_tlp_serr_dis_attr                                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_mmio_access_ctrl_grant_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_opcode_ctrl_lock_attr                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_bar0_k_cvp_bar_0_attr                                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_bar1_k_cvp_bar_1_attr                                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctl_k_cvp_bar_mode_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctl_k_cvp_bar_type_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctl_k_cvp_bar_used_attr                                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl0_k_compressed_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl0_k_encrypted_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl1_k_devbrd_type_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl1_k_vsec_next_offset_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_irq_ctrl_k_cvp_irq_en_attr                                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_irq_ctrl_k_gpio_irq_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_jtagid0_k_jtag_id_0_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_ctrl0_k_dfd_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_ctrl0_k_patcntr_en_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_0_attr                                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_1_attr                                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_2_attr                                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_3_attr                                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_trig_sel_0_attr                                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_trig_sel_1_attr                                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_0_attr                                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_1_attr                                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_2_attr                                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_3_attr                                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_pld_crs_en_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_rx_lane_flip_en_attr                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_sris_mode_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_tx_lane_flip_en_attr                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ehp_ctrl0_k_ehp_control_reg_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ehp_ctrl1_k_outstanding_crd_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ehp_ctrl1_k_tx_rd_th_attr                                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff0_k_exvf_msixpba_bir_pf0_attr                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff0_k_exvf_msixpba_offset_pf0_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff1_k_exvf_msixpba_bir_pf1_attr                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff1_k_exvf_msixpba_offset_pf1_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff2_k_exvf_msixpba_bir_pf2_attr                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff2_k_exvf_msixpba_offset_pf2_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff3_k_exvf_msixpba_bir_pf3_attr                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff3_k_exvf_msixpba_offset_pf3_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff4_k_exvf_msixpba_bir_pf4_attr                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff4_k_exvf_msixpba_offset_pf4_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff5_k_exvf_msixpba_bir_pf5_attr                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff5_k_exvf_msixpba_offset_pf5_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff6_k_exvf_msixpba_bir_pf6_attr                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff6_k_exvf_msixpba_offset_pf6_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff7_k_exvf_msixpba_bir_pf7_attr                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff7_k_exvf_msixpba_offset_pf7_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff0_k_exvf_msixtable_bir_pf0_attr                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff0_k_exvf_msixtable_offset_pf0_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff1_k_exvf_msixtable_bir_pf1_attr                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff1_k_exvf_msixtable_offset_pf1_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff2_k_exvf_msixtable_bir_pf2_attr                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff2_k_exvf_msixtable_offset_pf2_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff3_k_exvf_msixtable_bir_pf3_attr                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff3_k_exvf_msixtable_offset_pf3_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff4_k_exvf_msixtable_bir_pf4_attr                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff4_k_exvf_msixtable_offset_pf4_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff5_k_exvf_msixtable_bir_pf5_attr                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff5_k_exvf_msixtable_offset_pf5_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff6_k_exvf_msixtable_bir_pf6_attr                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff6_k_exvf_msixtable_offset_pf6_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff7_k_exvf_msixtable_bir_pf7_attr                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff7_k_exvf_msixtable_offset_pf7_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize0_k_exvf_msix_tablesize_pf0_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize0_k_exvf_msix_tablesize_pf1_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize1_k_exvf_msix_tablesize_pf2_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize1_k_exvf_msix_tablesize_pf3_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize2_k_exvf_msix_tablesize_pf4_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize2_k_exvf_msix_tablesize_pf5_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize3_k_exvf_msix_tablesize_pf6_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize3_k_exvf_msix_tablesize_pf7_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_cvp_cfg_err_en_attr                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_dbi_access_err_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr                                                                  = "false",

parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sd_eq_control1_reg_eval_interval_time = 0,

parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_multi_lane_control_off_upconfigure_support = "true",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                    = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                         = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                       = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req                                                             = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_reg_bar0_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_reg_bar0_type                                                                                     = "pf0_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar1_reg_bar1_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_reg_bar2_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_reg_bar2_type                                                                                     = "pf0_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_reg_bar3_mem_io                                                                                   = "pf0_bar3_mem",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_reg_bar3_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_reg_bar4_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_reg_bar4_type                                                                                     = "pf0_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar5_reg_bar5_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_id_nxt_ptr_reg_aux_curr                                                                            = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_id_nxt_ptr_reg_dsi                                                                                 = "pf0_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_id_nxt_ptr_reg_pme_support                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_reg_ari_acs_fun_grp_cap                                                                            = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_base_class_code                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_program_interface                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_revision_id                                                                     = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_subclass_code                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_con_status_reg_no_soft_rst                                                                             = "pf0_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                   = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap                                                               = "pf0_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id                                                            = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id                                                            = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_exp_rom_bar_mask_reg_rom_mask                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen2_ctrl_off_config_phy_tx_change                                                                     = "pf0_full_swing",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen2_ctrl_off_support_mod_ts                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable                                                           = "pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4                                                      = "gen4_pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5                                                      = "gen5_pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode                                                          = "pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4                                                     = "gen4_pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5                                                     = "gen5_pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec                                                               = 2047,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4                                                          = 927,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5                                                          = 927,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable                                                     = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4                                                = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5                                                = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_eieos_cnt                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_phase_2_3                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_phase_2_3_atg4                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_phase_2_3_atg5                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_redo                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_redo_atg4                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_redo_atg5                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_gen3_equalization_disable                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_ph01_en                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts                                                                    = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4                                                               = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5                                                               = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1_substates_off_l1sub_t_l1_2                                                                          = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1_substates_off_l1sub_t_power_off                                                                     = 2,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_comm_mode_support                                                                 = 10,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_pwr_on_scale_support                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_pwr_on_value_support                                                              = 5,

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_1_aspm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_2_aspm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support = "true",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_1_aspm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_aspm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_l1_1sub_cap_enable = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_l1_2sub_cap_enable = "disable",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_th_sca                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_th_val                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_t_common_mode                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                        = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency                                                         = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_port_num                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                 = "pf0_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                     = "pf0_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                         = "pf0_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_table_offset_reg_pci_msix_bir                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_table_offset_reg_pci_msix_table_offset                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported                                                       = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported                                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                  = "pf0_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp                                               = "pf0_not_implemented",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pipe_loopback_control_off_pipe_loopback                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset4                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset5                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset6                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset7                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset4                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset5                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset6                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset7                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset10                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset11                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset8                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset9                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset10                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset11                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset8                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset9                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset12                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset13                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset14                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset15                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset12                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset13                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset14                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset15                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset4                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset5                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset6                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset7                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset4                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset5                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset6                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset7                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset10                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset11                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset8                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset9                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset10                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset11                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset8                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset9                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset12                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset13                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset14                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset15                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset12                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset13                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset14                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset15                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_capability_reg_no_eq_needed_support                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_rsvdp_11                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_tx_precode_req                                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_tx_precoding_on                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_port_link_ctrl_off_fast_link_mode                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint4                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint5                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset4                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset5                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint4                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint5                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset4                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset5                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint6                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint7                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset6                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset7                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint6                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint7                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset6                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset7                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_rx_preset_hint8                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_rx_preset_hint9                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_tx_preset8                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_tx_preset9                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_rx_preset_hint8                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_rx_preset_hint9                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_tx_preset8                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_tx_preset9                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_rx_preset_hint10                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_rx_preset_hint11                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_tx_preset10                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_tx_preset11                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_rx_preset_hint10                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_rx_preset_hint11                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_tx_preset10                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_tx_preset11                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_rx_preset_hint12                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_rx_preset_hint13                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_tx_preset12                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_tx_preset13                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_rx_preset_hint12                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_rx_preset_hint13                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_tx_preset12                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_tx_preset13                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_rx_preset_hint14                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_rx_preset_hint15                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_tx_preset14                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_tx_preset15                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_rx_preset_hint14                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_rx_preset_hint15                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_tx_preset14                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_tx_preset15                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_type                                                                      = "pf0_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_type                                                                      = "pf0_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_type                                                                      = "pf0_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_vf_offset_position_sriov_vf_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_vf_offset_position_sriov_vf_stride                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sup_page_sizes_reg_sriov_sup_page_size                                                                 = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                         = "pf0_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_vf_device_id_reg_sriov_vf_device_id                                                                    = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_at_block                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                    = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                         = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                       = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_src_valid                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ats_capabilities_ctrl_reg_invalidate_q_depth                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ats_capabilities_ctrl_reg_page_aligned_req                                                             = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_mask_reg_pci_type0_bar0_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_mask_reg_pci_type0_bar0_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_reg_bar0_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_reg_bar0_type                                                                                     = "pf1_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar1_mask_reg_pci_type0_bar1_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar1_mask_reg_pci_type0_bar1_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar1_reg_bar1_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_mask_reg_pci_type0_bar2_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_mask_reg_pci_type0_bar2_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_reg_bar2_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_reg_bar2_type                                                                                     = "pf1_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar3_mask_reg_pci_type0_bar3_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar3_mask_reg_pci_type0_bar3_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar3_reg_bar3_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_mask_reg_pci_type0_bar4_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_mask_reg_pci_type0_bar4_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_reg_bar4_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_reg_bar4_type                                                                                     = "pf1_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar5_mask_reg_pci_type0_bar5_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar5_mask_reg_pci_type0_bar5_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar5_reg_bar5_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cap_id_nxt_ptr_reg_aux_curr                                                                            = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cap_id_nxt_ptr_reg_dsi                                                                                 = "pf1_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cap_id_nxt_ptr_reg_pme_support                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_base_class_code                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_program_interface                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_revision_id                                                                     = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_subclass_code                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_con_status_reg_no_soft_rst                                                                             = "pf1_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                   = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_capabilities_reg_pcie_cap_flr_cap                                                               = "pf1_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_control_device_status_pcie_cap_ext_tag_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_id_vendor_id_reg_pci_type0_device_id                                                            = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_id_vendor_id_reg_pci_type0_vendor_id                                                            = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_bar_mask_reg_rom_bar_enabled                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_bar_mask_reg_rom_mask                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_base_addr_reg_exp_rom_base_address                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_base_addr_reg_rom_bar_enable                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                        = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_capabilities_reg_pcie_cap_l1_exit_latency                                                         = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_capabilities_reg_pcie_cap_port_num                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                 = "pf1_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                     = "pf1_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_control_link_status_reg_pcie_cap_slot_clk_config                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                         = "pf1_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_pba_offset_reg_pci_msix_pba_bir                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_pba_offset_reg_pci_msix_pba_offset                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_table_offset_reg_pci_msix_bir                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_table_offset_reg_pci_msix_table_offset                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pasid_cap_cntrl_reg_execute_permission_supported                                                       = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pasid_cap_cntrl_reg_max_pasid_width                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pasid_cap_cntrl_reg_privileged_mode_supported                                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                  = "pf1_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                  = "pf1_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_type                                                                      = "pf1_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_type                                                                      = "pf1_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_type                                                                      = "pf1_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_vf_offset_position_sriov_vf_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_vf_offset_position_sriov_vf_stride                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sup_page_sizes_reg_sriov_sup_page_size                                                                 = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                         = "pf1_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_device_spec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_vf_device_id_reg_sriov_vf_device_id                                                                    = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_at_block                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                    = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                         = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                       = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_src_valid                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ats_capabilities_ctrl_reg_invalidate_q_depth                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ats_capabilities_ctrl_reg_page_aligned_req                                                             = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_mask_reg_pci_type0_bar0_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_mask_reg_pci_type0_bar0_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_reg_bar0_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_reg_bar0_type                                                                                     = "pf2_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar1_mask_reg_pci_type0_bar1_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar1_mask_reg_pci_type0_bar1_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar1_reg_bar1_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_mask_reg_pci_type0_bar2_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_mask_reg_pci_type0_bar2_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_reg_bar2_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_reg_bar2_type                                                                                     = "pf2_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar3_mask_reg_pci_type0_bar3_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar3_mask_reg_pci_type0_bar3_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar3_reg_bar3_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_mask_reg_pci_type0_bar4_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_mask_reg_pci_type0_bar4_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_reg_bar4_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_reg_bar4_type                                                                                     = "pf2_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar5_mask_reg_pci_type0_bar5_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar5_mask_reg_pci_type0_bar5_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar5_reg_bar5_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cap_id_nxt_ptr_reg_aux_curr                                                                            = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cap_id_nxt_ptr_reg_dsi                                                                                 = "pf2_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cap_id_nxt_ptr_reg_pme_support                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_base_class_code                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_program_interface                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_revision_id                                                                     = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_subclass_code                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_con_status_reg_no_soft_rst                                                                             = "pf2_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                   = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_capabilities_reg_pcie_cap_flr_cap                                                               = "pf2_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_control_device_status_pcie_cap_ext_tag_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_id_vendor_id_reg_pci_type0_device_id                                                            = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_id_vendor_id_reg_pci_type0_vendor_id                                                            = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_bar_mask_reg_rom_bar_enabled                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_bar_mask_reg_rom_mask                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_base_addr_reg_exp_rom_base_address                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_base_addr_reg_rom_bar_enable                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                        = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_capabilities_reg_pcie_cap_l1_exit_latency                                                         = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_capabilities_reg_pcie_cap_port_num                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                 = "pf2_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                     = "pf2_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_control_link_status_reg_pcie_cap_slot_clk_config                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                         = "pf2_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_pba_offset_reg_pci_msix_pba_bir                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_pba_offset_reg_pci_msix_pba_offset                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_table_offset_reg_pci_msix_bir                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_table_offset_reg_pci_msix_table_offset                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pasid_cap_cntrl_reg_execute_permission_supported                                                       = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pasid_cap_cntrl_reg_max_pasid_width                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pasid_cap_cntrl_reg_privileged_mode_supported                                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                  = "pf2_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                  = "pf2_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_type                                                                      = "pf2_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_type                                                                      = "pf2_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_type                                                                      = "pf2_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_vf_offset_position_sriov_vf_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_vf_offset_position_sriov_vf_stride                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sup_page_sizes_reg_sriov_sup_page_size                                                                 = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                         = "pf2_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_device_spec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_vf_device_id_reg_sriov_vf_device_id                                                                    = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_at_block                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                    = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                         = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                       = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_src_valid                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ats_capabilities_ctrl_reg_invalidate_q_depth                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ats_capabilities_ctrl_reg_page_aligned_req                                                             = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_mask_reg_pci_type0_bar0_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_mask_reg_pci_type0_bar0_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_reg_bar0_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_reg_bar0_type                                                                                     = "pf3_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar1_mask_reg_pci_type0_bar1_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar1_mask_reg_pci_type0_bar1_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar1_reg_bar1_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_mask_reg_pci_type0_bar2_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_mask_reg_pci_type0_bar2_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_reg_bar2_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_reg_bar2_type                                                                                     = "pf3_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar3_mask_reg_pci_type0_bar3_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar3_mask_reg_pci_type0_bar3_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar3_reg_bar3_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_mask_reg_pci_type0_bar4_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_mask_reg_pci_type0_bar4_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_reg_bar4_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_reg_bar4_type                                                                                     = "pf3_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar5_mask_reg_pci_type0_bar5_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar5_mask_reg_pci_type0_bar5_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar5_reg_bar5_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cap_id_nxt_ptr_reg_aux_curr                                                                            = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cap_id_nxt_ptr_reg_dsi                                                                                 = "pf3_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cap_id_nxt_ptr_reg_pme_support                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_base_class_code                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_program_interface                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_revision_id                                                                     = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_subclass_code                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_con_status_reg_no_soft_rst                                                                             = "pf3_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                   = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_capabilities_reg_pcie_cap_flr_cap                                                               = "pf3_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_control_device_status_pcie_cap_ext_tag_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_id_vendor_id_reg_pci_type0_device_id                                                            = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_id_vendor_id_reg_pci_type0_vendor_id                                                            = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_bar_mask_reg_rom_bar_enabled                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_bar_mask_reg_rom_mask                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_base_addr_reg_exp_rom_base_address                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_base_addr_reg_rom_bar_enable                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                        = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_capabilities_reg_pcie_cap_l1_exit_latency                                                         = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_capabilities_reg_pcie_cap_port_num                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                 = "pf3_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                     = "pf3_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_control_link_status_reg_pcie_cap_slot_clk_config                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                         = "pf3_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_pba_offset_reg_pci_msix_pba_bir                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_pba_offset_reg_pci_msix_pba_offset                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_table_offset_reg_pci_msix_bir                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_table_offset_reg_pci_msix_table_offset                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pasid_cap_cntrl_reg_execute_permission_supported                                                       = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pasid_cap_cntrl_reg_max_pasid_width                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pasid_cap_cntrl_reg_privileged_mode_supported                                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                  = "pf3_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                  = "pf3_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_type                                                                      = "pf3_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_type                                                                      = "pf3_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_type                                                                      = "pf3_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_vf_offset_position_sriov_vf_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_vf_offset_position_sriov_vf_stride                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sup_page_sizes_reg_sriov_sup_page_size                                                                 = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                         = "pf3_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_device_spec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_vf_device_id_reg_sriov_vf_device_id                                                                    = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_at_block                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                    = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                         = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                       = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_src_valid                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ats_capabilities_ctrl_reg_invalidate_q_depth                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ats_capabilities_ctrl_reg_page_aligned_req                                                             = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_mask_reg_pci_type0_bar0_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_mask_reg_pci_type0_bar0_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_reg_bar0_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_reg_bar0_type                                                                                     = "pf4_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar1_mask_reg_pci_type0_bar1_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar1_mask_reg_pci_type0_bar1_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar1_reg_bar1_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_mask_reg_pci_type0_bar2_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_mask_reg_pci_type0_bar2_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_reg_bar2_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_reg_bar2_type                                                                                     = "pf4_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar3_mask_reg_pci_type0_bar3_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar3_mask_reg_pci_type0_bar3_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar3_reg_bar3_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_mask_reg_pci_type0_bar4_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_mask_reg_pci_type0_bar4_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_reg_bar4_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_reg_bar4_type                                                                                     = "pf4_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar5_mask_reg_pci_type0_bar5_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar5_mask_reg_pci_type0_bar5_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar5_reg_bar5_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cap_id_nxt_ptr_reg_aux_curr                                                                            = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cap_id_nxt_ptr_reg_dsi                                                                                 = "pf4_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cap_id_nxt_ptr_reg_pme_support                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_base_class_code                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_program_interface                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_revision_id                                                                     = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_subclass_code                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_con_status_reg_no_soft_rst                                                                             = "pf4_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                   = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_capabilities_reg_pcie_cap_flr_cap                                                               = "pf4_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_control_device_status_pcie_cap_ext_tag_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_id_vendor_id_reg_pci_type0_device_id                                                            = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_id_vendor_id_reg_pci_type0_vendor_id                                                            = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_bar_mask_reg_rom_bar_enabled                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_bar_mask_reg_rom_mask                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_base_addr_reg_exp_rom_base_address                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_base_addr_reg_rom_bar_enable                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                        = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_capabilities_reg_pcie_cap_l1_exit_latency                                                         = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_capabilities_reg_pcie_cap_port_num                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                 = "pf4_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                     = "pf4_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_control_link_status_reg_pcie_cap_slot_clk_config                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                         = "pf4_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_pba_offset_reg_pci_msix_pba_bir                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_pba_offset_reg_pci_msix_pba_offset                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_table_offset_reg_pci_msix_bir                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_table_offset_reg_pci_msix_table_offset                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pasid_cap_cntrl_reg_execute_permission_supported                                                       = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pasid_cap_cntrl_reg_max_pasid_width                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pasid_cap_cntrl_reg_privileged_mode_supported                                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                  = "pf4_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                  = "pf4_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_type                                                                      = "pf4_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_type                                                                      = "pf4_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_type                                                                      = "pf4_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_vf_offset_position_sriov_vf_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_vf_offset_position_sriov_vf_stride                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sup_page_sizes_reg_sriov_sup_page_size                                                                 = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                         = "pf4_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_device_spec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_vf_device_id_reg_sriov_vf_device_id                                                                    = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_at_block                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                    = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                         = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                       = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_src_valid                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ats_capabilities_ctrl_reg_invalidate_q_depth                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ats_capabilities_ctrl_reg_page_aligned_req                                                             = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_mask_reg_pci_type0_bar0_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_mask_reg_pci_type0_bar0_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_reg_bar0_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_reg_bar0_type                                                                                     = "pf5_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar1_mask_reg_pci_type0_bar1_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar1_mask_reg_pci_type0_bar1_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar1_reg_bar1_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_mask_reg_pci_type0_bar2_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_mask_reg_pci_type0_bar2_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_reg_bar2_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_reg_bar2_type                                                                                     = "pf5_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar3_mask_reg_pci_type0_bar3_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar3_mask_reg_pci_type0_bar3_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar3_reg_bar3_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_mask_reg_pci_type0_bar4_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_mask_reg_pci_type0_bar4_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_reg_bar4_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_reg_bar4_type                                                                                     = "pf5_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar5_mask_reg_pci_type0_bar5_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar5_mask_reg_pci_type0_bar5_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar5_reg_bar5_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cap_id_nxt_ptr_reg_aux_curr                                                                            = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cap_id_nxt_ptr_reg_dsi                                                                                 = "pf5_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cap_id_nxt_ptr_reg_pme_support                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_base_class_code                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_program_interface                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_revision_id                                                                     = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_subclass_code                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_con_status_reg_no_soft_rst                                                                             = "pf5_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                   = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_capabilities_reg_pcie_cap_flr_cap                                                               = "pf5_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_control_device_status_pcie_cap_ext_tag_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_id_vendor_id_reg_pci_type0_device_id                                                            = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_id_vendor_id_reg_pci_type0_vendor_id                                                            = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_bar_mask_reg_rom_bar_enabled                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_bar_mask_reg_rom_mask                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_base_addr_reg_exp_rom_base_address                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_base_addr_reg_rom_bar_enable                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                        = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_capabilities_reg_pcie_cap_l1_exit_latency                                                         = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_capabilities_reg_pcie_cap_port_num                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                 = "pf5_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                     = "pf5_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_control_link_status_reg_pcie_cap_slot_clk_config                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                         = "pf5_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_pba_offset_reg_pci_msix_pba_bir                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_pba_offset_reg_pci_msix_pba_offset                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_table_offset_reg_pci_msix_bir                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_table_offset_reg_pci_msix_table_offset                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pasid_cap_cntrl_reg_execute_permission_supported                                                       = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pasid_cap_cntrl_reg_max_pasid_width                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pasid_cap_cntrl_reg_privileged_mode_supported                                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                  = "pf5_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                  = "pf5_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_type                                                                      = "pf5_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_type                                                                      = "pf5_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_type                                                                      = "pf5_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_vf_offset_position_sriov_vf_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_vf_offset_position_sriov_vf_stride                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sup_page_sizes_reg_sriov_sup_page_size                                                                 = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                         = "pf5_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_device_spec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_vf_device_id_reg_sriov_vf_device_id                                                                    = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_at_block                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                    = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                         = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                       = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_src_valid                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ats_capabilities_ctrl_reg_invalidate_q_depth                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ats_capabilities_ctrl_reg_page_aligned_req                                                             = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_mask_reg_pci_type0_bar0_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_mask_reg_pci_type0_bar0_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_reg_bar0_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_reg_bar0_type                                                                                     = "pf6_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar1_mask_reg_pci_type0_bar1_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar1_mask_reg_pci_type0_bar1_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar1_reg_bar1_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_mask_reg_pci_type0_bar2_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_mask_reg_pci_type0_bar2_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_reg_bar2_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_reg_bar2_type                                                                                     = "pf6_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar3_mask_reg_pci_type0_bar3_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar3_mask_reg_pci_type0_bar3_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar3_reg_bar3_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_mask_reg_pci_type0_bar4_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_mask_reg_pci_type0_bar4_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_reg_bar4_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_reg_bar4_type                                                                                     = "pf6_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar5_mask_reg_pci_type0_bar5_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar5_mask_reg_pci_type0_bar5_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar5_reg_bar5_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cap_id_nxt_ptr_reg_aux_curr                                                                            = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cap_id_nxt_ptr_reg_dsi                                                                                 = "pf6_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cap_id_nxt_ptr_reg_pme_support                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_base_class_code                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_program_interface                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_revision_id                                                                     = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_subclass_code                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_con_status_reg_no_soft_rst                                                                             = "pf6_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                   = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_capabilities_reg_pcie_cap_flr_cap                                                               = "pf6_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_control_device_status_pcie_cap_ext_tag_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_id_vendor_id_reg_pci_type0_device_id                                                            = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_id_vendor_id_reg_pci_type0_vendor_id                                                            = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_bar_mask_reg_rom_bar_enabled                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_bar_mask_reg_rom_mask                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_base_addr_reg_exp_rom_base_address                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_base_addr_reg_rom_bar_enable                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                        = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_capabilities_reg_pcie_cap_l1_exit_latency                                                         = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_capabilities_reg_pcie_cap_port_num                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                 = "pf6_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                     = "pf6_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_control_link_status_reg_pcie_cap_slot_clk_config                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                         = "pf6_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_pba_offset_reg_pci_msix_pba_bir                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_pba_offset_reg_pci_msix_pba_offset                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_table_offset_reg_pci_msix_bir                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_table_offset_reg_pci_msix_table_offset                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pasid_cap_cntrl_reg_execute_permission_supported                                                       = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pasid_cap_cntrl_reg_max_pasid_width                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pasid_cap_cntrl_reg_privileged_mode_supported                                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                  = "pf6_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                  = "pf6_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_type                                                                      = "pf6_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_type                                                                      = "pf6_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_type                                                                      = "pf6_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_vf_offset_position_sriov_vf_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_vf_offset_position_sriov_vf_stride                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sup_page_sizes_reg_sriov_sup_page_size                                                                 = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                         = "pf6_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_device_spec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_vf_device_id_reg_sriov_vf_device_id                                                                    = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_at_block                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                    = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                         = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                       = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                         = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_src_valid                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ats_capabilities_ctrl_reg_invalidate_q_depth                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ats_capabilities_ctrl_reg_page_aligned_req                                                             = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_mask_reg_pci_type0_bar0_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_mask_reg_pci_type0_bar0_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_reg_bar0_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_reg_bar0_type                                                                                     = "pf7_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar1_mask_reg_pci_type0_bar1_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar1_mask_reg_pci_type0_bar1_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar1_reg_bar1_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_mask_reg_pci_type0_bar2_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_mask_reg_pci_type0_bar2_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_reg_bar2_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_reg_bar2_type                                                                                     = "pf7_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar3_mask_reg_pci_type0_bar3_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar3_mask_reg_pci_type0_bar3_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar3_reg_bar3_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_mask_reg_pci_type0_bar4_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_mask_reg_pci_type0_bar4_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_reg_bar4_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_reg_bar4_type                                                                                     = "pf7_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar5_mask_reg_pci_type0_bar5_enabled                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar5_mask_reg_pci_type0_bar5_mask                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar5_reg_bar5_prefetch                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cap_id_nxt_ptr_reg_aux_curr                                                                            = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cap_id_nxt_ptr_reg_dsi                                                                                 = "pf7_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cap_id_nxt_ptr_reg_pme_support                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_base_class_code                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_program_interface                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_revision_id                                                                     = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_subclass_code                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_con_status_reg_no_soft_rst                                                                             = "pf7_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                   = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_capabilities_reg_pcie_cap_flr_cap                                                               = "pf7_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_control_device_status_pcie_cap_ext_tag_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_id_vendor_id_reg_pci_type0_device_id                                                            = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_id_vendor_id_reg_pci_type0_vendor_id                                                            = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_bar_mask_reg_rom_bar_enabled                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_bar_mask_reg_rom_mask                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_base_addr_reg_exp_rom_base_address                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_base_addr_reg_rom_bar_enable                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                        = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_capabilities_reg_pcie_cap_l1_exit_latency                                                         = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_capabilities_reg_pcie_cap_port_num                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                 = "pf7_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                     = "pf7_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_control_link_status_reg_pcie_cap_slot_clk_config                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                         = "pf7_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_pba_offset_reg_pci_msix_pba_bir                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_pba_offset_reg_pci_msix_pba_offset                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_table_offset_reg_pci_msix_bir                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_table_offset_reg_pci_msix_table_offset                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pasid_cap_cntrl_reg_execute_permission_supported                                                       = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pasid_cap_cntrl_reg_max_pasid_width                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pasid_cap_cntrl_reg_privileged_mode_supported                                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                  = "pf7_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                 = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                  = "pf7_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_type                                                                      = "pf7_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_type                                                                      = "pf7_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_type                                                                      = "pf7_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_vf_offset_position_sriov_vf_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_vf_offset_position_sriov_vf_stride                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sup_page_sizes_reg_sriov_sup_page_size                                                                 = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                         = "pf7_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_device_spec                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_vf_device_id_reg_sriov_vf_device_id                                                                    = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pfvf_sel_vsec_enable_attr                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_phy_rxelecidle_k_rxelecidle_disable_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_phy_rxtermination_k_rxtermination_attr                                                                     = 127,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ptm_ctrl_k_cfg_ptm_auto_update_signal_attr                                                                 = "false",

parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ptm_adj_lsb_k_cfg_ptm_local_clock_adj_lsb_attr = 0,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ptm_adj_msb_k_cfg_ptm_local_clock_adj_msb_attr = 0,

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_reset_ctrl0_k_cvp_intf_reset_ctl_attr                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_err_en_correct_err_en_attr                                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_err_en_fatal_err_en_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_err_en_nonfatal_err_en_attr                                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_bw_mgt_int_en_attr                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_link_eq_req_int_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_pme_int_en_attr                                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_hp_int_en_attr                                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_hp_pme_en_attr                                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_inta_en_attr                                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_intb_en_attr                                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_intc_en_attr                                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_intd_en_attr                                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_sriov_misc_ctrl_k_nonsriov_mode_attr                                                                       = 255,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_stagger_control_k_stag_dlycnt_attr                                                                         = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_stagger_control_k_stag_mode_attr                                                                           = 5,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id0_k_exvf_subsysid_pf0_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id0_k_exvf_subsysid_pf1_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id1_k_exvf_subsysid_pf2_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id1_k_exvf_subsysid_pf3_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id2_k_exvf_subsysid_pf4_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id2_k_exvf_subsysid_pf5_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id3_k_exvf_subsysid_pf6_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id3_k_exvf_subsysid_pf7_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf0_attr                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf1_attr                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablesize_pf0_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablesize_pf1_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf2_attr                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf3_attr                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablesize_pf2_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablesize_pf3_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf4_attr                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf5_attr                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablesize_pf4_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablesize_pf5_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf6_attr                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf7_attr                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablesize_pf6_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablesize_pf7_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tx_common_mode_k_txcommonmode_disable_attr                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_100_k_pf4_virtio_offset_cfg3_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_102_k_pf4_virtio_offset_cfg4_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_103_k_pf4_virtio_offset_cfg4_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_104_k_pf4_virtio_offset_cfg4_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_106_k_pf4_virtio_offset_cfg5_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_107_k_pf4_virtio_offset_cfg5_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_108_k_pf4_virtio_offset_cfg5_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_109_k_pf4_virtio_offset_cfg5_cfg_data_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_111_k_pf5_virtio_offset_cfg1_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_112_k_pf5_virtio_offset_cfg1_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_113_k_pf5_virtio_offset_cfg1_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_115_k_pf5_virtio_offset_cfg2_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_116_k_pf5_virtio_offset_cfg2_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_117_k_pf5_virtio_offset_cfg2_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_118_k_pf5_virtio_offset_cfg2_notify_off_multiplier_attr                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_120_k_pf5_virtio_offset_cfg3_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_121_k_pf5_virtio_offset_cfg3_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_122_k_pf5_virtio_offset_cfg3_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_124_k_pf5_virtio_offset_cfg4_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_125_k_pf5_virtio_offset_cfg4_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_126_k_pf5_virtio_offset_cfg4_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_128_k_pf5_virtio_offset_cfg5_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_129_k_pf5_virtio_offset_cfg5_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_130_k_pf5_virtio_offset_cfg5_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_131_k_pf5_virtio_offset_cfg5_cfg_data_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_133_k_pf6_virtio_offset_cfg1_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_134_k_pf6_virtio_offset_cfg1_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_135_k_pf6_virtio_offset_cfg1_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_137_k_pf6_virtio_offset_cfg2_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_138_k_pf6_virtio_offset_cfg2_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_139_k_pf6_virtio_offset_cfg2_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_140_k_pf6_virtio_offset_cfg2_notify_off_multiplier_attr                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_142_k_pf6_virtio_offset_cfg3_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_143_k_pf6_virtio_offset_cfg3_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_144_k_pf6_virtio_offset_cfg3_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_146_k_pf6_virtio_offset_cfg4_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_147_k_pf6_virtio_offset_cfg4_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_148_k_pf6_virtio_offset_cfg4_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_150_k_pf6_virtio_offset_cfg5_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_151_k_pf6_virtio_offset_cfg5_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_152_k_pf6_virtio_offset_cfg5_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_153_k_pf6_virtio_offset_cfg5_cfg_data_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_155_k_pf7_virtio_offset_cfg1_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_156_k_pf7_virtio_offset_cfg1_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_157_k_pf7_virtio_offset_cfg1_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_159_k_pf7_virtio_offset_cfg2_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_160_k_pf7_virtio_offset_cfg2_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_161_k_pf7_virtio_offset_cfg2_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_162_k_pf7_virtio_offset_cfg2_notify_off_multiplier_attr                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_164_k_pf7_virtio_offset_cfg3_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_165_k_pf7_virtio_offset_cfg3_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_166_k_pf7_virtio_offset_cfg3_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_168_k_pf7_virtio_offset_cfg4_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_169_k_pf7_virtio_offset_cfg4_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_170_k_pf7_virtio_offset_cfg4_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_172_k_pf7_virtio_offset_cfg5_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_173_k_pf7_virtio_offset_cfg5_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_174_k_pf7_virtio_offset_cfg5_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_175_k_pf7_virtio_offset_cfg5_cfg_data_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_23_k_pf1_virtio_offset_cfg1_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_24_k_pf1_virtio_offset_cfg1_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_25_k_pf1_virtio_offset_cfg1_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_27_k_pf1_virtio_offset_cfg2_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_28_k_pf1_virtio_offset_cfg2_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_29_k_pf1_virtio_offset_cfg2_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_30_k_pf1_virtio_offset_cfg2_notify_off_multiplier_attr                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_32_k_pf1_virtio_offset_cfg3_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_33_k_pf1_virtio_offset_cfg3_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_34_k_pf1_virtio_offset_cfg3_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_36_k_pf1_virtio_offset_cfg4_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_37_k_pf1_virtio_offset_cfg4_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_38_k_pf1_virtio_offset_cfg4_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_40_k_pf1_virtio_offset_cfg5_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_41_k_pf1_virtio_offset_cfg5_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_42_k_pf1_virtio_offset_cfg5_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_43_k_pf1_virtio_offset_cfg5_cfg_data_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_45_k_pf2_virtio_offset_cfg1_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_46_k_pf2_virtio_offset_cfg1_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_47_k_pf2_virtio_offset_cfg1_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_49_k_pf2_virtio_offset_cfg2_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_50_k_pf2_virtio_offset_cfg2_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_51_k_pf2_virtio_offset_cfg2_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_52_k_pf2_virtio_offset_cfg2_notify_off_multiplier_attr                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_54_k_pf2_virtio_offset_cfg3_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_55_k_pf2_virtio_offset_cfg3_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_56_k_pf2_virtio_offset_cfg3_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_58_k_pf2_virtio_offset_cfg4_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_59_k_pf2_virtio_offset_cfg4_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_60_k_pf2_virtio_offset_cfg4_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_62_k_pf2_virtio_offset_cfg5_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_63_k_pf2_virtio_offset_cfg5_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_64_k_pf2_virtio_offset_cfg5_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_65_k_pf2_virtio_offset_cfg5_cfg_data_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_67_k_pf3_virtio_offset_cfg1_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_68_k_pf3_virtio_offset_cfg1_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_69_k_pf3_virtio_offset_cfg1_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_71_k_pf3_virtio_offset_cfg2_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_72_k_pf3_virtio_offset_cfg2_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_73_k_pf3_virtio_offset_cfg2_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_74_k_pf3_virtio_offset_cfg2_notify_off_multiplier_attr                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_76_k_pf3_virtio_offset_cfg3_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_77_k_pf3_virtio_offset_cfg3_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_78_k_pf3_virtio_offset_cfg3_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_80_k_pf3_virtio_offset_cfg4_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_81_k_pf3_virtio_offset_cfg4_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_82_k_pf3_virtio_offset_cfg4_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_84_k_pf3_virtio_offset_cfg5_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_85_k_pf3_virtio_offset_cfg5_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_86_k_pf3_virtio_offset_cfg5_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_87_k_pf3_virtio_offset_cfg5_cfg_data_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_89_k_pf4_virtio_offset_cfg1_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_90_k_pf4_virtio_offset_cfg1_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_91_k_pf4_virtio_offset_cfg1_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_93_k_pf4_virtio_offset_cfg2_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_94_k_pf4_virtio_offset_cfg2_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_95_k_pf4_virtio_offset_cfg2_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_96_k_pf4_virtio_offset_cfg2_notify_off_multiplier_attr                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_98_k_pf4_virtio_offset_cfg3_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_99_k_pf4_virtio_offset_cfg3_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_cii_ctrl_k_cfg_update_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_cii_ctrl_k_cii_en_attr                                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_cvp_mode                                                                                           = "cvp_disabled",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_drop_vendor0_msg                                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_drop_vendor1_msg                                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_ep_native                                                                                          = "native",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_maxpayload_size                                                                                    = "max_payload_128",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_num_of_lanes                                                                                       = "num_16",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_acs_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_ats_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_bar1_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_bar3_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_bar5_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_dlink_cap_enable                                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_acs_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_ats_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_msix_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_tph_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_virtio_en                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_io_decode                                                                                      = "io32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_ltr_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_msi_enable                                                                                     = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_msix_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_pasid_cap_enable                                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_prefetch_decode                                                                                = "pref64",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_prs_ext_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_ras_des_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sn_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_num_vf_non_ari                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar0_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar1_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar2_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar3_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar4_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar5_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_tph_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_user_vsec_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_virtio_dev_specific_conf_en                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_virtio_en                                                                                      = "pf0_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_vsecras_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_acs_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_ats_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_bar1_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_bar3_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_bar5_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_enable                                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_acs_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_ats_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_msix_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_tph_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_virtio_en                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_msi_enable                                                                                     = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_msix_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_pasid_cap_enable                                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_prs_ext_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_ras_des_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sn_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_num_vf_non_ari                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar0_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar1_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar2_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar3_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar4_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar5_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_tph_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_user_vsec_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_user_vsec_offset                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_virtio_dev_specific_conf_en                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_virtio_en                                                                                      = "pf1_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_vsecras_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_acs_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_ats_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_bar1_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_bar3_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_bar5_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_enable                                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_acs_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_ats_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_msix_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_tph_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_virtio_en                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_msi_enable                                                                                     = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_msix_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_pasid_cap_enable                                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_prs_ext_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_ras_des_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sn_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_num_vf_non_ari                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar0_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar1_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar2_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar3_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar4_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar5_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_tph_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_user_vsec_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_user_vsec_offset                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_virtio_dev_specific_conf_en                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_virtio_en                                                                                      = "pf2_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_vsecras_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_acs_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_ats_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_bar1_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_bar3_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_bar5_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_enable                                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_acs_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_ats_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_msix_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_tph_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_virtio_en                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_msi_enable                                                                                     = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_msix_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_pasid_cap_enable                                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_prs_ext_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_ras_des_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sn_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_num_vf_non_ari                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar0_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar1_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar2_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar3_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar4_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar5_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_tph_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_user_vsec_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_user_vsec_offset                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_virtio_dev_specific_conf_en                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_virtio_en                                                                                      = "pf3_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_vsecras_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_acs_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_ats_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_bar1_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_bar3_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_bar5_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_enable                                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_acs_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_ats_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_msix_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_tph_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_virtio_en                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_msi_enable                                                                                     = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_msix_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_pasid_cap_enable                                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_prs_ext_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_ras_des_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sn_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_num_vf_non_ari                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar0_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar1_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar2_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar3_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar4_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar5_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_tph_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_user_vsec_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_user_vsec_offset                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_virtio_dev_specific_conf_en                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_virtio_en                                                                                      = "pf4_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_vsecras_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_acs_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_ats_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_bar1_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_bar3_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_bar5_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_enable                                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_acs_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_ats_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_msix_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_tph_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_virtio_en                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_msi_enable                                                                                     = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_msix_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_pasid_cap_enable                                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_prs_ext_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_ras_des_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sn_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_num_vf_non_ari                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar0_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar1_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar2_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar3_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar4_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar5_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_tph_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_user_vsec_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_user_vsec_offset                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_virtio_dev_specific_conf_en                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_virtio_en                                                                                      = "pf5_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_vsecras_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_acs_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_ats_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_bar1_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_bar3_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_bar5_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_enable                                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_acs_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_ats_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_msix_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_tph_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_virtio_en                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_msi_enable                                                                                     = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_msix_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_pasid_cap_enable                                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_prs_ext_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_ras_des_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sn_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_num_vf_non_ari                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar0_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar1_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar2_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar3_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar4_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar5_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_tph_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_user_vsec_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_user_vsec_offset                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_virtio_dev_specific_conf_en                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_virtio_en                                                                                      = "pf6_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_vsecras_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_acs_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_ats_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_bar1_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_bar3_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_bar5_mask_bit0                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_enable                                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_acs_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_ats_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_msix_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_tph_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_virtio_en                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_msi_enable                                                                                     = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_msix_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_pasid_cap_enable                                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_prs_ext_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_ras_des_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sn_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_num_vf_non_ari                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar0_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar1_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar2_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar3_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar4_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar5_enabled                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_tph_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_user_vsec_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_user_vsec_offset                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_virtio_dev_specific_conf_en                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_virtio_en                                                                                      = "pf7_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_vsecras_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_ptm_autoupdate                                                                                     = "autoupdate_10ms",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_addr_size0_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_pf_en0_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_start_addr0_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_addr_size1_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_pf_en1_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_start_addr1_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_addr_size2_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_pf_en2_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_start_addr2_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_addr_size3_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_pf_en3_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_start_addr3_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_addr_size4_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_pf_en4_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_start_addr4_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_addr_size5_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_pf_en5_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_start_addr5_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_addr_size6_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_pf_en6_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_start_addr6_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_addr_size7_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_pf_en7_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_start_addr7_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_fixedcred_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_mcred_attr                                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_reloadcred_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_tlp_serr_dis_attr                                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_mmio_access_ctrl_grant_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_opcode_ctrl_lock_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_compressed_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_encrypted_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_devbrd_type_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_vsec_next_offset_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_cvp_irq_en_attr                                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_gpio_irq_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid0_k_jtag_id_0_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid1_k_jtag_id_1_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid2_k_jtag_id_2_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid3_k_jtag_id_3_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_dfd_en_attr                                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_patcntr_en_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_0_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_1_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_2_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_3_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_trig_sel_0_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_trig_sel_1_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_0_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_1_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_2_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_3_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_crs_en_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_rx_lane_flip_en_attr                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_sris_mode_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_tx_lane_flip_en_attr                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_ehp_ctrl0_k_ehp_control_reg_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_outstanding_crd_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_tx_rd_th_attr                                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cvp_cfg_err_en_attr                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dbi_access_err_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr                                                                 = "false",

parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_sd_eq_control1_reg_eval_interval_time = 0,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_multi_lane_control_off_upconfigure_support = "true",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                        = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req                                                            = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_type                                                                                    = "pf0_bar0_mem64",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar1_reg_bar1_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_type                                                                                    = "pf0_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_mem_io                                                                                  = "pf0_bar3_mem",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_type                                                                                    = "pf0_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar5_reg_bar5_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bist_header_type_latency_cache_line_size_reg_multi_func                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_aux_curr                                                                           = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_dsi                                                                                = "pf0_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_pme_support                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_reg_ari_acs_fun_grp_cap                                                                           = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_base_class_code                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_program_interface                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_revision_id                                                                    = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_subclass_code                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_con_status_reg_no_soft_rst                                                                            = "pf0_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                 = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ext_tag_supp                                                         = "pf0_supported",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap                                                              = "pf0_not_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id                                                           = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id                                                           = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_mask                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_config_phy_tx_change                                                                    = "pf0_full_swing",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_select_deemph_var_mux                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_selectable_deemph_bit_mux                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_support_mod_ts                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable                                                          = "pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4                                                     = "gen4_pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5                                                     = "gen5_pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode                                                         = "pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4                                                    = "gen4_pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5                                                    = "gen5_pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec                                                              = 2047,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4                                                         = 927,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5                                                         = 927,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable                                                    = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4                                               = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5                                               = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg4                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg5                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo                                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg4                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg5                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4                                                              = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5                                                              = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_l1_2                                                                         = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_power_off                                                                    = 2,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_comm_mode_support                                                                = 10,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_scale_support                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_value_support                                                             = 5,

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_aspm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_aspm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support = "true",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_aspm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_aspm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_1sub_cap_enable = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_2sub_cap_enable = "disable",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_sca                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_val                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_t_common_mode                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                       = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency                                                        = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_port_num                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                = "pf0_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                    = "pf0_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                        = "pf0_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_misc_control_1_off_port_logic_wr_disable                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_bir                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_table_offset                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported                                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                 = "pf0_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp                                              = "pf0_not_implemented",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pipe_loopback_control_off_pipe_loopback                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_capability_reg_no_eq_needed_support                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rsvdp_11                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precode_req                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precoding_on                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_port_force_off_support_part_lanes_rxei_exit                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_port_link_ctrl_off_fast_link_mode                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                 = "pf0_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                        = "pf0_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_device_spec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pfvf_sel_vsec_enable_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_phy_rxelecidle_k_rxelecidle_disable_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_phy_rxtermination_k_rxtermination_attr                                                                    = 127,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_err_en_correct_err_en_attr                                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_err_en_fatal_err_en_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_err_en_nonfatal_err_en_attr                                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_bw_mgt_int_en_attr                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_eq_req_int_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_pme_int_en_attr                                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_int_en_attr                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_pme_en_attr                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_inta_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_intb_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_intc_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_intd_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_dlycnt_attr                                                                        = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_mode_attr                                                                          = 5,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_dllp_err_sts_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_tlp_err_sts_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_corrected_internal_err_sts_attr                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_dl_protocol_err_sts_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_ecrc_err_sts_attr                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_fc_protocol_err_sts_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_mlf_tlp_err_sts_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_err_sts_attr                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_overflow_err_sts_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_number_rollover_err_sts_attr                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_timer_timeout_err_sts_attr                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_surprise_down_err_sts_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_uncor_internal_err_sts_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tx_common_mode_k_txcommonmode_disable_attr                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cfg_update_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cii_en_attr                                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_cvp_mode                                                                                          = "cvp_disabled",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_drop_vendor0_msg                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_drop_vendor1_msg                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_ep_native                                                                                         = "native",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_maxpayload_size                                                                                   = "max_payload_128",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_num_of_lanes                                                                                      = "num_4",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_acs_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_ats_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_bar1_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_bar3_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_bar5_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_dlink_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_acs_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_ats_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_msix_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_tph_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_io_decode                                                                                     = "io32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_ltr_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_msi_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_msix_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_pasid_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_prefetch_decode                                                                               = "pref64",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_prs_ext_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_ras_des_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_sn_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_tph_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_user_vsec_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_dev_specific_conf_en                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_en                                                                                     = "pf0_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_vsecras_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_ptm_autoupdate                                                                                    = "autoupdate_10ms",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr                                                         = "false",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf0_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf1_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf2_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf3_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf4_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf5_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf6_attr = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf7_attr = "false",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_0_k_cii_addr_size0_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_0_k_cii_pf_en0_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_0_k_cii_start_addr0_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_1_k_cii_addr_size1_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_1_k_cii_pf_en1_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_1_k_cii_start_addr1_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_2_k_cii_addr_size2_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_2_k_cii_pf_en2_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_2_k_cii_start_addr2_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_3_k_cii_addr_size3_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_3_k_cii_pf_en3_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_3_k_cii_start_addr3_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_4_k_cii_addr_size4_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_4_k_cii_pf_en4_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_4_k_cii_start_addr4_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_5_k_cii_addr_size5_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_5_k_cii_pf_en5_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_5_k_cii_start_addr5_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_6_k_cii_addr_size6_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_6_k_cii_pf_en6_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_6_k_cii_start_addr6_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_7_k_cii_addr_size7_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_7_k_cii_pf_en7_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_7_k_cii_start_addr7_attr                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_fixedcred_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_mcred_attr                                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_reloadcred_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_tlp_serr_dis_attr                                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_mmio_access_ctrl_grant_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_opcode_ctrl_lock_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl0_k_compressed_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl0_k_encrypted_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl1_k_devbrd_type_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl1_k_vsec_next_offset_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_irq_ctrl_k_cvp_irq_en_attr                                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_irq_ctrl_k_gpio_irq_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid0_k_jtag_id_0_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid1_k_jtag_id_1_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid2_k_jtag_id_2_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid3_k_jtag_id_3_attr                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_ctrl0_k_dfd_en_attr                                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_ctrl0_k_patcntr_en_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_0_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_1_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_2_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_3_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_trig_sel_0_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_trig_sel_1_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_0_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_1_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_2_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_3_attr                                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_pld_crs_en_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_rx_lane_flip_en_attr                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_sris_mode_attr                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_tx_lane_flip_en_attr                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ehp_ctrl0_k_ehp_control_reg_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ehp_ctrl1_k_outstanding_crd_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ehp_ctrl1_k_tx_rd_th_attr                                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff0_k_exvf_msixpba_bir_pf0_attr                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff0_k_exvf_msixpba_offset_pf0_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff1_k_exvf_msixpba_bir_pf1_attr                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff1_k_exvf_msixpba_offset_pf1_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff2_k_exvf_msixpba_bir_pf2_attr                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff2_k_exvf_msixpba_offset_pf2_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff3_k_exvf_msixpba_bir_pf3_attr                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff3_k_exvf_msixpba_offset_pf3_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff4_k_exvf_msixpba_bir_pf4_attr                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff4_k_exvf_msixpba_offset_pf4_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff5_k_exvf_msixpba_bir_pf5_attr                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff5_k_exvf_msixpba_offset_pf5_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff6_k_exvf_msixpba_bir_pf6_attr                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff6_k_exvf_msixpba_offset_pf6_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff7_k_exvf_msixpba_bir_pf7_attr                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff7_k_exvf_msixpba_offset_pf7_attr                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff0_k_exvf_msixtable_bir_pf0_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff0_k_exvf_msixtable_offset_pf0_attr                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff1_k_exvf_msixtable_bir_pf1_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff1_k_exvf_msixtable_offset_pf1_attr                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff2_k_exvf_msixtable_bir_pf2_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff2_k_exvf_msixtable_offset_pf2_attr                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff3_k_exvf_msixtable_bir_pf3_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff3_k_exvf_msixtable_offset_pf3_attr                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff4_k_exvf_msixtable_bir_pf4_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff4_k_exvf_msixtable_offset_pf4_attr                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff5_k_exvf_msixtable_bir_pf5_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff5_k_exvf_msixtable_offset_pf5_attr                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff6_k_exvf_msixtable_bir_pf6_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff6_k_exvf_msixtable_offset_pf6_attr                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff7_k_exvf_msixtable_bir_pf7_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff7_k_exvf_msixtable_offset_pf7_attr                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize0_k_exvf_msix_tablesize_pf0_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize0_k_exvf_msix_tablesize_pf1_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize1_k_exvf_msix_tablesize_pf2_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize1_k_exvf_msix_tablesize_pf3_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize2_k_exvf_msix_tablesize_pf4_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize2_k_exvf_msix_tablesize_pf5_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize3_k_exvf_msix_tablesize_pf6_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize3_k_exvf_msix_tablesize_pf7_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_cvp_cfg_err_en_attr                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_dbi_access_err_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr                                                                 = "false",

parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sd_eq_control1_reg_eval_interval_time = 0,
parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sd_eq_control1_reg_eval_interval_time = 0,

parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_multi_lane_control_off_upconfigure_support = "true",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                        = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req                                                            = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_reg_bar0_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_reg_bar0_type                                                                                    = "pf0_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar1_reg_bar1_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_reg_bar2_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_reg_bar2_type                                                                                    = "pf0_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_reg_bar3_mem_io                                                                                  = "pf0_bar3_mem",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_reg_bar3_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_reg_bar4_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_reg_bar4_type                                                                                    = "pf0_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar5_reg_bar5_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_id_nxt_ptr_reg_aux_curr                                                                           = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_id_nxt_ptr_reg_dsi                                                                                = "pf0_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_id_nxt_ptr_reg_pme_support                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_reg_ari_acs_fun_grp_cap                                                                           = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_base_class_code                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_program_interface                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_revision_id                                                                    = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_subclass_code                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_con_status_reg_no_soft_rst                                                                            = "pf0_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                 = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_ext_tag_supp                                                         = "pf0_not_supported",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap                                                              = "pf0_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id                                                           = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id                                                           = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_exp_rom_bar_mask_reg_rom_mask                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_config_phy_tx_change                                                                    = "pf0_full_swing",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_select_deemph_var_mux                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_selectable_deemph_bit_mux                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_support_mod_ts                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable                                                          = "pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4                                                     = "gen4_pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5                                                     = "gen5_pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode                                                         = "pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4                                                    = "gen4_pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5                                                    = "gen5_pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec                                                              = 2047,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4                                                         = 927,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5                                                         = 927,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable                                                    = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4                                               = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5                                               = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_eieos_cnt                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_phase_2_3                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_phase_2_3_atg4                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_phase_2_3_atg5                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_redo                                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_redo_atg4                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_redo_atg5                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_gen3_equalization_disable                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_ph01_en                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts                                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4                                                              = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5                                                              = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1_substates_off_l1sub_t_l1_2                                                                         = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1_substates_off_l1sub_t_power_off                                                                    = 2,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_comm_mode_support                                                                = 10,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_pwr_on_scale_support                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_pwr_on_value_support                                                             = 5,

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_1_aspm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_2_aspm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support = "true",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_1_aspm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_aspm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_l1_1sub_cap_enable = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_l1_2sub_cap_enable = "disable",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_th_sca                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_th_val                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_t_common_mode                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                       = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency                                                        = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_port_num                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                = "pf0_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                    = "pf0_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                        = "pf0_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_table_offset_reg_pci_msix_bir                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_table_offset_reg_pci_msix_table_offset                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported                                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                 = "pf0_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp                                              = "pf0_not_implemented",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pipe_loopback_control_off_pipe_loopback                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset4                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset5                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset6                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset7                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset4                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset5                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset6                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset7                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset4                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset5                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset6                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset7                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset4                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset5                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset6                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset7                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_capability_reg_no_eq_needed_support                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_rsvdp_11                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_tx_precode_req                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_tx_precoding_on                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_port_force_off_support_part_lanes_rxei_exit                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_port_link_ctrl_off_fast_link_mode                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                 = "pf0_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint4                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint5                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset4                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset5                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint4                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint5                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset4                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset5                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint6                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint7                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset6                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset7                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint6                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint7                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset6                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset7                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_type                                                                     = "pf0_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_type                                                                     = "pf0_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_type                                                                     = "pf0_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_vf_offset_position_sriov_vf_offset                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_vf_offset_position_sriov_vf_stride                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sup_page_sizes_reg_sriov_sup_page_size                                                                = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                        = "pf0_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_device_spec                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_vf_device_id_reg_sriov_vf_device_id                                                                   = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_at_block                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                        = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_src_valid                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ats_capabilities_ctrl_reg_invalidate_q_depth                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ats_capabilities_ctrl_reg_page_aligned_req                                                            = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_mask_reg_pci_type0_bar0_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_mask_reg_pci_type0_bar0_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_reg_bar0_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_reg_bar0_type                                                                                    = "pf1_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar1_mask_reg_pci_type0_bar1_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar1_mask_reg_pci_type0_bar1_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar1_reg_bar1_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_mask_reg_pci_type0_bar2_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_mask_reg_pci_type0_bar2_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_reg_bar2_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_reg_bar2_type                                                                                    = "pf1_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar3_mask_reg_pci_type0_bar3_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar3_mask_reg_pci_type0_bar3_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar3_reg_bar3_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_mask_reg_pci_type0_bar4_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_mask_reg_pci_type0_bar4_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_reg_bar4_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_reg_bar4_type                                                                                    = "pf1_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar5_mask_reg_pci_type0_bar5_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar5_mask_reg_pci_type0_bar5_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar5_reg_bar5_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cap_id_nxt_ptr_reg_aux_curr                                                                           = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cap_id_nxt_ptr_reg_dsi                                                                                = "pf1_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cap_id_nxt_ptr_reg_pme_support                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_base_class_code                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_program_interface                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_revision_id                                                                    = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_subclass_code                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_con_status_reg_no_soft_rst                                                                            = "pf1_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                 = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_ext_tag_supp                                                         = "pf1_supported",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_flr_cap                                                              = "pf1_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_control_device_status_pcie_cap_ext_tag_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_id_vendor_id_reg_pci_type0_device_id                                                           = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_id_vendor_id_reg_pci_type0_vendor_id                                                           = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_exp_rom_bar_mask_reg_rom_bar_enabled                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_exp_rom_bar_mask_reg_rom_mask                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_exp_rom_base_addr_reg_rom_bar_enable                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                       = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_capabilities_reg_pcie_cap_l1_exit_latency                                                        = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_capabilities_reg_pcie_cap_port_num                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                = "pf1_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                    = "pf1_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_control_link_status_reg_pcie_cap_slot_clk_config                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                        = "pf1_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_pba_offset_reg_pci_msix_pba_bir                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_pba_offset_reg_pci_msix_pba_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_table_offset_reg_pci_msix_bir                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_table_offset_reg_pci_msix_table_offset                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pasid_cap_cntrl_reg_execute_permission_supported                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pasid_cap_cntrl_reg_max_pasid_width                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pasid_cap_cntrl_reg_privileged_mode_supported                                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                 = "pf1_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                 = "pf1_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_type                                                                     = "pf1_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_type                                                                     = "pf1_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_type                                                                     = "pf1_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_vf_offset_position_sriov_vf_offset                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_vf_offset_position_sriov_vf_stride                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sup_page_sizes_reg_sriov_sup_page_size                                                                = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                        = "pf1_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_device_spec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_vf_device_id_reg_sriov_vf_device_id                                                                   = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_at_block                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                        = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_src_valid                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ats_capabilities_ctrl_reg_invalidate_q_depth                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ats_capabilities_ctrl_reg_page_aligned_req                                                            = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_mask_reg_pci_type0_bar0_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_mask_reg_pci_type0_bar0_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_reg_bar0_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_reg_bar0_type                                                                                    = "pf2_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar1_mask_reg_pci_type0_bar1_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar1_mask_reg_pci_type0_bar1_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar1_reg_bar1_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_mask_reg_pci_type0_bar2_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_mask_reg_pci_type0_bar2_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_reg_bar2_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_reg_bar2_type                                                                                    = "pf2_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar3_mask_reg_pci_type0_bar3_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar3_mask_reg_pci_type0_bar3_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar3_reg_bar3_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_mask_reg_pci_type0_bar4_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_mask_reg_pci_type0_bar4_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_reg_bar4_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_reg_bar4_type                                                                                    = "pf2_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar5_mask_reg_pci_type0_bar5_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar5_mask_reg_pci_type0_bar5_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar5_reg_bar5_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cap_id_nxt_ptr_reg_aux_curr                                                                           = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cap_id_nxt_ptr_reg_dsi                                                                                = "pf2_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cap_id_nxt_ptr_reg_pme_support                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_base_class_code                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_program_interface                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_revision_id                                                                    = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_subclass_code                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_con_status_reg_no_soft_rst                                                                            = "pf2_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                 = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_ext_tag_supp                                                         = "pf2_supported",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_flr_cap                                                              = "pf2_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_control_device_status_pcie_cap_ext_tag_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_id_vendor_id_reg_pci_type0_device_id                                                           = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_id_vendor_id_reg_pci_type0_vendor_id                                                           = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_exp_rom_bar_mask_reg_rom_bar_enabled                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_exp_rom_bar_mask_reg_rom_mask                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_exp_rom_base_addr_reg_rom_bar_enable                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                       = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_capabilities_reg_pcie_cap_l1_exit_latency                                                        = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_capabilities_reg_pcie_cap_port_num                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                = "pf2_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                    = "pf2_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_control_link_status_reg_pcie_cap_slot_clk_config                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                        = "pf2_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_pba_offset_reg_pci_msix_pba_bir                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_pba_offset_reg_pci_msix_pba_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_table_offset_reg_pci_msix_bir                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_table_offset_reg_pci_msix_table_offset                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pasid_cap_cntrl_reg_execute_permission_supported                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pasid_cap_cntrl_reg_max_pasid_width                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pasid_cap_cntrl_reg_privileged_mode_supported                                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                 = "pf2_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                 = "pf2_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_type                                                                     = "pf2_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_type                                                                     = "pf2_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_type                                                                     = "pf2_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_vf_offset_position_sriov_vf_offset                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_vf_offset_position_sriov_vf_stride                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sup_page_sizes_reg_sriov_sup_page_size                                                                = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                        = "pf2_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_device_spec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_vf_device_id_reg_sriov_vf_device_id                                                                   = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_at_block                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                        = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_src_valid                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ats_capabilities_ctrl_reg_invalidate_q_depth                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ats_capabilities_ctrl_reg_page_aligned_req                                                            = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_mask_reg_pci_type0_bar0_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_mask_reg_pci_type0_bar0_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_reg_bar0_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_reg_bar0_type                                                                                    = "pf3_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar1_mask_reg_pci_type0_bar1_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar1_mask_reg_pci_type0_bar1_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar1_reg_bar1_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_mask_reg_pci_type0_bar2_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_mask_reg_pci_type0_bar2_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_reg_bar2_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_reg_bar2_type                                                                                    = "pf3_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar3_mask_reg_pci_type0_bar3_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar3_mask_reg_pci_type0_bar3_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar3_reg_bar3_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_mask_reg_pci_type0_bar4_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_mask_reg_pci_type0_bar4_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_reg_bar4_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_reg_bar4_type                                                                                    = "pf3_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar5_mask_reg_pci_type0_bar5_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar5_mask_reg_pci_type0_bar5_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar5_reg_bar5_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cap_id_nxt_ptr_reg_aux_curr                                                                           = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cap_id_nxt_ptr_reg_dsi                                                                                = "pf3_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cap_id_nxt_ptr_reg_pme_support                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_base_class_code                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_program_interface                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_revision_id                                                                    = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_subclass_code                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_con_status_reg_no_soft_rst                                                                            = "pf3_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                 = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_ext_tag_supp                                                         = "pf3_supported",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_flr_cap                                                              = "pf3_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_control_device_status_pcie_cap_ext_tag_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_id_vendor_id_reg_pci_type0_device_id                                                           = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_id_vendor_id_reg_pci_type0_vendor_id                                                           = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_exp_rom_bar_mask_reg_rom_bar_enabled                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_exp_rom_bar_mask_reg_rom_mask                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_exp_rom_base_addr_reg_rom_bar_enable                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                       = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_capabilities_reg_pcie_cap_l1_exit_latency                                                        = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_capabilities_reg_pcie_cap_port_num                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                = "pf3_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                    = "pf3_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_control_link_status_reg_pcie_cap_slot_clk_config                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                        = "pf3_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_pba_offset_reg_pci_msix_pba_bir                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_pba_offset_reg_pci_msix_pba_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_table_offset_reg_pci_msix_bir                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_table_offset_reg_pci_msix_table_offset                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pasid_cap_cntrl_reg_execute_permission_supported                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pasid_cap_cntrl_reg_max_pasid_width                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pasid_cap_cntrl_reg_privileged_mode_supported                                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                 = "pf3_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                 = "pf3_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_type                                                                     = "pf3_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_type                                                                     = "pf3_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_type                                                                     = "pf3_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_vf_offset_position_sriov_vf_offset                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_vf_offset_position_sriov_vf_stride                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sup_page_sizes_reg_sriov_sup_page_size                                                                = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                        = "pf3_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_device_spec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_vf_device_id_reg_sriov_vf_device_id                                                                   = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_at_block                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                        = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_src_valid                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ats_capabilities_ctrl_reg_invalidate_q_depth                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ats_capabilities_ctrl_reg_page_aligned_req                                                            = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_mask_reg_pci_type0_bar0_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_mask_reg_pci_type0_bar0_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_reg_bar0_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_reg_bar0_type                                                                                    = "pf4_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar1_mask_reg_pci_type0_bar1_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar1_mask_reg_pci_type0_bar1_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar1_reg_bar1_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_mask_reg_pci_type0_bar2_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_mask_reg_pci_type0_bar2_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_reg_bar2_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_reg_bar2_type                                                                                    = "pf4_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar3_mask_reg_pci_type0_bar3_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar3_mask_reg_pci_type0_bar3_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar3_reg_bar3_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_mask_reg_pci_type0_bar4_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_mask_reg_pci_type0_bar4_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_reg_bar4_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_reg_bar4_type                                                                                    = "pf4_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar5_mask_reg_pci_type0_bar5_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar5_mask_reg_pci_type0_bar5_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar5_reg_bar5_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cap_id_nxt_ptr_reg_aux_curr                                                                           = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cap_id_nxt_ptr_reg_dsi                                                                                = "pf4_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cap_id_nxt_ptr_reg_pme_support                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_base_class_code                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_program_interface                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_revision_id                                                                    = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_subclass_code                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_con_status_reg_no_soft_rst                                                                            = "pf4_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                 = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_ext_tag_supp                                                         = "pf4_supported",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_flr_cap                                                              = "pf4_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_control_device_status_pcie_cap_ext_tag_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_id_vendor_id_reg_pci_type0_device_id                                                           = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_id_vendor_id_reg_pci_type0_vendor_id                                                           = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_exp_rom_bar_mask_reg_rom_bar_enabled                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_exp_rom_bar_mask_reg_rom_mask                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_exp_rom_base_addr_reg_rom_bar_enable                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                       = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_capabilities_reg_pcie_cap_l1_exit_latency                                                        = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_capabilities_reg_pcie_cap_port_num                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                = "pf4_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                    = "pf4_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_control_link_status_reg_pcie_cap_slot_clk_config                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                        = "pf4_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_pba_offset_reg_pci_msix_pba_bir                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_pba_offset_reg_pci_msix_pba_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_table_offset_reg_pci_msix_bir                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_table_offset_reg_pci_msix_table_offset                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pasid_cap_cntrl_reg_execute_permission_supported                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pasid_cap_cntrl_reg_max_pasid_width                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pasid_cap_cntrl_reg_privileged_mode_supported                                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                 = "pf4_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                 = "pf4_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_type                                                                     = "pf4_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_type                                                                     = "pf4_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_type                                                                     = "pf4_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_vf_offset_position_sriov_vf_offset                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_vf_offset_position_sriov_vf_stride                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sup_page_sizes_reg_sriov_sup_page_size                                                                = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                        = "pf4_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_device_spec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_vf_device_id_reg_sriov_vf_device_id                                                                   = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_at_block                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                        = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_src_valid                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ats_capabilities_ctrl_reg_invalidate_q_depth                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ats_capabilities_ctrl_reg_page_aligned_req                                                            = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_mask_reg_pci_type0_bar0_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_mask_reg_pci_type0_bar0_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_reg_bar0_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_reg_bar0_type                                                                                    = "pf5_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar1_mask_reg_pci_type0_bar1_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar1_mask_reg_pci_type0_bar1_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar1_reg_bar1_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_mask_reg_pci_type0_bar2_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_mask_reg_pci_type0_bar2_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_reg_bar2_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_reg_bar2_type                                                                                    = "pf5_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar3_mask_reg_pci_type0_bar3_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar3_mask_reg_pci_type0_bar3_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar3_reg_bar3_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_mask_reg_pci_type0_bar4_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_mask_reg_pci_type0_bar4_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_reg_bar4_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_reg_bar4_type                                                                                    = "pf5_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar5_mask_reg_pci_type0_bar5_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar5_mask_reg_pci_type0_bar5_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar5_reg_bar5_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cap_id_nxt_ptr_reg_aux_curr                                                                           = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cap_id_nxt_ptr_reg_dsi                                                                                = "pf5_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cap_id_nxt_ptr_reg_pme_support                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_base_class_code                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_program_interface                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_revision_id                                                                    = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_subclass_code                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_con_status_reg_no_soft_rst                                                                            = "pf5_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                 = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_ext_tag_supp                                                         = "pf5_supported",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_flr_cap                                                              = "pf5_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_control_device_status_pcie_cap_ext_tag_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_id_vendor_id_reg_pci_type0_device_id                                                           = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_id_vendor_id_reg_pci_type0_vendor_id                                                           = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_exp_rom_bar_mask_reg_rom_bar_enabled                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_exp_rom_bar_mask_reg_rom_mask                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_exp_rom_base_addr_reg_rom_bar_enable                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                       = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_capabilities_reg_pcie_cap_l1_exit_latency                                                        = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_capabilities_reg_pcie_cap_port_num                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                = "pf5_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                    = "pf5_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_control_link_status_reg_pcie_cap_slot_clk_config                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                        = "pf5_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_pba_offset_reg_pci_msix_pba_bir                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_pba_offset_reg_pci_msix_pba_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_table_offset_reg_pci_msix_bir                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_table_offset_reg_pci_msix_table_offset                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pasid_cap_cntrl_reg_execute_permission_supported                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pasid_cap_cntrl_reg_max_pasid_width                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pasid_cap_cntrl_reg_privileged_mode_supported                                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                 = "pf5_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                 = "pf5_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_type                                                                     = "pf5_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_type                                                                     = "pf5_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_type                                                                     = "pf5_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_vf_offset_position_sriov_vf_offset                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_vf_offset_position_sriov_vf_stride                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sup_page_sizes_reg_sriov_sup_page_size                                                                = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                        = "pf5_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_device_spec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_vf_device_id_reg_sriov_vf_device_id                                                                   = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_at_block                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                        = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_src_valid                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ats_capabilities_ctrl_reg_invalidate_q_depth                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ats_capabilities_ctrl_reg_page_aligned_req                                                            = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_mask_reg_pci_type0_bar0_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_mask_reg_pci_type0_bar0_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_reg_bar0_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_reg_bar0_type                                                                                    = "pf6_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar1_mask_reg_pci_type0_bar1_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar1_mask_reg_pci_type0_bar1_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar1_reg_bar1_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_mask_reg_pci_type0_bar2_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_mask_reg_pci_type0_bar2_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_reg_bar2_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_reg_bar2_type                                                                                    = "pf6_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar3_mask_reg_pci_type0_bar3_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar3_mask_reg_pci_type0_bar3_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar3_reg_bar3_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_mask_reg_pci_type0_bar4_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_mask_reg_pci_type0_bar4_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_reg_bar4_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_reg_bar4_type                                                                                    = "pf6_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar5_mask_reg_pci_type0_bar5_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar5_mask_reg_pci_type0_bar5_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar5_reg_bar5_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cap_id_nxt_ptr_reg_aux_curr                                                                           = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cap_id_nxt_ptr_reg_dsi                                                                                = "pf6_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cap_id_nxt_ptr_reg_pme_support                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_base_class_code                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_program_interface                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_revision_id                                                                    = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_subclass_code                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_con_status_reg_no_soft_rst                                                                            = "pf6_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                 = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_ext_tag_supp                                                         = "pf6_supported",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_flr_cap                                                              = "pf6_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_control_device_status_pcie_cap_ext_tag_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_id_vendor_id_reg_pci_type0_device_id                                                           = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_id_vendor_id_reg_pci_type0_vendor_id                                                           = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_exp_rom_bar_mask_reg_rom_bar_enabled                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_exp_rom_bar_mask_reg_rom_mask                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_exp_rom_base_addr_reg_rom_bar_enable                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                       = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_capabilities_reg_pcie_cap_l1_exit_latency                                                        = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_capabilities_reg_pcie_cap_port_num                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                = "pf6_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                    = "pf6_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_control_link_status_reg_pcie_cap_slot_clk_config                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                        = "pf6_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_pba_offset_reg_pci_msix_pba_bir                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_pba_offset_reg_pci_msix_pba_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_table_offset_reg_pci_msix_bir                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_table_offset_reg_pci_msix_table_offset                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pasid_cap_cntrl_reg_execute_permission_supported                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pasid_cap_cntrl_reg_max_pasid_width                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pasid_cap_cntrl_reg_privileged_mode_supported                                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                 = "pf6_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                 = "pf6_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_type                                                                     = "pf6_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_type                                                                     = "pf6_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_type                                                                     = "pf6_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_vf_offset_position_sriov_vf_offset                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_vf_offset_position_sriov_vf_stride                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sup_page_sizes_reg_sriov_sup_page_size                                                                = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                        = "pf6_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_device_spec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_vf_device_id_reg_sriov_vf_device_id                                                                   = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_at_block                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                   = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                        = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_src_valid                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ats_capabilities_ctrl_reg_invalidate_q_depth                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ats_capabilities_ctrl_reg_page_aligned_req                                                            = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_mask_reg_pci_type0_bar0_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_mask_reg_pci_type0_bar0_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_reg_bar0_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_reg_bar0_type                                                                                    = "pf7_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar1_mask_reg_pci_type0_bar1_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar1_mask_reg_pci_type0_bar1_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar1_reg_bar1_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_mask_reg_pci_type0_bar2_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_mask_reg_pci_type0_bar2_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_reg_bar2_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_reg_bar2_type                                                                                    = "pf7_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar3_mask_reg_pci_type0_bar3_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar3_mask_reg_pci_type0_bar3_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar3_reg_bar3_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_mask_reg_pci_type0_bar4_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_mask_reg_pci_type0_bar4_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_reg_bar4_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_reg_bar4_type                                                                                    = "pf7_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar5_mask_reg_pci_type0_bar5_enabled                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar5_mask_reg_pci_type0_bar5_mask                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar5_reg_bar5_prefetch                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cap_id_nxt_ptr_reg_aux_curr                                                                           = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cap_id_nxt_ptr_reg_dsi                                                                                = "pf7_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cap_id_nxt_ptr_reg_pme_support                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cardbus_cis_ptr_reg_cardbus_cis_pointer                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_base_class_code                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_program_interface                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_revision_id                                                                    = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_subclass_code                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_con_status_reg_no_soft_rst                                                                            = "pf7_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                 = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                  = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_ext_tag_supp                                                         = "pf7_supported",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_flr_cap                                                              = "pf7_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_control_device_status_pcie_cap_ext_tag_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_id_vendor_id_reg_pci_type0_device_id                                                           = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_id_vendor_id_reg_pci_type0_vendor_id                                                           = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_exp_rom_bar_mask_reg_rom_bar_enabled                                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_exp_rom_bar_mask_reg_rom_mask                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_exp_rom_base_addr_reg_rom_bar_enable                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                       = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_capabilities_reg_pcie_cap_l1_exit_latency                                                        = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_capabilities_reg_pcie_cap_port_num                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                = "pf7_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                    = "pf7_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_control_link_status_reg_pcie_cap_slot_clk_config                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                        = "pf7_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_pba_offset_reg_pci_msix_pba_bir                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_pba_offset_reg_pci_msix_pba_offset                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_table_offset_reg_pci_msix_bir                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_table_offset_reg_pci_msix_table_offset                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pasid_cap_cntrl_reg_execute_permission_supported                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pasid_cap_cntrl_reg_max_pasid_width                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pasid_cap_cntrl_reg_privileged_mode_supported                                                         = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                  = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                 = "pf7_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride                                                = 256,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                 = "pf7_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar0_mask_reg_pci_sriov_bar0_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_type                                                                     = "pf7_sriov_vf_bar0_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar1_mask_reg_pci_sriov_bar1_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar1_reg_sriov_vf_bar1_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar2_mask_reg_pci_sriov_bar2_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_type                                                                     = "pf7_sriov_vf_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar3_mask_reg_pci_sriov_bar3_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar3_reg_sriov_vf_bar3_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar4_mask_reg_pci_sriov_bar4_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_type                                                                     = "pf7_sriov_vf_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar5_mask_reg_pci_sriov_bar5_mask                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar5_reg_sriov_vf_bar5_prefetch                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_vf_offset_position_sriov_vf_offset                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_vf_offset_position_sriov_vf_stride                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sup_page_sizes_reg_sriov_sup_page_size                                                                = 1363,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                        = "pf7_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_device_spec                                                               = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_vf_device_id_reg_sriov_vf_device_id                                                                   = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pfvf_sel_vsec_enable_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_phy_rxelecidle_k_rxelecidle_disable_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_phy_rxtermination_k_rxtermination_attr                                                                    = 127,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ptm_ctrl_k_cfg_ptm_auto_update_signal_attr                                                                = "false",

parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ptm_adj_lsb_k_cfg_ptm_local_clock_adj_lsb_attr = 0,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ptm_adj_msb_k_cfg_ptm_local_clock_adj_msb_attr = 0,

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_err_en_correct_err_en_attr                                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_err_en_fatal_err_en_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_err_en_nonfatal_err_en_attr                                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_bw_mgt_int_en_attr                                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_link_eq_req_int_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_pme_int_en_attr                                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_hp_int_en_attr                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_hp_pme_en_attr                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_inta_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_intb_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_intc_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_intd_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_sriov_misc_ctrl_k_nonsriov_mode_attr                                                                      = 255,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_stagger_control_k_stag_dlycnt_attr                                                                        = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_stagger_control_k_stag_mode_attr                                                                          = 5,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id0_k_exvf_subsysid_pf0_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id0_k_exvf_subsysid_pf1_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id1_k_exvf_subsysid_pf2_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id1_k_exvf_subsysid_pf3_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id2_k_exvf_subsysid_pf4_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id2_k_exvf_subsysid_pf5_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id3_k_exvf_subsysid_pf6_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id3_k_exvf_subsysid_pf7_attr                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf0_attr                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf1_attr                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablesize_pf0_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablesize_pf1_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf2_attr                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf3_attr                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablesize_pf2_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablesize_pf3_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf4_attr                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf5_attr                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablesize_pf4_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablesize_pf5_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf6_attr                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf7_attr                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablesize_pf6_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablesize_pf7_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tx_common_mode_k_txcommonmode_disable_attr                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_100_k_pf4_virtio_offset_cfg3_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_102_k_pf4_virtio_offset_cfg4_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_103_k_pf4_virtio_offset_cfg4_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_104_k_pf4_virtio_offset_cfg4_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_106_k_pf4_virtio_offset_cfg5_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_107_k_pf4_virtio_offset_cfg5_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_108_k_pf4_virtio_offset_cfg5_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_109_k_pf4_virtio_offset_cfg5_cfg_data_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_111_k_pf5_virtio_offset_cfg1_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_112_k_pf5_virtio_offset_cfg1_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_113_k_pf5_virtio_offset_cfg1_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_115_k_pf5_virtio_offset_cfg2_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_116_k_pf5_virtio_offset_cfg2_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_117_k_pf5_virtio_offset_cfg2_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_118_k_pf5_virtio_offset_cfg2_notify_off_multiplier_attr                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_120_k_pf5_virtio_offset_cfg3_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_121_k_pf5_virtio_offset_cfg3_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_122_k_pf5_virtio_offset_cfg3_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_124_k_pf5_virtio_offset_cfg4_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_125_k_pf5_virtio_offset_cfg4_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_126_k_pf5_virtio_offset_cfg4_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_128_k_pf5_virtio_offset_cfg5_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_129_k_pf5_virtio_offset_cfg5_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_130_k_pf5_virtio_offset_cfg5_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_131_k_pf5_virtio_offset_cfg5_cfg_data_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_133_k_pf6_virtio_offset_cfg1_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_134_k_pf6_virtio_offset_cfg1_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_135_k_pf6_virtio_offset_cfg1_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_137_k_pf6_virtio_offset_cfg2_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_138_k_pf6_virtio_offset_cfg2_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_139_k_pf6_virtio_offset_cfg2_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_140_k_pf6_virtio_offset_cfg2_notify_off_multiplier_attr                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_142_k_pf6_virtio_offset_cfg3_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_143_k_pf6_virtio_offset_cfg3_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_144_k_pf6_virtio_offset_cfg3_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_146_k_pf6_virtio_offset_cfg4_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_147_k_pf6_virtio_offset_cfg4_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_148_k_pf6_virtio_offset_cfg4_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_150_k_pf6_virtio_offset_cfg5_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_151_k_pf6_virtio_offset_cfg5_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_152_k_pf6_virtio_offset_cfg5_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_153_k_pf6_virtio_offset_cfg5_cfg_data_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_155_k_pf7_virtio_offset_cfg1_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_156_k_pf7_virtio_offset_cfg1_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_157_k_pf7_virtio_offset_cfg1_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_159_k_pf7_virtio_offset_cfg2_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_160_k_pf7_virtio_offset_cfg2_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_161_k_pf7_virtio_offset_cfg2_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_162_k_pf7_virtio_offset_cfg2_notify_off_multiplier_attr                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_164_k_pf7_virtio_offset_cfg3_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_165_k_pf7_virtio_offset_cfg3_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_166_k_pf7_virtio_offset_cfg3_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_168_k_pf7_virtio_offset_cfg4_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_169_k_pf7_virtio_offset_cfg4_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_170_k_pf7_virtio_offset_cfg4_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_172_k_pf7_virtio_offset_cfg5_cap_bar_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_173_k_pf7_virtio_offset_cfg5_cap_offset_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_174_k_pf7_virtio_offset_cfg5_cap_length_attr                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_175_k_pf7_virtio_offset_cfg5_cfg_data_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_23_k_pf1_virtio_offset_cfg1_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_24_k_pf1_virtio_offset_cfg1_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_25_k_pf1_virtio_offset_cfg1_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_27_k_pf1_virtio_offset_cfg2_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_28_k_pf1_virtio_offset_cfg2_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_29_k_pf1_virtio_offset_cfg2_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_30_k_pf1_virtio_offset_cfg2_notify_off_multiplier_attr                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_32_k_pf1_virtio_offset_cfg3_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_33_k_pf1_virtio_offset_cfg3_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_34_k_pf1_virtio_offset_cfg3_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_36_k_pf1_virtio_offset_cfg4_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_37_k_pf1_virtio_offset_cfg4_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_38_k_pf1_virtio_offset_cfg4_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_40_k_pf1_virtio_offset_cfg5_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_41_k_pf1_virtio_offset_cfg5_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_42_k_pf1_virtio_offset_cfg5_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_43_k_pf1_virtio_offset_cfg5_cfg_data_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_45_k_pf2_virtio_offset_cfg1_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_46_k_pf2_virtio_offset_cfg1_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_47_k_pf2_virtio_offset_cfg1_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_49_k_pf2_virtio_offset_cfg2_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_50_k_pf2_virtio_offset_cfg2_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_51_k_pf2_virtio_offset_cfg2_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_52_k_pf2_virtio_offset_cfg2_notify_off_multiplier_attr                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_54_k_pf2_virtio_offset_cfg3_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_55_k_pf2_virtio_offset_cfg3_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_56_k_pf2_virtio_offset_cfg3_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_58_k_pf2_virtio_offset_cfg4_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_59_k_pf2_virtio_offset_cfg4_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_60_k_pf2_virtio_offset_cfg4_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_62_k_pf2_virtio_offset_cfg5_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_63_k_pf2_virtio_offset_cfg5_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_64_k_pf2_virtio_offset_cfg5_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_65_k_pf2_virtio_offset_cfg5_cfg_data_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_67_k_pf3_virtio_offset_cfg1_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_68_k_pf3_virtio_offset_cfg1_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_69_k_pf3_virtio_offset_cfg1_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_71_k_pf3_virtio_offset_cfg2_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_72_k_pf3_virtio_offset_cfg2_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_73_k_pf3_virtio_offset_cfg2_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_74_k_pf3_virtio_offset_cfg2_notify_off_multiplier_attr                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_76_k_pf3_virtio_offset_cfg3_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_77_k_pf3_virtio_offset_cfg3_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_78_k_pf3_virtio_offset_cfg3_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_80_k_pf3_virtio_offset_cfg4_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_81_k_pf3_virtio_offset_cfg4_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_82_k_pf3_virtio_offset_cfg4_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_84_k_pf3_virtio_offset_cfg5_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_85_k_pf3_virtio_offset_cfg5_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_86_k_pf3_virtio_offset_cfg5_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_87_k_pf3_virtio_offset_cfg5_cfg_data_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_89_k_pf4_virtio_offset_cfg1_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_90_k_pf4_virtio_offset_cfg1_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_91_k_pf4_virtio_offset_cfg1_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_93_k_pf4_virtio_offset_cfg2_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_94_k_pf4_virtio_offset_cfg2_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_95_k_pf4_virtio_offset_cfg2_cap_length_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_96_k_pf4_virtio_offset_cfg2_notify_off_multiplier_attr                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_98_k_pf4_virtio_offset_cfg3_cap_bar_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_99_k_pf4_virtio_offset_cfg3_cap_offset_attr                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_cii_ctrl_k_cfg_update_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_cii_ctrl_k_cii_en_attr                                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_cvp_mode                                                                                          = "cvp_disabled",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_drop_vendor0_msg                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_drop_vendor1_msg                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_ep_native                                                                                         = "native",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_maxpayload_size                                                                                   = "max_payload_128",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_num_of_lanes                                                                                      = "num_8",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_acs_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_ats_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_bar1_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_bar3_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_bar5_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_dlink_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_acs_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_ats_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_msix_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_tph_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_virtio_en                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_io_decode                                                                                     = "io32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_ltr_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_msi_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_msix_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_pasid_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_prefetch_decode                                                                               = "pref64",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_prs_ext_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_ras_des_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sn_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_num_vf_non_ari                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar0_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar1_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar2_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar3_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar4_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar5_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_tph_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_user_vsec_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_virtio_dev_specific_conf_en                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_virtio_en                                                                                     = "pf0_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_vsecras_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_acs_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_ats_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_bar1_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_bar3_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_bar5_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_enable                                                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_acs_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_ats_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_msix_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_tph_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_virtio_en                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_msi_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_msix_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_pasid_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_prs_ext_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_ras_des_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sn_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_num_vf_non_ari                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar0_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar1_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar2_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar3_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar4_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar5_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_tph_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_user_vsec_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_user_vsec_offset                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_virtio_dev_specific_conf_en                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_virtio_en                                                                                     = "pf1_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_vsecras_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_acs_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_ats_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_bar1_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_bar3_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_bar5_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_enable                                                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_acs_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_ats_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_msix_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_tph_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_virtio_en                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_msi_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_msix_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_pasid_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_prs_ext_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_ras_des_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sn_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_num_vf_non_ari                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar0_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar1_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar2_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar3_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar4_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar5_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_tph_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_user_vsec_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_user_vsec_offset                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_virtio_dev_specific_conf_en                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_virtio_en                                                                                     = "pf2_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_vsecras_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_acs_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_ats_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_bar1_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_bar3_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_bar5_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_enable                                                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_acs_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_ats_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_msix_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_tph_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_virtio_en                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_msi_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_msix_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_pasid_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_prs_ext_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_ras_des_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sn_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_num_vf_non_ari                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar0_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar1_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar2_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar3_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar4_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar5_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_tph_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_user_vsec_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_user_vsec_offset                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_virtio_dev_specific_conf_en                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_virtio_en                                                                                     = "pf3_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_vsecras_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_acs_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_ats_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_bar1_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_bar3_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_bar5_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_enable                                                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_acs_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_ats_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_msix_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_tph_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_virtio_en                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_msi_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_msix_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_pasid_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_prs_ext_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_ras_des_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sn_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_num_vf_non_ari                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar0_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar1_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar2_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar3_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar4_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar5_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_tph_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_user_vsec_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_user_vsec_offset                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_virtio_dev_specific_conf_en                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_virtio_en                                                                                     = "pf4_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_vsecras_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_acs_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_ats_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_bar1_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_bar3_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_bar5_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_enable                                                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_acs_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_ats_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_msix_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_tph_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_virtio_en                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_msi_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_msix_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_pasid_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_prs_ext_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_ras_des_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sn_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_num_vf_non_ari                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar0_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar1_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar2_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar3_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar4_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar5_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_tph_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_user_vsec_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_user_vsec_offset                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_virtio_dev_specific_conf_en                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_virtio_en                                                                                     = "pf5_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_vsecras_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_acs_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_ats_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_bar1_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_bar3_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_bar5_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_enable                                                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_acs_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_ats_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_msix_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_tph_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_virtio_en                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_msi_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_msix_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_pasid_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_prs_ext_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_ras_des_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sn_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_num_vf_non_ari                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar0_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar1_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar2_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar3_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar4_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar5_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_tph_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_user_vsec_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_user_vsec_offset                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_virtio_dev_specific_conf_en                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_virtio_en                                                                                     = "pf6_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_vsecras_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_acs_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_ats_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_bar1_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_bar3_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_bar5_mask_bit0                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_enable                                                                                        = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_acs_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_ats_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_msix_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_tph_cap_enable                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_virtio_en                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_msi_enable                                                                                    = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_msix_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_pasid_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_prs_ext_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_ras_des_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sn_cap_enable                                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_num_vf_non_ari                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar0_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar1_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar2_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar3_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar4_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar5_enabled                                                                         = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_tph_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_user_vsec_cap_enable                                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_user_vsec_offset                                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_virtio_dev_specific_conf_en                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_virtio_en                                                                                     = "pf7_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_vsecras_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_ptm_autoupdate                                                                                    = "autoupdate_10ms",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_addr_size0_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_pf_en0_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_start_addr0_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_addr_size1_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_pf_en1_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_start_addr1_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_addr_size2_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_pf_en2_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_start_addr2_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_addr_size3_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_pf_en3_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_start_addr3_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_addr_size4_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_pf_en4_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_start_addr4_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_addr_size5_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_pf_en5_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_start_addr5_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_addr_size6_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_pf_en6_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_start_addr6_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_addr_size7_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_pf_en7_attr                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_start_addr7_attr                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_fixedcred_attr                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_mcred_attr                                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_reloadcred_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_tlp_serr_dis_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_mmio_access_ctrl_grant_attr                                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_opcode_ctrl_lock_attr                                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_compressed_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_encrypted_attr                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_devbrd_type_attr                                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_vsec_next_offset_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_cvp_irq_en_attr                                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_gpio_irq_attr                                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid0_k_jtag_id_0_attr                                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid1_k_jtag_id_1_attr                                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid2_k_jtag_id_2_attr                                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid3_k_jtag_id_3_attr                                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_dfd_en_attr                                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_patcntr_en_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_0_attr                                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_1_attr                                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_2_attr                                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_3_attr                                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_trig_sel_0_attr                                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_trig_sel_1_attr                                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_0_attr                                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_1_attr                                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_2_attr                                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_3_attr                                                                                         = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr                                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_crs_en_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_rx_lane_flip_en_attr                                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_sris_mode_attr                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_tx_lane_flip_en_attr                                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_ehp_ctrl0_k_ehp_control_reg_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_outstanding_crd_attr                                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_tx_rd_th_attr                                                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cvp_cfg_err_en_attr                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dbi_access_err_en_attr                                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr                                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr                                                                   = "false",

parameter [1:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_sd_eq_control1_reg_eval_interval_time = 0,
parameter [31:0] hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_multi_lane_control_off_upconfigure_support = "true",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                                                     = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                                                          = 8,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                                                          = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req                                                              = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_prefetch                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_type                                                                                      = "pf0_bar0_mem64",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar1_reg_bar1_prefetch                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_prefetch                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_type                                                                                      = "pf0_bar2_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_mem_io                                                                                    = "pf0_bar3_mem",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_prefetch                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_prefetch                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_type                                                                                      = "pf0_bar4_mem32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask                                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar5_reg_bar5_prefetch                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bist_header_type_latency_cache_line_size_reg_multi_func                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_aux_curr                                                                             = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_dsi                                                                                  = "pf0_not_required",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_pme_support                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_reg_ari_acs_fun_grp_cap                                                                             = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_base_class_code                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_program_interface                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_revision_id                                                                      = 1,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_subclass_code                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_con_status_reg_no_soft_rst                                                                              = "pf0_not_internally_reset",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                                                   = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                                                    = 7,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ext_tag_supp                                                           = "pf0_supported",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap                                                                = "pf0_not_capable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id                                                             = 4466,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id                                                             = 32902,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled                                                                    = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_mask                                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en                                                                    = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_config_phy_tx_change                                                                      = "pf0_full_swing",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_select_deemph_var_mux                                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_selectable_deemph_bit_mux                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_support_mod_ts                                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable                                                            = "pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4                                                       = "gen4_pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5                                                       = "gen5_pf0_continue",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode                                                           = "pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4                                                      = "gen4_pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5                                                      = "gen5_pf0_next_rec_equal",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec                                                                = 2047,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4                                                           = 927,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5                                                           = 927,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable                                                      = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4                                                 = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5                                                 = "enable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg4                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg5                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo                                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg4                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg5                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts                                                                     = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4                                                                = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5                                                                = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_l1_2                                                                           = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_power_off                                                                      = 2,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_comm_mode_support                                                                  = 10,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_scale_support                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_value_support                                                               = 5,

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_aspm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_aspm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support = "true",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_aspm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_aspm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_1sub_cap_enable = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_2sub_cap_enable = "disable",

parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_sca                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_val                                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_t_common_mode                                                                        = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency                                                         = 3,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency                                                          = 4,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_port_num                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis                                                  = "pf0_minus_6db",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control                                      = "pf0_aspm_dis",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin                                          = "pf0_inta",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_misc_control_1_off_port_logic_wr_disable                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset                                                                 = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_bir                                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_table_offset                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported                                                        = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width                                                                     = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported                                                           = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                                                    = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                                                   = "pf0_msi_vec_1",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                       = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp                                                = "pf0_not_implemented",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pipe_loopback_control_off_pipe_loopback                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3                                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_capability_reg_no_eq_needed_support                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rsvdp_11                                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precode_req                                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precoding_on                                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_port_force_off_support_part_lanes_rxei_exit                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_port_link_ctrl_off_fast_link_mode                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility                                           = "true",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                   = "pf0_not_in_msix_table_vf",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec                                                          = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator                                                          = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3                                                               = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                                                      = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                                                   = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                                                          = "pf0_not_in_msix_table",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_device_spec                                                                 = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pfvf_sel_vsec_enable_attr                                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_phy_rxelecidle_k_rxelecidle_disable_attr                                                                    = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_phy_rxtermination_k_rxtermination_attr                                                                      = 127,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_err_en_correct_err_en_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_err_en_fatal_err_en_attr                                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_err_en_nonfatal_err_en_attr                                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr                                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_bw_mgt_int_en_attr                                                                            = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_eq_req_int_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_pme_int_en_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_int_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_pme_en_attr                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_inta_en_attr                                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_intb_en_attr                                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_intc_en_attr                                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_intd_en_attr                                                                                      = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_dlycnt_attr                                                                          = 6,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_mode_attr                                                                            = 5,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr                                                                   = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr                                                                = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr                                                     = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr                                                              = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_dllp_err_sts_attr                                                                       = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_tlp_err_sts_attr                                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_corrected_internal_err_sts_attr                                                             = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_dl_protocol_err_sts_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_ecrc_err_sts_attr                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_fc_protocol_err_sts_attr                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_mlf_tlp_err_sts_attr                                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_err_sts_attr                                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_overflow_err_sts_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_number_rollover_err_sts_attr                                                         = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_timer_timeout_err_sts_attr                                                           = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_surprise_down_err_sts_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_uncor_internal_err_sts_attr                                                                 = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tx_common_mode_k_txcommonmode_disable_attr                                                                  = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr                                                             = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr                                                          = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr                                                            = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr                                                              = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr                                                           = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr                                                = 0,
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cfg_update_en_attr                                                                        = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cii_en_attr                                                                               = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_cvp_mode                                                                                            = "cvp_disabled",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_drop_vendor0_msg                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_drop_vendor1_msg                                                                                    = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_ep_native                                                                                           = "native",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_maxpayload_size                                                                                     = "max_payload_128",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_num_of_lanes                                                                                        = "num_4",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_acs_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_ats_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_bar1_mask_bit0                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_bar3_mask_bit0                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_bar5_mask_bit0                                                                                  = "false",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_dlink_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_acs_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_ats_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_msix_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_tph_cap_enable                                                                             = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_io_decode                                                                                       = "io32",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_ltr_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_msi_enable                                                                                      = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_msix_enable                                                                                     = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_pasid_cap_enable                                                                                = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_prefetch_decode                                                                                 = "pref64",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_prs_ext_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_ras_des_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_sn_cap_enable                                                                                   = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_tph_cap_enable                                                                                  = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_user_vsec_cap_enable                                                                            = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_dev_specific_conf_en                                                                     = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_en                                                                                       = "pf0_virtio_disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_vsecras_cap_enable                                                                              = "disable",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_ptm_autoupdate                                                                                      = "autoupdate_10ms",
parameter hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr                                                           = "false",
parameter hssi_ctr_u_pcie_top_sim_mode                                                                                                                                           = "disable",
parameter hssi_ctr_u_pcie_top_sup_mode                                                                                                                                           = "user_mode",
parameter hssi_ctr_u_pcie_top_virtual_dmwr_support                                                                                                                               = "false",
parameter hssi_ctr_u_pcie_top_virtual_l1sub_support                                                                                                                              = "false",
parameter hssi_ctr_u_phy_top_pcie_capable_octet0                                                                                                                                 = "octet0_gen5_capable",
parameter hssi_ctr_u_phy_top_pcie_capable_octet1                                                                                                                                 = "octet1_gen5_capable",
parameter hssi_ctr_u_phy_top_u_phy_octet0_powerdown_mode                                                                                                                         = "true",
parameter hssi_ctr_u_phy_top_u_phy_octet1_powerdown_mode                                                                                                                         = "true",
parameter hssi_ctr_u_rnr_aibaux_top_wrp_powerdown_mode                                                                                                                           = "true",
parameter hssi_aib_ssm_silicon_rev                                                                                                                                               = "UNUSED",
parameter hssi_aibnd_rx_0_silicon_rev                                                                                                                                            = "UNUSED",
parameter hssi_aibnd_rx_13_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_aibnd_rx_15_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_aibnd_rx_23_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_aibnd_tx_0_silicon_rev                                                                                                                                            = "UNUSED",
parameter hssi_aibnd_tx_13_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_aibnd_tx_15_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_aibnd_tx_23_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_avmm1_if_0_silicon_rev                                                                                                                                            = "UNUSED",
parameter hssi_avmm1_if_13_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_avmm1_if_15_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_avmm1_if_23_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_avmm2_if_0_silicon_rev                                                                                                                                            = "UNUSED",
parameter hssi_avmm2_if_13_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_avmm2_if_15_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_avmm2_if_23_silicon_rev                                                                                                                                           = "UNUSED",
parameter hssi_pldadapt_rx_0_silicon_rev                                                                                                                                         = "UNUSED",
parameter hssi_pldadapt_rx_13_silicon_rev                                                                                                                                        = "UNUSED",
parameter hssi_pldadapt_rx_15_silicon_rev                                                                                                                                        = "UNUSED",
parameter hssi_pldadapt_rx_23_silicon_rev                                                                                                                                        = "UNUSED",
parameter hssi_pldadapt_tx_0_silicon_rev                                                                                                                                         = "UNUSED",
parameter hssi_pldadapt_tx_13_silicon_rev                                                                                                                                        = "UNUSED",
parameter hssi_pldadapt_tx_15_silicon_rev                                                                                                                                        = "UNUSED",
parameter hssi_pldadapt_tx_23_silicon_rev                                                                                                                                        = "UNUSED" 
)
(// TOP_PORTS_HERE
   // Clocks
   output wire         coreclkout_hip,                //      coreclkout_hip.clk, Check User Guide for details
   output wire         side_clk,                //      side_clk, Check User Guide for details
   input  wire         refclk0,                       //             refclk0.clk, Check User Guide for details
   input  wire         refclk1,                       //             refclk1.clk, Check User Guide for details
   // Resets
   input  wire         pin_perst_n,                   //   i pin_perst.pin_perst, Check User Guide for details
   input  wire         ninit_done,                    //   ninit_done.ninit_done, Its a Init_done signal should be connected to Reset release IP
   output wire         p0_reset_status_n,
   // P0 Avalon-ST RX Interface 
   input  wire         p0_rx_st_ready_i,                                    //PORT_NAME_CHANGE p0_rx_st_ready
   output wire         p0_rx_st_par_err_o,                                  //PORT_NAME_CHANGE p0_rx_st_par_err
   // P0 Avalon-ST0 RX Interface 
   output wire [255:0] p0_rx_st0_data_o,                                    //PORT_NAME_CHANGE p0_rx_st0_data
   output wire [127:0] p0_rx_st0_hdr_o,                                     //PORT_NAME_CHANGE p0_rx_st0_hdr
   output wire [31:0]  p0_rx_st0_prefix_o,                                  //PORT_NAME_CHANGE p0_rx_st0_prefix
   output wire         p0_rx_st0_sop_o,                                     //PORT_NAME_CHANGE p0_rx_st0_sop
   output wire         p0_rx_st0_eop_o,                                     //PORT_NAME_CHANGE p0_rx_st0_eop
   output wire         p0_rx_st0_dvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st0_dvalid
   output wire         p0_rx_st0_hvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st0_hvalid
   output wire [1:0]   p0_rx_st0_pvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st0_pvalid
   output wire [7:0]   p0_rx_st0_data_par_o,                                //PORT_NAME_CHANGE p0_rx_st0_data_par
   output wire [3:0]   p0_rx_st0_hdr_par_o,                                 //PORT_NAME_CHANGE p0_rx_st0_hdr_par
   output wire         p0_rx_st0_prefix_par_o,                              //PORT_NAME_CHANGE p0_rx_st0_prefix_par
   output wire         p0_rx_st0_passthrough_o,                             //PORT_NAME_CHANGE p0_rx_st0_passthrough
   output wire [2:0]   p0_rx_st0_bar_o,                                     //PORT_NAME_CHANGE p0_rx_st0_bar
   output wire         p0_rx_st0_vfactive_o,                                //PORT_NAME_CHANGE p0_rx_st0_vfactive
   output wire [10:0]  p0_rx_st0_vfnum_o,                                   //PORT_NAME_CHANGE p0_rx_st0_vfnum
   output wire [2:0]   p0_rx_st0_pfnum_o,                                   //PORT_NAME_CHANGE p0_rx_st0_pfnum
   output wire [11:0]  p0_rx_st0_rssai_prefix_o,                            //PORT_NAME_CHANGE p0_rx_st0_rssai_prefix
   output wire         p0_rx_st0_rssai_prefix_par_o,                        //PORT_NAME_CHANGE p0_rx_st0_rssai_prefix_par
   output wire         p0_rx_st0_misc_par_o,                                //PORT_NAME_CHANGE p0_rx_st0_misc_par
   output wire [2:0]   p0_rx_st0_empty_o,                                   //PORT_NAME_CHANGE p0_rx_st0_empty
   // P0 Avalon-ST1 RX Interface 
   output wire [255:0] p0_rx_st1_data_o,                                    //PORT_NAME_CHANGE p0_rx_st1_data
   output wire [127:0] p0_rx_st1_hdr_o,                                     //PORT_NAME_CHANGE p0_rx_st1_hdr
   output wire [31:0]  p0_rx_st1_prefix_o,                                  //PORT_NAME_CHANGE p0_rx_st1_prefix
   output wire         p0_rx_st1_sop_o,                                     //PORT_NAME_CHANGE p0_rx_st1_sop
   output wire         p0_rx_st1_eop_o,                                     //PORT_NAME_CHANGE p0_rx_st1_eop
   output wire         p0_rx_st1_dvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st1_dvalid
   output wire         p0_rx_st1_hvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st1_hvalid
   output wire [1:0]   p0_rx_st1_pvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st1_pvalid
   output wire [7:0]   p0_rx_st1_data_par_o,                                //PORT_NAME_CHANGE p0_rx_st1_data_par
   output wire [3:0]   p0_rx_st1_hdr_par_o,                                 //PORT_NAME_CHANGE p0_rx_st1_hdr_par
   output wire         p0_rx_st1_prefix_par_o,                              //PORT_NAME_CHANGE p0_rx_st1_prefix_par
   output wire         p0_rx_st1_passthrough_o,                             //PORT_NAME_CHANGE p0_rx_st1_passthrough
   output wire [2:0]   p0_rx_st1_bar_o,                                     //PORT_NAME_CHANGE p0_rx_st1_bar
   output wire         p0_rx_st1_vfactive_o,                                //PORT_NAME_CHANGE p0_rx_st1_vfactive
   output wire [10:0]  p0_rx_st1_vfnum_o,                                   //PORT_NAME_CHANGE p0_rx_st1_vfnum
   output wire [2:0]   p0_rx_st1_pfnum_o,                                   //PORT_NAME_CHANGE p0_rx_st1_pfnum
   output wire [11:0]  p0_rx_st1_rssai_prefix_o,                            //PORT_NAME_CHANGE p0_rx_st1_rssai_prefix
   output wire         p0_rx_st1_rssai_prefix_par_o,                        //PORT_NAME_CHANGE p0_rx_st1_rssai_prefix_par
   output wire         p0_rx_st1_misc_par_o,                                //PORT_NAME_CHANGE p0_rx_st1_misc_par
   output wire [2:0]   p0_rx_st1_empty_o,                                   //PORT_NAME_CHANGE p0_rx_st1_empty
   // P0 Avalon-ST2 RX Interface 
   output wire [255:0] p0_rx_st2_data_o,                                    //PORT_NAME_CHANGE p0_rx_st2_data
   output wire [127:0] p0_rx_st2_hdr_o,                                     //PORT_NAME_CHANGE p0_rx_st2_hdr
   output wire [31:0]  p0_rx_st2_prefix_o,                                  //PORT_NAME_CHANGE p0_rx_st2_prefix
   output wire         p0_rx_st2_sop_o,                                     //PORT_NAME_CHANGE p0_rx_st2_sop
   output wire         p0_rx_st2_eop_o,                                     //PORT_NAME_CHANGE p0_rx_st2_eop
   output wire         p0_rx_st2_dvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st2_dvalid
   output wire         p0_rx_st2_hvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st2_hvalid
   output wire [1:0]   p0_rx_st2_pvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st2_pvalid
   output wire [7:0]   p0_rx_st2_data_par_o,                                //PORT_NAME_CHANGE p0_rx_st2_data_par
   output wire [3:0]   p0_rx_st2_hdr_par_o,                                 //PORT_NAME_CHANGE p0_rx_st2_hdr_par
   output wire         p0_rx_st2_prefix_par_o,                              //PORT_NAME_CHANGE p0_rx_st2_prefix_par
   output wire         p0_rx_st2_passthrough_o,                             //PORT_NAME_CHANGE p0_rx_st2_passthrough
   output wire [2:0]   p0_rx_st2_bar_o,                                     //PORT_NAME_CHANGE p0_rx_st2_bar
   output wire         p0_rx_st2_vfactive_o,                                //PORT_NAME_CHANGE p0_rx_st2_vfactive
   output wire [10:0]  p0_rx_st2_vfnum_o,                                   //PORT_NAME_CHANGE p0_rx_st2_vfnum
   output wire [2:0]   p0_rx_st2_pfnum_o,                                   //PORT_NAME_CHANGE p0_rx_st2_pfnum
   output wire [11:0]  p0_rx_st2_rssai_prefix_o,                            //PORT_NAME_CHANGE p0_rx_st2_rssai_prefix
   output wire         p0_rx_st2_rssai_prefix_par_o,                        //PORT_NAME_CHANGE p0_rx_st2_rssai_prefix_par
   output wire         p0_rx_st2_misc_par_o,                                //PORT_NAME_CHANGE p0_rx_st2_misc_par
   output wire [2:0]   p0_rx_st2_empty_o,                                   //PORT_NAME_CHANGE p0_rx_st2_empty
   // P0 Avalon-ST3 RX Interface 
   output wire [255:0] p0_rx_st3_data_o,                                    //PORT_NAME_CHANGE p0_rx_st3_data
   output wire [127:0] p0_rx_st3_hdr_o,                                     //PORT_NAME_CHANGE p0_rx_st3_hdr
   output wire [31:0]  p0_rx_st3_prefix_o,                                  //PORT_NAME_CHANGE p0_rx_st3_prefix
   output wire         p0_rx_st3_sop_o,                                     //PORT_NAME_CHANGE p0_rx_st3_sop
   output wire         p0_rx_st3_eop_o,                                     //PORT_NAME_CHANGE p0_rx_st3_eop
   output wire         p0_rx_st3_dvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st3_dvalid
   output wire         p0_rx_st3_hvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st3_hvalid
   output wire [1:0]   p0_rx_st3_pvalid_o,                                  //PORT_NAME_CHANGE p0_rx_st3_pvalid
   output wire [7:0]   p0_rx_st3_data_par_o,                                //PORT_NAME_CHANGE p0_rx_st3_data_par
   output wire [3:0]   p0_rx_st3_hdr_par_o,                                 //PORT_NAME_CHANGE p0_rx_st3_hdr_par
   output wire         p0_rx_st3_prefix_par_o,                              //PORT_NAME_CHANGE p0_rx_st3_prefix_par
   output wire         p0_rx_st3_passthrough_o,                             //PORT_NAME_CHANGE p0_rx_st3_passthrough
   output wire [2:0]   p0_rx_st3_bar_o,                                     //PORT_NAME_CHANGE p0_rx_st3_bar
   output wire         p0_rx_st3_vfactive_o,                                //PORT_NAME_CHANGE p0_rx_st3_vfactive
   output wire [10:0]  p0_rx_st3_vfnum_o,                                   //PORT_NAME_CHANGE p0_rx_st3_vfnum
   output wire [2:0]   p0_rx_st3_pfnum_o,                                   //PORT_NAME_CHANGE p0_rx_st3_pfnum
   output wire [11:0]  p0_rx_st3_rssai_prefix_o,                            //PORT_NAME_CHANGE p0_rx_st3_rssai_prefix
   output wire         p0_rx_st3_rssai_prefix_par_o,                        //PORT_NAME_CHANGE p0_rx_st3_rssai_prefix_par
   output wire         p0_rx_st3_misc_par_o,                                //PORT_NAME_CHANGE p0_rx_st3_misc_par
   output wire [2:0]   p0_rx_st3_empty_o,                                   //PORT_NAME_CHANGE p0_rx_st3_empty
   // P0 Avalon-ST RX Credit Interface 
   input  wire [2:0]   p0_rx_st_hcrd_ch_i,                                  //PORT_NAME_CHANGE p0_rx_st_Hcrd_ch
   input  wire [2:0]   p0_rx_st_hcrd_init_i,                                //PORT_NAME_CHANGE p0_rx_st_Hcrd_init
   input  wire [2:0]   p0_rx_st_hcrd_update_i,                              //PORT_NAME_CHANGE p0_rx_st_Hcrd_update
   input  wire [5:0]   p0_rx_st_hcrd_update_cnt_i,                          //PORT_NAME_CHANGE p0_rx_st_Hcrd_update_cnt
   output wire [2:0]   p0_rx_st_hcrd_init_ack_o,                            //PORT_NAME_CHANGE p0_rx_st_Hcrd_init_ack
   input  wire [2:0]   p0_rx_st_dcrd_ch_i,                                  //PORT_NAME_CHANGE p0_rx_st_Dcrd_ch
   input  wire [2:0]   p0_rx_st_dcrd_init_i,                                //PORT_NAME_CHANGE p0_rx_st_Dcrd_init
   input  wire [2:0]   p0_rx_st_dcrd_update_i,                              //PORT_NAME_CHANGE p0_rx_st_Dcrd_update
   input  wire [11:0]  p0_rx_st_dcrd_update_cnt_i,                          //PORT_NAME_CHANGE p0_rx_st_Dcrd_update_cnt
   output wire [2:0]   p0_rx_st_dcrd_init_ack_o,                            //PORT_NAME_CHANGE p0_rx_st_Dcrd_init_ack
   // Avalon-ST0 TX Credit Interface 
   output wire [2:0]   p0_tx_st_hcrd_ch_o,                                  //PORT_NAME_CHANGE p0_tx_st_Hcrd_ch
   output wire [2:0]   p0_tx_st_hcrd_init_o,                                //PORT_NAME_CHANGE p0_tx_st_Hcrd_init
   output wire [2:0]   p0_tx_st_hcrd_update_o,                              //PORT_NAME_CHANGE p0_tx_st_Hcrd_update
   output wire [5:0]   p0_tx_st_hcrd_update_cnt_o,                          //PORT_NAME_CHANGE p0_tx_st_Hcrd_update_cnt
   input  wire [2:0]   p0_tx_st_hcrd_init_ack_i,                            //PORT_NAME_CHANGE p0_tx_st_Hcrd_init_ack
   output wire [2:0]   p0_tx_st_dcrd_ch_o,                                  //PORT_NAME_CHANGE p0_tx_st_Dcrd_ch
   output wire [2:0]   p0_tx_st_dcrd_init_o,                                //PORT_NAME_CHANGE p0_tx_st_Dcrd_init
   output wire [2:0]   p0_tx_st_dcrd_update_o,                              //PORT_NAME_CHANGE p0_tx_st_Dcrd_update
   output wire [11:0]  p0_tx_st_dcrd_update_cnt_o,                          //PORT_NAME_CHANGE p0_tx_st_Dcrd_update_cnt
   input  wire [2:0]   p0_tx_st_dcrd_init_ack_i,                            //PORT_NAME_CHANGE p0_tx_st_Dcrd_init_ack
   // Avalon-ST TX Interface 
   output wire         p0_tx_st_ready_o,                                    //PORT_NAME_CHANGE p0_tx_st_ready
   output wire         p0_tx_st_par_err_o,                                  //PORT_NAME_CHANGE p0_tx_st_par_err        // Not Implemented
   // Avalon-ST0 TX Interface 
   input  wire [255:0] p0_tx_st0_data_i,                                    //PORT_NAME_CHANGE p0_tx_st0_data
   input  wire [127:0] p0_tx_st0_hdr_i,                                     //PORT_NAME_CHANGE p0_tx_st0_hdr
   input  wire [31:0]  p0_tx_st0_prefix_i,                                  //PORT_NAME_CHANGE p0_tx_st0_prefix
   input  wire         p0_tx_st0_sop_i,                                     //PORT_NAME_CHANGE p0_tx_st0_sop
   input  wire         p0_tx_st0_eop_i,                                     //PORT_NAME_CHANGE p0_tx_st0_eop
   input  wire         p0_tx_st0_dvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st0_dvalid
   input  wire         p0_tx_st0_hvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st0_hvalid
   input  wire [1:0]   p0_tx_st0_pvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st0_pvalid
   input  wire         p0_tx_st0_passthrough_i,                             //PORT_NAME_CHANGE p0_tx_st0_passthrough
   input  wire [7:0]   p0_tx_st0_data_par_i,                                //PORT_NAME_CHANGE p0_tx_st0_data_par
   input  wire [3:0]   p0_tx_st0_hdr_par_i,                                 //PORT_NAME_CHANGE p0_tx_st0_hdr_par
   input  wire         p0_tx_st0_prefix_par_i,                              //PORT_NAME_CHANGE p0_tx_st0_prefix_par
   input  wire [2:0]   p0_tx_st0_empty_i,                                   //PORT_NAME_CHANGE p0_tx_st0_empty
   input  wire [11:0]  p0_tx_st0_rssai_prefix_i,                            //PORT_NAME_CHANGE p0_tx_st0_rssai_prefix
   input  wire         p0_tx_st0_rssai_prefix_par_i,                        //PORT_NAME_CHANGE p0_tx_st0_rssai_prefix_par
   // Avalon-ST1 TX Interface 
   input  wire [255:0] p0_tx_st1_data_i,                                    //PORT_NAME_CHANGE p0_tx_st1_data
   input  wire [127:0] p0_tx_st1_hdr_i,                                     //PORT_NAME_CHANGE p0_tx_st1_hdr
   input  wire [31:0]  p0_tx_st1_prefix_i,                                  //PORT_NAME_CHANGE p0_tx_st1_prefix
   input  wire         p0_tx_st1_sop_i,                                     //PORT_NAME_CHANGE p0_tx_st1_sop
   input  wire         p0_tx_st1_eop_i,                                     //PORT_NAME_CHANGE p0_tx_st1_eop
   input  wire         p0_tx_st1_dvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st1_dvalid
   input  wire         p0_tx_st1_hvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st1_hvalid
   input  wire [1:0]   p0_tx_st1_pvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st1_pvalid
   input  wire         p0_tx_st1_passthrough_i,                             //PORT_NAME_CHANGE p0_tx_st1_passthrough
   input  wire [7:0]   p0_tx_st1_data_par_i,                                //PORT_NAME_CHANGE p0_tx_st1_data_par
   input  wire [3:0]   p0_tx_st1_hdr_par_i,                                 //PORT_NAME_CHANGE p0_tx_st1_hdr_par
   input  wire         p0_tx_st1_prefix_par_i,                              //PORT_NAME_CHANGE p0_tx_st1_prefix_par
   input  wire [2:0]   p0_tx_st1_empty_i,                                   //PORT_NAME_CHANGE p0_tx_st1_empty
   input  wire [11:0]  p0_tx_st1_rssai_prefix_i,                            //PORT_NAME_CHANGE p0_tx_st1_rssai_prefix
   input  wire         p0_tx_st1_rssai_prefix_par_i,                        //PORT_NAME_CHANGE p0_tx_st1_rssai_prefix_par
   // Avalon-ST2 TX Interface 
   input  wire [255:0] p0_tx_st2_data_i,                                    //PORT_NAME_CHANGE p0_tx_st2_data
   input  wire [127:0] p0_tx_st2_hdr_i,                                     //PORT_NAME_CHANGE p0_tx_st2_hdr
   input  wire [31:0]  p0_tx_st2_prefix_i,                                  //PORT_NAME_CHANGE p0_tx_st2_prefix
   input  wire         p0_tx_st2_sop_i,                                     //PORT_NAME_CHANGE p0_tx_st2_sop
   input  wire         p0_tx_st2_eop_i,                                     //PORT_NAME_CHANGE p0_tx_st2_eop
   input  wire         p0_tx_st2_dvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st2_dvalid
   input  wire         p0_tx_st2_hvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st2_hvalid
   input  wire [1:0]   p0_tx_st2_pvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st2_pvalid
   input  wire         p0_tx_st2_passthrough_i,                             //PORT_NAME_CHANGE p0_tx_st2_passthrough
   input  wire [7:0]   p0_tx_st2_data_par_i,                                //PORT_NAME_CHANGE p0_tx_st2_data_par
   input  wire [3:0]   p0_tx_st2_hdr_par_i,                                 //PORT_NAME_CHANGE p0_tx_st2_hdr_par
   input  wire         p0_tx_st2_prefix_par_i,                              //PORT_NAME_CHANGE p0_tx_st2_prefix_par
   input  wire [2:0]   p0_tx_st2_empty_i,                                   //PORT_NAME_CHANGE p0_tx_st2_empty
   input  wire [11:0]  p0_tx_st2_rssai_prefix_i,                            //PORT_NAME_CHANGE p0_tx_st2_rssai_prefix
   input  wire         p0_tx_st2_rssai_prefix_par_i,                        //PORT_NAME_CHANGE p0_tx_st2_rssai_prefix_par
   // Avalon-ST3 TX Interface 
   input  wire [255:0] p0_tx_st3_data_i,                                    //PORT_NAME_CHANGE p0_tx_st3_data
   input  wire [127:0] p0_tx_st3_hdr_i,                                     //PORT_NAME_CHANGE p0_tx_st3_hdr
   input  wire [31:0]  p0_tx_st3_prefix_i,                                  //PORT_NAME_CHANGE p0_tx_st3_prefix
   input  wire         p0_tx_st3_sop_i,                                     //PORT_NAME_CHANGE p0_tx_st3_sop
   input  wire         p0_tx_st3_eop_i,                                     //PORT_NAME_CHANGE p0_tx_st3_eop
   input  wire         p0_tx_st3_dvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st3_dvalid
   input  wire         p0_tx_st3_hvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st3_hvalid
   input  wire [1:0]   p0_tx_st3_pvalid_i,                                  //PORT_NAME_CHANGE p0_tx_st3_pvalid
   input  wire         p0_tx_st3_passthrough_i,                             //PORT_NAME_CHANGE p0_tx_st3_passthrough
   input  wire [7:0]   p0_tx_st3_data_par_i,                                //PORT_NAME_CHANGE p0_tx_st3_data_par
   input  wire [3:0]   p0_tx_st3_hdr_par_i,                                 //PORT_NAME_CHANGE p0_tx_st3_hdr_par
   input  wire         p0_tx_st3_prefix_par_i,                              //PORT_NAME_CHANGE p0_tx_st3_prefix_par
   input  wire [2:0]   p0_tx_st3_empty_i,                                   //PORT_NAME_CHANGE p0_tx_st3_empty
   input  wire [11:0]  p0_tx_st3_rssai_prefix_i,                            //PORT_NAME_CHANGE p0_tx_st3_rssai_prefix
   input  wire         p0_tx_st3_rssai_prefix_par_i,                        //PORT_NAME_CHANGE p0_tx_st3_rssai_prefix_par
   // Hot Plug Interface
   input  wire         p0_sys_eml_interlock_engaged_i,                     //PORT_NAME_CHANGE sys_eml_interlock_engaged,
   input  wire         p0_sys_cmd_cpled_int_i,                             //PORT_NAME_CHANGE sys_cmd_cpled_int,
   input  wire         p0_sys_pwr_fault_det_i,                             //PORT_NAME_CHANGE sys_pwr_fault_det,
   input  wire         p0_sys_mrl_sensor_state_i,                          //PORT_NAME_CHANGE sys_mrl_sensor_state,
   input  wire         p0_sys_pre_det_state_i,                             //PORT_NAME_CHANGE sys_pre_det_state,
   input  wire         p0_sys_atten_button_pressed_i,                      //PORT_NAME_CHANGE sys_atten_button_pressed,
   input  wire         p0_sys_aux_pwr_det_i,                               //PORT_NAME_CHANGE sys_aux_pwr_det,
   // Hard IP Status Interface
   output wire         p0_link_up_o,                                       //PORT_NAME_CHANGE p0_link_up,
   output wire         p0_dl_up_o,                                         //PORT_NAME_CHANGE p0_dl_up,
   // Power Management
   output wire [7:0]   p0_pm_curnt_state_o,                                //PORT_NAME_CHANGE p0_pm_curnt_state,
   output wire [31:0]  p0_pm_dstate_o,                                     //PORT_NAME_CHANGE p0_pm_dstate,
   input  wire         p0_app_init_rst_i,                                  //PORT_NAME_CHANGE p0_app_init_rst,
   input  wire [7:0]   p0_app_req_retry_en_i,                              //PORT_NAME_CHANGE p0_app_req_retry_en,
   input  wire         p0_app_xfer_pending_i,                              //PORT_NAME_CHANGE p0_app_xfer_pending,
   // CXL.mem and CXL.Cache RX
   // union
   //output cxl_cache_mem_rx_intf  cxl_cache_mem_rx_frame0, // inlcude 3-bit Prot ID
   //output cxl_cache_mem_rx_intf  cxl_cache_mem_rx_frame1, // include 3-bit Prot ID
   //interfaces_cxl_mem_rx
   output wire [3-1:0]     frame0_cxl_mem_port_id_o,
   output wire [1-1:0]     frame0_cxl_mem_m2s_rwd0_valid_o,
   output wire [1-1:0]     frame0_cxl_mem_m2s_rwd0_poison_o,
   output wire [4-1:0]     frame0_cxl_mem_m2s_rwd0_beparity_o,
   output wire [8-1:0]     frame0_cxl_mem_m2s_rwd0_dataparity_o,
   output wire [4-1:0]     frame0_cxl_mem_m2s_rwd0_memopcode_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_rwd0_metafield_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_rwd0_metavalue_o,
   output wire [3-1:0]     frame0_cxl_mem_m2s_rwd0_snptype_o,
   output wire [16-1:0]    frame0_cxl_mem_m2s_rwd0_tag_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_rwd0_tc_o,
   output wire [1-1:0]     frame0_cxl_mem_m2s_req1_valid_o,
   output wire [4-1:0]     frame0_cxl_mem_m2s_req1_memopcode_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_req1_metafield_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_req1_metavalue_o,
   output wire [3-1:0]     frame0_cxl_mem_m2s_req1_snptype_o,
   output wire [16-1:0]    frame0_cxl_mem_m2s_req1_tag_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_req1_tc_o,
   output wire [5-1:0]     frame0_cxl_mem_m2s_req1_rsvd_h_o,
   output wire [47-1:0]    frame0_cxl_mem_m2s_req1_address_o,
   output wire [5-1:0]     frame0_cxl_mem_m2s_req1_rsvd_l_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_req1_parity_o,
   output wire [3-1:0]     frame0_cxl_mem_not_mapped_2_o,
   output wire [1-1:0]     frame0_cxl_mem_m2s_req0_valid_o,
   output wire [4-1:0]     frame0_cxl_mem_m2s_req0_memopcode_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_req0_metafield_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_req0_metavalue_o,
   output wire [3-1:0]     frame0_cxl_mem_m2s_req0_snptype_o,
   output wire [16-1:0]    frame0_cxl_mem_m2s_req0_tag_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_req0_tc_o,
   output wire [5-1:0]     frame0_cxl_mem_m2s_req0_rsvd_h_o,
   output wire [47-1:0]    frame0_cxl_mem_m2s_req0_address_o,
   output wire [5-1:0]     frame0_cxl_mem_m2s_req0_rsvd_l_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_req0_parity_o,
   output wire [5-1:0]     frame0_cxl_mem_m2s_rwd0_rsvd_h_o,
   output wire [46-1:0]    frame0_cxl_mem_m2s_rwd0_address_o,
   output wire [5-1:0]     frame0_cxl_mem_m2s_rwd0_rsvd_l_o,
   output wire [2-1:0]     frame0_cxl_mem_not_mapped_1_o,
   output wire [6-1:0]     frame0_cxl_mem_m2s_datahdr1_o,
   output wire [32-1:0]    frame0_cxl_mem_m2s_rwd0_byteen_h_o,
   output wire [256-1:0]   frame0_cxl_mem_m2s_rwd0_data_h_o,
   output wire [4-1:0]     frame0_cxl_mem_not_mapped_0_o,
   output wire [2-1:0]     frame0_cxl_mem_m2s_rwd0_hdrparity_o,
   output wire [32-1:0]    frame0_cxl_mem_m2s_rwd0_byteen_l_o,
   output wire [256-1:0]   frame0_cxl_mem_m2s_rwd0_data_l_o,
   output wire [3-1:0]     frame1_cxl_mem_port_id_o,
   output wire [1-1:0]     frame1_cxl_mem_m2s_rwd0_valid_o,
   output wire [1-1:0]     frame1_cxl_mem_m2s_rwd0_poison_o,
   output wire [4-1:0]     frame1_cxl_mem_m2s_rwd0_beparity_o,
   output wire [8-1:0]     frame1_cxl_mem_m2s_rwd0_dataparity_o,
   output wire [4-1:0]     frame1_cxl_mem_m2s_rwd0_memopcode_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_rwd0_metafield_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_rwd0_metavalue_o,
   output wire [3-1:0]     frame1_cxl_mem_m2s_rwd0_snptype_o,
   output wire [16-1:0]    frame1_cxl_mem_m2s_rwd0_tag_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_rwd0_tc_o,
   output wire [1-1:0]     frame1_cxl_mem_m2s_req1_valid_o,
   output wire [4-1:0]     frame1_cxl_mem_m2s_req1_memopcode_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_req1_metafield_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_req1_metavalue_o,
   output wire [3-1:0]     frame1_cxl_mem_m2s_req1_snptype_o,
   output wire [16-1:0]    frame1_cxl_mem_m2s_req1_tag_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_req1_tc_o,
   output wire [5-1:0]     frame1_cxl_mem_m2s_req1_rsvd_h_o,
   output wire [47-1:0]    frame1_cxl_mem_m2s_req1_address_o,
   output wire [5-1:0]     frame1_cxl_mem_m2s_req1_rsvd_l_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_req1_parity_o,
   output wire [3-1:0]     frame1_cxl_mem_not_mapped_2_o,
   output wire [1-1:0]     frame1_cxl_mem_m2s_req0_valid_o,
   output wire [4-1:0]     frame1_cxl_mem_m2s_req0_memopcode_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_req0_metafield_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_req0_metavalue_o,
   output wire [3-1:0]     frame1_cxl_mem_m2s_req0_snptype_o,
   output wire [16-1:0]    frame1_cxl_mem_m2s_req0_tag_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_req0_tc_o,
   output wire [5-1:0]     frame1_cxl_mem_m2s_req0_rsvd_h_o,
   output wire [47-1:0]    frame1_cxl_mem_m2s_req0_address_o,
   output wire [5-1:0]     frame1_cxl_mem_m2s_req0_rsvd_l_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_req0_parity_o,
   output wire [5-1:0]     frame1_cxl_mem_m2s_rwd0_rsvd_h_o,
   output wire [46-1:0]    frame1_cxl_mem_m2s_rwd0_address_o,
   output wire [5-1:0]     frame1_cxl_mem_m2s_rwd0_rsvd_l_o,
   output wire [2-1:0]     frame1_cxl_mem_not_mapped_1_o,
   output wire [6-1:0]     frame1_cxl_mem_m2s_datahdr1_o,
   output wire [32-1:0]    frame1_cxl_mem_m2s_rwd0_byteen_h_o,
   output wire [256-1:0]   frame1_cxl_mem_m2s_rwd0_data_h_o,
   output wire [4-1:0]     frame1_cxl_mem_not_mapped_0_o,
   output wire [2-1:0]     frame1_cxl_mem_m2s_rwd0_hdrparity_o,
   output wire [32-1:0]    frame1_cxl_mem_m2s_rwd0_byteen_l_o,
   output wire [256-1:0]   frame1_cxl_mem_m2s_rwd0_data_l_o,
   //interfaces_cxl_cache_rx
   output wire [2:0]       frame0_cxl_cache_port_id_o,
   output wire [29:7]      frame0_cxl_cache_not_mapped_2_o,
   output wire             frame0_cxl_cache_h2d_rsp3_valid_o,
   output wire             frame0_cxl_cache_h2d_rsp3_rsvd_o,
   output wire [1:0]       frame0_cxl_cache_h2d_rsp3_parity_o,
   output wire [1:0]       frame0_cxl_cache_h2d_rsp3_pre_o,
   output wire [3:0]       frame0_cxl_cache_h2d_rsp3_opcode_o,
   output wire [11:0]      frame0_cxl_cache_h2d_rsp3_cqid_o,
   output wire [11:0]      frame0_cxl_cache_h2d_rsp3_data_o,
   output wire [6:1]       frame0_cxl_cache_not_mapped_1_o,
   output wire [11:0]      frame0_cxl_cache_h2d_data1_cqid_o,
   output wire             frame0_cxl_cache_h2d_req1_valid_o,
   output wire [1:0]       frame0_cxl_cache_h2d_req1_rsvd_o,
   output wire [2:0]       frame0_cxl_cache_h2d_req1_opcode_o,
   output wire [1:0]       frame0_cxl_cache_h2d_req1_parity_o,
   output wire [11:0]      frame0_cxl_cache_h2d_req1_uqid_o,
   output wire [45:0]      frame0_cxl_cache_h2d_req1_address_o,
   output wire             frame0_cxl_cache_h2d_rsp2_valid_o,
   output wire             frame0_cxl_cache_h2d_rsp2_rsvd_o,
   output wire [1:0]       frame0_cxl_cache_h2d_rsp2_parity_o,
   output wire [1:0]       frame0_cxl_cache_h2d_rsp2_pre_o,
   output wire [3:0]       frame0_cxl_cache_h2d_rsp2_opcode_o,
   output wire [11:0]      frame0_cxl_cache_h2d_rsp2_cqid_o,
   output wire [11:0]      frame0_cxl_cache_h2d_rsp2_data_o,
   output wire             frame0_cxl_cache_h2d_req0_valid_o,
   output wire [1:0]       frame0_cxl_cache_h2d_req0_rsvd_o,
   output wire [2:0]       frame0_cxl_cache_h2d_req0_opcode_o,
   output wire [1:0]       frame0_cxl_cache_h2d_req0_parity_o,
   output wire [11:0]      frame0_cxl_cache_h2d_req0_uqid_o,
   output wire [45:0]      frame0_cxl_cache_h2d_req0_address_o,
   output wire [1:0]       frame0_cxl_cache_h2d_datahdr1_parity_o,
   output wire             frame0_cxl_cache_not_mapped_0_o,
   output wire             frame0_cxl_cache_h2d_rsp1_valid_o,
   output wire             frame0_cxl_cache_h2d_rsp1_rsvd_o,
   output wire [1:0]       frame0_cxl_cache_h2d_rsp1_parity_o,
   output wire [1:0]       frame0_cxl_cache_h2d_rsp1_pre_o,
   output wire [3:0]       frame0_cxl_cache_h2d_rsp1_opcode_o,
   output wire [11:0]      frame0_cxl_cache_h2d_rsp1_cqid_o,
   output wire [11:0]      frame0_cxl_cache_h2d_rsp1_data_o,
   output wire [7:0]       frame0_cxl_cache_h2d_data1_rsvd_o,
   output wire             frame0_cxl_cache_h2d_rsp0_valid_o,
   output wire             frame0_cxl_cache_h2d_rsp0_rsvd_o,
   output wire [1:0]       frame0_cxl_cache_h2d_rsp0_parity_o,
   output wire [1:0]       frame0_cxl_cache_h2d_rsp0_pre_o,
   output wire [3:0]       frame0_cxl_cache_h2d_rsp0_opcode_o,
   output wire [11:0]      frame0_cxl_cache_h2d_rsp0_cqid_o,
   output wire [11:0]      frame0_cxl_cache_h2d_rsp0_data_o,
   output wire [511:256]   frame0_cxl_cache_h2d_data0_data_h_o,
   output wire             frame0_cxl_cache_h2d_data1_valid_o,
   output wire             frame0_cxl_cache_h2d_data1_chunkvalid_o,
   output wire             frame0_cxl_cache_h2d_data0_valid_o,
   output wire             frame0_cxl_cache_h2d_data0_chunkvalid_o,
   output wire             frame0_cxl_cache_h2d_data0_poison_o,
   output wire             frame0_cxl_cache_h2d_data0_goerr_o,
   output wire [1:0]       frame0_cxl_cache_h2d_datahdr0_parity_o,
   output wire [7:0]       frame0_cxl_cache_h2d_data0_dataparity_o,
   output wire [7:0]       frame0_cxl_cache_h2d_data0_rsvd_o,
   output wire             frame0_cxl_cache_h2d_data1_poison_o,
   output wire             frame0_cxl_cache_h2d_data1_goerr_o,
   output wire [11:0]      frame0_cxl_cache_h2d_data0_cqid_o,
   output wire [255:0]     frame0_cxl_cache_h2d_data0_data_l_o,
   output wire [2:0]       frame1_cxl_cache_port_id_o,
   output wire [29:7]      frame1_cxl_cache_not_mapped_2_o,
   output wire             frame1_cxl_cache_h2d_rsp3_valid_o,
   output wire             frame1_cxl_cache_h2d_rsp3_rsvd_o,
   output wire [1:0]       frame1_cxl_cache_h2d_rsp3_parity_o,
   output wire [1:0]       frame1_cxl_cache_h2d_rsp3_pre_o,
   output wire [3:0]       frame1_cxl_cache_h2d_rsp3_opcode_o,
   output wire [11:0]      frame1_cxl_cache_h2d_rsp3_cqid_o,
   output wire [11:0]      frame1_cxl_cache_h2d_rsp3_data_o,
   output wire [6:1]       frame1_cxl_cache_not_mapped_1_o,
   output wire [11:0]      frame1_cxl_cache_h2d_data1_cqid_o,
   output wire             frame1_cxl_cache_h2d_req1_valid_o,
   output wire [1:0]       frame1_cxl_cache_h2d_req1_rsvd_o,
   output wire [2:0]       frame1_cxl_cache_h2d_req1_opcode_o,
   output wire [1:0]       frame1_cxl_cache_h2d_req1_parity_o,
   output wire [11:0]      frame1_cxl_cache_h2d_req1_uqid_o,
   output wire [45:0]      frame1_cxl_cache_h2d_req1_address_o,
   output wire             frame1_cxl_cache_h2d_rsp2_valid_o,
   output wire             frame1_cxl_cache_h2d_rsp2_rsvd_o,
   output wire [1:0]       frame1_cxl_cache_h2d_rsp2_parity_o,
   output wire [1:0]       frame1_cxl_cache_h2d_rsp2_pre_o,
   output wire [3:0]       frame1_cxl_cache_h2d_rsp2_opcode_o,
   output wire [11:0]      frame1_cxl_cache_h2d_rsp2_cqid_o,
   output wire [11:0]      frame1_cxl_cache_h2d_rsp2_data_o,
   output wire             frame1_cxl_cache_h2d_req0_valid_o,
   output wire [1:0]       frame1_cxl_cache_h2d_req0_rsvd_o,
   output wire [2:0]       frame1_cxl_cache_h2d_req0_opcode_o,
   output wire [1:0]       frame1_cxl_cache_h2d_req0_parity_o,
   output wire [11:0]      frame1_cxl_cache_h2d_req0_uqid_o,
   output wire [45:0]      frame1_cxl_cache_h2d_req0_address_o,
   output wire [1:0]       frame1_cxl_cache_h2d_datahdr1_parity_o,
   output wire             frame1_cxl_cache_not_mapped_0_o,
   output wire             frame1_cxl_cache_h2d_rsp1_valid_o,
   output wire             frame1_cxl_cache_h2d_rsp1_rsvd_o,
   output wire [1:0]       frame1_cxl_cache_h2d_rsp1_parity_o,
   output wire [1:0]       frame1_cxl_cache_h2d_rsp1_pre_o,
   output wire [3:0]       frame1_cxl_cache_h2d_rsp1_opcode_o,
   output wire [11:0]      frame1_cxl_cache_h2d_rsp1_cqid_o,
   output wire [11:0]      frame1_cxl_cache_h2d_rsp1_data_o,
   output wire [7:0]       frame1_cxl_cache_h2d_data1_rsvd_o,
   output wire             frame1_cxl_cache_h2d_rsp0_valid_o,
   output wire             frame1_cxl_cache_h2d_rsp0_rsvd_o,
   output wire [1:0]       frame1_cxl_cache_h2d_rsp0_parity_o,
   output wire [1:0]       frame1_cxl_cache_h2d_rsp0_pre_o,
   output wire [3:0]       frame1_cxl_cache_h2d_rsp0_opcode_o,
   output wire [11:0]      frame1_cxl_cache_h2d_rsp0_cqid_o,
   output wire [11:0]      frame1_cxl_cache_h2d_rsp0_data_o,
   output wire [511:256]   frame1_cxl_cache_h2d_data0_data_h_o,
   output wire             frame1_cxl_cache_h2d_data1_valid_o,
   output wire             frame1_cxl_cache_h2d_data1_chunkvalid_o,
   output wire             frame1_cxl_cache_h2d_data0_valid_o,
   output wire             frame1_cxl_cache_h2d_data0_chunkvalid_o,
   output wire             frame1_cxl_cache_h2d_data0_poison_o,
   output wire             frame1_cxl_cache_h2d_data0_goerr_o,
   output wire [1:0]       frame1_cxl_cache_h2d_datahdr0_parity_o,
   output wire [7:0]       frame1_cxl_cache_h2d_data0_dataparity_o,
   output wire [7:0]       frame1_cxl_cache_h2d_data0_rsvd_o,
   output wire             frame1_cxl_cache_h2d_data1_poison_o,
   output wire             frame1_cxl_cache_h2d_data1_goerr_o,
   output wire [11:0]      frame1_cxl_cache_h2d_data0_cqid_o,
   output wire [255:0]     frame1_cxl_cache_h2d_data0_data_l_o,

   // CXL.mem and CXL.Cache TX
   //input  cxl_mem_s2m_tx_intf          cxl_mem_s2m_tx_frame0, // no ProtID, 1 ready
   //input                               cxl_mem_s2m_tx_frame0_valid,
   //output                              cxl_mem_s2m_tx_frame0_ready,
   //input  cxl_mem_s2m_tx_intf          cxl_mem_s2m_tx_frame1, // no ProtID, 1 ready
   //input                               cxl_mem_s2m_tx_frame1_valid,
   //output                              cxl_mem_s2m_tx_frame1_ready,
   //interfaces_cxl_mem_s2m_tx
   input  wire [1:0]       frame0_cxl_mem_s2m_ndr1_devload_i,
   input  wire             frame0_cxl_mem_s2m_ndr1_valid_i,
   input  wire [2:0]       frame0_cxl_mem_s2m_ndr1_opcode_i,
   input  wire [1:0]       frame0_cxl_mem_s2m_ndr1_metafield_i,
   input  wire [1:0]       frame0_cxl_mem_s2m_ndr1_metavalue_i,
   input  wire [1:0]       frame0_cxl_mem_s2m_ndr1_parity_i,
   input  wire [3:0]       frame0_cxl_mem_s2m_ndr1_rsvd_i,
   input  wire [15:0]      frame0_cxl_mem_s2m_ndr1_tag_i,
   input  wire [1:0]       frame0_cxl_mem_s2m_ndr0_devload_i,
   input  wire             frame0_cxl_mem_s2m_ndr0_valid_i,
   input  wire [2:0]       frame0_cxl_mem_s2m_ndr0_opcode_i,
   input  wire [1:0]       frame0_cxl_mem_s2m_ndr0_metafield_i,
   input  wire [1:0]       frame0_cxl_mem_s2m_ndr0_metavalue_i,
   input  wire [1:0]       frame0_cxl_mem_s2m_ndr0_parity_i,
   input  wire [3:0]       frame0_cxl_mem_s2m_ndr0_rsvd_i,
   input  wire [15:0]      frame0_cxl_mem_s2m_ndr0_tag_i,
   input  wire [54:0]      frame0_cxl_mem_s2m_drs_hdr1_i,
   input  wire             frame0_cxl_mem_s2m_drs0_valid_i,
   input  wire             frame0_cxl_mem_s2m_drs0_poison_i,
   input  wire [2:0]       frame0_cxl_mem_s2m_drs0_opcode_i,
   input  wire [1:0]       frame0_cxl_mem_s2m_drs0_metafield_i,
   input  wire [1:0]       frame0_cxl_mem_s2m_drs0_metavalue_i,
   input  wire [14:0]      frame0_cxl_mem_s2m_drs0_rsvd_i,
   input  wire [8:0]       frame0_cxl_mem_s2m_drs0_rsvd_field1_i, // revb 
   input  wire [1:0]       frame0_cxl_mem_s2m_drs0_devload_i,
   input  wire [3:0]       frame0_cxl_mem_s2m_drs0_rsvd_field0_i,
   input  wire [1:0]       frame0_cxl_mem_s2m_drs0_hdrparity_i,
   input  wire [7:0]       frame0_cxl_mem_s2m_drs0_dataparity_i,
   input  wire [15:0]      frame0_cxl_mem_s2m_drs0_tag_i,
   input  wire [511:0]     frame0_cxl_mem_s2m_drs0_data_i,
   input  wire             frame0_cxl_mem_s2m_valid_i,
   output wire             frame0_cxl_mem_s2m_ready_o,
   input  wire [1:0]       frame1_cxl_mem_s2m_ndr1_devload_i,
   input  wire             frame1_cxl_mem_s2m_ndr1_valid_i,
   input  wire [2:0]       frame1_cxl_mem_s2m_ndr1_opcode_i,
   input  wire [1:0]       frame1_cxl_mem_s2m_ndr1_metafield_i,
   input  wire [1:0]       frame1_cxl_mem_s2m_ndr1_metavalue_i,
   input  wire [1:0]       frame1_cxl_mem_s2m_ndr1_parity_i,
   input  wire [3:0]       frame1_cxl_mem_s2m_ndr1_rsvd_i,
   input  wire [15:0]      frame1_cxl_mem_s2m_ndr1_tag_i,
   input  wire [1:0]       frame1_cxl_mem_s2m_ndr0_devload_i,
   input  wire             frame1_cxl_mem_s2m_ndr0_valid_i,
   input  wire [2:0]       frame1_cxl_mem_s2m_ndr0_opcode_i,
   input  wire [1:0]       frame1_cxl_mem_s2m_ndr0_metafield_i,
   input  wire [1:0]       frame1_cxl_mem_s2m_ndr0_metavalue_i,
   input  wire [1:0]       frame1_cxl_mem_s2m_ndr0_parity_i,
   input  wire [3:0]       frame1_cxl_mem_s2m_ndr0_rsvd_i,
   input  wire [15:0]      frame1_cxl_mem_s2m_ndr0_tag_i,
   input  wire [54:0]      frame1_cxl_mem_s2m_drs_hdr1_i,
   input  wire             frame1_cxl_mem_s2m_drs0_valid_i,
   input  wire             frame1_cxl_mem_s2m_drs0_poison_i,
   input  wire [2:0]       frame1_cxl_mem_s2m_drs0_opcode_i,
   input  wire [1:0]       frame1_cxl_mem_s2m_drs0_metafield_i,
   input  wire [1:0]       frame1_cxl_mem_s2m_drs0_metavalue_i,
   input  wire [14:0]      frame1_cxl_mem_s2m_drs0_rsvd_i,
   input  wire [8:0]       frame1_cxl_mem_s2m_drs0_rsvd_field1_i, // revb 
   input  wire [1:0]       frame1_cxl_mem_s2m_drs0_devload_i,
   input  wire [3:0]       frame1_cxl_mem_s2m_drs0_rsvd_field0_i,

   input  wire [1:0]       frame1_cxl_mem_s2m_drs0_hdrparity_i,
   input  wire [7:0]       frame1_cxl_mem_s2m_drs0_dataparity_i,
   input  wire [15:0]      frame1_cxl_mem_s2m_drs0_tag_i,
   input  wire [511:0]     frame1_cxl_mem_s2m_drs0_data_i,
   input  wire             frame1_cxl_mem_s2m_valid_i,
   output wire             frame1_cxl_mem_s2m_ready_o,

   //input  cxl_cache_d2h_req_tx_intf    cxl_d2h_req_frame0, // 0 - 3, 1 ready
   //input  [3:0]                        cxl_d2h_req_frame0_valid,
   //output [3:0]                        cxl_d2h_req_frame0_ready,
   //input  cxl_cache_d2h_req_tx_intf    cxl_d2h_req_frame1, // 4 - 7, 1 ready
   //input  [3:0]                        cxl_d2h_req_frame1_valid,
   //output [3:0]                        cxl_d2h_req_frame1_ready,
   //interfaces_cxl_cache_d2h_req_tx
   input  wire [45:0]     frame0_cxl_cache_d2h_req3_address_i,
   input  wire [1:0]      frame0_cxl_cache_d2h_req3_parity_i,
   input  wire [11:0]     frame0_cxl_cache_d2h_req3_cqid_i,
   input  wire [1:0]      frame0_cxl_cache_d2h_req3_clos_i,
   input  wire [3:0]      frame0_cxl_cache_d2h_req3_secid_i,
   input  wire            frame0_cxl_cache_d2h_req3_nontemporal_i,
   input  wire            frame0_cxl_cache_d2h_req3_cachenear_i,
   input  wire            frame0_cxl_cache_d2h_req3_pushwrite_i,
   input  wire [2:0]      frame0_cxl_cache_d2h_req3_strmid_i,
   input  wire [6:0]      frame0_cxl_cache_d2h_req3_rsvd_i,
   input  wire [4:0]      frame0_cxl_cache_d2h_req3_opcode_i,
   input  wire            frame0_cxl_cache_d2h_req3_valid_i,
   input  wire [45:0]     frame0_cxl_cache_d2h_req2_address_i,
   input  wire [1:0]      frame0_cxl_cache_d2h_req2_parity_i,
   input  wire [11:0]     frame0_cxl_cache_d2h_req2_cqid_i,
   input  wire [1:0]      frame0_cxl_cache_d2h_req2_clos_i,
   input  wire [3:0]      frame0_cxl_cache_d2h_req2_secid_i,
   input  wire            frame0_cxl_cache_d2h_req2_nontemporal_i,
   input  wire            frame0_cxl_cache_d2h_req2_cachenear_i,
   input  wire            frame0_cxl_cache_d2h_req2_pushwrite_i,
   input  wire [2:0]      frame0_cxl_cache_d2h_req2_strmid_i,
   input  wire [6:0]      frame0_cxl_cache_d2h_req2_rsvd_i,
   input  wire [4:0]      frame0_cxl_cache_d2h_req2_opcode_i,
   input  wire            frame0_cxl_cache_d2h_req2_valid_i,
   input  wire [45:0]     frame0_cxl_cache_d2h_req1_address_i,
   input  wire [1:0]      frame0_cxl_cache_d2h_req1_parity_i,
   input  wire [11:0]     frame0_cxl_cache_d2h_req1_cqid_i,
   input  wire [1:0]      frame0_cxl_cache_d2h_req1_clos_i,
   input  wire [3:0]      frame0_cxl_cache_d2h_req1_secid_i,
   input  wire            frame0_cxl_cache_d2h_req1_nontemporal_i,
   input  wire            frame0_cxl_cache_d2h_req1_cachenear_i,
   input  wire            frame0_cxl_cache_d2h_req1_pushwrite_i,
   input  wire [2:0]      frame0_cxl_cache_d2h_req1_strmid_i,
   input  wire [6:0]      frame0_cxl_cache_d2h_req1_rsvd_i,
   input  wire [4:0]      frame0_cxl_cache_d2h_req1_opcode_i,
   input  wire            frame0_cxl_cache_d2h_req1_valid_i,
   input  wire [45:0]     frame0_cxl_cache_d2h_req0_address_i,
   input  wire [1:0]      frame0_cxl_cache_d2h_req0_parity_i,
   input  wire [11:0]     frame0_cxl_cache_d2h_req0_cqid_i,
   input  wire [1:0]      frame0_cxl_cache_d2h_req0_clos_i,
   input  wire [3:0]      frame0_cxl_cache_d2h_req0_secid_i,
   input  wire            frame0_cxl_cache_d2h_req0_nontemporal_i,
   input  wire            frame0_cxl_cache_d2h_req0_cachenear_i,
   input  wire            frame0_cxl_cache_d2h_req0_pushwrite_i,
   input  wire [2:0]      frame0_cxl_cache_d2h_req0_strmid_i,
   input  wire [6:0]      frame0_cxl_cache_d2h_req0_rsvd_i,
   input  wire [4:0]      frame0_cxl_cache_d2h_req0_opcode_i,
   input  wire            frame0_cxl_cache_d2h_req0_valid_i,
   input  wire [3:0]      frame0_cxl_cache_d2h_req_valid_i,
   output wire [3:0]      frame0_cxl_cache_d2h_req_ready_o,
   input  wire [45:0]     frame1_cxl_cache_d2h_req3_address_i,
   input  wire [1:0]      frame1_cxl_cache_d2h_req3_parity_i,
   input  wire [11:0]     frame1_cxl_cache_d2h_req3_cqid_i,
   input  wire [1:0]      frame1_cxl_cache_d2h_req3_clos_i,
   input  wire [3:0]      frame1_cxl_cache_d2h_req3_secid_i,
   input  wire            frame1_cxl_cache_d2h_req3_nontemporal_i,
   input  wire            frame1_cxl_cache_d2h_req3_cachenear_i,
   input  wire            frame1_cxl_cache_d2h_req3_pushwrite_i,
   input  wire [2:0]      frame1_cxl_cache_d2h_req3_strmid_i,
   input  wire [6:0]      frame1_cxl_cache_d2h_req3_rsvd_i,
   input  wire [4:0]      frame1_cxl_cache_d2h_req3_opcode_i,
   input  wire            frame1_cxl_cache_d2h_req3_valid_i,
   input  wire [45:0]     frame1_cxl_cache_d2h_req2_address_i,
   input  wire [1:0]      frame1_cxl_cache_d2h_req2_parity_i,
   input  wire [11:0]     frame1_cxl_cache_d2h_req2_cqid_i,
   input  wire [1:0]      frame1_cxl_cache_d2h_req2_clos_i,
   input  wire [3:0]      frame1_cxl_cache_d2h_req2_secid_i,
   input  wire            frame1_cxl_cache_d2h_req2_nontemporal_i,
   input  wire            frame1_cxl_cache_d2h_req2_cachenear_i,
   input  wire            frame1_cxl_cache_d2h_req2_pushwrite_i,
   input  wire [2:0]      frame1_cxl_cache_d2h_req2_strmid_i,
   input  wire [6:0]      frame1_cxl_cache_d2h_req2_rsvd_i,
   input  wire [4:0]      frame1_cxl_cache_d2h_req2_opcode_i,
   input  wire            frame1_cxl_cache_d2h_req2_valid_i,
   input  wire [45:0]     frame1_cxl_cache_d2h_req1_address_i,
   input  wire [1:0]      frame1_cxl_cache_d2h_req1_parity_i,
   input  wire [11:0]     frame1_cxl_cache_d2h_req1_cqid_i,
   input  wire [1:0]      frame1_cxl_cache_d2h_req1_clos_i,
   input  wire [3:0]      frame1_cxl_cache_d2h_req1_secid_i,
   input  wire            frame1_cxl_cache_d2h_req1_nontemporal_i,
   input  wire            frame1_cxl_cache_d2h_req1_cachenear_i,
   input  wire            frame1_cxl_cache_d2h_req1_pushwrite_i,
   input  wire [2:0]      frame1_cxl_cache_d2h_req1_strmid_i,
   input  wire [6:0]      frame1_cxl_cache_d2h_req1_rsvd_i,
   input  wire [4:0]      frame1_cxl_cache_d2h_req1_opcode_i,
   input  wire            frame1_cxl_cache_d2h_req1_valid_i,
   input  wire [45:0]     frame1_cxl_cache_d2h_req0_address_i,
   input  wire [1:0]      frame1_cxl_cache_d2h_req0_parity_i,
   input  wire [11:0]     frame1_cxl_cache_d2h_req0_cqid_i,
   input  wire [1:0]      frame1_cxl_cache_d2h_req0_clos_i,
   input  wire [3:0]      frame1_cxl_cache_d2h_req0_secid_i,
   input  wire            frame1_cxl_cache_d2h_req0_nontemporal_i,
   input  wire            frame1_cxl_cache_d2h_req0_cachenear_i,
   input  wire            frame1_cxl_cache_d2h_req0_pushwrite_i,
   input  wire [2:0]      frame1_cxl_cache_d2h_req0_strmid_i,
   input  wire [6:0]      frame1_cxl_cache_d2h_req0_rsvd_i,
   input  wire [4:0]      frame1_cxl_cache_d2h_req0_opcode_i,
   input  wire            frame1_cxl_cache_d2h_req0_valid_i,
   input  wire [3:0]      frame1_cxl_cache_d2h_req_valid_i,
   output wire [3:0]      frame1_cxl_cache_d2h_req_ready_o,

   //input  cxl_cache_d2h_rsp_tx_intf    cxl_d2h_rsp_frame0, // 0 - 1, 1 ready
   //input  [1:0]                        cxl_d2h_rsp_frame0_valid,
   //output [1:0]                        cxl_d2h_rsp_frame0_ready,
   //input  cxl_cache_d2h_rsp_tx_intf    cxl_d2h_rsp_frame1, // 2 - 3, 1 ready
   //input  [1:0]                        cxl_d2h_rsp_frame1_valid,
   //output [1:0]                        cxl_d2h_rsp_frame1_ready,
   //interfaces_cxl_cache_d2h_rsp_tx
   input  wire [1-1:0]     frame0_cxl_cache_d2h_rsp1_valid_i,
   input  wire [5-1:0]     frame0_cxl_cache_d2h_rsp1_opcode_i,
   input  wire [2-1:0]     frame0_cxl_cache_d2h_rsp1_parity_i,
   input  wire [2-1:0]     frame0_cxl_cache_d2h_rsp1_rsvd_i,
   input  wire [12-1:0]    frame0_cxl_cache_d2h_rsp1_uqid_i,
   input  wire [1-1:0]     frame0_cxl_cache_d2h_rsp0_valid_i,
   input  wire [5-1:0]     frame0_cxl_cache_d2h_rsp0_opcode_i,
   input  wire [2-1:0]     frame0_cxl_cache_d2h_rsp0_parity_i,
   input  wire [2-1:0]     frame0_cxl_cache_d2h_rsp0_rsvd_i,
   input  wire [12-1:0]    frame0_cxl_cache_d2h_rsp0_uqid_i,
   input  wire [2-1:0]     frame0_cxl_cache_d2h_rsp_valid_i,
   output wire [2-1:0]     frame0_cxl_cache_d2h_rsp_ready_o,
   input  wire [1-1:0]     frame1_cxl_cache_d2h_rsp1_valid_i,
   input  wire [5-1:0]     frame1_cxl_cache_d2h_rsp1_opcode_i,
   input  wire [2-1:0]     frame1_cxl_cache_d2h_rsp1_parity_i,
   input  wire [2-1:0]     frame1_cxl_cache_d2h_rsp1_rsvd_i,
   input  wire [12-1:0]    frame1_cxl_cache_d2h_rsp1_uqid_i,
   input  wire [1-1:0]     frame1_cxl_cache_d2h_rsp0_valid_i,
   input  wire [5-1:0]     frame1_cxl_cache_d2h_rsp0_opcode_i,
   input  wire [2-1:0]     frame1_cxl_cache_d2h_rsp0_parity_i,
   input  wire [2-1:0]     frame1_cxl_cache_d2h_rsp0_rsvd_i,
   input  wire [12-1:0]    frame1_cxl_cache_d2h_rsp0_uqid_i,
   input  wire [2-1:0]     frame1_cxl_cache_d2h_rsp_valid_i,
   output wire [2-1:0]     frame1_cxl_cache_d2h_rsp_ready_o,

   //input  cxl_cache_d2h_data_tx_intf   cxl_d2h_data_frame0, // 0, 1 ready
   //input                               cxl_d2h_data_frame0_valid,
   //output                              cxl_d2h_data_frame0_ready,
   //input  cxl_cache_d2h_data_tx_intf   cxl_d2h_data_frame1, // 1, 1 ready
   //input                               cxl_d2h_data_frame1_valid,
   //output                              cxl_d2h_data_frame1_ready,
   //interfaces_cxl_cache_d2h_data_tx
   input  wire [1-1:0]     frame0_cxl_cache_d2h_data_pushwrite_i,
   input  wire [12-1:0]    frame0_cxl_cache_d2h_data_uqid_i,
   input  wire [3-1:0]     frame0_cxl_cache_d2h_data_strmid_i,
   input  wire [2-1:0]     frame0_cxl_cache_d2h_data_hdrparity_i,
   input  wire [1-1:0]     frame0_cxl_cache_d2h_data_valid_i,
   input  wire [1-1:0]     frame0_cxl_cache_d2h_data_bogus_i,
   input  wire [1-1:0]     frame0_cxl_cache_d2h_data_poison_i,
   input  wire [8-1:0]     frame0_cxl_cache_d2h_data_dataparity_i,
   input  wire [1-1:0]     frame0_cxl_cache_d2h_data_rsvd_i,
   input  wire [4-1:0]     frame0_cxl_cache_d2h_data_beparity_i,
   input  wire [64-1:0]    frame0_cxl_cache_d2h_data_byteen_i,
   input  wire [512-1:0]   frame0_cxl_cache_d2h_data_data_i,
   input  wire [1-1:0]     frame0_cxl_cache_d2h_valid_i,
   output wire [1-1:0]     frame0_cxl_cache_d2h_data_ready_o,
   input  wire [1-1:0]     frame1_cxl_cache_d2h_data_pushwrite_i,
   input  wire [12-1:0]    frame1_cxl_cache_d2h_data_uqid_i,
   input  wire [3-1:0]     frame1_cxl_cache_d2h_data_strmid_i,
   input  wire [2-1:0]     frame1_cxl_cache_d2h_data_hdrparity_i,
   input  wire [1-1:0]     frame1_cxl_cache_d2h_data_valid_i,
   input  wire [1-1:0]     frame1_cxl_cache_d2h_data_bogus_i,
   input  wire [1-1:0]     frame1_cxl_cache_d2h_data_poison_i,
   input  wire [8-1:0]     frame1_cxl_cache_d2h_data_dataparity_i,
   input  wire [1-1:0]     frame1_cxl_cache_d2h_data_rsvd_i,
   input  wire [4-1:0]     frame1_cxl_cache_d2h_data_beparity_i,
   input  wire [64-1:0]    frame1_cxl_cache_d2h_data_byteen_i,
   input  wire [512-1:0]   frame1_cxl_cache_d2h_data_data_i,
   input  wire [1-1:0]     frame1_cxl_cache_d2h_valid_i,
   output wire [1-1:0]     frame1_cxl_cache_d2h_data_ready_o,

   //E2E Credit
   output wire             cxl_cache_d2h_data0_crdrtn_o,
   output wire             cxl_cache_d2h_req_crdrtn_o,
   output wire             cxl_cache_d2h_rsp_crdrtn_o,
   output wire             cxl_cache_d2h_pushwr_crdrtn_o,
   output wire             cxl_mem_s2m_drs0_crdrtn_o,
   output wire             cxl_mem_s2m_drs1_crdrtn_o,
   output wire             cxl_mem_s2m_ndr_crdrtn_o,
   input  wire             cxl_cache_h2d_data0_crdrtn_i,
   input  wire             cxl_cache_h2d_data1_crdrtn_i,
   input  wire             cxl_cache_h2d_req_crdrtn_i,
   input  wire             cxl_cache_h2d_rsp_crdrtn_i,
   input  wire             cxl_mem_m2s_req_crdrtn_i,
   input  wire             cxl_mem_m2s_rwd0_crdrtn_i,
   input  wire             cxl_mem_m2s_rwd1_crdrtn_i,
   input  wire             cxl_cache_h2d_rsp_crdrtn_fr0_i,
   input  wire             cxl_cache_h2d_rsp_crdrtn_fr1_i,
   input  wire             cxl_cache_h2d_req_crdrtn_fr0_i,
   input  wire             cxl_cache_h2d_req_crdrtn_fr1_i,
   input  wire             cxl_cache_h2d_data_crdrtn_fr0_i,
   input  wire             cxl_cache_h2d_data_crdrtn_fr1_i,
   input  wire             cxl_mem_m2s_rwd_crdrtn_fr0_i,
   input  wire             cxl_mem_m2s_rwd_crdrtn_fr1_i,
   input  wire             cxl_mem_m2s_req_crdrtn_fr0_i,
   input  wire             cxl_mem_m2s_req_crdrtn_fr1_i,

   output wire             cxl_mem_m2s_viral_o,
   output wire             cxl_cache_h2d_viral_o,
   input  wire             cxl_mem_s2m_viral_i,
   input  wire             cxl_cache_d2h_viral_i,

   output wire             pipe_direct_pld_tx_clk_out_o, // ch13_pipe_direct_pld_pcs_rx_clk_out1_dcm;
   output wire             ln0_pipe_direct_pld_rx_clk_out_o, // ch15_pipe_direct_pld_pcs_rx_clk_out1_dcm;
   output wire             ln1_pipe_direct_pld_rx_clk_out_o, // ch16_pipe_direct_pld_pcs_rx_clk_out1_dcm;
   output wire             ln2_pipe_direct_pld_rx_clk_out_o, // ch17_pipe_direct_pld_pcs_rx_clk_out1_dcm;
   output wire             ln3_pipe_direct_pld_rx_clk_out_o, // ch18_pipe_direct_pld_pcs_rx_clk_out1_dcm;
   output wire             ln4_pipe_direct_pld_rx_clk_out_o, // ch19_pipe_direct_pld_pcs_rx_clk_out1_dcm;
   output wire             ln5_pipe_direct_pld_rx_clk_out_o, // ch20_pipe_direct_pld_pcs_rx_clk_out1_dcm;
   output wire             ln6_pipe_direct_pld_rx_clk_out_o, // ch21_pipe_direct_pld_pcs_rx_clk_out1_dcm;
   output wire             ln7_pipe_direct_pld_rx_clk_out_o, // ch22_pipe_direct_pld_pcs_rx_clk_out1_dcm;
   // PIPE Direct Signals : Async Direc TX
   output wire  [7:0]     ln_pipe_direct_reset_status_n_o,
   
   // PIPE Direct Signals : Async Direc RX
   output wire       octet1_pipe_direct_synthfast_lockstatus_o,
   output wire       octet1_pipe_direct_synthfast_ready_o,
   output wire       octet1_pipe_direct_synthslow_lockstatus_o,
   output wire       octet1_pipe_direct_synthslow_ready_o,
   //output wire       o_ln0_pipe_direct_RXElecIdle,
   //output wire       o_ln1_pipe_direct_RXElecIdle,
   //output wire       o_ln2_pipe_direct_RXElecIdle,
   //output wire       o_ln3_pipe_direct_RXElecIdle,
   //output wire       o_ln4_pipe_direct_RXElecIdle,
   //output wire       o_ln5_pipe_direct_RXElecIdle,
   //output wire       o_ln6_pipe_direct_RXElecIdle,
   //output wire       o_ln7_pipe_direct_RXElecIdle,
   output wire       ln0_pipe_direct_cdrlockstatus_o,
   output wire       ln1_pipe_direct_cdrlockstatus_o,
   output wire       ln2_pipe_direct_cdrlockstatus_o,
   output wire       ln3_pipe_direct_cdrlockstatus_o,
   output wire       ln4_pipe_direct_cdrlockstatus_o,
   output wire       ln5_pipe_direct_cdrlockstatus_o,
   output wire       ln6_pipe_direct_cdrlockstatus_o,
   output wire       ln7_pipe_direct_cdrlockstatus_o,
   output wire       ln0_pipe_direct_cdrlock2data_o,
   output wire       ln1_pipe_direct_cdrlock2data_o,
   output wire       ln2_pipe_direct_cdrlock2data_o,
   output wire       ln3_pipe_direct_cdrlock2data_o,
   output wire       ln4_pipe_direct_cdrlock2data_o,
   output wire       ln5_pipe_direct_cdrlock2data_o,
   output wire       ln6_pipe_direct_cdrlock2data_o,
   output wire       ln7_pipe_direct_cdrlock2data_o,

   // PIPE Direct Signals : Ch 13 TX Deskew Channel
   input  wire       ln0_pipe_direct_rxtermination_i,
   input  wire       ln1_pipe_direct_rxtermination_i,
   input  wire       ln2_pipe_direct_rxtermination_i,
   input  wire       ln3_pipe_direct_rxtermination_i,
   input  wire       ln4_pipe_direct_rxtermination_i,
   input  wire       ln5_pipe_direct_rxtermination_i,
   input  wire       ln6_pipe_direct_rxtermination_i,
   input  wire       ln7_pipe_direct_rxtermination_i,

   input  wire       ln0_pipe_direct_pclkchangeack_i,
   input  wire       ln1_pipe_direct_pclkchangeack_i,
   input  wire       ln2_pipe_direct_pclkchangeack_i,
   input  wire       ln3_pipe_direct_pclkchangeack_i,
   input  wire       ln4_pipe_direct_pclkchangeack_i,
   input  wire       ln5_pipe_direct_pclkchangeack_i,
   input  wire       ln6_pipe_direct_pclkchangeack_i,
   input  wire       ln7_pipe_direct_pclkchangeack_i,
   input  wire       octet1_pipe_direct_deskew_clear_3_i,
   input  wire       octet1_pipe_direct_deskew_clear_2_i,
   input  wire       octet1_pipe_direct_deskew_clear_1_i,
   input  wire       octet1_pipe_direct_deskew_clear_0_i,
   //
   // PIPE Direct Signals : Ch 13 RX Deskew Channel

   output wire       ln0_pipe_direct_rxstandbystatus_o,
   output wire       ln1_pipe_direct_rxstandbystatus_o,
   output wire       ln2_pipe_direct_rxstandbystatus_o,
   output wire       ln3_pipe_direct_rxstandbystatus_o,
   output wire       ln4_pipe_direct_rxstandbystatus_o,
   output wire       ln5_pipe_direct_rxstandbystatus_o,
   output wire       ln6_pipe_direct_rxstandbystatus_o,
   output wire       ln7_pipe_direct_rxstandbystatus_o,
   output wire       ln0_pipe_direct_pclkchangeok_o,
   output wire       ln1_pipe_direct_pclkchangeok_o,
   output wire       ln2_pipe_direct_pclkchangeok_o,
   output wire       ln3_pipe_direct_pclkchangeok_o,
   output wire       ln4_pipe_direct_pclkchangeok_o,
   output wire       ln5_pipe_direct_pclkchangeok_o,
   output wire       ln6_pipe_direct_pclkchangeok_o,
   output wire       ln7_pipe_direct_pclkchangeok_o,
   output wire       ln0_pipe_direct_rxstatus_o,
   output wire       ln1_pipe_direct_rxstatus_o,
   output wire       ln2_pipe_direct_rxstatus_o,
   output wire       ln3_pipe_direct_rxstatus_o,
   output wire       ln4_pipe_direct_rxstatus_o,
   output wire       ln5_pipe_direct_rxstatus_o,
   output wire       ln6_pipe_direct_rxstatus_o,
   output wire       ln7_pipe_direct_rxstatus_o,
   output wire       ln0_pipe_direct_phystatus_o,
   output wire       ln1_pipe_direct_phystatus_o,
   output wire       ln2_pipe_direct_phystatus_o,
   output wire       ln3_pipe_direct_phystatus_o,
   output wire       ln4_pipe_direct_phystatus_o,
   output wire       ln5_pipe_direct_phystatus_o,
   output wire       ln6_pipe_direct_phystatus_o,
   output wire       ln7_pipe_direct_phystatus_o,
   output wire [7:0] octet1_pipe_direct_phy_dsk_active_chans_o,
   output wire [7:0] octet1_pipe_direct_phy_dsk_monitor_err_o,
   output wire       octet1_pipe_direct_phy_dsk_monitor_err_status_3_o,
   output wire [2:0] octet1_pipe_direct_phy_dsk_status_3_o,
   output wire       octet1_pipe_direct_phy_dsk_valid_3_o,
   output wire       octet1_pipe_direct_phy_dsk_eval_done_3_o,
   output wire       octet1_pipe_direct_phy_dsk_monitor_err_status_2_o,
   output wire [2:0] octet1_pipe_direct_phy_dsk_status_2_o,
   output wire       octet1_pipe_direct_phy_dsk_valid_2_o,
   output wire       octet1_pipe_direct_phy_dsk_eval_done_2_o,
   output wire       octet1_pipe_direct_phy_dsk_monitor_err_status_1_o,
   output wire [2:0] octet1_pipe_direct_phy_dsk_status_1_o,
   output wire       octet1_pipe_direct_phy_dsk_valid_1_o,
   output wire       octet1_pipe_direct_phy_dsk_eval_done_1_o,
   output wire       octet1_pipe_direct_phy_dsk_monitor_err_status_0_o,
   output wire [2:0] octet1_pipe_direct_phy_dsk_status_0_o,
   output wire       octet1_pipe_direct_phy_dsk_valid_0_o,
   output wire       octet1_pipe_direct_phy_dsk_eval_done_0_o,

   // PIPE Direct Signals : Ch 14 TX MsgBus
   input  wire [7:0] ln0_m2p_messagebus_i,
   input  wire [7:0] ln1_m2p_messagebus_i,
   input  wire [7:0] ln2_m2p_messagebus_i,
   input  wire [7:0] ln3_m2p_messagebus_i,
   input  wire [7:0] ln4_m2p_messagebus_i,
   input  wire [7:0] ln5_m2p_messagebus_i,
   input  wire [7:0] ln6_m2p_messagebus_i,
   input  wire [7:0] ln7_m2p_messagebus_i,
   //
   // PIPE Direct Signals : Ch 14 RX MsgBus
   output wire [7:0] ln0_p2m_messagebus_o,
   output wire [7:0] ln1_p2m_messagebus_o,
   output wire [7:0] ln2_p2m_messagebus_o,
   output wire [7:0] ln3_p2m_messagebus_o,
   output wire [7:0] ln4_p2m_messagebus_o,
   output wire [7:0] ln5_p2m_messagebus_o,
   output wire [7:0] ln6_p2m_messagebus_o,
   output wire [7:0] ln7_p2m_messagebus_o,

   // PIPE Direct Signals : Ch 15 TX
   input  wire             ln0_pipe_direct_txdeskewmarker_i,
   input  wire             ln0_pipe_direct_rxstandby_i,
   input  wire [3:0]       ln0_pipe_direct_txelecidle_i,
   input  wire [1:0]       ln0_pipe_direct_powerdown_i,
   input  wire [2:0]       ln0_pipe_direct_rate_i,
   input  wire             ln0_pipe_direct_txdetectrx_i,
   input  wire             ln0_pipe_direct_txdatavalid1_i,
   input  wire             ln0_pipe_direct_txdatavalid0_i,
   input  wire [63:0]      ln0_pipe_direct_txdata_i,
   input  wire             ln0_pipe_direct_pld_pcs_rst_n_i,
   // PIPE Direct Signals : Ch 15 RX
   output wire [11:0]      ln0_pipe_direct_reserved_o,
   output wire             ln0_pipe_direct_rxdatavalid1_o,
   output wire             ln0_pipe_direct_rxdatavalid0_o,
   output wire [63:0]      ln0_pipe_direct_rxdata_o,
   output wire             ln0_pipe_direct_rxelecidle_o,

   // PIPE Direct Signals : Ch 16
   input  wire             ln1_pipe_direct_txdeskewmarker_i,
   input  wire             ln1_pipe_direct_rxstandby_i,
   input  wire [3:0]       ln1_pipe_direct_txelecidle_i,
   input  wire [1:0]       ln1_pipe_direct_powerdown_i,
   input  wire [2:0]       ln1_pipe_direct_rate_i,
   input  wire             ln1_pipe_direct_txdetectrx_i,
   input  wire             ln1_pipe_direct_txdatavalid1_i,
   input  wire             ln1_pipe_direct_txdatavalid0_i,
   input  wire [63:0]      ln1_pipe_direct_txdata_i,
   input  wire             ln1_pipe_direct_pld_pcs_rst_n_i,
   output wire [11:0]      ln1_pipe_direct_reserved_o,
   output wire             ln1_pipe_direct_rxdatavalid1_o,
   output wire             ln1_pipe_direct_rxdatavalid0_o,
   output wire [63:0]      ln1_pipe_direct_rxdata_o,
   output wire             ln1_pipe_direct_rxelecidle_o,

   // PIPE Direct Signals : Ch 17
   input  wire             ln2_pipe_direct_txdeskewmarker_i,
   input  wire             ln2_pipe_direct_rxstandby_i,
   input  wire [3:0]       ln2_pipe_direct_txelecidle_i,
   input  wire [1:0]       ln2_pipe_direct_powerdown_i,
   input  wire [2:0]       ln2_pipe_direct_rate_i,
   input  wire             ln2_pipe_direct_txdetectrx_i,
   input  wire             ln2_pipe_direct_txdatavalid1_i,
   input  wire             ln2_pipe_direct_txdatavalid0_i,
   input  wire [63:0]      ln2_pipe_direct_txdata_i,
   input  wire             ln2_pipe_direct_pld_pcs_rst_n_i,
   output wire [11:0]      ln2_pipe_direct_reserved_o,
   output wire             ln2_pipe_direct_rxdatavalid1_o,
   output wire             ln2_pipe_direct_rxdatavalid0_o,
   output wire [63:0]      ln2_pipe_direct_rxdata_o,
   output wire             ln2_pipe_direct_rxelecidle_o,

   // PIPE Direct Signals : Ch 18
   input  wire             ln3_pipe_direct_txdeskewmarker_i,
   input  wire             ln3_pipe_direct_rxstandby_i,
   input  wire [3:0]       ln3_pipe_direct_txelecidle_i,
   input  wire [1:0]       ln3_pipe_direct_powerdown_i,
   input  wire [2:0]       ln3_pipe_direct_rate_i,
   input  wire             ln3_pipe_direct_txdetectrx_i,
   input  wire             ln3_pipe_direct_txdatavalid1_i,
   input  wire             ln3_pipe_direct_txdatavalid0_i,
   input  wire [63:0]      ln3_pipe_direct_txdata_i,
   input  wire             ln3_pipe_direct_pld_pcs_rst_n_i,
   output wire [11:0]      ln3_pipe_direct_reserved_o,
   output wire             ln3_pipe_direct_rxdatavalid1_o,
   output wire             ln3_pipe_direct_rxdatavalid0_o,
   output wire [63:0]      ln3_pipe_direct_rxdata_o,
   output wire             ln3_pipe_direct_rxelecidle_o,

   // PIPE Direct Signals : Ch 19
   input  wire             ln4_pipe_direct_txdeskewmarker_i,
   input  wire             ln4_pipe_direct_rxstandby_i,
   input  wire [3:0]       ln4_pipe_direct_txelecidle_i,
   input  wire [1:0]       ln4_pipe_direct_powerdown_i,
   input  wire [2:0]       ln4_pipe_direct_rate_i,
   input  wire             ln4_pipe_direct_txdetectrx_i,
   input  wire             ln4_pipe_direct_txdatavalid1_i,
   input  wire             ln4_pipe_direct_txdatavalid0_i,
   input  wire [63:0]      ln4_pipe_direct_txdata_i,
   input  wire             ln4_pipe_direct_pld_pcs_rst_n_i,
   output wire [11:0]      ln4_pipe_direct_reserved_o,
   output wire             ln4_pipe_direct_rxdatavalid1_o,
   output wire             ln4_pipe_direct_rxdatavalid0_o,
   output wire [63:0]      ln4_pipe_direct_rxdata_o,
   output wire             ln4_pipe_direct_rxelecidle_o,

   // PIPE Direct Signals : Ch 20
   input  wire             ln5_pipe_direct_txdeskewmarker_i,
   input  wire             ln5_pipe_direct_rxstandby_i,
   input  wire [3:0]       ln5_pipe_direct_txelecidle_i,
   input  wire [1:0]       ln5_pipe_direct_powerdown_i,
   input  wire [2:0]       ln5_pipe_direct_rate_i,
   input  wire             ln5_pipe_direct_txdetectrx_i,
   input  wire             ln5_pipe_direct_txdatavalid1_i,
   input  wire             ln5_pipe_direct_txdatavalid0_i,
   input  wire [63:0]      ln5_pipe_direct_txdata_i,
   input  wire             ln5_pipe_direct_pld_pcs_rst_n_i,
   output wire [11:0]      ln5_pipe_direct_reserved_o,
   output wire             ln5_pipe_direct_rxdatavalid1_o,
   output wire             ln5_pipe_direct_rxdatavalid0_o,
   output wire [63:0]      ln5_pipe_direct_rxdata_o,
   output wire             ln5_pipe_direct_rxelecidle_o,

   // PIPE Direct Signals : Ch 21
   input  wire             ln6_pipe_direct_txdeskewmarker_i,
   input  wire             ln6_pipe_direct_rxstandby_i,
   input  wire [3:0]       ln6_pipe_direct_txelecidle_i,
   input  wire [1:0]       ln6_pipe_direct_powerdown_i,
   input  wire [2:0]       ln6_pipe_direct_rate_i,
   input  wire             ln6_pipe_direct_txdetectrx_i,
   input  wire             ln6_pipe_direct_txdatavalid1_i,
   input  wire             ln6_pipe_direct_txdatavalid0_i,
   input  wire [63:0]      ln6_pipe_direct_txdata_i,
   input  wire             ln6_pipe_direct_pld_pcs_rst_n_i,
   output wire [11:0]      ln6_pipe_direct_reserved_o,
   output wire             ln6_pipe_direct_rxdatavalid1_o,
   output wire             ln6_pipe_direct_rxdatavalid0_o,
   output wire [63:0]      ln6_pipe_direct_rxdata_o,
   output wire             ln6_pipe_direct_rxelecidle_o,

   // PIPE Direct Signals : Ch 22
   input  wire             ln7_pipe_direct_txdeskewmarker_i,
   input  wire             ln7_pipe_direct_rxstandby_i,
   input  wire [3:0]       ln7_pipe_direct_txelecidle_i,
   input  wire [1:0]       ln7_pipe_direct_powerdown_i,
   input  wire [2:0]       ln7_pipe_direct_rate_i,
   input  wire             ln7_pipe_direct_txdetectrx_i,
   input  wire             ln7_pipe_direct_txdatavalid1_i,
   input  wire             ln7_pipe_direct_txdatavalid0_i,
   input  wire [63:0]      ln7_pipe_direct_txdata_i,
   input  wire             ln7_pipe_direct_pld_pcs_rst_n_i,
   output wire [11:0]      ln7_pipe_direct_reserved_o,
   output wire             ln7_pipe_direct_rxdatavalid1_o,
   output wire             ln7_pipe_direct_rxdatavalid0_o,
   output wire [63:0]      ln7_pipe_direct_rxdata_o,
   output wire             ln7_pipe_direct_rxelecidle_o,

   // Serial RX Data Interface
   input  wire         rx_n_in0,                      //          hip_serial.rx_n_in0,              Check User Guide for details
   input  wire         rx_n_in1,                      //                    .rx_n_in1,              Check User Guide for details
   input  wire         rx_n_in2,                      //                    .rx_n_in2,              Check User Guide for details
   input  wire         rx_n_in3,                      //                    .rx_n_in3,              Check User Guide for details
   input  wire         rx_n_in4,                      //                    .rx_n_in4,              Check User Guide for details
   input  wire         rx_n_in5,                      //                    .rx_n_in5,              Check User Guide for details
   input  wire         rx_n_in6,                      //                    .rx_n_in6,              Check User Guide for details
   input  wire         rx_n_in7,                      //                    .rx_n_in7,              Check User Guide for details
   input  wire         rx_n_in8,                      //                    .rx_n_in8,              Check User Guide for details
   input  wire         rx_n_in9,                      //                    .rx_n_in9,              Check User Guide for details
   input  wire         rx_n_in10,                     //                    .rx_n_in10,             Check User Guide for details
   input  wire         rx_n_in11,                     //                    .rx_n_in11,             Check User Guide for details
   input  wire         rx_n_in12,                     //                    .rx_n_in12,             Check User Guide for details
   input  wire         rx_n_in13,                     //                    .rx_n_in13,             Check User Guide for details
   input  wire         rx_n_in14,                     //                    .rx_n_in14,             Check User Guide for details
   input  wire         rx_n_in15,                     //                    .rx_n_in15,             Check User Guide for details
   input  wire         rx_p_in0,                      //                    .rx_p_in0,              Check User Guide for details
   input  wire         rx_p_in1,                      //                    .rx_p_in1,              Check User Guide for details
   input  wire         rx_p_in2,                      //                    .rx_p_in2,              Check User Guide for details
   input  wire         rx_p_in3,                      //                    .rx_p_in3,              Check User Guide for details
   input  wire         rx_p_in4,                      //                    .rx_p_in4,              Check User Guide for details
   input  wire         rx_p_in5,                      //                    .rx_p_in5,              Check User Guide for details
   input  wire         rx_p_in6,                      //                    .rx_p_in6,              Check User Guide for details
   input  wire         rx_p_in7,                      //                    .rx_p_in7,              Check User Guide for details
   input  wire         rx_p_in8,                      //                    .rx_p_in8,              Check User Guide for details
   input  wire         rx_p_in9,                      //                    .rx_p_in9,              Check User Guide for details
   input  wire         rx_p_in10,                     //                    .rx_p_in10,             Check User Guide for details
   input  wire         rx_p_in11,                     //                    .rx_p_in11,             Check User Guide for details
   input  wire         rx_p_in12,                     //                    .rx_p_in12,             Check User Guide for details
   input  wire         rx_p_in13,                     //                    .rx_p_in13,             Check User Guide for details
   input  wire         rx_p_in14,                     //                    .rx_p_in14,             Check User Guide for details
   input  wire         rx_p_in15,                     //                    .rx_p_in15,             Check User Guide for details
   // Serial TX Data Interface
   output wire         tx_n_out0,                     //                    .tx_n_out0,             Check User Guide for details
   output wire         tx_n_out1,                     //                    .tx_n_out1,             Check User Guide for details
   output wire         tx_n_out2,                     //                    .tx_n_out2,             Check User Guide for details
   output wire         tx_n_out3,                     //                    .tx_n_out3,             Check User Guide for details
   output wire         tx_n_out4,                     //                    .tx_n_out4,             Check User Guide for details
   output wire         tx_n_out5,                     //                    .tx_n_out5,             Check User Guide for details
   output wire         tx_n_out6,                     //                    .tx_n_out6,             Check User Guide for details
   output wire         tx_n_out7,                     //                    .tx_n_out7,             Check User Guide for details
   output wire         tx_n_out8,                     //                    .tx_n_out8,             Check User Guide for details
   output wire         tx_n_out9,                     //                    .tx_n_out9,             Check User Guide for details
   output wire         tx_n_out10,                    //                    .tx_n_out10,            Check User Guide for details
   output wire         tx_n_out11,                    //                    .tx_n_out11,            Check User Guide for details
   output wire         tx_n_out12,                    //                    .tx_n_out12,            Check User Guide for details
   output wire         tx_n_out13,                    //                    .tx_n_out13,            Check User Guide for details
   output wire         tx_n_out14,                    //                    .tx_n_out14,            Check User Guide for details
   output wire         tx_n_out15,                    //                    .tx_n_out15,            Check User Guide for details
   output wire         tx_p_out0,                     //                    .tx_p_out0,             Check User Guide for details
   output wire         tx_p_out1,                     //                    .tx_p_out1,             Check User Guide for details
   output wire         tx_p_out2,                     //                    .tx_p_out2,             Check User Guide for details
   output wire         tx_p_out3,                     //                    .tx_p_out3,             Check User Guide for details
   output wire         tx_p_out4,                     //                    .tx_p_out4,             Check User Guide for details
   output wire         tx_p_out5,                     //                    .tx_p_out5,             Check User Guide for details
   output wire         tx_p_out6,                     //                    .tx_p_out6,             Check User Guide for details
   output wire         tx_p_out7,                     //                    .tx_p_out7,             Check User Guide for details
   output wire         tx_p_out8,                     //                    .tx_p_out8,             Check User Guide for details
   output wire         tx_p_out9,                     //                    .tx_p_out9,             Check User Guide for details
   output wire         tx_p_out10,                    //                    .tx_p_out10,            Check User Guide for details
   output wire         tx_p_out11,                    //                    .tx_p_out11,            Check User Guide for details
   output wire         tx_p_out12,                    //                    .tx_p_out12,            Check User Guide for details
   output wire         tx_p_out13,                    //                    .tx_p_out13,            Check User Guide for details
   output wire         tx_p_out14,                    //                    .tx_p_out14,            Check User Guide for details
   output wire         tx_p_out15,                    //                    .tx_p_out15,            Check User Guide for details
   // IOSF Interface
   output wire         p0_mnpput_o,                        // Non-Posted Put from master to target
   output wire         p0_mpcput_o,                        // Posted or Completion Put from master to target
   input  wire         p0_mnpcup_i,                        // Non-Posted Credit Update from target to master
   input  wire         p0_mpccup_i,                        // Posted or Completion Credit Update from target to master
   output wire         p0_meom_o,                          // End of Message from master to target
   output wire [15:0]  p0_mpayload_o,                      // Message Payload from master to target
   output wire         p0_mparity_o,                       // Parity for message payload
   input  wire [ 2:0]  p0_side_ism_fabric_i,               //
   input  wire         p0_tnpput_i,                        // Non-Posted Put from master to target
   input  wire         p0_tpcput_i,                        // Posted or Completion Put from master to target
   output wire         p0_tnpcup_o,                        // Non-Posted Credit Update from target to master
   output wire         p0_tpccup_o,                        // Posted or Completion Credit Update from target to master
   input  wire         p0_teom_i,                          // End of Message from master to target
   input  wire [15:0]  p0_tpayload_i,                      // Message Payload from master to target
   input  wire         p0_tparity_i,                       // Parity for message payload
   output wire [ 2:0]  p0_side_ism_agent_o,
   // PTM Signals
   output wire         p0_ptm_clk_updated_o,
   output wire         p0_ptm_context_valid_o,
   output wire [63:0]  p0_ptm_local_clock_o,
   input  wire         p0_ptm_manual_update_i,


   input  wire          p0_pld_warm_rst_rdy_i,       //PORT_NAME_CHANGE cxl_pld_warm_rst_rdy_i,
   output wire          p0_pld_link_req_rst_o,       //PORT_NAME_CHANGE cxl_pld_link_req_rst_o,
   output wire          p0_pld_core_cold_rst_n,      //PORT_NAME_CHANGE cxl_pld_core_cold_rst_n,
   output wire          p0_pld_core_warm_rst_n,      //PORT_NAME_CHANGE cxl_pld_core_warm_rst_n,

   // Reconfig Interface
   input  wire         reconfig_clk,
   input  wire [20:0]  reconfig_address,
   input  wire         reconfig_read,
   output wire [ 7:0]  reconfig_readdata,
   output wire         reconfig_readdatavalid,
   input  wire         reconfig_write,
   input  wire [ 7:0]  reconfig_writedata,
   output wire [ 4:0]  reconfig_reserved_out,
   output wire         reconfig_waitrequest,

    //p0_application error reporting
    input                 p0_app_err_valid_i,
    input [31:0]          p0_app_err_hdr_i,
    input [13:0]          p0_app_err_info_i,
    input [2:0]           p0_app_err_func_num_i,
    input                   p0_app_err_vfa_i,
    input [10:0]            p0_app_err_vf_num_i,
    output                p0_app_err_ready_o,
    // Completion timeout
    output                 p0_cpl_timeout_o,
    output [2:0]           p0_cpl_timeout_func_num_o,
    output [10:0]          p0_cpl_timeout_vfunc_num_o, 
    output                 p0_cpl_timeout_vfunc_active_o,
    output [2:0]           p0_cpl_timeout_cpl_tc_o, 
    output [1:0]           p0_cpl_timeout_cpl_attr_o, 
    output [11:0]          p0_cpl_timeout_cpl_len_o, 
    output [9:0]           p0_cpl_timeout_cpl_tag_o,
    // FLR
    output [7:0]           p0_flr_rcvd_pf_o,
    output                 p0_flr_rcvd_vf_o,
    output [2:0]           p0_flr_rcvd_pf_num_o,
    output [10:0]          p0_flr_rcvd_vf_num_o,
    input  [7:0]           p0_flr_completed_pf_i,
    input                  p0_flr_completed_vf_i,
    input  [2:0]           p0_flr_completed_pf_num_i,
    input  [10:0]          p0_flr_completed_vf_num_i,
    output                 p0_flr_completed_ready_o,
    // CII
    output                 p0_cii_req_o,
    output                 p0_cii_hdr_poisoned_o,
    output [3:0]           p0_cii_hdr_first_be_o,
    output [2:0]           p0_cii_func_num_o,
    output                 p0_cii_wr_vf_active_o,
    output [10:0]          p0_cii_vf_num_o,
    output                 p0_cii_wr_o,
    output [9:0]           p0_cii_addr_o,
    output [31:0]          p0_cii_dout_o,
    input                  p0_cii_override_en_i,
    input [31:0]           p0_cii_override_din_i,
    input                  p0_cii_halt_i,
    input                  p0_cii_convert_pfd_i,
    input [31:0]           p0_cii_conv_pfdata_i,
    //MMIO
    output                  p0_pci_cfg_req_o,
    output [2:0]            p0_pci_cfg_func_num_o,
    output [2:0]            p0_pci_cfg_len_o,
    output [7:0]            p0_pci_cfg_bar_o,
    output [31:0]           p0_pci_cfg_offset_o,
    output                  p0_pci_cfg_wr_o,
    output [31:0]           p0_pci_cfg_writedata_o,
    output [2:0]            p0_pci_cfg_tag_o,
    output [3:0]            p0_pci_cfg_be_o,
    input  [31:0]           p0_pci_cfg_readdata_i,
    input                   p0_pci_cfg_ack_i,
    input                   p0_pci_cfg_df_i,
    input [1:0]             p0_pci_cfg_status_i,
    
    // User AVMM using custom registercxl_access
    input   [31:0]         p0_hip_reconfig_address_i,
    input                  p0_hip_reconfig_write_i,
    input   [7:0]          p0_hip_reconfig_writedata_i,
    input                  p0_hip_reconfig_read_i,
    output                 p0_hip_reconfig_readdatavalid_o,
    output  [7:0]          p0_hip_reconfig_readdata_o,
    output                 p0_hip_reconfig_waitrequest_o,
    output  [1:0]          p0_hip_reconfig_resp_o,
    input                  p0_hip_reconfig_requesttype_i,
    // [Hidden] avmm interface for MMIO CSB to HIP 
////    input                  p0_dbg_mmio_rst_n,
////    input                  p0_dbg_mmio_clk,
////    input   [20:0]         p0_dbg_mmio_address,
////    input                  p0_dbg_mmio_write,
////    input   [7:0]          p0_dbg_mmio_writedata,
////    input                  p0_dbg_mmio_read,
////    output                 p0_dbg_mmio_readdatavalid,
////    output  [7:0]          p0_dbg_mmio_readdata,
////    output                 p0_dbg_mmio_waitrequest,

  //CXL pm
    output logic            p0_pm_valid_o,
    output logic [7:0]      p0_pm_opcode_o,
    output logic [3:0]      p0_pm_tag_o,
    output logic [2:0]      p0_pm_misc_o,
    output logic [127:0]    p0_pm_data_o,
    input                   p0_pm_valid_i,
    input [7:0]             p0_pm_opcode_i,
    input [3:0]             p0_pm_tag_i,
    input [2:0]             p0_pm_misc_i,
    input [127:0]           p0_pm_data_i,
    // CXL aer
    output logic            p0_aermsg_correctable_valid_o,
    output logic            p0_aermsg_uncorrectable_valid_o,
    output logic            p0_aermsg_res_o,
    output logic            p0_aermsg_bts_o,
    output logic            p0_aermsg_bds_o,
    output logic            p0_aermsg_rrs_o,
    output logic            p0_aermsg_rtts_o,
    output logic            p0_aermsg_anes_o,
    output logic            p0_aermsg_cies_o,
    output logic            p0_aermsg_hlos_o,
    output logic [1:0]      p0_aermsg_fmt_o,
    output logic [4:0]      p0_aermsg_type_o,
    output logic [2:0]      p0_aermsg_tc_o,
    output logic            p0_aermsg_ido_o,
    output logic            p0_aermsg_th_o,
    output logic            p0_aermsg_td_o,
    output logic            p0_aermsg_ep_o,
    output logic            p0_aermsg_ro_o,
    output logic            p0_aermsg_ns_o,
    output logic [1:0]      p0_aermsg_at_o,
    output logic [9:0]      p0_aermsg_length_o,
    output logic [95:0]     p0_aermsg_header_o,
    output logic            p0_aermsg_und_o,
    output logic            p0_aermsg_anf_o,
    output logic            p0_aermsg_dlpes_o,
    output logic            p0_aermsg_sdes_o,
    output logic [4:0]      p0_aermsg_fep_o,
    output logic            p0_aermsg_pts_o,
    output logic            p0_aermsg_fcpes_o,
    output logic            p0_aermsg_cts_o,
    output logic            p0_aermsg_cas_o,
    output logic            p0_aermsg_ucs_o,
    output logic            p0_aermsg_ros_o,
    output logic            p0_aermsg_mts_o,
    output logic            p0_aermsg_uies_o,
    output logic            p0_aermsg_mbts_o,
    output logic            p0_aermsg_aebs_o,
    output logic            p0_aermsg_tpbes_o,
    output logic            p0_aermsg_ees_o,
    output logic            p0_aermsg_ures_o,
    output logic            p0_aermsg_avs_o,
    //CXL cfgupdate
    output logic            p0_cfgupdate_valid_o,
    output logic [6:0]      p0_cfgupdate_regtype_o,
    output logic            p0_cfgupdate_vfa_o,
    output logic [2:0]      p0_cfgupdate_pfnum_o,
    output logic [10:0]     p0_cfgupdate_vfnum_o,
    output logic [31:0]     p0_cfgupdate_info_o,       // [47:32] Reserved
    // CXL HIP_ERR
    output logic            p0_hip_err_valid_o,
    output logic [31:0]     p0_hip_err_hdr_o,
    output logic [13:0]     p0_hip_err_info_o,
    output logic [2:0]      p0_hip_err_pf_num_o,
    output logic            p0_hip_err_vfa_o,
    output logic [10:0]     p0_hip_err_vf_num_o,
    output logic            cache_mem_crd_flow_err_o,
    //CXL sim time reduction
    output         phy_sys_ial_0__pipe_Reset_l,
    output         phy_sys_ial_1__pipe_Reset_l,
    output         phy_sys_ial_2__pipe_Reset_l,
    output         phy_sys_ial_3__pipe_Reset_l,
    output         phy_sys_ial_4__pipe_Reset_l,
    output         phy_sys_ial_5__pipe_Reset_l,
    output         phy_sys_ial_6__pipe_Reset_l,
    output         phy_sys_ial_7__pipe_Reset_l,
    output         phy_sys_ial_8__pipe_Reset_l,
    output         phy_sys_ial_9__pipe_Reset_l,
    output         phy_sys_ial_10__pipe_Reset_l,
    output         phy_sys_ial_11__pipe_Reset_l,
    output         phy_sys_ial_12__pipe_Reset_l,
    output         phy_sys_ial_13__pipe_Reset_l,
    output         phy_sys_ial_14__pipe_Reset_l,
    output         phy_sys_ial_15__pipe_Reset_l,	
    output 	o_phy_0_pipe_TxDataValid,
    output [39:0]	o_phy_0_pipe_TxData,
    output	o_phy_0_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_0_pipe_TxElecIdle,
    output [3:0]	o_phy_0_pipe_PowerDown,
    output [2:0]	o_phy_0_pipe_Rate,
    output 	o_phy_0_pipe_PclkChangeAck,
    output [2:0]	o_phy_0_pipe_PCLKRate,
    output [1:0]	o_phy_0_pipe_Width,
    output	o_phy_0_pipe_PCLK,
    output	o_phy_0_pipe_rxelecidle_disable,
    output	o_phy_0_pipe_txcmnmode_disable,
    output	o_phy_0_pipe_srisenable,
    input		i_phy_0_pipe_RxClk,
    input		i_phy_0_pipe_RxValid,
    input	[39:0]	i_phy_0_pipe_RxData,
    input		i_phy_0_pipe_RxElecIdle,
    input	[2:0]	i_phy_0_pipe_RxStatus,
    input		i_phy_0_pipe_RxStandbyStatus,
    output	o_phy_0_pipe_RxStandby,
    output	o_phy_0_pipe_RxTermination,
    output [1:0]	o_phy_0_pipe_RxWidth,
    input		i_phy_0_pipe_PhyStatus,
    input		i_phy_0_pipe_PclkChangeOk,
    output [7:0]	o_phy_0_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_0_pipe_P2M_MessageBus,
    output	o_phy_1_pipe_TxDataValid,
    output [39:0]	o_phy_1_pipe_TxData,
    output	o_phy_1_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_1_pipe_TxElecIdle,
    output [3:0]	o_phy_1_pipe_PowerDown,
    output [2:0]	o_phy_1_pipe_Rate,
    output 	o_phy_1_pipe_PclkChangeAck,
    output [2:0]	o_phy_1_pipe_PCLKRate,
    output [1:0]	o_phy_1_pipe_Width,
    output	o_phy_1_pipe_PCLK,
    output	o_phy_1_pipe_rxelecidle_disable,
    output	o_phy_1_pipe_txcmnmode_disable,
    output	o_phy_1_pipe_srisenable,
    input		i_phy_1_pipe_RxClk,
    input		i_phy_1_pipe_RxValid,
    input	 [39:0]	i_phy_1_pipe_RxData,
    input	 	i_phy_1_pipe_RxElecIdle,
    input	 [2:0]	i_phy_1_pipe_RxStatus,
    input		i_phy_1_pipe_RxStandbyStatus,
    output	o_phy_1_pipe_RxStandby,
    output	o_phy_1_pipe_RxTermination,
    output [1:0]	o_phy_1_pipe_RxWidth,
    input	 	i_phy_1_pipe_PhyStatus,
    input	 	i_phy_1_pipe_PclkChangeOk,
    output [7:0]	o_phy_1_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_1_pipe_P2M_MessageBus,
    output	o_phy_2_pipe_TxDataValid,
    output [39:0]	o_phy_2_pipe_TxData,
    output 	o_phy_2_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_2_pipe_TxElecIdle,
    output [3:0]	o_phy_2_pipe_PowerDown,
    output [2:0]	o_phy_2_pipe_Rate,
    output 	o_phy_2_pipe_PclkChangeAck,
    output [2:0]	o_phy_2_pipe_PCLKRate,
    output [1:0]	o_phy_2_pipe_Width,
    output	o_phy_2_pipe_PCLK,
    output	o_phy_2_pipe_rxelecidle_disable,
    output	o_phy_2_pipe_txcmnmode_disable,
    output	o_phy_2_pipe_srisenable,
    input		i_phy_2_pipe_RxClk,
    input		i_phy_2_pipe_RxValid,
    input	[39:0]	i_phy_2_pipe_RxData,
    input		i_phy_2_pipe_RxElecIdle,
    input	[2:0]	i_phy_2_pipe_RxStatus,
    input		i_phy_2_pipe_RxStandbyStatus,
    output	o_phy_2_pipe_RxStandby,
    output	o_phy_2_pipe_RxTermination,
    output [1:0]	o_phy_2_pipe_RxWidth,
    input		i_phy_2_pipe_PhyStatus,
    input		i_phy_2_pipe_PclkChangeOk,
    output [7:0]	o_phy_2_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_2_pipe_P2M_MessageBus,
    output	o_phy_3_pipe_TxDataValid,
    output [39:0]	o_phy_3_pipe_TxData,
    output 	o_phy_3_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_3_pipe_TxElecIdle,
    output [3:0]	o_phy_3_pipe_PowerDown,
    output [2:0]	o_phy_3_pipe_Rate,
    output 	o_phy_3_pipe_PclkChangeAck,
    output [2:0]	o_phy_3_pipe_PCLKRate,
    output [1:0]	o_phy_3_pipe_Width,
    output	o_phy_3_pipe_PCLK,
    output	o_phy_3_pipe_rxelecidle_disable,
    output	o_phy_3_pipe_txcmnmode_disable,
    output	o_phy_3_pipe_srisenable,
    input		i_phy_3_pipe_RxClk,
    input		i_phy_3_pipe_RxValid,
    input	 [39:0]	i_phy_3_pipe_RxData,
    input	 	i_phy_3_pipe_RxElecIdle,
    input	 [2:0]	i_phy_3_pipe_RxStatus,
    input		i_phy_3_pipe_RxStandbyStatus,
    output	o_phy_3_pipe_RxStandby,
    output	o_phy_3_pipe_RxTermination,
    output [1:0]	o_phy_3_pipe_RxWidth,
    input		i_phy_3_pipe_PhyStatus,
    input		i_phy_3_pipe_PclkChangeOk,
    output [7:0]	o_phy_3_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_3_pipe_P2M_MessageBus,
    output	o_phy_4_pipe_TxDataValid,
    output [39:0]	o_phy_4_pipe_TxData,
    output 	o_phy_4_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_4_pipe_TxElecIdle,
    output [3:0]	o_phy_4_pipe_PowerDown,
    output [2:0]	o_phy_4_pipe_Rate,
    output 	o_phy_4_pipe_PclkChangeAck,
    output [2:0]	o_phy_4_pipe_PCLKRate,
    output [1:0]	o_phy_4_pipe_Width,
    output	o_phy_4_pipe_PCLK,
    output	o_phy_4_pipe_rxelecidle_disable,
    output	o_phy_4_pipe_txcmnmode_disable,
    output	o_phy_4_pipe_srisenable,
    input		i_phy_4_pipe_RxClk,
    input		i_phy_4_pipe_RxValid,
    input	 [39:0]	i_phy_4_pipe_RxData,
    input	 	i_phy_4_pipe_RxElecIdle,
    input	 [2:0]	i_phy_4_pipe_RxStatus,
    input	 	i_phy_4_pipe_RxStandbyStatus,
    output 	o_phy_4_pipe_RxStandby,
    output 	o_phy_4_pipe_RxTermination,
    output [1:0]	o_phy_4_pipe_RxWidth,
    input	 	i_phy_4_pipe_PhyStatus,
    input	 	i_phy_4_pipe_PclkChangeOk,
    output [7:0]	o_phy_4_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_4_pipe_P2M_MessageBus,
    output 	o_phy_5_pipe_TxDataValid,
    output [39:0]	o_phy_5_pipe_TxData,
    output 	o_phy_5_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_5_pipe_TxElecIdle,
    output [3:0]	o_phy_5_pipe_PowerDown,
    output [2:0]	o_phy_5_pipe_Rate,
    output 	o_phy_5_pipe_PclkChangeAck,
    output [2:0]	o_phy_5_pipe_PCLKRate,
    output [1:0]	o_phy_5_pipe_Width,
    output 	o_phy_5_pipe_PCLK,
    output 	o_phy_5_pipe_rxelecidle_disable,
    output 	o_phy_5_pipe_txcmnmode_disable,
    output 	o_phy_5_pipe_srisenable,
    input	 	i_phy_5_pipe_RxClk,
    input	 	i_phy_5_pipe_RxValid,
    input	 [39:0]	i_phy_5_pipe_RxData,
    input	 	i_phy_5_pipe_RxElecIdle,
    input	 [2:0]	i_phy_5_pipe_RxStatus,
    input	 	i_phy_5_pipe_RxStandbyStatus,
    output 	o_phy_5_pipe_RxStandby,
    output 	o_phy_5_pipe_RxTermination,
    output [1:0]	o_phy_5_pipe_RxWidth,
    input	 	i_phy_5_pipe_PhyStatus,
    input	 	i_phy_5_pipe_PclkChangeOk,
    output [7:0]	o_phy_5_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_5_pipe_P2M_MessageBus,
    output 	o_phy_6_pipe_TxDataValid,
    output [39:0]	o_phy_6_pipe_TxData,
    output 	o_phy_6_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_6_pipe_TxElecIdle,
    output [3:0]	o_phy_6_pipe_PowerDown,
    output [2:0]	o_phy_6_pipe_Rate,
    output 	o_phy_6_pipe_PclkChangeAck,
    output [2:0]	o_phy_6_pipe_PCLKRate,
    output [1:0]	o_phy_6_pipe_Width,
    output 	o_phy_6_pipe_PCLK,
    output 	o_phy_6_pipe_rxelecidle_disable,
    output 	o_phy_6_pipe_txcmnmode_disable,
    output 	o_phy_6_pipe_srisenable,
    input	 	i_phy_6_pipe_RxClk,
    input	 	i_phy_6_pipe_RxValid,
    input	 [39:0]	i_phy_6_pipe_RxData,
    input	 	i_phy_6_pipe_RxElecIdle,
    input	 [2:0]	i_phy_6_pipe_RxStatus,
    input	 	i_phy_6_pipe_RxStandbyStatus,
    output 	o_phy_6_pipe_RxStandby,
    output 	o_phy_6_pipe_RxTermination,
    output [1:0]	o_phy_6_pipe_RxWidth,
    input	 	i_phy_6_pipe_PhyStatus,
    input	 	i_phy_6_pipe_PclkChangeOk,
    output [7:0]	o_phy_6_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_6_pipe_P2M_MessageBus,
    output 	o_phy_7_pipe_TxDataValid,
    output [39:0]	o_phy_7_pipe_TxData,
    output 	o_phy_7_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_7_pipe_TxElecIdle,
    output [3:0]	o_phy_7_pipe_PowerDown,
    output [2:0]	o_phy_7_pipe_Rate,
    output 	o_phy_7_pipe_PclkChangeAck,
    output [2:0]	o_phy_7_pipe_PCLKRate,
    output [1:0]	o_phy_7_pipe_Width,
    output 	o_phy_7_pipe_PCLK,
    output 	o_phy_7_pipe_rxelecidle_disable,
    output 	o_phy_7_pipe_txcmnmode_disable,
    output 	o_phy_7_pipe_srisenable,
    input	 	i_phy_7_pipe_RxClk,
    input	 	i_phy_7_pipe_RxValid,
    input	 [39:0]	i_phy_7_pipe_RxData,
    input	 	i_phy_7_pipe_RxElecIdle,
    input	 [2:0]	i_phy_7_pipe_RxStatus,
    input	 	i_phy_7_pipe_RxStandbyStatus,
    output 	o_phy_7_pipe_RxStandby,
    output 	o_phy_7_pipe_RxTermination,
    output [1:0]	o_phy_7_pipe_RxWidth,
    input	 	i_phy_7_pipe_PhyStatus,
    input	 	i_phy_7_pipe_PclkChangeOk,
    output [7:0]	o_phy_7_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_7_pipe_P2M_MessageBus,
    output 	o_phy_8_pipe_TxDataValid,
    output [39:0]	o_phy_8_pipe_TxData,
    output 	o_phy_8_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_8_pipe_TxElecIdle,
    output [3:0]	o_phy_8_pipe_PowerDown,
    output [2:0]	o_phy_8_pipe_Rate,
    output 	o_phy_8_pipe_PclkChangeAck,
    output [2:0]	o_phy_8_pipe_PCLKRate,
    output [1:0]	o_phy_8_pipe_Width,
    output 	o_phy_8_pipe_PCLK,
    output 	o_phy_8_pipe_rxelecidle_disable,
    output 	o_phy_8_pipe_txcmnmode_disable,
    output 	o_phy_8_pipe_srisenable,
    input	 	i_phy_8_pipe_RxClk,
    input	 	i_phy_8_pipe_RxValid,
    input	 [39:0]	i_phy_8_pipe_RxData,
    input	 	i_phy_8_pipe_RxElecIdle,
    input	 [2:0]	i_phy_8_pipe_RxStatus,
    input	 	i_phy_8_pipe_RxStandbyStatus,
    output 	o_phy_8_pipe_RxStandby,
    output 	o_phy_8_pipe_RxTermination,
    output [1:0]	o_phy_8_pipe_RxWidth,
    input	 	i_phy_8_pipe_PhyStatus,
    input	 	i_phy_8_pipe_PclkChangeOk,
    output [7:0]	o_phy_8_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_8_pipe_P2M_MessageBus,
    output 	o_phy_9_pipe_TxDataValid,
    output [39:0]	o_phy_9_pipe_TxData,
    output 	o_phy_9_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_9_pipe_TxElecIdle,
    output [3:0]	o_phy_9_pipe_PowerDown,
    output [2:0]	o_phy_9_pipe_Rate,
    output 	o_phy_9_pipe_PclkChangeAck,
    output [2:0]	o_phy_9_pipe_PCLKRate,
    output [1:0]	o_phy_9_pipe_Width,
    output 	o_phy_9_pipe_PCLK,
    output 	o_phy_9_pipe_rxelecidle_disable,
    output 	o_phy_9_pipe_txcmnmode_disable,
    output 	o_phy_9_pipe_srisenable,
    input	 	i_phy_9_pipe_RxClk,
    input	 	i_phy_9_pipe_RxValid,
    input	 [39:0]	i_phy_9_pipe_RxData,
    input	 	i_phy_9_pipe_RxElecIdle,
    input	 [2:0]	i_phy_9_pipe_RxStatus,
    input	 	i_phy_9_pipe_RxStandbyStatus,
    output 	o_phy_9_pipe_RxStandby,
    output 	o_phy_9_pipe_RxTermination,
    output [1:0]	o_phy_9_pipe_RxWidth,
    input	 	i_phy_9_pipe_PhyStatus,
    input	 	i_phy_9_pipe_PclkChangeOk,
    output [7:0]	o_phy_9_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_9_pipe_P2M_MessageBus,
    output 	o_phy_10_pipe_TxDataValid,
    output [39:0]	o_phy_10_pipe_TxData,
    output 	o_phy_10_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_10_pipe_TxElecIdle,
    output [3:0]	o_phy_10_pipe_PowerDown,
    output [2:0]	o_phy_10_pipe_Rate,
    output 	o_phy_10_pipe_PclkChangeAck,
    output [2:0]	o_phy_10_pipe_PCLKRate,
    output [1:0]	o_phy_10_pipe_Width,
    output 	o_phy_10_pipe_PCLK,
    output 	o_phy_10_pipe_rxelecidle_disable,
    output 	o_phy_10_pipe_txcmnmode_disable,
    output 	o_phy_10_pipe_srisenable,
    input	 	i_phy_10_pipe_RxClk,
    input	 	i_phy_10_pipe_RxValid,
    input	 [39:0]	i_phy_10_pipe_RxData,
    input	 	i_phy_10_pipe_RxElecIdle,
    input	 [2:0]	i_phy_10_pipe_RxStatus,
    input	 	i_phy_10_pipe_RxStandbyStatus,
    output 	o_phy_10_pipe_RxStandby,
    output 	o_phy_10_pipe_RxTermination,
    output [1:0]	o_phy_10_pipe_RxWidth,
    input	 	i_phy_10_pipe_PhyStatus,
    input	 	i_phy_10_pipe_PclkChangeOk,
    output [7:0]	o_phy_10_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_10_pipe_P2M_MessageBus,
    output 	o_phy_11_pipe_TxDataValid,
    output [39:0]	o_phy_11_pipe_TxData,
    output 	o_phy_11_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_11_pipe_TxElecIdle,
    output [3:0]	o_phy_11_pipe_PowerDown,
    output [2:0]	o_phy_11_pipe_Rate,
    output 	o_phy_11_pipe_PclkChangeAck,
    output [2:0]	o_phy_11_pipe_PCLKRate,
    output [1:0]	o_phy_11_pipe_Width,
    output 	o_phy_11_pipe_PCLK,
    output 	o_phy_11_pipe_rxelecidle_disable,
    output 	o_phy_11_pipe_txcmnmode_disable,
    output 	o_phy_11_pipe_srisenable,
    input	 	i_phy_11_pipe_RxClk,
    input	 	i_phy_11_pipe_RxValid,
    input	 [39:0]	i_phy_11_pipe_RxData,
    input	 	i_phy_11_pipe_RxElecIdle,
    input	 [2:0]	i_phy_11_pipe_RxStatus,
    input	 	i_phy_11_pipe_RxStandbyStatus,
    output 	o_phy_11_pipe_RxStandby,
    output 	o_phy_11_pipe_RxTermination,
    output [1:0]	o_phy_11_pipe_RxWidth,
    input	 	i_phy_11_pipe_PhyStatus,
    input	 	i_phy_11_pipe_PclkChangeOk,
    output [7:0]	o_phy_11_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_11_pipe_P2M_MessageBus,
    output 	o_phy_12_pipe_TxDataValid,
    output [39:0]	o_phy_12_pipe_TxData,
    output 	o_phy_12_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_12_pipe_TxElecIdle,
    output [3:0]	o_phy_12_pipe_PowerDown,
    output [2:0]	o_phy_12_pipe_Rate,
    output 	o_phy_12_pipe_PclkChangeAck,
    output [2:0]	o_phy_12_pipe_PCLKRate,
    output [1:0]	o_phy_12_pipe_Width,
    output 	o_phy_12_pipe_PCLK,
    output 	o_phy_12_pipe_rxelecidle_disable,
    output 	o_phy_12_pipe_txcmnmode_disable,
    output 	o_phy_12_pipe_srisenable,
    input	 	i_phy_12_pipe_RxClk,
    input	 	i_phy_12_pipe_RxValid,
    input	 [39:0]	i_phy_12_pipe_RxData,
    input	 	i_phy_12_pipe_RxElecIdle,
    input	 [2:0]	i_phy_12_pipe_RxStatus,
    input	 	i_phy_12_pipe_RxStandbyStatus,
    output 	o_phy_12_pipe_RxStandby,
    output 	o_phy_12_pipe_RxTermination,
    output [1:0]	o_phy_12_pipe_RxWidth,
    input	 	i_phy_12_pipe_PhyStatus,
    input	 	i_phy_12_pipe_PclkChangeOk,
    output [7:0]	o_phy_12_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_12_pipe_P2M_MessageBus,
    output 	o_phy_13_pipe_TxDataValid,
    output [39:0]	o_phy_13_pipe_TxData,
    output 	o_phy_13_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_13_pipe_TxElecIdle,
    output [3:0]	o_phy_13_pipe_PowerDown,
    output [2:0]	o_phy_13_pipe_Rate,
    output 	o_phy_13_pipe_PclkChangeAck,
    output [2:0]	o_phy_13_pipe_PCLKRate,
    output [1:0]	o_phy_13_pipe_Width,
    output 	o_phy_13_pipe_PCLK,
    output 	o_phy_13_pipe_rxelecidle_disable,
    output 	o_phy_13_pipe_txcmnmode_disable,
    output 	o_phy_13_pipe_srisenable,
    input	 	i_phy_13_pipe_RxClk,
    input	 	i_phy_13_pipe_RxValid,
    input	 [39:0]	i_phy_13_pipe_RxData,
    input	 	i_phy_13_pipe_RxElecIdle,
    input	 [2:0]	i_phy_13_pipe_RxStatus,
    input	 	i_phy_13_pipe_RxStandbyStatus,
    output 	o_phy_13_pipe_RxStandby,
    output 	o_phy_13_pipe_RxTermination,
    output [1:0]	o_phy_13_pipe_RxWidth,
    input	 	i_phy_13_pipe_PhyStatus,
    input	 	i_phy_13_pipe_PclkChangeOk,
    output [7:0]	o_phy_13_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_13_pipe_P2M_MessageBus,
    output 	o_phy_14_pipe_TxDataValid,
    output [39:0]	o_phy_14_pipe_TxData,
    output 	o_phy_14_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_14_pipe_TxElecIdle,
    output [3:0]	o_phy_14_pipe_PowerDown,
    output [2:0]	o_phy_14_pipe_Rate,
    output 	o_phy_14_pipe_PclkChangeAck,
    output [2:0]	o_phy_14_pipe_PCLKRate,
    output [1:0]	o_phy_14_pipe_Width,
    output 	o_phy_14_pipe_PCLK,
    output 	o_phy_14_pipe_rxelecidle_disable,
    output 	o_phy_14_pipe_txcmnmode_disable,
    output 	o_phy_14_pipe_srisenable,
    input	 	i_phy_14_pipe_RxClk,
    input	 	i_phy_14_pipe_RxValid,
    input	 [39:0]	i_phy_14_pipe_RxData,
    input	 	i_phy_14_pipe_RxElecIdle,
    input	 [2:0]	i_phy_14_pipe_RxStatus,
    input	 	i_phy_14_pipe_RxStandbyStatus,
    output 	o_phy_14_pipe_RxStandby,
    output 	o_phy_14_pipe_RxTermination,
    output [1:0]	o_phy_14_pipe_RxWidth,
    input	 	i_phy_14_pipe_PhyStatus,
    input	 	i_phy_14_pipe_PclkChangeOk,
    output [7:0]	o_phy_14_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_14_pipe_P2M_MessageBus,
    output 	o_phy_15_pipe_TxDataValid,
    output [39:0]	o_phy_15_pipe_TxData,
    output 	o_phy_15_pipe_TxDetRxLpbk,
    output [3:0]	o_phy_15_pipe_TxElecIdle,
    output [3:0]	o_phy_15_pipe_PowerDown,
    output [2:0]	o_phy_15_pipe_Rate,
    output 	o_phy_15_pipe_PclkChangeAck,
    output [2:0]	o_phy_15_pipe_PCLKRate,
    output [1:0]	o_phy_15_pipe_Width,
    output 	o_phy_15_pipe_PCLK,
    output 	o_phy_15_pipe_rxelecidle_disable,
    output 	o_phy_15_pipe_txcmnmode_disable,
    output 	o_phy_15_pipe_srisenable,
    input	 	i_phy_15_pipe_RxClk,
    input	 	i_phy_15_pipe_RxValid,
    input	 [39:0]	i_phy_15_pipe_RxData,
    input	 	i_phy_15_pipe_RxElecIdle,
    input	 [2:0]	i_phy_15_pipe_RxStatus,
    input	 	i_phy_15_pipe_RxStandbyStatus,
    output 	o_phy_15_pipe_RxStandby,
    output 	o_phy_15_pipe_RxTermination,
    output [1:0]	o_phy_15_pipe_RxWidth,
    input	 	i_phy_15_pipe_PhyStatus,
    input	 	i_phy_15_pipe_PclkChangeOk,
    output [7:0]	o_phy_15_pipe_M2P_MessageBus,
    input	 [7:0]	i_phy_15_pipe_P2M_MessageBus,
    output	o_phy_0_pipe_rxbitslip_req,
    output [4:0]	o_phy_0_pipe_rxbitslip_va,
    input	 	i_phy_0_pipe_RxBitSlip_Ack,
    output 	o_phy_1_pipe_rxbitslip_req,
    output [4:0]	o_phy_1_pipe_rxbitslip_va,
    input	 	i_phy_1_pipe_RxBitSlip_Ack,
    output 	o_phy_2_pipe_rxbitslip_req,
    output [4:0]	o_phy_2_pipe_rxbitslip_va,
    input	 	i_phy_2_pipe_RxBitSlip_Ack,
    output 	o_phy_3_pipe_rxbitslip_req,
    output [4:0]	o_phy_3_pipe_rxbitslip_va,
    input	 	i_phy_3_pipe_RxBitSlip_Ack,
    output 	o_phy_4_pipe_rxbitslip_req,
    output [4:0]	o_phy_4_pipe_rxbitslip_va,
    input	 	i_phy_4_pipe_RxBitSlip_Ack,
    output 	o_phy_5_pipe_rxbitslip_req,
    output [4:0]	o_phy_5_pipe_rxbitslip_va,
    input	 	i_phy_5_pipe_RxBitSlip_Ack,
    output 	o_phy_6_pipe_rxbitslip_req,
    output [4:0]	o_phy_6_pipe_rxbitslip_va,
    input	 	i_phy_6_pipe_RxBitSlip_Ack,
    output 	o_phy_7_pipe_rxbitslip_req,
    output [4:0]	o_phy_7_pipe_rxbitslip_va,
    input	 	i_phy_7_pipe_RxBitSlip_Ack,
    output 	o_phy_8_pipe_rxbitslip_req,
    output [4:0]	o_phy_8_pipe_rxbitslip_va,
    input	 	i_phy_8_pipe_RxBitSlip_Ack,
    output 	o_phy_9_pipe_rxbitslip_req,
    output [4:0]	o_phy_9_pipe_rxbitslip_va,
    input	 	i_phy_9_pipe_RxBitSlip_Ack,
    output 	o_phy_10_pipe_rxbitslip_req,
    output [4:0]	o_phy_10_pipe_rxbitslip_va,
    input	 	i_phy_10_pipe_RxBitSlip_Ack,
    output 	o_phy_11_pipe_rxbitslip_req,
    output [4:0]	o_phy_11_pipe_rxbitslip_va,
    input	 	i_phy_11_pipe_RxBitSlip_Ack,
    output 	o_phy_12_pipe_rxbitslip_req,
    output [4:0]	o_phy_12_pipe_rxbitslip_va,
    input	 	i_phy_12_pipe_RxBitSlip_Ack,
    output 	o_phy_13_pipe_rxbitslip_req,
    output [4:0]	o_phy_13_pipe_rxbitslip_va,
    input	 	i_phy_13_pipe_RxBitSlip_Ack,
    output 	o_phy_14_pipe_rxbitslip_req,
    output [4:0]	o_phy_14_pipe_rxbitslip_va,
    input	 	i_phy_14_pipe_RxBitSlip_Ack,
    output 	o_phy_15_pipe_rxbitslip_req,
    output [4:0]	o_phy_15_pipe_rxbitslip_va,
    input		i_phy_15_pipe_RxBitSlip_Ack
);

  ////  localparam REVB            = (hssi_ctr_silicon_rev == "10nm6arnrb" || hssi_ctr_silicon_rev == "10nm8arnrb") ? 1 : 0;
localparam REV_B0                  = (hssi_ctr_silicon_rev == "10nm8arnrb" || hssi_ctr_silicon_rev == "10nm7arnrb" || hssi_ctr_silicon_rev == "10nm8parnrb" || hssi_ctr_silicon_rev == "10nm4arnrb") ? 1 : 0;
localparam REV_C0                  = (hssi_ctr_silicon_rev == "10nm4arnrc") ? 1 : 0;

   wire cxl_reset_status_n;
  rnr_cxl_pkg::cxl_cache_mem_rx_intf         cxl_cache_mem_rx_frame0;            // inlcude 3-bit Prot ID
  rnr_cxl_pkg::cxl_cache_mem_rx_intf         cxl_cache_mem_rx_frame1;            // include 3-bit Prot ID
   wire        o_D2H_Data0_CrdRtn;
   wire        o_D2H_Req_CrdRtn;
   wire        o_D2H_Rsp_CrdRtn;
   wire        o_S2M_DRS0_CrdRtn;
   wire        o_S2M_DRS1_CrdRtn;
   wire        o_S2M_NDR_CrdRtn;
   wire        o_D2HPushWrCrdRtn;
   wire        i_H2D_Data0_CrdRtn;
   wire        i_H2D_Data1_CrdRtn;
   wire        i_H2D_Req_CrdRtn;
   wire        i_H2D_Rsp_CrdRtn;
   wire        i_M2S_Req_CrdRtn;
   wire        i_M2S_RwD0_CrdRtn;
   wire        i_M2S_RwD1_CrdRtn;
   wire        i_H2D_Rsp_CrdRtn_fr0;
   wire        i_H2D_Rsp_CrdRtn_fr1;
   wire        i_H2D_Req_CrdRtn_fr0;
   wire        i_H2D_Req_CrdRtn_fr1;
   wire        i_H2D_Data0_CrdRtn_fr0;
   wire        i_H2D_Data0_CrdRtn_fr1;
   wire        i_M2S_RwD0_CrdRtn_fr0;
   wire        i_M2S_RwD0_CrdRtn_fr1;
   wire        i_M2S_Req_CrdRtn_fr0;
   wire        i_M2S_Req_CrdRtn_fr1;

   //------------------------------------CXL Sim Time Reduction start--------------------------------------------------------------//
  
    `define MYZPATH u_rtile_mdx1.u_z1578a_MD.inst_quartus.z1578a
    `ifdef RTILE_PIPE_MODE
    logic phy_sys_ial_0__pipe_Reset_l;
    logic phy_sys_ial_1__pipe_Reset_l;
    logic phy_sys_ial_2__pipe_Reset_l;
    logic phy_sys_ial_3__pipe_Reset_l;
    logic phy_sys_ial_4__pipe_Reset_l;
    logic phy_sys_ial_5__pipe_Reset_l;
    logic phy_sys_ial_6__pipe_Reset_l;
    logic phy_sys_ial_7__pipe_Reset_l;
    logic phy_sys_ial_8__pipe_Reset_l;
    logic phy_sys_ial_9__pipe_Reset_l;
    logic phy_sys_ial_10__pipe_Reset_l;
    logic phy_sys_ial_11__pipe_Reset_l;
    logic phy_sys_ial_12__pipe_Reset_l;
    logic phy_sys_ial_13__pipe_Reset_l;
    logic phy_sys_ial_14__pipe_Reset_l;
    logic phy_sys_ial_15__pipe_Reset_l;	
    logic o_phy_0_pipe_TxDataValid;
    logic [39:0]	o_phy_0_pipe_TxData;
    logic o_phy_0_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_0_pipe_TxElecIdle;
    logic [3:0]	o_phy_0_pipe_PowerDown;
    logic [2:0]	o_phy_0_pipe_Rate;
    logic o_phy_0_pipe_PclkChangeAck;
    logic [2:0]	o_phy_0_pipe_PCLKRate;
    logic [1:0]	o_phy_0_pipe_Width;
    logic o_phy_0_pipe_PCLK;
    logic o_phy_0_pipe_rxelecidle_disable;
    logic o_phy_0_pipe_txcmnmode_disable;
    logic o_phy_0_pipe_srisenable;
    logic i_phy_0_pipe_RxClk;
    logic i_phy_0_pipe_RxValid;
    logic [39:0]	i_phy_0_pipe_RxData;
    logic i_phy_0_pipe_RxElecIdle;
    logic [2:0]	i_phy_0_pipe_RxStatus;
    logic i_phy_0_pipe_RxStandbyStatus;
    logic o_phy_0_pipe_RxStandby;
    logic o_phy_0_pipe_RxTermination;
    logic [1:0]	o_phy_0_pipe_RxWidth;
    logic i_phy_0_pipe_PhyStatus;
    logic i_phy_0_pipe_PclkChangeOk;
    logic [7:0]	o_phy_0_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_0_pipe_P2M_MessageBus;
    logic o_phy_1_pipe_TxDataValid;
    logic [39:0]	o_phy_1_pipe_TxData;
    logic o_phy_1_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_1_pipe_TxElecIdle;
    logic [3:0]	o_phy_1_pipe_PowerDown;
    logic [2:0]	o_phy_1_pipe_Rate;
    logic o_phy_1_pipe_PclkChangeAck;
    logic [2:0]	o_phy_1_pipe_PCLKRate;
    logic [1:0]	o_phy_1_pipe_Width;
    logic o_phy_1_pipe_PCLK;
    logic o_phy_1_pipe_rxelecidle_disable;
    logic o_phy_1_pipe_txcmnmode_disable;
    logic o_phy_1_pipe_srisenable;
    logic i_phy_1_pipe_RxClk;
    logic i_phy_1_pipe_RxValid;
    logic [39:0]	i_phy_1_pipe_RxData;
    logic i_phy_1_pipe_RxElecIdle;
    logic [2:0]	i_phy_1_pipe_RxStatus;
    logic i_phy_1_pipe_RxStandbyStatus;
    logic o_phy_1_pipe_RxStandby;
    logic o_phy_1_pipe_RxTermination;
    logic [1:0]	o_phy_1_pipe_RxWidth;
    logic i_phy_1_pipe_PhyStatus;
    logic i_phy_1_pipe_PclkChangeOk;
    logic [7:0]	o_phy_1_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_1_pipe_P2M_MessageBus;
    logic o_phy_2_pipe_TxDataValid;
    logic [39:0]	o_phy_2_pipe_TxData;
    logic o_phy_2_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_2_pipe_TxElecIdle;
    logic [3:0]	o_phy_2_pipe_PowerDown;
    logic [2:0]	o_phy_2_pipe_Rate;
    logic o_phy_2_pipe_PclkChangeAck;
    logic [2:0]	o_phy_2_pipe_PCLKRate;
    logic [1:0]	o_phy_2_pipe_Width;
    logic o_phy_2_pipe_PCLK;
    logic o_phy_2_pipe_rxelecidle_disable;
    logic o_phy_2_pipe_txcmnmode_disable;
    logic o_phy_2_pipe_srisenable;
    logic i_phy_2_pipe_RxClk;
    logic i_phy_2_pipe_RxValid;
    logic [39:0]	i_phy_2_pipe_RxData;
    logic i_phy_2_pipe_RxElecIdle;
    logic [2:0]	i_phy_2_pipe_RxStatus;
    logic i_phy_2_pipe_RxStandbyStatus;
    logic o_phy_2_pipe_RxStandby;
    logic o_phy_2_pipe_RxTermination;
    logic [1:0]	o_phy_2_pipe_RxWidth;
    logic i_phy_2_pipe_PhyStatus;
    logic i_phy_2_pipe_PclkChangeOk;
    logic [7:0]	o_phy_2_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_2_pipe_P2M_MessageBus;
    logic o_phy_3_pipe_TxDataValid;
    logic [39:0]	o_phy_3_pipe_TxData;
    logic o_phy_3_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_3_pipe_TxElecIdle;
    logic [3:0]	o_phy_3_pipe_PowerDown;
    logic [2:0]	o_phy_3_pipe_Rate;
    logic o_phy_3_pipe_PclkChangeAck;
    logic [2:0]	o_phy_3_pipe_PCLKRate;
    logic [1:0]	o_phy_3_pipe_Width;
    logic o_phy_3_pipe_PCLK;
    logic o_phy_3_pipe_rxelecidle_disable;
    logic o_phy_3_pipe_txcmnmode_disable;
    logic o_phy_3_pipe_srisenable;
    logic i_phy_3_pipe_RxClk;
    logic i_phy_3_pipe_RxValid;
    logic [39:0]	i_phy_3_pipe_RxData;
    logic i_phy_3_pipe_RxElecIdle;
    logic [2:0]	i_phy_3_pipe_RxStatus;
    logic i_phy_3_pipe_RxStandbyStatus;
    logic o_phy_3_pipe_RxStandby;
    logic o_phy_3_pipe_RxTermination;
    logic [1:0]	o_phy_3_pipe_RxWidth;
    logic i_phy_3_pipe_PhyStatus;
    logic i_phy_3_pipe_PclkChangeOk;
    logic [7:0]	o_phy_3_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_3_pipe_P2M_MessageBus;
    logic o_phy_4_pipe_TxDataValid;
    logic [39:0]	o_phy_4_pipe_TxData;
    logic o_phy_4_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_4_pipe_TxElecIdle;
    logic [3:0]	o_phy_4_pipe_PowerDown;
    logic [2:0]	o_phy_4_pipe_Rate;
    logic o_phy_4_pipe_PclkChangeAck;
    logic [2:0]	o_phy_4_pipe_PCLKRate;
    logic [1:0]	o_phy_4_pipe_Width;
    logic o_phy_4_pipe_PCLK;
    logic o_phy_4_pipe_rxelecidle_disable;
    logic o_phy_4_pipe_txcmnmode_disable;
    logic o_phy_4_pipe_srisenable;
    logic i_phy_4_pipe_RxClk;
    logic i_phy_4_pipe_RxValid;
    logic [39:0]	i_phy_4_pipe_RxData;
    logic i_phy_4_pipe_RxElecIdle;
    logic [2:0]	i_phy_4_pipe_RxStatus;
    logic i_phy_4_pipe_RxStandbyStatus;
    logic o_phy_4_pipe_RxStandby;
    logic o_phy_4_pipe_RxTermination;
    logic [1:0]	o_phy_4_pipe_RxWidth;
    logic i_phy_4_pipe_PhyStatus;
    logic i_phy_4_pipe_PclkChangeOk;
    logic [7:0]	o_phy_4_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_4_pipe_P2M_MessageBus;
    logic o_phy_5_pipe_TxDataValid;
    logic [39:0]	o_phy_5_pipe_TxData;
    logic o_phy_5_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_5_pipe_TxElecIdle;
    logic [3:0]	o_phy_5_pipe_PowerDown;
    logic [2:0]	o_phy_5_pipe_Rate;
    logic o_phy_5_pipe_PclkChangeAck;
    logic [2:0]	o_phy_5_pipe_PCLKRate;
    logic [1:0]	o_phy_5_pipe_Width;
    logic o_phy_5_pipe_PCLK;
    logic o_phy_5_pipe_rxelecidle_disable;
    logic o_phy_5_pipe_txcmnmode_disable;
    logic o_phy_5_pipe_srisenable;
    logic i_phy_5_pipe_RxClk;
    logic i_phy_5_pipe_RxValid;
    logic [39:0]	i_phy_5_pipe_RxData;
    logic i_phy_5_pipe_RxElecIdle;
    logic [2:0]	i_phy_5_pipe_RxStatus;
    logic i_phy_5_pipe_RxStandbyStatus;
    logic o_phy_5_pipe_RxStandby;
    logic o_phy_5_pipe_RxTermination;
    logic [1:0]	o_phy_5_pipe_RxWidth;
    logic i_phy_5_pipe_PhyStatus;
    logic i_phy_5_pipe_PclkChangeOk;
    logic [7:0]	o_phy_5_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_5_pipe_P2M_MessageBus;
    logic o_phy_6_pipe_TxDataValid;
    logic [39:0]	o_phy_6_pipe_TxData;
    logic o_phy_6_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_6_pipe_TxElecIdle;
    logic [3:0]	o_phy_6_pipe_PowerDown;
    logic [2:0]	o_phy_6_pipe_Rate;
    logic o_phy_6_pipe_PclkChangeAck;
    logic [2:0]	o_phy_6_pipe_PCLKRate;
    logic [1:0]	o_phy_6_pipe_Width;
    logic o_phy_6_pipe_PCLK;
    logic o_phy_6_pipe_rxelecidle_disable;
    logic o_phy_6_pipe_txcmnmode_disable;
    logic o_phy_6_pipe_srisenable;
    logic i_phy_6_pipe_RxClk;
    logic i_phy_6_pipe_RxValid;
    logic [39:0]	i_phy_6_pipe_RxData;
    logic i_phy_6_pipe_RxElecIdle;
    logic [2:0]	i_phy_6_pipe_RxStatus;
    logic i_phy_6_pipe_RxStandbyStatus;
    logic o_phy_6_pipe_RxStandby;
    logic o_phy_6_pipe_RxTermination;
    logic [1:0]	o_phy_6_pipe_RxWidth;
    logic i_phy_6_pipe_PhyStatus;
    logic i_phy_6_pipe_PclkChangeOk;
    logic [7:0]	o_phy_6_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_6_pipe_P2M_MessageBus;
    logic o_phy_7_pipe_TxDataValid;
    logic [39:0]	o_phy_7_pipe_TxData;
    logic o_phy_7_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_7_pipe_TxElecIdle;
    logic [3:0]	o_phy_7_pipe_PowerDown;
    logic [2:0]	o_phy_7_pipe_Rate;
    logic o_phy_7_pipe_PclkChangeAck;
    logic [2:0]	o_phy_7_pipe_PCLKRate;
    logic [1:0]	o_phy_7_pipe_Width;
    logic o_phy_7_pipe_PCLK;
    logic o_phy_7_pipe_rxelecidle_disable;
    logic o_phy_7_pipe_txcmnmode_disable;
    logic o_phy_7_pipe_srisenable;
    logic i_phy_7_pipe_RxClk;
    logic i_phy_7_pipe_RxValid;
    logic [39:0]	i_phy_7_pipe_RxData;
    logic i_phy_7_pipe_RxElecIdle;
    logic [2:0]	i_phy_7_pipe_RxStatus;
    logic i_phy_7_pipe_RxStandbyStatus;
    logic o_phy_7_pipe_RxStandby;
    logic o_phy_7_pipe_RxTermination;
    logic [1:0]	o_phy_7_pipe_RxWidth;
    logic i_phy_7_pipe_PhyStatus;
    logic i_phy_7_pipe_PclkChangeOk;
    logic [7:0]	o_phy_7_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_7_pipe_P2M_MessageBus;
    logic o_phy_8_pipe_TxDataValid;
    logic [39:0]	o_phy_8_pipe_TxData;
    logic o_phy_8_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_8_pipe_TxElecIdle;
    logic [3:0]	o_phy_8_pipe_PowerDown;
    logic [2:0]	o_phy_8_pipe_Rate;
    logic o_phy_8_pipe_PclkChangeAck;
    logic [2:0]	o_phy_8_pipe_PCLKRate;
    logic [1:0]	o_phy_8_pipe_Width;
    logic o_phy_8_pipe_PCLK;
    logic o_phy_8_pipe_rxelecidle_disable;
    logic o_phy_8_pipe_txcmnmode_disable;
    logic o_phy_8_pipe_srisenable;
    logic i_phy_8_pipe_RxClk;
    logic i_phy_8_pipe_RxValid;
    logic [39:0]	i_phy_8_pipe_RxData;
    logic i_phy_8_pipe_RxElecIdle;
    logic [2:0]	i_phy_8_pipe_RxStatus;
    logic i_phy_8_pipe_RxStandbyStatus;
    logic o_phy_8_pipe_RxStandby;
    logic o_phy_8_pipe_RxTermination;
    logic [1:0]	o_phy_8_pipe_RxWidth;
    logic i_phy_8_pipe_PhyStatus;
    logic i_phy_8_pipe_PclkChangeOk;
    logic [7:0]	o_phy_8_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_8_pipe_P2M_MessageBus;
    logic o_phy_9_pipe_TxDataValid;
    logic [39:0]	o_phy_9_pipe_TxData;
    logic o_phy_9_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_9_pipe_TxElecIdle;
    logic [3:0]	o_phy_9_pipe_PowerDown;
    logic [2:0]	o_phy_9_pipe_Rate;
    logic o_phy_9_pipe_PclkChangeAck;
    logic [2:0]	o_phy_9_pipe_PCLKRate;
    logic [1:0]	o_phy_9_pipe_Width;
    logic o_phy_9_pipe_PCLK;
    logic o_phy_9_pipe_rxelecidle_disable;
    logic o_phy_9_pipe_txcmnmode_disable;
    logic o_phy_9_pipe_srisenable;
    logic i_phy_9_pipe_RxClk;
    logic i_phy_9_pipe_RxValid;
    logic [39:0]	i_phy_9_pipe_RxData;
    logic i_phy_9_pipe_RxElecIdle;
    logic [2:0]	i_phy_9_pipe_RxStatus;
    logic i_phy_9_pipe_RxStandbyStatus;
    logic o_phy_9_pipe_RxStandby;
    logic o_phy_9_pipe_RxTermination;
    logic [1:0]	o_phy_9_pipe_RxWidth;
    logic i_phy_9_pipe_PhyStatus;
    logic i_phy_9_pipe_PclkChangeOk;
    logic [7:0]	o_phy_9_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_9_pipe_P2M_MessageBus;
    logic o_phy_10_pipe_TxDataValid;
    logic [39:0]	o_phy_10_pipe_TxData;
    logic o_phy_10_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_10_pipe_TxElecIdle;
    logic [3:0]	o_phy_10_pipe_PowerDown;
    logic [2:0]	o_phy_10_pipe_Rate;
    logic o_phy_10_pipe_PclkChangeAck;
    logic [2:0]	o_phy_10_pipe_PCLKRate;
    logic [1:0]	o_phy_10_pipe_Width;
    logic o_phy_10_pipe_PCLK;
    logic o_phy_10_pipe_rxelecidle_disable;
    logic o_phy_10_pipe_txcmnmode_disable;
    logic o_phy_10_pipe_srisenable;
    logic i_phy_10_pipe_RxClk;
    logic i_phy_10_pipe_RxValid;
    logic [39:0]	i_phy_10_pipe_RxData;
    logic i_phy_10_pipe_RxElecIdle;
    logic [2:0]	i_phy_10_pipe_RxStatus;
    logic i_phy_10_pipe_RxStandbyStatus;
    logic o_phy_10_pipe_RxStandby;
    logic o_phy_10_pipe_RxTermination;
    logic [1:0]	o_phy_10_pipe_RxWidth;
    logic i_phy_10_pipe_PhyStatus;
    logic i_phy_10_pipe_PclkChangeOk;
    logic [7:0]	o_phy_10_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_10_pipe_P2M_MessageBus;
    logic o_phy_11_pipe_TxDataValid;
    logic [39:0]	o_phy_11_pipe_TxData;
    logic o_phy_11_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_11_pipe_TxElecIdle;
    logic [3:0]	o_phy_11_pipe_PowerDown;
    logic [2:0]	o_phy_11_pipe_Rate;
    logic o_phy_11_pipe_PclkChangeAck;
    logic [2:0]	o_phy_11_pipe_PCLKRate;
    logic [1:0]	o_phy_11_pipe_Width;
    logic o_phy_11_pipe_PCLK;
    logic o_phy_11_pipe_rxelecidle_disable;
    logic o_phy_11_pipe_txcmnmode_disable;
    logic o_phy_11_pipe_srisenable;
    logic i_phy_11_pipe_RxClk;
    logic i_phy_11_pipe_RxValid;
    logic [39:0]	i_phy_11_pipe_RxData;
    logic i_phy_11_pipe_RxElecIdle;
    logic [2:0]	i_phy_11_pipe_RxStatus;
    logic i_phy_11_pipe_RxStandbyStatus;
    logic o_phy_11_pipe_RxStandby;
    logic o_phy_11_pipe_RxTermination;
    logic [1:0]	o_phy_11_pipe_RxWidth;
    logic i_phy_11_pipe_PhyStatus;
    logic i_phy_11_pipe_PclkChangeOk;
    logic [7:0]	o_phy_11_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_11_pipe_P2M_MessageBus;
    logic o_phy_12_pipe_TxDataValid;
    logic [39:0]	o_phy_12_pipe_TxData;
    logic o_phy_12_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_12_pipe_TxElecIdle;
    logic [3:0]	o_phy_12_pipe_PowerDown;
    logic [2:0]	o_phy_12_pipe_Rate;
    logic o_phy_12_pipe_PclkChangeAck;
    logic [2:0]	o_phy_12_pipe_PCLKRate;
    logic [1:0]	o_phy_12_pipe_Width;
    logic o_phy_12_pipe_PCLK;
    logic o_phy_12_pipe_rxelecidle_disable;
    logic o_phy_12_pipe_txcmnmode_disable;
    logic o_phy_12_pipe_srisenable;
    logic i_phy_12_pipe_RxClk;
    logic i_phy_12_pipe_RxValid;
    logic [39:0]	i_phy_12_pipe_RxData;
    logic i_phy_12_pipe_RxElecIdle;
    logic [2:0]	i_phy_12_pipe_RxStatus;
    logic i_phy_12_pipe_RxStandbyStatus;
    logic o_phy_12_pipe_RxStandby;
    logic o_phy_12_pipe_RxTermination;
    logic [1:0]	o_phy_12_pipe_RxWidth;
    logic i_phy_12_pipe_PhyStatus;
    logic i_phy_12_pipe_PclkChangeOk;
    logic [7:0]	o_phy_12_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_12_pipe_P2M_MessageBus;
    logic o_phy_13_pipe_TxDataValid;
    logic [39:0]	o_phy_13_pipe_TxData;
    logic o_phy_13_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_13_pipe_TxElecIdle;
    logic [3:0]	o_phy_13_pipe_PowerDown;
    logic [2:0]	o_phy_13_pipe_Rate;
    logic o_phy_13_pipe_PclkChangeAck;
    logic [2:0]	o_phy_13_pipe_PCLKRate;
    logic [1:0]	o_phy_13_pipe_Width;
    logic o_phy_13_pipe_PCLK;
    logic o_phy_13_pipe_rxelecidle_disable;
    logic o_phy_13_pipe_txcmnmode_disable;
    logic o_phy_13_pipe_srisenable;
    logic i_phy_13_pipe_RxClk;
    logic i_phy_13_pipe_RxValid;
    logic [39:0]	i_phy_13_pipe_RxData;
    logic i_phy_13_pipe_RxElecIdle;
    logic [2:0]	i_phy_13_pipe_RxStatus;
    logic i_phy_13_pipe_RxStandbyStatus;
    logic o_phy_13_pipe_RxStandby;
    logic o_phy_13_pipe_RxTermination;
    logic [1:0]	o_phy_13_pipe_RxWidth;
    logic i_phy_13_pipe_PhyStatus;
    logic i_phy_13_pipe_PclkChangeOk;
    logic [7:0]	o_phy_13_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_13_pipe_P2M_MessageBus;
    logic o_phy_14_pipe_TxDataValid;
    logic [39:0]	o_phy_14_pipe_TxData;
    logic o_phy_14_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_14_pipe_TxElecIdle;
    logic [3:0]	o_phy_14_pipe_PowerDown;
    logic [2:0]	o_phy_14_pipe_Rate;
    logic o_phy_14_pipe_PclkChangeAck;
    logic [2:0]	o_phy_14_pipe_PCLKRate;
    logic [1:0]	o_phy_14_pipe_Width;
    logic o_phy_14_pipe_PCLK;
    logic o_phy_14_pipe_rxelecidle_disable;
    logic o_phy_14_pipe_txcmnmode_disable;
    logic o_phy_14_pipe_srisenable;
    logic i_phy_14_pipe_RxClk;
    logic i_phy_14_pipe_RxValid;
    logic [39:0]	i_phy_14_pipe_RxData;
    logic i_phy_14_pipe_RxElecIdle;
    logic [2:0]	i_phy_14_pipe_RxStatus;
    logic i_phy_14_pipe_RxStandbyStatus;
    logic o_phy_14_pipe_RxStandby;
    logic o_phy_14_pipe_RxTermination;
    logic [1:0]	o_phy_14_pipe_RxWidth;
    logic i_phy_14_pipe_PhyStatus;
    logic i_phy_14_pipe_PclkChangeOk;
    logic [7:0]	o_phy_14_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_14_pipe_P2M_MessageBus;
    logic o_phy_15_pipe_TxDataValid;
    logic [39:0]	o_phy_15_pipe_TxData;
    logic o_phy_15_pipe_TxDetRxLpbk;
    logic [3:0]	o_phy_15_pipe_TxElecIdle;
    logic [3:0]	o_phy_15_pipe_PowerDown;
    logic [2:0]	o_phy_15_pipe_Rate;
    logic o_phy_15_pipe_PclkChangeAck;
    logic [2:0]	o_phy_15_pipe_PCLKRate;
    logic [1:0]	o_phy_15_pipe_Width;
    logic o_phy_15_pipe_PCLK;
    logic o_phy_15_pipe_rxelecidle_disable;
    logic o_phy_15_pipe_txcmnmode_disable;
    logic o_phy_15_pipe_srisenable;
    logic i_phy_15_pipe_RxClk;
    logic i_phy_15_pipe_RxValid;
    logic [39:0]	i_phy_15_pipe_RxData;
    logic i_phy_15_pipe_RxElecIdle;
    logic [2:0]	i_phy_15_pipe_RxStatus;
    logic i_phy_15_pipe_RxStandbyStatus;
    logic o_phy_15_pipe_RxStandby;
    logic o_phy_15_pipe_RxTermination;
    logic [1:0]	o_phy_15_pipe_RxWidth;
    logic i_phy_15_pipe_PhyStatus;
    logic i_phy_15_pipe_PclkChangeOk;
    logic [7:0]	o_phy_15_pipe_M2P_MessageBus;
    logic [7:0]	i_phy_15_pipe_P2M_MessageBus;
    logic o_phy_0_pipe_rxbitslip_req;
    logic [4:0]	o_phy_0_pipe_rxbitslip_va;
    logic i_phy_0_pipe_RxBitSlip_Ack;
    logic o_phy_1_pipe_rxbitslip_req;
    logic [4:0]	o_phy_1_pipe_rxbitslip_va;
    logic i_phy_1_pipe_RxBitSlip_Ack;
    logic o_phy_2_pipe_rxbitslip_req;
    logic [4:0]	o_phy_2_pipe_rxbitslip_va;
    logic i_phy_2_pipe_RxBitSlip_Ack;
    logic o_phy_3_pipe_rxbitslip_req;
    logic [4:0]	o_phy_3_pipe_rxbitslip_va;
    logic i_phy_3_pipe_RxBitSlip_Ack;
    logic o_phy_4_pipe_rxbitslip_req;
    logic [4:0]	o_phy_4_pipe_rxbitslip_va;
    logic i_phy_4_pipe_RxBitSlip_Ack;
    logic o_phy_5_pipe_rxbitslip_req;
    logic [4:0]	o_phy_5_pipe_rxbitslip_va;
    logic i_phy_5_pipe_RxBitSlip_Ack;
    logic o_phy_6_pipe_rxbitslip_req;
    logic [4:0]	o_phy_6_pipe_rxbitslip_va;
    logic i_phy_6_pipe_RxBitSlip_Ack;
    logic o_phy_7_pipe_rxbitslip_req;
    logic [4:0]	o_phy_7_pipe_rxbitslip_va;
    logic i_phy_7_pipe_RxBitSlip_Ack;
    logic o_phy_8_pipe_rxbitslip_req;
    logic [4:0]	o_phy_8_pipe_rxbitslip_va;
    logic i_phy_8_pipe_RxBitSlip_Ack;
    logic o_phy_9_pipe_rxbitslip_req;
    logic [4:0]	o_phy_9_pipe_rxbitslip_va;
    logic i_phy_9_pipe_RxBitSlip_Ack;
    logic o_phy_10_pipe_rxbitslip_req;
    logic [4:0]	o_phy_10_pipe_rxbitslip_va;
    logic i_phy_10_pipe_RxBitSlip_Ack;
    logic o_phy_11_pipe_rxbitslip_req;
    logic [4:0]	o_phy_11_pipe_rxbitslip_va;
    logic i_phy_11_pipe_RxBitSlip_Ack;
    logic o_phy_12_pipe_rxbitslip_req;
    logic [4:0]	o_phy_12_pipe_rxbitslip_va;
    logic i_phy_12_pipe_RxBitSlip_Ack;
    logic o_phy_13_pipe_rxbitslip_req;
    logic [4:0]	o_phy_13_pipe_rxbitslip_va;
    logic i_phy_13_pipe_RxBitSlip_Ack;
    logic o_phy_14_pipe_rxbitslip_req;
    logic [4:0]	o_phy_14_pipe_rxbitslip_va;
    logic i_phy_14_pipe_RxBitSlip_Ack;
    logic o_phy_15_pipe_rxbitslip_req;
    logic [4:0]	o_phy_15_pipe_rxbitslip_va;
    logic i_phy_15_pipe_RxBitSlip_Ack;

    //-------------------------------------------------CXL Sim Time Reduction Assignment---------------------------------------------//
    
    assign phy_sys_ial_0__pipe_Reset_l         =       `MYZPATH.phy_sys_ial_0__pipe_Reset_l;
    assign phy_sys_ial_1__pipe_Reset_l         =       `MYZPATH.phy_sys_ial_1__pipe_Reset_l;
    assign phy_sys_ial_2__pipe_Reset_l         =       `MYZPATH.phy_sys_ial_2__pipe_Reset_l;
    assign phy_sys_ial_3__pipe_Reset_l         =       `MYZPATH.phy_sys_ial_3__pipe_Reset_l;
    assign phy_sys_ial_4__pipe_Reset_l         =       `MYZPATH.phy_sys_ial_4__pipe_Reset_l;
    assign phy_sys_ial_5__pipe_Reset_l         =       `MYZPATH.phy_sys_ial_5__pipe_Reset_l;
    assign phy_sys_ial_6__pipe_Reset_l         =       `MYZPATH.phy_sys_ial_6__pipe_Reset_l;
    assign phy_sys_ial_7__pipe_Reset_l         =       `MYZPATH.phy_sys_ial_7__pipe_Reset_l;
    assign phy_sys_ial_8__pipe_Reset_l         =       `MYZPATH.phy_sys_ial_8__pipe_Reset_l;
    assign phy_sys_ial_9__pipe_Reset_l         =       `MYZPATH.phy_sys_ial_9__pipe_Reset_l;
    assign phy_sys_ial_10__pipe_Reset_l        =       `MYZPATH.phy_sys_ial_10__pipe_Reset_l;
    assign phy_sys_ial_11__pipe_Reset_l        =       `MYZPATH.phy_sys_ial_11__pipe_Reset_l;
    assign phy_sys_ial_12__pipe_Reset_l        =       `MYZPATH.phy_sys_ial_12__pipe_Reset_l;
    assign phy_sys_ial_13__pipe_Reset_l        =       `MYZPATH.phy_sys_ial_13__pipe_Reset_l;
    assign phy_sys_ial_14__pipe_Reset_l        =       `MYZPATH.phy_sys_ial_14__pipe_Reset_l;
    assign phy_sys_ial_15__pipe_Reset_l	       =       `MYZPATH.phy_sys_ial_15__pipe_Reset_l;
    assign o_phy_0_pipe_TxDataValid            =       `MYZPATH.o_phy_0_pipe_TxDataValid;
    assign o_phy_0_pipe_TxData                 =       `MYZPATH.o_phy_0_pipe_TxData;
    assign o_phy_0_pipe_TxDetRxLpbk            =       `MYZPATH.o_phy_0_pipe_TxDetRxLpbk;
    assign o_phy_0_pipe_TxElecIdle             =       `MYZPATH.o_phy_0_pipe_TxElecIdle;
    assign o_phy_0_pipe_PowerDown              =       `MYZPATH.o_phy_0_pipe_PowerDown;
    assign o_phy_0_pipe_Rate                   =       `MYZPATH.o_phy_0_pipe_Rate;
    assign o_phy_0_pipe_PclkChangeAck          =       `MYZPATH.o_phy_0_pipe_PclkChangeAck;
    assign o_phy_0_pipe_PCLKRate               =       `MYZPATH.o_phy_0_pipe_PCLKRate;
    assign o_phy_0_pipe_Width                  =       `MYZPATH.o_phy_0_pipe_Width;
    assign o_phy_0_pipe_PCLK                   =       `MYZPATH.o_phy_0_pipe_PCLK;
    assign o_phy_0_pipe_rxelecidle_disable     =       `MYZPATH.o_phy_0_pipe_rxelecidle_disable;
    assign o_phy_0_pipe_txcmnmode_disable      =       `MYZPATH.o_phy_0_pipe_txcmnmode_disable;
    assign o_phy_0_pipe_srisenable             =       `MYZPATH.o_phy_0_pipe_srisenable;
    assign o_phy_0_pipe_RxStandby              =       `MYZPATH.o_phy_0_pipe_RxStandby;
    assign o_phy_0_pipe_RxTermination          =       `MYZPATH.o_phy_0_pipe_RxTermination;
    assign o_phy_0_pipe_RxWidth                =       `MYZPATH.o_phy_0_pipe_RxWidth;
    assign o_phy_0_pipe_M2P_MessageBus         =       `MYZPATH.o_phy_0_pipe_M2P_MessageBus;
    assign o_phy_1_pipe_TxDataValid            =       `MYZPATH.o_phy_1_pipe_TxDataValid;
    assign o_phy_1_pipe_TxData                 =       `MYZPATH.o_phy_1_pipe_TxData;
    assign o_phy_1_pipe_TxDetRxLpbk            =       `MYZPATH.o_phy_1_pipe_TxDetRxLpbk;
    assign o_phy_1_pipe_TxElecIdle             =       `MYZPATH.o_phy_1_pipe_TxElecIdle;
    assign o_phy_1_pipe_PowerDown              =       `MYZPATH.o_phy_1_pipe_PowerDown;
    assign o_phy_1_pipe_Rate                   =       `MYZPATH.o_phy_1_pipe_Rate;
    assign o_phy_1_pipe_PclkChangeAck          =       `MYZPATH.o_phy_1_pipe_PclkChangeAck;
    assign o_phy_1_pipe_PCLKRate               =       `MYZPATH.o_phy_1_pipe_PCLKRate;
    assign o_phy_1_pipe_Width                  =       `MYZPATH.o_phy_1_pipe_Width;
    assign o_phy_1_pipe_PCLK                   =       `MYZPATH.o_phy_1_pipe_PCLK;
    assign o_phy_1_pipe_rxelecidle_disable     =       `MYZPATH.o_phy_1_pipe_rxelecidle_disable;
    assign o_phy_1_pipe_txcmnmode_disable      =       `MYZPATH.o_phy_1_pipe_txcmnmode_disable;
    assign o_phy_1_pipe_srisenable             =       `MYZPATH.o_phy_1_pipe_srisenable;
    assign o_phy_1_pipe_RxStandby              =       `MYZPATH.o_phy_1_pipe_RxStandby;
    assign o_phy_1_pipe_RxTermination          =       `MYZPATH.o_phy_1_pipe_RxTermination;
    assign o_phy_1_pipe_RxWidth                =       `MYZPATH.o_phy_1_pipe_RxWidth;
    assign o_phy_1_pipe_M2P_MessageBus         =       `MYZPATH.o_phy_1_pipe_M2P_MessageBus;
    assign o_phy_2_pipe_TxDataValid            =       `MYZPATH.o_phy_2_pipe_TxDataValid;
    assign o_phy_2_pipe_TxData                 =       `MYZPATH.o_phy_2_pipe_TxData;
    assign o_phy_2_pipe_TxDetRxLpbk            =       `MYZPATH.o_phy_2_pipe_TxDetRxLpbk;
    assign o_phy_2_pipe_TxElecIdle             =       `MYZPATH.o_phy_2_pipe_TxElecIdle;
    assign o_phy_2_pipe_PowerDown              =       `MYZPATH.o_phy_2_pipe_PowerDown;
    assign o_phy_2_pipe_Rate                   =       `MYZPATH.o_phy_2_pipe_Rate;
    assign o_phy_2_pipe_PclkChangeAck          =       `MYZPATH.o_phy_2_pipe_PclkChangeAck;
    assign o_phy_2_pipe_PCLKRate               =       `MYZPATH.o_phy_2_pipe_PCLKRate;
    assign o_phy_2_pipe_Width                  =       `MYZPATH.o_phy_2_pipe_Width;
    assign o_phy_2_pipe_PCLK                   =       `MYZPATH.o_phy_2_pipe_PCLK;
    assign o_phy_2_pipe_rxelecidle_disable     =       `MYZPATH.o_phy_2_pipe_rxelecidle_disable;
    assign o_phy_2_pipe_txcmnmode_disable      =       `MYZPATH.o_phy_2_pipe_txcmnmode_disable;
    assign o_phy_2_pipe_srisenable             =       `MYZPATH.o_phy_2_pipe_srisenable;
    assign o_phy_2_pipe_RxStandby              =       `MYZPATH.o_phy_2_pipe_RxStandby;
    assign o_phy_2_pipe_RxTermination          =       `MYZPATH.o_phy_2_pipe_RxTermination;
    assign o_phy_2_pipe_RxWidth                =       `MYZPATH.o_phy_2_pipe_RxWidth;
    assign o_phy_2_pipe_M2P_MessageBus         =       `MYZPATH.o_phy_2_pipe_M2P_MessageBus;
    assign o_phy_3_pipe_TxDataValid            =       `MYZPATH.o_phy_3_pipe_TxDataValid;
    assign o_phy_3_pipe_TxData                 =       `MYZPATH.o_phy_3_pipe_TxData;
    assign o_phy_3_pipe_TxDetRxLpbk            =       `MYZPATH.o_phy_3_pipe_TxDetRxLpbk;
    assign o_phy_3_pipe_TxElecIdle             =       `MYZPATH.o_phy_3_pipe_TxElecIdle;
    assign o_phy_3_pipe_PowerDown              =       `MYZPATH.o_phy_3_pipe_PowerDown;
    assign o_phy_3_pipe_Rate                   =       `MYZPATH.o_phy_3_pipe_Rate;
    assign o_phy_3_pipe_PclkChangeAck          =       `MYZPATH.o_phy_3_pipe_PclkChangeAck;
    assign o_phy_3_pipe_PCLKRate               =       `MYZPATH.o_phy_3_pipe_PCLKRate;
    assign o_phy_3_pipe_Width                  =       `MYZPATH.o_phy_3_pipe_Width;
    assign o_phy_3_pipe_PCLK                   =       `MYZPATH.o_phy_3_pipe_PCLK;
    assign o_phy_3_pipe_rxelecidle_disable     =       `MYZPATH.o_phy_3_pipe_rxelecidle_disable;
    assign o_phy_3_pipe_txcmnmode_disable      =       `MYZPATH.o_phy_3_pipe_txcmnmode_disable;
    assign o_phy_3_pipe_srisenable             =       `MYZPATH.o_phy_3_pipe_srisenable;
    assign o_phy_3_pipe_RxStandby              =       `MYZPATH.o_phy_3_pipe_RxStandby;
    assign o_phy_3_pipe_RxTermination          =       `MYZPATH.o_phy_3_pipe_RxTermination;
    assign o_phy_3_pipe_RxWidth                =       `MYZPATH.o_phy_3_pipe_RxWidth;
    assign o_phy_3_pipe_M2P_MessageBus         =       `MYZPATH.o_phy_3_pipe_M2P_MessageBus;
    assign o_phy_4_pipe_TxDataValid            =       `MYZPATH.o_phy_4_pipe_TxDataValid;
    assign o_phy_4_pipe_TxData                 =       `MYZPATH.o_phy_4_pipe_TxData;
    assign o_phy_4_pipe_TxDetRxLpbk            =       `MYZPATH.o_phy_4_pipe_TxDetRxLpbk;
    assign o_phy_4_pipe_TxElecIdle             =       `MYZPATH.o_phy_4_pipe_TxElecIdle;
    assign o_phy_4_pipe_PowerDown              =       `MYZPATH.o_phy_4_pipe_PowerDown;
    assign o_phy_4_pipe_Rate                   =       `MYZPATH.o_phy_4_pipe_Rate;
    assign o_phy_4_pipe_PclkChangeAck          =       `MYZPATH.o_phy_4_pipe_PclkChangeAck;
    assign o_phy_4_pipe_PCLKRate               =       `MYZPATH.o_phy_4_pipe_PCLKRate;
    assign o_phy_4_pipe_Width                  =       `MYZPATH.o_phy_4_pipe_Width;
    assign o_phy_4_pipe_PCLK                   =       `MYZPATH.o_phy_4_pipe_PCLK;
    assign o_phy_4_pipe_rxelecidle_disable     =       `MYZPATH.o_phy_4_pipe_rxelecidle_disable;
    assign o_phy_4_pipe_txcmnmode_disable      =       `MYZPATH.o_phy_4_pipe_txcmnmode_disable;
    assign o_phy_4_pipe_srisenable             =       `MYZPATH.o_phy_4_pipe_srisenable;
    assign o_phy_4_pipe_RxStandby              =       `MYZPATH.o_phy_4_pipe_RxStandby;
    assign o_phy_4_pipe_RxTermination          =       `MYZPATH.o_phy_4_pipe_RxTermination;
    assign o_phy_4_pipe_RxWidth                =       `MYZPATH.o_phy_4_pipe_RxWidth;
    assign o_phy_4_pipe_M2P_MessageBus         =       `MYZPATH.o_phy_4_pipe_M2P_MessageBus;
    assign o_phy_5_pipe_TxDataValid            =       `MYZPATH.o_phy_5_pipe_TxDataValid;
    assign o_phy_5_pipe_TxData                 =       `MYZPATH.o_phy_5_pipe_TxData;
    assign o_phy_5_pipe_TxDetRxLpbk            =       `MYZPATH.o_phy_5_pipe_TxDetRxLpbk;
    assign o_phy_5_pipe_TxElecIdle             =       `MYZPATH.o_phy_5_pipe_TxElecIdle;
    assign o_phy_5_pipe_PowerDown              =       `MYZPATH.o_phy_5_pipe_PowerDown;
    assign o_phy_5_pipe_Rate                   =       `MYZPATH.o_phy_5_pipe_Rate;
    assign o_phy_5_pipe_PclkChangeAck          =       `MYZPATH.o_phy_5_pipe_PclkChangeAck;
    assign o_phy_5_pipe_PCLKRate               =       `MYZPATH.o_phy_5_pipe_PCLKRate;
    assign o_phy_5_pipe_Width                  =       `MYZPATH.o_phy_5_pipe_Width;
    assign o_phy_5_pipe_PCLK                   =       `MYZPATH.o_phy_5_pipe_PCLK;
    assign o_phy_5_pipe_rxelecidle_disable     =       `MYZPATH.o_phy_5_pipe_rxelecidle_disable;
    assign o_phy_5_pipe_txcmnmode_disable      =       `MYZPATH.o_phy_5_pipe_txcmnmode_disable;
    assign o_phy_5_pipe_srisenable             =       `MYZPATH.o_phy_5_pipe_srisenable;
    assign o_phy_5_pipe_RxStandby              =       `MYZPATH.o_phy_5_pipe_RxStandby;
    assign o_phy_5_pipe_RxTermination          =       `MYZPATH.o_phy_5_pipe_RxTermination;
    assign o_phy_5_pipe_RxWidth                =       `MYZPATH.o_phy_5_pipe_RxWidth;
    assign o_phy_5_pipe_M2P_MessageBus         =       `MYZPATH.o_phy_5_pipe_M2P_MessageBus;
    assign o_phy_6_pipe_TxDataValid            =       `MYZPATH.o_phy_6_pipe_TxDataValid;
    assign o_phy_6_pipe_TxData                 =       `MYZPATH.o_phy_6_pipe_TxData;
    assign o_phy_6_pipe_TxDetRxLpbk            =       `MYZPATH.o_phy_6_pipe_TxDetRxLpbk;
    assign o_phy_6_pipe_TxElecIdle             =       `MYZPATH.o_phy_6_pipe_TxElecIdle;
    assign o_phy_6_pipe_PowerDown              =       `MYZPATH.o_phy_6_pipe_PowerDown;
    assign o_phy_6_pipe_Rate                   =       `MYZPATH.o_phy_6_pipe_Rate;
    assign o_phy_6_pipe_PclkChangeAck          =       `MYZPATH.o_phy_6_pipe_PclkChangeAck;
    assign o_phy_6_pipe_PCLKRate               =       `MYZPATH.o_phy_6_pipe_PCLKRate;
    assign o_phy_6_pipe_Width                  =       `MYZPATH.o_phy_6_pipe_Width;
    assign o_phy_6_pipe_PCLK                   =       `MYZPATH.o_phy_6_pipe_PCLK;
    assign o_phy_6_pipe_rxelecidle_disable     =       `MYZPATH.o_phy_6_pipe_rxelecidle_disable;
    assign o_phy_6_pipe_txcmnmode_disable      =       `MYZPATH.o_phy_6_pipe_txcmnmode_disable;
    assign o_phy_6_pipe_srisenable             =       `MYZPATH.o_phy_6_pipe_srisenable;
    assign o_phy_6_pipe_RxStandby              =       `MYZPATH.o_phy_6_pipe_RxStandby;
    assign o_phy_6_pipe_RxTermination          =       `MYZPATH.o_phy_6_pipe_RxTermination;
    assign o_phy_6_pipe_RxWidth                =       `MYZPATH.o_phy_6_pipe_RxWidth;
    assign o_phy_6_pipe_M2P_MessageBus         =       `MYZPATH.o_phy_6_pipe_M2P_MessageBus;
    assign o_phy_7_pipe_TxDataValid            =       `MYZPATH.o_phy_7_pipe_TxDataValid;
    assign o_phy_7_pipe_TxData                 =       `MYZPATH.o_phy_7_pipe_TxData;
    assign o_phy_7_pipe_TxDetRxLpbk            =       `MYZPATH.o_phy_7_pipe_TxDetRxLpbk;
    assign o_phy_7_pipe_TxElecIdle             =       `MYZPATH.o_phy_7_pipe_TxElecIdle;
    assign o_phy_7_pipe_PowerDown              =       `MYZPATH.o_phy_7_pipe_PowerDown;
    assign o_phy_7_pipe_Rate                   =       `MYZPATH.o_phy_7_pipe_Rate;
    assign o_phy_7_pipe_PclkChangeAck          =       `MYZPATH.o_phy_7_pipe_PclkChangeAck;
    assign o_phy_7_pipe_PCLKRate               =       `MYZPATH.o_phy_7_pipe_PCLKRate;
    assign o_phy_7_pipe_Width                  =       `MYZPATH.o_phy_7_pipe_Width;
    assign o_phy_7_pipe_PCLK                   =       `MYZPATH.o_phy_7_pipe_PCLK;
    assign o_phy_7_pipe_rxelecidle_disable     =       `MYZPATH.o_phy_7_pipe_rxelecidle_disable;
    assign o_phy_7_pipe_txcmnmode_disable      =       `MYZPATH.o_phy_7_pipe_txcmnmode_disable;
    assign o_phy_7_pipe_srisenable             =       `MYZPATH.o_phy_7_pipe_srisenable;
    assign o_phy_7_pipe_RxStandby              =       `MYZPATH.o_phy_7_pipe_RxStandby;
    assign o_phy_7_pipe_RxTermination          =       `MYZPATH.o_phy_7_pipe_RxTermination;
    assign o_phy_7_pipe_RxWidth                =       `MYZPATH.o_phy_7_pipe_RxWidth;
    assign o_phy_7_pipe_M2P_MessageBus         =       `MYZPATH.o_phy_7_pipe_M2P_MessageBus;
    assign o_phy_8_pipe_TxDataValid            =       `MYZPATH.o_phy_8_pipe_TxDataValid;
    assign o_phy_8_pipe_TxData                 =       `MYZPATH.o_phy_8_pipe_TxData;
    assign o_phy_8_pipe_TxDetRxLpbk            =       `MYZPATH.o_phy_8_pipe_TxDetRxLpbk;
    assign o_phy_8_pipe_TxElecIdle             =       `MYZPATH.o_phy_8_pipe_TxElecIdle;
    assign o_phy_8_pipe_PowerDown              =       `MYZPATH.o_phy_8_pipe_PowerDown;
    assign o_phy_8_pipe_Rate                   =       `MYZPATH.o_phy_8_pipe_Rate;
    assign o_phy_8_pipe_PclkChangeAck          =       `MYZPATH.o_phy_8_pipe_PclkChangeAck;
    assign o_phy_8_pipe_PCLKRate               =       `MYZPATH.o_phy_8_pipe_PCLKRate;
    assign o_phy_8_pipe_Width                  =       `MYZPATH.o_phy_8_pipe_Width;
    assign o_phy_8_pipe_PCLK                   =       `MYZPATH.o_phy_8_pipe_PCLK;
    assign o_phy_8_pipe_rxelecidle_disable     =       `MYZPATH.o_phy_8_pipe_rxelecidle_disable;
    assign o_phy_8_pipe_txcmnmode_disable      =       `MYZPATH.o_phy_8_pipe_txcmnmode_disable;
    assign o_phy_8_pipe_srisenable             =       `MYZPATH.o_phy_8_pipe_srisenable;
    assign o_phy_8_pipe_RxStandby              =       `MYZPATH.o_phy_8_pipe_RxStandby;
    assign o_phy_8_pipe_RxTermination          =       `MYZPATH.o_phy_8_pipe_RxTermination;
    assign o_phy_8_pipe_RxWidth                =       `MYZPATH.o_phy_8_pipe_RxWidth;
    assign o_phy_8_pipe_M2P_MessageBus         =       `MYZPATH.o_phy_8_pipe_M2P_MessageBus;
    assign o_phy_9_pipe_TxDataValid            =       `MYZPATH.o_phy_9_pipe_TxDataValid;
    assign o_phy_9_pipe_TxData                 =       `MYZPATH.o_phy_9_pipe_TxData;
    assign o_phy_9_pipe_TxDetRxLpbk            =       `MYZPATH.o_phy_9_pipe_TxDetRxLpbk;
    assign o_phy_9_pipe_TxElecIdle             =       `MYZPATH.o_phy_9_pipe_TxElecIdle;
    assign o_phy_9_pipe_PowerDown              =       `MYZPATH.o_phy_9_pipe_PowerDown;
    assign o_phy_9_pipe_Rate                   =       `MYZPATH.o_phy_9_pipe_Rate;
    assign o_phy_9_pipe_PclkChangeAck          =       `MYZPATH.o_phy_9_pipe_PclkChangeAck;
    assign o_phy_9_pipe_PCLKRate               =       `MYZPATH.o_phy_9_pipe_PCLKRate;
    assign o_phy_9_pipe_Width                  =       `MYZPATH.o_phy_9_pipe_Width;
    assign o_phy_9_pipe_PCLK                   =       `MYZPATH.o_phy_9_pipe_PCLK;
    assign o_phy_9_pipe_rxelecidle_disable     =       `MYZPATH.o_phy_9_pipe_rxelecidle_disable;
    assign o_phy_9_pipe_txcmnmode_disable      =       `MYZPATH.o_phy_9_pipe_txcmnmode_disable;
    assign o_phy_9_pipe_srisenable             =       `MYZPATH.o_phy_9_pipe_srisenable;
    assign o_phy_9_pipe_RxStandby              =       `MYZPATH.o_phy_9_pipe_RxStandby;
    assign o_phy_9_pipe_RxTermination          =       `MYZPATH.o_phy_9_pipe_RxTermination;
    assign o_phy_9_pipe_RxWidth                =       `MYZPATH.o_phy_9_pipe_RxWidth;
    assign o_phy_9_pipe_M2P_MessageBus         =       `MYZPATH.o_phy_9_pipe_M2P_MessageBus;
    assign o_phy_10_pipe_TxDataValid           =       `MYZPATH.o_phy_10_pipe_TxDataValid;
    assign o_phy_10_pipe_TxData                =       `MYZPATH.o_phy_10_pipe_TxData;
    assign o_phy_10_pipe_TxDetRxLpbk           =       `MYZPATH.o_phy_10_pipe_TxDetRxLpbk;
    assign o_phy_10_pipe_TxElecIdle            =       `MYZPATH.o_phy_10_pipe_TxElecIdle;
    assign o_phy_10_pipe_PowerDown             =       `MYZPATH.o_phy_10_pipe_PowerDown;
    assign o_phy_10_pipe_Rate                  =       `MYZPATH.o_phy_10_pipe_Rate;
    assign o_phy_10_pipe_PclkChangeAck         =       `MYZPATH.o_phy_10_pipe_PclkChangeAck;
    assign o_phy_10_pipe_PCLKRate              =       `MYZPATH.o_phy_10_pipe_PCLKRate;
    assign o_phy_10_pipe_Width                 =       `MYZPATH.o_phy_10_pipe_Width;
    assign o_phy_10_pipe_PCLK                  =       `MYZPATH.o_phy_10_pipe_PCLK;
    assign o_phy_10_pipe_rxelecidle_disable    =       `MYZPATH.o_phy_10_pipe_rxelecidle_disable;
    assign o_phy_10_pipe_txcmnmode_disable     =       `MYZPATH.o_phy_10_pipe_txcmnmode_disable;
    assign o_phy_10_pipe_srisenable            =       `MYZPATH.o_phy_10_pipe_srisenable;
    assign o_phy_10_pipe_RxStandby             =       `MYZPATH.o_phy_10_pipe_RxStandby;
    assign o_phy_10_pipe_RxTermination         =       `MYZPATH.o_phy_10_pipe_RxTermination;
    assign o_phy_10_pipe_RxWidth               =       `MYZPATH.o_phy_10_pipe_RxWidth;
    assign o_phy_10_pipe_M2P_MessageBus        =       `MYZPATH.o_phy_10_pipe_M2P_MessageBus;
    assign o_phy_11_pipe_TxDataValid           =       `MYZPATH.o_phy_11_pipe_TxDataValid;
    assign o_phy_11_pipe_TxData                =       `MYZPATH.o_phy_11_pipe_TxData;
    assign o_phy_11_pipe_TxDetRxLpbk           =       `MYZPATH.o_phy_11_pipe_TxDetRxLpbk;
    assign o_phy_11_pipe_TxElecIdle            =       `MYZPATH.o_phy_11_pipe_TxElecIdle;
    assign o_phy_11_pipe_PowerDown             =       `MYZPATH.o_phy_11_pipe_PowerDown;
    assign o_phy_11_pipe_Rate                  =       `MYZPATH.o_phy_11_pipe_Rate;
    assign o_phy_11_pipe_PclkChangeAck         =       `MYZPATH.o_phy_11_pipe_PclkChangeAck;
    assign o_phy_11_pipe_PCLKRate              =       `MYZPATH.o_phy_11_pipe_PCLKRate;
    assign o_phy_11_pipe_Width                 =       `MYZPATH.o_phy_11_pipe_Width;
    assign o_phy_11_pipe_PCLK                  =       `MYZPATH.o_phy_11_pipe_PCLK;
    assign o_phy_11_pipe_rxelecidle_disable    =       `MYZPATH.o_phy_11_pipe_rxelecidle_disable;
    assign o_phy_11_pipe_txcmnmode_disable     =       `MYZPATH.o_phy_11_pipe_txcmnmode_disable;
    assign o_phy_11_pipe_srisenable            =       `MYZPATH.o_phy_11_pipe_srisenable;
    assign o_phy_11_pipe_RxStandby             =       `MYZPATH.o_phy_11_pipe_RxStandby;
    assign o_phy_11_pipe_RxTermination         =       `MYZPATH.o_phy_11_pipe_RxTermination;
    assign o_phy_11_pipe_RxWidth               =       `MYZPATH.o_phy_11_pipe_RxWidth;
    assign o_phy_11_pipe_M2P_MessageBus        =       `MYZPATH.o_phy_11_pipe_M2P_MessageBus;
    assign o_phy_12_pipe_TxDataValid           =       `MYZPATH.o_phy_12_pipe_TxDataValid;
    assign o_phy_12_pipe_TxData                =       `MYZPATH.o_phy_12_pipe_TxData;
    assign o_phy_12_pipe_TxDetRxLpbk           =       `MYZPATH.o_phy_12_pipe_TxDetRxLpbk;
    assign o_phy_12_pipe_TxElecIdle            =       `MYZPATH.o_phy_12_pipe_TxElecIdle;
    assign o_phy_12_pipe_PowerDown             =       `MYZPATH.o_phy_12_pipe_PowerDown;
    assign o_phy_12_pipe_Rate                  =       `MYZPATH.o_phy_12_pipe_Rate;
    assign o_phy_12_pipe_PclkChangeAck         =       `MYZPATH.o_phy_12_pipe_PclkChangeAck;
    assign o_phy_12_pipe_PCLKRate              =       `MYZPATH.o_phy_12_pipe_PCLKRate;
    assign o_phy_12_pipe_Width                 =       `MYZPATH.o_phy_12_pipe_Width;
    assign o_phy_12_pipe_PCLK                  =       `MYZPATH.o_phy_12_pipe_PCLK;
    assign o_phy_12_pipe_rxelecidle_disable    =       `MYZPATH.o_phy_12_pipe_rxelecidle_disable;
    assign o_phy_12_pipe_txcmnmode_disable     =       `MYZPATH.o_phy_12_pipe_txcmnmode_disable;
    assign o_phy_12_pipe_srisenable            =       `MYZPATH.o_phy_12_pipe_srisenable;
    assign o_phy_12_pipe_RxStandby             =       `MYZPATH.o_phy_12_pipe_RxStandby;
    assign o_phy_12_pipe_RxTermination         =       `MYZPATH.o_phy_12_pipe_RxTermination;
    assign o_phy_12_pipe_RxWidth               =       `MYZPATH.o_phy_12_pipe_RxWidth;
    assign o_phy_12_pipe_M2P_MessageBus        =       `MYZPATH.o_phy_12_pipe_M2P_MessageBus;
    assign o_phy_13_pipe_TxDataValid           =       `MYZPATH.o_phy_13_pipe_TxDataValid;
    assign o_phy_13_pipe_TxData                =       `MYZPATH.o_phy_13_pipe_TxData;
    assign o_phy_13_pipe_TxDetRxLpbk           =       `MYZPATH.o_phy_13_pipe_TxDetRxLpbk;
    assign o_phy_13_pipe_TxElecIdle            =       `MYZPATH.o_phy_13_pipe_TxElecIdle;
    assign o_phy_13_pipe_PowerDown             =       `MYZPATH.o_phy_13_pipe_PowerDown;
    assign o_phy_13_pipe_Rate                  =       `MYZPATH.o_phy_13_pipe_Rate;
    assign o_phy_13_pipe_PclkChangeAck         =       `MYZPATH.o_phy_13_pipe_PclkChangeAck;
    assign o_phy_13_pipe_PCLKRate              =       `MYZPATH.o_phy_13_pipe_PCLKRate;
    assign o_phy_13_pipe_Width                 =       `MYZPATH.o_phy_13_pipe_Width;
    assign o_phy_13_pipe_PCLK                  =       `MYZPATH.o_phy_13_pipe_PCLK;
    assign o_phy_13_pipe_rxelecidle_disable    =       `MYZPATH.o_phy_13_pipe_rxelecidle_disable;
    assign o_phy_13_pipe_txcmnmode_disable     =       `MYZPATH.o_phy_13_pipe_txcmnmode_disable;
    assign o_phy_13_pipe_srisenable            =       `MYZPATH.o_phy_13_pipe_srisenable;
    assign o_phy_13_pipe_RxStandby             =       `MYZPATH.o_phy_13_pipe_RxStandby;
    assign o_phy_13_pipe_RxTermination         =       `MYZPATH.o_phy_13_pipe_RxTermination;
    assign o_phy_13_pipe_RxWidth               =       `MYZPATH.o_phy_13_pipe_RxWidth;
    assign o_phy_13_pipe_M2P_MessageBus        =       `MYZPATH.o_phy_13_pipe_M2P_MessageBus;
    assign o_phy_14_pipe_TxDataValid           =       `MYZPATH.o_phy_14_pipe_TxDataValid;
    assign o_phy_14_pipe_TxData                =       `MYZPATH.o_phy_14_pipe_TxData;
    assign o_phy_14_pipe_TxDetRxLpbk           =       `MYZPATH.o_phy_14_pipe_TxDetRxLpbk;
    assign o_phy_14_pipe_TxElecIdle            =       `MYZPATH.o_phy_14_pipe_TxElecIdle;
    assign o_phy_14_pipe_PowerDown             =       `MYZPATH.o_phy_14_pipe_PowerDown;
    assign o_phy_14_pipe_Rate                  =       `MYZPATH.o_phy_14_pipe_Rate;
    assign o_phy_14_pipe_PclkChangeAck         =       `MYZPATH.o_phy_14_pipe_PclkChangeAck;
    assign o_phy_14_pipe_PCLKRate              =       `MYZPATH.o_phy_14_pipe_PCLKRate;
    assign o_phy_14_pipe_Width                 =       `MYZPATH.o_phy_14_pipe_Width;
    assign o_phy_14_pipe_PCLK                  =       `MYZPATH.o_phy_14_pipe_PCLK;
    assign o_phy_14_pipe_rxelecidle_disable    =       `MYZPATH.o_phy_14_pipe_rxelecidle_disable;
    assign o_phy_14_pipe_txcmnmode_disable     =       `MYZPATH.o_phy_14_pipe_txcmnmode_disable;
    assign o_phy_14_pipe_srisenable            =       `MYZPATH.o_phy_14_pipe_srisenable;
    assign o_phy_14_pipe_RxStandby             =       `MYZPATH.o_phy_14_pipe_RxStandby;
    assign o_phy_14_pipe_RxTermination         =       `MYZPATH.o_phy_14_pipe_RxTermination;
    assign o_phy_14_pipe_RxWidth               =       `MYZPATH.o_phy_14_pipe_RxWidth;
    assign o_phy_14_pipe_M2P_MessageBus        =       `MYZPATH.o_phy_14_pipe_M2P_MessageBus;
    assign o_phy_15_pipe_TxDataValid           =       `MYZPATH.o_phy_15_pipe_TxDataValid;
    assign o_phy_15_pipe_TxData                =       `MYZPATH.o_phy_15_pipe_TxData;
    assign o_phy_15_pipe_TxDetRxLpbk           =       `MYZPATH.o_phy_15_pipe_TxDetRxLpbk;
    assign o_phy_15_pipe_TxElecIdle            =       `MYZPATH.o_phy_15_pipe_TxElecIdle;
    assign o_phy_15_pipe_PowerDown             =       `MYZPATH.o_phy_15_pipe_PowerDown;
    assign o_phy_15_pipe_Rate                  =       `MYZPATH.o_phy_15_pipe_Rate;
    assign o_phy_15_pipe_PclkChangeAck         =       `MYZPATH.o_phy_15_pipe_PclkChangeAck;
    assign o_phy_15_pipe_PCLKRate              =       `MYZPATH.o_phy_15_pipe_PCLKRate;
    assign o_phy_15_pipe_Width                 =       `MYZPATH.o_phy_15_pipe_Width;
    assign o_phy_15_pipe_PCLK                  =       `MYZPATH.o_phy_15_pipe_PCLK;
    assign o_phy_15_pipe_rxelecidle_disable    =       `MYZPATH.o_phy_15_pipe_rxelecidle_disable;
    assign o_phy_15_pipe_txcmnmode_disable     =       `MYZPATH.o_phy_15_pipe_txcmnmode_disable;
    assign o_phy_15_pipe_srisenable            =       `MYZPATH.o_phy_15_pipe_srisenable;
    assign o_phy_15_pipe_RxStandby             =       `MYZPATH.o_phy_15_pipe_RxStandby;
    assign o_phy_15_pipe_RxTermination         =       `MYZPATH.o_phy_15_pipe_RxTermination;
    assign o_phy_15_pipe_RxWidth               =       `MYZPATH.o_phy_15_pipe_RxWidth;
    assign o_phy_15_pipe_M2P_MessageBus        =       `MYZPATH.o_phy_15_pipe_M2P_MessageBus;
    assign o_phy_0_pipe_rxbitslip_req          =       `MYZPATH.o_phy_0_pipe_rxbitslip_req;
    assign o_phy_0_pipe_rxbitslip_va           =       `MYZPATH.o_phy_0_pipe_rxbitslip_va;
    assign o_phy_1_pipe_rxbitslip_req          =       `MYZPATH.o_phy_1_pipe_rxbitslip_req;
    assign o_phy_1_pipe_rxbitslip_va           =       `MYZPATH.o_phy_1_pipe_rxbitslip_va;
    assign o_phy_2_pipe_rxbitslip_req          =       `MYZPATH.o_phy_2_pipe_rxbitslip_req;
    assign o_phy_2_pipe_rxbitslip_va           =       `MYZPATH.o_phy_2_pipe_rxbitslip_va;
    assign o_phy_3_pipe_rxbitslip_req          =       `MYZPATH.o_phy_3_pipe_rxbitslip_req;
    assign o_phy_3_pipe_rxbitslip_va           =       `MYZPATH.o_phy_3_pipe_rxbitslip_va;
    assign o_phy_4_pipe_rxbitslip_req          =       `MYZPATH.o_phy_4_pipe_rxbitslip_req;
    assign o_phy_4_pipe_rxbitslip_va           =       `MYZPATH.o_phy_4_pipe_rxbitslip_va;
    assign o_phy_5_pipe_rxbitslip_req          =       `MYZPATH.o_phy_5_pipe_rxbitslip_req;
    assign o_phy_5_pipe_rxbitslip_va           =       `MYZPATH.o_phy_5_pipe_rxbitslip_va;
    assign o_phy_6_pipe_rxbitslip_req          =       `MYZPATH.o_phy_6_pipe_rxbitslip_req;
    assign o_phy_6_pipe_rxbitslip_va           =       `MYZPATH.o_phy_6_pipe_rxbitslip_va;
    assign o_phy_7_pipe_rxbitslip_req          =       `MYZPATH.o_phy_7_pipe_rxbitslip_req;
    assign o_phy_7_pipe_rxbitslip_va           =       `MYZPATH.o_phy_7_pipe_rxbitslip_va;
    assign o_phy_8_pipe_rxbitslip_req          =       `MYZPATH.o_phy_8_pipe_rxbitslip_req;
    assign o_phy_8_pipe_rxbitslip_va           =       `MYZPATH.o_phy_8_pipe_rxbitslip_va;
    assign o_phy_9_pipe_rxbitslip_req          =       `MYZPATH.o_phy_9_pipe_rxbitslip_req;
    assign o_phy_9_pipe_rxbitslip_va           =       `MYZPATH.o_phy_9_pipe_rxbitslip_va;
    assign o_phy_10_pipe_rxbitslip_req         =       `MYZPATH.o_phy_10_pipe_rxbitslip_req;
    assign o_phy_10_pipe_rxbitslip_va          =       `MYZPATH.o_phy_10_pipe_rxbitslip_va;
    assign o_phy_11_pipe_rxbitslip_req         =       `MYZPATH.o_phy_11_pipe_rxbitslip_req;
    assign o_phy_11_pipe_rxbitslip_va          =       `MYZPATH.o_phy_11_pipe_rxbitslip_va;
    assign o_phy_12_pipe_rxbitslip_req         =       `MYZPATH.o_phy_12_pipe_rxbitslip_req;
    assign o_phy_12_pipe_rxbitslip_va          =       `MYZPATH.o_phy_12_pipe_rxbitslip_va;
    assign o_phy_13_pipe_rxbitslip_req         =       `MYZPATH.o_phy_13_pipe_rxbitslip_req;
    assign o_phy_13_pipe_rxbitslip_va          =       `MYZPATH.o_phy_13_pipe_rxbitslip_va;
    assign o_phy_14_pipe_rxbitslip_req         =       `MYZPATH.o_phy_14_pipe_rxbitslip_req;
    assign o_phy_14_pipe_rxbitslip_va          =       `MYZPATH.o_phy_14_pipe_rxbitslip_va;
    assign o_phy_15_pipe_rxbitslip_req         =       `MYZPATH.o_phy_15_pipe_rxbitslip_req;
    assign o_phy_15_pipe_rxbitslip_va          =       `MYZPATH.o_phy_15_pipe_rxbitslip_va;
    assign `MYZPATH.i_phy_0_pipe_RxClk                  =       i_phy_0_pipe_RxClk;
    assign `MYZPATH.i_phy_0_pipe_RxValid                =       i_phy_0_pipe_RxValid;
    assign `MYZPATH.i_phy_0_pipe_RxData                 =       i_phy_0_pipe_RxData;
    assign `MYZPATH.i_phy_0_pipe_RxElecIdle             =       i_phy_0_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_0_pipe_RxStatus               =       i_phy_0_pipe_RxStatus;
    assign `MYZPATH.i_phy_0_pipe_RxStandbyStatus        =       i_phy_0_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_0_pipe_PhyStatus              =       i_phy_0_pipe_PhyStatus;
    assign `MYZPATH.i_phy_0_pipe_PclkChangeOk           =       i_phy_0_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_0_pipe_P2M_MessageBus         =       i_phy_0_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_1_pipe_RxClk                  =       i_phy_1_pipe_RxClk;
    assign `MYZPATH.i_phy_1_pipe_RxValid                =       i_phy_1_pipe_RxValid;
    assign `MYZPATH.i_phy_1_pipe_RxData                 =       i_phy_1_pipe_RxData;
    assign `MYZPATH.i_phy_1_pipe_RxElecIdle             =       i_phy_1_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_1_pipe_RxStatus               =       i_phy_1_pipe_RxStatus;
    assign `MYZPATH.i_phy_1_pipe_RxStandbyStatus        =       i_phy_1_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_1_pipe_PhyStatus              =       i_phy_1_pipe_PhyStatus;
    assign `MYZPATH.i_phy_1_pipe_PclkChangeOk           =       i_phy_1_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_1_pipe_P2M_MessageBus         =       i_phy_1_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_2_pipe_RxClk                  =       i_phy_2_pipe_RxClk;
    assign `MYZPATH.i_phy_2_pipe_RxValid                =       i_phy_2_pipe_RxValid;
    assign `MYZPATH.i_phy_2_pipe_RxData                 =       i_phy_2_pipe_RxData;
    assign `MYZPATH.i_phy_2_pipe_RxElecIdle             =       i_phy_2_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_2_pipe_RxStatus               =       i_phy_2_pipe_RxStatus;
    assign `MYZPATH.i_phy_2_pipe_RxStandbyStatus        =       i_phy_2_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_2_pipe_PhyStatus              =       i_phy_2_pipe_PhyStatus;
    assign `MYZPATH.i_phy_2_pipe_PclkChangeOk           =       i_phy_2_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_2_pipe_P2M_MessageBus         =       i_phy_2_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_3_pipe_RxClk                  =       i_phy_3_pipe_RxClk;
    assign `MYZPATH.i_phy_3_pipe_RxValid                =       i_phy_3_pipe_RxValid;
    assign `MYZPATH.i_phy_3_pipe_RxData                 =       i_phy_3_pipe_RxData;
    assign `MYZPATH.i_phy_3_pipe_RxElecIdle             =       i_phy_3_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_3_pipe_RxStatus               =       i_phy_3_pipe_RxStatus;
    assign `MYZPATH.i_phy_3_pipe_RxStandbyStatus        =       i_phy_3_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_3_pipe_PhyStatus              =       i_phy_3_pipe_PhyStatus;
    assign `MYZPATH.i_phy_3_pipe_PclkChangeOk           =       i_phy_3_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_3_pipe_P2M_MessageBus         =       i_phy_3_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_4_pipe_RxClk                  =       i_phy_4_pipe_RxClk;
    assign `MYZPATH.i_phy_4_pipe_RxValid                =       i_phy_4_pipe_RxValid;
    assign `MYZPATH.i_phy_4_pipe_RxData                 =       i_phy_4_pipe_RxData;
    assign `MYZPATH.i_phy_4_pipe_RxElecIdle             =       i_phy_4_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_4_pipe_RxStatus               =       i_phy_4_pipe_RxStatus;
    assign `MYZPATH.i_phy_4_pipe_RxStandbyStatus        =       i_phy_4_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_4_pipe_PhyStatus              =       i_phy_4_pipe_PhyStatus;
    assign `MYZPATH.i_phy_4_pipe_PclkChangeOk           =       i_phy_4_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_4_pipe_P2M_MessageBus         =       i_phy_4_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_5_pipe_RxClk                  =       i_phy_5_pipe_RxClk;
    assign `MYZPATH.i_phy_5_pipe_RxValid                =       i_phy_5_pipe_RxValid;
    assign `MYZPATH.i_phy_5_pipe_RxData                 =       i_phy_5_pipe_RxData;
    assign `MYZPATH.i_phy_5_pipe_RxElecIdle             =       i_phy_5_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_5_pipe_RxStatus               =       i_phy_5_pipe_RxStatus;
    assign `MYZPATH.i_phy_5_pipe_RxStandbyStatus        =       i_phy_5_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_5_pipe_PhyStatus              =       i_phy_5_pipe_PhyStatus;
    assign `MYZPATH.i_phy_5_pipe_PclkChangeOk           =       i_phy_5_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_5_pipe_P2M_MessageBus         =       i_phy_5_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_6_pipe_RxClk                  =       i_phy_6_pipe_RxClk;
    assign `MYZPATH.i_phy_6_pipe_RxValid                =       i_phy_6_pipe_RxValid;
    assign `MYZPATH.i_phy_6_pipe_RxData                 =       i_phy_6_pipe_RxData;
    assign `MYZPATH.i_phy_6_pipe_RxElecIdle             =       i_phy_6_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_6_pipe_RxStatus               =       i_phy_6_pipe_RxStatus;
    assign `MYZPATH.i_phy_6_pipe_RxStandbyStatus        =       i_phy_6_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_6_pipe_PhyStatus              =       i_phy_6_pipe_PhyStatus;
    assign `MYZPATH.i_phy_6_pipe_PclkChangeOk           =       i_phy_6_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_6_pipe_P2M_MessageBus         =       i_phy_6_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_7_pipe_RxClk                  =       i_phy_7_pipe_RxClk;
    assign `MYZPATH.i_phy_7_pipe_RxValid                =       i_phy_7_pipe_RxValid;
    assign `MYZPATH.i_phy_7_pipe_RxData                 =       i_phy_7_pipe_RxData;
    assign `MYZPATH.i_phy_7_pipe_RxElecIdle             =       i_phy_7_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_7_pipe_RxStatus               =       i_phy_7_pipe_RxStatus;
    assign `MYZPATH.i_phy_7_pipe_RxStandbyStatus        =       i_phy_7_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_7_pipe_PhyStatus              =       i_phy_7_pipe_PhyStatus;
    assign `MYZPATH.i_phy_7_pipe_PclkChangeOk           =       i_phy_7_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_7_pipe_P2M_MessageBus         =       i_phy_7_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_8_pipe_RxClk                  =       i_phy_8_pipe_RxClk;
    assign `MYZPATH.i_phy_8_pipe_RxValid                =       i_phy_8_pipe_RxValid;
    assign `MYZPATH.i_phy_8_pipe_RxData                 =       i_phy_8_pipe_RxData;
    assign `MYZPATH.i_phy_8_pipe_RxElecIdle             =       i_phy_8_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_8_pipe_RxStatus               =       i_phy_8_pipe_RxStatus;
    assign `MYZPATH.i_phy_8_pipe_RxStandbyStatus        =       i_phy_8_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_8_pipe_PhyStatus              =       i_phy_8_pipe_PhyStatus;
    assign `MYZPATH.i_phy_8_pipe_PclkChangeOk           =       i_phy_8_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_8_pipe_P2M_MessageBus         =       i_phy_8_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_9_pipe_RxClk                  =       i_phy_9_pipe_RxClk;
    assign `MYZPATH.i_phy_9_pipe_RxValid                =       i_phy_9_pipe_RxValid;
    assign `MYZPATH.i_phy_9_pipe_RxData                 =       i_phy_9_pipe_RxData;
    assign `MYZPATH.i_phy_9_pipe_RxElecIdle             =       i_phy_9_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_9_pipe_RxStatus               =       i_phy_9_pipe_RxStatus;
    assign `MYZPATH.i_phy_9_pipe_RxStandbyStatus        =       i_phy_9_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_9_pipe_PhyStatus              =       i_phy_9_pipe_PhyStatus;
    assign `MYZPATH.i_phy_9_pipe_PclkChangeOk           =       i_phy_9_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_9_pipe_P2M_MessageBus         =       i_phy_9_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_10_pipe_RxClk                 =       i_phy_10_pipe_RxClk;
    assign `MYZPATH.i_phy_10_pipe_RxValid               =       i_phy_10_pipe_RxValid;
    assign `MYZPATH.i_phy_10_pipe_RxData                =       i_phy_10_pipe_RxData;
    assign `MYZPATH.i_phy_10_pipe_RxElecIdle            =       i_phy_10_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_10_pipe_RxStatus              =       i_phy_10_pipe_RxStatus;
    assign `MYZPATH.i_phy_10_pipe_RxStandbyStatus       =       i_phy_10_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_10_pipe_PhyStatus             =       i_phy_10_pipe_PhyStatus;
    assign `MYZPATH.i_phy_10_pipe_PclkChangeOk          =       i_phy_10_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_10_pipe_P2M_MessageBus        =       i_phy_10_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_11_pipe_RxClk                 =       i_phy_11_pipe_RxClk;
    assign `MYZPATH.i_phy_11_pipe_RxValid               =       i_phy_11_pipe_RxValid;
    assign `MYZPATH.i_phy_11_pipe_RxData                =       i_phy_11_pipe_RxData;
    assign `MYZPATH.i_phy_11_pipe_RxElecIdle            =       i_phy_11_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_11_pipe_RxStatus              =       i_phy_11_pipe_RxStatus;
    assign `MYZPATH.i_phy_11_pipe_RxStandbyStatus       =       i_phy_11_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_11_pipe_PhyStatus             =       i_phy_11_pipe_PhyStatus;
    assign `MYZPATH.i_phy_11_pipe_PclkChangeOk          =       i_phy_11_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_11_pipe_P2M_MessageBus        =       i_phy_11_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_12_pipe_RxClk                 =       i_phy_12_pipe_RxClk;
    assign `MYZPATH.i_phy_12_pipe_RxValid               =       i_phy_12_pipe_RxValid;
    assign `MYZPATH.i_phy_12_pipe_RxData                =       i_phy_12_pipe_RxData;
    assign `MYZPATH.i_phy_12_pipe_RxElecIdle            =       i_phy_12_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_12_pipe_RxStatus              =       i_phy_12_pipe_RxStatus;
    assign `MYZPATH.i_phy_12_pipe_RxStandbyStatus       =       i_phy_12_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_12_pipe_PhyStatus             =       i_phy_12_pipe_PhyStatus;
    assign `MYZPATH.i_phy_12_pipe_PclkChangeOk          =       i_phy_12_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_12_pipe_P2M_MessageBus        =       i_phy_12_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_13_pipe_RxClk                 =       i_phy_13_pipe_RxClk;
    assign `MYZPATH.i_phy_13_pipe_RxValid               =       i_phy_13_pipe_RxValid;
    assign `MYZPATH.i_phy_13_pipe_RxData                =       i_phy_13_pipe_RxData;
    assign `MYZPATH.i_phy_13_pipe_RxElecIdle            =       i_phy_13_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_13_pipe_RxStatus              =       i_phy_13_pipe_RxStatus;
    assign `MYZPATH.i_phy_13_pipe_RxStandbyStatus       =       i_phy_13_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_13_pipe_PhyStatus             =       i_phy_13_pipe_PhyStatus;
    assign `MYZPATH.i_phy_13_pipe_PclkChangeOk          =       i_phy_13_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_13_pipe_P2M_MessageBus        =       i_phy_13_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_14_pipe_RxClk                 =       i_phy_14_pipe_RxClk;
    assign `MYZPATH.i_phy_14_pipe_RxValid               =       i_phy_14_pipe_RxValid;
    assign `MYZPATH.i_phy_14_pipe_RxData                =       i_phy_14_pipe_RxData;
    assign `MYZPATH.i_phy_14_pipe_RxElecIdle            =       i_phy_14_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_14_pipe_RxStatus              =       i_phy_14_pipe_RxStatus;
    assign `MYZPATH.i_phy_14_pipe_RxStandbyStatus       =       i_phy_14_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_14_pipe_PhyStatus             =       i_phy_14_pipe_PhyStatus;
    assign `MYZPATH.i_phy_14_pipe_PclkChangeOk          =       i_phy_14_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_14_pipe_P2M_MessageBus        =       i_phy_14_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_15_pipe_RxClk                 =       i_phy_15_pipe_RxClk;
    assign `MYZPATH.i_phy_15_pipe_RxValid               =       i_phy_15_pipe_RxValid;
    assign `MYZPATH.i_phy_15_pipe_RxData                =       i_phy_15_pipe_RxData;
    assign `MYZPATH.i_phy_15_pipe_RxElecIdle            =       i_phy_15_pipe_RxElecIdle;
    assign `MYZPATH.i_phy_15_pipe_RxStatus              =       i_phy_15_pipe_RxStatus;
    assign `MYZPATH.i_phy_15_pipe_RxStandbyStatus       =       i_phy_15_pipe_RxStandbyStatus;
    assign `MYZPATH.i_phy_15_pipe_PhyStatus             =       i_phy_15_pipe_PhyStatus;
    assign `MYZPATH.i_phy_15_pipe_PclkChangeOk          =       i_phy_15_pipe_PclkChangeOk;
    assign `MYZPATH.i_phy_15_pipe_P2M_MessageBus        =       i_phy_15_pipe_P2M_MessageBus;
    assign `MYZPATH.i_phy_0_pipe_RxBitSlip_Ack          =       i_phy_0_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_1_pipe_RxBitSlip_Ack          =       i_phy_1_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_2_pipe_RxBitSlip_Ack          =       i_phy_2_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_3_pipe_RxBitSlip_Ack          =       i_phy_3_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_4_pipe_RxBitSlip_Ack          =       i_phy_4_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_5_pipe_RxBitSlip_Ack          =       i_phy_5_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_6_pipe_RxBitSlip_Ack          =       i_phy_6_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_7_pipe_RxBitSlip_Ack          =       i_phy_7_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_8_pipe_RxBitSlip_Ack          =       i_phy_8_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_9_pipe_RxBitSlip_Ack          =       i_phy_9_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_10_pipe_RxBitSlip_Ack         =       i_phy_10_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_11_pipe_RxBitSlip_Ack         =       i_phy_11_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_12_pipe_RxBitSlip_Ack         =       i_phy_12_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_13_pipe_RxBitSlip_Ack         =       i_phy_13_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_14_pipe_RxBitSlip_Ack         =       i_phy_14_pipe_RxBitSlip_Ack;
    assign `MYZPATH.i_phy_15_pipe_RxBitSlip_Ack         =       i_phy_15_pipe_RxBitSlip_Ack;
    `endif
    //-------------------------------------------------CXL Sim Time Reduction Assignment---------------------------------------------//

    //------------------------------------CXL Sim Time Reduction end----------------------------------------------------------------//

   // CXL Credit Signals
   assign cxl_cache_d2h_data0_crdrtn_o                = o_D2H_Data0_CrdRtn;
   assign cxl_cache_d2h_req_crdrtn_o                  = o_D2H_Req_CrdRtn;
   assign cxl_cache_d2h_rsp_crdrtn_o                  = o_D2H_Rsp_CrdRtn;

   assign  cxl_mem_s2m_drs0_crdrtn_o                  = o_S2M_DRS0_CrdRtn;
   assign  cxl_mem_s2m_drs1_crdrtn_o                  = o_S2M_DRS1_CrdRtn;
   assign  cxl_mem_s2m_ndr_crdrtn_o                   = o_S2M_NDR_CrdRtn;
   assign  cxl_cache_d2h_pushwr_crdrtn_o              = o_D2HPushWrCrdRtn;

   assign i_H2D_Data0_CrdRtn                          = cxl_cache_h2d_data0_crdrtn_i;
   assign i_H2D_Data1_CrdRtn                          = cxl_cache_h2d_data1_crdrtn_i;
   assign i_H2D_Req_CrdRtn                            = cxl_cache_h2d_req_crdrtn_i;
   assign i_H2D_Rsp_CrdRtn                            = cxl_cache_h2d_rsp_crdrtn_i;

   assign i_M2S_Req_CrdRtn                            = cxl_mem_m2s_req_crdrtn_i;
   assign i_M2S_RwD0_CrdRtn                           = cxl_mem_m2s_rwd0_crdrtn_i;
   assign i_M2S_RwD1_CrdRtn                           = cxl_mem_m2s_rwd1_crdrtn_i;

   assign  i_H2D_Rsp_CrdRtn_fr0                       = cxl_cache_h2d_rsp_crdrtn_fr0_i;
   assign  i_H2D_Rsp_CrdRtn_fr1                       = cxl_cache_h2d_rsp_crdrtn_fr1_i;
   assign  i_H2D_Req_CrdRtn_fr0                       = cxl_cache_h2d_req_crdrtn_fr0_i;
   assign  i_H2D_Req_CrdRtn_fr1                       = cxl_cache_h2d_req_crdrtn_fr1_i;
   assign  i_H2D_Data0_CrdRtn_fr0                     = cxl_cache_h2d_data_crdrtn_fr0_i;
   assign  i_H2D_Data0_CrdRtn_fr1                     = cxl_cache_h2d_data_crdrtn_fr1_i;
   assign   i_M2S_RwD0_CrdRtn_fr0                     = cxl_mem_m2s_rwd_crdrtn_fr0_i;
   assign  i_M2S_RwD0_CrdRtn_fr1                      = cxl_mem_m2s_rwd_crdrtn_fr1_i;
   assign  i_M2S_Req_CrdRtn_fr0                       = cxl_mem_m2s_req_crdrtn_fr0_i;
   assign  i_M2S_Req_CrdRtn_fr1                       = cxl_mem_m2s_req_crdrtn_fr1_i;


   //  //interfaces_cxl_mem_rx
   assign frame0_cxl_mem_port_id_o                      = cxl_cache_mem_rx_frame0.cxl_mem.prot_id;
   assign frame0_cxl_mem_m2s_rwd0_valid_o               = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_Valid;
   assign frame0_cxl_mem_m2s_rwd0_poison_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_Poison;
   assign frame0_cxl_mem_m2s_rwd0_beparity_o            = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_BEParity;
   assign frame0_cxl_mem_m2s_rwd0_dataparity_o          = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_DataParity;
   assign frame0_cxl_mem_m2s_rwd0_memopcode_o           = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_MemOpcode;
   assign frame0_cxl_mem_m2s_rwd0_metafield_o           = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_MetaField;
   assign frame0_cxl_mem_m2s_rwd0_metavalue_o           = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_MetaValue;
   assign frame0_cxl_mem_m2s_rwd0_snptype_o             = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_SnpType;
   assign frame0_cxl_mem_m2s_rwd0_tag_o                 = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_Tag;
   assign frame0_cxl_mem_m2s_rwd0_tc_o                  = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_TC;
   assign frame0_cxl_mem_m2s_req1_valid_o               = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_Valid;
   assign frame0_cxl_mem_m2s_req1_memopcode_o           = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_MemOpcode;
   assign frame0_cxl_mem_m2s_req1_metafield_o           = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_MetaField;
   assign frame0_cxl_mem_m2s_req1_metavalue_o           = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_MetaValue;
   assign frame0_cxl_mem_m2s_req1_snptype_o             = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_SnpType;
   assign frame0_cxl_mem_m2s_req1_tag_o                 = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_Tag;
   assign frame0_cxl_mem_m2s_req1_tc_o                  = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_TC;
   assign frame0_cxl_mem_m2s_req1_rsvd_h_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_Rsvd_H;
   assign frame0_cxl_mem_m2s_req1_address_o             = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_Address;
   assign frame0_cxl_mem_m2s_req1_rsvd_l_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_Rsvd_L;
   assign frame0_cxl_mem_m2s_req1_parity_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req1_Parity;
   assign frame0_cxl_mem_not_mapped_2_o                 = cxl_cache_mem_rx_frame0.cxl_mem.NOT_MAPPED_2;
   assign frame0_cxl_mem_m2s_req0_valid_o               = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_Valid;
   assign frame0_cxl_mem_m2s_req0_memopcode_o           = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_MemOpcode;
   assign frame0_cxl_mem_m2s_req0_metafield_o           = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_MetaField;
   assign frame0_cxl_mem_m2s_req0_metavalue_o           = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_MetaValue;
   assign frame0_cxl_mem_m2s_req0_snptype_o             = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_SnpType;
   assign frame0_cxl_mem_m2s_req0_tag_o                 = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_Tag;
   assign frame0_cxl_mem_m2s_req0_tc_o                  = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_TC;
   assign frame0_cxl_mem_m2s_req0_rsvd_h_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_Rsvd_H;
   assign frame0_cxl_mem_m2s_req0_address_o             = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_Address;
   assign frame0_cxl_mem_m2s_req0_rsvd_l_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_Rsvd_L;
   assign frame0_cxl_mem_m2s_req0_parity_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_Req0_Parity;
   assign frame0_cxl_mem_m2s_rwd0_rsvd_h_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_Rsvd_H;
   assign frame0_cxl_mem_m2s_rwd0_address_o             = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_Address;
   assign frame0_cxl_mem_m2s_rwd0_rsvd_l_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_Rsvd_L;
   assign frame0_cxl_mem_not_mapped_1_o                 = cxl_cache_mem_rx_frame0.cxl_mem.NOT_MAPPED_1;
   assign frame0_cxl_mem_m2s_datahdr1_o                 = cxl_cache_mem_rx_frame0.cxl_mem.M2SDataHdr1;
   assign frame0_cxl_mem_m2s_rwd0_byteen_h_o            = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_ByteEn_H;
   assign frame0_cxl_mem_m2s_rwd0_data_h_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_Data_H;
   assign frame0_cxl_mem_not_mapped_0_o                 = cxl_cache_mem_rx_frame0.cxl_mem.NOT_MAPPED_0;
   assign frame0_cxl_mem_m2s_rwd0_hdrparity_o           = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_HdrParity;
   assign frame0_cxl_mem_m2s_rwd0_byteen_l_o            = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_ByteEn_L;
   assign frame0_cxl_mem_m2s_rwd0_data_l_o              = cxl_cache_mem_rx_frame0.cxl_mem.M2S_RwD0_Data_L;
   assign frame1_cxl_mem_port_id_o                      = cxl_cache_mem_rx_frame1.cxl_mem.prot_id;
   assign frame1_cxl_mem_m2s_rwd0_valid_o               = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_Valid;
   assign frame1_cxl_mem_m2s_rwd0_poison_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_Poison;
   assign frame1_cxl_mem_m2s_rwd0_beparity_o            = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_BEParity;
   assign frame1_cxl_mem_m2s_rwd0_dataparity_o          = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_DataParity;
   assign frame1_cxl_mem_m2s_rwd0_memopcode_o           = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_MemOpcode;
   assign frame1_cxl_mem_m2s_rwd0_metafield_o           = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_MetaField;
   assign frame1_cxl_mem_m2s_rwd0_metavalue_o           = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_MetaValue;
   assign frame1_cxl_mem_m2s_rwd0_snptype_o             = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_SnpType;
   assign frame1_cxl_mem_m2s_rwd0_tag_o                 = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_Tag;
   assign frame1_cxl_mem_m2s_rwd0_tc_o                  = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_TC;
   assign frame1_cxl_mem_m2s_req1_valid_o               = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_Valid;
   assign frame1_cxl_mem_m2s_req1_memopcode_o           = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_MemOpcode;
   assign frame1_cxl_mem_m2s_req1_metafield_o           = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_MetaField;
   assign frame1_cxl_mem_m2s_req1_metavalue_o           = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_MetaValue;
   assign frame1_cxl_mem_m2s_req1_snptype_o             = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_SnpType;
   assign frame1_cxl_mem_m2s_req1_tag_o                 = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_Tag;
   assign frame1_cxl_mem_m2s_req1_tc_o                  = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_TC;
   assign frame1_cxl_mem_m2s_req1_rsvd_h_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_Rsvd_H;
   assign frame1_cxl_mem_m2s_req1_address_o             = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_Address;
   assign frame1_cxl_mem_m2s_req1_rsvd_l_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_Rsvd_L;
   assign frame1_cxl_mem_m2s_req1_parity_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req1_Parity;
   assign frame1_cxl_mem_not_mapped_2_o                 = cxl_cache_mem_rx_frame1.cxl_mem.NOT_MAPPED_2;
   assign frame1_cxl_mem_m2s_req0_valid_o               = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_Valid;
   assign frame1_cxl_mem_m2s_req0_memopcode_o           = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_MemOpcode;
   assign frame1_cxl_mem_m2s_req0_metafield_o           = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_MetaField;
   assign frame1_cxl_mem_m2s_req0_metavalue_o           = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_MetaValue;
   assign frame1_cxl_mem_m2s_req0_snptype_o             = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_SnpType;
   assign frame1_cxl_mem_m2s_req0_tag_o                 = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_Tag;
   assign frame1_cxl_mem_m2s_req0_tc_o                  = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_TC;
   assign frame1_cxl_mem_m2s_req0_rsvd_h_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_Rsvd_H;
   assign frame1_cxl_mem_m2s_req0_address_o             = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_Address;
   assign frame1_cxl_mem_m2s_req0_rsvd_l_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_Rsvd_L;
   assign frame1_cxl_mem_m2s_req0_parity_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_Req0_Parity;
   assign frame1_cxl_mem_m2s_rwd0_rsvd_h_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_Rsvd_H;
   assign frame1_cxl_mem_m2s_rwd0_address_o             = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_Address;
   assign frame1_cxl_mem_m2s_rwd0_rsvd_l_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_Rsvd_L;
   assign frame1_cxl_mem_not_mapped_1_o                 = cxl_cache_mem_rx_frame1.cxl_mem.NOT_MAPPED_1;
   assign frame1_cxl_mem_m2s_datahdr1_o                  = cxl_cache_mem_rx_frame1.cxl_mem.M2SDataHdr1;
   assign frame1_cxl_mem_m2s_rwd0_byteen_h_o            = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_ByteEn_H;
   assign frame1_cxl_mem_m2s_rwd0_data_h_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_Data_H;
   assign frame1_cxl_mem_not_mapped_0_o                 = cxl_cache_mem_rx_frame1.cxl_mem.NOT_MAPPED_0;
   assign frame1_cxl_mem_m2s_rwd0_hdrparity_o           = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_HdrParity;
   assign frame1_cxl_mem_m2s_rwd0_byteen_l_o            = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_ByteEn_L;
   assign frame1_cxl_mem_m2s_rwd0_data_l_o              = cxl_cache_mem_rx_frame1.cxl_mem.M2S_RwD0_Data_L;
   //interfaces_cxl_cache_rx
   assign frame0_cxl_cache_port_id_o                    = cxl_cache_mem_rx_frame0.cxl_cache.prot_id;
   assign frame0_cxl_cache_not_mapped_2_o               = cxl_cache_mem_rx_frame0.cxl_cache.NOT_MAPPED_2;
   assign frame0_cxl_cache_h2d_rsp3_valid_o             = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp3_Valid;
   assign frame0_cxl_cache_h2d_rsp3_rsvd_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp3_Rsvd;
   assign frame0_cxl_cache_h2d_rsp3_parity_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp3_Parity;
   assign frame0_cxl_cache_h2d_rsp3_pre_o               = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp3_PRE;
   assign frame0_cxl_cache_h2d_rsp3_opcode_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp3_Opcode;
   assign frame0_cxl_cache_h2d_rsp3_cqid_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp3_CqID;
   assign frame0_cxl_cache_h2d_rsp3_data_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp3_Data;
   assign frame0_cxl_cache_not_mapped_1_o               = cxl_cache_mem_rx_frame0.cxl_cache.NOT_MAPPED_1;
   assign frame0_cxl_cache_h2d_data1_cqid_o             = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data1_CqID;
   assign frame0_cxl_cache_h2d_req1_valid_o             = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req1_Valid;
   assign frame0_cxl_cache_h2d_req1_rsvd_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req1_Rsvd;
   assign frame0_cxl_cache_h2d_req1_opcode_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req1_Opcode;
   assign frame0_cxl_cache_h2d_req1_parity_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req1_Parity;
   assign frame0_cxl_cache_h2d_req1_uqid_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req1_UqID;
   assign frame0_cxl_cache_h2d_req1_address_o           = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req1_Address;
   assign frame0_cxl_cache_h2d_rsp2_valid_o             = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp2_Valid;
   assign frame0_cxl_cache_h2d_rsp2_rsvd_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp2_Rsvd;
   assign frame0_cxl_cache_h2d_rsp2_parity_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp2_Parity;
   assign frame0_cxl_cache_h2d_rsp2_pre_o               = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp2_PRE;
   assign frame0_cxl_cache_h2d_rsp2_opcode_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp2_Opcode;
   assign frame0_cxl_cache_h2d_rsp2_cqid_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp2_CqID;
   assign frame0_cxl_cache_h2d_rsp2_data_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp2_Data;
   assign frame0_cxl_cache_h2d_req0_valid_o             = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req0_Valid;
   assign frame0_cxl_cache_h2d_req0_rsvd_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req0_Rsvd;
   assign frame0_cxl_cache_h2d_req0_opcode_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req0_Opcode;
   assign frame0_cxl_cache_h2d_req0_parity_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req0_Parity;
   assign frame0_cxl_cache_h2d_req0_uqid_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req0_UqID;
   assign frame0_cxl_cache_h2d_req0_address_o           = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Req0_Address;
   assign frame0_cxl_cache_h2d_datahdr1_parity_o        = cxl_cache_mem_rx_frame0.cxl_cache.H2D_DataHdr1_Parity;
   assign frame0_cxl_cache_not_mapped_0_o               = cxl_cache_mem_rx_frame0.cxl_cache.NOT_MAPPED_0;
   assign frame0_cxl_cache_h2d_rsp1_valid_o             = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp1_Valid;
   assign frame0_cxl_cache_h2d_rsp1_rsvd_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp1_Rsvd;
   assign frame0_cxl_cache_h2d_rsp1_parity_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp1_Parity;
   assign frame0_cxl_cache_h2d_rsp1_pre_o               = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp1_PRE;
   assign frame0_cxl_cache_h2d_rsp1_opcode_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp1_Opcode;
   assign frame0_cxl_cache_h2d_rsp1_cqid_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp1_CqID;
   assign frame0_cxl_cache_h2d_rsp1_data_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp1_Data;
   assign frame0_cxl_cache_h2d_data1_rsvd_o             = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data1_Rsvd;
   assign frame0_cxl_cache_h2d_rsp0_valid_o             = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp0_Valid;
   assign frame0_cxl_cache_h2d_rsp0_rsvd_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp0_Rsvd;
   assign frame0_cxl_cache_h2d_rsp0_parity_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp0_Parity;
   assign frame0_cxl_cache_h2d_rsp0_pre_o               = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp0_PRE;
   assign frame0_cxl_cache_h2d_rsp0_opcode_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp0_Opcode;
   assign frame0_cxl_cache_h2d_rsp0_cqid_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp0_CqID;
   assign frame0_cxl_cache_h2d_rsp0_data_o              = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Rsp0_Data;
   assign frame0_cxl_cache_h2d_data0_data_h_o           = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data0_Data_H;
   assign frame0_cxl_cache_h2d_data1_valid_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data1_Valid;
   assign frame0_cxl_cache_h2d_data1_chunkvalid_o       = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data1_ChunkValid;
   assign frame0_cxl_cache_h2d_data0_valid_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data0_Valid;
   assign frame0_cxl_cache_h2d_data0_chunkvalid_o       = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data0_ChunkValid;
   assign frame0_cxl_cache_h2d_data0_poison_o           = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data0_Poison;
   assign frame0_cxl_cache_h2d_data0_goerr_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data0_GoErr;
   assign frame0_cxl_cache_h2d_datahdr0_parity_o        = cxl_cache_mem_rx_frame0.cxl_cache.H2D_DataHdr0_Parity;
   assign frame0_cxl_cache_h2d_data0_dataparity_o       = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data0_DataParity;
   assign frame0_cxl_cache_h2d_data0_rsvd_o             = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data0_Rsvd;
   assign frame0_cxl_cache_h2d_data1_poison_o           = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data1_Poison;
   assign frame0_cxl_cache_h2d_data1_goerr_o            = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data1_GoErr;
   assign frame0_cxl_cache_h2d_data0_cqid_o             = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data0_CqID;
   assign frame0_cxl_cache_h2d_data0_data_l_o           = cxl_cache_mem_rx_frame0.cxl_cache.H2D_Data0_Data_L;
   assign frame1_cxl_cache_port_id_o                    = cxl_cache_mem_rx_frame1.cxl_cache.prot_id;
   assign frame1_cxl_cache_not_mapped_2_o               = cxl_cache_mem_rx_frame1.cxl_cache.NOT_MAPPED_2;
   assign frame1_cxl_cache_h2d_rsp3_valid_o             = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp3_Valid;
   assign frame1_cxl_cache_h2d_rsp3_rsvd_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp3_Rsvd;
   assign frame1_cxl_cache_h2d_rsp3_parity_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp3_Parity;
   assign frame1_cxl_cache_h2d_rsp3_pre_o               = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp3_PRE;
   assign frame1_cxl_cache_h2d_rsp3_opcode_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp3_Opcode;
   assign frame1_cxl_cache_h2d_rsp3_cqid_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp3_CqID;
   assign frame1_cxl_cache_h2d_rsp3_data_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp3_Data;
   assign frame1_cxl_cache_not_mapped_1_o               = cxl_cache_mem_rx_frame1.cxl_cache.NOT_MAPPED_1;
   assign frame1_cxl_cache_h2d_data1_cqid_o             = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data1_CqID;
   assign frame1_cxl_cache_h2d_req1_valid_o             = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req1_Valid;
   assign frame1_cxl_cache_h2d_req1_rsvd_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req1_Rsvd;
   assign frame1_cxl_cache_h2d_req1_opcode_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req1_Opcode;
   assign frame1_cxl_cache_h2d_req1_parity_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req1_Parity;
   assign frame1_cxl_cache_h2d_req1_uqid_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req1_UqID;
   assign frame1_cxl_cache_h2d_req1_address_o           = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req1_Address;
   assign frame1_cxl_cache_h2d_rsp2_valid_o             = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp2_Valid;
   assign frame1_cxl_cache_h2d_rsp2_rsvd_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp2_Rsvd;
   assign frame1_cxl_cache_h2d_rsp2_parity_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp2_Parity;
   assign frame1_cxl_cache_h2d_rsp2_pre_o               = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp2_PRE;
   assign frame1_cxl_cache_h2d_rsp2_opcode_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp2_Opcode;
   assign frame1_cxl_cache_h2d_rsp2_cqid_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp2_CqID;
   assign frame1_cxl_cache_h2d_rsp2_data_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp2_Data;
   assign frame1_cxl_cache_h2d_req0_valid_o             = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req0_Valid;
   assign frame1_cxl_cache_h2d_req0_rsvd_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req0_Rsvd;
   assign frame1_cxl_cache_h2d_req0_opcode_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req0_Opcode;
   assign frame1_cxl_cache_h2d_req0_parity_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req0_Parity;
   assign frame1_cxl_cache_h2d_req0_uqid_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req0_UqID;
   assign frame1_cxl_cache_h2d_req0_address_o           = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Req0_Address;
   assign frame1_cxl_cache_h2d_datahdr1_parity_o        = cxl_cache_mem_rx_frame1.cxl_cache.H2D_DataHdr1_Parity;
   assign frame1_cxl_cache_not_mapped_0_o               = cxl_cache_mem_rx_frame1.cxl_cache.NOT_MAPPED_0;
   assign frame1_cxl_cache_h2d_rsp1_valid_o             = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp1_Valid;
   assign frame1_cxl_cache_h2d_rsp1_rsvd_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp1_Rsvd;
   assign frame1_cxl_cache_h2d_rsp1_parity_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp1_Parity;
   assign frame1_cxl_cache_h2d_rsp1_pre_o               = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp1_PRE;
   assign frame1_cxl_cache_h2d_rsp1_opcode_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp1_Opcode;
   assign frame1_cxl_cache_h2d_rsp1_cqid_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp1_CqID;
   assign frame1_cxl_cache_h2d_rsp1_data_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp1_Data;
   assign frame1_cxl_cache_h2d_data1_rsvd_o             = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data1_Rsvd;
   assign frame1_cxl_cache_h2d_rsp0_valid_o             = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp0_Valid;
   assign frame1_cxl_cache_h2d_rsp0_rsvd_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp0_Rsvd;
   assign frame1_cxl_cache_h2d_rsp0_parity_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp0_Parity;
   assign frame1_cxl_cache_h2d_rsp0_pre_o               = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp0_PRE;
   assign frame1_cxl_cache_h2d_rsp0_opcode_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp0_Opcode;
   assign frame1_cxl_cache_h2d_rsp0_cqid_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp0_CqID;
   assign frame1_cxl_cache_h2d_rsp0_data_o              = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Rsp0_Data;
   assign frame1_cxl_cache_h2d_data0_data_h_o           = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data0_Data_H;
   assign frame1_cxl_cache_h2d_data1_valid_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data1_Valid;
   assign frame1_cxl_cache_h2d_data1_chunkvalid_o       = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data1_ChunkValid;
   assign frame1_cxl_cache_h2d_data0_valid_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data0_Valid;
   assign frame1_cxl_cache_h2d_data0_chunkvalid_o       = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data0_ChunkValid;
   assign frame1_cxl_cache_h2d_data0_poison_o           = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data0_Poison;
   assign frame1_cxl_cache_h2d_data0_goerr_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data0_GoErr;
   assign frame1_cxl_cache_h2d_datahdr0_parity_o        = cxl_cache_mem_rx_frame1.cxl_cache.H2D_DataHdr0_Parity;
   assign frame1_cxl_cache_h2d_data0_dataparity_o       = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data0_DataParity;
   assign frame1_cxl_cache_h2d_data0_rsvd_o             = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data0_Rsvd;
   assign frame1_cxl_cache_h2d_data1_poison_o           = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data1_Poison;
   assign frame1_cxl_cache_h2d_data1_goerr_o            = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data1_GoErr;
   assign frame1_cxl_cache_h2d_data0_cqid_o             = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data0_CqID;
   assign frame1_cxl_cache_h2d_data0_data_l_o           = cxl_cache_mem_rx_frame1.cxl_cache.H2D_Data0_Data_L;

   // CXL.mem and CXL.Cache TX
   rnr_cxl_pkg::cxl_mem_s2m_tx_intf          cxl_mem_s2m_tx_frame0;
   logic                        cxl_mem_s2m_tx_frame0_ready;
   rnr_cxl_pkg::cxl_mem_s2m_tx_intf          cxl_mem_s2m_tx_frame1;
   logic                        cxl_mem_s2m_tx_frame1_ready;
   //interfaces_cxl_mem_s2m_tx
////  if  (hssi_ctr_silicon_rev == "10nm6arnrb" || hssi_ctr_silicon_rev == "10nm8arnrb") begin
  assign cxl_mem_s2m_tx_frame0.S2M_NDR1_DevLoad = frame0_cxl_mem_s2m_ndr1_devload_i; //B0 only
  assign cxl_mem_s2m_tx_frame0.S2M_NDR0_DevLoad = frame0_cxl_mem_s2m_ndr0_devload_i; //B0 only
  assign cxl_mem_s2m_tx_frame1.S2M_NDR1_DevLoad = frame1_cxl_mem_s2m_ndr1_devload_i; //B0 only
  assign cxl_mem_s2m_tx_frame1.S2M_NDR0_DevLoad = frame1_cxl_mem_s2m_ndr0_devload_i;
////  end
////  else begin
////   assign cxl_mem_s2m_tx_frame0.S2M_NDR1_DevLoad = 'h0; //B0 only
////   assign cxl_mem_s2m_tx_frame0.S2M_NDR0_DevLoad = 'h0; //B0 only
////   assign cxl_mem_s2m_tx_frame1.S2M_NDR1_DevLoad = 'h0; //B0 only
////   assign cxl_mem_s2m_tx_frame1.S2M_NDR0_DevLoad = 'h0;
////  end
   assign cxl_mem_s2m_tx_frame0.S2M_NDR1_Valid        =   frame0_cxl_mem_s2m_ndr1_valid_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR1_Opcode       =   frame0_cxl_mem_s2m_ndr1_opcode_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR1_MetaField    =   frame0_cxl_mem_s2m_ndr1_metafield_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR1_MetaValue    =   frame0_cxl_mem_s2m_ndr1_metavalue_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR1_Parity       =   frame0_cxl_mem_s2m_ndr1_parity_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR1_Rsvd         =   frame0_cxl_mem_s2m_ndr1_rsvd_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR1_Tag          =   frame0_cxl_mem_s2m_ndr1_tag_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR0_Valid        =   frame0_cxl_mem_s2m_ndr0_valid_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR0_Opcode       =   frame0_cxl_mem_s2m_ndr0_opcode_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR0_MetaField    =   frame0_cxl_mem_s2m_ndr0_metafield_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR0_MetaValue    =   frame0_cxl_mem_s2m_ndr0_metavalue_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR0_Parity       =   frame0_cxl_mem_s2m_ndr0_parity_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR0_Rsvd         =   frame0_cxl_mem_s2m_ndr0_rsvd_i;
   assign cxl_mem_s2m_tx_frame0.S2M_NDR0_Tag          =   frame0_cxl_mem_s2m_ndr0_tag_i;
   assign cxl_mem_s2m_tx_frame0.S2MDRSHdr1            =   frame0_cxl_mem_s2m_drs_hdr1_i;
   assign cxl_mem_s2m_tx_frame0.S2M_DRS0_Valid        =   frame0_cxl_mem_s2m_drs0_valid_i;
   assign cxl_mem_s2m_tx_frame0.S2M_DRS0_Poison       =   frame0_cxl_mem_s2m_drs0_poison_i;
   assign cxl_mem_s2m_tx_frame0.S2M_DRS0_Opcode       =   frame0_cxl_mem_s2m_drs0_opcode_i;
   assign cxl_mem_s2m_tx_frame0.S2M_DRS0_MetaField    =   frame0_cxl_mem_s2m_drs0_metafield_i;
   assign cxl_mem_s2m_tx_frame0.S2M_DRS0_MetaValue    =   frame0_cxl_mem_s2m_drs0_metavalue_i;
   assign cxl_mem_s2m_tx_frame0.S2M_DRS0_HdrParity    =   frame0_cxl_mem_s2m_drs0_hdrparity_i;
   assign cxl_mem_s2m_tx_frame0.S2M_DRS0_DataParity   =   frame0_cxl_mem_s2m_drs0_dataparity_i;
   assign cxl_mem_s2m_tx_frame0.S2M_DRS0_Tag          =   frame0_cxl_mem_s2m_drs0_tag_i;
   assign cxl_mem_s2m_tx_frame0.S2M_DRS0_Data         =   frame0_cxl_mem_s2m_drs0_data_i;
   assign cxl_mem_s2m_tx_frame0_valid                 =   frame0_cxl_mem_s2m_valid_i;
   assign frame0_cxl_mem_s2m_ready_o                  =   cxl_mem_s2m_tx_frame0_ready;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR1_Valid        =   frame1_cxl_mem_s2m_ndr1_valid_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR1_Opcode       =   frame1_cxl_mem_s2m_ndr1_opcode_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR1_MetaField    =   frame1_cxl_mem_s2m_ndr1_metafield_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR1_MetaValue    =   frame1_cxl_mem_s2m_ndr1_metavalue_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR1_Parity       =   frame1_cxl_mem_s2m_ndr1_parity_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR1_Rsvd         =   frame1_cxl_mem_s2m_ndr1_rsvd_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR1_Tag          =   frame1_cxl_mem_s2m_ndr1_tag_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR0_Valid        =   frame1_cxl_mem_s2m_ndr0_valid_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR0_Opcode       =   frame1_cxl_mem_s2m_ndr0_opcode_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR0_MetaField    =   frame1_cxl_mem_s2m_ndr0_metafield_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR0_MetaValue    =   frame1_cxl_mem_s2m_ndr0_metavalue_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR0_Parity       =   frame1_cxl_mem_s2m_ndr0_parity_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR0_Rsvd         =   frame1_cxl_mem_s2m_ndr0_rsvd_i;
   assign cxl_mem_s2m_tx_frame1.S2M_NDR0_Tag          =   frame1_cxl_mem_s2m_ndr0_tag_i;
   assign cxl_mem_s2m_tx_frame1.S2MDRSHdr1            =   frame1_cxl_mem_s2m_drs_hdr1_i;
   assign cxl_mem_s2m_tx_frame1.S2M_DRS0_Valid        =   frame1_cxl_mem_s2m_drs0_valid_i;
   assign cxl_mem_s2m_tx_frame1.S2M_DRS0_Poison       =   frame1_cxl_mem_s2m_drs0_poison_i;
   assign cxl_mem_s2m_tx_frame1.S2M_DRS0_Opcode       =   frame1_cxl_mem_s2m_drs0_opcode_i;
   assign cxl_mem_s2m_tx_frame1.S2M_DRS0_MetaField    =   frame1_cxl_mem_s2m_drs0_metafield_i;
   assign cxl_mem_s2m_tx_frame1.S2M_DRS0_MetaValue    =   frame1_cxl_mem_s2m_drs0_metavalue_i;
   assign cxl_mem_s2m_tx_frame1.S2M_DRS0_HdrParity    =   frame1_cxl_mem_s2m_drs0_hdrparity_i;
   assign cxl_mem_s2m_tx_frame1.S2M_DRS0_DataParity   =   frame1_cxl_mem_s2m_drs0_dataparity_i;
   assign cxl_mem_s2m_tx_frame1.S2M_DRS0_Tag          =   frame1_cxl_mem_s2m_drs0_tag_i;
   assign cxl_mem_s2m_tx_frame1.S2M_DRS0_Data         =   frame1_cxl_mem_s2m_drs0_data_i;
   assign cxl_mem_s2m_tx_frame1_valid                 =   frame1_cxl_mem_s2m_valid_i;
   assign frame1_cxl_mem_s2m_ready_o                  =   cxl_mem_s2m_tx_frame1_ready;

   if(REV_B0 == 1 || REV_C0 == 1) begin 
     assign cxl_mem_s2m_tx_frame0.S2M_DRS0_Rsvd         =   {frame0_cxl_mem_s2m_drs0_rsvd_field1_i,frame0_cxl_mem_s2m_drs0_devload_i,frame0_cxl_mem_s2m_drs0_rsvd_field0_i};
     assign cxl_mem_s2m_tx_frame1.S2M_DRS0_Rsvd         =   {frame1_cxl_mem_s2m_drs0_rsvd_field1_i,frame1_cxl_mem_s2m_drs0_devload_i,frame1_cxl_mem_s2m_drs0_rsvd_field0_i};
   end 
   else begin
     assign cxl_mem_s2m_tx_frame0.S2M_DRS0_Rsvd         =   frame0_cxl_mem_s2m_drs0_rsvd_i;
     assign cxl_mem_s2m_tx_frame1.S2M_DRS0_Rsvd         =   frame1_cxl_mem_s2m_drs0_rsvd_i;
   end 
   rnr_cxl_pkg::cxl_cache_d2h_req_tx_intf    cxl_d2h_req_frame0;
   logic [3:0]                  cxl_d2h_req_frame0_valid;
   logic [3:0]                  cxl_d2h_req_frame0_ready;
   rnr_cxl_pkg::cxl_cache_d2h_req_tx_intf    cxl_d2h_req_frame1;
   logic [3:0]                  cxl_d2h_req_frame1_valid;
   logic [3:0]                  cxl_d2h_req_frame1_ready;

   //interfaces_cxl_cache_d2h_req_tx
   assign cxl_d2h_req_frame0.D2H_Req3_Address         =   frame0_cxl_cache_d2h_req3_address_i;
   assign cxl_d2h_req_frame0.D2H_Req3_Parity          =   frame0_cxl_cache_d2h_req3_parity_i;
   assign cxl_d2h_req_frame0.D2H_Req3_CqID            =   frame0_cxl_cache_d2h_req3_cqid_i;
   assign cxl_d2h_req_frame0.D2H_Req3_Clos            =   frame0_cxl_cache_d2h_req3_clos_i;
   assign cxl_d2h_req_frame0.D2H_Req3_SecID           =   frame0_cxl_cache_d2h_req3_secid_i;
   assign cxl_d2h_req_frame0.D2H_Req3_NonTemporal     =   frame0_cxl_cache_d2h_req3_nontemporal_i;
   assign cxl_d2h_req_frame0.D2H_Req3_CacheNear       =   frame0_cxl_cache_d2h_req3_cachenear_i;
   assign cxl_d2h_req_frame0.D2H_Req3_PushWrite       =   frame0_cxl_cache_d2h_req3_pushwrite_i;
   assign cxl_d2h_req_frame0.D2H_Req3_StrmID          =   frame0_cxl_cache_d2h_req3_strmid_i;
   assign cxl_d2h_req_frame0.D2H_Req3_Rsvd            =   frame0_cxl_cache_d2h_req3_rsvd_i;
   assign cxl_d2h_req_frame0.D2H_Req3_Opcode          =   frame0_cxl_cache_d2h_req3_opcode_i;
   assign cxl_d2h_req_frame0.D2H_Req3_Valid           =   frame0_cxl_cache_d2h_req3_valid_i;
   assign cxl_d2h_req_frame0.D2H_Req2_Address         =   frame0_cxl_cache_d2h_req2_address_i;
   assign cxl_d2h_req_frame0.D2H_Req2_Parity          =   frame0_cxl_cache_d2h_req2_parity_i;
   assign cxl_d2h_req_frame0.D2H_Req2_CqID            =   frame0_cxl_cache_d2h_req2_cqid_i;
   assign cxl_d2h_req_frame0.D2H_Req2_Clos            =   frame0_cxl_cache_d2h_req2_clos_i;
   assign cxl_d2h_req_frame0.D2H_Req2_SecID           =   frame0_cxl_cache_d2h_req2_secid_i;
   assign cxl_d2h_req_frame0.D2H_Req2_NonTemporal     =   frame0_cxl_cache_d2h_req2_nontemporal_i;
   assign cxl_d2h_req_frame0.D2H_Req2_CacheNear       =   frame0_cxl_cache_d2h_req2_cachenear_i;
   assign cxl_d2h_req_frame0.D2H_Req2_PushWrite       =   frame0_cxl_cache_d2h_req2_pushwrite_i;
   assign cxl_d2h_req_frame0.D2H_Req2_StrmID          =   frame0_cxl_cache_d2h_req2_strmid_i;
   assign cxl_d2h_req_frame0.D2H_Req2_Rsvd            =   frame0_cxl_cache_d2h_req2_rsvd_i;
   assign cxl_d2h_req_frame0.D2H_Req2_Opcode          =   frame0_cxl_cache_d2h_req2_opcode_i;
   assign cxl_d2h_req_frame0.D2H_Req2_Valid           =   frame0_cxl_cache_d2h_req2_valid_i;
   assign cxl_d2h_req_frame0.D2H_Req1_Address         =   frame0_cxl_cache_d2h_req1_address_i;
   assign cxl_d2h_req_frame0.D2H_Req1_Parity          =   frame0_cxl_cache_d2h_req1_parity_i;
   assign cxl_d2h_req_frame0.D2H_Req1_CqID            =   frame0_cxl_cache_d2h_req1_cqid_i;
   assign cxl_d2h_req_frame0.D2H_Req1_Clos            =   frame0_cxl_cache_d2h_req1_clos_i;
   assign cxl_d2h_req_frame0.D2H_Req1_SecID           =   frame0_cxl_cache_d2h_req1_secid_i;
   assign cxl_d2h_req_frame0.D2H_Req1_NonTemporal     =   frame0_cxl_cache_d2h_req1_nontemporal_i;
   assign cxl_d2h_req_frame0.D2H_Req1_CacheNear       =   frame0_cxl_cache_d2h_req1_cachenear_i;
   assign cxl_d2h_req_frame0.D2H_Req1_PushWrite       =   frame0_cxl_cache_d2h_req1_pushwrite_i;
   assign cxl_d2h_req_frame0.D2H_Req1_StrmID          =   frame0_cxl_cache_d2h_req1_strmid_i;
   assign cxl_d2h_req_frame0.D2H_Req1_Rsvd            =   frame0_cxl_cache_d2h_req1_rsvd_i;
   assign cxl_d2h_req_frame0.D2H_Req1_Opcode          =   frame0_cxl_cache_d2h_req1_opcode_i;
   assign cxl_d2h_req_frame0.D2H_Req1_Valid           =   frame0_cxl_cache_d2h_req1_valid_i;
   assign cxl_d2h_req_frame0.D2H_Req0_Address         =   frame0_cxl_cache_d2h_req0_address_i;
   assign cxl_d2h_req_frame0.D2H_Req0_Parity          =   frame0_cxl_cache_d2h_req0_parity_i;
   assign cxl_d2h_req_frame0.D2H_Req0_CqID            =   frame0_cxl_cache_d2h_req0_cqid_i;
   assign cxl_d2h_req_frame0.D2H_Req0_Clos            =   frame0_cxl_cache_d2h_req0_clos_i;
   assign cxl_d2h_req_frame0.D2H_Req0_SecID           =   frame0_cxl_cache_d2h_req0_secid_i;
   assign cxl_d2h_req_frame0.D2H_Req0_NonTemporal     =   frame0_cxl_cache_d2h_req0_nontemporal_i;
   assign cxl_d2h_req_frame0.D2H_Req0_CacheNear       =   frame0_cxl_cache_d2h_req0_cachenear_i;
   assign cxl_d2h_req_frame0.D2H_Req0_PushWrite       =   frame0_cxl_cache_d2h_req0_pushwrite_i;
   assign cxl_d2h_req_frame0.D2H_Req0_StrmID          =   frame0_cxl_cache_d2h_req0_strmid_i;
   assign cxl_d2h_req_frame0.D2H_Req0_Rsvd            =   frame0_cxl_cache_d2h_req0_rsvd_i;
   assign cxl_d2h_req_frame0.D2H_Req0_Opcode          =   frame0_cxl_cache_d2h_req0_opcode_i;
   assign cxl_d2h_req_frame0.D2H_Req0_Valid           =   frame0_cxl_cache_d2h_req0_valid_i;
   if (opt_d2h_req23_en_hwtcl ==1 || opt_cache_formatb_en_hwtcl ==1)
    assign cxl_d2h_req_frame0_valid                   =   frame0_cxl_cache_d2h_req_valid_i;
   else
    assign cxl_d2h_req_frame0_valid                   =  {2'b0,frame0_cxl_cache_d2h_req_valid_i[1:0]};

   assign frame0_cxl_cache_d2h_req_ready_o                    =   cxl_d2h_req_frame0_ready;
   assign cxl_d2h_req_frame1.D2H_Req3_Address         =   frame1_cxl_cache_d2h_req3_address_i;
   assign cxl_d2h_req_frame1.D2H_Req3_Parity          =   frame1_cxl_cache_d2h_req3_parity_i;
   assign cxl_d2h_req_frame1.D2H_Req3_CqID            =   frame1_cxl_cache_d2h_req3_cqid_i;
   assign cxl_d2h_req_frame1.D2H_Req3_Clos            =   frame1_cxl_cache_d2h_req3_clos_i;
   assign cxl_d2h_req_frame1.D2H_Req3_SecID           =   frame1_cxl_cache_d2h_req3_secid_i;
   assign cxl_d2h_req_frame1.D2H_Req3_NonTemporal     =   frame1_cxl_cache_d2h_req3_nontemporal_i;
   assign cxl_d2h_req_frame1.D2H_Req3_CacheNear       =   frame1_cxl_cache_d2h_req3_cachenear_i;
   assign cxl_d2h_req_frame1.D2H_Req3_PushWrite       =   frame1_cxl_cache_d2h_req3_pushwrite_i;
   assign cxl_d2h_req_frame1.D2H_Req3_StrmID          =   frame1_cxl_cache_d2h_req3_strmid_i;
   assign cxl_d2h_req_frame1.D2H_Req3_Rsvd            =   frame1_cxl_cache_d2h_req3_rsvd_i;
   assign cxl_d2h_req_frame1.D2H_Req3_Opcode          =   frame1_cxl_cache_d2h_req3_opcode_i;
   assign cxl_d2h_req_frame1.D2H_Req3_Valid           =   frame1_cxl_cache_d2h_req3_valid_i;
   assign cxl_d2h_req_frame1.D2H_Req2_Address         =   frame1_cxl_cache_d2h_req2_address_i;
   assign cxl_d2h_req_frame1.D2H_Req2_Parity          =   frame1_cxl_cache_d2h_req2_parity_i;
   assign cxl_d2h_req_frame1.D2H_Req2_CqID            =   frame1_cxl_cache_d2h_req2_cqid_i;
   assign cxl_d2h_req_frame1.D2H_Req2_Clos            =   frame1_cxl_cache_d2h_req2_clos_i;
   assign cxl_d2h_req_frame1.D2H_Req2_SecID           =   frame1_cxl_cache_d2h_req2_secid_i;
   assign cxl_d2h_req_frame1.D2H_Req2_NonTemporal     =   frame1_cxl_cache_d2h_req2_nontemporal_i;
   assign cxl_d2h_req_frame1.D2H_Req2_CacheNear       =   frame1_cxl_cache_d2h_req2_cachenear_i;
   assign cxl_d2h_req_frame1.D2H_Req2_PushWrite       =   frame1_cxl_cache_d2h_req2_pushwrite_i;
   assign cxl_d2h_req_frame1.D2H_Req2_StrmID          =   frame1_cxl_cache_d2h_req2_strmid_i;
   assign cxl_d2h_req_frame1.D2H_Req2_Rsvd            =   frame1_cxl_cache_d2h_req2_rsvd_i;
   assign cxl_d2h_req_frame1.D2H_Req2_Opcode          =   frame1_cxl_cache_d2h_req2_opcode_i;
   assign cxl_d2h_req_frame1.D2H_Req2_Valid           =   frame1_cxl_cache_d2h_req2_valid_i;
   assign cxl_d2h_req_frame1.D2H_Req1_Address         =   frame1_cxl_cache_d2h_req1_address_i;
   assign cxl_d2h_req_frame1.D2H_Req1_Parity          =   frame1_cxl_cache_d2h_req1_parity_i;
   assign cxl_d2h_req_frame1.D2H_Req1_CqID            =   frame1_cxl_cache_d2h_req1_cqid_i;
   assign cxl_d2h_req_frame1.D2H_Req1_Clos            =   frame1_cxl_cache_d2h_req1_clos_i;
   assign cxl_d2h_req_frame1.D2H_Req1_SecID           =   frame1_cxl_cache_d2h_req1_secid_i;
   assign cxl_d2h_req_frame1.D2H_Req1_NonTemporal     =   frame1_cxl_cache_d2h_req1_nontemporal_i;
   assign cxl_d2h_req_frame1.D2H_Req1_CacheNear       =   frame1_cxl_cache_d2h_req1_cachenear_i;
   assign cxl_d2h_req_frame1.D2H_Req1_PushWrite       =   frame1_cxl_cache_d2h_req1_pushwrite_i;
   assign cxl_d2h_req_frame1.D2H_Req1_StrmID          =   frame1_cxl_cache_d2h_req1_strmid_i;
   assign cxl_d2h_req_frame1.D2H_Req1_Rsvd            =   frame1_cxl_cache_d2h_req1_rsvd_i;
   assign cxl_d2h_req_frame1.D2H_Req1_Opcode          =   frame1_cxl_cache_d2h_req1_opcode_i;
   assign cxl_d2h_req_frame1.D2H_Req1_Valid           =   frame1_cxl_cache_d2h_req1_valid_i;
   assign cxl_d2h_req_frame1.D2H_Req0_Address         =   frame1_cxl_cache_d2h_req0_address_i;
   assign cxl_d2h_req_frame1.D2H_Req0_Parity          =   frame1_cxl_cache_d2h_req0_parity_i;
   assign cxl_d2h_req_frame1.D2H_Req0_CqID            =   frame1_cxl_cache_d2h_req0_cqid_i;
   assign cxl_d2h_req_frame1.D2H_Req0_Clos            =   frame1_cxl_cache_d2h_req0_clos_i;
   assign cxl_d2h_req_frame1.D2H_Req0_SecID           =   frame1_cxl_cache_d2h_req0_secid_i;
   assign cxl_d2h_req_frame1.D2H_Req0_NonTemporal     =   frame1_cxl_cache_d2h_req0_nontemporal_i;
   assign cxl_d2h_req_frame1.D2H_Req0_CacheNear       =   frame1_cxl_cache_d2h_req0_cachenear_i;
   assign cxl_d2h_req_frame1.D2H_Req0_PushWrite       =   frame1_cxl_cache_d2h_req0_pushwrite_i;
   assign cxl_d2h_req_frame1.D2H_Req0_StrmID          =   frame1_cxl_cache_d2h_req0_strmid_i;
   assign cxl_d2h_req_frame1.D2H_Req0_Rsvd            =   frame1_cxl_cache_d2h_req0_rsvd_i;
   assign cxl_d2h_req_frame1.D2H_Req0_Opcode          =   frame1_cxl_cache_d2h_req0_opcode_i;
   assign cxl_d2h_req_frame1.D2H_Req0_Valid           =   frame1_cxl_cache_d2h_req0_valid_i;
  if (opt_d2h_req23_en_hwtcl ==1 || opt_cache_formatb_en_hwtcl ==1)
    assign cxl_d2h_req_frame1_valid                   =   frame1_cxl_cache_d2h_req_valid_i;
   else
    assign cxl_d2h_req_frame1_valid                   =   {2'b0,frame1_cxl_cache_d2h_req_valid_i[1:0]};

   assign frame1_cxl_cache_d2h_req_ready_o                    =   cxl_d2h_req_frame1_ready;

   rnr_cxl_pkg::cxl_cache_d2h_rsp_tx_intf     cxl_d2h_rsp_frame0;                 // 0 - 1;           1 ready
   wire [1:0]                    cxl_d2h_rsp_frame0_valid;
   wire [1:0]                    cxl_d2h_rsp_frame0_ready;
   rnr_cxl_pkg::cxl_cache_d2h_rsp_tx_intf     cxl_d2h_rsp_frame1;                 // 2 - 3;           1 ready
   wire [1:0]                    cxl_d2h_rsp_frame1_valid;
   wire [1:0]                    cxl_d2h_rsp_frame1_ready;

   //interfaces_cxl_cache_d2h_rsp_tx
   assign cxl_d2h_rsp_frame0.D2H_Rsp1_Valid           = frame0_cxl_cache_d2h_rsp1_valid_i;
   assign cxl_d2h_rsp_frame0.D2H_Rsp1_Opcode          = frame0_cxl_cache_d2h_rsp1_opcode_i;
   assign cxl_d2h_rsp_frame0.D2H_Rsp1_Parity          = frame0_cxl_cache_d2h_rsp1_parity_i;
   assign cxl_d2h_rsp_frame0.D2H_Rsp1_Rsvd            = frame0_cxl_cache_d2h_rsp1_rsvd_i;
   assign cxl_d2h_rsp_frame0.D2H_Rsp1_UqID            = frame0_cxl_cache_d2h_rsp1_uqid_i;
   assign cxl_d2h_rsp_frame0.D2H_Rsp0_Valid           = frame0_cxl_cache_d2h_rsp0_valid_i;
   assign cxl_d2h_rsp_frame0.D2H_Rsp0_Opcode          = frame0_cxl_cache_d2h_rsp0_opcode_i;
   assign cxl_d2h_rsp_frame0.D2H_Rsp0_Parity          = frame0_cxl_cache_d2h_rsp0_parity_i;
   assign cxl_d2h_rsp_frame0.D2H_Rsp0_Rsvd            = frame0_cxl_cache_d2h_rsp0_rsvd_i;
   assign cxl_d2h_rsp_frame0.D2H_Rsp0_UqID            = frame0_cxl_cache_d2h_rsp0_uqid_i;
   assign cxl_d2h_rsp_frame0_valid                    = frame0_cxl_cache_d2h_rsp_valid_i;
   assign frame0_cxl_cache_d2h_rsp_ready_o                    = cxl_d2h_rsp_frame0_ready;
   assign cxl_d2h_rsp_frame1.D2H_Rsp1_Valid           = frame1_cxl_cache_d2h_rsp1_valid_i;
   assign cxl_d2h_rsp_frame1.D2H_Rsp1_Opcode          = frame1_cxl_cache_d2h_rsp1_opcode_i;
   assign cxl_d2h_rsp_frame1.D2H_Rsp1_Parity          = frame1_cxl_cache_d2h_rsp1_parity_i;
   assign cxl_d2h_rsp_frame1.D2H_Rsp1_Rsvd            = frame1_cxl_cache_d2h_rsp1_rsvd_i;
   assign cxl_d2h_rsp_frame1.D2H_Rsp1_UqID            = frame1_cxl_cache_d2h_rsp1_uqid_i;
   assign cxl_d2h_rsp_frame1.D2H_Rsp0_Valid           = frame1_cxl_cache_d2h_rsp0_valid_i;
   assign cxl_d2h_rsp_frame1.D2H_Rsp0_Opcode          = frame1_cxl_cache_d2h_rsp0_opcode_i;
   assign cxl_d2h_rsp_frame1.D2H_Rsp0_Parity          = frame1_cxl_cache_d2h_rsp0_parity_i;
   assign cxl_d2h_rsp_frame1.D2H_Rsp0_Rsvd            = frame1_cxl_cache_d2h_rsp0_rsvd_i;
   assign cxl_d2h_rsp_frame1.D2H_Rsp0_UqID            = frame1_cxl_cache_d2h_rsp0_uqid_i;
   assign cxl_d2h_rsp_frame1_valid                    = frame1_cxl_cache_d2h_rsp_valid_i;
   assign frame1_cxl_cache_d2h_rsp_ready_o                    = cxl_d2h_rsp_frame1_ready;

   rnr_cxl_pkg::cxl_cache_d2h_data_tx_intf    cxl_d2h_data_frame0;                // 0                           = cxl_cache_mem_rx_frame0.cxl_mem. 1 ready
   wire                          cxl_d2h_data_frame0_valid;
   wire                          cxl_d2h_data_frame0_ready;
   rnr_cxl_pkg::cxl_cache_d2h_data_tx_intf    cxl_d2h_data_frame1;                // 1                           = cxl_cache_mem_rx_frame0.cxl_mem. 1 ready
   wire                          cxl_d2h_data_frame1_valid;
   wire                          cxl_d2h_data_frame1_ready;

   //interfaces_cxl_cache_d2h_data_tx
   assign cxl_d2h_data_frame0_valid                   = frame0_cxl_cache_d2h_valid_i;
   assign frame0_cxl_cache_d2h_data_ready_o                   = cxl_d2h_data_frame0_ready;
   assign cxl_d2h_data_frame0.D2H_Data_PushWrite      = frame0_cxl_cache_d2h_data_pushwrite_i;
   assign cxl_d2h_data_frame0.D2H_Data_UqID           = frame0_cxl_cache_d2h_data_uqid_i;
   assign cxl_d2h_data_frame0.D2H_Data_StrmID         = frame0_cxl_cache_d2h_data_strmid_i;
   assign cxl_d2h_data_frame0.D2H_Data_HdrParity      = frame0_cxl_cache_d2h_data_hdrparity_i;
   assign cxl_d2h_data_frame0.D2H_Data_Valid          = frame0_cxl_cache_d2h_data_valid_i;
   assign cxl_d2h_data_frame0.D2H_Data_Bogus          = frame0_cxl_cache_d2h_data_bogus_i;
   assign cxl_d2h_data_frame0.D2H_Data_Poison         = frame0_cxl_cache_d2h_data_poison_i;
   assign cxl_d2h_data_frame0.D2H_Data_DataParity     = frame0_cxl_cache_d2h_data_dataparity_i;
   assign cxl_d2h_data_frame0.D2H_Data_Rsvd           = frame0_cxl_cache_d2h_data_rsvd_i;
   assign cxl_d2h_data_frame0.D2H_Data_BEParity       = frame0_cxl_cache_d2h_data_beparity_i;
   assign cxl_d2h_data_frame0.D2H_Data_ByteEn         = frame0_cxl_cache_d2h_data_byteen_i;
   assign cxl_d2h_data_frame0.D2H_Data_Data           = frame0_cxl_cache_d2h_data_data_i;
   assign cxl_d2h_data_frame1_valid                   = frame1_cxl_cache_d2h_valid_i;
   assign frame1_cxl_cache_d2h_data_ready_o                   = cxl_d2h_data_frame1_ready;
   assign cxl_d2h_data_frame1.D2H_Data_PushWrite      = frame1_cxl_cache_d2h_data_pushwrite_i;
   assign cxl_d2h_data_frame1.D2H_Data_UqID           = frame1_cxl_cache_d2h_data_uqid_i;
   assign cxl_d2h_data_frame1.D2H_Data_StrmID         = frame1_cxl_cache_d2h_data_strmid_i;
   assign cxl_d2h_data_frame1.D2H_Data_HdrParity      = frame1_cxl_cache_d2h_data_hdrparity_i;
   assign cxl_d2h_data_frame1.D2H_Data_Valid          = frame1_cxl_cache_d2h_data_valid_i;
   assign cxl_d2h_data_frame1.D2H_Data_Bogus          = frame1_cxl_cache_d2h_data_bogus_i;
   assign cxl_d2h_data_frame1.D2H_Data_Poison         = frame1_cxl_cache_d2h_data_poison_i;
   assign cxl_d2h_data_frame1.D2H_Data_DataParity     = frame1_cxl_cache_d2h_data_dataparity_i;
   assign cxl_d2h_data_frame1.D2H_Data_Rsvd           = frame1_cxl_cache_d2h_data_rsvd_i;
   assign cxl_d2h_data_frame1.D2H_Data_BEParity       = frame1_cxl_cache_d2h_data_beparity_i;
   assign cxl_d2h_data_frame1.D2H_Data_ByteEn         = frame1_cxl_cache_d2h_data_byteen_i;
   assign cxl_d2h_data_frame1.D2H_Data_Data           = frame1_cxl_cache_d2h_data_data_i;


 // Declare Signals In Top Module
/* output */ logic          p1_reset_status_n;
/* input  */ logic          p1_pld_warm_rst_rdy_i;
/* output */ logic          p1_pld_link_req_rst_o;
/* input  */ logic          p2_pld_warm_rst_rdy_i;
/* output */ logic          p2_pld_link_req_rst_o;
/* output */ logic          p2_reset_status_n;
/* input  */ logic          p3_pld_warm_rst_rdy_i;
/* output */ logic          p3_pld_link_req_rst_o;
/* output */ logic          p3_reset_status_n;
/* input  */ logic          p0_app_rst_n;
/* input  */ logic          p1_app_rst_n;
/* input  */ logic          p2_app_rst_n;
/* input  */ logic          p3_app_rst_n;
/* input  */ logic          cxl_app_rst_n;
/* input  */ logic          cxl_pll_locked_i;
/* input  */ logic          i_clk;
/* input  */ logic          i_rst_n;
/* input  */ logic          i_rx_dsk_clear;
/* input  */ logic          i_tx_dsk_clear;
/* output */ logic          rx_deskew_valid;
/* output */ logic          rx_deskew_done;
/* output */ logic          rx_deskew_lock_err;
/* output */ logic [31:0]   rx_dsk_monitor_err;
/* output */ logic          o_ptm_clk_updated;
/* output */ logic          o_ptm_context_valid;
/* output */ logic [63:0]   o_ptm_local_clock;
/* input  */ logic          i_ptm_manual_update;
/* output */ logic          rx_st0_dvalid;
/* output */ logic          rx_st1_dvalid;
/* output */ logic          rx_st2_dvalid;
/* output */ logic          rx_st3_dvalid;
/* output */ logic          rx_st0_sop;
/* output */ logic          rx_st1_sop;
/* output */ logic          rx_st2_sop;
/* output */ logic          rx_st3_sop;
/* output */ logic          rx_st0_eop;
/* output */ logic          rx_st1_eop;
/* output */ logic          rx_st2_eop;
/* output */ logic          rx_st3_eop;
/* output */ logic          rx_st0_passthrough;
/* output */ logic          rx_st1_passthrough;
/* output */ logic          rx_st2_passthrough;
/* output */ logic          rx_st3_passthrough;
/* output */ logic [255:0]  rx_st0_data;
/* output */ logic [255:0]  rx_st1_data;
/* output */ logic [255:0]  rx_st2_data;
/* output */ logic [255:0]  rx_st3_data;
/* output */ logic [7:0]    rx_st0_data_parity;
/* output */ logic [7:0]    rx_st1_data_parity;
/* output */ logic [7:0]    rx_st2_data_parity;
/* output */ logic [7:0]    rx_st3_data_parity;
/* output */ logic [127:0]  rx_st0_hdr;
/* output */ logic [127:0]  rx_st1_hdr;
/* output */ logic [127:0]  rx_st2_hdr;
/* output */ logic [127:0]  rx_st3_hdr;
/* output */ logic [3:0]    rx_st0_hdr_parity;
/* output */ logic [3:0]    rx_st1_hdr_parity;
/* output */ logic [3:0]    rx_st2_hdr_parity;
/* output */ logic [3:0]    rx_st3_hdr_parity;
/* output */ logic          rx_st0_hvalid;
/* output */ logic          rx_st1_hvalid;
/* output */ logic          rx_st2_hvalid;
/* output */ logic          rx_st3_hvalid;
/* output */ logic [31:0]   rx_st0_prefix;
/* output */ logic [31:0]   rx_st1_prefix;
/* output */ logic [31:0]   rx_st2_prefix;
/* output */ logic [31:0]   rx_st3_prefix;
/* output */ logic          rx_st0_prefix_parity;
/* output */ logic          rx_st1_prefix_parity;
/* output */ logic          rx_st2_prefix_parity;
/* output */ logic          rx_st3_prefix_parity;
/* output */ logic [11:0]   rx_st0_rssai_prefix;
/* output */ logic [11:0]   rx_st1_rssai_prefix;
/* output */ logic [11:0]   rx_st2_rssai_prefix;
/* output */ logic [11:0]   rx_st3_rssai_prefix;
/* output */ logic          rx_st0_rssai_prefix_parity;
/* output */ logic          rx_st1_rssai_prefix_parity;
/* output */ logic          rx_st2_rssai_prefix_parity;
/* output */ logic          rx_st3_rssai_prefix_parity;
/* output */ logic [1:0]    rx_st0_pvalid;
/* output */ logic [1:0]    rx_st1_pvalid;
/* output */ logic [1:0]    rx_st2_pvalid;
/* output */ logic [1:0]    rx_st3_pvalid;
/* output */ logic [2:0]    rx_st0_bar;
/* output */ logic [2:0]    rx_st1_bar;
/* output */ logic [2:0]    rx_st2_bar;
/* output */ logic [2:0]    rx_st3_bar;
/* output */ logic          rx_st0_vfactive;
/* output */ logic          rx_st1_vfactive;
/* output */ logic          rx_st2_vfactive;
/* output */ logic          rx_st3_vfactive;
/* output */ logic [10:0]   rx_st0_vfnum;
/* output */ logic [10:0]   rx_st1_vfnum;
/* output */ logic [10:0]   rx_st2_vfnum;
/* output */ logic [10:0]   rx_st3_vfnum;
/* output */ logic [2:0]    rx_st0_pfnum;
/* output */ logic [2:0]    rx_st1_pfnum;
/* output */ logic [2:0]    rx_st2_pfnum;
/* output */ logic [2:0]    rx_st3_pfnum;
/* output */ logic          rx_st0_chnum;
/* output */ logic          rx_st1_chnum;
/* output */ logic          rx_st2_chnum;
/* output */ logic          rx_st3_chnum;
/* output */ logic          rx_st0_misc_parity;
/* output */ logic          rx_st1_misc_parity;
/* output */ logic          rx_st2_misc_parity;
/* output */ logic          rx_st3_misc_parity;
/* output */ logic [2:0]    rx_st0_empty;
/* output */ logic [2:0]    rx_st1_empty;
/* output */ logic [2:0]    rx_st2_empty;
/* output */ logic [2:0]    rx_st3_empty;
/* input  */ logic [2:0]    rx_st_Hcrdt_update;
/* input  */ logic [2:0]    rx_st_Hcrdt_ch;
/* input  */ logic [5:0]    rx_st_Hcrdt_update_cnt;
/* input  */ logic [2:0]    rx_st_Hcrdt_init;
/* output */ logic [2:0]    rx_st_Hcrdt_init_ack;
/* input  */ logic [2:0]    rx_st_Dcrdt_update;
/* input  */ logic [2:0]    rx_st_Dcrdt_ch;
/* input  */ logic [11:0]   rx_st_Dcrdt_update_cnt;
/* input  */ logic [2:0]    rx_st_Dcrdt_init;
/* output */ logic [2:0]    rx_st_Dcrdt_init_ack;
/* output */ logic          tx_st_ready;
/* input  */ logic          tx_st0_dvalid;
/* input  */ logic          tx_st1_dvalid;
/* input  */ logic          tx_st2_dvalid;
/* input  */ logic          tx_st3_dvalid;
/* input  */ logic          tx_st0_sop;
/* input  */ logic          tx_st1_sop;
/* input  */ logic          tx_st2_sop;
/* input  */ logic          tx_st3_sop;
/* input  */ logic          tx_st0_eop;
/* input  */ logic          tx_st1_eop;
/* input  */ logic          tx_st2_eop;
/* input  */ logic          tx_st3_eop;
/* input  */ logic          tx_st0_passthrough;
/* input  */ logic          tx_st1_passthrough;
/* input  */ logic          tx_st2_passthrough;
/* input  */ logic          tx_st3_passthrough;
/* input  */ logic [255:0]  tx_st0_data;
/* input  */ logic [255:0]  tx_st1_data;
/* input  */ logic [255:0]  tx_st2_data;
/* input  */ logic [255:0]  tx_st3_data;
/* input  */ logic [7:0]    tx_st0_data_parity;
/* input  */ logic [7:0]    tx_st1_data_parity;
/* input  */ logic [7:0]    tx_st2_data_parity;
/* input  */ logic [7:0]    tx_st3_data_parity;
/* input  */ logic [127:0]  tx_st0_hdr;
/* input  */ logic [127:0]  tx_st1_hdr;
/* input  */ logic [127:0]  tx_st2_hdr;
/* input  */ logic [127:0]  tx_st3_hdr;
/* input  */ logic [3:0]    tx_st0_hdr_parity;
/* input  */ logic [3:0]    tx_st1_hdr_parity;
/* input  */ logic [3:0]    tx_st2_hdr_parity;
/* input  */ logic [3:0]    tx_st3_hdr_parity;
/* input  */ logic          tx_st0_hvalid;
/* input  */ logic          tx_st1_hvalid;
/* input  */ logic          tx_st2_hvalid;
/* input  */ logic          tx_st3_hvalid;
/* input  */ logic [31:0]   tx_st0_prefix;
/* input  */ logic [31:0]   tx_st1_prefix;
/* input  */ logic [31:0]   tx_st2_prefix;
/* input  */ logic [31:0]   tx_st3_prefix;
/* input  */ logic          tx_st0_prefix_parity;
/* input  */ logic          tx_st1_prefix_parity;
/* input  */ logic          tx_st2_prefix_parity;
/* input  */ logic          tx_st3_prefix_parity;
/* input  */ logic [11:0]   tx_st0_rssai_prefix;
/* input  */ logic [11:0]   tx_st1_rssai_prefix;
/* input  */ logic [11:0]   tx_st2_rssai_prefix;
/* input  */ logic [11:0]   tx_st3_rssai_prefix;
/* input  */ logic          tx_st0_rssai_prefix_parity;
/* input  */ logic          tx_st1_rssai_prefix_parity;
/* input  */ logic          tx_st2_rssai_prefix_parity;
/* input  */ logic          tx_st3_rssai_prefix_parity;
/* input  */ logic [1:0]    tx_st0_pvalid;
/* input  */ logic [1:0]    tx_st1_pvalid;
/* input  */ logic [1:0]    tx_st2_pvalid;
/* input  */ logic [1:0]    tx_st3_pvalid;
/* input  */ logic [2:0]    tx_st0_empty;
/* input  */ logic [2:0]    tx_st1_empty;
/* input  */ logic [2:0]    tx_st2_empty;
/* input  */ logic [2:0]    tx_st3_empty;
/* output */ logic [2:0]    tx_st_Hcrdt_update;
/* output */ logic [2:0]    tx_st_Hcrdt_vc;
/* output */ logic [5:0]    tx_st_Hcrdt_update_cnt;
/* output */ logic [2:0]    tx_st_Hcrdt_init;
/* input  */ logic [2:0]    tx_st_Hcrdt_init_ack;
/* output */ logic [2:0]    tx_st_Dcrdt_update;
/* output */ logic [2:0]    tx_st_Dcrdt_vc;
/* output */ logic [11:0]   tx_st_Dcrdt_update_cnt;
/* output */ logic [2:0]    tx_st_Dcrdt_init;
/* input  */ logic [2:0]    tx_st_Dcrdt_init_ack;
/* output */ logic [3:0]    o_ial_ch18_ext_fsr;
/* output */ logic [7:0]    o_ial_ch18_ext_ssr;
/* output */ logic [2:0]    o_ial_ch18_fsr;
/* output */ logic [64:0]   o_ial_ch18_ssr;
/* output */ logic [3:0]    o_ial_ch19_ext_fsr;
/* output */ logic [7:0]    o_ial_ch19_ext_ssr;
/* output */ logic [2:0]    o_ial_ch19_fsr;
/* output */ logic [64:0]   o_ial_ch19_ssr;
/* output */ logic [5:0]    o_ial_ch1_async_direct;
/* output */ logic [3:0]    o_ial_ch20_ext_fsr;
/* output */ logic [7:0]    o_ial_ch20_ext_ssr;
/* output */ logic [2:0]    o_ial_ch20_fsr;
/* output */ logic [64:0]   o_ial_ch20_ssr;
/* output */ logic [3:0]    o_ial_ch21_ext_fsr;
/* output */ logic [7:0]    o_ial_ch21_ext_ssr;
/* output */ logic [2:0]    o_ial_ch21_fsr;
/* output */ logic [64:0]   o_ial_ch21_ssr;
/* output */ logic [3:0]    o_ial_ch22_ext_fsr;
/* output */ logic [7:0]    o_ial_ch22_ext_ssr;
/* output */ logic [2:0]    o_ial_ch22_fsr;
/* output */ logic [64:0]   o_ial_ch22_ssr;
/* output */ logic [3:0]    o_ial_ch23_ext_fsr;
/* output */ logic [7:0]    o_ial_ch23_ext_ssr;
/* output */ logic [2:0]    o_ial_ch23_fsr;
/* output */ logic [64:0]   o_ial_ch23_ssr;
/* output */ logic [5:0]    o_ial_ch2_async_direct;
/* output */ logic [5:0]    o_ial_ch3_async_direct;
/* input  */ logic [3:0]    i_ial_ch19_ext_fsr;
/* input  */ logic [39:0]   i_ial_ch19_ext_ssr;
/* input  */ logic [2:0]    i_ial_ch19_fsr;
/* input  */ logic [60:0]   i_ial_ch19_ssr;
/* input  */ logic [3:0]    i_ial_ch20_ext_fsr;
/* input  */ logic [39:0]   i_ial_ch20_ext_ssr;
/* input  */ logic [2:0]    i_ial_ch20_fsr;
/* input  */ logic [60:0]   i_ial_ch20_ssr;
/* input  */ logic [3:0]    i_ial_ch21_ext_fsr;
/* input  */ logic [39:0]   i_ial_ch21_ext_ssr;
/* input  */ logic [2:0]    i_ial_ch21_fsr;
/* input  */ logic [60:0]   i_ial_ch21_ssr;
/* input  */ logic [7:0]    i_ial_ch22_async_direct;
/* input  */ logic [3:0]    i_ial_ch22_ext_fsr;
/* input  */ logic [39:0]   i_ial_ch22_ext_ssr;
/* input  */ logic [2:0]    i_ial_ch22_fsr;
/* input  */ logic [60:0]   i_ial_ch22_ssr;
/* input  */ logic [7:0]    i_ial_ch23_async_direct;
/* input  */ logic [3:0]    i_ial_ch23_ext_fsr;
/* input  */ logic [39:0]   i_ial_ch23_ext_ssr;
/* input  */ logic [2:0]    i_ial_ch23_fsr;
/* input  */ logic [60:0]   i_ial_ch23_ssr;
/* output */ logic [5:0]    o_ch0_async_direct_aib2pld;
/* output */ logic [5:0]    o_ch1_async_direct_aib2pld;
/* output */ logic [5:0]    o_ch2_async_direct_aib2pld;
/* output */ logic [5:0]    o_ch3_async_direct_aib2pld;
/* output */ logic [5:0]    o_ch4_async_direct_aib2pld;
/* output */ logic [5:0]    o_ch5_async_direct_aib2pld;
/* output */ logic [5:0]    o_ch6_async_direct_aib2pld;
/* output */ logic [4:0]    o_ch7_async_direct_aib2pld;
/* output */ logic [6:0]    o_ch11_fsr_aib2pld;
/* output */ logic [6:0]    o_ch9_fsr_aib2pld;
/* input  */ logic [7:0]    i_ch0_async_direct_pld2aib;
/* input  */ logic [7:0]    i_ch1_async_direct_pld2aib;
/* input  */ logic [7:0]    i_ch2_async_direct_pld2aib;
/* input  */ logic [7:0]    i_ch3_async_direct_pld2aib;
/* input  */ logic [7:0]    i_ch4_async_direct_pld2aib;
/* input  */ logic [7:0]    i_ch5_async_direct_pld2aib;
/* input  */ logic [7:0]    i_ch6_async_direct_pld2aib;
/* input  */ logic [7:0]    i_ch7_async_direct_pld2aib;
/* input  */ logic [6:0]    i_ch11_fsr_pld2aib;
/* input  */ logic [6:0]    i_ch9_fsr_pld2aib;
//* output */ logic [7:0]    o_user_avmm_readdata;
//* output */ logic          o_user_avmm_readdatavalid;
//* output */ logic          o_user_avmm_writedone;
//* input  */ logic          i_user_avmm2_clk_rowclk;
//* input  */ logic          i_ch0_user_avmm1_clk_rowclk;
//* input  */ logic          i_user_avmm_read;
//* input  */ logic [20:0]   i_user_avmm_reg_addr;
//* input  */ logic          i_user_avmm_write;
//* input  */ logic [7:0]    i_user_avmm_writedata;
/* input  */ logic [77:0]   ch13_pipe_direct_tx_octet1;
/* input  */ logic [77:0]   ch14_pipe_direct_tx_octet1;
/* input  */ logic [77:0]   ch15_pipe_direct_tx_octet1;
/* input  */ logic [77:0]   ch16_pipe_direct_tx_octet1;
/* input  */ logic [77:0]   ch17_pipe_direct_tx_octet1;
/* input  */ logic [77:0]   ch18_pipe_direct_tx_octet1;
/* input  */ logic [77:0]   ch19_pipe_direct_tx_octet1;
/* input  */ logic [77:0]   ch20_pipe_direct_tx_octet1;
/* input  */ logic [77:0]   ch21_pipe_direct_tx_octet1;
/* input  */ logic [77:0]   ch22_pipe_direct_tx_octet1;
/* output */ logic [77:0]   ch13_pipe_direct_rx_octet1;
/* output */ logic [77:0]   ch14_pipe_direct_rx_octet1;
/* output */ logic [77:0]   ch15_pipe_direct_rx_octet1;
/* output */ logic [77:0]   ch16_pipe_direct_rx_octet1;
/* output */ logic [77:0]   ch17_pipe_direct_rx_octet1;
/* output */ logic [77:0]   ch18_pipe_direct_rx_octet1;
/* output */ logic [77:0]   ch19_pipe_direct_rx_octet1;
/* output */ logic [77:0]   ch20_pipe_direct_rx_octet1;
/* output */ logic [77:0]   ch21_pipe_direct_rx_octet1;
/* output */ logic [77:0]   ch22_pipe_direct_rx_octet1;
/* output */ logic          ch15_pipe_direct_tx_octet1_pwrdwn_status_l8;
/* output */ logic          ch16_pipe_direct_tx_octet1_pwrdwn_status_l9;
/* output */ logic          ch17_pipe_direct_tx_octet1_pwrdwn_status_l10;
/* output */ logic          ch18_pipe_direct_tx_octet1_pwrdwn_status_l11;
/* output */ logic          ch19_pipe_direct_tx_octet1_pwrdwn_status_l12;
/* output */ logic          ch20_pipe_direct_tx_octet1_pwrdwn_status_l13;
/* output */ logic          ch21_pipe_direct_tx_octet1_pwrdwn_status_l14;
/* output */ logic          ch22_pipe_direct_tx_octet1_pwrdwn_status_l15;
/* input  */ logic          ch15_pipe_direct_tx_octet1_PLD_PCS_rst_n_l8;
/* input  */ logic          ch16_pipe_direct_tx_octet1_PLD_PCS_rst_n_l9;
/* input  */ logic          ch17_pipe_direct_tx_octet1_PLD_PCS_rst_n_l10;
/* input  */ logic          ch18_pipe_direct_tx_octet1_PLD_PCS_rst_n_l11;
/* input  */ logic          ch19_pipe_direct_tx_octet1_PLD_PCS_rst_n_l12;
/* input  */ logic          ch20_pipe_direct_tx_octet1_PLD_PCS_rst_n_l13;
/* input  */ logic          ch21_pipe_direct_tx_octet1_PLD_PCS_rst_n_l14;
/* input  */ logic          ch22_pipe_direct_tx_octet1_PLD_PCS_rst_n_l15;
/* output */ logic          ch15_pipe_direct_rx_octet1_RXElecIdle_l8;
/* output */ logic          ch16_pipe_direct_rx_octet1_RXElecIdle_l9;
/* output */ logic          ch17_pipe_direct_rx_octet1_RXElecIdle_l10;
/* output */ logic          ch18_pipe_direct_rx_octet1_RXElecIdle_l11;
/* output */ logic          ch19_pipe_direct_rx_octet1_RXElecIdle_l12;
/* output */ logic          ch20_pipe_direct_rx_octet1_RXElecIdle_l13;
/* output */ logic          ch21_pipe_direct_rx_octet1_RXElecIdle_l14;
/* output */ logic          ch22_pipe_direct_rx_octet1_RXElecIdle_l15;
/* output */ logic          ch15_pipe_direct_rx_octet1_rx_cdrlock2data_l8;
/* output */ logic          ch16_pipe_direct_rx_octet1_rx_cdrlock2data_l9;
/* output */ logic          ch17_pipe_direct_rx_octet1_rx_cdrlock2data_l10;
/* output */ logic          ch18_pipe_direct_rx_octet1_rx_cdrlock2data_l11;
/* output */ logic          ch19_pipe_direct_rx_octet1_rx_cdrlock2data_l12;
/* output */ logic          ch20_pipe_direct_rx_octet1_rx_cdrlock2data_l13;
/* output */ logic          ch21_pipe_direct_rx_octet1_rx_cdrlock2data_l14;
/* output */ logic          ch22_pipe_direct_rx_octet1_rx_cdrlock2data_l15;
/* output */ logic          ch15_pipe_direct_rx_octet1_rx_cdrlockstatus_l8;
/* output */ logic          ch16_pipe_direct_rx_octet1_rx_cdrlockstatus_l9;
/* output */ logic          ch17_pipe_direct_rx_octet1_rx_cdrlockstatus_l10;
/* output */ logic          ch18_pipe_direct_rx_octet1_rx_cdrlockstatus_l11;
/* output */ logic          ch19_pipe_direct_rx_octet1_rx_cdrlockstatus_l12;
/* output */ logic          ch20_pipe_direct_rx_octet1_rx_cdrlockstatus_l13;
/* output */ logic          ch21_pipe_direct_rx_octet1_rx_cdrlockstatus_l14;
/* output */ logic          ch22_pipe_direct_rx_octet1_rx_cdrlockstatus_l15;
/* output */ logic          pipe_direct_rx_octet1_synthfast_lockstatus1;
/* output */ logic          pipe_direct_rx_octet1_synthfast_ready1;
/* output */ logic          pipe_direct_rx_octet1_synthslow_lockstatus1;
/* output */ logic          pipe_direct_rx_octet1_synthslow_ready1;
/* output */ logic          ch13_pipe_direct_pld_fabric_tx_transfer_en;
/* output */ logic          ch13_pipe_direct_pld_hssi_osc_transfer_en;
/* output */ logic          ch13_pipe_direct_pld_hssi_rx_transfer_en;
/* input  */ logic          ch13_pipe_direct_pld_adapter_rx_pld_rst_n;
/* input  */ logic          ch13_pipe_direct_pld_rx_dll_lock_req;
/* input  */ logic          ch13_pipe_direct_pld_adapter_tx_pld_rst_n;
/* input  */ logic          ch13_pipe_direct_pld_tx_dll_lock_req;
/* output */ logic          ch14_pipe_direct_pld_fabric_tx_transfer_en;
/* output */ logic          ch14_pipe_direct_pld_hssi_osc_transfer_en;
/* output */ logic          ch14_pipe_direct_pld_hssi_rx_transfer_en;
/* input  */ logic          ch14_pipe_direct_pld_adapter_rx_pld_rst_n;
/* input  */ logic          ch14_pipe_direct_pld_rx_dll_lock_req;
/* input  */ logic          ch14_pipe_direct_pld_adapter_tx_pld_rst_n;
/* input  */ logic          ch14_pipe_direct_pld_tx_dll_lock_req;
/* output */ logic          ch15_pipe_direct_pld_fabric_tx_transfer_en;
/* output */ logic          ch15_pipe_direct_pld_hssi_osc_transfer_en;
/* output */ logic          ch15_pipe_direct_pld_hssi_rx_transfer_en;
/* input  */ logic          ch15_pipe_direct_pld_adapter_rx_pld_rst_n;
/* input  */ logic          ch15_pipe_direct_pld_rx_dll_lock_req;
/* input  */ logic          ch15_pipe_direct_pld_adapter_tx_pld_rst_n;
/* input  */ logic          ch15_pipe_direct_pld_tx_dll_lock_req;
/* output */ logic          ch16_pipe_direct_pld_fabric_tx_transfer_en;
/* output */ logic          ch16_pipe_direct_pld_hssi_osc_transfer_en;
/* output */ logic          ch16_pipe_direct_pld_hssi_rx_transfer_en;
/* input  */ logic          ch16_pipe_direct_pld_adapter_rx_pld_rst_n;
/* input  */ logic          ch16_pipe_direct_pld_rx_dll_lock_req;
/* input  */ logic          ch16_pipe_direct_pld_adapter_tx_pld_rst_n;
/* input  */ logic          ch16_pipe_direct_pld_tx_dll_lock_req;
/* output */ logic          ch17_pipe_direct_pld_fabric_tx_transfer_en;
/* output */ logic          ch17_pipe_direct_pld_hssi_osc_transfer_en;
/* output */ logic          ch17_pipe_direct_pld_hssi_rx_transfer_en;
/* input  */ logic          ch17_pipe_direct_pld_adapter_rx_pld_rst_n;
/* input  */ logic          ch17_pipe_direct_pld_rx_dll_lock_req;
/* input  */ logic          ch17_pipe_direct_pld_adapter_tx_pld_rst_n;
/* input  */ logic          ch17_pipe_direct_pld_tx_dll_lock_req;
/* output */ logic          ch18_pipe_direct_pld_fabric_tx_transfer_en;
/* output */ logic          ch18_pipe_direct_pld_hssi_osc_transfer_en;
/* output */ logic          ch18_pipe_direct_pld_hssi_rx_transfer_en;
/* input  */ logic          ch18_pipe_direct_pld_adapter_rx_pld_rst_n;
/* input  */ logic          ch18_pipe_direct_pld_rx_dll_lock_req;
/* input  */ logic          ch18_pipe_direct_pld_adapter_tx_pld_rst_n;
/* input  */ logic          ch18_pipe_direct_pld_tx_dll_lock_req;
/* output */ logic          ch19_pipe_direct_pld_fabric_tx_transfer_en;
/* output */ logic          ch19_pipe_direct_pld_hssi_osc_transfer_en;
/* output */ logic          ch19_pipe_direct_pld_hssi_rx_transfer_en;
/* input  */ logic          ch19_pipe_direct_pld_adapter_rx_pld_rst_n;
/* input  */ logic          ch19_pipe_direct_pld_rx_dll_lock_req;
/* input  */ logic          ch19_pipe_direct_pld_adapter_tx_pld_rst_n;
/* input  */ logic          ch19_pipe_direct_pld_tx_dll_lock_req;
/* output */ logic          ch20_pipe_direct_pld_fabric_tx_transfer_en;
/* output */ logic          ch20_pipe_direct_pld_hssi_osc_transfer_en;
/* output */ logic          ch20_pipe_direct_pld_hssi_rx_transfer_en;
/* input  */ logic          ch20_pipe_direct_pld_adapter_rx_pld_rst_n;
/* input  */ logic          ch20_pipe_direct_pld_rx_dll_lock_req;
/* input  */ logic          ch20_pipe_direct_pld_adapter_tx_pld_rst_n;
/* input  */ logic          ch20_pipe_direct_pld_tx_dll_lock_req;
/* output */ logic          ch21_pipe_direct_pld_fabric_tx_transfer_en;
/* output */ logic          ch21_pipe_direct_pld_hssi_osc_transfer_en;
/* output */ logic          ch21_pipe_direct_pld_hssi_rx_transfer_en;
/* input  */ logic          ch21_pipe_direct_pld_adapter_rx_pld_rst_n;
/* input  */ logic          ch21_pipe_direct_pld_rx_dll_lock_req;
/* input  */ logic          ch21_pipe_direct_pld_adapter_tx_pld_rst_n;
/* input  */ logic          ch21_pipe_direct_pld_tx_dll_lock_req;
/* output */ logic          ch22_pipe_direct_pld_fabric_tx_transfer_en;
/* output */ logic          ch22_pipe_direct_pld_hssi_osc_transfer_en;
/* output */ logic          ch22_pipe_direct_pld_hssi_rx_transfer_en;
/* input  */ logic          ch22_pipe_direct_pld_adapter_rx_pld_rst_n;
/* input  */ logic          ch22_pipe_direct_pld_rx_dll_lock_req;
/* input  */ logic          ch22_pipe_direct_pld_adapter_tx_pld_rst_n;
/* input  */ logic          ch22_pipe_direct_pld_tx_dll_lock_req;
/* output */ logic          ch13_pipe_direct_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          ch13_pipe_direct_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          ch14_pipe_direct_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          ch14_pipe_direct_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          ch15_pipe_direct_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          ch15_pipe_direct_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          ch16_pipe_direct_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          ch16_pipe_direct_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          ch17_pipe_direct_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          ch17_pipe_direct_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          ch18_pipe_direct_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          ch18_pipe_direct_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          ch19_pipe_direct_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          ch19_pipe_direct_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          ch20_pipe_direct_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          ch20_pipe_direct_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          ch21_pipe_direct_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          ch21_pipe_direct_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          ch22_pipe_direct_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          ch22_pipe_direct_pld_pcs_tx_clk_out1_dcm;
/* input  */ logic          ch13_pipe_direct_pld_rx_clk1_dcm;
/* input  */ logic          ch13_pipe_direct_pld_tx_clk1_dcm;
/* input  */ logic          ch14_pipe_direct_pld_rx_clk1_dcm;
/* input  */ logic          ch14_pipe_direct_pld_tx_clk1_dcm;
/* input  */ logic          ch15_pipe_direct_pld_rx_clk1_dcm;
/* input  */ logic          ch15_pipe_direct_pld_tx_clk1_dcm;
/* input  */ logic          ch16_pipe_direct_pld_rx_clk1_dcm;
/* input  */ logic          ch16_pipe_direct_pld_tx_clk1_dcm;
/* input  */ logic          ch17_pipe_direct_pld_rx_clk1_dcm;
/* input  */ logic          ch17_pipe_direct_pld_tx_clk1_dcm;
/* input  */ logic          ch18_pipe_direct_pld_rx_clk1_dcm;
/* input  */ logic          ch18_pipe_direct_pld_tx_clk1_dcm;
/* input  */ logic          ch19_pipe_direct_pld_rx_clk1_dcm;
/* input  */ logic          ch19_pipe_direct_pld_tx_clk1_dcm;
/* input  */ logic          ch20_pipe_direct_pld_rx_clk1_dcm;
/* input  */ logic          ch20_pipe_direct_pld_tx_clk1_dcm;
/* input  */ logic          ch21_pipe_direct_pld_rx_clk1_dcm;
/* input  */ logic          ch21_pipe_direct_pld_tx_clk1_dcm;
/* input  */ logic          ch22_pipe_direct_pld_rx_clk1_dcm;
/* input  */ logic          ch22_pipe_direct_pld_tx_clk1_dcm;
/* input  */ logic [2:0]    ial_phy_tx_fsr_0__tx_chnl_fsr;
/* input  */ logic [3:0]    ial_phy_tx_fsr_0__tx_ext_fsr;
/* input  */ logic [2:0]    ial_phy_tx_fsr_1__tx_chnl_fsr;
/* input  */ logic [3:0]    ial_phy_tx_fsr_1__tx_ext_fsr;
/* input  */ logic [2:0]    ial_phy_tx_fsr_2__tx_chnl_fsr;
/* input  */ logic [3:0]    ial_phy_tx_fsr_2__tx_ext_fsr;
/* input  */ logic [2:0]    ial_phy_tx_fsr_3__tx_chnl_fsr;
/* input  */ logic [3:0]    ial_phy_tx_fsr_3__tx_ext_fsr;
/* input  */ logic [2:0]    ial_phy_tx_fsr_4__tx_chnl_fsr;
/* input  */ logic [3:0]    ial_phy_tx_fsr_4__tx_ext_fsr;
/* input  */ logic [2:0]    ial_phy_tx_fsr_5__tx_chnl_fsr;
/* input  */ logic [3:0]    ial_phy_tx_fsr_5__tx_ext_fsr;
/* input  */ logic [2:0]    pcie_phy_tx_fsr_10__tx_chnl_fsr;
/* input  */ logic [3:0]    pcie_phy_tx_fsr_10__tx_ext_fsr;
/* input  */ logic [2:0]    pcie_phy_tx_fsr_11__tx_chnl_fsr;
/* input  */ logic [3:0]    pcie_phy_tx_fsr_11__tx_ext_fsr;
/* output */ logic          o_ch0_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch0_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch0_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch0_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch0_pld_pma_hclk_hioint;
/* output */ logic          o_ch0_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch0_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch10_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch10_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch10_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch10_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch10_pld_pma_hclk_hioint;
/* output */ logic          o_ch10_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch10_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch11_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch11_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch11_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch11_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch11_pld_pma_hclk_hioint;
/* output */ logic          o_ch11_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch11_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch12_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch12_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch12_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch12_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch12_pld_pma_hclk_hioint;
/* output */ logic          o_ch12_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch12_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch13_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch13_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch13_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch13_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch13_pld_pma_hclk_hioint;
/* output */ logic          o_ch13_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch13_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch14_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch14_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch14_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch14_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch14_pld_pma_hclk_hioint;
/* output */ logic          o_ch14_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch14_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch15_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch15_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch15_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch15_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch15_pld_pma_hclk_hioint;
/* output */ logic          o_ch15_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch15_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch16_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch16_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch16_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch16_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch16_pld_pma_hclk_hioint;
/* output */ logic          o_ch16_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch16_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch17_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch17_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch17_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch17_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch17_pld_pma_hclk_hioint;
/* output */ logic          o_ch17_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch17_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch18_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch18_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch18_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch18_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch18_pld_pma_hclk_hioint;
/* output */ logic          o_ch18_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch18_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch19_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch19_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch19_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch19_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch19_pld_pma_hclk_hioint;
/* output */ logic          o_ch19_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch19_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch1_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch1_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch1_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch1_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch1_pld_pma_hclk_hioint;
/* output */ logic          o_ch1_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch1_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch20_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch20_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch20_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch20_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch20_pld_pma_hclk_hioint;
/* output */ logic          o_ch20_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch20_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch21_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch21_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch21_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch21_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch21_pld_pma_hclk_hioint;
/* output */ logic          o_ch21_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch21_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch22_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch22_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch22_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch22_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch22_pld_pma_hclk_hioint;
/* output */ logic          o_ch22_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch22_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch23_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch23_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch23_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch23_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch23_pld_pma_hclk_hioint;
/* output */ logic          o_ch23_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch23_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch2_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch2_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch2_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch2_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch2_pld_pma_hclk_hioint;
/* output */ logic          o_ch2_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch2_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch3_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch3_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch3_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch3_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch3_pld_pma_hclk_hioint;
/* output */ logic          o_ch3_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch3_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch4_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch4_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch4_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch4_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch4_pld_pma_hclk_hioint;
/* output */ logic          o_ch4_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch4_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch5_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch5_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch5_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch5_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch5_pld_pma_hclk_hioint;
/* output */ logic          o_ch5_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch5_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch6_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch6_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch6_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch6_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch6_pld_pma_hclk_hioint;
/* output */ logic          o_ch6_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch6_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch7_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch7_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch7_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch7_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch7_pld_pma_hclk_hioint;
/* output */ logic          o_ch7_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch7_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch8_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch8_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch8_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch8_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch8_pld_pma_hclk_hioint;
/* output */ logic          o_ch8_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch8_pld_pma_internal_clk2_hioint;
/* output */ logic          o_ch9_pld_pcs_rx_clk_out1_hioint;
/* output */ logic          o_ch9_pld_pcs_rx_clk_out2_hioint;
/* output */ logic          o_ch9_pld_pcs_tx_clk_out1_hioint;
/* output */ logic          o_ch9_pld_pcs_tx_clk_out2_hioint;
/* output */ logic          o_ch9_pld_pma_hclk_hioint;
/* output */ logic          o_ch9_pld_pma_internal_clk1_hioint;
/* output */ logic          o_ch9_pld_pma_internal_clk2_hioint;
/* input  */ logic          i_ch0_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch0_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch0_pld_sclk1_rowclk;
/* input  */ logic          i_ch0_pld_sclk2_rowclk;
/* input  */ logic          i_ch10_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch10_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch10_pld_sclk1_rowclk;
/* input  */ logic          i_ch10_pld_sclk2_rowclk;
/* input  */ logic          i_ch10_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch10_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch11_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch11_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch11_pld_sclk1_rowclk;
/* input  */ logic          i_ch11_pld_sclk2_rowclk;
/* input  */ logic          i_ch11_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch11_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch12_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch12_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch12_pld_sclk1_rowclk;
/* input  */ logic          i_ch12_pld_sclk2_rowclk;
/* input  */ logic          i_ch12_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch12_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch13_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch13_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch13_pld_sclk1_rowclk;
/* input  */ logic          i_ch13_pld_sclk2_rowclk;
/* input  */ logic          i_ch13_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch13_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch14_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch14_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch14_pld_sclk1_rowclk;
/* input  */ logic          i_ch14_pld_sclk2_rowclk;
/* input  */ logic          i_ch14_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch14_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch15_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch15_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch15_pld_sclk1_rowclk;
/* input  */ logic          i_ch15_pld_sclk2_rowclk;
/* input  */ logic          i_ch15_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch15_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch16_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch16_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch16_pld_sclk1_rowclk;
/* input  */ logic          i_ch16_pld_sclk2_rowclk;
/* input  */ logic          i_ch16_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch16_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch17_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch17_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch17_pld_sclk1_rowclk;
/* input  */ logic          i_ch17_pld_sclk2_rowclk;
/* input  */ logic          i_ch17_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch17_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch18_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch18_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch18_pld_sclk1_rowclk;
/* input  */ logic          i_ch18_pld_sclk2_rowclk;
/* input  */ logic          i_ch18_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch18_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch19_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch19_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch19_pld_sclk1_rowclk;
/* input  */ logic          i_ch19_pld_sclk2_rowclk;
/* input  */ logic          i_ch19_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch19_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch1_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch1_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch1_pld_sclk1_rowclk;
/* input  */ logic          i_ch1_pld_sclk2_rowclk;
/* input  */ logic          i_ch1_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch1_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch20_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch20_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch20_pld_sclk1_rowclk;
/* input  */ logic          i_ch20_pld_sclk2_rowclk;
/* input  */ logic          i_ch20_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch20_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch21_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch21_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch21_pld_sclk1_rowclk;
/* input  */ logic          i_ch21_pld_sclk2_rowclk;
/* input  */ logic          i_ch21_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch21_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch22_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch22_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch22_pld_sclk1_rowclk;
/* input  */ logic          i_ch22_pld_sclk2_rowclk;
/* input  */ logic          i_ch22_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch22_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch23_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch23_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch23_pld_sclk1_rowclk;
/* input  */ logic          i_ch23_pld_sclk2_rowclk;
/* input  */ logic          i_ch23_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch23_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch2_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch2_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch2_pld_sclk1_rowclk;
/* input  */ logic          i_ch2_pld_sclk2_rowclk;
/* input  */ logic          i_ch2_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch2_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch3_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch3_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch3_pld_sclk1_rowclk;
/* input  */ logic          i_ch3_pld_sclk2_rowclk;
/* input  */ logic          i_ch3_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch3_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch4_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch4_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch4_pld_sclk1_rowclk;
/* input  */ logic          i_ch4_pld_sclk2_rowclk;
/* input  */ logic          i_ch4_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch4_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch5_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch5_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch5_pld_sclk1_rowclk;
/* input  */ logic          i_ch5_pld_sclk2_rowclk;
/* input  */ logic          i_ch5_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch5_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch6_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch6_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch6_pld_sclk1_rowclk;
/* input  */ logic          i_ch6_pld_sclk2_rowclk;
/* input  */ logic          i_ch6_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch6_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch7_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch7_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch7_pld_sclk1_rowclk;
/* input  */ logic          i_ch7_pld_sclk2_rowclk;
/* input  */ logic          i_ch7_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch7_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch8_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch8_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch8_pld_sclk1_rowclk;
/* input  */ logic          i_ch8_pld_sclk2_rowclk;
/* input  */ logic          i_ch8_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch8_user_avmm2_clk_rowclk;
/* input  */ logic          i_ch9_pld_pma_coreclkin_rowclk;
/* input  */ logic          i_ch9_pld_rx_clk2_rowclk;
/* input  */ logic          i_ch9_pld_sclk1_rowclk;
/* input  */ logic          i_ch9_pld_sclk2_rowclk;
/* input  */ logic          i_ch9_user_avmm1_clk_rowclk;
/* input  */ logic          i_ch9_user_avmm2_clk_rowclk;
/* output */ logic [2:0]    o_ch0_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch0_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch0_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch0_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch0_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch10_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch10_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch10_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch10_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch10_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch11_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch11_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch11_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch11_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch11_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch12_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch12_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch12_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch12_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch12_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch13_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch13_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch13_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch13_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch13_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch14_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch14_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch14_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch14_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch14_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch15_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch15_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch15_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch15_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch16_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch16_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch16_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch16_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch16_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch17_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch17_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch17_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch17_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch17_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch18_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch18_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch18_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch18_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch18_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch19_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch19_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch19_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch19_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch19_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch1_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch1_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch1_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch1_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch1_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch20_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch20_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch20_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch20_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch20_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch21_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch21_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch21_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch21_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch21_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch22_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch22_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch22_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch22_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch22_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch23_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch23_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch23_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch23_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch23_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch2_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch2_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch2_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch2_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch2_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch3_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch3_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch3_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch3_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch3_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch4_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch4_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch4_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch4_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch4_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch5_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch5_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch5_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch5_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch5_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch6_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch6_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch6_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch6_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch6_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch7_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch7_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch7_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch7_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch7_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch8_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch8_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch8_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch8_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch8_pld_pcs_tx_clk_out2_dcm;
/* output */ logic [2:0]    o_ch9_pld_fpll_shared_direct_async_out_dcm;
/* output */ logic          o_ch9_pld_pcs_rx_clk_out1_dcm;
/* output */ logic          o_ch9_pld_pcs_rx_clk_out2_dcm;
/* output */ logic          o_ch9_pld_pcs_tx_clk_out1_dcm;
/* output */ logic          o_ch9_pld_pcs_tx_clk_out2_dcm;
/* input  */ logic [1:0]    i_ch0_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch0_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch10_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch10_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch11_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch11_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch12_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch12_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch13_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch13_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch14_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch14_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch15_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch15_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch16_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch16_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch17_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch17_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch18_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch18_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch19_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch19_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch1_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch1_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch20_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch20_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch21_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch21_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch22_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch22_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch23_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch23_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch2_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch2_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch3_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch3_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch4_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch4_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch5_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch5_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch6_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch6_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch7_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch7_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch8_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch8_pld_rx_clk2_dcm;
/* input  */ logic [1:0]    i_ch9_pld_fpll_shared_direct_async_in_dcm;
/* input  */ logic          i_ch9_pld_rx_clk2_dcm;
/* input  */ logic          i_aux_por_vccl_ovr;
/* input  */ logic [3:0]    i_id;
/* input  */ logic          i_jtag_hijack;
/* input  */ logic          i_jtag_tck;
/* input  */ logic          i_jtag_tdi;
/* output */ logic          io_jtag_tdo;
/* input  */ logic          i_jtag_tms;
/* input  */ logic          i_jtag_trst;
/* input  */ logic          i_sens_therm;
/* input  */ logic          i_strap_spare_in0;
/* input  */ logic          i_strap_spare_in1;
/* input  */ logic          i_edm_in;
/* output */ logic          o_edm_out;
/* output */ logic          o_sens_therm;
/* input  */ logic          s0_0_1__maib_rotate__maib_rotate;
/* input  */ logic          s0_187_1__aib_jtag_return__tdo;
/* input  */ logic          s1_0_1__aib_jtag_out__tck;
/* input  */ logic          s1_0_1__aib_jtag_out__tdi;
/* input  */ logic          s1_0_1__aib_jtag_out__tms;
/* input  */ logic          s1_0_1__dts_temptrip__temptrip;
/* input  */ logic          s2_0_1__aib_jtag_out__tck;
/* input  */ logic          s2_0_1__aib_jtag_out__tdi;
/* input  */ logic          s2_0_1__aib_jtag_out__tms;
/* input  */ logic          s2_187_1__aib_jtag_return__tdo;
/* input  */ logic [3:0]    s4_0_1__aib_cjtag_ctrl_id__cjtag_id;
/* input  */ logic          s5_187_1__cnoc__abort;
/* input  */ logic          s5_187_1__cnoc__clk;
/* input  */ logic          s5_187_1__cnoc__clk_n;
/* input  */ logic [32:0]   s5_187_1__cnoc__data;
/* input  */ logic          s5_187_1__cnoc__end_of_packet;
/* input  */ logic          s5_187_1__cnoc__nonsecure_interrupt;
/* input  */ logic          s5_187_1__cnoc__por;
/* input  */ logic          s5_187_1__cnoc__por_n;
/* input  */ logic          s5_187_1__cnoc__secure_interrupt;
/* input  */ logic          s5_187_1__cnoc__start_of_packet;
/* input  */ logic          s5_187_1__cnoc__sync;
/* input  */ logic          s5_187_1__cnoc__valid;
/* input  */ logic          s5_187_1__cnoc__warm_reset_n;
/* input  */ logic          s8_187_1__aib_jtag_return__tdo;
/* input  */ logic          s9_0_1__aib_jtag_out__tck;
/* input  */ logic          s9_0_1__aib_jtag_out__tdi;
/* input  */ logic          s9_0_1__aib_jtag_out__tms;
/* input  */ logic          s11_187_1__aib_jtag_out__tck;
/* input  */ logic          s11_187_1__aib_jtag_out__tdi;
/* input  */ logic          s11_187_1__aib_jtag_out__tms;
/* input  */ logic          s12_187_1__aib_jtag_out__tck;
/* input  */ logic          s12_187_1__aib_jtag_out__tdi;
/* input  */ logic          s12_187_1__aib_jtag_out__tms;
/* input  */ logic          s13_0_1__aib_jtag_return__tdo;
/* input  */ logic          s14_0_1__cjtag__tck;
/* input  */ logic          s14_0_1__cjtag__tdi;
/* input  */ logic          s14_0_1__cjtag__tms;
/* input  */ logic [3:0]    s14_187_1__aib_cjtag_ctrl_id__cjtag_id;
/* input  */ logic          s15_187_1__cjtag__tck;
/* input  */ logic          s15_187_1__cjtag__tdi;
/* input  */ logic          s15_187_1__cjtag__tms;
/* input  */ logic          s16_0_1__aib_jtag_return__tdo;
/* input  */ logic          s17_187_1__cjtag_return__tdo;
/* input  */ logic          s18_0_1__aib_jtag_return__tdo;
/* input  */ logic          s19_187_1__aib_jtag_out__tck;
/* input  */ logic          s19_187_1__aib_jtag_out__tdi;
/* input  */ logic          s19_187_1__aib_jtag_out__tms;
/* input  */ logic          s20_187_1__cnoc__abort;
/* input  */ logic          s20_187_1__cnoc__clk;
/* input  */ logic          s20_187_1__cnoc__clk_n;
/* input  */ logic [32:0]   s20_187_1__cnoc__data;
/* input  */ logic          s20_187_1__cnoc__end_of_packet;
/* input  */ logic          s20_187_1__cnoc__nonsecure_interrupt;
/* input  */ logic          s20_187_1__cnoc__por;
/* input  */ logic          s20_187_1__cnoc__por_n;
/* input  */ logic          s20_187_1__cnoc__secure_interrupt;
/* input  */ logic          s20_187_1__cnoc__start_of_packet;
/* input  */ logic          s20_187_1__cnoc__sync;
/* input  */ logic          s20_187_1__cnoc__valid;
/* input  */ logic          s20_187_1__cnoc__warm_reset_n;
/* input  */ logic          s21_0_1__cjtag_return__tdo;
/* input  */ logic          s23_0_1__cnoc__abort;
/* input  */ logic          s23_0_1__cnoc__clk;
/* input  */ logic          s23_0_1__cnoc__clk_n;
/* input  */ logic [32:0]   s23_0_1__cnoc__data;
/* input  */ logic          s23_0_1__cnoc__end_of_packet;
/* input  */ logic          s23_0_1__cnoc__nonsecure_interrupt;
/* input  */ logic          s23_0_1__cnoc__por;
/* input  */ logic          s23_0_1__cnoc__por_n;
/* input  */ logic          s23_0_1__cnoc__secure_interrupt;
/* input  */ logic          s23_0_1__cnoc__start_of_packet;
/* input  */ logic          s23_0_1__cnoc__sync;
/* input  */ logic          s23_0_1__cnoc__valid;
/* input  */ logic          s23_0_1__cnoc__warm_reset_n;
/* input  */ logic          s23_187_1__include_aib_jtag_segment__include_aib_jtag_segment;
/* input  */ logic          s25_187_1__include_aib_jtag_segment__include_aib_jtag_segment;
/* input  */ logic          s27_187_1__include_aib_jtag_segment__include_aib_jtag_segment;
/* input  */ logic          s28_187_1__dts_temptrip__temptrip;
/* input  */ logic          s30_0_1__dc_bsc_sdata__s_data;
/* input  */ logic          s30_187_1__dc_bsc_sdata__s_data;
/* input  */ logic          s32_187_1__sdm_mission_bus__clk;
/* input  */ logic [31:0]   s32_187_1__sdm_mission_bus__data;
/* input  */ logic          s32_187_1__sdm_mission_bus__valid;
/* input  */ logic [27:0]   s33_187_1__sdm_test_bus__data;
/* input  */ logic [15:0]   s34_0_1__sdm_testmode_ctrl__test_io_ctrl;
/* input  */ logic [15:0]   s37_0_1__test_return__data;
/* input  */ logic          s37_0_1__test_return__valid;
/* input  */ logic [4:0]    s38_0_1__scan_sdm_so__scan_out;
/* input  */ logic [3:0]    s39_0_1__cr_ctrl__muxsel_avst;
/* input  */ logic          s39_0_1__cr_ctrl__muxsel_test_cnoc;
/* input  */ logic          s124_0_1__include_aib_jtag_segment__include_aib_jtag_segment;
/* input  */ logic          s126_0_1__include_aib_jtag_segment__include_aib_jtag_segment;
/* input  */ logic          s128_0_1__include_aib_jtag_segment__include_aib_jtag_segment;
/* output */ logic [107:0]  o_s0_23_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_44_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_45_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_46_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_47_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_48_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_49_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_70_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_91_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_92_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_93_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_94_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_95_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_96_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_117_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_138_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_139_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_140_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_141_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_142_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_143_1__core_periphery__data_to_core;
/* output */ logic [107:0]  o_s0_164_1__core_periphery__data_to_core;
/* output */ logic [65:0]   s0_100_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_101_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_105_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_106_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_107_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_108_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_111_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_112_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_113_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_114_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_11_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_120_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_121_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_122_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_126_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_127_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_128_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_12_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_133_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_134_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_135_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_13_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_145_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_146_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_147_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_14_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_152_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_153_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_154_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_158_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_159_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_160_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_167_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_168_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_169_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_173_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_174_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_175_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_17_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_180_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_181_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_182_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_183_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_18_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_19_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_20_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_26_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_27_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_28_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_29_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_32_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_33_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_34_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_35_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_39_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_40_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_41_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_42_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_4_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_51_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_52_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_53_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_54_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_58_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_59_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_5_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_60_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_61_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_64_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_65_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_66_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_67_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_6_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_73_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_74_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_75_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_76_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_79_1__core_periphery__data_to_core_unused;
/* output */ logic [85:0]   s0_7_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_80_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_81_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_82_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_86_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_87_1__core_periphery__data_to_core_unused;
/* output */ logic [65:0]   s0_88_1__core_periphery__data_to_core_unused;
/* output */ logic [95:0]   s0_89_1__core_periphery__data_to_core_unused;
/* output */ logic [39:0]   s0_98_1__core_periphery__data_to_core_unused;
/* output */ logic [53:0]   s0_99_1__core_periphery__data_to_core_unused;
/* input  */ logic [15:0]   i_s0_3_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_8_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_9_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_10_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_15_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_16_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_21_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_22_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_23_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_24_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_25_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_30_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_31_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_36_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_37_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_38_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_43_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_44_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_45_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_46_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_47_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_48_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_49_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_50_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_55_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_56_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_57_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_62_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_63_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_68_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_69_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_70_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_71_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_72_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_77_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_78_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_83_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_84_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_85_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_90_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_91_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_92_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_93_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_94_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_95_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_96_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_97_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_102_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_103_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_104_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_109_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_110_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_115_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_116_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_117_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_118_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_119_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_124_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_125_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_130_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_131_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_132_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_137_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_138_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_139_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_140_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_141_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_142_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_143_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_144_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_149_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_150_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_151_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_156_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_157_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_162_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_163_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_164_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_165_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_166_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_171_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_172_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_177_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_178_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_179_1__core_periphery__clock_from_core;
/* input  */ logic [15:0]   i_s0_184_1__core_periphery__clock_from_core;
/* input  */ logic [95:0]   i_s0_3_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_9_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_10_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_15_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_16_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_21_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_22_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_23_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_24_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_25_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_30_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_31_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_36_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_37_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_38_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_43_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_44_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_45_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_46_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_47_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_48_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_49_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_50_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_55_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_56_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_57_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_62_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_63_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_68_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_69_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_70_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_71_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_72_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_77_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_78_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_83_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_84_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_90_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_91_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_92_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_93_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_94_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_95_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_96_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_97_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_102_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_103_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_104_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_109_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_110_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_115_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_116_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_117_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_118_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_119_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_124_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_125_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_130_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_131_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_132_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_137_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_138_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_139_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_140_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_141_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_142_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_143_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_144_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_149_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_150_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_151_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_156_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_157_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_162_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_163_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_164_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_165_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_166_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_171_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_172_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_177_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_178_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_179_1__core_periphery__data_from_core;
/* input  */ logic [95:0]   i_s0_184_1__core_periphery__data_from_core;
/* input  */ logic [13:0]   s0_100_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_100_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_101_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_101_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_105_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_105_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_106_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_106_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_107_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_107_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_108_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_108_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_111_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_111_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_112_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_112_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_113_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_113_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_114_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_114_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_11_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_11_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_120_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_120_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_121_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_121_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_122_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_122_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_123_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_123_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_126_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_126_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_127_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_127_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_128_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_128_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_129_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_129_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_12_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_12_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_133_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_133_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_134_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_134_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_135_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_135_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_136_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_136_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_13_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_13_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_145_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_145_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_146_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_146_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_147_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_147_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_148_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_148_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_14_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_14_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_152_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_152_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_153_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_153_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_154_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_154_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_155_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_155_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_158_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_158_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_159_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_159_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_160_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_160_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_161_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_161_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_167_1__core_periphery__clock_from_core_unused;
/* input  */ logic [72:0]   s0_167_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_168_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_168_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_169_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_169_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_170_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_170_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_173_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_173_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_174_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_174_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_175_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_175_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_176_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_176_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_17_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_17_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_180_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_180_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_181_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_181_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_182_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_182_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_183_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_183_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_18_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_18_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_19_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_19_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_20_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_20_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_26_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_26_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_27_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_27_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_28_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_28_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_29_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_29_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_32_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_32_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_33_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_33_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_34_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_34_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_35_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_35_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_39_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_39_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_40_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_40_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_41_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_41_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_42_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_42_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_4_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_4_1__core_periphery__data_from_core_unused; //;
/* input  */ logic [14:0]   s0_51_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_51_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_52_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_52_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_53_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_53_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_54_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_54_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_58_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_58_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_59_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_59_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_5_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_5_1__core_periphery__data_from_core_unused; //;
/* input  */ logic [13:0]   s0_60_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_60_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_61_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_61_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_64_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_64_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_65_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_65_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_66_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_66_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_67_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_67_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_6_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_6_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_73_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_73_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_74_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_74_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_75_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_75_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_76_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_76_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_79_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_79_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_7_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_7_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_80_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_80_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_81_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_81_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_82_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_82_1__core_periphery__data_from_core_unused;
/* input  */ logic [93:0]   s0_85_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_86_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_86_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_87_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_87_1__core_periphery__data_from_core_unused;
/* input  */ logic [13:0]   s0_88_1__core_periphery__clock_from_core_unused;
/* input  */ logic [21:0]   s0_88_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_89_1__core_periphery__clock_from_core_unused;
/* input  */ logic [66:0]   s0_89_1__core_periphery__data_from_core_unused;
/* input  */ logic [64:0]   s0_8_1__core_periphery__data_from_core_unused;
/* input  */ logic [14:0]   s0_98_1__core_periphery__clock_from_core_unused;
/* input  */ logic [59:0]   s0_98_1__core_periphery__data_from_core_unused;
/* input  */ logic [9:0]    s0_99_1__core_periphery__clock_from_core_unused;
/* input  */ logic [34:0]   s0_99_1__core_periphery__data_from_core_unused;
/* input  */ logic          vcc_dts_ref;
/* input  */ logic          vcce_pll_ref;

 // Assign Ports 
 // AVST Ports 
 assign  p0_rx_st_par_err_o = 1'b0;
 assign  p0_tx_st_par_err_o = 1'b0;
/* output */ assign p0_ptm_clk_updated_o                                    = o_ptm_clk_updated;
/* output */ assign p0_ptm_context_valid_o                                  = o_ptm_context_valid;
/* output */ assign p0_ptm_local_clock_o                                    = o_ptm_local_clock;
/* input  */ assign i_ptm_manual_update                                  = p0_ptm_manual_update_i;
/* output */ assign p0_rx_st0_dvalid_o                                   = rx_st0_dvalid;
/* output */ assign p0_rx_st1_dvalid_o                                   = rx_st1_dvalid;
/* output */ assign p0_rx_st2_dvalid_o                                   = rx_st2_dvalid;
/* output */ assign p0_rx_st3_dvalid_o                                   = rx_st3_dvalid;
/* output */ assign p0_rx_st0_sop_o                                      = rx_st0_sop;
/* output */ assign p0_rx_st1_sop_o                                      = rx_st1_sop;
/* output */ assign p0_rx_st2_sop_o                                      = rx_st2_sop;
/* output */ assign p0_rx_st3_sop_o                                      = rx_st3_sop;
/* output */ assign p0_rx_st0_eop_o                                      = rx_st0_eop;
/* output */ assign p0_rx_st1_eop_o                                      = rx_st1_eop;
/* output */ assign p0_rx_st2_eop_o                                      = rx_st2_eop;
/* output */ assign p0_rx_st3_eop_o                                      = rx_st3_eop;
/* output */ assign p0_rx_st0_passthrough_o                              = rx_st0_passthrough;
/* output */ assign p0_rx_st1_passthrough_o                              = rx_st1_passthrough;
/* output */ assign p0_rx_st2_passthrough_o                              = rx_st2_passthrough;
/* output */ assign p0_rx_st3_passthrough_o                              = rx_st3_passthrough;
/* output */ assign p0_rx_st0_data_o                                     = rx_st0_data;
/* output */ assign p0_rx_st1_data_o                                     = rx_st1_data;
/* output */ assign p0_rx_st2_data_o                                     = rx_st2_data;
/* output */ assign p0_rx_st3_data_o                                     = rx_st3_data;
/* output */ assign p0_rx_st0_data_par_o                                 = rx_st0_data_parity;
/* output */ assign p0_rx_st1_data_par_o                                 = rx_st1_data_parity;
/* output */ assign p0_rx_st2_data_par_o                                 = rx_st2_data_parity;
/* output */ assign p0_rx_st3_data_par_o                                 = rx_st3_data_parity;
/* output */ assign p0_rx_st0_hdr_o                                      = rx_st0_hdr;
/* output */ assign p0_rx_st1_hdr_o                                      = rx_st1_hdr;
/* output */ assign p0_rx_st2_hdr_o                                      = rx_st2_hdr;
/* output */ assign p0_rx_st3_hdr_o                                      = rx_st3_hdr;
/* output */ assign p0_rx_st0_hdr_par_o                                  = rx_st0_hdr_parity;
/* output */ assign p0_rx_st1_hdr_par_o                                  = rx_st1_hdr_parity;
/* output */ assign p0_rx_st2_hdr_par_o                                  = rx_st2_hdr_parity;
/* output */ assign p0_rx_st3_hdr_par_o                                  = rx_st3_hdr_parity;
/* output */ assign p0_rx_st0_hvalid_o                                   = rx_st0_hvalid;
/* output */ assign p0_rx_st1_hvalid_o                                   = rx_st1_hvalid;
/* output */ assign p0_rx_st2_hvalid_o                                   = rx_st2_hvalid;
/* output */ assign p0_rx_st3_hvalid_o                                   = rx_st3_hvalid;
/* output */ assign p0_rx_st0_prefix_o                                   = rx_st0_prefix;
/* output */ assign p0_rx_st1_prefix_o                                   = rx_st1_prefix;
/* output */ assign p0_rx_st2_prefix_o                                   = rx_st2_prefix;
/* output */ assign p0_rx_st3_prefix_o                                   = rx_st3_prefix;
/* output */ assign p0_rx_st0_prefix_par_o                               = rx_st0_prefix_parity;
/* output */ assign p0_rx_st1_prefix_par_o                               = rx_st1_prefix_parity;
/* output */ assign p0_rx_st2_prefix_par_o                               = rx_st2_prefix_parity;
/* output */ assign p0_rx_st3_prefix_par_o                               = rx_st3_prefix_parity;
/* output */ assign p0_rx_st0_rssai_prefix_o                             = rx_st0_rssai_prefix;
/* output */ assign p0_rx_st1_rssai_prefix_o                             = rx_st1_rssai_prefix;
/* output */ assign p0_rx_st2_rssai_prefix_o                             = rx_st2_rssai_prefix;
/* output */ assign p0_rx_st3_rssai_prefix_o                             = rx_st3_rssai_prefix;
/* output */ assign p0_rx_st0_rssai_prefix_par_o                         = rx_st0_rssai_prefix_parity;
/* output */ assign p0_rx_st1_rssai_prefix_par_o                         = rx_st1_rssai_prefix_parity;
/* output */ assign p0_rx_st2_rssai_prefix_par_o                         = rx_st2_rssai_prefix_parity;
/* output */ assign p0_rx_st3_rssai_prefix_par_o                         = rx_st3_rssai_prefix_parity;
/* output */ assign p0_rx_st0_pvalid_o                                   = rx_st0_pvalid;
/* output */ assign p0_rx_st1_pvalid_o                                   = rx_st1_pvalid;
/* output */ assign p0_rx_st2_pvalid_o                                   = rx_st2_pvalid;
/* output */ assign p0_rx_st3_pvalid_o                                   = rx_st3_pvalid;
/* output */ assign p0_rx_st0_bar_o                                      = rx_st0_bar;
/* output */ assign p0_rx_st1_bar_o                                      = rx_st1_bar;
/* output */ assign p0_rx_st2_bar_o                                      = rx_st2_bar;
/* output */ assign p0_rx_st3_bar_o                                      = rx_st3_bar;
/* output */ assign p0_rx_st0_vfactive_o                                 = rx_st0_vfactive;
/* output */ assign p0_rx_st1_vfactive_o                                 = rx_st1_vfactive;
/* output */ assign p0_rx_st2_vfactive_o                                 = rx_st2_vfactive;
/* output */ assign p0_rx_st3_vfactive_o                                 = rx_st3_vfactive;
/* output */ assign p0_rx_st0_vfnum_o                                    = rx_st0_vfnum;
/* output */ assign p0_rx_st1_vfnum_o                                    = rx_st1_vfnum;
/* output */ assign p0_rx_st2_vfnum_o                                    = rx_st2_vfnum;
/* output */ assign p0_rx_st3_vfnum_o                                    = rx_st3_vfnum;
/* output */ assign p0_rx_st0_pfnum_o                                    = rx_st0_pfnum;
/* output */ assign p0_rx_st1_pfnum_o                                    = rx_st1_pfnum;
/* output */ assign p0_rx_st2_pfnum_o                                    = rx_st2_pfnum;
/* output */ assign p0_rx_st3_pfnum_o                                    = rx_st3_pfnum;
/* output */ assign p0_rx_st0_chnum_o                                    = rx_st0_chnum;
/* output */ assign p0_rx_st1_chnum_o                                    = rx_st1_chnum;
/* output */ assign p0_rx_st2_chnum_o                                    = rx_st2_chnum;
/* output */ assign p0_rx_st3_chnum_o                                    = rx_st3_chnum;
/* output */ assign p0_rx_st0_misc_par_o                                 = rx_st0_misc_parity;
/* output */ assign p0_rx_st1_misc_par_o                                 = rx_st1_misc_parity;
/* output */ assign p0_rx_st2_misc_par_o                                 = rx_st2_misc_parity;
/* output */ assign p0_rx_st3_misc_par_o                                 = rx_st3_misc_parity;
/* output */ assign p0_rx_st0_empty_o                                    = rx_st0_empty;
/* output */ assign p0_rx_st1_empty_o                                    = rx_st1_empty;
/* output */ assign p0_rx_st2_empty_o                                    = rx_st2_empty;
/* output */ assign p0_rx_st3_empty_o                                    = rx_st3_empty;
/* input  */ assign rx_st_Hcrdt_update                                   = p0_rx_st_hcrd_update_i;
/* input  */ assign rx_st_Hcrdt_ch                                       = p0_rx_st_hcrd_ch_i;
/* input  */ assign rx_st_Hcrdt_update_cnt                               = p0_rx_st_hcrd_update_cnt_i;
/* input  */ assign rx_st_Hcrdt_init                                     = p0_rx_st_hcrd_init_i;
/* output */ assign p0_rx_st_hcrd_init_ack_o                             = rx_st_Hcrdt_init_ack;
/* input  */ assign rx_st_Dcrdt_update                                   = p0_rx_st_dcrd_update_i;
/* input  */ assign rx_st_Dcrdt_ch                                       = p0_rx_st_dcrd_ch_i;
/* input  */ assign rx_st_Dcrdt_update_cnt                               = p0_rx_st_dcrd_update_cnt_i;
/* input  */ assign rx_st_Dcrdt_init                                     = p0_rx_st_dcrd_init_i;
/* output */ assign p0_rx_st_dcrd_init_ack_o                             = rx_st_Dcrdt_init_ack;
/* output */ assign p0_tx_st_ready_o                                     = tx_st_ready;
/* input  */ assign tx_st0_dvalid                                        = p0_tx_st0_dvalid_i;
/* input  */ assign tx_st1_dvalid                                        = p0_tx_st1_dvalid_i;
/* input  */ assign tx_st2_dvalid                                        = p0_tx_st2_dvalid_i;
/* input  */ assign tx_st3_dvalid                                        = p0_tx_st3_dvalid_i;
/* input  */ assign tx_st0_sop                                           = p0_tx_st0_sop_i;
/* input  */ assign tx_st1_sop                                           = p0_tx_st1_sop_i;
/* input  */ assign tx_st2_sop                                           = p0_tx_st2_sop_i;
/* input  */ assign tx_st3_sop                                           = p0_tx_st3_sop_i;
/* input  */ assign tx_st0_eop                                           = p0_tx_st0_eop_i;
/* input  */ assign tx_st1_eop                                           = p0_tx_st1_eop_i;
/* input  */ assign tx_st2_eop                                           = p0_tx_st2_eop_i;
/* input  */ assign tx_st3_eop                                           = p0_tx_st3_eop_i;
/* input  */ assign tx_st0_passthrough                                   = p0_tx_st0_passthrough_i;
/* input  */ assign tx_st1_passthrough                                   = p0_tx_st1_passthrough_i;
/* input  */ assign tx_st2_passthrough                                   = p0_tx_st2_passthrough_i;
/* input  */ assign tx_st3_passthrough                                   = p0_tx_st3_passthrough_i;
/* input  */ assign tx_st0_data                                          = p0_tx_st0_data_i;
/* input  */ assign tx_st1_data                                          = p0_tx_st1_data_i;
/* input  */ assign tx_st2_data                                          = p0_tx_st2_data_i;
/* input  */ assign tx_st3_data                                          = p0_tx_st3_data_i;
/* input  */ assign tx_st0_data_parity                                   = p0_tx_st0_data_par_i;
/* input  */ assign tx_st1_data_parity                                   = p0_tx_st1_data_par_i;
/* input  */ assign tx_st2_data_parity                                   = p0_tx_st2_data_par_i;
/* input  */ assign tx_st3_data_parity                                   = p0_tx_st3_data_par_i;
/* input  */ assign tx_st0_hdr                                           = p0_tx_st0_hdr_i;
/* input  */ assign tx_st1_hdr                                           = p0_tx_st1_hdr_i;
/* input  */ assign tx_st2_hdr                                           = p0_tx_st2_hdr_i;
/* input  */ assign tx_st3_hdr                                           = p0_tx_st3_hdr_i;
/* input  */ assign tx_st0_hdr_parity                                    = p0_tx_st0_hdr_par_i;
/* input  */ assign tx_st1_hdr_parity                                    = p0_tx_st1_hdr_par_i;
/* input  */ assign tx_st2_hdr_parity                                    = p0_tx_st2_hdr_par_i;
/* input  */ assign tx_st3_hdr_parity                                    = p0_tx_st3_hdr_par_i;
/* input  */ assign tx_st0_hvalid                                        = p0_tx_st0_hvalid_i;
/* input  */ assign tx_st1_hvalid                                        = p0_tx_st1_hvalid_i;
/* input  */ assign tx_st2_hvalid                                        = p0_tx_st2_hvalid_i;
/* input  */ assign tx_st3_hvalid                                        = p0_tx_st3_hvalid_i;
/* input  */ assign tx_st0_prefix                                        = p0_tx_st0_prefix_i;
/* input  */ assign tx_st1_prefix                                        = p0_tx_st1_prefix_i;
/* input  */ assign tx_st2_prefix                                        = p0_tx_st2_prefix_i;
/* input  */ assign tx_st3_prefix                                        = p0_tx_st3_prefix_i;
/* input  */ assign tx_st0_prefix_parity                                 = p0_tx_st0_prefix_par_i;
/* input  */ assign tx_st1_prefix_parity                                 = p0_tx_st1_prefix_par_i;
/* input  */ assign tx_st2_prefix_parity                                 = p0_tx_st2_prefix_par_i;
/* input  */ assign tx_st3_prefix_parity                                 = p0_tx_st3_prefix_par_i;
/* input  */ assign tx_st0_rssai_prefix                                  = p0_tx_st0_rssai_prefix_i;
/* input  */ assign tx_st1_rssai_prefix                                  = p0_tx_st1_rssai_prefix_i;
/* input  */ assign tx_st2_rssai_prefix                                  = p0_tx_st2_rssai_prefix_i;
/* input  */ assign tx_st3_rssai_prefix                                  = p0_tx_st3_rssai_prefix_i;
/* input  */ assign tx_st0_rssai_prefix_parity                           = p0_tx_st0_rssai_prefix_par_i;
/* input  */ assign tx_st1_rssai_prefix_parity                           = p0_tx_st1_rssai_prefix_par_i;
/* input  */ assign tx_st2_rssai_prefix_parity                           = p0_tx_st2_rssai_prefix_par_i;
/* input  */ assign tx_st3_rssai_prefix_parity                           = p0_tx_st3_rssai_prefix_par_i;
/* input  */ assign tx_st0_pvalid                                        = p0_tx_st0_pvalid_i;
/* input  */ assign tx_st1_pvalid                                        = p0_tx_st1_pvalid_i;
/* input  */ assign tx_st2_pvalid                                        = p0_tx_st2_pvalid_i;
/* input  */ assign tx_st3_pvalid                                        = p0_tx_st3_pvalid_i;
/* input  */ assign tx_st0_empty                                         = p0_tx_st0_empty_i;
/* input  */ assign tx_st1_empty                                         = p0_tx_st1_empty_i;
/* input  */ assign tx_st2_empty                                         = p0_tx_st2_empty_i;
/* input  */ assign tx_st3_empty                                         = p0_tx_st3_empty_i;
/* output */ assign p0_tx_st_hcrd_update_o                               = tx_st_Hcrdt_update;
/* output */ assign p0_tx_st_hcrd_ch_o                                   = tx_st_Hcrdt_vc;
/* output */ assign p0_tx_st_hcrd_update_cnt_o                           = tx_st_Hcrdt_update_cnt;
/* output */ assign p0_tx_st_hcrd_init_o                                 = tx_st_Hcrdt_init;
/* input  */ assign tx_st_Hcrdt_init_ack                                 = p0_tx_st_hcrd_init_ack_i;
/* output */ assign p0_tx_st_dcrd_update_o                               = tx_st_Dcrdt_update;
/* output */ assign p0_tx_st_dcrd_ch_o                                   = tx_st_Dcrdt_vc;
/* output */ assign p0_tx_st_dcrd_update_cnt_o                           = tx_st_Dcrdt_update_cnt;
/* output */ assign p0_tx_st_dcrd_init_o                                 = tx_st_Dcrdt_init;
/* input  */ assign tx_st_Dcrdt_init_ack                                 = p0_tx_st_dcrd_init_ack_i;
/* input  */ assign i_ch0_pld_sclk1_rowclk                               = o_ch0_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch0_pld_sclk2_rowclk                               = o_ch0_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch10_pld_sclk1_rowclk                              = o_ch10_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch10_pld_sclk2_rowclk                              = o_ch10_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch11_pld_sclk1_rowclk                              = o_ch11_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch11_pld_sclk2_rowclk                              = o_ch11_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch12_pld_sclk1_rowclk                              = o_ch12_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch12_pld_sclk2_rowclk                              = o_ch12_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch13_pld_sclk1_rowclk                              = o_ch13_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch13_pld_sclk2_rowclk                              = o_ch13_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch14_pld_sclk1_rowclk                              = o_ch14_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch14_pld_sclk2_rowclk                              = o_ch14_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch15_pld_sclk1_rowclk                              = o_ch15_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch15_pld_sclk2_rowclk                              = o_ch15_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch16_pld_sclk1_rowclk                              = o_ch16_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch16_pld_sclk2_rowclk                              = o_ch16_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch17_pld_sclk1_rowclk                              = o_ch17_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch17_pld_sclk2_rowclk                              = o_ch17_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch18_pld_sclk1_rowclk                              = o_ch18_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch18_pld_sclk2_rowclk                              = o_ch18_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch19_pld_sclk1_rowclk                              = o_ch19_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch19_pld_sclk2_rowclk                              = o_ch19_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch1_pld_sclk1_rowclk                               = o_ch1_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch1_pld_sclk2_rowclk                               = o_ch1_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch20_pld_sclk1_rowclk                              = o_ch20_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch20_pld_sclk2_rowclk                              = o_ch20_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch21_pld_sclk1_rowclk                              = o_ch21_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch21_pld_sclk2_rowclk                              = o_ch21_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch22_pld_sclk1_rowclk                              = o_ch22_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch22_pld_sclk2_rowclk                              = o_ch22_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch23_pld_sclk1_rowclk                              = o_ch23_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch23_pld_sclk2_rowclk                              = o_ch23_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch2_pld_sclk1_rowclk                               = o_ch2_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch2_pld_sclk2_rowclk                               = o_ch2_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch3_pld_sclk1_rowclk                               = o_ch3_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch3_pld_sclk2_rowclk                               = o_ch3_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch4_pld_sclk1_rowclk                               = o_ch4_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch4_pld_sclk2_rowclk                               = o_ch4_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch5_pld_sclk1_rowclk                               = o_ch5_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch5_pld_sclk2_rowclk                               = o_ch5_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch6_pld_sclk1_rowclk                               = o_ch6_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch6_pld_sclk2_rowclk                               = o_ch6_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch7_pld_sclk1_rowclk                               = o_ch7_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch7_pld_sclk2_rowclk                               = o_ch7_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch8_pld_sclk1_rowclk                               = o_ch8_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch8_pld_sclk2_rowclk                               = o_ch8_pld_pcs_tx_clk_out2_dcm;
/* input  */ assign i_ch9_pld_sclk1_rowclk                               = o_ch9_pld_pcs_tx_clk_out1_dcm;
/* input  */ assign i_ch9_pld_sclk2_rowclk                               = o_ch9_pld_pcs_tx_clk_out2_dcm;
   // Reconfig Interface
/* input  */ assign i_jtag_hijack                                      = 1'b0;
/* input  */ assign s0_5_1__core_periphery__data_from_core_unused[33]  =  1'b0;  //adapter_scan_rst_n
/* input  */ assign s0_5_1__core_periphery__data_from_core_unused[13]  =  1'b1;  //adapter_scan_mode_n
/* input  */ assign s0_5_1__core_periphery__data_from_core_unused[14]  =  1'b1;  //adapter_scan_shift_n
/* input  */ assign s0_5_1__core_periphery__data_from_core_unused[24]  =  1'b1;  //adapter_clk_sel_n
/* input  */ assign s0_5_1__core_periphery__data_from_core_unused[25]  =  1'b0;  //adapter_occ_enable
/* input  */ assign s0_5_1__core_periphery__data_from_core_unused[26]  =  1'b1;  //adapter_global_pipe_se
/* input  */ assign s0_4_1__core_periphery__data_from_core_unused[37]  =  1'b1;  //hvqk_mode_in
/* input  */ assign cxl_pll_locked_i                                   =  1'b1;
//SJ
wire i_clk0;
wire i_clk1;
assign i_clk                                              =  i_clk0;
//// tennm_sdm_oscillator #(
////// Parameters
//// .sim_clkout_period_ps(5000)
////) u_src_clk(
////       // Input Ports
////       // Output Ports
////       .clkout(i_clk0 ),
////       .clkout1(i_clk1)
////);

altera_s10_configuration_clock s10_configuration_clock_0 (
             .clkout (i_clk0)  //  output,  width = 1, clkout.clk
);



/* input  */ assign i_rst_n                                            =  1'b1;
/* input  */ assign i_rx_dsk_clear                                     =  1'b0;
/* input  */ assign i_tx_dsk_clear                                     =  1'b0;
/* input  */ assign i_ch0_async_direct_pld2aib[0]                      =  1'b1;  // assign pld_superrst_n = i_ch0_async_direct_pld2aib[0];
/* input  */ assign i_ch1_async_direct_pld2aib[0]                      =  1'b1;  // assign pld_fullrst_n = i_ch1_async_direct_pld2aib[0];
/* input  */ assign i_ch0_async_direct_pld2aib[5]                      =  1'b1;  // assign pld_cxl_ipxrst_n = i_ch0_async_direct_pld2aib[5];
/* input  */ assign i_ch1_async_direct_pld2aib[5]                      =  1'b1;  // assign pld_cxl_ipxprst_n = i_ch1_async_direct_pld2aib[5];
/* input  */ assign p0_reset_status_n                                  =  cxl_reset_status_n; // PORT_NAME_CHANGE_REMOVED

/* input  */ assign s0_5_1__core_periphery__data_from_core_unused[27]  =  1'b1;  //adapter_occ_scan_in
/* input  */ assign s0_52_1__core_periphery__data_from_core_unused[27] =  1'b1;  //adapter_occ_scan_in
/* input  */ assign s0_99_1__core_periphery__data_from_core_unused[27] =  1'b1;  //adapter_occ_scan_in
/* input  */ assign s0_146_1__core_periphery__data_from_core_unused[27]=  1'b1;  //adapter_occ_scan_in

  localparam  MAX_CONVERSION_SIZE = 128;
  localparam  MAX_STRING_CHARS    = 64;

  function [MAX_CONVERSION_SIZE-1:0] str_2_bin;
     input [MAX_STRING_CHARS*8-1:0] instring;

     integer this_char;
     integer i;
     begin
        this_char = 0;
        i = 0;
        // Initialize accumulator
        str_2_bin = {MAX_CONVERSION_SIZE{1'b0}};
        for(i=MAX_STRING_CHARS-1;i>=0;i=i-1) begin
           this_char = instring[i*8+:8];
           // Add value of this digit
           if(this_char >= 48 && this_char <= 57)
              str_2_bin = (str_2_bin * 10) + (this_char - 48);
        end
     end
  endfunction

// user_avmm_interface user_avmm_if();
//
///* input  */ assign user_avmm_if.app_user_avmm_clk                    =  reconfig_clk;
///* input  */ assign user_avmm_if.app_user_avmm_address                =  reconfig_address;
///* input  */ assign user_avmm_if.app_user_avmm_read                   =  reconfig_read;
///* input  */ assign user_avmm_if.app_user_avmm_write                  =  reconfig_write;
///* input  */ assign user_avmm_if.app_user_avmm_writedata              =  reconfig_writedata;
///* output */ assign reconfig_readdata                                 =  user_avmm_if.app_user_avmm_readdata;
///* output */ assign reconfig_readdatavalid                            =  user_avmm_if.app_user_avmm_readdatavalid;
///* output */ assign reconfig_waitrequest                              =  user_avmm_if.app_user_avmm_waitrequest;
///* output */ assign reconfig_reserved_out                             =  5'h00; //Need to be updated
//
//             assign i_user_avmm2_clk_rowclk                           =  user_avmm_if.user_avmm_clk;
//             assign i_user_avmm_reg_addr                              =  user_avmm_if.user_avmm_address;
//             assign i_user_avmm_read                                  =  user_avmm_if.user_avmm_read;
//             assign i_user_avmm_write                                 =  user_avmm_if.user_avmm_write;
//             assign i_user_avmm_writedata                             =  user_avmm_if.user_avmm_writedata;
//             assign user_avmm_if.user_avmm_readdata                   =  o_user_avmm_readdata;
//             assign user_avmm_if.user_avmm_readdatavalid              =  o_user_avmm_readdatavalid;
//             assign user_avmm_if.user_avmm_writedone                  =  o_user_avmm_writedone;
// 
// rnr_cxl_user_avmm_adapter user_avmm(
//                  .rst_n(p0_reset_status_n),
//                  .avmm_user_ports(user_avmm_if.app_user_avmm_ports),  // user interface
//                  .avmm_maib_ports(user_avmm_if.pld_user_avmm_ports)   // maib interface 
//               );

//SJ  assign user_avmm_if.app_phyq_sel[4:0] = '0; 
//assign p0_pld_warm_rst_rdy_i = '0; 
assign p1_pld_warm_rst_rdy_i = '0; 
assign p2_pld_warm_rst_rdy_i = '0; 
assign p3_pld_warm_rst_rdy_i = '0; 
assign p0_app_rst_n = '0; 
assign p1_app_rst_n = '0; 
assign p2_app_rst_n = '0; 
assign p3_app_rst_n = '0; 
assign cxl_app_rst_n = '0; 
assign i_ial_ch19_ext_fsr[3:0] = '0; 
assign i_ial_ch19_ext_ssr[39:0] = '0; 
assign i_ial_ch19_fsr[2:0] = '0; 
assign i_ial_ch19_ssr[60:0] = '0; 
assign i_ial_ch20_ext_fsr[3:0] = '0; 
assign i_ial_ch20_ext_ssr[39:0] = '0; 
assign i_ial_ch20_fsr[2:0] = '0; 
assign i_ial_ch20_ssr[60:0] = '0; 
assign i_ial_ch21_ext_fsr[3:0] = '0; 
assign i_ial_ch21_ext_ssr[39:0] = '0; 
assign i_ial_ch21_fsr[2:0] = '0; 
assign i_ial_ch21_ssr[60:0] = '0; 
assign i_ial_ch22_async_direct[7:0] = '0; 
assign i_ial_ch22_ext_fsr[3:0] = '0; 
assign i_ial_ch22_ext_ssr[39:0] = '0; 
assign i_ial_ch22_fsr[2:0] = '0; 
assign i_ial_ch22_ssr[60:0] = '0; 
assign i_ial_ch23_async_direct[7:0] = '0; 
assign i_ial_ch23_ext_fsr[3:0] = '0; 
assign i_ial_ch23_ext_ssr[39:0] = '0; 
assign i_ial_ch23_fsr[2:0] = '0; 
assign i_ial_ch23_ssr[60:0] = '0; 
assign i_ch0_async_direct_pld2aib[7:6] = '0; 
assign i_ch0_async_direct_pld2aib[4:1] = '0; 
assign i_ch1_async_direct_pld2aib[7:6] = '0; 
assign i_ch1_async_direct_pld2aib[4:1] = '0; 
assign i_ch2_async_direct_pld2aib[7:0] = '0; 
assign i_ch3_async_direct_pld2aib[7:0] = '0; 
assign i_ch4_async_direct_pld2aib[7:0] = '0; 
assign i_ch5_async_direct_pld2aib[7:0] = '0; 
assign i_ch6_async_direct_pld2aib[7:0] = '0; 
assign i_ch7_async_direct_pld2aib[7:0] = '0; 
assign i_ch11_fsr_pld2aib[6:0] = '0; 
assign i_ch9_fsr_pld2aib[6:0] = '0; 
assign ial_phy_tx_fsr_0__tx_chnl_fsr[2:0] = '0; 
assign ial_phy_tx_fsr_0__tx_ext_fsr[3:0] = '0; 
assign ial_phy_tx_fsr_1__tx_chnl_fsr[2:0] = '0; 
assign ial_phy_tx_fsr_1__tx_ext_fsr[3:0] = '0; 
assign ial_phy_tx_fsr_2__tx_chnl_fsr[2:0] = '0; 
assign ial_phy_tx_fsr_2__tx_ext_fsr[3:0] = '0; 
assign ial_phy_tx_fsr_3__tx_chnl_fsr[2:0] = '0; 
assign ial_phy_tx_fsr_3__tx_ext_fsr[3:0] = '0; 
assign ial_phy_tx_fsr_4__tx_chnl_fsr[2:0] = '0; 
assign ial_phy_tx_fsr_4__tx_ext_fsr[3:0] = '0; 
assign ial_phy_tx_fsr_5__tx_chnl_fsr[2:0] = '0; 
assign ial_phy_tx_fsr_5__tx_ext_fsr[3:0] = '0; 
assign pcie_phy_tx_fsr_10__tx_chnl_fsr[2:0] = '0; 
assign pcie_phy_tx_fsr_10__tx_ext_fsr[3:0] = '0; 
assign pcie_phy_tx_fsr_11__tx_chnl_fsr[2:0] = '0; 
assign pcie_phy_tx_fsr_11__tx_ext_fsr[3:0] = '0; 
assign i_ch0_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch10_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch11_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch12_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch13_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch14_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch15_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch16_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch17_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch18_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch19_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch1_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch20_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch21_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch22_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch23_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch2_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch3_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch4_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch5_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch6_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch7_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch8_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch9_pld_pma_coreclkin_rowclk = 1'b1; 
assign i_ch0_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch0_pld_rx_clk2_dcm = '0; 
assign i_ch10_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch10_pld_rx_clk2_dcm = '0; 
assign i_ch11_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch11_pld_rx_clk2_dcm = '0; 
assign i_ch12_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch12_pld_rx_clk2_dcm = '0; 
assign i_ch13_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch13_pld_rx_clk2_dcm = '0; 
assign i_ch14_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch14_pld_rx_clk2_dcm = '0; 
assign i_ch15_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch15_pld_rx_clk2_dcm = '0; 
assign i_ch16_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch16_pld_rx_clk2_dcm = '0; 
assign i_ch17_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch17_pld_rx_clk2_dcm = '0; 
assign i_ch18_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch18_pld_rx_clk2_dcm = '0; 
assign i_ch19_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch19_pld_rx_clk2_dcm = '0; 
assign i_ch1_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch1_pld_rx_clk2_dcm = '0; 
assign i_ch20_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch20_pld_rx_clk2_dcm = '0; 
assign i_ch21_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch21_pld_rx_clk2_dcm = '0; 
assign i_ch22_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch22_pld_rx_clk2_dcm = '0; 
assign i_ch23_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch23_pld_rx_clk2_dcm = '0; 
assign i_ch2_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch2_pld_rx_clk2_dcm = '0; 
assign i_ch3_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch3_pld_rx_clk2_dcm = '0; 
assign i_ch4_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch4_pld_rx_clk2_dcm = '0; 
assign i_ch5_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch5_pld_rx_clk2_dcm = '0; 
assign i_ch6_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch6_pld_rx_clk2_dcm = '0; 
assign i_ch7_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch7_pld_rx_clk2_dcm = '0; 
assign i_ch8_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch8_pld_rx_clk2_dcm = '0; 
assign i_ch9_pld_fpll_shared_direct_async_in_dcm[1:0] = '0; 
assign i_ch9_pld_rx_clk2_dcm = '0; 
assign i_aux_por_vccl_ovr = '0; 
assign i_id[3:0] = '0; 
assign i_jtag_tck = '0; 
assign i_jtag_tdi = '0; 
assign i_jtag_tms = '0; 
assign i_jtag_trst = '0; 
assign i_sens_therm = '0; 
assign i_strap_spare_in0 = '0; 
assign i_strap_spare_in1 = '0; 
assign i_edm_in = '0; 
assign s0_0_1__maib_rotate__maib_rotate = '0; 
assign s0_187_1__aib_jtag_return__tdo = '0; 
assign s1_0_1__aib_jtag_out__tck = '0; 
assign s1_0_1__aib_jtag_out__tdi = '0; 
assign s1_0_1__aib_jtag_out__tms = '0; 
assign s1_0_1__dts_temptrip__temptrip = '0; 
assign s2_0_1__aib_jtag_out__tck = '0; 
assign s2_0_1__aib_jtag_out__tdi = '0; 
assign s2_0_1__aib_jtag_out__tms = '0; 
assign s2_187_1__aib_jtag_return__tdo = '0; 
assign s4_0_1__aib_cjtag_ctrl_id__cjtag_id[3:0] = '0; 
assign s5_187_1__cnoc__abort = '0; 
assign s5_187_1__cnoc__clk = '0; 
assign s5_187_1__cnoc__clk_n = '0; 
assign s5_187_1__cnoc__data[32:0] = '0; 
assign s5_187_1__cnoc__end_of_packet = '0; 
assign s5_187_1__cnoc__nonsecure_interrupt = '0; 
assign s5_187_1__cnoc__por = '0; 
assign s5_187_1__cnoc__por_n = '0; 
assign s5_187_1__cnoc__secure_interrupt = '0; 
assign s5_187_1__cnoc__start_of_packet = '0; 
assign s5_187_1__cnoc__sync = '0; 
assign s5_187_1__cnoc__valid = '0; 
assign s5_187_1__cnoc__warm_reset_n = '0; 
assign s8_187_1__aib_jtag_return__tdo = '0; 
assign s9_0_1__aib_jtag_out__tck = '0; 
assign s9_0_1__aib_jtag_out__tdi = '0; 
assign s9_0_1__aib_jtag_out__tms = '0; 
assign s11_187_1__aib_jtag_out__tck = '0; 
assign s11_187_1__aib_jtag_out__tdi = '0; 
assign s11_187_1__aib_jtag_out__tms = '0; 
assign s12_187_1__aib_jtag_out__tck = '0; 
assign s12_187_1__aib_jtag_out__tdi = '0; 
assign s12_187_1__aib_jtag_out__tms = '0; 
assign s13_0_1__aib_jtag_return__tdo = '0; 
assign s14_0_1__cjtag__tck = '0; 
assign s14_0_1__cjtag__tdi = '0; 
assign s14_0_1__cjtag__tms = '0; 
assign s14_187_1__aib_cjtag_ctrl_id__cjtag_id[3:0] = '0; 
assign s15_187_1__cjtag__tck = '0; 
assign s15_187_1__cjtag__tdi = '0; 
assign s15_187_1__cjtag__tms = '0; 
assign s16_0_1__aib_jtag_return__tdo = '0; 
assign s17_187_1__cjtag_return__tdo = '0; 
assign s18_0_1__aib_jtag_return__tdo = '0; 
assign s19_187_1__aib_jtag_out__tck = '0; 
assign s19_187_1__aib_jtag_out__tdi = '0; 
assign s19_187_1__aib_jtag_out__tms = '0; 
assign s20_187_1__cnoc__abort = '0; 
assign s20_187_1__cnoc__clk = '0; 
assign s20_187_1__cnoc__clk_n = '0; 
assign s20_187_1__cnoc__data[32:0] = '0; 
assign s20_187_1__cnoc__end_of_packet = '0; 
assign s20_187_1__cnoc__nonsecure_interrupt = '0; 
assign s20_187_1__cnoc__por = '0; 
assign s20_187_1__cnoc__por_n = '0; 
assign s20_187_1__cnoc__secure_interrupt = '0; 
assign s20_187_1__cnoc__start_of_packet = '0; 
assign s20_187_1__cnoc__sync = '0; 
assign s20_187_1__cnoc__valid = '0; 
assign s20_187_1__cnoc__warm_reset_n = '0; 
assign s21_0_1__cjtag_return__tdo = '0; 
assign s23_0_1__cnoc__abort = '0; 
assign s23_0_1__cnoc__clk = '0; 
assign s23_0_1__cnoc__clk_n = '0; 
assign s23_0_1__cnoc__data[32:0] = '0; 
assign s23_0_1__cnoc__end_of_packet = '0; 
assign s23_0_1__cnoc__nonsecure_interrupt = '0; 
assign s23_0_1__cnoc__por = '0; 
assign s23_0_1__cnoc__por_n = '0; 
assign s23_0_1__cnoc__secure_interrupt = '0; 
assign s23_0_1__cnoc__start_of_packet = '0; 
assign s23_0_1__cnoc__sync = '0; 
assign s23_0_1__cnoc__valid = '0; 
assign s23_0_1__cnoc__warm_reset_n = '0; 
assign s23_187_1__include_aib_jtag_segment__include_aib_jtag_segment = '0; 
assign s25_187_1__include_aib_jtag_segment__include_aib_jtag_segment = '0; 
assign s27_187_1__include_aib_jtag_segment__include_aib_jtag_segment = '0; 
assign s28_187_1__dts_temptrip__temptrip = '0; 
assign s30_0_1__dc_bsc_sdata__s_data = '0; 
assign s30_187_1__dc_bsc_sdata__s_data = '0; 
assign s32_187_1__sdm_mission_bus__clk = '0; 
assign s32_187_1__sdm_mission_bus__data[31:0] = '0; 
assign s32_187_1__sdm_mission_bus__valid = '0; 
assign s33_187_1__sdm_test_bus__data[27:0] = '0; 
assign s34_0_1__sdm_testmode_ctrl__test_io_ctrl[15:0] = '0; 
assign s37_0_1__test_return__data[15:0] = '0; 
assign s37_0_1__test_return__valid = '0; 
assign s38_0_1__scan_sdm_so__scan_out[4:0] = '0; 
assign s39_0_1__cr_ctrl__muxsel_avst[3:0] = '0; 
assign s39_0_1__cr_ctrl__muxsel_test_cnoc = '0; 
assign s124_0_1__include_aib_jtag_segment__include_aib_jtag_segment = '0; 
assign s126_0_1__include_aib_jtag_segment__include_aib_jtag_segment = '0; 
assign s128_0_1__include_aib_jtag_segment__include_aib_jtag_segment = '0; 
assign i_s0_3_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_8_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_9_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_10_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_15_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_16_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_21_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_22_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_23_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_24_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_25_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_30_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_31_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_36_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_37_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_38_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_43_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_44_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_45_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_46_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_47_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_48_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_49_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_50_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_55_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_56_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_57_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_62_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_63_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_68_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_69_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_70_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_71_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_72_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_77_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_78_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_83_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_84_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_85_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_90_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_91_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_92_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_93_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_94_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_95_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_96_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_97_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_102_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_103_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_104_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_109_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_110_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_115_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_116_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_117_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_118_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_119_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_124_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_125_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_130_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_131_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_132_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_137_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_138_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_139_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_140_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_141_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_142_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_143_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_144_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_149_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_150_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_151_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_156_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_157_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_162_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_163_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_164_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_165_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_166_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_171_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_172_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_177_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_178_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_179_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_184_1__core_periphery__clock_from_core[15:0] = '0; 
assign i_s0_3_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_9_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_10_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_15_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_16_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_21_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_22_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_23_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_24_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_25_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_30_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_31_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_36_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_37_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_38_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_43_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_44_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_45_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_46_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_47_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_48_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_49_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_50_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_55_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_56_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_57_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_62_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_63_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_68_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_69_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_70_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_71_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_72_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_77_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_78_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_83_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_84_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_90_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_91_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_92_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_93_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_94_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_95_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_96_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_97_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_102_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_103_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_104_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_109_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_110_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_115_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_116_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_117_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_118_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_119_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_124_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_125_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_130_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_131_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_132_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_137_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_138_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_139_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_140_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_141_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_142_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_143_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_144_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_149_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_150_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_151_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_156_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_157_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_162_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_163_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_164_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_165_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_166_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_171_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_172_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_177_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_178_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_179_1__core_periphery__data_from_core[95:0] = '0; 
assign i_s0_184_1__core_periphery__data_from_core[95:0] = '0; 
assign s0_4_1__core_periphery__data_from_core_unused[59:38] = '0; 
assign s0_4_1__core_periphery__data_from_core_unused[36:0] = '0; 
assign s0_5_1__core_periphery__data_from_core_unused[34] = '0; 
assign s0_5_1__core_periphery__data_from_core_unused[32:28] = '0; 
assign s0_5_1__core_periphery__data_from_core_unused[23:15] = '0; 
assign s0_5_1__core_periphery__data_from_core_unused[12:0] = '0; 
assign vcc_dts_ref = '0; 
assign vcce_pll_ref = '0; 
assign i_ch0_user_avmm1_clk_rowclk = '0; 
assign i_ch0_pld_rx_clk2_rowclk = '0; 
assign i_ch10_pld_rx_clk2_rowclk = '0; 
assign i_ch10_user_avmm1_clk_rowclk = '0; 
assign i_ch10_user_avmm2_clk_rowclk = '0; 
assign i_ch11_pld_rx_clk2_rowclk = '0; 
assign i_ch11_user_avmm1_clk_rowclk = '0; 
assign i_ch11_user_avmm2_clk_rowclk = '0; 
assign i_ch12_pld_rx_clk2_rowclk = '0; 
assign i_ch12_user_avmm1_clk_rowclk = '0; 
assign i_ch12_user_avmm2_clk_rowclk = '0; 
assign i_ch13_pld_rx_clk2_rowclk = '0; 
assign i_ch13_user_avmm1_clk_rowclk = '0; 
assign i_ch13_user_avmm2_clk_rowclk = '0; 
assign i_ch14_pld_rx_clk2_rowclk = '0; 
assign i_ch14_user_avmm1_clk_rowclk = '0; 
assign i_ch14_user_avmm2_clk_rowclk = '0; 
assign i_ch15_pld_rx_clk2_rowclk = '0; 
assign i_ch15_user_avmm1_clk_rowclk = '0; 
assign i_ch15_user_avmm2_clk_rowclk = '0; 
assign i_ch16_pld_rx_clk2_rowclk = '0; 
assign i_ch16_user_avmm1_clk_rowclk = '0; 
assign i_ch16_user_avmm2_clk_rowclk = '0; 
assign i_ch17_pld_rx_clk2_rowclk = '0; 
assign i_ch17_user_avmm1_clk_rowclk = '0; 
assign i_ch17_user_avmm2_clk_rowclk = '0; 
assign i_ch18_pld_rx_clk2_rowclk = '0; 
assign i_ch18_user_avmm1_clk_rowclk = '0; 
assign i_ch18_user_avmm2_clk_rowclk = '0; 
assign i_ch19_pld_rx_clk2_rowclk = '0; 
assign i_ch19_user_avmm1_clk_rowclk = '0; 
assign i_ch19_user_avmm2_clk_rowclk = '0; 
assign i_ch1_pld_rx_clk2_rowclk = '0; 
assign i_ch1_user_avmm1_clk_rowclk = '0; 
assign i_ch1_user_avmm2_clk_rowclk = '0; 
assign i_ch20_pld_rx_clk2_rowclk = '0; 
assign i_ch20_user_avmm1_clk_rowclk = '0; 
assign i_ch20_user_avmm2_clk_rowclk = '0; 
assign i_ch21_pld_rx_clk2_rowclk = '0; 
assign i_ch21_user_avmm1_clk_rowclk = '0; 
assign i_ch21_user_avmm2_clk_rowclk = '0; 
assign i_ch22_pld_rx_clk2_rowclk = '0; 
assign i_ch22_user_avmm1_clk_rowclk = '0; 
assign i_ch22_user_avmm2_clk_rowclk = '0; 
assign i_ch23_pld_rx_clk2_rowclk = '0; 
assign i_ch23_user_avmm1_clk_rowclk = '0; 
assign i_ch23_user_avmm2_clk_rowclk = '0; 
assign i_ch2_pld_rx_clk2_rowclk = '0; 
assign i_ch2_user_avmm1_clk_rowclk = '0; 
assign i_ch2_user_avmm2_clk_rowclk = '0; 
assign i_ch3_pld_rx_clk2_rowclk = '0; 
assign i_ch3_user_avmm1_clk_rowclk = '0; 
assign i_ch3_user_avmm2_clk_rowclk = '0; 
assign i_ch4_pld_rx_clk2_rowclk = '0; 
assign i_ch4_user_avmm1_clk_rowclk = '0; 
assign i_ch4_user_avmm2_clk_rowclk = '0; 
assign i_ch5_pld_rx_clk2_rowclk = '0; 
assign i_ch5_user_avmm1_clk_rowclk = '0; 
assign i_ch5_user_avmm2_clk_rowclk = '0; 
assign i_ch6_pld_rx_clk2_rowclk = '0; 
assign i_ch6_user_avmm1_clk_rowclk = '0; 
assign i_ch6_user_avmm2_clk_rowclk = '0; 
assign i_ch7_pld_rx_clk2_rowclk = '0; 
assign i_ch7_user_avmm1_clk_rowclk = '0; 
assign i_ch7_user_avmm2_clk_rowclk = '0; 
assign i_ch8_pld_rx_clk2_rowclk = '0; 
assign i_ch8_user_avmm1_clk_rowclk = '0; 
assign i_ch8_user_avmm2_clk_rowclk = '0; 
assign i_ch9_pld_rx_clk2_rowclk = '0; 
assign i_ch9_user_avmm1_clk_rowclk = '0; 
assign i_ch9_user_avmm2_clk_rowclk = '0; 
assign s0_100_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_100_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_101_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_101_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_105_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_105_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_106_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_106_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_107_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_107_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_108_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_108_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_111_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_111_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_112_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_112_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_113_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_113_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_114_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_114_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_11_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_11_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_120_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_120_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_121_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_121_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_122_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_122_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_123_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_123_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_126_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_126_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_127_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_127_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_128_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_128_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_129_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_129_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_12_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_12_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_133_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_133_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_134_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_134_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_135_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_135_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_136_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_136_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_13_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_13_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_145_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_145_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_146_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_146_1__core_periphery__data_from_core_unused[34:28] = '0; 
assign s0_146_1__core_periphery__data_from_core_unused[26:0] = '0; 
assign s0_147_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_147_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_148_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_148_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_14_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_14_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_152_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_152_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_153_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_153_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_154_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_154_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_155_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_155_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_158_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_158_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_159_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_159_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_160_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_160_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_161_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_161_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_167_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_167_1__core_periphery__data_from_core_unused[72:0] = '0; 
assign s0_168_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_168_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_169_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_169_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_170_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_170_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_173_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_173_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_174_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_174_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_175_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_175_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_176_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_176_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_17_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_17_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_180_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_180_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_181_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_181_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_182_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_182_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_183_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_183_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_18_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_18_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_19_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_19_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_20_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_20_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_26_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_26_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_27_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_27_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_28_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_28_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_29_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_29_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_32_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_32_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_33_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_33_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_34_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_34_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_35_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_35_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_39_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_39_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_40_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_40_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_41_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_41_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_42_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_42_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_4_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_51_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_51_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_52_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_52_1__core_periphery__data_from_core_unused[34:28] = '0; 
assign s0_52_1__core_periphery__data_from_core_unused[26:0] = '0; 
assign s0_53_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_53_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_54_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_54_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_58_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_58_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_59_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_59_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_5_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_60_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_60_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_61_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_61_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_64_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_64_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_65_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_65_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_66_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_66_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_67_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_67_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_6_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_6_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_73_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_73_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_74_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_74_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_75_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_75_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_76_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_76_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_79_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_79_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_7_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_7_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_80_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_80_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_81_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_81_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_82_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_82_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_85_1__core_periphery__data_from_core_unused[93:0] = '0; 
assign s0_86_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_86_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_87_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_87_1__core_periphery__data_from_core_unused[34:0] = '0; 
assign s0_88_1__core_periphery__clock_from_core_unused[13:0] = '0; 
assign s0_88_1__core_periphery__data_from_core_unused[21:0] = '0; 
assign s0_89_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_89_1__core_periphery__data_from_core_unused[66:0] = '0; 
assign s0_8_1__core_periphery__data_from_core_unused[64:0] = '0; 
assign s0_98_1__core_periphery__clock_from_core_unused[14:0] = '0; 
assign s0_98_1__core_periphery__data_from_core_unused[59:0] = '0; 
assign s0_99_1__core_periphery__clock_from_core_unused[9:0] = '0; 
assign s0_99_1__core_periphery__data_from_core_unused[34:28] = '0; 
assign s0_99_1__core_periphery__data_from_core_unused[26:0] = '0; 
assign p0_link_up_o = '0; 
assign p0_dl_up_o = '0; 
assign p0_pm_curnt_state_o[7:0] = '0; 
assign p0_pm_dstate_o[31:0] = '0; 

assign ch13_pipe_direct_pld_rx_clk1_dcm = '0; 
assign ch13_pipe_direct_pld_tx_clk1_dcm = '0; 
assign ch14_pipe_direct_pld_rx_clk1_dcm = '0; 
assign ch14_pipe_direct_pld_tx_clk1_dcm = '0; 
assign ch15_pipe_direct_pld_rx_clk1_dcm = '0; 
assign ch15_pipe_direct_pld_tx_clk1_dcm = '0; 
assign ch16_pipe_direct_pld_rx_clk1_dcm = '0; 
assign ch16_pipe_direct_pld_tx_clk1_dcm = '0; 
assign ch17_pipe_direct_pld_rx_clk1_dcm = '0; 
assign ch17_pipe_direct_pld_tx_clk1_dcm = '0; 
assign ch18_pipe_direct_pld_rx_clk1_dcm = '0; 
assign ch18_pipe_direct_pld_tx_clk1_dcm = '0; 
assign ch19_pipe_direct_pld_rx_clk1_dcm = '0; 
assign ch19_pipe_direct_pld_tx_clk1_dcm = '0; 
assign ch20_pipe_direct_pld_rx_clk1_dcm = '0; 
assign ch20_pipe_direct_pld_tx_clk1_dcm = '0; 
assign ch21_pipe_direct_pld_rx_clk1_dcm = '0; 
assign ch21_pipe_direct_pld_tx_clk1_dcm = '0; 
assign ch22_pipe_direct_pld_rx_clk1_dcm = '0; 
assign ch22_pipe_direct_pld_tx_clk1_dcm = '0; 

assign ch13_pipe_direct_pld_adapter_rx_pld_rst_n = '0; 
assign ch13_pipe_direct_pld_rx_dll_lock_req = '0; 
assign ch13_pipe_direct_pld_adapter_tx_pld_rst_n = '0; 
assign ch13_pipe_direct_pld_tx_dll_lock_req = '0; 
assign ch14_pipe_direct_pld_adapter_rx_pld_rst_n = '0; 
assign ch14_pipe_direct_pld_rx_dll_lock_req = '0; 
assign ch14_pipe_direct_pld_adapter_tx_pld_rst_n = '0; 
assign ch14_pipe_direct_pld_tx_dll_lock_req = '0; 
assign ch15_pipe_direct_pld_adapter_rx_pld_rst_n = '0; 
assign ch15_pipe_direct_pld_rx_dll_lock_req = '0; 
assign ch15_pipe_direct_pld_adapter_tx_pld_rst_n = '0; 
assign ch15_pipe_direct_pld_tx_dll_lock_req = '0; 
assign ch16_pipe_direct_pld_adapter_rx_pld_rst_n = '0; 
assign ch16_pipe_direct_pld_rx_dll_lock_req = '0; 
assign ch16_pipe_direct_pld_adapter_tx_pld_rst_n = '0; 
assign ch16_pipe_direct_pld_tx_dll_lock_req = '0; 
assign ch17_pipe_direct_pld_adapter_rx_pld_rst_n = '0; 
assign ch17_pipe_direct_pld_rx_dll_lock_req = '0; 
assign ch17_pipe_direct_pld_adapter_tx_pld_rst_n = '0; 
assign ch17_pipe_direct_pld_tx_dll_lock_req = '0; 
assign ch18_pipe_direct_pld_adapter_rx_pld_rst_n = '0; 
assign ch18_pipe_direct_pld_rx_dll_lock_req = '0; 
assign ch18_pipe_direct_pld_adapter_tx_pld_rst_n = '0; 
assign ch18_pipe_direct_pld_tx_dll_lock_req = '0; 
assign ch19_pipe_direct_pld_adapter_rx_pld_rst_n = '0; 
assign ch19_pipe_direct_pld_rx_dll_lock_req = '0; 
assign ch19_pipe_direct_pld_adapter_tx_pld_rst_n = '0; 
assign ch19_pipe_direct_pld_tx_dll_lock_req = '0; 
assign ch20_pipe_direct_pld_adapter_rx_pld_rst_n = '0; 
assign ch20_pipe_direct_pld_rx_dll_lock_req = '0; 
assign ch20_pipe_direct_pld_adapter_tx_pld_rst_n = '0; 
assign ch20_pipe_direct_pld_tx_dll_lock_req = '0; 
assign ch21_pipe_direct_pld_adapter_rx_pld_rst_n = '0; 
assign ch21_pipe_direct_pld_rx_dll_lock_req = '0; 
assign ch21_pipe_direct_pld_adapter_tx_pld_rst_n = '0; 
assign ch21_pipe_direct_pld_tx_dll_lock_req = '0; 
assign ch22_pipe_direct_pld_adapter_rx_pld_rst_n = '0; 
assign ch22_pipe_direct_pld_rx_dll_lock_req = '0; 
assign ch22_pipe_direct_pld_adapter_tx_pld_rst_n = '0; 
assign ch22_pipe_direct_pld_tx_dll_lock_req = '0; 

generate 
   if (hssi_ctr_topology == "pipe_direct_cxl_x8") begin : pipe_direct_cxl_x8
      // PIPE Direct Signals 
      assign octet1_pipe_direct_synthfast_lockstatus_o                     = pipe_direct_rx_octet1_synthfast_lockstatus1;
      assign octet1_pipe_direct_synthfast_ready_o                          = pipe_direct_rx_octet1_synthfast_ready1;
      assign octet1_pipe_direct_synthslow_lockstatus_o                     = pipe_direct_rx_octet1_synthslow_lockstatus1;
      assign octet1_pipe_direct_synthslow_ready_o                          = pipe_direct_rx_octet1_synthslow_ready1;
      assign pipe_direct_pld_tx_clk_out_o                            = ch15_pipe_direct_pld_pcs_tx_clk_out1_dcm;
      assign ln0_pipe_direct_pld_rx_clk_out_o                        = ch15_pipe_direct_pld_pcs_rx_clk_out1_dcm;
      assign ln1_pipe_direct_pld_rx_clk_out_o                        = ch16_pipe_direct_pld_pcs_rx_clk_out1_dcm;
      assign ln2_pipe_direct_pld_rx_clk_out_o                        = ch17_pipe_direct_pld_pcs_rx_clk_out1_dcm;
      assign ln3_pipe_direct_pld_rx_clk_out_o                        = ch18_pipe_direct_pld_pcs_rx_clk_out1_dcm;
      assign ln4_pipe_direct_pld_rx_clk_out_o                        = ch19_pipe_direct_pld_pcs_rx_clk_out1_dcm;
      assign ln5_pipe_direct_pld_rx_clk_out_o                        = ch20_pipe_direct_pld_pcs_rx_clk_out1_dcm;
      assign ln6_pipe_direct_pld_rx_clk_out_o                        = ch21_pipe_direct_pld_pcs_rx_clk_out1_dcm;
      assign ln7_pipe_direct_pld_rx_clk_out_o                        = ch22_pipe_direct_pld_pcs_rx_clk_out1_dcm;
      assign ln0_pipe_direct_reserved_o = 12'h000;
      assign ln1_pipe_direct_reserved_o = 12'h000;
      assign ln2_pipe_direct_reserved_o = 12'h000;
      assign ln3_pipe_direct_reserved_o = 12'h000;
      assign ln4_pipe_direct_reserved_o = 12'h000;
      assign ln5_pipe_direct_reserved_o = 12'h000;
      assign ln6_pipe_direct_reserved_o = 12'h000;
      assign ln7_pipe_direct_reserved_o = 12'h000;
      //
      // CH13 TX : Deskew
      assign ch13_pipe_direct_tx_octet1[77:20]                       = '1;
      assign ch13_pipe_direct_tx_octet1[19]                          = ln7_pipe_direct_rxtermination_i;
      assign ch13_pipe_direct_tx_octet1[18]                          = ln6_pipe_direct_rxtermination_i;
      assign ch13_pipe_direct_tx_octet1[17]                          = ln5_pipe_direct_rxtermination_i;
      assign ch13_pipe_direct_tx_octet1[16]                          = ln4_pipe_direct_rxtermination_i;
      assign ch13_pipe_direct_tx_octet1[15]                          = ln3_pipe_direct_rxtermination_i;
      assign ch13_pipe_direct_tx_octet1[14]                          = ln2_pipe_direct_rxtermination_i;
      assign ch13_pipe_direct_tx_octet1[13]                          = ln1_pipe_direct_rxtermination_i;
      assign ch13_pipe_direct_tx_octet1[12]                          = ln0_pipe_direct_rxtermination_i;
      assign ch13_pipe_direct_tx_octet1[11]                          = ln7_pipe_direct_pclkchangeack_i;
      assign ch13_pipe_direct_tx_octet1[10]                          = ln6_pipe_direct_pclkchangeack_i;
      assign ch13_pipe_direct_tx_octet1[9]                           = ln5_pipe_direct_pclkchangeack_i;
      assign ch13_pipe_direct_tx_octet1[8]                           = ln4_pipe_direct_pclkchangeack_i;
      assign ch13_pipe_direct_tx_octet1[7]                           = ln3_pipe_direct_pclkchangeack_i;
      assign ch13_pipe_direct_tx_octet1[6]                           = ln2_pipe_direct_pclkchangeack_i;
      assign ch13_pipe_direct_tx_octet1[5]                           = ln1_pipe_direct_pclkchangeack_i;
      assign ch13_pipe_direct_tx_octet1[4]                           = ln0_pipe_direct_pclkchangeack_i;
      assign ch13_pipe_direct_tx_octet1[3]                           = octet1_pipe_direct_deskew_clear_3_i;
      assign ch13_pipe_direct_tx_octet1[2]                           = octet1_pipe_direct_deskew_clear_2_i;
      assign ch13_pipe_direct_tx_octet1[1]                           = octet1_pipe_direct_deskew_clear_1_i;
      assign ch13_pipe_direct_tx_octet1[0]                           = octet1_pipe_direct_deskew_clear_0_i;
      // CH13 RX : Deskew
      assign ln7_pipe_direct_rxstandbystatus_o                       = ch13_pipe_direct_rx_octet1[71];
      assign ln6_pipe_direct_rxstandbystatus_o                       = ch13_pipe_direct_rx_octet1[70];
      assign ln5_pipe_direct_rxstandbystatus_o                       = ch13_pipe_direct_rx_octet1[69];
      assign ln4_pipe_direct_rxstandbystatus_o                       = ch13_pipe_direct_rx_octet1[68];
      assign ln3_pipe_direct_rxstandbystatus_o                       = ch13_pipe_direct_rx_octet1[67];
      assign ln2_pipe_direct_rxstandbystatus_o                       = ch13_pipe_direct_rx_octet1[66];
      assign ln1_pipe_direct_rxstandbystatus_o                       = ch13_pipe_direct_rx_octet1[65];
      assign ln0_pipe_direct_rxstandbystatus_o                       = ch13_pipe_direct_rx_octet1[64];
      assign ln7_pipe_direct_pclkchangeok_o                          = ch13_pipe_direct_rx_octet1[63];
      assign ln6_pipe_direct_pclkchangeok_o                          = ch13_pipe_direct_rx_octet1[62];
      assign ln5_pipe_direct_pclkchangeok_o                          = ch13_pipe_direct_rx_octet1[61];
      assign ln4_pipe_direct_pclkchangeok_o                          = ch13_pipe_direct_rx_octet1[60];
      assign ln3_pipe_direct_pclkchangeok_o                          = ch13_pipe_direct_rx_octet1[59];
      assign ln2_pipe_direct_pclkchangeok_o                          = ch13_pipe_direct_rx_octet1[58];
      assign ln1_pipe_direct_pclkchangeok_o                          = ch13_pipe_direct_rx_octet1[57];
      assign ln0_pipe_direct_pclkchangeok_o                          = ch13_pipe_direct_rx_octet1[56];
      assign ln7_pipe_direct_rxstatus_o                              = ch13_pipe_direct_rx_octet1[55];
      assign ln6_pipe_direct_rxstatus_o                              = ch13_pipe_direct_rx_octet1[54];
      assign ln5_pipe_direct_rxstatus_o                              = ch13_pipe_direct_rx_octet1[53];
      assign ln4_pipe_direct_rxstatus_o                              = ch13_pipe_direct_rx_octet1[52];
      assign ln3_pipe_direct_rxstatus_o                              = ch13_pipe_direct_rx_octet1[51];
      assign ln2_pipe_direct_rxstatus_o                              = ch13_pipe_direct_rx_octet1[50];
      assign ln1_pipe_direct_rxstatus_o                              = ch13_pipe_direct_rx_octet1[49];
      assign ln0_pipe_direct_rxstatus_o                              = ch13_pipe_direct_rx_octet1[48];
      assign ln7_pipe_direct_phystatus_o                             = ch13_pipe_direct_rx_octet1[47];
      assign ln6_pipe_direct_phystatus_o                             = ch13_pipe_direct_rx_octet1[46];
      assign ln5_pipe_direct_phystatus_o                             = ch13_pipe_direct_rx_octet1[45];
      assign ln4_pipe_direct_phystatus_o                             = ch13_pipe_direct_rx_octet1[44];
      assign ln3_pipe_direct_phystatus_o                             = ch13_pipe_direct_rx_octet1[43];
      assign ln2_pipe_direct_phystatus_o                             = ch13_pipe_direct_rx_octet1[42];
      assign ln1_pipe_direct_phystatus_o                             = ch13_pipe_direct_rx_octet1[41];
      assign ln0_pipe_direct_phystatus_o                             = ch13_pipe_direct_rx_octet1[40];
      assign octet1_pipe_direct_phy_dsk_active_chans_o[7:0]          = ch13_pipe_direct_rx_octet1[39:32];
      assign octet1_pipe_direct_phy_dsk_monitor_err_o[7:0]           = ch13_pipe_direct_rx_octet1[31:24];
      assign octet1_pipe_direct_phy_dsk_monitor_err_status_3_o       = ch13_pipe_direct_rx_octet1[23];
      assign octet1_pipe_direct_phy_dsk_status_3_o[2:0]              = ch13_pipe_direct_rx_octet1[22:20];
      assign octet1_pipe_direct_phy_dsk_valid_3_o                    = ch13_pipe_direct_rx_octet1[19];
      assign octet1_pipe_direct_phy_dsk_eval_done_3_o                = ch13_pipe_direct_rx_octet1[18];
      assign octet1_pipe_direct_phy_dsk_monitor_err_status_2_o       = ch13_pipe_direct_rx_octet1[17];
      assign octet1_pipe_direct_phy_dsk_status_2_o[2:0]              = ch13_pipe_direct_rx_octet1[16:14];
      assign octet1_pipe_direct_phy_dsk_valid_2_o                    = ch13_pipe_direct_rx_octet1[13];
      assign octet1_pipe_direct_phy_dsk_eval_done_2_o                = ch13_pipe_direct_rx_octet1[12];
      assign octet1_pipe_direct_phy_dsk_monitor_err_status_1_o       = ch13_pipe_direct_rx_octet1[11];
      assign octet1_pipe_direct_phy_dsk_status_1_o[2:0]              = ch13_pipe_direct_rx_octet1[10:8];
      assign octet1_pipe_direct_phy_dsk_valid_1_o                    = ch13_pipe_direct_rx_octet1[7];
      assign octet1_pipe_direct_phy_dsk_eval_done_1_o                = ch13_pipe_direct_rx_octet1[6];
      assign octet1_pipe_direct_phy_dsk_monitor_err_status_0_o       = ch13_pipe_direct_rx_octet1[5];
      assign octet1_pipe_direct_phy_dsk_status_0_o[2:0]              = ch13_pipe_direct_rx_octet1[4:2];
      assign octet1_pipe_direct_phy_dsk_valid_0_o                    = ch13_pipe_direct_rx_octet1[1];
      assign octet1_pipe_direct_phy_dsk_eval_done_0_o                = ch13_pipe_direct_rx_octet1[0];
      // CH14 TX : MSG Channel
      assign ch14_pipe_direct_tx_octet1[77:64]                       = '1;
      assign ch14_pipe_direct_tx_octet1[63:56]                       = ln7_m2p_messagebus_i;
      assign ch14_pipe_direct_tx_octet1[55:48]                       = ln6_m2p_messagebus_i;
      assign ch14_pipe_direct_tx_octet1[47:40]                       = ln5_m2p_messagebus_i;
      assign ch14_pipe_direct_tx_octet1[39:32]                       = ln4_m2p_messagebus_i;
      assign ch14_pipe_direct_tx_octet1[31:24]                       = ln3_m2p_messagebus_i;
      assign ch14_pipe_direct_tx_octet1[23:16]                       = ln2_m2p_messagebus_i;
      assign ch14_pipe_direct_tx_octet1[15:8]                        = ln1_m2p_messagebus_i;
      assign ch14_pipe_direct_tx_octet1[7:0]                         = ln0_m2p_messagebus_i;
      // CH14 RX : MSG Channel
      assign ln7_p2m_messagebus_o                                    = ch14_pipe_direct_rx_octet1[63:56];
      assign ln6_p2m_messagebus_o                                    = ch14_pipe_direct_rx_octet1[55:48];
      assign ln5_p2m_messagebus_o                                    = ch14_pipe_direct_rx_octet1[47:40];
      assign ln4_p2m_messagebus_o                                    = ch14_pipe_direct_rx_octet1[39:32];
      assign ln3_p2m_messagebus_o                                    = ch14_pipe_direct_rx_octet1[31:24];
      assign ln2_p2m_messagebus_o                                    = ch14_pipe_direct_rx_octet1[23:16];
      assign ln1_p2m_messagebus_o                                    = ch14_pipe_direct_rx_octet1[15:8];
      assign ln0_p2m_messagebus_o                                    = ch14_pipe_direct_rx_octet1[7:0];
      
      // CH15 TX : PIPE DIRECT 
      assign ch15_pipe_direct_tx_octet1[77]                          = ln0_pipe_direct_txdeskewmarker_i;
      assign ch15_pipe_direct_tx_octet1[76]                          = ln0_pipe_direct_rxstandby_i;
      assign ch15_pipe_direct_tx_octet1[75:72]                       = ln0_pipe_direct_txelecidle_i;
      assign ch15_pipe_direct_tx_octet1[71:70]                       = ln0_pipe_direct_powerdown_i;
      assign ch15_pipe_direct_tx_octet1[69:67]                       = ln0_pipe_direct_rate_i;
      assign ch15_pipe_direct_tx_octet1[66]                          = ln0_pipe_direct_txdetectrx_i;
      assign ch15_pipe_direct_tx_octet1[65]                          = ln0_pipe_direct_txdatavalid1_i;
      assign ch15_pipe_direct_tx_octet1[64]                          = ln0_pipe_direct_txdatavalid0_i;
      assign ch15_pipe_direct_tx_octet1[63:0]                        = ln0_pipe_direct_txdata_i;
      assign ch15_pipe_direct_tx_octet1_PLD_PCS_rst_n_l8             = ln0_pipe_direct_pld_pcs_rst_n_i;
      // CH15 RX : PIPE DIRECT 
      assign ln0_pipe_direct_rxdatavalid1_o                                      = ch15_pipe_direct_rx_octet1[65];
      assign ln0_pipe_direct_rxdatavalid0_o                                      = ch15_pipe_direct_rx_octet1[64];
      assign ln0_pipe_direct_rxdata_o                                            = ch15_pipe_direct_rx_octet1[63:0];
      assign ln0_pipe_direct_rxelecidle_o                                        = ch15_pipe_direct_rx_octet1_RXElecIdle_l8;
      assign ln0_pipe_direct_cdrlockstatus_o                      = ch15_pipe_direct_rx_octet1_rx_cdrlockstatus_l8;
      assign ln0_pipe_direct_cdrlock2data_o                       = ch15_pipe_direct_rx_octet1_rx_cdrlock2data_l8;
      
      // CH16 TX : PIPE DIRECT 
      assign ch16_pipe_direct_tx_octet1[77]                          = ln1_pipe_direct_txdeskewmarker_i;
      assign ch16_pipe_direct_tx_octet1[76]                          = ln1_pipe_direct_rxstandby_i;
      assign ch16_pipe_direct_tx_octet1[75:72]                       = ln1_pipe_direct_txelecidle_i;
      assign ch16_pipe_direct_tx_octet1[71:70]                       = ln1_pipe_direct_powerdown_i;
      assign ch16_pipe_direct_tx_octet1[69:67]                       = ln1_pipe_direct_rate_i;
      assign ch16_pipe_direct_tx_octet1[66]                          = ln1_pipe_direct_txdetectrx_i;
      assign ch16_pipe_direct_tx_octet1[65]                          = ln1_pipe_direct_txdatavalid1_i;
      assign ch16_pipe_direct_tx_octet1[64]                          = ln1_pipe_direct_txdatavalid0_i;
      assign ch16_pipe_direct_tx_octet1[63:0]                        = ln1_pipe_direct_txdata_i;
      assign ch16_pipe_direct_tx_octet1_PLD_PCS_rst_n_l9             = ln1_pipe_direct_pld_pcs_rst_n_i;
      // CH16 RX : PIPE DIRECT 
      assign ln1_pipe_direct_rxdatavalid1_o                                      = ch16_pipe_direct_rx_octet1[65];
      assign ln1_pipe_direct_rxdatavalid0_o                                      = ch16_pipe_direct_rx_octet1[64];
      assign ln1_pipe_direct_rxdata_o                                            = ch16_pipe_direct_rx_octet1[63:0];
      assign ln1_pipe_direct_rxelecidle_o                                        = ch16_pipe_direct_rx_octet1_RXElecIdle_l9;
      assign ln1_pipe_direct_cdrlockstatus_o                      = ch16_pipe_direct_rx_octet1_rx_cdrlockstatus_l9;
      assign ln1_pipe_direct_cdrlock2data_o                       = ch16_pipe_direct_rx_octet1_rx_cdrlock2data_l9;
      
      // CH17 TX : PIPE DIRECT 
      assign ch17_pipe_direct_tx_octet1[77]                          = ln2_pipe_direct_txdeskewmarker_i;
      assign ch17_pipe_direct_tx_octet1[76]                          = ln2_pipe_direct_rxstandby_i;
      assign ch17_pipe_direct_tx_octet1[75:72]                       = ln2_pipe_direct_txelecidle_i;
      assign ch17_pipe_direct_tx_octet1[71:70]                       = ln2_pipe_direct_powerdown_i;
      assign ch17_pipe_direct_tx_octet1[69:67]                       = ln2_pipe_direct_rate_i;
      assign ch17_pipe_direct_tx_octet1[66]                          = ln2_pipe_direct_txdetectrx_i;
      assign ch17_pipe_direct_tx_octet1[65]                          = ln2_pipe_direct_txdatavalid1_i;
      assign ch17_pipe_direct_tx_octet1[64]                          = ln2_pipe_direct_txdatavalid0_i;
      assign ch17_pipe_direct_tx_octet1[63:0]                        = ln2_pipe_direct_txdata_i;
      assign ch17_pipe_direct_tx_octet1_PLD_PCS_rst_n_l10            = ln2_pipe_direct_pld_pcs_rst_n_i;
      // CH17 RX : PIPE DIRECT 
      assign ln2_pipe_direct_rxdatavalid1_o                                      = ch17_pipe_direct_rx_octet1[65];
      assign ln2_pipe_direct_rxdatavalid0_o                                      = ch17_pipe_direct_rx_octet1[64];
      assign ln2_pipe_direct_rxdata_o                                            = ch17_pipe_direct_rx_octet1[63:0];
      assign ln2_pipe_direct_rxelecidle_o                                        = ch17_pipe_direct_rx_octet1_RXElecIdle_l10;
      assign ln2_pipe_direct_cdrlockstatus_o                      = ch17_pipe_direct_rx_octet1_rx_cdrlockstatus_l10;
      assign ln2_pipe_direct_cdrlock2data_o                       = ch17_pipe_direct_rx_octet1_rx_cdrlock2data_l10;
      
      // CH18 TX : PIPE DIRECT 
      assign ch18_pipe_direct_tx_octet1[77]                          = ln3_pipe_direct_txdeskewmarker_i;
      assign ch18_pipe_direct_tx_octet1[76]                          = ln3_pipe_direct_rxstandby_i;
      assign ch18_pipe_direct_tx_octet1[75:72]                       = ln3_pipe_direct_txelecidle_i;
      assign ch18_pipe_direct_tx_octet1[71:70]                       = ln3_pipe_direct_powerdown_i;
      assign ch18_pipe_direct_tx_octet1[69:67]                       = ln3_pipe_direct_rate_i;
      assign ch18_pipe_direct_tx_octet1[66]                          = ln3_pipe_direct_txdetectrx_i;
      assign ch18_pipe_direct_tx_octet1[65]                          = ln3_pipe_direct_txdatavalid1_i;
      assign ch18_pipe_direct_tx_octet1[64]                          = ln3_pipe_direct_txdatavalid0_i;
      assign ch18_pipe_direct_tx_octet1[63:0]                        = ln3_pipe_direct_txdata_i;
      assign ch18_pipe_direct_tx_octet1_PLD_PCS_rst_n_l11            = ln3_pipe_direct_pld_pcs_rst_n_i;
      // CH18 RX : PIPE DIRECT 
      assign ln3_pipe_direct_rxdatavalid1_o                                      = ch18_pipe_direct_rx_octet1[65];
      assign ln3_pipe_direct_rxdatavalid0_o                                      = ch18_pipe_direct_rx_octet1[64];
      assign ln3_pipe_direct_rxdata_o                                            = ch18_pipe_direct_rx_octet1[63:0];
      assign ln3_pipe_direct_rxelecidle_o                                        = ch18_pipe_direct_rx_octet1_RXElecIdle_l11;
      assign ln3_pipe_direct_cdrlockstatus_o                      = ch18_pipe_direct_rx_octet1_rx_cdrlockstatus_l11;
      assign ln3_pipe_direct_cdrlock2data_o                       = ch18_pipe_direct_rx_octet1_rx_cdrlock2data_l11;
      
      // CH19 TX : PIPE DIRECT 
      assign ch19_pipe_direct_tx_octet1[77]                          = ln4_pipe_direct_txdeskewmarker_i;
      assign ch19_pipe_direct_tx_octet1[76]                          = ln4_pipe_direct_rxstandby_i;
      assign ch19_pipe_direct_tx_octet1[75:72]                       = ln4_pipe_direct_txelecidle_i;
      assign ch19_pipe_direct_tx_octet1[71:70]                       = ln4_pipe_direct_powerdown_i;
      assign ch19_pipe_direct_tx_octet1[69:67]                       = ln4_pipe_direct_rate_i;
      assign ch19_pipe_direct_tx_octet1[66]                          = ln4_pipe_direct_txdetectrx_i;
      assign ch19_pipe_direct_tx_octet1[65]                          = ln4_pipe_direct_txdatavalid1_i;
      assign ch19_pipe_direct_tx_octet1[64]                          = ln4_pipe_direct_txdatavalid0_i;
      assign ch19_pipe_direct_tx_octet1[63:0]                        = ln4_pipe_direct_txdata_i;
      assign ch19_pipe_direct_tx_octet1_PLD_PCS_rst_n_l12            = ln4_pipe_direct_pld_pcs_rst_n_i;
      // CH19 RX : PIPE DIRECT 
      assign ln4_pipe_direct_rxdatavalid1_o                                      = ch19_pipe_direct_rx_octet1[65];
      assign ln4_pipe_direct_rxdatavalid0_o                                      = ch19_pipe_direct_rx_octet1[64];
      assign ln4_pipe_direct_rxdata_o                                            = ch19_pipe_direct_rx_octet1[63:0];
      assign ln4_pipe_direct_rxelecidle_o                                        = ch19_pipe_direct_rx_octet1_RXElecIdle_l12;
      assign ln4_pipe_direct_cdrlockstatus_o                      = ch19_pipe_direct_rx_octet1_rx_cdrlockstatus_l12;
      assign ln4_pipe_direct_cdrlock2data_o                       = ch19_pipe_direct_rx_octet1_rx_cdrlock2data_l12;
      
      // CH20 TX : PIPE DIRECT 
      assign ch20_pipe_direct_tx_octet1[77]                          = ln5_pipe_direct_txdeskewmarker_i;
      assign ch20_pipe_direct_tx_octet1[76]                          = ln5_pipe_direct_rxstandby_i;
      assign ch20_pipe_direct_tx_octet1[75:72]                       = ln5_pipe_direct_txelecidle_i;
      assign ch20_pipe_direct_tx_octet1[71:70]                       = ln5_pipe_direct_powerdown_i;
      assign ch20_pipe_direct_tx_octet1[69:67]                       = ln5_pipe_direct_rate_i;
      assign ch20_pipe_direct_tx_octet1[66]                          = ln5_pipe_direct_txdetectrx_i;
      assign ch20_pipe_direct_tx_octet1[65]                          = ln5_pipe_direct_txdatavalid1_i;
      assign ch20_pipe_direct_tx_octet1[64]                          = ln5_pipe_direct_txdatavalid0_i;
      assign ch20_pipe_direct_tx_octet1[63:0]                        = ln5_pipe_direct_txdata_i;
      assign ch20_pipe_direct_tx_octet1_PLD_PCS_rst_n_l13            = ln5_pipe_direct_pld_pcs_rst_n_i;
      // CH20 RX : PIPE DIRECT 
      assign ln5_pipe_direct_rxdatavalid1_o                                      = ch20_pipe_direct_rx_octet1[65];
      assign ln5_pipe_direct_rxdatavalid0_o                                      = ch20_pipe_direct_rx_octet1[64];
      assign ln5_pipe_direct_rxdata_o                                            = ch20_pipe_direct_rx_octet1[63:0];
      assign ln5_pipe_direct_rxelecidle_o                                        = ch20_pipe_direct_rx_octet1_RXElecIdle_l13;
      assign ln5_pipe_direct_cdrlockstatus_o                      = ch20_pipe_direct_rx_octet1_rx_cdrlockstatus_l13;
      assign ln5_pipe_direct_cdrlock2data_o                       = ch20_pipe_direct_rx_octet1_rx_cdrlock2data_l13;
      
      // CH21 TX : PIPE DIRECT 
      assign ch21_pipe_direct_tx_octet1[77]                          = ln6_pipe_direct_txdeskewmarker_i;
      assign ch21_pipe_direct_tx_octet1[76]                          = ln6_pipe_direct_rxstandby_i;
      assign ch21_pipe_direct_tx_octet1[75:72]                       = ln6_pipe_direct_txelecidle_i;
      assign ch21_pipe_direct_tx_octet1[71:70]                       = ln6_pipe_direct_powerdown_i;
      assign ch21_pipe_direct_tx_octet1[69:67]                       = ln6_pipe_direct_rate_i;
      assign ch21_pipe_direct_tx_octet1[66]                          = ln6_pipe_direct_txdetectrx_i;
      assign ch21_pipe_direct_tx_octet1[65]                          = ln6_pipe_direct_txdatavalid1_i;
      assign ch21_pipe_direct_tx_octet1[64]                          = ln6_pipe_direct_txdatavalid0_i;
      assign ch21_pipe_direct_tx_octet1[63:0]                        = ln6_pipe_direct_txdata_i;
      assign ch21_pipe_direct_tx_octet1_PLD_PCS_rst_n_l14            = ln6_pipe_direct_pld_pcs_rst_n_i;
      // CH21 RX : PIPE DIRECT 
      assign ln6_pipe_direct_rxdatavalid1_o                                      = ch21_pipe_direct_rx_octet1[65];
      assign ln6_pipe_direct_rxdatavalid0_o                                      = ch21_pipe_direct_rx_octet1[64];
      assign ln6_pipe_direct_rxdata_o                                            = ch21_pipe_direct_rx_octet1[63:0];
      assign ln6_pipe_direct_rxelecidle_o                                        = ch21_pipe_direct_rx_octet1_RXElecIdle_l14;
      assign ln6_pipe_direct_cdrlockstatus_o                      = ch21_pipe_direct_rx_octet1_rx_cdrlockstatus_l14;
      assign ln6_pipe_direct_cdrlock2data_o                       = ch21_pipe_direct_rx_octet1_rx_cdrlock2data_l14;
      
      // CH22 TX : PIPE DIRECT 
      assign ch22_pipe_direct_tx_octet1[77]                          = ln7_pipe_direct_txdeskewmarker_i;
      assign ch22_pipe_direct_tx_octet1[76]                          = ln7_pipe_direct_rxstandby_i;
      assign ch22_pipe_direct_tx_octet1[75:72]                       = ln7_pipe_direct_txelecidle_i;
      assign ch22_pipe_direct_tx_octet1[71:70]                       = ln7_pipe_direct_powerdown_i;
      assign ch22_pipe_direct_tx_octet1[69:67]                       = ln7_pipe_direct_rate_i;
      assign ch22_pipe_direct_tx_octet1[66]                          = ln7_pipe_direct_txdetectrx_i;
      assign ch22_pipe_direct_tx_octet1[65]                          = ln7_pipe_direct_txdatavalid1_i;
      assign ch22_pipe_direct_tx_octet1[64]                          = ln7_pipe_direct_txdatavalid0_i;
      assign ch22_pipe_direct_tx_octet1[63:0]                        = ln7_pipe_direct_txdata_i;
      assign ch22_pipe_direct_tx_octet1_PLD_PCS_rst_n_l15            = ln7_pipe_direct_pld_pcs_rst_n_i;
      // CH22 RX : PIPE DIRECT 
      assign ln7_pipe_direct_rxdatavalid1_o                                      = ch22_pipe_direct_rx_octet1[65];
      assign ln7_pipe_direct_rxdatavalid0_o                                      = ch22_pipe_direct_rx_octet1[64];
      assign ln7_pipe_direct_rxdata_o                                            = ch22_pipe_direct_rx_octet1[63:0];
      assign ln7_pipe_direct_rxelecidle_o                                        = ch22_pipe_direct_rx_octet1_RXElecIdle_l15;
      assign ln7_pipe_direct_cdrlockstatus_o                      = ch22_pipe_direct_rx_octet1_rx_cdrlockstatus_l15;
      assign ln7_pipe_direct_cdrlock2data_o                       = ch22_pipe_direct_rx_octet1_rx_cdrlock2data_l15;
   // TODO end
   // TODO else begin
   // TODO    assign ch13_pipe_direct_tx_octet1[77:0]                        = '0;
   // TODO    assign ch14_pipe_direct_tx_octet1[77:0]                        = '0;
   // TODO    assign ch15_pipe_direct_tx_octet1[77:0]                        = '0;
   // TODO    assign ch16_pipe_direct_tx_octet1[77:0]                        = '0;
   // TODO    assign ch17_pipe_direct_tx_octet1[77:0]                        = '0;
   // TODO    assign ch18_pipe_direct_tx_octet1[77:0]                        = '0;
   // TODO    assign ch19_pipe_direct_tx_octet1[77:0]                        = '0;
   // TODO    assign ch20_pipe_direct_tx_octet1[77:0]                        = '0;
   // TODO    assign ch21_pipe_direct_tx_octet1[77:0]                        = '0;
   // TODO    assign ch22_pipe_direct_tx_octet1[77:0]                        = '0;
   // TODO end
   end else begin : cxl_x16
      assign ch13_pipe_direct_tx_octet1[77:0] = '0; 
      assign ch14_pipe_direct_tx_octet1[77:0] = '0; 
      assign ch15_pipe_direct_tx_octet1[77:0] = '0; 
      assign ch16_pipe_direct_tx_octet1[77:0] = '0; 
      assign ch17_pipe_direct_tx_octet1[77:0] = '0; 
      assign ch18_pipe_direct_tx_octet1[77:0] = '0; 
      assign ch19_pipe_direct_tx_octet1[77:0] = '0; 
      assign ch20_pipe_direct_tx_octet1[77:0] = '0; 
      assign ch21_pipe_direct_tx_octet1[77:0] = '0; 
      assign ch22_pipe_direct_tx_octet1[77:0] = '0; 
      assign ch15_pipe_direct_tx_octet1_PLD_PCS_rst_n_l8 = '0; 
      assign ch16_pipe_direct_tx_octet1_PLD_PCS_rst_n_l9 = '0; 
      assign ch17_pipe_direct_tx_octet1_PLD_PCS_rst_n_l10 = '0; 
      assign ch18_pipe_direct_tx_octet1_PLD_PCS_rst_n_l11 = '0; 
      assign ch19_pipe_direct_tx_octet1_PLD_PCS_rst_n_l12 = '0; 
      assign ch20_pipe_direct_tx_octet1_PLD_PCS_rst_n_l13 = '0; 
      assign ch21_pipe_direct_tx_octet1_PLD_PCS_rst_n_l14 = '0; 
      assign ch22_pipe_direct_tx_octet1_PLD_PCS_rst_n_l15 = '0; 
   end
endgenerate

// assign s0_182_1__core_periphery__data_from_core[71] = '0; 
// assign fifo_out[609:0] = '0; 
// assign fifo_out[561:0] = '0; 
 z1578a_mdx1 # (
   .qhip_csb2wire_en_hwtcl                                                                                                              (qhip_csb2wire_en_hwtcl),
   .qhip_mmio_enable_hwtcl                                                                                                              (qhip_mmio_enable_hwtcl),
   .opt_tx_big_buffer_hwtcl                                                                                                             (opt_tx_big_buffer_hwtcl),
   .opt_csb_pll_en_hwtcl                                                                                                                (opt_csb_pll_en_hwtcl),
   .opt_cache_formatb_en_hwtcl                                                                                                          (opt_cache_formatb_en_hwtcl),
   .opt_chemem_flow_err_det_en_hwtcl                                                                                                    (opt_chemem_flow_err_det_en_hwtcl),
   .hssi_aib_ssm_silicon_rev                                                                                                            ( hssi_aib_ssm_silicon_rev),
   .hssi_aibnd_rx_0_aib_ber_margining_ctrl                                                                                              ( hssi_aibnd_rx_0_aib_ber_margining_ctrl),
   .hssi_aibnd_rx_0_aib_datasel_gr0                                                                                                     ( hssi_aibnd_rx_0_aib_datasel_gr0),
   .hssi_aibnd_rx_0_aib_datasel_gr1                                                                                                     ( hssi_aibnd_rx_0_aib_datasel_gr1),
   .hssi_aibnd_rx_0_aib_datasel_gr2                                                                                                     ( hssi_aibnd_rx_0_aib_datasel_gr2),
   .hssi_aibnd_rx_0_aib_dllstr_align_clkdiv                                                                                             ( hssi_aibnd_rx_0_aib_dllstr_align_clkdiv),
   .hssi_aibnd_rx_0_aib_dllstr_align_dly_pst                                                                                            ( hssi_aibnd_rx_0_aib_dllstr_align_dly_pst),
   .hssi_aibnd_rx_0_aib_dllstr_align_dy_ctl_static                                                                                      ( hssi_aibnd_rx_0_aib_dllstr_align_dy_ctl_static),
   .hssi_aibnd_rx_0_aib_dllstr_align_dy_ctlsel                                                                                          ( hssi_aibnd_rx_0_aib_dllstr_align_dy_ctlsel),
   .hssi_aibnd_rx_0_aib_dllstr_align_entest                                                                                             ( hssi_aibnd_rx_0_aib_dllstr_align_entest),
   .hssi_aibnd_rx_0_aib_dllstr_align_halfcode                                                                                           ( hssi_aibnd_rx_0_aib_dllstr_align_halfcode),
   .hssi_aibnd_rx_0_aib_dllstr_align_selflock                                                                                           ( hssi_aibnd_rx_0_aib_dllstr_align_selflock),
   .hssi_aibnd_rx_0_aib_dllstr_align_st_core_dn_prgmnvrt                                                                                ( hssi_aibnd_rx_0_aib_dllstr_align_st_core_dn_prgmnvrt),
   .hssi_aibnd_rx_0_aib_dllstr_align_st_core_up_prgmnvrt                                                                                ( hssi_aibnd_rx_0_aib_dllstr_align_st_core_up_prgmnvrt),
   .hssi_aibnd_rx_0_aib_dllstr_align_st_core_updnen                                                                                     ( hssi_aibnd_rx_0_aib_dllstr_align_st_core_updnen),
   .hssi_aibnd_rx_0_aib_dllstr_align_st_dftmuxsel                                                                                       ( hssi_aibnd_rx_0_aib_dllstr_align_st_dftmuxsel),
   .hssi_aibnd_rx_0_aib_dllstr_align_st_en                                                                                              ( hssi_aibnd_rx_0_aib_dllstr_align_st_en),
   .hssi_aibnd_rx_0_aib_dllstr_align_st_hps_ctrl_en                                                                                     ( hssi_aibnd_rx_0_aib_dllstr_align_st_hps_ctrl_en),
   .hssi_aibnd_rx_0_aib_dllstr_align_st_lockreq_muxsel                                                                                  ( hssi_aibnd_rx_0_aib_dllstr_align_st_lockreq_muxsel),
   .hssi_aibnd_rx_0_aib_dllstr_align_st_new_dll                                                                                         ( hssi_aibnd_rx_0_aib_dllstr_align_st_new_dll),
   .hssi_aibnd_rx_0_aib_dllstr_align_st_rst                                                                                             ( hssi_aibnd_rx_0_aib_dllstr_align_st_rst),
   .hssi_aibnd_rx_0_aib_dllstr_align_st_rst_prgmnvrt                                                                                    ( hssi_aibnd_rx_0_aib_dllstr_align_st_rst_prgmnvrt),
   .hssi_aibnd_rx_0_aib_dllstr_align_test_clk_pll_en_n                                                                                  ( hssi_aibnd_rx_0_aib_dllstr_align_test_clk_pll_en_n),
   .hssi_aibnd_rx_0_aib_inctrl_gr0                                                                                                      ( hssi_aibnd_rx_0_aib_inctrl_gr0),
   .hssi_aibnd_rx_0_aib_inctrl_gr1                                                                                                      ( hssi_aibnd_rx_0_aib_inctrl_gr1),
   .hssi_aibnd_rx_0_aib_inctrl_gr2                                                                                                      ( hssi_aibnd_rx_0_aib_inctrl_gr2),
   .hssi_aibnd_rx_0_aib_inctrl_gr3                                                                                                      ( hssi_aibnd_rx_0_aib_inctrl_gr3),
   .hssi_aibnd_rx_0_aib_outctrl_gr0                                                                                                     ( hssi_aibnd_rx_0_aib_outctrl_gr0),
   .hssi_aibnd_rx_0_aib_outctrl_gr1                                                                                                     ( hssi_aibnd_rx_0_aib_outctrl_gr1),
   .hssi_aibnd_rx_0_aib_outctrl_gr2                                                                                                     ( hssi_aibnd_rx_0_aib_outctrl_gr2),
   .hssi_aibnd_rx_0_aib_outndrv_r12                                                                                                     ( hssi_aibnd_rx_0_aib_outndrv_r12),
   .hssi_aibnd_rx_0_aib_outndrv_r34                                                                                                     ( hssi_aibnd_rx_0_aib_outndrv_r34),
   .hssi_aibnd_rx_0_aib_outndrv_r56                                                                                                     ( hssi_aibnd_rx_0_aib_outndrv_r56),
   .hssi_aibnd_rx_0_aib_outndrv_r78                                                                                                     ( hssi_aibnd_rx_0_aib_outndrv_r78),
   .hssi_aibnd_rx_0_aib_outpdrv_r12                                                                                                     ( hssi_aibnd_rx_0_aib_outpdrv_r12),
   .hssi_aibnd_rx_0_aib_outpdrv_r34                                                                                                     ( hssi_aibnd_rx_0_aib_outpdrv_r34),
   .hssi_aibnd_rx_0_aib_outpdrv_r56                                                                                                     ( hssi_aibnd_rx_0_aib_outpdrv_r56),
   .hssi_aibnd_rx_0_aib_outpdrv_r78                                                                                                     ( hssi_aibnd_rx_0_aib_outpdrv_r78),
   .hssi_aibnd_rx_0_aib_red_shift_en                                                                                                    ( hssi_aibnd_rx_0_aib_red_shift_en),
   .hssi_aibnd_rx_0_dft_hssitestip_dll_dcc_en                                                                                           ( hssi_aibnd_rx_0_dft_hssitestip_dll_dcc_en),
   .hssi_aibnd_rx_0_op_mode                                                                                                             ( hssi_aibnd_rx_0_op_mode),
   .hssi_aibnd_rx_0_powerdown_mode                                                                                                      ( hssi_aibnd_rx_0_powerdown_mode),
   .hssi_aibnd_rx_0_powermode_ac                                                                                                        ( hssi_aibnd_rx_0_powermode_ac),
   .hssi_aibnd_rx_0_powermode_dc                                                                                                        ( hssi_aibnd_rx_0_powermode_dc),
   .hssi_aibnd_rx_0_powermode_freq_hz_aib_hssi_rx_transfer_clk                                                                          ( hssi_aibnd_rx_0_powermode_freq_hz_aib_hssi_rx_transfer_clk),
   .hssi_aibnd_rx_0_redundancy_en                                                                                                       ( hssi_aibnd_rx_0_redundancy_en),
   .hssi_aibnd_rx_0_sup_mode                                                                                                            ( hssi_aibnd_rx_0_sup_mode),
   .hssi_aibnd_rx_0_silicon_rev                                                                                                         ( hssi_aibnd_rx_0_silicon_rev),
   .hssi_aibnd_tx_0_aib_datasel_gr0                                                                                                     ( hssi_aibnd_tx_0_aib_datasel_gr0),
   .hssi_aibnd_tx_0_aib_datasel_gr1                                                                                                     ( hssi_aibnd_tx_0_aib_datasel_gr1),
   .hssi_aibnd_tx_0_aib_datasel_gr2                                                                                                     ( hssi_aibnd_tx_0_aib_datasel_gr2),
   .hssi_aibnd_tx_0_aib_datasel_gr3                                                                                                     ( hssi_aibnd_tx_0_aib_datasel_gr3),
   .hssi_aibnd_tx_0_aib_ddrctrl_gr0                                                                                                     ( hssi_aibnd_tx_0_aib_ddrctrl_gr0),
   .hssi_aibnd_tx_0_aib_hssi_tx_transfer_clk_hz                                                                                         ( hssi_aibnd_tx_0_aib_hssi_tx_transfer_clk_hz),
   .hssi_aibnd_tx_0_aib_iinasyncen                                                                                                      ( hssi_aibnd_tx_0_aib_iinasyncen),
   .hssi_aibnd_tx_0_aib_iinclken                                                                                                        ( hssi_aibnd_tx_0_aib_iinclken),
   .hssi_aibnd_tx_0_aib_outctrl_gr0                                                                                                     ( hssi_aibnd_tx_0_aib_outctrl_gr0),
   .hssi_aibnd_tx_0_aib_outctrl_gr1                                                                                                     ( hssi_aibnd_tx_0_aib_outctrl_gr1),
   .hssi_aibnd_tx_0_aib_outctrl_gr2                                                                                                     ( hssi_aibnd_tx_0_aib_outctrl_gr2),
   .hssi_aibnd_tx_0_aib_outctrl_gr3                                                                                                     ( hssi_aibnd_tx_0_aib_outctrl_gr3),
   .hssi_aibnd_tx_0_aib_outndrv_r34                                                                                                     ( hssi_aibnd_tx_0_aib_outndrv_r34),
   .hssi_aibnd_tx_0_aib_outndrv_r56                                                                                                     ( hssi_aibnd_tx_0_aib_outndrv_r56),
   .hssi_aibnd_tx_0_aib_outpdrv_r34                                                                                                     ( hssi_aibnd_tx_0_aib_outpdrv_r34),
   .hssi_aibnd_tx_0_aib_outpdrv_r56                                                                                                     ( hssi_aibnd_tx_0_aib_outpdrv_r56),
   .hssi_aibnd_tx_0_aib_red_dirclkn_shiften                                                                                             ( hssi_aibnd_tx_0_aib_red_dirclkn_shiften),
   .hssi_aibnd_tx_0_aib_red_dirclkp_shiften                                                                                             ( hssi_aibnd_tx_0_aib_red_dirclkp_shiften),
   .hssi_aibnd_tx_0_aib_red_drx_shiften                                                                                                 ( hssi_aibnd_tx_0_aib_red_drx_shiften),
   .hssi_aibnd_tx_0_aib_red_dtx_shiften                                                                                                 ( hssi_aibnd_tx_0_aib_red_dtx_shiften),
   .hssi_aibnd_tx_0_aib_red_pout_shiften                                                                                                ( hssi_aibnd_tx_0_aib_red_pout_shiften),
   .hssi_aibnd_tx_0_aib_red_rx_shiften                                                                                                  ( hssi_aibnd_tx_0_aib_red_rx_shiften),
   .hssi_aibnd_tx_0_aib_red_tx_shiften                                                                                                  ( hssi_aibnd_tx_0_aib_red_tx_shiften),
   .hssi_aibnd_tx_0_aib_red_txferclkout_shiften                                                                                         ( hssi_aibnd_tx_0_aib_red_txferclkout_shiften),
   .hssi_aibnd_tx_0_aib_red_txferclkoutn_shiften                                                                                        ( hssi_aibnd_tx_0_aib_red_txferclkoutn_shiften),
   .hssi_aibnd_tx_0_aib_tx_clkdiv                                                                                                       ( hssi_aibnd_tx_0_aib_tx_clkdiv),
   .hssi_aibnd_tx_0_aib_tx_dcc_byp                                                                                                      ( hssi_aibnd_tx_0_aib_tx_dcc_byp),
   .hssi_aibnd_tx_0_aib_tx_dcc_byp_iocsr_unused                                                                                         ( hssi_aibnd_tx_0_aib_tx_dcc_byp_iocsr_unused),
   .hssi_aibnd_tx_0_aib_tx_dcc_cont_cal                                                                                                 ( hssi_aibnd_tx_0_aib_tx_dcc_cont_cal),
   .hssi_aibnd_tx_0_aib_tx_dcc_cont_cal_iocsr_unused                                                                                    ( hssi_aibnd_tx_0_aib_tx_dcc_cont_cal_iocsr_unused),
   .hssi_aibnd_tx_0_aib_tx_dcc_dft                                                                                                      ( hssi_aibnd_tx_0_aib_tx_dcc_dft),
   .hssi_aibnd_tx_0_aib_tx_dcc_dft_sel                                                                                                  ( hssi_aibnd_tx_0_aib_tx_dcc_dft_sel),
   .hssi_aibnd_tx_0_aib_tx_dcc_dll_dft_sel                                                                                              ( hssi_aibnd_tx_0_aib_tx_dcc_dll_dft_sel),
   .hssi_aibnd_tx_0_aib_tx_dcc_dll_entest                                                                                               ( hssi_aibnd_tx_0_aib_tx_dcc_dll_entest),
   .hssi_aibnd_tx_0_aib_tx_dcc_dy_ctl_static                                                                                            ( hssi_aibnd_tx_0_aib_tx_dcc_dy_ctl_static),
   .hssi_aibnd_tx_0_aib_tx_dcc_dy_ctlsel                                                                                                ( hssi_aibnd_tx_0_aib_tx_dcc_dy_ctlsel),
   .hssi_aibnd_tx_0_aib_tx_dcc_en                                                                                                       ( hssi_aibnd_tx_0_aib_tx_dcc_en),
   .hssi_aibnd_tx_0_aib_tx_dcc_en_iocsr_unused                                                                                          ( hssi_aibnd_tx_0_aib_tx_dcc_en_iocsr_unused),
   .hssi_aibnd_tx_0_aib_tx_dcc_manual_dn                                                                                                ( hssi_aibnd_tx_0_aib_tx_dcc_manual_dn),
   .hssi_aibnd_tx_0_aib_tx_dcc_manual_up                                                                                                ( hssi_aibnd_tx_0_aib_tx_dcc_manual_up),
   .hssi_aibnd_tx_0_aib_tx_dcc_rst_prgmnvrt                                                                                             ( hssi_aibnd_tx_0_aib_tx_dcc_rst_prgmnvrt),
   .hssi_aibnd_tx_0_aib_tx_dcc_st_core_dn_prgmnvrt                                                                                      ( hssi_aibnd_tx_0_aib_tx_dcc_st_core_dn_prgmnvrt),
   .hssi_aibnd_tx_0_aib_tx_dcc_st_core_up_prgmnvrt                                                                                      ( hssi_aibnd_tx_0_aib_tx_dcc_st_core_up_prgmnvrt),
   .hssi_aibnd_tx_0_aib_tx_dcc_st_core_updnen                                                                                           ( hssi_aibnd_tx_0_aib_tx_dcc_st_core_updnen),
   .hssi_aibnd_tx_0_aib_tx_dcc_st_dftmuxsel                                                                                             ( hssi_aibnd_tx_0_aib_tx_dcc_st_dftmuxsel),
   .hssi_aibnd_tx_0_aib_tx_dcc_st_dly_pst                                                                                               ( hssi_aibnd_tx_0_aib_tx_dcc_st_dly_pst),
   .hssi_aibnd_tx_0_aib_tx_dcc_st_en                                                                                                    ( hssi_aibnd_tx_0_aib_tx_dcc_st_en),
   .hssi_aibnd_tx_0_aib_tx_dcc_st_hps_ctrl_en                                                                                           ( hssi_aibnd_tx_0_aib_tx_dcc_st_hps_ctrl_en),
   .hssi_aibnd_tx_0_aib_tx_dcc_st_lockreq_muxsel                                                                                        ( hssi_aibnd_tx_0_aib_tx_dcc_st_lockreq_muxsel),
   .hssi_aibnd_tx_0_aib_tx_dcc_st_new_dll                                                                                               ( hssi_aibnd_tx_0_aib_tx_dcc_st_new_dll),
   .hssi_aibnd_tx_0_aib_tx_dcc_st_rst                                                                                                   ( hssi_aibnd_tx_0_aib_tx_dcc_st_rst),
   .hssi_aibnd_tx_0_aib_tx_dcc_test_clk_pll_en_n                                                                                        ( hssi_aibnd_tx_0_aib_tx_dcc_test_clk_pll_en_n),
   .hssi_aibnd_tx_0_aib_tx_halfcode                                                                                                     ( hssi_aibnd_tx_0_aib_tx_halfcode),
   .hssi_aibnd_tx_0_aib_tx_selflock                                                                                                     ( hssi_aibnd_tx_0_aib_tx_selflock),
   .hssi_aibnd_tx_0_dfd_dll_dcc_en                                                                                                      ( hssi_aibnd_tx_0_dfd_dll_dcc_en),
   .hssi_aibnd_tx_0_dft_hssitestip_dll_dcc_en                                                                                           ( hssi_aibnd_tx_0_dft_hssitestip_dll_dcc_en),
   .hssi_aibnd_tx_0_op_mode                                                                                                             ( hssi_aibnd_tx_0_op_mode),
   .hssi_aibnd_tx_0_powerdown_mode                                                                                                      ( hssi_aibnd_tx_0_powerdown_mode),
   .hssi_aibnd_tx_0_powermode_ac                                                                                                        ( hssi_aibnd_tx_0_powermode_ac),
   .hssi_aibnd_tx_0_powermode_dc                                                                                                        ( hssi_aibnd_tx_0_powermode_dc),
   .hssi_aibnd_tx_0_powermode_freq_hz_aib_hssi_tx_transfer_clk                                                                          ( hssi_aibnd_tx_0_powermode_freq_hz_aib_hssi_tx_transfer_clk),
   .hssi_aibnd_tx_0_redundancy_en                                                                                                       ( hssi_aibnd_tx_0_redundancy_en),
   .hssi_aibnd_tx_0_sup_mode                                                                                                            ( hssi_aibnd_tx_0_sup_mode),
   .hssi_aibnd_tx_0_silicon_rev                                                                                                         ( hssi_aibnd_tx_0_silicon_rev),
   .hssi_pldadapt_tx_0_aib_clk1_sel                                                                                                     ( hssi_pldadapt_tx_0_aib_clk1_sel),
   .hssi_pldadapt_tx_0_aib_clk2_sel                                                                                                     ( hssi_pldadapt_tx_0_aib_clk2_sel),
   .hssi_pldadapt_tx_0_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                            ( hssi_pldadapt_tx_0_hdpldadapt_aib_fabric_pld_pma_hclk_hz),
   .hssi_pldadapt_tx_0_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz                                                                          ( hssi_pldadapt_tx_0_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz),
   .hssi_pldadapt_tx_0_hdpldadapt_aib_fabric_tx_sr_clk_in_hz                                                                            ( hssi_pldadapt_tx_0_hdpldadapt_aib_fabric_tx_sr_clk_in_hz),
   .hssi_pldadapt_tx_0_bonding_dft_en                                                                                                   ( hssi_pldadapt_tx_0_bonding_dft_en),
   .hssi_pldadapt_tx_0_bonding_dft_val                                                                                                  ( hssi_pldadapt_tx_0_bonding_dft_val),
   .hssi_pldadapt_tx_0_chnl_bonding                                                                                                     ( hssi_pldadapt_tx_0_chnl_bonding),
   .hssi_pldadapt_tx_0_comp_cnt                                                                                                         ( hssi_pldadapt_tx_0_comp_cnt),
   .hssi_pldadapt_tx_0_compin_sel                                                                                                       ( hssi_pldadapt_tx_0_compin_sel),
   .hssi_pldadapt_tx_0_hdpldadapt_csr_clk_hz                                                                                            ( hssi_pldadapt_tx_0_hdpldadapt_csr_clk_hz),
   .hssi_pldadapt_tx_0_ctrl_plane_bonding                                                                                               ( hssi_pldadapt_tx_0_ctrl_plane_bonding),
   .hssi_pldadapt_tx_0_ds_bypass_pipeln                                                                                                 ( hssi_pldadapt_tx_0_ds_bypass_pipeln),
   .hssi_pldadapt_tx_0_ds_last_chnl                                                                                                     ( hssi_pldadapt_tx_0_ds_last_chnl),
   .hssi_pldadapt_tx_0_ds_master                                                                                                        ( hssi_pldadapt_tx_0_ds_master),
   .hssi_pldadapt_tx_0_duplex_mode                                                                                                      ( hssi_pldadapt_tx_0_duplex_mode),
   .hssi_pldadapt_tx_0_dv_bond                                                                                                          ( hssi_pldadapt_tx_0_dv_bond),
   .hssi_pldadapt_tx_0_dv_gen                                                                                                           ( hssi_pldadapt_tx_0_dv_gen),
   .hssi_pldadapt_tx_0_fifo_double_write                                                                                                ( hssi_pldadapt_tx_0_fifo_double_write),
   .hssi_pldadapt_tx_0_fifo_mode                                                                                                        ( hssi_pldadapt_tx_0_fifo_mode),
   .hssi_pldadapt_tx_0_fifo_rd_clk_frm_gen_scg_en                                                                                       ( hssi_pldadapt_tx_0_fifo_rd_clk_frm_gen_scg_en),
   .hssi_pldadapt_tx_0_fifo_rd_clk_scg_en                                                                                               ( hssi_pldadapt_tx_0_fifo_rd_clk_scg_en),
   .hssi_pldadapt_tx_0_fifo_rd_clk_sel                                                                                                  ( hssi_pldadapt_tx_0_fifo_rd_clk_sel),
   .hssi_pldadapt_tx_0_fifo_stop_rd                                                                                                     ( hssi_pldadapt_tx_0_fifo_stop_rd),
   .hssi_pldadapt_tx_0_fifo_stop_wr                                                                                                     ( hssi_pldadapt_tx_0_fifo_stop_wr),
   .hssi_pldadapt_tx_0_fifo_width                                                                                                       ( hssi_pldadapt_tx_0_fifo_width),
   .hssi_pldadapt_tx_0_fifo_wr_clk_scg_en                                                                                               ( hssi_pldadapt_tx_0_fifo_wr_clk_scg_en),
   .hssi_pldadapt_tx_0_fpll_shared_direct_async_in_sel                                                                                  ( hssi_pldadapt_tx_0_fpll_shared_direct_async_in_sel),
   .hssi_pldadapt_tx_0_frmgen_burst                                                                                                     ( hssi_pldadapt_tx_0_frmgen_burst),
   .hssi_pldadapt_tx_0_frmgen_bypass                                                                                                    ( hssi_pldadapt_tx_0_frmgen_bypass),
   .hssi_pldadapt_tx_0_frmgen_mfrm_length                                                                                               ( hssi_pldadapt_tx_0_frmgen_mfrm_length),
   .hssi_pldadapt_tx_0_frmgen_pipeln                                                                                                    ( hssi_pldadapt_tx_0_frmgen_pipeln),
   .hssi_pldadapt_tx_0_frmgen_pyld_ins                                                                                                  ( hssi_pldadapt_tx_0_frmgen_pyld_ins),
   .hssi_pldadapt_tx_0_frmgen_wordslip                                                                                                  ( hssi_pldadapt_tx_0_frmgen_wordslip),
   .hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit0_rst_val                                                                                      ( hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit0_rst_val),
   .hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit1_rst_val                                                                                      ( hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit1_rst_val),
   .hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit2_rst_val                                                                                      ( hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit2_rst_val),
   .hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit3_rst_val                                                                                      ( hssi_pldadapt_tx_0_fsr_hip_fsr_in_bit3_rst_val),
   .hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit0_rst_val                                                                                     ( hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit0_rst_val),
   .hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit1_rst_val                                                                                     ( hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit1_rst_val),
   .hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit2_rst_val                                                                                     ( hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit2_rst_val),
   .hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit3_rst_val                                                                                     ( hssi_pldadapt_tx_0_fsr_hip_fsr_out_bit3_rst_val),
   .hssi_pldadapt_tx_0_fsr_mask_tx_pll_rst_val                                                                                          ( hssi_pldadapt_tx_0_fsr_mask_tx_pll_rst_val),
   .hssi_pldadapt_tx_0_fsr_pld_txelecidle_rst_val                                                                                       ( hssi_pldadapt_tx_0_fsr_pld_txelecidle_rst_val),
   .hssi_pldadapt_tx_0_gb_tx_idwidth                                                                                                    ( hssi_pldadapt_tx_0_gb_tx_idwidth),
   .hssi_pldadapt_tx_0_gb_tx_odwidth                                                                                                    ( hssi_pldadapt_tx_0_gb_tx_odwidth),
   .hssi_pldadapt_tx_0_hip_mode                                                                                                         ( hssi_pldadapt_tx_0_hip_mode),
   .hssi_pldadapt_tx_0_hip_osc_clk_scg_en                                                                                               ( hssi_pldadapt_tx_0_hip_osc_clk_scg_en),
   .hssi_pldadapt_tx_0_hrdrst_dcd_cal_done_bypass                                                                                       ( hssi_pldadapt_tx_0_hrdrst_dcd_cal_done_bypass),
   .hssi_pldadapt_tx_0_hrdrst_rst_sm_dis                                                                                                ( hssi_pldadapt_tx_0_hrdrst_rst_sm_dis),
   .hssi_pldadapt_tx_0_hrdrst_rx_osc_clk_scg_en                                                                                         ( hssi_pldadapt_tx_0_hrdrst_rx_osc_clk_scg_en),
   .hssi_pldadapt_tx_0_hrdrst_user_ctl_en                                                                                               ( hssi_pldadapt_tx_0_hrdrst_user_ctl_en),
   .hssi_pldadapt_tx_0_indv                                                                                                             ( hssi_pldadapt_tx_0_indv),
   .hssi_pldadapt_tx_0_is_paired_with                                                                                                   ( hssi_pldadapt_tx_0_is_paired_with),
   .hssi_pldadapt_tx_0_loopback_mode                                                                                                    ( hssi_pldadapt_tx_0_loopback_mode),
   .hssi_pldadapt_tx_0_low_latency_en                                                                                                   ( hssi_pldadapt_tx_0_low_latency_en),
   .hssi_pldadapt_tx_0_osc_clk_scg_en                                                                                                   ( hssi_pldadapt_tx_0_osc_clk_scg_en),
   .hssi_pldadapt_tx_0_phcomp_rd_del                                                                                                    ( hssi_pldadapt_tx_0_phcomp_rd_del),
   .hssi_pldadapt_tx_0_pipe_mode                                                                                                        ( hssi_pldadapt_tx_0_pipe_mode),
   .hssi_pldadapt_tx_0_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                               ( hssi_pldadapt_tx_0_hdpldadapt_pld_avmm1_clk_rowclk_hz),
   .hssi_pldadapt_tx_0_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                               ( hssi_pldadapt_tx_0_hdpldadapt_pld_avmm2_clk_rowclk_hz),
   .hssi_pldadapt_tx_0_pld_clk1_delay_en                                                                                                ( hssi_pldadapt_tx_0_pld_clk1_delay_en),
   .hssi_pldadapt_tx_0_pld_clk1_delay_sel                                                                                               ( hssi_pldadapt_tx_0_pld_clk1_delay_sel),
   .hssi_pldadapt_tx_0_pld_clk1_inv_en                                                                                                  ( hssi_pldadapt_tx_0_pld_clk1_inv_en),
   .hssi_pldadapt_tx_0_pld_clk1_sel                                                                                                     ( hssi_pldadapt_tx_0_pld_clk1_sel),
   .hssi_pldadapt_tx_0_pld_clk2_sel                                                                                                     ( hssi_pldadapt_tx_0_pld_clk2_sel),
   .hssi_pldadapt_tx_0_hdpldadapt_pld_sclk1_rowclk_hz                                                                                   ( hssi_pldadapt_tx_0_hdpldadapt_pld_sclk1_rowclk_hz),
   .hssi_pldadapt_tx_0_hdpldadapt_pld_sclk2_rowclk_hz                                                                                   ( hssi_pldadapt_tx_0_hdpldadapt_pld_sclk2_rowclk_hz),
   .hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk1_dcm_hz                                                                                    ( hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk1_dcm_hz),
   .hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk1_rowclk_hz                                                                                 ( hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk1_rowclk_hz),
   .hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk2_dcm_hz                                                                                    ( hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk2_dcm_hz),
   .hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk2_rowclk_hz                                                                                 ( hssi_pldadapt_tx_0_hdpldadapt_pld_tx_clk2_rowclk_hz),
   .hssi_pldadapt_tx_0_pma_aib_tx_clk_expected_setting                                                                                  ( hssi_pldadapt_tx_0_pma_aib_tx_clk_expected_setting),
   .hssi_pldadapt_tx_0_powerdown_mode                                                                                                   ( hssi_pldadapt_tx_0_powerdown_mode),
   .hssi_pldadapt_tx_0_powermode_dc                                                                                                     ( hssi_pldadapt_tx_0_powermode_dc),
   .hssi_pldadapt_tx_0_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                        ( hssi_pldadapt_tx_0_powermode_freq_hz_aib_fabric_rx_sr_clk_in),
   .hssi_pldadapt_tx_0_powermode_freq_hz_pld_tx_clk1_dcm                                                                                ( hssi_pldadapt_tx_0_powermode_freq_hz_pld_tx_clk1_dcm),
   .hssi_pldadapt_tx_0_sh_err                                                                                                           ( hssi_pldadapt_tx_0_sh_err),
   .hssi_pldadapt_tx_0_hdpldadapt_speed_grade                                                                                           ( hssi_pldadapt_tx_0_hdpldadapt_speed_grade),
   .hssi_pldadapt_tx_0_hdpldadapt_sr_sr_testbus_sel                                                                                     ( hssi_pldadapt_tx_0_hdpldadapt_sr_sr_testbus_sel),
   .hssi_pldadapt_tx_0_stretch_num_stages                                                                                               ( hssi_pldadapt_tx_0_stretch_num_stages),
   .hssi_pldadapt_tx_0_sup_mode                                                                                                         ( hssi_pldadapt_tx_0_sup_mode),
   .hssi_pldadapt_tx_0_tx_datapath_tb_sel                                                                                               ( hssi_pldadapt_tx_0_tx_datapath_tb_sel),
   .hssi_pldadapt_tx_0_tx_fastbond_rden                                                                                                 ( hssi_pldadapt_tx_0_tx_fastbond_rden),
   .hssi_pldadapt_tx_0_tx_fastbond_wren                                                                                                 ( hssi_pldadapt_tx_0_tx_fastbond_wren),
   .hssi_pldadapt_tx_0_tx_fifo_power_mode                                                                                               ( hssi_pldadapt_tx_0_tx_fifo_power_mode),
   .hssi_pldadapt_tx_0_tx_fifo_read_latency_adjust                                                                                      ( hssi_pldadapt_tx_0_tx_fifo_read_latency_adjust),
   .hssi_pldadapt_tx_0_tx_fifo_write_latency_adjust                                                                                     ( hssi_pldadapt_tx_0_tx_fifo_write_latency_adjust),
   .hssi_pldadapt_tx_0_tx_hip_aib_ssr_in_polling_bypass                                                                                 ( hssi_pldadapt_tx_0_tx_hip_aib_ssr_in_polling_bypass),
   .hssi_pldadapt_tx_0_tx_osc_clock_setting                                                                                             ( hssi_pldadapt_tx_0_tx_osc_clock_setting),
   .hssi_pldadapt_tx_0_tx_pld_10g_tx_bitslip_polling_bypass                                                                             ( hssi_pldadapt_tx_0_tx_pld_10g_tx_bitslip_polling_bypass),
   .hssi_pldadapt_tx_0_tx_pld_8g_tx_boundary_sel_polling_bypass                                                                         ( hssi_pldadapt_tx_0_tx_pld_8g_tx_boundary_sel_polling_bypass),
   .hssi_pldadapt_tx_0_tx_pld_pma_fpll_cnt_sel_polling_bypass                                                                           ( hssi_pldadapt_tx_0_tx_pld_pma_fpll_cnt_sel_polling_bypass),
   .hssi_pldadapt_tx_0_tx_pld_pma_fpll_num_phase_shifts_polling_bypass                                                                  ( hssi_pldadapt_tx_0_tx_pld_pma_fpll_num_phase_shifts_polling_bypass),
   .hssi_pldadapt_tx_0_tx_usertest_sel                                                                                                  ( hssi_pldadapt_tx_0_tx_usertest_sel),
   .hssi_pldadapt_tx_0_txfifo_empty                                                                                                     ( hssi_pldadapt_tx_0_txfifo_empty),
   .hssi_pldadapt_tx_0_txfifo_full                                                                                                      ( hssi_pldadapt_tx_0_txfifo_full),
   .hssi_pldadapt_tx_0_txfifo_mode                                                                                                      ( hssi_pldadapt_tx_0_txfifo_mode),
   .hssi_pldadapt_tx_0_txfifo_pempty                                                                                                    ( hssi_pldadapt_tx_0_txfifo_pempty),
   .hssi_pldadapt_tx_0_txfifo_pfull                                                                                                     ( hssi_pldadapt_tx_0_txfifo_pfull),
   .hssi_pldadapt_tx_0_us_bypass_pipeln                                                                                                 ( hssi_pldadapt_tx_0_us_bypass_pipeln),
   .hssi_pldadapt_tx_0_us_last_chnl                                                                                                     ( hssi_pldadapt_tx_0_us_last_chnl),
   .hssi_pldadapt_tx_0_us_master                                                                                                        ( hssi_pldadapt_tx_0_us_master),
   .hssi_pldadapt_tx_0_word_align_enable                                                                                                ( hssi_pldadapt_tx_0_word_align_enable),
   .hssi_pldadapt_tx_0_word_mark                                                                                                        ( hssi_pldadapt_tx_0_word_mark),
   .hssi_pldadapt_tx_0_silicon_rev                                                                                                      ( hssi_pldadapt_tx_0_silicon_rev),
   .hssi_pldadapt_tx_0_reconfig_settings                                                                                                ( hssi_pldadapt_tx_0_reconfig_settings),
   .hssi_pldadapt_rx_0_aib_clk1_sel                                                                                                     ( hssi_pldadapt_rx_0_aib_clk1_sel),
   .hssi_pldadapt_rx_0_aib_clk2_sel                                                                                                     ( hssi_pldadapt_rx_0_aib_clk2_sel),
   .hssi_pldadapt_rx_0_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                            ( hssi_pldadapt_rx_0_hdpldadapt_aib_fabric_pld_pma_hclk_hz),
   .hssi_pldadapt_rx_0_hdpldadapt_aib_fabric_rx_sr_clk_in_hz                                                                            ( hssi_pldadapt_rx_0_hdpldadapt_aib_fabric_rx_sr_clk_in_hz),
   .hssi_pldadapt_rx_0_hdpldadapt_aib_fabric_rx_transfer_clk_hz                                                                         ( hssi_pldadapt_rx_0_hdpldadapt_aib_fabric_rx_transfer_clk_hz),
   .hssi_pldadapt_rx_0_asn_bypass_pma_pcie_sw_done                                                                                      ( hssi_pldadapt_rx_0_asn_bypass_pma_pcie_sw_done),
   .hssi_pldadapt_rx_0_asn_en                                                                                                           ( hssi_pldadapt_rx_0_asn_en),
   .hssi_pldadapt_rx_0_asn_wait_for_dll_reset_cnt                                                                                       ( hssi_pldadapt_rx_0_asn_wait_for_dll_reset_cnt),
   .hssi_pldadapt_rx_0_asn_wait_for_fifo_flush_cnt                                                                                      ( hssi_pldadapt_rx_0_asn_wait_for_fifo_flush_cnt),
   .hssi_pldadapt_rx_0_asn_wait_for_pma_pcie_sw_done_cnt                                                                                ( hssi_pldadapt_rx_0_asn_wait_for_pma_pcie_sw_done_cnt),
   .hssi_pldadapt_rx_0_bonding_dft_en                                                                                                   ( hssi_pldadapt_rx_0_bonding_dft_en),
   .hssi_pldadapt_rx_0_bonding_dft_val                                                                                                  ( hssi_pldadapt_rx_0_bonding_dft_val),
   .hssi_pldadapt_rx_0_chnl_bonding                                                                                                     ( hssi_pldadapt_rx_0_chnl_bonding),
   .hssi_pldadapt_rx_0_clock_del_measure_enable                                                                                         ( hssi_pldadapt_rx_0_clock_del_measure_enable),
   .hssi_pldadapt_rx_0_comp_cnt                                                                                                         ( hssi_pldadapt_rx_0_comp_cnt),
   .hssi_pldadapt_rx_0_compin_sel                                                                                                       ( hssi_pldadapt_rx_0_compin_sel),
   .hssi_pldadapt_rx_0_hdpldadapt_csr_clk_hz                                                                                            ( hssi_pldadapt_rx_0_hdpldadapt_csr_clk_hz),
   .hssi_pldadapt_rx_0_ctrl_plane_bonding                                                                                               ( hssi_pldadapt_rx_0_ctrl_plane_bonding),
   .hssi_pldadapt_rx_0_ds_bypass_pipeln                                                                                                 ( hssi_pldadapt_rx_0_ds_bypass_pipeln),
   .hssi_pldadapt_rx_0_ds_last_chnl                                                                                                     ( hssi_pldadapt_rx_0_ds_last_chnl),
   .hssi_pldadapt_rx_0_ds_master                                                                                                        ( hssi_pldadapt_rx_0_ds_master),
   .hssi_pldadapt_rx_0_duplex_mode                                                                                                      ( hssi_pldadapt_rx_0_duplex_mode),
   .hssi_pldadapt_rx_0_dv_mode                                                                                                          ( hssi_pldadapt_rx_0_dv_mode),
   .hssi_pldadapt_rx_0_fifo_double_read                                                                                                 ( hssi_pldadapt_rx_0_fifo_double_read),
   .hssi_pldadapt_rx_0_fifo_mode                                                                                                        ( hssi_pldadapt_rx_0_fifo_mode),
   .hssi_pldadapt_rx_0_fifo_rd_clk_ins_sm_scg_en                                                                                        ( hssi_pldadapt_rx_0_fifo_rd_clk_ins_sm_scg_en),
   .hssi_pldadapt_rx_0_fifo_rd_clk_scg_en                                                                                               ( hssi_pldadapt_rx_0_fifo_rd_clk_scg_en),
   .hssi_pldadapt_rx_0_fifo_rd_clk_sel                                                                                                  ( hssi_pldadapt_rx_0_fifo_rd_clk_sel),
   .hssi_pldadapt_rx_0_fifo_stop_rd                                                                                                     ( hssi_pldadapt_rx_0_fifo_stop_rd),
   .hssi_pldadapt_rx_0_fifo_stop_wr                                                                                                     ( hssi_pldadapt_rx_0_fifo_stop_wr),
   .hssi_pldadapt_rx_0_fifo_width                                                                                                       ( hssi_pldadapt_rx_0_fifo_width),
   .hssi_pldadapt_rx_0_fifo_wr_clk_del_sm_scg_en                                                                                        ( hssi_pldadapt_rx_0_fifo_wr_clk_del_sm_scg_en),
   .hssi_pldadapt_rx_0_fifo_wr_clk_scg_en                                                                                               ( hssi_pldadapt_rx_0_fifo_wr_clk_scg_en),
   .hssi_pldadapt_rx_0_fifo_wr_clk_sel                                                                                                  ( hssi_pldadapt_rx_0_fifo_wr_clk_sel),
   .hssi_pldadapt_rx_0_free_run_div_clk                                                                                                 ( hssi_pldadapt_rx_0_free_run_div_clk),
   .hssi_pldadapt_rx_0_fsr_pld_10g_rx_crc32_err_rst_val                                                                                 ( hssi_pldadapt_rx_0_fsr_pld_10g_rx_crc32_err_rst_val),
   .hssi_pldadapt_rx_0_fsr_pld_8g_sigdet_out_rst_val                                                                                    ( hssi_pldadapt_rx_0_fsr_pld_8g_sigdet_out_rst_val),
   .hssi_pldadapt_rx_0_fsr_pld_ltd_b_rst_val                                                                                            ( hssi_pldadapt_rx_0_fsr_pld_ltd_b_rst_val),
   .hssi_pldadapt_rx_0_fsr_pld_ltr_rst_val                                                                                              ( hssi_pldadapt_rx_0_fsr_pld_ltr_rst_val),
   .hssi_pldadapt_rx_0_fsr_pld_rx_fifo_align_clr_rst_val                                                                                ( hssi_pldadapt_rx_0_fsr_pld_rx_fifo_align_clr_rst_val),
   .hssi_pldadapt_rx_0_gb_rx_idwidth                                                                                                    ( hssi_pldadapt_rx_0_gb_rx_idwidth),
   .hssi_pldadapt_rx_0_gb_rx_odwidth                                                                                                    ( hssi_pldadapt_rx_0_gb_rx_odwidth),
   .hssi_pldadapt_rx_0_hip_mode                                                                                                         ( hssi_pldadapt_rx_0_hip_mode),
   .hssi_pldadapt_rx_0_hrdrst_align_bypass                                                                                              ( hssi_pldadapt_rx_0_hrdrst_align_bypass),
   .hssi_pldadapt_rx_0_hrdrst_dll_lock_bypass                                                                                           ( hssi_pldadapt_rx_0_hrdrst_dll_lock_bypass),
   .hssi_pldadapt_rx_0_hrdrst_rst_sm_dis                                                                                                ( hssi_pldadapt_rx_0_hrdrst_rst_sm_dis),
   .hssi_pldadapt_rx_0_hrdrst_rx_osc_clk_scg_en                                                                                         ( hssi_pldadapt_rx_0_hrdrst_rx_osc_clk_scg_en),
   .hssi_pldadapt_rx_0_hrdrst_user_ctl_en                                                                                               ( hssi_pldadapt_rx_0_hrdrst_user_ctl_en),
   .hssi_pldadapt_rx_0_indv                                                                                                             ( hssi_pldadapt_rx_0_indv),
   .hssi_pldadapt_rx_0_internal_clk1_sel1                                                                                               ( hssi_pldadapt_rx_0_internal_clk1_sel1),
   .hssi_pldadapt_rx_0_internal_clk1_sel2                                                                                               ( hssi_pldadapt_rx_0_internal_clk1_sel2),
   .hssi_pldadapt_rx_0_internal_clk2_sel1                                                                                               ( hssi_pldadapt_rx_0_internal_clk2_sel1),
   .hssi_pldadapt_rx_0_internal_clk2_sel2                                                                                               ( hssi_pldadapt_rx_0_internal_clk2_sel2),
   .hssi_pldadapt_rx_0_is_paired_with                                                                                                   ( hssi_pldadapt_rx_0_is_paired_with),
   .hssi_pldadapt_rx_0_loopback_mode                                                                                                    ( hssi_pldadapt_rx_0_loopback_mode),
   .hssi_pldadapt_rx_0_low_latency_en                                                                                                   ( hssi_pldadapt_rx_0_low_latency_en),
   .hssi_pldadapt_rx_0_lpbk_mode                                                                                                        ( hssi_pldadapt_rx_0_lpbk_mode),
   .hssi_pldadapt_rx_0_osc_clk_scg_en                                                                                                   ( hssi_pldadapt_rx_0_osc_clk_scg_en),
   .hssi_pldadapt_rx_0_phcomp_rd_del                                                                                                    ( hssi_pldadapt_rx_0_phcomp_rd_del),
   .hssi_pldadapt_rx_0_pipe_enable                                                                                                      ( hssi_pldadapt_rx_0_pipe_enable),
   .hssi_pldadapt_rx_0_pipe_mode                                                                                                        ( hssi_pldadapt_rx_0_pipe_mode),
   .hssi_pldadapt_rx_0_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                               ( hssi_pldadapt_rx_0_hdpldadapt_pld_avmm1_clk_rowclk_hz),
   .hssi_pldadapt_rx_0_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                               ( hssi_pldadapt_rx_0_hdpldadapt_pld_avmm2_clk_rowclk_hz),
   .hssi_pldadapt_rx_0_pld_clk1_delay_en                                                                                                ( hssi_pldadapt_rx_0_pld_clk1_delay_en),
   .hssi_pldadapt_rx_0_pld_clk1_delay_sel                                                                                               ( hssi_pldadapt_rx_0_pld_clk1_delay_sel),
   .hssi_pldadapt_rx_0_pld_clk1_inv_en                                                                                                  ( hssi_pldadapt_rx_0_pld_clk1_inv_en),
   .hssi_pldadapt_rx_0_pld_clk1_sel                                                                                                     ( hssi_pldadapt_rx_0_pld_clk1_sel),
   .hssi_pldadapt_rx_0_hdpldadapt_pld_rx_clk1_dcm_hz                                                                                    ( hssi_pldadapt_rx_0_hdpldadapt_pld_rx_clk1_dcm_hz),
   .hssi_pldadapt_rx_0_hdpldadapt_pld_rx_clk1_rowclk_hz                                                                                 ( hssi_pldadapt_rx_0_hdpldadapt_pld_rx_clk1_rowclk_hz),
   .hssi_pldadapt_rx_0_hdpldadapt_pld_sclk1_rowclk_hz                                                                                   ( hssi_pldadapt_rx_0_hdpldadapt_pld_sclk1_rowclk_hz),
   .hssi_pldadapt_rx_0_hdpldadapt_pld_sclk2_rowclk_hz                                                                                   ( hssi_pldadapt_rx_0_hdpldadapt_pld_sclk2_rowclk_hz),
   .hssi_pldadapt_rx_0_pma_hclk_scg_en                                                                                                  ( hssi_pldadapt_rx_0_pma_hclk_scg_en),
   .hssi_pldadapt_rx_0_powerdown_mode                                                                                                   ( hssi_pldadapt_rx_0_powerdown_mode),
   .hssi_pldadapt_rx_0_powermode_dc                                                                                                     ( hssi_pldadapt_rx_0_powermode_dc),
   .hssi_pldadapt_rx_0_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                        ( hssi_pldadapt_rx_0_powermode_freq_hz_aib_fabric_rx_sr_clk_in),
   .hssi_pldadapt_rx_0_powermode_freq_hz_pld_rx_clk1_dcm                                                                                ( hssi_pldadapt_rx_0_powermode_freq_hz_pld_rx_clk1_dcm),
   .hssi_pldadapt_rx_0_rx_datapath_tb_sel                                                                                               ( hssi_pldadapt_rx_0_rx_datapath_tb_sel),
   .hssi_pldadapt_rx_0_rx_fastbond_rden                                                                                                 ( hssi_pldadapt_rx_0_rx_fastbond_rden),
   .hssi_pldadapt_rx_0_rx_fastbond_wren                                                                                                 ( hssi_pldadapt_rx_0_rx_fastbond_wren),
   .hssi_pldadapt_rx_0_rx_fifo_power_mode                                                                                               ( hssi_pldadapt_rx_0_rx_fifo_power_mode),
   .hssi_pldadapt_rx_0_rx_fifo_read_latency_adjust                                                                                      ( hssi_pldadapt_rx_0_rx_fifo_read_latency_adjust),
   .hssi_pldadapt_rx_0_rx_fifo_write_ctrl                                                                                               ( hssi_pldadapt_rx_0_rx_fifo_write_ctrl),
   .hssi_pldadapt_rx_0_rx_fifo_write_latency_adjust                                                                                     ( hssi_pldadapt_rx_0_rx_fifo_write_latency_adjust),
   .hssi_pldadapt_rx_0_rx_osc_clock_setting                                                                                             ( hssi_pldadapt_rx_0_rx_osc_clock_setting),
   .hssi_pldadapt_rx_0_rx_pld_8g_eidleinfersel_polling_bypass                                                                           ( hssi_pldadapt_rx_0_rx_pld_8g_eidleinfersel_polling_bypass),
   .hssi_pldadapt_rx_0_rx_pld_pma_eye_monitor_polling_bypass                                                                            ( hssi_pldadapt_rx_0_rx_pld_pma_eye_monitor_polling_bypass),
   .hssi_pldadapt_rx_0_rx_pld_pma_pcie_switch_polling_bypass                                                                            ( hssi_pldadapt_rx_0_rx_pld_pma_pcie_switch_polling_bypass),
   .hssi_pldadapt_rx_0_rx_pld_pma_reser_out_polling_bypass                                                                              ( hssi_pldadapt_rx_0_rx_pld_pma_reser_out_polling_bypass),
   .hssi_pldadapt_rx_0_rx_prbs_flags_sr_enable                                                                                          ( hssi_pldadapt_rx_0_rx_prbs_flags_sr_enable),
   .hssi_pldadapt_rx_0_rx_true_b2b                                                                                                      ( hssi_pldadapt_rx_0_rx_true_b2b),
   .hssi_pldadapt_rx_0_rx_usertest_sel                                                                                                  ( hssi_pldadapt_rx_0_rx_usertest_sel),
   .hssi_pldadapt_rx_0_rxfifo_empty                                                                                                     ( hssi_pldadapt_rx_0_rxfifo_empty),
   .hssi_pldadapt_rx_0_rxfifo_full                                                                                                      ( hssi_pldadapt_rx_0_rxfifo_full),
   .hssi_pldadapt_rx_0_rxfifo_mode                                                                                                      ( hssi_pldadapt_rx_0_rxfifo_mode),
   .hssi_pldadapt_rx_0_rxfifo_pempty                                                                                                    ( hssi_pldadapt_rx_0_rxfifo_pempty),
   .hssi_pldadapt_rx_0_rxfifo_pfull                                                                                                     ( hssi_pldadapt_rx_0_rxfifo_pfull),
   .hssi_pldadapt_rx_0_rxfiford_post_ct_sel                                                                                             ( hssi_pldadapt_rx_0_rxfiford_post_ct_sel),
   .hssi_pldadapt_rx_0_rxfifowr_post_ct_sel                                                                                             ( hssi_pldadapt_rx_0_rxfifowr_post_ct_sel),
   .hssi_pldadapt_rx_0_sclk_sel                                                                                                         ( hssi_pldadapt_rx_0_sclk_sel),
   .hssi_pldadapt_rx_0_hdpldadapt_speed_grade                                                                                           ( hssi_pldadapt_rx_0_hdpldadapt_speed_grade),
   .hssi_pldadapt_rx_0_hdpldadapt_sr_sr_testbus_sel                                                                                     ( hssi_pldadapt_rx_0_hdpldadapt_sr_sr_testbus_sel),
   .hssi_pldadapt_rx_0_stretch_num_stages                                                                                               ( hssi_pldadapt_rx_0_stretch_num_stages),
   .hssi_pldadapt_rx_0_sup_mode                                                                                                         ( hssi_pldadapt_rx_0_sup_mode),
   .hssi_pldadapt_rx_0_txfiford_post_ct_sel                                                                                             ( hssi_pldadapt_rx_0_txfiford_post_ct_sel),
   .hssi_pldadapt_rx_0_txfifowr_post_ct_sel                                                                                             ( hssi_pldadapt_rx_0_txfifowr_post_ct_sel),
   .hssi_pldadapt_rx_0_us_bypass_pipeln                                                                                                 ( hssi_pldadapt_rx_0_us_bypass_pipeln),
   .hssi_pldadapt_rx_0_us_last_chnl                                                                                                     ( hssi_pldadapt_rx_0_us_last_chnl),
   .hssi_pldadapt_rx_0_us_master                                                                                                        ( hssi_pldadapt_rx_0_us_master),
   .hssi_pldadapt_rx_0_word_align                                                                                                       ( hssi_pldadapt_rx_0_word_align),
   .hssi_pldadapt_rx_0_word_align_enable                                                                                                ( hssi_pldadapt_rx_0_word_align_enable),
   .hssi_pldadapt_rx_0_silicon_rev                                                                                                      ( hssi_pldadapt_rx_0_silicon_rev),
   .hssi_pldadapt_rx_0_reconfig_settings                                                                                                ( hssi_pldadapt_rx_0_reconfig_settings),
   .hssi_avmm1_if_0_pcs_arbiter_ctrl                                                                                                    ( hssi_avmm1_if_0_pcs_arbiter_ctrl),
   .hssi_avmm1_if_0_hssiadapt_avmm_clk_dcg_en                                                                                           ( hssi_avmm1_if_0_hssiadapt_avmm_clk_dcg_en),
   .hssi_avmm1_if_0_hssiadapt_avmm_clk_scg_en                                                                                           ( hssi_avmm1_if_0_hssiadapt_avmm_clk_scg_en),
   .hssi_avmm1_if_0_pldadapt_avmm_clk_scg_en                                                                                            ( hssi_avmm1_if_0_pldadapt_avmm_clk_scg_en),
   .hssi_avmm1_if_0_pcs_cal_done                                                                                                        ( hssi_avmm1_if_0_pcs_cal_done),
   .hssi_avmm1_if_0_pcs_cal_reserved                                                                                                    ( hssi_avmm1_if_0_pcs_cal_reserved),
   .hssi_avmm1_if_0_pcs_calibration_feature_en                                                                                          ( hssi_avmm1_if_0_pcs_calibration_feature_en),
   .hssi_avmm1_if_0_pldadapt_gate_dis                                                                                                   ( hssi_avmm1_if_0_pldadapt_gate_dis),
   .hssi_avmm1_if_0_pcs_hip_cal_en                                                                                                      ( hssi_avmm1_if_0_pcs_hip_cal_en),
   .hssi_avmm1_if_0_hssiadapt_nfhssi_calibratio_feature_en                                                                              ( hssi_avmm1_if_0_hssiadapt_nfhssi_calibratio_feature_en),
   .hssi_avmm1_if_0_pldadapt_nfhssi_calibratio_feature_en                                                                               ( hssi_avmm1_if_0_pldadapt_nfhssi_calibratio_feature_en),
   .hssi_avmm1_if_0_hssiadapt_osc_clk_scg_en                                                                                            ( hssi_avmm1_if_0_hssiadapt_osc_clk_scg_en),
   .hssi_avmm1_if_0_pldadapt_osc_clk_scg_en                                                                                             ( hssi_avmm1_if_0_pldadapt_osc_clk_scg_en),
   .hssi_avmm1_if_0_hssiadapt_read_blocking_enable                                                                                      ( hssi_avmm1_if_0_hssiadapt_read_blocking_enable),
   .hssi_avmm1_if_0_pldadapt_read_blocking_enable                                                                                       ( hssi_avmm1_if_0_pldadapt_read_blocking_enable),
   .hssi_avmm1_if_0_hssiadapt_uc_blocking_enable                                                                                        ( hssi_avmm1_if_0_hssiadapt_uc_blocking_enable),
   .hssi_avmm1_if_0_pldadapt_uc_blocking_enable                                                                                         ( hssi_avmm1_if_0_pldadapt_uc_blocking_enable),
   .hssi_avmm1_if_0_hssiadapt_write_resp_en                                                                                             ( hssi_avmm1_if_0_hssiadapt_write_resp_en),
   .hssi_avmm1_if_0_hssiadapt_avmm_osc_clock_setting                                                                                    ( hssi_avmm1_if_0_hssiadapt_avmm_osc_clock_setting),
   .hssi_avmm1_if_0_pldadapt_avmm_osc_clock_setting                                                                                     ( hssi_avmm1_if_0_pldadapt_avmm_osc_clock_setting),
   .hssi_avmm1_if_0_hssiadapt_avmm_testbus_sel                                                                                          ( hssi_avmm1_if_0_hssiadapt_avmm_testbus_sel),
   .hssi_avmm1_if_0_pldadapt_avmm_testbus_sel                                                                                           ( hssi_avmm1_if_0_pldadapt_avmm_testbus_sel),
   .hssi_avmm1_if_0_func_mode                                                                                                           ( hssi_avmm1_if_0_func_mode),
   .hssi_avmm1_if_0_hssiadapt_sr_hip_mode                                                                                               ( hssi_avmm1_if_0_hssiadapt_sr_hip_mode),
   .hssi_avmm1_if_0_hssiadapt_hip_mode                                                                                                  ( hssi_avmm1_if_0_hssiadapt_hip_mode),
   .hssi_avmm1_if_0_pldadapt_hip_mode                                                                                                   ( hssi_avmm1_if_0_pldadapt_hip_mode),
   .hssi_avmm1_if_0_hssiadapt_sr_powerdown_mode                                                                                         ( hssi_avmm1_if_0_hssiadapt_sr_powerdown_mode),
   .hssi_avmm1_if_0_hssiadapt_sr_sr_free_run_div_clk                                                                                    ( hssi_avmm1_if_0_hssiadapt_sr_sr_free_run_div_clk),
   .hssi_avmm1_if_0_hssiadapt_sr_sr_hip_en                                                                                              ( hssi_avmm1_if_0_hssiadapt_sr_sr_hip_en),
   .hssi_avmm1_if_0_hssiadapt_sr_sr_osc_clk_div_sel                                                                                     ( hssi_avmm1_if_0_hssiadapt_sr_sr_osc_clk_div_sel),
   .hssi_avmm1_if_0_hssiadapt_sr_sr_osc_clk_scg_en                                                                                      ( hssi_avmm1_if_0_hssiadapt_sr_sr_osc_clk_scg_en),
   .hssi_avmm1_if_0_hssiadapt_sr_sr_parity_en                                                                                           ( hssi_avmm1_if_0_hssiadapt_sr_sr_parity_en),
   .hssi_avmm1_if_0_hssiadapt_sr_sr_reserved_in_en                                                                                      ( hssi_avmm1_if_0_hssiadapt_sr_sr_reserved_in_en),
   .hssi_avmm1_if_0_hssiadapt_sr_sr_reserved_out_en                                                                                     ( hssi_avmm1_if_0_hssiadapt_sr_sr_reserved_out_en),
   .hssi_avmm1_if_0_hssiadapt_sr_sup_mode                                                                                               ( hssi_avmm1_if_0_hssiadapt_sr_sup_mode),
   .hssi_avmm1_if_0_topology                                                                                                            ( hssi_avmm1_if_0_topology),
   .hssi_avmm1_if_0_silicon_rev                                                                                                         ( hssi_avmm1_if_0_silicon_rev),
   .hssi_avmm1_if_0_calibration_type                                                                                                    ( hssi_avmm1_if_0_calibration_type),
   .hssi_avmm2_if_0_pcs_arbiter_ctrl                                                                                                    ( hssi_avmm2_if_0_pcs_arbiter_ctrl),
   .hssi_avmm2_if_0_hssiadapt_avmm_clk_dcg_en                                                                                           ( hssi_avmm2_if_0_hssiadapt_avmm_clk_dcg_en),
   .hssi_avmm2_if_0_hssiadapt_avmm_clk_scg_en                                                                                           ( hssi_avmm2_if_0_hssiadapt_avmm_clk_scg_en),
   .hssi_avmm2_if_0_pldadapt_avmm_clk_scg_en                                                                                            ( hssi_avmm2_if_0_pldadapt_avmm_clk_scg_en),
   .hssi_avmm2_if_0_pcs_cal_done                                                                                                        ( hssi_avmm2_if_0_pcs_cal_done),
   .hssi_avmm2_if_0_pcs_cal_reserved                                                                                                    ( hssi_avmm2_if_0_pcs_cal_reserved),
   .hssi_avmm2_if_0_pcs_calibration_feature_en                                                                                          ( hssi_avmm2_if_0_pcs_calibration_feature_en),
   .hssi_avmm2_if_0_pldadapt_gate_dis                                                                                                   ( hssi_avmm2_if_0_pldadapt_gate_dis),
   .hssi_avmm2_if_0_pcs_hip_cal_en                                                                                                      ( hssi_avmm2_if_0_pcs_hip_cal_en),
   .hssi_avmm2_if_0_hssiadapt_osc_clk_scg_en                                                                                            ( hssi_avmm2_if_0_hssiadapt_osc_clk_scg_en),
   .hssi_avmm2_if_0_pldadapt_osc_clk_scg_en                                                                                             ( hssi_avmm2_if_0_pldadapt_osc_clk_scg_en),
   .hssi_avmm2_if_0_hssiadapt_avmm_osc_clock_setting                                                                                    ( hssi_avmm2_if_0_hssiadapt_avmm_osc_clock_setting),
   .hssi_avmm2_if_0_pldadapt_avmm_osc_clock_setting                                                                                     ( hssi_avmm2_if_0_pldadapt_avmm_osc_clock_setting),
   .hssi_avmm2_if_0_hssiadapt_avmm_testbus_sel                                                                                          ( hssi_avmm2_if_0_hssiadapt_avmm_testbus_sel),
   .hssi_avmm2_if_0_pldadapt_avmm_testbus_sel                                                                                           ( hssi_avmm2_if_0_pldadapt_avmm_testbus_sel),
   .hssi_avmm2_if_0_func_mode                                                                                                           ( hssi_avmm2_if_0_func_mode),
   .hssi_avmm2_if_0_hssiadapt_hip_mode                                                                                                  ( hssi_avmm2_if_0_hssiadapt_hip_mode),
   .hssi_avmm2_if_0_pldadapt_hip_mode                                                                                                   ( hssi_avmm2_if_0_pldadapt_hip_mode),
   .hssi_avmm2_if_0_topology                                                                                                            ( hssi_avmm2_if_0_topology),
   .hssi_avmm2_if_0_silicon_rev                                                                                                         ( hssi_avmm2_if_0_silicon_rev),
   .hssi_avmm2_if_0_calibration_type                                                                                                    ( hssi_avmm2_if_0_calibration_type),
   .hssi_aibnd_rx_13_aib_ber_margining_ctrl                                                                                             ( hssi_aibnd_rx_13_aib_ber_margining_ctrl),
   .hssi_aibnd_rx_13_aib_datasel_gr0                                                                                                    ( hssi_aibnd_rx_13_aib_datasel_gr0),
   .hssi_aibnd_rx_13_aib_datasel_gr1                                                                                                    ( hssi_aibnd_rx_13_aib_datasel_gr1),
   .hssi_aibnd_rx_13_aib_datasel_gr2                                                                                                    ( hssi_aibnd_rx_13_aib_datasel_gr2),
   .hssi_aibnd_rx_13_aib_dllstr_align_clkdiv                                                                                            ( hssi_aibnd_rx_13_aib_dllstr_align_clkdiv),
   .hssi_aibnd_rx_13_aib_dllstr_align_dly_pst                                                                                           ( hssi_aibnd_rx_13_aib_dllstr_align_dly_pst),
   .hssi_aibnd_rx_13_aib_dllstr_align_dy_ctl_static                                                                                     ( hssi_aibnd_rx_13_aib_dllstr_align_dy_ctl_static),
   .hssi_aibnd_rx_13_aib_dllstr_align_dy_ctlsel                                                                                         ( hssi_aibnd_rx_13_aib_dllstr_align_dy_ctlsel),
   .hssi_aibnd_rx_13_aib_dllstr_align_entest                                                                                            ( hssi_aibnd_rx_13_aib_dllstr_align_entest),
   .hssi_aibnd_rx_13_aib_dllstr_align_halfcode                                                                                          ( hssi_aibnd_rx_13_aib_dllstr_align_halfcode),
   .hssi_aibnd_rx_13_aib_dllstr_align_selflock                                                                                          ( hssi_aibnd_rx_13_aib_dllstr_align_selflock),
   .hssi_aibnd_rx_13_aib_dllstr_align_st_core_dn_prgmnvrt                                                                               ( hssi_aibnd_rx_13_aib_dllstr_align_st_core_dn_prgmnvrt),
   .hssi_aibnd_rx_13_aib_dllstr_align_st_core_up_prgmnvrt                                                                               ( hssi_aibnd_rx_13_aib_dllstr_align_st_core_up_prgmnvrt),
   .hssi_aibnd_rx_13_aib_dllstr_align_st_core_updnen                                                                                    ( hssi_aibnd_rx_13_aib_dllstr_align_st_core_updnen),
   .hssi_aibnd_rx_13_aib_dllstr_align_st_dftmuxsel                                                                                      ( hssi_aibnd_rx_13_aib_dllstr_align_st_dftmuxsel),
   .hssi_aibnd_rx_13_aib_dllstr_align_st_en                                                                                             ( hssi_aibnd_rx_13_aib_dllstr_align_st_en),
   .hssi_aibnd_rx_13_aib_dllstr_align_st_hps_ctrl_en                                                                                    ( hssi_aibnd_rx_13_aib_dllstr_align_st_hps_ctrl_en),
   .hssi_aibnd_rx_13_aib_dllstr_align_st_lockreq_muxsel                                                                                 ( hssi_aibnd_rx_13_aib_dllstr_align_st_lockreq_muxsel),
   .hssi_aibnd_rx_13_aib_dllstr_align_st_new_dll                                                                                        ( hssi_aibnd_rx_13_aib_dllstr_align_st_new_dll),
   .hssi_aibnd_rx_13_aib_dllstr_align_st_rst                                                                                            ( hssi_aibnd_rx_13_aib_dllstr_align_st_rst),
   .hssi_aibnd_rx_13_aib_dllstr_align_st_rst_prgmnvrt                                                                                   ( hssi_aibnd_rx_13_aib_dllstr_align_st_rst_prgmnvrt),
   .hssi_aibnd_rx_13_aib_dllstr_align_test_clk_pll_en_n                                                                                 ( hssi_aibnd_rx_13_aib_dllstr_align_test_clk_pll_en_n),
   .hssi_aibnd_rx_13_aib_inctrl_gr0                                                                                                     ( hssi_aibnd_rx_13_aib_inctrl_gr0),
   .hssi_aibnd_rx_13_aib_inctrl_gr1                                                                                                     ( hssi_aibnd_rx_13_aib_inctrl_gr1),
   .hssi_aibnd_rx_13_aib_inctrl_gr2                                                                                                     ( hssi_aibnd_rx_13_aib_inctrl_gr2),
   .hssi_aibnd_rx_13_aib_inctrl_gr3                                                                                                     ( hssi_aibnd_rx_13_aib_inctrl_gr3),
   .hssi_aibnd_rx_13_aib_outctrl_gr0                                                                                                    ( hssi_aibnd_rx_13_aib_outctrl_gr0),
   .hssi_aibnd_rx_13_aib_outctrl_gr1                                                                                                    ( hssi_aibnd_rx_13_aib_outctrl_gr1),
   .hssi_aibnd_rx_13_aib_outctrl_gr2                                                                                                    ( hssi_aibnd_rx_13_aib_outctrl_gr2),
   .hssi_aibnd_rx_13_aib_outndrv_r12                                                                                                    ( hssi_aibnd_rx_13_aib_outndrv_r12),
   .hssi_aibnd_rx_13_aib_outndrv_r34                                                                                                    ( hssi_aibnd_rx_13_aib_outndrv_r34),
   .hssi_aibnd_rx_13_aib_outndrv_r56                                                                                                    ( hssi_aibnd_rx_13_aib_outndrv_r56),
   .hssi_aibnd_rx_13_aib_outndrv_r78                                                                                                    ( hssi_aibnd_rx_13_aib_outndrv_r78),
   .hssi_aibnd_rx_13_aib_outpdrv_r12                                                                                                    ( hssi_aibnd_rx_13_aib_outpdrv_r12),
   .hssi_aibnd_rx_13_aib_outpdrv_r34                                                                                                    ( hssi_aibnd_rx_13_aib_outpdrv_r34),
   .hssi_aibnd_rx_13_aib_outpdrv_r56                                                                                                    ( hssi_aibnd_rx_13_aib_outpdrv_r56),
   .hssi_aibnd_rx_13_aib_outpdrv_r78                                                                                                    ( hssi_aibnd_rx_13_aib_outpdrv_r78),
   .hssi_aibnd_rx_13_aib_red_shift_en                                                                                                   ( hssi_aibnd_rx_13_aib_red_shift_en),
   .hssi_aibnd_rx_13_dft_hssitestip_dll_dcc_en                                                                                          ( hssi_aibnd_rx_13_dft_hssitestip_dll_dcc_en),
   .hssi_aibnd_rx_13_op_mode                                                                                                            ( hssi_aibnd_rx_13_op_mode),
   .hssi_aibnd_rx_13_powerdown_mode                                                                                                     ( hssi_aibnd_rx_13_powerdown_mode),
   .hssi_aibnd_rx_13_powermode_ac                                                                                                       ( hssi_aibnd_rx_13_powermode_ac),
   .hssi_aibnd_rx_13_powermode_dc                                                                                                       ( hssi_aibnd_rx_13_powermode_dc),
   .hssi_aibnd_rx_13_powermode_freq_hz_aib_hssi_rx_transfer_clk                                                                         ( hssi_aibnd_rx_13_powermode_freq_hz_aib_hssi_rx_transfer_clk),
   .hssi_aibnd_rx_13_redundancy_en                                                                                                      ( hssi_aibnd_rx_13_redundancy_en),
   .hssi_aibnd_rx_13_sup_mode                                                                                                           ( hssi_aibnd_rx_13_sup_mode),
   .hssi_aibnd_rx_13_silicon_rev                                                                                                        ( hssi_aibnd_rx_13_silicon_rev),
   .hssi_aibnd_tx_13_aib_datasel_gr0                                                                                                    ( hssi_aibnd_tx_13_aib_datasel_gr0),
   .hssi_aibnd_tx_13_aib_datasel_gr1                                                                                                    ( hssi_aibnd_tx_13_aib_datasel_gr1),
   .hssi_aibnd_tx_13_aib_datasel_gr2                                                                                                    ( hssi_aibnd_tx_13_aib_datasel_gr2),
   .hssi_aibnd_tx_13_aib_datasel_gr3                                                                                                    ( hssi_aibnd_tx_13_aib_datasel_gr3),
   .hssi_aibnd_tx_13_aib_ddrctrl_gr0                                                                                                    ( hssi_aibnd_tx_13_aib_ddrctrl_gr0),
   .hssi_aibnd_tx_13_aib_hssi_tx_transfer_clk_hz                                                                                        ( hssi_aibnd_tx_13_aib_hssi_tx_transfer_clk_hz),
   .hssi_aibnd_tx_13_aib_iinasyncen                                                                                                     ( hssi_aibnd_tx_13_aib_iinasyncen),
   .hssi_aibnd_tx_13_aib_iinclken                                                                                                       ( hssi_aibnd_tx_13_aib_iinclken),
   .hssi_aibnd_tx_13_aib_outctrl_gr0                                                                                                    ( hssi_aibnd_tx_13_aib_outctrl_gr0),
   .hssi_aibnd_tx_13_aib_outctrl_gr1                                                                                                    ( hssi_aibnd_tx_13_aib_outctrl_gr1),
   .hssi_aibnd_tx_13_aib_outctrl_gr2                                                                                                    ( hssi_aibnd_tx_13_aib_outctrl_gr2),
   .hssi_aibnd_tx_13_aib_outctrl_gr3                                                                                                    ( hssi_aibnd_tx_13_aib_outctrl_gr3),
   .hssi_aibnd_tx_13_aib_outndrv_r34                                                                                                    ( hssi_aibnd_tx_13_aib_outndrv_r34),
   .hssi_aibnd_tx_13_aib_outndrv_r56                                                                                                    ( hssi_aibnd_tx_13_aib_outndrv_r56),
   .hssi_aibnd_tx_13_aib_outpdrv_r34                                                                                                    ( hssi_aibnd_tx_13_aib_outpdrv_r34),
   .hssi_aibnd_tx_13_aib_outpdrv_r56                                                                                                    ( hssi_aibnd_tx_13_aib_outpdrv_r56),
   .hssi_aibnd_tx_13_aib_red_dirclkn_shiften                                                                                            ( hssi_aibnd_tx_13_aib_red_dirclkn_shiften),
   .hssi_aibnd_tx_13_aib_red_dirclkp_shiften                                                                                            ( hssi_aibnd_tx_13_aib_red_dirclkp_shiften),
   .hssi_aibnd_tx_13_aib_red_drx_shiften                                                                                                ( hssi_aibnd_tx_13_aib_red_drx_shiften),
   .hssi_aibnd_tx_13_aib_red_dtx_shiften                                                                                                ( hssi_aibnd_tx_13_aib_red_dtx_shiften),
   .hssi_aibnd_tx_13_aib_red_pout_shiften                                                                                               ( hssi_aibnd_tx_13_aib_red_pout_shiften),
   .hssi_aibnd_tx_13_aib_red_rx_shiften                                                                                                 ( hssi_aibnd_tx_13_aib_red_rx_shiften),
   .hssi_aibnd_tx_13_aib_red_tx_shiften                                                                                                 ( hssi_aibnd_tx_13_aib_red_tx_shiften),
   .hssi_aibnd_tx_13_aib_red_txferclkout_shiften                                                                                        ( hssi_aibnd_tx_13_aib_red_txferclkout_shiften),
   .hssi_aibnd_tx_13_aib_red_txferclkoutn_shiften                                                                                       ( hssi_aibnd_tx_13_aib_red_txferclkoutn_shiften),
   .hssi_aibnd_tx_13_aib_tx_clkdiv                                                                                                      ( hssi_aibnd_tx_13_aib_tx_clkdiv),
   .hssi_aibnd_tx_13_aib_tx_dcc_byp                                                                                                     ( hssi_aibnd_tx_13_aib_tx_dcc_byp),
   .hssi_aibnd_tx_13_aib_tx_dcc_byp_iocsr_unused                                                                                        ( hssi_aibnd_tx_13_aib_tx_dcc_byp_iocsr_unused),
   .hssi_aibnd_tx_13_aib_tx_dcc_cont_cal                                                                                                ( hssi_aibnd_tx_13_aib_tx_dcc_cont_cal),
   .hssi_aibnd_tx_13_aib_tx_dcc_cont_cal_iocsr_unused                                                                                   ( hssi_aibnd_tx_13_aib_tx_dcc_cont_cal_iocsr_unused),
   .hssi_aibnd_tx_13_aib_tx_dcc_dft                                                                                                     ( hssi_aibnd_tx_13_aib_tx_dcc_dft),
   .hssi_aibnd_tx_13_aib_tx_dcc_dft_sel                                                                                                 ( hssi_aibnd_tx_13_aib_tx_dcc_dft_sel),
   .hssi_aibnd_tx_13_aib_tx_dcc_dll_dft_sel                                                                                             ( hssi_aibnd_tx_13_aib_tx_dcc_dll_dft_sel),
   .hssi_aibnd_tx_13_aib_tx_dcc_dll_entest                                                                                              ( hssi_aibnd_tx_13_aib_tx_dcc_dll_entest),
   .hssi_aibnd_tx_13_aib_tx_dcc_dy_ctl_static                                                                                           ( hssi_aibnd_tx_13_aib_tx_dcc_dy_ctl_static),
   .hssi_aibnd_tx_13_aib_tx_dcc_dy_ctlsel                                                                                               ( hssi_aibnd_tx_13_aib_tx_dcc_dy_ctlsel),
   .hssi_aibnd_tx_13_aib_tx_dcc_en                                                                                                      ( hssi_aibnd_tx_13_aib_tx_dcc_en),
   .hssi_aibnd_tx_13_aib_tx_dcc_en_iocsr_unused                                                                                         ( hssi_aibnd_tx_13_aib_tx_dcc_en_iocsr_unused),
   .hssi_aibnd_tx_13_aib_tx_dcc_manual_dn                                                                                               ( hssi_aibnd_tx_13_aib_tx_dcc_manual_dn),
   .hssi_aibnd_tx_13_aib_tx_dcc_manual_up                                                                                               ( hssi_aibnd_tx_13_aib_tx_dcc_manual_up),
   .hssi_aibnd_tx_13_aib_tx_dcc_rst_prgmnvrt                                                                                            ( hssi_aibnd_tx_13_aib_tx_dcc_rst_prgmnvrt),
   .hssi_aibnd_tx_13_aib_tx_dcc_st_core_dn_prgmnvrt                                                                                     ( hssi_aibnd_tx_13_aib_tx_dcc_st_core_dn_prgmnvrt),
   .hssi_aibnd_tx_13_aib_tx_dcc_st_core_up_prgmnvrt                                                                                     ( hssi_aibnd_tx_13_aib_tx_dcc_st_core_up_prgmnvrt),
   .hssi_aibnd_tx_13_aib_tx_dcc_st_core_updnen                                                                                          ( hssi_aibnd_tx_13_aib_tx_dcc_st_core_updnen),
   .hssi_aibnd_tx_13_aib_tx_dcc_st_dftmuxsel                                                                                            ( hssi_aibnd_tx_13_aib_tx_dcc_st_dftmuxsel),
   .hssi_aibnd_tx_13_aib_tx_dcc_st_dly_pst                                                                                              ( hssi_aibnd_tx_13_aib_tx_dcc_st_dly_pst),
   .hssi_aibnd_tx_13_aib_tx_dcc_st_en                                                                                                   ( hssi_aibnd_tx_13_aib_tx_dcc_st_en),
   .hssi_aibnd_tx_13_aib_tx_dcc_st_hps_ctrl_en                                                                                          ( hssi_aibnd_tx_13_aib_tx_dcc_st_hps_ctrl_en),
   .hssi_aibnd_tx_13_aib_tx_dcc_st_lockreq_muxsel                                                                                       ( hssi_aibnd_tx_13_aib_tx_dcc_st_lockreq_muxsel),
   .hssi_aibnd_tx_13_aib_tx_dcc_st_new_dll                                                                                              ( hssi_aibnd_tx_13_aib_tx_dcc_st_new_dll),
   .hssi_aibnd_tx_13_aib_tx_dcc_st_rst                                                                                                  ( hssi_aibnd_tx_13_aib_tx_dcc_st_rst),
   .hssi_aibnd_tx_13_aib_tx_dcc_test_clk_pll_en_n                                                                                       ( hssi_aibnd_tx_13_aib_tx_dcc_test_clk_pll_en_n),
   .hssi_aibnd_tx_13_aib_tx_halfcode                                                                                                    ( hssi_aibnd_tx_13_aib_tx_halfcode),
   .hssi_aibnd_tx_13_aib_tx_selflock                                                                                                    ( hssi_aibnd_tx_13_aib_tx_selflock),
   .hssi_aibnd_tx_13_dfd_dll_dcc_en                                                                                                     ( hssi_aibnd_tx_13_dfd_dll_dcc_en),
   .hssi_aibnd_tx_13_dft_hssitestip_dll_dcc_en                                                                                          ( hssi_aibnd_tx_13_dft_hssitestip_dll_dcc_en),
   .hssi_aibnd_tx_13_op_mode                                                                                                            ( hssi_aibnd_tx_13_op_mode),
   .hssi_aibnd_tx_13_powerdown_mode                                                                                                     ( hssi_aibnd_tx_13_powerdown_mode),
   .hssi_aibnd_tx_13_powermode_ac                                                                                                       ( hssi_aibnd_tx_13_powermode_ac),
   .hssi_aibnd_tx_13_powermode_dc                                                                                                       ( hssi_aibnd_tx_13_powermode_dc),
   .hssi_aibnd_tx_13_powermode_freq_hz_aib_hssi_tx_transfer_clk                                                                         ( hssi_aibnd_tx_13_powermode_freq_hz_aib_hssi_tx_transfer_clk),
   .hssi_aibnd_tx_13_redundancy_en                                                                                                      ( hssi_aibnd_tx_13_redundancy_en),
   .hssi_aibnd_tx_13_sup_mode                                                                                                           ( hssi_aibnd_tx_13_sup_mode),
   .hssi_aibnd_tx_13_silicon_rev                                                                                                        ( hssi_aibnd_tx_13_silicon_rev),
   .hssi_pldadapt_tx_13_aib_clk1_sel                                                                                                    ( hssi_pldadapt_tx_13_aib_clk1_sel),
   .hssi_pldadapt_tx_13_aib_clk2_sel                                                                                                    ( hssi_pldadapt_tx_13_aib_clk2_sel),
   .hssi_pldadapt_tx_13_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                           ( hssi_pldadapt_tx_13_hdpldadapt_aib_fabric_pld_pma_hclk_hz),
   .hssi_pldadapt_tx_13_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz                                                                         ( hssi_pldadapt_tx_13_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz),
   .hssi_pldadapt_tx_13_hdpldadapt_aib_fabric_tx_sr_clk_in_hz                                                                           ( hssi_pldadapt_tx_13_hdpldadapt_aib_fabric_tx_sr_clk_in_hz),
   .hssi_pldadapt_tx_13_bonding_dft_en                                                                                                  ( hssi_pldadapt_tx_13_bonding_dft_en),
   .hssi_pldadapt_tx_13_bonding_dft_val                                                                                                 ( hssi_pldadapt_tx_13_bonding_dft_val),
   .hssi_pldadapt_tx_13_chnl_bonding                                                                                                    ( hssi_pldadapt_tx_13_chnl_bonding),
   .hssi_pldadapt_tx_13_comp_cnt                                                                                                        ( hssi_pldadapt_tx_13_comp_cnt),
   .hssi_pldadapt_tx_13_compin_sel                                                                                                      ( hssi_pldadapt_tx_13_compin_sel),
   .hssi_pldadapt_tx_13_hdpldadapt_csr_clk_hz                                                                                           ( hssi_pldadapt_tx_13_hdpldadapt_csr_clk_hz),
   .hssi_pldadapt_tx_13_ctrl_plane_bonding                                                                                              ( hssi_pldadapt_tx_13_ctrl_plane_bonding),
   .hssi_pldadapt_tx_13_ds_bypass_pipeln                                                                                                ( hssi_pldadapt_tx_13_ds_bypass_pipeln),
   .hssi_pldadapt_tx_13_ds_last_chnl                                                                                                    ( hssi_pldadapt_tx_13_ds_last_chnl),
   .hssi_pldadapt_tx_13_ds_master                                                                                                       ( hssi_pldadapt_tx_13_ds_master),
   .hssi_pldadapt_tx_13_duplex_mode                                                                                                     ( hssi_pldadapt_tx_13_duplex_mode),
   .hssi_pldadapt_tx_13_dv_bond                                                                                                         ( hssi_pldadapt_tx_13_dv_bond),
   .hssi_pldadapt_tx_13_dv_gen                                                                                                          ( hssi_pldadapt_tx_13_dv_gen),
   .hssi_pldadapt_tx_13_fifo_double_write                                                                                               ( hssi_pldadapt_tx_13_fifo_double_write),
   .hssi_pldadapt_tx_13_fifo_mode                                                                                                       ( hssi_pldadapt_tx_13_fifo_mode),
   .hssi_pldadapt_tx_13_fifo_rd_clk_frm_gen_scg_en                                                                                      ( hssi_pldadapt_tx_13_fifo_rd_clk_frm_gen_scg_en),
   .hssi_pldadapt_tx_13_fifo_rd_clk_scg_en                                                                                              ( hssi_pldadapt_tx_13_fifo_rd_clk_scg_en),
   .hssi_pldadapt_tx_13_fifo_rd_clk_sel                                                                                                 ( hssi_pldadapt_tx_13_fifo_rd_clk_sel),
   .hssi_pldadapt_tx_13_fifo_stop_rd                                                                                                    ( hssi_pldadapt_tx_13_fifo_stop_rd),
   .hssi_pldadapt_tx_13_fifo_stop_wr                                                                                                    ( hssi_pldadapt_tx_13_fifo_stop_wr),
   .hssi_pldadapt_tx_13_fifo_width                                                                                                      ( hssi_pldadapt_tx_13_fifo_width),
   .hssi_pldadapt_tx_13_fifo_wr_clk_scg_en                                                                                              ( hssi_pldadapt_tx_13_fifo_wr_clk_scg_en),
   .hssi_pldadapt_tx_13_fpll_shared_direct_async_in_sel                                                                                 ( hssi_pldadapt_tx_13_fpll_shared_direct_async_in_sel),
   .hssi_pldadapt_tx_13_frmgen_burst                                                                                                    ( hssi_pldadapt_tx_13_frmgen_burst),
   .hssi_pldadapt_tx_13_frmgen_bypass                                                                                                   ( hssi_pldadapt_tx_13_frmgen_bypass),
   .hssi_pldadapt_tx_13_frmgen_mfrm_length                                                                                              ( hssi_pldadapt_tx_13_frmgen_mfrm_length),
   .hssi_pldadapt_tx_13_frmgen_pipeln                                                                                                   ( hssi_pldadapt_tx_13_frmgen_pipeln),
   .hssi_pldadapt_tx_13_frmgen_pyld_ins                                                                                                 ( hssi_pldadapt_tx_13_frmgen_pyld_ins),
   .hssi_pldadapt_tx_13_frmgen_wordslip                                                                                                 ( hssi_pldadapt_tx_13_frmgen_wordslip),
   .hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit0_rst_val                                                                                     ( hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit0_rst_val),
   .hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit1_rst_val                                                                                     ( hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit1_rst_val),
   .hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit2_rst_val                                                                                     ( hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit2_rst_val),
   .hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit3_rst_val                                                                                     ( hssi_pldadapt_tx_13_fsr_hip_fsr_in_bit3_rst_val),
   .hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit0_rst_val                                                                                    ( hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit0_rst_val),
   .hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit1_rst_val                                                                                    ( hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit1_rst_val),
   .hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit2_rst_val                                                                                    ( hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit2_rst_val),
   .hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit3_rst_val                                                                                    ( hssi_pldadapt_tx_13_fsr_hip_fsr_out_bit3_rst_val),
   .hssi_pldadapt_tx_13_fsr_mask_tx_pll_rst_val                                                                                         ( hssi_pldadapt_tx_13_fsr_mask_tx_pll_rst_val),
   .hssi_pldadapt_tx_13_fsr_pld_txelecidle_rst_val                                                                                      ( hssi_pldadapt_tx_13_fsr_pld_txelecidle_rst_val),
   .hssi_pldadapt_tx_13_gb_tx_idwidth                                                                                                   ( hssi_pldadapt_tx_13_gb_tx_idwidth),
   .hssi_pldadapt_tx_13_gb_tx_odwidth                                                                                                   ( hssi_pldadapt_tx_13_gb_tx_odwidth),
   .hssi_pldadapt_tx_13_hip_mode                                                                                                        ( hssi_pldadapt_tx_13_hip_mode),
   .hssi_pldadapt_tx_13_hip_osc_clk_scg_en                                                                                              ( hssi_pldadapt_tx_13_hip_osc_clk_scg_en),
   .hssi_pldadapt_tx_13_hrdrst_dcd_cal_done_bypass                                                                                      ( hssi_pldadapt_tx_13_hrdrst_dcd_cal_done_bypass),
   .hssi_pldadapt_tx_13_hrdrst_rst_sm_dis                                                                                               ( hssi_pldadapt_tx_13_hrdrst_rst_sm_dis),
   .hssi_pldadapt_tx_13_hrdrst_rx_osc_clk_scg_en                                                                                        ( hssi_pldadapt_tx_13_hrdrst_rx_osc_clk_scg_en),
   .hssi_pldadapt_tx_13_hrdrst_user_ctl_en                                                                                              ( hssi_pldadapt_tx_13_hrdrst_user_ctl_en),
   .hssi_pldadapt_tx_13_indv                                                                                                            ( hssi_pldadapt_tx_13_indv),
   .hssi_pldadapt_tx_13_is_paired_with                                                                                                  ( hssi_pldadapt_tx_13_is_paired_with),
   .hssi_pldadapt_tx_13_loopback_mode                                                                                                   ( hssi_pldadapt_tx_13_loopback_mode),
   .hssi_pldadapt_tx_13_low_latency_en                                                                                                  ( hssi_pldadapt_tx_13_low_latency_en),
   .hssi_pldadapt_tx_13_osc_clk_scg_en                                                                                                  ( hssi_pldadapt_tx_13_osc_clk_scg_en),
   .hssi_pldadapt_tx_13_phcomp_rd_del                                                                                                   ( hssi_pldadapt_tx_13_phcomp_rd_del),
   .hssi_pldadapt_tx_13_pipe_mode                                                                                                       ( hssi_pldadapt_tx_13_pipe_mode),
   .hssi_pldadapt_tx_13_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                              ( hssi_pldadapt_tx_13_hdpldadapt_pld_avmm1_clk_rowclk_hz),
   .hssi_pldadapt_tx_13_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                              ( hssi_pldadapt_tx_13_hdpldadapt_pld_avmm2_clk_rowclk_hz),
   .hssi_pldadapt_tx_13_pld_clk1_delay_en                                                                                               ( hssi_pldadapt_tx_13_pld_clk1_delay_en),
   .hssi_pldadapt_tx_13_pld_clk1_delay_sel                                                                                              ( hssi_pldadapt_tx_13_pld_clk1_delay_sel),
   .hssi_pldadapt_tx_13_pld_clk1_inv_en                                                                                                 ( hssi_pldadapt_tx_13_pld_clk1_inv_en),
   .hssi_pldadapt_tx_13_pld_clk1_sel                                                                                                    ( hssi_pldadapt_tx_13_pld_clk1_sel),
   .hssi_pldadapt_tx_13_pld_clk2_sel                                                                                                    ( hssi_pldadapt_tx_13_pld_clk2_sel),
   .hssi_pldadapt_tx_13_hdpldadapt_pld_sclk1_rowclk_hz                                                                                  ( hssi_pldadapt_tx_13_hdpldadapt_pld_sclk1_rowclk_hz),
   .hssi_pldadapt_tx_13_hdpldadapt_pld_sclk2_rowclk_hz                                                                                  ( hssi_pldadapt_tx_13_hdpldadapt_pld_sclk2_rowclk_hz),
   .hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk1_dcm_hz                                                                                   ( hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk1_dcm_hz),
   .hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk1_rowclk_hz                                                                                ( hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk1_rowclk_hz),
   .hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk2_dcm_hz                                                                                   ( hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk2_dcm_hz),
   .hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk2_rowclk_hz                                                                                ( hssi_pldadapt_tx_13_hdpldadapt_pld_tx_clk2_rowclk_hz),
   .hssi_pldadapt_tx_13_pma_aib_tx_clk_expected_setting                                                                                 ( hssi_pldadapt_tx_13_pma_aib_tx_clk_expected_setting),
   .hssi_pldadapt_tx_13_powerdown_mode                                                                                                  ( hssi_pldadapt_tx_13_powerdown_mode),
   .hssi_pldadapt_tx_13_powermode_dc                                                                                                    ( hssi_pldadapt_tx_13_powermode_dc),
   .hssi_pldadapt_tx_13_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                       ( hssi_pldadapt_tx_13_powermode_freq_hz_aib_fabric_rx_sr_clk_in),
   .hssi_pldadapt_tx_13_powermode_freq_hz_pld_tx_clk1_dcm                                                                               ( hssi_pldadapt_tx_13_powermode_freq_hz_pld_tx_clk1_dcm),
   .hssi_pldadapt_tx_13_sh_err                                                                                                          ( hssi_pldadapt_tx_13_sh_err),
   .hssi_pldadapt_tx_13_hdpldadapt_speed_grade                                                                                          ( hssi_pldadapt_tx_13_hdpldadapt_speed_grade),
   .hssi_pldadapt_tx_13_hdpldadapt_sr_sr_testbus_sel                                                                                    ( hssi_pldadapt_tx_13_hdpldadapt_sr_sr_testbus_sel),
   .hssi_pldadapt_tx_13_stretch_num_stages                                                                                              ( hssi_pldadapt_tx_13_stretch_num_stages),
   .hssi_pldadapt_tx_13_sup_mode                                                                                                        ( hssi_pldadapt_tx_13_sup_mode),
   .hssi_pldadapt_tx_13_tx_datapath_tb_sel                                                                                              ( hssi_pldadapt_tx_13_tx_datapath_tb_sel),
   .hssi_pldadapt_tx_13_tx_fastbond_rden                                                                                                ( hssi_pldadapt_tx_13_tx_fastbond_rden),
   .hssi_pldadapt_tx_13_tx_fastbond_wren                                                                                                ( hssi_pldadapt_tx_13_tx_fastbond_wren),
   .hssi_pldadapt_tx_13_tx_fifo_power_mode                                                                                              ( hssi_pldadapt_tx_13_tx_fifo_power_mode),
   .hssi_pldadapt_tx_13_tx_fifo_read_latency_adjust                                                                                     ( hssi_pldadapt_tx_13_tx_fifo_read_latency_adjust),
   .hssi_pldadapt_tx_13_tx_fifo_write_latency_adjust                                                                                    ( hssi_pldadapt_tx_13_tx_fifo_write_latency_adjust),
   .hssi_pldadapt_tx_13_tx_hip_aib_ssr_in_polling_bypass                                                                                ( hssi_pldadapt_tx_13_tx_hip_aib_ssr_in_polling_bypass),
   .hssi_pldadapt_tx_13_tx_osc_clock_setting                                                                                            ( hssi_pldadapt_tx_13_tx_osc_clock_setting),
   .hssi_pldadapt_tx_13_tx_pld_10g_tx_bitslip_polling_bypass                                                                            ( hssi_pldadapt_tx_13_tx_pld_10g_tx_bitslip_polling_bypass),
   .hssi_pldadapt_tx_13_tx_pld_8g_tx_boundary_sel_polling_bypass                                                                        ( hssi_pldadapt_tx_13_tx_pld_8g_tx_boundary_sel_polling_bypass),
   .hssi_pldadapt_tx_13_tx_pld_pma_fpll_cnt_sel_polling_bypass                                                                          ( hssi_pldadapt_tx_13_tx_pld_pma_fpll_cnt_sel_polling_bypass),
   .hssi_pldadapt_tx_13_tx_pld_pma_fpll_num_phase_shifts_polling_bypass                                                                 ( hssi_pldadapt_tx_13_tx_pld_pma_fpll_num_phase_shifts_polling_bypass),
   .hssi_pldadapt_tx_13_tx_usertest_sel                                                                                                 ( hssi_pldadapt_tx_13_tx_usertest_sel),
   .hssi_pldadapt_tx_13_txfifo_empty                                                                                                    ( hssi_pldadapt_tx_13_txfifo_empty),
   .hssi_pldadapt_tx_13_txfifo_full                                                                                                     ( hssi_pldadapt_tx_13_txfifo_full),
   .hssi_pldadapt_tx_13_txfifo_mode                                                                                                     ( hssi_pldadapt_tx_13_txfifo_mode),
   .hssi_pldadapt_tx_13_txfifo_pempty                                                                                                   ( hssi_pldadapt_tx_13_txfifo_pempty),
   .hssi_pldadapt_tx_13_txfifo_pfull                                                                                                    ( hssi_pldadapt_tx_13_txfifo_pfull),
   .hssi_pldadapt_tx_13_us_bypass_pipeln                                                                                                ( hssi_pldadapt_tx_13_us_bypass_pipeln),
   .hssi_pldadapt_tx_13_us_last_chnl                                                                                                    ( hssi_pldadapt_tx_13_us_last_chnl),
   .hssi_pldadapt_tx_13_us_master                                                                                                       ( hssi_pldadapt_tx_13_us_master),
   .hssi_pldadapt_tx_13_word_align_enable                                                                                               ( hssi_pldadapt_tx_13_word_align_enable),
   .hssi_pldadapt_tx_13_word_mark                                                                                                       ( hssi_pldadapt_tx_13_word_mark),
   .hssi_pldadapt_tx_13_silicon_rev                                                                                                     ( hssi_pldadapt_tx_13_silicon_rev),
   .hssi_pldadapt_tx_13_reconfig_settings                                                                                               ( hssi_pldadapt_tx_13_reconfig_settings),
   .hssi_pldadapt_rx_13_aib_clk1_sel                                                                                                    ( hssi_pldadapt_rx_13_aib_clk1_sel),
   .hssi_pldadapt_rx_13_aib_clk2_sel                                                                                                    ( hssi_pldadapt_rx_13_aib_clk2_sel),
   .hssi_pldadapt_rx_13_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                           ( hssi_pldadapt_rx_13_hdpldadapt_aib_fabric_pld_pma_hclk_hz),
   .hssi_pldadapt_rx_13_hdpldadapt_aib_fabric_rx_sr_clk_in_hz                                                                           ( hssi_pldadapt_rx_13_hdpldadapt_aib_fabric_rx_sr_clk_in_hz),
   .hssi_pldadapt_rx_13_hdpldadapt_aib_fabric_rx_transfer_clk_hz                                                                        ( hssi_pldadapt_rx_13_hdpldadapt_aib_fabric_rx_transfer_clk_hz),
   .hssi_pldadapt_rx_13_asn_bypass_pma_pcie_sw_done                                                                                     ( hssi_pldadapt_rx_13_asn_bypass_pma_pcie_sw_done),
   .hssi_pldadapt_rx_13_asn_en                                                                                                          ( hssi_pldadapt_rx_13_asn_en),
   .hssi_pldadapt_rx_13_asn_wait_for_dll_reset_cnt                                                                                      ( hssi_pldadapt_rx_13_asn_wait_for_dll_reset_cnt),
   .hssi_pldadapt_rx_13_asn_wait_for_fifo_flush_cnt                                                                                     ( hssi_pldadapt_rx_13_asn_wait_for_fifo_flush_cnt),
   .hssi_pldadapt_rx_13_asn_wait_for_pma_pcie_sw_done_cnt                                                                               ( hssi_pldadapt_rx_13_asn_wait_for_pma_pcie_sw_done_cnt),
   .hssi_pldadapt_rx_13_bonding_dft_en                                                                                                  ( hssi_pldadapt_rx_13_bonding_dft_en),
   .hssi_pldadapt_rx_13_bonding_dft_val                                                                                                 ( hssi_pldadapt_rx_13_bonding_dft_val),
   .hssi_pldadapt_rx_13_chnl_bonding                                                                                                    ( hssi_pldadapt_rx_13_chnl_bonding),
   .hssi_pldadapt_rx_13_clock_del_measure_enable                                                                                        ( hssi_pldadapt_rx_13_clock_del_measure_enable),
   .hssi_pldadapt_rx_13_comp_cnt                                                                                                        ( hssi_pldadapt_rx_13_comp_cnt),
   .hssi_pldadapt_rx_13_compin_sel                                                                                                      ( hssi_pldadapt_rx_13_compin_sel),
   .hssi_pldadapt_rx_13_hdpldadapt_csr_clk_hz                                                                                           ( hssi_pldadapt_rx_13_hdpldadapt_csr_clk_hz),
   .hssi_pldadapt_rx_13_ctrl_plane_bonding                                                                                              ( hssi_pldadapt_rx_13_ctrl_plane_bonding),
   .hssi_pldadapt_rx_13_ds_bypass_pipeln                                                                                                ( hssi_pldadapt_rx_13_ds_bypass_pipeln),
   .hssi_pldadapt_rx_13_ds_last_chnl                                                                                                    ( hssi_pldadapt_rx_13_ds_last_chnl),
   .hssi_pldadapt_rx_13_ds_master                                                                                                       ( hssi_pldadapt_rx_13_ds_master),
   .hssi_pldadapt_rx_13_duplex_mode                                                                                                     ( hssi_pldadapt_rx_13_duplex_mode),
   .hssi_pldadapt_rx_13_dv_mode                                                                                                         ( hssi_pldadapt_rx_13_dv_mode),
   .hssi_pldadapt_rx_13_fifo_double_read                                                                                                ( hssi_pldadapt_rx_13_fifo_double_read),
   .hssi_pldadapt_rx_13_fifo_mode                                                                                                       ( hssi_pldadapt_rx_13_fifo_mode),
   .hssi_pldadapt_rx_13_fifo_rd_clk_ins_sm_scg_en                                                                                       ( hssi_pldadapt_rx_13_fifo_rd_clk_ins_sm_scg_en),
   .hssi_pldadapt_rx_13_fifo_rd_clk_scg_en                                                                                              ( hssi_pldadapt_rx_13_fifo_rd_clk_scg_en),
   .hssi_pldadapt_rx_13_fifo_rd_clk_sel                                                                                                 ( hssi_pldadapt_rx_13_fifo_rd_clk_sel),
   .hssi_pldadapt_rx_13_fifo_stop_rd                                                                                                    ( hssi_pldadapt_rx_13_fifo_stop_rd),
   .hssi_pldadapt_rx_13_fifo_stop_wr                                                                                                    ( hssi_pldadapt_rx_13_fifo_stop_wr),
   .hssi_pldadapt_rx_13_fifo_width                                                                                                      ( hssi_pldadapt_rx_13_fifo_width),
   .hssi_pldadapt_rx_13_fifo_wr_clk_del_sm_scg_en                                                                                       ( hssi_pldadapt_rx_13_fifo_wr_clk_del_sm_scg_en),
   .hssi_pldadapt_rx_13_fifo_wr_clk_scg_en                                                                                              ( hssi_pldadapt_rx_13_fifo_wr_clk_scg_en),
   .hssi_pldadapt_rx_13_fifo_wr_clk_sel                                                                                                 ( hssi_pldadapt_rx_13_fifo_wr_clk_sel),
   .hssi_pldadapt_rx_13_free_run_div_clk                                                                                                ( hssi_pldadapt_rx_13_free_run_div_clk),
   .hssi_pldadapt_rx_13_fsr_pld_10g_rx_crc32_err_rst_val                                                                                ( hssi_pldadapt_rx_13_fsr_pld_10g_rx_crc32_err_rst_val),
   .hssi_pldadapt_rx_13_fsr_pld_8g_sigdet_out_rst_val                                                                                   ( hssi_pldadapt_rx_13_fsr_pld_8g_sigdet_out_rst_val),
   .hssi_pldadapt_rx_13_fsr_pld_ltd_b_rst_val                                                                                           ( hssi_pldadapt_rx_13_fsr_pld_ltd_b_rst_val),
   .hssi_pldadapt_rx_13_fsr_pld_ltr_rst_val                                                                                             ( hssi_pldadapt_rx_13_fsr_pld_ltr_rst_val),
   .hssi_pldadapt_rx_13_fsr_pld_rx_fifo_align_clr_rst_val                                                                               ( hssi_pldadapt_rx_13_fsr_pld_rx_fifo_align_clr_rst_val),
   .hssi_pldadapt_rx_13_gb_rx_idwidth                                                                                                   ( hssi_pldadapt_rx_13_gb_rx_idwidth),
   .hssi_pldadapt_rx_13_gb_rx_odwidth                                                                                                   ( hssi_pldadapt_rx_13_gb_rx_odwidth),
   .hssi_pldadapt_rx_13_hip_mode                                                                                                        ( hssi_pldadapt_rx_13_hip_mode),
   .hssi_pldadapt_rx_13_hrdrst_align_bypass                                                                                             ( hssi_pldadapt_rx_13_hrdrst_align_bypass),
   .hssi_pldadapt_rx_13_hrdrst_dll_lock_bypass                                                                                          ( hssi_pldadapt_rx_13_hrdrst_dll_lock_bypass),
   .hssi_pldadapt_rx_13_hrdrst_rst_sm_dis                                                                                               ( hssi_pldadapt_rx_13_hrdrst_rst_sm_dis),
   .hssi_pldadapt_rx_13_hrdrst_rx_osc_clk_scg_en                                                                                        ( hssi_pldadapt_rx_13_hrdrst_rx_osc_clk_scg_en),
   .hssi_pldadapt_rx_13_hrdrst_user_ctl_en                                                                                              ( hssi_pldadapt_rx_13_hrdrst_user_ctl_en),
   .hssi_pldadapt_rx_13_indv                                                                                                            ( hssi_pldadapt_rx_13_indv),
   .hssi_pldadapt_rx_13_internal_clk1_sel1                                                                                              ( hssi_pldadapt_rx_13_internal_clk1_sel1),
   .hssi_pldadapt_rx_13_internal_clk1_sel2                                                                                              ( hssi_pldadapt_rx_13_internal_clk1_sel2),
   .hssi_pldadapt_rx_13_internal_clk2_sel1                                                                                              ( hssi_pldadapt_rx_13_internal_clk2_sel1),
   .hssi_pldadapt_rx_13_internal_clk2_sel2                                                                                              ( hssi_pldadapt_rx_13_internal_clk2_sel2),
   .hssi_pldadapt_rx_13_is_paired_with                                                                                                  ( hssi_pldadapt_rx_13_is_paired_with),
   .hssi_pldadapt_rx_13_loopback_mode                                                                                                   ( hssi_pldadapt_rx_13_loopback_mode),
   .hssi_pldadapt_rx_13_low_latency_en                                                                                                  ( hssi_pldadapt_rx_13_low_latency_en),
   .hssi_pldadapt_rx_13_lpbk_mode                                                                                                       ( hssi_pldadapt_rx_13_lpbk_mode),
   .hssi_pldadapt_rx_13_osc_clk_scg_en                                                                                                  ( hssi_pldadapt_rx_13_osc_clk_scg_en),
   .hssi_pldadapt_rx_13_phcomp_rd_del                                                                                                   ( hssi_pldadapt_rx_13_phcomp_rd_del),
   .hssi_pldadapt_rx_13_pipe_enable                                                                                                     ( hssi_pldadapt_rx_13_pipe_enable),
   .hssi_pldadapt_rx_13_pipe_mode                                                                                                       ( hssi_pldadapt_rx_13_pipe_mode),
   .hssi_pldadapt_rx_13_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                              ( hssi_pldadapt_rx_13_hdpldadapt_pld_avmm1_clk_rowclk_hz),
   .hssi_pldadapt_rx_13_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                              ( hssi_pldadapt_rx_13_hdpldadapt_pld_avmm2_clk_rowclk_hz),
   .hssi_pldadapt_rx_13_pld_clk1_delay_en                                                                                               ( hssi_pldadapt_rx_13_pld_clk1_delay_en),
   .hssi_pldadapt_rx_13_pld_clk1_delay_sel                                                                                              ( hssi_pldadapt_rx_13_pld_clk1_delay_sel),
   .hssi_pldadapt_rx_13_pld_clk1_inv_en                                                                                                 ( hssi_pldadapt_rx_13_pld_clk1_inv_en),
   .hssi_pldadapt_rx_13_pld_clk1_sel                                                                                                    ( hssi_pldadapt_rx_13_pld_clk1_sel),
   .hssi_pldadapt_rx_13_hdpldadapt_pld_rx_clk1_dcm_hz                                                                                   ( hssi_pldadapt_rx_13_hdpldadapt_pld_rx_clk1_dcm_hz),
   .hssi_pldadapt_rx_13_hdpldadapt_pld_rx_clk1_rowclk_hz                                                                                ( hssi_pldadapt_rx_13_hdpldadapt_pld_rx_clk1_rowclk_hz),
   .hssi_pldadapt_rx_13_hdpldadapt_pld_sclk1_rowclk_hz                                                                                  ( hssi_pldadapt_rx_13_hdpldadapt_pld_sclk1_rowclk_hz),
   .hssi_pldadapt_rx_13_hdpldadapt_pld_sclk2_rowclk_hz                                                                                  ( hssi_pldadapt_rx_13_hdpldadapt_pld_sclk2_rowclk_hz),
   .hssi_pldadapt_rx_13_pma_hclk_scg_en                                                                                                 ( hssi_pldadapt_rx_13_pma_hclk_scg_en),
   .hssi_pldadapt_rx_13_powerdown_mode                                                                                                  ( hssi_pldadapt_rx_13_powerdown_mode),
   .hssi_pldadapt_rx_13_powermode_dc                                                                                                    ( hssi_pldadapt_rx_13_powermode_dc),
   .hssi_pldadapt_rx_13_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                       ( hssi_pldadapt_rx_13_powermode_freq_hz_aib_fabric_rx_sr_clk_in),
   .hssi_pldadapt_rx_13_powermode_freq_hz_pld_rx_clk1_dcm                                                                               ( hssi_pldadapt_rx_13_powermode_freq_hz_pld_rx_clk1_dcm),
   .hssi_pldadapt_rx_13_rx_datapath_tb_sel                                                                                              ( hssi_pldadapt_rx_13_rx_datapath_tb_sel),
   .hssi_pldadapt_rx_13_rx_fastbond_rden                                                                                                ( hssi_pldadapt_rx_13_rx_fastbond_rden),
   .hssi_pldadapt_rx_13_rx_fastbond_wren                                                                                                ( hssi_pldadapt_rx_13_rx_fastbond_wren),
   .hssi_pldadapt_rx_13_rx_fifo_power_mode                                                                                              ( hssi_pldadapt_rx_13_rx_fifo_power_mode),
   .hssi_pldadapt_rx_13_rx_fifo_read_latency_adjust                                                                                     ( hssi_pldadapt_rx_13_rx_fifo_read_latency_adjust),
   .hssi_pldadapt_rx_13_rx_fifo_write_ctrl                                                                                              ( hssi_pldadapt_rx_13_rx_fifo_write_ctrl),
   .hssi_pldadapt_rx_13_rx_fifo_write_latency_adjust                                                                                    ( hssi_pldadapt_rx_13_rx_fifo_write_latency_adjust),
   .hssi_pldadapt_rx_13_rx_osc_clock_setting                                                                                            ( hssi_pldadapt_rx_13_rx_osc_clock_setting),
   .hssi_pldadapt_rx_13_rx_pld_8g_eidleinfersel_polling_bypass                                                                          ( hssi_pldadapt_rx_13_rx_pld_8g_eidleinfersel_polling_bypass),
   .hssi_pldadapt_rx_13_rx_pld_pma_eye_monitor_polling_bypass                                                                           ( hssi_pldadapt_rx_13_rx_pld_pma_eye_monitor_polling_bypass),
   .hssi_pldadapt_rx_13_rx_pld_pma_pcie_switch_polling_bypass                                                                           ( hssi_pldadapt_rx_13_rx_pld_pma_pcie_switch_polling_bypass),
   .hssi_pldadapt_rx_13_rx_pld_pma_reser_out_polling_bypass                                                                             ( hssi_pldadapt_rx_13_rx_pld_pma_reser_out_polling_bypass),
   .hssi_pldadapt_rx_13_rx_prbs_flags_sr_enable                                                                                         ( hssi_pldadapt_rx_13_rx_prbs_flags_sr_enable),
   .hssi_pldadapt_rx_13_rx_true_b2b                                                                                                     ( hssi_pldadapt_rx_13_rx_true_b2b),
   .hssi_pldadapt_rx_13_rx_usertest_sel                                                                                                 ( hssi_pldadapt_rx_13_rx_usertest_sel),
   .hssi_pldadapt_rx_13_rxfifo_empty                                                                                                    ( hssi_pldadapt_rx_13_rxfifo_empty),
   .hssi_pldadapt_rx_13_rxfifo_full                                                                                                     ( hssi_pldadapt_rx_13_rxfifo_full),
   .hssi_pldadapt_rx_13_rxfifo_mode                                                                                                     ( hssi_pldadapt_rx_13_rxfifo_mode),
   .hssi_pldadapt_rx_13_rxfifo_pempty                                                                                                   ( hssi_pldadapt_rx_13_rxfifo_pempty),
   .hssi_pldadapt_rx_13_rxfifo_pfull                                                                                                    ( hssi_pldadapt_rx_13_rxfifo_pfull),
   .hssi_pldadapt_rx_13_rxfiford_post_ct_sel                                                                                            ( hssi_pldadapt_rx_13_rxfiford_post_ct_sel),
   .hssi_pldadapt_rx_13_rxfifowr_post_ct_sel                                                                                            ( hssi_pldadapt_rx_13_rxfifowr_post_ct_sel),
   .hssi_pldadapt_rx_13_sclk_sel                                                                                                        ( hssi_pldadapt_rx_13_sclk_sel),
   .hssi_pldadapt_rx_13_hdpldadapt_speed_grade                                                                                          ( hssi_pldadapt_rx_13_hdpldadapt_speed_grade),
   .hssi_pldadapt_rx_13_hdpldadapt_sr_sr_testbus_sel                                                                                    ( hssi_pldadapt_rx_13_hdpldadapt_sr_sr_testbus_sel),
   .hssi_pldadapt_rx_13_stretch_num_stages                                                                                              ( hssi_pldadapt_rx_13_stretch_num_stages),
   .hssi_pldadapt_rx_13_sup_mode                                                                                                        ( hssi_pldadapt_rx_13_sup_mode),
   .hssi_pldadapt_rx_13_txfiford_post_ct_sel                                                                                            ( hssi_pldadapt_rx_13_txfiford_post_ct_sel),
   .hssi_pldadapt_rx_13_txfifowr_post_ct_sel                                                                                            ( hssi_pldadapt_rx_13_txfifowr_post_ct_sel),
   .hssi_pldadapt_rx_13_us_bypass_pipeln                                                                                                ( hssi_pldadapt_rx_13_us_bypass_pipeln),
   .hssi_pldadapt_rx_13_us_last_chnl                                                                                                    ( hssi_pldadapt_rx_13_us_last_chnl),
   .hssi_pldadapt_rx_13_us_master                                                                                                       ( hssi_pldadapt_rx_13_us_master),
   .hssi_pldadapt_rx_13_word_align                                                                                                      ( hssi_pldadapt_rx_13_word_align),
   .hssi_pldadapt_rx_13_word_align_enable                                                                                               ( hssi_pldadapt_rx_13_word_align_enable),
   .hssi_pldadapt_rx_13_silicon_rev                                                                                                     ( hssi_pldadapt_rx_13_silicon_rev),
   .hssi_pldadapt_rx_13_reconfig_settings                                                                                               ( hssi_pldadapt_rx_13_reconfig_settings),
   .hssi_avmm1_if_13_pcs_arbiter_ctrl                                                                                                   ( hssi_avmm1_if_13_pcs_arbiter_ctrl),
   .hssi_avmm1_if_13_hssiadapt_avmm_clk_dcg_en                                                                                          ( hssi_avmm1_if_13_hssiadapt_avmm_clk_dcg_en),
   .hssi_avmm1_if_13_hssiadapt_avmm_clk_scg_en                                                                                          ( hssi_avmm1_if_13_hssiadapt_avmm_clk_scg_en),
   .hssi_avmm1_if_13_pldadapt_avmm_clk_scg_en                                                                                           ( hssi_avmm1_if_13_pldadapt_avmm_clk_scg_en),
   .hssi_avmm1_if_13_pcs_cal_done                                                                                                       ( hssi_avmm1_if_13_pcs_cal_done),
   .hssi_avmm1_if_13_pcs_cal_reserved                                                                                                   ( hssi_avmm1_if_13_pcs_cal_reserved),
   .hssi_avmm1_if_13_pcs_calibration_feature_en                                                                                         ( hssi_avmm1_if_13_pcs_calibration_feature_en),
   .hssi_avmm1_if_13_pldadapt_gate_dis                                                                                                  ( hssi_avmm1_if_13_pldadapt_gate_dis),
   .hssi_avmm1_if_13_pcs_hip_cal_en                                                                                                     ( hssi_avmm1_if_13_pcs_hip_cal_en),
   .hssi_avmm1_if_13_hssiadapt_nfhssi_calibratio_feature_en                                                                             ( hssi_avmm1_if_13_hssiadapt_nfhssi_calibratio_feature_en),
   .hssi_avmm1_if_13_pldadapt_nfhssi_calibratio_feature_en                                                                              ( hssi_avmm1_if_13_pldadapt_nfhssi_calibratio_feature_en),
   .hssi_avmm1_if_13_hssiadapt_osc_clk_scg_en                                                                                           ( hssi_avmm1_if_13_hssiadapt_osc_clk_scg_en),
   .hssi_avmm1_if_13_pldadapt_osc_clk_scg_en                                                                                            ( hssi_avmm1_if_13_pldadapt_osc_clk_scg_en),
   .hssi_avmm1_if_13_hssiadapt_read_blocking_enable                                                                                     ( hssi_avmm1_if_13_hssiadapt_read_blocking_enable),
   .hssi_avmm1_if_13_pldadapt_read_blocking_enable                                                                                      ( hssi_avmm1_if_13_pldadapt_read_blocking_enable),
   .hssi_avmm1_if_13_hssiadapt_uc_blocking_enable                                                                                       ( hssi_avmm1_if_13_hssiadapt_uc_blocking_enable),
   .hssi_avmm1_if_13_pldadapt_uc_blocking_enable                                                                                        ( hssi_avmm1_if_13_pldadapt_uc_blocking_enable),
   .hssi_avmm1_if_13_hssiadapt_write_resp_en                                                                                            ( hssi_avmm1_if_13_hssiadapt_write_resp_en),
   .hssi_avmm1_if_13_hssiadapt_avmm_osc_clock_setting                                                                                   ( hssi_avmm1_if_13_hssiadapt_avmm_osc_clock_setting),
   .hssi_avmm1_if_13_pldadapt_avmm_osc_clock_setting                                                                                    ( hssi_avmm1_if_13_pldadapt_avmm_osc_clock_setting),
   .hssi_avmm1_if_13_hssiadapt_avmm_testbus_sel                                                                                         ( hssi_avmm1_if_13_hssiadapt_avmm_testbus_sel),
   .hssi_avmm1_if_13_pldadapt_avmm_testbus_sel                                                                                          ( hssi_avmm1_if_13_pldadapt_avmm_testbus_sel),
   .hssi_avmm1_if_13_func_mode                                                                                                          ( hssi_avmm1_if_13_func_mode),
   .hssi_avmm1_if_13_hssiadapt_sr_hip_mode                                                                                              ( hssi_avmm1_if_13_hssiadapt_sr_hip_mode),
   .hssi_avmm1_if_13_hssiadapt_hip_mode                                                                                                 ( hssi_avmm1_if_13_hssiadapt_hip_mode),
   .hssi_avmm1_if_13_pldadapt_hip_mode                                                                                                  ( hssi_avmm1_if_13_pldadapt_hip_mode),
   .hssi_avmm1_if_13_hssiadapt_sr_powerdown_mode                                                                                        ( hssi_avmm1_if_13_hssiadapt_sr_powerdown_mode),
   .hssi_avmm1_if_13_hssiadapt_sr_sr_free_run_div_clk                                                                                   ( hssi_avmm1_if_13_hssiadapt_sr_sr_free_run_div_clk),
   .hssi_avmm1_if_13_hssiadapt_sr_sr_hip_en                                                                                             ( hssi_avmm1_if_13_hssiadapt_sr_sr_hip_en),
   .hssi_avmm1_if_13_hssiadapt_sr_sr_osc_clk_div_sel                                                                                    ( hssi_avmm1_if_13_hssiadapt_sr_sr_osc_clk_div_sel),
   .hssi_avmm1_if_13_hssiadapt_sr_sr_osc_clk_scg_en                                                                                     ( hssi_avmm1_if_13_hssiadapt_sr_sr_osc_clk_scg_en),
   .hssi_avmm1_if_13_hssiadapt_sr_sr_parity_en                                                                                          ( hssi_avmm1_if_13_hssiadapt_sr_sr_parity_en),
   .hssi_avmm1_if_13_hssiadapt_sr_sr_reserved_in_en                                                                                     ( hssi_avmm1_if_13_hssiadapt_sr_sr_reserved_in_en),
   .hssi_avmm1_if_13_hssiadapt_sr_sr_reserved_out_en                                                                                    ( hssi_avmm1_if_13_hssiadapt_sr_sr_reserved_out_en),
   .hssi_avmm1_if_13_hssiadapt_sr_sup_mode                                                                                              ( hssi_avmm1_if_13_hssiadapt_sr_sup_mode),
   .hssi_avmm1_if_13_topology                                                                                                           ( hssi_avmm1_if_13_topology),
   .hssi_avmm1_if_13_silicon_rev                                                                                                        ( hssi_avmm1_if_13_silicon_rev),
   .hssi_avmm1_if_13_calibration_type                                                                                                   ( hssi_avmm1_if_13_calibration_type),
   .hssi_avmm2_if_13_pcs_arbiter_ctrl                                                                                                   ( hssi_avmm2_if_13_pcs_arbiter_ctrl),
   .hssi_avmm2_if_13_hssiadapt_avmm_clk_dcg_en                                                                                          ( hssi_avmm2_if_13_hssiadapt_avmm_clk_dcg_en),
   .hssi_avmm2_if_13_hssiadapt_avmm_clk_scg_en                                                                                          ( hssi_avmm2_if_13_hssiadapt_avmm_clk_scg_en),
   .hssi_avmm2_if_13_pldadapt_avmm_clk_scg_en                                                                                           ( hssi_avmm2_if_13_pldadapt_avmm_clk_scg_en),
   .hssi_avmm2_if_13_pcs_cal_done                                                                                                       ( hssi_avmm2_if_13_pcs_cal_done),
   .hssi_avmm2_if_13_pcs_cal_reserved                                                                                                   ( hssi_avmm2_if_13_pcs_cal_reserved),
   .hssi_avmm2_if_13_pcs_calibration_feature_en                                                                                         ( hssi_avmm2_if_13_pcs_calibration_feature_en),
   .hssi_avmm2_if_13_pldadapt_gate_dis                                                                                                  ( hssi_avmm2_if_13_pldadapt_gate_dis),
   .hssi_avmm2_if_13_pcs_hip_cal_en                                                                                                     ( hssi_avmm2_if_13_pcs_hip_cal_en),
   .hssi_avmm2_if_13_hssiadapt_osc_clk_scg_en                                                                                           ( hssi_avmm2_if_13_hssiadapt_osc_clk_scg_en),
   .hssi_avmm2_if_13_pldadapt_osc_clk_scg_en                                                                                            ( hssi_avmm2_if_13_pldadapt_osc_clk_scg_en),
   .hssi_avmm2_if_13_hssiadapt_avmm_osc_clock_setting                                                                                   ( hssi_avmm2_if_13_hssiadapt_avmm_osc_clock_setting),
   .hssi_avmm2_if_13_pldadapt_avmm_osc_clock_setting                                                                                    ( hssi_avmm2_if_13_pldadapt_avmm_osc_clock_setting),
   .hssi_avmm2_if_13_hssiadapt_avmm_testbus_sel                                                                                         ( hssi_avmm2_if_13_hssiadapt_avmm_testbus_sel),
   .hssi_avmm2_if_13_pldadapt_avmm_testbus_sel                                                                                          ( hssi_avmm2_if_13_pldadapt_avmm_testbus_sel),
   .hssi_avmm2_if_13_func_mode                                                                                                          ( hssi_avmm2_if_13_func_mode),
   .hssi_avmm2_if_13_hssiadapt_hip_mode                                                                                                 ( hssi_avmm2_if_13_hssiadapt_hip_mode),
   .hssi_avmm2_if_13_pldadapt_hip_mode                                                                                                  ( hssi_avmm2_if_13_pldadapt_hip_mode),
   .hssi_avmm2_if_13_topology                                                                                                           ( hssi_avmm2_if_13_topology),
   .hssi_avmm2_if_13_silicon_rev                                                                                                        ( hssi_avmm2_if_13_silicon_rev),
   .hssi_avmm2_if_13_calibration_type                                                                                                   ( hssi_avmm2_if_13_calibration_type),
   .hssi_aibnd_rx_15_aib_ber_margining_ctrl                                                                                             ( hssi_aibnd_rx_15_aib_ber_margining_ctrl),
   .hssi_aibnd_rx_15_aib_datasel_gr0                                                                                                    ( hssi_aibnd_rx_15_aib_datasel_gr0),
   .hssi_aibnd_rx_15_aib_datasel_gr1                                                                                                    ( hssi_aibnd_rx_15_aib_datasel_gr1),
   .hssi_aibnd_rx_15_aib_datasel_gr2                                                                                                    ( hssi_aibnd_rx_15_aib_datasel_gr2),
   .hssi_aibnd_rx_15_aib_dllstr_align_clkdiv                                                                                            ( hssi_aibnd_rx_15_aib_dllstr_align_clkdiv),
   .hssi_aibnd_rx_15_aib_dllstr_align_dly_pst                                                                                           ( hssi_aibnd_rx_15_aib_dllstr_align_dly_pst),
   .hssi_aibnd_rx_15_aib_dllstr_align_dy_ctl_static                                                                                     ( hssi_aibnd_rx_15_aib_dllstr_align_dy_ctl_static),
   .hssi_aibnd_rx_15_aib_dllstr_align_dy_ctlsel                                                                                         ( hssi_aibnd_rx_15_aib_dllstr_align_dy_ctlsel),
   .hssi_aibnd_rx_15_aib_dllstr_align_entest                                                                                            ( hssi_aibnd_rx_15_aib_dllstr_align_entest),
   .hssi_aibnd_rx_15_aib_dllstr_align_halfcode                                                                                          ( hssi_aibnd_rx_15_aib_dllstr_align_halfcode),
   .hssi_aibnd_rx_15_aib_dllstr_align_selflock                                                                                          ( hssi_aibnd_rx_15_aib_dllstr_align_selflock),
   .hssi_aibnd_rx_15_aib_dllstr_align_st_core_dn_prgmnvrt                                                                               ( hssi_aibnd_rx_15_aib_dllstr_align_st_core_dn_prgmnvrt),
   .hssi_aibnd_rx_15_aib_dllstr_align_st_core_up_prgmnvrt                                                                               ( hssi_aibnd_rx_15_aib_dllstr_align_st_core_up_prgmnvrt),
   .hssi_aibnd_rx_15_aib_dllstr_align_st_core_updnen                                                                                    ( hssi_aibnd_rx_15_aib_dllstr_align_st_core_updnen),
   .hssi_aibnd_rx_15_aib_dllstr_align_st_dftmuxsel                                                                                      ( hssi_aibnd_rx_15_aib_dllstr_align_st_dftmuxsel),
   .hssi_aibnd_rx_15_aib_dllstr_align_st_en                                                                                             ( hssi_aibnd_rx_15_aib_dllstr_align_st_en),
   .hssi_aibnd_rx_15_aib_dllstr_align_st_hps_ctrl_en                                                                                    ( hssi_aibnd_rx_15_aib_dllstr_align_st_hps_ctrl_en),
   .hssi_aibnd_rx_15_aib_dllstr_align_st_lockreq_muxsel                                                                                 ( hssi_aibnd_rx_15_aib_dllstr_align_st_lockreq_muxsel),
   .hssi_aibnd_rx_15_aib_dllstr_align_st_new_dll                                                                                        ( hssi_aibnd_rx_15_aib_dllstr_align_st_new_dll),
   .hssi_aibnd_rx_15_aib_dllstr_align_st_rst                                                                                            ( hssi_aibnd_rx_15_aib_dllstr_align_st_rst),
   .hssi_aibnd_rx_15_aib_dllstr_align_st_rst_prgmnvrt                                                                                   ( hssi_aibnd_rx_15_aib_dllstr_align_st_rst_prgmnvrt),
   .hssi_aibnd_rx_15_aib_dllstr_align_test_clk_pll_en_n                                                                                 ( hssi_aibnd_rx_15_aib_dllstr_align_test_clk_pll_en_n),
   .hssi_aibnd_rx_15_aib_inctrl_gr0                                                                                                     ( hssi_aibnd_rx_15_aib_inctrl_gr0),
   .hssi_aibnd_rx_15_aib_inctrl_gr1                                                                                                     ( hssi_aibnd_rx_15_aib_inctrl_gr1),
   .hssi_aibnd_rx_15_aib_inctrl_gr2                                                                                                     ( hssi_aibnd_rx_15_aib_inctrl_gr2),
   .hssi_aibnd_rx_15_aib_inctrl_gr3                                                                                                     ( hssi_aibnd_rx_15_aib_inctrl_gr3),
   .hssi_aibnd_rx_15_aib_outctrl_gr0                                                                                                    ( hssi_aibnd_rx_15_aib_outctrl_gr0),
   .hssi_aibnd_rx_15_aib_outctrl_gr1                                                                                                    ( hssi_aibnd_rx_15_aib_outctrl_gr1),
   .hssi_aibnd_rx_15_aib_outctrl_gr2                                                                                                    ( hssi_aibnd_rx_15_aib_outctrl_gr2),
   .hssi_aibnd_rx_15_aib_outndrv_r12                                                                                                    ( hssi_aibnd_rx_15_aib_outndrv_r12),
   .hssi_aibnd_rx_15_aib_outndrv_r34                                                                                                    ( hssi_aibnd_rx_15_aib_outndrv_r34),
   .hssi_aibnd_rx_15_aib_outndrv_r56                                                                                                    ( hssi_aibnd_rx_15_aib_outndrv_r56),
   .hssi_aibnd_rx_15_aib_outndrv_r78                                                                                                    ( hssi_aibnd_rx_15_aib_outndrv_r78),
   .hssi_aibnd_rx_15_aib_outpdrv_r12                                                                                                    ( hssi_aibnd_rx_15_aib_outpdrv_r12),
   .hssi_aibnd_rx_15_aib_outpdrv_r34                                                                                                    ( hssi_aibnd_rx_15_aib_outpdrv_r34),
   .hssi_aibnd_rx_15_aib_outpdrv_r56                                                                                                    ( hssi_aibnd_rx_15_aib_outpdrv_r56),
   .hssi_aibnd_rx_15_aib_outpdrv_r78                                                                                                    ( hssi_aibnd_rx_15_aib_outpdrv_r78),
   .hssi_aibnd_rx_15_aib_red_shift_en                                                                                                   ( hssi_aibnd_rx_15_aib_red_shift_en),
   .hssi_aibnd_rx_15_dft_hssitestip_dll_dcc_en                                                                                          ( hssi_aibnd_rx_15_dft_hssitestip_dll_dcc_en),
   .hssi_aibnd_rx_15_op_mode                                                                                                            ( hssi_aibnd_rx_15_op_mode),
   .hssi_aibnd_rx_15_powerdown_mode                                                                                                     ( hssi_aibnd_rx_15_powerdown_mode),
   .hssi_aibnd_rx_15_powermode_ac                                                                                                       ( hssi_aibnd_rx_15_powermode_ac),
   .hssi_aibnd_rx_15_powermode_dc                                                                                                       ( hssi_aibnd_rx_15_powermode_dc),
   .hssi_aibnd_rx_15_powermode_freq_hz_aib_hssi_rx_transfer_clk                                                                         ( hssi_aibnd_rx_15_powermode_freq_hz_aib_hssi_rx_transfer_clk),
   .hssi_aibnd_rx_15_redundancy_en                                                                                                      ( hssi_aibnd_rx_15_redundancy_en),
   .hssi_aibnd_rx_15_sup_mode                                                                                                           ( hssi_aibnd_rx_15_sup_mode),
   .hssi_aibnd_rx_15_silicon_rev                                                                                                        ( hssi_aibnd_rx_15_silicon_rev),
   .hssi_aibnd_tx_15_aib_datasel_gr0                                                                                                    ( hssi_aibnd_tx_15_aib_datasel_gr0),
   .hssi_aibnd_tx_15_aib_datasel_gr1                                                                                                    ( hssi_aibnd_tx_15_aib_datasel_gr1),
   .hssi_aibnd_tx_15_aib_datasel_gr2                                                                                                    ( hssi_aibnd_tx_15_aib_datasel_gr2),
   .hssi_aibnd_tx_15_aib_datasel_gr3                                                                                                    ( hssi_aibnd_tx_15_aib_datasel_gr3),
   .hssi_aibnd_tx_15_aib_ddrctrl_gr0                                                                                                    ( hssi_aibnd_tx_15_aib_ddrctrl_gr0),
   .hssi_aibnd_tx_15_aib_hssi_tx_transfer_clk_hz                                                                                        ( hssi_aibnd_tx_15_aib_hssi_tx_transfer_clk_hz),
   .hssi_aibnd_tx_15_aib_iinasyncen                                                                                                     ( hssi_aibnd_tx_15_aib_iinasyncen),
   .hssi_aibnd_tx_15_aib_iinclken                                                                                                       ( hssi_aibnd_tx_15_aib_iinclken),
   .hssi_aibnd_tx_15_aib_outctrl_gr0                                                                                                    ( hssi_aibnd_tx_15_aib_outctrl_gr0),
   .hssi_aibnd_tx_15_aib_outctrl_gr1                                                                                                    ( hssi_aibnd_tx_15_aib_outctrl_gr1),
   .hssi_aibnd_tx_15_aib_outctrl_gr2                                                                                                    ( hssi_aibnd_tx_15_aib_outctrl_gr2),
   .hssi_aibnd_tx_15_aib_outctrl_gr3                                                                                                    ( hssi_aibnd_tx_15_aib_outctrl_gr3),
   .hssi_aibnd_tx_15_aib_outndrv_r34                                                                                                    ( hssi_aibnd_tx_15_aib_outndrv_r34),
   .hssi_aibnd_tx_15_aib_outndrv_r56                                                                                                    ( hssi_aibnd_tx_15_aib_outndrv_r56),
   .hssi_aibnd_tx_15_aib_outpdrv_r34                                                                                                    ( hssi_aibnd_tx_15_aib_outpdrv_r34),
   .hssi_aibnd_tx_15_aib_outpdrv_r56                                                                                                    ( hssi_aibnd_tx_15_aib_outpdrv_r56),
   .hssi_aibnd_tx_15_aib_red_dirclkn_shiften                                                                                            ( hssi_aibnd_tx_15_aib_red_dirclkn_shiften),
   .hssi_aibnd_tx_15_aib_red_dirclkp_shiften                                                                                            ( hssi_aibnd_tx_15_aib_red_dirclkp_shiften),
   .hssi_aibnd_tx_15_aib_red_drx_shiften                                                                                                ( hssi_aibnd_tx_15_aib_red_drx_shiften),
   .hssi_aibnd_tx_15_aib_red_dtx_shiften                                                                                                ( hssi_aibnd_tx_15_aib_red_dtx_shiften),
   .hssi_aibnd_tx_15_aib_red_pout_shiften                                                                                               ( hssi_aibnd_tx_15_aib_red_pout_shiften),
   .hssi_aibnd_tx_15_aib_red_rx_shiften                                                                                                 ( hssi_aibnd_tx_15_aib_red_rx_shiften),
   .hssi_aibnd_tx_15_aib_red_tx_shiften                                                                                                 ( hssi_aibnd_tx_15_aib_red_tx_shiften),
   .hssi_aibnd_tx_15_aib_red_txferclkout_shiften                                                                                        ( hssi_aibnd_tx_15_aib_red_txferclkout_shiften),
   .hssi_aibnd_tx_15_aib_red_txferclkoutn_shiften                                                                                       ( hssi_aibnd_tx_15_aib_red_txferclkoutn_shiften),
   .hssi_aibnd_tx_15_aib_tx_clkdiv                                                                                                      ( hssi_aibnd_tx_15_aib_tx_clkdiv),
   .hssi_aibnd_tx_15_aib_tx_dcc_byp                                                                                                     ( hssi_aibnd_tx_15_aib_tx_dcc_byp),
   .hssi_aibnd_tx_15_aib_tx_dcc_byp_iocsr_unused                                                                                        ( hssi_aibnd_tx_15_aib_tx_dcc_byp_iocsr_unused),
   .hssi_aibnd_tx_15_aib_tx_dcc_cont_cal                                                                                                ( hssi_aibnd_tx_15_aib_tx_dcc_cont_cal),
   .hssi_aibnd_tx_15_aib_tx_dcc_cont_cal_iocsr_unused                                                                                   ( hssi_aibnd_tx_15_aib_tx_dcc_cont_cal_iocsr_unused),
   .hssi_aibnd_tx_15_aib_tx_dcc_dft                                                                                                     ( hssi_aibnd_tx_15_aib_tx_dcc_dft),
   .hssi_aibnd_tx_15_aib_tx_dcc_dft_sel                                                                                                 ( hssi_aibnd_tx_15_aib_tx_dcc_dft_sel),
   .hssi_aibnd_tx_15_aib_tx_dcc_dll_dft_sel                                                                                             ( hssi_aibnd_tx_15_aib_tx_dcc_dll_dft_sel),
   .hssi_aibnd_tx_15_aib_tx_dcc_dll_entest                                                                                              ( hssi_aibnd_tx_15_aib_tx_dcc_dll_entest),
   .hssi_aibnd_tx_15_aib_tx_dcc_dy_ctl_static                                                                                           ( hssi_aibnd_tx_15_aib_tx_dcc_dy_ctl_static),
   .hssi_aibnd_tx_15_aib_tx_dcc_dy_ctlsel                                                                                               ( hssi_aibnd_tx_15_aib_tx_dcc_dy_ctlsel),
   .hssi_aibnd_tx_15_aib_tx_dcc_en                                                                                                      ( hssi_aibnd_tx_15_aib_tx_dcc_en),
   .hssi_aibnd_tx_15_aib_tx_dcc_en_iocsr_unused                                                                                         ( hssi_aibnd_tx_15_aib_tx_dcc_en_iocsr_unused),
   .hssi_aibnd_tx_15_aib_tx_dcc_manual_dn                                                                                               ( hssi_aibnd_tx_15_aib_tx_dcc_manual_dn),
   .hssi_aibnd_tx_15_aib_tx_dcc_manual_up                                                                                               ( hssi_aibnd_tx_15_aib_tx_dcc_manual_up),
   .hssi_aibnd_tx_15_aib_tx_dcc_rst_prgmnvrt                                                                                            ( hssi_aibnd_tx_15_aib_tx_dcc_rst_prgmnvrt),
   .hssi_aibnd_tx_15_aib_tx_dcc_st_core_dn_prgmnvrt                                                                                     ( hssi_aibnd_tx_15_aib_tx_dcc_st_core_dn_prgmnvrt),
   .hssi_aibnd_tx_15_aib_tx_dcc_st_core_up_prgmnvrt                                                                                     ( hssi_aibnd_tx_15_aib_tx_dcc_st_core_up_prgmnvrt),
   .hssi_aibnd_tx_15_aib_tx_dcc_st_core_updnen                                                                                          ( hssi_aibnd_tx_15_aib_tx_dcc_st_core_updnen),
   .hssi_aibnd_tx_15_aib_tx_dcc_st_dftmuxsel                                                                                            ( hssi_aibnd_tx_15_aib_tx_dcc_st_dftmuxsel),
   .hssi_aibnd_tx_15_aib_tx_dcc_st_dly_pst                                                                                              ( hssi_aibnd_tx_15_aib_tx_dcc_st_dly_pst),
   .hssi_aibnd_tx_15_aib_tx_dcc_st_en                                                                                                   ( hssi_aibnd_tx_15_aib_tx_dcc_st_en),
   .hssi_aibnd_tx_15_aib_tx_dcc_st_hps_ctrl_en                                                                                          ( hssi_aibnd_tx_15_aib_tx_dcc_st_hps_ctrl_en),
   .hssi_aibnd_tx_15_aib_tx_dcc_st_lockreq_muxsel                                                                                       ( hssi_aibnd_tx_15_aib_tx_dcc_st_lockreq_muxsel),
   .hssi_aibnd_tx_15_aib_tx_dcc_st_new_dll                                                                                              ( hssi_aibnd_tx_15_aib_tx_dcc_st_new_dll),
   .hssi_aibnd_tx_15_aib_tx_dcc_st_rst                                                                                                  ( hssi_aibnd_tx_15_aib_tx_dcc_st_rst),
   .hssi_aibnd_tx_15_aib_tx_dcc_test_clk_pll_en_n                                                                                       ( hssi_aibnd_tx_15_aib_tx_dcc_test_clk_pll_en_n),
   .hssi_aibnd_tx_15_aib_tx_halfcode                                                                                                    ( hssi_aibnd_tx_15_aib_tx_halfcode),
   .hssi_aibnd_tx_15_aib_tx_selflock                                                                                                    ( hssi_aibnd_tx_15_aib_tx_selflock),
   .hssi_aibnd_tx_15_dfd_dll_dcc_en                                                                                                     ( hssi_aibnd_tx_15_dfd_dll_dcc_en),
   .hssi_aibnd_tx_15_dft_hssitestip_dll_dcc_en                                                                                          ( hssi_aibnd_tx_15_dft_hssitestip_dll_dcc_en),
   .hssi_aibnd_tx_15_op_mode                                                                                                            ( hssi_aibnd_tx_15_op_mode),
   .hssi_aibnd_tx_15_powerdown_mode                                                                                                     ( hssi_aibnd_tx_15_powerdown_mode),
   .hssi_aibnd_tx_15_powermode_ac                                                                                                       ( hssi_aibnd_tx_15_powermode_ac),
   .hssi_aibnd_tx_15_powermode_dc                                                                                                       ( hssi_aibnd_tx_15_powermode_dc),
   .hssi_aibnd_tx_15_powermode_freq_hz_aib_hssi_tx_transfer_clk                                                                         ( hssi_aibnd_tx_15_powermode_freq_hz_aib_hssi_tx_transfer_clk),
   .hssi_aibnd_tx_15_redundancy_en                                                                                                      ( hssi_aibnd_tx_15_redundancy_en),
   .hssi_aibnd_tx_15_sup_mode                                                                                                           ( hssi_aibnd_tx_15_sup_mode),
   .hssi_aibnd_tx_15_silicon_rev                                                                                                        ( hssi_aibnd_tx_15_silicon_rev),
   .hssi_pldadapt_tx_15_aib_clk1_sel                                                                                                    ( hssi_pldadapt_tx_15_aib_clk1_sel),
   .hssi_pldadapt_tx_15_aib_clk2_sel                                                                                                    ( hssi_pldadapt_tx_15_aib_clk2_sel),
   .hssi_pldadapt_tx_15_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                           ( hssi_pldadapt_tx_15_hdpldadapt_aib_fabric_pld_pma_hclk_hz),
   .hssi_pldadapt_tx_15_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz                                                                         ( hssi_pldadapt_tx_15_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz),
   .hssi_pldadapt_tx_15_hdpldadapt_aib_fabric_tx_sr_clk_in_hz                                                                           ( hssi_pldadapt_tx_15_hdpldadapt_aib_fabric_tx_sr_clk_in_hz),
   .hssi_pldadapt_tx_15_bonding_dft_en                                                                                                  ( hssi_pldadapt_tx_15_bonding_dft_en),
   .hssi_pldadapt_tx_15_bonding_dft_val                                                                                                 ( hssi_pldadapt_tx_15_bonding_dft_val),
   .hssi_pldadapt_tx_15_chnl_bonding                                                                                                    ( hssi_pldadapt_tx_15_chnl_bonding),
   .hssi_pldadapt_tx_15_comp_cnt                                                                                                        ( hssi_pldadapt_tx_15_comp_cnt),
   .hssi_pldadapt_tx_15_compin_sel                                                                                                      ( hssi_pldadapt_tx_15_compin_sel),
   .hssi_pldadapt_tx_15_hdpldadapt_csr_clk_hz                                                                                           ( hssi_pldadapt_tx_15_hdpldadapt_csr_clk_hz),
   .hssi_pldadapt_tx_15_ctrl_plane_bonding                                                                                              ( hssi_pldadapt_tx_15_ctrl_plane_bonding),
   .hssi_pldadapt_tx_15_ds_bypass_pipeln                                                                                                ( hssi_pldadapt_tx_15_ds_bypass_pipeln),
   .hssi_pldadapt_tx_15_ds_last_chnl                                                                                                    ( hssi_pldadapt_tx_15_ds_last_chnl),
   .hssi_pldadapt_tx_15_ds_master                                                                                                       ( hssi_pldadapt_tx_15_ds_master),
   .hssi_pldadapt_tx_15_duplex_mode                                                                                                     ( hssi_pldadapt_tx_15_duplex_mode),
   .hssi_pldadapt_tx_15_dv_bond                                                                                                         ( hssi_pldadapt_tx_15_dv_bond),
   .hssi_pldadapt_tx_15_dv_gen                                                                                                          ( hssi_pldadapt_tx_15_dv_gen),
   .hssi_pldadapt_tx_15_fifo_double_write                                                                                               ( hssi_pldadapt_tx_15_fifo_double_write),
   .hssi_pldadapt_tx_15_fifo_mode                                                                                                       ( hssi_pldadapt_tx_15_fifo_mode),
   .hssi_pldadapt_tx_15_fifo_rd_clk_frm_gen_scg_en                                                                                      ( hssi_pldadapt_tx_15_fifo_rd_clk_frm_gen_scg_en),
   .hssi_pldadapt_tx_15_fifo_rd_clk_scg_en                                                                                              ( hssi_pldadapt_tx_15_fifo_rd_clk_scg_en),
   .hssi_pldadapt_tx_15_fifo_rd_clk_sel                                                                                                 ( hssi_pldadapt_tx_15_fifo_rd_clk_sel),
   .hssi_pldadapt_tx_15_fifo_stop_rd                                                                                                    ( hssi_pldadapt_tx_15_fifo_stop_rd),
   .hssi_pldadapt_tx_15_fifo_stop_wr                                                                                                    ( hssi_pldadapt_tx_15_fifo_stop_wr),
   .hssi_pldadapt_tx_15_fifo_width                                                                                                      ( hssi_pldadapt_tx_15_fifo_width),
   .hssi_pldadapt_tx_15_fifo_wr_clk_scg_en                                                                                              ( hssi_pldadapt_tx_15_fifo_wr_clk_scg_en),
   .hssi_pldadapt_tx_15_fpll_shared_direct_async_in_sel                                                                                 ( hssi_pldadapt_tx_15_fpll_shared_direct_async_in_sel),
   .hssi_pldadapt_tx_15_frmgen_burst                                                                                                    ( hssi_pldadapt_tx_15_frmgen_burst),
   .hssi_pldadapt_tx_15_frmgen_bypass                                                                                                   ( hssi_pldadapt_tx_15_frmgen_bypass),
   .hssi_pldadapt_tx_15_frmgen_mfrm_length                                                                                              ( hssi_pldadapt_tx_15_frmgen_mfrm_length),
   .hssi_pldadapt_tx_15_frmgen_pipeln                                                                                                   ( hssi_pldadapt_tx_15_frmgen_pipeln),
   .hssi_pldadapt_tx_15_frmgen_pyld_ins                                                                                                 ( hssi_pldadapt_tx_15_frmgen_pyld_ins),
   .hssi_pldadapt_tx_15_frmgen_wordslip                                                                                                 ( hssi_pldadapt_tx_15_frmgen_wordslip),
   .hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit0_rst_val                                                                                     ( hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit0_rst_val),
   .hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit1_rst_val                                                                                     ( hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit1_rst_val),
   .hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit2_rst_val                                                                                     ( hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit2_rst_val),
   .hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit3_rst_val                                                                                     ( hssi_pldadapt_tx_15_fsr_hip_fsr_in_bit3_rst_val),
   .hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit0_rst_val                                                                                    ( hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit0_rst_val),
   .hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit1_rst_val                                                                                    ( hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit1_rst_val),
   .hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit2_rst_val                                                                                    ( hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit2_rst_val),
   .hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit3_rst_val                                                                                    ( hssi_pldadapt_tx_15_fsr_hip_fsr_out_bit3_rst_val),
   .hssi_pldadapt_tx_15_fsr_mask_tx_pll_rst_val                                                                                         ( hssi_pldadapt_tx_15_fsr_mask_tx_pll_rst_val),
   .hssi_pldadapt_tx_15_fsr_pld_txelecidle_rst_val                                                                                      ( hssi_pldadapt_tx_15_fsr_pld_txelecidle_rst_val),
   .hssi_pldadapt_tx_15_gb_tx_idwidth                                                                                                   ( hssi_pldadapt_tx_15_gb_tx_idwidth),
   .hssi_pldadapt_tx_15_gb_tx_odwidth                                                                                                   ( hssi_pldadapt_tx_15_gb_tx_odwidth),
   .hssi_pldadapt_tx_15_hip_mode                                                                                                        ( hssi_pldadapt_tx_15_hip_mode),
   .hssi_pldadapt_tx_15_hip_osc_clk_scg_en                                                                                              ( hssi_pldadapt_tx_15_hip_osc_clk_scg_en),
   .hssi_pldadapt_tx_15_hrdrst_dcd_cal_done_bypass                                                                                      ( hssi_pldadapt_tx_15_hrdrst_dcd_cal_done_bypass),
   .hssi_pldadapt_tx_15_hrdrst_rst_sm_dis                                                                                               ( hssi_pldadapt_tx_15_hrdrst_rst_sm_dis),
   .hssi_pldadapt_tx_15_hrdrst_rx_osc_clk_scg_en                                                                                        ( hssi_pldadapt_tx_15_hrdrst_rx_osc_clk_scg_en),
   .hssi_pldadapt_tx_15_hrdrst_user_ctl_en                                                                                              ( hssi_pldadapt_tx_15_hrdrst_user_ctl_en),
   .hssi_pldadapt_tx_15_indv                                                                                                            ( hssi_pldadapt_tx_15_indv),
   .hssi_pldadapt_tx_15_is_paired_with                                                                                                  ( hssi_pldadapt_tx_15_is_paired_with),
   .hssi_pldadapt_tx_15_loopback_mode                                                                                                   ( hssi_pldadapt_tx_15_loopback_mode),
   .hssi_pldadapt_tx_15_low_latency_en                                                                                                  ( hssi_pldadapt_tx_15_low_latency_en),
   .hssi_pldadapt_tx_15_osc_clk_scg_en                                                                                                  ( hssi_pldadapt_tx_15_osc_clk_scg_en),
   .hssi_pldadapt_tx_15_phcomp_rd_del                                                                                                   ( hssi_pldadapt_tx_15_phcomp_rd_del),
   .hssi_pldadapt_tx_15_pipe_mode                                                                                                       ( hssi_pldadapt_tx_15_pipe_mode),
   .hssi_pldadapt_tx_15_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                              ( hssi_pldadapt_tx_15_hdpldadapt_pld_avmm1_clk_rowclk_hz),
   .hssi_pldadapt_tx_15_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                              ( hssi_pldadapt_tx_15_hdpldadapt_pld_avmm2_clk_rowclk_hz),
   .hssi_pldadapt_tx_15_pld_clk1_delay_en                                                                                               ( hssi_pldadapt_tx_15_pld_clk1_delay_en),
   .hssi_pldadapt_tx_15_pld_clk1_delay_sel                                                                                              ( hssi_pldadapt_tx_15_pld_clk1_delay_sel),
   .hssi_pldadapt_tx_15_pld_clk1_inv_en                                                                                                 ( hssi_pldadapt_tx_15_pld_clk1_inv_en),
   .hssi_pldadapt_tx_15_pld_clk1_sel                                                                                                    ( hssi_pldadapt_tx_15_pld_clk1_sel),
   .hssi_pldadapt_tx_15_pld_clk2_sel                                                                                                    ( hssi_pldadapt_tx_15_pld_clk2_sel),
   .hssi_pldadapt_tx_15_hdpldadapt_pld_sclk1_rowclk_hz                                                                                  ( hssi_pldadapt_tx_15_hdpldadapt_pld_sclk1_rowclk_hz),
   .hssi_pldadapt_tx_15_hdpldadapt_pld_sclk2_rowclk_hz                                                                                  ( hssi_pldadapt_tx_15_hdpldadapt_pld_sclk2_rowclk_hz),
   .hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk1_dcm_hz                                                                                   ( hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk1_dcm_hz),
   .hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk1_rowclk_hz                                                                                ( hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk1_rowclk_hz),
   .hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk2_dcm_hz                                                                                   ( hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk2_dcm_hz),
   .hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk2_rowclk_hz                                                                                ( hssi_pldadapt_tx_15_hdpldadapt_pld_tx_clk2_rowclk_hz),
   .hssi_pldadapt_tx_15_pma_aib_tx_clk_expected_setting                                                                                 ( hssi_pldadapt_tx_15_pma_aib_tx_clk_expected_setting),
   .hssi_pldadapt_tx_15_powerdown_mode                                                                                                  ( hssi_pldadapt_tx_15_powerdown_mode),
   .hssi_pldadapt_tx_15_powermode_dc                                                                                                    ( hssi_pldadapt_tx_15_powermode_dc),
   .hssi_pldadapt_tx_15_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                       ( hssi_pldadapt_tx_15_powermode_freq_hz_aib_fabric_rx_sr_clk_in),
   .hssi_pldadapt_tx_15_powermode_freq_hz_pld_tx_clk1_dcm                                                                               ( hssi_pldadapt_tx_15_powermode_freq_hz_pld_tx_clk1_dcm),
   .hssi_pldadapt_tx_15_sh_err                                                                                                          ( hssi_pldadapt_tx_15_sh_err),
   .hssi_pldadapt_tx_15_hdpldadapt_speed_grade                                                                                          ( hssi_pldadapt_tx_15_hdpldadapt_speed_grade),
   .hssi_pldadapt_tx_15_hdpldadapt_sr_sr_testbus_sel                                                                                    ( hssi_pldadapt_tx_15_hdpldadapt_sr_sr_testbus_sel),
   .hssi_pldadapt_tx_15_stretch_num_stages                                                                                              ( hssi_pldadapt_tx_15_stretch_num_stages),
   .hssi_pldadapt_tx_15_sup_mode                                                                                                        ( hssi_pldadapt_tx_15_sup_mode),
   .hssi_pldadapt_tx_15_tx_datapath_tb_sel                                                                                              ( hssi_pldadapt_tx_15_tx_datapath_tb_sel),
   .hssi_pldadapt_tx_15_tx_fastbond_rden                                                                                                ( hssi_pldadapt_tx_15_tx_fastbond_rden),
   .hssi_pldadapt_tx_15_tx_fastbond_wren                                                                                                ( hssi_pldadapt_tx_15_tx_fastbond_wren),
   .hssi_pldadapt_tx_15_tx_fifo_power_mode                                                                                              ( hssi_pldadapt_tx_15_tx_fifo_power_mode),
   .hssi_pldadapt_tx_15_tx_fifo_read_latency_adjust                                                                                     ( hssi_pldadapt_tx_15_tx_fifo_read_latency_adjust),
   .hssi_pldadapt_tx_15_tx_fifo_write_latency_adjust                                                                                    ( hssi_pldadapt_tx_15_tx_fifo_write_latency_adjust),
   .hssi_pldadapt_tx_15_tx_hip_aib_ssr_in_polling_bypass                                                                                ( hssi_pldadapt_tx_15_tx_hip_aib_ssr_in_polling_bypass),
   .hssi_pldadapt_tx_15_tx_osc_clock_setting                                                                                            ( hssi_pldadapt_tx_15_tx_osc_clock_setting),
   .hssi_pldadapt_tx_15_tx_pld_10g_tx_bitslip_polling_bypass                                                                            ( hssi_pldadapt_tx_15_tx_pld_10g_tx_bitslip_polling_bypass),
   .hssi_pldadapt_tx_15_tx_pld_8g_tx_boundary_sel_polling_bypass                                                                        ( hssi_pldadapt_tx_15_tx_pld_8g_tx_boundary_sel_polling_bypass),
   .hssi_pldadapt_tx_15_tx_pld_pma_fpll_cnt_sel_polling_bypass                                                                          ( hssi_pldadapt_tx_15_tx_pld_pma_fpll_cnt_sel_polling_bypass),
   .hssi_pldadapt_tx_15_tx_pld_pma_fpll_num_phase_shifts_polling_bypass                                                                 ( hssi_pldadapt_tx_15_tx_pld_pma_fpll_num_phase_shifts_polling_bypass),
   .hssi_pldadapt_tx_15_tx_usertest_sel                                                                                                 ( hssi_pldadapt_tx_15_tx_usertest_sel),
   .hssi_pldadapt_tx_15_txfifo_empty                                                                                                    ( hssi_pldadapt_tx_15_txfifo_empty),
   .hssi_pldadapt_tx_15_txfifo_full                                                                                                     ( hssi_pldadapt_tx_15_txfifo_full),
   .hssi_pldadapt_tx_15_txfifo_mode                                                                                                     ( hssi_pldadapt_tx_15_txfifo_mode),
   .hssi_pldadapt_tx_15_txfifo_pempty                                                                                                   ( hssi_pldadapt_tx_15_txfifo_pempty),
   .hssi_pldadapt_tx_15_txfifo_pfull                                                                                                    ( hssi_pldadapt_tx_15_txfifo_pfull),
   .hssi_pldadapt_tx_15_us_bypass_pipeln                                                                                                ( hssi_pldadapt_tx_15_us_bypass_pipeln),
   .hssi_pldadapt_tx_15_us_last_chnl                                                                                                    ( hssi_pldadapt_tx_15_us_last_chnl),
   .hssi_pldadapt_tx_15_us_master                                                                                                       ( hssi_pldadapt_tx_15_us_master),
   .hssi_pldadapt_tx_15_word_align_enable                                                                                               ( hssi_pldadapt_tx_15_word_align_enable),
   .hssi_pldadapt_tx_15_word_mark                                                                                                       ( hssi_pldadapt_tx_15_word_mark),
   .hssi_pldadapt_tx_15_silicon_rev                                                                                                     ( hssi_pldadapt_tx_15_silicon_rev),
   .hssi_pldadapt_tx_15_reconfig_settings                                                                                               ( hssi_pldadapt_tx_15_reconfig_settings),
   .hssi_pldadapt_rx_15_aib_clk1_sel                                                                                                    ( hssi_pldadapt_rx_15_aib_clk1_sel),
   .hssi_pldadapt_rx_15_aib_clk2_sel                                                                                                    ( hssi_pldadapt_rx_15_aib_clk2_sel),
   .hssi_pldadapt_rx_15_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                           ( hssi_pldadapt_rx_15_hdpldadapt_aib_fabric_pld_pma_hclk_hz),
   .hssi_pldadapt_rx_15_hdpldadapt_aib_fabric_rx_sr_clk_in_hz                                                                           ( hssi_pldadapt_rx_15_hdpldadapt_aib_fabric_rx_sr_clk_in_hz),
   .hssi_pldadapt_rx_15_hdpldadapt_aib_fabric_rx_transfer_clk_hz                                                                        ( hssi_pldadapt_rx_15_hdpldadapt_aib_fabric_rx_transfer_clk_hz),
   .hssi_pldadapt_rx_15_asn_bypass_pma_pcie_sw_done                                                                                     ( hssi_pldadapt_rx_15_asn_bypass_pma_pcie_sw_done),
   .hssi_pldadapt_rx_15_asn_en                                                                                                          ( hssi_pldadapt_rx_15_asn_en),
   .hssi_pldadapt_rx_15_asn_wait_for_dll_reset_cnt                                                                                      ( hssi_pldadapt_rx_15_asn_wait_for_dll_reset_cnt),
   .hssi_pldadapt_rx_15_asn_wait_for_fifo_flush_cnt                                                                                     ( hssi_pldadapt_rx_15_asn_wait_for_fifo_flush_cnt),
   .hssi_pldadapt_rx_15_asn_wait_for_pma_pcie_sw_done_cnt                                                                               ( hssi_pldadapt_rx_15_asn_wait_for_pma_pcie_sw_done_cnt),
   .hssi_pldadapt_rx_15_bonding_dft_en                                                                                                  ( hssi_pldadapt_rx_15_bonding_dft_en),
   .hssi_pldadapt_rx_15_bonding_dft_val                                                                                                 ( hssi_pldadapt_rx_15_bonding_dft_val),
   .hssi_pldadapt_rx_15_chnl_bonding                                                                                                    ( hssi_pldadapt_rx_15_chnl_bonding),
   .hssi_pldadapt_rx_15_clock_del_measure_enable                                                                                        ( hssi_pldadapt_rx_15_clock_del_measure_enable),
   .hssi_pldadapt_rx_15_comp_cnt                                                                                                        ( hssi_pldadapt_rx_15_comp_cnt),
   .hssi_pldadapt_rx_15_compin_sel                                                                                                      ( hssi_pldadapt_rx_15_compin_sel),
   .hssi_pldadapt_rx_15_hdpldadapt_csr_clk_hz                                                                                           ( hssi_pldadapt_rx_15_hdpldadapt_csr_clk_hz),
   .hssi_pldadapt_rx_15_ctrl_plane_bonding                                                                                              ( hssi_pldadapt_rx_15_ctrl_plane_bonding),
   .hssi_pldadapt_rx_15_ds_bypass_pipeln                                                                                                ( hssi_pldadapt_rx_15_ds_bypass_pipeln),
   .hssi_pldadapt_rx_15_ds_last_chnl                                                                                                    ( hssi_pldadapt_rx_15_ds_last_chnl),
   .hssi_pldadapt_rx_15_ds_master                                                                                                       ( hssi_pldadapt_rx_15_ds_master),
   .hssi_pldadapt_rx_15_duplex_mode                                                                                                     ( hssi_pldadapt_rx_15_duplex_mode),
   .hssi_pldadapt_rx_15_dv_mode                                                                                                         ( hssi_pldadapt_rx_15_dv_mode),
   .hssi_pldadapt_rx_15_fifo_double_read                                                                                                ( hssi_pldadapt_rx_15_fifo_double_read),
   .hssi_pldadapt_rx_15_fifo_mode                                                                                                       ( hssi_pldadapt_rx_15_fifo_mode),
   .hssi_pldadapt_rx_15_fifo_rd_clk_ins_sm_scg_en                                                                                       ( hssi_pldadapt_rx_15_fifo_rd_clk_ins_sm_scg_en),
   .hssi_pldadapt_rx_15_fifo_rd_clk_scg_en                                                                                              ( hssi_pldadapt_rx_15_fifo_rd_clk_scg_en),
   .hssi_pldadapt_rx_15_fifo_rd_clk_sel                                                                                                 ( hssi_pldadapt_rx_15_fifo_rd_clk_sel),
   .hssi_pldadapt_rx_15_fifo_stop_rd                                                                                                    ( hssi_pldadapt_rx_15_fifo_stop_rd),
   .hssi_pldadapt_rx_15_fifo_stop_wr                                                                                                    ( hssi_pldadapt_rx_15_fifo_stop_wr),
   .hssi_pldadapt_rx_15_fifo_width                                                                                                      ( hssi_pldadapt_rx_15_fifo_width),
   .hssi_pldadapt_rx_15_fifo_wr_clk_del_sm_scg_en                                                                                       ( hssi_pldadapt_rx_15_fifo_wr_clk_del_sm_scg_en),
   .hssi_pldadapt_rx_15_fifo_wr_clk_scg_en                                                                                              ( hssi_pldadapt_rx_15_fifo_wr_clk_scg_en),
   .hssi_pldadapt_rx_15_fifo_wr_clk_sel                                                                                                 ( hssi_pldadapt_rx_15_fifo_wr_clk_sel),
   .hssi_pldadapt_rx_15_free_run_div_clk                                                                                                ( hssi_pldadapt_rx_15_free_run_div_clk),
   .hssi_pldadapt_rx_15_fsr_pld_10g_rx_crc32_err_rst_val                                                                                ( hssi_pldadapt_rx_15_fsr_pld_10g_rx_crc32_err_rst_val),
   .hssi_pldadapt_rx_15_fsr_pld_8g_sigdet_out_rst_val                                                                                   ( hssi_pldadapt_rx_15_fsr_pld_8g_sigdet_out_rst_val),
   .hssi_pldadapt_rx_15_fsr_pld_ltd_b_rst_val                                                                                           ( hssi_pldadapt_rx_15_fsr_pld_ltd_b_rst_val),
   .hssi_pldadapt_rx_15_fsr_pld_ltr_rst_val                                                                                             ( hssi_pldadapt_rx_15_fsr_pld_ltr_rst_val),
   .hssi_pldadapt_rx_15_fsr_pld_rx_fifo_align_clr_rst_val                                                                               ( hssi_pldadapt_rx_15_fsr_pld_rx_fifo_align_clr_rst_val),
   .hssi_pldadapt_rx_15_gb_rx_idwidth                                                                                                   ( hssi_pldadapt_rx_15_gb_rx_idwidth),
   .hssi_pldadapt_rx_15_gb_rx_odwidth                                                                                                   ( hssi_pldadapt_rx_15_gb_rx_odwidth),
   .hssi_pldadapt_rx_15_hip_mode                                                                                                        ( hssi_pldadapt_rx_15_hip_mode),
   .hssi_pldadapt_rx_15_hrdrst_align_bypass                                                                                             ( hssi_pldadapt_rx_15_hrdrst_align_bypass),
   .hssi_pldadapt_rx_15_hrdrst_dll_lock_bypass                                                                                          ( hssi_pldadapt_rx_15_hrdrst_dll_lock_bypass),
   .hssi_pldadapt_rx_15_hrdrst_rst_sm_dis                                                                                               ( hssi_pldadapt_rx_15_hrdrst_rst_sm_dis),
   .hssi_pldadapt_rx_15_hrdrst_rx_osc_clk_scg_en                                                                                        ( hssi_pldadapt_rx_15_hrdrst_rx_osc_clk_scg_en),
   .hssi_pldadapt_rx_15_hrdrst_user_ctl_en                                                                                              ( hssi_pldadapt_rx_15_hrdrst_user_ctl_en),
   .hssi_pldadapt_rx_15_indv                                                                                                            ( hssi_pldadapt_rx_15_indv),
   .hssi_pldadapt_rx_15_internal_clk1_sel1                                                                                              ( hssi_pldadapt_rx_15_internal_clk1_sel1),
   .hssi_pldadapt_rx_15_internal_clk1_sel2                                                                                              ( hssi_pldadapt_rx_15_internal_clk1_sel2),
   .hssi_pldadapt_rx_15_internal_clk2_sel1                                                                                              ( hssi_pldadapt_rx_15_internal_clk2_sel1),
   .hssi_pldadapt_rx_15_internal_clk2_sel2                                                                                              ( hssi_pldadapt_rx_15_internal_clk2_sel2),
   .hssi_pldadapt_rx_15_is_paired_with                                                                                                  ( hssi_pldadapt_rx_15_is_paired_with),
   .hssi_pldadapt_rx_15_loopback_mode                                                                                                   ( hssi_pldadapt_rx_15_loopback_mode),
   .hssi_pldadapt_rx_15_low_latency_en                                                                                                  ( hssi_pldadapt_rx_15_low_latency_en),
   .hssi_pldadapt_rx_15_lpbk_mode                                                                                                       ( hssi_pldadapt_rx_15_lpbk_mode),
   .hssi_pldadapt_rx_15_osc_clk_scg_en                                                                                                  ( hssi_pldadapt_rx_15_osc_clk_scg_en),
   .hssi_pldadapt_rx_15_phcomp_rd_del                                                                                                   ( hssi_pldadapt_rx_15_phcomp_rd_del),
   .hssi_pldadapt_rx_15_pipe_enable                                                                                                     ( hssi_pldadapt_rx_15_pipe_enable),
   .hssi_pldadapt_rx_15_pipe_mode                                                                                                       ( hssi_pldadapt_rx_15_pipe_mode),
   .hssi_pldadapt_rx_15_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                              ( hssi_pldadapt_rx_15_hdpldadapt_pld_avmm1_clk_rowclk_hz),
   .hssi_pldadapt_rx_15_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                              ( hssi_pldadapt_rx_15_hdpldadapt_pld_avmm2_clk_rowclk_hz),
   .hssi_pldadapt_rx_15_pld_clk1_delay_en                                                                                               ( hssi_pldadapt_rx_15_pld_clk1_delay_en),
   .hssi_pldadapt_rx_15_pld_clk1_delay_sel                                                                                              ( hssi_pldadapt_rx_15_pld_clk1_delay_sel),
   .hssi_pldadapt_rx_15_pld_clk1_inv_en                                                                                                 ( hssi_pldadapt_rx_15_pld_clk1_inv_en),
   .hssi_pldadapt_rx_15_pld_clk1_sel                                                                                                    ( hssi_pldadapt_rx_15_pld_clk1_sel),
   .hssi_pldadapt_rx_15_hdpldadapt_pld_rx_clk1_dcm_hz                                                                                   ( hssi_pldadapt_rx_15_hdpldadapt_pld_rx_clk1_dcm_hz),
   .hssi_pldadapt_rx_15_hdpldadapt_pld_rx_clk1_rowclk_hz                                                                                ( hssi_pldadapt_rx_15_hdpldadapt_pld_rx_clk1_rowclk_hz),
   .hssi_pldadapt_rx_15_hdpldadapt_pld_sclk1_rowclk_hz                                                                                  ( hssi_pldadapt_rx_15_hdpldadapt_pld_sclk1_rowclk_hz),
   .hssi_pldadapt_rx_15_hdpldadapt_pld_sclk2_rowclk_hz                                                                                  ( hssi_pldadapt_rx_15_hdpldadapt_pld_sclk2_rowclk_hz),
   .hssi_pldadapt_rx_15_pma_hclk_scg_en                                                                                                 ( hssi_pldadapt_rx_15_pma_hclk_scg_en),
   .hssi_pldadapt_rx_15_powerdown_mode                                                                                                  ( hssi_pldadapt_rx_15_powerdown_mode),
   .hssi_pldadapt_rx_15_powermode_dc                                                                                                    ( hssi_pldadapt_rx_15_powermode_dc),
   .hssi_pldadapt_rx_15_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                       ( hssi_pldadapt_rx_15_powermode_freq_hz_aib_fabric_rx_sr_clk_in),
   .hssi_pldadapt_rx_15_powermode_freq_hz_pld_rx_clk1_dcm                                                                               ( hssi_pldadapt_rx_15_powermode_freq_hz_pld_rx_clk1_dcm),
   .hssi_pldadapt_rx_15_rx_datapath_tb_sel                                                                                              ( hssi_pldadapt_rx_15_rx_datapath_tb_sel),
   .hssi_pldadapt_rx_15_rx_fastbond_rden                                                                                                ( hssi_pldadapt_rx_15_rx_fastbond_rden),
   .hssi_pldadapt_rx_15_rx_fastbond_wren                                                                                                ( hssi_pldadapt_rx_15_rx_fastbond_wren),
   .hssi_pldadapt_rx_15_rx_fifo_power_mode                                                                                              ( hssi_pldadapt_rx_15_rx_fifo_power_mode),
   .hssi_pldadapt_rx_15_rx_fifo_read_latency_adjust                                                                                     ( hssi_pldadapt_rx_15_rx_fifo_read_latency_adjust),
   .hssi_pldadapt_rx_15_rx_fifo_write_ctrl                                                                                              ( hssi_pldadapt_rx_15_rx_fifo_write_ctrl),
   .hssi_pldadapt_rx_15_rx_fifo_write_latency_adjust                                                                                    ( hssi_pldadapt_rx_15_rx_fifo_write_latency_adjust),
   .hssi_pldadapt_rx_15_rx_osc_clock_setting                                                                                            ( hssi_pldadapt_rx_15_rx_osc_clock_setting),
   .hssi_pldadapt_rx_15_rx_pld_8g_eidleinfersel_polling_bypass                                                                          ( hssi_pldadapt_rx_15_rx_pld_8g_eidleinfersel_polling_bypass),
   .hssi_pldadapt_rx_15_rx_pld_pma_eye_monitor_polling_bypass                                                                           ( hssi_pldadapt_rx_15_rx_pld_pma_eye_monitor_polling_bypass),
   .hssi_pldadapt_rx_15_rx_pld_pma_pcie_switch_polling_bypass                                                                           ( hssi_pldadapt_rx_15_rx_pld_pma_pcie_switch_polling_bypass),
   .hssi_pldadapt_rx_15_rx_pld_pma_reser_out_polling_bypass                                                                             ( hssi_pldadapt_rx_15_rx_pld_pma_reser_out_polling_bypass),
   .hssi_pldadapt_rx_15_rx_prbs_flags_sr_enable                                                                                         ( hssi_pldadapt_rx_15_rx_prbs_flags_sr_enable),
   .hssi_pldadapt_rx_15_rx_true_b2b                                                                                                     ( hssi_pldadapt_rx_15_rx_true_b2b),
   .hssi_pldadapt_rx_15_rx_usertest_sel                                                                                                 ( hssi_pldadapt_rx_15_rx_usertest_sel),
   .hssi_pldadapt_rx_15_rxfifo_empty                                                                                                    ( hssi_pldadapt_rx_15_rxfifo_empty),
   .hssi_pldadapt_rx_15_rxfifo_full                                                                                                     ( hssi_pldadapt_rx_15_rxfifo_full),
   .hssi_pldadapt_rx_15_rxfifo_mode                                                                                                     ( hssi_pldadapt_rx_15_rxfifo_mode),
   .hssi_pldadapt_rx_15_rxfifo_pempty                                                                                                   ( hssi_pldadapt_rx_15_rxfifo_pempty),
   .hssi_pldadapt_rx_15_rxfifo_pfull                                                                                                    ( hssi_pldadapt_rx_15_rxfifo_pfull),
   .hssi_pldadapt_rx_15_rxfiford_post_ct_sel                                                                                            ( hssi_pldadapt_rx_15_rxfiford_post_ct_sel),
   .hssi_pldadapt_rx_15_rxfifowr_post_ct_sel                                                                                            ( hssi_pldadapt_rx_15_rxfifowr_post_ct_sel),
   .hssi_pldadapt_rx_15_sclk_sel                                                                                                        ( hssi_pldadapt_rx_15_sclk_sel),
   .hssi_pldadapt_rx_15_hdpldadapt_speed_grade                                                                                          ( hssi_pldadapt_rx_15_hdpldadapt_speed_grade),
   .hssi_pldadapt_rx_15_hdpldadapt_sr_sr_testbus_sel                                                                                    ( hssi_pldadapt_rx_15_hdpldadapt_sr_sr_testbus_sel),
   .hssi_pldadapt_rx_15_stretch_num_stages                                                                                              ( hssi_pldadapt_rx_15_stretch_num_stages),
   .hssi_pldadapt_rx_15_sup_mode                                                                                                        ( hssi_pldadapt_rx_15_sup_mode),
   .hssi_pldadapt_rx_15_txfiford_post_ct_sel                                                                                            ( hssi_pldadapt_rx_15_txfiford_post_ct_sel),
   .hssi_pldadapt_rx_15_txfifowr_post_ct_sel                                                                                            ( hssi_pldadapt_rx_15_txfifowr_post_ct_sel),
   .hssi_pldadapt_rx_15_us_bypass_pipeln                                                                                                ( hssi_pldadapt_rx_15_us_bypass_pipeln),
   .hssi_pldadapt_rx_15_us_last_chnl                                                                                                    ( hssi_pldadapt_rx_15_us_last_chnl),
   .hssi_pldadapt_rx_15_us_master                                                                                                       ( hssi_pldadapt_rx_15_us_master),
   .hssi_pldadapt_rx_15_word_align                                                                                                      ( hssi_pldadapt_rx_15_word_align),
   .hssi_pldadapt_rx_15_word_align_enable                                                                                               ( hssi_pldadapt_rx_15_word_align_enable),
   .hssi_pldadapt_rx_15_silicon_rev                                                                                                     ( hssi_pldadapt_rx_15_silicon_rev),
   .hssi_pldadapt_rx_15_reconfig_settings                                                                                               ( hssi_pldadapt_rx_15_reconfig_settings),
   .hssi_avmm1_if_15_pcs_arbiter_ctrl                                                                                                   ( hssi_avmm1_if_15_pcs_arbiter_ctrl),
   .hssi_avmm1_if_15_hssiadapt_avmm_clk_dcg_en                                                                                          ( hssi_avmm1_if_15_hssiadapt_avmm_clk_dcg_en),
   .hssi_avmm1_if_15_hssiadapt_avmm_clk_scg_en                                                                                          ( hssi_avmm1_if_15_hssiadapt_avmm_clk_scg_en),
   .hssi_avmm1_if_15_pldadapt_avmm_clk_scg_en                                                                                           ( hssi_avmm1_if_15_pldadapt_avmm_clk_scg_en),
   .hssi_avmm1_if_15_pcs_cal_done                                                                                                       ( hssi_avmm1_if_15_pcs_cal_done),
   .hssi_avmm1_if_15_pcs_cal_reserved                                                                                                   ( hssi_avmm1_if_15_pcs_cal_reserved),
   .hssi_avmm1_if_15_pcs_calibration_feature_en                                                                                         ( hssi_avmm1_if_15_pcs_calibration_feature_en),
   .hssi_avmm1_if_15_pldadapt_gate_dis                                                                                                  ( hssi_avmm1_if_15_pldadapt_gate_dis),
   .hssi_avmm1_if_15_pcs_hip_cal_en                                                                                                     ( hssi_avmm1_if_15_pcs_hip_cal_en),
   .hssi_avmm1_if_15_hssiadapt_nfhssi_calibratio_feature_en                                                                             ( hssi_avmm1_if_15_hssiadapt_nfhssi_calibratio_feature_en),
   .hssi_avmm1_if_15_pldadapt_nfhssi_calibratio_feature_en                                                                              ( hssi_avmm1_if_15_pldadapt_nfhssi_calibratio_feature_en),
   .hssi_avmm1_if_15_hssiadapt_osc_clk_scg_en                                                                                           ( hssi_avmm1_if_15_hssiadapt_osc_clk_scg_en),
   .hssi_avmm1_if_15_pldadapt_osc_clk_scg_en                                                                                            ( hssi_avmm1_if_15_pldadapt_osc_clk_scg_en),
   .hssi_avmm1_if_15_hssiadapt_read_blocking_enable                                                                                     ( hssi_avmm1_if_15_hssiadapt_read_blocking_enable),
   .hssi_avmm1_if_15_pldadapt_read_blocking_enable                                                                                      ( hssi_avmm1_if_15_pldadapt_read_blocking_enable),
   .hssi_avmm1_if_15_hssiadapt_uc_blocking_enable                                                                                       ( hssi_avmm1_if_15_hssiadapt_uc_blocking_enable),
   .hssi_avmm1_if_15_pldadapt_uc_blocking_enable                                                                                        ( hssi_avmm1_if_15_pldadapt_uc_blocking_enable),
   .hssi_avmm1_if_15_hssiadapt_write_resp_en                                                                                            ( hssi_avmm1_if_15_hssiadapt_write_resp_en),
   .hssi_avmm1_if_15_hssiadapt_avmm_osc_clock_setting                                                                                   ( hssi_avmm1_if_15_hssiadapt_avmm_osc_clock_setting),
   .hssi_avmm1_if_15_pldadapt_avmm_osc_clock_setting                                                                                    ( hssi_avmm1_if_15_pldadapt_avmm_osc_clock_setting),
   .hssi_avmm1_if_15_hssiadapt_avmm_testbus_sel                                                                                         ( hssi_avmm1_if_15_hssiadapt_avmm_testbus_sel),
   .hssi_avmm1_if_15_pldadapt_avmm_testbus_sel                                                                                          ( hssi_avmm1_if_15_pldadapt_avmm_testbus_sel),
   .hssi_avmm1_if_15_func_mode                                                                                                          ( hssi_avmm1_if_15_func_mode),
   .hssi_avmm1_if_15_hssiadapt_sr_hip_mode                                                                                              ( hssi_avmm1_if_15_hssiadapt_sr_hip_mode),
   .hssi_avmm1_if_15_hssiadapt_hip_mode                                                                                                 ( hssi_avmm1_if_15_hssiadapt_hip_mode),
   .hssi_avmm1_if_15_pldadapt_hip_mode                                                                                                  ( hssi_avmm1_if_15_pldadapt_hip_mode),
   .hssi_avmm1_if_15_hssiadapt_sr_powerdown_mode                                                                                        ( hssi_avmm1_if_15_hssiadapt_sr_powerdown_mode),
   .hssi_avmm1_if_15_hssiadapt_sr_sr_free_run_div_clk                                                                                   ( hssi_avmm1_if_15_hssiadapt_sr_sr_free_run_div_clk),
   .hssi_avmm1_if_15_hssiadapt_sr_sr_hip_en                                                                                             ( hssi_avmm1_if_15_hssiadapt_sr_sr_hip_en),
   .hssi_avmm1_if_15_hssiadapt_sr_sr_osc_clk_div_sel                                                                                    ( hssi_avmm1_if_15_hssiadapt_sr_sr_osc_clk_div_sel),
   .hssi_avmm1_if_15_hssiadapt_sr_sr_osc_clk_scg_en                                                                                     ( hssi_avmm1_if_15_hssiadapt_sr_sr_osc_clk_scg_en),
   .hssi_avmm1_if_15_hssiadapt_sr_sr_parity_en                                                                                          ( hssi_avmm1_if_15_hssiadapt_sr_sr_parity_en),
   .hssi_avmm1_if_15_hssiadapt_sr_sr_reserved_in_en                                                                                     ( hssi_avmm1_if_15_hssiadapt_sr_sr_reserved_in_en),
   .hssi_avmm1_if_15_hssiadapt_sr_sr_reserved_out_en                                                                                    ( hssi_avmm1_if_15_hssiadapt_sr_sr_reserved_out_en),
   .hssi_avmm1_if_15_hssiadapt_sr_sup_mode                                                                                              ( hssi_avmm1_if_15_hssiadapt_sr_sup_mode),
   .hssi_avmm1_if_15_topology                                                                                                           ( hssi_avmm1_if_15_topology),
   .hssi_avmm1_if_15_silicon_rev                                                                                                        ( hssi_avmm1_if_15_silicon_rev),
   .hssi_avmm1_if_15_calibration_type                                                                                                   ( hssi_avmm1_if_15_calibration_type),
   .hssi_avmm2_if_15_pcs_arbiter_ctrl                                                                                                   ( hssi_avmm2_if_15_pcs_arbiter_ctrl),
   .hssi_avmm2_if_15_hssiadapt_avmm_clk_dcg_en                                                                                          ( hssi_avmm2_if_15_hssiadapt_avmm_clk_dcg_en),
   .hssi_avmm2_if_15_hssiadapt_avmm_clk_scg_en                                                                                          ( hssi_avmm2_if_15_hssiadapt_avmm_clk_scg_en),
   .hssi_avmm2_if_15_pldadapt_avmm_clk_scg_en                                                                                           ( hssi_avmm2_if_15_pldadapt_avmm_clk_scg_en),
   .hssi_avmm2_if_15_pcs_cal_done                                                                                                       ( hssi_avmm2_if_15_pcs_cal_done),
   .hssi_avmm2_if_15_pcs_cal_reserved                                                                                                   ( hssi_avmm2_if_15_pcs_cal_reserved),
   .hssi_avmm2_if_15_pcs_calibration_feature_en                                                                                         ( hssi_avmm2_if_15_pcs_calibration_feature_en),
   .hssi_avmm2_if_15_pldadapt_gate_dis                                                                                                  ( hssi_avmm2_if_15_pldadapt_gate_dis),
   .hssi_avmm2_if_15_pcs_hip_cal_en                                                                                                     ( hssi_avmm2_if_15_pcs_hip_cal_en),
   .hssi_avmm2_if_15_hssiadapt_osc_clk_scg_en                                                                                           ( hssi_avmm2_if_15_hssiadapt_osc_clk_scg_en),
   .hssi_avmm2_if_15_pldadapt_osc_clk_scg_en                                                                                            ( hssi_avmm2_if_15_pldadapt_osc_clk_scg_en),
   .hssi_avmm2_if_15_hssiadapt_avmm_osc_clock_setting                                                                                   ( hssi_avmm2_if_15_hssiadapt_avmm_osc_clock_setting),
   .hssi_avmm2_if_15_pldadapt_avmm_osc_clock_setting                                                                                    ( hssi_avmm2_if_15_pldadapt_avmm_osc_clock_setting),
   .hssi_avmm2_if_15_hssiadapt_avmm_testbus_sel                                                                                         ( hssi_avmm2_if_15_hssiadapt_avmm_testbus_sel),
   .hssi_avmm2_if_15_pldadapt_avmm_testbus_sel                                                                                          ( hssi_avmm2_if_15_pldadapt_avmm_testbus_sel),
   .hssi_avmm2_if_15_func_mode                                                                                                          ( hssi_avmm2_if_15_func_mode),
   .hssi_avmm2_if_15_hssiadapt_hip_mode                                                                                                 ( hssi_avmm2_if_15_hssiadapt_hip_mode),
   .hssi_avmm2_if_15_pldadapt_hip_mode                                                                                                  ( hssi_avmm2_if_15_pldadapt_hip_mode),
   .hssi_avmm2_if_15_topology                                                                                                           ( hssi_avmm2_if_15_topology),
   .hssi_avmm2_if_15_silicon_rev                                                                                                        ( hssi_avmm2_if_15_silicon_rev),
   .hssi_avmm2_if_15_calibration_type                                                                                                   ( hssi_avmm2_if_15_calibration_type),
   .hssi_aibnd_rx_23_aib_ber_margining_ctrl                                                                                             ( hssi_aibnd_rx_23_aib_ber_margining_ctrl),
   .hssi_aibnd_rx_23_aib_datasel_gr0                                                                                                    ( hssi_aibnd_rx_23_aib_datasel_gr0),
   .hssi_aibnd_rx_23_aib_datasel_gr1                                                                                                    ( hssi_aibnd_rx_23_aib_datasel_gr1),
   .hssi_aibnd_rx_23_aib_datasel_gr2                                                                                                    ( hssi_aibnd_rx_23_aib_datasel_gr2),
   .hssi_aibnd_rx_23_aib_dllstr_align_clkdiv                                                                                            ( hssi_aibnd_rx_23_aib_dllstr_align_clkdiv),
   .hssi_aibnd_rx_23_aib_dllstr_align_dly_pst                                                                                           ( hssi_aibnd_rx_23_aib_dllstr_align_dly_pst),
   .hssi_aibnd_rx_23_aib_dllstr_align_dy_ctl_static                                                                                     ( hssi_aibnd_rx_23_aib_dllstr_align_dy_ctl_static),
   .hssi_aibnd_rx_23_aib_dllstr_align_dy_ctlsel                                                                                         ( hssi_aibnd_rx_23_aib_dllstr_align_dy_ctlsel),
   .hssi_aibnd_rx_23_aib_dllstr_align_entest                                                                                            ( hssi_aibnd_rx_23_aib_dllstr_align_entest),
   .hssi_aibnd_rx_23_aib_dllstr_align_halfcode                                                                                          ( hssi_aibnd_rx_23_aib_dllstr_align_halfcode),
   .hssi_aibnd_rx_23_aib_dllstr_align_selflock                                                                                          ( hssi_aibnd_rx_23_aib_dllstr_align_selflock),
   .hssi_aibnd_rx_23_aib_dllstr_align_st_core_dn_prgmnvrt                                                                               ( hssi_aibnd_rx_23_aib_dllstr_align_st_core_dn_prgmnvrt),
   .hssi_aibnd_rx_23_aib_dllstr_align_st_core_up_prgmnvrt                                                                               ( hssi_aibnd_rx_23_aib_dllstr_align_st_core_up_prgmnvrt),
   .hssi_aibnd_rx_23_aib_dllstr_align_st_core_updnen                                                                                    ( hssi_aibnd_rx_23_aib_dllstr_align_st_core_updnen),
   .hssi_aibnd_rx_23_aib_dllstr_align_st_dftmuxsel                                                                                      ( hssi_aibnd_rx_23_aib_dllstr_align_st_dftmuxsel),
   .hssi_aibnd_rx_23_aib_dllstr_align_st_en                                                                                             ( hssi_aibnd_rx_23_aib_dllstr_align_st_en),
   .hssi_aibnd_rx_23_aib_dllstr_align_st_hps_ctrl_en                                                                                    ( hssi_aibnd_rx_23_aib_dllstr_align_st_hps_ctrl_en),
   .hssi_aibnd_rx_23_aib_dllstr_align_st_lockreq_muxsel                                                                                 ( hssi_aibnd_rx_23_aib_dllstr_align_st_lockreq_muxsel),
   .hssi_aibnd_rx_23_aib_dllstr_align_st_new_dll                                                                                        ( hssi_aibnd_rx_23_aib_dllstr_align_st_new_dll),
   .hssi_aibnd_rx_23_aib_dllstr_align_st_rst                                                                                            ( hssi_aibnd_rx_23_aib_dllstr_align_st_rst),
   .hssi_aibnd_rx_23_aib_dllstr_align_st_rst_prgmnvrt                                                                                   ( hssi_aibnd_rx_23_aib_dllstr_align_st_rst_prgmnvrt),
   .hssi_aibnd_rx_23_aib_dllstr_align_test_clk_pll_en_n                                                                                 ( hssi_aibnd_rx_23_aib_dllstr_align_test_clk_pll_en_n),
   .hssi_aibnd_rx_23_aib_inctrl_gr0                                                                                                     ( hssi_aibnd_rx_23_aib_inctrl_gr0),
   .hssi_aibnd_rx_23_aib_inctrl_gr1                                                                                                     ( hssi_aibnd_rx_23_aib_inctrl_gr1),
   .hssi_aibnd_rx_23_aib_inctrl_gr2                                                                                                     ( hssi_aibnd_rx_23_aib_inctrl_gr2),
   .hssi_aibnd_rx_23_aib_inctrl_gr3                                                                                                     ( hssi_aibnd_rx_23_aib_inctrl_gr3),
   .hssi_aibnd_rx_23_aib_outctrl_gr0                                                                                                    ( hssi_aibnd_rx_23_aib_outctrl_gr0),
   .hssi_aibnd_rx_23_aib_outctrl_gr1                                                                                                    ( hssi_aibnd_rx_23_aib_outctrl_gr1),
   .hssi_aibnd_rx_23_aib_outctrl_gr2                                                                                                    ( hssi_aibnd_rx_23_aib_outctrl_gr2),
   .hssi_aibnd_rx_23_aib_outndrv_r12                                                                                                    ( hssi_aibnd_rx_23_aib_outndrv_r12),
   .hssi_aibnd_rx_23_aib_outndrv_r34                                                                                                    ( hssi_aibnd_rx_23_aib_outndrv_r34),
   .hssi_aibnd_rx_23_aib_outndrv_r56                                                                                                    ( hssi_aibnd_rx_23_aib_outndrv_r56),
   .hssi_aibnd_rx_23_aib_outndrv_r78                                                                                                    ( hssi_aibnd_rx_23_aib_outndrv_r78),
   .hssi_aibnd_rx_23_aib_outpdrv_r12                                                                                                    ( hssi_aibnd_rx_23_aib_outpdrv_r12),
   .hssi_aibnd_rx_23_aib_outpdrv_r34                                                                                                    ( hssi_aibnd_rx_23_aib_outpdrv_r34),
   .hssi_aibnd_rx_23_aib_outpdrv_r56                                                                                                    ( hssi_aibnd_rx_23_aib_outpdrv_r56),
   .hssi_aibnd_rx_23_aib_outpdrv_r78                                                                                                    ( hssi_aibnd_rx_23_aib_outpdrv_r78),
   .hssi_aibnd_rx_23_aib_red_shift_en                                                                                                   ( hssi_aibnd_rx_23_aib_red_shift_en),
   .hssi_aibnd_rx_23_dft_hssitestip_dll_dcc_en                                                                                          ( hssi_aibnd_rx_23_dft_hssitestip_dll_dcc_en),
   .hssi_aibnd_rx_23_op_mode                                                                                                            ( hssi_aibnd_rx_23_op_mode),
   .hssi_aibnd_rx_23_powerdown_mode                                                                                                     ( hssi_aibnd_rx_23_powerdown_mode),
   .hssi_aibnd_rx_23_powermode_ac                                                                                                       ( hssi_aibnd_rx_23_powermode_ac),
   .hssi_aibnd_rx_23_powermode_dc                                                                                                       ( hssi_aibnd_rx_23_powermode_dc),
   .hssi_aibnd_rx_23_powermode_freq_hz_aib_hssi_rx_transfer_clk                                                                         ( hssi_aibnd_rx_23_powermode_freq_hz_aib_hssi_rx_transfer_clk),
   .hssi_aibnd_rx_23_redundancy_en                                                                                                      ( hssi_aibnd_rx_23_redundancy_en),
   .hssi_aibnd_rx_23_sup_mode                                                                                                           ( hssi_aibnd_rx_23_sup_mode),
   .hssi_aibnd_rx_23_silicon_rev                                                                                                        ( hssi_aibnd_rx_23_silicon_rev),
   .hssi_aibnd_tx_23_aib_datasel_gr0                                                                                                    ( hssi_aibnd_tx_23_aib_datasel_gr0),
   .hssi_aibnd_tx_23_aib_datasel_gr1                                                                                                    ( hssi_aibnd_tx_23_aib_datasel_gr1),
   .hssi_aibnd_tx_23_aib_datasel_gr2                                                                                                    ( hssi_aibnd_tx_23_aib_datasel_gr2),
   .hssi_aibnd_tx_23_aib_datasel_gr3                                                                                                    ( hssi_aibnd_tx_23_aib_datasel_gr3),
   .hssi_aibnd_tx_23_aib_ddrctrl_gr0                                                                                                    ( hssi_aibnd_tx_23_aib_ddrctrl_gr0),
   .hssi_aibnd_tx_23_aib_hssi_tx_transfer_clk_hz                                                                                        ( hssi_aibnd_tx_23_aib_hssi_tx_transfer_clk_hz),
   .hssi_aibnd_tx_23_aib_iinasyncen                                                                                                     ( hssi_aibnd_tx_23_aib_iinasyncen),
   .hssi_aibnd_tx_23_aib_iinclken                                                                                                       ( hssi_aibnd_tx_23_aib_iinclken),
   .hssi_aibnd_tx_23_aib_outctrl_gr0                                                                                                    ( hssi_aibnd_tx_23_aib_outctrl_gr0),
   .hssi_aibnd_tx_23_aib_outctrl_gr1                                                                                                    ( hssi_aibnd_tx_23_aib_outctrl_gr1),
   .hssi_aibnd_tx_23_aib_outctrl_gr2                                                                                                    ( hssi_aibnd_tx_23_aib_outctrl_gr2),
   .hssi_aibnd_tx_23_aib_outctrl_gr3                                                                                                    ( hssi_aibnd_tx_23_aib_outctrl_gr3),
   .hssi_aibnd_tx_23_aib_outndrv_r34                                                                                                    ( hssi_aibnd_tx_23_aib_outndrv_r34),
   .hssi_aibnd_tx_23_aib_outndrv_r56                                                                                                    ( hssi_aibnd_tx_23_aib_outndrv_r56),
   .hssi_aibnd_tx_23_aib_outpdrv_r34                                                                                                    ( hssi_aibnd_tx_23_aib_outpdrv_r34),
   .hssi_aibnd_tx_23_aib_outpdrv_r56                                                                                                    ( hssi_aibnd_tx_23_aib_outpdrv_r56),
   .hssi_aibnd_tx_23_aib_red_dirclkn_shiften                                                                                            ( hssi_aibnd_tx_23_aib_red_dirclkn_shiften),
   .hssi_aibnd_tx_23_aib_red_dirclkp_shiften                                                                                            ( hssi_aibnd_tx_23_aib_red_dirclkp_shiften),
   .hssi_aibnd_tx_23_aib_red_drx_shiften                                                                                                ( hssi_aibnd_tx_23_aib_red_drx_shiften),
   .hssi_aibnd_tx_23_aib_red_dtx_shiften                                                                                                ( hssi_aibnd_tx_23_aib_red_dtx_shiften),
   .hssi_aibnd_tx_23_aib_red_pout_shiften                                                                                               ( hssi_aibnd_tx_23_aib_red_pout_shiften),
   .hssi_aibnd_tx_23_aib_red_rx_shiften                                                                                                 ( hssi_aibnd_tx_23_aib_red_rx_shiften),
   .hssi_aibnd_tx_23_aib_red_tx_shiften                                                                                                 ( hssi_aibnd_tx_23_aib_red_tx_shiften),
   .hssi_aibnd_tx_23_aib_red_txferclkout_shiften                                                                                        ( hssi_aibnd_tx_23_aib_red_txferclkout_shiften),
   .hssi_aibnd_tx_23_aib_red_txferclkoutn_shiften                                                                                       ( hssi_aibnd_tx_23_aib_red_txferclkoutn_shiften),
   .hssi_aibnd_tx_23_aib_tx_clkdiv                                                                                                      ( hssi_aibnd_tx_23_aib_tx_clkdiv),
   .hssi_aibnd_tx_23_aib_tx_dcc_byp                                                                                                     ( hssi_aibnd_tx_23_aib_tx_dcc_byp),
   .hssi_aibnd_tx_23_aib_tx_dcc_byp_iocsr_unused                                                                                        ( hssi_aibnd_tx_23_aib_tx_dcc_byp_iocsr_unused),
   .hssi_aibnd_tx_23_aib_tx_dcc_cont_cal                                                                                                ( hssi_aibnd_tx_23_aib_tx_dcc_cont_cal),
   .hssi_aibnd_tx_23_aib_tx_dcc_cont_cal_iocsr_unused                                                                                   ( hssi_aibnd_tx_23_aib_tx_dcc_cont_cal_iocsr_unused),
   .hssi_aibnd_tx_23_aib_tx_dcc_dft                                                                                                     ( hssi_aibnd_tx_23_aib_tx_dcc_dft),
   .hssi_aibnd_tx_23_aib_tx_dcc_dft_sel                                                                                                 ( hssi_aibnd_tx_23_aib_tx_dcc_dft_sel),
   .hssi_aibnd_tx_23_aib_tx_dcc_dll_dft_sel                                                                                             ( hssi_aibnd_tx_23_aib_tx_dcc_dll_dft_sel),
   .hssi_aibnd_tx_23_aib_tx_dcc_dll_entest                                                                                              ( hssi_aibnd_tx_23_aib_tx_dcc_dll_entest),
   .hssi_aibnd_tx_23_aib_tx_dcc_dy_ctl_static                                                                                           ( hssi_aibnd_tx_23_aib_tx_dcc_dy_ctl_static),
   .hssi_aibnd_tx_23_aib_tx_dcc_dy_ctlsel                                                                                               ( hssi_aibnd_tx_23_aib_tx_dcc_dy_ctlsel),
   .hssi_aibnd_tx_23_aib_tx_dcc_en                                                                                                      ( hssi_aibnd_tx_23_aib_tx_dcc_en),
   .hssi_aibnd_tx_23_aib_tx_dcc_en_iocsr_unused                                                                                         ( hssi_aibnd_tx_23_aib_tx_dcc_en_iocsr_unused),
   .hssi_aibnd_tx_23_aib_tx_dcc_manual_dn                                                                                               ( hssi_aibnd_tx_23_aib_tx_dcc_manual_dn),
   .hssi_aibnd_tx_23_aib_tx_dcc_manual_up                                                                                               ( hssi_aibnd_tx_23_aib_tx_dcc_manual_up),
   .hssi_aibnd_tx_23_aib_tx_dcc_rst_prgmnvrt                                                                                            ( hssi_aibnd_tx_23_aib_tx_dcc_rst_prgmnvrt),
   .hssi_aibnd_tx_23_aib_tx_dcc_st_core_dn_prgmnvrt                                                                                     ( hssi_aibnd_tx_23_aib_tx_dcc_st_core_dn_prgmnvrt),
   .hssi_aibnd_tx_23_aib_tx_dcc_st_core_up_prgmnvrt                                                                                     ( hssi_aibnd_tx_23_aib_tx_dcc_st_core_up_prgmnvrt),
   .hssi_aibnd_tx_23_aib_tx_dcc_st_core_updnen                                                                                          ( hssi_aibnd_tx_23_aib_tx_dcc_st_core_updnen),
   .hssi_aibnd_tx_23_aib_tx_dcc_st_dftmuxsel                                                                                            ( hssi_aibnd_tx_23_aib_tx_dcc_st_dftmuxsel),
   .hssi_aibnd_tx_23_aib_tx_dcc_st_dly_pst                                                                                              ( hssi_aibnd_tx_23_aib_tx_dcc_st_dly_pst),
   .hssi_aibnd_tx_23_aib_tx_dcc_st_en                                                                                                   ( hssi_aibnd_tx_23_aib_tx_dcc_st_en),
   .hssi_aibnd_tx_23_aib_tx_dcc_st_hps_ctrl_en                                                                                          ( hssi_aibnd_tx_23_aib_tx_dcc_st_hps_ctrl_en),
   .hssi_aibnd_tx_23_aib_tx_dcc_st_lockreq_muxsel                                                                                       ( hssi_aibnd_tx_23_aib_tx_dcc_st_lockreq_muxsel),
   .hssi_aibnd_tx_23_aib_tx_dcc_st_new_dll                                                                                              ( hssi_aibnd_tx_23_aib_tx_dcc_st_new_dll),
   .hssi_aibnd_tx_23_aib_tx_dcc_st_rst                                                                                                  ( hssi_aibnd_tx_23_aib_tx_dcc_st_rst),
   .hssi_aibnd_tx_23_aib_tx_dcc_test_clk_pll_en_n                                                                                       ( hssi_aibnd_tx_23_aib_tx_dcc_test_clk_pll_en_n),
   .hssi_aibnd_tx_23_aib_tx_halfcode                                                                                                    ( hssi_aibnd_tx_23_aib_tx_halfcode),
   .hssi_aibnd_tx_23_aib_tx_selflock                                                                                                    ( hssi_aibnd_tx_23_aib_tx_selflock),
   .hssi_aibnd_tx_23_dfd_dll_dcc_en                                                                                                     ( hssi_aibnd_tx_23_dfd_dll_dcc_en),
   .hssi_aibnd_tx_23_dft_hssitestip_dll_dcc_en                                                                                          ( hssi_aibnd_tx_23_dft_hssitestip_dll_dcc_en),
   .hssi_aibnd_tx_23_op_mode                                                                                                            ( hssi_aibnd_tx_23_op_mode),
   .hssi_aibnd_tx_23_powerdown_mode                                                                                                     ( hssi_aibnd_tx_23_powerdown_mode),
   .hssi_aibnd_tx_23_powermode_ac                                                                                                       ( hssi_aibnd_tx_23_powermode_ac),
   .hssi_aibnd_tx_23_powermode_dc                                                                                                       ( hssi_aibnd_tx_23_powermode_dc),
   .hssi_aibnd_tx_23_powermode_freq_hz_aib_hssi_tx_transfer_clk                                                                         ( hssi_aibnd_tx_23_powermode_freq_hz_aib_hssi_tx_transfer_clk),
   .hssi_aibnd_tx_23_redundancy_en                                                                                                      ( hssi_aibnd_tx_23_redundancy_en),
   .hssi_aibnd_tx_23_sup_mode                                                                                                           ( hssi_aibnd_tx_23_sup_mode),
   .hssi_aibnd_tx_23_silicon_rev                                                                                                        ( hssi_aibnd_tx_23_silicon_rev),
   .hssi_pldadapt_tx_23_aib_clk1_sel                                                                                                    ( hssi_pldadapt_tx_23_aib_clk1_sel),
   .hssi_pldadapt_tx_23_aib_clk2_sel                                                                                                    ( hssi_pldadapt_tx_23_aib_clk2_sel),
   .hssi_pldadapt_tx_23_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                           ( hssi_pldadapt_tx_23_hdpldadapt_aib_fabric_pld_pma_hclk_hz),
   .hssi_pldadapt_tx_23_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz                                                                         ( hssi_pldadapt_tx_23_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz),
   .hssi_pldadapt_tx_23_hdpldadapt_aib_fabric_tx_sr_clk_in_hz                                                                           ( hssi_pldadapt_tx_23_hdpldadapt_aib_fabric_tx_sr_clk_in_hz),
   .hssi_pldadapt_tx_23_bonding_dft_en                                                                                                  ( hssi_pldadapt_tx_23_bonding_dft_en),
   .hssi_pldadapt_tx_23_bonding_dft_val                                                                                                 ( hssi_pldadapt_tx_23_bonding_dft_val),
   .hssi_pldadapt_tx_23_chnl_bonding                                                                                                    ( hssi_pldadapt_tx_23_chnl_bonding),
   .hssi_pldadapt_tx_23_comp_cnt                                                                                                        ( hssi_pldadapt_tx_23_comp_cnt),
   .hssi_pldadapt_tx_23_compin_sel                                                                                                      ( hssi_pldadapt_tx_23_compin_sel),
   .hssi_pldadapt_tx_23_hdpldadapt_csr_clk_hz                                                                                           ( hssi_pldadapt_tx_23_hdpldadapt_csr_clk_hz),
   .hssi_pldadapt_tx_23_ctrl_plane_bonding                                                                                              ( hssi_pldadapt_tx_23_ctrl_plane_bonding),
   .hssi_pldadapt_tx_23_ds_bypass_pipeln                                                                                                ( hssi_pldadapt_tx_23_ds_bypass_pipeln),
   .hssi_pldadapt_tx_23_ds_last_chnl                                                                                                    ( hssi_pldadapt_tx_23_ds_last_chnl),
   .hssi_pldadapt_tx_23_ds_master                                                                                                       ( hssi_pldadapt_tx_23_ds_master),
   .hssi_pldadapt_tx_23_duplex_mode                                                                                                     ( hssi_pldadapt_tx_23_duplex_mode),
   .hssi_pldadapt_tx_23_dv_bond                                                                                                         ( hssi_pldadapt_tx_23_dv_bond),
   .hssi_pldadapt_tx_23_dv_gen                                                                                                          ( hssi_pldadapt_tx_23_dv_gen),
   .hssi_pldadapt_tx_23_fifo_double_write                                                                                               ( hssi_pldadapt_tx_23_fifo_double_write),
   .hssi_pldadapt_tx_23_fifo_mode                                                                                                       ( hssi_pldadapt_tx_23_fifo_mode),
   .hssi_pldadapt_tx_23_fifo_rd_clk_frm_gen_scg_en                                                                                      ( hssi_pldadapt_tx_23_fifo_rd_clk_frm_gen_scg_en),
   .hssi_pldadapt_tx_23_fifo_rd_clk_scg_en                                                                                              ( hssi_pldadapt_tx_23_fifo_rd_clk_scg_en),
   .hssi_pldadapt_tx_23_fifo_rd_clk_sel                                                                                                 ( hssi_pldadapt_tx_23_fifo_rd_clk_sel),
   .hssi_pldadapt_tx_23_fifo_stop_rd                                                                                                    ( hssi_pldadapt_tx_23_fifo_stop_rd),
   .hssi_pldadapt_tx_23_fifo_stop_wr                                                                                                    ( hssi_pldadapt_tx_23_fifo_stop_wr),
   .hssi_pldadapt_tx_23_fifo_width                                                                                                      ( hssi_pldadapt_tx_23_fifo_width),
   .hssi_pldadapt_tx_23_fifo_wr_clk_scg_en                                                                                              ( hssi_pldadapt_tx_23_fifo_wr_clk_scg_en),
   .hssi_pldadapt_tx_23_fpll_shared_direct_async_in_sel                                                                                 ( hssi_pldadapt_tx_23_fpll_shared_direct_async_in_sel),
   .hssi_pldadapt_tx_23_frmgen_burst                                                                                                    ( hssi_pldadapt_tx_23_frmgen_burst),
   .hssi_pldadapt_tx_23_frmgen_bypass                                                                                                   ( hssi_pldadapt_tx_23_frmgen_bypass),
   .hssi_pldadapt_tx_23_frmgen_mfrm_length                                                                                              ( hssi_pldadapt_tx_23_frmgen_mfrm_length),
   .hssi_pldadapt_tx_23_frmgen_pipeln                                                                                                   ( hssi_pldadapt_tx_23_frmgen_pipeln),
   .hssi_pldadapt_tx_23_frmgen_pyld_ins                                                                                                 ( hssi_pldadapt_tx_23_frmgen_pyld_ins),
   .hssi_pldadapt_tx_23_frmgen_wordslip                                                                                                 ( hssi_pldadapt_tx_23_frmgen_wordslip),
   .hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit0_rst_val                                                                                     ( hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit0_rst_val),
   .hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit1_rst_val                                                                                     ( hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit1_rst_val),
   .hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit2_rst_val                                                                                     ( hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit2_rst_val),
   .hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit3_rst_val                                                                                     ( hssi_pldadapt_tx_23_fsr_hip_fsr_in_bit3_rst_val),
   .hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit0_rst_val                                                                                    ( hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit0_rst_val),
   .hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit1_rst_val                                                                                    ( hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit1_rst_val),
   .hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit2_rst_val                                                                                    ( hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit2_rst_val),
   .hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit3_rst_val                                                                                    ( hssi_pldadapt_tx_23_fsr_hip_fsr_out_bit3_rst_val),
   .hssi_pldadapt_tx_23_fsr_mask_tx_pll_rst_val                                                                                         ( hssi_pldadapt_tx_23_fsr_mask_tx_pll_rst_val),
   .hssi_pldadapt_tx_23_fsr_pld_txelecidle_rst_val                                                                                      ( hssi_pldadapt_tx_23_fsr_pld_txelecidle_rst_val),
   .hssi_pldadapt_tx_23_gb_tx_idwidth                                                                                                   ( hssi_pldadapt_tx_23_gb_tx_idwidth),
   .hssi_pldadapt_tx_23_gb_tx_odwidth                                                                                                   ( hssi_pldadapt_tx_23_gb_tx_odwidth),
   .hssi_pldadapt_tx_23_hip_mode                                                                                                        ( hssi_pldadapt_tx_23_hip_mode),
   .hssi_pldadapt_tx_23_hip_osc_clk_scg_en                                                                                              ( hssi_pldadapt_tx_23_hip_osc_clk_scg_en),
   .hssi_pldadapt_tx_23_hrdrst_dcd_cal_done_bypass                                                                                      ( hssi_pldadapt_tx_23_hrdrst_dcd_cal_done_bypass),
   .hssi_pldadapt_tx_23_hrdrst_rst_sm_dis                                                                                               ( hssi_pldadapt_tx_23_hrdrst_rst_sm_dis),
   .hssi_pldadapt_tx_23_hrdrst_rx_osc_clk_scg_en                                                                                        ( hssi_pldadapt_tx_23_hrdrst_rx_osc_clk_scg_en),
   .hssi_pldadapt_tx_23_hrdrst_user_ctl_en                                                                                              ( hssi_pldadapt_tx_23_hrdrst_user_ctl_en),
   .hssi_pldadapt_tx_23_indv                                                                                                            ( hssi_pldadapt_tx_23_indv),
   .hssi_pldadapt_tx_23_is_paired_with                                                                                                  ( hssi_pldadapt_tx_23_is_paired_with),
   .hssi_pldadapt_tx_23_loopback_mode                                                                                                   ( hssi_pldadapt_tx_23_loopback_mode),
   .hssi_pldadapt_tx_23_low_latency_en                                                                                                  ( hssi_pldadapt_tx_23_low_latency_en),
   .hssi_pldadapt_tx_23_osc_clk_scg_en                                                                                                  ( hssi_pldadapt_tx_23_osc_clk_scg_en),
   .hssi_pldadapt_tx_23_phcomp_rd_del                                                                                                   ( hssi_pldadapt_tx_23_phcomp_rd_del),
   .hssi_pldadapt_tx_23_pipe_mode                                                                                                       ( hssi_pldadapt_tx_23_pipe_mode),
   .hssi_pldadapt_tx_23_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                              ( hssi_pldadapt_tx_23_hdpldadapt_pld_avmm1_clk_rowclk_hz),
   .hssi_pldadapt_tx_23_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                              ( hssi_pldadapt_tx_23_hdpldadapt_pld_avmm2_clk_rowclk_hz),
   .hssi_pldadapt_tx_23_pld_clk1_delay_en                                                                                               ( hssi_pldadapt_tx_23_pld_clk1_delay_en),
   .hssi_pldadapt_tx_23_pld_clk1_delay_sel                                                                                              ( hssi_pldadapt_tx_23_pld_clk1_delay_sel),
   .hssi_pldadapt_tx_23_pld_clk1_inv_en                                                                                                 ( hssi_pldadapt_tx_23_pld_clk1_inv_en),
   .hssi_pldadapt_tx_23_pld_clk1_sel                                                                                                    ( hssi_pldadapt_tx_23_pld_clk1_sel),
   .hssi_pldadapt_tx_23_pld_clk2_sel                                                                                                    ( hssi_pldadapt_tx_23_pld_clk2_sel),
   .hssi_pldadapt_tx_23_hdpldadapt_pld_sclk1_rowclk_hz                                                                                  ( hssi_pldadapt_tx_23_hdpldadapt_pld_sclk1_rowclk_hz),
   .hssi_pldadapt_tx_23_hdpldadapt_pld_sclk2_rowclk_hz                                                                                  ( hssi_pldadapt_tx_23_hdpldadapt_pld_sclk2_rowclk_hz),
   .hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk1_dcm_hz                                                                                   ( hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk1_dcm_hz),
   .hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk1_rowclk_hz                                                                                ( hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk1_rowclk_hz),
   .hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk2_dcm_hz                                                                                   ( hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk2_dcm_hz),
   .hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk2_rowclk_hz                                                                                ( hssi_pldadapt_tx_23_hdpldadapt_pld_tx_clk2_rowclk_hz),
   .hssi_pldadapt_tx_23_pma_aib_tx_clk_expected_setting                                                                                 ( hssi_pldadapt_tx_23_pma_aib_tx_clk_expected_setting),
   .hssi_pldadapt_tx_23_powerdown_mode                                                                                                  ( hssi_pldadapt_tx_23_powerdown_mode),
   .hssi_pldadapt_tx_23_powermode_dc                                                                                                    ( hssi_pldadapt_tx_23_powermode_dc),
   .hssi_pldadapt_tx_23_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                       ( hssi_pldadapt_tx_23_powermode_freq_hz_aib_fabric_rx_sr_clk_in),
   .hssi_pldadapt_tx_23_powermode_freq_hz_pld_tx_clk1_dcm                                                                               ( hssi_pldadapt_tx_23_powermode_freq_hz_pld_tx_clk1_dcm),
   .hssi_pldadapt_tx_23_sh_err                                                                                                          ( hssi_pldadapt_tx_23_sh_err),
   .hssi_pldadapt_tx_23_hdpldadapt_speed_grade                                                                                          ( hssi_pldadapt_tx_23_hdpldadapt_speed_grade),
   .hssi_pldadapt_tx_23_hdpldadapt_sr_sr_testbus_sel                                                                                    ( hssi_pldadapt_tx_23_hdpldadapt_sr_sr_testbus_sel),
   .hssi_pldadapt_tx_23_stretch_num_stages                                                                                              ( hssi_pldadapt_tx_23_stretch_num_stages),
   .hssi_pldadapt_tx_23_sup_mode                                                                                                        ( hssi_pldadapt_tx_23_sup_mode),
   .hssi_pldadapt_tx_23_tx_datapath_tb_sel                                                                                              ( hssi_pldadapt_tx_23_tx_datapath_tb_sel),
   .hssi_pldadapt_tx_23_tx_fastbond_rden                                                                                                ( hssi_pldadapt_tx_23_tx_fastbond_rden),
   .hssi_pldadapt_tx_23_tx_fastbond_wren                                                                                                ( hssi_pldadapt_tx_23_tx_fastbond_wren),
   .hssi_pldadapt_tx_23_tx_fifo_power_mode                                                                                              ( hssi_pldadapt_tx_23_tx_fifo_power_mode),
   .hssi_pldadapt_tx_23_tx_fifo_read_latency_adjust                                                                                     ( hssi_pldadapt_tx_23_tx_fifo_read_latency_adjust),
   .hssi_pldadapt_tx_23_tx_fifo_write_latency_adjust                                                                                    ( hssi_pldadapt_tx_23_tx_fifo_write_latency_adjust),
   .hssi_pldadapt_tx_23_tx_hip_aib_ssr_in_polling_bypass                                                                                ( hssi_pldadapt_tx_23_tx_hip_aib_ssr_in_polling_bypass),
   .hssi_pldadapt_tx_23_tx_osc_clock_setting                                                                                            ( hssi_pldadapt_tx_23_tx_osc_clock_setting),
   .hssi_pldadapt_tx_23_tx_pld_10g_tx_bitslip_polling_bypass                                                                            ( hssi_pldadapt_tx_23_tx_pld_10g_tx_bitslip_polling_bypass),
   .hssi_pldadapt_tx_23_tx_pld_8g_tx_boundary_sel_polling_bypass                                                                        ( hssi_pldadapt_tx_23_tx_pld_8g_tx_boundary_sel_polling_bypass),
   .hssi_pldadapt_tx_23_tx_pld_pma_fpll_cnt_sel_polling_bypass                                                                          ( hssi_pldadapt_tx_23_tx_pld_pma_fpll_cnt_sel_polling_bypass),
   .hssi_pldadapt_tx_23_tx_pld_pma_fpll_num_phase_shifts_polling_bypass                                                                 ( hssi_pldadapt_tx_23_tx_pld_pma_fpll_num_phase_shifts_polling_bypass),
   .hssi_pldadapt_tx_23_tx_usertest_sel                                                                                                 ( hssi_pldadapt_tx_23_tx_usertest_sel),
   .hssi_pldadapt_tx_23_txfifo_empty                                                                                                    ( hssi_pldadapt_tx_23_txfifo_empty),
   .hssi_pldadapt_tx_23_txfifo_full                                                                                                     ( hssi_pldadapt_tx_23_txfifo_full),
   .hssi_pldadapt_tx_23_txfifo_mode                                                                                                     ( hssi_pldadapt_tx_23_txfifo_mode),
   .hssi_pldadapt_tx_23_txfifo_pempty                                                                                                   ( hssi_pldadapt_tx_23_txfifo_pempty),
   .hssi_pldadapt_tx_23_txfifo_pfull                                                                                                    ( hssi_pldadapt_tx_23_txfifo_pfull),
   .hssi_pldadapt_tx_23_us_bypass_pipeln                                                                                                ( hssi_pldadapt_tx_23_us_bypass_pipeln),
   .hssi_pldadapt_tx_23_us_last_chnl                                                                                                    ( hssi_pldadapt_tx_23_us_last_chnl),
   .hssi_pldadapt_tx_23_us_master                                                                                                       ( hssi_pldadapt_tx_23_us_master),
   .hssi_pldadapt_tx_23_word_align_enable                                                                                               ( hssi_pldadapt_tx_23_word_align_enable),
   .hssi_pldadapt_tx_23_word_mark                                                                                                       ( hssi_pldadapt_tx_23_word_mark),
   .hssi_pldadapt_tx_23_silicon_rev                                                                                                     ( hssi_pldadapt_tx_23_silicon_rev),
   .hssi_pldadapt_tx_23_reconfig_settings                                                                                               ( hssi_pldadapt_tx_23_reconfig_settings),
   .hssi_pldadapt_rx_23_aib_clk1_sel                                                                                                    ( hssi_pldadapt_rx_23_aib_clk1_sel),
   .hssi_pldadapt_rx_23_aib_clk2_sel                                                                                                    ( hssi_pldadapt_rx_23_aib_clk2_sel),
   .hssi_pldadapt_rx_23_hdpldadapt_aib_fabric_pld_pma_hclk_hz                                                                           ( hssi_pldadapt_rx_23_hdpldadapt_aib_fabric_pld_pma_hclk_hz),
   .hssi_pldadapt_rx_23_hdpldadapt_aib_fabric_rx_sr_clk_in_hz                                                                           ( hssi_pldadapt_rx_23_hdpldadapt_aib_fabric_rx_sr_clk_in_hz),
   .hssi_pldadapt_rx_23_hdpldadapt_aib_fabric_rx_transfer_clk_hz                                                                        ( hssi_pldadapt_rx_23_hdpldadapt_aib_fabric_rx_transfer_clk_hz),
   .hssi_pldadapt_rx_23_asn_bypass_pma_pcie_sw_done                                                                                     ( hssi_pldadapt_rx_23_asn_bypass_pma_pcie_sw_done),
   .hssi_pldadapt_rx_23_asn_en                                                                                                          ( hssi_pldadapt_rx_23_asn_en),
   .hssi_pldadapt_rx_23_asn_wait_for_dll_reset_cnt                                                                                      ( hssi_pldadapt_rx_23_asn_wait_for_dll_reset_cnt),
   .hssi_pldadapt_rx_23_asn_wait_for_fifo_flush_cnt                                                                                     ( hssi_pldadapt_rx_23_asn_wait_for_fifo_flush_cnt),
   .hssi_pldadapt_rx_23_asn_wait_for_pma_pcie_sw_done_cnt                                                                               ( hssi_pldadapt_rx_23_asn_wait_for_pma_pcie_sw_done_cnt),
   .hssi_pldadapt_rx_23_bonding_dft_en                                                                                                  ( hssi_pldadapt_rx_23_bonding_dft_en),
   .hssi_pldadapt_rx_23_bonding_dft_val                                                                                                 ( hssi_pldadapt_rx_23_bonding_dft_val),
   .hssi_pldadapt_rx_23_chnl_bonding                                                                                                    ( hssi_pldadapt_rx_23_chnl_bonding),
   .hssi_pldadapt_rx_23_clock_del_measure_enable                                                                                        ( hssi_pldadapt_rx_23_clock_del_measure_enable),
   .hssi_pldadapt_rx_23_comp_cnt                                                                                                        ( hssi_pldadapt_rx_23_comp_cnt),
   .hssi_pldadapt_rx_23_compin_sel                                                                                                      ( hssi_pldadapt_rx_23_compin_sel),
   .hssi_pldadapt_rx_23_hdpldadapt_csr_clk_hz                                                                                           ( hssi_pldadapt_rx_23_hdpldadapt_csr_clk_hz),
   .hssi_pldadapt_rx_23_ctrl_plane_bonding                                                                                              ( hssi_pldadapt_rx_23_ctrl_plane_bonding),
   .hssi_pldadapt_rx_23_ds_bypass_pipeln                                                                                                ( hssi_pldadapt_rx_23_ds_bypass_pipeln),
   .hssi_pldadapt_rx_23_ds_last_chnl                                                                                                    ( hssi_pldadapt_rx_23_ds_last_chnl),
   .hssi_pldadapt_rx_23_ds_master                                                                                                       ( hssi_pldadapt_rx_23_ds_master),
   .hssi_pldadapt_rx_23_duplex_mode                                                                                                     ( hssi_pldadapt_rx_23_duplex_mode),
   .hssi_pldadapt_rx_23_dv_mode                                                                                                         ( hssi_pldadapt_rx_23_dv_mode),
   .hssi_pldadapt_rx_23_fifo_double_read                                                                                                ( hssi_pldadapt_rx_23_fifo_double_read),
   .hssi_pldadapt_rx_23_fifo_mode                                                                                                       ( hssi_pldadapt_rx_23_fifo_mode),
   .hssi_pldadapt_rx_23_fifo_rd_clk_ins_sm_scg_en                                                                                       ( hssi_pldadapt_rx_23_fifo_rd_clk_ins_sm_scg_en),
   .hssi_pldadapt_rx_23_fifo_rd_clk_scg_en                                                                                              ( hssi_pldadapt_rx_23_fifo_rd_clk_scg_en),
   .hssi_pldadapt_rx_23_fifo_rd_clk_sel                                                                                                 ( hssi_pldadapt_rx_23_fifo_rd_clk_sel),
   .hssi_pldadapt_rx_23_fifo_stop_rd                                                                                                    ( hssi_pldadapt_rx_23_fifo_stop_rd),
   .hssi_pldadapt_rx_23_fifo_stop_wr                                                                                                    ( hssi_pldadapt_rx_23_fifo_stop_wr),
   .hssi_pldadapt_rx_23_fifo_width                                                                                                      ( hssi_pldadapt_rx_23_fifo_width),
   .hssi_pldadapt_rx_23_fifo_wr_clk_del_sm_scg_en                                                                                       ( hssi_pldadapt_rx_23_fifo_wr_clk_del_sm_scg_en),
   .hssi_pldadapt_rx_23_fifo_wr_clk_scg_en                                                                                              ( hssi_pldadapt_rx_23_fifo_wr_clk_scg_en),
   .hssi_pldadapt_rx_23_fifo_wr_clk_sel                                                                                                 ( hssi_pldadapt_rx_23_fifo_wr_clk_sel),
   .hssi_pldadapt_rx_23_free_run_div_clk                                                                                                ( hssi_pldadapt_rx_23_free_run_div_clk),
   .hssi_pldadapt_rx_23_fsr_pld_10g_rx_crc32_err_rst_val                                                                                ( hssi_pldadapt_rx_23_fsr_pld_10g_rx_crc32_err_rst_val),
   .hssi_pldadapt_rx_23_fsr_pld_8g_sigdet_out_rst_val                                                                                   ( hssi_pldadapt_rx_23_fsr_pld_8g_sigdet_out_rst_val),
   .hssi_pldadapt_rx_23_fsr_pld_ltd_b_rst_val                                                                                           ( hssi_pldadapt_rx_23_fsr_pld_ltd_b_rst_val),
   .hssi_pldadapt_rx_23_fsr_pld_ltr_rst_val                                                                                             ( hssi_pldadapt_rx_23_fsr_pld_ltr_rst_val),
   .hssi_pldadapt_rx_23_fsr_pld_rx_fifo_align_clr_rst_val                                                                               ( hssi_pldadapt_rx_23_fsr_pld_rx_fifo_align_clr_rst_val),
   .hssi_pldadapt_rx_23_gb_rx_idwidth                                                                                                   ( hssi_pldadapt_rx_23_gb_rx_idwidth),
   .hssi_pldadapt_rx_23_gb_rx_odwidth                                                                                                   ( hssi_pldadapt_rx_23_gb_rx_odwidth),
   .hssi_pldadapt_rx_23_hip_mode                                                                                                        ( hssi_pldadapt_rx_23_hip_mode),
   .hssi_pldadapt_rx_23_hrdrst_align_bypass                                                                                             ( hssi_pldadapt_rx_23_hrdrst_align_bypass),
   .hssi_pldadapt_rx_23_hrdrst_dll_lock_bypass                                                                                          ( hssi_pldadapt_rx_23_hrdrst_dll_lock_bypass),
   .hssi_pldadapt_rx_23_hrdrst_rst_sm_dis                                                                                               ( hssi_pldadapt_rx_23_hrdrst_rst_sm_dis),
   .hssi_pldadapt_rx_23_hrdrst_rx_osc_clk_scg_en                                                                                        ( hssi_pldadapt_rx_23_hrdrst_rx_osc_clk_scg_en),
   .hssi_pldadapt_rx_23_hrdrst_user_ctl_en                                                                                              ( hssi_pldadapt_rx_23_hrdrst_user_ctl_en),
   .hssi_pldadapt_rx_23_indv                                                                                                            ( hssi_pldadapt_rx_23_indv),
   .hssi_pldadapt_rx_23_internal_clk1_sel1                                                                                              ( hssi_pldadapt_rx_23_internal_clk1_sel1),
   .hssi_pldadapt_rx_23_internal_clk1_sel2                                                                                              ( hssi_pldadapt_rx_23_internal_clk1_sel2),
   .hssi_pldadapt_rx_23_internal_clk2_sel1                                                                                              ( hssi_pldadapt_rx_23_internal_clk2_sel1),
   .hssi_pldadapt_rx_23_internal_clk2_sel2                                                                                              ( hssi_pldadapt_rx_23_internal_clk2_sel2),
   .hssi_pldadapt_rx_23_is_paired_with                                                                                                  ( hssi_pldadapt_rx_23_is_paired_with),
   .hssi_pldadapt_rx_23_loopback_mode                                                                                                   ( hssi_pldadapt_rx_23_loopback_mode),
   .hssi_pldadapt_rx_23_low_latency_en                                                                                                  ( hssi_pldadapt_rx_23_low_latency_en),
   .hssi_pldadapt_rx_23_lpbk_mode                                                                                                       ( hssi_pldadapt_rx_23_lpbk_mode),
   .hssi_pldadapt_rx_23_osc_clk_scg_en                                                                                                  ( hssi_pldadapt_rx_23_osc_clk_scg_en),
   .hssi_pldadapt_rx_23_phcomp_rd_del                                                                                                   ( hssi_pldadapt_rx_23_phcomp_rd_del),
   .hssi_pldadapt_rx_23_pipe_enable                                                                                                     ( hssi_pldadapt_rx_23_pipe_enable),
   .hssi_pldadapt_rx_23_pipe_mode                                                                                                       ( hssi_pldadapt_rx_23_pipe_mode),
   .hssi_pldadapt_rx_23_hdpldadapt_pld_avmm1_clk_rowclk_hz                                                                              ( hssi_pldadapt_rx_23_hdpldadapt_pld_avmm1_clk_rowclk_hz),
   .hssi_pldadapt_rx_23_hdpldadapt_pld_avmm2_clk_rowclk_hz                                                                              ( hssi_pldadapt_rx_23_hdpldadapt_pld_avmm2_clk_rowclk_hz),
   .hssi_pldadapt_rx_23_pld_clk1_delay_en                                                                                               ( hssi_pldadapt_rx_23_pld_clk1_delay_en),
   .hssi_pldadapt_rx_23_pld_clk1_delay_sel                                                                                              ( hssi_pldadapt_rx_23_pld_clk1_delay_sel),
   .hssi_pldadapt_rx_23_pld_clk1_inv_en                                                                                                 ( hssi_pldadapt_rx_23_pld_clk1_inv_en),
   .hssi_pldadapt_rx_23_pld_clk1_sel                                                                                                    ( hssi_pldadapt_rx_23_pld_clk1_sel),
   .hssi_pldadapt_rx_23_hdpldadapt_pld_rx_clk1_dcm_hz                                                                                   ( hssi_pldadapt_rx_23_hdpldadapt_pld_rx_clk1_dcm_hz),
   .hssi_pldadapt_rx_23_hdpldadapt_pld_rx_clk1_rowclk_hz                                                                                ( hssi_pldadapt_rx_23_hdpldadapt_pld_rx_clk1_rowclk_hz),
   .hssi_pldadapt_rx_23_hdpldadapt_pld_sclk1_rowclk_hz                                                                                  ( hssi_pldadapt_rx_23_hdpldadapt_pld_sclk1_rowclk_hz),
   .hssi_pldadapt_rx_23_hdpldadapt_pld_sclk2_rowclk_hz                                                                                  ( hssi_pldadapt_rx_23_hdpldadapt_pld_sclk2_rowclk_hz),
   .hssi_pldadapt_rx_23_pma_hclk_scg_en                                                                                                 ( hssi_pldadapt_rx_23_pma_hclk_scg_en),
   .hssi_pldadapt_rx_23_powerdown_mode                                                                                                  ( hssi_pldadapt_rx_23_powerdown_mode),
   .hssi_pldadapt_rx_23_powermode_dc                                                                                                    ( hssi_pldadapt_rx_23_powermode_dc),
   .hssi_pldadapt_rx_23_powermode_freq_hz_aib_fabric_rx_sr_clk_in                                                                       ( hssi_pldadapt_rx_23_powermode_freq_hz_aib_fabric_rx_sr_clk_in),
   .hssi_pldadapt_rx_23_powermode_freq_hz_pld_rx_clk1_dcm                                                                               ( hssi_pldadapt_rx_23_powermode_freq_hz_pld_rx_clk1_dcm),
   .hssi_pldadapt_rx_23_rx_datapath_tb_sel                                                                                              ( hssi_pldadapt_rx_23_rx_datapath_tb_sel),
   .hssi_pldadapt_rx_23_rx_fastbond_rden                                                                                                ( hssi_pldadapt_rx_23_rx_fastbond_rden),
   .hssi_pldadapt_rx_23_rx_fastbond_wren                                                                                                ( hssi_pldadapt_rx_23_rx_fastbond_wren),
   .hssi_pldadapt_rx_23_rx_fifo_power_mode                                                                                              ( hssi_pldadapt_rx_23_rx_fifo_power_mode),
   .hssi_pldadapt_rx_23_rx_fifo_read_latency_adjust                                                                                     ( hssi_pldadapt_rx_23_rx_fifo_read_latency_adjust),
   .hssi_pldadapt_rx_23_rx_fifo_write_ctrl                                                                                              ( hssi_pldadapt_rx_23_rx_fifo_write_ctrl),
   .hssi_pldadapt_rx_23_rx_fifo_write_latency_adjust                                                                                    ( hssi_pldadapt_rx_23_rx_fifo_write_latency_adjust),
   .hssi_pldadapt_rx_23_rx_osc_clock_setting                                                                                            ( hssi_pldadapt_rx_23_rx_osc_clock_setting),
   .hssi_pldadapt_rx_23_rx_pld_8g_eidleinfersel_polling_bypass                                                                          ( hssi_pldadapt_rx_23_rx_pld_8g_eidleinfersel_polling_bypass),
   .hssi_pldadapt_rx_23_rx_pld_pma_eye_monitor_polling_bypass                                                                           ( hssi_pldadapt_rx_23_rx_pld_pma_eye_monitor_polling_bypass),
   .hssi_pldadapt_rx_23_rx_pld_pma_pcie_switch_polling_bypass                                                                           ( hssi_pldadapt_rx_23_rx_pld_pma_pcie_switch_polling_bypass),
   .hssi_pldadapt_rx_23_rx_pld_pma_reser_out_polling_bypass                                                                             ( hssi_pldadapt_rx_23_rx_pld_pma_reser_out_polling_bypass),
   .hssi_pldadapt_rx_23_rx_prbs_flags_sr_enable                                                                                         ( hssi_pldadapt_rx_23_rx_prbs_flags_sr_enable),
   .hssi_pldadapt_rx_23_rx_true_b2b                                                                                                     ( hssi_pldadapt_rx_23_rx_true_b2b),
   .hssi_pldadapt_rx_23_rx_usertest_sel                                                                                                 ( hssi_pldadapt_rx_23_rx_usertest_sel),
   .hssi_pldadapt_rx_23_rxfifo_empty                                                                                                    ( hssi_pldadapt_rx_23_rxfifo_empty),
   .hssi_pldadapt_rx_23_rxfifo_full                                                                                                     ( hssi_pldadapt_rx_23_rxfifo_full),
   .hssi_pldadapt_rx_23_rxfifo_mode                                                                                                     ( hssi_pldadapt_rx_23_rxfifo_mode),
   .hssi_pldadapt_rx_23_rxfifo_pempty                                                                                                   ( hssi_pldadapt_rx_23_rxfifo_pempty),
   .hssi_pldadapt_rx_23_rxfifo_pfull                                                                                                    ( hssi_pldadapt_rx_23_rxfifo_pfull),
   .hssi_pldadapt_rx_23_rxfiford_post_ct_sel                                                                                            ( hssi_pldadapt_rx_23_rxfiford_post_ct_sel),
   .hssi_pldadapt_rx_23_rxfifowr_post_ct_sel                                                                                            ( hssi_pldadapt_rx_23_rxfifowr_post_ct_sel),
   .hssi_pldadapt_rx_23_sclk_sel                                                                                                        ( hssi_pldadapt_rx_23_sclk_sel),
   .hssi_pldadapt_rx_23_hdpldadapt_speed_grade                                                                                          ( hssi_pldadapt_rx_23_hdpldadapt_speed_grade),
   .hssi_pldadapt_rx_23_hdpldadapt_sr_sr_testbus_sel                                                                                    ( hssi_pldadapt_rx_23_hdpldadapt_sr_sr_testbus_sel),
   .hssi_pldadapt_rx_23_stretch_num_stages                                                                                              ( hssi_pldadapt_rx_23_stretch_num_stages),
   .hssi_pldadapt_rx_23_sup_mode                                                                                                        ( hssi_pldadapt_rx_23_sup_mode),
   .hssi_pldadapt_rx_23_txfiford_post_ct_sel                                                                                            ( hssi_pldadapt_rx_23_txfiford_post_ct_sel),
   .hssi_pldadapt_rx_23_txfifowr_post_ct_sel                                                                                            ( hssi_pldadapt_rx_23_txfifowr_post_ct_sel),
   .hssi_pldadapt_rx_23_us_bypass_pipeln                                                                                                ( hssi_pldadapt_rx_23_us_bypass_pipeln),
   .hssi_pldadapt_rx_23_us_last_chnl                                                                                                    ( hssi_pldadapt_rx_23_us_last_chnl),
   .hssi_pldadapt_rx_23_us_master                                                                                                       ( hssi_pldadapt_rx_23_us_master),
   .hssi_pldadapt_rx_23_word_align                                                                                                      ( hssi_pldadapt_rx_23_word_align),
   .hssi_pldadapt_rx_23_word_align_enable                                                                                               ( hssi_pldadapt_rx_23_word_align_enable),
   .hssi_pldadapt_rx_23_silicon_rev                                                                                                     ( hssi_pldadapt_rx_23_silicon_rev),
   .hssi_pldadapt_rx_23_reconfig_settings                                                                                               ( hssi_pldadapt_rx_23_reconfig_settings),
   .hssi_avmm1_if_23_pcs_arbiter_ctrl                                                                                                   ( hssi_avmm1_if_23_pcs_arbiter_ctrl),
   .hssi_avmm1_if_23_hssiadapt_avmm_clk_dcg_en                                                                                          ( hssi_avmm1_if_23_hssiadapt_avmm_clk_dcg_en),
   .hssi_avmm1_if_23_hssiadapt_avmm_clk_scg_en                                                                                          ( hssi_avmm1_if_23_hssiadapt_avmm_clk_scg_en),
   .hssi_avmm1_if_23_pldadapt_avmm_clk_scg_en                                                                                           ( hssi_avmm1_if_23_pldadapt_avmm_clk_scg_en),
   .hssi_avmm1_if_23_pcs_cal_done                                                                                                       ( hssi_avmm1_if_23_pcs_cal_done),
   .hssi_avmm1_if_23_pcs_cal_reserved                                                                                                   ( hssi_avmm1_if_23_pcs_cal_reserved),
   .hssi_avmm1_if_23_pcs_calibration_feature_en                                                                                         ( hssi_avmm1_if_23_pcs_calibration_feature_en),
   .hssi_avmm1_if_23_pldadapt_gate_dis                                                                                                  ( hssi_avmm1_if_23_pldadapt_gate_dis),
   .hssi_avmm1_if_23_pcs_hip_cal_en                                                                                                     ( hssi_avmm1_if_23_pcs_hip_cal_en),
   .hssi_avmm1_if_23_hssiadapt_nfhssi_calibratio_feature_en                                                                             ( hssi_avmm1_if_23_hssiadapt_nfhssi_calibratio_feature_en),
   .hssi_avmm1_if_23_pldadapt_nfhssi_calibratio_feature_en                                                                              ( hssi_avmm1_if_23_pldadapt_nfhssi_calibratio_feature_en),
   .hssi_avmm1_if_23_hssiadapt_osc_clk_scg_en                                                                                           ( hssi_avmm1_if_23_hssiadapt_osc_clk_scg_en),
   .hssi_avmm1_if_23_pldadapt_osc_clk_scg_en                                                                                            ( hssi_avmm1_if_23_pldadapt_osc_clk_scg_en),
   .hssi_avmm1_if_23_hssiadapt_read_blocking_enable                                                                                     ( hssi_avmm1_if_23_hssiadapt_read_blocking_enable),
   .hssi_avmm1_if_23_pldadapt_read_blocking_enable                                                                                      ( hssi_avmm1_if_23_pldadapt_read_blocking_enable),
   .hssi_avmm1_if_23_hssiadapt_uc_blocking_enable                                                                                       ( hssi_avmm1_if_23_hssiadapt_uc_blocking_enable),
   .hssi_avmm1_if_23_pldadapt_uc_blocking_enable                                                                                        ( hssi_avmm1_if_23_pldadapt_uc_blocking_enable),
   .hssi_avmm1_if_23_hssiadapt_write_resp_en                                                                                            ( hssi_avmm1_if_23_hssiadapt_write_resp_en),
   .hssi_avmm1_if_23_hssiadapt_avmm_osc_clock_setting                                                                                   ( hssi_avmm1_if_23_hssiadapt_avmm_osc_clock_setting),
   .hssi_avmm1_if_23_pldadapt_avmm_osc_clock_setting                                                                                    ( hssi_avmm1_if_23_pldadapt_avmm_osc_clock_setting),
   .hssi_avmm1_if_23_hssiadapt_avmm_testbus_sel                                                                                         ( hssi_avmm1_if_23_hssiadapt_avmm_testbus_sel),
   .hssi_avmm1_if_23_pldadapt_avmm_testbus_sel                                                                                          ( hssi_avmm1_if_23_pldadapt_avmm_testbus_sel),
   .hssi_avmm1_if_23_func_mode                                                                                                          ( hssi_avmm1_if_23_func_mode),
   .hssi_avmm1_if_23_hssiadapt_sr_hip_mode                                                                                              ( hssi_avmm1_if_23_hssiadapt_sr_hip_mode),
   .hssi_avmm1_if_23_hssiadapt_hip_mode                                                                                                 ( hssi_avmm1_if_23_hssiadapt_hip_mode),
   .hssi_avmm1_if_23_pldadapt_hip_mode                                                                                                  ( hssi_avmm1_if_23_pldadapt_hip_mode),
   .hssi_avmm1_if_23_hssiadapt_sr_powerdown_mode                                                                                        ( hssi_avmm1_if_23_hssiadapt_sr_powerdown_mode),
   .hssi_avmm1_if_23_hssiadapt_sr_sr_free_run_div_clk                                                                                   ( hssi_avmm1_if_23_hssiadapt_sr_sr_free_run_div_clk),
   .hssi_avmm1_if_23_hssiadapt_sr_sr_hip_en                                                                                             ( hssi_avmm1_if_23_hssiadapt_sr_sr_hip_en),
   .hssi_avmm1_if_23_hssiadapt_sr_sr_osc_clk_div_sel                                                                                    ( hssi_avmm1_if_23_hssiadapt_sr_sr_osc_clk_div_sel),
   .hssi_avmm1_if_23_hssiadapt_sr_sr_osc_clk_scg_en                                                                                     ( hssi_avmm1_if_23_hssiadapt_sr_sr_osc_clk_scg_en),
   .hssi_avmm1_if_23_hssiadapt_sr_sr_parity_en                                                                                          ( hssi_avmm1_if_23_hssiadapt_sr_sr_parity_en),
   .hssi_avmm1_if_23_hssiadapt_sr_sr_reserved_in_en                                                                                     ( hssi_avmm1_if_23_hssiadapt_sr_sr_reserved_in_en),
   .hssi_avmm1_if_23_hssiadapt_sr_sr_reserved_out_en                                                                                    ( hssi_avmm1_if_23_hssiadapt_sr_sr_reserved_out_en),
   .hssi_avmm1_if_23_hssiadapt_sr_sup_mode                                                                                              ( hssi_avmm1_if_23_hssiadapt_sr_sup_mode),
   .hssi_avmm1_if_23_topology                                                                                                           ( hssi_avmm1_if_23_topology),
   .hssi_avmm1_if_23_silicon_rev                                                                                                        ( hssi_avmm1_if_23_silicon_rev),
   .hssi_avmm1_if_23_calibration_type                                                                                                   ( hssi_avmm1_if_23_calibration_type),
   .hssi_avmm2_if_23_pcs_arbiter_ctrl                                                                                                   ( hssi_avmm2_if_23_pcs_arbiter_ctrl),
   .hssi_avmm2_if_23_hssiadapt_avmm_clk_dcg_en                                                                                          ( hssi_avmm2_if_23_hssiadapt_avmm_clk_dcg_en),
   .hssi_avmm2_if_23_hssiadapt_avmm_clk_scg_en                                                                                          ( hssi_avmm2_if_23_hssiadapt_avmm_clk_scg_en),
   .hssi_avmm2_if_23_pldadapt_avmm_clk_scg_en                                                                                           ( hssi_avmm2_if_23_pldadapt_avmm_clk_scg_en),
   .hssi_avmm2_if_23_pcs_cal_done                                                                                                       ( hssi_avmm2_if_23_pcs_cal_done),
   .hssi_avmm2_if_23_pcs_cal_reserved                                                                                                   ( hssi_avmm2_if_23_pcs_cal_reserved),
   .hssi_avmm2_if_23_pcs_calibration_feature_en                                                                                         ( hssi_avmm2_if_23_pcs_calibration_feature_en),
   .hssi_avmm2_if_23_pldadapt_gate_dis                                                                                                  ( hssi_avmm2_if_23_pldadapt_gate_dis),
   .hssi_avmm2_if_23_pcs_hip_cal_en                                                                                                     ( hssi_avmm2_if_23_pcs_hip_cal_en),
   .hssi_avmm2_if_23_hssiadapt_osc_clk_scg_en                                                                                           ( hssi_avmm2_if_23_hssiadapt_osc_clk_scg_en),
   .hssi_avmm2_if_23_pldadapt_osc_clk_scg_en                                                                                            ( hssi_avmm2_if_23_pldadapt_osc_clk_scg_en),
   .hssi_avmm2_if_23_hssiadapt_avmm_osc_clock_setting                                                                                   ( hssi_avmm2_if_23_hssiadapt_avmm_osc_clock_setting),
   .hssi_avmm2_if_23_pldadapt_avmm_osc_clock_setting                                                                                    ( hssi_avmm2_if_23_pldadapt_avmm_osc_clock_setting),
   .hssi_avmm2_if_23_hssiadapt_avmm_testbus_sel                                                                                         ( hssi_avmm2_if_23_hssiadapt_avmm_testbus_sel),
   .hssi_avmm2_if_23_pldadapt_avmm_testbus_sel                                                                                          ( hssi_avmm2_if_23_pldadapt_avmm_testbus_sel),
   .hssi_avmm2_if_23_func_mode                                                                                                          ( hssi_avmm2_if_23_func_mode),
   .hssi_avmm2_if_23_hssiadapt_hip_mode                                                                                                 ( hssi_avmm2_if_23_hssiadapt_hip_mode),
   .hssi_avmm2_if_23_pldadapt_hip_mode                                                                                                  ( hssi_avmm2_if_23_pldadapt_hip_mode),
   .hssi_avmm2_if_23_topology                                                                                                           ( hssi_avmm2_if_23_topology),
   .hssi_avmm2_if_23_silicon_rev                                                                                                        ( hssi_avmm2_if_23_silicon_rev),
   .hssi_avmm2_if_23_calibration_type                                                                                                   ( hssi_avmm2_if_23_calibration_type),
   .hssi_ctr_active_lane_octet0                                                                                                         ( hssi_ctr_active_lane_octet0),
   .hssi_ctr_active_lane_octet1                                                                                                         ( hssi_ctr_active_lane_octet1),
   .hssi_ctr_htol                                                                                                                       ( hssi_ctr_htol),
   .hssi_ctr_independent_pcie_x8x8                                                                                                      ( hssi_ctr_independent_pcie_x8x8),
   .hssi_ctr_iopads_powerdown_mode                                                                                                      ( hssi_ctr_iopads_powerdown_mode),
   .hssi_ctr_is_cvp_enable                                                                                                              ( hssi_ctr_is_cvp_enable),
   .hssi_ctr_pcie_capable                                                                                                               ( hssi_ctr_pcie_capable),
   .hssi_ctr_pcie_p0_config                                                                                                             ( hssi_ctr_pcie_p0_config),
   .hssi_ctr_pcie_p1_config                                                                                                             ( hssi_ctr_pcie_p1_config),
   .hssi_ctr_pcie_p2_config                                                                                                             ( hssi_ctr_pcie_p2_config),
   .hssi_ctr_pcie_p3_config                                                                                                             ( hssi_ctr_pcie_p3_config),
   .hssi_ctr_pcie_pld_data_width                                                                                                        ( hssi_ctr_pcie_pld_data_width),
   .hssi_ctr_pcie_virt_aspm                                                                                                             ( hssi_ctr_pcie_virt_aspm),
   .hssi_ctr_pipe_direct_octet0                                                                                                         ( hssi_ctr_pipe_direct_octet0),
   .hssi_ctr_pipe_direct_octet1                                                                                                         ( hssi_ctr_pipe_direct_octet1),
   .hssi_ctr_pld_txrx_clk_hz                                                                                                            ( hssi_ctr_pld_txrx_clk_hz),
   .hssi_ctr_powerdown_mode                                                                                                             ( hssi_ctr_powerdown_mode),
   .hssi_ctr_sup_mode                                                                                                                   ( hssi_ctr_sup_mode),
   .hssi_ctr_topology                                                                                                                   ( hssi_ctr_topology),
   .hssi_ctr_u_aib_top_powerdown_mode                                                                                                   ( hssi_ctr_u_aib_top_powerdown_mode),
   .hssi_ctr_u_aib_top_sup_mode                                                                                                         ( hssi_ctr_u_aib_top_sup_mode),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp0                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp1                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp2                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp3                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_reset_n                                                                     ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp1                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp2                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp3                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger1_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_0_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_10_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_11_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_12_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_13_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_14_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_15_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_16_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_17_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_18_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_19_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp0                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp1                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp2                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp3                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_reset_n                                                                     ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp1                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp2                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp3                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger1_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_1_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_20_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_21_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_22_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                             ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                 ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp0                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp1                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp2                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp3                                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_reset_n                                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp1                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp2                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp3                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger1_sel_grp0                                                          ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_23_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp0                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp1                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp2                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp3                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_reset_n                                                                     ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp1                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp2                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp3                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger1_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_2_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp0                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp1                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp2                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp3                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_reset_n                                                                     ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp1                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp2                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp3                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger1_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_3_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp0                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp1                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp2                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp3                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_reset_n                                                                     ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp1                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp2                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp3                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger1_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_4_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp0                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp1                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp2                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp3                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_reset_n                                                                     ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp1                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp2                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp3                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger1_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_5_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp0                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp1                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp2                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp3                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_reset_n                                                                     ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp1                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp2                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp3                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger1_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_6_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp0                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp1                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp2                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp3                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_reset_n                                                                     ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp1                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp2                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp3                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger1_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_7_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp0                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp1                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp2                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp3                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_reset_n                                                                     ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp1                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp2                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp3                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger1_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_8_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_avmm_avmm_testbus_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_avmm_avmm_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_internal_clk1_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel                                                ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_internal_clk2_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_pcs_testbus_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel                                              ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_pma_div2_clk_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_ssr_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel                                                  ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_rx_usertest_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_rxchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel                                                   ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_sr_sr_osc_clk_div_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_hrdrst_user_ctl_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_phcomp_rd_del                                                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_phcomp_rd_del),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_stretch_num_stages                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_stretch_num_stages),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_adapter_txchnl_tx_datapath_tb_sel),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp0                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp1                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp2                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp3                                                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_data_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_reset_n                                                                     ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp1                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp1),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp2                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp2),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp3                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger0_sel_grp3),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger1_sel_grp0                                                           ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibadapter_dfd_trigger1_sel_grp0),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibchl_top_wrp_xrnr_aibchl_top_xrxdatapath_rx_dft_hssitestip_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en                               ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dfd_dll_dcc_en),
   .hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en                    ( hssi_ctr_u_aib_top_u_aibadapt_wrap_9_rnr_aibchl_top_wrp_xrnr_aibchl_top_xtxdatapath_tx_dft_hssitestip_dll_dcc_en),
   
   .hssi_ctr_true_independent_support_mode ( hssi_ctr_true_independent_support_mode),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_disable_phy_timer ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_disable_phy_timer),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_enable_phy_status ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_enable_phy_status),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_octet_cfg_en ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_octet_cfg_en),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pin_perst0_is_fullrst ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pin_perst0_is_fullrst),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pin_perst1_is_fullrst ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pin_perst1_is_fullrst),
   
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_async_direct_rx_sel                                                                  ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_async_direct_rx_sel),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_byp_mode                                                                             ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_byp_mode),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_ctrl_0_control                                                                ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_ctrl_0_control)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_ctrl_1_control                                                                ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_ctrl_1_control)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_ctrl_2_control                                                                ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_ctrl_2_control)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_irq_msk                                                                       ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_bypass_irq_msk)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_pldpll_disable                                                                   ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_pldpll_disable),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_second_pipepll_en                                                                ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_second_pipepll_en),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_sel_reset_assert                                                                 ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_sel_reset_assert),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_sel_reset_deassert                                                               ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cfg_sel_reset_deassert),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cold_reset_time                                                                      ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cold_reset_time),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_core_rst_width                                                                       ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_core_rst_width),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cpll_post_rls_quiet_time                                                             ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cpll_post_rls_quiet_time),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cpll_post_rst_quiet_time                                                             ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_cpll_post_rst_quiet_time),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_adpt_0to7                                                                    ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_adpt_0to7)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_adpt_16to23                                                                  ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_adpt_16to23)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_adpt_8to15                                                                   ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_adpt_8to15)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_hrc                                                                          ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_mux_hrc),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_pattern_cntr_data_sel                                                            ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_pattern_cntr_data_sel),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_reset_n                                                                          ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dfd_reset_n),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dis_chkplllock_b4_corerst                                                            ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dis_chkplllock_b4_corerst),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dis_phystatchk_b4_partialrst                                                         ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_dis_phystatchk_b4_partialrst),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_error_irq_msk                                                                        ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_error_irq_msk)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp0_sel                                                                     ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp0_sel)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp1_sel                                                                     ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp1_sel)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp2_sel                                                                     ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp2_sel)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp3_sel                                                                     ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_hrc_dfd_grp3_sel)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_lane_rls_quiet_time                                                                  ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_lane_rls_quiet_time),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_lane_stagger_disable                                                                 ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_lane_stagger_disable),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_lane_stagger_interval                                                                ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_lane_stagger_interval),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_linkreq_fullrst                                                                      ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_linkreq_fullrst),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_linkreq_partialrst                                                                   ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_linkreq_partialrst),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_perst_hi_filt_time                                                                   ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_perst_hi_filt_time),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_perst_lo_filt_time                                                                   ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_perst_lo_filt_time),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_phy_lane_rst_width                                                                   ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_phy_lane_rst_width),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_phy_post_lane_rst_quiet_time                                                         ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_phy_post_lane_rst_quiet_time),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pin_perst_is_full_rst                                                                ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pin_perst_is_full_rst),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pipepll_error_timeout                                                                ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pipepll_error_timeout)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pldpll_error_timeout                                                                 ( str_2_bin(hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pldpll_error_timeout)),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pldpll_rsten_warm                                                                    ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_pldpll_rsten_warm),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_post_core_rst_quiet_time                                                             ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_post_core_rst_quiet_time),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_sideband_clksel                                                                      ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_sideband_clksel),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_warm_rst_timeout                                                                     ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_warm_rst_timeout),
   .hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_warm_rst_timeout_prescaler                                                           ( hssi_ctr_u_aib_top_u_rnr_aib_cmn_u_rnr_hrc_top_warm_rst_timeout_prescaler),
   .hssi_ctr_u_ctrl_powerdown_mode                                                                                                      ( hssi_ctr_u_ctrl_powerdown_mode),
   
   .hssi_ctr_u_ctrl_toolkit_debug_mode ( hssi_ctr_u_ctrl_toolkit_debug_mode),
   
   .hssi_ctr_u_ial_top_cxl_op_mode                                                                                                      ( hssi_ctr_u_ial_top_cxl_op_mode),
   .hssi_ctr_u_ial_top_r_credit_return_scheme                                                                                           ( hssi_ctr_u_ial_top_r_credit_return_scheme),
   .hssi_ctr_u_ial_top_r_cxlio_dphy_send_lidl_en_dis                                                                                    ( hssi_ctr_u_ial_top_r_cxlio_dphy_send_lidl_en_dis),
   .hssi_ctr_u_ial_top_r_flp_phy_rcvd_ts2_all_lanes_dis                                                                                 ( hssi_ctr_u_ial_top_r_flp_phy_rcvd_ts2_all_lanes_dis),
   .hssi_ctr_u_ial_top_r_s2m_drs_bypass_disrepflithdr                                                                                   ( hssi_ctr_u_ial_top_r_s2m_drs_bypass_disrepflithdr),
   .hssi_ctr_u_ial_top_r_wptr_delay                                                                                                     ( hssi_ctr_u_ial_top_r_wptr_delay),
   .hssi_ctr_u_ial_top_rnr_ialup_flp_inst_flxbusptctl_driftbuf_en                                                                       ( hssi_ctr_u_ial_top_rnr_ialup_flp_inst_flxbusptctl_driftbuf_en),
   .hssi_ctr_u_ial_top_rnr_ialup_flp_inst_hybrid_x4_width                                                                               ( hssi_ctr_u_ial_top_rnr_ialup_flp_inst_hybrid_x4_width),
   .hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl2_ialinvratelnkdn                                                                       ( hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl2_ialinvratelnkdn),
   .hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl2_vid                                                                                   ( hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl2_vid),
   .hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl_comclk                                                                                 ( hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl_comclk),
   .hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl_force_ial                                                                              ( hssi_ctr_u_ial_top_rnr_ialup_flp_inst_iapctl_force_ial),
   .hssi_ctr_u_ial_top_rnr_ialup_flp_inst_sosctl_srisen                                                                                 ( hssi_ctr_u_ial_top_rnr_ialup_flp_inst_sosctl_srisen),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_cxl_ldid_en                                                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_cxl_ldid_en),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_ialpmmctl_vid                                                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_ialpmmctl_vid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_ialpmmctl_vmeb15                                                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_ialpmmctl_vmeb15),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rcrbbar_en                                                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rcrbbar_en),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cfg_avmm_csr_k_partial_bypass_configload                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cfg_avmm_csr_k_partial_bypass_configload),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_chemem_ctrl_k_perframe_addr_steer_opt                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_chemem_ctrl_k_perframe_addr_steer_opt),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_chemem_ctrl_k_perframe_cqid_steer_opt                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_chemem_ctrl_k_perframe_cqid_steer_opt),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_chemem_ctrl_k_perframe_slice_en                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_chemem_ctrl_k_perframe_slice_en),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_clk_csr_k_clkreq_hysterisis                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_clk_csr_k_clkreq_hysterisis),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_clk_csr_k_clock_control                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_clk_csr_k_clock_control),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_clk_csr_k_osc_clk_dis                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_clk_csr_k_osc_clk_dis),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_2_k_compressed                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_2_k_compressed),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_2_k_devbrd_type                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_2_k_devbrd_type),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_2_k_encryped                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_2_k_encryped),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_3_k_jtag_id_3                                                        ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_3_k_jtag_id_3)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_4_k_jtag_id_2                                                        ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_4_k_jtag_id_2)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_5_k_jtag_id_1                                                        ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_5_k_jtag_id_1)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_6_k_jtag_id_0                                                        ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_6_k_jtag_id_0)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_7_k_cvp_irq_en                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_7_k_cvp_irq_en),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_7_k_cvp_write_mask_ctl                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_7_k_cvp_write_mask_ctl),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_7_k_gpio_irq                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_cvp_ctrl_7_k_gpio_irq),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_h2d_arb_ctrl_k_h2drsp_throttle_en                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_h2d_arb_ctrl_k_h2drsp_throttle_en),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_ica_ctrl_k_ica_dbg_stepthrumode                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_ica_ctrl_k_ica_dbg_stepthrumode),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_opcode_lock_k_opcode_lock                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_opcode_lock_k_opcode_lock),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_aer_cntrl_reg_aer_ecrc_chk_capable                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_aer_cntrl_reg_aer_ecrc_chk_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_aer_cntrl_reg_aer_ecrc_gen_capable                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_aer_cntrl_reg_aer_ecrc_gen_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_global_inval_suppport                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_global_inval_suppport),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_inval_queue_dep                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_inval_queue_dep),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_page_aglign_req                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_page_aglign_req),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_ro_support                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ats_reg_ro_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg2_cpl_to_dis_support                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg2_cpl_to_dis_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg2_ee_tlp_prefix_support                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg2_ee_tlp_prefix_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg2_tph_cpl_support                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg2_tph_cpl_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_ep_l0_acc_lat                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_ep_l0_acc_lat),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_ep_l1_acc_lat                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_ep_l1_acc_lat),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_flr_cap                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_flr_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_rb_err_rptr                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devcapreg_rb_err_rptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devvendid_deviceid                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devvendid_deviceid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devvendid_vendorid                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_devvendid_vendorid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_high_memory_range1_size_high                   ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_high_memory_range1_size_high)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_desired_interleave_range1                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_desired_interleave_range1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_media_type_range1                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_media_type_range1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_active_range1                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_active_range1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_class_range1                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_class_range1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_info_valid_range1                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_info_valid_range1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_range1_size_low                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range1_size_low_memory_range1_size_low),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_high_memory_range2_size_high                   ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_high_memory_range2_size_high)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_desired_interleave_range2                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_desired_interleave_range2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_media_type_range2                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_media_type_range2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_active_range2                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_active_range2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_class_range2                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_class_range2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_info_valid_range2                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_info_valid_range2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_range2_size_low                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_flex_bus_range2_size_low_memory_range2_size_low),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_dvsecid                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_dvsecid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_hdm_count                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_hdm_count),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_mem_hwinit_mode                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_mem_hwinit_mode),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_viral_capable                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_dvsec_head2_cap_viral_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msi_cap_reg_extnd_msg_data_capable                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msi_cap_reg_extnd_msg_data_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msi_cap_reg_mul_msg_cap                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msi_cap_reg_mul_msg_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msi_cap_reg_per_vector_msk_cap                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msi_cap_reg_per_vector_msk_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_cap_reg_table_sz                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_cap_reg_table_sz),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_pba_ptr_pba_bir                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_pba_ptr_pba_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_pba_ptr_pba_offset                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_pba_ptr_pba_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_table_ptr_table_bir                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_table_ptr_table_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_table_ptr_table_offset                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_msix_table_ptr_table_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_pasid_reg_exec_permi_supp                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_pasid_reg_exec_permi_supp),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_pasid_reg_pasid_max_width                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_pasid_reg_pasid_max_width),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_pasid_reg_privil_mode_supp                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_pasid_reg_privil_mode_supp),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ptm_cap_reg_local_clock_granularity                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ptm_cap_reg_local_clock_granularity),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ptm_cap_reg_ptm_rqstr_capable                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_ptm_cap_reg_ptm_rqstr_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_reset_entry_bypass_reset_entry_bypass_idle_check                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_reset_entry_bypass_reset_entry_bypass_idle_check),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_revclasscode_class_codes                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_revclasscode_class_codes),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_revclasscode_rid                                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_revclasscode_rid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_siov_dvsec_flags_h                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_siov_dvsec_flags_h),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_siov_dvsec_funtion_dependency_link                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_siov_dvsec_funtion_dependency_link),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_siov_reg3_ims_support                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_siov_reg3_ims_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_sriov_cap_vf_mig_cap                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_sriov_cap_vf_mig_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_sriov_cap_vf_mig_int                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_sriov_cap_vf_mig_int),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_subsystemid_subsystemid                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_subsystemid_subsystemid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_subsystemid_subsystemvendorid                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_subsystemid_subsystemvendorid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_dev_spec_mode_supd                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_dev_spec_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_etph_req_supd                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_etph_req_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_int_vct_mode_supd                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_int_vct_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_st_table_loc                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_st_table_loc),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_tph_st_tab_size                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_tph_req_cap_reg_tph_st_tab_size),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_0_vf_ats_globalinv_support_0                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_0_vf_ats_globalinv_support_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_0_vf_ats_invqueue_depth_0                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_0_vf_ats_invqueue_depth_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_0_vf_ats_pagealignedreq_0                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_0_vf_ats_pagealignedreq_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_1_vf_ats_globalinv_support_1                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_1_vf_ats_globalinv_support_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_1_vf_ats_invqueue_depth_1                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_1_vf_ats_invqueue_depth_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_1_vf_ats_pagealignedreq_1                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_1_vf_ats_pagealignedreq_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_2_vf_ats_globalinv_support_2                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_2_vf_ats_globalinv_support_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_2_vf_ats_invqueue_depth_2                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_2_vf_ats_invqueue_depth_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_2_vf_ats_pagealignedreq_2                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_2_vf_ats_pagealignedreq_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_3_vf_ats_globalinv_support_3                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_3_vf_ats_globalinv_support_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_3_vf_ats_invqueue_depth_3                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_3_vf_ats_invqueue_depth_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_3_vf_ats_pagealignedreq_3                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_3_vf_ats_pagealignedreq_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_4_vf_ats_globalinv_support_4                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_4_vf_ats_globalinv_support_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_4_vf_ats_invqueue_depth_4                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_4_vf_ats_invqueue_depth_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_4_vf_ats_pagealignedreq_4                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_4_vf_ats_pagealignedreq_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_5_vf_ats_globalinv_support_5                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_5_vf_ats_globalinv_support_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_5_vf_ats_invqueue_depth_5                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_5_vf_ats_invqueue_depth_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_5_vf_ats_pagealignedreq_5                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_5_vf_ats_pagealignedreq_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_6_vf_ats_globalinv_support_6                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_6_vf_ats_globalinv_support_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_6_vf_ats_invqueue_depth_6                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_6_vf_ats_invqueue_depth_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_6_vf_ats_pagealignedreq_6                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_6_vf_ats_pagealignedreq_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_7_vf_ats_globalinv_support_7                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_7_vf_ats_globalinv_support_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_7_vf_ats_invqueue_depth_7                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_7_vf_ats_invqueue_depth_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_7_vf_ats_pagealignedreq_7                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_atscap_7_vf_ats_pagealignedreq_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_device_id_vf_device_id                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_device_id_vf_device_id),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_0_vf_msix_pba_bir_0                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_0_vf_msix_pba_bir_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_0_vf_msix_pba_offset_0                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_0_vf_msix_pba_offset_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_1_vf_msix_pba_bir_1                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_1_vf_msix_pba_bir_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_1_vf_msix_pba_offset_1                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_1_vf_msix_pba_offset_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_2_vf_msix_pba_bir_2                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_2_vf_msix_pba_bir_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_2_vf_msix_pba_offset_2                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_2_vf_msix_pba_offset_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_3_vf_msix_pba_bir_3                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_3_vf_msix_pba_bir_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_3_vf_msix_pba_offset_3                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_3_vf_msix_pba_offset_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_4_vf_msix_pba_bir_4                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_4_vf_msix_pba_bir_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_4_vf_msix_pba_offset_4                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_4_vf_msix_pba_offset_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_5_vf_msix_pba_bir_5                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_5_vf_msix_pba_bir_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_5_vf_msix_pba_offset_5                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_5_vf_msix_pba_offset_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_6_vf_msix_pba_bir_6                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_6_vf_msix_pba_bir_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_6_vf_msix_pba_offset_6                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_6_vf_msix_pba_offset_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_7_vf_msix_pba_bir_7                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_7_vf_msix_pba_bir_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_7_vf_msix_pba_offset_7                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_pba_7_vf_msix_pba_offset_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_0_vf_msix_table_bir_0                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_0_vf_msix_table_bir_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_0_vf_msix_table_offset_0                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_0_vf_msix_table_offset_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_1_vf_msix_table_bir_1                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_1_vf_msix_table_bir_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_1_vf_msix_table_offset_1                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_1_vf_msix_table_offset_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_2_vf_msix_table_bir_2                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_2_vf_msix_table_bir_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_2_vf_msix_table_offset_2                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_2_vf_msix_table_offset_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_3_vf_msix_table_bir_3                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_3_vf_msix_table_bir_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_3_vf_msix_table_offset_3                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_3_vf_msix_table_offset_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_4_vf_msix_table_bir_4                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_4_vf_msix_table_bir_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_4_vf_msix_table_offset_4                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_4_vf_msix_table_offset_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_5_vf_msix_table_bir_5                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_5_vf_msix_table_bir_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_5_vf_msix_table_offset_5                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_5_vf_msix_table_offset_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_6_vf_msix_table_bir_6                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_6_vf_msix_table_bir_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_6_vf_msix_table_offset_6                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_6_vf_msix_table_offset_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_7_vf_msix_table_bir_7                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_7_vf_msix_table_bir_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_7_vf_msix_table_offset_7                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_msix_table_7_vf_msix_table_offset_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_offset_stride_first_vf_off                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_offset_stride_first_vf_off),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_0_vf_msix_tablesz_0                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_0_vf_msix_tablesz_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_1_vf_msix_tablesz_1                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_1_vf_msix_tablesz_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_2_vf_msix_tablesz_2                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_2_vf_msix_tablesz_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_3_vf_msix_tablesz_3                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_3_vf_msix_tablesz_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_4_vf_msix_tablesz_4                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_4_vf_msix_tablesz_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_5_vf_msix_tablesz_5                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_5_vf_msix_tablesz_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_6_vf_msix_tablesz_6                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_6_vf_msix_tablesz_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_7_vf_msix_tablesz_7                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_capabilities_7_vf_msix_tablesz_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_0_vf_revision_id_0                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_0_vf_revision_id_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_0_vf_subysystem_id_0                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_0_vf_subysystem_id_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_1_vf_revision_id_1                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_1_vf_revision_id_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_1_vf_subysystem_id_1                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_1_vf_subysystem_id_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_2_vf_revision_id_2                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_2_vf_revision_id_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_2_vf_subysystem_id_2                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_2_vf_subysystem_id_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_3_vf_revision_id_3                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_3_vf_revision_id_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_3_vf_subysystem_id_3                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_3_vf_subysystem_id_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_4_vf_revision_id_4                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_4_vf_revision_id_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_4_vf_subysystem_id_4                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_4_vf_subysystem_id_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_5_vf_revision_id_5                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_5_vf_revision_id_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_5_vf_subysystem_id_5                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_5_vf_subysystem_id_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_6_vf_revision_id_6                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_6_vf_revision_id_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_6_vf_subysystem_id_6                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_6_vf_subysystem_id_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_7_vf_revision_id_7                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_7_vf_revision_id_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_7_vf_subysystem_id_7                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_pci_cfg_7_vf_subysystem_id_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_devspecific_mode_0                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_devspecific_mode_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_exttphreq_0                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_exttphreq_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_intvec_mode_0                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_intvec_mode_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_sttable_loc_0                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_sttable_loc_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_sttable_size_0                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_0_vf_tph_sttable_size_0),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_devspecific_mode_1                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_devspecific_mode_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_exttphreq_1                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_exttphreq_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_intvec_mode_1                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_intvec_mode_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_sttable_loc_1                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_sttable_loc_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_sttable_size_1                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_1_vf_tph_sttable_size_1),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_devspecific_mode_2                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_devspecific_mode_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_exttphreq_2                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_exttphreq_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_intvec_mode_2                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_intvec_mode_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_sttable_loc_2                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_sttable_loc_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_sttable_size_2                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_2_vf_tph_sttable_size_2),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_devspecific_mode_3                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_devspecific_mode_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_exttphreq_3                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_exttphreq_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_intvec_mode_3                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_intvec_mode_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_sttable_loc_3                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_sttable_loc_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_sttable_size_3                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_3_vf_tph_sttable_size_3),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_devspecific_mode_4                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_devspecific_mode_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_exttphreq_4                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_exttphreq_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_intvec_mode_4                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_intvec_mode_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_sttable_loc_4                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_sttable_loc_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_sttable_size_4                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_4_vf_tph_sttable_size_4),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_devspecific_mode_5                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_devspecific_mode_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_exttphreq_5                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_exttphreq_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_intvec_mode_5                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_intvec_mode_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_sttable_loc_5                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_sttable_loc_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_sttable_size_5                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_5_vf_tph_sttable_size_5),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_devspecific_mode_6                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_devspecific_mode_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_exttphreq_6                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_exttphreq_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_intvec_mode_6                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_intvec_mode_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_sttable_loc_6                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_sttable_loc_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_sttable_size_6                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_6_vf_tph_sttable_size_6),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_devspecific_mode_7                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_devspecific_mode_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_exttphreq_7                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_exttphreq_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_intvec_mode_7                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_intvec_mode_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_sttable_loc_7                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_sttable_loc_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_sttable_size_7                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf0_vf_tphcap_7_vf_tph_sttable_size_7),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_global_inval_suppport                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_global_inval_suppport),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_inval_queue_dep                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_inval_queue_dep),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_page_aglign_req                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_page_aglign_req),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_ro_support                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_ats_reg_ro_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_devcapreg2_tph_cpl_support                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_devcapreg2_tph_cpl_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_devvendid_deviceid                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_devvendid_deviceid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msi_cap_reg_extnd_msg_data_capable                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msi_cap_reg_extnd_msg_data_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msi_cap_reg_mul_msg_cap                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msi_cap_reg_mul_msg_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msi_cap_reg_per_vector_msk_cap                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msi_cap_reg_per_vector_msk_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_cap_reg_function_mask                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_cap_reg_function_mask),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_cap_reg_table_sz                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_cap_reg_table_sz),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_pba_ptr_pba_bir                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_pba_ptr_pba_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_pba_ptr_pba_offset                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_pba_ptr_pba_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_table_ptr_table_bir                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_table_ptr_table_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_table_ptr_table_offset                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_msix_table_ptr_table_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_revclasscode_class_codes                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_revclasscode_class_codes),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_revclasscode_rid                                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_revclasscode_rid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_siov_dvsec_flags_h                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_siov_dvsec_flags_h),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_siov_dvsec_funtion_dependency_link                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_siov_dvsec_funtion_dependency_link),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_siov_reg3_ims_support                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_siov_reg3_ims_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_sriov_cap_vf_mig_cap                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_sriov_cap_vf_mig_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_sriov_cap_vf_mig_int                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_sriov_cap_vf_mig_int),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_dev_spec_mode_supd                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_dev_spec_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_etph_req_supd                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_etph_req_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_int_vct_mode_supd                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_int_vct_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_st_table_loc                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_st_table_loc),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_tph_st_tab_size                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_tph_req_cap_reg_tph_st_tab_size),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_vf_device_id_vf_device_id                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_vf_device_id_vf_device_id),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_vf_offset_stride_first_vf_off                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf1_vf_offset_stride_first_vf_off),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_global_inval_suppport                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_global_inval_suppport),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_inval_queue_dep                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_inval_queue_dep),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_page_aglign_req                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_page_aglign_req),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_ro_support                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_ats_reg_ro_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_devcapreg2_tph_cpl_support                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_devcapreg2_tph_cpl_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_devvendid_deviceid                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_devvendid_deviceid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msi_cap_reg_extnd_msg_data_capable                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msi_cap_reg_extnd_msg_data_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msi_cap_reg_mul_msg_cap                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msi_cap_reg_mul_msg_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msi_cap_reg_per_vector_msk_cap                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msi_cap_reg_per_vector_msk_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_cap_reg_function_mask                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_cap_reg_function_mask),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_cap_reg_table_sz                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_cap_reg_table_sz),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_pba_ptr_pba_bir                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_pba_ptr_pba_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_pba_ptr_pba_offset                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_pba_ptr_pba_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_table_ptr_table_bir                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_table_ptr_table_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_table_ptr_table_offset                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_msix_table_ptr_table_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_revclasscode_class_codes                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_revclasscode_class_codes),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_revclasscode_rid                                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_revclasscode_rid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_siov_dvsec_flags_h                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_siov_dvsec_flags_h),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_siov_dvsec_funtion_dependency_link                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_siov_dvsec_funtion_dependency_link),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_siov_reg3_ims_support                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_siov_reg3_ims_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_sriov_cap_vf_mig_cap                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_sriov_cap_vf_mig_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_sriov_cap_vf_mig_int                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_sriov_cap_vf_mig_int),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_dev_spec_mode_supd                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_dev_spec_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_etph_req_supd                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_etph_req_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_int_vct_mode_supd                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_int_vct_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_st_table_loc                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_st_table_loc),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_tph_st_tab_size                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_tph_req_cap_reg_tph_st_tab_size),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_vf_device_id_vf_device_id                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_vf_device_id_vf_device_id),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_vf_offset_stride_first_vf_off                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf2_vf_offset_stride_first_vf_off),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_global_inval_suppport                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_global_inval_suppport),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_inval_queue_dep                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_inval_queue_dep),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_page_aglign_req                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_page_aglign_req),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_ro_support                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_ats_reg_ro_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_devcapreg2_tph_cpl_support                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_devcapreg2_tph_cpl_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_devvendid_deviceid                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_devvendid_deviceid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msi_cap_reg_extnd_msg_data_capable                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msi_cap_reg_extnd_msg_data_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msi_cap_reg_mul_msg_cap                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msi_cap_reg_mul_msg_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msi_cap_reg_per_vector_msk_cap                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msi_cap_reg_per_vector_msk_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_cap_reg_function_mask                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_cap_reg_function_mask),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_cap_reg_table_sz                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_cap_reg_table_sz),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_pba_ptr_pba_bir                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_pba_ptr_pba_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_pba_ptr_pba_offset                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_pba_ptr_pba_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_table_ptr_table_bir                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_table_ptr_table_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_table_ptr_table_offset                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_msix_table_ptr_table_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_revclasscode_class_codes                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_revclasscode_class_codes),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_revclasscode_rid                                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_revclasscode_rid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_siov_dvsec_flags_h                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_siov_dvsec_flags_h),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_siov_dvsec_funtion_dependency_link                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_siov_dvsec_funtion_dependency_link),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_siov_reg3_ims_support                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_siov_reg3_ims_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_sriov_cap_vf_mig_cap                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_sriov_cap_vf_mig_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_sriov_cap_vf_mig_int                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_sriov_cap_vf_mig_int),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_dev_spec_mode_supd                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_dev_spec_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_etph_req_supd                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_etph_req_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_int_vct_mode_supd                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_int_vct_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_st_table_loc                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_st_table_loc),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_tph_st_tab_size                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_tph_req_cap_reg_tph_st_tab_size),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_vf_device_id_vf_device_id                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_vf_device_id_vf_device_id),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_vf_offset_stride_first_vf_off                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf3_vf_offset_stride_first_vf_off),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_global_inval_suppport                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_global_inval_suppport),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_inval_queue_dep                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_inval_queue_dep),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_page_aglign_req                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_page_aglign_req),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_ro_support                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_ats_reg_ro_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_devcapreg2_tph_cpl_support                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_devcapreg2_tph_cpl_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_devvendid_deviceid                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_devvendid_deviceid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msi_cap_reg_extnd_msg_data_capable                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msi_cap_reg_extnd_msg_data_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msi_cap_reg_mul_msg_cap                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msi_cap_reg_mul_msg_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msi_cap_reg_per_vector_msk_cap                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msi_cap_reg_per_vector_msk_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_cap_reg_function_mask                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_cap_reg_function_mask),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_cap_reg_table_sz                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_cap_reg_table_sz),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_pba_ptr_pba_bir                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_pba_ptr_pba_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_pba_ptr_pba_offset                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_pba_ptr_pba_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_table_ptr_table_bir                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_table_ptr_table_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_table_ptr_table_offset                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_msix_table_ptr_table_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_revclasscode_class_codes                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_revclasscode_class_codes),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_revclasscode_rid                                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_revclasscode_rid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_siov_dvsec_flags_h                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_siov_dvsec_flags_h),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_siov_dvsec_funtion_dependency_link                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_siov_dvsec_funtion_dependency_link),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_siov_reg3_ims_support                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_siov_reg3_ims_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_sriov_cap_vf_mig_cap                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_sriov_cap_vf_mig_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_sriov_cap_vf_mig_int                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_sriov_cap_vf_mig_int),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_dev_spec_mode_supd                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_dev_spec_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_etph_req_supd                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_etph_req_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_int_vct_mode_supd                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_int_vct_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_st_table_loc                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_st_table_loc),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_tph_st_tab_size                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_tph_req_cap_reg_tph_st_tab_size),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_vf_device_id_vf_device_id                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_vf_device_id_vf_device_id),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_vf_offset_stride_first_vf_off                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf4_vf_offset_stride_first_vf_off),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_global_inval_suppport                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_global_inval_suppport),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_inval_queue_dep                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_inval_queue_dep),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_page_aglign_req                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_page_aglign_req),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_ro_support                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_ats_reg_ro_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_devcapreg2_tph_cpl_support                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_devcapreg2_tph_cpl_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_devvendid_deviceid                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_devvendid_deviceid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msi_cap_reg_extnd_msg_data_capable                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msi_cap_reg_extnd_msg_data_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msi_cap_reg_mul_msg_cap                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msi_cap_reg_mul_msg_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msi_cap_reg_per_vector_msk_cap                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msi_cap_reg_per_vector_msk_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_cap_reg_function_mask                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_cap_reg_function_mask),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_cap_reg_table_sz                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_cap_reg_table_sz),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_pba_ptr_pba_bir                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_pba_ptr_pba_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_pba_ptr_pba_offset                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_pba_ptr_pba_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_table_ptr_table_bir                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_table_ptr_table_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_table_ptr_table_offset                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_msix_table_ptr_table_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_revclasscode_class_codes                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_revclasscode_class_codes),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_revclasscode_rid                                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_revclasscode_rid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_siov_dvsec_flags_h                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_siov_dvsec_flags_h),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_siov_dvsec_funtion_dependency_link                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_siov_dvsec_funtion_dependency_link),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_siov_reg3_ims_support                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_siov_reg3_ims_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_sriov_cap_vf_mig_cap                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_sriov_cap_vf_mig_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_sriov_cap_vf_mig_int                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_sriov_cap_vf_mig_int),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_dev_spec_mode_supd                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_dev_spec_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_etph_req_supd                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_etph_req_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_int_vct_mode_supd                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_int_vct_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_st_table_loc                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_st_table_loc),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_tph_st_tab_size                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_tph_req_cap_reg_tph_st_tab_size),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_vf_device_id_vf_device_id                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_vf_device_id_vf_device_id),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_vf_offset_stride_first_vf_off                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf5_vf_offset_stride_first_vf_off),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_global_inval_suppport                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_global_inval_suppport),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_inval_queue_dep                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_inval_queue_dep),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_page_aglign_req                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_page_aglign_req),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_ro_support                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_ats_reg_ro_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_devcapreg2_tph_cpl_support                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_devcapreg2_tph_cpl_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_devvendid_deviceid                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_devvendid_deviceid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msi_cap_reg_extnd_msg_data_capable                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msi_cap_reg_extnd_msg_data_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msi_cap_reg_mul_msg_cap                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msi_cap_reg_mul_msg_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msi_cap_reg_per_vector_msk_cap                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msi_cap_reg_per_vector_msk_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_cap_reg_function_mask                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_cap_reg_function_mask),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_cap_reg_table_sz                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_cap_reg_table_sz),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_pba_ptr_pba_bir                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_pba_ptr_pba_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_pba_ptr_pba_offset                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_pba_ptr_pba_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_table_ptr_table_bir                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_table_ptr_table_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_table_ptr_table_offset                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_msix_table_ptr_table_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_revclasscode_class_codes                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_revclasscode_class_codes),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_revclasscode_rid                                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_revclasscode_rid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_siov_dvsec_flags_h                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_siov_dvsec_flags_h),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_siov_dvsec_funtion_dependency_link                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_siov_dvsec_funtion_dependency_link),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_siov_reg3_ims_support                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_siov_reg3_ims_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_sriov_cap_vf_mig_cap                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_sriov_cap_vf_mig_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_sriov_cap_vf_mig_int                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_sriov_cap_vf_mig_int),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_dev_spec_mode_supd                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_dev_spec_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_etph_req_supd                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_etph_req_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_int_vct_mode_supd                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_int_vct_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_st_table_loc                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_st_table_loc),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_tph_st_tab_size                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_tph_req_cap_reg_tph_st_tab_size),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_vf_device_id_vf_device_id                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_vf_device_id_vf_device_id),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_vf_offset_stride_first_vf_off                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf6_vf_offset_stride_first_vf_off),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_global_inval_suppport                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_global_inval_suppport),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_inval_queue_dep                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_inval_queue_dep),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_page_aglign_req                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_page_aglign_req),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_ro_support                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_ats_reg_ro_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_devcapreg2_tph_cpl_support                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_devcapreg2_tph_cpl_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_devvendid_deviceid                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_devvendid_deviceid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msi_cap_reg_extnd_msg_data_capable                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msi_cap_reg_extnd_msg_data_capable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msi_cap_reg_mul_msg_cap                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msi_cap_reg_mul_msg_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msi_cap_reg_per_vector_msk_cap                                            ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msi_cap_reg_per_vector_msk_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_cap_reg_function_mask                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_cap_reg_function_mask),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_cap_reg_table_sz                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_cap_reg_table_sz),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_pba_ptr_pba_bir                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_pba_ptr_pba_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_pba_ptr_pba_offset                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_pba_ptr_pba_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_table_ptr_table_bir                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_table_ptr_table_bir),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_table_ptr_table_offset                                               ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_msix_table_ptr_table_offset),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_revclasscode_class_codes                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_revclasscode_class_codes),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_revclasscode_rid                                                          ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_revclasscode_rid),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_siov_dvsec_flags_h                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_siov_dvsec_flags_h),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_siov_dvsec_funtion_dependency_link                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_siov_dvsec_funtion_dependency_link),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_siov_reg3_ims_support                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_siov_reg3_ims_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_sriov_cap_vf_mig_cap                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_sriov_cap_vf_mig_cap),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_sriov_cap_vf_mig_int                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_sriov_cap_vf_mig_int),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_dev_spec_mode_supd                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_dev_spec_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_etph_req_supd                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_etph_req_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_int_vct_mode_supd                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_int_vct_mode_supd),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_st_table_loc                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_st_table_loc),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_tph_st_tab_size                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_tph_req_cap_reg_tph_st_tab_size),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_vf_device_id_vf_device_id                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_vf_device_id_vf_device_id),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_vf_offset_stride_first_vf_off                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pf7_vf_offset_stride_first_vf_off),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pld_sbep_portid_k_pld_sbep_id                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_pld_sbep_portid_k_pld_sbep_id),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_powerdown_mode                                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_powerdown_mode),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_r_spare_ctl2_k_r_spare_ctl2                                                   ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_r_spare_ctl2_k_r_spare_ctl2)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_reset_csr_k_pld_crs_en                                                        ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_reset_csr_k_pld_crs_en),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_sup_mode                                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_sup_mode),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_addr_a2a3_data_pack                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_addr_a2a3_data_pack),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_acs_next_ptr                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_acs_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_aer_next_ptr                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_aer_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_ats_next_ptr                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_ats_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_cxl_next_ptr                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_cxl_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_ltr_next_ptr                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_ltr_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_msi_next_ptr                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_msi_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_msix_next_ptr                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_msix_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pasid_next_ptr                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pasid_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pcie_next_ptr                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pcie_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pm_next_ptr                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pm_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pri_next_ptr                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_pri_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_ptm_next_ptr                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_ptm_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_siov_next_ptr                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_siov_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_sriov_next_ptr                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_sriov_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_tph_next_ptr                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_tph_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_vc_next_ptr                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cfg_ext_vc_next_ptr),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cvp_bar_num                                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cvp_bar_num),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cvp_mode                                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_cvp_mode),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_functional_mode                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_functional_mode),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_maxpayload_size                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_maxpayload_size),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_num_of_pf                                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_num_of_pf),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_acs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_aer_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_aer_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_ats_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar1_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar1_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar1_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar3_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar3_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar3_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar5_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar5_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar5_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_cxl_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_cxl_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_expansion_rom_enable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_expansion_rom_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_expansion_rom_mask                                                ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_expansion_rom_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_ltr_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_ltr_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_msi_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_msi_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_msix_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_num_of_vf                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_num_of_vf),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_pasid_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_pasid_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_prs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_prs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_ptm_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_ptm_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_siov_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_siov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_sriov_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_sriov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_tph_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vc_cap_enable                                                     ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vc_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_acs_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_ats_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar1_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar1_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar1_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar3_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar3_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar3_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar5_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar5_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar5_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_msix_cap_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_tph_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf0_vf_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_acs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_aer_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_aer_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_ats_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar1_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar1_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar1_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar3_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar3_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar3_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar5_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar5_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar5_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_msi_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_msi_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_msix_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_num_of_vf                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_num_of_vf),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_pasid_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_pasid_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_prs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_prs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_siov_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_siov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_sriov_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_sriov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_tph_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_acs_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_ats_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar1_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar1_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar1_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar3_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar3_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar3_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar5_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar5_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar5_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_msix_cap_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_tph_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf1_vf_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_acs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_aer_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_aer_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_ats_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar1_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar1_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar1_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar3_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar3_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar3_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar5_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar5_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar5_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_msi_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_msi_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_msix_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_num_of_vf                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_num_of_vf),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_pasid_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_pasid_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_prs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_prs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_siov_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_siov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_sriov_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_sriov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_tph_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_acs_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_ats_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar1_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar1_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar1_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar3_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar3_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar3_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar5_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar5_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar5_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_msix_cap_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_tph_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf2_vf_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_acs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_aer_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_aer_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_ats_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar1_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar1_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar1_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar3_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar3_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar3_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar5_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar5_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar5_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_msi_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_msi_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_msix_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_num_of_vf                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_num_of_vf),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_pasid_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_pasid_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_prs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_prs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_siov_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_siov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_sriov_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_sriov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_tph_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_acs_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_ats_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar1_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar1_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar1_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar3_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar3_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar3_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar5_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar5_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar5_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_msix_cap_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_tph_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf3_vf_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_acs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_aer_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_aer_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_ats_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar1_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar1_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar1_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar3_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar3_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar3_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar5_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar5_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar5_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_msi_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_msi_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_msix_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_num_of_vf                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_num_of_vf),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_pasid_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_pasid_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_prs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_prs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_siov_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_siov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_sriov_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_sriov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_tph_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_acs_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_ats_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar1_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar1_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar1_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar3_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar3_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar3_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar5_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar5_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar5_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_msix_cap_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_tph_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf4_vf_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_acs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_aer_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_aer_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_ats_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar1_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar1_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar1_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar3_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar3_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar3_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar5_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar5_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar5_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_msi_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_msi_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_msix_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_num_of_vf                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_num_of_vf),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_pasid_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_pasid_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_prs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_prs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_siov_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_siov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_sriov_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_sriov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_tph_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_acs_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_ats_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar1_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar1_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar1_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar3_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar3_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar3_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar5_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar5_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar5_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_msix_cap_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_tph_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf5_vf_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_acs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_aer_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_aer_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_ats_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar1_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar1_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar1_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar3_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar3_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar3_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar5_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar5_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar5_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_msi_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_msi_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_msix_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_num_of_vf                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_num_of_vf),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_pasid_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_pasid_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_prs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_prs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_siov_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_siov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_sriov_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_sriov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_tph_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_acs_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_ats_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar1_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar1_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar1_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar3_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar3_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar3_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar5_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar5_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar5_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_msix_cap_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_tph_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf6_vf_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_acs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_aer_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_aer_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_ats_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar1_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar1_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar1_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar3_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar3_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar3_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_64b_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar5_enable                                                       ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar5_mask                                                         ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar5_prefetchable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_msi_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_msi_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_msix_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_num_of_vf                                                         ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_num_of_vf),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_pasid_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_pasid_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_prs_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_prs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_siov_cap_enable                                                   ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_siov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_sriov_cap_enable                                                  ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_sriov_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_tph_cap_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_acs_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_acs_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_ats_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_ats_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar0_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar1_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar1_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar1_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar1_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar1_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar1_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar2_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar3_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar3_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar3_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar3_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar3_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar3_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_64b_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_64b_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar4_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar5_enable                                                    ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar5_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar5_mask                                                      ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar5_mask)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar5_prefetchable                                              ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_bar5_prefetchable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_msix_cap_enable                                                ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_msix_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_tph_cap_enable                                                 ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pf7_vf_tph_cap_enable),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pri_out_pagereq_capacity                                              ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_pri_out_pagereq_capacity)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_ptile_header_fmt                                                      ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_ptile_header_fmt),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_supported_page_size                                                   ( str_2_bin(hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_supported_page_size)),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_tag_support                                                           ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_rnr_pialup_inst_virtual_tag_support),
   .hssi_ctr_u_ial_top_rnr_ialup_icm_inst_target_link_speed                                                                             ( hssi_ctr_u_ial_top_rnr_ialup_icm_inst_target_link_speed),
   .hssi_ctr_u_ial_top_sup_mode                                                                                                         ( hssi_ctr_u_ial_top_sup_mode),
   .hssi_ctr_u_pcie_top_powerdown_mode                                                                                                  ( hssi_ctr_u_pcie_top_powerdown_mode),
   .hssi_ctr_u_pcie_top_ptm_enable                                                                                                      ( hssi_ctr_u_pcie_top_ptm_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_avmm_ctrl_k_rstrdy_resp_en_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_avmm_ctrl_k_rstrdy_resp_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_avmm_ctrl_k_security_bypass_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_avmm_ctrl_k_security_bypass_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p0_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p1_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p2_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p3_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_deskew_ctrl_k_dskw_force_done_p3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_dfd_en_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_dfd_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_dfd_patcntr_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_dfd_patcntr_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar0_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar0_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar1_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar1_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar2_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar2_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar3_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl1_k_xbar3_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane0_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane0_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane1_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane1_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane2_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane2_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane3_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl2_k_lane3_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl3_k_trig0_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl3_k_trig0_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl3_k_trig1_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl3_k_trig1_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q0_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q0_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q1_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q1_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q2_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q2_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q3_sel_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_dfdmux_ctrl_k_dfd_q3_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_aib_sel_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_aib_sel_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_error_mask_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_error_mask_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_sts_cor_en_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_sts_cor_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_sts_uc_en_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_ecc_sts_uc_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_nparity_ecc_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_nparity_ecc_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_par_sts_uc_en_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_ecc_ctrl_k_par_sts_uc_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_hw_mode_override_en                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_cfgtop_inst_hw_mode_override_en),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf0_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf1_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf2_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf3_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf4_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf5_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf6_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf7_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf7_attr),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_0_k_cii_addr_size0_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_0_k_cii_addr_size0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_0_k_cii_pf_en0_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_0_k_cii_pf_en0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_0_k_cii_start_addr0_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_0_k_cii_start_addr0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_1_k_cii_addr_size1_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_1_k_cii_addr_size1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_1_k_cii_pf_en1_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_1_k_cii_pf_en1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_1_k_cii_start_addr1_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_1_k_cii_start_addr1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_2_k_cii_addr_size2_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_2_k_cii_addr_size2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_2_k_cii_pf_en2_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_2_k_cii_pf_en2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_2_k_cii_start_addr2_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_2_k_cii_start_addr2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_3_k_cii_addr_size3_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_3_k_cii_addr_size3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_3_k_cii_pf_en3_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_3_k_cii_pf_en3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_3_k_cii_start_addr3_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_3_k_cii_start_addr3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_4_k_cii_addr_size4_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_4_k_cii_addr_size4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_4_k_cii_pf_en4_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_4_k_cii_pf_en4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_4_k_cii_start_addr4_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_4_k_cii_start_addr4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_5_k_cii_addr_size5_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_5_k_cii_addr_size5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_5_k_cii_pf_en5_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_5_k_cii_pf_en5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_5_k_cii_start_addr5_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_5_k_cii_start_addr5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_6_k_cii_addr_size6_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_6_k_cii_addr_size6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_6_k_cii_pf_en6_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_6_k_cii_pf_en6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_6_k_cii_start_addr6_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_6_k_cii_start_addr6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_7_k_cii_addr_size7_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_7_k_cii_addr_size7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_7_k_cii_pf_en7_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_7_k_cii_pf_en7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_7_k_cii_start_addr7_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cii_range_7_k_cii_start_addr7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_fixedcred_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_fixedcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_mcred_attr                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_mcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_reloadcred_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_reloadcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_tlp_serr_dis_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_ctrl0_k_tlp_serr_dis_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_mmio_access_ctrl_grant_attr                                         ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_mmio_access_ctrl_grant_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_opcode_ctrl_lock_attr                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_csb_opcode_ctrl_lock_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_bar0_k_cvp_bar_0_attr                                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_bar0_k_cvp_bar_0_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_bar1_k_cvp_bar_1_attr                                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_bar1_k_cvp_bar_1_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctl_k_cvp_bar_mode_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctl_k_cvp_bar_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctl_k_cvp_bar_type_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctl_k_cvp_bar_type_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctl_k_cvp_bar_used_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctl_k_cvp_bar_used_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl0_k_compressed_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl0_k_compressed_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl0_k_encrypted_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl0_k_encrypted_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl1_k_devbrd_type_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl1_k_devbrd_type_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl1_k_vsec_next_offset_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_ctrl1_k_vsec_next_offset_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_irq_ctrl_k_cvp_irq_en_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_irq_ctrl_k_cvp_irq_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_irq_ctrl_k_gpio_irq_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_irq_ctrl_k_gpio_irq_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_jtagid0_k_jtag_id_0_attr                                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_cvp_jtagid0_k_jtag_id_0_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_ctrl0_k_dfd_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_ctrl0_k_dfd_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_ctrl0_k_patcntr_en_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_ctrl0_k_patcntr_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_0_attr                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_1_attr                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_2_attr                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_3_attr                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_data_sel_3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_trig_sel_0_attr                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_trig_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_trig_sel_1_attr                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_trig_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_0_attr                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_1_attr                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_2_attr                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_3_attr                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dfd_xbar_sel_3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_pld_crs_en_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_pld_crs_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_rx_lane_flip_en_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_rx_lane_flip_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_sris_mode_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_sris_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_tx_lane_flip_en_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_dwc_ctrl0_k_tx_lane_flip_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ehp_ctrl0_k_ehp_control_reg_attr                                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ehp_ctrl0_k_ehp_control_reg_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ehp_ctrl1_k_outstanding_crd_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ehp_ctrl1_k_outstanding_crd_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ehp_ctrl1_k_tx_rd_th_attr                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ehp_ctrl1_k_tx_rd_th_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff0_k_exvf_msixpba_bir_pf0_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff0_k_exvf_msixpba_bir_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff0_k_exvf_msixpba_offset_pf0_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff0_k_exvf_msixpba_offset_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff1_k_exvf_msixpba_bir_pf1_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff1_k_exvf_msixpba_bir_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff1_k_exvf_msixpba_offset_pf1_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff1_k_exvf_msixpba_offset_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff2_k_exvf_msixpba_bir_pf2_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff2_k_exvf_msixpba_bir_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff2_k_exvf_msixpba_offset_pf2_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff2_k_exvf_msixpba_offset_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff3_k_exvf_msixpba_bir_pf3_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff3_k_exvf_msixpba_bir_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff3_k_exvf_msixpba_offset_pf3_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff3_k_exvf_msixpba_offset_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff4_k_exvf_msixpba_bir_pf4_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff4_k_exvf_msixpba_bir_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff4_k_exvf_msixpba_offset_pf4_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff4_k_exvf_msixpba_offset_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff5_k_exvf_msixpba_bir_pf5_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff5_k_exvf_msixpba_bir_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff5_k_exvf_msixpba_offset_pf5_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff5_k_exvf_msixpba_offset_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff6_k_exvf_msixpba_bir_pf6_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff6_k_exvf_msixpba_bir_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff6_k_exvf_msixpba_offset_pf6_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff6_k_exvf_msixpba_offset_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff7_k_exvf_msixpba_bir_pf7_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff7_k_exvf_msixpba_bir_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff7_k_exvf_msixpba_offset_pf7_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_poff7_k_exvf_msixpba_offset_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff0_k_exvf_msixtable_bir_pf0_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff0_k_exvf_msixtable_bir_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff0_k_exvf_msixtable_offset_pf0_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff0_k_exvf_msixtable_offset_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff1_k_exvf_msixtable_bir_pf1_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff1_k_exvf_msixtable_bir_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff1_k_exvf_msixtable_offset_pf1_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff1_k_exvf_msixtable_offset_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff2_k_exvf_msixtable_bir_pf2_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff2_k_exvf_msixtable_bir_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff2_k_exvf_msixtable_offset_pf2_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff2_k_exvf_msixtable_offset_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff3_k_exvf_msixtable_bir_pf3_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff3_k_exvf_msixtable_bir_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff3_k_exvf_msixtable_offset_pf3_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff3_k_exvf_msixtable_offset_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff4_k_exvf_msixtable_bir_pf4_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff4_k_exvf_msixtable_bir_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff4_k_exvf_msixtable_offset_pf4_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff4_k_exvf_msixtable_offset_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff5_k_exvf_msixtable_bir_pf5_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff5_k_exvf_msixtable_bir_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff5_k_exvf_msixtable_offset_pf5_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff5_k_exvf_msixtable_offset_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff6_k_exvf_msixtable_bir_pf6_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff6_k_exvf_msixtable_bir_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff6_k_exvf_msixtable_offset_pf6_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff6_k_exvf_msixtable_offset_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff7_k_exvf_msixtable_bir_pf7_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff7_k_exvf_msixtable_bir_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff7_k_exvf_msixtable_offset_pf7_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_toff7_k_exvf_msixtable_offset_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize0_k_exvf_msix_tablesize_pf0_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize0_k_exvf_msix_tablesize_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize0_k_exvf_msix_tablesize_pf1_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize0_k_exvf_msix_tablesize_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize1_k_exvf_msix_tablesize_pf2_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize1_k_exvf_msix_tablesize_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize1_k_exvf_msix_tablesize_pf3_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize1_k_exvf_msix_tablesize_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize2_k_exvf_msix_tablesize_pf4_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize2_k_exvf_msix_tablesize_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize2_k_exvf_msix_tablesize_pf5_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize2_k_exvf_msix_tablesize_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize3_k_exvf_msix_tablesize_pf6_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize3_k_exvf_msix_tablesize_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize3_k_exvf_msix_tablesize_pf7_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_m6_tsize3_k_exvf_msix_tablesize_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_cvp_cfg_err_en_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_cvp_cfg_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_dbi_access_err_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_dbi_access_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sd_eq_control1_reg_eval_interval_time),
   
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_multi_lane_control_off_upconfigure_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_multi_lane_control_off_upconfigure_support),
   
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_reg_bar0_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_reg_bar0_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar1_reg_bar1_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_reg_bar2_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_reg_bar2_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_reg_bar3_mem_io                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_reg_bar3_mem_io),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_reg_bar3_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_reg_bar4_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_reg_bar4_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar5_reg_bar5_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_id_nxt_ptr_reg_aux_curr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_id_nxt_ptr_reg_dsi                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_id_nxt_ptr_reg_pme_support                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_reg_ari_acs_fun_grp_cap                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_cap_reg_ari_acs_fun_grp_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_base_class_code                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_program_interface                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_revision_id                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_subclass_code                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_con_status_reg_no_soft_rst                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_exp_rom_bar_mask_reg_rom_mask                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen2_ctrl_off_config_phy_tx_change                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen2_ctrl_off_config_phy_tx_change),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen2_ctrl_off_support_mod_ts                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen2_ctrl_off_support_mod_ts),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_eieos_cnt                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_eieos_cnt),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_phase_2_3                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_phase_2_3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_phase_2_3_atg4                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_phase_2_3_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_phase_2_3_atg5                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_phase_2_3_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_redo                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_redo),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_redo_atg4                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_redo_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_redo_atg5                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_eq_redo_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_gen3_equalization_disable                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_gen3_equalization_disable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_ph01_en                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_ph01_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1_substates_off_l1sub_t_l1_2                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1_substates_off_l1sub_t_l1_2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1_substates_off_l1sub_t_power_off                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1_substates_off_l1sub_t_power_off),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_comm_mode_support                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_comm_mode_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_pwr_on_scale_support                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_pwr_on_scale_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_pwr_on_value_support                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_pwr_on_value_support),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_1_aspm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_1_aspm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_2_aspm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_2_aspm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_1_aspm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_1_aspm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_aspm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_aspm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_l1_1sub_cap_enable ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_l1_1sub_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_l1_2sub_cap_enable ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_l1_2sub_cap_enable),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_th_sca                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_th_sca),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_th_val                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_l1_2_th_val),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_t_common_mode                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_l1sub_control1_reg_t_common_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_port_num                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_table_offset_reg_pci_msix_bir                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_table_offset_reg_pci_msix_table_offset                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pipe_loopback_control_off_pipe_loopback                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pipe_loopback_control_off_pipe_loopback),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset4                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset5                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset6                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset7                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset4                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset5                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset6                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset7                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset10                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset10),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset11                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset8                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset8),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset9                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_dsp_16g_tx_preset9),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset10                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset10),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset11                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset8                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset8),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset9                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_28h_reg_usp_16g_tx_preset9),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset12                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset12),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset13                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset13),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset14                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset14),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset15                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_dsp_16g_tx_preset15),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset12                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset12),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset13                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset13),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset14                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset14),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset15                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl16g_cap_off_2ch_reg_usp_16g_tx_preset15),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset4                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset5                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset6                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset7                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset4                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset5                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset6                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset7                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset10                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset10),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset11                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset8                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset8),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset9                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_dsp_32g_tx_preset9),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset10                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset10),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset11                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset8                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset8),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset9                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_28h_reg_usp_32g_tx_preset9),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset12                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset12),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset13                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset13),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset14                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset14),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset15                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_dsp_32g_tx_preset15),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset12                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset12),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset13                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset13),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset14                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset14),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset15                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_cap_off_2ch_reg_usp_32g_tx_preset15),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_capability_reg_no_eq_needed_support                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_capability_reg_no_eq_needed_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_rsvdp_11                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_rsvdp_11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_tx_precode_req                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_tx_precode_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_tx_precoding_on                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_pl32g_status_reg_tx_precoding_on),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_port_link_ctrl_off_fast_link_mode                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_port_link_ctrl_off_fast_link_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint4                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint5                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset4                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset5                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint4                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint5                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset4                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset5                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint6                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint7                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset6                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset7                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint6                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint7                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset6                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset7                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_rx_preset_hint8                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_rx_preset_hint8),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_rx_preset_hint9                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_rx_preset_hint9),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_tx_preset8                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_tx_preset8),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_tx_preset9                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_dsp_tx_preset9),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_rx_preset_hint8                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_rx_preset_hint8),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_rx_preset_hint9                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_rx_preset_hint9),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_tx_preset8                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_tx_preset8),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_tx_preset9                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_1ch_reg_usp_tx_preset9),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_rx_preset_hint10                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_rx_preset_hint10),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_rx_preset_hint11                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_rx_preset_hint11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_tx_preset10                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_tx_preset10),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_tx_preset11                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_dsp_tx_preset11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_rx_preset_hint10                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_rx_preset_hint10),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_rx_preset_hint11                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_rx_preset_hint11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_tx_preset10                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_tx_preset10),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_tx_preset11                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_20h_reg_usp_tx_preset11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_rx_preset_hint12                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_rx_preset_hint12),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_rx_preset_hint13                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_rx_preset_hint13),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_tx_preset12                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_tx_preset12),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_tx_preset13                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_dsp_tx_preset13),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_rx_preset_hint12                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_rx_preset_hint12),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_rx_preset_hint13                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_rx_preset_hint13),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_tx_preset12                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_tx_preset12),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_tx_preset13                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_24h_reg_usp_tx_preset13),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_rx_preset_hint14                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_rx_preset_hint14),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_rx_preset_hint15                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_rx_preset_hint15),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_tx_preset14                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_tx_preset14),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_tx_preset15                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_dsp_tx_preset15),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_rx_preset_hint14                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_rx_preset_hint14),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_rx_preset_hint15                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_rx_preset_hint15),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_tx_preset14                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_tx_preset14),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_tx_preset15                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_spcie_cap_off_28h_reg_usp_tx_preset15),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar0_mask_reg_pci_sriov_bar0_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar1_mask_reg_pci_sriov_bar1_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar1_reg_sriov_vf_bar1_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar2_mask_reg_pci_sriov_bar2_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar3_mask_reg_pci_sriov_bar3_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar3_reg_sriov_vf_bar3_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar4_mask_reg_pci_sriov_bar4_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar5_mask_reg_pci_sriov_bar5_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar5_reg_sriov_vf_bar5_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_vf_offset_position_sriov_vf_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_vf_offset_position_sriov_vf_stride                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sup_page_sizes_reg_sriov_sup_page_size                              ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_vf_device_id_reg_sriov_vf_device_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf0_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_at_block                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_egress_control                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_src_valid                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_usp_forwarding                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ats_capabilities_ctrl_reg_invalidate_q_depth                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ats_capabilities_ctrl_reg_page_aligned_req                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_mask_reg_pci_type0_bar0_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_mask_reg_pci_type0_bar0_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_reg_bar0_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_reg_bar0_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar1_mask_reg_pci_type0_bar1_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar1_mask_reg_pci_type0_bar1_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar1_reg_bar1_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_mask_reg_pci_type0_bar2_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_mask_reg_pci_type0_bar2_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_reg_bar2_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_reg_bar2_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar3_mask_reg_pci_type0_bar3_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar3_mask_reg_pci_type0_bar3_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar3_reg_bar3_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_mask_reg_pci_type0_bar4_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_mask_reg_pci_type0_bar4_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_reg_bar4_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_reg_bar4_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar5_mask_reg_pci_type0_bar5_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar5_mask_reg_pci_type0_bar5_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar5_reg_bar5_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cap_id_nxt_ptr_reg_aux_curr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cap_id_nxt_ptr_reg_dsi                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cap_id_nxt_ptr_reg_pme_support                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cardbus_cis_ptr_reg_cardbus_cis_pointer                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_base_class_code                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_program_interface                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_revision_id                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_subclass_code                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_con_status_reg_no_soft_rst                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_capabilities_reg_pcie_cap_flr_cap                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_control_device_status_pcie_cap_ext_tag_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_id_vendor_id_reg_pci_type0_device_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_id_vendor_id_reg_pci_type0_vendor_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_bar_mask_reg_rom_bar_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_bar_mask_reg_rom_mask                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_base_addr_reg_exp_rom_base_address                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_base_addr_reg_exp_rom_base_address),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_base_addr_reg_rom_bar_enable                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_capabilities_reg_pcie_cap_l0s_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_capabilities_reg_pcie_cap_l1_exit_latency                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_capabilities_reg_pcie_cap_port_num                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_control2_link_status2_reg_pcie_cap_sel_deemphasis              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_control_link_status_reg_pcie_cap_active_state_link_pm_control  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_control_link_status_reg_pcie_cap_slot_clk_config               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_pba_offset_reg_pci_msix_pba_bir                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_pba_offset_reg_pci_msix_pba_offset                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_table_offset_reg_pci_msix_bir                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_table_offset_reg_pci_msix_table_offset                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pasid_cap_cntrl_reg_execute_permission_supported                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pasid_cap_cntrl_reg_max_pasid_width                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pasid_cap_cntrl_reg_privileged_mode_supported                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_device_spec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar0_mask_reg_pci_sriov_bar0_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar1_mask_reg_pci_sriov_bar1_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar1_reg_sriov_vf_bar1_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar2_mask_reg_pci_sriov_bar2_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar3_mask_reg_pci_sriov_bar3_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar3_reg_sriov_vf_bar3_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar4_mask_reg_pci_sriov_bar4_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar5_mask_reg_pci_sriov_bar5_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar5_reg_sriov_vf_bar5_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_vf_offset_position_sriov_vf_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_vf_offset_position_sriov_vf_stride                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sup_page_sizes_reg_sriov_sup_page_size                              ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_int_vec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_size                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_device_spec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_vf_device_id_reg_sriov_vf_device_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf1_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_at_block                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_egress_control                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_src_valid                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_usp_forwarding                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ats_capabilities_ctrl_reg_invalidate_q_depth                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ats_capabilities_ctrl_reg_page_aligned_req                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_mask_reg_pci_type0_bar0_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_mask_reg_pci_type0_bar0_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_reg_bar0_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_reg_bar0_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar1_mask_reg_pci_type0_bar1_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar1_mask_reg_pci_type0_bar1_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar1_reg_bar1_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_mask_reg_pci_type0_bar2_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_mask_reg_pci_type0_bar2_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_reg_bar2_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_reg_bar2_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar3_mask_reg_pci_type0_bar3_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar3_mask_reg_pci_type0_bar3_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar3_reg_bar3_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_mask_reg_pci_type0_bar4_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_mask_reg_pci_type0_bar4_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_reg_bar4_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_reg_bar4_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar5_mask_reg_pci_type0_bar5_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar5_mask_reg_pci_type0_bar5_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar5_reg_bar5_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cap_id_nxt_ptr_reg_aux_curr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cap_id_nxt_ptr_reg_dsi                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cap_id_nxt_ptr_reg_pme_support                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cardbus_cis_ptr_reg_cardbus_cis_pointer                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_base_class_code                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_program_interface                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_revision_id                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_subclass_code                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_con_status_reg_no_soft_rst                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_capabilities_reg_pcie_cap_flr_cap                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_control_device_status_pcie_cap_ext_tag_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_id_vendor_id_reg_pci_type0_device_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_id_vendor_id_reg_pci_type0_vendor_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_bar_mask_reg_rom_bar_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_bar_mask_reg_rom_mask                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_base_addr_reg_exp_rom_base_address                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_base_addr_reg_exp_rom_base_address),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_base_addr_reg_rom_bar_enable                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_capabilities_reg_pcie_cap_l0s_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_capabilities_reg_pcie_cap_l1_exit_latency                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_capabilities_reg_pcie_cap_port_num                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_control2_link_status2_reg_pcie_cap_sel_deemphasis              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_control_link_status_reg_pcie_cap_active_state_link_pm_control  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_control_link_status_reg_pcie_cap_slot_clk_config               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_pba_offset_reg_pci_msix_pba_bir                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_pba_offset_reg_pci_msix_pba_offset                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_table_offset_reg_pci_msix_bir                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_table_offset_reg_pci_msix_table_offset                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pasid_cap_cntrl_reg_execute_permission_supported                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pasid_cap_cntrl_reg_max_pasid_width                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pasid_cap_cntrl_reg_privileged_mode_supported                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_device_spec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar0_mask_reg_pci_sriov_bar0_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar1_mask_reg_pci_sriov_bar1_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar1_reg_sriov_vf_bar1_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar2_mask_reg_pci_sriov_bar2_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar3_mask_reg_pci_sriov_bar3_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar3_reg_sriov_vf_bar3_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar4_mask_reg_pci_sriov_bar4_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar5_mask_reg_pci_sriov_bar5_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar5_reg_sriov_vf_bar5_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_vf_offset_position_sriov_vf_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_vf_offset_position_sriov_vf_stride                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sup_page_sizes_reg_sriov_sup_page_size                              ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_int_vec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_size                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_device_spec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_vf_device_id_reg_sriov_vf_device_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf2_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_at_block                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_egress_control                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_src_valid                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_usp_forwarding                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ats_capabilities_ctrl_reg_invalidate_q_depth                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ats_capabilities_ctrl_reg_page_aligned_req                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_mask_reg_pci_type0_bar0_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_mask_reg_pci_type0_bar0_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_reg_bar0_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_reg_bar0_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar1_mask_reg_pci_type0_bar1_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar1_mask_reg_pci_type0_bar1_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar1_reg_bar1_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_mask_reg_pci_type0_bar2_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_mask_reg_pci_type0_bar2_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_reg_bar2_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_reg_bar2_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar3_mask_reg_pci_type0_bar3_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar3_mask_reg_pci_type0_bar3_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar3_reg_bar3_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_mask_reg_pci_type0_bar4_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_mask_reg_pci_type0_bar4_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_reg_bar4_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_reg_bar4_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar5_mask_reg_pci_type0_bar5_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar5_mask_reg_pci_type0_bar5_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar5_reg_bar5_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cap_id_nxt_ptr_reg_aux_curr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cap_id_nxt_ptr_reg_dsi                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cap_id_nxt_ptr_reg_pme_support                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cardbus_cis_ptr_reg_cardbus_cis_pointer                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_base_class_code                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_program_interface                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_revision_id                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_subclass_code                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_con_status_reg_no_soft_rst                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_capabilities_reg_pcie_cap_flr_cap                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_control_device_status_pcie_cap_ext_tag_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_id_vendor_id_reg_pci_type0_device_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_id_vendor_id_reg_pci_type0_vendor_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_bar_mask_reg_rom_bar_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_bar_mask_reg_rom_mask                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_base_addr_reg_exp_rom_base_address                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_base_addr_reg_exp_rom_base_address),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_base_addr_reg_rom_bar_enable                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_capabilities_reg_pcie_cap_l0s_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_capabilities_reg_pcie_cap_l1_exit_latency                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_capabilities_reg_pcie_cap_port_num                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_control2_link_status2_reg_pcie_cap_sel_deemphasis              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_control_link_status_reg_pcie_cap_active_state_link_pm_control  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_control_link_status_reg_pcie_cap_slot_clk_config               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_pba_offset_reg_pci_msix_pba_bir                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_pba_offset_reg_pci_msix_pba_offset                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_table_offset_reg_pci_msix_bir                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_table_offset_reg_pci_msix_table_offset                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pasid_cap_cntrl_reg_execute_permission_supported                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pasid_cap_cntrl_reg_max_pasid_width                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pasid_cap_cntrl_reg_privileged_mode_supported                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_device_spec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar0_mask_reg_pci_sriov_bar0_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar1_mask_reg_pci_sriov_bar1_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar1_reg_sriov_vf_bar1_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar2_mask_reg_pci_sriov_bar2_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar3_mask_reg_pci_sriov_bar3_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar3_reg_sriov_vf_bar3_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar4_mask_reg_pci_sriov_bar4_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar5_mask_reg_pci_sriov_bar5_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar5_reg_sriov_vf_bar5_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_vf_offset_position_sriov_vf_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_vf_offset_position_sriov_vf_stride                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sup_page_sizes_reg_sriov_sup_page_size                              ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_int_vec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_size                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_device_spec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_vf_device_id_reg_sriov_vf_device_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf3_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_at_block                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_egress_control                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_src_valid                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_usp_forwarding                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ats_capabilities_ctrl_reg_invalidate_q_depth                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ats_capabilities_ctrl_reg_page_aligned_req                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_mask_reg_pci_type0_bar0_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_mask_reg_pci_type0_bar0_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_reg_bar0_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_reg_bar0_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar1_mask_reg_pci_type0_bar1_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar1_mask_reg_pci_type0_bar1_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar1_reg_bar1_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_mask_reg_pci_type0_bar2_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_mask_reg_pci_type0_bar2_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_reg_bar2_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_reg_bar2_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar3_mask_reg_pci_type0_bar3_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar3_mask_reg_pci_type0_bar3_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar3_reg_bar3_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_mask_reg_pci_type0_bar4_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_mask_reg_pci_type0_bar4_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_reg_bar4_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_reg_bar4_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar5_mask_reg_pci_type0_bar5_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar5_mask_reg_pci_type0_bar5_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar5_reg_bar5_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cap_id_nxt_ptr_reg_aux_curr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cap_id_nxt_ptr_reg_dsi                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cap_id_nxt_ptr_reg_pme_support                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cardbus_cis_ptr_reg_cardbus_cis_pointer                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_base_class_code                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_program_interface                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_revision_id                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_subclass_code                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_con_status_reg_no_soft_rst                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_capabilities_reg_pcie_cap_flr_cap                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_control_device_status_pcie_cap_ext_tag_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_id_vendor_id_reg_pci_type0_device_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_id_vendor_id_reg_pci_type0_vendor_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_bar_mask_reg_rom_bar_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_bar_mask_reg_rom_mask                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_base_addr_reg_exp_rom_base_address                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_base_addr_reg_exp_rom_base_address),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_base_addr_reg_rom_bar_enable                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_capabilities_reg_pcie_cap_l0s_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_capabilities_reg_pcie_cap_l1_exit_latency                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_capabilities_reg_pcie_cap_port_num                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_control2_link_status2_reg_pcie_cap_sel_deemphasis              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_control_link_status_reg_pcie_cap_active_state_link_pm_control  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_control_link_status_reg_pcie_cap_slot_clk_config               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_pba_offset_reg_pci_msix_pba_bir                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_pba_offset_reg_pci_msix_pba_offset                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_table_offset_reg_pci_msix_bir                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_table_offset_reg_pci_msix_table_offset                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pasid_cap_cntrl_reg_execute_permission_supported                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pasid_cap_cntrl_reg_max_pasid_width                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pasid_cap_cntrl_reg_privileged_mode_supported                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_device_spec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar0_mask_reg_pci_sriov_bar0_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar1_mask_reg_pci_sriov_bar1_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar1_reg_sriov_vf_bar1_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar2_mask_reg_pci_sriov_bar2_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar3_mask_reg_pci_sriov_bar3_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar3_reg_sriov_vf_bar3_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar4_mask_reg_pci_sriov_bar4_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar5_mask_reg_pci_sriov_bar5_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar5_reg_sriov_vf_bar5_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_vf_offset_position_sriov_vf_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_vf_offset_position_sriov_vf_stride                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sup_page_sizes_reg_sriov_sup_page_size                              ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_int_vec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_size                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_device_spec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_vf_device_id_reg_sriov_vf_device_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf4_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_at_block                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_egress_control                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_src_valid                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_usp_forwarding                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ats_capabilities_ctrl_reg_invalidate_q_depth                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ats_capabilities_ctrl_reg_page_aligned_req                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_mask_reg_pci_type0_bar0_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_mask_reg_pci_type0_bar0_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_reg_bar0_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_reg_bar0_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar1_mask_reg_pci_type0_bar1_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar1_mask_reg_pci_type0_bar1_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar1_reg_bar1_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_mask_reg_pci_type0_bar2_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_mask_reg_pci_type0_bar2_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_reg_bar2_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_reg_bar2_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar3_mask_reg_pci_type0_bar3_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar3_mask_reg_pci_type0_bar3_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar3_reg_bar3_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_mask_reg_pci_type0_bar4_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_mask_reg_pci_type0_bar4_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_reg_bar4_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_reg_bar4_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar5_mask_reg_pci_type0_bar5_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar5_mask_reg_pci_type0_bar5_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar5_reg_bar5_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cap_id_nxt_ptr_reg_aux_curr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cap_id_nxt_ptr_reg_dsi                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cap_id_nxt_ptr_reg_pme_support                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cardbus_cis_ptr_reg_cardbus_cis_pointer                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_base_class_code                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_program_interface                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_revision_id                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_subclass_code                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_con_status_reg_no_soft_rst                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_capabilities_reg_pcie_cap_flr_cap                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_control_device_status_pcie_cap_ext_tag_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_id_vendor_id_reg_pci_type0_device_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_id_vendor_id_reg_pci_type0_vendor_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_bar_mask_reg_rom_bar_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_bar_mask_reg_rom_mask                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_base_addr_reg_exp_rom_base_address                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_base_addr_reg_exp_rom_base_address),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_base_addr_reg_rom_bar_enable                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_capabilities_reg_pcie_cap_l0s_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_capabilities_reg_pcie_cap_l1_exit_latency                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_capabilities_reg_pcie_cap_port_num                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_control2_link_status2_reg_pcie_cap_sel_deemphasis              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_control_link_status_reg_pcie_cap_active_state_link_pm_control  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_control_link_status_reg_pcie_cap_slot_clk_config               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_pba_offset_reg_pci_msix_pba_bir                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_pba_offset_reg_pci_msix_pba_offset                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_table_offset_reg_pci_msix_bir                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_table_offset_reg_pci_msix_table_offset                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pasid_cap_cntrl_reg_execute_permission_supported                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pasid_cap_cntrl_reg_max_pasid_width                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pasid_cap_cntrl_reg_privileged_mode_supported                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_device_spec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar0_mask_reg_pci_sriov_bar0_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar1_mask_reg_pci_sriov_bar1_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar1_reg_sriov_vf_bar1_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar2_mask_reg_pci_sriov_bar2_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar3_mask_reg_pci_sriov_bar3_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar3_reg_sriov_vf_bar3_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar4_mask_reg_pci_sriov_bar4_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar5_mask_reg_pci_sriov_bar5_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar5_reg_sriov_vf_bar5_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_vf_offset_position_sriov_vf_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_vf_offset_position_sriov_vf_stride                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sup_page_sizes_reg_sriov_sup_page_size                              ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_int_vec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_size                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_device_spec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_vf_device_id_reg_sriov_vf_device_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf5_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_at_block                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_egress_control                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_src_valid                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_usp_forwarding                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ats_capabilities_ctrl_reg_invalidate_q_depth                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ats_capabilities_ctrl_reg_page_aligned_req                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_mask_reg_pci_type0_bar0_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_mask_reg_pci_type0_bar0_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_reg_bar0_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_reg_bar0_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar1_mask_reg_pci_type0_bar1_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar1_mask_reg_pci_type0_bar1_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar1_reg_bar1_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_mask_reg_pci_type0_bar2_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_mask_reg_pci_type0_bar2_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_reg_bar2_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_reg_bar2_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar3_mask_reg_pci_type0_bar3_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar3_mask_reg_pci_type0_bar3_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar3_reg_bar3_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_mask_reg_pci_type0_bar4_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_mask_reg_pci_type0_bar4_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_reg_bar4_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_reg_bar4_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar5_mask_reg_pci_type0_bar5_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar5_mask_reg_pci_type0_bar5_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar5_reg_bar5_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cap_id_nxt_ptr_reg_aux_curr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cap_id_nxt_ptr_reg_dsi                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cap_id_nxt_ptr_reg_pme_support                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cardbus_cis_ptr_reg_cardbus_cis_pointer                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_base_class_code                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_program_interface                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_revision_id                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_subclass_code                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_con_status_reg_no_soft_rst                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_capabilities_reg_pcie_cap_flr_cap                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_control_device_status_pcie_cap_ext_tag_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_id_vendor_id_reg_pci_type0_device_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_id_vendor_id_reg_pci_type0_vendor_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_bar_mask_reg_rom_bar_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_bar_mask_reg_rom_mask                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_base_addr_reg_exp_rom_base_address                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_base_addr_reg_exp_rom_base_address),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_base_addr_reg_rom_bar_enable                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_capabilities_reg_pcie_cap_l0s_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_capabilities_reg_pcie_cap_l1_exit_latency                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_capabilities_reg_pcie_cap_port_num                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_control2_link_status2_reg_pcie_cap_sel_deemphasis              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_control_link_status_reg_pcie_cap_active_state_link_pm_control  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_control_link_status_reg_pcie_cap_slot_clk_config               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_pba_offset_reg_pci_msix_pba_bir                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_pba_offset_reg_pci_msix_pba_offset                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_table_offset_reg_pci_msix_bir                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_table_offset_reg_pci_msix_table_offset                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pasid_cap_cntrl_reg_execute_permission_supported                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pasid_cap_cntrl_reg_max_pasid_width                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pasid_cap_cntrl_reg_privileged_mode_supported                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_device_spec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar0_mask_reg_pci_sriov_bar0_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar1_mask_reg_pci_sriov_bar1_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar1_reg_sriov_vf_bar1_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar2_mask_reg_pci_sriov_bar2_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar3_mask_reg_pci_sriov_bar3_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar3_reg_sriov_vf_bar3_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar4_mask_reg_pci_sriov_bar4_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar5_mask_reg_pci_sriov_bar5_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar5_reg_sriov_vf_bar5_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_vf_offset_position_sriov_vf_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_vf_offset_position_sriov_vf_stride                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sup_page_sizes_reg_sriov_sup_page_size                              ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_int_vec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_size                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_device_spec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_vf_device_id_reg_sriov_vf_device_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf6_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_at_block                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_egress_control                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_src_valid                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_usp_forwarding                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ats_capabilities_ctrl_reg_invalidate_q_depth                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ats_capabilities_ctrl_reg_page_aligned_req                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_mask_reg_pci_type0_bar0_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_mask_reg_pci_type0_bar0_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_reg_bar0_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_reg_bar0_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar1_mask_reg_pci_type0_bar1_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar1_mask_reg_pci_type0_bar1_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar1_reg_bar1_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_mask_reg_pci_type0_bar2_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_mask_reg_pci_type0_bar2_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_reg_bar2_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_reg_bar2_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar3_mask_reg_pci_type0_bar3_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar3_mask_reg_pci_type0_bar3_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar3_reg_bar3_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_mask_reg_pci_type0_bar4_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_mask_reg_pci_type0_bar4_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_reg_bar4_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_reg_bar4_type                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar5_mask_reg_pci_type0_bar5_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar5_mask_reg_pci_type0_bar5_mask                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar5_reg_bar5_prefetch                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cap_id_nxt_ptr_reg_aux_curr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cap_id_nxt_ptr_reg_dsi                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cap_id_nxt_ptr_reg_pme_support                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cardbus_cis_ptr_reg_cardbus_cis_pointer                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_base_class_code                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_program_interface                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_revision_id                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_subclass_code                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_con_status_reg_no_soft_rst                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_capabilities_reg_pcie_cap_flr_cap                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_control_device_status_pcie_cap_ext_tag_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_id_vendor_id_reg_pci_type0_device_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_id_vendor_id_reg_pci_type0_vendor_id                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_bar_mask_reg_rom_bar_enabled                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_bar_mask_reg_rom_mask                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_base_addr_reg_exp_rom_base_address                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_base_addr_reg_exp_rom_base_address),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_base_addr_reg_rom_bar_enable                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_capabilities_reg_pcie_cap_l0s_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_capabilities_reg_pcie_cap_l1_exit_latency                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_capabilities_reg_pcie_cap_port_num                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_control2_link_status2_reg_pcie_cap_sel_deemphasis              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_control_link_status_reg_pcie_cap_active_state_link_pm_control  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_control_link_status_reg_pcie_cap_slot_clk_config               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_pba_offset_reg_pci_msix_pba_bir                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_pba_offset_reg_pci_msix_pba_offset                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_table_offset_reg_pci_msix_bir                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_table_offset_reg_pci_msix_table_offset                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pasid_cap_cntrl_reg_execute_permission_supported                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pasid_cap_cntrl_reg_max_pasid_width                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pasid_cap_cntrl_reg_privileged_mode_supported                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_device_spec                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar0_mask_reg_pci_sriov_bar0_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar1_mask_reg_pci_sriov_bar1_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar1_reg_sriov_vf_bar1_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar2_mask_reg_pci_sriov_bar2_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar3_mask_reg_pci_sriov_bar3_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar3_reg_sriov_vf_bar3_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar4_mask_reg_pci_sriov_bar4_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_type                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar5_mask_reg_pci_sriov_bar5_mask                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar5_reg_sriov_vf_bar5_prefetch                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_vf_offset_position_sriov_vf_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_vf_offset_position_sriov_vf_stride                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sup_page_sizes_reg_sriov_sup_page_size                              ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_int_vec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_size                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_device_spec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_vf_device_id_reg_sriov_vf_device_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pf7_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pfvf_sel_vsec_enable_attr                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_pfvf_sel_vsec_enable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_phy_rxelecidle_k_rxelecidle_disable_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_phy_rxelecidle_k_rxelecidle_disable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_phy_rxtermination_k_rxtermination_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_phy_rxtermination_k_rxtermination_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ptm_ctrl_k_cfg_ptm_auto_update_signal_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ptm_ctrl_k_cfg_ptm_auto_update_signal_attr),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ptm_adj_lsb_k_cfg_ptm_local_clock_adj_lsb_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ptm_adj_lsb_k_cfg_ptm_local_clock_adj_lsb_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ptm_adj_msb_k_cfg_ptm_local_clock_adj_msb_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_ptm_adj_msb_k_cfg_ptm_local_clock_adj_msb_attr),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_reset_ctrl0_k_cvp_intf_reset_ctl_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_reset_ctrl0_k_cvp_intf_reset_ctl_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_err_en_correct_err_en_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_err_en_correct_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_err_en_fatal_err_en_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_err_en_fatal_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_err_en_nonfatal_err_en_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_err_en_nonfatal_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_bw_mgt_int_en_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_bw_mgt_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_link_eq_req_int_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_link_eq_req_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_pme_int_en_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_cfg_pme_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_hp_int_en_attr                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_hp_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_hp_pme_en_attr                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_hp_pme_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_inta_en_attr                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_inta_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_intb_en_attr                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_intb_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_intc_en_attr                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_intc_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_intd_en_attr                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_rp_irq_en_intd_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_sriov_misc_ctrl_k_nonsriov_mode_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_sriov_misc_ctrl_k_nonsriov_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_stagger_control_k_stag_dlycnt_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_stagger_control_k_stag_dlycnt_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_stagger_control_k_stag_mode_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_stagger_control_k_stag_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id0_k_exvf_subsysid_pf0_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id0_k_exvf_subsysid_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id0_k_exvf_subsysid_pf1_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id0_k_exvf_subsysid_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id1_k_exvf_subsysid_pf2_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id1_k_exvf_subsysid_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id1_k_exvf_subsysid_pf3_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id1_k_exvf_subsysid_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id2_k_exvf_subsysid_pf4_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id2_k_exvf_subsysid_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id2_k_exvf_subsysid_pf5_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id2_k_exvf_subsysid_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id3_k_exvf_subsysid_pf6_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id3_k_exvf_subsysid_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id3_k_exvf_subsysid_pf7_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_subs_id3_k_exvf_subsysid_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf0_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf1_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablesize_pf0_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablesize_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablesize_pf1_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl0_k_exvf_tph_sttablesize_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf2_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf3_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablesize_pf2_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablesize_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablesize_pf3_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl1_k_exvf_tph_sttablesize_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf4_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf5_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablesize_pf4_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablesize_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablesize_pf5_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl2_k_exvf_tph_sttablesize_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf6_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf7_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablesize_pf6_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablesize_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablesize_pf7_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tph_ctl3_k_exvf_tph_sttablesize_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tx_common_mode_k_txcommonmode_disable_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_tx_common_mode_k_txcommonmode_disable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_100_k_pf4_virtio_offset_cfg3_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_100_k_pf4_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_102_k_pf4_virtio_offset_cfg4_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_102_k_pf4_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_103_k_pf4_virtio_offset_cfg4_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_103_k_pf4_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_104_k_pf4_virtio_offset_cfg4_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_104_k_pf4_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_106_k_pf4_virtio_offset_cfg5_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_106_k_pf4_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_107_k_pf4_virtio_offset_cfg5_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_107_k_pf4_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_108_k_pf4_virtio_offset_cfg5_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_108_k_pf4_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_109_k_pf4_virtio_offset_cfg5_cfg_data_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_109_k_pf4_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_111_k_pf5_virtio_offset_cfg1_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_111_k_pf5_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_112_k_pf5_virtio_offset_cfg1_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_112_k_pf5_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_113_k_pf5_virtio_offset_cfg1_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_113_k_pf5_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_115_k_pf5_virtio_offset_cfg2_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_115_k_pf5_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_116_k_pf5_virtio_offset_cfg2_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_116_k_pf5_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_117_k_pf5_virtio_offset_cfg2_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_117_k_pf5_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_118_k_pf5_virtio_offset_cfg2_notify_off_multiplier_attr          ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_118_k_pf5_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_120_k_pf5_virtio_offset_cfg3_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_120_k_pf5_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_121_k_pf5_virtio_offset_cfg3_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_121_k_pf5_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_122_k_pf5_virtio_offset_cfg3_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_122_k_pf5_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_124_k_pf5_virtio_offset_cfg4_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_124_k_pf5_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_125_k_pf5_virtio_offset_cfg4_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_125_k_pf5_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_126_k_pf5_virtio_offset_cfg4_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_126_k_pf5_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_128_k_pf5_virtio_offset_cfg5_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_128_k_pf5_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_129_k_pf5_virtio_offset_cfg5_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_129_k_pf5_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_130_k_pf5_virtio_offset_cfg5_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_130_k_pf5_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_131_k_pf5_virtio_offset_cfg5_cfg_data_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_131_k_pf5_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_133_k_pf6_virtio_offset_cfg1_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_133_k_pf6_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_134_k_pf6_virtio_offset_cfg1_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_134_k_pf6_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_135_k_pf6_virtio_offset_cfg1_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_135_k_pf6_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_137_k_pf6_virtio_offset_cfg2_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_137_k_pf6_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_138_k_pf6_virtio_offset_cfg2_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_138_k_pf6_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_139_k_pf6_virtio_offset_cfg2_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_139_k_pf6_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_140_k_pf6_virtio_offset_cfg2_notify_off_multiplier_attr          ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_140_k_pf6_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_142_k_pf6_virtio_offset_cfg3_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_142_k_pf6_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_143_k_pf6_virtio_offset_cfg3_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_143_k_pf6_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_144_k_pf6_virtio_offset_cfg3_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_144_k_pf6_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_146_k_pf6_virtio_offset_cfg4_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_146_k_pf6_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_147_k_pf6_virtio_offset_cfg4_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_147_k_pf6_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_148_k_pf6_virtio_offset_cfg4_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_148_k_pf6_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_150_k_pf6_virtio_offset_cfg5_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_150_k_pf6_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_151_k_pf6_virtio_offset_cfg5_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_151_k_pf6_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_152_k_pf6_virtio_offset_cfg5_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_152_k_pf6_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_153_k_pf6_virtio_offset_cfg5_cfg_data_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_153_k_pf6_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_155_k_pf7_virtio_offset_cfg1_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_155_k_pf7_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_156_k_pf7_virtio_offset_cfg1_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_156_k_pf7_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_157_k_pf7_virtio_offset_cfg1_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_157_k_pf7_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_159_k_pf7_virtio_offset_cfg2_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_159_k_pf7_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_160_k_pf7_virtio_offset_cfg2_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_160_k_pf7_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_161_k_pf7_virtio_offset_cfg2_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_161_k_pf7_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_162_k_pf7_virtio_offset_cfg2_notify_off_multiplier_attr          ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_162_k_pf7_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_164_k_pf7_virtio_offset_cfg3_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_164_k_pf7_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_165_k_pf7_virtio_offset_cfg3_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_165_k_pf7_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_166_k_pf7_virtio_offset_cfg3_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_166_k_pf7_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_168_k_pf7_virtio_offset_cfg4_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_168_k_pf7_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_169_k_pf7_virtio_offset_cfg4_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_169_k_pf7_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_170_k_pf7_virtio_offset_cfg4_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_170_k_pf7_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_172_k_pf7_virtio_offset_cfg5_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_172_k_pf7_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_173_k_pf7_virtio_offset_cfg5_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_173_k_pf7_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_174_k_pf7_virtio_offset_cfg5_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_174_k_pf7_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_175_k_pf7_virtio_offset_cfg5_cfg_data_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_175_k_pf7_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_23_k_pf1_virtio_offset_cfg1_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_23_k_pf1_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_24_k_pf1_virtio_offset_cfg1_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_24_k_pf1_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_25_k_pf1_virtio_offset_cfg1_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_25_k_pf1_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_27_k_pf1_virtio_offset_cfg2_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_27_k_pf1_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_28_k_pf1_virtio_offset_cfg2_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_28_k_pf1_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_29_k_pf1_virtio_offset_cfg2_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_29_k_pf1_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_30_k_pf1_virtio_offset_cfg2_notify_off_multiplier_attr           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_30_k_pf1_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_32_k_pf1_virtio_offset_cfg3_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_32_k_pf1_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_33_k_pf1_virtio_offset_cfg3_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_33_k_pf1_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_34_k_pf1_virtio_offset_cfg3_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_34_k_pf1_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_36_k_pf1_virtio_offset_cfg4_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_36_k_pf1_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_37_k_pf1_virtio_offset_cfg4_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_37_k_pf1_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_38_k_pf1_virtio_offset_cfg4_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_38_k_pf1_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_40_k_pf1_virtio_offset_cfg5_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_40_k_pf1_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_41_k_pf1_virtio_offset_cfg5_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_41_k_pf1_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_42_k_pf1_virtio_offset_cfg5_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_42_k_pf1_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_43_k_pf1_virtio_offset_cfg5_cfg_data_attr                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_43_k_pf1_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_45_k_pf2_virtio_offset_cfg1_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_45_k_pf2_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_46_k_pf2_virtio_offset_cfg1_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_46_k_pf2_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_47_k_pf2_virtio_offset_cfg1_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_47_k_pf2_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_49_k_pf2_virtio_offset_cfg2_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_49_k_pf2_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_50_k_pf2_virtio_offset_cfg2_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_50_k_pf2_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_51_k_pf2_virtio_offset_cfg2_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_51_k_pf2_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_52_k_pf2_virtio_offset_cfg2_notify_off_multiplier_attr           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_52_k_pf2_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_54_k_pf2_virtio_offset_cfg3_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_54_k_pf2_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_55_k_pf2_virtio_offset_cfg3_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_55_k_pf2_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_56_k_pf2_virtio_offset_cfg3_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_56_k_pf2_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_58_k_pf2_virtio_offset_cfg4_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_58_k_pf2_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_59_k_pf2_virtio_offset_cfg4_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_59_k_pf2_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_60_k_pf2_virtio_offset_cfg4_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_60_k_pf2_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_62_k_pf2_virtio_offset_cfg5_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_62_k_pf2_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_63_k_pf2_virtio_offset_cfg5_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_63_k_pf2_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_64_k_pf2_virtio_offset_cfg5_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_64_k_pf2_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_65_k_pf2_virtio_offset_cfg5_cfg_data_attr                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_65_k_pf2_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_67_k_pf3_virtio_offset_cfg1_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_67_k_pf3_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_68_k_pf3_virtio_offset_cfg1_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_68_k_pf3_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_69_k_pf3_virtio_offset_cfg1_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_69_k_pf3_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_71_k_pf3_virtio_offset_cfg2_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_71_k_pf3_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_72_k_pf3_virtio_offset_cfg2_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_72_k_pf3_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_73_k_pf3_virtio_offset_cfg2_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_73_k_pf3_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_74_k_pf3_virtio_offset_cfg2_notify_off_multiplier_attr           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_74_k_pf3_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_76_k_pf3_virtio_offset_cfg3_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_76_k_pf3_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_77_k_pf3_virtio_offset_cfg3_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_77_k_pf3_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_78_k_pf3_virtio_offset_cfg3_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_78_k_pf3_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_80_k_pf3_virtio_offset_cfg4_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_80_k_pf3_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_81_k_pf3_virtio_offset_cfg4_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_81_k_pf3_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_82_k_pf3_virtio_offset_cfg4_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_82_k_pf3_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_84_k_pf3_virtio_offset_cfg5_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_84_k_pf3_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_85_k_pf3_virtio_offset_cfg5_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_85_k_pf3_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_86_k_pf3_virtio_offset_cfg5_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_86_k_pf3_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_87_k_pf3_virtio_offset_cfg5_cfg_data_attr                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_87_k_pf3_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_89_k_pf4_virtio_offset_cfg1_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_89_k_pf4_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_90_k_pf4_virtio_offset_cfg1_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_90_k_pf4_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_91_k_pf4_virtio_offset_cfg1_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_91_k_pf4_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_93_k_pf4_virtio_offset_cfg2_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_93_k_pf4_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_94_k_pf4_virtio_offset_cfg2_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_94_k_pf4_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_95_k_pf4_virtio_offset_cfg2_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_95_k_pf4_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_96_k_pf4_virtio_offset_cfg2_notify_off_multiplier_attr           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_96_k_pf4_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_98_k_pf4_virtio_offset_cfg3_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_98_k_pf4_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_99_k_pf4_virtio_offset_cfg3_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_99_k_pf4_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_cii_ctrl_k_cfg_update_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_cii_ctrl_k_cfg_update_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_cii_ctrl_k_cii_en_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_cii_ctrl_k_cii_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_cvp_mode                                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_cvp_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_drop_vendor0_msg                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_drop_vendor0_msg),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_drop_vendor1_msg                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_drop_vendor1_msg),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_ep_native                                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_ep_native),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_maxpayload_size                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_maxpayload_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_num_of_lanes                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_num_of_lanes),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_acs_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_ats_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_bar1_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_bar3_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_bar5_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_dlink_cap_enable                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_dlink_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_acs_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_ats_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_msix_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_tph_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_virtio_en                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_io_decode                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_io_decode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_ltr_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_ltr_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_msi_enable                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_msix_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_pasid_cap_enable                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_prefetch_decode                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_prefetch_decode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_prs_ext_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_ras_des_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sn_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_num_vf_non_ari                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar0_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar1_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar2_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar3_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar4_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar5_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_tph_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_user_vsec_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_virtio_dev_specific_conf_en                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_virtio_en                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_vsecras_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf0_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_acs_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_ats_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_bar1_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_bar3_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_bar5_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_enable                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_acs_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_ats_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_msix_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_tph_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_virtio_en                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_msi_enable                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_msix_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_pasid_cap_enable                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_prs_ext_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_ras_des_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sn_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_num_vf_non_ari                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar0_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar1_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar2_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar3_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar4_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar5_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_tph_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_user_vsec_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_user_vsec_offset                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_virtio_dev_specific_conf_en                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_virtio_en                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_vsecras_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf1_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_acs_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_ats_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_bar1_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_bar3_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_bar5_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_enable                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_acs_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_ats_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_msix_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_tph_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_virtio_en                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_msi_enable                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_msix_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_pasid_cap_enable                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_prs_ext_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_ras_des_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sn_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_num_vf_non_ari                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar0_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar1_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar2_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar3_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar4_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar5_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_tph_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_user_vsec_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_user_vsec_offset                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_virtio_dev_specific_conf_en                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_virtio_en                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_vsecras_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf2_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_acs_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_ats_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_bar1_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_bar3_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_bar5_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_enable                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_acs_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_ats_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_msix_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_tph_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_virtio_en                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_msi_enable                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_msix_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_pasid_cap_enable                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_prs_ext_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_ras_des_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sn_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_num_vf_non_ari                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar0_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar1_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar2_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar3_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar4_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar5_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_tph_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_user_vsec_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_user_vsec_offset                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_virtio_dev_specific_conf_en                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_virtio_en                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_vsecras_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf3_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_acs_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_ats_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_bar1_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_bar3_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_bar5_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_enable                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_acs_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_ats_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_msix_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_tph_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_virtio_en                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_msi_enable                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_msix_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_pasid_cap_enable                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_prs_ext_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_ras_des_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sn_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_num_vf_non_ari                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar0_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar1_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar2_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar3_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar4_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar5_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_tph_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_user_vsec_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_user_vsec_offset                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_virtio_dev_specific_conf_en                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_virtio_en                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_vsecras_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf4_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_acs_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_ats_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_bar1_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_bar3_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_bar5_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_enable                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_acs_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_ats_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_msix_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_tph_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_virtio_en                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_msi_enable                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_msix_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_pasid_cap_enable                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_prs_ext_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_ras_des_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sn_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_num_vf_non_ari                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar0_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar1_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar2_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar3_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar4_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar5_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_tph_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_user_vsec_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_user_vsec_offset                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_virtio_dev_specific_conf_en                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_virtio_en                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_vsecras_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf5_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_acs_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_ats_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_bar1_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_bar3_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_bar5_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_enable                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_acs_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_ats_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_msix_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_tph_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_virtio_en                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_msi_enable                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_msix_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_pasid_cap_enable                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_prs_ext_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_ras_des_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sn_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_num_vf_non_ari                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar0_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar1_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar2_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar3_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar4_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar5_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_tph_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_user_vsec_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_user_vsec_offset                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_virtio_dev_specific_conf_en                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_virtio_en                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_vsecras_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf6_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_acs_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_ats_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_bar1_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_bar3_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_bar5_mask_bit0                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_enable                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_acs_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_ats_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_msix_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_tph_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_virtio_en                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_msi_enable                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_msix_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_pasid_cap_enable                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_prs_ext_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_ras_des_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sn_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_num_vf_non_ari                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar0_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar1_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar2_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar3_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar4_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar5_enabled                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_tph_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_user_vsec_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_user_vsec_offset                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_virtio_dev_specific_conf_en                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_virtio_en                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_vsecras_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_pf7_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_ptm_autoupdate                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_ptm_autoupdate),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p0_inst_rnr_pcie_ip16_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_addr_size0_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_addr_size0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_pf_en0_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_pf_en0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_start_addr0_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_start_addr0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_addr_size1_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_addr_size1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_pf_en1_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_pf_en1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_start_addr1_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_start_addr1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_addr_size2_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_addr_size2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_pf_en2_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_pf_en2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_start_addr2_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_start_addr2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_addr_size3_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_addr_size3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_pf_en3_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_pf_en3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_start_addr3_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_start_addr3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_addr_size4_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_addr_size4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_pf_en4_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_pf_en4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_start_addr4_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_start_addr4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_addr_size5_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_addr_size5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_pf_en5_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_pf_en5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_start_addr5_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_start_addr5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_addr_size6_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_addr_size6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_pf_en6_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_pf_en6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_start_addr6_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_start_addr6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_addr_size7_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_addr_size7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_pf_en7_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_pf_en7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_start_addr7_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_start_addr7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_fixedcred_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_fixedcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_mcred_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_mcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_reloadcred_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_reloadcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_tlp_serr_dis_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_tlp_serr_dis_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_mmio_access_ctrl_grant_attr                                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_mmio_access_ctrl_grant_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_opcode_ctrl_lock_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_csb_opcode_ctrl_lock_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_compressed_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_compressed_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_encrypted_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_encrypted_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_devbrd_type_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_devbrd_type_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_vsec_next_offset_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_vsec_next_offset_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_cvp_irq_en_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_cvp_irq_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_gpio_irq_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_gpio_irq_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid0_k_jtag_id_0_attr                                           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid0_k_jtag_id_0_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid1_k_jtag_id_1_attr                                           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid1_k_jtag_id_1_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid2_k_jtag_id_2_attr                                           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid2_k_jtag_id_2_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid3_k_jtag_id_3_attr                                           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_cvp_jtagid3_k_jtag_id_3_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_dfd_en_attr                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_dfd_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_patcntr_en_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_patcntr_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_0_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_1_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_2_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_3_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_data_sel_3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_trig_sel_0_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_trig_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_trig_sel_1_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_trig_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_0_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_1_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_2_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_3_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_crs_en_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_crs_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_rx_lane_flip_en_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_rx_lane_flip_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_sris_mode_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_sris_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_tx_lane_flip_en_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_tx_lane_flip_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_ehp_ctrl0_k_ehp_control_reg_attr                                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_ehp_ctrl0_k_ehp_control_reg_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_outstanding_crd_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_outstanding_crd_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_tx_rd_th_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_tx_rd_th_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cvp_cfg_err_en_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cvp_cfg_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dbi_access_err_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dbi_access_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_multi_lane_control_off_upconfigure_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_multi_lane_control_off_upconfigure_support),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar1_reg_bar1_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_mem_io                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_mem_io),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar5_reg_bar5_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bist_header_type_latency_cache_line_size_reg_multi_func            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_bist_header_type_latency_cache_line_size_reg_multi_func),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_aux_curr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_dsi                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_pme_support                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_reg_ari_acs_fun_grp_cap                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_cap_reg_ari_acs_fun_grp_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_base_class_code                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_program_interface                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_revision_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_subclass_code                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_con_status_reg_no_soft_rst                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ext_tag_supp                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ext_tag_supp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_mask                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_config_phy_tx_change                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_config_phy_tx_change),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_select_deemph_var_mux                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_select_deemph_var_mux),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_selectable_deemph_bit_mux                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_selectable_deemph_bit_mux),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_support_mod_ts                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_support_mod_ts),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg4                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg5                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg4                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg5                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_l1_2                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_l1_2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_power_off                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_power_off),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_comm_mode_support                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_comm_mode_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_scale_support                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_scale_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_value_support                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_value_support),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_aspm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_aspm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_aspm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_aspm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_aspm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_aspm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_aspm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_aspm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_1sub_cap_enable ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_1sub_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_2sub_cap_enable ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_2sub_cap_enable),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_sca                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_sca),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_val                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_val),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_t_common_mode                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_t_common_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_port_num                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_misc_control_1_off_port_logic_wr_disable                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_misc_control_1_off_port_logic_wr_disable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_bir                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_table_offset                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pipe_loopback_control_off_pipe_loopback                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pipe_loopback_control_off_pipe_loopback),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_capability_reg_no_eq_needed_support                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_capability_reg_no_eq_needed_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rsvdp_11                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rsvdp_11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precode_req                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precode_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precoding_on                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precoding_on),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_port_force_off_support_part_lanes_rxei_exit                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_port_force_off_support_part_lanes_rxei_exit),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_port_link_ctrl_off_fast_link_mode                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_port_link_ctrl_off_fast_link_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_device_spec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pfvf_sel_vsec_enable_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_pfvf_sel_vsec_enable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_phy_rxelecidle_k_rxelecidle_disable_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_phy_rxelecidle_k_rxelecidle_disable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_phy_rxtermination_k_rxtermination_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_phy_rxtermination_k_rxtermination_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_err_en_correct_err_en_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_err_en_correct_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_err_en_fatal_err_en_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_err_en_fatal_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_err_en_nonfatal_err_en_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_err_en_nonfatal_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_bw_mgt_int_en_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_bw_mgt_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_eq_req_int_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_eq_req_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_pme_int_en_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_pme_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_int_en_attr                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_pme_en_attr                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_pme_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_inta_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_inta_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_intb_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_intb_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_intc_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_intc_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_intd_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_rp_irq_en_intd_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_dlycnt_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_dlycnt_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_mode_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_dllp_err_sts_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_dllp_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_tlp_err_sts_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_tlp_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_corrected_internal_err_sts_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_corrected_internal_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_dl_protocol_err_sts_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_dl_protocol_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_ecrc_err_sts_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_ecrc_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_fc_protocol_err_sts_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_fc_protocol_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_mlf_tlp_err_sts_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_mlf_tlp_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_err_sts_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_overflow_err_sts_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_overflow_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_number_rollover_err_sts_attr                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_number_rollover_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_timer_timeout_err_sts_attr                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_timer_timeout_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_surprise_down_err_sts_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_surprise_down_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_uncor_internal_err_sts_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_uncor_internal_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tx_common_mode_k_txcommonmode_disable_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_tx_common_mode_k_txcommonmode_disable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cfg_update_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cfg_update_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cii_en_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cii_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_cvp_mode                                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_cvp_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_drop_vendor0_msg                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_drop_vendor0_msg),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_drop_vendor1_msg                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_drop_vendor1_msg),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_ep_native                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_ep_native),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_maxpayload_size                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_maxpayload_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_num_of_lanes                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_num_of_lanes),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_acs_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_ats_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_bar1_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_bar3_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_bar5_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_dlink_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_dlink_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_acs_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_ats_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_msix_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_tph_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_io_decode                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_io_decode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_ltr_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_ltr_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_msi_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_msix_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_pasid_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_prefetch_decode                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_prefetch_decode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_prs_ext_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_ras_des_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_sn_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_tph_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_user_vsec_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_dev_specific_conf_en                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_en                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_vsecras_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_pf0_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_ptm_autoupdate                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_ptm_autoupdate),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip4_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr),
   
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf0_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf1_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf2_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf3_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl0_k_exvf_ats_pagealignreq_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf4_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf5_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf6_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf7_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ats_ctl1_k_exvf_ats_pagealignreq_pf7_attr),
   
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_0_k_cii_addr_size0_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_0_k_cii_addr_size0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_0_k_cii_pf_en0_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_0_k_cii_pf_en0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_0_k_cii_start_addr0_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_0_k_cii_start_addr0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_1_k_cii_addr_size1_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_1_k_cii_addr_size1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_1_k_cii_pf_en1_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_1_k_cii_pf_en1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_1_k_cii_start_addr1_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_1_k_cii_start_addr1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_2_k_cii_addr_size2_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_2_k_cii_addr_size2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_2_k_cii_pf_en2_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_2_k_cii_pf_en2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_2_k_cii_start_addr2_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_2_k_cii_start_addr2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_3_k_cii_addr_size3_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_3_k_cii_addr_size3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_3_k_cii_pf_en3_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_3_k_cii_pf_en3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_3_k_cii_start_addr3_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_3_k_cii_start_addr3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_4_k_cii_addr_size4_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_4_k_cii_addr_size4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_4_k_cii_pf_en4_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_4_k_cii_pf_en4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_4_k_cii_start_addr4_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_4_k_cii_start_addr4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_5_k_cii_addr_size5_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_5_k_cii_addr_size5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_5_k_cii_pf_en5_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_5_k_cii_pf_en5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_5_k_cii_start_addr5_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_5_k_cii_start_addr5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_6_k_cii_addr_size6_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_6_k_cii_addr_size6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_6_k_cii_pf_en6_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_6_k_cii_pf_en6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_6_k_cii_start_addr6_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_6_k_cii_start_addr6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_7_k_cii_addr_size7_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_7_k_cii_addr_size7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_7_k_cii_pf_en7_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_7_k_cii_pf_en7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_7_k_cii_start_addr7_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cii_range_7_k_cii_start_addr7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_fixedcred_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_fixedcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_mcred_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_mcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_reloadcred_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_reloadcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_tlp_serr_dis_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_ctrl0_k_tlp_serr_dis_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_mmio_access_ctrl_grant_attr                                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_mmio_access_ctrl_grant_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_opcode_ctrl_lock_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_csb_opcode_ctrl_lock_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl0_k_compressed_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl0_k_compressed_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl0_k_encrypted_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl0_k_encrypted_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl1_k_devbrd_type_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl1_k_devbrd_type_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl1_k_vsec_next_offset_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_ctrl1_k_vsec_next_offset_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_irq_ctrl_k_cvp_irq_en_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_irq_ctrl_k_cvp_irq_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_irq_ctrl_k_gpio_irq_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_irq_ctrl_k_gpio_irq_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid0_k_jtag_id_0_attr                                           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid0_k_jtag_id_0_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid1_k_jtag_id_1_attr                                           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid1_k_jtag_id_1_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid2_k_jtag_id_2_attr                                           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid2_k_jtag_id_2_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid3_k_jtag_id_3_attr                                           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_cvp_jtagid3_k_jtag_id_3_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_ctrl0_k_dfd_en_attr                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_ctrl0_k_dfd_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_ctrl0_k_patcntr_en_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_ctrl0_k_patcntr_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_0_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_1_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_2_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_3_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_data_sel_3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_trig_sel_0_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_trig_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_trig_sel_1_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_trig_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_0_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_1_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_2_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_3_attr                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dfd_xbar_sel_3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_pld_crs_en_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_pld_crs_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_rx_lane_flip_en_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_rx_lane_flip_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_sris_mode_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_sris_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_tx_lane_flip_en_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_dwc_ctrl0_k_tx_lane_flip_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ehp_ctrl0_k_ehp_control_reg_attr                                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ehp_ctrl0_k_ehp_control_reg_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ehp_ctrl1_k_outstanding_crd_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ehp_ctrl1_k_outstanding_crd_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ehp_ctrl1_k_tx_rd_th_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ehp_ctrl1_k_tx_rd_th_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff0_k_exvf_msixpba_bir_pf0_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff0_k_exvf_msixpba_bir_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff0_k_exvf_msixpba_offset_pf0_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff0_k_exvf_msixpba_offset_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff1_k_exvf_msixpba_bir_pf1_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff1_k_exvf_msixpba_bir_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff1_k_exvf_msixpba_offset_pf1_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff1_k_exvf_msixpba_offset_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff2_k_exvf_msixpba_bir_pf2_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff2_k_exvf_msixpba_bir_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff2_k_exvf_msixpba_offset_pf2_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff2_k_exvf_msixpba_offset_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff3_k_exvf_msixpba_bir_pf3_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff3_k_exvf_msixpba_bir_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff3_k_exvf_msixpba_offset_pf3_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff3_k_exvf_msixpba_offset_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff4_k_exvf_msixpba_bir_pf4_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff4_k_exvf_msixpba_bir_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff4_k_exvf_msixpba_offset_pf4_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff4_k_exvf_msixpba_offset_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff5_k_exvf_msixpba_bir_pf5_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff5_k_exvf_msixpba_bir_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff5_k_exvf_msixpba_offset_pf5_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff5_k_exvf_msixpba_offset_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff6_k_exvf_msixpba_bir_pf6_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff6_k_exvf_msixpba_bir_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff6_k_exvf_msixpba_offset_pf6_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff6_k_exvf_msixpba_offset_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff7_k_exvf_msixpba_bir_pf7_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff7_k_exvf_msixpba_bir_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff7_k_exvf_msixpba_offset_pf7_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_poff7_k_exvf_msixpba_offset_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff0_k_exvf_msixtable_bir_pf0_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff0_k_exvf_msixtable_bir_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff0_k_exvf_msixtable_offset_pf0_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff0_k_exvf_msixtable_offset_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff1_k_exvf_msixtable_bir_pf1_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff1_k_exvf_msixtable_bir_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff1_k_exvf_msixtable_offset_pf1_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff1_k_exvf_msixtable_offset_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff2_k_exvf_msixtable_bir_pf2_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff2_k_exvf_msixtable_bir_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff2_k_exvf_msixtable_offset_pf2_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff2_k_exvf_msixtable_offset_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff3_k_exvf_msixtable_bir_pf3_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff3_k_exvf_msixtable_bir_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff3_k_exvf_msixtable_offset_pf3_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff3_k_exvf_msixtable_offset_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff4_k_exvf_msixtable_bir_pf4_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff4_k_exvf_msixtable_bir_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff4_k_exvf_msixtable_offset_pf4_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff4_k_exvf_msixtable_offset_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff5_k_exvf_msixtable_bir_pf5_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff5_k_exvf_msixtable_bir_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff5_k_exvf_msixtable_offset_pf5_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff5_k_exvf_msixtable_offset_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff6_k_exvf_msixtable_bir_pf6_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff6_k_exvf_msixtable_bir_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff6_k_exvf_msixtable_offset_pf6_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff6_k_exvf_msixtable_offset_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff7_k_exvf_msixtable_bir_pf7_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff7_k_exvf_msixtable_bir_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff7_k_exvf_msixtable_offset_pf7_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_toff7_k_exvf_msixtable_offset_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize0_k_exvf_msix_tablesize_pf0_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize0_k_exvf_msix_tablesize_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize0_k_exvf_msix_tablesize_pf1_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize0_k_exvf_msix_tablesize_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize1_k_exvf_msix_tablesize_pf2_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize1_k_exvf_msix_tablesize_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize1_k_exvf_msix_tablesize_pf3_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize1_k_exvf_msix_tablesize_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize2_k_exvf_msix_tablesize_pf4_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize2_k_exvf_msix_tablesize_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize2_k_exvf_msix_tablesize_pf5_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize2_k_exvf_msix_tablesize_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize3_k_exvf_msix_tablesize_pf6_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize3_k_exvf_msix_tablesize_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize3_k_exvf_msix_tablesize_pf7_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_m6_tsize3_k_exvf_msix_tablesize_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_cvp_cfg_err_en_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_cvp_cfg_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_dbi_access_err_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_dbi_access_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sd_eq_control1_reg_eval_interval_time),
   
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_multi_lane_control_off_upconfigure_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_multi_lane_control_off_upconfigure_support),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_reg_bar0_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_reg_bar0_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar1_reg_bar1_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_reg_bar2_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_reg_bar2_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_reg_bar3_mem_io                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_reg_bar3_mem_io),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_reg_bar3_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_reg_bar4_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_reg_bar4_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar5_reg_bar5_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_id_nxt_ptr_reg_aux_curr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_id_nxt_ptr_reg_dsi                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_id_nxt_ptr_reg_pme_support                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_reg_ari_acs_fun_grp_cap                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_cap_reg_ari_acs_fun_grp_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_base_class_code                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_program_interface                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_revision_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_subclass_code                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_con_status_reg_no_soft_rst                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_ext_tag_supp                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_ext_tag_supp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_exp_rom_bar_mask_reg_rom_mask                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_config_phy_tx_change                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_config_phy_tx_change),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_select_deemph_var_mux                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_select_deemph_var_mux),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_selectable_deemph_bit_mux                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_selectable_deemph_bit_mux),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_support_mod_ts                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen2_ctrl_off_support_mod_ts),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_eieos_cnt                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_eieos_cnt),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_phase_2_3                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_phase_2_3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_phase_2_3_atg4                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_phase_2_3_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_phase_2_3_atg5                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_phase_2_3_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_redo                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_redo),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_redo_atg4                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_redo_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_redo_atg5                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_eq_redo_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_gen3_equalization_disable                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_gen3_equalization_disable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_ph01_en                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_ph01_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1_substates_off_l1sub_t_l1_2                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1_substates_off_l1sub_t_l1_2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1_substates_off_l1sub_t_power_off                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1_substates_off_l1sub_t_power_off),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_comm_mode_support                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_comm_mode_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_pwr_on_scale_support                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_pwr_on_scale_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_pwr_on_value_support                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_pwr_on_value_support),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_1_aspm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_1_aspm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_2_aspm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_2_aspm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_1_aspm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_1_aspm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_aspm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_aspm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_l1_1sub_cap_enable ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_l1_1sub_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_l1_2sub_cap_enable ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_l1_2sub_cap_enable),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_th_sca                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_th_sca),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_th_val                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_l1_2_th_val),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_t_common_mode                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_l1sub_control1_reg_t_common_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_port_num                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_table_offset_reg_pci_msix_bir                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_table_offset_reg_pci_msix_table_offset                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pipe_loopback_control_off_pipe_loopback                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pipe_loopback_control_off_pipe_loopback),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset4                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset5                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset6                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset7                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_dsp_16g_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset4                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset5                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset6                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset7                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl16g_cap_off_24h_reg_usp_16g_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset4                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset5                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset6                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset7                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_dsp_32g_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset4                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset5                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset6                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset7                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_cap_off_24h_reg_usp_32g_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_capability_reg_no_eq_needed_support                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_capability_reg_no_eq_needed_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_rsvdp_11                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_rsvdp_11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_tx_precode_req                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_tx_precode_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_tx_precoding_on                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_pl32g_status_reg_tx_precoding_on),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_port_force_off_support_part_lanes_rxei_exit                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_port_force_off_support_part_lanes_rxei_exit),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_port_link_ctrl_off_fast_link_mode                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_port_link_ctrl_off_fast_link_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint4                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint5                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_rx_preset_hint5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset4                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset5                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_dsp_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint4                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint5                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_rx_preset_hint5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset4                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset5                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_14h_reg_usp_tx_preset5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint6                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint7                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_rx_preset_hint7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset6                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset7                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_dsp_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint6                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint7                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_rx_preset_hint7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset6                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset6),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset7                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_spcie_cap_off_18h_reg_usp_tx_preset7),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar0_mask_reg_pci_sriov_bar0_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar1_mask_reg_pci_sriov_bar1_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar1_reg_sriov_vf_bar1_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar2_mask_reg_pci_sriov_bar2_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar3_mask_reg_pci_sriov_bar3_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar3_reg_sriov_vf_bar3_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar4_mask_reg_pci_sriov_bar4_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar5_mask_reg_pci_sriov_bar5_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar5_reg_sriov_vf_bar5_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_vf_offset_position_sriov_vf_offset                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_vf_offset_position_sriov_vf_stride                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sup_page_sizes_reg_sriov_sup_page_size                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_device_spec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_vf_device_id_reg_sriov_vf_device_id                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf0_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_at_block                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_egress_control                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_src_valid                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_usp_forwarding                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ats_capabilities_ctrl_reg_invalidate_q_depth                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ats_capabilities_ctrl_reg_page_aligned_req                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_mask_reg_pci_type0_bar0_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_mask_reg_pci_type0_bar0_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_reg_bar0_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_reg_bar0_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar1_mask_reg_pci_type0_bar1_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar1_mask_reg_pci_type0_bar1_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar1_reg_bar1_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_mask_reg_pci_type0_bar2_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_mask_reg_pci_type0_bar2_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_reg_bar2_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_reg_bar2_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar3_mask_reg_pci_type0_bar3_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar3_mask_reg_pci_type0_bar3_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar3_reg_bar3_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_mask_reg_pci_type0_bar4_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_mask_reg_pci_type0_bar4_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_reg_bar4_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_reg_bar4_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar5_mask_reg_pci_type0_bar5_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar5_mask_reg_pci_type0_bar5_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar5_reg_bar5_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cap_id_nxt_ptr_reg_aux_curr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cap_id_nxt_ptr_reg_dsi                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cap_id_nxt_ptr_reg_pme_support                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cardbus_cis_ptr_reg_cardbus_cis_pointer                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_base_class_code                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_program_interface                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_revision_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_subclass_code                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_con_status_reg_no_soft_rst                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_ext_tag_supp                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_ext_tag_supp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_flr_cap                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_control_device_status_pcie_cap_ext_tag_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_id_vendor_id_reg_pci_type0_device_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_id_vendor_id_reg_pci_type0_vendor_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_exp_rom_bar_mask_reg_rom_bar_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_exp_rom_bar_mask_reg_rom_mask                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_exp_rom_base_addr_reg_rom_bar_enable                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_capabilities_reg_pcie_cap_l0s_exit_latency                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_capabilities_reg_pcie_cap_l1_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_capabilities_reg_pcie_cap_port_num                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_control2_link_status2_reg_pcie_cap_sel_deemphasis             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_control_link_status_reg_pcie_cap_active_state_link_pm_control ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_control_link_status_reg_pcie_cap_slot_clk_config              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_pba_offset_reg_pci_msix_pba_bir                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_pba_offset_reg_pci_msix_pba_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_table_offset_reg_pci_msix_bir                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_table_offset_reg_pci_msix_table_offset                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pasid_cap_cntrl_reg_execute_permission_supported                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pasid_cap_cntrl_reg_max_pasid_width                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pasid_cap_cntrl_reg_privileged_mode_supported                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_device_spec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar0_mask_reg_pci_sriov_bar0_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar1_mask_reg_pci_sriov_bar1_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar1_reg_sriov_vf_bar1_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar2_mask_reg_pci_sriov_bar2_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar3_mask_reg_pci_sriov_bar3_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar3_reg_sriov_vf_bar3_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar4_mask_reg_pci_sriov_bar4_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar5_mask_reg_pci_sriov_bar5_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar5_reg_sriov_vf_bar5_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_vf_offset_position_sriov_vf_offset                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_vf_offset_position_sriov_vf_stride                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sup_page_sizes_reg_sriov_sup_page_size                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_int_vec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_device_spec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_vf_device_id_reg_sriov_vf_device_id                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf1_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_at_block                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_egress_control                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_src_valid                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_usp_forwarding                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ats_capabilities_ctrl_reg_invalidate_q_depth                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ats_capabilities_ctrl_reg_page_aligned_req                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_mask_reg_pci_type0_bar0_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_mask_reg_pci_type0_bar0_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_reg_bar0_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_reg_bar0_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar1_mask_reg_pci_type0_bar1_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar1_mask_reg_pci_type0_bar1_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar1_reg_bar1_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_mask_reg_pci_type0_bar2_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_mask_reg_pci_type0_bar2_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_reg_bar2_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_reg_bar2_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar3_mask_reg_pci_type0_bar3_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar3_mask_reg_pci_type0_bar3_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar3_reg_bar3_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_mask_reg_pci_type0_bar4_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_mask_reg_pci_type0_bar4_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_reg_bar4_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_reg_bar4_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar5_mask_reg_pci_type0_bar5_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar5_mask_reg_pci_type0_bar5_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar5_reg_bar5_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cap_id_nxt_ptr_reg_aux_curr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cap_id_nxt_ptr_reg_dsi                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cap_id_nxt_ptr_reg_pme_support                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cardbus_cis_ptr_reg_cardbus_cis_pointer                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_base_class_code                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_program_interface                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_revision_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_subclass_code                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_con_status_reg_no_soft_rst                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_ext_tag_supp                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_ext_tag_supp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_flr_cap                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_control_device_status_pcie_cap_ext_tag_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_id_vendor_id_reg_pci_type0_device_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_id_vendor_id_reg_pci_type0_vendor_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_exp_rom_bar_mask_reg_rom_bar_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_exp_rom_bar_mask_reg_rom_mask                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_exp_rom_base_addr_reg_rom_bar_enable                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_capabilities_reg_pcie_cap_l0s_exit_latency                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_capabilities_reg_pcie_cap_l1_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_capabilities_reg_pcie_cap_port_num                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_control2_link_status2_reg_pcie_cap_sel_deemphasis             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_control_link_status_reg_pcie_cap_active_state_link_pm_control ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_control_link_status_reg_pcie_cap_slot_clk_config              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_pba_offset_reg_pci_msix_pba_bir                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_pba_offset_reg_pci_msix_pba_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_table_offset_reg_pci_msix_bir                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_table_offset_reg_pci_msix_table_offset                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pasid_cap_cntrl_reg_execute_permission_supported                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pasid_cap_cntrl_reg_max_pasid_width                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pasid_cap_cntrl_reg_privileged_mode_supported                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_device_spec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar0_mask_reg_pci_sriov_bar0_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar1_mask_reg_pci_sriov_bar1_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar1_reg_sriov_vf_bar1_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar2_mask_reg_pci_sriov_bar2_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar3_mask_reg_pci_sriov_bar3_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar3_reg_sriov_vf_bar3_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar4_mask_reg_pci_sriov_bar4_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar5_mask_reg_pci_sriov_bar5_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar5_reg_sriov_vf_bar5_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_vf_offset_position_sriov_vf_offset                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_vf_offset_position_sriov_vf_stride                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sup_page_sizes_reg_sriov_sup_page_size                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_int_vec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_device_spec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_vf_device_id_reg_sriov_vf_device_id                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf2_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_at_block                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_egress_control                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_src_valid                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_usp_forwarding                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ats_capabilities_ctrl_reg_invalidate_q_depth                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ats_capabilities_ctrl_reg_page_aligned_req                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_mask_reg_pci_type0_bar0_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_mask_reg_pci_type0_bar0_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_reg_bar0_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_reg_bar0_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar1_mask_reg_pci_type0_bar1_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar1_mask_reg_pci_type0_bar1_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar1_reg_bar1_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_mask_reg_pci_type0_bar2_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_mask_reg_pci_type0_bar2_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_reg_bar2_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_reg_bar2_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar3_mask_reg_pci_type0_bar3_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar3_mask_reg_pci_type0_bar3_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar3_reg_bar3_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_mask_reg_pci_type0_bar4_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_mask_reg_pci_type0_bar4_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_reg_bar4_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_reg_bar4_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar5_mask_reg_pci_type0_bar5_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar5_mask_reg_pci_type0_bar5_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar5_reg_bar5_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cap_id_nxt_ptr_reg_aux_curr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cap_id_nxt_ptr_reg_dsi                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cap_id_nxt_ptr_reg_pme_support                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cardbus_cis_ptr_reg_cardbus_cis_pointer                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_base_class_code                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_program_interface                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_revision_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_subclass_code                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_con_status_reg_no_soft_rst                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_ext_tag_supp                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_ext_tag_supp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_flr_cap                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_control_device_status_pcie_cap_ext_tag_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_id_vendor_id_reg_pci_type0_device_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_id_vendor_id_reg_pci_type0_vendor_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_exp_rom_bar_mask_reg_rom_bar_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_exp_rom_bar_mask_reg_rom_mask                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_exp_rom_base_addr_reg_rom_bar_enable                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_capabilities_reg_pcie_cap_l0s_exit_latency                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_capabilities_reg_pcie_cap_l1_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_capabilities_reg_pcie_cap_port_num                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_control2_link_status2_reg_pcie_cap_sel_deemphasis             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_control_link_status_reg_pcie_cap_active_state_link_pm_control ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_control_link_status_reg_pcie_cap_slot_clk_config              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_pba_offset_reg_pci_msix_pba_bir                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_pba_offset_reg_pci_msix_pba_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_table_offset_reg_pci_msix_bir                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_table_offset_reg_pci_msix_table_offset                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pasid_cap_cntrl_reg_execute_permission_supported                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pasid_cap_cntrl_reg_max_pasid_width                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pasid_cap_cntrl_reg_privileged_mode_supported                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_device_spec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar0_mask_reg_pci_sriov_bar0_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar1_mask_reg_pci_sriov_bar1_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar1_reg_sriov_vf_bar1_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar2_mask_reg_pci_sriov_bar2_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar3_mask_reg_pci_sriov_bar3_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar3_reg_sriov_vf_bar3_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar4_mask_reg_pci_sriov_bar4_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar5_mask_reg_pci_sriov_bar5_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar5_reg_sriov_vf_bar5_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_vf_offset_position_sriov_vf_offset                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_vf_offset_position_sriov_vf_stride                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sup_page_sizes_reg_sriov_sup_page_size                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_int_vec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_device_spec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_vf_device_id_reg_sriov_vf_device_id                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf3_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_at_block                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_egress_control                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_src_valid                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_usp_forwarding                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ats_capabilities_ctrl_reg_invalidate_q_depth                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ats_capabilities_ctrl_reg_page_aligned_req                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_mask_reg_pci_type0_bar0_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_mask_reg_pci_type0_bar0_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_reg_bar0_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_reg_bar0_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar1_mask_reg_pci_type0_bar1_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar1_mask_reg_pci_type0_bar1_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar1_reg_bar1_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_mask_reg_pci_type0_bar2_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_mask_reg_pci_type0_bar2_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_reg_bar2_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_reg_bar2_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar3_mask_reg_pci_type0_bar3_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar3_mask_reg_pci_type0_bar3_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar3_reg_bar3_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_mask_reg_pci_type0_bar4_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_mask_reg_pci_type0_bar4_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_reg_bar4_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_reg_bar4_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar5_mask_reg_pci_type0_bar5_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar5_mask_reg_pci_type0_bar5_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar5_reg_bar5_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cap_id_nxt_ptr_reg_aux_curr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cap_id_nxt_ptr_reg_dsi                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cap_id_nxt_ptr_reg_pme_support                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cardbus_cis_ptr_reg_cardbus_cis_pointer                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_base_class_code                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_program_interface                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_revision_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_subclass_code                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_con_status_reg_no_soft_rst                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_ext_tag_supp                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_ext_tag_supp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_flr_cap                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_control_device_status_pcie_cap_ext_tag_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_id_vendor_id_reg_pci_type0_device_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_id_vendor_id_reg_pci_type0_vendor_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_exp_rom_bar_mask_reg_rom_bar_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_exp_rom_bar_mask_reg_rom_mask                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_exp_rom_base_addr_reg_rom_bar_enable                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_capabilities_reg_pcie_cap_l0s_exit_latency                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_capabilities_reg_pcie_cap_l1_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_capabilities_reg_pcie_cap_port_num                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_control2_link_status2_reg_pcie_cap_sel_deemphasis             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_control_link_status_reg_pcie_cap_active_state_link_pm_control ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_control_link_status_reg_pcie_cap_slot_clk_config              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_pba_offset_reg_pci_msix_pba_bir                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_pba_offset_reg_pci_msix_pba_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_table_offset_reg_pci_msix_bir                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_table_offset_reg_pci_msix_table_offset                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pasid_cap_cntrl_reg_execute_permission_supported                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pasid_cap_cntrl_reg_max_pasid_width                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pasid_cap_cntrl_reg_privileged_mode_supported                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_device_spec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar0_mask_reg_pci_sriov_bar0_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar1_mask_reg_pci_sriov_bar1_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar1_reg_sriov_vf_bar1_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar2_mask_reg_pci_sriov_bar2_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar3_mask_reg_pci_sriov_bar3_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar3_reg_sriov_vf_bar3_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar4_mask_reg_pci_sriov_bar4_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar5_mask_reg_pci_sriov_bar5_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar5_reg_sriov_vf_bar5_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_vf_offset_position_sriov_vf_offset                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_vf_offset_position_sriov_vf_stride                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sup_page_sizes_reg_sriov_sup_page_size                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_int_vec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_device_spec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_vf_device_id_reg_sriov_vf_device_id                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf4_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_at_block                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_egress_control                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_src_valid                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_usp_forwarding                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ats_capabilities_ctrl_reg_invalidate_q_depth                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ats_capabilities_ctrl_reg_page_aligned_req                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_mask_reg_pci_type0_bar0_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_mask_reg_pci_type0_bar0_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_reg_bar0_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_reg_bar0_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar1_mask_reg_pci_type0_bar1_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar1_mask_reg_pci_type0_bar1_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar1_reg_bar1_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_mask_reg_pci_type0_bar2_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_mask_reg_pci_type0_bar2_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_reg_bar2_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_reg_bar2_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar3_mask_reg_pci_type0_bar3_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar3_mask_reg_pci_type0_bar3_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar3_reg_bar3_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_mask_reg_pci_type0_bar4_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_mask_reg_pci_type0_bar4_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_reg_bar4_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_reg_bar4_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar5_mask_reg_pci_type0_bar5_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar5_mask_reg_pci_type0_bar5_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar5_reg_bar5_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cap_id_nxt_ptr_reg_aux_curr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cap_id_nxt_ptr_reg_dsi                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cap_id_nxt_ptr_reg_pme_support                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cardbus_cis_ptr_reg_cardbus_cis_pointer                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_base_class_code                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_program_interface                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_revision_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_subclass_code                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_con_status_reg_no_soft_rst                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_ext_tag_supp                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_ext_tag_supp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_flr_cap                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_control_device_status_pcie_cap_ext_tag_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_id_vendor_id_reg_pci_type0_device_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_id_vendor_id_reg_pci_type0_vendor_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_exp_rom_bar_mask_reg_rom_bar_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_exp_rom_bar_mask_reg_rom_mask                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_exp_rom_base_addr_reg_rom_bar_enable                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_capabilities_reg_pcie_cap_l0s_exit_latency                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_capabilities_reg_pcie_cap_l1_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_capabilities_reg_pcie_cap_port_num                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_control2_link_status2_reg_pcie_cap_sel_deemphasis             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_control_link_status_reg_pcie_cap_active_state_link_pm_control ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_control_link_status_reg_pcie_cap_slot_clk_config              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_pba_offset_reg_pci_msix_pba_bir                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_pba_offset_reg_pci_msix_pba_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_table_offset_reg_pci_msix_bir                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_table_offset_reg_pci_msix_table_offset                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pasid_cap_cntrl_reg_execute_permission_supported                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pasid_cap_cntrl_reg_max_pasid_width                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pasid_cap_cntrl_reg_privileged_mode_supported                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_device_spec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar0_mask_reg_pci_sriov_bar0_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar1_mask_reg_pci_sriov_bar1_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar1_reg_sriov_vf_bar1_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar2_mask_reg_pci_sriov_bar2_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar3_mask_reg_pci_sriov_bar3_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar3_reg_sriov_vf_bar3_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar4_mask_reg_pci_sriov_bar4_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar5_mask_reg_pci_sriov_bar5_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar5_reg_sriov_vf_bar5_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_vf_offset_position_sriov_vf_offset                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_vf_offset_position_sriov_vf_stride                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sup_page_sizes_reg_sriov_sup_page_size                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_int_vec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_device_spec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_vf_device_id_reg_sriov_vf_device_id                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf5_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_at_block                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_egress_control                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_src_valid                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_usp_forwarding                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ats_capabilities_ctrl_reg_invalidate_q_depth                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ats_capabilities_ctrl_reg_page_aligned_req                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_mask_reg_pci_type0_bar0_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_mask_reg_pci_type0_bar0_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_reg_bar0_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_reg_bar0_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar1_mask_reg_pci_type0_bar1_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar1_mask_reg_pci_type0_bar1_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar1_reg_bar1_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_mask_reg_pci_type0_bar2_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_mask_reg_pci_type0_bar2_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_reg_bar2_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_reg_bar2_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar3_mask_reg_pci_type0_bar3_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar3_mask_reg_pci_type0_bar3_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar3_reg_bar3_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_mask_reg_pci_type0_bar4_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_mask_reg_pci_type0_bar4_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_reg_bar4_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_reg_bar4_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar5_mask_reg_pci_type0_bar5_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar5_mask_reg_pci_type0_bar5_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar5_reg_bar5_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cap_id_nxt_ptr_reg_aux_curr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cap_id_nxt_ptr_reg_dsi                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cap_id_nxt_ptr_reg_pme_support                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cardbus_cis_ptr_reg_cardbus_cis_pointer                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_base_class_code                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_program_interface                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_revision_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_subclass_code                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_con_status_reg_no_soft_rst                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_ext_tag_supp                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_ext_tag_supp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_flr_cap                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_control_device_status_pcie_cap_ext_tag_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_id_vendor_id_reg_pci_type0_device_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_id_vendor_id_reg_pci_type0_vendor_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_exp_rom_bar_mask_reg_rom_bar_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_exp_rom_bar_mask_reg_rom_mask                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_exp_rom_base_addr_reg_rom_bar_enable                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_capabilities_reg_pcie_cap_l0s_exit_latency                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_capabilities_reg_pcie_cap_l1_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_capabilities_reg_pcie_cap_port_num                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_control2_link_status2_reg_pcie_cap_sel_deemphasis             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_control_link_status_reg_pcie_cap_active_state_link_pm_control ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_control_link_status_reg_pcie_cap_slot_clk_config              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_pba_offset_reg_pci_msix_pba_bir                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_pba_offset_reg_pci_msix_pba_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_table_offset_reg_pci_msix_bir                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_table_offset_reg_pci_msix_table_offset                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pasid_cap_cntrl_reg_execute_permission_supported                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pasid_cap_cntrl_reg_max_pasid_width                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pasid_cap_cntrl_reg_privileged_mode_supported                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_device_spec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar0_mask_reg_pci_sriov_bar0_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar1_mask_reg_pci_sriov_bar1_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar1_reg_sriov_vf_bar1_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar2_mask_reg_pci_sriov_bar2_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar3_mask_reg_pci_sriov_bar3_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar3_reg_sriov_vf_bar3_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar4_mask_reg_pci_sriov_bar4_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar5_mask_reg_pci_sriov_bar5_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar5_reg_sriov_vf_bar5_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_vf_offset_position_sriov_vf_offset                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_vf_offset_position_sriov_vf_stride                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sup_page_sizes_reg_sriov_sup_page_size                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_int_vec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_device_spec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_vf_device_id_reg_sriov_vf_device_id                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf6_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_at_block                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_egress_control                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_src_valid                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_usp_forwarding                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ats_capabilities_ctrl_reg_invalidate_q_depth                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ats_capabilities_ctrl_reg_page_aligned_req                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_mask_reg_pci_type0_bar0_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_mask_reg_pci_type0_bar0_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_reg_bar0_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_reg_bar0_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar1_mask_reg_pci_type0_bar1_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar1_mask_reg_pci_type0_bar1_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar1_reg_bar1_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_mask_reg_pci_type0_bar2_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_mask_reg_pci_type0_bar2_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_reg_bar2_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_reg_bar2_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar3_mask_reg_pci_type0_bar3_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar3_mask_reg_pci_type0_bar3_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar3_reg_bar3_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_mask_reg_pci_type0_bar4_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_mask_reg_pci_type0_bar4_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_reg_bar4_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_reg_bar4_type                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar5_mask_reg_pci_type0_bar5_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar5_mask_reg_pci_type0_bar5_mask                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar5_reg_bar5_prefetch                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cap_id_nxt_ptr_reg_aux_curr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cap_id_nxt_ptr_reg_dsi                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cap_id_nxt_ptr_reg_pme_support                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cardbus_cis_ptr_reg_cardbus_cis_pointer                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_cardbus_cis_ptr_reg_cardbus_cis_pointer)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_base_class_code                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_program_interface                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_revision_id                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_subclass_code                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_con_status_reg_no_soft_rst                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_ext_tag_supp                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_ext_tag_supp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_flr_cap                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_control_device_status_pcie_cap_ext_tag_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_id_vendor_id_reg_pci_type0_device_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_id_vendor_id_reg_pci_type0_vendor_id                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_exp_rom_bar_mask_reg_rom_bar_enabled                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_exp_rom_bar_mask_reg_rom_mask                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_exp_rom_base_addr_reg_rom_bar_enable                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_capabilities_reg_pcie_cap_l0s_exit_latency                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_capabilities_reg_pcie_cap_l1_exit_latency                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_capabilities_reg_pcie_cap_port_num                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_control2_link_status2_reg_pcie_cap_sel_deemphasis             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_control_link_status_reg_pcie_cap_active_state_link_pm_control ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_control_link_status_reg_pcie_cap_slot_clk_config              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_pba_offset_reg_pci_msix_pba_bir                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_pba_offset_reg_pci_msix_pba_offset                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_table_offset_reg_pci_msix_bir                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_table_offset_reg_pci_msix_table_offset                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pasid_cap_cntrl_reg_execute_permission_supported                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pasid_cap_cntrl_reg_max_pasid_width                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pasid_cap_cntrl_reg_privileged_mode_supported                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                               ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_sriov_vf_offset_position_shadow_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_device_spec                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar0_mask_reg_pci_sriov_bar0_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar0_mask_reg_pci_sriov_bar0_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar0_reg_sriov_vf_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar1_mask_reg_pci_sriov_bar1_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar1_mask_reg_pci_sriov_bar1_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar1_reg_sriov_vf_bar1_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar1_reg_sriov_vf_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar2_mask_reg_pci_sriov_bar2_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar2_mask_reg_pci_sriov_bar2_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar2_reg_sriov_vf_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar3_mask_reg_pci_sriov_bar3_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar3_mask_reg_pci_sriov_bar3_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar3_reg_sriov_vf_bar3_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar3_reg_sriov_vf_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar4_mask_reg_pci_sriov_bar4_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar4_mask_reg_pci_sriov_bar4_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_type                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar4_reg_sriov_vf_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar5_mask_reg_pci_sriov_bar5_mask                            ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar5_mask_reg_pci_sriov_bar5_mask)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar5_reg_sriov_vf_bar5_prefetch                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_bar5_reg_sriov_vf_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_vf_offset_position_sriov_vf_offset                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_vf_offset_position_sriov_vf_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_vf_offset_position_sriov_vf_stride                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sriov_vf_offset_position_sriov_vf_stride),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sup_page_sizes_reg_sriov_sup_page_size                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_sup_page_sizes_reg_sriov_sup_page_size)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_int_vec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_size                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_device_spec                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_vf_device_id_reg_sriov_vf_device_id                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pf7_vf_device_id_reg_sriov_vf_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pfvf_sel_vsec_enable_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_pfvf_sel_vsec_enable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_phy_rxelecidle_k_rxelecidle_disable_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_phy_rxelecidle_k_rxelecidle_disable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_phy_rxtermination_k_rxtermination_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_phy_rxtermination_k_rxtermination_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ptm_ctrl_k_cfg_ptm_auto_update_signal_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ptm_ctrl_k_cfg_ptm_auto_update_signal_attr),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ptm_adj_lsb_k_cfg_ptm_local_clock_adj_lsb_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ptm_adj_lsb_k_cfg_ptm_local_clock_adj_lsb_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ptm_adj_msb_k_cfg_ptm_local_clock_adj_msb_attr ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_ptm_adj_msb_k_cfg_ptm_local_clock_adj_msb_attr),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_err_en_correct_err_en_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_err_en_correct_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_err_en_fatal_err_en_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_err_en_fatal_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_err_en_nonfatal_err_en_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_err_en_nonfatal_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_bw_mgt_int_en_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_bw_mgt_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_link_eq_req_int_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_link_eq_req_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_pme_int_en_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_cfg_pme_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_hp_int_en_attr                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_hp_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_hp_pme_en_attr                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_hp_pme_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_inta_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_inta_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_intb_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_intb_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_intc_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_intc_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_intd_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_rp_irq_en_intd_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_sriov_misc_ctrl_k_nonsriov_mode_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_sriov_misc_ctrl_k_nonsriov_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_stagger_control_k_stag_dlycnt_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_stagger_control_k_stag_dlycnt_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_stagger_control_k_stag_mode_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_stagger_control_k_stag_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id0_k_exvf_subsysid_pf0_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id0_k_exvf_subsysid_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id0_k_exvf_subsysid_pf1_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id0_k_exvf_subsysid_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id1_k_exvf_subsysid_pf2_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id1_k_exvf_subsysid_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id1_k_exvf_subsysid_pf3_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id1_k_exvf_subsysid_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id2_k_exvf_subsysid_pf4_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id2_k_exvf_subsysid_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id2_k_exvf_subsysid_pf5_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id2_k_exvf_subsysid_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id3_k_exvf_subsysid_pf6_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id3_k_exvf_subsysid_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id3_k_exvf_subsysid_pf7_attr                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_subs_id3_k_exvf_subsysid_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf0_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf1_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablelocation_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablesize_pf0_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablesize_pf0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablesize_pf1_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl0_k_exvf_tph_sttablesize_pf1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf2_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf3_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablelocation_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablesize_pf2_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablesize_pf2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablesize_pf3_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl1_k_exvf_tph_sttablesize_pf3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf4_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf5_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablelocation_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablesize_pf4_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablesize_pf4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablesize_pf5_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl2_k_exvf_tph_sttablesize_pf5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf6_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf7_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablelocation_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablesize_pf6_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablesize_pf6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablesize_pf7_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tph_ctl3_k_exvf_tph_sttablesize_pf7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tx_common_mode_k_txcommonmode_disable_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_tx_common_mode_k_txcommonmode_disable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_100_k_pf4_virtio_offset_cfg3_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_100_k_pf4_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_102_k_pf4_virtio_offset_cfg4_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_102_k_pf4_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_103_k_pf4_virtio_offset_cfg4_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_103_k_pf4_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_104_k_pf4_virtio_offset_cfg4_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_104_k_pf4_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_106_k_pf4_virtio_offset_cfg5_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_106_k_pf4_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_107_k_pf4_virtio_offset_cfg5_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_107_k_pf4_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_108_k_pf4_virtio_offset_cfg5_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_108_k_pf4_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_109_k_pf4_virtio_offset_cfg5_cfg_data_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_109_k_pf4_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_111_k_pf5_virtio_offset_cfg1_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_111_k_pf5_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_112_k_pf5_virtio_offset_cfg1_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_112_k_pf5_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_113_k_pf5_virtio_offset_cfg1_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_113_k_pf5_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_115_k_pf5_virtio_offset_cfg2_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_115_k_pf5_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_116_k_pf5_virtio_offset_cfg2_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_116_k_pf5_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_117_k_pf5_virtio_offset_cfg2_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_117_k_pf5_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_118_k_pf5_virtio_offset_cfg2_notify_off_multiplier_attr         ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_118_k_pf5_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_120_k_pf5_virtio_offset_cfg3_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_120_k_pf5_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_121_k_pf5_virtio_offset_cfg3_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_121_k_pf5_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_122_k_pf5_virtio_offset_cfg3_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_122_k_pf5_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_124_k_pf5_virtio_offset_cfg4_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_124_k_pf5_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_125_k_pf5_virtio_offset_cfg4_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_125_k_pf5_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_126_k_pf5_virtio_offset_cfg4_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_126_k_pf5_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_128_k_pf5_virtio_offset_cfg5_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_128_k_pf5_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_129_k_pf5_virtio_offset_cfg5_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_129_k_pf5_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_130_k_pf5_virtio_offset_cfg5_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_130_k_pf5_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_131_k_pf5_virtio_offset_cfg5_cfg_data_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_131_k_pf5_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_133_k_pf6_virtio_offset_cfg1_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_133_k_pf6_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_134_k_pf6_virtio_offset_cfg1_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_134_k_pf6_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_135_k_pf6_virtio_offset_cfg1_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_135_k_pf6_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_137_k_pf6_virtio_offset_cfg2_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_137_k_pf6_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_138_k_pf6_virtio_offset_cfg2_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_138_k_pf6_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_139_k_pf6_virtio_offset_cfg2_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_139_k_pf6_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_140_k_pf6_virtio_offset_cfg2_notify_off_multiplier_attr         ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_140_k_pf6_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_142_k_pf6_virtio_offset_cfg3_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_142_k_pf6_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_143_k_pf6_virtio_offset_cfg3_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_143_k_pf6_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_144_k_pf6_virtio_offset_cfg3_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_144_k_pf6_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_146_k_pf6_virtio_offset_cfg4_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_146_k_pf6_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_147_k_pf6_virtio_offset_cfg4_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_147_k_pf6_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_148_k_pf6_virtio_offset_cfg4_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_148_k_pf6_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_150_k_pf6_virtio_offset_cfg5_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_150_k_pf6_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_151_k_pf6_virtio_offset_cfg5_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_151_k_pf6_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_152_k_pf6_virtio_offset_cfg5_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_152_k_pf6_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_153_k_pf6_virtio_offset_cfg5_cfg_data_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_153_k_pf6_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_155_k_pf7_virtio_offset_cfg1_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_155_k_pf7_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_156_k_pf7_virtio_offset_cfg1_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_156_k_pf7_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_157_k_pf7_virtio_offset_cfg1_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_157_k_pf7_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_159_k_pf7_virtio_offset_cfg2_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_159_k_pf7_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_160_k_pf7_virtio_offset_cfg2_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_160_k_pf7_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_161_k_pf7_virtio_offset_cfg2_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_161_k_pf7_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_162_k_pf7_virtio_offset_cfg2_notify_off_multiplier_attr         ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_162_k_pf7_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_164_k_pf7_virtio_offset_cfg3_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_164_k_pf7_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_165_k_pf7_virtio_offset_cfg3_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_165_k_pf7_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_166_k_pf7_virtio_offset_cfg3_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_166_k_pf7_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_168_k_pf7_virtio_offset_cfg4_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_168_k_pf7_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_169_k_pf7_virtio_offset_cfg4_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_169_k_pf7_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_170_k_pf7_virtio_offset_cfg4_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_170_k_pf7_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_172_k_pf7_virtio_offset_cfg5_cap_bar_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_172_k_pf7_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_173_k_pf7_virtio_offset_cfg5_cap_offset_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_173_k_pf7_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_174_k_pf7_virtio_offset_cfg5_cap_length_attr                    ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_174_k_pf7_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_175_k_pf7_virtio_offset_cfg5_cfg_data_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_175_k_pf7_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_23_k_pf1_virtio_offset_cfg1_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_23_k_pf1_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_24_k_pf1_virtio_offset_cfg1_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_24_k_pf1_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_25_k_pf1_virtio_offset_cfg1_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_25_k_pf1_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_27_k_pf1_virtio_offset_cfg2_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_27_k_pf1_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_28_k_pf1_virtio_offset_cfg2_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_28_k_pf1_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_29_k_pf1_virtio_offset_cfg2_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_29_k_pf1_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_30_k_pf1_virtio_offset_cfg2_notify_off_multiplier_attr          ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_30_k_pf1_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_32_k_pf1_virtio_offset_cfg3_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_32_k_pf1_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_33_k_pf1_virtio_offset_cfg3_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_33_k_pf1_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_34_k_pf1_virtio_offset_cfg3_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_34_k_pf1_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_36_k_pf1_virtio_offset_cfg4_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_36_k_pf1_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_37_k_pf1_virtio_offset_cfg4_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_37_k_pf1_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_38_k_pf1_virtio_offset_cfg4_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_38_k_pf1_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_40_k_pf1_virtio_offset_cfg5_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_40_k_pf1_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_41_k_pf1_virtio_offset_cfg5_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_41_k_pf1_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_42_k_pf1_virtio_offset_cfg5_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_42_k_pf1_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_43_k_pf1_virtio_offset_cfg5_cfg_data_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_43_k_pf1_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_45_k_pf2_virtio_offset_cfg1_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_45_k_pf2_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_46_k_pf2_virtio_offset_cfg1_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_46_k_pf2_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_47_k_pf2_virtio_offset_cfg1_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_47_k_pf2_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_49_k_pf2_virtio_offset_cfg2_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_49_k_pf2_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_50_k_pf2_virtio_offset_cfg2_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_50_k_pf2_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_51_k_pf2_virtio_offset_cfg2_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_51_k_pf2_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_52_k_pf2_virtio_offset_cfg2_notify_off_multiplier_attr          ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_52_k_pf2_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_54_k_pf2_virtio_offset_cfg3_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_54_k_pf2_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_55_k_pf2_virtio_offset_cfg3_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_55_k_pf2_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_56_k_pf2_virtio_offset_cfg3_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_56_k_pf2_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_58_k_pf2_virtio_offset_cfg4_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_58_k_pf2_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_59_k_pf2_virtio_offset_cfg4_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_59_k_pf2_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_60_k_pf2_virtio_offset_cfg4_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_60_k_pf2_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_62_k_pf2_virtio_offset_cfg5_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_62_k_pf2_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_63_k_pf2_virtio_offset_cfg5_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_63_k_pf2_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_64_k_pf2_virtio_offset_cfg5_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_64_k_pf2_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_65_k_pf2_virtio_offset_cfg5_cfg_data_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_65_k_pf2_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_67_k_pf3_virtio_offset_cfg1_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_67_k_pf3_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_68_k_pf3_virtio_offset_cfg1_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_68_k_pf3_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_69_k_pf3_virtio_offset_cfg1_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_69_k_pf3_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_71_k_pf3_virtio_offset_cfg2_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_71_k_pf3_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_72_k_pf3_virtio_offset_cfg2_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_72_k_pf3_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_73_k_pf3_virtio_offset_cfg2_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_73_k_pf3_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_74_k_pf3_virtio_offset_cfg2_notify_off_multiplier_attr          ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_74_k_pf3_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_76_k_pf3_virtio_offset_cfg3_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_76_k_pf3_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_77_k_pf3_virtio_offset_cfg3_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_77_k_pf3_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_78_k_pf3_virtio_offset_cfg3_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_78_k_pf3_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr                      ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_80_k_pf3_virtio_offset_cfg4_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_80_k_pf3_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_81_k_pf3_virtio_offset_cfg4_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_81_k_pf3_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_82_k_pf3_virtio_offset_cfg4_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_82_k_pf3_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_84_k_pf3_virtio_offset_cfg5_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_84_k_pf3_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_85_k_pf3_virtio_offset_cfg5_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_85_k_pf3_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_86_k_pf3_virtio_offset_cfg5_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_86_k_pf3_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_87_k_pf3_virtio_offset_cfg5_cfg_data_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_87_k_pf3_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_89_k_pf4_virtio_offset_cfg1_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_89_k_pf4_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr           ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_90_k_pf4_virtio_offset_cfg1_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_90_k_pf4_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_91_k_pf4_virtio_offset_cfg1_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_91_k_pf4_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_93_k_pf4_virtio_offset_cfg2_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_93_k_pf4_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_94_k_pf4_virtio_offset_cfg2_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_94_k_pf4_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_95_k_pf4_virtio_offset_cfg2_cap_length_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_95_k_pf4_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_96_k_pf4_virtio_offset_cfg2_notify_off_multiplier_attr          ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_96_k_pf4_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_98_k_pf4_virtio_offset_cfg3_cap_bar_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_98_k_pf4_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_99_k_pf4_virtio_offset_cfg3_cap_offset_attr                     ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_99_k_pf4_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_cii_ctrl_k_cfg_update_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_cii_ctrl_k_cfg_update_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_cii_ctrl_k_cii_en_attr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_cii_ctrl_k_cii_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_cvp_mode                                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_cvp_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_drop_vendor0_msg                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_drop_vendor0_msg),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_drop_vendor1_msg                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_drop_vendor1_msg),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_ep_native                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_ep_native),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_maxpayload_size                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_maxpayload_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_num_of_lanes                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_num_of_lanes),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_acs_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_ats_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_bar1_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_bar3_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_bar5_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_dlink_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_dlink_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_acs_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_ats_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_msix_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_tph_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_virtio_en                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_io_decode                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_io_decode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_ltr_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_ltr_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_msi_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_msix_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_pasid_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_prefetch_decode                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_prefetch_decode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_prs_ext_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_ras_des_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sn_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_num_vf_non_ari                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar0_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar1_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar2_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar3_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar4_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar5_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_tph_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_user_vsec_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_virtio_dev_specific_conf_en                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_virtio_en                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_vsecras_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf0_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_acs_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_ats_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_bar1_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_bar3_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_bar5_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_enable                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_acs_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_ats_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_msix_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_tph_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_virtio_en                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_msi_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_msix_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_pasid_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_prs_ext_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_ras_des_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sn_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_num_vf_non_ari                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar0_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar1_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar2_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar3_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar4_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar5_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_tph_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_user_vsec_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_user_vsec_offset                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_virtio_dev_specific_conf_en                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_virtio_en                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_vsecras_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf1_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_acs_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_ats_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_bar1_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_bar3_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_bar5_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_enable                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_acs_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_ats_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_msix_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_tph_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_virtio_en                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_msi_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_msix_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_pasid_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_prs_ext_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_ras_des_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sn_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_num_vf_non_ari                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar0_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar1_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar2_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar3_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar4_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar5_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_tph_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_user_vsec_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_user_vsec_offset                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_virtio_dev_specific_conf_en                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_virtio_en                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_vsecras_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf2_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_acs_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_ats_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_bar1_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_bar3_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_bar5_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_enable                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_acs_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_ats_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_msix_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_tph_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_virtio_en                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_msi_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_msix_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_pasid_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_prs_ext_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_ras_des_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sn_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_num_vf_non_ari                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar0_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar1_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar2_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar3_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar4_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar5_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_tph_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_user_vsec_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_user_vsec_offset                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_virtio_dev_specific_conf_en                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_virtio_en                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_vsecras_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf3_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_acs_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_ats_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_bar1_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_bar3_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_bar5_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_enable                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_acs_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_ats_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_msix_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_tph_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_virtio_en                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_msi_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_msix_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_pasid_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_prs_ext_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_ras_des_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sn_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_num_vf_non_ari                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar0_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar1_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar2_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar3_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar4_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar5_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_tph_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_user_vsec_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_user_vsec_offset                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_virtio_dev_specific_conf_en                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_virtio_en                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_vsecras_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf4_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_acs_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_ats_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_bar1_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_bar3_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_bar5_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_enable                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_acs_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_ats_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_msix_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_tph_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_virtio_en                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_msi_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_msix_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_pasid_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_prs_ext_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_ras_des_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sn_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_num_vf_non_ari                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar0_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar1_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar2_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar3_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar4_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar5_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_tph_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_user_vsec_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_user_vsec_offset                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_virtio_dev_specific_conf_en                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_virtio_en                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_vsecras_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf5_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_acs_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_ats_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_bar1_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_bar3_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_bar5_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_enable                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_acs_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_ats_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_msix_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_tph_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_virtio_en                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_msi_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_msix_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_pasid_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_prs_ext_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_ras_des_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sn_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_num_vf_non_ari                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar0_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar1_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar2_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar3_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar4_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar5_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_tph_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_user_vsec_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_user_vsec_offset                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_virtio_dev_specific_conf_en                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_virtio_en                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_vsecras_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf6_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_acs_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_ats_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_bar1_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_bar3_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_bar5_mask_bit0                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_enable                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_acs_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_ats_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_msix_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_tph_cap_enable                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_virtio_en                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_exvf_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_msi_enable                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_msix_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_pasid_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_prs_ext_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_ras_des_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sn_cap_enable                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_num_vf_non_ari                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_num_vf_non_ari),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar0_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar1_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar2_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar3_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar4_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar5_enabled                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_sriov_vf_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_tph_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_user_vsec_cap_enable                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_user_vsec_offset                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_user_vsec_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_virtio_dev_specific_conf_en                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_virtio_en                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_vsecras_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_pf7_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_ptm_autoupdate                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_ptm_autoupdate),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p1p3_inst_rnr_pcie_ip8_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_addr_size0_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_addr_size0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_pf_en0_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_pf_en0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_start_addr0_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_0_k_cii_start_addr0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_addr_size1_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_addr_size1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_pf_en1_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_pf_en1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_start_addr1_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_1_k_cii_start_addr1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_addr_size2_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_addr_size2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_pf_en2_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_pf_en2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_start_addr2_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_2_k_cii_start_addr2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_addr_size3_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_addr_size3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_pf_en3_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_pf_en3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_start_addr3_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_3_k_cii_start_addr3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_addr_size4_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_addr_size4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_pf_en4_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_pf_en4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_start_addr4_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_4_k_cii_start_addr4_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_addr_size5_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_addr_size5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_pf_en5_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_pf_en5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_start_addr5_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_5_k_cii_start_addr5_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_addr_size6_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_addr_size6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_pf_en6_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_pf_en6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_start_addr6_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_6_k_cii_start_addr6_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_addr_size7_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_addr_size7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_pf_en7_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_pf_en7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_start_addr7_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cii_range_7_k_cii_start_addr7_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_cfg_sys_serr_dis_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_fixedcred_attr                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_fixedcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_mcred_attr                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_mcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_reloadcred_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_reloadcred_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_tlp_serr_dis_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_ctrl0_k_tlp_serr_dis_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_mmio_access_ctrl_grant_attr                                          ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_mmio_access_ctrl_grant_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_opcode_ctrl_lock_attr                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_csb_opcode_ctrl_lock_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_compressed_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_compressed_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_encrypted_attr                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl0_k_encrypted_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_devbrd_type_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_devbrd_type_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_vsec_next_offset_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_ctrl1_k_vsec_next_offset_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_cvp_irq_en_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_cvp_irq_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_gpio_irq_attr                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_gpio_irq_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_irq_ctrl_k_irq_misc_ctrl_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid0_k_jtag_id_0_attr                                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid0_k_jtag_id_0_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid1_k_jtag_id_1_attr                                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid1_k_jtag_id_1_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid2_k_jtag_id_2_attr                                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid2_k_jtag_id_2_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid3_k_jtag_id_3_attr                                             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_cvp_jtagid3_k_jtag_id_3_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_dfd_en_attr                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_dfd_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_patcntr_en_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_ctrl0_k_patcntr_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_0_attr                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_1_attr                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_2_attr                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_3_attr                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_data_sel_3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_trig_sel_0_attr                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_trig_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_trig_sel_1_attr                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_trig_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_0_attr                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_0_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_1_attr                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_1_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_2_attr                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_2_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_3_attr                                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dfd_xbar_sel_3_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_aib_loopback_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_crs_en_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_pld_crs_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_rx_lane_flip_en_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_rx_lane_flip_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_sris_mode_attr                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_sris_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_tx_lane_flip_en_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_dwc_ctrl0_k_tx_lane_flip_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_ehp_ctrl0_k_ehp_control_reg_attr                                         ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_ehp_ctrl0_k_ehp_control_reg_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_outstanding_crd_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_outstanding_crd_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_tx_rd_th_attr                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_ehp_ctrl1_k_tx_rd_th_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cfg_ram_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_csb_msg_dropped_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cvp_cfg_err_en_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_cvp_cfg_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dbi_access_err_en_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dbi_access_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_rx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_dwc_tx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_rx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_ehp_tx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_pipe_msgbuf_overflow_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_to_ack_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_irq_en_k_rcvd_pm_turnoff_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cfg_ram_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_csb_msg_dropped_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_cvp_cfg_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dbi_access_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_rx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_dwc_tx_parity_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_rx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_correctable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_ehp_tx_uncorrectable_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_pipe_msgbuf_overflow_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_to_ack_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_misc_ssm_irq_en_k_rcvd_pm_turnoff_en_attr),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_sd_eq_control1_reg_eval_interval_time ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_sd_eq_control1_reg_eval_interval_time),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_prs_req_capacity_reg_prs_outstanding_capacity),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_multi_lane_control_off_upconfigure_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_multi_lane_control_off_upconfigure_support),
   
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_at_block),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_direct_translated_p2p),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_egress_ctrl_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_cpl_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_egress_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_p2p_req_redirect),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_src_valid),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_acs_capabilities_ctrl_reg_acs_usp_forwarding),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_invalidate_q_depth),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ats_capabilities_ctrl_reg_page_aligned_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_mask_reg_pci_type0_bar0_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_prefetch                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_type                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar0_reg_bar0_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar1_mask_reg_pci_type0_bar1_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar1_reg_bar1_prefetch                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar1_reg_bar1_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_mask_reg_pci_type0_bar2_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_prefetch                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_type                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar2_reg_bar2_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_mask_reg_pci_type0_bar3_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_mem_io                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_mem_io),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_prefetch                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar3_reg_bar3_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_mask_reg_pci_type0_bar4_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_prefetch                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_type                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar4_reg_bar4_type),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar5_mask_reg_pci_type0_bar5_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar5_reg_bar5_prefetch                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bar5_reg_bar5_prefetch),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bist_header_type_latency_cache_line_size_reg_multi_func              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_bist_header_type_latency_cache_line_size_reg_multi_func),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_aux_curr                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_aux_curr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_dsi                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_dsi),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_pme_support                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_id_nxt_ptr_reg_pme_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_reg_ari_acs_fun_grp_cap                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_cap_reg_ari_acs_fun_grp_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_base_class_code                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_base_class_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_program_interface                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_program_interface),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_revision_id                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_revision_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_subclass_code                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_class_code_revision_id_subclass_code),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_con_status_reg_no_soft_rst                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_con_status_reg_no_soft_rst),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_dev3_ext_cap_device_control3_reg_dev3_cap_dmwr_egress_blk),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l0s_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ep_l1_accpt_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ext_tag_supp                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_ext_tag_supp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_capabilities_reg_pcie_cap_flr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_control_device_status_pcie_cap_ext_tag_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_device_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_device_id_vendor_id_reg_pci_type0_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_bar_enabled),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_mask                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_exp_rom_bar_mask_reg_rom_mask),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_exp_rom_base_addr_reg_rom_bar_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_auto_lane_flip_ctrl_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_config_phy_tx_change                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_config_phy_tx_change),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_select_deemph_var_mux                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_select_deemph_var_mux),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_selectable_deemph_bit_mux                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_selectable_deemph_bit_mux),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_support_mod_ts                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen2_ctrl_off_support_mod_ts),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_eval_2ms_disable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_phase23_exit_mode_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_eq_pset_req_vec_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_eq_control_off_gen3_lower_rate_eq_redo_enable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_eieos_cnt_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg4                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg5                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_phase_2_3_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg4                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg5                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_eq_redo_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_gen3_equalization_disable_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_ph01_en_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg4),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_gen3_related_off_rxeq_rgrdless_rxts_atg5),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_l1_2                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_l1_2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_power_off                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1_substates_off_l1sub_t_power_off),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_comm_mode_support                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_comm_mode_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_scale_support                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_scale_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_value_support                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_pwr_on_value_support),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_aspm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_aspm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_aspm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_aspm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_1_pcipm_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_capability_reg_l1_2_pcipm_support),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_aspm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_aspm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_1_pcipm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_aspm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_aspm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_pcipm_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_1sub_cap_enable ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_1sub_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_2sub_cap_enable ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_l1_2sub_cap_enable),

   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_sca                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_sca),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_val                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_l1_2_th_val),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_t_common_mode                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_l1sub_control1_reg_t_common_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l0s_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_l1_exit_latency),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_port_num                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_port_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_capabilities_reg_pcie_cap_surprise_down_err_rep_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control2_link_status2_reg_pcie_cap_sel_deemphasis),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_active_state_link_pm_control),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_auto_bw_int_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_link_bw_man_int_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_link_control_link_status_reg_pcie_cap_slot_clk_config),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_max_latency_min_grant_interrupt_pin_interrupt_line_reg_int_pin),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_misc_control_1_off_port_logic_wr_disable                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_misc_control_1_off_port_logic_wr_disable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_pba_offset_reg_pci_msix_pba_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_bir                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_bir),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_table_offset                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_msix_table_offset_reg_pci_msix_table_offset),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_execute_permission_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_max_pasid_width),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pasid_cap_cntrl_reg_privileged_mode_supported),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_64_bit_addr_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_ext_data_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msi_cap_id_next_ctrl_reg_pci_msi_multiple_msg_cap),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_int_msg_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pcie_cap_id_pcie_next_cap_ptr_pcie_cap_reg_pcie_slot_imp),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pipe_loopback_control_off_pipe_loopback                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pipe_loopback_control_off_pipe_loopback),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_dsp_16g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl16g_cap_off_20h_reg_usp_16g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_dsp_32g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_cap_off_20h_reg_usp_32g_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_capability_reg_no_eq_needed_support                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_capability_reg_no_eq_needed_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_no_eq_needed_rcvd),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rsvdp_11                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rsvdp_11),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_rx_enh_link_behavior_ctrl),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precode_req                                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precode_req),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precoding_on                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_pl32g_status_reg_tx_precoding_on),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_port_force_off_support_part_lanes_rxei_exit                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_port_force_off_support_part_lanes_rxei_exit),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_port_link_ctrl_off_fast_link_mode                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_port_link_ctrl_off_fast_link_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_root_control_root_capabilities_reg_pcie_cap_crs_sw_visibility),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw                                 ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_1_sn_ser_num_reg_1_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw                                 ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_ser_num_reg_dw_2_sn_ser_num_reg_2_dw)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_pci_msix_cap_id_next_ctrl_reg_pci_msix_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_shadow_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_attention_indicator_button),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_electromech_interlock),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_capable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_hot_plug_surprise),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_mrl_sensor),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_no_cmd_cpl_support),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_phy_slot_num),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_controller),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_power_indicator),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_scale),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_slot_capabilities_reg_pcie_cap_slot_power_limit_value),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_rx_preset_hint1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_dsp_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_rx_preset_hint1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_0ch_reg_usp_tx_preset1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_rx_preset_hint3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_dsp_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_rx_preset_hint3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset2),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_spcie_cap_off_10h_reg_usp_tx_preset3),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_dev_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_subsystem_id_subsystem_vendor_id_reg_subsys_vendor_id),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_int_vec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_loc_1),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_cap_st_table_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_device_spec                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pf0_tph_req_cap_reg_reg_tph_req_device_spec),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pfvf_sel_vsec_enable_attr                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_pfvf_sel_vsec_enable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_phy_rxelecidle_k_rxelecidle_disable_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_phy_rxelecidle_k_rxelecidle_disable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_phy_rxtermination_k_rxtermination_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_phy_rxtermination_k_rxtermination_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_reset_ctrl1_k_clrhip_not_rst_sticky_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_err_en_correct_err_en_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_err_en_correct_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_err_en_fatal_err_en_attr                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_err_en_fatal_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_err_en_nonfatal_err_en_attr                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_err_en_nonfatal_err_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_aer_rc_err_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_bw_mgt_int_en_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_bw_mgt_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_auto_bw_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_eq_req_int_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_link_eq_req_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_pme_int_en_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_cfg_pme_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_int_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_int_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_pme_en_attr                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_hp_pme_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_inta_en_attr                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_inta_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_intb_en_attr                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_intb_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_intc_en_attr                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_intc_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_intd_en_attr                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_rp_irq_en_intd_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_dlycnt_attr                                       ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_dlycnt_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_mode_attr                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_stagger_control_k_stag_mode_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_dllp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_bad_tlp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_corrected_internal_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_dl_protocol_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_ecrc_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_fc_protocol_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_mlf_tlp_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_rcvr_overflow_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_number_rollover_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_replay_timer_timeout_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_surprise_down_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_en_k_cfg_uncor_internal_err_sts_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_dllp_err_sts_attr                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_dllp_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_tlp_err_sts_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_bad_tlp_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_corrected_internal_err_sts_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_corrected_internal_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_dl_protocol_err_sts_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_dl_protocol_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_ecrc_err_sts_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_ecrc_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_fc_protocol_err_sts_attr                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_fc_protocol_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_mlf_tlp_err_sts_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_mlf_tlp_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_err_sts_attr                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_overflow_err_sts_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_rcvr_overflow_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_number_rollover_err_sts_attr                      ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_number_rollover_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_timer_timeout_err_sts_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_replay_timer_timeout_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_surprise_down_err_sts_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_surprise_down_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_uncor_internal_err_sts_attr                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tlb_err_sts_cfg_uncor_internal_err_sts_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tx_common_mode_k_txcommonmode_disable_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_tx_common_mode_k_txcommonmode_disable_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_10_k_pf0_virtio_offset_cfg3_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_11_k_pf0_virtio_offset_cfg3_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_12_k_pf0_virtio_offset_cfg3_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_14_k_pf0_virtio_offset_cfg4_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_15_k_pf0_virtio_offset_cfg4_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_16_k_pf0_virtio_offset_cfg4_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_18_k_pf0_virtio_offset_cfg5_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_19_k_pf0_virtio_offset_cfg5_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_1_k_pf0_virtio_offset_cfg1_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr                       ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_20_k_pf0_virtio_offset_cfg5_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr                         ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_21_k_pf0_virtio_offset_cfg5_cfg_data_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_2_k_pf0_virtio_offset_cfg1_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_3_k_pf0_virtio_offset_cfg1_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_5_k_pf0_virtio_offset_cfg2_cap_bar_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_6_k_pf0_virtio_offset_cfg2_cap_offset_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr                        ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_7_k_pf0_virtio_offset_cfg2_cap_length_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr             ( str_2_bin(hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_8_k_pf0_virtio_offset_cfg2_notify_off_multiplier_attr)),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cfg_update_en_attr                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cfg_update_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cii_en_attr                                            ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_cii_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtio_cii_ctrl_k_pfdata_vf_virtio_en_attr),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_cvp_mode                                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_cvp_mode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_drop_vendor0_msg                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_drop_vendor0_msg),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_drop_vendor1_msg                                                 ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_drop_vendor1_msg),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_ep_native                                                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_ep_native),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_maxpayload_size                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_maxpayload_size),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_num_of_lanes                                                     ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_num_of_lanes),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_acs_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_ats_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_bar1_mask_bit0                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_bar1_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_bar3_mask_bit0                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_bar3_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_bar5_mask_bit0                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_bar5_mask_bit0),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_dlink_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_dlink_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_acs_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_acs_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_ats_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_ats_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_msix_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_msix_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_tph_cap_enable                                          ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_exvf_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_io_decode                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_io_decode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_ltr_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_ltr_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_msi_enable                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_msi_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_msix_enable                                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_msix_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_pasid_cap_enable                                             ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_pasid_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_prefetch_decode                                              ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_prefetch_decode),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_prs_ext_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_prs_ext_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_ras_des_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_ras_des_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_sn_cap_enable                                                ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_sn_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_tph_cap_enable                                               ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_tph_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_user_vsec_cap_enable                                         ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_user_vsec_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_dev_specific_conf_en                                  ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_dev_specific_conf_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_en                                                    ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_virtio_en),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_vsecras_cap_enable                                           ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_pf0_vsecras_cap_enable),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_ptm_autoupdate                                                   ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_ptm_autoupdate),
   .hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr                        ( hssi_ctr_u_pcie_top_rnr_pcie_par_p2_inst_rnr_pcie_ip4_inst_virtual_tlp_bypass_en_dwc_ctrl0_k_ecrc_strip_attr),
   .hssi_ctr_u_pcie_top_sim_mode                                                                                                        ( hssi_ctr_u_pcie_top_sim_mode),
   .hssi_ctr_u_pcie_top_sup_mode                                                                                                        ( hssi_ctr_u_pcie_top_sup_mode),
   .hssi_ctr_u_pcie_top_virtual_dmwr_support                                                                                            ( hssi_ctr_u_pcie_top_virtual_dmwr_support),
   .hssi_ctr_u_pcie_top_virtual_l1sub_support                                                                                           ( hssi_ctr_u_pcie_top_virtual_l1sub_support),
   .hssi_ctr_u_phy_top_pcie_capable_octet0                                                                                              ( hssi_ctr_u_phy_top_pcie_capable_octet0),
   .hssi_ctr_u_phy_top_pcie_capable_octet1                                                                                              ( hssi_ctr_u_phy_top_pcie_capable_octet1),
   .hssi_ctr_u_phy_top_u_phy_octet0_powerdown_mode                                                                                      ( hssi_ctr_u_phy_top_u_phy_octet0_powerdown_mode),
   .hssi_ctr_u_phy_top_u_phy_octet1_powerdown_mode                                                                                      ( hssi_ctr_u_phy_top_u_phy_octet1_powerdown_mode),
   .hssi_ctr_u_rnr_aibaux_top_wrp_powerdown_mode                                                                                        ( hssi_ctr_u_rnr_aibaux_top_wrp_powerdown_mode),
   .hssi_ctr_silicon_rev                                                                                                                ( hssi_ctr_silicon_rev)
)
u_rtile_mdx1 (
/* input         */ .refclk0                                                         (refclk0),
/* input         */ .refclk1                                                         (refclk1),
/* output        */ .coreclkout_hip                                                  (coreclkout_hip),
/* output        */ .side_clk                                                        (side_clk),
/* input         */ .pin_perst_n                                                     (pin_perst_n),
/* input         */ .ninit_done                                                      (ninit_done),
/* output        */ .p0_pin_perst_n                                                  (p0_pin_perst_n),
/* output        */ .p1_pin_perst_n                                                  (p1_pin_perst_n),
/* output        */ .p2_pin_perst_n                                                  (p2_pin_perst_n),
/* output        */ .p3_pin_perst_n                                                  (p3_pin_perst_n),
/* output        */ .cxl_pin_perst_n                                                 (cxl_pin_perst_n),
/* output        */ .p0_reset_status_n                                               ( ),
/* input         */ .p0_pld_warm_rst_rdy_i                                           (p0_pld_warm_rst_rdy_i),
/* output        */ .p0_pld_link_req_rst_o                                           (),
/* output        */ .p1_reset_status_n                                               ( ),
/* input         */ .p1_pld_warm_rst_rdy_i                                           (p1_pld_warm_rst_rdy_i),
/* output        */ .p1_pld_link_req_rst_o                                           (p1_pld_link_req_rst_o),
/* input         */ .p2_pld_warm_rst_rdy_i                                           (p2_pld_warm_rst_rdy_i),
/* output        */ .p2_pld_link_req_rst_o                                           (p2_pld_link_req_rst_o),
/* output        */ .p2_reset_status_n                                               ( ),
/* input         */ .p3_pld_warm_rst_rdy_i                                           (p3_pld_warm_rst_rdy_i),
/* output        */ .p3_pld_link_req_rst_o                                           (p3_pld_link_req_rst_o),
/* output        */ .p3_reset_status_n                                               ( ),
/* input         */ .cxl_pld_warm_rst_rdy_i                                          (p0_pld_warm_rst_rdy_i),
/* output        */ .cxl_pld_link_req_rst_o                                          (p0_pld_link_req_rst_o),
/* output        */ .cxl_reset_status_n                                              (cxl_reset_status_n),
/* output        */ .cxl_pld_core_cold_rst_n                                         (p0_pld_core_cold_rst_n),
/* output        */ .cxl_pld_core_warm_rst_n                                         (p0_pld_core_warm_rst_n),
/* input         */ .p0_app_rst_n                                                    (p0_app_rst_n),
/* input         */ .p1_app_rst_n                                                    (p1_app_rst_n),
/* input         */ .p2_app_rst_n                                                    (p2_app_rst_n),
/* input         */ .p3_app_rst_n                                                    (p3_app_rst_n),
/* input         */ .cxl_app_rst_n                                                   (cxl_app_rst_n),
/* input         */ .cxl_pll_locked_i                                                (cxl_pll_locked_i),
/* input         */ .i_clk                                                           (i_clk),
/* input         */ .i_rst_n                                                         (i_rst_n),
/* input         */ .i_rx_dsk_clear                                                  (i_rx_dsk_clear),
/* input         */ .i_tx_dsk_clear                                                  (i_tx_dsk_clear),
/* output        */ .rx_deskew_valid                                                 (rx_deskew_valid),
/* output        */ .rx_deskew_done                                                  (rx_deskew_done),
/* output        */ .rx_deskew_lock_err                                              (rx_deskew_lock_err),
/* output [31:0] */ .rx_dsk_monitor_err                                              (rx_dsk_monitor_err),
/* output        */ .o_ptm_clk_updated                                               (o_ptm_clk_updated),
/* output        */ .o_ptm_context_valid                                             (o_ptm_context_valid),
/* output        */ .o_ptm_local_clock                                               (o_ptm_local_clock),
/* input         */ .i_ptm_manual_update                                             (i_ptm_manual_update),
/* output        */ .rx_st0_dvalid                                                   (rx_st0_dvalid),
/* output        */ .rx_st1_dvalid                                                   (rx_st1_dvalid),
/* output        */ .rx_st2_dvalid                                                   (rx_st2_dvalid),
/* output        */ .rx_st3_dvalid                                                   (rx_st3_dvalid),
/* output        */ .rx_st0_sop                                                      (rx_st0_sop),
/* output        */ .rx_st1_sop                                                      (rx_st1_sop),
/* output        */ .rx_st2_sop                                                      (rx_st2_sop),
/* output        */ .rx_st3_sop                                                      (rx_st3_sop),
/* output        */ .rx_st0_eop                                                      (rx_st0_eop),
/* output        */ .rx_st1_eop                                                      (rx_st1_eop),
/* output        */ .rx_st2_eop                                                      (rx_st2_eop),
/* output        */ .rx_st3_eop                                                      (rx_st3_eop),
/* output        */ .rx_st0_passthrough                                              (rx_st0_passthrough),
/* output        */ .rx_st1_passthrough                                              (rx_st1_passthrough),
/* output        */ .rx_st2_passthrough                                              (rx_st2_passthrough),
/* output        */ .rx_st3_passthrough                                              (rx_st3_passthrough),
/* output [255:0]*/ .rx_st0_data                                                     (rx_st0_data),
/* output [255:0]*/ .rx_st1_data                                                     (rx_st1_data),
/* output [255:0]*/ .rx_st2_data                                                     (rx_st2_data),
/* output [255:0]*/ .rx_st3_data                                                     (rx_st3_data),
/* output [7:0]  */ .rx_st0_data_parity                                              (rx_st0_data_parity),
/* output [7:0]  */ .rx_st1_data_parity                                              (rx_st1_data_parity),
/* output [7:0]  */ .rx_st2_data_parity                                              (rx_st2_data_parity),
/* output [7:0]  */ .rx_st3_data_parity                                              (rx_st3_data_parity),
/* output [127:0]*/ .rx_st0_hdr                                                      (rx_st0_hdr),
/* output [127:0]*/ .rx_st1_hdr                                                      (rx_st1_hdr),
/* output [127:0]*/ .rx_st2_hdr                                                      (rx_st2_hdr),
/* output [127:0]*/ .rx_st3_hdr                                                      (rx_st3_hdr),
/* output [3:0]  */ .rx_st0_hdr_parity                                               (rx_st0_hdr_parity),
/* output [3:0]  */ .rx_st1_hdr_parity                                               (rx_st1_hdr_parity),
/* output [3:0]  */ .rx_st2_hdr_parity                                               (rx_st2_hdr_parity),
/* output [3:0]  */ .rx_st3_hdr_parity                                               (rx_st3_hdr_parity),
/* output        */ .rx_st0_hvalid                                                   (rx_st0_hvalid),
/* output        */ .rx_st1_hvalid                                                   (rx_st1_hvalid),
/* output        */ .rx_st2_hvalid                                                   (rx_st2_hvalid),
/* output        */ .rx_st3_hvalid                                                   (rx_st3_hvalid),
/* output [31:0] */ .rx_st0_prefix                                                   (rx_st0_prefix),
/* output [31:0] */ .rx_st1_prefix                                                   (rx_st1_prefix),
/* output [31:0] */ .rx_st2_prefix                                                   (rx_st2_prefix),
/* output [31:0] */ .rx_st3_prefix                                                   (rx_st3_prefix),
/* output        */ .rx_st0_prefix_parity                                            (rx_st0_prefix_parity),
/* output        */ .rx_st1_prefix_parity                                            (rx_st1_prefix_parity),
/* output        */ .rx_st2_prefix_parity                                            (rx_st2_prefix_parity),
/* output        */ .rx_st3_prefix_parity                                            (rx_st3_prefix_parity),
/* output [11:0] */ .rx_st0_rssai_prefix                                             (rx_st0_rssai_prefix),
/* output [11:0] */ .rx_st1_rssai_prefix                                             (rx_st1_rssai_prefix),
/* output [11:0] */ .rx_st2_rssai_prefix                                             (rx_st2_rssai_prefix),
/* output [11:0] */ .rx_st3_rssai_prefix                                             (rx_st3_rssai_prefix),
/* output        */ .rx_st0_rssai_prefix_parity                                      (rx_st0_rssai_prefix_parity),
/* output        */ .rx_st1_rssai_prefix_parity                                      (rx_st1_rssai_prefix_parity),
/* output        */ .rx_st2_rssai_prefix_parity                                      (rx_st2_rssai_prefix_parity),
/* output        */ .rx_st3_rssai_prefix_parity                                      (rx_st3_rssai_prefix_parity),
/* output [1:0]  */ .rx_st0_pvalid                                                   (rx_st0_pvalid),
/* output [1:0]  */ .rx_st1_pvalid                                                   (rx_st1_pvalid),
/* output [1:0]  */ .rx_st2_pvalid                                                   (rx_st2_pvalid),
/* output [1:0]  */ .rx_st3_pvalid                                                   (rx_st3_pvalid),
/* output [2:0]  */ .rx_st0_bar                                                      (rx_st0_bar),
/* output [2:0]  */ .rx_st1_bar                                                      (rx_st1_bar),
/* output [2:0]  */ .rx_st2_bar                                                      (rx_st2_bar),
/* output [2:0]  */ .rx_st3_bar                                                      (rx_st3_bar),
/* output        */ .rx_st0_vfactive                                                 (rx_st0_vfactive),
/* output        */ .rx_st1_vfactive                                                 (rx_st1_vfactive),
/* output        */ .rx_st2_vfactive                                                 (rx_st2_vfactive),
/* output        */ .rx_st3_vfactive                                                 (rx_st3_vfactive),
/* output [10:0] */ .rx_st0_vfnum                                                    (rx_st0_vfnum),
/* output [10:0] */ .rx_st1_vfnum                                                    (rx_st1_vfnum),
/* output [10:0] */ .rx_st2_vfnum                                                    (rx_st2_vfnum),
/* output [10:0] */ .rx_st3_vfnum                                                    (rx_st3_vfnum),
/* output [2:0]  */ .rx_st0_pfnum                                                    (rx_st0_pfnum),
/* output [2:0]  */ .rx_st1_pfnum                                                    (rx_st1_pfnum),
/* output [2:0]  */ .rx_st2_pfnum                                                    (rx_st2_pfnum),
/* output [2:0]  */ .rx_st3_pfnum                                                    (rx_st3_pfnum),
/* output        */ .rx_st0_chnum                                                    (rx_st0_chnum),
/* output        */ .rx_st1_chnum                                                    (rx_st1_chnum),
/* output        */ .rx_st2_chnum                                                    (rx_st2_chnum),
/* output        */ .rx_st3_chnum                                                    (rx_st3_chnum),
/* output        */ .rx_st0_misc_parity                                              (rx_st0_misc_parity),
/* output        */ .rx_st1_misc_parity                                              (rx_st1_misc_parity),
/* output        */ .rx_st2_misc_parity                                              (rx_st2_misc_parity),
/* output        */ .rx_st3_misc_parity                                              (rx_st3_misc_parity),
/* output [2:0]  */ .rx_st0_empty                                                    (rx_st0_empty),
/* output [2:0]  */ .rx_st1_empty                                                    (rx_st1_empty),
/* output [2:0]  */ .rx_st2_empty                                                    (rx_st2_empty),
/* output [2:0]  */ .rx_st3_empty                                                    (rx_st3_empty),
/* input  [2:0]  */ .rx_st_Hcrdt_update                                              (rx_st_Hcrdt_update),
/* input  [2:0]  */ .rx_st_Hcrdt_ch                                                  (rx_st_Hcrdt_ch),
/* input  [5:0]  */ .rx_st_Hcrdt_update_cnt                                          (rx_st_Hcrdt_update_cnt),
/* input  [2:0]  */ .rx_st_Hcrdt_init                                                (rx_st_Hcrdt_init),
/* output [2:0]  */ .rx_st_Hcrdt_init_ack                                            (rx_st_Hcrdt_init_ack),
/* input  [2:0]  */ .rx_st_Dcrdt_update                                              (rx_st_Dcrdt_update),
/* input  [2:0]  */ .rx_st_Dcrdt_ch                                                  (rx_st_Dcrdt_ch),
/* input  [11:0] */ .rx_st_Dcrdt_update_cnt                                          (rx_st_Dcrdt_update_cnt),
/* input  [2:0]  */ .rx_st_Dcrdt_init                                                (rx_st_Dcrdt_init),
/* output [2:0]  */ .rx_st_Dcrdt_init_ack                                            (rx_st_Dcrdt_init_ack),
/* output        */ .tx_st_ready                                                     (tx_st_ready),
/* input         */ .tx_st0_dvalid                                                   (tx_st0_dvalid),
/* input         */ .tx_st1_dvalid                                                   (tx_st1_dvalid),
/* input         */ .tx_st2_dvalid                                                   (tx_st2_dvalid),
/* input         */ .tx_st3_dvalid                                                   (tx_st3_dvalid),
/* input         */ .tx_st0_sop                                                      (tx_st0_sop),
/* input         */ .tx_st1_sop                                                      (tx_st1_sop),
/* input         */ .tx_st2_sop                                                      (tx_st2_sop),
/* input         */ .tx_st3_sop                                                      (tx_st3_sop),
/* input         */ .tx_st0_eop                                                      (tx_st0_eop),
/* input         */ .tx_st1_eop                                                      (tx_st1_eop),
/* input         */ .tx_st2_eop                                                      (tx_st2_eop),
/* input         */ .tx_st3_eop                                                      (tx_st3_eop),
/* input         */ .tx_st0_passthrough                                              (tx_st0_passthrough),
/* input         */ .tx_st1_passthrough                                              (tx_st1_passthrough),
/* input         */ .tx_st2_passthrough                                              (tx_st2_passthrough),
/* input         */ .tx_st3_passthrough                                              (tx_st3_passthrough),
/* input  [255:0]*/ .tx_st0_data                                                     (tx_st0_data),
/* input  [255:0]*/ .tx_st1_data                                                     (tx_st1_data),
/* input  [255:0]*/ .tx_st2_data                                                     (tx_st2_data),
/* input  [255:0]*/ .tx_st3_data                                                     (tx_st3_data),
/* input  [7:0]  */ .tx_st0_data_parity                                              (tx_st0_data_parity),
/* input  [7:0]  */ .tx_st1_data_parity                                              (tx_st1_data_parity),
/* input  [7:0]  */ .tx_st2_data_parity                                              (tx_st2_data_parity),
/* input  [7:0]  */ .tx_st3_data_parity                                              (tx_st3_data_parity),
/* input  [127:0]*/ .tx_st0_hdr                                                      (tx_st0_hdr),
/* input  [127:0]*/ .tx_st1_hdr                                                      (tx_st1_hdr),
/* input  [127:0]*/ .tx_st2_hdr                                                      (tx_st2_hdr),
/* input  [127:0]*/ .tx_st3_hdr                                                      (tx_st3_hdr),
/* input  [3:0]  */ .tx_st0_hdr_parity                                               (tx_st0_hdr_parity),
/* input  [3:0]  */ .tx_st1_hdr_parity                                               (tx_st1_hdr_parity),
/* input  [3:0]  */ .tx_st2_hdr_parity                                               (tx_st2_hdr_parity),
/* input  [3:0]  */ .tx_st3_hdr_parity                                               (tx_st3_hdr_parity),
/* input         */ .tx_st0_hvalid                                                   (tx_st0_hvalid),
/* input         */ .tx_st1_hvalid                                                   (tx_st1_hvalid),
/* input         */ .tx_st2_hvalid                                                   (tx_st2_hvalid),
/* input         */ .tx_st3_hvalid                                                   (tx_st3_hvalid),
/* input  [31:0] */ .tx_st0_prefix                                                   (tx_st0_prefix),
/* input  [31:0] */ .tx_st1_prefix                                                   (tx_st1_prefix),
/* input  [31:0] */ .tx_st2_prefix                                                   (tx_st2_prefix),
/* input  [31:0] */ .tx_st3_prefix                                                   (tx_st3_prefix),
/* input         */ .tx_st0_prefix_parity                                            (tx_st0_prefix_parity),
/* input         */ .tx_st1_prefix_parity                                            (tx_st1_prefix_parity),
/* input         */ .tx_st2_prefix_parity                                            (tx_st2_prefix_parity),
/* input         */ .tx_st3_prefix_parity                                            (tx_st3_prefix_parity),
/* input  [11:0] */ .tx_st0_rssai_prefix                                             (tx_st0_rssai_prefix),
/* input  [11:0] */ .tx_st1_rssai_prefix                                             (tx_st1_rssai_prefix),
/* input  [11:0] */ .tx_st2_rssai_prefix                                             (tx_st2_rssai_prefix),
/* input  [11:0] */ .tx_st3_rssai_prefix                                             (tx_st3_rssai_prefix),
/* input         */ .tx_st0_rssai_prefix_parity                                      (tx_st0_rssai_prefix_parity),
/* input         */ .tx_st1_rssai_prefix_parity                                      (tx_st1_rssai_prefix_parity),
/* input         */ .tx_st2_rssai_prefix_parity                                      (tx_st2_rssai_prefix_parity),
/* input         */ .tx_st3_rssai_prefix_parity                                      (tx_st3_rssai_prefix_parity),
/* input  [1:0]  */ .tx_st0_pvalid                                                   (tx_st0_pvalid),
/* input  [1:0]  */ .tx_st1_pvalid                                                   (tx_st1_pvalid),
/* input  [1:0]  */ .tx_st2_pvalid                                                   (tx_st2_pvalid),
/* input  [1:0]  */ .tx_st3_pvalid                                                   (tx_st3_pvalid),
/* input  [2:0]  */ .tx_st0_empty                                                    (tx_st0_empty),
/* input  [2:0]  */ .tx_st1_empty                                                    (tx_st1_empty),
/* input  [2:0]  */ .tx_st2_empty                                                    (tx_st2_empty),
/* input  [2:0]  */ .tx_st3_empty                                                    (tx_st3_empty),
/* output [2:0]  */ .tx_st_Hcrdt_update                                              (tx_st_Hcrdt_update),
/* output [2:0]  */ .tx_st_Hcrdt_vc                                                  (tx_st_Hcrdt_vc),
/* output [5:0]  */ .tx_st_Hcrdt_update_cnt                                          (tx_st_Hcrdt_update_cnt),
/* output [2:0]  */ .tx_st_Hcrdt_init                                                (tx_st_Hcrdt_init),
/* input  [2:0]  */ .tx_st_Hcrdt_init_ack                                            (tx_st_Hcrdt_init_ack),
/* output [2:0]  */ .tx_st_Dcrdt_update                                              (tx_st_Dcrdt_update),
/* output [2:0]  */ .tx_st_Dcrdt_vc                                                  (tx_st_Dcrdt_vc),
/* output [11:0] */ .tx_st_Dcrdt_update_cnt                                          (tx_st_Dcrdt_update_cnt),
/* output [2:0]  */ .tx_st_Dcrdt_init                                                (tx_st_Dcrdt_init),
/* input  [2:0]  */ .tx_st_Dcrdt_init_ack                                            (tx_st_Dcrdt_init_ack),
/* output        */ .mnpput                                                          (p0_mnpput_o),
/* output        */ .mpcput                                                          (p0_mpcput_o),
/* input         */ .mnpcup                                                          (p0_mnpcup_i),
/* input         */ .mpccup                                                          (p0_mpccup_i),
/* output        */ .meom                                                            (p0_meom_o),
/* output [15:0] */ .mpayload                                                        (p0_mpayload_o),
/* output        */ .mparity                                                         (p0_mparity_o),
/* input  [2:0]  */ .side_ism_fabric                                                 (p0_side_ism_fabric_i),
/* input         */ .tnpput                                                          (p0_tnpput_i),
/* input         */ .tpcput                                                          (p0_tpcput_i),
/* output        */ .tnpcup                                                          (p0_tnpcup_o),
/* output        */ .tpccup                                                          (p0_tpccup_o),
/* input         */ .teom                                                            (p0_teom_i),
/* input  [15:0] */ .tpayload                                                        (p0_tpayload_i),
/* input         */ .tparity                                                         (p0_tparity_i),
/* output [2:0]  */ .side_ism_agent                                                  (p0_side_ism_agent_o),
/* output        */ .cxl_cache_mem_rx_frame0                                         (cxl_cache_mem_rx_frame0),
/* output        */ .cxl_cache_mem_rx_frame1                                         (cxl_cache_mem_rx_frame1),
/* input         */ .cxl_mem_s2m_tx_frame0                                           (cxl_mem_s2m_tx_frame0),
/* input         */ .cxl_mem_s2m_tx_frame0_valid                                     (cxl_mem_s2m_tx_frame0_valid),
/* output        */ .cxl_mem_s2m_tx_frame0_ready                                     (cxl_mem_s2m_tx_frame0_ready),
/* input         */ .cxl_mem_s2m_tx_frame1                                           (cxl_mem_s2m_tx_frame1),
/* input         */ .cxl_mem_s2m_tx_frame1_valid                                     (cxl_mem_s2m_tx_frame1_valid),
/* output        */ .cxl_mem_s2m_tx_frame1_ready                                     (cxl_mem_s2m_tx_frame1_ready),
/* input         */ .cxl_d2h_req_frame0                                              (cxl_d2h_req_frame0),
/* input  [3:0]  */ .cxl_d2h_req_frame0_valid                                        (cxl_d2h_req_frame0_valid),
/* output [3:0]  */ .cxl_d2h_req_frame0_ready                                        (cxl_d2h_req_frame0_ready),
/* input         */ .cxl_d2h_req_frame1                                              (cxl_d2h_req_frame1),
/* input  [3:0]  */ .cxl_d2h_req_frame1_valid                                        (cxl_d2h_req_frame1_valid),
/* output [3:0]  */ .cxl_d2h_req_frame1_ready                                        (cxl_d2h_req_frame1_ready),
/* input         */ .cxl_d2h_rsp_frame0                                              (cxl_d2h_rsp_frame0),
/* input  [1:0]  */ .cxl_d2h_rsp_frame0_valid                                        (cxl_d2h_rsp_frame0_valid),
/* output [1:0]  */ .cxl_d2h_rsp_frame0_ready                                        (cxl_d2h_rsp_frame0_ready),
/* input         */ .cxl_d2h_rsp_frame1                                              (cxl_d2h_rsp_frame1),
/* input  [1:0]  */ .cxl_d2h_rsp_frame1_valid                                        (cxl_d2h_rsp_frame1_valid),
/* output [1:0]  */ .cxl_d2h_rsp_frame1_ready                                        (cxl_d2h_rsp_frame1_ready),
/* input         */ .cxl_d2h_data_frame0                                             (cxl_d2h_data_frame0),
/* input         */ .cxl_d2h_data_frame0_valid                                       (cxl_d2h_data_frame0_valid),
/* output        */ .cxl_d2h_data_frame0_ready                                       (cxl_d2h_data_frame0_ready),
/* input         */ .cxl_d2h_data_frame1                                             (cxl_d2h_data_frame1),
/* input         */ .cxl_d2h_data_frame1_valid                                       (cxl_d2h_data_frame1_valid),
/* output        */ .cxl_d2h_data_frame1_ready                                       (cxl_d2h_data_frame1_ready),
/* output        */ .o_D2H_Data0_CrdRtn                                              (o_D2H_Data0_CrdRtn),
/* output        */ .o_D2H_Req_CrdRtn                                                (o_D2H_Req_CrdRtn),
/* output        */ .o_D2H_Rsp_CrdRtn                                                (o_D2H_Rsp_CrdRtn),
/* output        */ .o_S2M_DRS0_CrdRtn                                               (o_S2M_DRS0_CrdRtn),
/* output        */ .o_S2M_DRS1_CrdRtn                                               (o_S2M_DRS1_CrdRtn),
/* output        */ .o_S2M_NDR_CrdRtn                                                (o_S2M_NDR_CrdRtn),
/* output        */ .o_D2HPushWrCrdRtn                                               (o_D2HPushWrCrdRtn),
/* input         */ .i_H2D_Data0_CrdRtn                                              (i_H2D_Data0_CrdRtn),
/* input         */ .i_H2D_Data1_CrdRtn                                              (i_H2D_Data1_CrdRtn),
/* input         */ .i_H2D_Req_CrdRtn                                                (i_H2D_Req_CrdRtn),
/* input         */ .i_H2D_Rsp_CrdRtn                                                (i_H2D_Rsp_CrdRtn),
/* input         */ .i_M2S_Req_CrdRtn                                                (i_M2S_Req_CrdRtn),
/* input         */ .i_M2S_RwD0_CrdRtn                                               (i_M2S_RwD0_CrdRtn),
/* input         */ .i_M2S_RwD1_CrdRtn                                               (i_M2S_RwD1_CrdRtn),
		   .i_H2D_Rsp_CrdRtn_fr0       (i_H2D_Rsp_CrdRtn_fr0   ),
		   .i_H2D_Rsp_CrdRtn_fr1       (i_H2D_Rsp_CrdRtn_fr1   ),
		   .i_H2D_Req_CrdRtn_fr0       (i_H2D_Req_CrdRtn_fr0   ),
		   .i_H2D_Req_CrdRtn_fr1       (i_H2D_Req_CrdRtn_fr1   ),
		   .i_H2D_Data0_CrdRtn_fr0     (i_H2D_Data0_CrdRtn_fr0 ),
		   .i_H2D_Data0_CrdRtn_fr1     (i_H2D_Data0_CrdRtn_fr1 ),
		   .i_M2S_RwD0_CrdRtn_fr0      (i_M2S_RwD0_CrdRtn_fr0  ),
		   .i_M2S_RwD0_CrdRtn_fr1      (i_M2S_RwD0_CrdRtn_fr1  ),
		   .i_M2S_Req_CrdRtn_fr0       (i_M2S_Req_CrdRtn_fr0   ),
		   .i_M2S_Req_CrdRtn_fr1       (i_M2S_Req_CrdRtn_fr1   ),

/* output        */ .o_M2S_viral                                                     (cxl_mem_m2s_viral_o    ),
/* output        */ .o_H2D_viral                                                     (cxl_cache_h2d_viral_o  ),
/* input         */ .i_S2M_viral                                                     (cxl_mem_s2m_viral_i    ),
/* input         */ .i_D2H_viral                                                     (cxl_cache_d2h_viral_i  ),
/* output [3:0]  */ .o_ial_ch18_ext_fsr                                              (o_ial_ch18_ext_fsr),
/* output [7:0]  */ .o_ial_ch18_ext_ssr                                              (o_ial_ch18_ext_ssr),
/* output [2:0]  */ .o_ial_ch18_fsr                                                  (o_ial_ch18_fsr),
/* output [64:0] */ .o_ial_ch18_ssr                                                  (o_ial_ch18_ssr),
/* output [3:0]  */ .o_ial_ch19_ext_fsr                                              (o_ial_ch19_ext_fsr),
/* output [7:0]  */ .o_ial_ch19_ext_ssr                                              (o_ial_ch19_ext_ssr),
/* output [2:0]  */ .o_ial_ch19_fsr                                                  (o_ial_ch19_fsr),
/* output [64:0] */ .o_ial_ch19_ssr                                                  (o_ial_ch19_ssr),
/* output [5:0]  */ .o_ial_ch1_async_direct                                          (o_ial_ch1_async_direct),
/* output [3:0]  */ .o_ial_ch20_ext_fsr                                              (o_ial_ch20_ext_fsr),
/* output [7:0]  */ .o_ial_ch20_ext_ssr                                              (o_ial_ch20_ext_ssr),
/* output [2:0]  */ .o_ial_ch20_fsr                                                  (o_ial_ch20_fsr),
/* output [64:0] */ .o_ial_ch20_ssr                                                  (o_ial_ch20_ssr),
/* output [3:0]  */ .o_ial_ch21_ext_fsr                                              (o_ial_ch21_ext_fsr),
/* output [7:0]  */ .o_ial_ch21_ext_ssr                                              (o_ial_ch21_ext_ssr),
/* output [2:0]  */ .o_ial_ch21_fsr                                                  (o_ial_ch21_fsr),
/* output [64:0] */ .o_ial_ch21_ssr                                                  (o_ial_ch21_ssr),
/* output [3:0]  */ .o_ial_ch22_ext_fsr                                              (o_ial_ch22_ext_fsr),
/* output [7:0]  */ .o_ial_ch22_ext_ssr                                              (o_ial_ch22_ext_ssr),
/* output [2:0]  */ .o_ial_ch22_fsr                                                  (o_ial_ch22_fsr),
/* output [64:0] */ .o_ial_ch22_ssr                                                  (o_ial_ch22_ssr),
/* output [3:0]  */ .o_ial_ch23_ext_fsr                                              (o_ial_ch23_ext_fsr),
/* output [7:0]  */ .o_ial_ch23_ext_ssr                                              (o_ial_ch23_ext_ssr),
/* output [2:0]  */ .o_ial_ch23_fsr                                                  (o_ial_ch23_fsr),
/* output [64:0] */ .o_ial_ch23_ssr                                                  (o_ial_ch23_ssr),
/* output [5:0]  */ .o_ial_ch2_async_direct                                          (o_ial_ch2_async_direct),
/* output [5:0]  */ .o_ial_ch3_async_direct                                          (o_ial_ch3_async_direct),
/* input  [3:0]  */ .i_ial_ch19_ext_fsr                                              (i_ial_ch19_ext_fsr),
/* input  [39:0] */ .i_ial_ch19_ext_ssr                                              (i_ial_ch19_ext_ssr),
/* input  [2:0]  */ .i_ial_ch19_fsr                                                  (i_ial_ch19_fsr),
/* input  [60:0] */ .i_ial_ch19_ssr                                                  (i_ial_ch19_ssr),
/* input  [3:0]  */ .i_ial_ch20_ext_fsr                                              (i_ial_ch20_ext_fsr),
/* input  [39:0] */ .i_ial_ch20_ext_ssr                                              (i_ial_ch20_ext_ssr),
/* input  [2:0]  */ .i_ial_ch20_fsr                                                  (i_ial_ch20_fsr),
/* input  [60:0] */ .i_ial_ch20_ssr                                                  (i_ial_ch20_ssr),
/* input  [3:0]  */ .i_ial_ch21_ext_fsr                                              (i_ial_ch21_ext_fsr),
/* input  [39:0] */ .i_ial_ch21_ext_ssr                                              (i_ial_ch21_ext_ssr),
/* input  [2:0]  */ .i_ial_ch21_fsr                                                  (i_ial_ch21_fsr),
/* input  [60:0] */ .i_ial_ch21_ssr                                                  (i_ial_ch21_ssr),
/* input  [7:0]  */ .i_ial_ch22_async_direct                                         (i_ial_ch22_async_direct),
/* input  [3:0]  */ .i_ial_ch22_ext_fsr                                              (i_ial_ch22_ext_fsr),
/* input  [39:0] */ .i_ial_ch22_ext_ssr                                              (i_ial_ch22_ext_ssr),
/* input  [2:0]  */ .i_ial_ch22_fsr                                                  (i_ial_ch22_fsr),
/* input  [60:0] */ .i_ial_ch22_ssr                                                  (i_ial_ch22_ssr),
/* input  [7:0]  */ .i_ial_ch23_async_direct                                         (i_ial_ch23_async_direct),
/* input  [3:0]  */ .i_ial_ch23_ext_fsr                                              (i_ial_ch23_ext_fsr),
/* input  [39:0] */ .i_ial_ch23_ext_ssr                                              (i_ial_ch23_ext_ssr),
/* input  [2:0]  */ .i_ial_ch23_fsr                                                  (i_ial_ch23_fsr),
/* input  [60:0] */ .i_ial_ch23_ssr                                                  (i_ial_ch23_ssr),
/* output [5:0]  */ .o_ch0_async_direct_aib2pld                                      (o_ch0_async_direct_aib2pld),
/* output [5:0]  */ .o_ch1_async_direct_aib2pld                                      (o_ch1_async_direct_aib2pld),
/* output [5:0]  */ .o_ch2_async_direct_aib2pld                                      (o_ch2_async_direct_aib2pld),
/* output [5:0]  */ .o_ch3_async_direct_aib2pld                                      (o_ch3_async_direct_aib2pld),
/* output [5:0]  */ .o_ch4_async_direct_aib2pld                                      (o_ch4_async_direct_aib2pld),
/* output [5:0]  */ .o_ch5_async_direct_aib2pld                                      (o_ch5_async_direct_aib2pld),
/* output [5:0]  */ .o_ch6_async_direct_aib2pld                                      (o_ch6_async_direct_aib2pld),
/* output [4:0]  */ .o_ch7_async_direct_aib2pld                                      (o_ch7_async_direct_aib2pld),
/* output [6:0]  */ .o_ch11_fsr_aib2pld                                              (o_ch11_fsr_aib2pld),
/* output [6:0]  */ .o_ch9_fsr_aib2pld                                               (o_ch9_fsr_aib2pld),
/* input  [7:0]  */ .i_ch0_async_direct_pld2aib                                      (i_ch0_async_direct_pld2aib),
/* input  [7:0]  */ .i_ch1_async_direct_pld2aib                                      (i_ch1_async_direct_pld2aib),
/* input  [7:0]  */ .i_ch2_async_direct_pld2aib                                      (i_ch2_async_direct_pld2aib),
/* input  [7:0]  */ .i_ch3_async_direct_pld2aib                                      (i_ch3_async_direct_pld2aib),
/* input  [7:0]  */ .i_ch4_async_direct_pld2aib                                      (i_ch4_async_direct_pld2aib),
/* input  [7:0]  */ .i_ch5_async_direct_pld2aib                                      (i_ch5_async_direct_pld2aib),
/* input  [7:0]  */ .i_ch6_async_direct_pld2aib                                      (i_ch6_async_direct_pld2aib),
/* input  [7:0]  */ .i_ch7_async_direct_pld2aib                                      (i_ch7_async_direct_pld2aib),
/* input  [6:0]  */ .i_ch11_fsr_pld2aib                                              (i_ch11_fsr_pld2aib),
/* input  [6:0]  */ .i_ch9_fsr_pld2aib                                               (i_ch9_fsr_pld2aib),
//* output [7:0]  */ .o_user_avmm_readdata                                            (o_user_avmm_readdata),
//* output        */ .o_user_avmm_readdatavalid                                       (o_user_avmm_readdatavalid),
//* output        */ .o_user_avmm_writedone                                           (o_user_avmm_writedone),
//* input         */ .i_user_avmm2_clk_rowclk                                         (i_user_avmm2_clk_rowclk),
//* input         */ .i_ch0_user_avmm1_clk_rowclk                                     (i_ch0_user_avmm1_clk_rowclk),
//* input         */ .i_user_avmm_read                                                (i_user_avmm_read),
//* input  [20:0] */ .i_user_avmm_reg_addr                                            (i_user_avmm_reg_addr),
//* input         */ .i_user_avmm_write                                               (i_user_avmm_write),
//* input  [7:0]  */ .i_user_avmm_writedata                                           (i_user_avmm_writedata),
/* input         */ .reconfig_clk                                                    (reconfig_clk),
/* input  [20:0] */ .reconfig_address                                                (reconfig_address),
/* input         */ .reconfig_read                                                   (reconfig_read),
/* output [ 7:0] */ .reconfig_readdata                                               (reconfig_readdata),
/* output        */ .reconfig_readdatavalid                                          (reconfig_readdatavalid),
/* input         */ .reconfig_write                                                  (reconfig_write),
/* input  [ 7:0] */ .reconfig_writedata                                              (reconfig_writedata),
/* output [ 4:0] */ .reconfig_reserved_out                                           (reconfig_reserved_out),
/* output        */ .reconfig_waitrequest                                            (reconfig_waitrequest),
/* output [ 7:0] */ .ln_reset_status_n                                               (ln_pipe_direct_reset_status_n_o),
/* input  [77:0] */ .ch13_pipe_direct_tx_octet1                                      (ch13_pipe_direct_tx_octet1),
/* input  [77:0] */ .ch14_pipe_direct_tx_octet1                                      (ch14_pipe_direct_tx_octet1),
/* input  [77:0] */ .ch15_pipe_direct_tx_octet1                                      (ch15_pipe_direct_tx_octet1),
/* input  [77:0] */ .ch16_pipe_direct_tx_octet1                                      (ch16_pipe_direct_tx_octet1),
/* input  [77:0] */ .ch17_pipe_direct_tx_octet1                                      (ch17_pipe_direct_tx_octet1),
/* input  [77:0] */ .ch18_pipe_direct_tx_octet1                                      (ch18_pipe_direct_tx_octet1),
/* input  [77:0] */ .ch19_pipe_direct_tx_octet1                                      (ch19_pipe_direct_tx_octet1),
/* input  [77:0] */ .ch20_pipe_direct_tx_octet1                                      (ch20_pipe_direct_tx_octet1),
/* input  [77:0] */ .ch21_pipe_direct_tx_octet1                                      (ch21_pipe_direct_tx_octet1),
/* input  [77:0] */ .ch22_pipe_direct_tx_octet1                                      (ch22_pipe_direct_tx_octet1),
/* output [77:0] */ .ch13_pipe_direct_rx_octet1                                      (ch13_pipe_direct_rx_octet1),
/* output [77:0] */ .ch14_pipe_direct_rx_octet1                                      (ch14_pipe_direct_rx_octet1),
/* output [77:0] */ .ch15_pipe_direct_rx_octet1                                      (ch15_pipe_direct_rx_octet1),
/* output [77:0] */ .ch16_pipe_direct_rx_octet1                                      (ch16_pipe_direct_rx_octet1),
/* output [77:0] */ .ch17_pipe_direct_rx_octet1                                      (ch17_pipe_direct_rx_octet1),
/* output [77:0] */ .ch18_pipe_direct_rx_octet1                                      (ch18_pipe_direct_rx_octet1),
/* output [77:0] */ .ch19_pipe_direct_rx_octet1                                      (ch19_pipe_direct_rx_octet1),
/* output [77:0] */ .ch20_pipe_direct_rx_octet1                                      (ch20_pipe_direct_rx_octet1),
/* output [77:0] */ .ch21_pipe_direct_rx_octet1                                      (ch21_pipe_direct_rx_octet1),
/* output [77:0] */ .ch22_pipe_direct_rx_octet1                                      (ch22_pipe_direct_rx_octet1),
/* output        */ .ch15_pipe_direct_tx_octet1_pwrdwn_status_l8                     (ch15_pipe_direct_tx_octet1_pwrdwn_status_l8),
/* output        */ .ch16_pipe_direct_tx_octet1_pwrdwn_status_l9                     (ch16_pipe_direct_tx_octet1_pwrdwn_status_l9),
/* output        */ .ch17_pipe_direct_tx_octet1_pwrdwn_status_l10                    (ch17_pipe_direct_tx_octet1_pwrdwn_status_l10),
/* output        */ .ch18_pipe_direct_tx_octet1_pwrdwn_status_l11                    (ch18_pipe_direct_tx_octet1_pwrdwn_status_l11),
/* output        */ .ch19_pipe_direct_tx_octet1_pwrdwn_status_l12                    (ch19_pipe_direct_tx_octet1_pwrdwn_status_l12),
/* output        */ .ch20_pipe_direct_tx_octet1_pwrdwn_status_l13                    (ch20_pipe_direct_tx_octet1_pwrdwn_status_l13),
/* output        */ .ch21_pipe_direct_tx_octet1_pwrdwn_status_l14                    (ch21_pipe_direct_tx_octet1_pwrdwn_status_l14),
/* output        */ .ch22_pipe_direct_tx_octet1_pwrdwn_status_l15                    (ch22_pipe_direct_tx_octet1_pwrdwn_status_l15),
/* input         */ .ch15_pipe_direct_tx_octet1_PLD_PCS_rst_n_l8                     (ch15_pipe_direct_tx_octet1_PLD_PCS_rst_n_l8),
/* input         */ .ch16_pipe_direct_tx_octet1_PLD_PCS_rst_n_l9                     (ch16_pipe_direct_tx_octet1_PLD_PCS_rst_n_l9),
/* input         */ .ch17_pipe_direct_tx_octet1_PLD_PCS_rst_n_l10                    (ch17_pipe_direct_tx_octet1_PLD_PCS_rst_n_l10),
/* input         */ .ch18_pipe_direct_tx_octet1_PLD_PCS_rst_n_l11                    (ch18_pipe_direct_tx_octet1_PLD_PCS_rst_n_l11),
/* input         */ .ch19_pipe_direct_tx_octet1_PLD_PCS_rst_n_l12                    (ch19_pipe_direct_tx_octet1_PLD_PCS_rst_n_l12),
/* input         */ .ch20_pipe_direct_tx_octet1_PLD_PCS_rst_n_l13                    (ch20_pipe_direct_tx_octet1_PLD_PCS_rst_n_l13),
/* input         */ .ch21_pipe_direct_tx_octet1_PLD_PCS_rst_n_l14                    (ch21_pipe_direct_tx_octet1_PLD_PCS_rst_n_l14),
/* input         */ .ch22_pipe_direct_tx_octet1_PLD_PCS_rst_n_l15                    (ch22_pipe_direct_tx_octet1_PLD_PCS_rst_n_l15),
/* output        */ .ch15_pipe_direct_rx_octet1_RXElecIdle_l8                        (ch15_pipe_direct_rx_octet1_RXElecIdle_l8),
/* output        */ .ch16_pipe_direct_rx_octet1_RXElecIdle_l9                        (ch16_pipe_direct_rx_octet1_RXElecIdle_l9),
/* output        */ .ch17_pipe_direct_rx_octet1_RXElecIdle_l10                       (ch17_pipe_direct_rx_octet1_RXElecIdle_l10),
/* output        */ .ch18_pipe_direct_rx_octet1_RXElecIdle_l11                       (ch18_pipe_direct_rx_octet1_RXElecIdle_l11),
/* output        */ .ch19_pipe_direct_rx_octet1_RXElecIdle_l12                       (ch19_pipe_direct_rx_octet1_RXElecIdle_l12),
/* output        */ .ch20_pipe_direct_rx_octet1_RXElecIdle_l13                       (ch20_pipe_direct_rx_octet1_RXElecIdle_l13),
/* output        */ .ch21_pipe_direct_rx_octet1_RXElecIdle_l14                       (ch21_pipe_direct_rx_octet1_RXElecIdle_l14),
/* output        */ .ch22_pipe_direct_rx_octet1_RXElecIdle_l15                       (ch22_pipe_direct_rx_octet1_RXElecIdle_l15),
/* output        */ .ch15_pipe_direct_rx_octet1_rx_cdrlock2data_l8                   (ch15_pipe_direct_rx_octet1_rx_cdrlock2data_l8),
/* output        */ .ch16_pipe_direct_rx_octet1_rx_cdrlock2data_l9                   (ch16_pipe_direct_rx_octet1_rx_cdrlock2data_l9),
/* output        */ .ch17_pipe_direct_rx_octet1_rx_cdrlock2data_l10                  (ch17_pipe_direct_rx_octet1_rx_cdrlock2data_l10),
/* output        */ .ch18_pipe_direct_rx_octet1_rx_cdrlock2data_l11                  (ch18_pipe_direct_rx_octet1_rx_cdrlock2data_l11),
/* output        */ .ch19_pipe_direct_rx_octet1_rx_cdrlock2data_l12                  (ch19_pipe_direct_rx_octet1_rx_cdrlock2data_l12),
/* output        */ .ch20_pipe_direct_rx_octet1_rx_cdrlock2data_l13                  (ch20_pipe_direct_rx_octet1_rx_cdrlock2data_l13),
/* output        */ .ch21_pipe_direct_rx_octet1_rx_cdrlock2data_l14                  (ch21_pipe_direct_rx_octet1_rx_cdrlock2data_l14),
/* output        */ .ch22_pipe_direct_rx_octet1_rx_cdrlock2data_l15                  (ch22_pipe_direct_rx_octet1_rx_cdrlock2data_l15),
/* output        */ .ch15_pipe_direct_rx_octet1_rx_cdrlockstatus_l8                  (ch15_pipe_direct_rx_octet1_rx_cdrlockstatus_l8),
/* output        */ .ch16_pipe_direct_rx_octet1_rx_cdrlockstatus_l9                  (ch16_pipe_direct_rx_octet1_rx_cdrlockstatus_l9),
/* output        */ .ch17_pipe_direct_rx_octet1_rx_cdrlockstatus_l10                 (ch17_pipe_direct_rx_octet1_rx_cdrlockstatus_l10),
/* output        */ .ch18_pipe_direct_rx_octet1_rx_cdrlockstatus_l11                 (ch18_pipe_direct_rx_octet1_rx_cdrlockstatus_l11),
/* output        */ .ch19_pipe_direct_rx_octet1_rx_cdrlockstatus_l12                 (ch19_pipe_direct_rx_octet1_rx_cdrlockstatus_l12),
/* output        */ .ch20_pipe_direct_rx_octet1_rx_cdrlockstatus_l13                 (ch20_pipe_direct_rx_octet1_rx_cdrlockstatus_l13),
/* output        */ .ch21_pipe_direct_rx_octet1_rx_cdrlockstatus_l14                 (ch21_pipe_direct_rx_octet1_rx_cdrlockstatus_l14),
/* output        */ .ch22_pipe_direct_rx_octet1_rx_cdrlockstatus_l15                 (ch22_pipe_direct_rx_octet1_rx_cdrlockstatus_l15),
/* output        */ .pipe_direct_rx_octet1_synthfast_lockstatus1                     (pipe_direct_rx_octet1_synthfast_lockstatus1),
/* output        */ .pipe_direct_rx_octet1_synthfast_ready1                          (pipe_direct_rx_octet1_synthfast_ready1),
/* output        */ .pipe_direct_rx_octet1_synthslow_lockstatus1                     (pipe_direct_rx_octet1_synthslow_lockstatus1),
/* output        */ .pipe_direct_rx_octet1_synthslow_ready1                          (pipe_direct_rx_octet1_synthslow_ready1),
/* output        */ .ch13_pipe_direct_pld_fabric_tx_transfer_en                      (ch13_pipe_direct_pld_fabric_tx_transfer_en),
/* output        */ .ch13_pipe_direct_pld_hssi_osc_transfer_en                       (ch13_pipe_direct_pld_hssi_osc_transfer_en),
/* output        */ .ch13_pipe_direct_pld_hssi_rx_transfer_en                        (ch13_pipe_direct_pld_hssi_rx_transfer_en),
/* input         */ .ch13_pipe_direct_pld_adapter_rx_pld_rst_n                       (ch13_pipe_direct_pld_adapter_rx_pld_rst_n),
/* input         */ .ch13_pipe_direct_pld_rx_dll_lock_req                            (ch13_pipe_direct_pld_rx_dll_lock_req),
/* input         */ .ch13_pipe_direct_pld_adapter_tx_pld_rst_n                       (ch13_pipe_direct_pld_adapter_tx_pld_rst_n),
/* input         */ .ch13_pipe_direct_pld_tx_dll_lock_req                            (ch13_pipe_direct_pld_tx_dll_lock_req),
/* output        */ .ch14_pipe_direct_pld_fabric_tx_transfer_en                      (ch14_pipe_direct_pld_fabric_tx_transfer_en),
/* output        */ .ch14_pipe_direct_pld_hssi_osc_transfer_en                       (ch14_pipe_direct_pld_hssi_osc_transfer_en),
/* output        */ .ch14_pipe_direct_pld_hssi_rx_transfer_en                        (ch14_pipe_direct_pld_hssi_rx_transfer_en),
/* input         */ .ch14_pipe_direct_pld_adapter_rx_pld_rst_n                       (ch14_pipe_direct_pld_adapter_rx_pld_rst_n),
/* input         */ .ch14_pipe_direct_pld_rx_dll_lock_req                            (ch14_pipe_direct_pld_rx_dll_lock_req),
/* input         */ .ch14_pipe_direct_pld_adapter_tx_pld_rst_n                       (ch14_pipe_direct_pld_adapter_tx_pld_rst_n),
/* input         */ .ch14_pipe_direct_pld_tx_dll_lock_req                            (ch14_pipe_direct_pld_tx_dll_lock_req),
/* output        */ .ch15_pipe_direct_pld_fabric_tx_transfer_en                      (ch15_pipe_direct_pld_fabric_tx_transfer_en),
/* output        */ .ch15_pipe_direct_pld_hssi_osc_transfer_en                       (ch15_pipe_direct_pld_hssi_osc_transfer_en),
/* output        */ .ch15_pipe_direct_pld_hssi_rx_transfer_en                        (ch15_pipe_direct_pld_hssi_rx_transfer_en),
/* input         */ .ch15_pipe_direct_pld_adapter_rx_pld_rst_n                       (ch15_pipe_direct_pld_adapter_rx_pld_rst_n),
/* input         */ .ch15_pipe_direct_pld_rx_dll_lock_req                            (ch15_pipe_direct_pld_rx_dll_lock_req),
/* input         */ .ch15_pipe_direct_pld_adapter_tx_pld_rst_n                       (ch15_pipe_direct_pld_adapter_tx_pld_rst_n),
/* input         */ .ch15_pipe_direct_pld_tx_dll_lock_req                            (ch15_pipe_direct_pld_tx_dll_lock_req),
/* output        */ .ch16_pipe_direct_pld_fabric_tx_transfer_en                      (ch16_pipe_direct_pld_fabric_tx_transfer_en),
/* output        */ .ch16_pipe_direct_pld_hssi_osc_transfer_en                       (ch16_pipe_direct_pld_hssi_osc_transfer_en),
/* output        */ .ch16_pipe_direct_pld_hssi_rx_transfer_en                        (ch16_pipe_direct_pld_hssi_rx_transfer_en),
/* input         */ .ch16_pipe_direct_pld_adapter_rx_pld_rst_n                       (ch16_pipe_direct_pld_adapter_rx_pld_rst_n),
/* input         */ .ch16_pipe_direct_pld_rx_dll_lock_req                            (ch16_pipe_direct_pld_rx_dll_lock_req),
/* input         */ .ch16_pipe_direct_pld_adapter_tx_pld_rst_n                       (ch16_pipe_direct_pld_adapter_tx_pld_rst_n),
/* input         */ .ch16_pipe_direct_pld_tx_dll_lock_req                            (ch16_pipe_direct_pld_tx_dll_lock_req),
/* output        */ .ch17_pipe_direct_pld_fabric_tx_transfer_en                      (ch17_pipe_direct_pld_fabric_tx_transfer_en),
/* output        */ .ch17_pipe_direct_pld_hssi_osc_transfer_en                       (ch17_pipe_direct_pld_hssi_osc_transfer_en),
/* output        */ .ch17_pipe_direct_pld_hssi_rx_transfer_en                        (ch17_pipe_direct_pld_hssi_rx_transfer_en),
/* input         */ .ch17_pipe_direct_pld_adapter_rx_pld_rst_n                       (ch17_pipe_direct_pld_adapter_rx_pld_rst_n),
/* input         */ .ch17_pipe_direct_pld_rx_dll_lock_req                            (ch17_pipe_direct_pld_rx_dll_lock_req),
/* input         */ .ch17_pipe_direct_pld_adapter_tx_pld_rst_n                       (ch17_pipe_direct_pld_adapter_tx_pld_rst_n),
/* input         */ .ch17_pipe_direct_pld_tx_dll_lock_req                            (ch17_pipe_direct_pld_tx_dll_lock_req),
/* output        */ .ch18_pipe_direct_pld_fabric_tx_transfer_en                      (ch18_pipe_direct_pld_fabric_tx_transfer_en),
/* output        */ .ch18_pipe_direct_pld_hssi_osc_transfer_en                       (ch18_pipe_direct_pld_hssi_osc_transfer_en),
/* output        */ .ch18_pipe_direct_pld_hssi_rx_transfer_en                        (ch18_pipe_direct_pld_hssi_rx_transfer_en),
/* input         */ .ch18_pipe_direct_pld_adapter_rx_pld_rst_n                       (ch18_pipe_direct_pld_adapter_rx_pld_rst_n),
/* input         */ .ch18_pipe_direct_pld_rx_dll_lock_req                            (ch18_pipe_direct_pld_rx_dll_lock_req),
/* input         */ .ch18_pipe_direct_pld_adapter_tx_pld_rst_n                       (ch18_pipe_direct_pld_adapter_tx_pld_rst_n),
/* input         */ .ch18_pipe_direct_pld_tx_dll_lock_req                            (ch18_pipe_direct_pld_tx_dll_lock_req),
/* output        */ .ch19_pipe_direct_pld_fabric_tx_transfer_en                      (ch19_pipe_direct_pld_fabric_tx_transfer_en),
/* output        */ .ch19_pipe_direct_pld_hssi_osc_transfer_en                       (ch19_pipe_direct_pld_hssi_osc_transfer_en),
/* output        */ .ch19_pipe_direct_pld_hssi_rx_transfer_en                        (ch19_pipe_direct_pld_hssi_rx_transfer_en),
/* input         */ .ch19_pipe_direct_pld_adapter_rx_pld_rst_n                       (ch19_pipe_direct_pld_adapter_rx_pld_rst_n),
/* input         */ .ch19_pipe_direct_pld_rx_dll_lock_req                            (ch19_pipe_direct_pld_rx_dll_lock_req),
/* input         */ .ch19_pipe_direct_pld_adapter_tx_pld_rst_n                       (ch19_pipe_direct_pld_adapter_tx_pld_rst_n),
/* input         */ .ch19_pipe_direct_pld_tx_dll_lock_req                            (ch19_pipe_direct_pld_tx_dll_lock_req),
/* output        */ .ch20_pipe_direct_pld_fabric_tx_transfer_en                      (ch20_pipe_direct_pld_fabric_tx_transfer_en),
/* output        */ .ch20_pipe_direct_pld_hssi_osc_transfer_en                       (ch20_pipe_direct_pld_hssi_osc_transfer_en),
/* output        */ .ch20_pipe_direct_pld_hssi_rx_transfer_en                        (ch20_pipe_direct_pld_hssi_rx_transfer_en),
/* input         */ .ch20_pipe_direct_pld_adapter_rx_pld_rst_n                       (ch20_pipe_direct_pld_adapter_rx_pld_rst_n),
/* input         */ .ch20_pipe_direct_pld_rx_dll_lock_req                            (ch20_pipe_direct_pld_rx_dll_lock_req),
/* input         */ .ch20_pipe_direct_pld_adapter_tx_pld_rst_n                       (ch20_pipe_direct_pld_adapter_tx_pld_rst_n),
/* input         */ .ch20_pipe_direct_pld_tx_dll_lock_req                            (ch20_pipe_direct_pld_tx_dll_lock_req),
/* output        */ .ch21_pipe_direct_pld_fabric_tx_transfer_en                      (ch21_pipe_direct_pld_fabric_tx_transfer_en),
/* output        */ .ch21_pipe_direct_pld_hssi_osc_transfer_en                       (ch21_pipe_direct_pld_hssi_osc_transfer_en),
/* output        */ .ch21_pipe_direct_pld_hssi_rx_transfer_en                        (ch21_pipe_direct_pld_hssi_rx_transfer_en),
/* input         */ .ch21_pipe_direct_pld_adapter_rx_pld_rst_n                       (ch21_pipe_direct_pld_adapter_rx_pld_rst_n),
/* input         */ .ch21_pipe_direct_pld_rx_dll_lock_req                            (ch21_pipe_direct_pld_rx_dll_lock_req),
/* input         */ .ch21_pipe_direct_pld_adapter_tx_pld_rst_n                       (ch21_pipe_direct_pld_adapter_tx_pld_rst_n),
/* input         */ .ch21_pipe_direct_pld_tx_dll_lock_req                            (ch21_pipe_direct_pld_tx_dll_lock_req),
/* output        */ .ch22_pipe_direct_pld_fabric_tx_transfer_en                      (ch22_pipe_direct_pld_fabric_tx_transfer_en),
/* output        */ .ch22_pipe_direct_pld_hssi_osc_transfer_en                       (ch22_pipe_direct_pld_hssi_osc_transfer_en),
/* output        */ .ch22_pipe_direct_pld_hssi_rx_transfer_en                        (ch22_pipe_direct_pld_hssi_rx_transfer_en),
/* input         */ .ch22_pipe_direct_pld_adapter_rx_pld_rst_n                       (ch22_pipe_direct_pld_adapter_rx_pld_rst_n),
/* input         */ .ch22_pipe_direct_pld_rx_dll_lock_req                            (ch22_pipe_direct_pld_rx_dll_lock_req),
/* input         */ .ch22_pipe_direct_pld_adapter_tx_pld_rst_n                       (ch22_pipe_direct_pld_adapter_tx_pld_rst_n),
/* input         */ .ch22_pipe_direct_pld_tx_dll_lock_req                            (ch22_pipe_direct_pld_tx_dll_lock_req),
/* output        */ .ch13_pipe_direct_pld_pcs_rx_clk_out1_dcm                        (ch13_pipe_direct_pld_pcs_rx_clk_out1_dcm),
/* output        */ .ch13_pipe_direct_pld_pcs_tx_clk_out1_dcm                        (ch13_pipe_direct_pld_pcs_tx_clk_out1_dcm),
/* output        */ .ch14_pipe_direct_pld_pcs_rx_clk_out1_dcm                        (ch14_pipe_direct_pld_pcs_rx_clk_out1_dcm),
/* output        */ .ch14_pipe_direct_pld_pcs_tx_clk_out1_dcm                        (ch14_pipe_direct_pld_pcs_tx_clk_out1_dcm),
/* output        */ .ch15_pipe_direct_pld_pcs_rx_clk_out1_dcm                        (ch15_pipe_direct_pld_pcs_rx_clk_out1_dcm),
/* output        */ .ch15_pipe_direct_pld_pcs_tx_clk_out1_dcm                        (ch15_pipe_direct_pld_pcs_tx_clk_out1_dcm),
/* output        */ .ch16_pipe_direct_pld_pcs_rx_clk_out1_dcm                        (ch16_pipe_direct_pld_pcs_rx_clk_out1_dcm),
/* output        */ .ch16_pipe_direct_pld_pcs_tx_clk_out1_dcm                        (ch16_pipe_direct_pld_pcs_tx_clk_out1_dcm),
/* output        */ .ch17_pipe_direct_pld_pcs_rx_clk_out1_dcm                        (ch17_pipe_direct_pld_pcs_rx_clk_out1_dcm),
/* output        */ .ch17_pipe_direct_pld_pcs_tx_clk_out1_dcm                        (ch17_pipe_direct_pld_pcs_tx_clk_out1_dcm),
/* output        */ .ch18_pipe_direct_pld_pcs_rx_clk_out1_dcm                        (ch18_pipe_direct_pld_pcs_rx_clk_out1_dcm),
/* output        */ .ch18_pipe_direct_pld_pcs_tx_clk_out1_dcm                        (ch18_pipe_direct_pld_pcs_tx_clk_out1_dcm),
/* output        */ .ch19_pipe_direct_pld_pcs_rx_clk_out1_dcm                        (ch19_pipe_direct_pld_pcs_rx_clk_out1_dcm),
/* output        */ .ch19_pipe_direct_pld_pcs_tx_clk_out1_dcm                        (ch19_pipe_direct_pld_pcs_tx_clk_out1_dcm),
/* output        */ .ch20_pipe_direct_pld_pcs_rx_clk_out1_dcm                        (ch20_pipe_direct_pld_pcs_rx_clk_out1_dcm),
/* output        */ .ch20_pipe_direct_pld_pcs_tx_clk_out1_dcm                        (ch20_pipe_direct_pld_pcs_tx_clk_out1_dcm),
/* output        */ .ch21_pipe_direct_pld_pcs_rx_clk_out1_dcm                        (ch21_pipe_direct_pld_pcs_rx_clk_out1_dcm),
/* output        */ .ch21_pipe_direct_pld_pcs_tx_clk_out1_dcm                        (ch21_pipe_direct_pld_pcs_tx_clk_out1_dcm),
/* output        */ .ch22_pipe_direct_pld_pcs_rx_clk_out1_dcm                        (ch22_pipe_direct_pld_pcs_rx_clk_out1_dcm),
/* output        */ .ch22_pipe_direct_pld_pcs_tx_clk_out1_dcm                        (ch22_pipe_direct_pld_pcs_tx_clk_out1_dcm),
/* input         */ .ch13_pipe_direct_pld_rx_clk1_dcm                                (ch13_pipe_direct_pld_rx_clk1_dcm),
/* input         */ .ch13_pipe_direct_pld_tx_clk1_dcm                                (ch13_pipe_direct_pld_tx_clk1_dcm),
/* input         */ .ch14_pipe_direct_pld_rx_clk1_dcm                                (ch14_pipe_direct_pld_rx_clk1_dcm),
/* input         */ .ch14_pipe_direct_pld_tx_clk1_dcm                                (ch14_pipe_direct_pld_tx_clk1_dcm),
/* input         */ .ch15_pipe_direct_pld_rx_clk1_dcm                                (ch15_pipe_direct_pld_rx_clk1_dcm),
/* input         */ .ch15_pipe_direct_pld_tx_clk1_dcm                                (ch15_pipe_direct_pld_tx_clk1_dcm),
/* input         */ .ch16_pipe_direct_pld_rx_clk1_dcm                                (ch16_pipe_direct_pld_rx_clk1_dcm),
/* input         */ .ch16_pipe_direct_pld_tx_clk1_dcm                                (ch16_pipe_direct_pld_tx_clk1_dcm),
/* input         */ .ch17_pipe_direct_pld_rx_clk1_dcm                                (ch17_pipe_direct_pld_rx_clk1_dcm),
/* input         */ .ch17_pipe_direct_pld_tx_clk1_dcm                                (ch17_pipe_direct_pld_tx_clk1_dcm),
/* input         */ .ch18_pipe_direct_pld_rx_clk1_dcm                                (ch18_pipe_direct_pld_rx_clk1_dcm),
/* input         */ .ch18_pipe_direct_pld_tx_clk1_dcm                                (ch18_pipe_direct_pld_tx_clk1_dcm),
/* input         */ .ch19_pipe_direct_pld_rx_clk1_dcm                                (ch19_pipe_direct_pld_rx_clk1_dcm),
/* input         */ .ch19_pipe_direct_pld_tx_clk1_dcm                                (ch19_pipe_direct_pld_tx_clk1_dcm),
/* input         */ .ch20_pipe_direct_pld_rx_clk1_dcm                                (ch20_pipe_direct_pld_rx_clk1_dcm),
/* input         */ .ch20_pipe_direct_pld_tx_clk1_dcm                                (ch20_pipe_direct_pld_tx_clk1_dcm),
/* input         */ .ch21_pipe_direct_pld_rx_clk1_dcm                                (ch21_pipe_direct_pld_rx_clk1_dcm),
/* input         */ .ch21_pipe_direct_pld_tx_clk1_dcm                                (ch21_pipe_direct_pld_tx_clk1_dcm),
/* input         */ .ch22_pipe_direct_pld_rx_clk1_dcm                                (ch22_pipe_direct_pld_rx_clk1_dcm),
/* input         */ .ch22_pipe_direct_pld_tx_clk1_dcm                                (ch22_pipe_direct_pld_tx_clk1_dcm),
/* input  [2:0]  */ .ial_phy_tx_fsr_0__tx_chnl_fsr                                   (ial_phy_tx_fsr_0__tx_chnl_fsr),
/* input  [3:0]  */ .ial_phy_tx_fsr_0__tx_ext_fsr                                    (ial_phy_tx_fsr_0__tx_ext_fsr),
/* input  [2:0]  */ .ial_phy_tx_fsr_1__tx_chnl_fsr                                   (ial_phy_tx_fsr_1__tx_chnl_fsr),
/* input  [3:0]  */ .ial_phy_tx_fsr_1__tx_ext_fsr                                    (ial_phy_tx_fsr_1__tx_ext_fsr),
/* input  [2:0]  */ .ial_phy_tx_fsr_2__tx_chnl_fsr                                   (ial_phy_tx_fsr_2__tx_chnl_fsr),
/* input  [3:0]  */ .ial_phy_tx_fsr_2__tx_ext_fsr                                    (ial_phy_tx_fsr_2__tx_ext_fsr),
/* input  [2:0]  */ .ial_phy_tx_fsr_3__tx_chnl_fsr                                   (ial_phy_tx_fsr_3__tx_chnl_fsr),
/* input  [3:0]  */ .ial_phy_tx_fsr_3__tx_ext_fsr                                    (ial_phy_tx_fsr_3__tx_ext_fsr),
/* input  [2:0]  */ .ial_phy_tx_fsr_4__tx_chnl_fsr                                   (ial_phy_tx_fsr_4__tx_chnl_fsr),
/* input  [3:0]  */ .ial_phy_tx_fsr_4__tx_ext_fsr                                    (ial_phy_tx_fsr_4__tx_ext_fsr),
/* input  [2:0]  */ .ial_phy_tx_fsr_5__tx_chnl_fsr                                   (ial_phy_tx_fsr_5__tx_chnl_fsr),
/* input  [3:0]  */ .ial_phy_tx_fsr_5__tx_ext_fsr                                    (ial_phy_tx_fsr_5__tx_ext_fsr),
/* input  [2:0]  */ .pcie_phy_tx_fsr_10__tx_chnl_fsr                                 (pcie_phy_tx_fsr_10__tx_chnl_fsr),
/* input  [3:0]  */ .pcie_phy_tx_fsr_10__tx_ext_fsr                                  (pcie_phy_tx_fsr_10__tx_ext_fsr),
/* input  [2:0]  */ .pcie_phy_tx_fsr_11__tx_chnl_fsr                                 (pcie_phy_tx_fsr_11__tx_chnl_fsr),
/* input  [3:0]  */ .pcie_phy_tx_fsr_11__tx_ext_fsr                                  (pcie_phy_tx_fsr_11__tx_ext_fsr),
/* output        */ .tx_n_out0                                                       (tx_n_out0),
/* output        */ .tx_n_out1                                                       (tx_n_out1),
/* output        */ .tx_n_out2                                                       (tx_n_out2),
/* output        */ .tx_n_out3                                                       (tx_n_out3),
/* output        */ .tx_n_out4                                                       (tx_n_out4),
/* output        */ .tx_n_out5                                                       (tx_n_out5),
/* output        */ .tx_n_out6                                                       (tx_n_out6),
/* output        */ .tx_n_out7                                                       (tx_n_out7),
/* output        */ .tx_n_out8                                                       (tx_n_out8),
/* output        */ .tx_n_out9                                                       (tx_n_out9),
/* output        */ .tx_n_out10                                                      (tx_n_out10),
/* output        */ .tx_n_out11                                                      (tx_n_out11),
/* output        */ .tx_n_out12                                                      (tx_n_out12),
/* output        */ .tx_n_out13                                                      (tx_n_out13),
/* output        */ .tx_n_out14                                                      (tx_n_out14),
/* output        */ .tx_n_out15                                                      (tx_n_out15),
/* output        */ .tx_p_out0                                                       (tx_p_out0),
/* output        */ .tx_p_out1                                                       (tx_p_out1),
/* output        */ .tx_p_out2                                                       (tx_p_out2),
/* output        */ .tx_p_out3                                                       (tx_p_out3),
/* output        */ .tx_p_out4                                                       (tx_p_out4),
/* output        */ .tx_p_out5                                                       (tx_p_out5),
/* output        */ .tx_p_out6                                                       (tx_p_out6),
/* output        */ .tx_p_out7                                                       (tx_p_out7),
/* output        */ .tx_p_out8                                                       (tx_p_out8),
/* output        */ .tx_p_out9                                                       (tx_p_out9),
/* output        */ .tx_p_out10                                                      (tx_p_out10),
/* output        */ .tx_p_out11                                                      (tx_p_out11),
/* output        */ .tx_p_out12                                                      (tx_p_out12),
/* output        */ .tx_p_out13                                                      (tx_p_out13),
/* output        */ .tx_p_out14                                                      (tx_p_out14),
/* output        */ .tx_p_out15                                                      (tx_p_out15),
/* input         */ .rx_n_in0                                                        (rx_n_in0),
/* input         */ .rx_n_in1                                                        (rx_n_in1),
/* input         */ .rx_n_in2                                                        (rx_n_in2),
/* input         */ .rx_n_in3                                                        (rx_n_in3),
/* input         */ .rx_n_in4                                                        (rx_n_in4),
/* input         */ .rx_n_in5                                                        (rx_n_in5),
/* input         */ .rx_n_in6                                                        (rx_n_in6),
/* input         */ .rx_n_in7                                                        (rx_n_in7),
/* input         */ .rx_n_in8                                                        (rx_n_in8),
/* input         */ .rx_n_in9                                                        (rx_n_in9),
/* input         */ .rx_n_in10                                                       (rx_n_in10),
/* input         */ .rx_n_in11                                                       (rx_n_in11),
/* input         */ .rx_n_in12                                                       (rx_n_in12),
/* input         */ .rx_n_in13                                                       (rx_n_in13),
/* input         */ .rx_n_in14                                                       (rx_n_in14),
/* input         */ .rx_n_in15                                                       (rx_n_in15),
/* input         */ .rx_p_in0                                                        (rx_p_in0),
/* input         */ .rx_p_in1                                                        (rx_p_in1),
/* input         */ .rx_p_in2                                                        (rx_p_in2),
/* input         */ .rx_p_in3                                                        (rx_p_in3),
/* input         */ .rx_p_in4                                                        (rx_p_in4),
/* input         */ .rx_p_in5                                                        (rx_p_in5),
/* input         */ .rx_p_in6                                                        (rx_p_in6),
/* input         */ .rx_p_in7                                                        (rx_p_in7),
/* input         */ .rx_p_in8                                                        (rx_p_in8),
/* input         */ .rx_p_in9                                                        (rx_p_in9),
/* input         */ .rx_p_in10                                                       (rx_p_in10),
/* input         */ .rx_p_in11                                                       (rx_p_in11),
/* input         */ .rx_p_in12                                                       (rx_p_in12),
/* input         */ .rx_p_in13                                                       (rx_p_in13),
/* input         */ .rx_p_in14                                                       (rx_p_in14),
/* input         */ .rx_p_in15                                                       (rx_p_in15),
/* output        */ .o_ch0_pld_pcs_rx_clk_out1_hioint                                (o_ch0_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch0_pld_pcs_rx_clk_out2_hioint                                (o_ch0_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch0_pld_pcs_tx_clk_out1_hioint                                (o_ch0_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch0_pld_pcs_tx_clk_out2_hioint                                (o_ch0_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch0_pld_pma_hclk_hioint                                       (o_ch0_pld_pma_hclk_hioint),
/* output        */ .o_ch0_pld_pma_internal_clk1_hioint                              (o_ch0_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch0_pld_pma_internal_clk2_hioint                              (o_ch0_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch10_pld_pcs_rx_clk_out1_hioint                               (o_ch10_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch10_pld_pcs_rx_clk_out2_hioint                               (o_ch10_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch10_pld_pcs_tx_clk_out1_hioint                               (o_ch10_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch10_pld_pcs_tx_clk_out2_hioint                               (o_ch10_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch10_pld_pma_hclk_hioint                                      (o_ch10_pld_pma_hclk_hioint),
/* output        */ .o_ch10_pld_pma_internal_clk1_hioint                             (o_ch10_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch10_pld_pma_internal_clk2_hioint                             (o_ch10_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch11_pld_pcs_rx_clk_out1_hioint                               (o_ch11_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch11_pld_pcs_rx_clk_out2_hioint                               (o_ch11_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch11_pld_pcs_tx_clk_out1_hioint                               (o_ch11_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch11_pld_pcs_tx_clk_out2_hioint                               (o_ch11_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch11_pld_pma_hclk_hioint                                      (o_ch11_pld_pma_hclk_hioint),
/* output        */ .o_ch11_pld_pma_internal_clk1_hioint                             (o_ch11_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch11_pld_pma_internal_clk2_hioint                             (o_ch11_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch12_pld_pcs_rx_clk_out1_hioint                               (o_ch12_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch12_pld_pcs_rx_clk_out2_hioint                               (o_ch12_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch12_pld_pcs_tx_clk_out1_hioint                               (o_ch12_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch12_pld_pcs_tx_clk_out2_hioint                               (o_ch12_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch12_pld_pma_hclk_hioint                                      (o_ch12_pld_pma_hclk_hioint),
/* output        */ .o_ch12_pld_pma_internal_clk1_hioint                             (o_ch12_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch12_pld_pma_internal_clk2_hioint                             (o_ch12_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch13_pld_pcs_rx_clk_out1_hioint                               (o_ch13_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch13_pld_pcs_rx_clk_out2_hioint                               (o_ch13_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch13_pld_pcs_tx_clk_out1_hioint                               (o_ch13_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch13_pld_pcs_tx_clk_out2_hioint                               (o_ch13_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch13_pld_pma_hclk_hioint                                      (o_ch13_pld_pma_hclk_hioint),
/* output        */ .o_ch13_pld_pma_internal_clk1_hioint                             (o_ch13_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch13_pld_pma_internal_clk2_hioint                             (o_ch13_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch14_pld_pcs_rx_clk_out1_hioint                               (o_ch14_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch14_pld_pcs_rx_clk_out2_hioint                               (o_ch14_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch14_pld_pcs_tx_clk_out1_hioint                               (o_ch14_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch14_pld_pcs_tx_clk_out2_hioint                               (o_ch14_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch14_pld_pma_hclk_hioint                                      (o_ch14_pld_pma_hclk_hioint),
/* output        */ .o_ch14_pld_pma_internal_clk1_hioint                             (o_ch14_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch14_pld_pma_internal_clk2_hioint                             (o_ch14_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch15_pld_pcs_rx_clk_out1_hioint                               (o_ch15_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch15_pld_pcs_rx_clk_out2_hioint                               (o_ch15_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch15_pld_pcs_tx_clk_out1_hioint                               (o_ch15_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch15_pld_pcs_tx_clk_out2_hioint                               (o_ch15_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch15_pld_pma_hclk_hioint                                      (o_ch15_pld_pma_hclk_hioint),
/* output        */ .o_ch15_pld_pma_internal_clk1_hioint                             (o_ch15_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch15_pld_pma_internal_clk2_hioint                             (o_ch15_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch16_pld_pcs_rx_clk_out1_hioint                               (o_ch16_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch16_pld_pcs_rx_clk_out2_hioint                               (o_ch16_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch16_pld_pcs_tx_clk_out1_hioint                               (o_ch16_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch16_pld_pcs_tx_clk_out2_hioint                               (o_ch16_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch16_pld_pma_hclk_hioint                                      (o_ch16_pld_pma_hclk_hioint),
/* output        */ .o_ch16_pld_pma_internal_clk1_hioint                             (o_ch16_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch16_pld_pma_internal_clk2_hioint                             (o_ch16_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch17_pld_pcs_rx_clk_out1_hioint                               (o_ch17_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch17_pld_pcs_rx_clk_out2_hioint                               (o_ch17_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch17_pld_pcs_tx_clk_out1_hioint                               (o_ch17_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch17_pld_pcs_tx_clk_out2_hioint                               (o_ch17_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch17_pld_pma_hclk_hioint                                      (o_ch17_pld_pma_hclk_hioint),
/* output        */ .o_ch17_pld_pma_internal_clk1_hioint                             (o_ch17_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch17_pld_pma_internal_clk2_hioint                             (o_ch17_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch18_pld_pcs_rx_clk_out1_hioint                               (o_ch18_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch18_pld_pcs_rx_clk_out2_hioint                               (o_ch18_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch18_pld_pcs_tx_clk_out1_hioint                               (o_ch18_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch18_pld_pcs_tx_clk_out2_hioint                               (o_ch18_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch18_pld_pma_hclk_hioint                                      (o_ch18_pld_pma_hclk_hioint),
/* output        */ .o_ch18_pld_pma_internal_clk1_hioint                             (o_ch18_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch18_pld_pma_internal_clk2_hioint                             (o_ch18_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch19_pld_pcs_rx_clk_out1_hioint                               (o_ch19_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch19_pld_pcs_rx_clk_out2_hioint                               (o_ch19_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch19_pld_pcs_tx_clk_out1_hioint                               (o_ch19_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch19_pld_pcs_tx_clk_out2_hioint                               (o_ch19_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch19_pld_pma_hclk_hioint                                      (o_ch19_pld_pma_hclk_hioint),
/* output        */ .o_ch19_pld_pma_internal_clk1_hioint                             (o_ch19_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch19_pld_pma_internal_clk2_hioint                             (o_ch19_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch1_pld_pcs_rx_clk_out1_hioint                                (o_ch1_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch1_pld_pcs_rx_clk_out2_hioint                                (o_ch1_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch1_pld_pcs_tx_clk_out1_hioint                                (o_ch1_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch1_pld_pcs_tx_clk_out2_hioint                                (o_ch1_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch1_pld_pma_hclk_hioint                                       (o_ch1_pld_pma_hclk_hioint),
/* output        */ .o_ch1_pld_pma_internal_clk1_hioint                              (o_ch1_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch1_pld_pma_internal_clk2_hioint                              (o_ch1_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch20_pld_pcs_rx_clk_out1_hioint                               (o_ch20_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch20_pld_pcs_rx_clk_out2_hioint                               (o_ch20_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch20_pld_pcs_tx_clk_out1_hioint                               (o_ch20_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch20_pld_pcs_tx_clk_out2_hioint                               (o_ch20_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch20_pld_pma_hclk_hioint                                      (o_ch20_pld_pma_hclk_hioint),
/* output        */ .o_ch20_pld_pma_internal_clk1_hioint                             (o_ch20_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch20_pld_pma_internal_clk2_hioint                             (o_ch20_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch21_pld_pcs_rx_clk_out1_hioint                               (o_ch21_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch21_pld_pcs_rx_clk_out2_hioint                               (o_ch21_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch21_pld_pcs_tx_clk_out1_hioint                               (o_ch21_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch21_pld_pcs_tx_clk_out2_hioint                               (o_ch21_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch21_pld_pma_hclk_hioint                                      (o_ch21_pld_pma_hclk_hioint),
/* output        */ .o_ch21_pld_pma_internal_clk1_hioint                             (o_ch21_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch21_pld_pma_internal_clk2_hioint                             (o_ch21_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch22_pld_pcs_rx_clk_out1_hioint                               (o_ch22_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch22_pld_pcs_rx_clk_out2_hioint                               (o_ch22_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch22_pld_pcs_tx_clk_out1_hioint                               (o_ch22_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch22_pld_pcs_tx_clk_out2_hioint                               (o_ch22_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch22_pld_pma_hclk_hioint                                      (o_ch22_pld_pma_hclk_hioint),
/* output        */ .o_ch22_pld_pma_internal_clk1_hioint                             (o_ch22_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch22_pld_pma_internal_clk2_hioint                             (o_ch22_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch23_pld_pcs_rx_clk_out1_hioint                               (o_ch23_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch23_pld_pcs_rx_clk_out2_hioint                               (o_ch23_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch23_pld_pcs_tx_clk_out1_hioint                               (o_ch23_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch23_pld_pcs_tx_clk_out2_hioint                               (o_ch23_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch23_pld_pma_hclk_hioint                                      (o_ch23_pld_pma_hclk_hioint),
/* output        */ .o_ch23_pld_pma_internal_clk1_hioint                             (o_ch23_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch23_pld_pma_internal_clk2_hioint                             (o_ch23_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch2_pld_pcs_rx_clk_out1_hioint                                (o_ch2_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch2_pld_pcs_rx_clk_out2_hioint                                (o_ch2_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch2_pld_pcs_tx_clk_out1_hioint                                (o_ch2_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch2_pld_pcs_tx_clk_out2_hioint                                (o_ch2_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch2_pld_pma_hclk_hioint                                       (o_ch2_pld_pma_hclk_hioint),
/* output        */ .o_ch2_pld_pma_internal_clk1_hioint                              (o_ch2_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch2_pld_pma_internal_clk2_hioint                              (o_ch2_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch3_pld_pcs_rx_clk_out1_hioint                                (o_ch3_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch3_pld_pcs_rx_clk_out2_hioint                                (o_ch3_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch3_pld_pcs_tx_clk_out1_hioint                                (o_ch3_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch3_pld_pcs_tx_clk_out2_hioint                                (o_ch3_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch3_pld_pma_hclk_hioint                                       (o_ch3_pld_pma_hclk_hioint),
/* output        */ .o_ch3_pld_pma_internal_clk1_hioint                              (o_ch3_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch3_pld_pma_internal_clk2_hioint                              (o_ch3_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch4_pld_pcs_rx_clk_out1_hioint                                (o_ch4_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch4_pld_pcs_rx_clk_out2_hioint                                (o_ch4_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch4_pld_pcs_tx_clk_out1_hioint                                (o_ch4_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch4_pld_pcs_tx_clk_out2_hioint                                (o_ch4_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch4_pld_pma_hclk_hioint                                       (o_ch4_pld_pma_hclk_hioint),
/* output        */ .o_ch4_pld_pma_internal_clk1_hioint                              (o_ch4_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch4_pld_pma_internal_clk2_hioint                              (o_ch4_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch5_pld_pcs_rx_clk_out1_hioint                                (o_ch5_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch5_pld_pcs_rx_clk_out2_hioint                                (o_ch5_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch5_pld_pcs_tx_clk_out1_hioint                                (o_ch5_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch5_pld_pcs_tx_clk_out2_hioint                                (o_ch5_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch5_pld_pma_hclk_hioint                                       (o_ch5_pld_pma_hclk_hioint),
/* output        */ .o_ch5_pld_pma_internal_clk1_hioint                              (o_ch5_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch5_pld_pma_internal_clk2_hioint                              (o_ch5_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch6_pld_pcs_rx_clk_out1_hioint                                (o_ch6_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch6_pld_pcs_rx_clk_out2_hioint                                (o_ch6_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch6_pld_pcs_tx_clk_out1_hioint                                (o_ch6_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch6_pld_pcs_tx_clk_out2_hioint                                (o_ch6_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch6_pld_pma_hclk_hioint                                       (o_ch6_pld_pma_hclk_hioint),
/* output        */ .o_ch6_pld_pma_internal_clk1_hioint                              (o_ch6_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch6_pld_pma_internal_clk2_hioint                              (o_ch6_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch7_pld_pcs_rx_clk_out1_hioint                                (o_ch7_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch7_pld_pcs_rx_clk_out2_hioint                                (o_ch7_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch7_pld_pcs_tx_clk_out1_hioint                                (o_ch7_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch7_pld_pcs_tx_clk_out2_hioint                                (o_ch7_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch7_pld_pma_hclk_hioint                                       (o_ch7_pld_pma_hclk_hioint),
/* output        */ .o_ch7_pld_pma_internal_clk1_hioint                              (o_ch7_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch7_pld_pma_internal_clk2_hioint                              (o_ch7_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch8_pld_pcs_rx_clk_out1_hioint                                (o_ch8_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch8_pld_pcs_rx_clk_out2_hioint                                (o_ch8_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch8_pld_pcs_tx_clk_out1_hioint                                (o_ch8_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch8_pld_pcs_tx_clk_out2_hioint                                (o_ch8_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch8_pld_pma_hclk_hioint                                       (o_ch8_pld_pma_hclk_hioint),
/* output        */ .o_ch8_pld_pma_internal_clk1_hioint                              (o_ch8_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch8_pld_pma_internal_clk2_hioint                              (o_ch8_pld_pma_internal_clk2_hioint),
/* output        */ .o_ch9_pld_pcs_rx_clk_out1_hioint                                (o_ch9_pld_pcs_rx_clk_out1_hioint),
/* output        */ .o_ch9_pld_pcs_rx_clk_out2_hioint                                (o_ch9_pld_pcs_rx_clk_out2_hioint),
/* output        */ .o_ch9_pld_pcs_tx_clk_out1_hioint                                (o_ch9_pld_pcs_tx_clk_out1_hioint),
/* output        */ .o_ch9_pld_pcs_tx_clk_out2_hioint                                (o_ch9_pld_pcs_tx_clk_out2_hioint),
/* output        */ .o_ch9_pld_pma_hclk_hioint                                       (o_ch9_pld_pma_hclk_hioint),
/* output        */ .o_ch9_pld_pma_internal_clk1_hioint                              (o_ch9_pld_pma_internal_clk1_hioint),
/* output        */ .o_ch9_pld_pma_internal_clk2_hioint                              (o_ch9_pld_pma_internal_clk2_hioint),
/* input         */ .i_ch0_pld_pma_coreclkin_rowclk                                  (i_ch0_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch0_pld_rx_clk2_rowclk                                        (i_ch0_pld_rx_clk2_rowclk),
/* input         */ .i_ch0_pld_sclk1_rowclk                                          (i_ch0_pld_sclk1_rowclk),
/* input         */ .i_ch0_pld_sclk2_rowclk                                          (i_ch0_pld_sclk2_rowclk),
/* input         */ .i_ch10_pld_pma_coreclkin_rowclk                                 (i_ch10_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch10_pld_rx_clk2_rowclk                                       (i_ch10_pld_rx_clk2_rowclk),
/* input         */ .i_ch10_pld_sclk1_rowclk                                         (i_ch10_pld_sclk1_rowclk),
/* input         */ .i_ch10_pld_sclk2_rowclk                                         (i_ch10_pld_sclk2_rowclk),
/* input         */ .i_ch10_user_avmm1_clk_rowclk                                    (i_ch10_user_avmm1_clk_rowclk),
/* input         */ .i_ch10_user_avmm2_clk_rowclk                                    (i_ch10_user_avmm2_clk_rowclk),
/* input         */ .i_ch11_pld_pma_coreclkin_rowclk                                 (i_ch11_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch11_pld_rx_clk2_rowclk                                       (i_ch11_pld_rx_clk2_rowclk),
/* input         */ .i_ch11_pld_sclk1_rowclk                                         (i_ch11_pld_sclk1_rowclk),
/* input         */ .i_ch11_pld_sclk2_rowclk                                         (i_ch11_pld_sclk2_rowclk),
/* input         */ .i_ch11_user_avmm1_clk_rowclk                                    (i_ch11_user_avmm1_clk_rowclk),
/* input         */ .i_ch11_user_avmm2_clk_rowclk                                    (i_ch11_user_avmm2_clk_rowclk),
/* input         */ .i_ch12_pld_pma_coreclkin_rowclk                                 (i_ch12_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch12_pld_rx_clk2_rowclk                                       (i_ch12_pld_rx_clk2_rowclk),
/* input         */ .i_ch12_pld_sclk1_rowclk                                         (i_ch12_pld_sclk1_rowclk),
/* input         */ .i_ch12_pld_sclk2_rowclk                                         (i_ch12_pld_sclk2_rowclk),
/* input         */ .i_ch12_user_avmm1_clk_rowclk                                    (i_ch12_user_avmm1_clk_rowclk),
/* input         */ .i_ch12_user_avmm2_clk_rowclk                                    (i_ch12_user_avmm2_clk_rowclk),
/* input         */ .i_ch13_pld_pma_coreclkin_rowclk                                 (i_ch13_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch13_pld_rx_clk2_rowclk                                       (i_ch13_pld_rx_clk2_rowclk),
/* input         */ .i_ch13_pld_sclk1_rowclk                                         (i_ch13_pld_sclk1_rowclk),
/* input         */ .i_ch13_pld_sclk2_rowclk                                         (i_ch13_pld_sclk2_rowclk),
/* input         */ .i_ch13_user_avmm1_clk_rowclk                                    (i_ch13_user_avmm1_clk_rowclk),
/* input         */ .i_ch13_user_avmm2_clk_rowclk                                    (i_ch13_user_avmm2_clk_rowclk),
/* input         */ .i_ch14_pld_pma_coreclkin_rowclk                                 (i_ch14_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch14_pld_rx_clk2_rowclk                                       (i_ch14_pld_rx_clk2_rowclk),
/* input         */ .i_ch14_pld_sclk1_rowclk                                         (i_ch14_pld_sclk1_rowclk),
/* input         */ .i_ch14_pld_sclk2_rowclk                                         (i_ch14_pld_sclk2_rowclk),
/* input         */ .i_ch14_user_avmm1_clk_rowclk                                    (i_ch14_user_avmm1_clk_rowclk),
/* input         */ .i_ch14_user_avmm2_clk_rowclk                                    (i_ch14_user_avmm2_clk_rowclk),
/* input         */ .i_ch15_pld_pma_coreclkin_rowclk                                 (i_ch15_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch15_pld_rx_clk2_rowclk                                       (i_ch15_pld_rx_clk2_rowclk),
/* input         */ .i_ch15_pld_sclk1_rowclk                                         (i_ch15_pld_sclk1_rowclk),
/* input         */ .i_ch15_pld_sclk2_rowclk                                         (i_ch15_pld_sclk2_rowclk),
/* input         */ .i_ch15_user_avmm1_clk_rowclk                                    (i_ch15_user_avmm1_clk_rowclk),
/* input         */ .i_ch15_user_avmm2_clk_rowclk                                    (i_ch15_user_avmm2_clk_rowclk),
/* input         */ .i_ch16_pld_pma_coreclkin_rowclk                                 (i_ch16_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch16_pld_rx_clk2_rowclk                                       (i_ch16_pld_rx_clk2_rowclk),
/* input         */ .i_ch16_pld_sclk1_rowclk                                         (i_ch16_pld_sclk1_rowclk),
/* input         */ .i_ch16_pld_sclk2_rowclk                                         (i_ch16_pld_sclk2_rowclk),
/* input         */ .i_ch16_user_avmm1_clk_rowclk                                    (i_ch16_user_avmm1_clk_rowclk),
/* input         */ .i_ch16_user_avmm2_clk_rowclk                                    (i_ch16_user_avmm2_clk_rowclk),
/* input         */ .i_ch17_pld_pma_coreclkin_rowclk                                 (i_ch17_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch17_pld_rx_clk2_rowclk                                       (i_ch17_pld_rx_clk2_rowclk),
/* input         */ .i_ch17_pld_sclk1_rowclk                                         (i_ch17_pld_sclk1_rowclk),
/* input         */ .i_ch17_pld_sclk2_rowclk                                         (i_ch17_pld_sclk2_rowclk),
/* input         */ .i_ch17_user_avmm1_clk_rowclk                                    (i_ch17_user_avmm1_clk_rowclk),
/* input         */ .i_ch17_user_avmm2_clk_rowclk                                    (i_ch17_user_avmm2_clk_rowclk),
/* input         */ .i_ch18_pld_pma_coreclkin_rowclk                                 (i_ch18_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch18_pld_rx_clk2_rowclk                                       (i_ch18_pld_rx_clk2_rowclk),
/* input         */ .i_ch18_pld_sclk1_rowclk                                         (i_ch18_pld_sclk1_rowclk),
/* input         */ .i_ch18_pld_sclk2_rowclk                                         (i_ch18_pld_sclk2_rowclk),
/* input         */ .i_ch18_user_avmm1_clk_rowclk                                    (i_ch18_user_avmm1_clk_rowclk),
/* input         */ .i_ch18_user_avmm2_clk_rowclk                                    (i_ch18_user_avmm2_clk_rowclk),
/* input         */ .i_ch19_pld_pma_coreclkin_rowclk                                 (i_ch19_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch19_pld_rx_clk2_rowclk                                       (i_ch19_pld_rx_clk2_rowclk),
/* input         */ .i_ch19_pld_sclk1_rowclk                                         (i_ch19_pld_sclk1_rowclk),
/* input         */ .i_ch19_pld_sclk2_rowclk                                         (i_ch19_pld_sclk2_rowclk),
/* input         */ .i_ch19_user_avmm1_clk_rowclk                                    (i_ch19_user_avmm1_clk_rowclk),
/* input         */ .i_ch19_user_avmm2_clk_rowclk                                    (i_ch19_user_avmm2_clk_rowclk),
/* input         */ .i_ch1_pld_pma_coreclkin_rowclk                                  (i_ch1_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch1_pld_rx_clk2_rowclk                                        (i_ch1_pld_rx_clk2_rowclk),
/* input         */ .i_ch1_pld_sclk1_rowclk                                          (i_ch1_pld_sclk1_rowclk),
/* input         */ .i_ch1_pld_sclk2_rowclk                                          (i_ch1_pld_sclk2_rowclk),
/* input         */ .i_ch1_user_avmm1_clk_rowclk                                     (i_ch1_user_avmm1_clk_rowclk),
/* input         */ .i_ch1_user_avmm2_clk_rowclk                                     (i_ch1_user_avmm2_clk_rowclk),
/* input         */ .i_ch20_pld_pma_coreclkin_rowclk                                 (i_ch20_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch20_pld_rx_clk2_rowclk                                       (i_ch20_pld_rx_clk2_rowclk),
/* input         */ .i_ch20_pld_sclk1_rowclk                                         (i_ch20_pld_sclk1_rowclk),
/* input         */ .i_ch20_pld_sclk2_rowclk                                         (i_ch20_pld_sclk2_rowclk),
/* input         */ .i_ch20_user_avmm1_clk_rowclk                                    (i_ch20_user_avmm1_clk_rowclk),
/* input         */ .i_ch20_user_avmm2_clk_rowclk                                    (i_ch20_user_avmm2_clk_rowclk),
/* input         */ .i_ch21_pld_pma_coreclkin_rowclk                                 (i_ch21_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch21_pld_rx_clk2_rowclk                                       (i_ch21_pld_rx_clk2_rowclk),
/* input         */ .i_ch21_pld_sclk1_rowclk                                         (i_ch21_pld_sclk1_rowclk),
/* input         */ .i_ch21_pld_sclk2_rowclk                                         (i_ch21_pld_sclk2_rowclk),
/* input         */ .i_ch21_user_avmm1_clk_rowclk                                    (i_ch21_user_avmm1_clk_rowclk),
/* input         */ .i_ch21_user_avmm2_clk_rowclk                                    (i_ch21_user_avmm2_clk_rowclk),
/* input         */ .i_ch22_pld_pma_coreclkin_rowclk                                 (i_ch22_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch22_pld_rx_clk2_rowclk                                       (i_ch22_pld_rx_clk2_rowclk),
/* input         */ .i_ch22_pld_sclk1_rowclk                                         (i_ch22_pld_sclk1_rowclk),
/* input         */ .i_ch22_pld_sclk2_rowclk                                         (i_ch22_pld_sclk2_rowclk),
/* input         */ .i_ch22_user_avmm1_clk_rowclk                                    (i_ch22_user_avmm1_clk_rowclk),
/* input         */ .i_ch22_user_avmm2_clk_rowclk                                    (i_ch22_user_avmm2_clk_rowclk),
/* input         */ .i_ch23_pld_pma_coreclkin_rowclk                                 (i_ch23_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch23_pld_rx_clk2_rowclk                                       (i_ch23_pld_rx_clk2_rowclk),
/* input         */ .i_ch23_pld_sclk1_rowclk                                         (i_ch23_pld_sclk1_rowclk),
/* input         */ .i_ch23_pld_sclk2_rowclk                                         (i_ch23_pld_sclk2_rowclk),
/* input         */ .i_ch23_user_avmm1_clk_rowclk                                    (i_ch23_user_avmm1_clk_rowclk),
/* input         */ .i_ch23_user_avmm2_clk_rowclk                                    (i_ch23_user_avmm2_clk_rowclk),
/* input         */ .i_ch2_pld_pma_coreclkin_rowclk                                  (i_ch2_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch2_pld_rx_clk2_rowclk                                        (i_ch2_pld_rx_clk2_rowclk),
/* input         */ .i_ch2_pld_sclk1_rowclk                                          (i_ch2_pld_sclk1_rowclk),
/* input         */ .i_ch2_pld_sclk2_rowclk                                          (i_ch2_pld_sclk2_rowclk),
/* input         */ .i_ch2_user_avmm1_clk_rowclk                                     (i_ch2_user_avmm1_clk_rowclk),
/* input         */ .i_ch2_user_avmm2_clk_rowclk                                     (i_ch2_user_avmm2_clk_rowclk),
/* input         */ .i_ch3_pld_pma_coreclkin_rowclk                                  (i_ch3_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch3_pld_rx_clk2_rowclk                                        (i_ch3_pld_rx_clk2_rowclk),
/* input         */ .i_ch3_pld_sclk1_rowclk                                          (i_ch3_pld_sclk1_rowclk),
/* input         */ .i_ch3_pld_sclk2_rowclk                                          (i_ch3_pld_sclk2_rowclk),
/* input         */ .i_ch3_user_avmm1_clk_rowclk                                     (i_ch3_user_avmm1_clk_rowclk),
/* input         */ .i_ch3_user_avmm2_clk_rowclk                                     (i_ch3_user_avmm2_clk_rowclk),
/* input         */ .i_ch4_pld_pma_coreclkin_rowclk                                  (i_ch4_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch4_pld_rx_clk2_rowclk                                        (i_ch4_pld_rx_clk2_rowclk),
/* input         */ .i_ch4_pld_sclk1_rowclk                                          (i_ch4_pld_sclk1_rowclk),
/* input         */ .i_ch4_pld_sclk2_rowclk                                          (i_ch4_pld_sclk2_rowclk),
/* input         */ .i_ch4_user_avmm1_clk_rowclk                                     (i_ch4_user_avmm1_clk_rowclk),
/* input         */ .i_ch4_user_avmm2_clk_rowclk                                     (i_ch4_user_avmm2_clk_rowclk),
/* input         */ .i_ch5_pld_pma_coreclkin_rowclk                                  (i_ch5_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch5_pld_rx_clk2_rowclk                                        (i_ch5_pld_rx_clk2_rowclk),
/* input         */ .i_ch5_pld_sclk1_rowclk                                          (i_ch5_pld_sclk1_rowclk),
/* input         */ .i_ch5_pld_sclk2_rowclk                                          (i_ch5_pld_sclk2_rowclk),
/* input         */ .i_ch5_user_avmm1_clk_rowclk                                     (i_ch5_user_avmm1_clk_rowclk),
/* input         */ .i_ch5_user_avmm2_clk_rowclk                                     (i_ch5_user_avmm2_clk_rowclk),
/* input         */ .i_ch6_pld_pma_coreclkin_rowclk                                  (i_ch6_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch6_pld_rx_clk2_rowclk                                        (i_ch6_pld_rx_clk2_rowclk),
/* input         */ .i_ch6_pld_sclk1_rowclk                                          (i_ch6_pld_sclk1_rowclk),
/* input         */ .i_ch6_pld_sclk2_rowclk                                          (i_ch6_pld_sclk2_rowclk),
/* input         */ .i_ch6_user_avmm1_clk_rowclk                                     (i_ch6_user_avmm1_clk_rowclk),
/* input         */ .i_ch6_user_avmm2_clk_rowclk                                     (i_ch6_user_avmm2_clk_rowclk),
/* input         */ .i_ch7_pld_pma_coreclkin_rowclk                                  (i_ch7_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch7_pld_rx_clk2_rowclk                                        (i_ch7_pld_rx_clk2_rowclk),
/* input         */ .i_ch7_pld_sclk1_rowclk                                          (i_ch7_pld_sclk1_rowclk),
/* input         */ .i_ch7_pld_sclk2_rowclk                                          (i_ch7_pld_sclk2_rowclk),
/* input         */ .i_ch7_user_avmm1_clk_rowclk                                     (i_ch7_user_avmm1_clk_rowclk),
/* input         */ .i_ch7_user_avmm2_clk_rowclk                                     (i_ch7_user_avmm2_clk_rowclk),
/* input         */ .i_ch8_pld_pma_coreclkin_rowclk                                  (i_ch8_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch8_pld_rx_clk2_rowclk                                        (i_ch8_pld_rx_clk2_rowclk),
/* input         */ .i_ch8_pld_sclk1_rowclk                                          (i_ch8_pld_sclk1_rowclk),
/* input         */ .i_ch8_pld_sclk2_rowclk                                          (i_ch8_pld_sclk2_rowclk),
/* input         */ .i_ch8_user_avmm1_clk_rowclk                                     (i_ch8_user_avmm1_clk_rowclk),
/* input         */ .i_ch8_user_avmm2_clk_rowclk                                     (i_ch8_user_avmm2_clk_rowclk),
/* input         */ .i_ch9_pld_pma_coreclkin_rowclk                                  (i_ch9_pld_pma_coreclkin_rowclk),
/* input         */ .i_ch9_pld_rx_clk2_rowclk                                        (i_ch9_pld_rx_clk2_rowclk),
/* input         */ .i_ch9_pld_sclk1_rowclk                                          (i_ch9_pld_sclk1_rowclk),
/* input         */ .i_ch9_pld_sclk2_rowclk                                          (i_ch9_pld_sclk2_rowclk),
/* input         */ .i_ch9_user_avmm1_clk_rowclk                                     (i_ch9_user_avmm1_clk_rowclk),
/* input         */ .i_ch9_user_avmm2_clk_rowclk                                     (i_ch9_user_avmm2_clk_rowclk),
/* output [2:0]  */ .o_ch0_pld_fpll_shared_direct_async_out_dcm                      (o_ch0_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch0_pld_pcs_rx_clk_out1_dcm                                   (o_ch0_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch0_pld_pcs_rx_clk_out2_dcm                                   (o_ch0_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch0_pld_pcs_tx_clk_out1_dcm                                   (o_ch0_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch0_pld_pcs_tx_clk_out2_dcm                                   (o_ch0_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch10_pld_fpll_shared_direct_async_out_dcm                     (o_ch10_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch10_pld_pcs_rx_clk_out1_dcm                                  (o_ch10_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch10_pld_pcs_rx_clk_out2_dcm                                  (o_ch10_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch10_pld_pcs_tx_clk_out1_dcm                                  (o_ch10_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch10_pld_pcs_tx_clk_out2_dcm                                  (o_ch10_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch11_pld_fpll_shared_direct_async_out_dcm                     (o_ch11_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch11_pld_pcs_rx_clk_out1_dcm                                  (o_ch11_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch11_pld_pcs_rx_clk_out2_dcm                                  (o_ch11_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch11_pld_pcs_tx_clk_out1_dcm                                  (o_ch11_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch11_pld_pcs_tx_clk_out2_dcm                                  (o_ch11_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch12_pld_fpll_shared_direct_async_out_dcm                     (o_ch12_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch12_pld_pcs_rx_clk_out1_dcm                                  (o_ch12_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch12_pld_pcs_rx_clk_out2_dcm                                  (o_ch12_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch12_pld_pcs_tx_clk_out1_dcm                                  (o_ch12_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch12_pld_pcs_tx_clk_out2_dcm                                  (o_ch12_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch13_pld_fpll_shared_direct_async_out_dcm                     (o_ch13_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch13_pld_pcs_rx_clk_out1_dcm                                  (o_ch13_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch13_pld_pcs_rx_clk_out2_dcm                                  (o_ch13_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch13_pld_pcs_tx_clk_out1_dcm                                  (o_ch13_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch13_pld_pcs_tx_clk_out2_dcm                                  (o_ch13_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch14_pld_fpll_shared_direct_async_out_dcm                     (o_ch14_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch14_pld_pcs_rx_clk_out1_dcm                                  (o_ch14_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch14_pld_pcs_rx_clk_out2_dcm                                  (o_ch14_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch14_pld_pcs_tx_clk_out1_dcm                                  (o_ch14_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch14_pld_pcs_tx_clk_out2_dcm                                  (o_ch14_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch15_pld_fpll_shared_direct_async_out_dcm                     (o_ch15_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch15_pld_pcs_rx_clk_out2_dcm                                  (o_ch15_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch15_pld_pcs_tx_clk_out1_dcm                                  (o_ch15_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch15_pld_pcs_tx_clk_out2_dcm                                  (o_ch15_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch16_pld_fpll_shared_direct_async_out_dcm                     (o_ch16_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch16_pld_pcs_rx_clk_out1_dcm                                  (o_ch16_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch16_pld_pcs_rx_clk_out2_dcm                                  (o_ch16_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch16_pld_pcs_tx_clk_out1_dcm                                  (o_ch16_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch16_pld_pcs_tx_clk_out2_dcm                                  (o_ch16_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch17_pld_fpll_shared_direct_async_out_dcm                     (o_ch17_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch17_pld_pcs_rx_clk_out1_dcm                                  (o_ch17_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch17_pld_pcs_rx_clk_out2_dcm                                  (o_ch17_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch17_pld_pcs_tx_clk_out1_dcm                                  (o_ch17_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch17_pld_pcs_tx_clk_out2_dcm                                  (o_ch17_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch18_pld_fpll_shared_direct_async_out_dcm                     (o_ch18_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch18_pld_pcs_rx_clk_out1_dcm                                  (o_ch18_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch18_pld_pcs_rx_clk_out2_dcm                                  (o_ch18_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch18_pld_pcs_tx_clk_out1_dcm                                  (o_ch18_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch18_pld_pcs_tx_clk_out2_dcm                                  (o_ch18_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch19_pld_fpll_shared_direct_async_out_dcm                     (o_ch19_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch19_pld_pcs_rx_clk_out1_dcm                                  (o_ch19_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch19_pld_pcs_rx_clk_out2_dcm                                  (o_ch19_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch19_pld_pcs_tx_clk_out1_dcm                                  (o_ch19_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch19_pld_pcs_tx_clk_out2_dcm                                  (o_ch19_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch1_pld_fpll_shared_direct_async_out_dcm                      (o_ch1_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch1_pld_pcs_rx_clk_out1_dcm                                   (o_ch1_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch1_pld_pcs_rx_clk_out2_dcm                                   (o_ch1_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch1_pld_pcs_tx_clk_out1_dcm                                   (o_ch1_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch1_pld_pcs_tx_clk_out2_dcm                                   (o_ch1_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch20_pld_fpll_shared_direct_async_out_dcm                     (o_ch20_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch20_pld_pcs_rx_clk_out1_dcm                                  (o_ch20_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch20_pld_pcs_rx_clk_out2_dcm                                  (o_ch20_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch20_pld_pcs_tx_clk_out1_dcm                                  (o_ch20_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch20_pld_pcs_tx_clk_out2_dcm                                  (o_ch20_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch21_pld_fpll_shared_direct_async_out_dcm                     (o_ch21_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch21_pld_pcs_rx_clk_out1_dcm                                  (o_ch21_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch21_pld_pcs_rx_clk_out2_dcm                                  (o_ch21_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch21_pld_pcs_tx_clk_out1_dcm                                  (o_ch21_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch21_pld_pcs_tx_clk_out2_dcm                                  (o_ch21_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch22_pld_fpll_shared_direct_async_out_dcm                     (o_ch22_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch22_pld_pcs_rx_clk_out1_dcm                                  (o_ch22_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch22_pld_pcs_rx_clk_out2_dcm                                  (o_ch22_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch22_pld_pcs_tx_clk_out1_dcm                                  (o_ch22_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch22_pld_pcs_tx_clk_out2_dcm                                  (o_ch22_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch23_pld_fpll_shared_direct_async_out_dcm                     (o_ch23_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch23_pld_pcs_rx_clk_out1_dcm                                  (o_ch23_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch23_pld_pcs_rx_clk_out2_dcm                                  (o_ch23_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch23_pld_pcs_tx_clk_out1_dcm                                  (o_ch23_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch23_pld_pcs_tx_clk_out2_dcm                                  (o_ch23_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch2_pld_fpll_shared_direct_async_out_dcm                      (o_ch2_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch2_pld_pcs_rx_clk_out1_dcm                                   (o_ch2_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch2_pld_pcs_rx_clk_out2_dcm                                   (o_ch2_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch2_pld_pcs_tx_clk_out1_dcm                                   (o_ch2_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch2_pld_pcs_tx_clk_out2_dcm                                   (o_ch2_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch3_pld_fpll_shared_direct_async_out_dcm                      (o_ch3_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch3_pld_pcs_rx_clk_out1_dcm                                   (o_ch3_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch3_pld_pcs_rx_clk_out2_dcm                                   (o_ch3_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch3_pld_pcs_tx_clk_out1_dcm                                   (o_ch3_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch3_pld_pcs_tx_clk_out2_dcm                                   (o_ch3_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch4_pld_fpll_shared_direct_async_out_dcm                      (o_ch4_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch4_pld_pcs_rx_clk_out1_dcm                                   (o_ch4_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch4_pld_pcs_rx_clk_out2_dcm                                   (o_ch4_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch4_pld_pcs_tx_clk_out1_dcm                                   (o_ch4_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch4_pld_pcs_tx_clk_out2_dcm                                   (o_ch4_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch5_pld_fpll_shared_direct_async_out_dcm                      (o_ch5_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch5_pld_pcs_rx_clk_out1_dcm                                   (o_ch5_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch5_pld_pcs_rx_clk_out2_dcm                                   (o_ch5_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch5_pld_pcs_tx_clk_out1_dcm                                   (o_ch5_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch5_pld_pcs_tx_clk_out2_dcm                                   (o_ch5_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch6_pld_fpll_shared_direct_async_out_dcm                      (o_ch6_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch6_pld_pcs_rx_clk_out1_dcm                                   (o_ch6_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch6_pld_pcs_rx_clk_out2_dcm                                   (o_ch6_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch6_pld_pcs_tx_clk_out1_dcm                                   (o_ch6_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch6_pld_pcs_tx_clk_out2_dcm                                   (o_ch6_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch7_pld_fpll_shared_direct_async_out_dcm                      (o_ch7_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch7_pld_pcs_rx_clk_out1_dcm                                   (o_ch7_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch7_pld_pcs_rx_clk_out2_dcm                                   (o_ch7_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch7_pld_pcs_tx_clk_out1_dcm                                   (o_ch7_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch7_pld_pcs_tx_clk_out2_dcm                                   (o_ch7_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch8_pld_fpll_shared_direct_async_out_dcm                      (o_ch8_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch8_pld_pcs_rx_clk_out1_dcm                                   (o_ch8_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch8_pld_pcs_rx_clk_out2_dcm                                   (o_ch8_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch8_pld_pcs_tx_clk_out1_dcm                                   (o_ch8_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch8_pld_pcs_tx_clk_out2_dcm                                   (o_ch8_pld_pcs_tx_clk_out2_dcm),
/* output [2:0]  */ .o_ch9_pld_fpll_shared_direct_async_out_dcm                      (o_ch9_pld_fpll_shared_direct_async_out_dcm),
/* output        */ .o_ch9_pld_pcs_rx_clk_out1_dcm                                   (o_ch9_pld_pcs_rx_clk_out1_dcm),
/* output        */ .o_ch9_pld_pcs_rx_clk_out2_dcm                                   (o_ch9_pld_pcs_rx_clk_out2_dcm),
/* output        */ .o_ch9_pld_pcs_tx_clk_out1_dcm                                   (o_ch9_pld_pcs_tx_clk_out1_dcm),
/* output        */ .o_ch9_pld_pcs_tx_clk_out2_dcm                                   (o_ch9_pld_pcs_tx_clk_out2_dcm),
/* input  [1:0]  */ .i_ch0_pld_fpll_shared_direct_async_in_dcm                       (i_ch0_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch0_pld_rx_clk2_dcm                                           (i_ch0_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch10_pld_fpll_shared_direct_async_in_dcm                      (i_ch10_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch10_pld_rx_clk2_dcm                                          (i_ch10_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch11_pld_fpll_shared_direct_async_in_dcm                      (i_ch11_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch11_pld_rx_clk2_dcm                                          (i_ch11_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch12_pld_fpll_shared_direct_async_in_dcm                      (i_ch12_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch12_pld_rx_clk2_dcm                                          (i_ch12_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch13_pld_fpll_shared_direct_async_in_dcm                      (i_ch13_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch13_pld_rx_clk2_dcm                                          (i_ch13_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch14_pld_fpll_shared_direct_async_in_dcm                      (i_ch14_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch14_pld_rx_clk2_dcm                                          (i_ch14_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch15_pld_fpll_shared_direct_async_in_dcm                      (i_ch15_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch15_pld_rx_clk2_dcm                                          (i_ch15_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch16_pld_fpll_shared_direct_async_in_dcm                      (i_ch16_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch16_pld_rx_clk2_dcm                                          (i_ch16_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch17_pld_fpll_shared_direct_async_in_dcm                      (i_ch17_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch17_pld_rx_clk2_dcm                                          (i_ch17_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch18_pld_fpll_shared_direct_async_in_dcm                      (i_ch18_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch18_pld_rx_clk2_dcm                                          (i_ch18_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch19_pld_fpll_shared_direct_async_in_dcm                      (i_ch19_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch19_pld_rx_clk2_dcm                                          (i_ch19_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch1_pld_fpll_shared_direct_async_in_dcm                       (i_ch1_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch1_pld_rx_clk2_dcm                                           (i_ch1_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch20_pld_fpll_shared_direct_async_in_dcm                      (i_ch20_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch20_pld_rx_clk2_dcm                                          (i_ch20_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch21_pld_fpll_shared_direct_async_in_dcm                      (i_ch21_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch21_pld_rx_clk2_dcm                                          (i_ch21_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch22_pld_fpll_shared_direct_async_in_dcm                      (i_ch22_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch22_pld_rx_clk2_dcm                                          (i_ch22_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch23_pld_fpll_shared_direct_async_in_dcm                      (i_ch23_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch23_pld_rx_clk2_dcm                                          (i_ch23_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch2_pld_fpll_shared_direct_async_in_dcm                       (i_ch2_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch2_pld_rx_clk2_dcm                                           (i_ch2_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch3_pld_fpll_shared_direct_async_in_dcm                       (i_ch3_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch3_pld_rx_clk2_dcm                                           (i_ch3_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch4_pld_fpll_shared_direct_async_in_dcm                       (i_ch4_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch4_pld_rx_clk2_dcm                                           (i_ch4_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch5_pld_fpll_shared_direct_async_in_dcm                       (i_ch5_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch5_pld_rx_clk2_dcm                                           (i_ch5_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch6_pld_fpll_shared_direct_async_in_dcm                       (i_ch6_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch6_pld_rx_clk2_dcm                                           (i_ch6_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch7_pld_fpll_shared_direct_async_in_dcm                       (i_ch7_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch7_pld_rx_clk2_dcm                                           (i_ch7_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch8_pld_fpll_shared_direct_async_in_dcm                       (i_ch8_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch8_pld_rx_clk2_dcm                                           (i_ch8_pld_rx_clk2_dcm),
/* input  [1:0]  */ .i_ch9_pld_fpll_shared_direct_async_in_dcm                       (i_ch9_pld_fpll_shared_direct_async_in_dcm),
/* input         */ .i_ch9_pld_rx_clk2_dcm                                           (i_ch9_pld_rx_clk2_dcm),
/* input         */ .i_aux_por_vccl_ovr                                              (i_aux_por_vccl_ovr),
/* input  [3:0]  */ .i_id                                                            (i_id),
/* input         */ .i_jtag_hijack                                                   (i_jtag_hijack),
/* input         */ .i_jtag_tck                                                      (i_jtag_tck),
/* input         */ .i_jtag_tdi                                                      (i_jtag_tdi),
/* output        */ .io_jtag_tdo                                                     (io_jtag_tdo),
/* input         */ .i_jtag_tms                                                      (i_jtag_tms),
/* input         */ .i_jtag_trst                                                     (i_jtag_trst),
/* input         */ .i_sens_therm                                                    (i_sens_therm),
/* input         */ .i_strap_spare_in0                                               (i_strap_spare_in0),
/* input         */ .i_strap_spare_in1                                               (i_strap_spare_in1),
/* inout         */ .io_aprobe2_0                                                    ( ),
/* inout         */ .io_aprobe2_1                                                    ( ),
/* inout         */ .io_aprobe_0                                                     ( ),
/* inout         */ .io_aprobe_1                                                     ( ),
/* inout  [23:0] */ .io_dfx                                                          ( ),
/* input         */ .i_edm_in                                                        (i_edm_in),
/* output        */ .o_edm_out                                                       (o_edm_out),
/* output        */ .o_sens_therm                                                    (o_sens_therm),
/* inout         */ .aprobe_dts_0                                                    ( ),
/* inout         */ .aprobe_dts_1                                                    ( ),
/* inout         */ .aprobe_pll_0                                                    ( ),
/* inout         */ .aprobe_pll_1                                                    ( ),
/* inout         */ .io_rcomp_n_0                                                    ( ),
/* inout         */ .io_rcomp_n_1                                                    ( ),
/* inout         */ .io_rcomp_p_0                                                    ( ),
/* inout         */ .io_rcomp_p_1                                                    ( ),
/* input         */ .s0_0_1__maib_rotate__maib_rotate                                (s0_0_1__maib_rotate__maib_rotate),
/* input         */ .s0_187_1__aib_jtag_return__tdo                                  (s0_187_1__aib_jtag_return__tdo),
/* input         */ .s1_0_1__aib_jtag_out__tck                                       (s1_0_1__aib_jtag_out__tck),
/* input         */ .s1_0_1__aib_jtag_out__tdi                                       (s1_0_1__aib_jtag_out__tdi),
/* input         */ .s1_0_1__aib_jtag_out__tms                                       (s1_0_1__aib_jtag_out__tms),
/* input         */ .s1_0_1__dts_temptrip__temptrip                                  (s1_0_1__dts_temptrip__temptrip),
/* input         */ .s2_0_1__aib_jtag_out__tck                                       (s2_0_1__aib_jtag_out__tck),
/* input         */ .s2_0_1__aib_jtag_out__tdi                                       (s2_0_1__aib_jtag_out__tdi),
/* input         */ .s2_0_1__aib_jtag_out__tms                                       (s2_0_1__aib_jtag_out__tms),
/* input         */ .s2_187_1__aib_jtag_return__tdo                                  (s2_187_1__aib_jtag_return__tdo),
/* input  [3:0]  */ .s4_0_1__aib_cjtag_ctrl_id__cjtag_id                             (s4_0_1__aib_cjtag_ctrl_id__cjtag_id),
/* input         */ .s5_187_1__cnoc__abort                                           (s5_187_1__cnoc__abort),
/* input         */ .s5_187_1__cnoc__clk                                             (s5_187_1__cnoc__clk),
/* input         */ .s5_187_1__cnoc__clk_n                                           (s5_187_1__cnoc__clk_n),
/* input  [32:0] */ .s5_187_1__cnoc__data                                            (s5_187_1__cnoc__data),
/* input         */ .s5_187_1__cnoc__end_of_packet                                   (s5_187_1__cnoc__end_of_packet),
/* input         */ .s5_187_1__cnoc__nonsecure_interrupt                             (s5_187_1__cnoc__nonsecure_interrupt),
/* input         */ .s5_187_1__cnoc__por                                             (s5_187_1__cnoc__por),
/* input         */ .s5_187_1__cnoc__por_n                                           (s5_187_1__cnoc__por_n),
/* input         */ .s5_187_1__cnoc__secure_interrupt                                (s5_187_1__cnoc__secure_interrupt),
/* input         */ .s5_187_1__cnoc__start_of_packet                                 (s5_187_1__cnoc__start_of_packet),
/* input         */ .s5_187_1__cnoc__sync                                            (s5_187_1__cnoc__sync),
/* input         */ .s5_187_1__cnoc__valid                                           (s5_187_1__cnoc__valid),
/* input         */ .s5_187_1__cnoc__warm_reset_n                                    (s5_187_1__cnoc__warm_reset_n),
/* input         */ .s8_187_1__aib_jtag_return__tdo                                  (s8_187_1__aib_jtag_return__tdo),
/* input         */ .s9_0_1__aib_jtag_out__tck                                       (s9_0_1__aib_jtag_out__tck),
/* input         */ .s9_0_1__aib_jtag_out__tdi                                       (s9_0_1__aib_jtag_out__tdi),
/* input         */ .s9_0_1__aib_jtag_out__tms                                       (s9_0_1__aib_jtag_out__tms),
/* input         */ .s11_187_1__aib_jtag_out__tck                                    (s11_187_1__aib_jtag_out__tck),
/* input         */ .s11_187_1__aib_jtag_out__tdi                                    (s11_187_1__aib_jtag_out__tdi),
/* input         */ .s11_187_1__aib_jtag_out__tms                                    (s11_187_1__aib_jtag_out__tms),
/* input         */ .s12_187_1__aib_jtag_out__tck                                    (s12_187_1__aib_jtag_out__tck),
/* input         */ .s12_187_1__aib_jtag_out__tdi                                    (s12_187_1__aib_jtag_out__tdi),
/* input         */ .s12_187_1__aib_jtag_out__tms                                    (s12_187_1__aib_jtag_out__tms),
/* input         */ .s13_0_1__aib_jtag_return__tdo                                   (s13_0_1__aib_jtag_return__tdo),
/* input         */ .s14_0_1__cjtag__tck                                             (s14_0_1__cjtag__tck),
/* input         */ .s14_0_1__cjtag__tdi                                             (s14_0_1__cjtag__tdi),
/* input         */ .s14_0_1__cjtag__tms                                             (s14_0_1__cjtag__tms),
/* input  [3:0]  */ .s14_187_1__aib_cjtag_ctrl_id__cjtag_id                          (s14_187_1__aib_cjtag_ctrl_id__cjtag_id),
/* input         */ .s15_187_1__cjtag__tck                                           (s15_187_1__cjtag__tck),
/* input         */ .s15_187_1__cjtag__tdi                                           (s15_187_1__cjtag__tdi),
/* input         */ .s15_187_1__cjtag__tms                                           (s15_187_1__cjtag__tms),
/* input         */ .s16_0_1__aib_jtag_return__tdo                                   (s16_0_1__aib_jtag_return__tdo),
/* input         */ .s17_187_1__cjtag_return__tdo                                    (s17_187_1__cjtag_return__tdo),
/* input         */ .s18_0_1__aib_jtag_return__tdo                                   (s18_0_1__aib_jtag_return__tdo),
/* input         */ .s19_187_1__aib_jtag_out__tck                                    (s19_187_1__aib_jtag_out__tck),
/* input         */ .s19_187_1__aib_jtag_out__tdi                                    (s19_187_1__aib_jtag_out__tdi),
/* input         */ .s19_187_1__aib_jtag_out__tms                                    (s19_187_1__aib_jtag_out__tms),
/* input         */ .s20_187_1__cnoc__abort                                          (s20_187_1__cnoc__abort),
/* input         */ .s20_187_1__cnoc__clk                                            (s20_187_1__cnoc__clk),
/* input         */ .s20_187_1__cnoc__clk_n                                          (s20_187_1__cnoc__clk_n),
/* input  [32:0] */ .s20_187_1__cnoc__data                                           (s20_187_1__cnoc__data),
/* input         */ .s20_187_1__cnoc__end_of_packet                                  (s20_187_1__cnoc__end_of_packet),
/* input         */ .s20_187_1__cnoc__nonsecure_interrupt                            (s20_187_1__cnoc__nonsecure_interrupt),
/* input         */ .s20_187_1__cnoc__por                                            (s20_187_1__cnoc__por),
/* input         */ .s20_187_1__cnoc__por_n                                          (s20_187_1__cnoc__por_n),
/* input         */ .s20_187_1__cnoc__secure_interrupt                               (s20_187_1__cnoc__secure_interrupt),
/* input         */ .s20_187_1__cnoc__start_of_packet                                (s20_187_1__cnoc__start_of_packet),
/* input         */ .s20_187_1__cnoc__sync                                           (s20_187_1__cnoc__sync),
/* input         */ .s20_187_1__cnoc__valid                                          (s20_187_1__cnoc__valid),
/* input         */ .s20_187_1__cnoc__warm_reset_n                                   (s20_187_1__cnoc__warm_reset_n),
/* input         */ .s21_0_1__cjtag_return__tdo                                      (s21_0_1__cjtag_return__tdo),
/* input         */ .s23_0_1__cnoc__abort                                            (s23_0_1__cnoc__abort),
/* input         */ .s23_0_1__cnoc__clk                                              (s23_0_1__cnoc__clk),
/* input         */ .s23_0_1__cnoc__clk_n                                            (s23_0_1__cnoc__clk_n),
/* input  [32:0] */ .s23_0_1__cnoc__data                                             (s23_0_1__cnoc__data),
/* input         */ .s23_0_1__cnoc__end_of_packet                                    (s23_0_1__cnoc__end_of_packet),
/* input         */ .s23_0_1__cnoc__nonsecure_interrupt                              (s23_0_1__cnoc__nonsecure_interrupt),
/* input         */ .s23_0_1__cnoc__por                                              (s23_0_1__cnoc__por),
/* input         */ .s23_0_1__cnoc__por_n                                            (s23_0_1__cnoc__por_n),
/* input         */ .s23_0_1__cnoc__secure_interrupt                                 (s23_0_1__cnoc__secure_interrupt),
/* input         */ .s23_0_1__cnoc__start_of_packet                                  (s23_0_1__cnoc__start_of_packet),
/* input         */ .s23_0_1__cnoc__sync                                             (s23_0_1__cnoc__sync),
/* input         */ .s23_0_1__cnoc__valid                                            (s23_0_1__cnoc__valid),
/* input         */ .s23_0_1__cnoc__warm_reset_n                                     (s23_0_1__cnoc__warm_reset_n),
/* input         */ .s23_187_1__include_aib_jtag_segment__include_aib_jtag_segment   (s23_187_1__include_aib_jtag_segment__include_aib_jtag_segment),
/* input         */ .s25_187_1__include_aib_jtag_segment__include_aib_jtag_segment   (s25_187_1__include_aib_jtag_segment__include_aib_jtag_segment),
/* input         */ .s27_187_1__include_aib_jtag_segment__include_aib_jtag_segment   (s27_187_1__include_aib_jtag_segment__include_aib_jtag_segment),
/* input         */ .s28_187_1__dts_temptrip__temptrip                               (s28_187_1__dts_temptrip__temptrip),
/* input         */ .s30_0_1__dc_bsc_sdata__s_data                                   (s30_0_1__dc_bsc_sdata__s_data),
/* input         */ .s30_187_1__dc_bsc_sdata__s_data                                 (s30_187_1__dc_bsc_sdata__s_data),
/* input         */ .s32_187_1__sdm_mission_bus__clk                                 (s32_187_1__sdm_mission_bus__clk),
/* input  [31:0] */ .s32_187_1__sdm_mission_bus__data                                (s32_187_1__sdm_mission_bus__data),
/* input         */ .s32_187_1__sdm_mission_bus__valid                               (s32_187_1__sdm_mission_bus__valid),
/* input  [27:0] */ .s33_187_1__sdm_test_bus__data                                   (s33_187_1__sdm_test_bus__data),
/* input  [15:0] */ .s34_0_1__sdm_testmode_ctrl__test_io_ctrl                        (s34_0_1__sdm_testmode_ctrl__test_io_ctrl),
/* input  [15:0] */ .s37_0_1__test_return__data                                      (s37_0_1__test_return__data),
/* input         */ .s37_0_1__test_return__valid                                     (s37_0_1__test_return__valid),
/* input  [4:0]  */ .s38_0_1__scan_sdm_so__scan_out                                  (s38_0_1__scan_sdm_so__scan_out),
/* input  [3:0]  */ .s39_0_1__cr_ctrl__muxsel_avst                                   (s39_0_1__cr_ctrl__muxsel_avst),
/* input         */ .s39_0_1__cr_ctrl__muxsel_test_cnoc                              (s39_0_1__cr_ctrl__muxsel_test_cnoc),
/* input         */ .s124_0_1__include_aib_jtag_segment__include_aib_jtag_segment    (s124_0_1__include_aib_jtag_segment__include_aib_jtag_segment),
/* input         */ .s126_0_1__include_aib_jtag_segment__include_aib_jtag_segment    (s126_0_1__include_aib_jtag_segment__include_aib_jtag_segment),
/* input         */ .s128_0_1__include_aib_jtag_segment__include_aib_jtag_segment    (s128_0_1__include_aib_jtag_segment__include_aib_jtag_segment),
/* output [107:0]*/ .o_s0_23_1__core_periphery__data_to_core                         (o_s0_23_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_44_1__core_periphery__data_to_core                         (o_s0_44_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_45_1__core_periphery__data_to_core                         (o_s0_45_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_46_1__core_periphery__data_to_core                         (o_s0_46_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_47_1__core_periphery__data_to_core                         (o_s0_47_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_48_1__core_periphery__data_to_core                         (o_s0_48_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_49_1__core_periphery__data_to_core                         (o_s0_49_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_70_1__core_periphery__data_to_core                         (o_s0_70_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_91_1__core_periphery__data_to_core                         (o_s0_91_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_92_1__core_periphery__data_to_core                         (o_s0_92_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_93_1__core_periphery__data_to_core                         (o_s0_93_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_94_1__core_periphery__data_to_core                         (o_s0_94_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_95_1__core_periphery__data_to_core                         (o_s0_95_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_96_1__core_periphery__data_to_core                         (o_s0_96_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_117_1__core_periphery__data_to_core                        (o_s0_117_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_138_1__core_periphery__data_to_core                        (o_s0_138_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_139_1__core_periphery__data_to_core                        (o_s0_139_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_140_1__core_periphery__data_to_core                        (o_s0_140_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_141_1__core_periphery__data_to_core                        (o_s0_141_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_142_1__core_periphery__data_to_core                        (o_s0_142_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_143_1__core_periphery__data_to_core                        (o_s0_143_1__core_periphery__data_to_core),
/* output [107:0]*/ .o_s0_164_1__core_periphery__data_to_core                        (o_s0_164_1__core_periphery__data_to_core),
/* output [65:0] */ .s0_100_1__core_periphery__data_to_core_unused                   (s0_100_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_101_1__core_periphery__data_to_core_unused                   (s0_101_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_105_1__core_periphery__data_to_core_unused                   (s0_105_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_106_1__core_periphery__data_to_core_unused                   (s0_106_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_107_1__core_periphery__data_to_core_unused                   (s0_107_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_108_1__core_periphery__data_to_core_unused                   (s0_108_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_111_1__core_periphery__data_to_core_unused                   (s0_111_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_112_1__core_periphery__data_to_core_unused                   (s0_112_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_113_1__core_periphery__data_to_core_unused                   (s0_113_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_114_1__core_periphery__data_to_core_unused                   (s0_114_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_11_1__core_periphery__data_to_core_unused                    (s0_11_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_120_1__core_periphery__data_to_core_unused                   (s0_120_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_121_1__core_periphery__data_to_core_unused                   (s0_121_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_122_1__core_periphery__data_to_core_unused                   (s0_122_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_126_1__core_periphery__data_to_core_unused                   (s0_126_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_127_1__core_periphery__data_to_core_unused                   (s0_127_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_128_1__core_periphery__data_to_core_unused                   (s0_128_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_12_1__core_periphery__data_to_core_unused                    (s0_12_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_133_1__core_periphery__data_to_core_unused                   (s0_133_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_134_1__core_periphery__data_to_core_unused                   (s0_134_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_135_1__core_periphery__data_to_core_unused                   (s0_135_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_13_1__core_periphery__data_to_core_unused                    (s0_13_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_145_1__core_periphery__data_to_core_unused                   (s0_145_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_146_1__core_periphery__data_to_core_unused                   (s0_146_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_147_1__core_periphery__data_to_core_unused                   (s0_147_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_14_1__core_periphery__data_to_core_unused                    (s0_14_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_152_1__core_periphery__data_to_core_unused                   (s0_152_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_153_1__core_periphery__data_to_core_unused                   (s0_153_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_154_1__core_periphery__data_to_core_unused                   (s0_154_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_158_1__core_periphery__data_to_core_unused                   (s0_158_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_159_1__core_periphery__data_to_core_unused                   (s0_159_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_160_1__core_periphery__data_to_core_unused                   (s0_160_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_167_1__core_periphery__data_to_core_unused                   (s0_167_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_168_1__core_periphery__data_to_core_unused                   (s0_168_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_169_1__core_periphery__data_to_core_unused                   (s0_169_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_173_1__core_periphery__data_to_core_unused                   (s0_173_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_174_1__core_periphery__data_to_core_unused                   (s0_174_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_175_1__core_periphery__data_to_core_unused                   (s0_175_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_17_1__core_periphery__data_to_core_unused                    (s0_17_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_180_1__core_periphery__data_to_core_unused                   (s0_180_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_181_1__core_periphery__data_to_core_unused                   (s0_181_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_182_1__core_periphery__data_to_core_unused                   (s0_182_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_183_1__core_periphery__data_to_core_unused                   (s0_183_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_18_1__core_periphery__data_to_core_unused                    (s0_18_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_19_1__core_periphery__data_to_core_unused                    (s0_19_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_20_1__core_periphery__data_to_core_unused                    (s0_20_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_26_1__core_periphery__data_to_core_unused                    (s0_26_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_27_1__core_periphery__data_to_core_unused                    (s0_27_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_28_1__core_periphery__data_to_core_unused                    (s0_28_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_29_1__core_periphery__data_to_core_unused                    (s0_29_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_32_1__core_periphery__data_to_core_unused                    (s0_32_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_33_1__core_periphery__data_to_core_unused                    (s0_33_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_34_1__core_periphery__data_to_core_unused                    (s0_34_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_35_1__core_periphery__data_to_core_unused                    (s0_35_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_39_1__core_periphery__data_to_core_unused                    (s0_39_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_40_1__core_periphery__data_to_core_unused                    (s0_40_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_41_1__core_periphery__data_to_core_unused                    (s0_41_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_42_1__core_periphery__data_to_core_unused                    (s0_42_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_4_1__core_periphery__data_to_core_unused                     (s0_4_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_51_1__core_periphery__data_to_core_unused                    (s0_51_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_52_1__core_periphery__data_to_core_unused                    (s0_52_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_53_1__core_periphery__data_to_core_unused                    (s0_53_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_54_1__core_periphery__data_to_core_unused                    (s0_54_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_58_1__core_periphery__data_to_core_unused                    (s0_58_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_59_1__core_periphery__data_to_core_unused                    (s0_59_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_5_1__core_periphery__data_to_core_unused                     (s0_5_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_60_1__core_periphery__data_to_core_unused                    (s0_60_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_61_1__core_periphery__data_to_core_unused                    (s0_61_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_64_1__core_periphery__data_to_core_unused                    (s0_64_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_65_1__core_periphery__data_to_core_unused                    (s0_65_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_66_1__core_periphery__data_to_core_unused                    (s0_66_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_67_1__core_periphery__data_to_core_unused                    (s0_67_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_6_1__core_periphery__data_to_core_unused                     (s0_6_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_73_1__core_periphery__data_to_core_unused                    (s0_73_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_74_1__core_periphery__data_to_core_unused                    (s0_74_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_75_1__core_periphery__data_to_core_unused                    (s0_75_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_76_1__core_periphery__data_to_core_unused                    (s0_76_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_79_1__core_periphery__data_to_core_unused                    (s0_79_1__core_periphery__data_to_core_unused),
/* output [85:0] */ .s0_7_1__core_periphery__data_to_core_unused                     (s0_7_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_80_1__core_periphery__data_to_core_unused                    (s0_80_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_81_1__core_periphery__data_to_core_unused                    (s0_81_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_82_1__core_periphery__data_to_core_unused                    (s0_82_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_86_1__core_periphery__data_to_core_unused                    (s0_86_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_87_1__core_periphery__data_to_core_unused                    (s0_87_1__core_periphery__data_to_core_unused),
/* output [65:0] */ .s0_88_1__core_periphery__data_to_core_unused                    (s0_88_1__core_periphery__data_to_core_unused),
/* output [95:0] */ .s0_89_1__core_periphery__data_to_core_unused                    (s0_89_1__core_periphery__data_to_core_unused),
/* output [39:0] */ .s0_98_1__core_periphery__data_to_core_unused                    (s0_98_1__core_periphery__data_to_core_unused),
/* output [53:0] */ .s0_99_1__core_periphery__data_to_core_unused                    (s0_99_1__core_periphery__data_to_core_unused),
/* input  [15:0] */ .i_s0_3_1__core_periphery__clock_from_core                       (i_s0_3_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_8_1__core_periphery__clock_from_core                       (i_s0_8_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_9_1__core_periphery__clock_from_core                       (i_s0_9_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_10_1__core_periphery__clock_from_core                      (i_s0_10_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_15_1__core_periphery__clock_from_core                      (i_s0_15_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_16_1__core_periphery__clock_from_core                      (i_s0_16_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_21_1__core_periphery__clock_from_core                      (i_s0_21_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_22_1__core_periphery__clock_from_core                      (i_s0_22_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_23_1__core_periphery__clock_from_core                      (i_s0_23_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_24_1__core_periphery__clock_from_core                      (i_s0_24_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_25_1__core_periphery__clock_from_core                      (i_s0_25_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_30_1__core_periphery__clock_from_core                      (i_s0_30_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_31_1__core_periphery__clock_from_core                      (i_s0_31_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_36_1__core_periphery__clock_from_core                      (i_s0_36_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_37_1__core_periphery__clock_from_core                      (i_s0_37_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_38_1__core_periphery__clock_from_core                      (i_s0_38_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_43_1__core_periphery__clock_from_core                      (i_s0_43_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_44_1__core_periphery__clock_from_core                      (i_s0_44_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_45_1__core_periphery__clock_from_core                      (i_s0_45_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_46_1__core_periphery__clock_from_core                      (i_s0_46_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_47_1__core_periphery__clock_from_core                      (i_s0_47_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_48_1__core_periphery__clock_from_core                      (i_s0_48_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_49_1__core_periphery__clock_from_core                      (i_s0_49_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_50_1__core_periphery__clock_from_core                      (i_s0_50_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_55_1__core_periphery__clock_from_core                      (i_s0_55_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_56_1__core_periphery__clock_from_core                      (i_s0_56_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_57_1__core_periphery__clock_from_core                      (i_s0_57_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_62_1__core_periphery__clock_from_core                      (i_s0_62_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_63_1__core_periphery__clock_from_core                      (i_s0_63_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_68_1__core_periphery__clock_from_core                      (i_s0_68_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_69_1__core_periphery__clock_from_core                      (i_s0_69_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_70_1__core_periphery__clock_from_core                      (i_s0_70_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_71_1__core_periphery__clock_from_core                      (i_s0_71_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_72_1__core_periphery__clock_from_core                      (i_s0_72_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_77_1__core_periphery__clock_from_core                      (i_s0_77_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_78_1__core_periphery__clock_from_core                      (i_s0_78_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_83_1__core_periphery__clock_from_core                      (i_s0_83_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_84_1__core_periphery__clock_from_core                      (i_s0_84_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_85_1__core_periphery__clock_from_core                      (i_s0_85_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_90_1__core_periphery__clock_from_core                      (i_s0_90_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_91_1__core_periphery__clock_from_core                      (i_s0_91_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_92_1__core_periphery__clock_from_core                      (i_s0_92_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_93_1__core_periphery__clock_from_core                      (i_s0_93_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_94_1__core_periphery__clock_from_core                      (i_s0_94_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_95_1__core_periphery__clock_from_core                      (i_s0_95_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_96_1__core_periphery__clock_from_core                      (i_s0_96_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_97_1__core_periphery__clock_from_core                      (i_s0_97_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_102_1__core_periphery__clock_from_core                     (i_s0_102_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_103_1__core_periphery__clock_from_core                     (i_s0_103_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_104_1__core_periphery__clock_from_core                     (i_s0_104_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_109_1__core_periphery__clock_from_core                     (i_s0_109_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_110_1__core_periphery__clock_from_core                     (i_s0_110_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_115_1__core_periphery__clock_from_core                     (i_s0_115_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_116_1__core_periphery__clock_from_core                     (i_s0_116_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_117_1__core_periphery__clock_from_core                     (i_s0_117_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_118_1__core_periphery__clock_from_core                     (i_s0_118_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_119_1__core_periphery__clock_from_core                     (i_s0_119_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_124_1__core_periphery__clock_from_core                     (i_s0_124_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_125_1__core_periphery__clock_from_core                     (i_s0_125_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_130_1__core_periphery__clock_from_core                     (i_s0_130_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_131_1__core_periphery__clock_from_core                     (i_s0_131_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_132_1__core_periphery__clock_from_core                     (i_s0_132_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_137_1__core_periphery__clock_from_core                     (i_s0_137_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_138_1__core_periphery__clock_from_core                     (i_s0_138_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_139_1__core_periphery__clock_from_core                     (i_s0_139_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_140_1__core_periphery__clock_from_core                     (i_s0_140_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_141_1__core_periphery__clock_from_core                     (i_s0_141_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_142_1__core_periphery__clock_from_core                     (i_s0_142_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_143_1__core_periphery__clock_from_core                     (i_s0_143_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_144_1__core_periphery__clock_from_core                     (i_s0_144_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_149_1__core_periphery__clock_from_core                     (i_s0_149_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_150_1__core_periphery__clock_from_core                     (i_s0_150_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_151_1__core_periphery__clock_from_core                     (i_s0_151_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_156_1__core_periphery__clock_from_core                     (i_s0_156_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_157_1__core_periphery__clock_from_core                     (i_s0_157_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_162_1__core_periphery__clock_from_core                     (i_s0_162_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_163_1__core_periphery__clock_from_core                     (i_s0_163_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_164_1__core_periphery__clock_from_core                     (i_s0_164_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_165_1__core_periphery__clock_from_core                     (i_s0_165_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_166_1__core_periphery__clock_from_core                     (i_s0_166_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_171_1__core_periphery__clock_from_core                     (i_s0_171_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_172_1__core_periphery__clock_from_core                     (i_s0_172_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_177_1__core_periphery__clock_from_core                     (i_s0_177_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_178_1__core_periphery__clock_from_core                     (i_s0_178_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_179_1__core_periphery__clock_from_core                     (i_s0_179_1__core_periphery__clock_from_core),
/* input  [15:0] */ .i_s0_184_1__core_periphery__clock_from_core                     (i_s0_184_1__core_periphery__clock_from_core),
/* input  [95:0] */ .i_s0_3_1__core_periphery__data_from_core                        (i_s0_3_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_9_1__core_periphery__data_from_core                        (i_s0_9_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_10_1__core_periphery__data_from_core                       (i_s0_10_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_15_1__core_periphery__data_from_core                       (i_s0_15_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_16_1__core_periphery__data_from_core                       (i_s0_16_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_21_1__core_periphery__data_from_core                       (i_s0_21_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_22_1__core_periphery__data_from_core                       (i_s0_22_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_23_1__core_periphery__data_from_core                       (i_s0_23_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_24_1__core_periphery__data_from_core                       (i_s0_24_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_25_1__core_periphery__data_from_core                       (i_s0_25_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_30_1__core_periphery__data_from_core                       (i_s0_30_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_31_1__core_periphery__data_from_core                       (i_s0_31_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_36_1__core_periphery__data_from_core                       (i_s0_36_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_37_1__core_periphery__data_from_core                       (i_s0_37_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_38_1__core_periphery__data_from_core                       (i_s0_38_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_43_1__core_periphery__data_from_core                       (i_s0_43_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_44_1__core_periphery__data_from_core                       (i_s0_44_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_45_1__core_periphery__data_from_core                       (i_s0_45_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_46_1__core_periphery__data_from_core                       (i_s0_46_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_47_1__core_periphery__data_from_core                       (i_s0_47_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_48_1__core_periphery__data_from_core                       (i_s0_48_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_49_1__core_periphery__data_from_core                       (i_s0_49_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_50_1__core_periphery__data_from_core                       (i_s0_50_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_55_1__core_periphery__data_from_core                       (i_s0_55_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_56_1__core_periphery__data_from_core                       (i_s0_56_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_57_1__core_periphery__data_from_core                       (i_s0_57_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_62_1__core_periphery__data_from_core                       (i_s0_62_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_63_1__core_periphery__data_from_core                       (i_s0_63_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_68_1__core_periphery__data_from_core                       (i_s0_68_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_69_1__core_periphery__data_from_core                       (i_s0_69_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_70_1__core_periphery__data_from_core                       (i_s0_70_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_71_1__core_periphery__data_from_core                       (i_s0_71_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_72_1__core_periphery__data_from_core                       (i_s0_72_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_77_1__core_periphery__data_from_core                       (i_s0_77_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_78_1__core_periphery__data_from_core                       (i_s0_78_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_83_1__core_periphery__data_from_core                       (i_s0_83_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_84_1__core_periphery__data_from_core                       (i_s0_84_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_90_1__core_periphery__data_from_core                       (i_s0_90_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_91_1__core_periphery__data_from_core                       (i_s0_91_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_92_1__core_periphery__data_from_core                       (i_s0_92_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_93_1__core_periphery__data_from_core                       (i_s0_93_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_94_1__core_periphery__data_from_core                       (i_s0_94_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_95_1__core_periphery__data_from_core                       (i_s0_95_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_96_1__core_periphery__data_from_core                       (i_s0_96_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_97_1__core_periphery__data_from_core                       (i_s0_97_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_102_1__core_periphery__data_from_core                      (i_s0_102_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_103_1__core_periphery__data_from_core                      (i_s0_103_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_104_1__core_periphery__data_from_core                      (i_s0_104_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_109_1__core_periphery__data_from_core                      (i_s0_109_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_110_1__core_periphery__data_from_core                      (i_s0_110_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_115_1__core_periphery__data_from_core                      (i_s0_115_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_116_1__core_periphery__data_from_core                      (i_s0_116_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_117_1__core_periphery__data_from_core                      (i_s0_117_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_118_1__core_periphery__data_from_core                      (i_s0_118_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_119_1__core_periphery__data_from_core                      (i_s0_119_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_124_1__core_periphery__data_from_core                      (i_s0_124_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_125_1__core_periphery__data_from_core                      (i_s0_125_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_130_1__core_periphery__data_from_core                      (i_s0_130_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_131_1__core_periphery__data_from_core                      (i_s0_131_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_132_1__core_periphery__data_from_core                      (i_s0_132_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_137_1__core_periphery__data_from_core                      (i_s0_137_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_138_1__core_periphery__data_from_core                      (i_s0_138_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_139_1__core_periphery__data_from_core                      (i_s0_139_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_140_1__core_periphery__data_from_core                      (i_s0_140_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_141_1__core_periphery__data_from_core                      (i_s0_141_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_142_1__core_periphery__data_from_core                      (i_s0_142_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_143_1__core_periphery__data_from_core                      (i_s0_143_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_144_1__core_periphery__data_from_core                      (i_s0_144_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_149_1__core_periphery__data_from_core                      (i_s0_149_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_150_1__core_periphery__data_from_core                      (i_s0_150_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_151_1__core_periphery__data_from_core                      (i_s0_151_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_156_1__core_periphery__data_from_core                      (i_s0_156_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_157_1__core_periphery__data_from_core                      (i_s0_157_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_162_1__core_periphery__data_from_core                      (i_s0_162_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_163_1__core_periphery__data_from_core                      (i_s0_163_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_164_1__core_periphery__data_from_core                      (i_s0_164_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_165_1__core_periphery__data_from_core                      (i_s0_165_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_166_1__core_periphery__data_from_core                      (i_s0_166_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_171_1__core_periphery__data_from_core                      (i_s0_171_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_172_1__core_periphery__data_from_core                      (i_s0_172_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_177_1__core_periphery__data_from_core                      (i_s0_177_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_178_1__core_periphery__data_from_core                      (i_s0_178_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_179_1__core_periphery__data_from_core                      (i_s0_179_1__core_periphery__data_from_core),
/* input  [95:0] */ .i_s0_184_1__core_periphery__data_from_core                      (i_s0_184_1__core_periphery__data_from_core),
/* input  [13:0] */ .s0_100_1__core_periphery__clock_from_core_unused                (s0_100_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_100_1__core_periphery__data_from_core_unused                 (s0_100_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_101_1__core_periphery__clock_from_core_unused                (s0_101_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_101_1__core_periphery__data_from_core_unused                 (s0_101_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_105_1__core_periphery__clock_from_core_unused                (s0_105_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_105_1__core_periphery__data_from_core_unused                 (s0_105_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_106_1__core_periphery__clock_from_core_unused                (s0_106_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_106_1__core_periphery__data_from_core_unused                 (s0_106_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_107_1__core_periphery__clock_from_core_unused                (s0_107_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_107_1__core_periphery__data_from_core_unused                 (s0_107_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_108_1__core_periphery__clock_from_core_unused                (s0_108_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_108_1__core_periphery__data_from_core_unused                 (s0_108_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_111_1__core_periphery__clock_from_core_unused                (s0_111_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_111_1__core_periphery__data_from_core_unused                 (s0_111_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_112_1__core_periphery__clock_from_core_unused                (s0_112_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_112_1__core_periphery__data_from_core_unused                 (s0_112_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_113_1__core_periphery__clock_from_core_unused                (s0_113_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_113_1__core_periphery__data_from_core_unused                 (s0_113_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_114_1__core_periphery__clock_from_core_unused                (s0_114_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_114_1__core_periphery__data_from_core_unused                 (s0_114_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_11_1__core_periphery__clock_from_core_unused                 (s0_11_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_11_1__core_periphery__data_from_core_unused                  (s0_11_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_120_1__core_periphery__clock_from_core_unused                (s0_120_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_120_1__core_periphery__data_from_core_unused                 (s0_120_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_121_1__core_periphery__clock_from_core_unused                (s0_121_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_121_1__core_periphery__data_from_core_unused                 (s0_121_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_122_1__core_periphery__clock_from_core_unused                (s0_122_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_122_1__core_periphery__data_from_core_unused                 (s0_122_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_123_1__core_periphery__clock_from_core_unused                (s0_123_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_123_1__core_periphery__data_from_core_unused                 (s0_123_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_126_1__core_periphery__clock_from_core_unused                (s0_126_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_126_1__core_periphery__data_from_core_unused                 (s0_126_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_127_1__core_periphery__clock_from_core_unused                (s0_127_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_127_1__core_periphery__data_from_core_unused                 (s0_127_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_128_1__core_periphery__clock_from_core_unused                (s0_128_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_128_1__core_periphery__data_from_core_unused                 (s0_128_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_129_1__core_periphery__clock_from_core_unused                (s0_129_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_129_1__core_periphery__data_from_core_unused                 (s0_129_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_12_1__core_periphery__clock_from_core_unused                 (s0_12_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_12_1__core_periphery__data_from_core_unused                  (s0_12_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_133_1__core_periphery__clock_from_core_unused                (s0_133_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_133_1__core_periphery__data_from_core_unused                 (s0_133_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_134_1__core_periphery__clock_from_core_unused                (s0_134_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_134_1__core_periphery__data_from_core_unused                 (s0_134_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_135_1__core_periphery__clock_from_core_unused                (s0_135_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_135_1__core_periphery__data_from_core_unused                 (s0_135_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_136_1__core_periphery__clock_from_core_unused                (s0_136_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_136_1__core_periphery__data_from_core_unused                 (s0_136_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_13_1__core_periphery__clock_from_core_unused                 (s0_13_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_13_1__core_periphery__data_from_core_unused                  (s0_13_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_145_1__core_periphery__clock_from_core_unused                (s0_145_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_145_1__core_periphery__data_from_core_unused                 (s0_145_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_146_1__core_periphery__clock_from_core_unused                (s0_146_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_146_1__core_periphery__data_from_core_unused                 (s0_146_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_147_1__core_periphery__clock_from_core_unused                (s0_147_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_147_1__core_periphery__data_from_core_unused                 (s0_147_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_148_1__core_periphery__clock_from_core_unused                (s0_148_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_148_1__core_periphery__data_from_core_unused                 (s0_148_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_14_1__core_periphery__clock_from_core_unused                 (s0_14_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_14_1__core_periphery__data_from_core_unused                  (s0_14_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_152_1__core_periphery__clock_from_core_unused                (s0_152_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_152_1__core_periphery__data_from_core_unused                 (s0_152_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_153_1__core_periphery__clock_from_core_unused                (s0_153_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_153_1__core_periphery__data_from_core_unused                 (s0_153_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_154_1__core_periphery__clock_from_core_unused                (s0_154_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_154_1__core_periphery__data_from_core_unused                 (s0_154_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_155_1__core_periphery__clock_from_core_unused                (s0_155_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_155_1__core_periphery__data_from_core_unused                 (s0_155_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_158_1__core_periphery__clock_from_core_unused                (s0_158_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_158_1__core_periphery__data_from_core_unused                 (s0_158_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_159_1__core_periphery__clock_from_core_unused                (s0_159_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_159_1__core_periphery__data_from_core_unused                 (s0_159_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_160_1__core_periphery__clock_from_core_unused                (s0_160_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_160_1__core_periphery__data_from_core_unused                 (s0_160_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_161_1__core_periphery__clock_from_core_unused                (s0_161_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_161_1__core_periphery__data_from_core_unused                 (s0_161_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_167_1__core_periphery__clock_from_core_unused                (s0_167_1__core_periphery__clock_from_core_unused),
/* input  [72:0] */ .s0_167_1__core_periphery__data_from_core_unused                 (s0_167_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_168_1__core_periphery__clock_from_core_unused                (s0_168_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_168_1__core_periphery__data_from_core_unused                 (s0_168_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_169_1__core_periphery__clock_from_core_unused                (s0_169_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_169_1__core_periphery__data_from_core_unused                 (s0_169_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_170_1__core_periphery__clock_from_core_unused                (s0_170_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_170_1__core_periphery__data_from_core_unused                 (s0_170_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_173_1__core_periphery__clock_from_core_unused                (s0_173_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_173_1__core_periphery__data_from_core_unused                 (s0_173_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_174_1__core_periphery__clock_from_core_unused                (s0_174_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_174_1__core_periphery__data_from_core_unused                 (s0_174_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_175_1__core_periphery__clock_from_core_unused                (s0_175_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_175_1__core_periphery__data_from_core_unused                 (s0_175_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_176_1__core_periphery__clock_from_core_unused                (s0_176_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_176_1__core_periphery__data_from_core_unused                 (s0_176_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_17_1__core_periphery__clock_from_core_unused                 (s0_17_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_17_1__core_periphery__data_from_core_unused                  (s0_17_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_180_1__core_periphery__clock_from_core_unused                (s0_180_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_180_1__core_periphery__data_from_core_unused                 (s0_180_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_181_1__core_periphery__clock_from_core_unused                (s0_181_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_181_1__core_periphery__data_from_core_unused                 (s0_181_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_182_1__core_periphery__clock_from_core_unused                (s0_182_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_182_1__core_periphery__data_from_core_unused                 (s0_182_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_183_1__core_periphery__clock_from_core_unused                (s0_183_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_183_1__core_periphery__data_from_core_unused                 (s0_183_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_18_1__core_periphery__clock_from_core_unused                 (s0_18_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_18_1__core_periphery__data_from_core_unused                  (s0_18_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_19_1__core_periphery__clock_from_core_unused                 (s0_19_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_19_1__core_periphery__data_from_core_unused                  (s0_19_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_20_1__core_periphery__clock_from_core_unused                 (s0_20_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_20_1__core_periphery__data_from_core_unused                  (s0_20_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_26_1__core_periphery__clock_from_core_unused                 (s0_26_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_26_1__core_periphery__data_from_core_unused                  (s0_26_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_27_1__core_periphery__clock_from_core_unused                 (s0_27_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_27_1__core_periphery__data_from_core_unused                  (s0_27_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_28_1__core_periphery__clock_from_core_unused                 (s0_28_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_28_1__core_periphery__data_from_core_unused                  (s0_28_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_29_1__core_periphery__clock_from_core_unused                 (s0_29_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_29_1__core_periphery__data_from_core_unused                  (s0_29_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_32_1__core_periphery__clock_from_core_unused                 (s0_32_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_32_1__core_periphery__data_from_core_unused                  (s0_32_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_33_1__core_periphery__clock_from_core_unused                 (s0_33_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_33_1__core_periphery__data_from_core_unused                  (s0_33_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_34_1__core_periphery__clock_from_core_unused                 (s0_34_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_34_1__core_periphery__data_from_core_unused                  (s0_34_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_35_1__core_periphery__clock_from_core_unused                 (s0_35_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_35_1__core_periphery__data_from_core_unused                  (s0_35_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_39_1__core_periphery__clock_from_core_unused                 (s0_39_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_39_1__core_periphery__data_from_core_unused                  (s0_39_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_40_1__core_periphery__clock_from_core_unused                 (s0_40_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_40_1__core_periphery__data_from_core_unused                  (s0_40_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_41_1__core_periphery__clock_from_core_unused                 (s0_41_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_41_1__core_periphery__data_from_core_unused                  (s0_41_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_42_1__core_periphery__clock_from_core_unused                 (s0_42_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_42_1__core_periphery__data_from_core_unused                  (s0_42_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_4_1__core_periphery__clock_from_core_unused                  (s0_4_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_4_1__core_periphery__data_from_core_unused                   (s0_4_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_51_1__core_periphery__clock_from_core_unused                 (s0_51_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_51_1__core_periphery__data_from_core_unused                  (s0_51_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_52_1__core_periphery__clock_from_core_unused                 (s0_52_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_52_1__core_periphery__data_from_core_unused                  (s0_52_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_53_1__core_periphery__clock_from_core_unused                 (s0_53_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_53_1__core_periphery__data_from_core_unused                  (s0_53_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_54_1__core_periphery__clock_from_core_unused                 (s0_54_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_54_1__core_periphery__data_from_core_unused                  (s0_54_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_58_1__core_periphery__clock_from_core_unused                 (s0_58_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_58_1__core_periphery__data_from_core_unused                  (s0_58_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_59_1__core_periphery__clock_from_core_unused                 (s0_59_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_59_1__core_periphery__data_from_core_unused                  (s0_59_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_5_1__core_periphery__clock_from_core_unused                  (s0_5_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_5_1__core_periphery__data_from_core_unused                   (s0_5_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_60_1__core_periphery__clock_from_core_unused                 (s0_60_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_60_1__core_periphery__data_from_core_unused                  (s0_60_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_61_1__core_periphery__clock_from_core_unused                 (s0_61_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_61_1__core_periphery__data_from_core_unused                  (s0_61_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_64_1__core_periphery__clock_from_core_unused                 (s0_64_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_64_1__core_periphery__data_from_core_unused                  (s0_64_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_65_1__core_periphery__clock_from_core_unused                 (s0_65_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_65_1__core_periphery__data_from_core_unused                  (s0_65_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_66_1__core_periphery__clock_from_core_unused                 (s0_66_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_66_1__core_periphery__data_from_core_unused                  (s0_66_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_67_1__core_periphery__clock_from_core_unused                 (s0_67_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_67_1__core_periphery__data_from_core_unused                  (s0_67_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_6_1__core_periphery__clock_from_core_unused                  (s0_6_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_6_1__core_periphery__data_from_core_unused                   (s0_6_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_73_1__core_periphery__clock_from_core_unused                 (s0_73_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_73_1__core_periphery__data_from_core_unused                  (s0_73_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_74_1__core_periphery__clock_from_core_unused                 (s0_74_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_74_1__core_periphery__data_from_core_unused                  (s0_74_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_75_1__core_periphery__clock_from_core_unused                 (s0_75_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_75_1__core_periphery__data_from_core_unused                  (s0_75_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_76_1__core_periphery__clock_from_core_unused                 (s0_76_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_76_1__core_periphery__data_from_core_unused                  (s0_76_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_79_1__core_periphery__clock_from_core_unused                 (s0_79_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_79_1__core_periphery__data_from_core_unused                  (s0_79_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_7_1__core_periphery__clock_from_core_unused                  (s0_7_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_7_1__core_periphery__data_from_core_unused                   (s0_7_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_80_1__core_periphery__clock_from_core_unused                 (s0_80_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_80_1__core_periphery__data_from_core_unused                  (s0_80_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_81_1__core_periphery__clock_from_core_unused                 (s0_81_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_81_1__core_periphery__data_from_core_unused                  (s0_81_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_82_1__core_periphery__clock_from_core_unused                 (s0_82_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_82_1__core_periphery__data_from_core_unused                  (s0_82_1__core_periphery__data_from_core_unused),
/* input  [93:0] */ .s0_85_1__core_periphery__data_from_core_unused                  (s0_85_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_86_1__core_periphery__clock_from_core_unused                 (s0_86_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_86_1__core_periphery__data_from_core_unused                  (s0_86_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_87_1__core_periphery__clock_from_core_unused                 (s0_87_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_87_1__core_periphery__data_from_core_unused                  (s0_87_1__core_periphery__data_from_core_unused),
/* input  [13:0] */ .s0_88_1__core_periphery__clock_from_core_unused                 (s0_88_1__core_periphery__clock_from_core_unused),
/* input  [21:0] */ .s0_88_1__core_periphery__data_from_core_unused                  (s0_88_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_89_1__core_periphery__clock_from_core_unused                 (s0_89_1__core_periphery__clock_from_core_unused),
/* input  [66:0] */ .s0_89_1__core_periphery__data_from_core_unused                  (s0_89_1__core_periphery__data_from_core_unused),
/* input  [64:0] */ .s0_8_1__core_periphery__data_from_core_unused                   (s0_8_1__core_periphery__data_from_core_unused),
/* input  [14:0] */ .s0_98_1__core_periphery__clock_from_core_unused                 (s0_98_1__core_periphery__clock_from_core_unused),
/* input  [59:0] */ .s0_98_1__core_periphery__data_from_core_unused                  (s0_98_1__core_periphery__data_from_core_unused),
/* input  [9:0]  */ .s0_99_1__core_periphery__clock_from_core_unused                 (s0_99_1__core_periphery__clock_from_core_unused),
/* input  [34:0] */ .s0_99_1__core_periphery__data_from_core_unused                  (s0_99_1__core_periphery__data_from_core_unused),
/* input         */ .vcc_dts_ref                                                     (vcc_dts_ref),
/* input         */ .vcce_pll_ref                                                    (vcce_pll_ref),


		.p0_app_err_valid_i		(p0_app_err_valid_i),
		.p0_app_err_hdr_i			(p0_app_err_hdr_i),
		.p0_app_err_info_i			(p0_app_err_info_i),
		.p0_app_err_func_num_i		(p0_app_err_func_num_i),
                .p0_app_err_vfa_i               (p0_app_err_vfa_i),
                .p0_app_err_vf_num_i            (p0_app_err_vf_num_i),

		.p0_app_err_ready_o		(p0_app_err_ready_o),
		.p0_cpl_timeout_o			(p0_cpl_timeout_o),
		.p0_cpl_timeout_func_num_o		(p0_cpl_timeout_func_num_o),
		.p0_cpl_timeout_vfunc_num_o	(p0_cpl_timeout_vfunc_num_o),
		.p0_cpl_timeout_vfunc_active_o	(p0_cpl_timeout_vfunc_active_o),
		.p0_cpl_timeout_cpl_tc_o		(p0_cpl_timeout_cpl_tc_o),
		.p0_cpl_timeout_cpl_attr_o		(p0_cpl_timeout_cpl_attr_o),
		.p0_cpl_timeout_cpl_len_o		(p0_cpl_timeout_cpl_len_o),
		.p0_cpl_timeout_cpl_tag_o		(p0_cpl_timeout_cpl_tag_o),
		.p0_flr_rcvd_pf_o			(p0_flr_rcvd_pf_o),
		.p0_flr_rcvd_vf_o			(p0_flr_rcvd_vf_o),
		.p0_flr_rcvd_pf_num_o		(p0_flr_rcvd_pf_num_o),
		.p0_flr_rcvd_vf_num_o		(p0_flr_rcvd_vf_num_o),
		.p0_flr_completed_pf_i		(p0_flr_completed_pf_i),
		.p0_flr_completed_vf_i		(p0_flr_completed_vf_i),
		.p0_flr_completed_pf_num_i		(p0_flr_completed_pf_num_i),
		.p0_flr_completed_vf_num_i		(p0_flr_completed_vf_num_i),
		.p0_flr_completed_ready_o		(p0_flr_completed_ready_o),
		.p0_cii_req_o			(p0_cii_req_o),
		.p0_cii_hdr_poisoned_o		(p0_cii_hdr_poisoned_o),
		.p0_cii_hdr_first_be_o		(p0_cii_hdr_first_be_o),
		.p0_cii_func_num_o			(p0_cii_func_num_o),
		.p0_cii_wr_vf_active_o		(p0_cii_wr_vf_active_o),
		.p0_cii_vf_num_o			(p0_cii_vf_num_o),
		.p0_cii_wr_o			(p0_cii_wr_o),
		.p0_cii_addr_o			(p0_cii_addr_o),
		.p0_cii_dout_o			(p0_cii_dout_o),
		.p0_cii_override_en_i		(p0_cii_override_en_i),
		.p0_cii_override_din_i		(p0_cii_override_din_i),
		.p0_cii_halt_i			(p0_cii_halt_i),
                .p0_cii_convert_pfd_i           (p0_cii_convert_pfd_i),
                .p0_cii_conv_pfdata_i           (p0_cii_conv_pfdata_i),
                .p0_pci_cfg_req_o              (p0_pci_cfg_req_o),
                .p0_pci_cfg_func_num_o         (p0_pci_cfg_func_num_o),
                .p0_pci_cfg_len_o              (p0_pci_cfg_len_o),
                .p0_pci_cfg_bar_o              (p0_pci_cfg_bar_o),
                .p0_pci_cfg_offset_o           (p0_pci_cfg_offset_o),
                .p0_pci_cfg_wr_o               (p0_pci_cfg_wr_o),
                .p0_pci_cfg_writedata_o        (p0_pci_cfg_writedata_o),
                .p0_pci_cfg_readdata_i         (p0_pci_cfg_readdata_i),
                .p0_pci_cfg_tag_o              (p0_pci_cfg_tag_o),
                .p0_pci_cfg_be_o               (p0_pci_cfg_be_o),
                .p0_pci_cfg_ack_i              (p0_pci_cfg_ack_i),
                .p0_pci_cfg_df_i               (p0_pci_cfg_df_i),
                .p0_pci_cfg_status_i           (p0_pci_cfg_status_i),
		.p0_hip_reconfig_address_i		(p0_hip_reconfig_address_i),
		.p0_hip_reconfig_write_i		(p0_hip_reconfig_write_i),
                .p0_hip_reconfig_writedata_i           (p0_hip_reconfig_writedata_i),
                .p0_hip_reconfig_read_i                 (p0_hip_reconfig_read_i),
                .p0_hip_reconfig_readdatavalid_o        (p0_hip_reconfig_readdatavalid_o),
                .p0_hip_reconfig_readdata_o             (p0_hip_reconfig_readdata_o),
                .p0_hip_reconfig_waitrequest_o          (p0_hip_reconfig_waitrequest_o),
                .p0_hip_reconfig_resp_o            (p0_hip_reconfig_resp_o),
                .p0_hip_reconfig_requesttype_i          (p0_hip_reconfig_requesttype_i),
////            .p0_dbg_mmio_address            (p0_dbg_mmio_address),
////            .p0_dbg_mmio_write                      (p0_dbg_mmio_write),
////            .p0_dbg_mmio_writedata          (p0_dbg_mmio_writedata),
////            .p0_dbg_mmio_read                       (p0_dbg_mmio_read),
////            .p0_dbg_mmio_readdatavalid              (p0_dbg_mmio_readdatavalid),
////            .p0_dbg_mmio_readdata           (p0_dbg_mmio_readdata),
////            .p0_dbg_mmio_waitrequest                (p0_dbg_mmio_waitrequest),
		.p0_pm_valid_i			(p0_pm_valid_i),
                .p0_pm_opcode_i		(p0_pm_opcode_i),
                .p0_pm_tag_i			(p0_pm_tag_i),
                .p0_pm_misc_i			(p0_pm_misc_i),
                .p0_pm_data_i			(p0_pm_data_i),
    		.p0_pm_valid_o			(p0_pm_valid_o),
    		.p0_pm_opcode_o		(p0_pm_opcode_o),
    		.p0_pm_tag_o			(p0_pm_tag_o),
    		.p0_pm_misc_o			(p0_pm_misc_o),
    		.p0_pm_data_o			(p0_pm_data_o),
    		.p0_aermsg_correctable_valid_o	(p0_aermsg_correctable_valid_o),
    		.p0_aermsg_uncorrectable_valid_o(p0_aermsg_uncorrectable_valid_o),
    		.p0_aermsg_res_o		(p0_aermsg_res_o),
    		.p0_aermsg_bts_o		(p0_aermsg_bts_o),
    		.p0_aermsg_bds_o		(p0_aermsg_bds_o),
    		.p0_aermsg_rrs_o		(p0_aermsg_rrs_o),
    		.p0_aermsg_rtts_o		(p0_aermsg_rtts_o),
    		.p0_aermsg_anes_o		(p0_aermsg_anes_o),
    		.p0_aermsg_cies_o		(p0_aermsg_cies_o),
    		.p0_aermsg_hlos_o		(p0_aermsg_hlos_o),
    		.p0_aermsg_fmt_o		(p0_aermsg_fmt_o),
    		.p0_aermsg_type_o		(p0_aermsg_type_o),
    		.p0_aermsg_tc_o		(p0_aermsg_tc_o),
    		.p0_aermsg_ido_o		(p0_aermsg_ido_o),
    		.p0_aermsg_th_o		(p0_aermsg_th_o),
    		.p0_aermsg_td_o		(p0_aermsg_td_o),
    		.p0_aermsg_ep_o		(p0_aermsg_ep_o),
    		.p0_aermsg_ro_o		(p0_aermsg_ro_o ),
    		.p0_aermsg_ns_o		(p0_aermsg_ns_o),
    		.p0_aermsg_at_o		(p0_aermsg_at_o),
    		.p0_aermsg_length_o		(p0_aermsg_length_o),
    		.p0_aermsg_header_o		(p0_aermsg_header_o),
    		.p0_aermsg_und_o		(p0_aermsg_und_o),
    		.p0_aermsg_anf_o		(p0_aermsg_anf_o),
    		.p0_aermsg_dlpes_o		(p0_aermsg_dlpes_o),
    		.p0_aermsg_sdes_o		(p0_aermsg_sdes_o),
    		.p0_aermsg_fep_o		(p0_aermsg_fep_o),
    		.p0_aermsg_pts_o		(p0_aermsg_pts_o),
    		.p0_aermsg_fcpes_o		(p0_aermsg_fcpes_o),
    		.p0_aermsg_cts_o		(p0_aermsg_cts_o),
    		.p0_aermsg_cas_o		(p0_aermsg_cas_o),
    		.p0_aermsg_ucs_o		(p0_aermsg_ucs_o),
    		.p0_aermsg_ros_o		(p0_aermsg_ros_o),
    		.p0_aermsg_mts_o		(p0_aermsg_mts_o),
    		.p0_aermsg_uies_o		(p0_aermsg_uies_o),
    		.p0_aermsg_mbts_o		(p0_aermsg_mbts_o),
    		.p0_aermsg_aebs_o		(p0_aermsg_aebs_o),
    		.p0_aermsg_tpbes_o		(p0_aermsg_tpbes_o),
    		.p0_aermsg_ees_o		(p0_aermsg_ees_o),
    		.p0_aermsg_ures_o		(p0_aermsg_ures_o),
    		.p0_aermsg_avs_o		(p0_aermsg_avs_o),
    		.p0_cfgupdate_valid_o		(p0_cfgupdate_valid_o),
    		.p0_cfgupdate_regtype_o	(p0_cfgupdate_regtype_o),
    		.p0_cfgupdate_vfa_o		(p0_cfgupdate_vfa_o),
    		.p0_cfgupdate_pfnum_o		(p0_cfgupdate_pfnum_o),
    		.p0_cfgupdate_vfnum_o		(p0_cfgupdate_vfnum_o),
    		.p0_cfgupdate_info_o		(p0_cfgupdate_info_o),
    		.p0_hip_err_valid_o		(p0_hip_err_valid_o),
    		.p0_hip_err_hdr_o		(p0_hip_err_hdr_o),
    		.p0_hip_err_info_o		(p0_hip_err_info_o),
    		.p0_hip_err_pf_num_o		(p0_hip_err_pf_num_o),
    		.p0_hip_err_vfa_o		(p0_hip_err_vfa_o),
    		.p0_hip_err_vf_num_o		(p0_hip_err_vf_num_o),
    		.cache_mem_crd_flow_err_o	(cache_mem_crd_flow_err_o)

);

// Simulation requires all params from lampas
`ifndef ALTERA_RESERVED_QIS
`include "./rtile_cxl_settings.svh"
`endif
endmodule
module  altera_s10_configuration_clock
     (
     clkout
     );
 
     parameter DEVICE_FAMILY   = " Stratix 10";
 
     output   clkout;
 
 
 
//synthesis read_comments_as_HDL on
//     wire  wire_clkout;
//     altera_config_clock_source_endpoint s10_config_clk_inst (
//         .clk        (wire_clkout)
//     );
//synthesis read_comments_as_HDL off

//synthesis translate_off 
    localparam CLOCK_PERIOD = 4;
    localparam HALF_CLOCK_PERIOD = CLOCK_PERIOD/2;                                                                                                                               
    reg  wire_clkout;
    initial begin
        wire_clkout <= 1'b1;
        forever #HALF_CLOCK_PERIOD wire_clkout <= ~wire_clkout; // most efficient method for sim speed      
    end
//synthesis translate_on 

     assign clkout = wire_clkout;
endmodule //altera_int_osc

