// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vRgucS1vE19aPhObcq5AFs183Ue8yVSNap5PIMqslPZggZNquVyxcCWaQdNl
Sbbm0+uutDt3ua1MlAVHuNg8vLxU0JiYnTGH0W9hW6zZ5w6y6uMQTA2pWSLV
t5/LnhbNvzGQe9tlXh3litxmaB7T5/c5By2fJkV7wMdHlBqIgMpnEusCftZl
GOv2uOHqaPMmR8/aeZ/gi/5Knnbz59kd5/CLl50jkQnvGgIA/9YDE3Uy+frz
A8pAEFQgyh+hug38yU5xmYmsYxHXQlIMq/3nS6J/i8PBLqb9hVT8edK6WmBf
IG9heCQ9L6jeg1Oqk5OTm907CSoiN4diuogbIFbgwg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I1SqZQ64BqPBu5U0of0rca361NWVQB3NzTP9yBW14w63fbObUw/xlV1kLj8R
cBBJoqDwCvpdTLJj4JK3YID7uh66WdTL6DJAaF+aCo3W0g2kY18JZ2XVAqCl
wV1FBRYyYVRQv7+1Ev55FhfXoUHQcTxq9wYGqenYz8DImBebsarw3A7RWw1R
Y0ZkPfUOtgt8L/+rutPYDTkm26fJaVyOIfnn/ypdmVacTjvxba/sH6QOh/KE
xqNJB/Q957GRyiPhTSn2FBIi438A5CGkIRRSVZ2Mjb5OoRLrUyl7N5R8m+NU
djpcNN6m59zqXRdh2JYF0AlKrA1TteFp/igujle8qA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aIug24uCoEC2JtYPICq4L80Y0s7cLJnCb+FHWQ3cY9Y8VJzqp+I/xRH7MHr/
8XslS7KpaN4Hbke/Ewse+JLiPeRdopSuF++5MR9UzmmOt7LP9ygC6+LjkyZC
hI+ADH8Lt5ctx8E7ys5DQWz8AVQhgMeXQG3GdRT7kCHazXhmRbRUZFEYAlcs
aUJ4TvXbi1yip/ve/NzY9HtosMb+Kb9xeZee5itLt7l34UJXBYYv4QIDmJ4n
87+gKbZ0nUXWRiy6LX/ybzwopCkhwpp7F+2wmJ443b+JX/LimergpHccFEpA
t2pMBxgvcpn3vFKwwzmJI0WuiNEGxlsaHRVACbVqTA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nUZeQWfC1qaFF5TRX8oTA8pkDSrG8CastjTvtWbquxvl8xxLlUcKOBfXZo1k
asEl+wv5EvfO21/mh1qjq9h7H/9OUGHtd6EnF0dVMvt2S3bBdMp3DmwZXejc
F3WcVCL3mwL0neH3Pvijt2T9e8Vh2t2V+GlfT7o104AEG3m0cv6C2It1vvZc
hrPU4kYKvzGHpyvRQOC0IY/zrYC52jszOEhJTY5gAm30pysfbAzo1xGleUTb
8T8BKOGJu67Vj32sVg5xaXnTRSXrApk3V5lZRLI1oyjkXZIF6j8P5e1/Qyaj
7V44An6TO01XRXDN6Lqv5O4AC6s7R6N3wFKxenqRnA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fzhZQmMlEVPBpCTvuphz0CGNwXgrCBAdtlngy3Qg0W+TQ5kpYYiYicoFhTRm
0QU/3zRaR/x9HklUbI7GOvexVj1uKqc28s147bK1iSf1R5jnyLi/fuUKuHoI
BLl9iIY+IbaF1spApNYCkLa0+eVHqain6LgcZHq2aAnaoq4Njbs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mKp+04454DlOujODjpSvOVyPrMfSUiYDWuS9HJ1oGDrpwmlKC24bKEU+PZq2
snSX2zRhbt1jvVbIWghz8nPNyCxZ7JBoD6MLzB1wSKBUsqJQt4DaiHYXFDbB
AGZ8advLhD4jcI5Z6dMjIAe6e/8PBBGhfxGJjgmTslaMVvYNXfjBw1S5SXUs
CGqgjr4ntm0vCW0yBH2ixXnEB8pU2Qsvc1NG0E/pi+ItfLJ7iHdAnR3kxOzp
q0sXIMbV3euPXz4pWI+SY9eNhNqBP5/4lNV789/i5F4/6crqUbAQjVnK9F10
Ah4Y20CXZA0EhPbOV+pAWY6eSI2BAwp2+MnNY3mrjDoFtP4S+sOQl72uxDg3
OFmgJwZwdQnee29OGO7EcCH0JgDcJvb4SCpFXmLUNR6etn41D82ofvkaiPJu
F1tjlNF94/s2iboCgC3saFHGjMoPfbk8rUiQcIYpAjH655ZAenzZiRAvZj47
w1sbtVCOanCdVd5nwaXzXmYmddLI68um


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aJSPWfOYwN4bsJVU3z+DRrP4biLd85su1cHFHsfIgkdsw9FB4k1ARSDz47s2
bazCbmO7AcJ0vq4UJvUhfolgRCw21PbTkcu56Wx9TQzwFJTDGkc6eLQNR2Yf
yxR+acj6gyqXo8a7FE+TVT0M1L8fG6IgfsyQCgqhFc4auqpYTV8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Qi+D/HM+LL/tweKf3eLiQ5U6taZM7iXUMyJrkJjW75ZayT1hsZOo+qU+npO9
oRMit7i4KKhNnTK3iFFmiuz4EzG0ej4KfkqqsQF1tW0aZx4qr9AmpaVCk2yW
faoeW+6Mc7++vLQAHXbGt3P9Hk4mZXfQVkZSK2hJO2p+TRdXvXk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12432)
`pragma protect data_block
bAkjaKPFLUny2EejdHcKycco7me+r/xHx3uebbiS4mcSuC79P0RmwV2LFiBR
p+e1wqeccfyDsUa/iyucMNhsAxPETrKv5WlG/oUhWuvKDJPd60vHOlyDajiX
d45Rv4jpI4GZ8JP1dGyzXhO32rRz78neUxErw0plXGU41/STN/tSgtwHWcTC
hqJ9Dkry0OH9WvG2FMO5W8S9Yoa2SEK2cL1lgDcEE8GLtBajb7LkBJhJYyRi
5crBrj8ytkkPaIHutuyZv8nJqTRB3ARcV36YQd3ezMmMxEFNVPOnCw25a164
/NqsWs985D1FMTDVInIlIUiWyWTzh7qx2oJMHrpSm9VQMQjVmnUUtcJuF7Oe
gaa7dZYu542ipa6QJi3RnP6/GHsh3CDfI5caeJANClD494MeOShOU5pSq0WG
N0yyz+tn1AEdsVgKqwh5jiwkjtkFDFLEVSJvDef2E0Bdi/UQs/CK31J5sZPt
QjCFuWx1yHp2mTsaDV8MiQAZMrIc6vrro4Rtw0PfPZJTx1EvZewQ4i0Jtbru
lz4iejzlH59YnEbql/UGVExuSNsecE0E+OfmTsz4WctjIGz3tjSY5MyBvbFv
66bhCp2fERBsV0KvQkH5dlCtYnagR2AG8LiXA9UbEfkUt+p2svfp4b8826Yp
Ymc7tvOFyZnN5VaY9/BoRSPEmOFk+1MkDYr9yzIssKhUAgmO7qNKZTW+00OC
bf/NUO45AOS6p5PLgPLFVnFtptkzsGfVTA+t0Hj4eQ0Phdf/Up1zKnurfnyj
Ma615Y6obRLx6cE8a8UCs44+bZLdxztkB/udPlcFrYfuHSO18Sq4EfOxx2uB
SCacbGQtmpFHTblnWQLB3n4C1pbkNaa42S4yaA0al39tqyRMxMQ6fwHJZ1Bp
bFu8KCqrssIdeD7JLCZTyHu271/nOnmx2p8HzpjKah6n8PmfUNfDpgPhQ2Yq
STletCHskQsE5tzoH72wvAHIrydidrtJyrpjizOa/wR76KuClA1bpXoDNez4
9l1cDp1FyxfZ+U9zD+3ZZ7AMx3UVWZfw9zYEwqgocyzprJGsMwZ2mTmd9NNp
4n8pR5T+LmsbEgeJQPMR/F8Q+SDapqbm4w4EqHV3OKPrHkk+Al0zyeBYv8aW
ntfE0Q5yOynDWdWWdiznRvt8n+z7DcpjS1iN5rwsPsWsTmCfzVsuyHoLTkO9
aAwg41TdUcwWfKEvqB+bgVaP4oQmrZmc6VHYaow2QQeS4KrjlOtcz/ckCxg9
kDqmkL72Vi7zYN1FNXsbTqIzl4eRiLPl9uNuKpxdZnbT3iI+PJrNxg5tZEly
UT74+57Xj6rQ9SL19qiK0xuEYBOwzCO7LPxJCipwzGNrl/aqXYZjX40rsLP0
GNxWO0O0m+MPucH8DJOlE7WS44dvOzItYJyXOav7GvkkhWaFfWwAamwg7lsV
/3sCpTIqr66z7ZLENMQNUrBg8JGLkeWJ1SatnubnF/wktui+L7Xnof4uCEUs
KGCwSE0J9vy3pHeWMjFpgIzb5YM+0yWth7T7Mx60edMmtCcp8NIIHvjcDgxt
tYaoOqVTlrOIEybK7wNuAQUVpanLG7i/KEonpvangMSTmX0Cw519rVLdIDc2
svghgT/2VeXv31h+2KSdfMowmvrGXw0nlvbd85Mzv+yRotMt/L7mV3yx7gL/
1pWOE7eV0jdf9lks+i8qHjE3gNjNYg20bdAOoIlozH3LeSvsrytcA3nVFjFW
asyajXVnAWeIJ/PYQUvxzof4cJEdgYe5UoN6tx+raNeFS69VRDwBWylH/7fs
oASSCR4J3EyS+CQhnRT5mVySUgvVXebi1HFFTe84W+ZwNOtmW1b/DIT8ipQB
SYvM+5825LDjFVdeareUnpYkM4HRsz2vnDEua+OgcrA1i0Ve/JOlMpLwJx76
DOIRFvVnMrRdk7y8uYLSw8e9ZNYj6MpE7IT2q4C1JgozQUKKcXpXeaCTzrNu
MeqkJrY7fUJALIUhNJU0Wyib0vesmkavVehfVMHHTu+TfsBNS73tiuU0RHNY
DOUdFTotQd/nKMCNFwE5JsB+jTb5Cldson/CntQ4572bINFelCLSqxSln9Bh
70CPeIE5AT2PaKMhr0l8HF6fPn1+m2xJK5FavrP+JNCdKPLGojqFQbR2VEPW
fcR+Lzf0MVsWLactQZJ+pu0hKCzC5CmnKALYbkRnZmGEjjXEZc2JNvbuu5t1
RYdRpPTDFnU8Td0hFQcQsOckABxedlsDd1qV+ZPjoSY3pm39hqmrq7jxOc/t
IsrtVQwQYrRMBW/cOWG/MAhbIa9iTFzay1wMzYFs9BOpaaFbagpgGnODWFCz
h/YX534zXsdN/4q6kEplNDg/hfQP42me879828AH+4GYeXbXFrEC9OodCn8w
AdknGSTvZjmakdaJZvm/dwXE1T6Ab/i2a4c4BAGi/Y28xFvIjM6bGG1TAdAh
d0VoXbrRtez2ZqlcMb8Xp/GBFNrdaZKafJUiNxAcON90lvy8VVgQjA6jZCpJ
4hP8ew+/VFKOPeNvocdWHLl6lVPifMKZc69/egRLWlPs0nkBMtCSTy4ixy3s
XlB/dbbGCtLyYLlWAiqwITqyVfVNVf946AxOiFBW8ypDtK1zZF0JQJAYtEDL
coN4ybBDD6SKoY8mEkMVHE+oBxBHFpL0MD0+W2ZU8MzgThRqJxakaS7R+8QR
lm1pudeBSFJKyWYrcxX+Gidy5rkJn9/irxPNrOk/TliFVGL+CejDwGrz7LgT
rvz/dMRxcKJ4OwnZOHSBV7d1iApLq+6uC69QD0BK5JGJk3hyq2aADd6+dtpb
w+FjesTrGje0/JvMWLlBoEA8Xo8saisYuN+0dK3Dy8ACBxvhauvy/ugpMFuV
l58JVe9JVLKhDQD+a7XX1zbNjbEw6PB13zBQJ6REtXpqI/8JcJr6n70La88V
15SKbpf0j6r9wLvIe17fQcrqFkCQG2Qx4MWGeYEx92LeKDypC3EO/KoUY6iZ
tJK5glKPx7vOMJkJE0FRsSiFjbb36HpWq+rnWkR092OSrUaghkCJL6vWdZPB
hsbJV336Apvldgaxq/HhlsPs2GQvQ4Cqldx50KuRYJIy4K5deow6rgOazOjj
CU6XfmQrmUtOfSw+y8Oyxspf4CDhmHDmRfe0HdFbxX3ipzoBgra9x7+DAOjY
WYKd0VZEeppM3YLkHQ9iarzhELW1UyQIz/kcTmBSASFeE2b3Gg7vPX0M35Jx
cFvAjwZ5RFJbvmLmfID5WJwKuwXTdrH0zhXGwkmb6P1ETz4Ncp8ENSAWuTtH
sw5L/yyP6SAEScZGyxM9meBsuFYnSsxY9ySY8ocPDU/13+mJb/RCNzEm+VNV
2lOTReCc5kgEgogaxPYwmry/R+Cd63bLZzlctRf2Ri4Y8BrQdayVj4dkeUus
OI7lMhLkc4ZUoD8dBGOwBx/xdN5mj+vpT8kMHR2HTl0VoK99Qj2GTn8b92X8
cxPxT3BubU0rbE6MqhEUlGsYIklavs3OoKS9qSkAtFfs0SlenS0CeuUu5nBf
F5UmfFEhfx6b9jzeQcGzBIYchdGzAxM8LsQFoenIoU3AFVVUFwddKv7oepmr
WCH53DXCSNgojGHS+NpoTA5CzPwLibmO6k4/aS2H/qfRSC0/UJcYGziU+HaA
2n0pqwcD+TOcjBLv/sDsg+xNjkz8O51ZjHUSPUBp9JHs5RWD9i0E4ZGUgwRn
ai1YUMB+zmrpVsi9CVDnAK/DbOrqAMqljbqsIqRuq7DPnLHt2u1Jt0vJJEqp
qCYU5tRGrY4X4wVOSg9N2IRcVBrzYs8b8dKey43XVG/etfh4q9Az97T227MX
L8dfOQdrXm2iBAWqabfFl79hrvboHGAb8uuojZ7huUQtqmTV/UfnPquxdRij
Ah2UyzgBzQUzKM76EH+Nj8BJb9JG/X67sZh26QCHt/AXVy7z/WSyouRTy4FZ
gel8UNt4Recl7vMxrzLZxR6DNE4nQGiFYCwoMJ3Bn6g1jYE7F+FfdQ1Jaz7s
7RPk01tWGL+2zveMfgfy7k47E4T9PwOBuAmqza0hSZjO3Lc2ri7wyagHDGjq
MR1z2bt1TxM2ei6PKPXoqF0MOBNwL+UldFNaOTsQUvnXpW5qInEgsqNS6k6+
/h1Ud3yMDb3ajZMTpVfQ6qhxu4NDppoI4jAhoHEleIC2/AOJG0I981pqm/eY
PZ/j3DPzbE2gvJ9FefInwT1OrWuc+RXTMVvku+Lr1o27Kkw22P06WE0pccK3
4i+7+1O7FGKKG+r1Ex3y82MN5KIr7uaE3u68PImdp2+iGgg+z5wfyd4Ujw0C
wkOi8iSBZRwBAd+X2FLBdyfYsysGh0wGjk8BDtqzmqIHOA0WyXUelBI56yap
6YPkNKlOpDHAC6IE3CgQXeuQa8Yfp5doObZ9w1y8ccHOxH3VNHo4eIIgvftT
2IEAi/jr3E86J/ysGvl7ho3VJ4GCxB0gToa/SXyP9BdyEJH9r11VyQ2YWemt
ORiDwZcak1zXSWPXGKskuOKlj87ms7EXEmH1duxJsMSnurGDSFUaIGomHxxF
YnDaivPq8m7W6GkMPCnyc6/sdPc3HUuYqdTSTB93gHtlC3ZbU9bxSu9wFU8J
cX57KftwK1OHtQyCJ6goHvyT1LAa1LRKTu2yNOFW+mqrePmqEA0kHQGlGrh6
gG3WV+YcUDIceKb9cIJcSm39CgDyOqiIgVadRIwSsOA5KRdnbVnv2aYFhsWt
8YDNfwEPNA1tAKjHOzMROFvvBkkS4yGEPPQw2IXKtqEX1YLSxRo3Nar+qPWW
mFK43juhTkNr+wxhX8Zuk6G63I3rvtGo1/EhVfmjAP0LLlbpfGipKnJ4uxe8
pfCT4rHxbW6VQycvNLDUrt2YDWGjYJwgSCMOgD/F/2mVLbYQHCdo5m0UVFiu
RrmgKO1t0Xna7UKqqrkMPc7eqJvD8ThWwt+K15cqrN7u59PoN4++2cpWOgRc
Tm1fJPrkOMGtecxZ8RuvzHCw1dNEBmw2VSrq6HTc277DjVdn6aXmMabkcIso
z1DCo3wc2mAnVQMdxp5eXggqOdGkgLfioDBD1xgb5eFOrTsANYeDm5Uv4qBu
NxeQ2IV8WsfLjp8Is5uqrmxVOi5cN6dDQWNfWOcWNHXIxxkCASZ1DonfCBb+
Q4tv6LjLfH8sXWu6DQodLYbs3MqwAEimPRMTdIKuFGhPksh9ZG5lZjzbwzKj
QBKCj5SHFF5eH6Wvju1rtO/ertDgF5kFU45+kHjxVGZ/sm2nm8aYH7Z+Lpay
lLm+N/T0Nq+SVPe1qMZHPkVDCJ9VGHHW4YBRH6rA7sUZWQnrohdiZbJKiSQd
S+G/ZxzUXGs3eqX/Si5Y2ra5gQOikqmwXrfkN13Wdc0DEYRxmIK7RafKrvzi
t2nDeBc+qouAiVr9bRpTzkaTmVVacDi+LUjByS14yUgDfcJToZAbNpK76SBW
cpHIaVrdMLhuIRRnP9UegzO0GDNppzAAUT8T6kp3phJ4B5VrsBcI+2zxcLiG
YsqCPxEAroD3NE3XnGa4jCvQVpOdwZQZlujJZ2Qysd+ciLDx6MmZSpPbkaFE
M5H1kKL5xWVb6mlB9/tjXU52+WozR8n2tk1vQSrDX+hekrTlc2rjZEnGxy9Y
n8Hbidu2Mwh9wycxfP1x3gSWCF18CFs/+tNyp4ZqhImdI8MVdnge7nXLfBrn
1bWR7t6H4BgQOr1UkjCE1AmbA12dB1EyaRmfRgz3XuFyLVGeQcl/aP+iqYne
uXXxX8JGXAw9UE8ihfFv1AYteTsZxv+sZouMYfPhwzrXisde9+N5QCknUibf
KlKjPUy8PF9r7PyZIYoyRebARadqV6Q4dJNkLhNaDuQnIG/LMQGNlZz853mP
7lql6LS5kaO1iFrkiiomrVstSOz9u12C4bywfe9Hw/QjJ1lgnF9rWnHJhDBG
jrbac1YI+lM1QesuqdO/+/xK3DZEgY+/GQdfajL0mz39sRT/eHQjJjnCKG/x
JwUDB0jaBr27KD66X1PcrlfTsMK6Fd0nZxHWQ5L8U4+CK4KS43yj1kJHYHqg
6jeAl8IwFmIq74ZiWBfQqwyVHTwPjj767mBpye9VNr7woK7Sv4gVkwWHrKgD
x0ZtzLkzD5GR2KVAiU+ac9pDk8KzxB83p37qQbjQ551BAi5CNja7100U5ulJ
tH+3W0IZApWF7zqY1I+MHwlAQG+liylJtd5kzqIkPibxSdoq5+8wBJjcALSZ
6YltQ9kQ/9atzZ7ekSd01y0NzaFEBL610IqwcWP0U3ouUjYlTg5SChGLlIE7
FyZCnbcLuWWRP3ANWWfVvKNMy9JXWb4DrlOqk/4KAjYCh0rY55lw4I20GO+W
dx1Ju/oISOWYpqhad1dlvY2cWeFxSbhkkF3x0f0BX7NagZh6UxRr7DgL3yDp
WkozYXslvH2cgdtngemMJfQDpSNXkhxA9fnK48E1I2r5YrcJDQbK2glFz7ub
H2N67Mki91oIZeivW8Hifo5VcJUypOrJGDHTOYFTmXv4A/o6l4x5y2LYty0e
V6mfqkFqkxvsKVrFkU06oXQjtYAucGm9MupSQIwRlACND4pJY07Qjdm8uFCA
lG+t0taV/RAj0gGfdi+iW+UNuhQYHOtqS8ahq/As9kqRS0vVHqZ+g20tptAv
4cDxrQVPKoMoKN9jg19m3xC4ZW5IVm9iEJdhIb1vBGAvw0ud49lxDgoSZS9E
hD+SI7W6J+fQknjaGz79IFXVkhbQJoSuFa3Phze/MCnCf2eliJK8quaBx/Pi
v5lFmtk+D53wOypH2XpLWyx868tZIsBz6u3VvmzDdDokXnu3aw1tSuf3K9gh
bEo7IWCnY08pk4CLtCC6Iof1lVCp8INI5fFeiV4twhA6TqV0MgDnDqiZKzGT
z3TVWYOtXz8imwss1IKSUbqfQ1DfyD7BkeBw+jMDdOUHdbJe84kAuNjEOxZz
XhYeRliToiTFe4/yIEQm/mYl07ckWlY17H4mlGdynRn1SpzcYcw58jLCB6M0
Nf4c6JhjjvlgKswDWaZrNjy29dARTv3FAGM9mrWhf3f6Vm6I3JYyTygb8jzW
Xx/R+5YFK/MBnpoGUhm96aOVLwg448LokTcrbWpP/yKyPpS3O75VlbwH8P0X
rYxHIE3fS+FfrmVCu/CDqQ0jMdPX7RFXjEyQXqlP3KPt1YHzSPD/lxhq2qlM
uwIDFwQKI8Gab74jDUWsqHI4ymDErYsTcKOdRyiiQw5rjIAEcF8qgNINCsJb
1o4c40qFmFQo6wBUiQE6Xs3DEaDfnQb1z0jLZutdUPlUgbgOoCApfaJ3KY5N
qcHtBcW2XDxEZ3GQk8rEQBGSpZuO0MGx2yJs+e3MtHo/CfjXRu99PbT/H9Wt
hkfA6Pxz3dIC+haUrfsozNis0axpDK/uqHxiG6HSBfySbhaW3/1jINjFhBwf
4y9MChD0oTTx27q1Aa9Dy7zBLgF4laiD3fvOvTl1KXiC1xrCz8P/HZ4B+ymX
mET7keJl3xCSMcOMBRVBADSbqolJXvfJS4LBcATLHd/uVgcjmVOvUBSjlddx
pTXcnntjsfvJvmkofPqyeKPOR8JYGY5XQYNhAeWvo9spAb2XeCOCzD0zqI9h
/NN7cVxE9oggAB7/Sdp0Xxf0LokXSPtS04fuEZaAaU2fyGyhFJJQN5ztg0ce
+ofGHbUHD9ROez06sXEqzDh9muhL6dzbPYO4OXRSPta8cjGFcSrJL1tVYw7d
IkzIA5nJmHP4D/2awztF5K3QbYk2JrFLn+74j3ZxSmQKkX3QBuyIP3yc4NV2
ITVfZ5y1Mh8whccRgup6UtOkH4CQF99aLI4U00rgPZa7uPhcjgD0CBjQjnzU
+PNMnHeIDnJxkQaaRDVsKJaqP7LDrABDAGjU7DJgUNW666XGS9TO6guo4mZy
59xUKiWf54HuO1enBpIfE8/vUZVj+Endf+vq6TV4DGGctEuBb0Us6hSZL8iF
Eixv8ITdNPOPEOX0zoSBTZJZoq7ehOc5fXDn0yrNeYldfBqassC1ag33Q4Kw
Z/62wyFWu4ApEMwyB7pt+GDmQtXKM6alBwPHq4EnxYcOjbUG6XHh2dc/IkbI
/UH2dsvT4BkXiUEfEJlNYgnlNkigbYjkNQKvwuatn5xstAfJsVUzeyo1GzQb
VDdarEIWpYC4Y04KM49aCJGambewvfLUeC4dIWX5wmhcLt8wF+1sqlLjBEhm
U1dhB6o4CrQ6VV3ozNNkE/bivBzITbnj3ipc7yvZthUklnWdvhG102HtWY9g
+AANOCmguFOcgGZDfmL8Kf/qxWS8kB5aiZtM895bmI0q9C6fWhQcBSd01xHz
XsseTTIn3V4iDWYeDRn5D1Dsbi9wOCBaF3/hluHd/1aackyzFfE4XWLYPW3v
5XGmTR1nCnq+e7FklUFlQHzkPkNSxGITmij58gzGMo145rVyKYLmg/S2QlVj
iN4qEds9rBhDVou0zIYnGx2kc+iszhzDGTpU/XnG7SlI1MyCIkknPgcU4IFV
Qee+rIJVrY5Qf6LC+MEbk9QO09Lb6uJJNq+UGxPA+WXevY8mtzrLK0ILT0+O
hgxNXK3VLeFW/JnJwqUB2jjVX+kIvVNSEMB9ByTdJcBquQ/ur0FvZts1t7iN
y26PBkKmgBO/c7gkcmt3WgTlOw4vA9NAcW1+dsA7LIeVPerzLo+L9zaFKQa2
/tqMGU7ZQbi6qR/iMiXeeYQokY2xu4rV83sU6+E4wRlXDRXfZJ5TUM4+ECpc
GQbh3VNjOHjlBkFqogSst3jo7FC68L+ttb35u4M1238ToCgGQFMMNmlIc06e
IM9iqy7D+sDEa48dASqe67WlqGMmFAeQPpsi8Qdr4T+jo2a5ckVSxfiE8qlv
+vY4nvZVA2Ss1FfKtphsFi+F+iYG/6gAHDVzULa5IRmmpuOnGyND386OXwog
AI6mlxv/gKyih+1zwxei38HCRlRQjIq5cK4QADYf38q9bok/lbXZQLTR8zvr
Zk2PGJINQ+nacPKntqQoM05iNjrUIT2hIObVDbxG0w4BEv8Fd93cBvII33+5
elNOrSpsxmG2tuoH0oHfkZaTkVznsUwDzq+IECCxtSrAhMsy0dzCqy4NFYsA
KYVINHqfz8unt3G7iS2zojbdSoTNJTfY/uRYDRFEhKN2THSGsZfW6uQHHx41
ihAn8LqXOV4MY+mjhyK22uRX0BVAQl5+fsh+bd1FAauX6/Xbj0gwcpIclIgE
+ZW0WdD8K8JI5DjQYikDm63zhLWhhMYKKdOj/BY3pfUxc4F2Y1ODvAi6x8Ot
fVR/ynCTIdqcWtw3DVlfVESW1jVzhYLgk1iBlPTiscewn144b1be1qaiEYkl
5n4wOwd6nR7+vo3NCnk/rNt5nsbh5fIu5wsf92nrPKNNE40zBTgnk8fwt322
vL2muYKoMaRWS+qJ6+KHEXi9LwJZUyqzNzlJIuyl1Jx7BWLkQ3/o2SoMeHNX
o9VipgcLocCepqZTaJgHCJM8pefwEPBye2KfdOc5aWif3EnVB4/E6CcUbAR5
7WTTOaRm9hC5u+AN7thMQnkLma9rluXvNoTOCZeZk/mUENpnXo13jjzbgILv
bBFlPJ+iTfbjzxiHgM31qUVSTeIJXm0bM9P4RPsk83YzM7mShSsIhuBD4spw
YPjtLQ9Nlkl4t0kUk+JUDORlUARvZgMtiDaJqCW5jSVRFyTfIQP10VBN1J71
IMUViVL0OWXdmxepFxmE0FUDvgGMxwjEb3YA3DSyUGziM35u8Cgl3Sw+wJlv
NndmIFWXLgoPEwXpoZEKuc+OVY9QHEXB7g0iTiglNtc2Bkyi7poetT95knoQ
c+cFnDLkv11ydLOn0jt4Z5A6lzOv8P8nRdNvKXr63ZUHL6OWTSXavGtlnuCq
++jM/JeYqLqKduD/iXEb4UM2057xfRmq7p7zuLRRyzMZfv/lmKg40bGA7GnW
Bnf+nZYEm0JfxD6bgOkaewVx0VMh3DLd5Zf14Bu8gH/ngAWLUveVDg2sxAyY
ap5o/UK9QAOIBDAfgSB0D7jGjbQ8B0nAbZX4rWpbwV7UJO293yQxQiRlUTg6
mk3j3g8iGoGkKYN5KuzdGux4rXOR7+lfUhIda/ByICnp4qOmnvJ1rQwUlT4E
mwCNZbUegWhRPnXVTDfjK8IGgQTaZf1SVq8B3sTalTF8t35eA8D7tPlneq5w
f8CO8zFlZkhSXRSU1XyslBVaJNCgBk5REM6kvzLmu4a08WTR8uL9Ij28FosO
1KN/QMskTVGXuiyo3yJwl2s6BnGYYyZN/x1t74xH8o5dwENDQXcK5x2JAFFj
atN2nzL/BMJ4P1BEiOz5B/nSZK2o2yefZ44x0pLYpbZKLSnTF61pVAS04E4u
GcgbMrqCa1CglsADFws70FwPyqowRTem9ZUi16qKLJReorc7mCNflWEK0HUU
9sVncU9N4zrqD5vbe22fCMvo1eS796Po0dDkDcxcHbeH5+Zm9fmuHr33UmWS
2tWoUS3cGUs1PqWe1+PWYD2OhD/6VkROXNMXHL0hcDqHVLpc1ZxoYnIg4Xcv
oAx//gyYnQ/baqOJwT281mdFf9qHmvSuothmBHuRVXfCZE/0FlvxIPy9DYud
tmaLhj6UXG8s6HAdto/1bPk1UL/BRGae61w3EZWEtMBs4OhTyINwMEsRUL35
vinqgd+6xmnEvcnF4W3kDRfwyu0gBlJ96U3rccrcmva0k+T28grPV518o6Zj
H6ELufDBn3r/v3Kr+Ve+eXZPq6nqDlkYk8CVK8iusNx3GiCPZXXTfNHLQJ2C
KkmWxzTAJdTn5iW0PEbmx5T7jUGmrwel/JA8TrBXl49sjM0EsaJtkuuMkvzj
MtC5nQCHDlQ12KHg1EE/Q6KapRgsyqikr7i4CQe8NU4asjUI2GU4sCs+IEf+
EuNKdcLQU5yNBmSfu9tqnv5h1hXhAfHxJWoEnLBf1FsX/QIxqSVqFGd7eiuA
NGFNt59vDQcJHbB7AYZhS/LUpCY9jo/N/UThEgf2kH+JgRYz7qBxRwAxKvnx
XJfiDMI0r/KpiJmGnRFgXvUUuK1FYhqVCroGsKSTpFqQibSkeDLsF0LLdV0u
bL06wstcGKuRI27C8CONpME6Ag9gJ0Wy56CJu4A+o84joB2o/0SMzMjvaJ+V
XYEDEuyJG9Ync9t5yOQrMEkRwidQIe/TNHPyGV0N1RoBSoiwbiP58PMmwO59
9lQO2gvxHkOQkUrWxz3PFKkkMBw3sSMLEZJRLYcf+2wupDLoZX81jHc6uOjB
6YuL62Lu5BMEachIwz/NJOtF/o3gAhsTZDA4evm4YiWSdtwndFFs4tERLO2y
5i0stVo5dHbpFWd2mpFDRPh5ND8IQo8sks9H+zrplZ1DkcnudGyRGPJdMZaY
KQDsz2eWF0i2b13s5TrK5KS6JEB0z5+w15UxwR8c4nNiY81/8Mxi6NWoMIfy
+7HuQgGChV/L8Kg0KZzoEbcDN6tDzy+rQKT9XDJpMnSbaIUyK8gLJAK/IXuo
da5CtO5yIOjZo7gg0W19zrOE9IXtGi/rfaSOPmY6gQIRZLyv8KOzJIYK/JBS
bp/JxJd4Jc4QWA4J+O02NJfSITsVaF+rNANhIzWI6xTzZNoko6UvM+lfLfHz
tsBv1rlAHUxyyQ52/ot3vEbhT4HfCogH+m8jo5bUJ7wRcMDkBxoyXTXgwT+p
2hLQoi0GxK5xMoVyRlJv63EzzRPSI2BfdROXex5pTBfpr0L/hCqnl9AuMZOx
8EpK0ggFjbIdGPHAOGE8GS5nhzk+qxrB3CDwVMO9MxWUO6SLCtJeXZDZWfvS
e8mR5bEz7tg0KB58d500TM8sN9YhkVgmz46Q017acJv5pwieClr1/9NwKgi+
Mu9dVPA4+IFKydoKR1pIJUmZqGWxArxgLmAHeKpaiCkWguDF6N+HlJre41u+
SxrHbzx4mmFZ9OAbviXCdfWiEW4EFkJq91y5zzWPbmTCCmp1o41ZvhxCICb/
O9B/qc5ldCyI67pPopAUir63ebR3oN85J9jui0bW2LypGELA1PnaA+Ve4bqo
q1EZqomSpDmrsDXVqS/yMQcJq58PnKDLU7aDnHvC0SIKBCgn42JwBFqpfN3N
iYzqMBAI1KXHo/v1tVp416P/fEVzoxu3TDO8pFWvBoSk6lAB0bo7V+K/Y+mI
h3VOB+OuwfzdwMKQ3xlXkryCZOvC5uCrmIJrXsVkbGI43VKvcze017os0u9l
rMB/pYyQ7kaqk38ZQItbONUEZdwqqpHI0/DQlsSwfZ0ClByyxja6mPVh5xf9
F+Lw9rbvRhFoRzWgfljlMhgHHAygphOYEJjG2rEJHwRiSxHeg6IRLnMtQsSl
Ihpe+uGYKlknT54gktyygugAB8qWNtn1bbXtoKdRqiMjZGdcQx9OXc0cGhqd
PrYf1Js1H50ffohQjla69Y3+5AWtzdiSY7syEGZ3oivUxjCGSrK4/JYzFaEW
3+9X4JdeWLhrhGTMYR+lGyGVj2TP1hf4bVwh6/68QIZBvdwQEY23YbKspdLQ
CLfg4bu1U5ZLBgaQnpfnXL6z4abIuyVjfWbxOEDiKHsDgSoArwVuw8LSq+/y
K4NApWBv8auR6nvqTkpWPvpo6HcmbE1K3ObvmLJ2iltNa0gwK97qrWqRbRBf
h3FEkTL/mVP0l5A/oQkmlt8uzDZjxTJG+O5nFgTxnMWFi67OEDjI9OrrxDVv
5EB7exJJtWOCn3MFwfsL5Fo4oet5dGzYJE2WYfKbzfaPMopvUwpVOy3MvwcD
IYzr6AxyCllETNnt4QuwRG4qyg9sXBbyylN163j0MrTAIUutoVvuGI6aY/jd
zoWhtbMrGSrLDoI1f7eyEV2UoWfMlc1s5tVpgW2snHefmiQUCGf02TLPODDH
ii+2CWz6IbuITyVJazPXxQfZVR9mQF/T7Ld3k/qWOz98SzdmvkParZzUkG5Y
anv3h+yxvhCDVQSJNyxx+pgzuUXCbwrMu1GSocZp7qhTGb4SZVHrpqBvaLH5
oVkruXGcVclpDPNt1TCbOB3gzpwWI0dsi7UoziS1bLsbEc4gf8rqsPiOqqCR
P4Rbww9gdin0QCfonVAKatAtAFTPeULWKpJTEii/8atc2NDeNRX1DBU9pkGQ
GF2FJknEP9kW0TxdUV7VKWgjnn1tiLgIyDhXfmz+9moUBa/0nsPY1qp7kl5e
5QlXIoojJecrZO/bex80pXDPKuYbFkeEbZGVKk073cFZVl5K5gPoJywh9vdc
e1AX28BNmK6N4MVbrlPKaj8+v3DpwmqhfFoW2hY7mUM/tNcEQ3HY1OXOQlf4
qZ9XUdGizzK1Cnia8KhZU9txsi5NalVnIFDfA3K+DJURZ6H3OeWi2pJynvbN
hKxpl4O0vaBlTj5v+yxnkitDq8ssQ3q6Z7CwvSHHLReKOq/aoIn0OquFm/yM
3vrqqSkowrV/lo0FM+0jcFg6Wk3bX+BLt3YGybt1uziXD9GQnDV2Mto7//jj
NBm6kf8QXWcGiweI7+EqXbuNocHabfVLhSTFkBYfEiriJOfoDbhk5HiMK7CP
ck2Z/NVRXEN1aHSG3SMMl2KG0PKgoc3835AKExKMPVxL8ycTEcf8b0uKaOTU
pCE+0PlSlKzBXxXJzEtu7TTrcOxBm9XfVQmZdsa+qZOMoynICQskN1hCFniE
icjeVEvpW4ni24iQhBzN5S/jNx3dBwaNMBzfUB1nx3HZZloeWWAcRT8HvQ0H
AALgpB//kR87616DJ9/ww82Rx6ktDYbXHCkTOIGyh4cVVcJGv0hoYVSDdF3g
x0hpPX3PvvkxEG3cIwL0SrC0jSCD3lmk264ejYeRrver8Dj1d7V2zdfA65qF
ZSX1klIYwSPOlx6z8s9kxjDgx50U8IbpgaQGFxpjPJpLUbbLwWFgW5N4bWZy
i+ot0hq5Ohm0ap7HU6jVxnQXlLEWLL+ke4mqjUcTujOO/DXfVkEC6k7Z6eVi
hp/9zXv9M3tVQdS7V0JZlsSRR+Aunpi008DYB+1sb0SdmMFDjZ4fMIngzgln
oamwprMGiBxDLDrkQ8S8QX1bwJlAFYXn7eNb6M2ABOJv4qt/4mdsxFlIGzJ5
iR4Hg6DXwDcSubhi7Hvebw0hc0QofMtaV9MY9oU4dO3aal+luDfjwzqFwT4A
KH4PRncd3jghe17551ojcHcYE8g+17t1O4lALpqJo83FHXwphhdRdczqE2qK
PQq4bqZ5aoa2NdHl/+fR1rynRFYLjrjab08g1CfIxBIf1zMlOdhPyL2gzBYt
cfTTRF4fbugWmTnkyQ0EvlhR1E3MhIja2yKXXSn5NnaKVNHcQ317T6JskNZo
xtQr90HW68QsJ3KUODkN3nyY7WWmXplEBgIo4D30KOceiaOcelzU0UPmghxC
9jj/FEiJokN23qQ5P/sj+oIMLPnVNu0Jrr54yBAB8Wd2CWeMNmqCHeVXdQMr
9fLScLj1tCWbOIWypykHb6B9qIrfj9cJ/HQgUXwKe1LoHwtwYDJdFYXNDQI7
NxqHrBNnVfW7MEvvOKP525Dm3hEYEE9PN0iAPcDCU7oN4y9M8IkyYJmc8uYw
EZlbvgyWxYamoTK4src88Z1GxoYoN3lnHtW1HUsb9g2xNvnrw/+3t2X/pvef
ZFY6cX76rum1g7lUJwBmlQxeAqd22wRIJvVhKCGqnNM6vNF+9+EL9iaw+iCi
S07ISFpwIFRL18hnacOyzgpolbqU5sJ17TZBFeK8MLv7Du433VPFp/rukID7
9PfJR5hYOcWr5b9CPw3DhnDVQCbOrF1Urhwpmnve9HgEWABps4Fa6aRdOCFI
IN9o/iKvKbaToxdMqQGOqIZxUbNRK2ss8L4CG8MNRYMBjEiMPg/XHZd2ec6U
K1ejJOGzBgSPdgpq8aRvhdM4tvd6PS4RJ5FeFMDKmZ1xLM+7uaMqoLoMByST
q4cavzwZ9CSvan22rUpJyQN3V81D2p1t2PVg7IujYwNZw/wTeP0dqGMlKydO
jviEiyCcng6h4o55R7KiDaDMJr6LWd4IEyp164MVobMjEMP4K5nuuwMfanX+
im9zkNw4pXaZwew0GXfjjNxEEwOBiF67AYC+WRaBZ6zmsFLWFMUUprEEuC+b
2dCyU8h9IVbX9j+Xkl/Lby2SfNsCgIhdlP6g0Lnkm57ANyZ+Ay/GI4UTlWsx
3JkZda+lf9HynnZ/kA4GuT+Y0fWpj+rshOChl4zSTVPszKFTrjckeVSVJGpy
9akxykLoXUOdGVZAAjygVpyQpI3xykL8W2VMRzLUAKZlltrqzEspJXUE5kUM
lrxDhuYoEEFLO1fU39MVeUn81Ct/H8AvHo4jLvTIdAFJwVXd6ZIQ4uOI8Qjs
IraQnVcoe9e+A9oIurvkNIqW8XMdqzlX/YZ/vJARhjvOcuJM64jzPqzJLYaA
EPl+DzMr7xGoaxdbHPFnUUOlIjJ47pa51JlQRfLHQ8jsPMmafNCCO6P1NHVE
cKe/AOhp6zwvbSWSU26t4Vc/EUA4zSfnJryd/Zyy9F1+UbW6aIsW5HhB5BD+
ynH6ng94a+sM2DyhOeH5dKz+pE9nBqLewcoc74neO8ngdHwIFiDQbF3Qy4aB
lsHHCyw/vxwlgx6ZgVr8z9cw//QV4WM17l8vTLSwKaufKeiMpZpQbfYwwa/Q
sM6BDVy8qRHUz2kFheHzHo55mylG5kNCKiExvF9iG07+h6z7ihkVBXcxxjNl
kKt0UUTTLDYhQhFJfsrQgZg3k38iTPZX6ZRPKsMC0i68r54vRo7gAG79Z1m0
K1FE7q5XzZLx1qOUsZBya93TgUyQ6aQdCjqAVEljGOSLf8K9quAsibeIH5zL
fDO8yGMNM0XCO7QqVOfEhr5i7Oj/FDnHqOPbOyeAq8nz2YWrubpYgAy2XVcx
IEd9rlXPWlRnMvbjhvfABfrLqJb2EbMjSroNu0r+vyW/WqNgi/wVbRxgn4ut
PIb9gM75vbFqhNVf3tNAEQvE9mLgolAw/ezMsE50EDvF841k2KB2LNtSDcwv
lj38nF0cCyLPYvrrJNqK1h4ag9ue5NqBNH1Ydi7Zvo3IPrw6q+sHtyKFwcGV
0eXN/5lpyAz8jsMeVCoGrybluJYnQpGpENwRBsUKiAS97tAT+NGcWPKEe1ZC
JrJkMlYRYcG7KbXEpO9T7Amqx7dG3crfU5LsIZUN+pQZwT8wMA9LanYgaigD
7glgfurbwK3LK0I94nheyzLWMjf7g/umi/djkPXkLWpRzjQhHV1V4PwhvfpR
dwEX0+0dL/fzhE9BIEBJ9D6rbRVI7N4zWavc/l436+CBaOt3QOfFB2LZ1IXP
YJlmaUj1t61d8S/RuIriKYvuKR6kXo66/2TVzc0cUkaBBeEaALfYGk/1+7hG
JnC2uSovMJK2BG+If7dbM87Woq21PMeMIxzfwgQSlID4kciHJa46acAnWboZ
XxprDWqeOYu2VLgjfrZHoUXg4R+4kMfWi5DXNfKEgNOnO0YhaOybPbFML0kw
mSNhUosQkZer3WStC4qZJNWs7FSjb0GyqDs8QLeZoO3DtIMnj6hYak0pV0Ur
U2Brwdz2h2773bPd

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1LLfdbr5brUILWcJtPP2/OEXLnB/J5HIIKN4pEBU13wEK4YJyB19gDz6CUrf3naXGeSmawvPmX+SDB3SwF90y4ch4FzfYaIrYsTaOvN4nQTzjhf2bxTNrE04LAN7BlKtmo24LgPtByhSOVKRdRUnC6vBK9SrZ1h9lBImRypoxnf1qoi3bZcO15xFKOqX76ZxxZDyNOggzIAzrsB8gLwXvAVidZdOOwbHbJxTnhn5mTZjVLRUw0/VlrS4RW1l+3TOFSMeEN6tSxI1HOHuFTdnBHAn4eJ4ZPYuxjeVK/NBj6ZnPF4ztXSqKq0tnPsU56pzbGWNeiv4hZInEw7z9lvBTh4dQsRQP8dZqQf6sCkQLcgR46pqwiKJdknonX3aiHu49o/g0d/vkYzcIlUqfnFvfruo0QZWty4dZ8JYhT7a93UZpIGEjC+VBmNXgnblCSxTJ3lEeqjKP6k8zusJXsG8txx/BlswK3Rw51rWOrer8c5oAMUxG0ceSlu7vl5695uCKfQIfEh34hEHx92V1+hAMDwY08skQrsUEfBcl/7WOLQENPfEXCBpo4ijtBhShzK10Uyp6wz3BgS2AyzmSuGdeXkd36k3ivGSqeg91M7r0O5U1pE1dtdOnU5XzokBmUjOYbi1WVFLTkYgqqWbPgBMORAvX1HAXq1l6XZ3BTMpsYdK7DFGhwPfHhzgA4XNvxbmAbMuFqsJW1xsP02CP+itaiw3BRDKSYSUIeoroQBXmx9hmdHCedJrMy2TimBUpB/GQTtyIOUaq/QXGUOxOkXUm1B"
`endif