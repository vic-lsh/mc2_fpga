// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Xbg64d9irMdQ3kghtD1ALq1JOqnsq4Jivl1ix0nnMTWLpTcaXA2CuZdYsk8A
UJk6W/otBUQga1n5fWgxf4j7ibaFbdkXhd7MjQYyI3nKyk4nhf1QNGHU3RaW
q/q9BWO0lZrPx+c/muNZMYgc+n2Qxkml9cHTsfPFC5AbyOMoVG2b/G366XxH
JCSe+y1/BI3oDH/rRyM0iMa33DCd1CNWE7eUYhOvivx7YaDmbfv5tXUbbwTm
WKnp9n2F7nIdWdbjk2UegNe/IOPhbqo8qBLzkDpIjtASXH6XL1/R5menemo/
RnbCGnED6sMspoAIez+jJYKB7GGa9iDXuHST7Qview==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PpHHSuVRrbaKvXBMSwWzSSMyzSf5OcCoV1+XpAcwvu/F24jnYR+GDrvLAmMN
/A+DuY5f63NIZnRF4Jsshv0SjFrM2jTE21x+15vOwSg9boFdcL3pghadcRcT
k4p+12st4M+5gyiA7bsQQIvbN6akvVw+Cx2gYENmgQS6xggjlMpBaN3j4Ol0
rxW7bemPtxbrAG70nQNpyxStHSQLrEbMvFkDvfe23ghFxuOfEJv+THLi8J4k
VH5rjOMgqnn6+F4WpPII2suk/ZNfuchm9yyQJbSTWtT/cpkoI9dWFtizVIFf
sLS7LqHS3xOJM1iX7CJDHdl7Y6b1s/8keOCIehUEFg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Dj8AD2RlDqezMMIUFvb2OqZ58DKX1r18lAQqZkKLYiiV7S70+pzhp0OOMz9Z
8eBSyxL0BpcYVNDE1G1VSiIOuuhZL6SwD/HzajbgVAG5ZitmmoFPLPn2BvqO
zWj9gzzsLi4V4fgNkbnmtRXTOnsVBKCo4i8bHbQaqIm9gp6ap6TeOxWK6qW3
lbJn7db9JEdnmsEJa5D78BcNOkq/akGsbSf5r4a42eFp89eJgpYGzMqduCSK
GsUWBIesEXLpekiaielKrWrcA1DgUGQzDW3+AiUe4MejRNVHmbq3EXdEEcXY
IDDYzxxK5byBKCp5YfQ+fmE8uNNxGvnSZ7/xZp2XIA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qAzMYhBAz3HGhY8OXbVRYaSgWRsc+JFrxD9XdcodDh+iyJcHqoEz0wo826FM
M7nxMXdJ4S5+/Z2ltayNLyBqwUC8B8XJoy9yOIp4PlVO63HCEb0P4xbMtlou
D5zfwHD0+Exs2j23hBtmaHHSv/n+OonKcVKd3zKyvihCZKm+RwDyQ4pZSHYE
JE+rmiKP0a8zEqdbwGJCftwcJFoQ7BSryBkiA3K/fQxVGoKHxl4rjtrxElh1
S6QiNRJjzDxlh021Q1rfY1TSq4KKKOp8Gh98EBRcIM0zwGp0b9IS2RPc8pNE
NApzIfkGqgeakOFM/VjTbAPlIck9qWJ4tzpZq/7vWA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fg3kN3I7X+zv2/3O8clc0g74ioIbWZ92mBFxtHhCrfdd1TEmlCl9b7HwGLaY
PkSwOTyouhCAIa7AbVFXreaTtnm6P7kPxxZ41O/0nO/2v4xPy3IWSBkF3+66
BMWUV0fynTcTskoLNPrKy4ACTifSON7wSxs9ngrOFtsfVep4WrQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
tHohi9mfsWR7XNm/5jGIVKAnA02M0+Gok+o4Mc0xSfBP7BKA5ThBWvRasu9l
RYuD38SKV5N0eYGoh69t2XwamZmx8Bs3xrjFmH/F5y0ICBl6CR5LHpEm+O6N
XCmZOg6ubpfKy/TmKSJbirGO05qKJUaYo5ckxkbYNc7npPLlKONwkYOoIyQc
Pq6di9ie6tRP6RnswSWMIRfiwRC/WPj7cDj7U6IdErxidc/6b8hNwgWAaTWL
YjjWC3IWUA5fjeEGTgrQZ++8IckBk7P6oxU1aN79DOW4OvdydIBU0Ciq+b2B
mNpAEQBf8ceP4zWAnZ6fvaI0FzrVSxI9REJXJKEn59yCjxSTuZ5zpW9XL7jN
EJ1/gkhSEGRPuHSEbYeDxKJuUj8Ga7QSad2YmwZdM6dWIY/wlfmOEY7KHzfJ
53qd4HqJ7IT6R7uzc1KrTxZJvmTPebyLwMmKNyaTJnBe69ipvFe8tBNvWn88
b4Tme2DyZqbFYmPaECQZI/CDSHm+5Zv6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZnuXjxGZrpKmBYMNfKq4RN57xR9zOXMoeZxATevExH1DikmqACmcfLYfZu8Q
4Zq70up21DK1LCM5o+iYcltHiewUAVZ6tbQKpDBuZyKcpky6Dl9tmkfNMRut
hIqM7pvh6885ds7Jsx/d2u1yCvNTxFudaEvHiXYg+wLyWq0wf6E=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ulkV7l/3Mu709KCwA2NG5+hD9DSE08cpCmee2awDZR5/xtWrBtf43ZAstYkQ
KwBU5KK7/C9Oy38gsyLJCra1od/yqWba0nkv1j5AKItKJ+PCgF6tR2sJlgVH
gclXw0Bog1x2PAnRf8ljtSRXq3RbDt7QPmtIgpTAxhGDcwERWsk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9680)
`pragma protect data_block
Hu0E0B1OCq6nIFq1KOjgyVagA6K0HX0mhAneo8OhlDT+a8PJjKQIG7LOn5Ta
wFybc17ck6K/OYhvba+R9B+PcUK58x29h1S2nbZkSPIEYjVdPLqGGuFCyMWO
gXgKIKpgQAg+cO0BsQElnqVkBH/2XDNhr/osxYXC6fAhfYXP5jB/ocTTh4xY
POAOUn3Hd3pRrXCusrsPCxh11CF3LcwAIVQhvmQrn9CNCMUDA7LYMvf8hsX3
eNU+5zPCcn7V3bM4Y9ZvR2LrnBQd/xXu5pq9MHbz0oYq00L0OM7WGITY3Apz
1nHYgd5rbQ+fNxEtJW/8sssJ8IWTgeTMRWigACUoJB1Jq866eESlYrFyea0R
Tl9nWgSykqAAS/jv3aVpLfR2rzTWICpjTNYPTPed3iJvD/EOw4/4tmWTUhdu
TB+vC/uBtXUKoevolQ/EVCB4F4P1S5sne0iDWND6IUjUSWy2zDMsKn68UlXC
1cdXpSPuZt+7wn1dpQ+O4n16944hpYxK82HDfuY7RdU+m+H3U3HJjs2RMDcf
Qwzs7CII4lFFmaGAP99epuBbFoQtU+avK1Uu1S597Y2bTpAuh+7Qke6UD7rN
IQThL4u3pnfeZuHdL3vd3HvH9vxM3OHBbukNZ3ebbHaSCqtD5hvBK1yOF84W
bHbtYUr8lS7qAYNNUcpXc4BEhNpO4HnHV16SXUF7/NUJ2qaN69GicUsj8A7e
XfS0AHCYnB0kIPNXNGZfu8VqM0oO5k2tjRayyGvkGliUBpbKIocrnYnpSInH
einvMjSByn6j/UYYlfp82WrhDanxxPUekn0o6HDREt/m+lAq4Kf9eBIHm2cx
KfrlbNtyNhEbyYGQrDSvDiWi+XDlRtFKxRJeFCZ98D03j+QiSacQahHhlAsI
TbJyR2ykKDGFbyYBXwhLmQP6U/DVTdaiN8V9XD4dTso+GhBEJI+LHkg807VN
hsKsfHrlp47345S8+IENYX6ZEPAMQGhy+fntFHU9TDR/HxRi4u/prwrh0vdJ
/RH08C3ODWyNq3YZ4IW6Oo4xihrsbMqsTlj24yDhIKJ/DqC5XQxGycshXlHz
FdQz9OGnHAM90bxKpmnseMB7v3e042C0ZtYuv4ROyeSXn/f2/1T2OTLwJiHb
ahfc5NzPSXdT6FPgm0oR6yrUvU5Xw3CQbE8LvIZkCyDpZZKjNanSY/A4pZJW
tlXtdtnIqhA3WvqHo4uJbptDrm58S4nvf301KhCJONI0U0iUEhaQGq1TX8/E
fga2Pam8jiG4Z2DC6TvOZWxVHZRlZP4HoPjT5Lq2xzZsaoJbVbTCUcs3keHe
nbmQqYAJhcnTVUKSC63Isu0762zMsFy37ZIyAb+zbCIkwCKQucpWJC+KSF10
NFbLSooLCV+ShPB16Nf7QBNbu+yGu2MG301kSMMp+Fz/SqmL2OzyGgzMvNoQ
slt3GUvFdlVgLVs+m/InHg6olRFe5vI4o1x6Mg9FiQouxzJtRissAy1kFCJD
MCjNEG1wUaVdKJexom4GCpTJMbx4+7V7geLG6VeREWtL0UhDaVVbvybkTMSj
lvkFATDMm9rsGSeqcWV0iEtrp1ITNJlRxaJF2+LsTYWgNF4pJgdpUyvdZU9G
3tuIIVkSWdm8K4DHy0hMx5cS1i/Uq1q99icSNn7VFVUKLTBJwTLtrzwYnMxz
OV6nEYUbUE2F0Awovp7ZmewmQGd+VueaHbcDtejIrU477Ddofj7QUeP44NDX
Hf8nVRlUc3Zb9K66SqRy3h9YwPPwTJl9+AC2++jPyIB3vteXhGpPBpd06XYj
j/1gwQmg20oH02qPhP0mUeMn0iLNwoj/k4DboQCL46LFNu5TRABOwYuSXBQZ
2Ea+SXNuHj0Qwcf9BZTIangLdCXhsZ7hdPSkDtel03hH/ayQANy7mmHOH66E
8AOgvp75iv7SXIOS+7NhDKR16M4/OfU6wLijEmnxKR/5KrCudYm/9qMsjdtR
m7GWZgh32bZru3C84PUIR7dsCZBufvxHpizkEASjxvAS0PsHAuGSLieJx/LP
bjNEPuH9nrccMtrY+fy+qCRmzBz9o6iuCyoZg6pw16TvcKfJG+0UF+MhGqrT
lp3IkIo6SmGEeOgUCUMNZpwgQsQVbG8MlfyyyPLumTCNXbJL+yedhCYR3rox
2q0ypt8/ubQfVZOSrxKqVkHzGipF33ecuITTktz3F5eoTilmOyWH1yHyzNqU
KNF8vF21oVDnyJ8Yes7WDFnzdPZlrjLxQ9nT72bnqSc2mooOA8wvSXqk6Uvc
jdlamYnbmAzO+rif6hEyVf3zsMcNzKGSPScNcQyoLA/HPmeIAzzhBt6iM1Yg
2dIFhgGMQpNb5rWUhwgXz3EnUsTcrqFp++USlxPcwCq7P9ndXFnz+HKYMEzr
dQEZW2ikNnLSZYHxGkgj0n39vPuKKT3/Tm4meNvQWwTUDn9wL3A8vsEIlHxd
MQqpq4mvKm6VYMZZbk5OO3BQgRDm59JQQHMPD4/LZJvDzlCicKcGsBsk6trV
a495PI3dU6LnsxvaOefMDyTe87Wqi+dVpCKtb27iSB/5yqMGPJFPmSQsrDrC
QahshqoIoQ3E/cKIoRfekeMjIN3ej9kmqKdRYf9VkVqIYG0/1Zn2MZoBHxPF
Eb8ayyKBDRL4qz1CIT/xl5EYVlfLU2u6dYodpyx1BuxJEaXNWW59/UtzDOyW
U1kwQObO45heih/Y1orIDRTlQtur1zssfbI79kaBOntwVjeGQljYlE/Rrwwq
XKVzOplUQN7bkOf7mi5d+zKCRae6JNDakBynQpBb8l2itGYt6z6qDiyM7IAb
8xNDSpvHVCEhtMLEahk8VWAcKc3guN+oiqNwDlpD+U1mv10f8UgHN+XrD6Zq
AqYjXT5A6dpPLJGLclM3cr/AweNC2pSE9evMq+JVYgf7rJHHIR5qF02CJfad
R6w25VAeePO/Wmwi1nnMnM0FEKwIhGMvkbxR4ms3Vw0CmtZPlvGobd6RlX3U
NIvNTHGCWUlAq6n2B66mlnXjILV5DTclyVNUrBeK1roSvS1ZZ9YINqVp42WX
yrsMqtEROza2gLy4N7pK3dOD5R0K1O8ramXxbC/Nn8ti35fA1MbVSdpPgmq0
xSfZ2uol2vVxQR1410SnshC2AIJd2NMJJurT9ug8RtYuuNjSy1UfaAS7SS1v
FughtBugcT3hMO4He5glcrOVyNXMruM33fBW5FIY8RqMmtvAKlUgd+yasMLi
wE6/wfcS116zcsB3cnWj8hWiwyzJ+wOSTEqHcxzUBM66S1QgD8zj+RckBIyx
f7E111/vRzxt7M4iD7Rg7R9P1YUo6K6UlhP60+UXZvTe5mKTlJdz7Q789O9C
BfixekaUXcYW1dUvio1uzUTyj/j2JI5fE3wUhA3wmvKEfG2JT+NSoMVLY4tW
7+u+Td3t9OmfJ7fXN/MQXQb/dP098KvXKn4uYt+zJybqO9f7KB+6hQOr+fpq
ic8dY0v812U/gxMJgWjhpsz30YyaAXxD2/7FW7dVJsCtTVGHeO71tJZlP2ID
ca+mJV+s+GAgxwd1Ct6GS40PVbEWLxYcTlkVZIHSMk4T8Z7fsV8dCnmylxD7
n0kRJoRBZaOhka1JRcYu8eStvm8IYUAPbg9xaEhz9+b18kvNFnqnU/o4xVtd
xpDqZrioh5NJmn+DA7Lt+63vCeEaoFUj7nsOM+YqGNaWx8/K9zR2KgHOaKMh
KAz3gebIjsFnvqzMd2xIfrBcq+wJdqwaK0ORD9KJHqvQxvgJVXTsQHaOlcR8
s7v0FnYfcmTA5dm22w+vCOQLRbsITaeDVXv66I5pg3oPW5tklPNrlJ0PA2/y
NiqbPevdMDm/zeI6s8Im9etxCivdwHLMZEjECJLmxE9z7fzar8qtTdMgQ2BO
zBdjAVS1aHxqrFbyhCieE8kP0JxxWP8RsG/dvvjWApoIjbXNRUMMdG4vWO1w
fJMd0+rwMM9P6IxT4Ip9GPbc4jifQzeTnhYD9RUP71azsNPU8q0/WcuE2oio
mUfEYVM3yoC9kKzFpp2pNK1RvTdiW0ICmViIILPuS1LOnCr28Yexj78r5pjp
IIbPK38SsKHS2gf6xnkVbiguOpa3j6EB5dUMN++cWKNjpS7tgnntCy0Aow3R
5JIJYWfNgT6TaVHD9ZMosprgzgRwQOVwPH6wyi8tGlBBeGJU1xKEA2dPY18l
nZTiR6gvQM1DrkZc8vANRynJ3S5wNSK+QTWoIUMVDdiUecpctjdYEUPmwvJx
T2AHa9OL6pvczjHeXn5c+E0+fA5ppkpRXE8T6jiVtw/U46Pf61os9Fe84EWo
ObQhnBeJBcmjARybYhJ3cRLFhNejHfZAuJZQJPGdp+IHDeNpKEz/LVofg1Aq
489oLdVB7kP/eUK5NVX56QDkGiDG8CvmggePlCBsLi/o10S5AfpA+q3+kMBp
3SulnpPGZ3fvG+7OO6I/sygCR4h65ivWqJKklCsY0pujw9m5swlBWWFp82hr
OMGwQKf1gsUI07kX1xHKrF8dX9ET67yepvQ7sBe5hEfHS5R3ZKWCLuScu2gC
t+HdzKj4hPl4zcQTAE05rETlX9e6bp5RZfQ//duyGC41jusRytBhRASWsDZM
ZtYoy/jSQrR8Fa1GovwkPGmNSU5uQlCHz51UhEe5FSvP8xeMwwZvI5Glx0vw
g7zK4pT8A8YcMPQ+uw6H56k5rwYjhulrHyxKhMn1Hl3tcjNBch/3tpgNZ+1A
cwfG5AZboY5dAqy37NgVP3EUfeetEphGYkgGadC5+UVI5rvlMNVzdRmhSh9r
AXQhaWWWsThXmh+RRyfIoadIGW+Bu6SHtVXRDCAF6wCH64m3ut/8FgyjbSbM
2hfeVsg02TE3UelZHpFYQ+lOLuY9TZZkQ6p62acmzIq4dFTnhe79POV/ZxoX
rsVhb7qw0QgAx6HPjHoJfFPIvb8gHrY4tb5lM2i9pJKfdU7cWfcJ1k95Lg8e
Ie2ZIrQU/cLA92TnBa8XaKtw21KC3qo9qSAsXLTievi1fQN1DQ9/CTeo+ZFL
IGN5sQnEJb24f54VaMPjW9VUnsusg2P2Ul8w4dpiAA9Wx7po1KXYEBYZcpb8
/p7PN4r/w5oyghw0UYozGhLEqbwUZNHin1JnYK6jL51wJPqh5nG+GZOFdBTo
AxpPHxs370NaKk+QUtbj8tfeE0DNlkmatSwXW5FnL4j+aEg3JodjgB2owXwG
KN+/on+L2cXZslAZY20RRSuRiFuiCAr0/tyPgyiQFIX6OQeJJ6ecZrGqg9H2
d9pUY5rkaqjCMHVtsK4ydUQ33bLYBxDWOpMiInr5S1a69dMe+RIUU31ihZxU
Mxvny7yMVhD9Bhg/hCRyCzmR7hDNwN1HWhb0t3tO/knPimX/xB0FnEj2zX5V
Y8CQT94xbBL7KA4Urut/M9A1oJ3WTMBtG9KL+1c7hcNOe4AwfpEzDvPsHFNp
Jj2UfJ8hYkEXXAi4BodeGUS43ZFr60RzcL+3T3XodKh+CTbuz8BZNdhbkb0h
eWZraCMfKffKBBkEpG8wr33srZep/689ePH+Z39Xbk609LORIpj8IzX7kG4/
WuDdw44gyk4u9i3XFDpP2XYl1Io4VBDofet7PL5++FUhdccK2YcNh2OAnyQn
/QMIPREJgrx9b4djT23QCTvQnUF/dPGRujJw4//97iUGSZ7i6U4gZmSCfbQz
T6a0Mg4DtZkwfdy00dTVum6gF8oN8EpVaedepruNP5DfxfzRWy0U3GncsSUg
jdsIcTauC9mUNbISqvqKZ2MrDd+OcRmTKhC2YJSD3AOnqHU+/g3Xjs5jImBK
LD2WtUK/fs4ymptCES8HFAXiZ0dKFsRl0okErf7aiGQklC5tTTQFNlATdtFF
nnIqC7bIRjqlRwyIlkB8+70KtRjcHXuJl/wfYhDUyO3Q87Rnm7driTyUDHmF
32t7FalDN98JFqJjpmV+f6AsoD/TOyQ8IE5MFJVBc90e5gmUmlDiO5OUtaxn
56xpkhaxCZePZ6LfZfpwZOboFL4V6h4y0MbQyLdCmZ2TaHcL+i0byfcPnv1n
1Pyqkpe0Pn2zRLr262/54yZXArXO0ZIQOHGOjTAT5ukYhy02rVaZrKHcZ8td
/uoRMcG4WZluyRWPQz+Klt2GHOk/7+JIKpovyIv4ngDqhB3CCCnnqlwVweGI
JCPIQP/HKh1bLT338er6C0Bj/zCMGyre7kslsRp1VPIl6R5OWlmn5z9KNiVF
RbfiMyJBU3CGYW50qIPX9OPhbjvCYbFdb84dxXly25z4lyQHjyC1+lAB+ghp
shouOZXj1U76XQd0Ic2rVsYREEHyaeNn7IfJaAzhT+KbDL99MB9cYBkk2+vH
LLvk+8jvLVsX+LyDnvvWjz5VIJRu6DGNN6Iok66kDiaO2KQMz76CHGztULQe
G/VNnCTnZJx41OK19xGqY1g49Jvzngd30WdwT4MxEmN0H6tnwHUgGzJkcWBb
DfLrNBrdyapbxMvstaHz3xPVc49vlWn5cVznAO7S/N4d1kbtuXIYHBm9pKrp
5EJXdL8nlMijvuAfLZHu5OF7Tjwnkns93i6OYNOtIJqm4Ae3KPgJ1X7pNmLb
pEYD5GZD+2NCdd/taGhUeFlzr4eF3fJEr5GcGcgLNYHYG1hBUWFcc3PfkSv+
FQoYvGjaTnzK251WNBKlIM21pmXD4FNSofys/KsnaPn1qP8FTrSSWcVK6vBJ
sYtZkeyTEZ689Qmg0twuFjg+7m84q4e+GuXcpdG2ak0INVk70e6AYhxwKqRA
cQcTgVCpuWrP4gBRE+JB/jmMLSjxb6O3Ckaf9ztacV+NH+ExTIbvHGxEgRhT
M0ClnHE2FjXlOUrHs84CrCywE0Td3oOWjSqPkfgqH48IiaRx/3PRqxmlEXrE
yezqnMgcPKm3Du8hllh3LjQwJNd3RMW3w7dE9NtLAPfazhBZFhNm9ua3mCpU
QXGSUMx4BEARrdN8qMc8ZQpDsgRVrksRvEIxgmyQkhSAS80Xn5cakwByu3Ug
oCcvZBkD7gwobvuzp2ApmL4MbeWzxqqFTMImvpYx4VvfAXq9zil5f56I3G9L
z/uYEDq8o9ODQR63Bwv5kTc1JxWiTXGi7aIaNjHE/CPv1k1N/7ahCQlOQc+D
puojqxa66/tALD/ARbKlSuv7SucESZHZmSFcFUk2ScWVeoLT0om7DaQdp/E8
MH11LR55jksm63Ax9j4AoLIAp2387eNv+WzY0JeCuLkqfU53755jbcitLYHz
cGghFtpIce8NQZLRI4BXVbaZbIWCn25wbuMpm5Ts+XqECkw0YKGKH+uWGz9v
k/XsSd5rEUMQiwzsh/Dyi4s8TH22lF2KJTI4pVUVjeGL1e7uzUgZNHiYpkyd
TvtYHiRi3oCVoJuvC3XDzy/0aGDQeWGQXoe1vWa4h3TLedbpZ0tRPGLPuZuH
FsemwFhhqvsRg4c75f1INZjCEook4iVdjKGwiH2H20d1Kjq74wD/gxRqZW4U
RFr8qt2+gXFnSzyzarQ72t1PFnYoEgPjaLSkkh6Q2WakskSMlaR6jf7bvZ0h
zmzEOeeVdCLulmNDAGyTgOFsQN0aU/ga7q0rL6fgX2q0vc1mIJ/A+GfMMW/Y
5nP0cwdeYEP/uK30Qa2RnGo0ISnza0wMrFaIYSWqv3h6biHScXDMelho66hO
hYLHmQMgmjHradVGOODhhMvmYF/UjiD4h/xjuj41C1LUrOBI6z+UTpxyLdwP
pu80OIj4Q+/A1KMVDljSgsIfPZZUbjVIHdMwKM9D21UIegPrqq9KM/YMEqF5
zeuJ3cq73r+aksD+hLxrMrQZoQLxWZ+s6YCQI77czR2740w+wAXrNIhM30Vr
Sg04Dy8z8bQT54ciHp3wLxOqTEIvkXrc3EM9RiR7Zu7SPzskxWXo9oNgjDdP
iKMPQva54muyEOUtgHWjby9obmQG5ynlYnJlGaot2pU0rdq07WnuCquFN138
TWxtwQelnwJJtmlNehJONC74Nk4pCzG6GaWQ6U9ZDB2czaA+lhw2n4+m7OyS
/ynZagJMKFzBpzbaIfJbMj0rHx7xRmAJEXf5HDNZjAXVwXGbFx7IpoVG/UCP
QJ2NJAcN7lXthwbKH4fg3EXnpzlTq7eqEd0ycHujXE9qEoP9RP/QRZ35BpRM
4OViG5W3IRbu+K8sNASzHXSw3RS9h1CnILtQO6r4yWvBDIYcaYMyOgHWQOC/
P1TXLvFf9stlRnhV/Umzg4N6bshhU7KUMKJwKb8Atj+p/g4VeSsJgSz1mjyH
eUFuWv2Rgb94ypvoe1z1y0TQgi1F7N5SBuz6Xi32XPCMmg3H+P0dq5Yp8F/O
A5XxeYIW/WAfdFiQEqUvcQOrnNvWfiLb1oa9RVQfoFMHmNP+trxQBPZ0h4hf
5sNwIl4qldlNP4LFl7fhKKR/kePiOnS+L42kjYhN2vyCE1dpODzHMFyz7C8F
2DCM1DQHrE2yyVU+cM67QdXW+dxnDbz39G2dItx7R82eYbW4y9vn8p7kIniC
hTXWAclfte8+eouEQzrvPVN+taMDq9m+tYkE0lHaI9vY3x5DIMNIN+Xf1rLv
Gn0DQydWTGN5sQZ8Fab2i7K3JTsKW++n4vQ0dcQtTxbFNZIzo+RTdAejKQni
ygCGjpvmEf+/ZVjA1A1XUpkEn3oCi7B+41izW+lzMzBfIgT2wcIljBOTgfzL
Um8qExnxPDIQhyhvKkQzsBUGaUq4kCe/8LJvjwFBrs488EaoSl1vsUiOoqCH
MePqKVnSNV55kEPuYleMQ7H7E3EW/i/x2EKpeUHc2zi93LFMUkbESshYu5Jq
NmIf0lbn5EuBZH0doiCQYD+ZueMkf4YRe8+XWmhfAf+d9crOTTEkg6EryX8h
8zDNk71vrE+6bwLoXfq2U1xVIXER/LwSauoOu4QSCeA7r9IVWw/3LO9hDzqR
tqizGpj/ERq7syhFJp8F7sxM35ubDfZhFJHjhjpGuxAyOQscWSnvLZ90D4Hl
bEyRNNTl1plNBTgOZl1AHnQPPegwYN3dr/hTPyacXwQGgksnrr3pTyw/2F1R
qkXQ0hGP+z5lxhIoRx9nQhSjGUnzjDBmo+tLnrImjd0erJSSx6danpzJD2Du
6vS09US65fD0y17ciwdWboPz7lVZL4nJ20+olSy5Q+aSE+WZJEuPkc+UwsSB
ffBz+qG+UhC1c+DHhSSeZZv8IzL/RHQnRjnkINQGOxa8iHK/3jvRgr/wvM2f
0ZBfX06QQPHXp1bIkEpSYOrRJv/tU7IyC6TYd8cdPcU0SOPYb1Lz8NHDZqX/
qB9ePa855679DHFCGGfGSwkre7bHOi6ap84vhaRmQIz/fKPtaTwltMkP2crX
zRScfkzTxsZo6er4BlmdUfZXR352Zq4qIFeurDTVEPWilLbL7nvTqlwFGJhM
FLW8liWw89hlf7dO82lbUBDQrrwqHiE5nilkZH+iWr2iJuA2iJ0kI4R4XakW
VFEpm1pTLlZZfTYpm9MjxQo0X9KkGBCV/sozKHJ6NNopuzTM7YNFGEwFTv9z
ENucDcOpp+hBjYxVz839P8rmm27UKwfKEVtV4NtQm7V5xiwqLhHsp1Q2oAxy
SvbJEudVwWCwhta8kp8T7RNe5/Z9CrtX6ozUZGn50s4UE/lEQTlInaLpOPFC
8ACgMVUyHN/35oMxg2dyHuOJ0wiF1r6GOAQ3vTrSFm8sYFIRMe2VmIG77pNv
dh6GX/xL7Z1jnb5LfW4Ri0QL0msjjgk42Rdlvd30WzHf9k5ndJfV+ga8nMsh
rrkAhkOmNDRS9vbDkrLvAsxNjvAzLq6ScnevE3DeLKeBsxnPAnqKPtWLnRY2
zlGAwrXn6ZxKYtkZWQxbMexsbIKgu40spJwQWzBQkXnDoMwz6XZFYj0thI2L
0DqIgeWq1b8eY6/kOXkDfE5MKVm4trluACAQrjgsq/QREs4UzrRaP3q5OJQv
3t+FlzRJOBa7Fs1VbsAGcHxXD0vHdx/NDlUHdLVE608l3Z3Ej+Jpw0NvCLEC
oZ7ZY2S50nAC8VUyL4mBW5MkkkTKfDsTLiNADYzg1K+ualhFtm9uZPAwqL0x
vLuZ5899S1wfSB7SdstJrpe0OIIy0pq8o9CmPuU5k6J2i+gCle9di0kGXyHW
Fg6QX9vSlVZiNKGECutsxA2KTL2iZxpnyguKCnozTtOHFvlffCDDrtnXVatm
RpiQkFspECoDhNTMKBGX7uVYutjABpUjQ3YjPFrGpNV4d5fQtCv/xxwQh270
OjuMzPni4+ilqKhW69C58sIwxhYZFD3eJwexYs1fN80hsZbZSBt8xxCoBNS6
HuJUcuhcG9/NpMGwTzWs1rErS4ayn9Qy47eLW2XON3sxREYO2KqlHvDGw6h0
l1tdKECMo8aihrDdqUdM3khfjht8xQK0+iin71S34ywqa27mvfEl1e3DeIMP
q0fxHmwZNyIgKDH1URYAU1b9EqJx1Yi7bwqAcS/ucLBw3g7CLIo4EFN6zU7K
wEVmPbM8zVYvAcukP2DzdczZJeVPzm4LSWCm/O0V3fePHc6jV6gglu7uNVzl
t+PXQPPDkP2GSPdWdOSDr9nq6FhxtB5EkMESUOSfxvAmSIKY0WJ/sHKUsGhW
AJhhmo1XAouWwYYFdfGAk6Ip6iqIw9oPdiYBD+/l7OeM2PT+78qqYIEpYmXJ
ZlVB/1Zc9eQ0V0z7i+xdOyvKjgNJIRnxtFT7wvz4b25cJ+24DnKNT6Fz7BwF
uEj7F7Wu5aHQcc/7WoC8UESzlqB9gX6VZvpEyDW0CKttO414JqM5SFK3Xl59
Ii+MxhxWLCsqGku6X9D9C+Robfsx5fM3riNix91KWy0cqrDyz2PojMCFhFMy
EjrIvliLBVxFZ344JebSSJlFiciRr/cisOAxZVuuYQFeuvD+ytBIdNXuaNWS
mmWIwga08EfBLDpl3icpv5jckjJSJUaG9vGNI1ngLLQsFcMPTzb+RuA5E94A
3dYX8gGn0R4BQO+FTWTWSP9o/qSNqThhZAcxHCHKcdD3Wqy3/eqvFrIJ3MXn
+dGVZV4anGRJtZSDXrmLmwwUT/KmvpveYSxeUymiT1AN5h4Q6keKaBFzjU45
m4Sp3xjQOjunKPGGsNMKvfWFqWd8fPVh0zF4z4Nu3nXLlncs0XMerK4TGUob
bozQz0IenliB9tHhDrmr4f/ab7tTtv8+PzzBNX1uftL093XozmzvzXZJlYUV
wYIdqvo2fF2oAojHOIwGVbs0Z5TAXdmUykTee2OH39HP0oeYoFec86HYJU0A
j1rk3okG+yDUE2Fd4GdCGXJh8uVSs+kfeAl+RkAwJJFs4akLCUkoIKZjCIiE
UuLID3/2KG3ybafEQzxlvfy/L49WTJVHfkea3RAioR+s1tb+gAEK1QCksueG
xMrns2BntF9Q6GzlJZChx0vBE1fgzGnmM3weDgStfYBEdLEHBERTMHY6ZI1Y
sZ6Ig/fF7rOq8rOn/KKgEqrIyANNQ0hwTsXLlLYkyHFkuBcVWyLy24BsTIBA
VcvmyNRAeNQODS4SzQ8oeNFxGBoFK09bSomuNaSaDr1vhuCXr3yqPREsHzfM
7Mu4IAiWyHfKJJ9f/aBzVaa/3oaYb6y139kVc3+8wTsDCp5XPR9fUY8i75UL
KmfvdkR3Xy2oZa440tHskLYeWX8CjhL5ycQd/nEIlDnIBv2bSpXreFjmbkm8
vYdRaTLe/wKVE+b4V43LEjcAoFHY5MxmGCfjFYPrZTkTLeXbV4CFuWMp+ehu
/VjdJ49bmroBUB+/C56/9xxHp3+/jifODO8+DPPxtf68XKxSCdOUQ4AWZvMM
wkzLsCvkz9HKmS8rQmrysKlLaNiM5O37tpHuy+fRdODxW0t03lUZf3v/bu3w
dQwl69nmswml27FpKGIztytmbwmmjsXnEPU47/XvXabeDIEoivjQ8qSAfTDU
/VvsHVfj6aH9bBC0pgvY9dRPai8ZMKB7uaVAneLhbBsXQU5lHNW4gk2VCLtj
tAhCV7TjUx8G6IyO9YiseyYSzgjd/OjBFgrpmMDaAikJACYqWt+9SpWfFi6b
TL4xaopfWDHMW3CWfBPYoINpOYDatrLz2haEz2H3fA5A9lprX36k5lX+OXUS
7iFU80YO46R5qt1stDUP2dKPmbEIf5/IrZ0OWvFLLI1EokiGxMuD6BOCLqBH
32/dWp7bkA5TeCO34pEbevcIklofyr/MljBFqf0nwklTV3X21QNQ4hQD22V5
ev7F2HC53wTFQ1xu184JwHcXZnIEmWQoZYNBNhcwskrbUs/lZOowc+RmpaNg
hbyCph6TdXof8F6Qgez30NqYRPuK3SZ7plVwsQiVzVM98Obc5PUihOE2he90
z8n3OIr8tWVQa2edb6+HeEtb9YkGRbxMBRHqIiYxSvW/b/OJZzlgIiuaQVkI
o7TkVVy1P/DADiTm9cV6LaYbj/AQtTmscOYMXrKNTkqiuvq7jVw3Nm0esLDS
I1lh1soHJMJbAhuV98fREoelgjtu4mTEwXdrp6t7cfcaTFjxCmGrxQbTNCQt
3EdXg4vvjqJqXl0gmXRoATkygs78CNSORLo7UXGOcPToEduCQTxnO9E27I+i
GcwxpVr1nuJCkYxVYUz99Lu6eGWGrO+DUYG4Vw+BrXZmcoK6k2I6IJEJJZZa
Xm/OgbvK6+OOnM162PvIxjNAlQllwbKGMpTTLp+TmqgIgwpPjhcvZ4z3nqH0
MOz4qJL+duB1Qc2Jou/pPSi04H0RRBjeu/YfHqw6A/f/gwS/v5dNVwkjMY2x
SIDxcun3vO5ueU3sKxLHICu9nV0IL9LN526OsOcQmM/FJjCnkdWnx6KV8ryu
9hD1G/UeIzdoaPG0dsQkHUMXz4uZDQrSOOB9cxk1c4+gMdxSYxMTegsNLPhj
hHi2la4=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qTSDP8mpcUCiwvaxwJcaPxzpz0z6aXrqeH0KZWrzQ7Gn0jpb/sp9lBtnCpYHuEg5kkVrI1xmgeju/3bdnqw7WIDXUFvBrgwY4CZ0jYLikmgk4ISEaL7xqZjwJUWbG4W10pjBBB3slX8LoMyS8ttLE5SYDHQh2L5xBn2Rh5ofmpW6aOO/u5ixzAxFhT2qk3kteq1bOhoq6021ryrHP6OCX2HgP0nFgQe29wa0whHG2W6SylndjOtedavpdQVFyPEP9PkChD+FrtjSEXxODFoli91vIRCXMiIwbqkIMwr+Xiyktw74ddu/AMtd6+9HJSa5BlBhnkS687VuZRSWI0Oy32+lEYFG444z7G80cDZSssL9CPd5zZfBBoaDXDaM32zcfWirVda66BN1b0rDF2Fly0rQgqsckb9Wa7aZEnYCtwPcAY5vkQ+3ona/tg2JykRQptrqUcY5NWFaLHI8G1NNh0BXWiVvvDJequrrk+Jt/9AgrFQOgor6DBPq92vjegfa8vi0PXBZjHqJolbsvmGWowSDrw+0fIz//2uscUGWfedv3BSrhCHYRGvl2q1wVe0IXnmNZwDc09I5OEogk3NEWQ7LQVrkp6vUtctgk+26nLO+AxPB5b+YiZW1CkXL8kTSrMb6KSBzkfHlJC8HG+W9zHrLwcn3EtiYLIBaDjxfr9FBHos9wNvpRlv2a/xuxUrTq6SwSDnvJlre1IHjuyj//5EB01AhkIzxqTdVvUghkpQJ4Ia0fOgL5vfHcI6Z51zwwDUwzOwP6gW/ABlO+LSsnRS"
`endif