// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0l9r1Bz/DfjZN0P8VqQTUSgYG1SUCKFHi6zvBhfcHLkKVE8vNrmftx/jlY0E
MLLdk67XYNbiY7rwO0YGgMUSGYOKGmLkleQ3WMzPEahQkgOKoqRlF17a0H3q
y3RUPJwCj1LQu6DCtBBzBtQYuxGdkznKJuL1ZApIlrDNUAjooJ5aSZfKMHzI
8EKqy4tjh9fa93u10f1V0BB5KUoOC757F9Xw4ifKZmh/NSL4lvw5AUOmkaU3
jPdk/wEpPcpVJrRAs9rb/2tzcHDCxjmtFOsKzq7s3QXbWAYd2/vrF3lYnzVS
pyh4MB++C/mwlLgca1gzgblN7sf0XsU+7YKCVQThEw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dreIKwMf+5Xlc/VL7j0JjJuqFtwOhGdnHNcTazEvo3m6MrFc3uXQ0T4N5tzV
XGP0oEzQzs6c5DZpujew2j0Q7URnj6CVpwl6X3XQVRHG8eu/K2bWbKQs53xr
pi5ddw9asAUNkBPwEwebVGlZpjWpq7VbABmYKvNO+zUqbcUjrU6BClTIOCEC
BkcCTATjYZ6CgQFaBHoBZyN8zGIUyakarR4hTzrgh2K9U5mh7wrqVig5MX9H
amF+uobktX6qScNjMsAbV2GkrGcq5/YzPlukQuPKC4g33wDFFq6z3ocGI4hh
QGokCIGkSyuvGa+lzE2dOd4kXYz2/HfKsN7pYo5mWA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ixx9iayETRYJ1Ayf5nc0Jjk6L17zyEMHpQbUv2/lR3kA5FxLAcfNQ1hAwf8y
ROfde8JOWK0eHelSKwSYeSRfGqjjcS6DNrllEmU0LBEnPd0yfpDfr2cap1h4
RyVUhLU7726YflU8drq+/czeMQF8B1ggvr1tBiz8ruBPy+N4SfRPEPlGiJrE
YQE4cWfA1T11dL/WwmUvJ0IFcfveBPvOHbY/Aa7GJlm23EVJpqwBS13ZaN8p
q+n5Ry6eh8pbaDuoHM3+WehcI+maOY9pk5IYQOcJrkZoWEMgZDSenHXDMkVG
jQ1l4hDMPqZ39Qo7Og6eZ5E8eO7RQZOxW7BYcd/tpg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rBMR8LFdNdn2FsaZuNLUyfopUteOG3bEwK8ReR8FEgj48Au5pRvE5YdoKtF7
iWjmk3m4tJk1IIFNFaJXJPtaRAXR0TJV6NpXN/OgZu5fNYtII/rLgOrhOH00
b6F8hQ6WYuT9pMWlPqGHerCcB7XC0wZk7QExEbW/B+IoDROGaQDT8TYYTNKx
Z873y2FNjTyQFdsvpRpaVUy6iWAbv3SvkB6nKjTPp1T9sGgOVK+pF41Hyrm2
Hc/IY+VuSW9HPcIoejrs55YGd5b2CbswlVUOsUl1zp0E7QrbPQ30zH3oZB54
NsUjPs+G3LDQ6sV6CeWPUQRaLu79ZQ+BpHAdKNr/bQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B2C0KhdDPfS/PByMLgozXGSS6BT5kIQXpifWgBL95AmXNIMC9tof48J+tKnp
2agkGAGsw23/bnGQaeXs1coycVccFuqFn1ErreJpn8Afo4QiPDgNejLJp5M6
It60qv+FCzpKSbEk58ENMpW+96krMGtiFsKuhWgOfybE1NPLS0c=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
faD21ufM11YhZqvCeFX0D+ME+12NCOVJvfTfNxX2yurhF4LeEGozxCs+N8RT
h1YFKIkBpRIsFsXXuKSiptLGEAyEYc5KZsCf5wDJJPFyGlWj6H33x2rDp3Lf
hjumUaRNX+FE61B5owD3uSoyVST4RKB7+lKthiqAd7Wc53ObkvLI8b5T2RNH
QzJFOTNwWKzFzgJKlS7oFcDO1+l03LzhadHHwkrK8MIfQZz/SD+FCtWXFmaM
Ttks+TUZhO4VJCU51UUGw6XiFPmNxK8G5r+4RxelBnn6U0WwNu8NbhIfmYlU
EPKPdEspWALTGxUI3khiQtzauBZYo/PYoBQOuqa9dnlDKQtKIhSfq/vyK1bm
cwbxwGD/QT07UMa7rjK1F7rAJkyYg7qV2+arqZ1LHlZaKVNcB0BMoOh8DeIs
dzyWpdEeK07PvAZ/rklrK5YBZi9pe8ZYK+qAr611xzr6l86XbQL0h75hUHDy
gTHcZUx25NuhhrNnQVlKDylPiJzdx3Kh


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VxhQy1wxPH2/geoQamEvsvBZLdX0bRI80Mqs6Eerw6XkxympGJM5KgoeHSTw
VcqvPQAcJOB2keQe37hpPLSeYiDd3b7Q3Qi1s5JRN367HEA3X5W8fVBgj9Zd
XEspjzX44TzX0mUcQUr18Gq2TOtLmcnFautzpfAF/Sc28lrdQt8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NKtO4WbFLC0JdzbVIMjtOS5apIHFrOAeyr3/fV1qJczOBBNtfKkItNG3fjSM
mcIIZoMXhczwFs9cdQO9d5akMkBKCK5RJ8ukHIhXtfumAJbws7C3T6htt+i0
GAUNlttdyMAjUiJ5sJEdcjyKqMxsk9vLTyXWFSAZAeLhcTcozqk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 84400)
`pragma protect data_block
veifpfo8xH+h6BPspS2/e7DVnVs6I07g/8fddOxyr2skTWT0EHEor2xPEV4U
Y+Nhzexs0ycs3++K1NrH2zHTTyVXWC3rnECO3zDjIsb9aUOgeKXpbLULIxgb
wTaXmrqGw3e212yUsWtDDDDEgVrC0AYxuAThyTY0jf2UomnCWc/5+nbFVhlG
PIQTninGIUw32Zumgd8gZw2kxkbFU41EYNFTdn/GJShk4AuqLEQgHYv/ADvT
qhNoygzufTw6ZlnskYLjZsRKE122dSWv+CX23qdPYjcorjNE+hT8miGm2Ez4
ZfPO63r05BDME8uRGf0gWfIXCHkC8cOlGHo3s0JVoPTnusqATuGVmQXjYINq
rxB7fej5QLQS35/i5PAPtJOet+qGV8fItB1JaiTtYuUR0ed+57IQo6Qyqq3w
mA2qSSv25/H8IW0jj+7B3+SMGc/wdPImq1qRRm8cihN8Tf5nLPGk3K6ylGNB
UjNF+lLS7EGCnL5w7f40Ep0+iOWs+zyRAd1UEYdz22WyjGNTHogJlWU4T0/q
pGtkf+2v0uAHis7PJ8Q6OUkL1kyMoQwtqh6g22ZVFRAKAG6XQ+eM6kCIVK7u
G6Tdzsu0qwnRIrEccXvsebrtIlLngPeoWJ23rF+5rEpeLivF026h2qypfGtn
elhnBhLngxeNx31/kqfCYVTyfQOmXY/iNtWDwCH8JbfPnRJiwK2kO+juIpp3
/4d52RXagFzcDT6zTPMi48Kn8ieCWlaF+ReUYOT19dE+dBsxywRzG1W6tkK1
ecLpoK/xp1dh7CPewsZNH4RftxW4cjAGLwoeprzktP15BeKnA4ZS6qGqjTvr
GL8QryOMlpwaPLz6B6irE468uu+AnH/7KuAy2nDpOZ+Oz/Jn3EwZ/Shuqxc3
sK0VfUekMCch7ShhArf2PsXJ5+PrdVA5mQ//WyQDeNGos+bSJ9c0CYIOSAGK
CWFYmCpz1igGG51e/e9ChR7N+psEtmKFbOOiRBt9MeMFb1mFAR7hVA7DCFWk
s/1dyiJIefiVk0WkNGEDZSSzPvgevBJ0nB8QzvPPJtka20mLZhsVayQIlGoR
/yUr8L6L7bqJUVlPBZ3InE4dvqz7pcHkFiIMrGhBKST1EAlXR3GQ/fBSs2QZ
TgmVBe9Pi4QYYs23CH9ioSMCKQmNgDzwb67Jd4UpjQIjz9HM6rZFiMNlDm6C
74KHMhVxaDDo3h049MHkk/vGfX0UFqsCxMxeWDvbboz0wTT7pQ/4vwWqRmpI
AzfT2hBtXhrVjE8tOs7ANutFk9aey4ZPOd0MEMzPBYx9h8JxQ+RMde/H934p
gbkOG/Uxr+83E1bkidpbo+ZSMyESVJITiITze8DmEhx5B4AlOV6iIwXwgXYj
i3Yh6FW3w0ElPpUnT8oKwnsL9nL7V7u/v0VOjhDS1EJfv4umAPRVfNKz4M9C
Zxs0HfxYssQvtKn0DbGeElzdGRU7IUGG6hZBqWh2Mmou7GIwEUgjfw+18BLn
FIPAJcbRpcC7an8XTQB5mAqxP9k2dPYJXHOYfvlxsY/y74YbA4IurXCngIDS
DM5757/yFbh71FjsYDrBkDXdSuZrOCb/BGuJJZ+DpG2oDjY1/f2aOZqWU8+a
zU6a/xofnzRVDVJfAxBcxUzDSHFUzh+9gSFw2d+8A7AUDf8AF5EkR0PxTshU
hfsWlf4NhWqEc/8vFL/MuXwf/FW2ThOibIqdbibNWEz6CnbcPU/4rf3Vitu4
sCODM2OttUcjc7Q/bKY7zzkTPPI+jMJ6OorbW0AB0qnPmvKYjxULgci+VvUu
5G8grWYQbdn4pzhZrTazIMtLY4jIBuCx5CBs1b6e3m7eRf7ok6r4oNNgx7gc
hvxrWAzIcOMbmT38pWHNZ9+hoKgDwvyUFDOJvEN5Bk1VHTlWX4WND8AHUfrp
tGg9+nqIV0irDq7gQO3/QoKreJP/dgxoXKvyq33gWmjYAsg/+ub6ix1B5mDu
hkt+mSA7FbH8D+vsWGYO+vwtYpxNeBmUwKSufKmoOoVU9JGMRGHsowYh8aGd
GLXZ60zmikBENoiYol0Q/KFGU1ZKP9P9hjwap42lb8he5qVUG8bAG376dJBE
mc48E40ZPVJISqi8e/Qu6QjVPGGbE0Qy2iatvBodf55dDY9tW6l5SWyOYjdT
pdQx1KT52HiQyhyXu3+DbEFFoKp+LxSuv8vXK3P8Kkh3zNcAsTuYbZfRIbHq
yh5UqChpXNHvKP0klR8eBwPOYwTGe1XdFbRU/vaRBzo8FzSecy7uG7oXOq+S
wXUhXPFeouOO9NM558VlHARb12GTlL3PQl4sLh8bGcrP9SDsWvWxZQ5DrS/t
a22t5WGC6bMfXFzObwU4r/wT5yNuNAoL0BPtg4KxXQncdegIYcka42+gCmjx
IqjN0rn25EdOyJnxuHvRch9tnbHjKfvgmfjf13JYD49A/YHrsjLE3AQUzL3l
5x6owc53H513N8pMBhY2fjjAZxMokigTof0as5UDC0hJxjUckbZMC1xVgI6K
HbZsvYsSz3OyFoGb5CI5jF9IcnTu7x+vCy5GI2w7kA9tdZX/xc2IumWlohOu
jdVidhWj6GuIQNoSr0Lnm44cY6i7rL5rKxFP6SbY4p0eS5HGfUaVVP0ZpiCB
wPfI6y4RwIzqxFq+85RdgEXMFkMs0OCYwvWx1ulkaQIQplqCkQDwPMsxLX+q
yV3hLvrocN4IzQj3fOsWfkuDexsZaV6hpD8Blzlu92SVXaHk89Et13m1asBY
TIPfwUUfYhrBsq89LRyip9erTJiJemDNgEnAvpHd4xIwAGpssTopf15W4kZ6
cIcRWJyWmHc+6D6Gv+vuD/rn0LMZPRj3KZOK5YaXHxkQS99zHj4/iMY16XDU
TGCqNudwJ0QxIlYbv4a3Czk9iOwaND4uO7VEsk/FZWs61BgNgGHi+xbVlEbk
wUYk3ShdLjzFDDaKRA79hU84fQAtYBbjnFuykN0/0t0LBXrtc/dvIL7SoZg7
wi7KbkBJdX8wYYtKiRsqC3t1OYEeoFWNRkQGQkerjlNaN+yuQnWes6/NE8K6
y4lt44Ii1imSeSts9e1k3PLnzXkDaooZj5WxgMQpFjGvRHKEjECEVU8AcIdd
vl4iSU7PCkTQdCVID+SqsB3adgNyxCaT1HsHYDY7muP991ddavODM8Si3/9i
qaxlPF2OUHpIE+d5ZSbMTYccF9DFdTVPyQHC5meyu5cnp8VsYE3NscGiW1JS
CZW0zT2jvpodYPF07ZC8zFiGqoKgDMMAN0jrJZvYwymap2uzTCSa1lv2X9Oo
VgGmp8Bh9uEJb/69WC7oql9qey4r4kxOWy18ZNWhzafpcebTRO5HEBlAs5m/
+5r/Ii0BdgoPDnIxKNV06P1hDB/HDTJCUyCSeE8FchRb++r/4IWMWoj2mqrd
xY8AlxeUT5SuJHK2rRFmN8jXTKsL7DpF6tpBnf4wsju02ey4aU1vcrKrD9oU
85QY9HEoTzH/NgEdxIq2LpCHucBvQz6cNa8E42Ag+Fjhxegf1vopt2zXNS5J
vc4I4qYmotkDsaUdCvdMqaNQ4FtIQllpb7SodaiW6Y8HkWXf8WR/+Dr2rxMk
wPcukS3Knaifnk/ZwnE1GmwByuKpzuG2XovAXF7xkzO9zR1Po3OqP4t+Ia/3
TpSp7RCD/EQnm/Q6IPK53VdhA/WW6mleKwIpVW4LAYZ2Rrb8KDFfSb2ZP0HL
QBT6B9wx/EhjvBVkb1DdH4pSFzSB6E0blhV6kUloP+mRVb3wOdVvydhINa4F
aTQRvMlt1TuVZV3ork0XsOfQW9T4lCJystB/78Q0fSVQLF268VVEXjBSoxZy
7u6U2L6LNhz/gmZzTNyZZzqAgJ+sLnOlozWuRRex+z/uPUZrN+pZL49xd8qm
zQxgkn5EaQkxPGsMgX8XJ79GKtSSBQ4WBZ71MGco1kpytRNVT8z1extOqpcM
uH4+hCTacR+4HFAGlyIczerCl6SlqWo4eCN3egNs+QosPI/mB3JbizZJSjpj
Mjj8ieSybwC7MaZxPdWw6K04Vcs71H+T1C7bootiQsh4veO9P7s26zuZ/o4a
TgOrb2Q98vmO3lf3QlySOr8Ivz/wkb6tzTHCINM1TexoXPGh6tXeCi+BEQHM
INLo8GAc8ReQ7tol5wh7lZSg4KLjgPf7BpfFk39mOIYZv2E/rtfSG8ZYaPxq
5lIDf2urwLWrWjDEPgfMakL8oJp3HqUQnc8k2y3UbfdMWeB+61JBbgXGgSvS
w/HRy7wN64L/Gc+OW6RK8wb4ZVAI5eipL6YOCxZnnyOwWjjQSLtRbV4WVkZd
LgjKX0BBJpcb5XPaFUSg8iKnvx4/7m666hBw6/yJ0QyqVuP3BOhGcySpYccI
yYXNf9aPkrtuABMZegatMVHeG1V9Vzt9PwZ8P2yGPJtKa5a/wlLm6EuB/eiR
MBfhHeZp1f7K5yCu/UXNCl6GEjHd4UQ3eK7hf8JkLYcAkHRX6kSIAWsLIXo1
VzGvtwsNGc55jVCZOhJ5BJ3tcMY9aRnsqQBbJQjHsH/Yk0F3CSlrPlz1jvpC
kVSRdYCZE0zcxv7y58vBao/6a+1KDS1b0NqPE4WROe6SGpJe5Y1mb8umd94W
KPrRsE5op78M07tOhi9OteaaeES9J0Owb1aZWw7DkGQjVepwYjsyCCQqRf40
6hGf+XFE6R7qGQ4MYYiOCbVJ9JE9PUJdvecoofTbGp24YmFQG4qaDWQ0i4ds
128XdPMpo/R1b4T7D1eqBc3469whHEyMAnSQu8cBvI5+8IjfNvlrDUPgf64S
tzTxYD6YSxo3BwO/Uuu+3AORSmmZBzlyoA5pmPtJSpCD3kN43l7nxc48vMMl
WGHSenFHSnZSib/qFIyXp7PULu1u19Wf9WI3bjqli1oB9GYzBjoLHjRiA844
WVMRQTNvlW+q0aq/MvieTQUTBPFA7v9YL7s+RtOBqRyVkYTf7VaBORZKkt+f
cYo7pXmz8UtqOfmUEa+iIa6sKg5THp3914OAjRO3Y/fKMTUs8pe9S6xURL+E
JAmSi7yhf1S0wpj8p2t6qVZPF/omlW2uxhWN05+/zV47/1BwDUWjnhoQisnv
X2pNvZbNiVKHvxh70WsQpoAPJX0N0XC1XmYkvSY39CF3CfT8I0QSMOXWZdw9
E7UpngMYjrTPcHYApE/qKXwyRiyuKn9kEd27dn+iXqp3ikdMTwfLJDrGQJ3I
0c62/f08AlKJxt/apbbH87IrxUZEsckfrMW5AaOwnPVPWBZRNznXbjEhyhP2
76oJreVgd/RKyeFFomeVPUULR5yXmcqfOMQv8uIGY4keCRkKtKCxvGUjRJ9K
jQnG+pE8yo3GmUfTKParOJ3DCqWRHC7b53nmaLzpJsi4VrydvFeusNt2V6O3
dAbMMkkSp9DVERkJj+kc5OAiT087YkxDV1+CkzI0sRqdYaoO4rzQZzFgb8UR
TuvmZay2FkJfAF+6qohv4aOGqzq+jqggCm5XG5iO4HCuTJJJRZfavrzeAsr4
kTOc8SKajfH6ag1jZMRlYumTMKs79aMUqXP26BSYy3Dmb6aBdRN8T5QxLX28
1oOOzXtInafimfidY5zsjLGm6ChkW3b7M99DKfxPxZJ1Sw8CKMX2titWAmYY
XDvaB3FJgyCeWzo6a782ArEMdOmU3TXs7aKShkKVoAkyNA23xvle96yOUVE1
oEgbCD2IqURcVm6vYcp/Z2bcGsYxPLuFhfOgFmsaGUSVjVvGtNRPgi/Wb3Vn
sVtsuf8D6jwLIY39V3lXbiq/M7WJmR8YOLoE7mrAKC/U8WtyiRvWaC1sSmFQ
Uvpgx30Zwg4HyuxJtFNOBA+Uhvpmeu8SoKouuA2jPXzcvTo+V1MD5KIz7g5N
EhRm258pB11wNWCkXoBZnib72nxpWfk0q/0Yc+wjacXTaoL/QQxZJRCzsm2l
y0gYwx0cVcnUHER8Eo4NJOAsiH8VzVG30Qr4ix+8PRl3fVr2hmAMAODvDyUJ
0ZpPey2R7kJO/zLNTwAwPh+jOg5LNx7EEm+kvtDgpWQxAs3ordiUc+tRG4bH
F5Vsp8of2kxWMEnkLZ7x31tXQCOSm2i/GaRfSVQ1flUljHtcswzDLS2EigYS
FM0VCgQlvmmIwK6/gvIzLY9HFbY9ICRGhV8bZH9o6i4xJBIm4+Lxqe9TzboG
TRJhmTlRJ1GLNWHxnJGDD8sDUYBC2imtMbbrWcrW96F7E1G/N/+Z5CVhnPyP
pLwJqAYOsnO4oZTHqCCupBZ6h0eKxtyg+3MIctIGkpS6rJuXvzVxRsYOpASc
KYsXexgXswIZaiZz+EfzwZiL2fAL2s6L3srkqVnaK7kTVE11m+xq6iLzc1Ts
8R9BKJeRM8Qf3kt1F1oahknw2cnjN6oqFqKMc8pfKOx/7H35OLfn+C6HKe0B
hC09tjGIlUNaUPbHNWAlry2YTYHG4Pmd+QGE5Im0dXCtmNZK98dzSE0kmgWM
91Vs8MAWcaVSrdcze+2dJbaVoYcdzfOMLHMvcwDae8Qhd88r7lioRV5rTBZV
CEWllMUdV7pPe1RglpfLSHnwWWTjaVn1/flMFDiYNni+53y+D8BULFDhXuGM
LH43Nvl0JljkPl4lYmsAD7XxHXGTAoqxIJYYV71ZDjQRX0rUczppHdT9PRq3
XuQGKf2Kr/mTL2bAS8uwVEeG0hDHCimq7HRydSTEDkdjop58vUWQx4+O+our
rlCp/RGE1bYIz6uq+49FmtmroAdt6KdZRNuic0AIR7ZPOcHj+0wMJ+Ja7+4C
vstsX8kEju7cAQlAImJwNgMKISnXX6ytqKewLJUHUqWAIk7uEauO8NN9flYW
RGyVO/ymm9qwgBMUam9OHcWmf4VkRUMrHbAV4mNNyxBs95bNC1ytC8hdERHp
ZPS8sapd5dnw37gltpfU4jlEUdDTjapCDl+JkvAcpTJHSesrzWLFY3d02JbR
XGvrNsrumN8v5EEAPClWONmwYtRlodt5yLks06XzcAYx98w86zWAUznyBbwC
v8wqDbt1cMoNmYiyrV8n9OrjvONX8dic6Ppotf4iMpvZW9l60Tv052fIhZTu
OvE44gqwPgFwWAgVrFFOPnuYEex56EPR5aRO9Ba8KkV5xYQq1rv0xXoEwpP2
C/0N7lD4Gm9eWf23l7SLtwIXq2cWHmjjedtXIc6hoaHhp8GYCswcYruRt6n7
Rj8esDQ22qYVyH01YVkzy7YtzqqJARn0B4Oc6b/n0JvK12IcHD5Lwop8Xq8h
dGxpk6ivdv2jlZCUkp5KGw+Ld+KadI0b7Ua3gKdnvAdzUHrYV4QjDb7mPNIW
8UEPueNAMz3TF6Gmz1UReY8SsyS7jnUJOLBC0qhrd5N0aUkoBQkpVoo9AH11
iJPK7Gww/3YkiV+aUhjBfJ+2sqopiX1VLR41QtvKEjlzOFVyWCMeNX2Li4Jg
0IYIEoHbaGPOFna8WqGdfKxxVR65T8gCaXHSq45FvSzShu7+5j1FFIs3Qu5f
0tc6oOucuVZu8cg+jcpc+9Kp2e3kDm2n96NG14iS2gUYHxxN+IJIrjzdBooD
wHef5O8/K/cBaPLdTrIv8LSphANPigW11DPTO9mp6cZQ37h0/X5XS167LV0g
BHG8CqE7qgEb2EXdWeVeXzCmDvpy0XT4378ZpFZzntCbqocPwO6os3laVy0J
+x5dKY5CsNdnyX243StayRiWU1U/N7xjVw9HXKz+rNQrxoDKhs/tv28ihnPA
j/kh+Lp9YFcTBocfqQctTfAF1plwV3+QShYfiY19wR16Fqz5xmgCefuB4WDl
M8OkJpCeHs25MW4dZUnPTN9LpWaWZTOnrJNs6sZo+Aivb4BpENKXbOrc0Ntv
OLcs8jJnrvrnNfD+KRIXP0Oi+dQFKCpdrmfATFXdlJndwwQ96aNp9LRRk1j8
6ysxy4qzyyYeBdKYc3GNI7iqUJOIrmCQBRnZFJE1fIvC9tcL/oFrN3oJ8B05
FZQIQ7MknO6zjm7vcN2kFpYB89vQya6srWfS8c/N2eX0aIO1WJvvcd6Vl1qv
Rx/iP5s3UPAH8aWmGVuxozv9q0fGrQP2RkLBDplJ4e5LtUzQcRaA1h+8Em30
Kaa2YpMjRfj6syOG/UKSPDA68d5qbXgsXkLrLKmYaRiSgRJJui/38KC4bKJE
OV57/fjnj6ccX6PCoZxwsivmt3GXwShkUGZQ0q4P7hlkMwUQ78IwqRUAhSYq
t7fRorFQ+/CnmyB4t2/4B9qhfdEvvj1G6KFI5rVFA4Lj0yslOon+IFCgR++B
OZ4Jtj9zypNXCichEr3XLkWgPWDJ/RpVWElTaqvG2FBLKtQ7Ys4jo7NOVsym
0JYAi372aKI/Z9uO4lEbauc9fFcdwmKuZRgPS06ffsXBU0/wupyBrxsUoMXd
ga/RNVDD+ze+bB19DMhl0koe8jjFduA0o+2oW7BWvxubFz43f6dM9CbcsVEK
3ps8IlRx3AwijvcCNIJWan/3ETfBM5abhHgLvijx1LTWDCPiteLiSBKDiK3T
JQLNXjlYPc3Y7G9kwp/ugk7aikUVpnh0ll4NewyLRuH2m2s9jWX+Y2ojiVsU
FzRc8hzK7VQ68eZPcxOTM3nrkoi81gTQaLGaBruor0LDsW7Uv9tkvDJ4NskF
qC04E0laZp7LoP8Jt0wt6nO6sl7CWG5jZQDikP0HCsDg22OUeEFgdv25gNwm
AlGQpLo8zfWnA9/cpmhhNGJFgHvnwmVg4yiQ7eErxa1lmcWTfYt5+YniEt/e
StOCOhUpOuMi71nUmG315huojAuTQMmfaaMtcNuHLDzLC84OyPtKyUat6ye6
TtCPtytWzwT7BNBL5B2hBJ4xXG6UWt7bBpoorbY7521SYKWpzheorJvU8Yjh
FoR1WuKY4SQoFckqk405sS3ZB9thbucrd5W3MyJxULk8EYMkPtW7bcGKDwym
08cXWsqukivE7fTI4VLnYnHF9RRfTjt4DGEajccCzO6s2B5T04kM/qTgEfdl
HQofscGGnNFDoDvp+AcekILfFKqFd/bSR97dw3egwMxuEo2pQvud8QF8ZSWv
oXaJqHAtd1M/d/ywIjx3xFgeZl8OYpVpUPYrmm6TvqX/duS2h6e8dZbSPvs9
elayrxhvR6x2pjUBDRkw+Hi8iWWV0u2/KWG4eX5hw3KHdU1qR6gU6c6b8zlb
hMLFWe/yZE4m8PB8uB24CX1I8knY5QFbBOaqsqCZr0WPrIDtdGa8/lOvsiJG
Eit2MLmF7GYWBA1Srv+SCRZGE5ls+okC5GP59ipbpl1NRiKUP5S8dfSsVFlk
5sVplg/ztMfigmXZIzgSFlyReDxvKS9xQiUPs2NkMgXIA2viqlAWkEgOfMDo
EQuEZyqSDTBCbWBAdOBaWqqRkpKuM0xRn48g7tgC3P2F2LdNA6ywNazPTZW7
zbMptkB1M7/3Lkq+zFooT8veaLXEk8gCyR71teGOobmHovGK/rbAWY5UyCoA
W53E3dmESyO+K0Tzwuo1v5oTc1Sx+laCQ9VX6U9EyvmTZ5FMfW/xksrZtdFL
WqdcgvQQOru+t3plG1sK+O4wFlFRvnW/t0BWYWpbe00LnmexQBRHQ5w8T8Kl
5w/ufPcBQFFkDpAnSB4vi4B5LNvzmkpzDBMZ92VI2sHaynLQudW/DgXpPkyy
Jg+K5X9E2i7OJGbX/iH87PFovn2GU4lrwudwQJTKRsMTB78Pg+XXFe6+ELk/
izX6cyza+5+jK39haa8Ce7doQundsS5NEJFONJGqrN9AN2xSDbWPYr1Alihl
NPaQ6XRFjLomm3O0kzWQhJY0PRClry0Cf8iJ+X/INdKBTiqG93ArGjiJe50J
8OBH+RiqxtRaad0SEg2vB35Q2leOAho5cc8/gHq/o+Rsjb2if3rVfPrnJhUs
+ZLOYGWm8i7lzBO8TNDIjKlVrKE8PyrSn5Fs78cHu3mKlZ1tQJHjEwqU8Rk7
tLpLuF3nedv6feOBCPaDjemkV1hhZyALwFE/Gy1Ry8iB35Ily4Edgq/f6iQ6
H6OuQMX0gpnXq5ojqLMDSQGd8xXJxfu5PNEE3OaqcsHLgfMEmy6Lk2/rpb7S
4Btvjv63U/0z5Lzwu2San+3DxCas9frK56fc2bGR1h/NaZvKv0+mWk2/XezF
b7vdUujXANybKcJ7bMbxRd0JZh3F3zqmMhN7BKVYNfICKrRk4EYIQuZyyG+G
oOTK4kcJj3atdczaRXRaNPO9ZjaaOM5ES3Qy4e38EgkRw0wJDorqW927bhHu
qx0TN7omRIZo5gDHP9STF1Zoq6eNdAKKSwKbOD9XODN2LyLYhegGS8gARj5D
zYqRJfLKKYGmbBa7VoF1CBugpux5D1GwpUgFGxRp016ApcDvxQFsJwR248Jp
qyXEEjtOqixYMNraeHm6VZJB47s/+VN9xaBU4vulZfMYrrXMJMczATme86eE
46XA495szZz63gIrW9j6UOj+6qwz6boy+fpPiatC4Ce5NSNEjh2N5QKNeLcN
9EsppPjVbW1SCCyld29Lcxm6IYQoP+uFICRv0drDeBsRCupJlAjodki9I6aM
GnJBoIwamSaldLfU+kg++2x4AfLNHv/PaGFwsYYTH3IrFN4AazABiX5lIDQP
K8XyjFr/I+KDEJuDyqljf3QBoTZvwW+ml6ralx9OVY4e6kYqKxuoio5qc14O
z3dntsKXE692KBoJP0pZGCIgGLI/FyEfq44F5kZetuXmPghWk5vuE5Gv0egQ
WnejBaTSOS40Fz5jkgy2ykQGOrquevP9m2kO4b1Y9U+mvjxzcfDQMt2XF/kM
GtOL/vWm1d016bVsbVFWXQhrp5i07GADNbxmm+bGWBUNMj0UqsFHfz4KWV+2
KkCrVl4l3qJI0nDHgEK5zvP5+quoUm5hPz94WSGBR+YRL7MsDduFvoieltll
mr9VgbLp1UWAtYPpq08cO5IqhhntoLvfDqmkyvD+xI9IXYkm9m7DqOHCNgKj
xQ82pRxqBwIQH9l1eRUWjge/HmJZqKc+kEw7E3LL9ZUz6OeIKdiOMdU0+L00
jKSRJs7WJ5RQ7KCJhsh4Nw4PKtPpmhjTDY4swbtl7N5DooRt0Qazt8C6v69r
KMFb5sI6xeRTJTCePDoOTV7fDPH75nbewJbQSX+FvAQjvdFK4NYmvsY99yBq
RzwiV1zCpC9kvudOqHAxu5d7jQkMrfy5ZpTmRqF3JQ6QPpzkj5d7KzYtyQlk
3RwKhfo3kDhyrkoBcKe3c4S93sUqG/VnXCZkA44kfrQFQz9pQfn83xzw3uEx
+6Cy987lWDnOBszumvyuCucN9v/A86BdFjrEgPX8U+u8V7iF+nhpawdnX240
5A2g6Cwty3ncwPmetF1wKCwxiX9gVMp3Wcqa35se2s4U/gktukznfPDg0+19
SChvaBytIZeVMmnvNy0R2yKT44IjmEfk04OdwYjuu3qhiSTqzIuS430dAiSk
GJTDTyZAZ5ZDDQZNIa74ZAMBtcjddGOariICDhEfInr+p2BbJrQyXIetD01Z
obyD8GtPiTMo0lcmMQ2U9arvVbWwJOwXiMrSHuxibVNNAhk1Gg7PwZo3/N3D
KI2EB6yRWHGInqDwKm5ibiDsgFLQXm86p5JMMHfxHwlGTgC3Z2W8CBQqDBzh
PSE5PeiruypmDAJ5jmLQ8OdrAX+ve5M6rsedJGuhu7Ed40/8T+/0FvMvjiwi
lZabpPYFT9xQfa1J/YJUFCWiq2vCebDZdkt7jh1DbWiSZt1qkdeb57XZ20AT
UEEz9HOLAgt7zARbyFn1f+nOxdwBdRWrQxTm5f1kzgkfdB2dOmcjoLxYGVk0
GVHCWQtZn9eEZD26HGRgbUDrHIWQ0zsSVBGZGa5eWftkxN/yeCl/CwvQzTYq
T8Tdl6smc/5gNRKcl8P1aDO+IsE9hLE/Eq3hffsPG3q//f++IbFHCdL1aXnn
ASzUYX6PzplVAmSbyQ8OECE4mnkCrHtSKF7zo/nbf23/trSQz5y6wQhDbkVs
ITOXuRhLJNbD3WC8rZVuM/s6d053YSpx8M2ar7goHbYzHwJDVavhMr0AqkeS
Ue0ryiJj6c126yOzahnPTHA14hbaK1otMjVfRMiqHKv9bLsieL7hDC68swG/
Dxj6UsQ8JdpB69xqERLRucNZnO2RNfxpPU2prwlwxbp4cmkTfqA0OPwD+IQP
1n+1PNU0HKDsLhysJCCPvD2DOV2CkcEtMPQhfpI476+Uoe0WsE7JSgMOVGfj
jZ4gEEHkcNst/cVwQb4P6/ZFSGHTIxxgLzI/+qZBumHdm701GaO3+GWsB1ZH
jQYJtR/1OAsYloykscxUw2wgzHXLv9sWiFeip+pzbMCHonbHHA5O9NCZTp4j
7bo0Z8rqok9gowald0AEef0uBs6y9Nf63OUKSwrfLZe+CVArlabYhzWSRzNQ
3ttJl6+Qh4RECaMVPjpMY+ZBjaubNbjw/mc02mrlc+HRb6miRjxat9rrlc6u
uygJ5XnEj20BKAXmhrVNeK3BbcXlnWmT10/vwuxGqVlgqlB2qlHIZj6QIcEZ
196l4YBdV0rOncE4kmWIsL8QGMOj0wRdpyzjzMttqw+Ogp7LyYV+5aUDJr0J
Uy56Tnm3pfDx96SEseN3Kh5b+jku2ICadeYT+yHyK1He0RjdRTPt2KHEdeun
okWVu9YoG+aANSmPCgrBW6Nyag5NOcBqbvmriu5jNeSlGWorRvw1C/r7GEXe
7ggYT3rcZFYXOWg+bFJQVniAJSem1862LjMEbRGpRZ6xxNi6dVFn+I3jEw8T
b0t0TeedPADzyN9OlDaTeNsfs2DJty+hYsJ8b/vAHTYLipf22RubsgUOWy3w
4QTZevIn80t3iUdkok0VFf2myc2EmrL/rLV6i86Ucq4fa3SoM7gf/hDjPGZk
6or50eJzKJAtygWOi4TMbQ1AcsuKl0nVMmR9b+Pzoak51p4OwH4lkMNumTgk
ffBzrA46+gj1ZwQTEe1yNQc33aeYvOw4fmieN+oms3axXnrebNgIeYfybvXa
LnSMEXv6rI1AknWmh0Nv1og1synkYl6VITP3fjTq1it/WuzOQ90l9RTWBEoA
iomVi4Qoz3UcOHQH4YiVSR8S5vMSAtYfM0W3HR3xkjh43Y493msZw3uDmgFq
PiS0yV6ULDMKPUDsWU17U3CuktigDKvzj/DgRwmkFVmjtjKXvPEcVK4XVzKb
NX15Tr32kdq6JOEUT02PoRb/PDOUMU1UKTiEgfo4mb1DLO5yuXbPZeztZUVM
A1neRmXtm56mQnQ37IR3BJaJJG9Y2nm7SgzEoW4G/gCwqtPK04JMot9aTxUN
GyNj/bseZVQPzhuMtCvdJ/S2bC2bVFN9FnKpApwRg88owq3Du6f2x88nZzVZ
02bc2TtnK8LmKXuRgWvtOwIjeG5qTMhyGUkKk41hCwYyMHyXUFCcOISH3Qer
pnC1CnAPOkmBqxhEh+HX4h5O+bE4YR7fVfCenokMtChiC01GXDKv4HXVJIN7
r9OJgIIS43hCMdAPA1WLmKAy6Shhg/M7Ei+FTDCN0K1223xkW7AbOAfNCEKb
CTG6441g59z4jW9AdI5XiadKxy1e5ceIoPi8203lsQ5zSK8Zoonw97+V0/Nw
wJwYG3PIiKhh+aFNn/SCTt13V/7BIDoiJPh+4FrW+KmEMJTxPiZblaoNWXVD
2Uq/1L+fTFLW/kXihW+7ZP1nLYpHGmdHAixfrXXMW3lIWt+vyj49vK+r/j7e
GERaCXKyKIPD1cY5FBxdyMlzOlXsp8YsTs1v7bUfOE8MsNQCE5mRm2bLXPBp
Tb8gvF7RPgf/PSBgq2eYPMCKtJccntRphdbFr4NxjZp1RU3pk909Cn+aKAua
ikB3/58Wbx0M1cyfKo2J57ixcfXIP+RgUllCPXbn+0wxTCnDEs3gW2I3Jlhm
bUOw5qCG0aFXlE8CFO6CIFuyQIAOroPurv2hyfTN1a+1bJ7n4hCg23gmXt3G
daodFcRD2K6y9Oawelk7iwGchDT6OwaxXTlwkkkhAYDXUUQSEjmULVBYqHwX
6Nl0wqbAhIHqSS4OCHEVcbT9zJEXwkzXfyB3CgYc1XirY5u4eLuIHGoT4NJo
T3wnhFnt9Kaxtqp4ogAyR4EZ5BZVmTpwAx27Wr77roGtVJsPRB/xOvmvtXb9
WbQv74bpIMbl70FxkO5vmVmH6LGbCkVYiUZgmUIUEk0N8Mja99OM6FA8Jiu0
mRiKL4MVejEtt/yEQ4y1i5UKRqAclcpvl9IAlV/SK5KsQly7iWmdV9SoVNcd
YEGQV5AXf4Ryk1LFdWQhusOlJwoeazmRRxvDaBq2TzO3h0tqWxi1uWMyBXiC
OdBHied6ipHYQK1OgGB7ZFuBjS2ogPC3YOTtn0u3htyxWETlBgVvFfq81tKH
Ngxf8Xn08e4bCwxgmFr17LnNVIZl4XhFsLMwdYwOoPj3Z1g5iex2Hd5dTsz0
EZtE5h8lfJRQDYhKN6aZcBFCY93DujheMR3eMtVOQUDxCWtXo0iv3rFEk5BO
qhd9aJJ6nn7/kG82otGoQZU8skGyppwHxZ2W0EOIGqve8AMaZQu+6IEwJsHa
KkRqI1l1RyqDuBhOEdM0EMLwKKQBtWz0eq8Gtrp9ki/ofdQjje7wIBMkHZlU
unZE/kRGb/7IJe8xrAB35yKnoVQtneSw081iCraNbnVjLkMwVf764N+OJMzh
q9xFfQBNjhI5BnEcjg8TJLDMKgBLgdBKD2B5H78Q0lE8UJzCvtokABP7/1lx
JnZjw3kIttHwGf3uryyeOVipQGRM70u71xknHjOIyK6JhFjpebrg22qkIDKl
JtikqEuwpz3KvKuKs6OjXYaYgv9VmkodvUuxPdEEw+mhGYVjicEjYuodAOtZ
13JI3JNesxFhd/kBEtKfJuaY5zLzzaLU8AhsHSpoBJ2gMSYcvl3236DtUGFr
3AAlbpjBpxWTdgVJq6zxmnT5FDmj95g30rKzQyKfPoObi7i0JfKopEYxgWVG
TpZ5LyMjehJKG+zXQuXrAxEuGaA2zm6NJySP130qzaLFTWXcF6L5kSwCWEI2
phRVsY7l1dsw9UAkI4mfKFTJojr316tHx7rY1dAETfSGZ9xRTbn/qWimMYZR
Q9K4R+uXM8x/T+yxXabu6Kg3q0ztM/DDMiB9trvboCpqF8HF/3ZRtdKq91WX
NU07NI+y1TRv0xRm4xQNOGeeJWeRUvT8/wVxGOTxpQm8+5tPtwXPDcmeVFBn
kHcP2lJrZ8T8Tn8PpIXiYPs5ghWNBP222J/3fIzSZvM8NQbBBWC0raJCUFII
aBQdUAJYGiiPu70ci806P4hC9xQWOk6WrHNZCLtmv8cWc/1nXWdbRkfM6lzk
7vr8mwIG4VfVSob2tjqoXfBg4Fo5ubI1dwgtrI6K1fjo+VnCSfs9VN64Qhqy
q6xEKorqzwghP+B/sYYmVv6j7q3rX4NZZSG3Y5aSe0mmWNpPV6NV9SpAlbHI
0PBXHL02vDb+ETOVOpdz9Ate7h/aAYwmCRC6jvOJV+lj8UXl4Efzrc1vJr6U
N8U71Y9aj1U4zsAyFFhBJJMyXfpA6lz5ceP/onqrqlGMk7ZhjWerFVIrbmgu
3yGDJsJDJ6oBKXLrZarPnI9NQzjj8MiaaJ/8VZGGT+vU/zs32fV4735w6Fvw
cOoONQmRXeXIad7m5jwWT+PFzBzeFFcb57ZSnk3RgYnIJWGaB5Snzyz3dVYf
B7LxlBly+Zum3/kCnsrn3IuEH9UnVFzysp5SI5/uIpOLQRJl8wHWNJkxlNoA
vB46raGfZ8moW7o0IEH+Cb9TfcehrlSMsNx8U+if5/MiIuLexuvJoPhzDFeq
pMODt/63eWj+tZIiwmFmwi1llann2Ip7RuhNQfyxGtw05/QfK/h0qXsrpQ/s
LtpJWZfhPrL1SoT2yQhRnYFQCAXdvDDIIo4t1Mhbfp1gen2rw0Yn7ddvGQ4l
rDf+nPOBNgqQGFr/fjAJON/sDW7tt7zdNMzG3d+w6n2ZM1q9QpYIr2tmmYIN
W5jyPBIx9d4J8rnfMFvF7Mpu84ay0HD17ntNYfu3mQBsYrqUuU+HdNuPlRoT
XM2c+SWl8288BM45goSvm2yNF+Nd5Z7UBsitycICoB2S8gX7Yn7Ozoxn2d5h
/su2c5IVjxAN271f/27dgM76qTvd2VOyGc5E6lKe/8k9BTfsUuMMrP8oKDgq
sHHJw7eCk3T284LvoynaOnfo6Qr2/O8bxUO8Zj/CM4OvG2R5xWKC/ssD+Fse
yUI5FzjQ4Dl9FoiHouxbE+rzkhkFqyZGSyBJuldBBibVXV/dLWnklrxcJkaX
9w3YAwxyvrpo3qlLdaRrPXl17PgU16c016EnmShyjXOzrn5sQ6tParWRPN1P
NZwJqmZNfmt+67nHkTAPZPwdUM1dhwZSTbw2pDhr1Wwq9Gq3fNW5bLL+Pd9F
t+XzXBGAkjEMx5xCoaKdmRt2+RsQuTAvtkXdxGMuJEdh5F8ET0d5qJh354fI
7nuMLUniA43qj64W/9q+0maZ4+LaH0JkTRXefqD0e93p8mDf0Y6Q4eJRUF5t
8uOzrcTA2Q8R0rYoZ5+tfOAmdtoHIT0rTVYdJLJGqxtfeb+qrx2/dOOkgCC6
jBmcs93T4IYp1f1qdFnN3jRp8aAzFo2Q29XCqU89/dpTtuN200toJREYY0TN
x/HrEY8vhHmnjpkY41Bec9N9ukjzAFE1P+FMBp1onuSEhDLF1oQzE/5P1u8j
IRMjSyMStwUic1hBJYXU/8VdSDTzdF4bhxK6BlfMaCpxWnOzWIwl/hoTDd8H
pO8LurLVzBSvW1nSc+A9zFDc1h+AUuLdesrA7SBqc+OITrLRQIPpBW9F96rG
Be1NnE2dmvOeqJvmFp396Hg6WOeQ6RMXK9gIOH6Zc4YxE6/C8YYURULGigtQ
PbAUSk//Ej2OptSmAVCM6ZoddhCi3PCPLpYIxEra49O7OBX58ayF3cB2SHqg
nPrKgCiHFFyBZCJgwL9kPNE43ptIgpnEtRPf0uBrafAN3hoX4W6kQuKSa7p7
FqWQvL2BeYF7LV45nheBlmjX3wKm3lf4xvWzX2v0ryFCsbGcERFiuzQxC7FO
hY/bu5O7rMOH6N+NLs1090r78unF9p2YSIndJmUjneyWyGMq0ZX+HoUseaQG
hykxHqq6kVGQN6yHMn9Yt7NECB1lfz5o1P+BZJ8wNl4xFEsct3RIpSyOZUNh
wW8+cCg4y4iPhv/ONxp0Rf+0bnpuVlWllWX6i1gXZx1ob2X2I50sER4FVZCq
IBIukcWmm2KrG7svHMWrotUk4CviVjFPcUt3fg92XZDLVtDY5HN7uKTYpCYB
yI2V8a4PnPRgBwao0QO+8h3q3UxZeRlSdqlqTofaIT69Azi+njDkHovJY0P3
Uj/XlPsoEfJ4nb1yZJUjJ3X6ttqHXZ1mexpsilhtsCusCODBgrx3FPeCY9s9
Vp9RfGRXTcf/Sq2+hfPRx3av6CydqU+pHiI697p5pKLbaSlc45va3wGmmBLc
lS7RIj7plLyUZryZVtUgcgu4SwyezlZXOzQuJhar/VbEiiRW42vai9FPyqb5
yVY7e7t+2IAOsC4CvEdSNkGM4aKKzOvcQvIXJxFGRGJk9PiUw99NM9BQdaKG
SkYQKKgIPyg7InMWHzVf9V3WsZkTceuELGFB30qzU16vlu+bFDKRWNkzWksV
tbxytSxHQcK3vUCz56DfY0zRYW96iCMV8uZo7F61VX7xx48f0EqEK/xIexvR
QOI7jX+lLW2Pc/5mmmlCR5qkTKCJEj4sPpzLJuFJOHjv4NY2XHVDsvyfS7aP
8f9vz5zl+00BSh8UeyejrbFMsQyBnyPbEqCcmI/TX73Z4lKZ3Ce7AE8fPq8x
X8EPRn4IyxOM/mUCYxH1SNS1LreMtzoHAEDBM20Lqcq6n/I+1DoI48k1ZUgG
T4NL0QCc+OrYT1zfQ5APn5+KTRbbdY5oJuqpRlIsSOPz+6LnSSv7tZbNUlL5
zSrtUjcrNuRyBgkb4wRvcEyQbd7bAevHf1CmkJcT6CGL04SDtlqi7N/4rOq4
oppuRzoAfdReaKx7yNqk20v7lDNXFSvu/oCIco8qmo8LU0pBabHztFAzH1PI
KYmXmbVEIbDftgAFm0CkWZbPlmsshBZc0J+R+06Jj2IHdz7INLz/goLUHQrB
LhXQGY41GMuWe4Keza3Cc9rWiQ6/ouprtmEkFHK/jbkCWxbcmbA51tpEhEeA
YOSWtAzB7AzmElGslmv4WHHS8o+j6uJNLsOVvz4wX2htHHlm3KVA3maBrAxh
zrt+T1/J4AJKI5STaYzEN3uJzCA7vNdIGtvFraRNc4mpPK9FjKTCShLGRI3A
+0YgJ+kN+B+m2zNtiBSds7hHOR7ySCrW9+0uWRIjVb4DlqtRyqxZRPZGWqCa
3/EjkDfi2THbnRzLtqdxhE3C89se1qKmX7Jn2BkSFyadpz9fmy7HfToS3E5H
3UB4wZBAGGNM7d2YDRQxbQCcGFyY7fUTuSWHatilPV+tCqmIYVfJqTnf5pVr
XKG8/CwjO4H24UbCutWlIBZk0ynhRnM5iX0+03srzwcDPSaezZikfycqOXWy
nn01Epq61F7YQNJ1/7e/l+glL+IyOZoh688eOH/+gKZYl+ES2gsvvHMWwXtT
xEf3cay78g/eywBDYCf4U7hxc17Dg0GDA/oBnBaZMECPbNvJjN2V5IHfx53W
OZvnYmUL95kPjeMFPECq7vMopgxt2qvgeqx1vAug56WszOGN/nhmoutq5l5z
d5pNMwVX/N925f8bO9OOp6MPQO1xqTl4kTfhm34ByB5gfpf419MnL90qwITn
7H/1ldJGZOn2KpWmxo1hV1HtoTyM5nnmVHPMxs/nya5yLS5mhW80+UqjT7MN
oKq1Wlas5Rb4eZUBOChQw2/Ny3qoX4OMc7noigKQVoTPQzwkbOUp24ErwnTK
JHHZjT9e124qFHOQdQDpja1iPMM5YGXSwpk0/uMyOCW68pbD4VChCTXOMEdM
sXl19vpVxY7g1PA+YOk4lFz8rJd8JAV3mKaP+IwD0E/oaFIwovtCWAfDoAHJ
pq6Uu/hs1ePQ8ZIrYflOJR5xB3S6JfAcgRkT94+8+81lpD+KYGYOv8gJsFGi
yEr++/112Khhe30YKdgsXo9m7wwq04/BcfhaP0MxcKdmlX90LQXimAw1kEUS
WwPZyyV0HDRhjdPry3SySJABkfJjTIoiVB2/SJPKPjYDINmGD54ExJ6SWhbD
vTFlzo/KPVs56H3TmhKj2xrljd/WSgCcu4qmR0bGrk3xD8soBwqu8FmZ+IoN
2KpXnURJLwOFipcebcpZn2iP86KCFyigeQEvbuAeCybY7Ggzgsy9UEF0CAe8
vpTNfAHO4UGW9cQRQqE1LY7kYtxnDU/XhYegKm0exTiwPHgv8Cw+jyXIKmv9
WwClTHFRGRcxEKRFCwpCzmcde2p1XLhWU584DaRicPoc79eNSO53n5Y9EZDk
RqLoKD1M5LVW0Hyg3lwqV7X2+VlToI8fUTFpWkOqO1iD02pb5Ro1Y2oKgBfx
TZVmDNHZyzHTro2s0LnvjwKePR+5r5HjlzkhjCH7hb71brSwTEAET6TWyHK2
Rt9AZJMOMjGjaLWID/ooG1mAhQfx8nrfvFjpO2sfFr0Qn4uRbPcB1rH/F4bd
16JA8MYvRENHzRyX4MphYhaBwgGPkli918wtA9DelUyOrXfnGNSypovjCgkl
/PECFFsl51z7jHZfDv0acGE58OMeLzfu9k2XiZK7uNYKVBJ77YVTslO52kJs
d903CBnrE3KSVfIPjB+hb4PXmOYIvTnyH8nq6/Tf7wBELzODcp4VyQORyky4
BmQNNetXhpxbOGRc71yb7J+XA3OlAovh/ka0wJJQyUgwJBiAMErXtP+AhXwI
g30R33RzuiZ49yMioiYSG8bDBXz0tDjBFvLmJid/WI1Dr8jWkHMrxdMeooca
6nxk0b8SHx/RdR+buMYy3fBIzh/HlLuaB+1ANfiJlLHEbPSqDTOLoSCzZ5AH
e7RyHS2YdzhRbHs9/5iCFKNFxegG2gISkI5PZVdvuDL376AI35wZ3xBvLktv
dRwZVpwrn4jP6k6TR7APXdbe7TvZRlj4Nm7fHGnUJOa46/Igv+SKP0R1YZTP
c4yFExZbWTU9x5d/R1/II+/VhCa+JSfgHU89g9QjSVu0RMvxwunsUrvCLQRg
fH/WAq5tlaggFUI1tGZwrjIDOHFew2QmghceidQsed0kuS2oFZ4OHrXBdGRN
C0RGLEj4hiQXsU673TKI1y2/0upqb+MVwCXuoiVwOnGDzo0Z6DfcLFTZnBBz
bDwRwTF4TnpuW5o3mXiOaORCY6R+kiDXP3cKnYTy0CVWcke1oXLaxrc806dR
YWYAoHQ61GEV8OGTTofE5J+XSwo1W1zg4G9Cw7KVgqMZ8APdJmZMyv2ERQnM
FdVf+q+2JFpxEJ7n+ReLi0OaX5Qjtqpwphg7OElq7gQxS27akJPm7qvBUWc1
MnDAg5bSiC9Po3ijIlZlL5+Bt7FpiqzH+SaYJ5YC18FCQ149cKHllhgpTuBe
cZiAbgsB7HCweUhUTkgyERIcfjL85Q262B/fvi3ucr1OnK/j/h/lZBiT6i/F
3n31Qk217VY2IDWfqKNPVz/0ndnr+XoDpsve2ZE8ocJ7eoOEOhV5QoPYOLHP
0If3Q67QUAVzhrt3bfWZcpr1Faj0yYWhJ/lSqKF142KMikbw9IYZUDbL/HdT
PJDj7u0FXVgYYGBxI6gInhagmhbXTcvwrQPRvqHfyPJbVtDPS4ztuhIrtGNd
B/yKnu6VK3XuuBkkNQPwsubp4a86zChgEXMMrfnTRl2/9sU+CQC2qJJij+rm
AowLzBxcBGOuzBXorfVqzztMzAO8cIOvOuw88eZTaxoDB9nQ7H9kFP99Kihg
qVokn++VOoYXQ8oJkpoh4RSh3GtP+Sm1pVZ2b3E8XA2PIVcRlbElgbdiZsOm
D0XMERoNx1+ncsK4ARDvpoJWJyGvBJyWYWYIJ97rxeyCZJbSF5QasE23u58m
rEMnGInoriQUNEU58ca5JhOpEnwUl93pMH3V/zyjlJu1pF5f1myb505HecW+
SLnoCasy6OSKLhIS1OSeEQ5wmrLwltbxEDps7fDRgF6hyrSnwOIO1iPqDPB0
ARcc9vcQp7wOoBnYUhA8Gcks9DBTr1saKH/sKsjHAl4OzsIOEA/DLr+tHeqK
cU8fG6hqo4OEzMCwWeI+87GJKwJprN5sHLe9K/FMbizkX84cwzW57Biv8ys5
ezWNhdMVKplYmXz43ug7zw3WcvV3xkVGEDNo4dDJSE1ahuav27hfxfYfUo8v
FBtFcdHtjqvW9i2t1GzC0G/HUu88dOypYe4Ffqz7JB5U/smOojFyAEN0KsLI
QmvWPevoaLNb4Zgl5rEHYxsL5xIlAkyVgHQEqr4g7K//a3bT6IfYgcTfbxzM
zQWtiYbTn7UqBm8kVubAixoDtE6XNxqqVv78stqZ1X8Re4s65+uSrFjcTTnd
Gc5fqSJVd5Snx1vqOKDkLr80nt+P+GZVc8BOdLvfaVtarW0w9OP/8WQqyjD3
1eeBj3tEVBSLqvpjwMEtMTgol/8esOqolXd+15SaoLeMO1SDn02OOZxyWB4s
znNCVAdSCgdbEz/xtY3GjmXT72N9UNM36vJYN6TMT5+zvUBWygdfMUFR2bNE
8oMtKMjzYPJDtlGhhScNMQewjI5N+ofCdtdXJRLow90kLeoCOC9xlWevpE22
k746L5xx0tvi/feeSKfcL9iaKB4fsDrE09ofi4l3hExgNUgUsaO4PeuVPiWc
Hielpj3ysjOvt5NxRpE/KqT4DIk/5FsOPx8ecqJV4hJ3tsL4RUIZ2TCoEdW6
LrCAgEOkSamnRzjuKYJvueVQKbRmFmUd/j2qz1+xKVsLrxlPo0ejpW/+QndN
7/OF0dwOCj61vc5do5v7QdpsMBXNvsKMV7+6Fy4yXt3P1z5xO9+T+YTpQRAh
EAsG/in86BLod9Y63tcfCZyjclEvASP2Y9PAjjN7MQSaNWj9oDSTQXzfT30Q
rKZOuRAY8XXVUt5TNb52ieXvbSx0uQd2nyX8o/W2Q0lBbnvhwWIy33qOjRiJ
bpN5YVvnvMoqEDfOJYf6Sr9AOVLhdEzKMJ/XylrY0ul3f1TpmVXLJkhztiHV
fte2pLpS8qnHt/ZVx/Rex6zHMzF6OuV4jeGoul/kls2RWwZrw3QNMhdH0Kwq
WJom1Ja3Vrw8bCCQAWw9vZgmzU2To3G5FXxJjeEQloAxenq6S/vwVCcp15Oy
ckdFwfyJI6mchpgt/mPraJnXHxoMO65oaiP9lQvV52FTb1HMV99Sux0s75Ne
dsgqFqTmRAB5Rh0najS0xUA8V1IoPxY9C9ZZxfq5ksDv4yNUyYgVSuuSB0tR
7+rl9OomPXDJODZQZufmDqkFdf7GONWFsMymAYUvUl2aM9ewd6QMtoJesfD9
Zve17kId08wpdVohrEtj+UyO0zRcXk9ddsVQ384584ENtmmE7LDZYnczhFGs
iPSrP8Ux0D9gEbUSzuBqmqBJz9D3ZO/6b70abglDtrkmc/bE285A+mbp5ZW5
pXGfl1X9l+F2SyonjnjTTrgYRJkYqLUx8rFokZoMfVY2VSSrOl23jSvRnRig
j1j8/v0oUeUGCR9SazOZK4WS5PntARqeAjTok8VJK+y1y1KLIDUgEKkLX1Jw
PUekMFbbCOf6XkH+OaaCe4luTJZxzVSItITrVDvyQDr8O/EAm0bzQyGl9awc
Ivbhcr5F+oYnIJXAFX2ABEj+tzSVDUcyIe6w4DP0wB6Mdba9f0dxeAzTgUBo
EXF0mM5i8vxlOyCdCDlf4c7B+FBLlSEz4is6MQaccMGntGdl/ktdyq5h9qkO
H4JdKsO97GNHJ6eRl4LxIM9U4a+zRp1wyYr1tLqmqLUUalWnwcpFu6MkhaPQ
hFxAknC5Whm9o4A1CDdz9FITeUEGkotZGp5CpHcjyWrSgbyRpAP3iPQCSuw+
shtgTUZYFt1dYBRy31as+HAHvutfXdlCYJcN+bvGlylp61DJ/eu2pMO7Qa8G
H1jzEFF7D/JXP/xjxK7FUNlsiUjVggfVWQ6T9HY82AeQg6NOVLhExLjDoqep
UyIS3n/OFO9qME28lnwA3SyE6TxKF83ckNcfzY0HAqlAyLJmh6UoBY4juqvt
JoX2PLmocHzKbX9Pkc6ZURzS8IBgUNQ3Qrtjjw+xC7LRJj86GZN0PDaRyL03
S9d/gdFdX7VhTu3DBPRgAkeTHp2j1J0qsUDJmQMxk8/zAJFtENJU4kUOvrlO
wKLN+ErEuC6vAFZxdSy3H6avUnPbEGc2x+51K0+naz55VLhTTn5qLow2pjHw
iCF5H5oTM/t2yi1uAy00LVrL3rwonxEP0AJY8iePKIPcVXFE/2O11YUT1W3G
ETY4s1w3vv8QbB3TwuiDF/B/42+lQfVpOf83TUnE8fOH6tnkUIGsP6z0mu+m
m5O702+9qThpdXFkYhjzQ4Jv8UdErJ775yzV1Kp+48ecLz7gra1f9hF7h6T5
Bt6XcMesNgerIIq9iOhdej4PgO2TI+wnVVgQgHzk8UYBjpWp6zvJmIS7Bfl1
D/vCODHJR0IyuskqXYnPN0ory9hxwVL5gWwYqYuHurmg4PA+UC6irUc3ve68
1uIHkZm8bdzCpYr+5tqSaCIAVNv/y86TGF1+94fwGYUx5/uUS0FUi22XUTB7
EFTF8EKU+v3zdvN35MJHI6yuopcoxBIOBHJj0agAEF7V2TZPzPB5N93ykE11
NAFzrwzU5oj8MvWHK+j+zrxRJofxFLjSzsVlHxc9PazZZsHqeM8qw1HR2ivl
sdtPyVS7H+xDOxlAwWMIJDRl0bb7oMMHLI0SAfOhQRhCV5WjBFSZE+qjBlZs
U0Mhk3l36swypWGzzkES7LHMVMNJV4T/yaWVlT6qHSoy6nPo/6JqWdzlj7mw
YclJZvWVHBmBlJFY242NyC6XK4YlnbsLM58pxB8YhiZ0MvcFRmIcg3eA2gB0
a3Up0m+o0EA57yFACvsnJb07LpcxvD3RRdyJSoVZg7wHRNeQwU1OjPhXO19V
OtQ1kdIUIS4aO4u8fHsnqpLKL48By6y6Vbf6pUrBQN3WwYyJW4FFZ6sZXt8M
7ot9V0VLfoHkOQ0LF+aIWj5/bO7o7h7eIPUO+EcnX5W3Bb8i8UknPn99zs4P
riweGVQS3U8aidn6A2/hSX1spLHjQLjL0QdaQOHKTZ21zDXLwTmxSEqngpYL
m2rzVLMgs08l/5mlTRtJ4CiTCPtJsr0uWwS3CPp3w2RK32r3UYPH1krVPqWm
QD41HTURoWDsoMe59OUilXG4ext3hUK/PqOxvyDKX3ChPWnONCjpzbgSouqA
WGA1f7PdmRoIpWLaDWG9UsjvuxCYczyon6QQS4iPpOClGuOIl76WvoEn/uSf
RpPVILNK83nwK+ZUd/CwJe77CrHqzlCuyVCIgjfjgKdl0+NzE5ViyWEMFs3M
FiCIlJ3j5Nl8Erom5VZ7IFKHgtKopdUrrAC6pu2whSlhJeA3HydMfeeopnKm
KrdOOn+5lNDe5r5DocmE2TVDInLlT4TRJdavHSiTPeB/EEB7Qpqe2wot4Q5R
ybso1p1Y5CVlRVlgba+/lPQGJgFZR3fKmuJNTCwLdYknKBHTQCGVtpVT1DGO
G5WfrppkXcyb38H3uXM0Toipz88tm/BJEvGx2Y8Pkid/cmyjb6apRHw/HKzb
ox8baSF6E/U5ZmrE8VG+WbK0x0T08OBRRSCoEf17FcN1iSYUS9UZUqhJKn/i
xvv6Ts0RLOJtep8XxvsCEvGANVIUj9If1sXGdAbRayaUTWbForYcwXNKSGJX
WHMWpoGjl2wNc2ky31RfIhJ8/cRUZmOgq0/CRv7mk05rX/WNJ7KPHcV0V+tv
eKyX8JFcPmXnKf2AR5Nurr+U5d+35vvIBl6pTWIdczkQM7yH6XKnMRglY0iK
Rva8WC2XbmrEr1rL8D3WH6f9tM6k4skPrPZbPLtncfoxAFqiMPXFiny7SXRo
hSqrpCisdNcCkWxVV5KH3pqPZX7hQf2LmD/2JA3SPeUmgAYGHYlsXpHADChg
5aXoa3AhDbE/7WQO4XC7d4hXX520DNwndfMUxGeeda0pMcFKn8l8sKMaW3M0
BfhPqE+/d0MkD1Od5OdvC1y1bZOZgOTTaJo/4NxiTAAEySu5q78cZksIKcz2
SHGJCqwapvZ9/AQ6+b7GzYwPVbgWYfdcr6RgUK0vHCb3uE2/TD+M6ZCyi8C5
+jZab0FW4kwDRyRkr8Vn0WdIZwgCOJuu8Rqh53T60ob33ivpck0OyCnbewm0
i00UhPx/ejcPvFCQKccucPfAcsQRljkRkBJLL5PbkfuhWcCvVpb9H+FISMcf
kh2Nk9vaUfduaN39Qav1hxaJe7jolCwe9JpYt3vGkP9JbUKWZsumciovriMN
BHVqVKAuKdKyVaHFmx/2PR7fQHGYFEyHrAoAXbGjgmjX8jc6YyXJtAm/ITHW
1X2uBzUlN+UodqXHLgQsQbb47K1b4ihn+dkbJEU9qJjjnyIsszihUPyBoT6K
A2s+JWwsvVbBypjLwGcF/nLHjPyn/toJXCKzHJWBPlaEX/c+zdLah/iMOubT
2ZxvzfvOQ6LP4l6OqCpfEXqIEnpwNilOS8e7pyxu3B9g6uX549wpwLOTxUtp
lk6Sa/PHGwq7NJKIzpNmczZPZ7lnz9rupIyj37ZE/P8R2hOpBXkNutwWeP1A
t0aEOMcw9bwF8ZlIF8DIZrw9whJ5raLoe/JdtH43WA1RABTY8DJmeReWvyAA
nxmOYAIBVB8d+euqBZj+mUhO8NilS8HgoaLk12Acr/bq6aJ4KvTDqUKG9Exw
gm1XcPeeJkZNo5fpz7Q/CcLKxUz3QMiWAyTGMNTEw8yq76tmfUKQa5aFs0t9
V9gO6RwxC+0FNYfsELYM0QMVBcAsF4338eQLnvYZZS0VVLWop4avsr7Py4gH
lXQjmsw4zatqtVkOlsFByIcK/DxzgKuAjPSw1bwJqQnYvmBCvIr71Cumkk3q
hD/ScLrT3IHwB8bR/Nqt3ta9ImxXyMGUQBuP8ZKjDGsXpT45VFdwQMPUUVMT
lft8ZVS4XHgDO4OTlsN1HYEuWeL4NLgZp46MVg5876DITYXCc4Gg89YhjBM8
X+ufeWsOcHaxmNIek3Ngk93th7c4Bi62Sr2oIRP8pfnoZaRY7pCqFkLca5mp
dIOpSarBsocROKXn5Wj0o8xxpN84usYpy+FJaKR3VyH5l29xW477B9hKsGwS
CxkFYPWjUc01ENRjAwf8nwfwxfV7STud/FdW5xzp29rvT0QuQ7JWVAhuM1l/
nSShCl0KwS5njsbW1RXhUfhgFAsfgdNbLyuFWK5eMLKX10+Oapx09tUBGvrO
LExyy+RDetQvUQnmpGEJSxA9jpwbW6bszuP0JrNip62+sC4Tw3rfza3w4rHx
IJeaT0RW2fa20Tj5KyDhNOjsc0i55KULIDjPRnck4JA+La7nOhIm8Ao6suM5
7Z3rsxMT3u6fZLsVkbtuxX+4sUQ9oD2IiW1SlH42ftK3f8SdwdSz4BZWLSRK
SE6WuVxQ488Q03yiSIjgGR720hR2beJTbeFTfx2fqUbvPklrlpk0Ufvt+DF1
EysyxGOtLgzT//xNDAYdIgWiK5D8JtqYrF9K+lzESGUppy1bwsGAj7VGcrqo
wwNz8TGunsVf42ZRh3CDhMhSp66ZKFvm7yOlToqdE4SxrUk9PoqrgIWKyC6f
/dgWPCo/+bjp4Y13Ta9D8otHrTppLV5yzvJeEPKFXnRMsV9Imp3+ib9ofSwm
On8ns9vbIiXRD50crob9qmbJuRn94xHoqnYkOJ1C3yCjvNz69wsMfTXirI3v
7VbA10Lktxxug/T8SffbEJhWaxTOinIvVzrmiIhxBPYfF6zkxK0dqJMjj857
2a14gYeNMlk432tGoqoUshFquJFlduMxpNQFw1cXeA2UkzlMiUjqF4f87S8f
LNL+NPogdkp11FAWPt/QazIS6S6OkR6i0V+x8VXYPCtbdQADK5TzdiZp/LNu
HW8ITxpcGyJCjv210QJlQiE7u3GbLvvHG1neAXgdOnKusof4W8nOXVt6XueB
BVs5K3zKa4WDi0DMjL25K0i9r+E1irtAjH31wNDhJLFYLQZR/AWKO3vzbi42
HtKnMj6iUTOtrtvuBMzL4GfgUrs7yra8oSAc6WfnDxa+2DLAaecOP9H44XkK
21e4Z381Z4vRTkR9Xc5HgWw/57kqTzgj3luSnK3d3nBSQr62o/lN0RY1/T5/
Pc1+Y0cuCh4SzrfT+DlPuN7eh7YG/wwNjd+Fn7xEsEIJpJi4dpu3co8ZPuPp
A71l+d7TYA21rZzeCVBgfaSneTAOkRuzJLsUn+1hLVAdE9asyBN6o2sjvLAZ
thov1iWfEGYYEfQjJVV037EcNxIxuoH45W6Hc34aVP+NciOdN+3SesvEmW9G
HtjwPiIT4LgXlXEMiX9LLoVWRsOvmCNaLMb1fRyCVjFAyiBDGplza6/KJIoc
84GBZYQXEMe+rr7bN7ZZ8A55vgBUvzyenFcQtCyLj14LxiUff6IR0XKdFhiP
yxgOxLG/UIEaFEbCOKMNgJaPbjtgKPcQd1tBYoyRFUSN5GI2Tp+IYgfnWYgG
vXyCjVrnIdVcwxzkN6Fsfstl892c7zMb4/HZDlhwqbWKZ0tgH9aNERlvp0k0
AUJIbvEBAZJEMvswj8XR/FadE6fNl3+xm9mP9/bUt0d19+/UEwXqDmrbQAhm
Rev2zu9FJOaZPVbYc5ce9wM0cCEGStj3q/906Ej112YkDG0x/AobgleFz79M
2OzSkwKghCjb0xg7QBXWPJ4J0LoTK7CzJ54u0SVYJQoyKao7gNGbwjqgONtb
FHa/U7oHvWZh6cgwmTmCoGwXXZbBr3FH7hb3kyCurYMS9H3r1jGpoF05Aiam
uJHJfNLodVGRruPkReC6Y0ZDlE1p/di16+o97S2GVhQqhqUAz8wCxp4fgurT
8vow7DdGZBV5e8iXVajrkDIG+GeJtx+gT1fmuucAgzRR0BzKdYEf8rJh4zRB
Yz8izhMy/oUrLgbPiWJsAVLauBbj9XnFwxH7uleYFOK9Eoko6LYE5ZcOFVpT
cMVdTPLFXxEcMg8R+eYrAvGbUQ0/ntig9I3lmmbN+8/WV5Gqe4h4OEOvnlYO
xgiixamRplJJbw42u1bSmZ8WiaLzgRVS3ku1yXNLoaa1VsXEdxzr9U4QrU7J
cRreKUdVLdbdzvemVH3uWEx48XsshviH5dBEIYc8bR5fzd+N3RNBmJVKaj5N
s/AbUJE6GAwQ8VpKrNVTlgN0oKoDqRBsyTxfHUVzGR/BtTinJ6nrHgTWMKk3
lZ5R0F4wzm8Lq5EnAz7rlTenxWlTCvhJco5Xb5Wc0LZACMbLHINnfNHQTAvY
1w7gP4lYnTjfu3oEgp3pvT/o8iRc1eD+WcZcwrkS9NeinSAoJj+zxINYlcFA
4AR0YJqHxkolVPJJbA7/C4VwnrrP/PCm0W4LSYPH0PyHO4MYkaxSQ3nnVhVk
gaHDiAwVWU55VnIlgKgVhghuHfh0y4jIkKGITohO1M2RDL14Lmb5w0NHMQDY
d/nEjyAV66cW7MS91vuEGPO2zYmXRFMnpsnL8Mk04ij0qagq5Z1u4wo916Co
DnwH1HFqRVJN/Rv+6qqvvEeAOvyVIZuIsABjkI58aiRQeNOFxv6PomxAh4Y2
IoS1zbNQP+SMLsk9mkPSFVl9IO8wkPjb2O7a6UFPjZ5yhhQgcRE3jbALk7kt
lFBovYVz335dETbNGJlC5+vLBU0EwZ3++opv2YBB/xhZxz7NQqb++1qHcbVD
eSv1YQ+lOwpJkxJrJoxfkHOnRsN37T0CF5p5e56VtfKROjdGTkuDUSSTjlmk
5BCbDX1+TtHw6Ot9RpLOlH16AvFoBCx5DQlI0a/6pQi53nkCYbEDbRVPxs+G
/ATe92FTNmO2KuN3YDXq8zCVAyyIcyrrolgHfmE07XGLTa6nMaKCdIw1QQOT
ZOc2HuhTWrRNxDMvCKlDkqXhUZFbsrXwrlgtws25Du62xcfna/YryjXrzXWo
tbkpLtF26yxlcGdiTyJ+f2w4OiVOszfRkSDcCituRVt7zgwTKHQ+O2/a9QOi
9z2P86qXdDcYvE9Ub9u16GPUiKZflsgXa4Quw/coym+7QzSG3XBi5FTifqJw
eJiIlpGY2CryR0QmoBizUAShx4IWnvpsm+yWUbK14qpRO+dlCPo+zrriYbz0
Bh+wYEQ6iKlI968VzyhW6ftLyKeyRlTh9nf4E4t4IKb6A0s5sjZuaLy0Nf89
sSM6IDbqHxvFlT1hioBndahhE1gK2hjK2tUYbazmMM74iRl8nfJ5EZfc3eX6
Fl1hAUnZCe+HKup4asYl7K3MYf3fWGhRB+aO5ErTIX7W8jm1LkvP610Llxxb
V/JTi1Mq/wCXRGbYsW4yxPqM90BYvzzoBuVpvlx1iB0RBrHpTiLYDZvoCLVs
04f6TswnYntngZesRot3vu1fbnr3s9Fl676UMGBD6SO22DcqzdPh22Y1EOvG
2CW9p6ouX/YKmna8GBf7+rr5I3h9UM/KqNFWQOhkUJUkvaqLFo3XNyGM4F5Z
IZTBjTbawHaykmcUdf/F5NAY6KLByrzvHcRFUjec8fnoh6dtZ91dcu6Oahfn
iR2Cqvs/QtsXVvhscdUUjqgc8r865+lPLCzRfGljmnIz9LY5BXgaed+bEgC3
HkzSYkfp9yNSTgJyyHHdWci1VL443giUf2eOmmLe7+FoUaU398o4qks4VAve
7Bsx8tSNk0zdi8uccZaRJt54IJcpXTywKcnmdg2XEvKwQG98g9IIq9s1BuK0
PVAJEaCKHIwt6A0KMPz1uW4MtBbcidXBApAUZaQfaRW4y/Gsqk/EiiiR2b6t
aXlxA4FxdUg88kORNJ3SvA9nOLUOl1b9f9Wq0ttUE46PSt4I4GTbk7W3cTHM
Kj/rjq1Xm+U1kZIaNdVK8NSDEI61oGSlYLj8nABixO/PHVOgnVfIuFEB6ZQx
ZTJaIOiVUDdkxuClFdQENoevygCgl5OeXjANjudvaUTJ22rx/Rk7wi+xvn1s
i/mIIHJrnsbut5ZSZoamIXf1UVXiJ30ew7s9KNtkNXhoTR9gWUvbnphdtJRC
RtT5Ls5+DDXESpbXpSWv66STZ6kMqnlzXGwjD1A3uvXtL672h7D+vKquZxiv
qIBKsrKNj1eUMGVAB+vljvW/is0nXdbPdrhnngh05zo3d+gcXff/s47SVVGr
aFh+yVgL9R7Dh0nK+aXYkKlkdQ3y2ZAT5Efj6WmgoqDa/mMRHCnMKHmElf1b
Kv8EEx+yiPfkxc+AGxEns1cl3/x0JhFaha91gONhrfkR6+bWHBqNylV9ExtY
bXMDhXBe/Tp2jyy/OUtei2NRrMFDlzq3aHh1lhwPgWfvhLVb+4IY9uqvPlCu
S3hU9jfzRgb4xi3J/kxjtaCeZvpZQMJ+py93fdgXG3Ew5te7anhpArQ4RJdV
HCYZopwiZUeT9cEd3k4mHVRApGKUDS0Ha4eQcp4DRENsDYYNs5emHmOy5eQq
9D9ghcKeuz5JkePz0vS00RldVgzyowQajg7Le2Q5SyHp2gwUOhblHQxPfWXr
b2cm6v5U21PLuujoOGbfXh1OHOVW1pO0qrHH26J7/rfxpo3xS0ax9JTMgb+f
mXhXU7EwbXJq9BD2jS14lV7+nY1YPf9quSWmu7Ss4QI8c3h0XWUwoU9UGGd6
M5Q6CJDtc/1wGbizkPyxE6K8vo7mViOvuu5qiqtXeRbnZBaf+AlNtOzX7f/e
iTHIjjb0hXvoyoM3deDnetZyfBrmjqmImsHeEsj/KgHxEegDSwzmVsKSwayD
/NFisT14AMREgiUtFDqx3pVEgdYTnwENFiDhvXGTLFA263XHOJR0rXp24TFu
wimik4my2Rrrf4WEoYI8L4ywgcrgG0IVFaR1ZjKArxCkOUa5/6aghAAiG9n0
dY7GnybCMbupKSVqmJGnwVTuha1eIHK4fv994U5xbvLIB5Tk1KlnK2VjLlr+
2acNaaABQQWXw4F5TUY8i8siIlEG69Uvr7pxYKiJH1El2XShovWSAPftIonn
SSRZD9uQzE7qztr+nwnofjle8e94IFZh9pG5a5MECI6J4DoZud8If3AliwZ+
xICo6fwOKW8sbOBaNapFZvbnOqKc5MtHHPq0e5J26Icm6CizGsXOHhUigefq
TKEY5pDbmUKrIZqVvABWIkaMuAjyw62EFuxTrHBK1u6VJFUkQXXtRXa7zYXn
7DhNaY3gMxbkHPVopJPoaiaJknLualx58B2QHytFHifbdo08T+Zawnwb5PMx
rSA9zq+35B+CwMB7RukxzURTHaKlmdQir9AK4tgvBviEok1Rk/8mdMYnpg5N
oB5/NR1kgK+0ILhvjck355YCZlwkb08uA2UARP/4hzqgYtpVSAEKClGQOxzh
GmM9i+ar3PiD+Z3hZtzYGM9MeA7wFMWVNArVpqO6ntYRJNai+AZ7xeVLMW+3
TfqaCye634as96uYpMDfewnfXdKxKzHS9Y4lEybyABS1ddvIA0JAyUxR9lPq
LZ+ikLgGNVywnjOgWpTTXqg1HriL2CHn2gccPIXtfOJiTo6p7GfIylalH+JS
7AJcKvTVgfJm2wY+h+qunrC+r7nJEF9wWsg83ZucCACP3qXtW/pUaBfNpOc9
Ix+8wdbXGyE7HV331K3XKHALZgXSlPDUJfPR7qcmrA8zkH4Reyj04Bflh1ia
ZeVk2HfZ6zkMwAO1MMYF5kSpWnB9kBo+Dfy7Od11NXSQpFn7yxg7mePHcuZx
nY1QOe/RgzYRqz7vzWJfnAu3bllwx4ho9oWSsGxytrOydnJMEw9soMKfn8Yc
C3dHdi75OlyQVsUeEplQ6cxhvk3p8kpnxhsd+zF99W13C5ZZnL9tJM0fDsqk
qs7R8OPeJBvWyaGREnFRm5kXcfsMscdhUZ/S5PQ3gq4kHbuYGc/x7isY9hRb
L1awATnmxYXElZqjaq8nKq8/WGW3rKwFQqGCrUrzPemedINhmRyfcb0dTD5+
52LkDUGE3r6QPk51m/itpom7XuUvCBP+7OmIMExSBKkDHLUTeC4a/zlzY4d1
V/hblUNkycDqEeS4pdU2G7FUpXY/wjHcQqGyiWXE9JwVWtzD3jf/kz4I6EA0
LXrl9vu9Ew229IL9mfb4+ccTCyLbl2YBRdYzffmHgqJMD1nqRI5wwF5Re5iQ
+QhGUJELhB0JaIqjK82EnaPRcAveb8b/wcBbZN3BqhuDkR8UMLQa/MY7U/JE
4KA9+9NVI+GUbSNQIdjt8rT0HbZ2ouR2ehXI9/6Z8veaY6NTQXfWklFQib33
drjoGw4X7GwzChjS7RRgf5epO79FxX2dep6hqg1vXsL+UsMlATuyhSBw3Gle
a76SC5UYQ9A3dZxgx3pr4XXw/OuVnFdw9Pwr/JtEWyXOfh66sgKfEXkSA+az
kG2B5K6IvLE+NWBeJMgSImnXJ0rXcFH0QR7IiOnUylvz5IXNVjBOP/rxLEpG
3fVcIODAdy/ShW2jW4Ysx0PHOPXbgqLe9P/aV2FcxHezbr2+beywkZGh2pxT
yJwUh/I6XkotFpHBEtfazB7O9LHDcynMzPZ9hPqKlSxAdiiGq3E4Rj43WzE/
XhJVZvS+CDcUFrIyF1y0/aN5GKoWFpV/2Ne9ddnKbMbAjIYicn21oIBJnr/d
y2p8mX9DPAST8SxPkK380G/TUm5YB71vvCaDveNRR6hXOr/KQ5FDOoxjDtUp
e3Z6GpWQRA57e+f6poKeieLFGctOBHSwu+m6cW2Tcrx/U02UeCwbjIbVazNd
AFLC5Pnbs3qu7iwv5no+6Zw0bnGni5og3g/UAFLjtK+emJKM3/OlMYyGCYpx
WrrUXZbZkZ9vhR2e7Mk+ns7NSWvWzvJ6cx+Cj8cdq2UcWqaway0c6ak2m1+N
KdmWlus7qLbaunhsnF3ji5ivMrreYf9fnzUa9e+ExtqO49cDS0N5SyVKDzK+
lJZj63RdRBHEnkwlO9f33megVlj2NjjkaV8TZk2Qi3nvNDynA7L7kkalUCm0
RtIVsgInjdnUYvKGsgqAPZfMqeXsBW2w9b2WhtkcuCy6hAh/jDOPfEe+WP/T
eoGZwPtX7f/i/V/U+YXBvk9LTZcLMSl+YpwssRBi4OesQd+2Tk4bv3HD/JKp
f9fpAb+A/kQy030UuEyM7045DJj9JYLJ/dVVIEuSPr2LNx5Z8VzEXbbARTme
HPWRNeoPBpqN3SPKf3UJTGzO+EJYT6Gj4IV8LlF5RLqfit8CKVrYt/gmqJ8+
p1Qg+xSsbDTM/TUnH9O5EF0uLuo31FwqFDwsytVz4SZigv7PrK0TtJ4TnLql
ia+hTO95yPXjB7N1XUezv/1GTEKYRDZiq93g0eYUAMu88YhwA6CXgjoO4Wdh
3TGeA4dEnnMCM4dDWismDAzYyUeULcXNVMUmgcE09y5C3ehxn4vObN0Yvr7H
JO0PkguaUBL3YUorp1AkjNPyGVpItYBfvA31I6lPugZluvMxucR9bWxM8U1N
NMXpcYxUeb4yllzRjPw+mwJGL/XMuUX8ZPC5KF+MNhxeXVAKnUPQ+aeLrvQO
e4IyNdMY6gaMpKCm7CcqyAgETTh/mJsKHDIGM1pZsM2Q9qcTlW/CHpG7aCyf
e96ktO6/RYJ8k3cZXuhVSrn5FFONOPYWgwrk2b6MQpieRIcbarMHfX5WmXX4
ZsParO9M6Y34fdootXAEJJ78q0kQDFXotlIHNm8l/TYunqSGIbSrCKwS0q4u
oYoM31IpNwA6F1+zxMg7N8hULuvnCAYKcfoW13+heaXIh3z76g5WbZAg2iTM
ot+tM6MLDvBmapU2NUGEVto+uCsVkh9YZkXrnD5/1bgTzv0UraJa3mRDKR8z
NPPVrqwI5TN6GNuHW8+oZGka5sXCLKM6zJ7yqj6FhpYgopVF6JWA9hkE1AXP
MsNXIi0KpkCaaX43S1xmyBdjjU+zQ01M2Kzcyp4ZMCiq1+OZ7XOLDdl1ucxV
9tEKPZ1+vrHdWzx//l5evbUZUcEY5cPHeUL11k37540RrqozEuM3nT2xBmJd
DauqZCP6kHtBlxCGHTri4BEVxFank9y/MP5w2hpRVNzWwNI1u3frg+hyhvoc
q3Ff47G6dzbDF0eG8+CHUGRldqtmPqfRKGODL35m60JZXxlIFzkHAn5CMqMT
saAi1udMbUOmJpCst+wUUN1K0iQ7+m4wlMWwyC74NlDlfzHOv4GbyEn5cTeV
DxFpf2ICCX+l68Y3oinAG1n6psjUaonq0hlBWdfNnaW0dOJwgCF2GJTKJBkx
f3YSzWQ6fzebbE4Mk/tPoqE9VGrGnbRaqlqQtjQkacW7jPzG1wmo75H+EGuN
C3IXWlJfi7mDQO2vd2A7HX8U6Bzp5pU9U9Vp0dWLD7kpnPkrrCn4wNU1FIsx
NL5tNzqdEgMqJWRoI9yCF3GIcjVoc6R/iCIr0aN9i447TN1/AP81UyGHT2Q0
e7eAUw58hl+h1QdXLRGf2ad1pFxJSNGMjcmQA3iaJlBuzz/N2jPmsvcKQVX+
mFSEuWw3HAwP+UNkmwKi7JWhBKoWzEEbUlgHA8xSPNJMCWN7+mfo94mu/1bw
Oe+ttFa+BIkPzTya+V8K8alwZDg/x8abqx/oZjnqLIGciOIBPnVqkvgS5LL1
oPUdXxJC6I4C16p93zb69bHh1gkO8T6/ZMlO9mdUPorYnClW7agsJz5Mgusm
EhPlbLZWlJxbk9N1phUBKevE3U/z/A/B/WmCI3nEmOA9iGcPU0qxXZBeOoa3
EoByLPFuoG2xi7B9OT7zmjgtJv7y6VvfL/uvp6FTZhdUosvnZULqC7j8puJL
ZF5MJkfBmv34eh0zn2g7NJu37cNLBOuqJ8bakvXpgSSxJm7mQSdBS8YDA4uq
Dx+Z86yafcoAM0JEGVT7FBStEPXRa3aeefEB4VtAO9kFFxGWfUxh2V0/R/cX
xCs2pgMp6Bl8shzH99ySwsvoald+Yi0e24qUAac2ilnK7jdANzxuV4Bh12g+
YCHSpcT61DARvSfwvWk6z9lYc4NObrgU1A6LtgbhQzDLpj7fJhwsbW6sITyk
d3vepCI3xUdFggyDRs/2EOh5nPyscyr0BKQ1JKVIGks8qGZkc0CBWsweP5GH
2z+J4OjGSmowgXlNKmf5T1qUiPt03VoGeGJ/+a1qsQU1P05wtv1o5IcQaWNW
sJBZkZ/mNtv66/Pz7Pgw4iZKFXgDTwpQmW1MVIqRApMsqFZp0dwXAC8aKRNt
KR8+R6dzEXU10y74hMSKjvUmH29adbFdQ1dNZCbVilVpcIVzlAJy/Fvaf4De
S/cHb3G3Q7zaKKEMED2J3zD3vQqlTJx9JRq88XVeRkjMFQgfQOHhqb9ojT06
Tm0inyZddGYWz0A8FwQqt3iSYCAI4TR8nTbyB7DRUE0ULnci1LmhMpTqR8Fd
eruFLpfVha+X8W+8FbLz55QH/VxF5ZxgAQHuJg5NV2/IiUEfQUHaZnhvN+B4
nqBmeDyre2XJESzon+vVf+tIjKUNozrDb7L4f2qP93Pbm2w1l1onKfCRr3qm
RBXD4vdPcpg0vJ9SEPrQTAYlAuOaYk9JAadjNupvrOC8KUaQL+6TenMx/xbJ
5bS48PAPhQYPLPUML/TYIkd11raDFL8GxhBIdpYv65i6PcWbd+d8CagAj8VE
/DE1PSzvj8qSGE/04lN4NpOU2HUJ9ozamHlgJW/xrm2XOkUvrCqHbaBdrTbE
vNFjgdlHMR4VhsH18XpnGlojUPfLkI8f6YyjyUJ/xDem1iOzNc0vRwskgJxE
d8f7fiB+6X29awzJwdtlvX7axSxcyUfadIf7rp5ca6xionipyxXtSlg+fC1m
R7elh9bENbIv5/ipj5X2rhT0cMRp12zz/3P8OkQ5kH7fhV2jfEu9XuB01oKu
Xn3+OqPxlcdH+EhsODZKW68lk93rpXuQY3d15wq/Lsr8eVbkJ8EpGznoO2ym
8j3vAgfR+mLuw0TXBNI/MJ7DpLhA44zvc5AhJ3hXEWDf4uv3f52H2uD/lJ/1
gp3JzgHe+tqVns8MePeNLZOooXYHb8+nJZcr47tQgYDFgWmPR0CaOkSBwsbm
t1rt1d+5t37Ny/mnBOIEktGuG3fD0j63jOCEXcNVpXJfOcdV3jh0uZq+saHw
h+v353ybOcosfpcOHk08/68cZcGoMXKIYFKgBjiQOR4ssS3Y+pZS9zW5DAMG
9BlwAn8ohx/iho4HN5l0bAZ0z+AYC/769k1O51grlwKTGzHe8FLJjizQLuya
3RwClSNxvsZcatgsXl5Hk3xNFkQL+Grqo1R1G1RPTt3ZP9lSARKVBIXVQXng
zcYZkj8Q7mvG93HoWLbWsDOTU2psu7mE3OU1lzNSTuASYBptH+LP0tmXzgj2
nDf9GMC23yhwTrK4eqYYUviCkt1ygCsjCVH9rU0Geut+LLwMmPhtzgDbXP5T
p90O5deFwNpxVYc/C+jiDHrAa0rSwGv1ILULOHaifTfm438qzsOWDes0i3Xq
OI1Ft212aHa39pvs/mIKO5e0uRyrrGlKX0JssJKtW6X85P1MOF13StkrJ8yM
Ekqm4wV3/55RjLhv3PE39JxEv5muOgqyTp3mBn8kh4lj6erppilKpeyc5H35
+fUaxXxUc4DgX0GYU4yYBl377h2s/RNovf82h7ODi+Zumk4XsNv0+JmNpv0G
gNto/0JiZmNe0EIhiviLxXPSYF99JhxO+0ym8SLGn+uP5yEnvU0zQhLq0v+q
/vEkoNVgaG501cljB4Xejd43IAN1WE/iowpgvSZzonRzRVbo73MHQexmXfUT
rO73n0XXTL5x8z65fj8/P2NZeWQqxPygq20aXCLeE2Lt/se8QnAnjl8AfZf9
hq0wwjnMxoFI80i9WohpFuwqJA5pTCuAs1FWAUFVbxRQ9ndPvoM4TUPhByku
+oKWIOQT7E6ehcMSkuxJbaDAomUvq58wkksmcXcO2FxXVYK6/fjYbBJ5BADm
MSGDFln/JNkx1Hen/zGvC+45eb9DFa7p8V9PtG/UtDP3CdPWV5oxMnPCNlyy
q8/hH82PoQTwXF29bxB2wDazt8ic+q2R/FJZTb7/dgUDUhAgivpZMxQbU1yt
g7cO62P0Bzg9DASLqLj8PATJLvxBKTG/JXKl2qsq1JcRrE9S6KtUbWKzFZts
McsKRq4WeEpNize8/pZYMKg5TwFAIqZbiNNNjpXPxnnaHuzKc9NVtPXFG2nx
BVLvuu/17+qRmXjdGXJMxyDXZYUsFEza8iLBaD4I43UdQpFY1rnObjgQWf0l
8/fj7TWEPP+0uCZwIjWEiy4dpI2veJsBVtkMmN2yyPO4+SXi/DlDY/vP3uxx
w/k9FRlku2aAG0fsScA8/cRUbkKvF0H97DTJXiiE8NCxMT9tofR3F4ThS2Fj
5I2ujpx4EJGPBnBc3LRj+7zZVOqDNZ5CAaiAgIp34DUD38m95MMU8rEsScgD
l08Qy5cnDsUYt/TaLTV1QEUVzf69eMnt2WpQC9JzM2ysGcsPE94GaYWIIXKQ
nbw1Vn/rBR4G1ghCAgvHOkRLruAUHdDwGHtkirTjWYIQJk+eT2E+TUWbHsSI
8QIfxgLV2KVFd5iiUlre5jh12gzJ4l8hLLCAccKPUNW9bgq2C6sp56xS5GVn
VX3JqGLZtbxqAeJJBjNccM7YgT0hrbdTVpUye9tGOX+4pGVsRAiU4T8I9E2K
g6RH7m7zrw75TvV97mW00SWcyYu6GSOgMQ6f65+kXG//tEQsOzT5dH115MOB
e9IGEy3sLZLdVxn/mKeCuteMs7lPrr/bhr28fNl11uN2di3bhsWzx0k3IIom
rFs9N7bQlg9+xc1jbtHyxhGwEVJVJPQ70LDG+0yASwI7mr7gGHiL16acXC3G
Qi84h6+fi8nj5L6ytd5HzAXX57QG6pzMFuVm32EVkhQkSPp3uM326h8emXlB
rwxv15QxbTLFHrjOi19i5IFJUleCX+v22hJIYvmuV9qx4Ujc+7lzMtGoSHy7
ARK4BH7XMuTH7uCug6nazXlB8IjPhjOX6SQtZKXN8heP9VO4NZ24YvvTlVs2
khPWDXrLZVh8wQFwJeBBg48sDxT4T6c4fOw/Eya3agPpY0DBGw7nYaqD/5WP
1AXhQ2my+qSDIhikqqb4MRF0oqR8kxGiWDtsIGdGUazd4+HFf8TrXtIdJoxT
Jmcb6Frw3caWAx13Fndr9rdrSbnh0I9fy22CAluJEnQGYAuo8cumFcvS+EMs
3xG8z7Kbe0roZP0wXZ7IGMPrrcOutIW/gfx8fPjlnub1fHPpdNEqDDN4mUdk
DJZZD6JvfQARgV55oRnvsYTfDTdxaO5hS4jUX1DiZ+DgzxkBO+WvkP8EPEQU
G4TSwKU6+LXf8pauhKjI8J5K7dIl2EnWpJl/Ls/OCG5r7YoUOMRWkyrKUope
pJLqOr+0FO4aUVwdYYbBuQhXnhY8GqrFJkkiJuRforzBrrbsN5FGn3ZfzzBu
wizip5Gq0OssmFnBZwOtpjdkmnD6QgcmPKost5QEahwMbMNNePZvR8xvbVqh
Tjnhe6ME3QzpnzMa6XJLOzpHaSTuZm8Ec7ms/g46rU6oLS+6n13z3H+Y35Tx
7SgyrvwpWik2guEcfzu5LKMv1Mk+5QrdJdb6xNimn/8XiBkcwXg9/yz9Bzm+
N0G4hQ7uH0yFZ/ESBuOh0xb04Xc3N95VUgwkQIUeXM4A2NtE7LYNmIwr0fQS
pVlfPDrMQAUyLBy4cgLJzumwsy6M5xhn80+7RJrmwgwspf8Eq9JPwVO4UvG1
U8gM1/LyixyLONeN53GRz3FG3+nF9s6gFiZEI8VolDjzPt1cbjNWG30S9Sg5
MecoGHUld+VemXtW9T9RRMvk/DsiGRVH91uO1At3XnjUmewVF+LurDN2vsDW
vhxXAZhvEL1WoBEy+E9nYDGHl5VfeDbEhsx8omLVhftRcQR0sR/TVTp0Ycsb
TK4R8UQrz3WzW2rpRKA3xUxWUn24HYY065Y2QE9Q2JlCkzjCGNTYCDd7Hjrt
li13KrW/MXskvMQzBglWxggfn/01OK7I2Qvcbor+yxXthg5YngW0rOGGwKkX
KKoSDdMfy0y+vw06SOS0jLa3b4IALW9V3SrvhC7gL2AxFWasZMdVsDbSX89u
ggKa7Zq4vtdTSLh9UVEDVid7iRDGErar3LdX+Oy41X8jQzcwmFXKzj6jTkQH
mBiccXiT3qgJtJuTDAg4e+pDTdXSJhNuy5gAxbj2gYiKXnUG4QdTxGFMcPod
occ5BPr82H76RMTmbjiC7XXyVDLtmjFR+CgdVboMH9ckGUSs81UFgdPjeXtQ
cvkilG2jDO7pdAK1PO8fq728a9eYkysv4+VeT9zeAK97NWyaAdLG/4tw9qOR
nFy8YAoA+zs2hExShsJL5T/yfbPWedMjvdVmqbicz3Vp30XMCwIaeOONWdkQ
6BlZlQlsXwrYP+nRhshIMV/PhxjG4x6TJY8eC+z52q9ep1y2aY5r3w4RhqlK
RKFN69QjO8TVhb2AZEKdu/2LAgN/93gRLD26rrJvNys9h0i0XnKgBIyRgeQO
bk9w7eKeqEXHJMvLPbttmFn3CYpLHdETRA0gik9sTsEel3+DNhUxth+33q56
rTY3psOvnsTckpjejoomedqbqwrFx4yBFxiJ9/xEGcQd+dC68FiQPTSChCWq
5lsOmpUuecUwM/x3pFVRB7XMPvhDVPiqP89xF8ftzAZAkt9jEee8atSObIoz
32odqe6PjGsnumsyOEuf/qbDMHBPcox+jtW63hPreUCwjnozN4JKHTjSUgnU
zPeAS/fgakdR4fEjy2dyFQKvCumAHp4kwuT4XoT+yzVcok8l7PNDraqb6Dcb
YpofSYhRl1XxhDE2ocrzlFoJoMFAwtO8JHsXBRooLoDkrUES0qvVUfy6lIcl
orOGblTkAGJ5PhJ5OvmMEOj7qkmvzWpksl7rwGj77fQfrKj7vow1eMiYAOnh
SH1KMi+d6SUIc484ThHJ7QqT1Fa2C2tJY2sZergmLluf+mE8I8apnJy/k7Y0
1488yql8PXZd9zMdE6hlrFk3foq8/Z0R7hdeWMdlv/haFpgaFTQrKMsyQegY
isQ4kU7IZi8xwY7KaXRYrbkArvj+qB1AH+endKNKMDYYeN/sFB8paUdc6tG1
2fxvKZqPAJeuaIlO0wrQ5DQlw5DiFXiqFBCa2+8DiiRYEXno2oAXdl5bFNt9
fQJsdzqlOAIVhVPbPP8QJ7MdN6+uzfXDv2qDTNGa8ymtzWuGiRg+9/9x3cTF
N0O5ay4VM4TtB4Uh0WuThKJGk3/o/FkMgHY0gJus7FN/z4HmXkg9Ylu20kZU
tF+cIw4Y1qbSU0PjSZydWambd9Ei3lw6WfLnYCiFwEgT/uF2lAx/7/y6XbMx
MTE5D2AhQFqgS+99Dr5uU+gR6keiJIWU0MUjscAaVZ0ws0L1elMaSxj8/DC8
RqkRN8BO19UrXyvpzkgls/zzylO/Cv/ck8IBpD+zoqrpSs4VmB+gtTjx5OO4
Q8pJgyi/77TvtyujJYA/UiXfM487w4rSGOHwqC6al7U+XjDQXWc2yU6PcCEJ
dhjQxQ2m3vkZ/GvrRY+YB2rhdsw36z+xsOPWsiuKkdhsXk2RqSC3SdErz8zV
RbBheZExGz6cC9J670X/NZjLbOFtbklYGbvaE7+quzFFC5/zV79J7yXy4f3J
/9FjYhh2mm2kVz5P/R0W0q4gx+JAjz49pNZuLEzBptvHtC9JALg4/oc3imJ8
Puw/WWDPnNmyWd5FvnfoSC8xiYTAHEM7f9/DIv734S7OhoXTk5bNxXXxkY3s
oTCE6X3QhgLzDGcHhg56bTyDKguW6MzJqE4sKBEiWo/oaMNycWcS/cYgqKhp
Gbv7c8vis7bzNrx9qlVhKksdG6zdN5Qa5eny+SJHV3jtdPCEqyGgaJE0vA60
Txr6Wk94rn8dpcLcowuwkbd3IOYWOC+9J08qvFBornrbfLOTjjDUH34EQHuT
5g2rHimx0wh6sSTmoqunsH2OVPS80JPlH+V2W6p7nTTihDYDX7oM6q1ZPXxl
E33Y4jL2Fps8xOMqra/Vu57nMhud/kXCFKq61DO1T1tnup5uSVkmOvi7m5z8
vIXZAgeQGWJpwK5SycwPwJbEsLwH6e2rDA85r8jd1tAlrRLFX7w0j4v4AMzk
gpCYkLBwIVREuwbCbvC5d44dlyCgT1Uep96vJt7c+XyoE6IslDbmQiI4eX7t
t4Q1A1TjJhj/R5yebzJ2yq+MQMFelmBpzLTIM0y2UeZTnlzEImW4/6RFyOAm
k9EkLlV2+5mQdJ0vZJ9P/rKpAvsJXHiG3kTNIK51htTEJFpKFoq2a9qh59RQ
QFg/eHtbLDLoodKf8hYa8pZZWFwiNIqCsx46Ebam4JyakI1MJOTku56kCjom
2T1b57EzmYaKlzZbW0UW24KYSl0QXBt32qJXxlW4QsS7TQKKFkfT8qwXE6Xr
+Ur/lhqPg7pZd/fkw8mCTuAyAnl+moD6MLSy/YbtdoiG2ZYH9ApOgLP0aTbN
oSv3iCGNGyuQoqxdWM/L7X4d8tklw8myobnU9gX2UhR4oYolIXMapHCmoDYs
LjhriTBlHVIQdoT1R3USGr+xEY6yW6J2Alj3iCB9oJm5K4VeHPq8ePdE2RhB
Ex/v3OfMtsYbVqNS5b/bOj9sr6lycikb3q9P9x5Et8Meqa0reqKvrK6fPt7Z
fyf1Q3Z6zD0MnJ5tIrlWEc4+GboCcyD4ThM3ADkQbt+1X36do3I1XiRuS2Wb
4xSz9ujN6m3KSRPu8cEyQO0ZRp9m4oR83jA9g6CVJY2CVH1137NHf0idYDwX
q3DuF5Ucz1K+z9o6ZCnby22dLTm0+cVU8j01ynQxeJiEWgiMb9fN5ZZGHJmH
YP6xwTuw1yZbTi6VQuk4tx6/T2+CP286sqWriBvniiPVIIys3pSA82dw0ZtR
926qlYsObSm0gvuSIao58hxzeQ/HBTHGUR8DG4tru2qf90i9WPjqPKRuCCOG
FGhZcQ8fDmz/7fP/oosfgA4VbOuhgRG2pg8PdD7nWbEchGUNL+byfLpJclLp
LG/iSGa/NaWHm+D4tgo4jYpwgpe8d+Kd5tdIqPc7FRAJC6BfzruN713NQvtJ
MY8TOKAE1K309Bv8Kh8g6/VnDbWZJpte0bfdeSRCmccFBfDXi82S/CPt6wDM
GEaMbV8CXezGJMmDCQbjJ/j+M7fknMOvouiOHPCYYDfR2BIwsxd3ofc4M1IC
CmEJHR0o7Tk96lLCWTRtRBHi+sdiDsBLyDx2+ZzgmMxtfuRWQiK6L6ccOG6K
9UrZr15XQSFxq/Sy6jc+7zYXci85oM12QVYiPic9ZzPndqQX/UDgAt68GSyf
aG/FfGokuVyH27H4W8cfQlYHwhaE9a9G0IAp1JLQFb+viPcQHQtmE6RP99CB
JQnwzJU8+tMRrWarmhtde23UkpARHbThRQWPkPuhlWtM024IoyMh4GpeCLdx
ntnWoeW/XyYtk5O8JAlAHtMNmllraMxTIovOQ8K0V9mwObQH31OAs3wBD/ki
8JHUNY1tJeKMuGnoUUzNFicoZoS4zzP4ZtaEsbS05pvnOo6ri4fdD2Z/uIcP
++GV1xOEPxrH7mU4RrxWzNMqdZ1ZetuT0WWQoWCcUhMDYCcjEe4YKGXz9H5z
uWDsJldfvmAoNPGRIHTRAS6uXUyn36EDVXeuCpIuyR6JM8+v+8ghL4qZy4zf
21Y+23DPsQMt/+qJ7fS3k8+vbXYWAuLaWAVcax0iY1952kCsYLPZ4R7kQgDK
8srKteSYAQl1XpmE7AY7xWYTOGbQVA6poMTKk/RQLZSPSgnfoVsZjT2G/e0E
FZuxktQT+j6sE9RcxKWrgmohNISpIbpTZEnR1XE2napmFN42xSXq/1TmcXmQ
ZSDooDNoQ6eMfskhsSIAn3OiH9T9kD1sjnLveKwUt1Z2VKbUpDtLTSR0FjBA
ze3q6oMOMuCw2wDvLNljnEI8uqJLFNtnG8aRZhh6pQ+OnDwhSO42qUns6O7c
2RDxECIJmS80D8AxAgC2DsK9ikMmTZqThrxHuLhMGflSR+Chnrlu3bkXE7y0
oiVfnuNZHbkDy8qsTkFM356TzivWtxsN9W3qZlTTNYqNnryXxIeabiOjhgX2
hHr5yCutWuZIbx1ZznwRhQlA93dG68nzGw1otmOJKIiiXhGWLaS6VWafXlvh
7s2LbDkwQXYMUGHH2WZe+n8IflWddzv1Siuw/s036PWpafWcOFvcfqq/Aq2d
54p9QB++4GzGblbyb0TSxYrlCjeV97yuUUmPRoo/mocEU4xh4APOlOGRXmnK
5tZXjU15XzM+nPjIWwH4T2hCNddom6sUxYAwg170B2YIkaT6H98k2iGFFhsy
FU33dryjEFUGYviF125GPzaY+cpOx0Kmo9YlwTcfdwr1wc6HP8NHj6VG+PMU
7vlzUVBiWuahtmA3toKwJbsrlSeAuo/ZV8K+VkM06Ivj0/Sha2P4FcPB4mRs
aQ3bRe7srwAeVRG0cr75S8AN3St034TYCMbDYNcFmyoAgOVa0js+WIxICHza
pdvdeBkyI0JqB9XP7JQbl60388wWTsIyqcUviFrNUmMBr+a0JAe7E3YsRcVh
QWFBhNL5SqqS7fq8XCGJJCrk8kpBxpH6QVoLDPtqEWg7ybXbl0qfn6xHkSck
LRLTdBPmxCkZSi+n9c79/KhXI2GV0/mrdTNOVVWRRcTQcv4Aat8+EM5an9DV
Gw1U6I9+oiJsuc9ODoHQYdXkhTWqthz0hkrwEbjRKXdcCYFCEKsOGtTJamYO
YVVoy5CFAiCH+QOzdjaY+5oTs8KBrDoBry9lwYiLpoDMbK6jC4KjLDv+GRug
x7zhrNE5X2H0FN9yVXKSMXzag+WgeUC79Flmn4AjBC0B5W3eIy8/kUr0Bl0H
jg2QfyqIKaBw3PPRA/j4JGrVk4ANehoW52gSDs7IoeqouwokgOblcLHpIHsl
5GU6lydbFXQCIRtUrfQiBtmyBNH8ianAm5oCvmXB7tH99MyRz9Us+bYJzjLa
zyROcKH5H8sPPvEOT/yMZeaf9hY71jSV9f581UuaVep/9GHPe9A9L9/jB2bB
83bm1s7ij69KI87O1UHbAkQ9Umf23fL3m6K3xRS6IhXlyxlPxS9b+TMbSsyW
n5G4ki0RBl+zkZhl2RI4CAGm+Ow4g9Qzljw5V3sRa5v1WOqN9qPzYa2zDKw0
D20L0WAww48duCoEdohJE4MCRL0rmv8qGlWQpYqm76iJTGrvRKWlYH0OBPd9
1YY38ptTVsCmAFBQungudQg3nPj7sdjIK9gkK+EFa8wyYP9dWlB0ACtyGr0G
QwmYvFkwsHj36Lm+k3ahUPus3/C1D1hXkJC8a42Xh0Zb5/7wcwIugNu4f1pd
Xnc5Cz7D208cLXl8U1rRP4JgwXzQjL3fBKdMpDMYHesNVIwkLP4IX1qk7Xtq
jCW+zweVeu4Do5NzfKbgwXHnihrLAOgL0WSPUyjIQW3SAg9cl7C4cqFeKvNP
H9+jT3k47LA/rUAXi9iOS5tA+7cmzRyET7fxbIHBheAWpiBJf/eSP45bmG4k
PMjZd6xTGBQpBMs3QzXeRjDhq7u2GMLYoYp93lLYpRuf7aHPmmHdqbQDagHQ
5/sKbdtIthgGAkuWxZXxqzXkL430RJLuy9hMdpPpH3fbm7+oWhVm8HbLwH9j
CH6/g1Boxq5V9PGx0/ECpTjvZSnD1UTkriEdPKGHyHJkijW8cUpEADaeJIEb
n/JrX9ePWj2C5+N2/W32lBJnt1/UbwDwabserdxwAF+QPikz0e6IIrPR5dni
DQYVj6TQlt2w9bv6ffJXESQ3/ViaehjPdkzpTK5I9/Ibn/8w6M6lZWpTXQpW
Sm8ZgB6oTVOjyNfF3OsEGo1Awg5t606DA+n60pL6zxBWeUFxXEvCBB7foQMn
+p7bgFs110TtubgJvKss/ma4zpPFCEuNe2aRmBvr9q1stT6WlZMOs1sOb9bS
9SfZT6+zgXLZ1FuOMsmhbSvchIQqJIgERduIfHQGHYJDhsvv6sIdVOUFzQJ+
D7YAoQvleTG9IAXNanDyxmREqDhOAjt1wskX3yQ3cmpfUwZ3XZgIBMurbuCg
OtMrHPyRemRIInJKkQsY5wJ1PRFCNMjKS0L4SsIzA+rfaiQaHt9TjVOmyc95
sGdOZANlDdbj1bj10w3UV3EF8alceLKlEYD4TwflnDAZoBSmc364iAKaFrkQ
MOj1B2K9riEWHjO3p+LdQFuOZrb3+DP672/gFlms7+3/xeD9dqXZD4uzpff+
1RcfdxCBCEyTjGzPtD/0Va8qFigMfPwtTzFQKjeyR03C0S55VCkkZ+6Dw01H
R/W0yzeK1uo6hvCFld2DoXahK2Ml8+6hfHGYa3fJP2B7LixtbeSVxv8LSVzl
mjICpii3AHXqxah6UIK0V8+8nTU56JtufpiY0XFNDq5xx4A47ofgYkz0w5qY
wyrZxQKIDGkrYYUU9OvfbftluZPI5El4vvx0mfw0H7oeQC4FsWEeAMdGiWhs
oT3XSmS24eblmZf59R/EKUqG5uqsS5vlYpy+A683hpXZtyzVhmS68iA5F8FK
dhu1r+F2b5KU7e5JNcNpYybHLXvkn5ktMEoZjCfJWLqXzGxFC57Z+g2hNQSV
IX+OQldG7lZ8SZDMFqPHjhYlTFw7aXMc3ki7rgTSC1Mk25Ca48RDqdyYjeFU
oJ26r0mdxYmGArD4OPQFXKZQ8fAZ3V7vk82YJaEinMBfr7MQXUimRjeNoZ/P
mE5swnzJultPuiZw/3yXSgRrtDBDeHpCvEjjCRCPoh4ml9iMXWc701YIpIV6
wxBlx8yUfwCeUrkI03eSxTzFbpsFH78jBMEHVs/eYTikB57L91tPSY/tBaLl
pk58lNoc/MiVP1IrHcfEtw0WlTtYTnpVnyjewrCn6WRfXwrtVFKgVLqL9H+O
//eXSRC+PIH73ZSfscNH9o3U+KfbIf82h9w/hCjVufye8c8NqvpI/vGbUmCa
SHU8zOG4Kut86byJtP7IxUhnFnmKwibpS3ajkHdCDTqe30Bc2flfmFmtTw7p
t1tcDRRMf3+LjrKdx7VtkvGBoPLysWPUGULPeOo6SlvHWUEztEZtaK6EYZJK
vIcfLJYzUUYPeMsFBRvWtqx6uNLfR9fPIy9iq8y+6xvi2QQY+dyFE+97JdeH
pQSVRHn/WbaCrckybvNsML+SbYfEkTgOX5liOsG+RYPCt3yUNsn5UYY945vp
epf/QoBaOjh77b+aEQ4JwzwdDmHaV7z5WxiieASPc5SOeQzAQe4qabsp/HVa
zl0auEWfxCdF0x3abb91Uw1zrunPPU9+0+lIMNkoC8ntdkrd0S+5fHgdZzbA
KZWBfjulPJQq/zSravhE81/Omjbq0+8FkAlBpS7LDOSf8m81h7ZD/tbPqhox
tJL9nDdGZqGozw9+7V0nljwEGU4Q/YlvzFDK3yDvRi2Rl0q56bHHD+2zEK7i
i18Uk3Ipg9+x+gxlolMM32P3MBB4iTUnonQU3+QDE6IWdCJWge1RtslK1Gcl
EFSjtrQSQZd47hYl8eazMXWSvsrzVluyvJVG59Cf4vZKwDAtJQqOL7Y4XXxY
NnmHnYFlyvQiaraMNjhFmySByLoYiHDGOzKq0RpOkmLlD/Z8Q+FHMUNtHcMu
gnZnqe4ILKwMZgWbw/RnUIqkLGnSRQOdeNoSLk/Ne3nS9FM5de4zP0KBlmBi
xEU8WR3AtSwZNdJobKiNex046SM33JM6/t7MHDiYU7LF0ngjI3yC6ig90O6c
NQT1Bl68B32Co3CZraDXFhisrfP1K7+NvcCtbkxe8jEcrKaYxZ73iBYHS6ut
0JodnfdXRx1D+qO3VWBTFd3QNsrl6eErd9+6pH6bFfN2pREhhGN6l9kUWEhh
YOFJGWEjV8Sqx3WopmvTL/Jz24Y/LNO0l9xlyoLhwubvwPLQk84pmeaZhh0/
o/kk9sWdQB2o/s1C4HQq6OVG+zro1RuIjGcHXM14bzx8cW6oUbuqyFye1URB
xmA0ye3yeUQchQlET4o80LWYRwyx/LiFcChp4V0LnSjiUf/bz1/uGZK9CE6C
QyFMIsdkiBLmhwR2bL8Cbto1pHI95HTlOV4PK2f0el/f7v5TO3StrNzz31uc
OV6PLbUc3gOQp9RiAccDg90mLVVj1NhAp6LNFS0orW5JpZ2fl8uHs+0yEfFo
0ZjvRdciFnku7w8Uc+Ue6inLye4XKfPMIqbunjM1CeXLRyNWEFR3SsAffr2g
7E1Y06wx8FCJY9YSQ9lzwLjJQXiaf3P4cVh+Txqzb02NFcJP5ean9dzOFzbD
El64cmon8hy/pxYPjkMiOgSzGRipjKPku4Zda0CRwZXrGuZNucZO7u9EnY+0
jlngdOvrJXNap+87dEf7+mLAZPqXa/CEddZoCewyuFgndFgmNvueR2hg+D2g
Bc7n07eVaMjA8g7Q1l5R+u8zTuerG7khe4DbL1LceICntWXYFv67bp3yrYbo
XKj/RaUTVqcjM7DCOF/yS5K2ds8LxOeqfywddk9MmVQgUStu23KKGj2x6J4h
VAc7rIx34rVK/E7LDFiUAW8+sKKXfWXUJO5bVgK7bRQ38tichFwuNoiifcIa
TVOhskV7kqbwe55uA28S+O6wWFrSxfuqcsDhA9YzCoLQxBQ+HCvXZbhlwi3W
NpXaWkYtcz98la+8lESwXB4tDSHV0T1n5je2C3wzxeEbJORUOHSqowBVfmHo
99BedFiWi6vU12RaaWLN+Jnxxc8KSUp74MXe0FIrpoGpsvB9yvCowpmONUIL
/910R+vZ5BZOccUwnbj5aWevezXLgLUkK3nqHpNr4SZgbEkTP3gz+TpaGgSB
Lv19eOXqJ7S8/TQX9YpNTRKEd9Ah07QlPUFVNjyGAiu7V7kTh1LdBpBrsTng
I54TZvc9Xr8DvNk8bHPwZ3jf2AYllyfkRF2THAZtQRcRxhSppZ9HgJxdvaFf
Giho8qAgrxwvWpmn+Ke2YwzCajyjNqGnHX1WZMnHlsmtgaHq7hMafBiyJF7t
Yf/nJbZImq/Ljjq/o6kkb1ENXcc/osIm4iJbSdSvq0OeOYM60JH2SuGZhD9b
6iudY9tSsVveRpTAmc5UlneRUA1499+7S/z3TGKUizFC6BAGIryiH8uAgPJL
p4SHM78i4i5VJby0GzqO7qRC52F2+laCFLogsfbspXChsTBfmBrdendYaRhe
3IbzQfPf2Tw34WR9qqZFCBVv5hkShiC9BaLcz1hYYVHjD63LlEKdmSClfEOc
uwumWsmZzA7IMc0B9zi4hndn/3ZYNnxjmy+H0Cc0bzH8zMwgVPNfquXb0TmH
EpRg3JkFntx+8WxQabysEeiQIEv+PKU7cJQjb5oP3/HEpQvN5cMoo02Ggf8x
mzcxTjtQPbeRMQWrUvuyU9kxG4rriUez6OK+spSu4JoI0dTkkhsbaClO+lQN
tloTbFc3krkdbofSUXgA0TIStaU5ZPOQ+qNF1V30jBW/obqdfghy5xD4osBw
exv7Jfr/hRYUpOgoKOUVhXm4T4J8I8iOaoCUmaqdtqml4uGpDIkJjWoqTQql
9KF06CSq3U6MfzFuECJVJLwLzPxXEDiwaZUT+wQgOFzpPlQ/TtaEN/jA/q5s
l34CmovSfrJNQf2uKKHZJa22eC5tf0jdVRpG5QJTeT0hzdWxgNG0Gw5VjJoi
7drwJTUpXSBtDSKtaxWhrhClP/eeS69hhqGrAOciw47df+JgTD7XwlicpIxo
PO83YO0A3smZ4PJK1AKNuE0nb13W0WPSi4HecMRs0x/B8lQMzhma1XHNtYPW
dKnvtKzf4vwZwOOVjPRPKFGdCUIPiOSIzbasxBk7hwNIgLAjiLaZjZpDjCAt
uEdMO435BCDEEo0pZOw9ipYS5qmaXa4+rDY5gu3voMbnl8o6gWYmluXzEsfO
k8I0/S+puG2aMFO6RaESAowa7Sj9TC+VKWC7yFj6lYIygY4okzpvbFaPnFih
gGHlV2acL4rjqcy/xdl5ZW/93iyK+noHSCVW4GUMOrBq5fYLvjcy97tmcQzu
xR7AkSoy5tI7dHXljvfOokJ8tV9Ku47MCS7lT8BZj6fNY9EszLBmKulNecAB
VVQ0q4IdBYdae1f8xS3C6AhGjx42NES5PeEWWHaZ7fXzEQ3R+P0itOYzbltS
RGbsntfoR6d92RCHr2T8RP0tZFAGCtE/2GWIxRB8DC5wGmho4Hqfv3YaDeLH
WiOpxbmDs3FLnghrZQ8mxJhq3MFDuW5ntVRdxnnl3Z678HUIcRNftEIKNMxB
SB2FLQ7mECldQ4WB7ItUwhP79igS5JjVzTN+cJ19jLopuepwp/NkT+saxR5w
5P7R8YuqSlNWkNFB7jdjFQBeLFXOwmVPfkdqHi4d/j51gP+KrznKrPNIeT8v
OHhwmXAXhLBj08u7RMK8ri+Vg/4omMoWVYeqyO06++0fLZk6uWc9gUkv/MW6
HRvOYMnSmR1oGFEjQSB31F5HHgj7HV4kjwx2VoKQ+FIBPoyoF47Gx1isC4FF
4U2IkhP2d+kNDj+B3HX3cWDLEojU7A/aWQ+L2fnHFIkF5IKhw+znlNYse4QW
AT2zb6MxJ8b9FqUesMQcU8EO18IPrX1+SQOacswFrMSrD1R+EDLBDPPzhv9/
A+f3q31Epv6lC7GflimqfWzuPBu6xw/aGXas3Z89Og7gGCwCYeR7ErhgPkYn
eD8yMR6lqoxn5T7DEUSGfRUk6oBIVafCNakI7Le1WckZvnlmN1hOtF03vdzn
To8kwPe1fihctj8/ArcbS9sv8hKmrMDRldCzdc+RXp92SwUMkjOHa9RO5w0y
IrA1ufYQ4xCA+MtTRpLi/7q9fD5ydh7nDgqfm3SUQZLlGDfroWtkfDgT9Dwq
DK4DrDwfAoCcmKV1ko5idCiOa8cIPwIMSB28h9QStyJTWJ/861n9H4Ex0ihl
fsqQq2omJ2Tld2j5yoo1d2J8cteWSHjLfX3HwHjAnsYyQdPu2sprEdo5iiv9
yhLDdhkh5Lt908wURJhv5l2gUlkjUxD5UGOywjrLzco6p4fKBRflVhr37/cS
hA+tbG5MG5Eqh+gVn4Fg4d+B6sKPCA/aCQsQrvvi6ksGVpW0A2hxWgpoKW7t
+AyS0zM5Vt/QPkiZvtz5ulV9uZM0lo6+JoSs2AnKDhA4pp1d93SdELgXQKL0
UCjgr1ZjPCrkRp6aUus2W2NFHQMwzCOx5EuKIxwgSDGJPYCkU6ACFozcevwy
NMP9iKbTniRkErs4hMgBAJKIVqUFM1Q5FOfndoi0wKoof/TVEp0P/FQI9pAN
R5XArjDxzV+mBqpUeTesHU9XXshW/S3Rf5mJcF1TYZfpjSgMdlRSsr1s+8pH
k5oRBHCqNgDpHJIPv7XFfvvo0M9b60HNTHdJfnyQKBHriObGZLXO9Rurc8eA
cAmGbYDIQiZI3CpM3oXCYyv+8lTrd+JS+NEZyERapfUCMcFLP820dxmtMpN7
/43wO6rIdmvBBWSU20vrW7UO6pSP47iTEVnw4zmO6kubJ955H5AteVBNosSE
YCof9YV4xxsufy+1OHd6ZgS1RFE85g4Mq2/oZTAovGiLipGlxHueoov/TCQm
+v1WbZCBBjeUvfbvB+UImL3rJTxuM4iE30EOMiS3V40P+Os2GQz+jR+rWb/z
JLcQN7Y05RhGpPOx5Xr0yLvUFp/64qLeTf+/ht9czpZTO+NesaImIR2aMB27
awMwM8XuNyF08yk94a4/9qGb/xHJ508eqrhTwRuIWTxrefSMW3E9juTfkwNJ
Igs7JGYOm/pXJ0VtCCHikBIpU6bkCICW+nxVtpMvlMqgHeu4NGW+RQK0ooDG
nkoiNYndT5K5aE7zLdMPoq/3Ah0/+DlvYavWJV9UrMzAkEP8ZtmEUMji5YmI
9nKo1k4YrhxhU4HMsnJdFsJjTasXsYFjNUybH9hLWQOMcjpAuksSeMsWq35A
O1VB9telAEwQjNqnZs8nMzmZYovJVx87xym4zvr6Qg9ULnFojk72Cf4rqiS1
lja4OafaV49pijJEnQ035dMs6fqrQT4nYWpChjj0msqIR2/eOBmRDzUxrTQ6
IQapgB5LrGIZkFy7cQS+wp0c0llZ2eewnsZVnk31yPTsWCJAarvy5TnAJ/tU
gPm2cT3By/VehAEVWpOoBx4GFUOmcwIzCwfZ1XOM6l7eadeSllJGo0sxdnDd
z01Pi7IhlJ3cu89p4C7GoBjHEGY+pmp/D0XmgoDwIKjMg8trjQSmgqjVvVMA
fIwYESUHDXCWkA1An88kcSv+IQSWPfQQJnPNOcP2rYJw8an9fXoFuLT3Hs8s
Llth+ehQ9N7h09EaLqsdkKqphBzsvw279CpV4CdbBXDMuOI8Ya/WccfO9MSc
eaYEV9triEZKKS/ZPA0ko53YsLPUUTNotOdak/EIgPG2y9sCoB/8f49nV2qS
CPDWr/KkI4CgnoAAdQ+WJTxeWwnth2LJKa5ATzlcC2e0W1u05eFeKjFWRwKQ
7+lVm7Tdz7tJQbY01TPGpgR+G1E5pjOtyUAK4gSapSJgTyKu3a/OMEIZx0EK
Qhds1qOoHjGyM63v0aYH9zwTsxfi+QFmteeYi+zlydxSQOM22v9+B+rKBu9j
x7D1+0TpJfjR00Ah8IWaYL4nAdYGj43PsRgqEjb4RKQRky5cty05Fpl8qpkS
KB8D9slu2FyDOoha7Vvn0J6G1GIhmwRrPneyrOc02hylQcYyVtjdzexHXCFM
j8F4cQFwIhQvh3CYPiSyPlUjb65FqTqWHcYkQNni+g8XyF2H1bgP6BFw8yYp
67JOAN3panFmD7zIPGcwG8ZiAyEvvcwQopE9bXtPJAkREoj0nKbrAksSPr5g
03x/Rtq7F2+ZAAvhXFwwjecSkBJBZa+QmiiiVNYBUtjt2Oy5Yb4GgiPtrplr
VJIgiNiLNSBDwx7RElWqwBvvd6CnXpup8ItV6D+4X86njbuPEotguG4PM7Zb
G7oHP0XKvOAt3WMNjCq6IARCAhx9+sZLhp6eMbeWbbK2H/vsPH9D0JKyDWow
wNEALFrH0l6G37BgjMPm+5e9sKdmHNOE+5Opx9Pag3XXnqj+WapvbbkgWPlz
PUmWUttI20f1/nPjHlZUxcyA8vWQt6odJ8h/UkvXy0mgxYxJwz+JN9ia3nyE
TyQ0cNSaldWrebr85Da0g/i6BtLwLniRuL8HqlzXcb4lBTSV+x/dntqhOBRf
MD0mhIzzPpd4+EUZfbIIzNRdjcC+Rk5twgoZop4HjL6/1uUrubdUGWdTQMw7
s0WgrsojR69QXVK2lvQXKsqvnnyUFdO+6SXq0JZxMYkZp5syMo7oIOc5/ShH
mokp/ALN88kJ4LQxnH8QnxC3IJ61+9u83nkkSkaBKqHTOn35QOJ+Nz5lzUoC
s48X34kWEoh6ets+jv5t+acy9d/ROwHNslMcoaf2qZ0ADPOJrOYXDQcHzjTf
9T6hy0TjseHrFmrQU6keoYBc6lL9UDlxuIpmtfv3gBOwVV8JkWyf6MHW4/he
TNozKksteS+HDSs/SEhgDeOeB/NwkFbEb5/03fvHti+lPcTLEHrRtErNzQRJ
65FnoDOZihZ8cT0GF6tuL4AbPELv6YWIiV9dtnJz1O8T8StwI9x9OV/MYNl3
GCM5YYoebGxRpiY67/xIyNN8g9gKICqrKpelRrj+vyAWuwM0+Jep2qb5wcpD
Pdss7A0jQoPsxXhuoLklvQViA2aRslK2xH691FFIg82rv+ujgXQCIO6MY4Wo
i0j03gI9FnrSZrKjfoDH0N/eJiOKT9Pbzoe2j78a3SVtPkDPoN3eYLM/7ARv
lKr9lpUxIdxXgbdYbVkwi4f4ZxQp5j1oUkN954xuN75HXRD7c2w0KRxh4+/a
5/DmfZxB+rhI61XXvJEd3EtyzDfRAxhwho6QcehhQ7WwHs+TcOcW+dz9dINN
T/c9fGPbG1brrd0M7qlC9u9RvaryCRDFfi+jartXRoQQcHI46gH+9rfN+41v
BLZnSFaIoPJPx1BixrQOC1xDi5x8fpWO8FUw1vK7WS2tXg7WwbqFzf/tdr5W
6RH5mpDlezOzxvPRDzZ7boRxTbIn+AC6C+Xg7Z+BbVrLMtR0HKy8WccQaHFf
ZmJF3kQO1eIz36I5UHh2tsCtKyAH8yE68G9h4I6F4WLnRlFQkYthJuleed9C
aOFnxbtjBWiqdwORRfegJ/NcUzVwN6Rnt4zMpGT8O4Gz5o+jBjZe1lmyIzy5
YQV3CEmiDk56cBRsYF1NJ5mkR4s4XczkoNiMnPXaEcQ7c08QE8q71rBK7HRf
5eHtqoXlZxoM1oY+BIzYehK2Ks7EEXkKVUcvia7kfugGxr/V9Ii5B86AP+v6
EpBGK860cITDipE6exBWrX8nTd1TORV8TFkDcXpabFy3bbziWX55gvo7IJM7
zU4gTiNqZ+8lQU8dXN3zzRCAe+SV64o/cTrrmQrIaaAdgxl2AsLHt1SMlRwW
zkV2YvcRYdFX0a8lbyRUcLIHgxzymuAb6Bhkn3rfoKlULNtYzJqnVSf1v40x
K3aFnushxqKXJ1OphQev6jgHW/0T0kz5IEVrfDSBhE7FtLescKwJm49EtMlT
ptkwu2r3DKY0fvMzbUmpI1xpHvSJx1I/Go5kJGvKwOx/NOkRK/Ha0r2lEtDS
DXoTTB7X1G2LxR1/EYG18acQ3x7r5iRzSrpy4pGcds1S6rm7a8S38nOhas9H
nfnI0c+ke6IU9HJXPtfDBpMe5AV3W8pO9dQqo8nC38MBoAG0l04pTWBazqZW
BocxUp3tzEb0wFBYKsQMzjjwTRInP3vlaDmBQridFfsC4nFgcHFETLC4oWE0
Xn0qJHwJpI2R3sZmFK5bB4h2z4ayJrTavcXYX5xQI4Uu5/rJcQhxlhK9fcoT
e5av7zLyBAcB0ZwKlFDlluEYEi0777Br4r9IJcstq81pMOcfEWosS+fu96aW
YS412F07i38mjNnX6vj0H3JAqfqxIduIGSepulpND5x/eQgGXLuiDqPPEaLj
tmJnfrTbE2mcj9dvKXdhvO8I9pi1dpoglpSaVPCKx+odzth1UP1dZsiBNlma
lKcq0uGDBQ6EBv/si/1dSsYb9ic3jJ/t3xzpMjAGgDqwxgz6S47mQsuFz0Dp
P0zarpoVl3QSwhGseDv1A6P6n5mcS4EBkLSxDeNRjDE+S4xqaiErtWiE1z7C
GzghdthhxuTLqavvYIQhXjcliZWzpVKZmCcz3D/jDnWl7Xzwm80ChSpfDIk0
CvKga6swcD4lJSd8MRbGKwwq0E6358762eWjpnzLUqywSW/txXrysJWBHmKw
+Tsn1+SohhUiiXKOKf+XW8tuYVdLF6nlvYN+NGPHhFSN1SviaruQj/+4DE6e
HzphT85EsDzIpJIKtYszlF6hNePf/BgQ/NRTVDWflVDG9ZECvr4pJyD5s5bz
NYnMgdpGTMVIQbApGNimQiOJTEhOgHsaSx89i8tRgWrmcQZXRT7f0Qk0OqkM
aeqljcYjvRAOPBmzWcQV5ADc8fLlvhp4tjd4af/FvG8aRHHZiwosxFCDyFQ9
KeVFlw38R0fscMU8xFShDtBI/ei3j/GO7Qk9NXkYW0RRJv/hcgM/76tiBisM
MxgErtBnYJPLg7BTw4+TnRWWbnXSbLAUuDIvV6peh0eSq9OE7fRQi4WLPFa/
9ZQhLoJx7+/VtuWqsq0RyyWOznEcumy4NXJd0d0lLB50VTfcCYUfv4Mx70hB
dn5JV4hSV0aL30SsaatLQoBbEbfTeSKisjLb77x//oh7fTIHykA03kS+7QiX
LVs/vg8jNqqN95D5Q9ddYpYU5v+5j2KUxfPzP41rk0FDXIuzceNyGSDePuyT
aEh72igtFnpDoidYYINpLR82cgHAUbf4Qh0665KiX4iuSvo6Pr4PyXPfkQFV
fcmG5oH+6urOCMxtIFdqTY7fWiYD9lp3Aw6t2+l52ZGcK6a5JNcG24GjMJbx
4nlkx+wTUEC9/huiBjuW+gB1Z6v5NIZ4/ZNx8026SIjEx3cqlR15zJJIvTko
1SjgkRhLSZfJ3c1ds7nRqAkFlFN7iABS+SjnL6tABoPq2y5fsft7dPDEL6PS
7f1L82NqBFjAPrvRqKrJBnyrIs8CtzkEXRbieq33CValZ+L1lIrFLY8V8QWh
JCUe9Swafqp07nAnAcBGZmIeDKnTl6BDeDZqPIxCRcS6KVLTZFVmNnHD+rar
gMUdLlt6Cr79g04TSnuRPvGPiep9kF1SNcnVuulbzBCe+WBPU7UiHcsAORSy
wvot6lQtgTtSJn8cl5cEWnaxKPXtAwudVcDoiEWg5C3l0JHxIgVzAPeHs7G5
fXr8OHqIlFxObUvrELzptKBZP6SFiiMP32oPMmYWPiJ6W8A5DTwBkWcI6jb3
aweROUTA/WQN4BdrTXXIHOVPaVCaN+nsHC9mOJeox/hgsVfSVawbeieK3CKo
Ojoc4nqfNEg+eoXm/b0soTDh5eJGzMtH4nXa4yLK6jPM2yAHcmx7zdOfb3k1
/W6xfP82spkCriQPqF4zU5clvYONhD+innhezjGAMcJ4NFcBpZnQFhEMplaW
aa7Vd6cQ79ZM1BAgd9e25FC9THAfS/rbv0ZovS4Wf0YtsmbauOBrYCUFe+zT
EnkvCXqyaIG3Knp8+cQSmcHH7leBa25SpC/rfYatMm0nm6roMITxhHS+vUcn
mbC3MA4rKkZPzoeZTswwmUw/jXC0YEJ1urn/FHaZgxarDxyRz1aHhj/844lC
3mn7KK/bsBPEq3CxvC0xP5joZyQF04v6eJAPX5fAMwiEzIkXOeohcQQ352yx
mmG/dC2KqBnIkP3awToXiBkKHAOrzO91HzcLxssyrSR1KNs0gcltdxjP8QNt
ETA2LG5Cv1uribfjsvn3dzr8pfK2p4mq39d6LSM8tjY/+SwhkTdSSghn4JKN
qgtrRlGlDuQO3koX0GJesUxO06SwE3NOyaybUn43ne6EM3v3we+DXZRRcLTM
ltb4RkithYZEg84Mh3KtNJ1nVBS3IIdKAhCCI9LQaNO2pgihhT2sZ9UyFIoj
XdZqVABHr6diE54yQjsyD6vgaBn2+uf8m/uHsm/fwTJIaF+256BWlNinHFfS
+sLxYXbNGZl5VGxRQRM81eoRafnblYL8KhYxQMRtvrjUkYTy4JGDvvSGLn8U
NdMq1IieDkrSjYlaDf4tPBTKy3fQJ/v2oCRJdJQ740UyG616vKiL97DB3aPn
TTMyre1MmjqnjiHcdLXm2bm1/sEG7HwDmqwgTCrTAmhDaGOAqjXaCIlWEzui
roBaIAflWAM1WnfjraV9Zr9kOKYnTpmUSMcphQuPARo/QEjj42eICxl5/cij
yu5RL1OJhCpivoTNOqwvZY3ZIFGQiMCfhKjDueYwm2tSeZ6xC1GV2SW1FAjF
iWlH6eNViRykbScha5QUDj+Q+TVKmFi7O5ayP2iOVSQnWHWrz5aSD3O4xGEe
YavLvZs9UeJlLmX0cpSu8JFtCQ0y1fhgqI8cTkNSybBfBcJBytsABeP5KzVN
60to5vb+RyqtYdaxUKsUVE+Y97+9nq3G83i2EkdZz++tF+Qqr0wDVH/BXB2l
kU8lzTR7PxkbljYlLE7AsfWVr7yEsWpwBmr719C6sJYCBQ+opymHdZvpvLLJ
enx56IVxrQWTMSLtYER1fG2+we7KHp54xfYARoyBEvCNSCj/gWTdEy2z5u2D
fAJnrnJliKJ9QpMG6GX2SQTfUXHmY7rvp0PSPi6GW/Pohf8CtzmCyf58gJjk
iSzo6Ei/wrOB1HCGokiYS2wBIV7dfxYCDcfyl0k0wU0r+jVdSFnl0TuMMV6S
6kweAojc3xrsu8gom3+cK005VfDhnjcjSjSCUsJBnAq7+M391bHAdd1K6Ssj
0U9emsQYCbeFTzCFV/73BVjN3nadP6q9qZxhIIuAJ7+mHzUaIpGoEAEv7ER+
O+rM5qG8xaQDV0dYlKMmiVp7OfW07ghCCJKH6aYV5vP8aJaGDG8/vTZc0Lu/
w2WTommJwFJcy3RrL9qGyrK1R2Iyc3b/kSZxV7R8fv37fsDKQlvKJAgwrDtX
CN4CwawhCYxpWqQ215kA3qQEhcoVgKi5cx8l3M0YmJwvTit1M7us80kskJO/
YA7fT2KrNfbcThkI7afaLzF3cYXgAwAxz/vse6RNMqcxSeCRzKUpSWZoELSB
lcUuUqQ6kaqYGWPbzAj4Ck722cFOS/WJkrjpjr8neo12tg4Q3HKUTfDY5oYw
wP+CzNQst7cORKB0ogUUveVDqXV/gAzDH1Z0W4FnZwNV+eir4XarWcEXKTos
rBYTNR8C9tVy0ixi2mWlMIdGunXGPvQrui95qCuxLOTzYIcLYmn6Hbdvwfj0
DUQ+82TbLIauiyH/j8Kr/kZH+6Xg0W7OQTMhW0/5eGYu9d2aMXE5GpK0arU7
H809AQ4ENngM+EKnY0ODpmrOML9i1wMV23LtkTis0ekLCVafw+II92d8HI0D
BjuuV44s9UeF6quMIGQw0MHu9TCSD4BK4oposE9pY/7eG90TjnngSfXy8D4k
VtLxd2ZQ5yp9C3bMgpewQmChBBNJKWTkiBjJTiXcFTJWPiWkfmusxnhLcl72
dpP0la8zUpdpHHyPTT632n1lHw2RdDAh1jL6uNq9RJ055kuDIEs633X9d1Qn
bHN2blXbAX0UZPKIuujG2tf2mSdGJyrW8a5z30onMl1l80i6qIVlpPevOa0C
cuS73UwGG8jhow+Ta8wwswNICbsoHzB3ksViQ9rKnXQyM7+IwBCpP09ERC+L
++vju1/7XwHrEXJuiHxwez228K54bKLDJi8YN1WFoj2tv79ZBgzPQGPn/Dlm
C5qhzJXaWZPKWcZ6zjAuCn04BGb09UT/2iyTURTaMZkpWz55QhuC1d5sJTr5
fe5G4Okb7JV9VOJCboyuO/SJ29LYiDAonuEZ7bosuglp7uCp/uo2hMR4Wou/
bma3OnswJwQrET4UUO0kpaU4GyoyDa8GCWvYTuo2e+0D812InN/IQZC555CT
5zd9tZl8K7mClWeoH/mQqEDPkG2ynUuBBBcvvYi3GYRAlI7DS6R8Rf4UnBr4
Z2SDOOt+vRj+a2jWrGaUSU3zD003rCRSFkCbXgMGeYOp37xT5WDtgfM7BpTV
7jNCQu1oopj34ct/duzqvM1ft5Ag/rEZ+JZ27pzhWEQpBVneeg7+fqhlwHKT
0JGLyXIbnvdXpMoTpoA6TCsO8eLstjO2/0WrKmIIHCctRgikLOOh0C7C1ADo
f8mxmSA+9slr9fuIehsnolqpBtDzeAp+bfvbQcyCCviJ1X0tI/jEWJsMiqQn
mSuVEvp+4+IYziv/t00mraM7aUdTgQKtLKwGv2vqtXIV5hE992Xz+cT/NFDu
6xzq7EBOZ+xjjq13fulPaKuLoEHax5Qyq8fTA5QtJnle8HitAbxzpASR70h+
jrKHWVxwuPX6sKDk3o0TYbb1o5q2e/VPdRgP84YMRN4z81ojQaIa9CdvegYn
WwcesGhJt5maqETWFFIi92XFKRWs1M934jB0jWDVY4ULwDuIn4Uf+1CGjCwt
KYU57eAsCWryc62sJ+UwW2D7MnN4crSd7Von/pVH7wuvj5z/KpUnXjwc6PG3
WubCi8w2bcklKJ5nOHXbXqk8m/2Q8cBbUoAi0Wyppm2qGO00RzbZYB9AzqcV
56qew7grph8vn3MB9/8mX9jZ9imfpStmyZNO9MI5Fc9U0H48f5mzqj3tdoMi
xfL+/oIlwbiWXQOAOtOZZtPXAg93z3DI2xVer44DBkf8vt+O9gupFdoLRydf
ILET9464cfZKOIi7FIDbPwoL+o5L7uMfJpz/h1MznZmmfBgDxplRYADx2+nX
+EhieAFC2l99SfXTBqdpyih3u60B+7pgMzf5vI9C8R8C7ydnruUhymUtTF5f
GoyLM2SgoJIXe+NtgukNQG+d1wmQ4UsNg2tE5cfPVKO5KZKnw1CAScZ6/FCY
Ao2NKbhPP9OQ6xMiJ96ghGT5CLygXzNy9zoBNz+60+eYNG5Yi+CxDhDzi4z2
GNBx8dX8apMNNuCtqRHYFochnZRkLzf3mnBoYMM0B/2BBw49n/9XKamkNWXL
MAXl052VBEfe3Wp28EMRMJjcvnjanJCONdHBxZbhqVBjpGNF9dMohVkDLSFO
p6mJEaxoYSQr6dNNTRdCh5dVvktbZ+eT7ouXRNUVPoKRgs5Cr0wSAq+kJ9Co
O7zA34tLlWv2+/hf70i/Rw7thGq77dP97hjIioXt6awszAnl08KenqiYikDd
vz3vvCqnCgtn9iEO9owC/EJ6FVXEMIGe1GHC8whJ9Q+jcunmTz7LzdcUPGzn
PBVP7GZWjRrWX2cREsH/Dfk4CxEmuC7b/YzpGDMAR1l36xA1P1flck6bSGji
zTsun4c9zgZev/mCXasuteirDEpR8dYRV+hjDvEoZJScaKX0gScWcOODEFoy
e/qsC7WnfdvwoZMncr2UB91xV0zULw+J1/LyM+jv4g7EPGcOBuB8erKXGvZP
ljFqAtKPeoP7DYvFfmnHEi++1CXQw41jzaXwu9KGYez3gW298ujHUkRajJF1
uWglLBYTZPPEUiIRMctKXUQzW1STO1kCAa1z24qWLVk/gdD94NhD4BDRre78
vesjA0ieb40sFOmuR3BBuQU6y4R/uNtM/LCVrsUl67P+rQQ3zpAU7YVvgUxs
A9wxvYYmDiDXH+UlZaiJ91uAmBAjlCb/b5BVJrjNoHJVFicmP6jZFVTbqeY7
U13OPNQDj0Mxj2jkXLr4PT03+rAzBBcd/4MnmfE2lEq6U1SoltFmDwwCccuD
t/rKgMhsZgDChUUpEbx0aQTx1ykPV/TowvX1XW2SoPghz/GYFJH7gCfptMHF
8u81Ocec4F/Dy6gIO4BtZVaxXQaaujiupam9W3o+aao5OVcIhEZeCImNw8aC
X/wMf0Y9mOGrxiCGh7b4BuR8atsixlTwC/aBK5+k6M8bbK7m/50yzQInVExd
SZWjTSftbekG5zYGXQ/RGWg1jMEDXJjblslUcapGtT0raRNWe1GsRfvMzxY/
xk/XIOyGuukCkNtqvBhN3DUYQM+JBP6A3XGcYIe7omTGs1c9LTXd/UyjLcKQ
5t4ZQnUUqvIrVtcpJbyDEg8JwG7oWEfQv2iZtSBmf2xvV0cv8vdRO5gbd/7T
DR6mjU+Y7aQqRWjkYfv0Wz3V+G9M292go1EZ4vAsVcFUeFcJVzsvPS4ECz7z
wln2DXolpi8BNsKajoAlMf9Ptk6e1exqTl06P9JqohSKV7qGQGqsrPc4AhjX
/JxHPY9JaiTIVj0J2Q0s3rTGX1x+AyDVQtKY8gOMNKDMcjVZGb3Ke4QSvq+p
q2Dc5CulBjYSqfbYWJGW8nIf9XnaA5C5FM7X1Wb6PodxZO0LIyOb24yhuqsZ
UE7KO9b/JBwblOBZJmApNWWeqIfOCP629UufyOLdd4wzE+IiizQsry2gf+77
m/JL9MNf3GkBFLup6MI8m385MtE//T5kGohrdMHDX+Wth3aePIc3YKtanPDF
FxJY9tpqcPmAc/t4b15kglr7B6mmzPErplZsnJLOx93xdhBcLQqkDW9q/acK
rQOonbBmzTmSjrRD6oeo0041kFr+Mdg4RDWunByzI0BXVtQXMh9U+umWqSnP
GvFDYxwpdebBZFGkUHlg0eWmhhtXZV4erqbHgieFddrkmAgHotrjIW07ECsQ
RTEEhtcXqxdDXwXjBIXBlJilp00vzAlk1odKRyBoAvFYb7ZFdhpX7TRBNQU4
aVMuTM09pccmFWa0Cib7USGKp6BtOuZJvw4t+motm3MKC3cU9nRqmDtl/OT2
p6sRPNld05dUyTq4ZTcF6FWUqjORfo0qaZFRtvpHop0cE2QGWrfpvsP9vn93
ny4opKKMIMqSzRkuQ4MEAJzVh+IgO8zN15a3yUhnNonH/qEP0oRlXTn+p5C2
3K0lKg/Z38znvVVMGvqzNwVJmaUdak2yi/92MskGhW0Hi70zhb968Rw4Zcgi
PVntPyC7ZZdK3uX3NJz+/m62cXvxvVCx8ZeKWmevPnYRMZZ9LI/IShgUcIAK
KPHHhvT1qAW5vUJS5fz5YBM/5H7zpqDGMqqWfSZRLxf37uYgx39rdTE3rLBI
Zj5dpFNuaRfjdt+TVYLYAjTMBsC8VGYrNqTFaFNbjjc75eIUvU+HfClIxkvu
Ex2GT6joI+OLdKwhcMI6jBQCYIuY0Hhoa6gp9EhE9Fg0nWed6yQcKsDJsksG
/olil3pZHq1XFF5lZVIxK5Kkn+0MJGqfxYevHRKx3ypcWboQCbZ9qdKS0PKc
LRg/BeQ0OGR3U3G4tq8rt9Ooc+1vYs2Qg6rcfVtG2Ex3YdmdiTxQW8kznyWU
TKhwOQnfugbWWhY7V0ed5Hew/FebnkcyvrjHCVml7nwWMFSdVzNoXVcRu0y8
JODZthh10y38T9QWO2Mrpzz2DIPIKsPDMrB6Ys6RT3mm9KW36vQ9JA5nx8sF
Bm521gvdWcmTCq3cWK3Lq1gYgTTPrgYwz3crUUkp0aFZ0QsaqFNL2LFoxsEd
64u4F3lpRFJ7XAegeeYYx+POt/Bj6kZ4Tpj24czksMGyEAx7o2yyWOqfbKF2
3tYn4Py62cwc+Ub/T+Y6pxmugetZ7pADgS/jTPQE3wHIrOdjySTAihd2Wt9J
dTOt3C00hopj54GO1rCz9JCM689zAWWSjumDhMZuWUfJTRINQEs5T0Ii5BaK
vMns0xgXkA84WxYVWbuJVb6VzZu83ejV9yn+1LGs5d8LlO+4+Tq1pZi+TulM
4H6PzAHoHKV6aTlVGxqrzDR3oXjFus2NxCARQhPfqGeOzU7eFZXxYlUyVhBm
x1CYoDkK+Vfx2mIqWZEfAwtO9g2Ht9sQtQCt1ugwWYIpDD70QFO8ZCoHT962
tPoJkawpf71BlaR9LSPYGfs7eO/WjIVfLB24GCVcRM/Yph77Oz0MB3f4G8aR
Dj9vPa+ITqwx1IeGtsmN3f4zdWLjHUvVtoT3wvh/8l6oMA1FrA1Oz5KhUBoi
mPAzsnepD3tJpameViKmS4jc5MPduaEQSdwXiD9bYP0TPg3CQz5ILx/VE6E/
u3on+R5AYXSNqSkUA0JjXOcB5xmScAVR16NucleTLTuQULPHh/NP2FpfuNH1
bnK7DoBfWurRIOG21gRK8Xh4Ch0eN54DC/zxgJh4cIVfP8IVDWTwCKbOZhJO
zh2oAAdGUirnTm71y22m1jrf9KJvzTLja2KNu0UWmiwLcfMAbKhM7fBekguf
yFezur/Eqo1RrkX9wRREBM9PoXpJCr2E1lNmSXHi6XADAGFVybe/Kgrdqh5i
ArWf0yzxs5jMD6M9SjaXjsbN204h6uYeF6ft1nb3X3NsIiFLk+kwtRS0V+s4
mVGvt4USwjh9j9U1jAjO8/kc3O1LFTZwC2EB6XxF1MyEAiSeEjOMNbszRCyJ
prZp9TU4FTVU6r8Sg6heeJL89Bpwm0tcRL0VpkLsroqgqBmaFKNd66GETGNe
mgcO29mk+feAaJHcjGxIOBSS8mll/64X1FA2xUiwCWTcQcKtGbCLM03QCpUr
K7RDcUbwpanqiX/Bo9voJBdclzjg1dBegfCSt2G7FMjap9V5NorPbT9Saj/P
pcxrujD8XNHmKtJKwRoemTUxtkq4bdZa9XGKuDSwkko97Wie6pXagrh4WQ5W
/YhZyBPthzJOws9LX/pxPArXp5NGiAcR0DpSQRrUyqzQKJPlhy9rptBFnu8j
H0YYi0xPPJTqyi8Ze1OzOEzROfWWCs5wREyexaL2qGP9M5K1J4SpipwHaoqL
LtGyP+shndfbIkPExzG54Rqucz7GdkVHXz1/QH3UwLgiBFawCoCMq9gwqqXe
Jx1nP2YEigEVpuYRuA1DYbW/RziNkYhOM/e4f27AFiXYnddRtErnMfU/1RGj
qQhRRADx4J9zfvNItu6V3ti8b9OzzELvDi+a/SLv4vLx1og/nNXUyGx5oFW+
KSurIYfumDGXkZ0JnAjt9zyw4j/L/0Twl+b7fU7/gjFJkwCHmyWjnWYDC+EU
Gobo5Wj1UJpfOxc+yuEut6mq4LxstEW0K1ljn9m2PsPqqNEvtOpbMF+V02yp
6BQMNLC0HPDm2pFGa5LuN9/Bmu1QdTnSjQJ0DXt0pGbdV8hq38PW2C5UZZ/S
xQoliN1PreqH3BnQfEoxo5gRi+nMBxdFgwrmTC8y2zduUtJpAkWwbJEoT7KA
MqN9gMsTJ92v6N4HwGEPjoBid+5/RzCUQL5Vg1/LUr68eM/fk2yohLhWpQkg
yo6oqH/NnZfd8fa7IYrL5KdxzJ2/yrt8/3CAYfPiL9zvoaayO9DNBmvnR6UQ
m6li16K6z4qqvEAng7glHPn3YpIdQtqPVE6Sj0K1Bfn/Mvgx0Z3ORzYUHbkm
tqJSpPsWJ/C4k2931xLN6HiHNeAYjo5A3jolewMA50B9teea/KempLUlzzr4
hhIGpUnLKQK41aphyIRtQbQV040pOqWAnN1qVhAT/w8wB0dLHtsx3J6DOaya
BC35ljX+LSAx+mmBSNoz30hz0v25fWyQoTKbsb/4YdW1azKhYAgnvs7/v4n2
cHhW8JsFzzMgMthS4gOVsY7pdEwSEgsGzDZOxrEDbIzuvGvB7kJh+/KQdG/x
XuCZFmDo2X9qgcVqzBBhBzaCngCc7KopPOjq4GDcdSK8M3VY6iKALQgTWLvF
/Cs8XxzxPy2xF7qut4rv6XhxCxOVBDi33x2oKJpmJ6M54zVM+oWIDt9sO+v1
dWDjm43WVVQYWx+DFHz7JxGufqzLjf4BjijhSpjCf76PBRXIpYWbzStVyqQ0
NaXD7asn26czY3gyfY/9sZv6rN9o4YwuzYO/h0sw1ilxL3Z90UQyBQ0ymOWp
FZStiyw4VXTrTDLkG3TL9EpCAZlcWHf+rcB8TPrvLTAu64BEBWT7hxsSaDHN
5LBqEj6Y6ea6JPC9XU9ev+D8tAZcF3cI2ayNY9K0i+SFoeo6567NvclMJzqX
51kcCTYbn7NT767gmVx595jN/h+oA1v87kcqBkmO5WdX75xs/9c8mOZQeMmc
MNvqyUcG5YoA6eiTemMZKXCVyU5DUCDWz1yDofq44k0PioJqwLd7BQj13EhT
6SmWk7QMXJIDoboVWRkliZNqt5r7gWan9i74gmRWUiP4s8Pk2tmVIOBYD38h
wBn2vhgRAZyaPNMJsVlAygLHHkrK0g0LJ2ZIc6uQdoyBNBuowbiVKhzF9NS7
DUzMHL3tWM+QPX/ugkUMZ9s8WvUMTsheWu8q2O7U2nuZlFjaCnLQ1CkW/43n
jahJeBz0d5/kReWjcSELKvbWOPvHuAQmbY/AUjGoL8bKP5TmJSnTpXhNRXAV
+F4uIqVlIgEkhA6srpypzIHkKk4uiFjJgGFiQOqtGVauFkES8WXXeU41Hvk2
P+hwcNmRzVXIBRX1C1nGFc2ohIOFzqu+6tnWJ0ctpcmua17qpff++S4B+QIM
h9sspUIWpq3lJmr79nnQQKG5VySECDAdYI0GOOGnfD+ITyzuBZGctuZBLU44
CBqpVTpHjqzvF29syXylOtndnapnn//+xsraraXtWXF7nRswsUpXIwcBBiT+
wIBs3xZamLcO1/qRrOs8l5EolT3WAPrFDy+OdURnghU5EtElJlFyICZBi5rt
zSODkBQM3CrfgWOmjZS5765WkMIrrdDglMuRSydXPQM/AFfaKRnqlpXP3ugf
prfw5jQcG+0djLRkP/IGFZUkDqXyRZBCjUMXT+I8RksH0qiqYDKc5RxdwjId
AzkIS0doAr3ZoHb3IaEAJcEuQQ+vsR713n/5EjvhvfnHxhOmpheRu333EVqD
RRWxQjKdvVbghb9Bcc55ns9pxKxCvCP+9LH/SI2YAoLvk2FfM4mkaY79rXJX
3w+/Ho6PTnRb/D1fTXSjI6v9DGFBu15LLK7gi1uIHB12Cv5b23522Jg5Y5e8
Tc6SHvpKM76nz+iipIEuE6nqe/Mo27yA1KB8VPsg9Q050UPKs2JtZ310lqWg
E80JtF5tM3U/0o2aI0AH9Wc1IVE9PjW0bt9ertQ5SdxVr9JvYxRuGv3fzGl7
nCzb2JRjhRvC5Od+X/1TcLfieL2GB6CbicxhlUedrIFn75mC6wxfeDL57CHQ
nqWSPBH3eSMaMYM54JQ3ibsQO9Pn8xY6uI0PaQgBW3PNxqzOvruqRYExw0Vb
qaeVDmqO2zj7kAsb8DrcgFQ06Z04GuHcfq4ewz2q16nWpwzBQpUtAJ6GcuIv
QCobkpfNHIZaNXe5IBUW+oNqmZdeZCFOh6ACN3jQUMaOeskdWwDXF+LY3Lup
vyOQvoCL8mU67QA03Nw9rM0BDOX8CIXy1tD/6pVc8Uk7QunLoCBetXCfT0z0
P+oyx0TwFY9xawKq6Xp34ymEKMRqRRpEFgzPLFXBwttboxPt5mh1TeTT0l8T
quhuqMqkaOpz4p4/nSaQuqZg9MwXlYjvZwNtXcO4NZ1NO67Bh5B/SzuKHFEM
8dpPMTU9gN5ViZ19Zjl+bAMvLAfIp/NOW3ZNh86MR+EzjYOoP3eJJiIW2X0/
NmlI/1dbbgfg3NWcWh9aXh/CCm9n+PkBgebigCW0TkZMs5Ys2EYAZptI5jER
TnqOCMSzaMcl6j7YgMbFXxyczen2xQTqwOWJ83fusX7VK2w+MzQuxHLrl4SO
iy5654Mss1Wzw7ADJ5kHjMynzIzzJF5ocyxWI0NsG5Fws+UIlcBS9G5tm1jr
5AwNCXdidnQ0J2KcyRAKOkGGylh7qcbNj/xF9vJG6I9oQUDNH5Rr+3FxGkiJ
2/cgB1ICF5889ponVwSla8EsZEg/AAJ44aQnHlnIwb7KqbF4eX08B5p1rb75
Z9YXws3Dbr3/sePSnxlIiy8sJS05mMeN4zkWoCvmMzGU+ppPwnldY1aAnFrY
ejoJCiqusC8mjr0p0JIYJcva4iQA/CLljjFmjMHLKGBMZ6AjAFWQPKw2x/NF
opjHKxG+oRK9NlTJ+fK5F8fXvYa7KHM6Rkw5GO7Hnebcmvc9uQMTL8AzRWlo
YL6esqIaRVzD7+P0REHN3nzUSXi/LlPqFeMznDVaiNk+P5DqdNfILkSpTkni
sYBikBfGQE/omJc9SNYe5eSXcsdL0gJEdUaFhUVg39pBBxA3lhMcMoxxhEF9
kPiE5BCJvpmFC6VDU+41D7jA52d/aGmjmQbJeCjQYl8khZxNspgY7aRV+01M
XwM+jscQQpsdibGACMDNn/SexDuXbWKRGn82RlgK9HkjPJP/YpAwYLTze52P
6rVhlV3xucCfDoPMmR5N983ZWv2xzP7WkyvCP+VI4v4ysIFoPNKpIO5aBk/d
GW7UcWaSiHAufOm6a0hnMPpAy0hcZAHLOEHRh/4hqpVrdN30iZ9bAjr74fdJ
hT8S5/ay4IW2ONsr4OW0gXKpY8q6fow/Bmmh22gVZDbypDReB9TBwZj0zKEd
PtrxUHNDHZxdqxE7MDs+sMmoUooCOibz2DdKo+Wa8I6naitVwoqCYA49RYTr
yMlBLLRu+odjIYZS+4wBB5ODr0nRvrpBqFJyv9qES2aJyS5HZ0A/utM0RIF2
xVSILRt58IMXGnOOZ091e91Vx+rwPGO4TkXY/Itz9yKzEl91EIVhNOvqBFbZ
02/ltPgIabkSTbttrKNAWcICLUGY5/mlhu9iG9zAnoIQXG1As7sXfmUdtZGy
pgZPYh3MQC5mN/AUpPVS2zKbEfwHw5huDMwnW0/69KdctO/zTmOdkwFB7Zj+
0Gifwks4wcV1rsnMMYM9kGxoj1RVLeKkRihe2n0SH83TVka1wcXmGSIH37p9
96XN3zXAwypVSQQgsbCCroTaNy/chSrQN6WZfWX9SWHF8kpF3IS5vrkejFWz
68iI7N+EnL+Zq24ET+wcp1rVFU3ItOcLXsp58oqVOV4kkg6WurDlBMwLLzVp
NPBweOM7VKYTTDHee0dzRMpGeA5fPM3C6B8P1nKYW8kD7dm0rt4cjK1QQ0Ip
SaVcYTm6T2tSK4nZPQ3O7/eAw+0fTgep23mvER9ufbj9+qXmV6rEFSSM8jHU
JMvrLOGHb3MXO1L/oNFxJJWc1Ytp+ixy18s76U2wbwkqA5S3wM594+ldFSCn
ua6iqluSsOYGEWu/zEK5DAMAyuxsPaouC7dVhzwOf9QBYBSN7cxm0pHq89g6
2tqs6F43my5BP/5GCGSH8J4AAG28JLmlqI+rpRoQPEy72h2yXpclOsdhPLyN
jg02nxG1Ci7PRX6BtRUq+gkJFEIf0c7AWBx2dhn6AAacCPoFLFC2R2kRKJTp
SpwO4R4ZDbTJudMVQYbNkOkupcAv7KW2fqfEzdEwCOhOifyTz9mCnkCTOuJ0
kitu943GKcSQb1SO/FNphsl2wGo6TXk8F2DAcgwVbpYZf9uURxfRn8fBRNiN
aYfEIwMUc+kU5x9RG105o4oFfahIKbxmwP4zswS72v72JQTAEJ0bw/pCTdPT
jqJ8YqoYwha4mWz9TMEEHXvz1Xgtax/y6MMCAnCpcokFQANkogGUGff9Xsxd
tTvJxjDw7KkXildFoHBe2Un2WBzTMydf6aWe6RuWWZ9gSu/MCwwRzwTo+Hzq
zCfXVX8FqER4v+Tzeww5QzHgUqPszVm4q+XLIPzYfctwoTI7O67AFBSoXIpe
cuoGByf5Bk2m3ALjjuzaSOM0lRWNmyfvx3BnWRWhg4m47hoxC8afJKjpusuW
rEzsCNpeiHTYMvGsz4n6yyq8fYFuc5Cg+1C+9lncUJFp1ZawCxBkK/wS4F5y
+GWxb8TZC/fDqC8KCiNe4GUWaElTeqxOOunwPlyL/8lbkjVGya8/VjlOPqPv
eYeLfeI/R1nKZjj1k580iN1/htVqzhJA9Dn1wxacCJtMCPuHTqIOIB+2pJRb
9AYJqB6WbC52SzwID/ohM0xIdI/guc4feAkXyerN8wdXbyDC7ylWGiC4DIIq
PT7xgW19/l76ptAaejb1W0Oa4RxyI4LmzWy9KULnW6ZnQyz89A2KME3nCjen
kFj6QSQGk0R1d4jpyqcw1IY6FcmPpw35P+rLo52pQTivxI8W7MqDF5nh8G6D
cfEuBQUl3FjizEi8BZQ/T0QhWN4ADfJIRwFzwtgpQ+fLSS3XHk5kJ7132IF6
ry1U7ub1kVmXvwFAhg10+DC4jaR9gvIjtgjlfD/48qGdCScXwsjvun+6QNBK
K8VlQoQZjhLFg0qO53Zs0CVA4ypsJ2i0GLEvGSkzl33hQMhQ/nIl83ngHEJy
PRrRmzRZsqcA+PoGoxDHgtMS6JgwVyjM7fqVpXkJEIokaXeiEG2G2dAFJj0h
A16eARdCXvwd+/EVz+WOAGrlYoAVQv0i63DNLGRS2rXnM23zDlDaZDGIUpzk
MlfhbMbTR8OX2i0KqYDnw3dXWVu2J3Nk1BD6/w3oCz018E+Crzm3gKXAl/E0
MEDJXZ12XvQODLtBWxtU9yikHlPmkWczBhXCJ5fX2H4gI5ovaaCazO5oR+JE
V5siqGXOaIaW1gXqyMK+vcQhOk726dJxzm71VWTe502W5sK2R45eSk28BQen
vN+DGSN6eojI0vAvWZDMzITOuduVUUw9fw2Bk483J6hA7Q5kwg7N+HAKIWqH
6/6aKiUo1pgca4R9hAGqoX0tqfJAZKz7Won0x6GPnKq6LtMZiOzlBsG9ybOn
Tjo9PmH5dkouP6qgfoAGlIFN2BTJt6JwptUlmxasYIaqJ8Il3dp+UFQei9Oq
Vijp9bGHy5W4ZrokMjLjo7oDqFXhjCv1qwutWGQXC0LcS+JK6JsGKROUYw4c
UGUBGNiei1N51lVroqWuek3jBatA+MuX289/MYsg+ovM3640Dju7DdeXQvYi
crovmNlJLb68aWKhKUYHHvPQEMUdIItVf8L6uhDJoEAjUuAEdre8eOWyadgE
SAVEAdMSzIYaph9PtWS4309yJufRin1PBtgzW5hNbltIqbY4wG6EwyP5g8Hk
97uIUoZos/uarkE4FSWUC5wdD2wueeraB3F2hyI5LX1aR6tHsGIdnx47wm8+
mZ9Jr3BZBwAIoW9P3Q4KVSBYbaoX9Z7NSwhtUsG0lFAz/wPyZ+0+yUOBnB4V
aYChA4GVo6GIiQKkxHdosbtuHWt47muk4Kx5v8sFpLQwbg2i8WjxM/3R/nb6
xsc4GKwkPCiEhpAY4CyXLgMPnBNb6HrRJLhwDVr2wjmA51iQLoB0WqtL/cnq
31eAaAreKUbEbHO013JSYsk0vdmpytY0qDgVilBfe9ycS5det3ze1Z0Go7AA
IQHMYVR18153kyaQiQWJ7642hTeKFN91G+Z3eSKVj/BT0UannJQJroD79szC
QwIKitas/cmJfcv81unUU5HmY6Rq/mNcQxHQywqhfEHzZtaZyf5mUVsWRUR3
Q9urGfy+xYt5BGBLiYqZe/i1p6LYVyhPiSWuN2BZt8qP5TsPSBO7kCcHSUzX
FkNaFkqSCHS0D/RGbUhDcU0d+lI4qQniir1heU4vzuDIPGwi5iISD5LQrPze
6hOS+zHDRN2NKVjoXNPOR77VYLeeKEi5yU77/tBPdX8U0mLhP1ctPvnDtdwT
StvkE04n/R0XBUJJJvbolOB114Akam9DxfeS6wnTfHa4OiGwYx5O0ZUEi3i7
tStpIT0j4FhRI3+4h5sKXWDzR4Bn6Xqm41rOMEIhWmXZyXFoII4c3F6+aVE9
CHDcdZ9bHQgzHzceduWZA3ITcka7Sf1DKbjYIi9nnJ28gh84bU+uQ61tW+4K
lnAA9CieOyX0homUfDb3qrrSAXlcI1bLGWstO3mGP7XVqksy9lR/hrS2tCxj
wCVo50srvLZSDSQbSjWik2hNFENMNi7af/TDsbeb9fZ+4c/ePQLhqWSVhWP0
hXCJ6rJOYjIX2jXpA5UaaZ1vKfftvSucUX3owKkYRGhvyndUIWAltUr3rF5a
0BBYf8pPrMqvteXLu/e8XCl6NoIBJxyHrlA+uTwEVfiW79Ra0UnU+6mStPDp
xLcAf5DPqE7WrdB691xe/MhG77ZetAVcPoBj+15hBIgWaJDJD9crHJgF2V3O
Yee1D4QT8JsEgqGnkpsPsmbcBhqSqF5ZaQnZjuvzHvbl6hrOG10x/aW87xEM
KCa3iGXwIvZLoGGLsYlLzp/WoeWL8JxHssHl/GFQ8jbGZoLeb4JDELwo8Hgc
ki9JZRdMhjWOkh/uEZ/+CrXVOnx96d25Tr2lhxTc9acXRgH+DnuU6axs/ZP2
KJcehJGtFZdlF8VM9EiggNjDDOLOzf6toxrCfe3Z2JaMeQK09dA9UhWyJMJB
w7zPMhnyhhfvSb0TOePvbno4u0YHLhZZd+8KaK1Egg0Zp0gDrpqY4voc7GT7
3TC4Pwhirp2XTNySi1eiBMxW3T06lM1lxRIy4ax7SEuDoGOmLUkkiPxZTOvS
O3W355QHweuAqTx1k/SpKgWpM7DeyGWwm13v8ss/1upkiLx/LQUP+kB2AP1k
oek7Ck9ltJt72RQn+9nyND+QGaGgazhzSstfP2mPE25mfIdCLw75Y3VRmo40
M/Hbet2xifEZOwgMvf39i1uEs/ddYlyqM9OqNydeCnkjSmu8r9wXdk3TIIq3
oPreVsq+PItrutMc6jDZnR7A7t7eNnDQXaQmHa6IFsQwGExezUigQutyNasx
fJCaOXBJKO/WrwIKlpkCpq3DVuuIKU/vbr5uAuLCKF9A1Nv2mnBenkms6dUh
MY4Ga7loUojQJ+w0l8vK+wrpmDbaDK9Sq6AxuX9hrpOPu6ieKS8ddmWEN0MN
PGTMZ08Qswq6iPy0lhW1oxMNL9ohSmtVxkzIDBVPPYRA7G+9fLVx39jEE7/A
cX5VY1RQiEY2knCz+J8sQwsC2tVFNjIboxR4ro7ykqnKkOCAxccwcd2UkcKw
RSueZGdJots7mqkaIs1FHw3xtUQ12DhLBXALdOOOvS1wjX6HgB4EBjxBCyp/
2lBQmshospT1/SGXePjNDuqohXIJtx8kcJnSQNneJoGdxXjMgHGLQkIiL4du
DKWjBeP+yWznEqBDlu9OYgHSB8TIMKx85BsKzCL28wkISBHISl7bs1FPMgvt
7beb7N3djoQgPvF99/NSP9xFyMedFvHQlqSGBnEkd6KF0CAPVcfQ/K7XgekY
Riz18YGiWuuRQsqqW5g9SIM7/k1Tg1c3NIHfMQ6w62ZnWXDlX18bRGQ+x+zG
VXSCwW4Dp+ULlttkXU3zR56vGFlMBDeuI8nbmzaFeUhblgxP6zo+lQYne3hD
QC2LAul1BhqlcHM+i77wSFplG+PRYGhABnMJIaB6iTBcU4I8i0RwoSxiQ0q8
nPiq1YIk/cCTwX8PJY11RVr0/S05cyF9bRHJtHxElH8pCHI7T+iOQzJsvCEZ
HD/tyV5ZzW7Z3QA+vqUY7tooaf/s5CNR2bWB5u7MNPVs1W/WVy9fMYBz6iJu
+p7TgQGm0jXLxb51STusIOGJAKMo4uVjeIdARNJXgF6tMq4QNrRIjYfqdN0m
PdxYK8NoY4MGXBo+Lep4RFTUCyW022vqOGJu4sCAeU3PRmfElMnF2Yv2s9RN
KJ39WhOro+TgtCNGGz6EHNomBVaDt48lBRi7j6Mef9fAL84tK+W9faWF6k0E
oZ2Zka4Sp/TpRxICcgReubfEKTAplIuyEi7Z5qpaPS5aYohnkwwOAFgpouyH
G3dp+isojS2K9VwbBzCP0XTbjsNca7mcg0/Pejy67ZiOwNfSCFhVRxM5yA8k
ibCiVrju7rmg6PwHLgldxX4fmNEm2BbLlE+TOD3EXfvrw43gy7XBt18D2q+a
JrLCtUbg3u0uAarHMvFBujRZgWp9cL4hSgrHKtQ+gOmgGRHYLVKPBgLajgp0
iqvC+BvAlgQEZQlCdO0XPV7G9UpjHUUwrmPBWV+9Mz0a86OF360h0aWooB4F
o5Dq0ZBHPwhThyLXT0pzDRSg7CVmcLkpcUq5CioLv2mg9wy3G3o0blexXbbn
wr4eyQXi0aSbaXZultJvFzga2V/kGc3nbq8Yb2THxza/YoFP2jYNcSTIj6by
td6cmf87XMqatnK4qAbLcZ/y2499bXJ86ePdZyJozzogOPcNvIi198ql/8Zs
VHRYcnCHhwbPdQiu+9r3QYjUJKOelapDZ5rMvsu48vCfliGtITaVFWorpNje
R05fejH2LckN5HChNjThCXpYhIrRwJ3Et/ecxwI5pQl6uu6t4qTbloeUWvx2
U/vDhAVEOE/KeDGaVjdTOvUx/LOnu4mwoneZFhS80xVdi1I76dTmaGeSwkiN
UGmES6xPDeB+9//VO2GN+woyb5tAEjl2whgJ2L3otmOM5/Qi+xSZC6M8YtLK
BT5O2qr0gNZvgBBGutvmEwyL6ioXmBKgJrC2Yc3KEyz+lcHGqiwrgr9+Mny7
brqBfdeqZlju9bcqsxMMumFiTLpLMrOuoWg6oeuaC4xNKDjk7jsE4AM+TwbX
mOMRr/sYW2VZy5W6s6H2jAphio0WX8EQYBo247wonRslQlXovJzHojGCYSw1
YDce9ALJQVBvzltHttQ8560+QpM8WmhMHdQMFWCt76jSVzuA0PrY3qDVDAY2
GKoC35hqAgNSkqnP4ia+RWiES1qrHar0SAd+Rsi2Ma8k4G3at/MDFwNyPz87
NsiAfceK/bMNXyaUb7HofiRRm90b0niLlA82wCGuwLqc9YbXzMHZnOPE34cf
AGSL0EtmJJ/c0aeRZGIGJNYtFD7IKL3z3RnsyWpyQNnE3Ve4sznLPxm0xCHd
4bdJyujy/hnDR0KQF8Bg1gcnV5NLdbpbpRe7DiyFLmF7jVb8spF7PsiJUxrN
S2rO6N+ocfdyel1j3USrXS0toYvvwB9a30Php6biQhjiKv7yZY5GkQ6zIRew
jEG7ynZd4kxtHFUdD6Gvllw/tNokkJlv91LxQGQ7FeZ3coFW4pYcuL1fD07S
U1J0Ejh05DF3btlqSnFWbBpBjrPEJNt+FiYGfuxnsGDFzJeFRjzA8wszMAGs
hUe5iveQBXRh3BvF+/nUOQhAbEGDxmRRDEtq7jcI6GdjX2DiYnRFdIodsmT+
LKmC2q/6wgHty09ZFaxKwW98eZW81Ztp39G5ULdlupvJFPTE06ri6QC7mEXR
KdwPi29zMQG2w4bfKPyJ2mWMhOJBqZYEsfwsYjCkMvCmqc+OqDfDEURI0cKc
uuUxQM+XghdFNm5ezRFO5S3Dc94Db8IiXiPW+zC7hsdYHVFPhC2VLi1yF1tG
m320UIHSfMAJUSYZF+Z8MrMFcWZp295c8x5lZkQXVqn6r+4xCXPhnDy4ZtvS
eNXehAYmcaqfq7ErMlgZdBkl8BYCvmOdVBIiP5LdylJPHJNB1nYPuCR0vkR7
s2CAiJn8yVu8B9VLXKAriD++B0cmrTcfCkeIIhnZGWTgOKMBiFVh/9dP+ln2
lpD2p+zMftIcAdp+6kAZOn5FvITGJLn2Oz9muRs6myhqUHTR9ySH/eglE2Lo
dNFEIQy0mxTa+lq1R9paqcbcVqlA8mRVrogCTVfPofiVDqZ0Fgb7VfCsYh++
8310//W7b2ufXaSq2dA4Ul7KGvN5QEctNLVivJ0/Mf78KQtNlgF82Z+vr6IM
RC668cpMuudKM68rAiFwV+QRTh9g81sdKFVPKqHEm00RmA/5tlG0Di6nHvfW
cWIzLhudIZSVWRfHjf2LVDMN6g1ns+igYnksILlc/oTKuoVtDoUJoDDp20fb
HSlm2dW8NLZH3WcSKrv9eAc6M0BepJY0iuf50KvZq4e2/c926CLdTSD6OaHY
JB4nQ96uFY4BiQyIDtVwiFgHpgAxHAWLXd9alQGGkbmibEFC2Cl7hD9Yfrhq
GeXNJnBN+9m4xgQPiS9p7cER6f1qLMk795Vq846s4eVfqbAFR79VV3F4nV3l
Ctb0e4ATYiO0XWluP1uHJ6P+YgL4q7541LazrvX+0j+80GPXLASF6sexIvtO
YnPiZgdPCulJ9xzt2VpY5SlxM5nhYyoKHIBhv4NPw1M7KNvCAQDu25l0mg3S
bezRTRwcpa8VUbv7gMxK5ZfKPoPKV4L8xtMbz7ChWa5iOvTynD0JDwPVW3xX
2tGzYhMDyRJ0/cGskRUrp+sQLlGZKPECu98qadqZQeGADciux8HNW94BQIF9
AF+eHw/dfE8MYghHywdtXi8gwB5Zo1LNzQF/TwUyDXaIdQsmqnPiUsEAs1az
xOUOD3qe8YgwchkdnSzNx6tUyiSD31iavWG2skVVSLQqLH+XmXhDXdXM3MCz
T0yfPC+rpzDlrGzOfZossXtlUB4DhG4djLnCmbgqXU0Fr5UP5ki4xl1z94gf
6jrSvacgCA87810J+mhz08n3BT9F0DPXOwu9CIiKNdxKRRlcIN9WYK+jfdLa
auoQcXTEBq48kMMQAQOEhuf/2qS073yUUlpP4xJhQIg7dksiTCNgV89u78n0
nIiaDZLknnryz8YEhbbZn8HQI2CZkZeJQmVCto1YhtRNKlvMJ7RxOp/hA0si
urLnwTTkQVFoi2Ru+WGX0U9S2S68MrSAcWxjiaOUHMdtOYnHFuIspKowo5aF
hqtv95Dn+Mbh38x/AS99V/Ioi5MLc13rKQnaUXj92q3Pjja4cyC3VizPe6iq
5b5km6lO22SPlu8ElcFRviU98+sXYOhhCPZV8YgRfuYNAGzTb1U3DMW/1pFT
/DRZR4INmLoEj3CpqTkSzzqu+/P78VyprAKroL6x9jpPbf9xf96OkogCWN5g
qZscdU4XmiqbjjOtrq2jWhj5gt/kqv24gAeMC6PG4WW4m+TG6y5GClIWciUt
0Gtn8iFbB8xN/aYBVja0LuEORnrXrmq6WZ5a+38dSARNbdJyFYRdkcnDUmHr
HtWH4jjsCEDxFhyrqdJvaoGPJgJDIQRp+64e5SJDBXXBUByTbXXWoup7MLR1
w2A6m6HnoqhR4tvwykTXPRwsm1dEiM35+UWltiV9iPNNSgyVf7Cdu04cVRCY
thlRFlJfkaUK2SknVLqSd/jhacmE1kFhL6ubApNUX5n9Ww7M0gEPPYudOIlq
5UfT5/eCctQbSTO4zRpZcPYxYCJOcCfrVvFgjkoCUPdgqDuJ/mYGmD+v2hqd
xkhevspxfMmbM5fPiGGR2gCwOKRNIDmgS0T7kHNG39C3u2uO5Xmr6T91ZgjL
SCJ/+Uln3WUb5W69tAQ9c9eeAyJ6NWfcXcrjRbgiUq7+tKZSMDcDqUaRnw46
Z4UgOYZPeLHF3SROXbEQ1u9eWKWQVwX/hEed+6Jp8PU+Np16ma9doZrRbCRX
s+LpUS0lR8vLWR2eO8FtZ1vHAQSB2CT0aSLrVCO9ZIlbTbkQd9Mk7SajtFJ0
/oY0M0bei/UNVdD9l54SD7lA3GuVzlMDB3qC0kfhKYNkHcU4BQ90cui8dUlZ
GUgmniV21rucmmiR2jL5udTTN3x5W1ZD2dekbmfKFhyykae+DJPd2IZzpv/W
Kq6QwUpXT5FgZrU8NK1/0HzzyQYYQR3BNRvaIdCqkVSs3wQ0D9y/Mhdk6Cnr
lon2lPaujCsxw4gMtoYiu+06kAWUJnKcRcHCk2ayt92N8UMXGBSjd/+dAQEZ
Jmrc6l/9NkztnaPLa7gxe9VtwbLoklKBN5P5YJ1UHTHHhWFuqjsPCvP95wfh
PF5nvBDr3J2NSW2CWHYJdjGH2BqccCR+1Lk+GHRfrucQesgrpoNei4Wr9zdX
B+5DcoI7IFhiBYhFe6fOuAvcKRgG/12aJ1ODR1aeBhYQPjhnXgG/ZUoCQTO6
HZMTYy4BQBbbPiew2ZeJ1OHVKHDwgag22AlX/xtyGnVu8tUgQgMQ8ZAOqYOq
EcHOeuDS6IEMqOzgPaXPuUoPNySCTBRBUYL5m1k+6HKwlMu95Uu3/95eRNMI
qiZcLNSVvE6gb9IovMlXVu9uhfCkIu0JwFIxSKKk48p5MYiuYCvZPQf7O5YF
79A7YQ9RQezNV6BWReJmciX6YLgdkmZZ1aoak4txfzRaBg/V9ZrN+s49NB5K
jQsOV+ieEE9rQfl0B6WISVc4OjbaAqMV4kVZGaEv6jzpPdj7JVRsNotyxqgY
Wsr8KQW87wclesfEbuItDyPMvQV759njU6LOgG/uzRe4CaooImCULrUYJd9d
bZeTNdstmmsMbCd+TYV+Gm0iGuCdetdUbADq6OvI+nBGUoWiSvuu5e5H9rgd
22jfT/G0Z9jqqAfisZ7bDgE+ublIr5GEyrLFX5H0bd5ZLNq6bfl+2qVrHCg7
Sd09sX/gF2i2I9T64rmQiihPXFy1Xq30s7WuXz1UU6lDiYF026xcLU0uwpHP
DnaVcTHhu83kVEhwoYdLQnglKI0RUR4kY8doRmdWxDTw2Vkrcl9cEdF4GxF3
0PBkpsnUr54QksNSYvLczzom0Ed/ZPiN++vPXaX5aWGvQ/3ge1ho2dvgibQT
1GlXgud5Ss9pFyzzQblvjicU4Kddeoo+NdARGhTzz+oNkEqrukJTXzJouQ//
WoQyVP6x+SB/x9ligXwRB/+9ngHiaBWVwmh27fWkDrFYnhnZZ1gnJZzsfqcr
ejZoQ8ahtNIAwet+pUmYMp+n8UJaCaipM9Hduz0E+N5sUoI39EpR358UlK6u
7+z0f8lHv1XMlezQcqfts1Q+wx1nTBYKvjHQbbgxPJWSXW+YuOWDdWE1SQ7m
28N7ljUuqFDn0QBVU1fkvSEW2pEgDguUax831q4nmvSIruxNlhSGH2q65kfX
UNhECNXx4wYQBN9dguVHmFBeJNe0cXQMDoHdYudHD2KbofiI1GyORHCgcodE
GWDCzr9BVKPNs7ipXK9O4bIsCExoTigUD3e1H0mMpCFdXtFKYDvtfkd2gW1Q
7TK/5Kz3xUwEmuVVplwPn+zBH15z+kxLQD/setC2BUGm6ag/xrH9xBARJdxm
TP7ceZz8e4VIPaEKgyE0YV9m+X1jqpydpZ6Xn+LBmcYf4e6+zcjRcqshSdRq
YZwHipRDgQXxIEcHdAY8ajXzsy3Unxj2w2Aw8e8mzXzTuriMTi4oYqrBTsK4
SxwO2oJspIWSEj73A59mhah6pJP/D+1hwWMO4Lc/GTg9Ll0Xjkr4899WdRoJ
m1o3zSyCD0e6zVhwSGepGpHmjxFGsHZSxVtcJcwgYREewaJilWwM5poGHkxm
MZDDRLYKU0XgufwUZrtflNvwylghaTK7n4uRkHlaJrmevPwKceDj6IAYWb73
loYkZFqVL6htUUml9isQLZc48OS97YL730qFB8HC+BPyRdO0sOIwO70DQCjL
DD1lSebTcTt3O9GpgOESgV+Bksm9cwmsmCqpoPb/yOwn6kSPCFeiEAVEVFfq
mu1tBlE2nDApeahesbaMV2cxBFhbU7sD2NTUgQpnpbXMZAn/fVuYrIkfHmwJ
zOeY1x2JWTgmWF6wtmFF9/gHJLyklGfStcBJCpsoF4xp7ZEp2qMrQVE3OZBw
Nvbi6uba0aSHOaAm+UKPYpR5LreU82i5extRwf+1GRiV3tX6skXiT2/7TbCF
vYdxHeoVRqBwXmMUNLczN2GOfHmqrr2UqVdYKVuVyzH0+2F+fbyl+8nm0/E/
8cXB08YuMNKsuQRskA7zwxWgdBObhc5kVG7bPEJSozStzinCi1INSYWc1q64
KGyGBnSJxfZoIeNroCKSe6CYur/nawqfhjJKDfOo7xDpIGO4Qk+Z4tkUpGS0
MO/n1i0Vw5Xb38NFeEKrNehrL94G3LdylsehbKewAUyS66pha+aTORMmBmzr
aQ0AEeb5dsdxgcJf7IzkKtMMzc1q0z9h4fdUoUb0l/k35VdOgXvjmUbvdyOm
dPjMkvqlhQtKbSf+G9sXQvBGWsRNvEOijD766IHbNhqzD8rqcw1JwNAFo0fO
NeOaXxU3ZOwz3OhPpl43g8PpkFXAV/qcryTcl9fXW/ZB5LeAKw+VXWvtbtlm
kDeiVouFJMSRgfJ2IeoD8rODQ+Rszx4nKTdnXEhI11QuxzP0C2x2U+6hq0fM
GsWHnHYume0mzUCtDmE72h6udgWN8MP7cydshj3iS+BwHxyAYpEsaCl2Ndmy
s0yhDcsF92tV+MF1ZR/vbOKQg5ai8NFRkPisA5wWScghbQM439sSeW8eZmuo
AVc7RoQeHo1u8hAgEaAxVoDMpWhuLyV/XqTgcD8bLU89mC+NUQHiB8+KrbCy
+cUNcdt3yVWOFI3uifaRcU3PRG+7yJbAnkuyV/bve2Y3qFnvZTqnHjqM+jjp
qnXqJQCBJav4zLzrRr9+H20ID6gE/A5dEuKQwdijghCyC1/lmyYgsuRY87fY
frAqWy5xMv9P1VHKEhXSr8r0PAZf95f4mS1UgWRZJY2beOkQwlIZ9gUAuDBr
KZZdaBe7t9HiTNIw5XvijsXBg8koQ9CBd667g8w31jbbqGxJomiOq1m5snP2
fh/WJQKzYzCMyjg2qSJEs6q6TQnagmF78ql3zLCI5fQZm5DhtPaqDpj/SN71
nX69qI0c1T0Zx8XqHhwtA0t11fOxjm7+iIykX1ZXlQr0vJ7A74RSxfDpmP7a
RgPhEEaMNlSyJiYbpt5t0bp90qkob1bnAn4vrzxKboIwqSPDjKUCU5x+KcL4
4GzDI1eU4Gpq9EGxrZGmWhPcMo38fBW7+McNcDZOtuWPPGquXY+xZYuCb7HD
G1TkGxMd53A29+WUNKfX4ApQLtBOUBe7TCyGsIRthb7mi9RiblFoeZ44ib6j
M00qUPRMYFANI1mJGNjtAKHDCYUmyt/G+mPCDDJpW5KtRxaae/KbCMte24Kc
aJU5Q/KZXxIDX9WZKosIuqMY/WPxkAa93SQ2vzScN3x/JQPTu395ycqgdRec
NjrAOqJ8LvD72e9xVg9ctf2H1OtZyqEPaeTc2P6i+xm0IspF6nPhqkBg6i8U
nAUrjTTt0Y/kRL/Qa9w9at8dxs/SrxgXLH89R7aHWnnZdL58BLf7h4TUIjVp
c7KZNk4Wrhb30ApAXCs6tuCvVTo1UGNKbBGyvRJKYuDPHoLO/JwCWIzce6Zs
/Law5U9L+KXnmvdLga9iCHEYebpPQVdjq4YqjuyIcbaibjaoQp3xkIWnYL53
QT/MOXOFpX3CA08mr/BOj5DCGtngo2eU+UyatiPAETt3sxYmziWkeuOm7F5K
WjqBBnyzUGuu1QkmONxV80XnF8PKNapyMjQEcGNfnpzEingsiRFf9iHJGB5c
7U4r25kUlKYOYgM0C+ijFsktZ/BtDO+/RMjcDRhhhxlZisLwPvS7oPAhJ9e8
FDNe+s0k01LTdPpg+KYb4YNp3CFmDKUcFIq+NsMSGSTY17TcZvHCDtf9rcA6
n10HW3x/5zcPM/hKuqgDXClMawt3akahkciDp+jxoSYgMEtnGCphmEMoWjQS
zS61BFUGEdjux3MqzjRrmkSsCEoZUT77PBIc75rkNpIL1lFvulCoVWfAXZR0
Gk6elKXhy5f6PhaVX2egn3Quk5yVtr5sNBDszDS3o05loFMw1OJGWdRYHR1A
Onw7cA32ZbOrhDKXJavnbsAagB0XU4OlxVeNz2rv/UUa0H8EtVqU9Mi9fOlx
T3dIwiMYv2JBkz9/PnPTZnVeToiqQGdwZzOBw0yGRHNw8ZdlcAkS2AXfyHOK
Hk+oi+dXPY+OQxwbmLBNRmOAr4wJUQebR7HlvJ/dmcREu4szz7AwFERg5Sx8
1ZWFdS2BaR3NPVw5rAQQDy2/yOS8O3iQhYOMtuOyNLhuhVdRMKkLcRhIRHib
46fWDsRR+4I6JTb3vnc5jXAVrOxI9y49GX5wgM9/AKHeRZ309P0Wc9hIDz+p
hBsDdd1/xeDNM67Ng5+cDopZK0Fbk8A06bKIFAmsKO4WG7sWjhkvF0CJP/FV
jtCS79XSZVzPrNcsYI98FP0SsUCnTlb50iBZh0uM5YonwJpp95DwK16YKtRI
ndLpMrZIAYJnDCWmJnMlBW2rbaCQh15TQgPbA25mssIXvYEV/GcH1XXvy2Ym
Cq7rs4eqZkFwg+Bi0Du1n0nKuv/z1fMl3sSHx4//GXWVHPSUuOG7nXI6DZxV
1AZZ2BtMtrVkxFTqmDceGNNbL2+fAPY+g9avZeMlHxHKpnhNVo/mfykPcZNb
X3XD7QHF5e2gIGc3LmdhFxfOcMwNN5PnBcUIVQtOgifPnoPqNLY3knHj3Qfm
OAzWH2CV/3CShf73RM3Z8kcjeChCJbYo246M8QVZf0zeubYIMOodGT+zDz5+
8v7vArv7/y27z74sfCSSsl8xGK1q5LsxER7hgYIc8fr9PZ5KJwVjrY4rGiK0
m2xgypg0Xv3SprWC0VFDTO7d1MsN1VIvABlge8NxQZgBn8gUWopU7RnpkCZ2
lYR0IugNxfqieiBgcYASz1rSeL0Guk2vbH8nilswQ1GjGdJPGpucX1rp9w1B
imcexrcQ1I4mSS4doyI7pZKX9fybXuzERpIRcKmtoiMEfks4dXndMH5XpCX0
uK9pdLUNnjpYOIGuHzDAjmoxN3oIdALuTtvwcy7LxBpkdoNGg5CFki0oVLnO
aUAlvKO3ixLelXV0hKjSsH0uu4Rs08EwXZZ/VmY6PaihfChjJw3l3XUQrwSv
x54jdbWOpUNG/ZEtvzsDKHf/Ux740w2Lml/9GDbFd2uvaGHHx1QK/UIY6hdZ
LqHKZ+I6TcdBRFq/T5PHtnpR9xisLKeRdE6U3O35ZNE8duLy4nV/tVrKZcfg
KM9AgTzjYEYIVj+y8e6qckS9ySEpdvqGGHb9ZGdcjKUXQ/NAovzB5uPiRPxL
dGypKhFIAP2P5Y+S7OOqHEgicJd33G43ZN02D35Vwv8q3Mm3Gy1kxRm44scS
VTh8Kdf+6XV/GArCZ2HedLYiX8zi9yxmVMYdGjKCqA0X3t1xinTFe/Fdc8ra
QZfaPRqJsBLjd+4uxsMHrbf5StjBfHo2z6tOhdCpjVHnzJRztwgZ6+lXT3FV
g/uwwZfwjr4wc2xpU9+r9SAO5J9FL4iyBM3N9e6YxMw07eY2FHhQbBMCeZRk
59tTJ46ZX3lkYAkDeNSJCSdCItwnDY7CtGBiK+qTRonpyUZLIlE7uNLN9DHV
Qk1v2dvvlOquii7tHrajyE1HtD7d/pTyRtPbGVpoUCiwnIcPxCaumIZBQP7s
xYEsIAvkqzUcHXeIgZ0JjLvuCbkF10PByeid1MdyFh2FQjhLGw3V8v2frrLZ
1SaUPaenIQ/ETkLO5zOt2GfO5uC848pOGP84Q4R7hQd0sLiUUtvG6T0q/aLz
rOKOdCWx+/zcrN8SbhxlVxESNon2Dmjt2ddAc6nw4gqyYK935vqsANj0Jj7k
vM3jF2q7EWVcwq+rgzuiyRhzNK5h6O7RDGCFTkKH0xOy0VR9jNpy21rDRTNh
m3sDC48/q/jPkXqhgOO0f8wDkZlDRKNsbBVcxVpkO9+ONTdpUGrVLjJRh+nB
nipSSfWC4JvMqQ9w7H6ZnxIgDj/RUfn7a+Uc4pX8JDXzUSU2hRYggwXDIpJj
uHihlWc33Op9K9rJOPAEU/wvIfNfWLnC4cVPghb2ZhUq9ucBkDuP6+HEOZV8
gfQQUyKjusEu80x9wiz1+ePC3SrL5VrrakaCdsHZtg6vyqMMt+i7/w8aFyya
trVQv5tHOZJRIAJ76CIve5jDZRfPLml0wKZlcOir29H50SQGyVbNUIotYDoP
xKSAiv1dmy8078NPZ+svVWXMeKrxs7/KSLExiRXPoRcofYTKqE8gZPfO7Bvy
C8Yza2SylIOYjjkOsYJc0hsyBSDA1KNd0hJf2p7fYi2VsNorH5FTwGchQVlD
mtmOTk2ssFKdiXYTECICct3RTO+jxl+ziEYEPLnAmUyzRRi8CtroIVrNY9GX
CbchyZNYin4EefIIwp9/Iontv9IvL9OVxhq+Rpe9Rphfqjhnr6iWzLMnC0sM
oy4aQAOqaMrYAkwyCiYmZ+hUpaViUtiq54lt9o6j5T3V/eciec5LTNwepbHi
mvVGtdDLUvImLyG5Fq05U0zF1fO4laTAibWN43+XbbnxynrEcjmUhkEA2olV
Ex9RPCywnbYqRBm6wU5u9PTt3ZlMayKnvfTI/D0gmknt4fRZwT7Cy6wKSJ6p
9Cp9qKd2gH3FhuqRQIEwwW5otRTsDjaxFfprP5Qef+597DUwZA27pcAAWlGV
Tjpd1xHOmEKqbYC0GKDwbFDsGvgy2EEYW0H91gKlh1fVJn7VFN5ID6yZfPQJ
gH4R7D/XYmZ+GMOn7PnA0W5v7hV8hbu9GI87ZtvC9UG/XOy8lyGdF9NVdxA8
IydIaaNEGSrK062G4aWga0KD557bFhglVqMPAwebRdEx0Ubz5d/LXsSvzsHC
IHyTjctExCtq1H9UpYrfc8ZykJF8qGhNgekUTAvGaYYUv1ozmRPxjzPYKwbB
QOqqBdRG8JLzra7zIm9Tt2BKArTzA9Ucs74YzPexJ2/CmqLCe7PLzNexcPOS
Sje7YxBozFUP9uGzaKzIsPlc1z1BcMIzY+1OYb+9pH3Lbuqc1NVWmicSRCiu
39/I/i3bbJDQC4Q/p1vTvsl8JIo5nnwMccCRArnkZU9RPldud+zEDza9TUiU
tc+9bPWwBXboi34Us6Kx2Bv/i7QlFMbzsKUwqP9pgxK7H0u0PXSyuHYiNJeR
6omRYCNB8vle6T8WW07Z9zN7Je7f8+GoFKds2jeY2NlPrC9pzl0YltfqbmD/
uCUzJrQh+k3WUIAqzMqOzKiDwYowrLsmIvD4gY5XZQIyrVWP1740xBEWd17I
CJaCWImldztnCubpKtStzHlfYZhSTh8SAt64mOAADuQAIA42AummyNynIUVT
UOHUiwG0s3F/INVoXx6kSHBuDlYgRP/Zu+F+tiaDa7SIADj8QyGrJgn8diay
Mj4ch8dLB5RMw3kHGWxhvdKXNH+RfdKaQAz9Jh4uirEG7cv7UGlTg6hjO8Sp
2zRewyGM48X//4XqpfNS0fngBGhK5AAWJhyHKumSW24kR7lCpF/byQMCxAgu
YesY6totzPTb8iu6yzEYGfh92V6NdTvjTWWsfiPUNVfbDl6Rs+R9z/Ro+LKs
sE5a/7xQdhovFutNNQAlHELu5RJqeI0Hcj2D+c8VBsM1fTao1lgSD3EZMOTE
WZlCvdU42k+d4gi9N7lZ52YcPWzpGH5Xho6nAa6xarz3iuBExKwzisQwBD32
K28B8zooDO3QfzMEA3MKRxvwPZY0nPmq409s7yHcUWxBOPsvckyxZR3uO1DA
JiC2hoTRj5hmff3oSLv3TqC7VEeZ/Gqr5tYWlANQtDFHRF/xHGvJvUDqYMWo
lwRAPSvi8b5UZ5FBb4oAe4B5es7MjqwFcyF0jw9d7uW8sOAP3TrSuk11Ux4J
MsERWkTg/IWp+a7lXuwdTJitjzi+l6v2s/RlUW7jsmS9o5fo3bdU6aEeMuCH
h/WVK+EDAkj2l0NYPS9DkWCUfqr3c9FLsv6P+xXWSAse/in/eB5hlyFcFSdc
qEuJ3aub+1SrCANNx7yUriEs/JLFe0x3VzSnMe6pXDZQClVUcRFFuAJ567Ck
hzw6bgEC3REvDGTJO+QNmkMP4bM/v37xcirEaiJ4xpPn0aX6vIxgDemuVvKM
r+wvTTqWI+U5rvwNnUZm2lBy7RfM7ObTtidy/fm6vc0u8kv8gras5kNWxP+H
6aTCL4SitmKrz334YotHnupPrb+lLsIIVKaYmicLfVwm71M7yvWIWQ7p9q2r
ATm6aWGt1SqEaUOWeE8YuYD588noLwXhyFEfOSTXkqcfgm+crWIf+veEAEmi
+d964vncU19Ucw5I7MSUYGrXqvRreUKmSZ7WQbGXRxF+rj6ApeD2MAOFbeRt
MLDsIaPzteSUh1EF+siDPZ40HzsB/3feQApYeLLeGnfyp8V6hyS3pvmvAi4U
L7Jdx5XVHUXK4769EMltipbEmlFZCfNcTSmBiz+2SkMhFGW1XI8WysHqxk/4
27dCHSOvukrKJzZgAH9LAcNf+frcRSKrXgMKpdttZjVfKxUSmAwYM4Iuulmw
+rnoLVqoBgsFubk59IUtP0JQfW98DcWRDwkVQt1urLuenr5ncYBHRu3mGVoR
rtz2u7ANtya1my1mwrAaVi9bE6Mn6DlGXHjdQkv3Up7AMEI9DJ3qeNKecUWK
SZ/HMd7zGICRAfU3icWoMVQ2oDFu65j3Hf6RMC/jS4OdUi07vPLErUnrGgl/
Q4UkqVjnMlBbvR4sT+NAuxcwhWHUHM80phlEmAtNH222CzymHua3qtpVxPOt
8BMFknLejcWx9o05rdja3EfLyB9ySxb0Q+0GTIk4gssJN0R9W+DDohhJIW/f
fY2gnE5LqrQjPY4CHg3p49g+BU9GLPqdHGGt9CD0BfzzJHlVGW2pH5SaXPRe
FoCLOyxKBeBAyXf6e4lYmWwLanQxxuEM2iffP0yQzBY7XwW3IGv8+X8TNDzw
wKg8RciLAOO6e0/33tKVL9phnQ7qIhd5Fe+MYvFr9IBAmq9lE4oHz68oaWQ/
qqgB+sN0kB98n3OxrQ5NIKquVKKs8jLDThGMZ5DDZlTfeukvHvbjkn4sirBL
YdlVbvXy1dlrXwjtZhaW6tb7BYwfNRZwRzBpZSVZxKmTKq6es0DiOIFN1Y5Y
O1I6pCGM2Zdspn0RPSZkd5JDa4QrKKyNdMd64OGWi1oxKoGe/4rjCvosYo7l
ZqAd+tD/ILgs443SF3kEPuO5jgg1HgvSNXfnTfVg/R2sBYyeJqi8K6oXmibY
/aDa9X+NReA8B71MquJiuvyev90pCeERsLqMCKgYdEUy8E8iFegfIKXC1Hi8
Yi7QnRhV1sq9azaFw4PiBmsHPSIAORHEOWZV/WXfEb50sAQd8bKJJwZfTReR
iWlkIVmbBDOIrmkUHncD4CIAcpZjP0PEldPZM5nYKR8VEMcZ0TS7Vo4GP3OD
vAxVQbE30Dyk7o6LX8Y1VaA5YNuKVoxIYxBDOhA1r30idA7TaDcKUSQK5Qf+
IXyGsHnE4SqPrp5ohnwOhLWA4ILgW1p9865aGGdHUjog9ALi+XsYiUqMAc0d
4lfGaGjEOZrTaAg8s2mHWty636McOGd2aN/gTr/DIOneynrfIc7LD182Zjsu
JKOsvmsd/e2SWuslWTiXgqHbvv23q5vlaFKoI5j67gJFe+BubLVhul8TfIz4
ALidovcnnlX5p6KB440CDNDWvEQ+m8MpUapurvNsnmvQp9bZU7CoA00ozn3p
mMBOIOF4SxqtdkBdlNEDFrABzL7vlvwTHhz9vRe+jZW+LTS+bCZD/7M34VEv
BLlGmCn/HtwUbne6Nz8a6mcr47l1IPSMYpv2ainO0tVmYpt6H7cKoYgH7ehD
h9c4Wk73G4d3+E4uqApBWVk0sxieWBhNgQH+TRwL3OmmOUMbzApEloDDH/pL
vm7NZ2JMht0LqI0hNNI7JzBcWzBBsgjVGmWvmUv5On51M8luuvLi+leyYMhp
EKMt+jRR2JBw4GBoQs5L1z4OBs2DXJ7c9NOzqYwo49Se1PIPFq/2FJYIyUMb
Yn/tzqKKU2aawL+szDhVeTyYpdloBWOmocbL1312v+x7/MPYesitQeW24anz
dSHh74N9FunTGrpQs6hu7zqoqJ6ZMvKtdaOCHStE6Ch6/PTY4i73siQqEa7w
h26Thze/ZUcv7MeSnaqEKwkhtS91ag+O6mdfLs1V9lDlHLm+VaT+eHoMGB0W
X47UydFj7syl5dkWem2Svg/EDAWzP1pTxvabP1rD+waFdyC/R8zxuvXOPiKI
+LO2d8HuyprrdbjDkNlDMA1JnZ2wdOuaRXWjxlrvjPkWs2eprmDHKpYGeq56
99aHiDbajixQLw5Fuzu5UCkWwF7ZiVVn20fydDrDrKiTCOWVSYCZ6o94H1/U
u/vnPx9IEp294iJBwVnNVKdgr6F9zeobqRxH51caiBL0DcgVunK3IxK6zkuD
y20KJusOLiXipxkAmONmDUAaAyc63JDC20fQLhJ2umHaUqopPAXuk3fiiYvD
5EG99358qzBo35++B2FLTUPuIG/GVnraDfuhyLXrWPkY+OUrJRL35taBSWq5
q/8uuDMqor3NV3SlHnmKvY5kxupFY5rDS9M2WHt4hT/vVD0tXIUIGJ5XTt1R
PEbWtEWuiuNSfmZOWOHBn40ZSMiszrtcEFbsCkbOEC46z+s3YvIjmKpIiPdz
5RvKAibNanZUMkStZYfHm9xZ1rFAdgozKnwgrNN32iSrD/Y+DvC9WpuHVKec
Gyzjh6l9J6s7NjrKv83GEOJs7GLOgbyb9zpkyJmUa8kVMeToOZuX8F9oFSzq
7YQLVlVKiFsXXU/2Fwfuhwuyd4gLC1aHvTFg+rKQNQSeB7r2R2mJISHn8xV3
Ie+hEsTONtXz9UXJpeIlro0aMD+2KmTYm4C+IELDKnDoVLULbn3TSgtS6Vlk
Bn6xi3n0teXjbeK6vgNCaQFOTiokK/HXTnhd7YpGDf5YBZ5/TRWvHgfUxmud
+8nabsLpQMrkNHzrZBhHLWBsLC6v5V5IwN9wd9HlBselrgTrq8JN6k0I0992
gfoMkaToaf6s1Hs6d3mGAkPIVNq1Oh0JEIOZccA8lME+AudznFqlzz4LRt0v
xp4/C/EJ6geo/dKHeFCWpuf2FNhuS7PMjkguJkU3Zm16Ew+24hZz3GE04zLN
QMZrCsaVEDx2h23V6MrAzG2RizeFsOG6VwA+UwXfpdWrWFAwMr/6MTVR1Hxj
fKpE8ZM00CSdw0Lu5RgrG1eMonVUMQ9m7t4PJqwptjP4N2uIWCsbFL1B5TW8
WShRsaU8/bA1G1SUmIzkIlOacFzL0SiO+viZ+Sa4QKYKBLcwb/UD1+Cef/Ld
1PaGYuZ+nw65jVyk0v8AH0Z8DhaUc/1RJySild0HGxX3kfF2Q2fOt9WQH9nx
79sDDc3QlGgTV73DhQKXobZ+8dbTK5uPHz+YAqiZ24E77WWLe4D5aCoWwDIj
ODQhjHfY8PzGNnIVbD+/iwHM4iKhCSfF07euP9lNHS2I8d+LzuAH74J5Y1Na
H5ZiHmHh0j04cSTPdI5zH0QD+y6VhkXo97tn3SpdtlQTlnK6a4+NQIgl5ChK
HL7O/17s0ERXGEVOTTyzIEoFX0Q5va4VIq7j40J0bL6XzqKSvI8ohob7YAos
ENccapy7ZHYecDTamAS8wG2AVIQoCJYfPLaWd8NlVsn6aQJPuNUK/W0MmJ5A
DGDDBbfFmnGqDq4WvrpBPt7cP1nL7X2H2fawWsJ+5DMxZUnmfjZj6XymBMuM
HlgzFSAxNmkCoxeuWq5AqOEZFwUn4quJwffinsf90WAzrtA/WIjv3gEcqoeX
lKyAgCObaUz1cshUB8OVGfXqz9aYdCBmnQ7MQOxTPL/Pd3NCeSCt7dyDkY6s
sq/Y7ybGbuKL9j67kkWVLTCumxyDvsrJKmzu6AR3ZFwoKcoJBFm5Wa7gyhRP
LEh/yTxPxfxF7nyKIQdJ7wWB7cvvvAZXA+MmusU31FGOfWrkzLhqeQmNnV6b
Gq1BYCLaX1ppHPn+dbY4JHxb/E1eTU5FLWrR9i0U5txsdtQEYhsQA3twgV8D
aOISvKIAvhXM9U3foxgejA9jPxvL5ce3R9L+IsIaSbwNit/QlFroI6nvlb6e
herUVnbN42Rk/HohiwsMcKXQEzrLND14w3kdFmDDYTDu8EKGIUzZVCbZZy/r
3H+MbTs+NmOq2R+73U+GPabJSdflOiTbVmWuCUwmzA8XDgWV4zmtej3fUQok
ceNzI8x1FcBDnwyeL7jYO5kMDHzMHf+y4ckkKCRgLptUctyAvuHXS+8Ixzb8
5uIOMQ9UkLxMd1eNMv1jTaO8jWA6lmiFAjIM2dpPrvdciP9B6nnt1Jo9NSBi
LgFaawYdcJ+soi/uSsaxgaVXzgbzsuZpiFfNn0KNGHFzg/e+c3gR0/rCxVMw
cfOrXJ6yms+eSRQEe6f7v3JE+v6kQfY9+Q0JLOsNxngN5eb32FBSTe246vRo
dzBZD0s6RMyZVdvz927Qodp/3/WmtPFFq8K9w57G2BVzxqfqXU8RgiSY0Mv7
XaRu/nraTnnAap3rMyIktDpTpGwkJ+BTyJKEnhr5OQ28WGaZSeTdYW3ALnYh
SBEzJnfI0tTnHxsDlrubJyGUVGGFV3TFApBdfpB7HtYuccwfNTmymA0IUnGX
uVSMOkWtREdzx7J1BwDtgQhDT7pput/bncxQRo1B0/OXJmoMaGx06Sh47kPN
50AU4FjKLJixUR+cYJoMu6Yqg+XEduYVCb5bgEBLLsSOVWu615F6zUm5wc/f
iO9vqMkLIW4qX3mQEWGNyzk5VZxW07CjMFPv01K2HLmVCm5TcKp3c9jV03iR
ZE3HfaPFsmIc2ec4+A0nBjrj4rzIYNmjPPhHRZRnxiSBXd4vvCjp+KYjhEZ7
ipZ8J3x0htAUIqCdWDz3VR3PMvZgrZAiJL7KF+5+2NIEXgmktdtqgYQJ3fUz
OgBo9oGsff0LW0oNePeGuLkbOgjJ8CeNBZ5SMd0eKJppHakmmIFsQ8YJ9mh7
82oOEQh1BmalV2x2N3qCj/dFg5w0QxEiwS9ZVyWiZzRXhbhWA1iq4XS4iAI6
wIloWI4pRCUkWYrerF/yJdgTsmZW8+9cbQsClv1lNsvDkkRPf+UOdJBMExBd
LkvvaMLY1mErz0/6oa4rmweKO5p3T/pVHykTtQcktVNNJwf0L8FVUZIMUNGH
Pq4is6H5rMQ+B7D/hZS8BLrzQuRgp7e4cY8hzKdEF2W49QePY7w2aU1e5MjP
7/Jf9ZW8lMSqCnlCbvnewd9e/okqRsyzGBJJXW51iUdVppCWdKnadW1WR/4v
Ywc48BZdSzaWsGOBH+dQArdcEGBT0IRRoVJzEqt+WyKiUBr8V/15VAN3aDrz
C3NYHprfP+D57gDc0E6kMCJKxdqIU9dqgCbGd+oWLIzJr+S9PKyBSm1S/p2m
s5GBEK7UJ9eZGk9qGN8Gva7C/j0w4+C/XIaYedKIEzsHAqkt/kItSgMJ8wYx
HZ1NN7KmP9NUV8e+ZddhESnG6ONMX13tEbNEi7Erj4gvyoUrvzMm1jPDH/qw
Ca3+gyVwP8igiwEXGAah8WFcQxZtoLhBpQ9sAQG0eKsU/gELvwOqS/aCN53f
GAWUka/0lt97UtKGL/PptZFsZ4J98xp6TaxUsuZPJ2EzlUg35OtkZEynqLU5
XHKya/QJVLlpt/x9NjdUhGJGdClCa2eD0Qs9ah09PVchKBVK+vkJiDQMpEf7
ZFVoD7/S9N7CFjKJ0kNKXP7D7wq6kbeDlEgIobDSSC9tWWBknBeRzjxCjVMz
J8li8A0Cc0BcJ9JNBa7Fn+Vn9wOnKFzdNNbnuXeUDo86Rl05YnbmucAF4v/v
JGTIAOEoWHRzBPqjfy5SZ1vBWdkzOJI8xGYeeLUWIdZd2oDwK6O5Ctn7rsjH
8THCrBb4HFeLY8uiYoVjVvG/I1y7m21r/vbSjf7ObM5ZtTz0Gl5qzUOn6Sy8
9I2/nUZEEW4dWsF9cqpkiN2VsFsfFaJ116lAVzoNPleJp0ab4K5OIS/xL8vq
Asz54qGvg98NZD+nJTbmvy9rrX3Mggy/pRZjefQlQRM4fxR0mOGWzPWYpcL4
giqd7M5wHT7qxUlPbBX5Pw42kkLcdbyUhLleFoIVLQ3cAxHABhpWfjizhXjC
HiLhMp9ovY75TZlXT8a/VBpjazdd5QSIcWJgPkAkmWAzTyY8S65QxGfmzZMW
AeLE4Okt/TKSsYKjDY1gvS+siOvMf2+dTXQtp72URt0K+wS926JqQ0HsSP5D
81PZCjNm8XCml7smlwtCk+EtbOiH8jRSzp/UVvA5YvlM9BJj/IX29HIiysHA
zkaFBuR098YIQZzBi0VadZaSnt7b34tAtjZjANgqyaOdczEqW+IHLYu2Ot2x
L9YuokZN3flkbupHoPiT+XOMuBkdyUyxYJWCk1Ct+WGbRbHPf646Tby+Ef6W
6ucZYgBfmeo9v5TpFT0kkwgzCUmjQK1Z9mS7d29jeI6qObfo4adNtNRO4x/A
DVRJ74sulGMT+7cC8XXfXEm6GETibdU+nTosgMNI4T9xe6+uIKE66LR+06XM
N1R92B9sMd3oV/e4zT0c/H3gRJySZZhO/P366UHc6gYbgk6YB9NcKOg8eF7I
1I+MC1uMm5Dhh2MJG9n5V8mpDZpW2RfEOKkpg53X9CEPfGoN75BalG+WMs/9
y6P/eng+IhNCw6T7cyU8v0SIGFA2zLXxZXZyfbsBljgvG2JAgTR3pAfJ4kGm
lzTmGLuhEh+nznLH3BWuW51tL/1ngJxa/aZgW+73M1FOkGOkgpyWKs/H1Vzt
PSZAOpKNDCmnn0udehyoEgVUNP2p9mg+nvWr8rLX6H+QDLhb8zv7esS7WoQD
1bxeLKPKg8V5A1zNaaiDufhlYBarLqngnFWnlKeTsKCVtGdHCgtiwLMBj+E1
QfKu9XaK6BjNjWnImLHU3Nr/AdkzTa8TUfDg5OjMKijtsYd5Bl5clOuWDenY
1Rwyu0SAPQ3tA0gARUKARnBdbDqlBaqBcmA9QvpIp9r6NXnMGNcBYgTm2htD
uKzCGs0SZnZBTOM5WF8FRlsTSDAyUjwg1xNYZq8/65y+TiZ6VTnmtl5oD/Bd
/PeEc01+WA6OAaj3RwIaN8SX3JWVKTAGib/zoKuIxx9UkzThNXZvG9b9y3pj
GFeGH2yQlHV/mcUS/L/LjjrZ6lfoQ9KCc7mOO+j2/C2sgAj/UpIAmZe0+ff4
r+sy/FOPo8B7O8//MG3tn982k77a72EG4GcEVa9gmT/qQmb3HVWm0Ct5D4EW
J5ztdXDWA0U1EeKeCtmDneMTJmzcWf7l6vRXhmmYsxorHc1QbIcsgVJd95x1
0xmOI5wAhnhVoF/tZ/2VyaE9Zg/0vdI0rug3J+pYJOyHLFz29uzKW6YfNH1W
xMAd6m1ERJ2UnGAfPAOiMdcr/Hu13cvK/FHWoLWYLCC4Z0iyYY3+sgShhBIh
QJ/KIMxgjWAyPm+2q0ZF31jOcAACE+UjbZBBJZRDhK6GR120xAuNbavDHk+D
jzWOIrEmA8j4ng2mdrD8szQRqXrZIJi6zsqs/YNSTqdBWg9a2515PyVB8M/5
L9ZCJRpl9cEfjBHMVA4YOVpZ1lMnRkOOTshmjlNURd3kJfM8tWvM1upHDWvo
LQpu2gEermD4NaY8oexTjVeVcmNniVVvDa6IGBZunrqaVVQemdy+f9S85w5J
cfqhlWjIfNYkt9H0el05yXwrt5LfSo9ajNCczQYI14B2ox9WNwA8uiNVuaM7
P7P2xSKIfIJ5bGdZS2IUQh4d2FT+uC98N4xVO/qgSxHNDQULU9oBOvrfB+ht
kPwJHVNJvwX7/epKAF+yabHe/OABnrkGAmp4FcaaV/Y+WhhA6eteUm6qKdXC
POIZwij7tVW1NBCSDbPRW+IGvoDZ6sj9Jk926UIP0mc6UycTdWJXAm5KBCjD
D/i5/0zEFsU/OnGNwTR/a8PF2lJykOZhMLg+d/7/j/PnFSVfIoqi9V0uK5Qd
qlQuanh8hu+30rnEbvblQfGoGmilnzfsT2yfjrFyhRLJdZguHAQP+9C/f2Ko
4F1OAsUUZN0IVmR43W+mRVstQKtyHMRFuH9gaCyZRmPTQwsluqIel2OIESQA
4wnrb8c3cm4fFgGPEf0OuljpB30+JjcsYpFgMxyJZl97OiPNx/mhCLMEw+QO
3Q0TALGGm8OjPlc4taPURtDkuprWMkUcbk9CZVq+BGV5e/oMpwVQA5zHddpC
i41RxmaROIH3xBaWBqmOmSd4BgkAybVL7begrF+xL4MH7NDAIx0vJDf+1Z/4
P8RENxGXpMIGUv5gf9RBHeXrQgpsshAbEgzV1/75wZth8hEpaLmisVorecSu
WNY1VdOqfuJ2D5WreIsemwKVfsOdSsgMdJJeu5aRdOb+j2mko9Jsntyt6uTZ
2HP3/Jl9r0WCJj2dZIFZRNoQwBiimRzd/l7NxJAJgEthoOT6w16fL61tugop
VOeoJ08+drtHkyFZgqbI7lCogzbVkqEJugAUZu6S7PU/z4cMrH8B7xifCFLz
iz/Xoqu78weGTfnbGYpdkfSf8PvCFFgvjFc59VMzjjS/7Wdv5rnlcsbJljtu
q+vPLG52m6IaeVdu8ilWv1y4ip388DghngZ7AB6hlHIEbUXas/Dhi30PHuFo
yfc0QL6SYlrulKM9Es3Qc5BIJvEaGAPEu88NK2dodb/5/SEWeLPprMgEEb8F
JPLtrhjR5jjiUFm+Xa7HfQiwgYVTi4/zfDjtsjXGaab/YGsH/ku4I65/NxWH
92vRauQjnYzIABqzkW3f+3p7OOu3gW3NgJsZFF5WGs78lo5lUyYxXR+5Vfe4
oUtahOT6wNbVudIujTtbhy5zKnS7d/STNgEW0kWvnaQl/FmhUsseuzpZVbsP
KQ+Q/YOkbyNnAfsg2skmA4TbYkTmTIoKIRTyYUEVBFfv7RVOwnuLjslK9zIV
GmQpENyM/Oea0fn+IW8t1DMgct3K5WrM+651f0eKpOkZD/1s3PjOn/Wcaqqo
GOMq6kQk5r6Tz0Aqtd6OLa25BvgwA/cKzF0jKvN7USfuJZjDco+8zD8iVsEz
r+dRxTmQD9PHbiYUuodC5U9cv1wKRYCyW47w7C0eysShssBLQAgnSjceFas1
dE9ZmYP4V/l8JreDW4Ysf9y0f6drAj+5lgz7tmEAxeTqOTJVJ9SYM6TaYrL7
G99mwfk/NBuJrlFbpaPyvHUzorOe5WYG3rocMZQUoyCFzsF48Y8nYZCl+GOl
skoXCHkY0VzR66PU+2VEKPf5WCbA0bQUJ7CuJb3mj+r/Z63sRJ3YGmHxT953
UbAKgEpXQq+jYXzNuHt4jm8XjOA8/1BO2ru/tKC2J2anEh2hd2elRxhSpcUI
NrawH0exozZYSSEX7xeBI8o+x/1kcXb4EG8hHO99fqLH+tamWrcQTyqqeXrs
MIgD+LCXrLk3dYFi20zFmwn1A7wpAoUMoX1jO1UkeXG84QAOaUeS9e7GzGix
/RC4/n9QzlTctoZCAc5fg9n5KZdAAOJ9PGFZOGuyn9AkMl9y8px24yPo0Fzh
EnoDk+CioO68gzcMAd3EB/HznmDVhm78A2zDjOYowlSVR2YufA6q08Zp0Tzw
S4Uwnl5Z7vr+U36hK3G98uRm//9o49PAEntMCM7uGpQzUKoZw27vOv+fpmw0
fOEf3fZHhvqefiSHi6ByZ4++JFKOaltlfE7aPvYtk9zDAfG0sxBlQTg8RBq7
xsrMFed57SSxo+ocgafNa+lg0n0OW0O8Nvv1LXYmtkuhOxMpVo//7GhDqrLb
F4vRUBj+nJJI1riN6Rx94nihCyUGQVI448iZ0b+qesPYvBWQSX8jk1msX3YX
TivFnaucS8o68mzTOYTAvQoxWeQMLpXt3rgEI3N+prLoB+bVVahqOqCCw1Ig
kux5BtVarAK9APG/JQEE7K9qewnQ1rrBAIFeB2euyWQzpee4dhWQ0CuPX7mD
y+QsA4HMQKVATzCNXfnl5bugZEEpWEgWos5b/SBwrN4VE9c+UXWNe5Llrulh
insZPCWVr8Vgo1c/Ig1UVF9b1bW09C8ciPI7dIX0GVFIaY0MFzyXgDSMpvLN
loAhQyLzSWORqZ0B18lzJUbdH8fxLlTm9XLuWqthtd5Ktt8M3XVrQ8cgwk79
pAl6JQ4niaD1xMFb9kWnD1FHoaWgEgJzUVHDXd3F4QkiDztHGBqg07cHYEsq
JnmkmJZOobXgHn92cjMZec4uvlccI+O2NA403irPxyFIjNQHLliRSSn1AlDm
VdW8kvwhBySAryqBUG7yCyB+qzk7+Kiut0Srz9HjU9GY1izbXPt7+6QUiot5
R8UBl2Sz+MPEjaV9I8Iv+J564v1D0bIqxzE++SGfJmxouJyzdg81pwO5xpyK
cKcfo5VyXKVjE5jTva81sS3Q3lH6bfs0U4WYdtcx5klNT2y9lCPX3uj5NoqM
gd6TbhSTfPnUWApig0JBsQ0kP6sgQVpUjJaIfmWgWoMiaHz+P1oRB+JyVYdT
fbFHSVjnABT7OlB7b2SzdfnYoW83F7M3KP6HlOZcaE5zHzUEKl1JiXVLE1OY
KWpKgtJc2xrGtMuL2H7fwI1/SjT3TeKrFaY0v/ikjwBdsI636TjhVMUHro1h
0u3CIbp2M2oKIKABSFI6m2dtEQUyLFpY2GXjLfd/WMKneqm8RTFEJSjP3PdI
lijTcemlDCHWL729JyWEmJX0/guu3U6zW6qHtgNKkWck+SSkaawVCV2/1hk8
uuNdKwZdgczz0AkDtvTZVu3fHgyeq0B75D7R+da/p1H2BwFDBsjx14cN8agC
1nmx085xLJgnFPv9yQO9bO8ppURpoe2nRBuGTJocfPm2X+VL/lY6+48B1s/b
AjY/L0+/TdQyom9Bt0QQWDyxkvT2522OsbVqNEf74snll9UdZT9WR7SFGJYp
OmYHRvHR081ol4l774xX5yemTmTtQI1FUdpu9b3/bFU17YUO0OT3fphtWbpf
m8feLtVWJ8N3FIP2RNuUCo2jTMutrGLuRDpg2v5CcauNygKbB5751PgUOmR2
/pewSuJlvoyeNhSjnGGEG0u/QGOUTt1VWp5KtoaO0OXmKIU3E9maryZhUMFB
kf2PDm/z64o/DD6TDCK0e0y4nRA3DXuEUUl++zZFeRFDWhV92XkgRrhoHBpy
BEF5IJX5kktyOoQFzIhHsNUB/EcAzT9FXVpPzNB4HzXM7R4AtyKAPxZz2Gs5
qrWjUQ4qgPhO9HT81tMFkjYAalXBlKQo8c9/gdvbgq1lXjWwMy//s2PrsDuG
lpSK1TmpNhJmBq6pXzpwz0HnsfcAUK99E1+I3EBOoef26GpOherxzbv7DTk9
N+nACKDg4jRXKkS5BX53nnU7egNDWoc3eT72vXVMvtmoN9YknhDBXTtB7MMa
eNMv5HPiLnl8iALd5xmiM790ro2R8wdTYFjSxuc8JJeLjCXSoYF1pKZ4N7IL
b+eI/N8AyvQD3tfy76KDUaHIlZB6JK4mQqn+fdtTOW4f5Z/obHSOEHJsEyD7
CN6DYvVlUHrXn7FWwr4B+NW+jY/R5pGqjV9EivMVfgPnzpltuCyNC7M0zeVG
diGmKhyGlNTcn5gobq1rMWTSsxDtmHSUJDu6NYOzGDstL4zzfi9+mUflCbct
fBrC/zn2sNZqAaaJTw6tShZ+P6kRUymCEgd89Tp1+xQHqqVEzJuR0nI26V3M
22ldgKUtHssranWTCzECAti50zTuL6HhfMUZYxfa0dkhkWfEhY4ueLJUxSxK
gB/DS85S8BCS13beA8yl8n5YX5Ut68UpCNPPzBgnrfX2lf8NTvcqJFJ6QUwd
y78poRNnq3Okd7Vnj1ydh5rclaBbgy1HbVGbDHBAHIWergVEIB5qouHb8IKZ
xS476nuMGn65S3l18BNgI99Fj4jKAhnVf6v19D/Nf5Sp9IQepPGR8zUR89bX
jzIVZR+hWPaTXWNRDkTJcUvaYoJhm+tIoOKtchy4JoCSpIh2RvbSQn/4jc9Y
rpEVQ1A3pEqFIuHoAcMiDNyk4YQokAeQ66xrcL1WXBWoo9EHl96DUk3yIxFZ
N/ws5eKPKwg0v1jJFdk9V6OBupr4z4qs84JvaOhIxoUyA7cWSvB+oPTGsbRH
4j6EKwWeuPxcKKCi/H2PkvaO210m09TC9GnaEP7X3xzuFPqwxU9pTY2giNHy
CLQFJh7CuHCiSNNWrHd9Do2MoQQPelUHQuHMqqnM45liF4zClUvUOTLv+eEY
Biz52PUscYH3rUbMCoNCX45EvmeMA+Fy3A4SyQ/sWs5QdSHQ6C5kJgL0o9Fq
7ylB+Wwo7MzK2adwVyglHtUWsikoUnWxromaqVeK3FLN5a+bCttcQ5l8uP48
Sxd0TBN/qRZawroXUQIPqJvSj0nWKNErSIxsDgTuQZwgYUuWr++x3JeNzuOY
317B4VX5LRwpEZkmPfsEi3DxhjSqsyOY4Ao3V2E36Hc8YvuHxmc2sYfmRDSY
K1bDdu6NLnZ4JClXDN9WRC6F9E2iD8Z5RfKk3/TaFPpCw1hP2ZKNj+B61Hfl
ZO8jLQKGpUWW7Vc/ADKwVf3K5jqn2OVcHAzXsXHQSHieXpXTqn3X5pMZTxG+
RGm3jixLG/sp/mXm282XCgr/CdXSQhs6DTsZ9ALTShwxQNQhLjfo/rzmdUjm
xmDreSVr9wyLcyDdQDVgx82n1fsTMZPZI9+MMuzzvx/kXEccmsRtv2/V2m9x
SvNGdwPBm3J/0PNyFiYRguofV2CTEoMFS6qltgOIMVFXTeUHfiElYSFWhx38
cy3mLUYvl4vaiiMAv6eGt694aTkg/tWm7aJcG5hTb4K8Ft9V98vOA9yy1zoI
4kSkQUlEX45HqzT9DX2mrH3t3RuS/bOQuk/3oiFj3VYQOsU+/BK+g2g3drrH
8RLFWjHORK5JzHyfrDJuGLXwmY+TcsE1gIr7inEmQ1uHmI42+EDH3mNfr8A9
J6TmB3DHUeI2DQARDuu+LWLO7oKQvN0EKk9LE4rDb7EtbElpQJ1IwZFsH/Qb
rAEfddMAw2EOdTu2PY1aQ/UTbCohvQ/qkLCUY0LYkssGxC6XkdNBcZoRfzN8
sdw7RpBwjcqYr0o9Zv98hylMdwwYQ1Cb/UyLeignjYjGMeTsUEe9p0qD/fvd
F8V3Ce/4YJuMr05U4X6IgT5QdZxELl5GV6CsCK5hUAFGi2SA9+MIOP5mOAz/
MkPQ3r2dBtiY2qZXMPjWWdr/M0CsDmlvri7A02TNd05pITw37llE1hutCqht
SUij6HfpA+fJ/5UO2IkrHgIXNwzk1JqsORVM3nQMJiCYfpNrMjNpKaJ5zWnE
VbFZPJNZqyV2vXYpmdS3GVS/glrjAckK3+VhsA4eKZxfYEY4AnknjZdyhG0J
amH21El5uCjeRHVFHdNL9V4BXHglMq6Ii53joL17zmMFF+iRwstybvyAl5gL
laWJUceXaJ39X4HmUw2R9l9MXMJlGkERsEQFDOFGt3d6Rnr81fA+MqtNUkga
OiXyUdG4u/i3N976QLqqufDSsKN4+vvty0FtPzi8wTybEw68+0PnBdknQk2+
JveZMsixGqoPvf9SKWHG04ZP+Tt2ykUk+dCAHjVL3MZoEU75rcf2Rr/rrcxQ
LHNpWJ3OClRwXZJT0JEzFmXpxzG2RAZlcc0LlrDsLubjcpHZZsJfVqq3SteC
FHfAzeGlhRW01/tsX5//MmNEnlpA43BThezsShB1A7tUrnp/7GPunqyxlzvJ
io9UCRyw7bVhBJof8vBhbDgFd5W8s3FBHETl36aOTRurlVCsHqufc9JVQ25l
1BY7HqZJlgNUSOroscbuBFhH2RGbnvdCp/JhWS4I0XhLhW16BXDNfI2pbbVZ
+YVIOo6gCNiSfLEjYUmoABNWzwHqlHgii1Xr506/ia6j8WpnzwUhqutSxWSh
F59ob8lZIArDUTvCKS5oyvRKEy9aPn+q1WyNjHcJoASkeeIMGbtWSD9HzcwM
ZZl/5kSq3+xwUnU7gjoLF4HHzI6hBmXaCgFlHWrngai/XEeRHibbyXDjG1fC
q3IVUV3q+FeZ0QI6sbLVj2Dg7AX4fmPE/wmmmepsCEsg4hFw6q8cdupwIsO8
6quEnLABUJ2+TQjlDUaCTTQ63m0imFyaStIY/jIZVvr9dKw1ItaD+wOAy19g
norLunLu/JPgHZVYsrtlA0hKFU5fjUqNOxSgj7i+sCjpvO0YOcT55hcMbefV
lY2m2HDKxuCWQH+vweUmnQzv3nhDU4pcguQDyM90jp+fC6eZ7SWDL7JCHBod
lnK+uxmeDAobAKjoxF0OxOi52zTmbi6QMODReuWRqwBXeA/zoB1187H7GYnN
8v0Q+RWM/rbeWWwXrhseFUC/Kl1LPAGwYA6hoYEdndqqbXzQyB/bat44L5Kn
ljg7ipa/2Ph38mZM95Tsc4QtK1N6xOfII0+vnKbUhf2ZaTj3ShbCf8+oov2f
NpJL4kZVZjrlnRZ7L6J/HrPWOSI9fKU0+EC9jg5brbFo2upiSXnCKO1Nq66i
3zFcnFWF57mncYZOExcvTT/qvdUOCLD7qr97ELCBPOYRB3Kj4GVX+NdKSHc/
ejRUvSiijNu2m3mxjzro6IUWw4CFlliPkZuz61v/YMLqeDeiFw3dL1psoTyi
mP1nnVpwGdJA5hty7B/fnOVAMHhqVz0E6M8guprvEIP4IaYSKlHyLWk3WSJb
VD6DR28CWi4kFN2eXHgwsfuGtIsRM7Pr30KkajPbD3bUzDNTbpLlEmPBz/IS
rEzG4Qbh89F/8OzOOI809ekfJjW1mmURGoSmeaYrelJr0vnsFfyMvmutWecx
wzvn9gg03FQ5m0ov+TXFn8RZCTCwTyHx/8oEKdB85N14SdBHsGhaOf//oYE6
M1b5SD8Gc9pupWB2hyN3zGqFRP8GrHR2+A50PaCPdHah7bCoQTTHtgKo7CM/
Vkgml6Ci0jcdtGk1j9qnLPxpp6L5JdF1MYoiVsEzDNa2SOAq52zbfq9rXsKV
unA5ntRtn8t+ggsniT66dTzgI58LLEwzEwfz7Tv78C5LHm1jiJU/nmiul9Hd
ccbZlGpuVAee5j7UM7yBI+YLXo0WZYVG3Z7qiZcBwIY4kQVVzkhSpXkBCNLg
z/kg1DcHF5kxq9A47mbGU44BVKD6REOSy929xpuvv77p+asf1Q0piGzwWOe7
IXbfn3KsM3n8TdRaR5j4t8/0M2Vle53n6j/Sohk+8mveicN96C9EnvMvDdJU
o1osI233rNprGFCcV29BLibMGN+PRIVst8q6SRn1oCVSSBJaREioG75lAWBM
Ms1mk/P+IXukcISUO0JPOa8RMvXLGEFIImsmZRFEF9KcerfRVI+cnQFHIkA4
6rCucOfXXbqtH8v9n0Qwzx3nlppRL9yoKR7JONPfjP6w1FyCZeirkm989gFR
h0w24Cxyrtbgi9ooSt9DjipxkMsKbXny343Vzhq8+S73GFZLry/E/yjxjCr9
q4r6kiGH/5pa/MfIVGQz0T3rfiQb/HjtIwffMLWH/K39+KKBaN8FzBz+Txst
P7WQ9HI7Vo1ijFGmMh/5P5eC/bYh1F59LGVNsMTL+hL2KMi5uE1N7z4Cg9e0
WdDvezUXYrc7vRhdsLnyCupxDyjAg3Al9iL03QyjD8wWyLP+jaWk/KSQNBRe
SQ0xdKDJvKqOcd2VgbVH0H4Nyity38w7B2Yh1oBYNAls0BvU1H+Pyle98CcB
zzCPdlM+sdz0dih4+wnNBc0XpxYqxZpofyEBOJGc9eQt6vsbN02d1tz73Z65
Afr2LrYuV6XcDN9UL2CmtKcr3coZZ9FVBUUI/Ga/E91zuo2WASgHcao6nSkS
4ImdbGRkNsMG2RBZ9fnPeWO9KxYe494tt4/nZ5Vh2zVkQdjSSriveY/vocPK
UzhFS2miKb4p+UCrziHcMZzUbHDSIUq0AZkEpBQIRSH5x/mLO7iI6iyJasi9
Ao+M7E2MyASelBuMLfcCDdkNAuTTiqVQNxuVCn0TH9tl3N5amqg3ecHj6Vjr
nPBFx2saqtJsBhBpsWZquahQIIufF8Wcgw1up1PK/PXE6QHUBxPv4LZAm/qS
oIc6yvSgF4XnfkQOc1VFUdguzJP9ksfooLVy98J42iNNP8T7B1uYt1xu6ber
aMckXqH411rXLumLItpbvcbe+RDRyN8kHbkLtS+q6KVu6RnIfPljzRgazFzf
8AQwz3Gtdmwt2UzI9LLBbtgxNUn+amz7njy0LW75EHfcHMW8Y7RAFwJjpqrV
+US1gJRX+t9lbsVZMrUh2+HC5frdN0Ernj1cBqi9mhe3AcjM1KBt55++6bb/
wPJTzzflSh9JVptrpCWsh9mZOPPmzzN+env6El2OHbCgayGlf+Z0Xw8dhYKB
uRX44e5Rn68v9qsGZdaDuj8AX7t6olIlAZFr0KjpkGPL67uobQ+detAWY4C1
ipdS4wXUBtt7W/dFvGA8WlJNo4kqpsI7wgUDmA3GDOFlOJ1oVZeYfREmDUQ1
XSKcNJziXGhDH0C5C9GdCHlIUBRssVYh8a+jiKyPI2cQx4rpvOqPJIF9ftrI
oYh7ikohAaQTG6o7b5812Hu35aKBleP0s9Zl7jvOgyxNSpW6aSKlnKH0z/Vu
9p177i8VoGh/ew3GITZnFBNI4+v4dnyA9mayu38xhkQjGGC443SupMJumtDs
+KaSyuluyiFqQY9u/dd3TRdyyndynp2CdwbM+Edf+fMnz9Mbna8zXQu9bfz6
+cqf60B7VxqrbKfdcRL3/55woWCbxhtYt5/C+Zhicpl/B2c4gkY+DmmSWjr9
wngWcxUC+kuODbRiJ3dDZQ6or4XDUeMGrNJmYyUb/d8AjvdHK/2PuH1mdcJT
c88CWcCML/0P4PM7Ge5iRRWmv1w0HsL+MXWxGe55Y4LUw+ln6qm+KameuGrR
m9oHF6obItNvxvEOvCj3QxDmvzPmx/a6gxWj+XSO1yP1VZJAUHquB2VsGSiu
kCrw8yFDiVqmy2vkDqexyQrf4Hcal39M5D0P6DfOoxt9wxQyFGozxdlR6dQ4
A0FuZDcjkLJcuSWpQwlVPCj0U24dAidEzg2C2/rNif2V1sEiZ7AIQTw4fijl
puS+b0RBRtHrqCnJYxLAfAcgIGx77YDBeg4+n0OLCv92gkIJWJtFcizqiwKj
0q4agnJNItQ7BIN0lxAjFMb1XX8fIsgBWVAmbS8pGcCXDfuvCxcP/EIpGTx8
5rcgy72gFZbdCe7Wt1lpfT4WUevOFbHnsmt1R4pRXKaUiMCrIbn3ZCAyEmrh
bSRn/64ipBXTfjj4dIJpLnu80eG4siwjQ2i9ZlElU6qAAlUFDmB8+Y5xE3l2
OLcHN70Gy8U6Vjs44QYHTSQU19kJwL5Cfc5+ycIZQ84b4hPx3D4Q+NGlx8GX
xkGHZLUdUbaxP0/UDBWFkbOZEiZ5pXCS6RuW+A8gxz3QzxwrQ1jl59oiRle2
VA8e/FMP4oJQI5EHFd5W2x2vOPJUroCYP9mYwM/tHLZeRLPFyK3l2i4zAvPV
CFpjcJ/zKNgRD/zpTSROflZg0vJMjIFmkp56deKZWxjluaV42fYnNNwU81k9
m0PxdyT29bYtBPEZ/MDpdCBBGRN+bOOiDWR997orUlODtokX4JCbH+MlggJs
WyI4M4LjRqn9TO50bCyUeEgadZ+AUBTz+MQCq0W96bmVlPohL2uWPzohTxPO
DtRr+p8Yxov6Tr9ATGAkB3Wc8zA7zTfUlBk4tE4Z7GFVy9yGOP0wFtokl8BZ
6KREZQI6aV8mDlFBuxNouq2+ZAmqKUPJakDKWpKYr3Zh4z9HK7BP8A3gk5LJ
t9GgapDPR8gsc0XLdrS95aqSjKidgR4fn3z9c/iPiy1dUr2WqhRUAUbAmbt9
PwVs+S07E/NwdSdBM05VnaiAINUq6P8sLTDffVPl4XtfWcRna9nexzAFBDqQ
7zp5VwvH2v6RGpxvWfuddS4KwRzFrLHeb/Zuh1s3L/oWgtf82pOf39hKO4Wd
smZXvu56z/9to/z6e3qy0dcKz89VK+jGLPQIaVynzrTv1UP8LynspTbbWtJm
9dcvpCp6Xkgk0mT1pzzLI4xkcqZ9eDTnyqNDSJ6VyjeKEvfB5upf1mKyFipd
OMExcCaNyzUDKqyZ5pUTesY/1Wm156QfibmjnbouuAPRwx8+P+7Avg4TWu67
qJqHe1cE1o2yVAeFzgRahobH5Z7bt68v6B+hH1mUPDIUw4DZUYnsDwUDvYGD
z5WVXWltTH0Jkm53BgPSdS7LMwzrlHJn5xn+1DiOS6URvO5v80M5/0O0LPV6
FDxRpcnSqxR3jHpk/9/dQZ2zwalcADCki8Qj7MyMfN93SvBUX19qdcf/0p6l
Nq29Nl84ltz63U/cGsFblFXJriakvO8ymK9/ReTbYli6aDNF/YQTYW5cH2Jq
XtLn/zg0JfGHE0qlp3nr6JQXS+27sgo/5q7y45OJ1tfVxcWW78NiM2y3UKNu
gNzPAQn9aJHLZI6yhlrRMjeK1iDIYk6N8I/zG9Fh7+RG+MpnAltiUIoLU9Gz
/X2UHz2Ht+Ds2wFO78gFGus72JU7UksjnZ/OAPekYO/AfwExJe/wiFbHItc1
SMjq7uCqXda0708DwuKSNGZpXmm7ARuXWrkKWD8QZs4yknmlLkYND5kGWlXI
g9rTh3/pGpevNoDynknY4DdA4fNHOnBm/pILF2DqOf87KtG2BQcb1+ZQApJ2
1WoZcZMcl+9kxgHvCR724H99mv0TT8K1/l+QLYNiDxNhcpx3oH0U/UNgm1Di
edHio8W7IiagsIKHRq4yyFDeZys5FN4OHylN0FiylBqZ1T6ip+NLhE3YLCsa
UTLsz7GV+EkTuf01W7aIVsbZwE41wHKcDcnYK9RKINZ5YzswYC2O5XD+3SA+
SMdkeXIuICzLsOB/11yXpWdOtQ98+cJkZ5TObeXcA6559OPbfWTzZaR4lDQY
aR6SnjcOxMwm4ozby8YqDUi8ZXWiuzH+8+JzHxnBw3YnIbG4OWQWoj1hwfLL
+CbAWbeC8hRvWyyRrrFrqphk+xL0FCBdk7Omn34wRras47EuGC5xDfeJjSKG
jZ2JNljJL/SMsLjFvtGh9IdxCGxF6TvTh8h6jMuvRMz9iYyd/yZwU1Pb2jig
1F6G/WKHV0n3zXanuKI8Y411WvBTwY11aqU2XT8o3PYtIvRhc6NwaFtvQWLO
3uT7WXnHzG4sWioPojZqPNxcrvUNI/iedRVXSo20Fej75ROnpAQ3xFvOPP/t
JeXhTJPeCZAVT0XXim/FoJaGdS4SXRljsaasdLZi/B5pYU26Savz6ZJftKAF
72WLiMBGIXDlsawJ7WnjgJLwKqyx0ktRi2x9GLamJTm6k2UtYYD74/AsE+aV
8LxNkNYg+5SfYy9X+a662rj9QJwbOTGtCdp0yOTGPm4UHjoxeMXzn8s6sIMs
MkpwvVLdPnhOZKg5iHpTi3MoPmOsWGzKd2eIrOAwSvlZc9e+jw0VMYjf7Aj5
zmjiqu3mLFQws3NsEZk2h0+d/Ndj1JKzadpNfqYnYFR+DI36YoaSijpph7IY
r0lpWRKp9e3Tg1NyR0J/mltTnE+k1+soUPwzhP/Q+YmmLgfdEA9+5JhBg2l+
pnQ7RxS+xCpoa1EvF/NToK4C/URQTYfmG5yc2CxxUDm9I/qs2ddKPKGduP42
tcDLNfKQcviUOwTMkDbIfCBfX04GNve3lAxbyxnbLxhSGh/PnGIJ4R/FruI4
rAXFSKb3sux7MaIAz8dvjZaezBG2m4Px8eawMNPI8T4gbtHzTVYsPIR7Kdbj
jnd5C2pLz6XB8yThhIzsaTc78AMhdQiHK5EbicMl0BdnffLL3X9xXASW90vj
xiLDVm1oYw309NuLj6IAF7jJaCPeH9UWVfv4tL9VMBME6/b3WNLeRENd3OFr
0FBalb48q/EAp1UQefT4YToEvgF2AAMebd+7B/YuyPrxhcJYmLnboJyql9F6
o9P3zRbAYIaYZuFScg2Ko2pHhUjD2I2EEB1o4f3eftIeFblkc8pHUwy+WL+V
x/P94Qvb5piKlQMuip65qtb+u2Kfc18oreBlNeDEIjDDgpq8WEPvpbpggoMZ
mT3xAiPPpAVEzyEg3HuBkjbRy+2QrABarJHUBZeItaT0z/pf+wv2FBYZP2pW
5LxcVj4X+40r5bqxeh+/aognroIKYhiB5Z9046LC3aY8/wBYDJYn49vrAP3V
7yzM2JMKX3eesIEsCh7NFErNXazCnhLJH7mSyle3gpyNfYDVl+lYgDIjDCrk
BBmgsLF6Ceg/LRRrjB8itkgqkC6GqjOfzKtT/eFlg+Ci4ulQidDF/yEvLlY3
UM0BKYtah9r7reILq9KWRXoZ9v0smM8EWB27JxAa8/nStk/mxCdQNV9CsiyH
Gih2ADqcIsxjmWWrkJ7SCGuet0uGThOiq0zf+dRcqx+TJt7hufw5ZTVpp4Yg
wmkShk49hEV6X3WQL9ybYMfet9brA9duRm+ta/bAIdL6ymKTeTGNyocrTOlf
mhwSa0qPWHLia9OVM3n5n9py3f0Z9m4y6bOMISUyKG820yIkQm/pmYXhzHDX
xKLhhWGob6yMezrp1LpgLJYSFXJTJ7PVZus36o3Z1YYofDDeRjzI2nSY6Z0I
AA/J6bkkn3Jy7T1YgoXnndk8rtN7CNG4FZ1L+Q+tlaCMzMhmRrb7QrZU7sj8
EtjfUJpHDTo5ENR6J1+gcxD86rSlrAuwWil4Zy0X/htU3awzCDiITVapBfm7
9hwRzb837fBW03VXM/qXvNPvMfHY22kFWrpZzTs3xcqk92p1gs18VymXgdmX
iKysfcQUMOfqjJRSDTl7jPbTAQYa3BDm3N2H2oMj54Ljw3f53boRtSSucSGQ
VSbqJuZNT+/vFVmmW2A/EKbtI4KpaXym2GgyrMVIQWZB6j9BAcyPMdijoG3f
l1FpavFD/ek4P+141AqdDuivbgGkJdAW7RT5zI+cE7HKhPVbBKA95OS9XkoW
JhHcgQW9itXGsujXgN/JYJTk4OAYEY5i0kcJaPlHQ99aG8HZi5J9Z1SMossk
wrP/3+PUw8mha+7VgB19sUwzzwNB1dSiO9AqFPVaMp4eDZCvl/As4b+p7E1u
XCcflxegfcX9n3wwqxdMS6enNraACowI/Wu5S45JrZWcWAFkYiY8OxPNgTe/
2WyKC92AHRbDoTfyFCCzANqsumDKZRyX7tlveddwP2uY+H+cN7YttIWFagx5
pYzFoqYmp0KN8iDFksJR2HU7x9VXXbd+11UQbkVxNskbAfNpFK9j/fqi6+RX
qCN7kITQXB57rmDCzzb1PUDSP2yVNVKBGlVG/UXvjEaemds9Q55AZ6vE0uCa
xmglczs5J6Y1cjauWiUB7Qb8Cs0Ewkf+BOGKSvDVTXR7W4YcuLl8emFvf3oW
BZDCDtwJAT8wF+p4XoeSneqoWaiE8mMIzk30n4b/CvzTqE/XhG8iJjknhgkL
q9DnfiRO9r6+u5Czl8HTasQZax3YtfwNy9VzSVbIcl6xhfx2GfeV93Dr3HNW
XfmB1tevTe3JuiKEyApKIDFkVLQLWbQctPraPFOMbRGw3bEZ7Zb63xV0sp/m
Tq6aoVhxP3QJ/prUfQ+CO7wqcceLZlwAEhpBq1mHU11EqKgyhp8RF2hbObEq
Qi9vgAuVnCGRUfTCNgzkY6YwoLTMpOFsZndUHwxzqhsWjgx/qjUHfRNyQWoL
WzwYO+Z8CYAJW2y1/LjSFOUlOD5cuBu8JLcEmuoz0Giviarx/Y1FuD2N2jxj
t68nQ5WKZuQCzJJkeZ3mxN0rnqLG8rH2wcEWW5Mvs+TOgvi1BcU6AXzWy5NX
/4ZGh5IGwGp/dREvk0AqPbJN2aDhXfRPsIf10r1iYupWYlSS6N2XJBDRfZTM
GqzQL5FyTKFk0bSg5wq3LRX8LG9+2vyeJp1wlcgQmOdHMyhIob9B2Di6gec0
zkBe0YnqsytHYkongPImF0K3l44eQt+LOVxVKgNBTAs+dvLbtd2UUb9dJZRZ
HN9t7Mx+2lizs5D6Iqitldy3NKgDpbFy/7xBknuWdUmzV7jngdFihQ1Dq95p
jSBb0otXeFpQUBvNe1Xp8B/144SNDGKV+F3lGoWVL+ZfD5moVsvQDOl2y8CD
Xb6k/RQRChDJnyi6KWNQ1IAzT+eX80FMd5IElhn5/7nmUNJulriF9Lq3a4AU
GhGBZY2ct3CighaPEJ3sUVmgMHNWgeucysrBe/8rrBmWW6ZP+GwD/+2AP/EJ
eh1O9RkLKc3mLVF2QafFNgjYzSvfeb6NShpacwYRyY92kKB5T9BKQQyt/qh+
RYx9qg2Q3+i0QevFQ6eQ6SuzepXswg0EhqgScXMIti1mk+wd1yhAZekLnpto
RCz9HQY9DcJpkkfWjriPP59SqpYxe2IxDWg5HqmK3QiwLtt9/V5ocgwjf2Fe
suBSROBg82kEmSU4b/AeXdHZTPFCSOrNBsJgFqASPcrfSoZWfWyksVcJJL6g
QV09NpCj+Zbaar0aovsIKBV5WmnIUMJBEpFWjdgF1Rh7diOP/dNlKAMjT+qt
GyQ7gxYRoDxOXSk69ikHRKGIanu/EWyXMdXGTl++ZrSgzelISN0rxOVaeJV+
TZhYffSJyvnTjJBp1o+8h0kWxwY4D1HfDjLYRiWn5LBERiXY7q6hcImhjr9T
PQWOprdekSelkG8mwrqAIWj2DmcqRXvgfuMC9oS8Lmz8B8UF56ZwWITF909P
YHLxnXI9Htjtf410T3OjkC5uJP1TD1BEaVK2lJ74b8hC8c3IfTAqaPtNfLOM
BjM7zhUZqyDmybrNLerDVy1JF30VxR8boMxcgXKZP2P3rhBMoqEyDCacfvGv
VYa1dMbNIvljVkIbCj7KQ3B8tT9ZiSkxUtb+I6xM0O6RnwiXmv9P7QtBbaE6
ur5br2U2SGZ72OL+J8x+dfreH/1+7m7Lc6d8lakYl/u/qqZBJ2DNKBhJ5Uys
L7gT2/QJngWZ2atQ4cSteOlgZOT3r6oD/gqC/uoZY08O2ZMIZnwSz2O5OCSx
dtxodMwDPi40upqN2ec4lGNCEljhvUPrHRigZ8MQWtxuKynRIOUK3UzfShgc
isQp/JD2pb46L1NklSR8ePGuPHfv8sByMf+drBm+bHz8/Tyuj17Rag5Nca2s
C141lEmsD6QhGqMrmOPCK2C0jT55YOemsXY/wyw3bMKPlxzcTAIU5I4S+g7u
3TUSsHPjyuTzS3jRGD4GF+k5g5zrXgxgAYPZwELJr00pJUkKgyD/CpH1VyDP
lGpr9mB2hai+D55F0xex7c+ggvATFMgUZjY2XsWJZh+Fxi/nTAIlEuxR9om1
yk2cOmWlW3s3ZprWXtWSQ2kwsGji1pXvJ/jQVMmwmo3BjFQXlYP3uiPEhwiC
Hbgx5U4blIWJOv5U8hSJLF4cRtkdNLohUPKcVZjl457ASrKXPDREU6hHtzvv
rSSaanLp/baWD3FnmFLDF9VwUBOpmV59CfGtJ1bisuU7hlrXVYa49bTGMm/G
R7y0OmQmoq/FGWhj+gG0PHv9IXTYoKCTNe8qqi/y8on70jjHRXK57hnM8J1z
zsX/bc0OSS5HYBzie01fkVhZGlFgwBQ2VF4LiSDvSsQNtv3+AdjCVdlnqrkC
aTxAssfpcXv+co6+wJVrtOBP8zwOrXBlSCJB/DsX+mxYDWCAVOHUrsw1LjVU
8axbXbsbX1lL9HnfGj8KhHZSmWLEIlbU23+4YxbBV0uQ83Xh2wRcNpH+hllI
Q3hXYhrtN5ZjUE4wRJmORo3YfwXFwiPEtPwN69Lp/aekYuIVL1l+wbTKHXec
gGPZw2lpPBOpdEK/1BUjXPowlC1Z04wjw6Tpp5M+qf3G+pgpB/Z8fQ6L9z8r
F2hdTrD2cvareXT7613NbjKvSib649Skn/VI5hDHOK9b2hkyG3ffepKn8//U
zW9UhtqOIYQQV7VLsH6MXobyb7Fx++dO53CEkLq6LdMwVd5aGws4hbre404p
lQEcKztNlOxW1X/n3YKxZn7+DUz4VhQheuOGUAXaT90gnqA67vwfwvyJs9O0
3Dfooi9xEjj4kjJii06n795mtvLMpsO8a/YF1sF7lp97V4AvnMT+AkRasyqO
EL/UD1k9ZAKoqBpBUj5iHJZSQCbyhq3MrJh9KYrPU8VselvZ2GLBerSRw6Ee
6hKbViUDwGAQXN0CmHfy66dT1h0bdcBRYTcJe59HbD6KMXnlCXAoIh2fNx4d
LsKaPiHhpe1gF/bgrRWnrJ0ORdISO0klJ5tkUlXdnwIenVZ37VT4Ct0OPDxE
u17o62o5wfe3Hn+CLs5kZX0mN0Ku8aodC/+mcuObp7M1ykZdyn4CL0tSv+OE
jQY5kgwQAE8F1lKHoeIiopB9S3/5IzYWdMQGk9aiEis5kirkfNAyiknssvS2
NOkGDGvw3Re0BT219dS+C7PqWFDW3huLgd71MUugVXYKPn7drk4F0e1MGItM
VLpxbYNtWP1A9oGAbhQl3mfB0NtxHyUBA+s2EQ1jFGid7EW13Q6gmPxZkPQ9
sojubctfudmR8YvPY7mb6LvXzPfI0aieWav8RxheraiPEwJj0MbD9GlgAmw9
Q/HJR/8Uv/ilRxG45eZBJaiBACuF9SRdPNnMV7WhkIBjUdCtDCJfo7dPx5qf
a+8xCOw9L1jaxuCRp7x1vCwlJ7COXoXbsfjrVJnb1DK4cSuJslVkiEGZLwn3
aJYnDCWJsXiuoPzEmm75zjTvhoZgJrvYjHYFsY9fLjWp3qGjaUN5L7FC2Yx1
KUNrY39J8zKHDTPHneGEJF1hz4UUGzPUguJ8chY+erpX3Kz0PQMyvyhyPRYe
gW6pFpowDxb+pcc9DNFpzgK4vKiHDi5xPLNv7PPbG6wmzdG68DT+Qppj8Buk
zrUdJcn+ZBs61t1f5wUsCvLZAKkZ818kljb+lYpb1g2g0G0OsWJRZz9Uycab
ceGwswIHVDcojj7lboQ1li/Nj5lQk2LBviRR5UtjPlZTQeX91KCpWfhj1h+6
ZvcgzVmKLx+jLeTmT7W0Sf28KFrWlOsKNNmSc02vSiVxwzhXBep7GKUMLjJb
yoYml5WEGGi/ovKQI1VoZf3pb27GsdHNiMLp5t9/JD4RwHMrPqL5bH+GFzsn
FHx0K4Q0VRYErslN205PqfeI8kdTzgAmQLGGmHqVK4rFXiioZuMazghJJ29A
NBHaChAKeQVPzsoQTwjn/b48Ydjy6cgkj7MN+IRhJx5vSYfQB5yez5dv3v0g
ns77Gza8Egh6fUmQPIw2GRDWd6xQGcTyPBz0bv9CgQImGk7VZNa9oPN5Y68K
95oBKI9KohsdI0IdZ19DSp5rIadvD2kg1HbKd4D/fjdESLWTMnppfZdBVu8O
8x825mdrepvO0iVG4RZD2eJmtiHE0AroeUKmDhF5PuY8bWpY5Eo2VsnNFCLb
WJBC8Td1Vjq3DiJzUlBWT2PfpRn0ShB1DHO9xcFUZF0Yb5oCgYuBPbp3iDA3
1gOQp5LXYBOYvOVJJyimT0BACXGYkPf1JQ0UQNN6kg/udFm34ZMqz7qoXtpE
9vJFw8dQQCOOj90AkR1DUBk6+iw1IxJ5B30J8RDEt7TAT6cjoLVSZuaQhccT
+R+VXDadgH6twE5ah99qNJPF1fB71ZBWUf1moUDYKeGpOyc7i1JY37UbqBUP
RvXVyd9WgOIOdLm0QOftHJ1IWtZYnWzOuBqSige0MO419FNyE/9WrzxB6ReD
cH/ZqZgyKWwQ3cbJ/UXFY0FvCkCzXUzq4dicMWFd2xqS16LhjIiSvPG6bvtH
XjSST+KqmXw+ygWbhbt9L62HkhMwGd64C8+6JrIVogCDpjN7Ka3Uiik4N4AY
H1QVv0QScaama0/FPWRb34QHkaU6H5T1+iybhFyrzYYbcQDQly4twNLkENIT
CtYu4xCiHqxy/dNeF9mJBdrLVa/BllMdF8zn4vIx7MjDOdBFGhuLPOx3oxGh
s/Pffs/cZEbr2xOAHiB+B6RCbYKsvlcA33UfItdg4aG4TPLSh+a1zgKWySdG
lz3OpExUPVWMujHifrsEVSQB17lbyC4ftqAwhiw4WMTezxnvjerrzB9J/U8p
gu4m66N3vU0cYQziR3HokLL4Z6M5z/ZjcoQ9NJ1yl9CmrU7i079zh712Qa7n
aHZ8GRc1zKu5WV4kdmOuAvZxOYd05w2q+/6eNEGVTylpYATGtTNsWdQKIXWS
wXbo2jLHUyEsCHjpeiR5+Nk73BZYlnV76IUoH6zYa/UeL1Y14NWE4ZQGmNhM
Ur0SuSIwHINDP5/UuEW1TMjQ+8IyoOVAOcKvrrNIYkzoDcbW8JxGdCfGcwT1
ienzDqrp16csHevR0NovTARfVdHt+n37PISTMwZrsz52f+PpzpqJyubftAlt
uotxnshdt3xgGMfdK8cNr7zS90K8ID+hmZyf01Kt20hr/uQx438bzhH8k9de
DZH5q4xlH8AYDF0DaLWnjbYjzSmtPwoOFRD3fJXy83BAqmXL5B90MS0DUG8/
n6zHRav9XqvuuRjW8UCZBcC1Dfz9L2nQdqpOA3G21arykT/VxFxEeGTnRwVq
lVJJewaXRD64HDEQ8umcuXqBgqqcTNnU5Tl57SlNGhXv+8mz+53NN1fZLWts
a1Rt992V7puR9syCpHl5ftOBN9lKu6DS7vXM9kKuMlIpSaTY0TVfPizYoaqA
LQFPAJGkNPlFn3vD3ht+03z4TtS8yttZAcD3X/9QlTJPU/1JzhRpc7kgQKId
RDsN8fs/yQunn23hkMKNhZKF5aJAYSuTr7bGy2HwnUUKs7XBCLAwtbGiauXA
n9txa8a+en0zjvkLlot3YcNuExZ1tYzZ5cECJYloKl2zKBNSZZiJ97D0qPN0
d7rUIurWA6l9iugY1NkNRTPCRS+QaOkF7W/yuI2gLiknSNDYZYgxrn/ag6jK
to++hz6K9eN7K8Q1TDlGcjlbdM2fcfSu2u4fAP4oZ1jla518WCx7mVyt+zJT
dvakue1zA8Vojy8tmQGCHzFve+Le1CPWGrSSVtU5ZxWqufu0afT7VfgMpaY7
E/mh0VrR7cSzNKkmKCNEG8xxi9h51iOwPCHFihv/LRzG6Os8YnZXUgoMprz3
WC+w51MmYzqghfbT/GuDUnHvJpurrwYE3fY8zWf5vF0zP0JJvErqNut+uorK
UiZWXyMIPSUrs7Zh9EByDblo7UpS2GH4tKq2PJQS9QSmu0HAfVaraKQcMguc
LM/B4Xy2MLIjXJHWpcBTBRq8c22fdXs24oOquUahsbEI6S9PtMw/M3Vuhv2c
Nz1DbuCRCHaSXWKcS4abu0DAbglifXuzHWRQAjbakK0dVbv6/o2ukh8XHECg
4lE4vb09xmB5VGESmwMHF3zsk99Y74CvjImspqGQwkHxca33UFftpTEtBfR8
JdDCl1WPpSEF84IgGLnIaEPtbUvvQRVpdbNLa322eM/K6xtrUhqg7Dqws9Kq
53kmpaubi6BOuaI9bqZZ6XFhYmLDbl8IoKmmM9AQvQmWjOdG9ymkY6ld3wmE
V8ZOBiM9UUDAlhiZu0+gQHzX5ahQ54tnJIIZjifZLhUfVYgXlux2LnGdkJVO
QlYftuKo7zp+ZLsR3C7GmSKillcaNysydbbm90ThbAylZjBZDSesHMLzRJbF
o/Ox8QJEOutm0+ESH045TgnklozSRNsg3yCA6OefPLSOMRZbg2pUwIDnPR2H
zzAtO+XHiDRf7bmTpkGkg0Ly9IltaouZ2S2RGoELFO5CsNjCD4vr6/+v3awO
b9ZIZk8wMfSni00aU9N/cRAfOrMVoe0SKvSIlUoZ070II9El/hCzXR/YLiGM
31Af9tdxUo1et96H6J4iPGQhvg6pddj7R/3S6S/Jolvxn4s8MXrSfIqvBfSO
/7GHl8t7W7+Dl8LYhr63M4kJE7c6auVl52UwfdrqE4IxRUzWej5+dSSnDGCN
qMc+NFj+kSyzXk4YwZG2CD4mYlvD69/xWoTUf+nVldEwGULWFwrY1rXppk3m
eZkEyu2IWHW9PIQ+/55FOwaWRQxIfErfkieMIEc/Y/LrsvAk9pOjIHC2Jreo
xsxkf3uJqBKHCYbs/8qYmNydKFATGOU5TBp2oqm+QXPIjAxslFfzGFEH7jCw
JJ+8v+hckbWQ12Br8++65eYbd6Y2O1TgLMxuxdA4mWK0a1k/MgOBHlrphC1w
727vDMzjv8X5JBXCWGBrtVZfbs2Y+DSB9VWQSZwFVLH3e8F0wEkEGMmDMdxY
bt7z/eP57LzoQAsaNp3AnmTjatgaRmv3U7gTp90v8ZJAhuDXkJ5eeRGvhf6J
j/i7KAnsypn02l28R3Iwvc8CtRVwhB6Br3FoHqLzQWeNLDhsCRUBSjMpX1zv
1YUqynY1WQVilo7Xxrs7+gXsMgEAGNiHXb4UYzTC8ZTun8S1vq+ZejMjJ+dI
c7ChB8JJqXZcsvSGt0rE8AOkDy29R65s+KyOic2RKBPv2zZ0P3UAiWuXp27h
PwRCWd2KKRQhBQ0F+lqY3RkbzVQkGIrnXzZ9tVfGSsDlYtpyj6W/5/5dDV45
ZALAd/Su8uSKZHUNPO4h/vi7hn1IE8r+aJkXzDG4+l6OvCZ3NXHUxqZfbIzd
+7U57DxRMNRoUPZydVANV2CguhbaTuvUlQwwZFz7YAQgausUrDl3mZbNFUUl
ouQAkg6tEQH6v7Otc7Htw1Eezbu+PsTav+h1I1H1Tow65OFCNGTe/8epbVM8
csJyo9BxnDTGoMl3te7LPSIUlI5m/S/+MQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EpDeueZifZzZsQIX8OXcLmcnSb3KV1uU3cy4+vo4byykLT3m4d65bwzFDfDNuYtJtjMWTHk55ljDRqNeLHwvuyybZlkIvHQst3X9i8AUniyL0CKFAZswtyFCbQWQOl7h9hM1c+QEtxJ14zpfDbnhH/Eo4992GHEipHR3QKJ14OwvDw2Jrn/fNwZmbq1fR4+YK3Hw4k1AgG8NQv6sCG1yuvQx5BuzzNXZ1Fz6b/NYNOeRqehRRt3ZsVcK8N1XhPcjq3yX8NSimMEofRmj8a2BWk8JztWOd0Yum2PzaXxjTvA5FwXz0ua0hrgOCXLpd+HHzvrWb+hAR8GX5wAEBZzBlC6fkjSC0Y9H9LKZ4S0JvOcXNadZq2OAh6oB+UspmVFspbECc1Eif/P/D5cpPVyYJ16gefzJQOWn0545tS0IkjdZXeKjbDg0djR3pWHADX/96zmuXdicOZAIvF+uirx9ij9BKN1XhHTD9SrpokIax6GfmPbnit4RcjsL58JlBc7TQSF+5Rnnbhcx5XVVBzsnPSKnChKid1KUByWU8e0GPkBC8CeS2uwlYgy9EymyegDwbPII+1rrI00kepyRiHr+NT4P40B1wgxMBvkDKbvnJvF1KfhZMq+D+LC6iJuRpeDB7xCKod9g3mJODUQIjoG4+L2ufjtt2NMvUWbYNboMq59WkFkhIM86HwjV3fSHwxcQm0R22LrXkGdJEl8W6y1ZFXXY1a4JDP4sNa23Sa1BlmzRKMUG2YxJWGplx9eXkZDXKSey9QHgUg8oZwEPZXLkQcI"
`endif