// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
icSKTPvvcacae3opUUOr72HU2QK/g1R5keWpoic1HwMcqusmCo9z2OBNnw0P
2m32xRaV9EALKLCnH8suAWmNfDjG4pJOCs4JFb9JE31cZZqEyt5CsjI3UHEO
M32rJETG3V91VHx6oaguy/r04ktLygI3XHR1CDmzr0Q8OBU0/8y/8PEzOVK9
3Maa49lk0xklCVboXEe7uNp34k+lOOEsK0xAPt7Ah1WEJJD4u2PQjcc0Mgo8
3pYtB8ebgOP2NUCioL9EvBE3u9nFLe5A6TSNhgDGQ0obY9YrHuOc70cJI4cz
NKlzIlEQKt/dbm/xXP6Xmxf5nDHbjHamFusPVtapJQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IFRoBFH9yWEc1KOlrmORnjZo6yfHz/Pk9pcoyuMysEw2vvwFviJTFCrAKiSq
ehm59a9cy7lw0L7qGTMMbuO97m+3SeTQU0LH6h6gq8KNOdRoexebBarhpjn0
S2r67+FZiS2TZSixAXYoYZT+cDKi7iGr0/GoCCd4MSj22IhkzKaj1hSsgGLq
l4pHj8F/RoJspxB2WzmtylvjIyVEfqaH0kOvoBzGeCkc+ipcRWhWYCPVWnxG
kk7fyISl6QsM/G8FUpxOyujW5Fjxiemhnt/YV/onKDMd1W+ZFWxnb6zNn8AD
ae+N7EI7mGk/15zdwysd+7lLDeJFOrwIlaEfzb5vAg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W9RQMt5ax+15xk4ySXehMWWv4eU8ej5e+Ei1EcBdRvLud99dbspAraJ5KQoq
cv6D35xi8aye43RoKXEV+vh8Ii3Y5bbNI9pv4gzzbj7CIFjsCBrOhwEn9J35
bPluXVMrG9GIOFRdSCXzAbJHE3Bxx9iVTgA8fYdLVPYOJbii8D6wKKzO79UL
VpzQk7O1MwcSQ+sCZnddOC3H+0IN2aHzkKjo7a9s9Fh++cxOH1sWSc9XVz0K
c5fxysSTvxhFvVxyE2KtQnHKAvVVoZaPwLq+5OW3xmQ9BNZktlmRk5ohup6F
HtBmmb9i45aWIXfwoeKF8HrfgzOllVQYOugwuYvnBA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V33iw1TRjM2uGLydLEYGGq8WehetoAIvh6lBsMd51bZdAirrYO7tfJoz33GK
WtHQtSxmY/F2NSvsMErJVMgJdqSIZKySvScIZR/Z/6O0rf5ug/OKUavJKk54
3MtMgaFa9bIz6AVdWlhzSO2eEMtGk/v1gbkx7jPcqCI9aqVI7ERUXGfAscNx
V12V4xu1PvdBlZRgA/Rw1Qu0iGAzOWihNLsjH9QTeAvLK+DMzO7Tn+sjSuSY
dBiAIaffYMiDeKDArAagjEtoT4YVEamhwF1awvSYUMORJBKxWgekgyqTzOex
S/EfRanude07f8/swxHjdHoru6aqj4rve/ZpNX4dhw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MTIgmc4rGfs5eeFwguAor/qA3i6X9iKq6mr/6OGIZT9oAL9ZUFZskgsongCc
2BLao/cnPyic6dbFnipzzADOOvi+zE10blRuC1wrUG2twtD+4HrSdeFaveRK
A3QMTWJ46+0ksPKHtV44K+8/82+5R+tabBr5Fedyc7DuHu7lVdQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
vcGDqK3z5ThVcOZdaPRq6KbleASXMPD3a2+9XQ+MQxe671e6bhPnwUFVoCQa
fWiuIJ3gvO+82m/+cKaVywZZVCO6cwk/odPXAByasrTKBBATYZrYBGne5xRq
6Kn8Sxgz1oanCC3KTARqQar0isHpZx68sEk16xdm/H57/k8g5MhhsH452dna
t5qnRDZ66y81jBqbM9eisq5i4y5fSMSCOznmRqi5fH+llxvnMPhVKu56Ppox
NgGCx7aKBvwwdVvNPmRs7aHLwS29aZlZH+OCoXdNM2989GIoc/fGtCr0R5N4
a33f6vXNJk86bHvilv4k9fDDoX2wlVDBOU40xUCkNlGA3KfWtn8I6CdW8CB/
Wf33CbGZv6S6s4p+ksjodhJyoVJf+fpucJiXUZ9/yod2ZCghgYAsM0ziPRnS
zTcaQGmBPV7IPDBmvEVh0mNUEqdJqroRerU2UzAXpFOVT8KCHeGZADmUfnoy
JDTyJHLPA4+ixNHRIeQjFsQC+hV7eDr/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UD5GC0NqfHl8+cgSjrOnX4dPMtEYx5Kbw3r+FJ4nzJdbpqiJQ3E0QRc6PBVP
p9PLFKWm1SIKhw7mZ0ztiFYDKFXGdBoDHyeDDdZw7RzxZGmTPf8lUEFA6dr2
b7uZMePgrX8V+nUfSQdYYQe7Ynbjpr64l+TJi57NPr4ZTc8vssM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
k1CMsoSlmEGFHX0xtd0ErMLv8MyJUpM1OOlJYVOfSlcgesHlkXsSSPCXGWli
ncc75EZBafU72KiKAe/rrQ+ytr/4oXhuOLBdXnakpJJdZfNRrGHdykig+ypm
pu4HA2Vah5Qp5dD+avNWt6WtIK4oUFRBfc0brkB6C/utq+SzJgA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16832)
`pragma protect data_block
zxPq05Nb5CV489MFY9HlFqE9YovmDTd9leCHH6WbppC0Od+hCnKY4SLpGk0e
fXI8Wl6snZFrpMYE8i+6MLe7EnrUJC/VSMXIGVpzcMesMCJHv/ligrOW9dOX
T6QO8DCPjsyZCrW0NFFQ4nfxkdBE+NySUkDbe0qMf92UyGJEnLgPUbM9ZZVY
OXiOec9wWtXwo3r/j5HM2xI8pin9Z+TmBg1f+AxGvhBjgKVENCGbDJRLpQKW
LrfO/e8KYjwWwka7joHgG4Vlgn5QhwhFLG/utyO4l6uaiGWesr5xgdR6lFR7
wyJSeydCd6BJLEEC3cYCxot7mRdWQtWnaeNa3kTGEpFpJ0oVl4LFxV2FCtMw
OfYJUnk4oPVdEbXUPUpsvuuxuULqmPydDtrJuMylhbtg/u0oXRMv4jiXLymN
QQ0fpyFL6BHriQ5MflPedPmqFoPhINiq5OqcJ+QO15uHWaj+faIVnIkIatXJ
BHWIQKG5Z0+zsdza6rPDJCb1miLc69rVhzMJPx6UCIyztud0r386QzCeoumE
xybbcoMFHBRgNRqGPG+LxKSHeEr22o+2ZB0qDL4+Xqhd2kx7gpzJS1RNmJpx
9J2q9ESdjVvXM3Z9taauz6O2TVEImlUM3ZG0gXPoNPm2Y2AqPRzU0SruRMFs
U6kKLiSj8ets1PIdR0WBgXhSskg9b9Ine9MUZabuu3YRiwyKwq8FUK2Cx8yY
arFgKvWOWE3Pf4DG6aKxS6xDg5Akhyc0BcSJrcTaQ7wT7zaHeSKYQ3w6ZuV5
8fZtyi0jP/RJ+zh/G934Vp3T6HisV49qlpavG12YQRBiIgeQfXrutBgh9z2g
fAchUeyWPcsyNRJwSlpTPkIUEgeun+hSTjmBfVlCY1QlWhMANdkrIYRwk92h
tfjyOh1YSwHnB2QiEACM30dq4UvWYI4r4Gc1/K10N+P54uuvoRvIIs/RrHpV
Tlg2nZiLUiIemmCw2bbW+j4GgKG5u7ZsB8HDWTUNOcU8nYcGlqAphZxbj0jc
52DDDW5BW8y3rn1jLGb/b10RtK4PDxDPqc1UEa8FxfO90kjRRh6dcJNrrJJN
NBYKNfnI4HeA5P8y5KAyznqnIkL9b3JaBUZGWj4lNTFP/waF0PfVhXfrLro8
TZVbcLXTsLZ2mQGvk93jszYuZuqjgriO+wf7SM3ocitJs5gwvNWLgL1vXMrf
ioZnpjgDNYFbgLRvz31istfjkC/U7GDM6+bthcYtJ7xuK5AsQvbUkoj1t4Ib
EzaHPwadbHAlIHB01cNWLPkTB4udBIoVCDawGJkTz7U3Q35cDixd3zBpMpHx
L2AGpknUXWg1gOzqVmRD5o2jAdJVp8/2cAUb7mEvxf01X7fTh310EW+7fBZt
0XZqgcw8x+sY2MV23AJpocuH1gSGK0eyfR7Q8FlUXvBkUdax7kszpL1vwpVr
JLm69Y7HCCIYydiGE/zZr7EXN6qJqMoHR9S+tU5eQeJjg0SmtqzZjn01NKAp
LpsMK8K06mOY90OOckP2S8GPdDs7AW7Jk6G/nYSA5k22O9oCyGkGLtGRoMLx
9THaZf4pZlKK4R4Ak5glSGJHONazkoaHpcVQ93FF2smI2u1cNGbY4tJGfClv
DHtwizNjbBhBHBuWC/fTx8lpOEPYcW9TUINLP+brHJThw86PDH383SLqaLuW
BXX8JSbXyXT41ObGEW1SwvCDttURGZBYbEnv0MRET9tw6ED259ZjZyApSzd7
Ec766vkriROKjIhzlHbd5tbBhtpqFedMkWTohPt2lya1Ui7/PQvxLvd9os+/
Y996Jm0hKYdsqUms60y1t/NiU6knbdG5pDBZrT4ae3gSAer6tMcJBskvHCm7
XRLU1Hqjg2uTv/sd5Stb22Q0c0PjnQX7eO+v1DNiL3OlIlKddFJ48L9Dgzky
bR2NZ1M51R1YYHoK7VT0FOvsC4A0Em35cJCLrrjxDslv8MMmOyuDoP7aqkhW
KIGovfs8pruB3pa6G3rwwbT6sFMOQUjzXzq8JbzbZ/G8yvp3Q44PhOFDE/T+
uIi/2yV4tY5OlLn/Mq+/XssCRkzCs6f2F8nQQLXzP9mMGtL6s4nA/xX4Krmm
TQ2GX5JJq5ukfam/y4LlKqlixIlcttNZhAHDI5Q9yQW5aVgPtxoEFBqyK6JT
7eC1GhogWWI8fqgIShjO2lHhL1I1RnJRENeD6GOC64uYBPCvfZomxVYM9tvm
hzMeO5gecE2zVINoE0293aDNmOUAnJjm/54gEdQTwGRhCq5tDTmkZniB700G
sIAc7w/5KzqD9eKQmIODAIsjjhBKW4kBrNJBXIMilBUN50bNloFVlxFoQ84n
iSDL1AXk8CBEviBEdZcylrk6TLfsreSNLvu8TK4D8u1NupJEhP6ljix52Lwq
m5A2HqCIwwabYovHHuvLS46jYK57T3Cml7X3XhNszJb1XOYpKbCYVEATHpM0
QH/CVcsiKuoWIqYTCwnKc1mlevllFtXhQ2Vx6Oz/bcCx2dh8Y0UyXAadf4P0
jRPv8sRN9J0rbwd/XECFPqtArNh8lvKbjeNXt+oAastwtsjBLpEPHUbwbvpo
lYeeE/8NYkMDdgx8Y0as100LJ5/ctpvXwAk+gFVHalQRGxPI5g+L/1uM4kuv
84633O14501h7IjRbzq+u5PmF6py0VzFiCXsD9FVriO1qUqLaysyr1zP90Tk
qGO9OPCi6dVwFHYsERkv0L5pAMjJMnIHyWMXdiHEuPtxjHuyS9NFYmx8fweO
gdG3jUMdtyhIRgMxFrHXwtaIHg5sSsZ2L+N0uomkX4Uocvh4C6X5Ez1i41o4
V+rbM+2oV2N69u9ZbD5Zy8jFwy/3Heud6zKlY9dFH1TV+slQF/wWCSAYiOpw
vtBeXyYDgHbTtb3qQMecWz5gvMGO9OG0XJbXkmj3oW3ps3NbPqG7xZv2ZeIl
/YmAT5B+e5gc0TZiiHyWSZnAKvySDBSaQv4rz92bUH8fCjaUPD0nMk/antoN
MoDeZ9uc2eueF1cwASJHMxRDFS+KLm6DiRS24GqsrY8YUKRA/l0DS4WGysLk
z2Bvx1rUICuWt8i3YBWBrS3XVUfleBp9c4mkgVnyJa8+hB4V4oV6GHvuVTFa
GGWdUxw9b5jYMQ7Bf+cKlovZwga3cou1pnPibeOx0/jX79ohB55Kd3LFd5An
37badOtFdALtvWobZIlBP+zbZIb+fr2oRyNkIsrHXTASZj0UyLCVzmIt/vF2
AeDqmXJuVCWTI8jEkaS0f2OA16l7FTZd8/UwUuKrS+6wBEehBIKhA0QXzH9g
uGNmAUdMQo80bksEX0Oz6T/sZR5OxKyzUkZuMOTlPb5jRrwQP7lXdRNhSyqv
wKyEWr2VJQqaTuKxmLA612tQwbUh09/+i0PIHlt71E3zNdnbHAwgPYsriMFJ
zUMqyRMzgsspNBhpfXV/rC5Y7SJsDnqH3PZGhgn+DxrISmk+kcz0g4VmJ8ly
wRgIEINB+5UOea7mq73th4v3KY3t/sgUg+BOP79JKw12/gZ6SY8+hM1iQITq
qlbsIopkYt9myY3QuoLH1013XXEhjxJDdzv5Kb04iW8hysClnDfjrHNwrF2e
u8/eFvjmDECC4p9oBrndYRmpQXAS6Oq3nFZYJ2ArZ1AUW+jf/CSIfkLsRVgx
2Ydv7+NE6LyrBdCYjctKeAyJHm0ORkAcSLVp7MuCCO12xmPDqgVYZYT5UQ+8
fecOaXblO3Maa4RoGTnioAg6T0JtuMCz8qPnEQIcA/w6HtRJIOQQ8NYVSA+6
TTSbU/Mzr2SQw8xqSDdwAf3lpHkUMgQaand/CDhbQ9LNf0QEZqcAC5axi7UP
fFhfEykTu/+VcjCcemdWGV+psaObwEG1iFEfslLJu7QYV+v0zWhN4XcfJJZs
MA6FTcelOkR418VwhPXaoNR/+VZ45WzOfqlav/14m6i2aZTLYEGj27Gy8L9y
uJxMJ+6CuonvtQPWCX7SoK0cGWWw8y07Uo2F4eJY9FTEkG3G8D3bAH39ia9P
vpGwQPJ/JOEJBt4Pj/TfRFc1NLKdJ2D38LbPQZX/qAllnrQP3kFJ7h50LmzP
vsx74kzbRqIR/4tMDjWPnxi2zJCfF3J5VQrYG6o+hwqBI1fiAvdGGZJgoV+6
AzuW3ffbXRk/l5PBIacZZJDBAwPZJWEB9HuDiz149URgMEWP6MKahDDRzgFe
yBzArT4saOoJic2RWX7fGGI+3d3fXyEcxACmZtpAommlOiMQK3cGGhwgQ2FH
k8Vk40I0OvUmbVyOgSE4AWYqKdUm4VCEE4vjVrFNcZJYqgR+s89AgOJaXQW2
jpYIAj6ODlLo6c56g0PylbTbsOYod5I+XySLyK+F6zfuNHRwQy9KTgr8H2Y+
y7k5cZLC1zg5ZXIZFMQp9KbrNk7CPyuUwneIt5Hxe3tw3u4zC7mJT0BKbRxd
op8aBzHVLE/MMfTMNFQWUWbwltreKUOobn6SXRRhQDGcpjgBPcHuan6DGBlm
jhypMRM/qdLlgdmZsK+MNW3oBS85vqEacw1rce+OL5/0PKPAdgfDG6yrkd+5
rR63u803PZqYbw0x87BXFn/Dq8fDgmkfAO8XmppQQnVbYHdLZHFIvPr/fbDW
wXlcTxMn8jf1Y6buL5B7QVoxakOBdxpBBg24RpFGySfbyqat5PwkOsNS3WGS
snnTx6H2UOb6KKo5MKSKEJgQEeepcEgAZI1It0UIH5Jn5i8Cjqo5qHkmRVH7
TivtMgvxqQmmT12ybfzPXAE3Z6sh9ASznW29guH3epgm3aH6epSDA1U2nQ0o
lXoJhUFjKGp+36rsyWjjlGSM9s54dfVYF6+RZbNWU8QyIoQPDT9+Gq7+UOoi
p4wjJT8GX5yX9j/xTQYUcW2dD4ALJV6RhIvhA2yJuJvWSPzzhQxRN140CCal
couy2G+qYV9hnvdjISdxrJ4ahgqV/emF0L/oOLAEBgDMpS733J1YUEJnCNT3
/X+BKC01I8c28TBWhwGLCT6abrRsnxMGTJ4MDM/XT+lrTW3PY5HeA7odIZi+
R5LpoFxfjPg5nz+pDMkeMZAHqcBFrpCTOXaK3qLOvhdDlv43+1dWeVxyKS3C
gxk+zcsfpoNCpRORCH8kRCP/IP44/8QhOiyJd1HntnRaP7s8muGTwi8Bjfi7
yz5hyzhU+wQzli5fT4HF/tm3GN+R3O8gZhacHqt8rF5fYPoiov2m6qUvWFZT
ATX8NZ445nMlZI3gG3qM/gVLXbLz+vOPOxRsuoYP6vkyuaZtAMZ+Irkyr/bs
AcGPBGDMKkEOwc3P06FQGGSrBqLbie3UAlOv2lvDVljOg4lQQ/fUDZn0E6oI
35t9izuB7scrKqh2Tc+S5FCabU243Q2cfx8+d2M5UYc9bJ6QcI9uz0dfur5S
Hn/lHdIN8/+wxnzBJPhhwqda0uh4FpDoppBJbhS4RxyuRwUEVr6Toho8otUB
KnMC65GZ06QU/26qoN6f9xowYqRAU5CVdqJYzci/D0M1ihJdH3JiXylbn6Xe
1LvuKd7AZcChHockZk75XRcXNFnMPLDLyC+12clnUeQnktYPrCXHN3OSRgUO
OotO7R1H8tgpOKXutINNrUGg/J1LvA5mLpSPX4vlygvepnkY0vOccP++dPio
v/iJWRWbSI05XnrfiyAxk3FdTeLwNQbew/ri5szB7ptxwFH/8fk0AEwqUpPJ
6ed03yzEr54r3toP/gFvrXWcgSI0xz4mWSJa7Vaa2wYo063vflZSeyZDTEnw
V1twiaM7TkAvu4qIqMNdE5DESnwBEflNsbmSwBelgdEikn8U6ameQkWWk8IQ
Wt57mQgZOmx3I/edhaPQEr1RCDqF2mUP90JugobmbHibmjCy4E7deByKG1Ia
I/FD2ryJuVqACat+8bbZxHWOxlnKiwUSrSJ5GfeY6VhnTYT+AWEiQM8vZrMK
STlVJRob+VJmAbqb66mCT4SH1fO555hrGW4k0ODQ0psC7TDSmjwDOYdJKBA6
rR2FoymWJiljZKuCORoyE2SprFBQ7ky5M2/S865P73FltZBmdWU9fSJgXtgT
4vQ0i/1Z6sWQXTrShH9N+JMWY6zvRUgXqOy+2lpZn8SZntwqe/2ZG/QGKIpM
qsF+DroPRkzifiRAB0ZMEtX08+bRtPpB4437op1RJSHPh89wKAKlYG+2xkQ8
RcamiFcYzgJIcCxDrHj/amWkWoh7xI3yX5p/gCWpTqa2N/J/U4l54TNhGLHf
tm9japaFlNuWFT0xUFIVknpz/TXL+c11kWKrd9XfCPV1Yt6WSxqRt9g7cEnd
tyT4QL8+QzlVfsUz6hquyJSFnKUyLQcblthmcSQprvHxmIk4LvvBrJdAIZAQ
u4N6RDqTW6/w4bI54ykhiTs8JJZqsnY5eaj1b0qt5WqTuhYsG0XDrIDvUNLf
bis7zoztsawZoC13QYOr5WSavjpO6bqg5VDJzhQONuCU3iPhxZIZO48JjRRL
UFOe0tkxsZbefTRAsTPtlJP03ug1jps7ZChtIHLn7cJ47/uN1+YKq+eTWUAn
2ac82ItkAU1xHqPnXFyfKQFPguwxOjcKCXU4Siu4GB/0PSm2/JqyH1PEduHJ
vDku1DrIhm3xqLKqHGyJWo/uUFayDIKhG7yGEy0pyvHDkl2kgfFKVnb7UBE/
LlTugbsqvbcLiF8Kr4iemhiHBYXQqkwP1VzxTOOqde6GnrzKFt/JTgYlDXri
RjCESAetOG63+XcOb8eXc0cHDbO/sb0mT2dexTEJynbos94+wVQNxAWiuc+k
L4cnE23hKFCnd9qb+9pLq3Q555atRnC+CuAkTOvGuYUnikheJPf5Wc5RXw1+
BdHA+rBO0eu6rVzXHEY7AifPBAtur6EkhbniPqAJtW4/mgq8wIkmXv2ZQZDn
kVLkc/o+2ISwogROzalsTUHA0sgssZIw5kjx2Q7mvVNZ55K+aARBUmvMPTsl
iDbmH3Cgv1D1+wzJXWnSXIP2azXmaNHgKPfS3K76CA5h8nmqfcLQCLXJgWp8
qSY+gbbwqLXAbInvw1ClqoagAdYaEgWSi9auVWgcXmtv3mymZjLFukVsvBgr
MFs9lN6PMKRxZd8WZxtxfg08GtJ/Py/hRY9KfHuL9DWMIzldpOpC17hug8gP
0Fuy7XfukGXnjSvp5JZq/nKgurUJR2GAXdUa9FQex2NkqE1EnnQ+aBuIwCda
RTshY1NMb2faDa2H4ghZD591rD7mnbgNml71VbKcV/0teeuVXCaic3jqT7RN
lmIck0DQcbPXvZyxGMAjE8nR2c8n72KI+//u9YfKo8O3B+GsMH3wpRPEw5cB
xW28TG1YvlBw08B3LfnRDrSoLP/waEH/N7JZfocw/EJIEOmjQJjqLXurHM9e
xNRtOlI22O8/AIec1xJsjbgBEBaejGlnuXsKA6qn8WimM+JqV0vqQ9HR3FA9
u2olVlIQCHaYLje98HjnDxt+Ied5urhfj1u9pKlXsmIrHWuFKa5AdldIY7i3
WtmeLlgLhRIJjeNTZVUjn+18L2OOXktO87P49UdF1UEGMJDRA3cwHtmG9IJK
KDk5OgDBKcXFTfk2iCSyDpYJX3axRQxsMDTRRz6jCXDOgXnUu/52OZqIEk1L
RxqYwJxCl7qtd8Wlc5FQDmBuGtIWriJIMaP1v7KAqV1aC6J5GfUoH/Ddlv42
ddT2nPdCPdMdh+Xfw0BIciaF2QpZVJEupoVmYuiGzwu4XD4e9fxHuhDbAaez
DfnfA+f9QsNrAiXwrua4d/+BVhI7AyE6N4kVfKg9fJAf884IhdE4o3jDvbpL
zAhR1UIptbfkBUsxkDA+g5ExIuMGt5FpC4747gRvSCaJVmAZNoqMBFJoi1QR
gmpUBP3Gt9bEvPuFUxCPISDR5DCblBY6cLVFRinW08q4lOqvWAKBo42JNXkE
cbf6b8+D4M1Ydrt/5UGk2KigcuXC8t1+9pnsNcmB+iSxLDTQ3GCGoyyZyQNf
g0JeERdYsR5kZbk/wCZXxB9Nxg+sWrEnd3Tfyif28SGYJvdGbzY9PxIs5xC/
NdbrbBhxjuCM4DayeuN9Qf+CnWQsGRYvZTXXP4gg7fNyvc2FX+p87ZLSnumC
/2gYYquOeZZeAzLtj5kqk02UTm9/zo2OnBtLVgtoPkrAqqTz2zT0qiRBLj/3
+MXr0Q0wp+eopVICJEVcgHcRlUwAop78FFeFa75pHvEGKOav8Tli0t9mwTtj
mGHWsH3e7xWMZzlVf+vD/y5ky33F9AuBsf11NSbH9oIoROAV73NvqVrtai4A
0LEuLPH+ciI4HRdRDfsBEJ/Gw9v9E8ruJRqq7zz2looMcnfSer8FJzT0C8uL
xzQ8NMRRR8jv+lmU7ZMZ+4ymWxOjiXM54n6+Ddlurh+Eg6QQIzLjw7XUihx+
Xf0An3Spt0VKdjAM6oosohL4wqpHWFLFsXJdtfLds7d7tUsW/1Qf6MsNMfv7
Sr4ngO1HmanOo8NzgmAIYe8kjCIJFm6zhzkF4M6mvml7r75iDUwMIO/u36Cq
HMDJNQZFiTTBHQwBVJzRVjEXA+frSd3STST3JmdAY5JllVBWxDJ4+WmbEJnR
8YubEhfdOQbli+rDAuWdmOTeGP76v0lXufcVOZex8kxioY9ndQrZpz7BbNK8
5EbkGU0TZ++Enk3OSQz6Tba5JW0cfNDd5Zezngdn892rdXkG0fugOKPHhCxR
URNl1Ajpi6rmg46auGf/bIT7s4orMlOQvMeaorNHokNCaR5f3dz0u9LdPfHo
Wz8Z/dqD9ps+iTuScifBlN0/1N5O9MqTrBhDuqnl1nWk+QHDSnhOeuUxEoVK
CEz1u+VRC7LJLTYVgJF/vN1zRPZhYOEN0ye6S176Xhr8g3WrbPdbK3IlBTVN
67p+glyWDBBPbsjXkZSADQFIM9A/2c8XdKj1C4Aed79a1rVnHaAq260QvglO
pvHaRw+NwNYhSzopY12daaJcPRGS4B4DlXoHjLUKlwrUoZGq3trdYSQjGBz5
IdjxYd5Zg/sjWbb9zvkCr/k+mFF+Zz/uwYyywarJTCmB0gdK7K8TtXk8GBT3
L7wqhDW8Kt3u/2L8e7p9/H5vrgpEoC1oFr/sD362oFgeI2PMqtc9G0Bc3rKI
V2ruVrmEpkupD9yA+KAz/rMGjmhNIUOBIH/qL2hJajCIBHQpG3erDZvYrMlO
IaA5qzWhZiccBT1vplblc2LeBiIzrpKOzuLd+Bt+8oU+h5AX1iRoONvenx6K
aDPvuA/rl40AIfJZxQdavf5RlSIYOFh8Hv9U1FIUUInu3a0gvfDc/9vUUorz
zdqSZAiwBWfNk5J5NMtSNISr5rXdhDkGfF+Mv/2CWFXuqXrWLzCSaHb63nRO
SKuJD8jIaIX8OVv+B/vT4E3I20B/rJbzTnGSCULSk60VTGEZjnV74RvONziH
rWx+zodOY0DMydZ3AQlH0APJ1uiTc/cjEhDZP/0cpjrRY63jFUe+jqNYj7Zn
I+eS9syAn26R/gBndhrQOhRppl+Ea/B8vTDPxlZyYtfo9eyfOHaoRT+9wIbi
QVgA4Tq2khJ2x5Rw56gc9vPjSui7drpsVJubGe2M2B50H1+9/6YMiM8Yc7AH
MNoYuwBLbFJVjqzBJjbPLZPLxUd8AozdDNw44XF0BCigXjlmWM6XZL5lvnqW
EO+aZvuFbzpqdPe+Cnka+6UwVZ/YsHmmMsDGrnHAAvnVi97/y6q/OTRn+N3u
wXRCYgHbUrr2ZDDHVkWN9FP5r/VFiwq/BxjLEFu9u3Fy6GwA1pxN2wjFlL8C
NuqFgkkl7dpfPpj13YqC2kHZCa3oehpRa/n8yfiLHwce7P6cnZbr/4UdANHU
Ro/2mfMUOPeJsI+CxFqyQF9siKY/YhyNSanfaPFeskuu9YHtVbqoyKdCxkOA
tIsQdsky4LOuFnlSpDry1JBqAzyO6nW5NZgGZM9qV0HgCbvKAqA0mWBMKh30
SOERUNe+hQLfA+twFAjs4nhDl7XyDLTkNgWPzfSXUIaeAR1H93wcthuXKL57
+plaoI+ZfNgTC6zmZlf3iF1M5iSHIGVDyyBSSDUFMnsGURqFdOe5CwG/Y5Dx
Axe91ADNuwyoGQhWuIV8nNAcDk7xA+uPW6glcH2irLkMIqqJAnNaJP//ybH1
Cluc1YKa03FqcEe5b2UBE3ZXo3oVBPUybqguvdikmDbHIQz22GfuY2k+Ekv5
vGPSokm9MOzLRZKsqsaPHUkGNoAFx5shBUrDBNVTb88P29mT/fDM5a1Bw88g
CK4uL76xptaEOZK98/hfrzFeiYeuP+9xRxh6kcSaWFgdod1PAsUSNPfOLjPi
IziJookIKPD2SF0RNQh2dx/hwQN8rGUNG0W2fd7JJPxFlfcSRR+a2PK/YW+G
iAjonweaUwyzdeSm7CzZPfsYH5maTf0fFiu0BqSKAuUjHcYN3l8rfsWLXF/l
HMnI1NcaNiV6xx0LWSEZuYFyfA5YfG5m7Zk7jGf65EWoKxffnWhMsRkla3nX
iDLeB4PIzsrdZMzw8FsGWDhdNNe9nhsK5wkfmdcP5dQEkno3qnOmXkF54oSN
+w+1Hh1iOaMlTpjAEFbZXgeMIioT3w8bLNVdCjzkQQHJGQtDuFjjb8ceKbzx
lY6i0+tcdWGK8uNwqGiUQx/G8QyhmPH8ugs0P9lEundT3IpUUTIn8fvkwwfN
SBr4z8YABEFJP337bq3rbSmSGtmrF5EKy3yYGL82suMxpL/18oKljujeXj1F
IXh9ScEgESC1/2SuzXU8i2NF/XUtxI9TBvf3MbozxK8yCT7heD/DwxJjMRnl
J5hYMvEWRwMzzJMU1tLdNCJTeapMBSlLe5qs6Alzj/TPMDdRYoOzAhk7h9kM
YVGFIrFvuLq4K2dcHk6267gKIm5E55Yxj7TYGg5ufLV4ofZcRcBa34gksrlI
qDldF7K6zT9pS9Yesel2guA+zkqr88AtbCYqDapw6DLDld9wAUzfwGf+czHU
dd+v6Giafuuh9x+Y+sjJnjZvfgjunv3VZQ8b//0/LnNzEw2c+0AbRytkB7uz
7pbVGuTFOPdi9MxQWCbFceEVXb8OSziV7No2o+5fH1hikt04OggMwbjCq49+
qJKUrYKHZ/CrV3aooZFNqAggiPpy1eWC1F+h4DWJbyHKkT9uuyjHtxtVO/fU
iqJ72Amw+0zmaZrJqxZfnMzt7mSltdJyZIUC/lFAcgwAt+GRYO7pI8XSeNvm
sDWUsawrxy/4XETtXZHwaF5tkCF5j67J1vXkmBJ94dkLcJWTjIrfhFrGXoVt
Pq9uRcgPl1WTl3zrp7Ml73uiyMCN6GwPsQjOK/Q7u0tRVXNbTHV/na7ijuUh
xckJe702swxyduMOQ0Xubcyo6Jqoi0v9SCk8+GCN3+DdKviKqKc1khuPdqnj
+tGtIvxXoGflfRcml0BNksQe693EJ1z1ywHpfcDLUVkvVbBj6P6zxgDmvrN8
KVMqIOtApEW0moK7XEF9J7bp/M8vvGQ7Rktn5B+eQrboK1jjqNIkeu4Vs+wi
IQbpECt3gVNUCETKw+GskPA1vIXzxzwNab9JYQHkK6FV8XCVXCs7WedtvVag
NDIpeq1/z2k1PcQR0opAyRmgenevsW4N/8WylDTvEuX6z8McLdapimK6rbbU
KlQVWrLsEQk+VvzbS0njjvOau4lQXk9OWGlp/GVfA+qcPuztSbB0nt9Zr/Ax
R8xcl6+1j7XUnuP7vAkkGR/lLkMtHyvYWrxNXMTpEs/dKkHe0Z5ryzB0/t0K
DS24oZkdIGGpCy/XAGV9aE0My+jNmHhIVORL9HwMn5L8Kd5H0tcLjQFIZcD+
KqV3XzjFMyhZ4pMqvQpc/4iZiXE8S+1hb0XCnhSJx6B35dKBaOXH348hmNTS
SFFmwGCyKm+71Y2Qf71jWng+C6iGovHvo7S7zKrN9/F50TwnzA2aYB46imk+
k2BBrA37qZl4Qr8QNpdmT9DwWw2DXPUOl3rbUsGzvjW2aMegVU2Hl9ee760l
ie1H2HYH9jE0RNRe3stiQpyT75OEyl4vXuc4pNyocNUH0RQ+C175J4XIbZio
ojkrfZsQg55LMFBaMeJ/LAw3wRr8r4IXAObD0SWiucyUCaj1X5Fx7yslfyX/
uQPGQdIrea0vjs3J5SZFL7bbcbxdxrgu1Y5srstZGC/nDAySCnp5zXxSXGT4
qA1FrDNRc0VgrydyspAppr9lr9+Tavui1uRO3Mroqx5L4MhA71EG9Yax/8ox
biFaoEh/+JQ7jnchvsEdj9Mt3w951V2ahbShFGw8lQ7EIqW5lwlf3wkqZ73m
HnU0yRJbvARDknLy+IxiRrp2FLeVlI4m03PbaadBN5xSbUydsQG3Nyd2qhpr
6ZOhTwyzsU4XkXb/6t8EfiSUNbzgVLwFMJNuS16JBfaKiyj/ih0CkXuhb3+w
FkNrOFmTe11TQEQtTzeFOlcc+TNJrrOpoRHB+ap0/K9uGIZi2hMmLbifjNM5
RuHJY9uKU7vlHcw7OWYcbZHIE5Qro0nYNaQR+0sBmI8W91DAOX767TKbuaNj
/cn1PsdtELnBWAnU8Rti3sSeJPyk0qhjQX7dS9fvJwVWUbr7KchpTZPg/NsR
wHHm9vx53GWln/QIT2pRXlnps4CDjq3N1lyujzXmv6Lr45rxgcMXLXzGFuBN
hhy6qTa9few16L4t0hOoBVZ+jULuQ05OuPlvinrFbQdlbOottKVLelQ8dDTk
YztcC8unHkNkEzibTeDRuduijyKzQOn3sO23T9CwkH1jFgS+wfVS177zSuyL
Gd5xmRUELKJHfL/uiuV6UqkOSmMGavCtNM2uQHRCyXLMXAVo5QuOASANg0NI
n17GNWpHBi6eyV5PI1hpcz4e4p8qnsbrKL9MwG2obv880/t5U8zwV0BWz43m
3VbH8IsWP4uVZlvI/BMJdJfZV/fxFHabb7tHLuVgDGEelcZe9huTyY2UYNYo
raso7VtqNEltWUYWj5PWidcMMtF4Jw9eC1dEn4HoziYlGl/2hX+TS+d6G1Ou
RBwC4/D6Bu6SiCfUWYltdorz0nVGYe9GFXu3p8fblC2q4N6y/BW6oE44O5y3
ODEmHjz9iGXXxGft58lMrqu7m4auog963lgBzhnknvrp+RUfXCvtSBIE0TOO
xFP5rVYk8k9WPQZkKVbLDBmUHMC8s1ZX+rDERbfG21BVzj7PYhO8yG3vDGMW
XzJKChO+zsh84hKZLz/c371z9aGonO7mFIcn7CjP9ZD2V2d4BxbKWLMaLXVX
ucntnaOotAFRbcRseTUzVsbZJmJxa8ZaXrOIcvqOjLMdh0L3wJbdGXRe5we4
sagWjzf2+cEU8aQkpJC+zo7gD5uAzHzT2O3EL5XzFpT4vN27+O+bGVQd4BcM
fjKuvSJx6HcVZMmOqr4tFrusFEahm48QlYp6ib02RsZyOGXotPJMCbyIIiXS
HBKk/ZSstCvjcUwTepFXXuZLo/4qwIauem2k15Ch3U6nhu64ktk0dfAqI7sf
6q4jbP//liZzevigXczwsmvXA59eUgTl2pKmbtN3j9XmbDEce5hItF80sHPh
UHuymToYwJo6UeaZbHYddXve/3h6MfvWq9oikCuxdHeGH3LPL/RNAfvbNCgd
7hYGThIUXHf7SEfh1aTcyvOOagyWYB07UGPlkgSKMopw7UVp8VYFvMDJ4V9d
/AFFP4XcYe0w6u98TvN9SX/yNm60If7ew4IQ+bfAYU+Q3wi54nwJT/MBYeTJ
awIFSzD8wCmTOKPjxgGyY0KzXPAGGVW1YUGHb1jCoVIckJzIJfpl+RlqI4EP
L7DG/90/SSqFgS6YEpIKeKwugqUV8N/dxEPSZto/Saut3O0yauI9mhbmJp09
PQO8Yt1uPquNsI0wf4f1Sho7t1bRllyBom/6YSEd4EA3+Wbmv6lGxzSkINUn
aAMnVK1c2EF0cV+oKfmf+OeQeTWo0JRshpInGO+A6yYwqZIY7QaBb9HpcZ0l
HYKlvdlrH5G3frt9hgoPyKBMCaCcY0WnEfhEgvuuKu77bjPguop3HCziw7Rx
bOjlsHfMihkXPSt8hYsz4yagWhzPT0IBLxSytZYN+YitclUDy2lWDegliQxs
eAgJu0ZK/PFHTADotOz6n2CE0FP+FP2txCEcXOqpYMTR3uqvvgLqRLnpqDZz
xvnDMiZrcurXzJqnMZxgX0iGyTFrZ9rQJM/As4D3wFesN5JZttQ6NVmSHnnE
uE+BAVVcVv5ya3I9MUweLcHOnJbDANNuTtlPN1ge1kGt0zFyKmfVvvs9dfib
14zNizUDxfwrBHotZfimXGZrZoENX7JtdQFG3hKD4ru9LZTuvWyYW6HDoKUW
GpStybqxuWaJZ0Evp6xzP99V3AQNZW0tQOv1IcJXaXCqmAeelujLOzqHSQzt
YnlwsSBTbj5zsDHgKhHivdVMM1mC1L+9cZY3MhKPthIU66MjJjm/YbKRENaW
CoFPWtnaKu0g6wvNPQ/spRNKp2Kkc66ZtsbC7SPO6w+c6zVw13VNVL/Tt9BI
MLYpcCYUIdIS0GUhLt4mrqBQ00zeqbyokutfaXBpf/Mg4WbqdyDma9mPP9/z
fOTP1+Yy85KRt4Wqob+LxvuybO9JxEiHMBui2+/FPjkfhdbvUVgB7AdSrCgy
AKgdZk7Kl73EZ9JeKwoDyC+xcMqtuuol/5kOYMpfNFqj5ZebAqrWpjut87+w
nnLvcUKvbcRZZAk1HeSilrsgBqrpEwUwJim1TG/T8JYdi7JundvsWtxrLE7Q
jFgXO4W+2pJifV7uLp60zta3YuO0JZNGZKAlyGgYLLdjkiVzSjYBusBLnuqu
vDP6Calrth+1zdbiy+tLxluZRC//vZZyFNAumSlcN3myxyI9p+8RIiO4p/kL
FGijJbUKInZA2l/rJX/V5ZREnJAu4JXg5oTBfm2juYvjLICX97fryHHxYbQU
gffuffRoZ1E4/4PmOmmZay6Gs9V4OHt9GCV0YxHWzovpHgnw5Rfcn83cPm4O
ccP7+kBV5x2ZijbSrBh1mFFjnUZ4cpJzx3+yrxeG3W6RZ9UQv5gq3Cw+poFD
8uBhxShEUo8ZQGddT305dAKgs3yYIKyECRPvh7S1jhEsmTU2nA/NsYJzXpIe
tERtwGprovYKJ8erEMRmKvk0ToHKQJ2RP8RUPB4ypy4L0q3tnTW/ZSj9a7xk
rCS0axN9DfYqD/yMWfYeZhgt75fWyGb99Tor9UMs6IvzQHdzvkn5GxTfxpAP
LZvYKwaiTo4zTSLEvIdTQ7O3Glqx5q0QbeU6n/vt1158agoA2mYPlxbFdRvj
ROU1clgb/SroZCPI+W84BIzb0eUZVGxqSxfU9A4RZcQypl7oLnAl+t3pg2Cf
8UFuUm7dx48ICDKjPCdnDniX0S7WhS7Ut/xA/KC2vFN1Cc+kZCAEYzy3NMg1
hmRHaxe6OI6k0qdrqkfEb7rZkQ0BOO7o1KIjzOpiXyS1Q3bwOrOUjbhbHGQI
3U2+pyHJ01Rbok5DVUwDpe1nEfyaVzc3HB1IRLkoPG5rDJx9KpAHCd+KQbmF
7Mvx3wGWdXpEVQzfleD22S7sfVw/rS1Td+qTM+xMXxoSG+uTjGQ6Lae/yIim
uaPuuP+ckcv8SRrXIoE+UhYr9XDRz4SspB6f5McGQpZU2xz75NXSEXt3ux7l
zp2yAGE7rYfKoZ865WqlkbPGeUpZjKN5HqWbsTToKLiEgtBNiLnTJHPecR7K
Y0RmjF5Q81jweXyyyNQinq1LI5rYXJYSxFtc613/k0WLdhfDZ1YrcnMNlWkQ
tF2/L6BuJM3G+ed1Z2D8vjI/WzD3Tm7WRBOQYZ6jTo9r5IKxdE4RvzD8li5G
Elp+FWetgj5WLlCI1spzSO24a8c11C8eIkwZOreTAXYqUjDEfXboK/BADza2
LdMB3DArZDYTiCsavmVjJUVbgR2+qljktkuA3WOZYn4FmAkqNFkmNOq7ooCN
/j/npnpPfdQlNEkHFZMWRHCDzzxxGJaCdIelPtRv2A+ehlGqbrtkGBkNvlvF
wWnuiJBlMvjlDlS7tu8r5lXyXGRl655+C3ou6d9wGFqg0ZTYv24EsfAbxRqM
3lNhmqy0iEoMRZnYINL5ntovuRfwECtSgQFo1eBuIrTh9Rks+G7XeAr7KsQI
5sV7qVpPyAzSnlIWCcX7lkXyqxgnfuYn84umNo2w8Qql0dlQnd5NGuc5ihvM
sXxPspmUoz2agyMARNxuQjPzrBg2BFPQGZqZF/CKTwrYn/q7rFu9qwOwCGtq
pv7W1RJV9dYFmJSemQrWt0NPDeAmQ3MXyhM1pguNw2UgjqIQNT5UyHez9SVf
xU1ME1cS4tnqcmZMwyTNFDlGNKC2KeX/BKlHpFItY4NB04PkjgPKOnMCHoQD
dRkf3THxnES62bmisHbslniwmZcyBMV7/c0CDXxX+tilvzrp1sjD3TjsXQSi
CuRboUsXDw+DxJVO2YZUMDiEi6cR2rG1CMadqz2qkEGk7v4s17NG7ZTMP51t
eHnYuw6pWu3P+jKsFqSEKtxEHRXLDrJlRdGGYkKO2/BWrOqjPHViAouA7d/m
FfE1Mj+u76aoClFcs51JkZUF8cwz8uf7QKKZNSBkrIPbYC2innA6RMtiaAmn
94/DhxVvC/ykPYNwN6fntskqPPaxBm6qzZjPVfu7cCaZQDYc+aJRM1QMRt6l
UqoFuAKE1bjdmwZCtJasgnYCigvjenlc9HLddBJaMejpxduZOzIQ5ESJtTgZ
Wc8P/U2ogp7BbIx7gLUexOfQw2a1/s3ZH64ulaNSareA2rrlIQceh269UUj+
+rY2cXQLn6qZz3EE5HZzEP1fZVzAjAgiQkKDi331o/YLw4vvR46Xuxfjg6ia
ljoBZ8hjherhll/iDusANokCO35NDb2ZkePIIY4CIcJHRC2SOWgVtHGG+qlc
+eDCF3m+gbnA7DHCNjBkK9J+iUwy1zDOq2mUWvhSnOrzPk30C+bb5+0EMwcC
1d87iAT4nTyC9yCi3Fu5fjSsZcDA4quf3gceVd7VqdRvhyH6pffDTMPOl7ux
sw2Cx0gRLbhGWo4tacTY6EgJKIjIdCmk2VYgAoaVXe0gUAmDDSDDTrHuqX7g
mgZQZGVDUl4OkGTaTQkpwy5ly3hJB/W5KY24fSFzK4Azf7DNbbeJ2om005OG
sZAocDL8CSrNPH/OfwcBTh+fOSANmK3z8odnK0Q8+ta/u4Gtmk+daLf50yTj
1YuDpDHGU2gZkwkm1TZcZixZfjmMOEGiKLPt+55WtQ5vY5I9tsmKBBEdNuUF
g6gQF3g523siZCNSttcD94r4XC7Qovf5NNoyJC9d2jZIeC9xci8YDK9HQDxm
ZnqNznHCSaw+EtXKw7WKIYTkoXIKy3b6vStveH5K4c9YiKESDj9iWAdN8g/R
eAWYWLDet9YcBIyGSOpmEDldRNAKjZfsJ8rejULp3IpQyogO0q/dyOavvNcu
3/laBLlT7CvB7/B6e1JV/hOOwkqWY3zIkAMGBZ4gvc8LUQZ+wBcqdPhZ5BkR
myRQMGo2oz278ieCBojmRUj3GeyMexKlXSQyXWadtveWS8NdVwsO7LABpz6s
rYhwe4JNhCTAEqUrRtv7c/9zYc4c1YtAA+EOrXOQRbqD9n2wTlAsDlMt8iRT
angR6yqznyR4cFYuTL8MRf8HYXQFL3XFAtmeUDjr9ClY6qo3OUQoNnwQHLDN
Y3YRiWC2zKm5EWhmIJcixg+6XwTWZfdj0kET0eJEmdSDF8V9w6+M828u2Qpg
Ngvwuk79gGAhyzmyGdp+yxxF7ubhWEdPB+1FIk4M5UnCXkHYCCe7ih1a/l48
ihRCylrLAQQLlNROon1jFOZjbhPy2aCzOfMIKpAf9fW99Gnrzie0PRm3LnaE
iCZaE8SI6Px9svQgChopLnLS/IhOULrcsyQtz6eDMv5kJ4Y9oRZRdXspZXhC
By4T+ao40rhy/Nk7x+LILaKUQR7445SaqGb8Dz8NgREOlfCgdEYH0yDz9io9
YFQu9yLscbP9lHPoHVBeMiI0Q5gVzGkLwe5bsM6RyJ2J559YulcOQqpOzC5l
8xWqhkevZ0pxaDyeigg+0XU6ta56BzDVqghezSJQ2eBj0bz9JenxI4k2Z+8a
GgJx9fsbTNTkP7vzuiXKkWAuhuRS7YuwTgbInKFgkUoaKGajqhT8CxkppQms
q6JXOB/5mQAV6AgC9LXODcCb+ZpaetQc8EhTKNdHktcScRM9t/QCFoPmaNgZ
VdSN94PWEmNg+9jvMk1XXX1VqJB06qFrKKB2TCGngJew7e2Uz+ueyW6QOt3d
NSFvH3bRY9jEAgiBev5EH3d2KMTOpyfKPQV8CpUY/YqF/oLl041wh++VHs+W
5NCtB8rdOavYqWqziURrJjlptyR3voG12Um3tauFGTyCeSkBlFDAoFMkdO1D
OvGY5APG61CztbQflBCWIlbR2x103ROhxICAG9ip0PY2fjceFIzl157EhO8w
C3DRTmvakeuysojQ6AQ0GwCn8onaH9eegkr8YyPGdwsWt6tOl/VPXKNhJMK2
MYLTkDKdE54lVbo67JmmDFUrj7O64bl+47+tLvBWjZioNRYjeUy7dPfnrJmn
EG01ULaNZNLVZrxGoch9vREoIcpc15kErKzyQQNUyH/61h3GFFXg5c3fCxE0
FbyFt6em197UDSqdyahp08l9VEfaw8nmCJHoppL2/EpSgim523m16+75mwks
oP/g1SKAs0vDvVxeOjDGe3UlGXD6Sh3VqJeUYYK6hQQUGjZuZZ3CtaVhsQFQ
f7lzeoq5S6rMTmzHVMf7g6CP0gnXOQKXEiMQxaHLWrV4eokPjzpM6QYB7FfF
NHFMvnnFPfzfKS23ZsX+DYfdungIkaDzKCE6JOdeKdndpeHJAcfEkR1CmtRQ
ySSw7Aias7U5m9SmgE1m1WlCm2TzTj07D1zqser1BT5vvyw8NLreySPmS7rt
30Z8K+l6yIuJqvZqyWNEaKziVt7s217Lle8heNsXGeYwByzmulVPyrqfztBu
a5ml2pTgAAuqKoAnoLKIcmkLwPz+e/miwEsaRWtCEcNx+L4lNI2rK0Sk4qjc
1BS+4sAHDZVkYj4BBwv43GTGPCYjsRclAAMmrdXxD2n3NlX22GzLCRvTbtb6
PBO4ppowaxtt/+7l++qoIKmougj4b5jyFPfEci1UDIzEoy4f8xmSGY7rBJmi
xq+bWpuP7CIMKYke0PX1ppum3e3LTIjQBvJnpfAyjFKMUgWj7IHbEWvL3cn4
PSQ2gPS1sd5fl0q9WRCKxJVRLTtj2upe5k/LywB3js7xkbgxPhJZBb7LpNVE
Z8IQ//4YY+2u5maxiXciX/zX/R0DdKtH5QaigZUBBZakBUc76C4aKs/UIg17
+gyZeFE5+bYKckhbIZt03t5iyMrwS0QAMzK5tT9PpXA+NRqjnZdnHrXvX3t5
x36MwKW3UF8BKKlNqRtOdaqaxRYsJvXNPzPIWuTsdmWkn04DEilRRdyDh1RI
czsbBCOETmYN3ip9vu4QAkZ3mALEY07lfaHr+SCVlMp3iVlg/S4vWaj/hUXL
xc2sN3rECZVLA5nUUhi48g9saZMt6MqhL4ikL3CkXZ7b6SMztOwT1X/1QPjs
HNbeCr4aAylRGQz/PjwDM1YSTGCf3BnvFYpIXX/6HRTB//VZaRibY+sUYaSl
76uigeiAKbSL7zuu3XhbfpUwmCYdyTqPVmbngIFZViWbsTViXyADo9SiX1uY
oEwJZ0uh1bOjaAIC3U32/QumLRyomLP9MoUsthk/OlJs1shyTotxaGTWJsxy
QV8NcuYL3LkjJ7bb0y+p4Nd2TU29W3kuyLemNqrSL69GRxNkJK3/bokoBL8t
0z+axRNmD1C2YfXwBTJV+VWdTlPLRHF9bmSmZNV4mWpiwUD68HYKrgxcE4i8
JC5gTlWkQcFLCsoidi3vso3IBi0GjqOJiqXk1cN5Pt5kuoc1ETaiQq4+nNcD
as5yW7dIQn9bqjMQwM+eCFDreWqD1lRBcznf5icCAJgGb6AymSgT/2i8qU/e
meDSddCezA2ChP9ETAtD6TXnAq8Ynfsk+FKQA+x178mPxfms5g/0b90zUkv/
wjHmCcC8saehC7kKBTxlIgdB1fdz6uliEFF/FCGlE83UzmKM4sjcllDJJuVe
hPu/X7Ip55FKmq/b5DXgj9iP8K1D6cm2ni2+mju8mjpDUFKpAQkO/VqWwS4y
Oatao50zodt/VpNK/MgC8+oThN5cp9D+owl81vWvhnRelYBvtghSQylqWsYT
QqC/eA2sJk5ia6A4tAE54tKmVl3wNIDMFbJLjhfXXf3ecAqo94YHZZiavPyw
hZ/kr/IoYVuP+nCGXdB1kDDImobcQhLHgx8QpevZjiVtWZycTWBCL3KYpkne
5sq5J2+dgNzeKbx4T37WVLiS2kwd3B07enHWN4LjF1i+D+UCBjwVUv9PinYS
zZ1MZJaSRv/uuE5WkYnoutzpM7oTH/ENBCElzU+BO8rmnuWPTIvU1FLDYIVA
h24xrqXIpbhEcHU5WNrZh64NvSf71Q8GcHorRtXQ2bsxeE17qZI+sIdAox85
qnJLsRH9pGHM5NNJWy+tRcRfhqVQ4RRkCXE1vieP0+/Jx//GpAKfTIJJ+9t3
tqe2KM6WGMQ9VwK1SLN4aqXEKbQvy1otKhHstFkbt3YjK3SVUwbcIITk+8HF
IzAqJ32I9iyRF2nDAxJiJQpHpCqwIyoDHBxboSO5KChME5aFEqZTfedJ6kB+
1MCNLeTD4B4pQf2T0VJ9jUfDj9qbbvcrkt/wuas3Fac1MHx/LLX8O145JZ4l
hGnJR2cTn2+iQ12yNenvt/qUEzta2rUJW0d4qjTK1g0ZhN6643QLwU3kjd+N
AZEJDNeVzX5e2ePMR0F94fSvcqnv2yO/Bs2yTYnirIvfoN+O3gGZuPs59Y3W
frqdrt1YXfjcwzz2DYqO7HpGHKa+qWN0u/5A3VYDo22H1irh797CRxf95KAa
aB1NqfIdfn6o3eWDo2BU4b7LJ7RR36MdEdDlnLZ0QV5ZAF0REVHwbBz+0wF0
jyt+N/aZMWo4ugDgSJpRsM5AC9Di8ZQFApptgcivjyUAnzVzBEQHvZNuzLqS
SOC2dQwCpdAd6IEf02sUesPlrFdoJn8jshKwf6/gd6XU2rJc1NFOkX1GTl2e
a4mJCTZg3XUBZvZEc1GPtw/9fWvcla4Blm+/gkzAd004Mg+OM4mO5JM64Q8a
gLPHiAE76RIIAg1ChATLpbTo2ua0jzh5r09W4HdFi8uD7nF+Cg3sv6QrDog/
oZAQEdPtbCUTLxTdsA2SajeUvu0XqBkjgUpKD0beetToBqCkm9dAwQPqpzev
V4MfuaON5vggfr72RrhnGqer2RtaM0g7x07l0040n0G6eB667W+b/SxCESNN
enh5N9tUEgoHCkZrtP6y2E7f1LhMUHPp3j10U2aTAwWUi+dsbvsCJSI26A/1
nuQOZXlq8MMSKPWXrGNAKuxeyAhNfX+QGc7zGS1O86V4eEZbk6EcW9Chtkpq
YiTHbO5XJgRgVqv6o2uVZ6WYPCLFEWXRcvaCkZEpiPzLg/Ou22xQH9B22VAK
fdc27q7F/kWua1yk68OY18IQNotQW720diizE5S2iH6b08/xBYXmahEkQQVo
NOYf29t8p9io2FfOnnDQ5PhSfYpvhWKxi7rkcQ2eHOeZI7M6UPTN8Lqs3ywp
Lf4Dgl1stizU5m6oHVi4tA7bAYpu3rwQsabtfR+k9g+/L9NypnbLg1r2M+tV
Ri7Vgtk0MwGoFTbDPtEQB/XMmx2Sg58E3v7mQMHjy8igJ8A2bud8mgtEFomE
Ueaks1TvauoL3Wxv/rsGAKDB1enAWjt/c3tifJMbZTkAc+0zTFTL2qBqGfzN
ghchQ/BLxZsTScHzEeaaG4+LqQJYTIyWw+WniDh1YthFuT6vuY9DQd6VcBM/
gayjjlH+QmuuRzalBD9qRBlivE4yDgN1mBjoc3ueMeLweTWRBRhke43j8dWG
qPubhCVV3fD+Y0KNZGCsLiJNXor4NzJa1UJyvUdFKNZhNd5e0tSakHNHG2rU
ZVOCODXnN2BhN5ftEP6Di+OHiVl5+6Zs6EKUEpNw1SPv1n6//xDcrk031H3E
WZ+X0/yWXoOVfKmCTtsNtNvnBwkualT4+WZr9VNnED8VbT4cZL/LptzR6KOV
5+w6Og9MWz2+6lCOktJZdEN21s1nDP3RZN8GrqlPVQ4qnzjIykANsIc2Hufz
/VZqMNqU63L5iVPEIUfPUK/dg4Qpo1s8jJR1J49h/WOfi1L4hxOio7hqvCzB
v4jigS3zY9AhhL2M+nsXWHOdJi9etyPraJrnrFbQXkQT9e6LjHLXfPIZD+6i
n04fMGuNOxiI39wDYEh6Wx7ckgxfEFAlzQFHvZoXCCyY4C0ffrbmZAm/YnkU
HiY=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+ErP0YWg0JDdSUgKXZqygAXXyYGaFbdeYbHuRBOYTxQe+5I49CDaggPrhsFJ8qYNFLVk80ertHMqbbLhO2cNcvIx/jgjV5n+J7gOYy/p5JkDrowEGGajr4tB4yId/oMyjJ/UQ133Mq80gQGDzR/mF6qX9lq9HLLeFuBaU35W5857kor2cf26/ckkiNCb7JbgWQHC/73pE8rhHmuO/Bry8V/Z3aCu2ESxyNsEtaijADea7dUie+8iPkYnJsSd+DcE9D/UrffbdKs7WTc976KftDQk6Mktt6SKqp9xpV28JVHImri05goFpAIglRWA5CtILf8fSbXTIfk2xKwGOlwGKLBs0f0DzPKTuk3FL88cIKdE9tR+6HXc6kwq1bOuyBELC4gouD1xHroGL0VFMVqXLL8Yk+XALSL58jHCSPMymMVYs+NbOFsQ1swEXwFMcsTw4sh9vAKU820TYe5XF7wNq6JGTvy4MTE9PQ8b+SG7DnBcwTEMG2u/FBL6P2HQgbWF7dX0QgvlTvnKsBzxjymqTRHL37F89v24ZHF7rKyJ/XSCqP+L7GU1Oxu510x2k3lGBc9FnX4sWGkS0O1Mbmzy7yDrmwiNTDnaVXGQ+NM4I9sO444zaXXKDxnVFlsDmYmteJT2D3u9VEsGzhzzRgFTXgcZHykj0tOD/UROaPIf4gSYbKFuG/iyURbDOTv19/hkuYHuF2i8Z8yp4J80cvCDOY3CXgyIWGLA6Tgeh3+J4sfMvWNAf4ytfk8LTDbIcv/TqWHMcyRh3iy1t6OBK822KlqR"
`endif