// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mBz6byiw4JGp6GevX1tibbcmL+VBMKvTYywgyZJJGg4T6jZcP7whPPj8mOuv
r8z7fqAVK2OxBN+vQgL/ZvtSJgZ3oWod1JLG3h6iCzjaGq5xJ0kJMNlr7Xe/
BAGdOtmJNCjJbcgcf/17fjMhuyrMcoeCpBz/fpzG3jj3QjIfCsyuJDo+StlN
HY7UlqLL52kyBBZAfnKcUXWkIhhH0NNycUUW80fx4NaYq0H3oqP1UjFLgIP+
rGo7DxQdUfm/d0H8CtOHDrJk930J0alcXeq7nil6+6AEqohtLLlbiTAtM58a
obRmQsVTGzBHJgi6Gp6K3c9TkKqQWCdDnzC+MWfjLQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R7/51t/9fKGApHHruMw6mFhpQA9vWNWrfXmlh3fBHwrIpYyiu8e/kV6XesX8
2zk7JfyLcr87I7XUHUzeKESdy1rvMHTvcnINp5SQpcouuAw/Fg/uQEJ1V1cK
xIVU9z2pigVquP1LykyuwS+p2UVJCXo2GeTUmea/vmKiI2bKoVse+ZEQRWjq
jH0L6XdENxosTsA4/hsw9CbPfvOZncwmmGyHTa44Fk8vLmQAnEATmpBplK4r
jZY0oM+cV4u0RjNXal/uU8+Vn16iyE/EhYSF+reGDYPXBCKuUl2h19ywh1e2
ZSD/MEm6NY37WHy9zOLecZzQdQM3i+TsFz5ypTJf3g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k/e+OuHdMGqSBRv+6xMVDzkssIJu7pziirN2OgzLsDiV9MsQ9mVZj+PmX57B
cVb4pHXIBA5/65kzsfRgLgHnYFr99QbDrWMeWcEGRc9scUORRSYhw8mULbBs
cE+OJAwVAzmX9fsV1eNpDigX19oUeJ9x1pzBe+n+OY+Ay7lWv4LlvFDMGAEG
TQSje/t7C4+WQXuzYrqWhcbKfAQK25xwhBOlWUXMRxlgclO465xnC51Er2WB
+mOAaULoF53oDF2itwzJ+Sx2g7kfdnJSrN5221f44ayb5DC29A5faFTdh1Ur
ln3nfgYT9fQ4P+YaJkeY48wD/MTFWu2wgfdQi7b7ww==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n1M9hvPSmVIheeQTGy1Q5NJb73o3wDNPZYV2IeMaz6FyLH8lgMe9c3j5vtW1
VmoD1khq5GtSzgVE+rgCIj8FChCvjPZWrvV/DwokVOenO4dFY9vYpOjd2HvO
lMjp+88mj6/BxqwZgDlF43xc0gLfdZ/NtqMxSvUR9nbwfry4UCryhjikmsTl
m0KSgEyDCcUHLC8JR3i6KnCJhT8YGdJk2MDhvcpD75XRfD+8J7B8pgFSE7YE
Zqd+q6kzF1XPdpALKZWw5xw2UkcLIsxyGpD43cGxkMAnyHVdJe9ih+DJA+8x
ViKY39V8OKwN0Cij+/VFFwkV/l7OOZTUYcBqqplYqA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ddWBTyWTQIeC2uVld7+QnvueTRWlwEAXwpBzHXEV/2MGxzuBLRHJdElZ1OU8
2DUs6Fjc29mt8RR24wCvHeCWxBh6h6IDJOzShpj+1x0dBr7c2vOQVINNTKpY
11Hv+6qezlOO5tOUaDJm6ykdWCP5MJ8If0PV/PYWW/VruPSNeXE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
aE3hG3zeGIbBlX9ULZVsRXhs6ajpXg44S3rvs/5/OE1Gw2fsPredD7hcCcTR
PW9QTWyFlsyu28Ozas/2sS65Ds0KU4mNebDLjmXGTq7GIi7VJn0Ngh5dyvU2
PqRcppHQRAPlnTLzA2y44DWrOcE8d1yOT5RijpML7ts2v1tL1FTMACY4Nzzc
YeldG5uGMI4l9Q7L333LT/pV/w7Jk3/6sh8DF307Sutclfsuxz5Uy6+p49Ei
KZCxW0MYlTkjdrggOyBoJaBjHlEcv1Z0LYLl0KvLvAUm1/ewnPMv8gCxBddi
QvqVxJQ4DfzxGJyZhNYdnZR4E+MZZbJlOjIG7QiqL5QdyfOhiP4gevHiL1Ki
DQ01/xcao7Zc/ed8OMWlOXLwIDlNx0g0WBb4L/Y29LBLGqMFwWYuknfjp33x
nQTBTHnNVrjM89Z0zlqv9v2ngZFVOvpsP5cCj9i0tIxafQWsp8EM6ayV6jnX
S5vSkEGRsSQLppzW5OPt+VN8UysKK5tz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JO1cJmYaXGTh8DuAd0h4z+lkuJMfrbofM2e2HDl+YbQstXXr0Ga/z2jKIuoh
LbNg3KaY0r/JOOyYSoUNMopmek3RNc16HqjZFS5qB3lUYZNu5n+BQmG99CLs
rD5rRaFkKH8VU8z5Y8oPZkFNwcqIi1z2hvaX+X5pjlQft6QC7cg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jdbDUIchjHEEGfh3qNsuQ52n81GqpYcrOtATEbZ4q0JAOzfQP3OxWsUUIczN
qN8IgFLxYMpeV43mLzFraHD+thmodKazOO3iggtpnFM5JA8hwN50nv2E+CK9
52jmGuCbhoZ82giOnprlMUxoCGMg0ikHCIye4VBmb6/BXXQaa5o=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15568)
`pragma protect data_block
OFKgazbz5vSyz5zh0wK0ZcXneOyiB5X7hkJVc5V6qo0SUGI90iw4kO5z8uQu
YAU0iy8fquTTbX6NDw/LV1IubeyYRUEzFal9e3za7xEqul2JB7xQNETLrMz9
Qz79hvdkRinUK0FlLQ7Hjx+aLqOkksAM05d6Rmzz8zLDpQ0HcdQ5IPXP+9pj
lKmchIXi/JbZhKkoeHNaXrLdjwqHH4fu994CInwQJMBaAgIVrSVATGtfAYLY
LAczlOe7BwBpgi+a54LAr9nhHt8rv7H5cWiXIQr0omsaZxq1Dl1VKZgyHiYV
4Zv8Z9COh0x2ZyIR4WGg5b5bWVz0IPgBZWSyBEwf332athqpvOZ4NjL9gptp
flNLvxIDqbylelnzjHRUwf7Ifk/salRBWn0FxP2tvq0kYOU9WUezuWwm78Li
E8cmOYuEmdwAyKaBm2X7OxaN7PjGhwGNr9NxW1Js59SeDMXQPSJfO8P+fZbV
ZdVyrF605wlUS7K9JCrvzCnfhpSdJjjOcmCWYMO1fUhATDbrD5BSEGqt4V7g
WrsCfroo37nNUn26p0hKNPiT901VYtEI/fZI/W9V5SIM50r4pgbn47pKqcXd
3uKx9pUl/mBk4A1LJoiZe2EGjaWFM/YDX96FN9Uj8lPOxJie/YpARL2Yqd/G
M0Awm/V+V2k1GavX0DXcnVVUWiPiXjIpP6UVYjDQBixuU1vXzThZT+zrbNdu
qBmegUSTkBH6vTnTGHD/IelAyvssNHzfT4Axz+A0MuWlb8O/XKTIJepETfI/
BtmUzmH7N5DcktdvG2jw2e69A/bt7NC6+toGgE8KQFikQ6xC02rXazcwU1A1
9nktE6qpA+atGzWwdA4abtOMSNP+6IhBWZKEsJmQECiwGF8Zcbtu4HTZkr8V
ACTG0ccMJaNFkmnzE43vWlL9L/PO0+ErUUAQvHpyBa9BgcAZjBiHjWrC9ziu
P7Qx3Z9W9yu/fRy31QSIxzJZgkdnMFHR+PgTpeySrooEaQicSsoiDY+unqsv
htNh+tbU5S3Lkha9PZmC9EjrKmgIt0s910pjeSl6uBvuAbK4iukADnmC/v6u
CT4ZdlJIMHW7uTIccmuHb716VSAHE20jiqrqVLAm2KDtlV3GyKjtgLHj+GTx
uAmh9l5KSq+Oph6HCAQDRVciafma5dMEFN7iDgB3qI28lwSp49zd8D5PxcVP
8DriiOecddVlBPbKOK3LoH/hnOvmVSSLL1tvSO6geEcS1qSDzE88lxThH2ZW
IndaLziO1gS7Pgg78PuPEloAGUE2bQRzyfW+Lxiugfi7Xop2utvEtdJr30++
vtpRbgi7K6a35APZprfNzp8EyhGY50e0fUKjrO+WY2nQx1mMw115nfqn0U9j
PJI4a4KvkW8sjgtnuMSTDwvtAAWzDqiOTy2V6KfoEtQW60r4v47LH56XHywQ
G0F8KglKarLedlclfta/s1AYUgeIG2KHR35X54IeLEneuIB2zUviP6+Xewq+
YVoNidNf9GdFKz1WcK6hkMmBuj11Tw0NI1IJYL/kPjw3OAiVfDCmmHwuZvIO
yFZQw5rAjIBv5Qwxoc5Yik/XMiHQpFJdxuTiluCOqvIxtLQO8MHVfHD6NLkV
ZSfnid1Gzw8CFlBYnnC8Ap0nm+52oplV10X86RB9EMUv6aZnJJtrheju145l
Ee1dT42H5dME3a8ZxS3X9lFN38Hu7/z58CXch3W2EU1OVjpWhd3Z85XsK5Pv
mdAQUloYaYsQky6cBGE9fVR/MBB2rG/cRyjHrcYTpQEmxxXGLNlRyS3Q1XQU
Vkr/Ln2rujcqUN2O6Giq1m+3NnkP8IijFblGuNC/cZqFBIOsryqZznq5e5BJ
dXPkN/zMbrG7xcRl4+JmLyA+umj6U2OqaHInviZrMCqB+AXpr2VZzlwTzOhR
ZmoN+2BBW/l6dnnlWTj4S9tyNNvZszD1NmGt4XwVosAsen6A4g/C8QV+uUjo
QxqoUajv45raTY5Dzt2VWDcnJlEswtu06Qa3t5S5DYy6tk+KH2i0e69K1r3H
tIHzLCqH7FpUE2Z1dJ7fbc6kt3FXx+F9NSV+2yCN8vVcIV6eBApau05/7eKi
U3N564DAeBVZUuUa0uma123z+YSV31lWbsYJzgmr/S5yOX0fsoYP4TyKzdF7
RnbWcPhQw+dcfV+FZ+SNUgdUksbOd35uXjzvT2epZAkrtSJ4va5DtEMCc2Sf
KPcdqs7nqAAK1gkBRe68Qn+2cH4cIntPsG9fLjwwOeHYRXIA+imARgwrSedc
xtn/C+BL31dtOJsU2svSfBCA8SD/shNOOFHtsolL2/5zUBpEF13EAopfBpWs
WCeyzMWfVJWowof1k0h+EgUy91B3J8Z86QXijl6cuCP4/+A19WT3IHoBRfDv
NKn28LqVtm4CKoPA7qmOArO7VcjBq8VqPkC9G7o0ITa4JURAs/z7TIoL2Krj
ysGU+8m8I4ZSKlzrbiM2wmrutstMRN68ybQhkmV7ZPS4yTffqJrZbZeDrlUh
3qfVQFwHyqGUrjhuKVEvXSxaWjgRnkACv7u8Sxh5D26aM259L4AJD44jsFOb
TIJhV0grb2iKpv1gY3E2bbbpT4E3Jpm8V0GN648IjzKQ1Ap56igLlfiUevEt
sHF3u0hK4fInTSFyeG15SRnSxgGIFUVYvmqfJbYB/07yVYQrlfh7306wLY2B
Dsv5zCE7758VrOXH2w/DruWzA1JG5Ydd0JZkRuQL7m49aH76Av89MVT9vTtG
vIn7IYzjy60KpxHwWQMiOcKyGCCvsEmOpitu0WkfU7rV+7oMFKhKoGB2XMbB
vL/lBzcZke+w8uy2YQ2sRLzQVYIjAOfqpYf9BuTTj0KVhm5PPGPyFKMD6U4I
brIxKMwkN0F32vGS0DxpJez+U1YO81wevBgiFQNXvQF+6j/qClEZow1MpQB3
DY6OoLCgiZ1+ynElm2i4P9c3GavuL8iCGzVQesRc2b5xW37ismmtf9yu7W4y
9XJVHqF8pbcPPyQWV4xmwNUuiCmEp82rPD3Qlw2Uqlh4ZFwY+2A7Ali9yxcU
3UlASLpS/skZYq3aYt/kcLk8jEkemf1gdlJbE48kmYjTQbXGs5Tn01RugEvj
//aQ9+VDJj6Nk8rKClwOt6Hse67Uy+dEl+MMrxmIv4uQWD+S+hjI2D2zmIJC
W4Vr3XaE4v75L8mgLqTNJ9Oobt4pfLsPvbU6+MnG7R8pHeIWTJHstn16dmgJ
JKZAr5wqMmZnE+WBIZyRy0ZSJ/UQKDkOh1fmfiwh+fohV7m3MiUFZ03IybyB
StwWC91QOOOqH3HtwuoEZdnEqTgzdr80/bK/5fdZVsJ2WYTlozQMTvUDhIts
+yw7z+z14+eQuR5VX60alIo+tHNcsmczM9Yq5hfQTS4WvHmwAgFoItOEvSO5
Rdd5Yt6vIzFQ/be6GlSnV6AWylavMl3XHveC7bsatY7sW7lZUfLT0rFh0mdt
cMwYpXPyTOtzmqTJEJJH197BpzpCPj4YLd2dSyYRVriMMsWCqGg55Rz4mLWz
FP5f/aIpqrEs15UAFoe7G/jyO+X9R2Wc0ceSg/VJQTvoK7pSOvAf7fWTakR4
VgGWu/dFmu0eSChSJqVURKpG4Ki3o/Mwes7YiDh4cH29mFubt/TtoqxtMr0w
1EvWiuKgrp4p8ph5tJ4B0PiFB6I5mi76Q0U6YTPj/aozexi356RMES5Y2yov
fn5iY2YvEya9GyZg1tBAVOvGd4aZxUiz7J6T4WWxh2hsQkGcEQIucAw6kKOn
xDiAnm81aBOTVBPoc7t4QNrHX8XWqsuLBL2sPqAR90BYwkATVsYIweHgMQ1+
mEBDbfS+KqV7OLTYDATjAFQE7AEhRZwOZuE5tyrnPimw8OPhYVhu/PVKKrXf
EQbeOUf1dzpGSIcTsfi9hKBezTnCIy62GgmiqwTAQeIGDaPspaQZ+svZLC9J
/EXTaAyF4Npr5YGhYpaEsu44OCYo5o7hNu554nzqRzrE7AKm1JdF6eKiuMeq
kI+1aV49l1v8578Zaz/UIWFQ1xPdjyiKKLvWsHpO2nUr3Iy+Hx7X7Dw1gzfS
9aCNstsQ1qE21RypMypcfruUb0gItiwaVu1tSsJZjzFe+haRk4p5jROTSw59
rJokEiTmeH92zvaCx9Aik50N5uiILr3sc0/mrtiukO/mIypysLLbrjrWAlYU
mulrPl/2edrQo2pRnyJGEeBFpdieMjuI9I8A7cqmkgT3AhqRQOihd/1XZvl9
zI48KBQeBL0pBVttSZyidO0vcf2Wg01sku0gtXNQXkYA9xz+ZsMQsiGQsWu/
ar97ecA/E9Y7JUm3pnowY95JpyytCy3O3Bzou+ipOrjbyr/X/+2AU7+xJDpc
EDiXJiRS7UXerBNR2NlBJEsXX0kYD1b6VHm9fL2oz0aHvinHgF0LVSb/io+y
HjNDkmwYXHTGdOkgl2IZJGn7fPYHOTU8bhrJOGq3a1rNhb93JQyUQNCTrFqa
lWOijZDaWBVurEU3QC/QlfQC5jz4dSyL90/myguvE2ChVnidDjDsV8ziYJSQ
H7cSC7/ZocxEazEz7LAt3zKVCrNsHomtO2vzLWIqCLKSZVV86qgwp4PJZ93p
Jrz1xlN4bSn8KANq5k0Ys4TOQyffJootfxUGnpKf9M8wBgGUEXne6ViWhtVa
kkBY50eTCUWxBg8NBy2A2OzaBhxYQtfPnhOf/tQq4bHrGBIDP10FulfyS5Xj
e2BBML1Yk7/D1Wy2J+JhaLlB4QE0Lq6ppeq20t2/q7e3HCFPalm5dXVk0C2Y
JxspE2D/vtdPcWZSAGCObqR+N82J/mKgyJAnNHWcWq5knOQUYpEshmImK8gq
Mu2cmuGJMlwGNQQOG5gK+Tf+phVYbK+zHkrUyYqTRC5HWTWx0DnIGz9F1BaW
WxhCqudGA3118xb7pOaCIhrLKFeaDXRycxhhZHzzujE3z60+0BwaDEDGt5Rv
5eNQjekc/bWuktMpIEkxBC76q4GIgsZjBlrqh1XRXDKBJR+pzw3oSynzxwbm
O/U2Uce1NUfpjs6TWqk/UeBNLHE/wTc+fXOTeOnrMmcFMDksMl+yNz8QCYct
PGxXzvQVb/BXKF7G8lzPud59jwHg83Jnx4sbtd7A6irZFyIKWBFK946KhFd3
a9voXbKEBK4T4TEqk1NxfNtCgdcQvDlTfVnpwwxdCx/bgeNpiyw3c8Vv0aFE
T3qiexjBc/zSMM/PKfO74tIaCuoety0E9jQnMzqHUPs25DA3RVVn44ZdN5ne
mUVFhgit2ZNtJbMPp1msDXxyfHemYfaXJOh1mxU23AQBdD96yGyK1BL+aB40
biW54/X55ia2gYPlvQqu+h2b6B6GdaMy+zXcNGVGMGyx1YMPFiKABoylWJiZ
Hu3/e8i/D8OFo53gxRFtVWhDLgJutetzi8tgD5CA42GtXXJvnlSADZCq8kCQ
InC54qvFb00ZRuCT1IXU0lhXOGCWQY2KMBl9dNJcHrVt7d8+nU/k2ePyZ7Ub
e1loY1kW1LmDoFw2Ep/OmIoA7uFAOYhhmRhIyR57z/MFRFfYP/ap28ASdMSe
PkFOlSJTEUzppgqPawwV4HWINvg2NRTjoKboW1XBJ0ZR/kvbbaa2g0VLOcMV
IqMyI/FVU0p3uCSuf7QpkzAeCi7HsG4vQlsiZMsJ7h6AD7rJAk66P2S4oh1r
TM/a3rZDzh5BGWtskaSU8gNLvghvtB/kYEgupz6wSNJBD3/V42ZGIEMjHbXG
BQYDP9D9sFrnHA/OYphFHgeAq8rTDReh2r+73IoWVGdL5K2+1zSKJ5xL56ne
ZXIOv/QloselDXb4mdlVGrcULuiNrMI1QaXDEvueBGBW1vv2sCLZNkjTKnE7
jNh2W4lgKat8m0t+DA3A/qZx6AXzab042JZywXDs2SYtLWNVJAuDj7sd/lOd
Y47EVJt0pdBODapCvan1YwsmKt9h17xRcQmF/mACvdT9s2F48yJYLEMbu9bT
knRa6wX9aMxbC6Pp4EJPd7WeREhGROP4ZJp/ZpND6Rw6eOOMr8ihJBMfjMSl
HgLZYeSYidSUoSIyd6FL6rL+Vb0fX9DZJQalvGjBUC7mdly5RRvZEzr5SHUl
wnwYhqJl1Z6VeAc/Mv0/5Ks2pRz5QNij/8eGDQcoJXA8FfmZBYVLjwrEGkQt
WJEkOm/QEVj9Nmu5EF7m63OUxn98om2U8HfcupPP5QXYn2oZBpUmGYbBEmNC
kfo1FH8Dab34OLw3bWHv8w4Kex3W6As0PChPG3GkS1ehAZfvNET1QJ6AiMuK
gtIxRDs+qLLoCE5rEKnyc0EZVAGn/LLwYg1wazRmVdVmGeeu+qbwUJ61OFyq
QBmK6Eqhg3eqD682zYsYRXRoQpws5csyAWfsfKaU16dLpy6Z+8//Q2QoDVVK
lEMfDPqnJ9MYhsNu8c+ITr+AyD9O6IJmtHhKesLITSk+M3vlUZPpo7xB6e88
ftyzjXCu7hoUubQBct91ENeQn+c9SycFjYpJCR69lKPXxdx7HVXT0CWP8M2q
J6Zs+ohUhC7FZc3aaZkf8qTfW0xHrwQFdo3JmpDF/ghq5s2dnldXIn8oZ6BD
hjYLDol9Zdb5/PXhzzYTMlVEJBVV6kdIAJugy421fl21T/f9mbz+yT85rXXl
FXkdHNyG/x2dIL1MfwYktT3dcPdYoG5gs28MfHSVEGRKXESGax+RE0SMmKGj
+mbuecQTKpn98yr+dtI5WOdoZTH6zJ+RKCZsSH6pioFN6bUN2nwLTYqPW0oo
nqCCNYB7TX26vf9OvZN8k4CCTAl9sPqv3min9ZFyFIQmHfDYg15Ba6adPE5z
FWYrgkc+P7k2WM8nFnZHXaXUl2cbskOh4BCS4HQ+yBbSO77LRw0bf6C4/VD4
c0UCejH58aTShDlreE3KokXDO7ZjSN2uNaF6cCAZuSx+qifvpQmCuqNszHsz
DMrDVI6Pp4sXKvJz3oFpQCZgq55bZWF+05pViFbuYE12q+aZbYA9rTf+22W/
aqIWKxmT/CPF/cHNRJeqQYkFCIgMi3U9VwYsY3ApdLjcbf6DV5F4qBMtWYRJ
FkNAs9nUODfwptkPrjSnlkZAcdsqxQHkfZKxLB/1THa32qr9edgtuFso7nF/
O9KxsTkTtnEhBr3Nua/gopeV6hdzBSs6ExjTJH9rMuQW41hZimVQ7urWKaVK
Uwm3q2k3eTCQeR/vFHTQwlG7rl6NNyl+jwWDDzC1NyYwYvPcX+YNs+Qy8Di/
UfjqC6asM5L0nfjqByx+FvBPQbkG/IJk+RywQ53V8nT5pgLkunzY559aarV6
j8d7oXzyKp2KPCL5VFUzajbgYKwl6ZhBk0CC0md1YcfaTIrF5E41xAi+Xqjp
JpdB6WNXA0fe8Qmdm+TEGBZnzY+XegpzLam7v2VcYYnCN0SlCA4yq/cGHF1T
Cd1OyYJ48hplhqadrGomiFKWeJNsTHIaxL+1hzHoM7rY9eZM/rt5bvjOztRm
i3IuSQV/L39QJ2QSaT4e3JErrqkMQ8JCMMso9xFKDEVnrk2MgcTZTh8Fb/OL
PtW7Iu+PGVid45pxw2ANIFqwOAEZ+DkNbuq+ReYnFdjGtcH1s7EkF8oz6wCp
CRXM6JD0cEKs6k1gIv/O6mM2TWSYMG+FoRAAYHteQPBcabDQUOwX25gHs3r9
SUv/hJfVz3tIIlH1QN+HqFf12L+lm9m79MhI3M710FKyJZUTfcPlo26wIuTq
tqjes7GH5y/DCKsvsO6he75g7f6PwYp3+gvSoGiceh6oV+jyW0ansVJGNtor
2ok2leX4RANxCmEUEjoi3RzbGHVOqNNBElk5roFwVORmAx4ucgFmHdechr2F
6Ygj8OcRxSZ9Clx4F+j+xcdvsqbts2PHnpuDtl9+hE0TVFDB1F7yX29spAyI
kqq/nAAk4bsaGfEqA/rNmRj4lacqqX+RiMjSIANrFSFj/lg2qtXyli9tS2YW
ijbVU2bsJTXTMuP3OAGYXClxKk82XPIzy0w5REo3v0c4KzUD2rFicHC3NJNl
qlACYdgbnsTh3rHdFe78OBvinmiYIiWcrPa46PD1IfsgqvmJjX4CTWLggefZ
FjzcFu57LV6WdFHXA9+qB/s78I2KSO+m+awJ20CS/yyzxwGEGjwDbSmHNMJM
llnZ0DlbNenlJiI6BCcgb0gr6LLrrsj0kmbZdWiH9Hx3Td+iGKZl72reMPsg
jl2OlKsg3/P4fmXW4e9PnkOjkA2fHMrRuKYL8/R6oyrHxhkRCCfLsMsOdVyJ
7flZ7gE6fMkmTSR5C438oottFIm7DdCSYqJCt+7VEixTXufh0vw/XWczKGZt
fz6dW/8ou7pi4YfhL7t4i/dz7VN+QUP8l8gWOZ/cjuND/CrRcuWVw2T0+9SE
bFmv1CLABtpW7l8GsuqbHQpJky15EVNJP2CSHBmTgcv2sqA+ue66PsTwbMS0
Ia/o5uPEi8flYS1lJOmuqhCWxVswRvcWyqZCI4et0Yw5P8QMZs3Hcm91cKGc
YRnJPwqj9pqSEGQ0yq/udp7GU4MrbJ8ss5rfoInAOcbxtyu5puVdy6ixAG6W
tsTqBf7yduIx+pqIA9OeYIb/QhLiWLxQJKHbbM6ffGrtk3+/P96IyCvb+mMv
xJ2MJyy+RndFqjcc9xrOvX8EfTpvPnFRh9MOMomgOL3kN39+D3GXNqP7hw5U
c4N6xE5WckVMioNKERzkOQSaUxEnpJfl7XQWPRqTCFDnjHvhq89y7vvNuOF0
bBfMrFhSq7bmuSDg3RbfoDnZk0Jjp0ANnoJ5spL3Cecg+akU4da97Nwd965p
7FxE8xFgsco/ZgGmZ/h1KjDIKLM4yaJ73HvIgrewE+d6TcKJifmfCt4GMYo5
DCYotIzgak+tfDFkUbTzOg4ZMrcvH4H19YYctqA66iXh9jUKiC+BrlRBlQtH
dMlry78/iAEfBng1y66+7GJx0/Byofps1jWQCTH8zSTr1FIIrWI+YnEV/EtC
rwHtpiZ9XebzRIla7J9PktqLe1gDBJWdzCFUm2f+r/Z6xV2rB2LfeoppM16K
MSnToOlF6Zp80NwQ1Y2p55w/kwNwgDe9nFhrDBFRr16mHSbIw8gV96qyp8n1
QpdmwAXnivlGULwOTCug2Y91KojungRbEBaWGzru5Ri7uV1flvQbsmobgOKj
ITi8RjfW/mhYahMQoChx6XVDMJsKnR2+8v+whCdi8mI/vydM+86/nwWw2An/
2cBFx1I80gIs9iXBXosyrPwvYNY2omfToPa0zmsi94TSIyXVx7W+g0UOKx1L
WcxGt/GEdcyJeTov/KdjO6A/L1XLQleSkBx1Etjim9jYyL7m+k3n/921+Udn
dpwxzIjtBqIgSCBElgPp0S3CRU3DsFQg9KgFy4/RiJTS9nEx1ZwVWpJxfQ9X
v1UypOMnl2I9lwU/cGEXK4pDR+yT371yNGxnAs28o7JUywR0gn+rU+1HAQbT
JyCmNebsbdnvOPFRz8TcIfk7D04PGPlJoAt0BWjKsHVYeUlFNTlpLgyItN5T
sk1db8RhauRXOqjpoNHXepq4mdk+WXKShB8sTlM13d1MdUzsx+NpZ8zYbjkI
vaYISbUAk4MFFyjZjiwGmZJaLO59PN+0HcbZ8+mK4+/p9830VjyyHvolIY8J
ORTj32HFidOL3FPIMMcIFxpZsRCeO0nQ7KQoXyHlIbW6JF8JHabxwmbP+QGr
Ae65VFwiDiNjSxrFmJZTT9jHfIveSVGEzSp5HC6WV7tv05r8v1NxAtAZG23/
/J9BFdkrBhKkSiDveJdU0OVlbQLY5vem8+He2XaYxrXdur1F5k4qyvpczQEN
JKNXsQtvSteq6A0V+2kkHMp3ONwyLsr+evvMF/XCaZxuKHGp5fo4q+9pKFPT
IVtO+urdCh0nh3SMKwvXawiMDLLBEYhdJgHB8wT5tUqlOp4PgfD7yoKOgRfi
WEFaisR5QIYetuHmqC9fyamXSyYn6NbBzX4lRVUxHrcgOE3Ll0mHjfS+tSE9
j7LQzuc3gHZ/tb7aTkkcmo8TMVy/J2sf/vwOqz42Gc8TxRsZW1V4VwKoO3Pc
M1wGSd2vCGfUj3YoJc7yHFEoat77A7AehTxQRgOxiA/aADV452/Ci8NwjeqG
f8pJuogEeR3gtpparpq40K0f6x2xdumvESmuOh/G76t/dQSkANVIwvZtxFPF
qU7sxJRn8nXB2I6ryoZAV9tTv9fo+KQp+lus1ueStNFm2pCHROqqOssVAW41
nDpIxlmvH0GKbo4js6aaLswwT886xjPSx+rtq+W+NA8YnKmh6STRYw9eiqRO
iP3+kN5kClOPiMGvC0f4cHimJ6gKQdzaG+V4s82WUSDJsS4EpPZYGWPYNQaS
yn2IjQIR3j2tWtwDt9IZp72ZrVNCnmI1BDPopX8kwWyAzbNb5RjYICqysRzA
ljFvEYUrNBGN5p6ev9jyPr23oAkevc+9FHQoszLBOBZ+rSeEEEaaf8N6mCR1
rOjVWnGMSG2Dz2hCidHMe9PokVrFbvpU/Rv+OqMhXCIX2q4qyDakm1vXBIqT
Ook+z79TX0NYMGRGZKeNf8C4M25WlS9vI2GKjtSxiVzUdXjmuXYb5kbvPSNk
/NocYAlSTFbV3wPQpKZm39nfI3/YD/KUUReeOeR20tLtrGxTn1JfPuTO0+IB
TyweN0dsmbXGoUFgDLph371oFmkXMe3fij4Ri+b6n//BI43Cr8MtKuHni1wF
HgZLvWICCMnJi5ZxqVYwdmlKjqDg3HUWFlGOT20stiFOllmhBdVvSFk0i+w+
g1hkyPtTX3AJlZph8VKSFZtzCsJCK2xXgVs1C9B9xuLfGWMWIs4mcI9qOow+
2zXf+94F0shiB8zXbK8dVxt0H+/c/xZ7UYBkVqgorkrAckFrlF1hJOyYdwfw
Uw7sBL1kifxg0n77+t6MGIKnZmJ0OxMuHNBPoZbZ4xev0xMzP7OMD6etm2gb
PZjEl+nhRyXla8KTzMig6hqzV0erpJiE/38uuLFqA4XhE+gpv2FFyVtTs2zT
EIgovUWkGtipIFHDa0vEwa3Akmb+hGxfB5UN9bSNS4QYlYb2HqHOEwSRcEQ1
za762r7tYoGqH0Wsz6SplE+PeAwQWCDQgRvH9flZPE791mEcLQNH/rL3kg1+
+n+2F9E1IC7UaHPfvHLKaoL2WOPMs2tl98Fm4c2dpBWEDKJR8MdcNzU4OlHV
nngZnEP0iSZgSJDpYZhDfCuDuYiHD1tbBERXV1dGw6sxk84m1klXb2+avIWT
lfeXLcsTtEPUwYkMDj9ncyNxP2FvH/aGOqhOnBuBA6L88UuKS2qN4mWvKn9A
x/6LOTsOG6Vwq8wgynOc3D0iAiBP4KTs/LcMN5gNG4GJ2q5YJAQLXiD4kAKO
yNvHOcSXSJ2/lN/1xXMB7f7HjIkT6h45csnyAnYJL4ye/78rPt9jhB2hOx01
h5+Cq9jencQ4xC9oHhvRaMqoP4BmttA6DzJnYowRvE4GFeTqvTOLMs83ETxG
doVk36OTah+4mhRQDlm2GshRWU9h0bYDbtmpS/rl5+1flLabK+o2SfyQRbgI
uQLaAAd3tylt0qroDFVobW7GSn3IbAucHM6aT8MUEOJFcr368ouyXo6bqTYi
lCAcpMXCqs5aMBvb2dAt/lVuHpfhmcNe1cwnFLB23v4EDi83PXnWfz2DuLtF
2VN5htwEx8cVfKSFBzT1irWAETyFvGnl7lXjMxEmv7+J33p9ajuPifIyoPp8
lbtF40c3cf0VNL41FsjcgzujGXEe86UkPZ9Qi75ui2Cljbiq+XgK97BxOp8x
Z2LKciCxb2BtPrG8ujwQpinH/0ld4EyT4rrzMPljY79FGi05K+JqCjXCQJ7g
ZLp0Un+VmycVebK1/xPD9EFLLL8/3bYT8rDMK71F8zrgHVdvOr7mg+yHM5hH
G+GPJWkAwT2mT7MD0R1fGBqIQSlDfF6Yheq9LguL8N+rlYcXzp/iQMivw6Kk
FjxY3R0h3ZM1GLC6eHNgSx8XuAMAYd6/7ubT8H1CDNMRqUEDGdXxlfpT2eme
Rddg5c0f2Ne8rqPiNl9+8BIBi9/7RsO8MlhlhUXbEJjudqSOTyYlKmVE/P9W
CCX9yvZkoZr6vv9ooIp1UxA/WEi+O0exlvaqxtNxsUcXp9TA7vmoswME/Wc4
gFpl6/wtD2nkrRO7qkUhJ7pAatWOgraskP5Ejo2riVXg47p5zAV1EcKhAezR
cC/dWtDpc47PKhxJ5n50IKOZILm5EX/3aAYtDfBncRPQNl2pCfsuFXMP9olf
+0NMwbABjygRHvZ+5PooZXb2g8U3IUrHTdrOZcxGdN5yugEIB1qWPCizwAR/
+ReT5X+pghnebQZaFImxpfF2DKYpdR5fvf1isKybm4bQ/UpBNvIgGSmEx/ac
UGd/qd8Sfe01vWwXv+0oXAw1QQp23vZHYoxQ88pub+EYqu5NOnOU2Ic5QTY9
tlouTomEU0VHC1U1Z0TFvMu+liSF4qAYRX2LUjFT6/5wMRK3HbTfad52hhv7
Evw9kOGFGlwlP1HPQhPSPekDGochkMvmipbmiO2bY6k4LVh/x7UzEyuZgCYi
a7sAtLnfYS1nhZs5NId8EDHoS8Nvy1DwOupkHpL9/k+CNUHh6SjDhE2gTg2j
m79Q4K/Z1ByO1rqbSBMtXj6WwdIk5S6riPRG1/ytEy/EkCO5c0zrQHEW0oTt
fAqh2yOwCXLKPuoMldkUK3Nz+HnG6BMkLXVeiuwPx8wLQ95yruooiGKDEG95
XMQY560yLHXqj5/mGuYHdXTVVUrByhya/rjyqGDOxGaNJIerINst+X3criRu
lqNxVDRYezrAAVVZA2MMdYkqbqvjwttmXPRKG8wGrKEQGJZf6wBZmR0rEyKb
HjunWd/7jYT53xb+Dy8mRC9ibBaAbqOqug0aOH+/7DvQuoUiyLUIJux1z4NA
SjHS3NbX7s8Bf+T2UjDsPyB73HDBFuIzA3HNOe1n63pkcskkw1nKinDP9mcO
Rvz3P4z4WA2d7EywHZHpzMjF2sl7VOjNtCAKZo1cyn1p6RSlZRafGOpY/c4s
f0CE2QkFkzNDrXX4pbYUmUQP7zNbG38599py382elF9o12Yg1uMzEAWqErcu
H2hYagNchFn12HRb41MDGaKD+4LXTirjCEcgZc6XY4Dbq6kUEheq6Pxx3XHY
wd/MHAycFM8y2ELDdRLuiwt0qjn7A0j+V+Ov2/aUgTeD5B/DICK3Fea9/ziu
7s1AUT/NaVQ2uc8fq7gvM6MpDYWTvVndVrEsy2CUaN7p7tWXK3okImWE7BnZ
4mHR3KY42xW+SmLsCQw+miKDuc0LrBVhA67369SMSH5FKnNLe25FnXqtS5x8
M7Z7izgmRbyoBesNK0bhG5PpZTjKpwnZe9TiwvMb8t98TJOLIOPOtLdnIyzx
zeJXJ3Ju/g2mOr1EWjwfSiMx+7VgwpKmX2/XmuQmoF0axpf3h7vS7IuGal8Z
OMH7nHUfhj6p4enlThdu7WMVMS/bpq1Hc2ZDv6fIZCPpMGKkMsGLVaEsVCQw
Vd4yxVypxk1WBtAqCPv/vxlbVPybOhmVE7ilVdrBM6RpntUte0JJNsveR4cj
q8ZNut20J3fVP5PVW3gqa9MilXZMKA5nCAeI0zmrBoC3tNQYxmbKUpbcVQrw
YSUcbFZp/xI+f/XmfRSo3o1K6WYsg1DSRRUXlYSrHWjGqAW+AY0BiEIGvxse
x/bdYSCj8/3qAst0C4pdyN/SiumGbxoOm6d3eeRD/ZpKv4XFJ311qlhpnl+d
hPyGei8ngP4YAoO9Teqt6J+Gfx1kbvyKR+NPFKT6fUEfZq2aDnMqSMAQKQl+
CR6A0d+LQbzhIuO7BVnaJx3CW2Q+43Q7BmZ3m2fK9talZzFPeGKikzxZXfWy
rB0fuS4UEJGrBr9OjCEExI3Fomzs6aCIB0NL+bmwUqRB0GlEoxQM0WNY4jgg
MLxY8b53qtYGNG1fS1fCdOIzuxGqrHBBmzg9WIY9afhkct1C8VN8cTSYpoTh
IB+FePLOQQbrzm4Wfg3bfsboNPC2EtdZmWxXczUfIja3515ci8qwb+GjXkUV
TJzwRnMJCDd5RgX1d3Y8gvebbZikbjlg1mWYqEZNO+AGi6TXQLexm7x0CWAh
A3EAY/TH6k5l11T0ZY6qlCvVMzF1XtwQZ9c70rL+tlbwNJqNi/T8i20pRBMM
3vX0OrdFsh1IpS+StDcjrZuEJakhAt4/FT7PuXGpk8HlFC5XX/ijv5ouxCon
6dNo6swHmZZlrY9Bb/p94xL9C0LewXlG/vDOslikUL6s8OudM9/haFpT9VgI
aBGPJALF5fLDqAlpr54hU8VN1j/av/SQiDUIAiFo967q8gtYFKT1zmDIQnUL
Yg4ZzaqxQm/WdmNN0H84IJRbe2HTBGMDjA4hCCZYxVp3nJ9lcbGKQuY4Ilwp
NeQ2bel0PKYxCzGetom6drEJiyjZMbTjVEKoAKCFATRsDmXqa/rdchrxQaVX
LuDre7ISlaDrTEEkRXxbV0liDVWbZ6cNwH9SEQ65fb8RPSl66yuMAXBHXqMD
mXwoQytCI4wFLtBy0AT+D7it7QNRuIf4N+wL3PmarpXxm9I+mVEOKbroLFF0
yuP+I4xveyuIqu0LJK0zPxwUlD1O4XrKpQtGP2kNdPEkD2SrIg0W1rR1LQMa
Z1PdKOGZt45WGzepwWc5Yn5/9iqug56txSYLEYDd/i4vOTlHTWTm947jZC98
V41fk/h52DkBM9lWNOdS0MbfD/9zqvCoqGyHA1AlZ5NdIq0j6kgFmelYgh1Z
/ccbgJ0yONteCfTya+1olSZfL9Fl68DAJMIL5MDJHI48r9ao/uhWGamiJxMX
kNKuVbp11FquFmkVXHfhJJWN6rSXlGqtAWZIbGvXszMsbQiwKo0T0Iyfsc8D
SDY991jAmCCdH5BZ8i3NTZRfNf/CrbEiv/yf6fId1UhRz7+L/MJmLMNUwSXy
m7Gcp0Waq3mS8/bbtZEkuFpcVhg8BlSRYMNYiQdvXBYqtL7bC+ArtMtBZuck
HyNm+PWilpowLqhVNO4qQY68jUDFMHo2ANqOXMcUQC6+D0KLJtESmexdJDGZ
aDHxmmOw3b0ln+9Psle9P7L+7kkue5T2l9E3fdzhLK1hIPgLhStMXZlTx2J6
8xoZXG+6HIlssUNvYrODEveMgHk6UHyZUi82Ru3v4G3/CO6su4h5/KCKmDdx
anaPBzqYqTT463QJctdj1aW3xoL0I9+UA1AZUzvzbVKklgEC2SbH2YAM4n2n
zWBz38eM/xTsMNP6Kq8Ns4A7yj1w69fW0zlXCJd7hw9L1nalKgQjjVhWpfWv
M+J/QpQtn4tqVLm10lA6BOqUDfFQRjinVVgfzdxNt+wU4QSpxSrb++YRxTa/
CV7n2PSUnJa+xNBMETR0qEUjHLDw1XiRnos3VxafuS85y/pSRnDX5PkhEALk
22F46u7kzW8VUG7ZAQIo4ka6xT+9tOF9fhMoCalM15iTiD4no51EPlvtx1R2
hgSI41YD2ij7K08wTsIIIX1tiHU2pXO64qm5sJ83qOOMXhP8tyJlF1DTn4wi
MzPiplS6fCdhVhkaPshzDNrrepBp5e2Q0H+rKXc2NrIp46tPSPaAsy917gq0
XK6YjCkT8PzfseOUaQwfYG6/mbs+Gqpp9c9SIdE6tvdzOiQ+xc/TINKTYNcr
OB5rztYFk7CgXlQ85vYvsE9RawayU7KmO7gbmJ/lYElJm6eKDcCFc+VajEhb
dRsuOQ++P62pVn4LMyHzM/m4/eGR8OYK0xHMZhS0OJIfuUOnV6+NaM99KohX
Ukp+vzcn4KlVXwpxPJwPIIe+i9lDByCQPBqgsvU6fAYmjPh6X+9KG+4Bxun/
E+zt/FWnKyKRtxandLU35prIyQwNDFU33P8FagudOWKXhjJzJvQScQ9hYff4
aKDAk7jRzqwSYGKsivVYKJn6jXvc1yqo+QC3BVzGu6e1Px/0Hdy6/AWypj5J
4LOE2IXwVZIzBlGeWtRPr3WvHQWgVXjyyQ87F0QCCwr9gyHy776iKojxqJd1
gMXpfNtFj19AF7NR5c+3d6S0gnvUjlETNjKcKQ+iseKqRKnkM2iWhXEfOCMq
nUFZ9mFGh6hIMDj5KGnFkXoyEJ7LPMxcXzmpvP2c+kaNjIKhm///wBDeZPS4
VN8wXE6rkyqJabwyzIy4StpnNL4If2bcW83ijGsC5X+IuKDkBKjk82KNDwue
qKLNmRrN7n0GQJPdn1PsgdnYVhREWd8ksGWVUMYgiR0ikd+Kvu6eQXkNgbxU
umtJKuVIUDxp8B08kGrmw+f1Of+z7+5W7rwx2rlGz8Kr/Hry5mvRjmTISKoj
/Pljt2ceCD5pshOew2CSXg/FTpUVc9igYriMwAX13YMF3WNGuxIF1YnYbSBv
GhuIWnhRS7dOPYCt2kaADafePTX4Nii2Bumck6/DpBMrXNuG3sayKWJlhNbZ
HxWwwZi4oHAKEfyI/ak8BuIH+5oKkkRAML1FM5fgWM90Uc/lDjqZt/3fIgol
EqDX9Ry2L2nZTKzffYOQ5YUANPH68R0hPZsFxpv4DPhHDMcrUq1dXf4ibgza
Le6IaFQvf/Pd42kd9nUEHvEErtkihSzjWwt8o/Mn75yaUtto0ugkJ4E7j7yL
mU69xpu3ogarev1+37ZwteLw/JsaHZx6vrAFxgEyOdlZibYCbbCZkGdbYlIz
KY9v/9r4exMcEMsXrjbj6V07NWj/7DJT4K7EE8Z8idgx6R+w7CjnzpDdD+QZ
dzebyGS4ektnycEKXmKtetDl2sDmTaJ+yxLtP1QehqDstyAtFi16ZVGMDBVP
blNmjcUAE2pE56y661e+A+AfrrFeVkfqfW6+/JWtoPR+V9Wh3Y6KOlHmgt0r
q0Rz/k0Hv/puAuVFHVsE6e6aDXeBPaJAHrL9O1Q+mGGym+6spWNswegxONVf
M6HMtrpMCpdoINUEZWq9D47ZHs9V71AZkoZ/4RRGS9QM1p65R4/2c6MQAAcl
40zuM5sJ6lc5BjpGn081rS4cY3meX2YUEwLlVhTlXgJFv3mxyQ5dhV5OSZwM
94UegV4B5GKGWvxHncQpEtt4RlupaqXQTO0HQ++/zR+II9e7xRRJPingGCj9
HEcvSqkyvw9qHa18a53MtuVUPNYG3VxL+DprsgkaHaduQJxqlpCwOb6qBZwz
sPOgu/BEPA1auE0iU/rHWnYlWFnVBE5WxKhgRrDxPd+iGs2/omXN86eJB2Vt
1rjbU+LPzjvo4AVmp4dIzpZiUOsP3oMRwlcy+lmS8BMVehWonhwKWTqZOiKk
mG2JVsP/knMiNsfaWHGLQ+Lakf+4qnMfIUTBzQ8XoAQIeXgXKjq16hen1+29
tojYnA0PTkXT5muCuAZuIEHrYG1crlPGag23ApM6R6OufleRbi9mt+OjkfNQ
nXBXi318/pKdW4XjAgO9GJ3rS63WBMV023cFWdG3V01wHmfJ3rO27fXpLYsV
y+CA7u1mT2pcUUcaZiRjA56QsAsgomu5fF4p+Ntv8niGf077FYVoKgvy3bav
xb4np8mT1PVqkX0Jimeu1lUgnUL+e1eMVHpyrA8v39W+P60ragqrO02rfQ/m
R6dhele0iqcjiz/emP8lxj/RzFSXKOIg692epNgqELv/V65rUDvhpANFX0wb
8ugS/yxPxjAd3n9SpynnsBfxPaBe7feyklE+n5UvTHzPkfj/kiU+IhhN4kSL
X+6BD1cji4vSi6tB0nDdjHL0l6oc4J9/ctfVq19IDEE3HM+QrSMFDGhnMlSx
nkuSJQ/sHB14mUIbQnvRsd4RduDwX5odk1ELyy0x9F2jbKLgxcxN9q0vFaRr
zszbDOXIFu7ysYQkHWaEePrVJixGpj/xP2CeV8yeQm6rT3BkzvRlBnzT9FwP
L5Wy0KXu377i+2GS7wiYs8YR5nZq/MmJvKpF2NeKiieVD/hzH7FUdj6CwBIo
vkPXGwU9Do63ZpbCXtIpvFrzoai5owtMIa0gsgnukC0XuVaYj8JLGTJMsXf2
G/f3WJIVfUJIfBccokQhJnYn5GqFLw65Qc88YwJBumGPfnysOupVgsUnkOhq
JabqB4Z7E+evilJWthlFmIXyqsDo4i0LPUqrlOH0Awrr8wLjxcfEjOIxBfyn
3h0GO7fTLVOMt1UwSeqU6ooRnkUqnalWO25bicjiL1MK6cESgTZlmiiIBNpZ
mKFbqlPDkvqu3FD5yPfXMf/kSSf2lA8L6Dx9FhM4bXmpWTER5M/ZSzTgtnyf
mbD6HpIFFp0Y+/r5jbj+ONBzHce/LKBOn0++D5yWmRSGen6p6bWImxqn+ZPK
uEXptF1lcD8k4oQQwslgVe7NTd8jR1Fa2tjOkTEeO7IQg4pGosOSSrHgdoB/
EfDVpmOhYCfE8869UccrG31PwOwL9RVKmnRFIE1QZVqXZTaAl+rm6lE3Bkih
hMb4rC29SI8zxEAGw6cr8wTCylahftaRC68aWMaq8S+mXILgPD8W2xpB8dWl
FSiOTmgzwvRfITx6jcoeKhJ72rNNSJuoHegsodCSvXPeZW1yViMs87pDwJEd
YiJ8ji2fN+afc5DQHvm3sqrLlyohSxTaC/0rVjuMqvV1xHljUaeVO08JNW13
ov59tYIuOf1tgxRPAXH7bO44bujjrATPXFNr/jCZtSME9MQ3Am7sIe14AzxE
fQS7TtM+6TQOa8OBjyJFNITBIU65nMwrW5pjJJI5TtdoUIXqlXKkRqbwDZLU
b/xbQzOU+oQsPLjyrh+7bXYXzLLXAjmApPkTUekSrjdnAoqUw/9l41JDfdPn
sSK4s4wWYyPNdLqZHpPWrEraTbAqav9MgHoSOjFY2hxyqKmSfHVrdmKeXTeC
UF9XjhkkS1B/D2kMZqd3Mte1kJDB7YIDH7oYGgmqi78A6MhMHCjs+nHvDKlw
Zf7kTVBQvhktHK+8X8Gjh+wUVoxX3q7etKHVaLuRJTML2lN4btu7aEuaeKzi
lHsJCpio+F7lTK69SZvupyzvBIglGUQaF8pGRgq2Z3OazbpzL1r/PaPN2/vk
qjmKl2rzVXeFxpKw37xFy5nEcLXcpo8BE2jd3DT88iAwFbnu2yxEWssyB+Vs
xio6UvfjsXboroHIuuFirN9qttQeMkPZ1iRiQnudug8wrg/p6N5Rxe7I3qPY
Kb5jey6GO3xIFFQdgYGuA1uevybzIThGG05xFMNNMEMbcEKLOWJhlc4S1+AO
sDfMTJRzdDCytbxYorFnWfqkPRZYVii++8pGbLfS/B9vwCLBtY1HJM8xfRSy
JzY+aw961aMr6bfo1uXr0LyyD2TGfYPJWRV6JKbqbyzDXjW2I1750184IoJr
yH05VzmF1jeXaCzH9FDzDzlxpSLPIqvH8fdihR1DTFySK/9SeV8UAut6Dqlk
R4eQhr6y92oZatoiJMlhaC8PE88v3U9hJBG2pjMdE2SJ6KQ4zl/CuVse4Llz
OTSKmPOBXE43+5A4Kvh/N3PUQPB7F5HVKkuoPaZ5+Qwez98y827C3RYTRZZT
J6avSv3/nfFTiznr7NnlUZoG/Wo8RuTjMwEKuIaMMiVzhU3o9XaRjnVh4Py4
5zUY802B/zw3/4zJJ6RKfAUjR0UQKFlmKDl5u6hYGidZxcl7Naz24g2j+Zjh
b27v1VgxwxjJ9J22RYtfwupwsOBuExWt+c4F+7V6Ung2vOQo2AmKxKA3d5j+
IJj7aPTbwKSUdCD3XeIk9VtsiDl7gMzz6XkrmrqPo3zPkGb3SKgKgpkYiVLh
hYuWixEl0RtPTv5nekenNoLoGioivX6C2GbK2rbV1XmXGJ3OJUuAziupmVGs
XEQHavRIclaSakaKtxf3mswYp5SQRr9qT6+1U5gFNR8qz8WLjK36E/TU3wjU
/a2WNg3hgbYO//NiZc70H2GdZejaytJhlJ31bJ+GqV8mGB+n5RhXbdgJHUgW
TSMnyKjOYgoVOoxn0OW4YTB7mfdM34DViQFtG4ONw3T6YqPokBkT55bqHfhI
QMz/xA4Yk+2ZeEIOIJk6fGZV/Wb2XMc/FeSHnxHo6mxlTvIelt5eMmO04MSQ
oHJ4E7yS5aXaWux1gZXRbJYzs+gvr4A82u3RJyWn2EDwzwoXW0dK5Jk5D2ue
BIerh7QLwuJtBF97ZbfxEvin3ImH1lwaqXTWFUm6+jz1kVHiAlLDHHYWD7Et
73jeTDPNHNNjARCbvfyaphex5bjh6GUX5DGRTeukryc5hYkhyPCYeGGH+WcC
/9tJBNNQm0wc47527agPnKmkf002sXKRQ/0VmIGKeT2CJIpoLtQPVxFVA5WP
uCUOaVWEf6nNdSwIex40/vuRl7yW6CKQH3g+3Y3hof81Y+1C8BYcsXroa0oe
Sj+mG2pFLdNTsXnYCxWA9W832A8EpDxLKA1ryZPvPzg1uDoVEzkIZHl/dJZD
EvOm9kKmLLiaQTKl1UIiDNVrVc4Kl6IrYsF2MUQua01Tm4uaDR4nFKNoU4ki
B/tHM5xnAxIhq1JcNB3/EexEod1Oqfni8r+WxisfLEpms/HEjt1p5HN4Rsly
kf8Vq/RPkQYl/FiCgE6tXsuaRoipazKlNvxQuufGrZgGvQp0qA+fAr5EXmYG
7Bn9yiu2Zqls0cIvNWk6Jj8Vx/KxRQTkvJAAef1GKpeFYWZidllyAVTKM4TI
xUGwHuoFMxobiCsO61/DEMEC8obQX7hbTTCk7pcMPi04cPp90kDDKqfZfQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Eq3BLFKKEgzQT20LWMYCAU6By/LyREMHCLEH/WL2f2MPkWF0VBkqNemI9VlUH5iWX4IURFlyVmIh5E/HQ/os9bJkSpgbrVRO/lhtwMTF/bsaLrUVm0P5/lyoif1rLBuP54PPIELikdE27b7yZS4Uq/ID+UoTWCUtIdcAM4ss5e/TepriEbKaqE/TJe9aYE5a12U29YdxwgXwFDGIzf7pALYcBa7Anu/qCgVgGoVZyzuw3u8TfSgMbCrxk1Su/fVdDAvABHVV4xM4rpIYpSMHcMPpls2SuHSaTZ7/0HUR9LKIcA9Zmqg8el3CrEmr/chw7TfHXv61vOOjFI1/X6bW/eaXadrLODkQw5ztCmGmTRiEqB0mR1xzOh1+DoDE2325XhiRUA+Q2O7LWFHSy/eNwZpPWEANi5ygnIoG5VGjXP1YywHFX9cxfLlVTuLNSzyMujZve/krz0OwR6DT0ILNEDz/3HBH18g/51Ey4RyJ8GUNWnnZ3vEE4O26+OkLKqDXFRITuf/9z2zVIpVhtuW5ygpxeK8aKOOSNel4BZpe43OyGXKtXaokvqkyZRk61qRT2zlEEK2zv0q9HraXflQus6rBVBPYdVzco1z2Ewp3v9X5zoJBuXJMC3hrqvLP5esrtZsqborf41RWTS4H8eGPE8qE5wiHQKgsz4C+OCA6cx/yK6BIV5BU3hG15/kn+8MSiZqy/XSIEZ9QNPtwCPsZ5o0OrAnkpAjeqoJ0r64zu5La6sQB4n6HccUrFGUfTaEmqSbvaUd9sMCv7ioFFERDgnv"
`endif