// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
X5lWkKIY2KrreQkGVkLiGM257WCHDb9qtz5vuwb9dKw3H0Cz+qSGoiV+cJuq
c0fYjagBYxKg5y2eEsMjBtRTxQbQQkBVu+tWppjn42ADj6PP1BwIoTApyoYX
M/CU/wKQYoh9qBFS0Ewh/DDavT31QrTIq/vIlAqLSnZoHMSNt4OhRLd/OudF
EXDlkW2k4289Q0IT28xOEoE2nmdNb2GB5spVPDI4pZWsBxGCYMR/NRI8/Yd5
oBRdpVeXld2QgIwD7Ny5yR0hRkF5nU4K0DaCjkwccwjUdwtTpyA1vfo8v7tG
2/+7cjFH0gR216lCo/+rb2ACK5QzS63ZfLgyIwdh0g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ahPSM2Jjgogf28YSEB6S9OlSPFx8iWVBhcw8sqEPvtUZPlOWDRGDnsAVIxkB
W2Uu1UXBqERUpzOKDyYVMQ3exFUbkRtB4K09WT0xT5rLxWraOryBnuqudTBC
Rm2SS8lMSmbMa/aNglTcXVKhQ0XVii2wViqSzpzrIOPaXFddDS/4qiJ1PPyj
gbxm9y28xg5Ztf6SZJjpfP0PUvJ1FnszzqqlrH0Na/0wTHUs4XOIrTTmnuWa
f0DBVJ4t3yNu3DiI4R88hGJgNS1z4BWSre4QbIdUBkre10P6hOvs7SU11cbF
K51ohu8PN9NIi2HXABumG43EcsbN2kt0OclJlzDDEw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
q9Te8HcoFuy3YXrMhCHtP8SmdOIbkoZ+9+AvbipNdBI7JvukNsBZc878O5k5
3xQAaUdsVZT3ky/ETa4Ac3kIYcA7HBss20srnRf0KoXrzyi65F3zfAg8+Cdv
vGmgo8Dp5jhp6ZWh5YW3nW7BdmNEp+mu12IczqJlW+qMqykMZEds8Rhh3Uqx
C0LQXBm82NSyb8siuZlPq3KgT6zQF5cFaWEaONwEJ3nLHnd92l1kVnr6nnPT
jM5KreCVYgmcIgXA/oJJaBGrApk/Qwbn94uSyAAJKqr2HEEWvG3XHRJ5PH6G
e5Rf1DCQDvbsFPr0Vru3Utbp+U9zafvSvFPusmNOhQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BiJvUPz/jNkoV+uuLGwUJwvvT7tpnwDHiCS3t4RcNXH1WXl15pVWN/qCUEqI
eX+Rw4y8WVRJzj6c1mvj6MPqLcz9ywKrhnWkodejE6fz7HhY2VCw9F8uqwqI
p7qr7yb7R6rz6L49K2Z3Y/mAhcBCxCZT7VbN8a4KO/7cMBQ9yhoJU11DVD+R
miBNe1Ou9s098uqqmmTVEnnBLqRi6yFyf/NIBgBmJwg6QomzWJcqilIKBFJD
EF1brybvjs4CGZg0vf5vCR7k8Anm74gIM/SJ8nf50ROJUGz2VceZuWfn/DtE
T43+72qsCqhE85A5X8WNxQUef3CCqid5THMg+y/wCg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
s2WilCBh6EqibUwzbWL81DowLx7w8TUP9S9UVA8u4pFm3ss3UC7PQWX1YSc5
extNjg4/kuL097h4cPUz4rQhhg1EarkXEeakH5bPUYY0jia6XIARyBKNe9kS
Zf2UA5ajVTNQ37eDMbC7yBJp8iRWwVZ9/cXqeMY+V9lrxpGyE2w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JJVfCon96/qIBQBuCSN7FseCw/ISRUZscPRtbLOV12XLgHkzsAgh7DD7jiDL
wlLckFJzmSTf8ngBZ2jfiOfDqfTJjaVtxhQP5/VGQ/MO/gCQ5fURZJ8YV4sp
pJJL9zaUpgI2EBnH3t0HEBYR4rah1oP8WvYjbnW60Ci9+bLVxfKOmlBoMIvP
e8RqGt5SpRC+awVl2perUj8Dk139Abq9huxe1fxnvaj4EntxBu14Opiz1omd
uHt5/8QYH4X+OhQTK2u52SeX4RmeEPkF/BiqR1jEvCZilq8k0wlT5twPqJ1S
ZH6iP6AZ/MkptvuhjjmANBc5zp/HgQXWsrTk4ylc2RhMKBoAggMfSRQN9lIz
bBAEOPaEoFeYs5RXjEbkvxK4UDd+uuBZQk67swCQhJSrPk1j0/rm5VlgKSct
DZ2shC3SnwCn5zJgJUlMcnsNRWSekO6GUvGIrM7tFq+HhMXxZgo8WkIi/9xZ
96e9qjNjCrzZ78ysyepECZhq9izUS/z4


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YyVneFXAVdW+JDZWdJ4Ag7ZvT5C3DtBV6JCmtRdppgrZNEGO11+nRgdjLH07
60MxiBOr0k6H6v1oF64y7+1xNoPXNA3pCa3y9ekhhevRBJGb2UDXna8mQJaI
LyGygpRqOjJ9iAL4nDS5P0NACjIXI10RuXzWlODdmFW07Xfjhw4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AGPb4JC0NZjlrYNABfHqDozAzn3pQogj85qhQLdfYxeE2hEfAQTAu0sawZr4
fq8Z4EMqzEP/LLnKjDryKJnzXjQTmXMidL+yFM+Cse1u49cQzzHdCuF+/gDp
4ksJcpwG3z+41cuscsgrv1+9Mekk/hCXfFYMohCLkF03EVSqCGM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7904)
`pragma protect data_block
S4QE4s8zLcCDQkhc67KrCa/uXenmBwjPfQH0+eEq52Soh7EWOsI6Pf3pyWDc
LoC8YkTiMFGyKKJI8TZoUfXxAm6a5yjpI4D+oWWG8GVHBSBYjr2s0Bt5Kaqs
+o0r0nptqwIj+DvcsaCwGfcxZB74BgqYcw37aLwgiejF6BC5LiB6+5SXIkJW
8pkWyb+FN+Rl1jS02E8DqgkiDM205Y7e2qEFRz4O22jMPstBZSaDl0jtOlgL
kAolOIEpkKoWVuKQavjgqnc2WE07ZonoWt++SNAjyWqDDWBj/tf66/Icd7PY
Axzn033jVnhQtGbTVbbTpgB/rXj2pq9uaCjXqbeYbzaLgbGJJRLP/aXMNBgn
AxKcx1koBJ1TxSXatcfqHo0WeMDoXPzt/4X8QyRzXJ+8zfKPxS+Nol4QjlfJ
y6FzRozLIaHf1AYvXwhnDxSz7rNzh1vTkc0jdnMoCPE6PiGfMFCMU/UFE5HQ
bjcXT3CUx3abwnJUSQtjqbLhIZKH2eodARtgNjt6rGtBKsHQ7OpebWvePVT5
PdRTpDCAkfCM/dLMbG5raFw0vNTfy/6lA4bttVByHFgEGWfaFaCndbIjj01y
Y1HF1kfIEyu7PeXpYkfNZuo2glcFplBsyabMnFYRCHOPcKO9ort2s0C6I04D
W6UGQw/02rSrN38VMGngkEL0/JIa4Y18cSPt9fiESLlIHH5xkItFNDYEgA3x
oBBThla0MvKAbXfQXTGpvj6hsj1kL5jteBrpHH7hvLYmi7cR3Zi4KQtJBNUk
1S/6yYazzBzJHmmdGto9JLb1R70qpISmsQ7eWd2gO2VZo2b5fjBiNM0r8/4J
erxBc8r/3YUuFoaFPoYn8rOJNcOswzHAIS+ViIFhcr4vgbx2Wcvj3QFkHKeN
wV2Zme7dP+/0TQwmBcIFhWrM3g77Jk+uBsNS6LLnz8DMn3bX/Wu4SYHnrx+s
27/7sJMyVju8HOdiYNpe+XxletMpy/mkZrcI2tJ+q1HWyHJwhgFphyiZ4gDC
D0jP/zpePZvv5xKuZQrbvYxvYFCOCuV8JRLjFHFna7OIhWC8zlrOlrbkNOuW
Lu+UqE6cw4DGY5UphGpwU+6I2Ny7Ud2K4BybuZNAaJEjhMNqkAUbEdp/t1Sx
++Iw5TF866jumdaaPG0UavXYfpME991bJowCMGk3fpQWQSQKa9X7oQr6THO8
BvLdTd64f27wC4qfTxOf5J8Bsl5h/ygLwBLzjgjqnI9zlXcQQf68ILMf2gG+
sRhbJSYzOnNHpmJ1n/r2fG5ehQmPf+ir+Jf4P9Dae/VBOoHcarPcadbzym2H
asz51EShm4FyRB1RvjYPRTI2NgMJTOKFpD0H4ggIWzSghjSqQ5okyHu21cEz
jRFYY1nyMcoedTpwo/exvB2LkWvTttbTjTXm4EpqQoEwDDFbH8JYmSP9FJPN
302NyMrXvupcZv48bfW+MmMawwulXkpR8pdC06se6FCLTSrq4KhqELloFdvM
U3Na2mJdMH1VQ+r2zUrcFqq2q+ash8pbnaXN1SbPg286xU2W2VOSETHvqtMp
FmC/zb2xj2lw5EGb7LKCsix7ynvXOryAp4oZfiISXJQQgUSOtYUCeDYYBhI5
QNFQJSGO9CoUrW8Sh/dy5QO0B5XbitdlY/BBSJ6LJQA8dnRClWhCnGi66Trd
PVvbBV30g1W3AM1rXILVKYZUWkns1mkCgyLkxHMNPsucHKJ/BkyQKWOV67OX
/af3jd20kJr4IH4M2mdBQjrjUQczsM1cFkgMFgjUIg6BScokiFwFvcSxkhh+
6Bzr1lZS90qI5SIft0j6pw1vGoCwIOiRxp/yTg+aTBGwBK97gVXXzZBlbyYv
5sUB+tNaAWHyK++36lvzeJSTg1graueZX2nyU+HBpicUnFcMFEncIwpL9rFx
s9nL348sIFCVM5dVSKuj6Kcs5ogH2Uhj0BqjjVwrzwn2e+id7BGhIHXOZ7VQ
mNcIv6Ok1vrSwudtDv3m+DMnzqYQyWrL2rIFiGi/sRRJ9nrLGWcsZCiDabxu
iBjs+YfkA3TV5/nA/n6afmhpUWNnCiFBwvY/c7VEDHaiu6GgMHZken6pujqD
ouS4x/iawKuIPxkE57zKRdH9DZvS1DxtrTRzbUmx3pym2mdk2WF0azWmYrkN
YGLI0ZQod0k7faSW/3Eh8fGcD4BA1CF6Almh+CAbHhXWGeOaWdIpd4EA86jX
QZ155uIQtB9hFcelvoWsypUy4xsi+Khk5hIs6cGE0q8N1poY0JveQFoTU2U/
DTVvunw9C8Z2D2XvMSepkFPVaMe1JbKkPznCTwR359GMvZX6a2RADbNGZ+hy
/wQ1dcfpkoMzwZuKouBFEM9guH2WFpLYwfGRlewd9ZY7/msjaUg3e+LHW9Lh
tZ/O5Wcn3EOitMfmnWTPCih4u5ASKx6m9jcNseIcfHRYputI7qE6+KMhjCAe
o2COgiBWYFa5IraV72no/KdWwuhBGzm9+w4dXSW4jq9cualUXM0bFAxCLZHj
VZzt01deE4Q74/RyJEypI+26hd4NzBFZ/LoQKt+8jZ4YX9Zy8UV/R9Hha+A9
w2njg5FlEexnqFJoeQpKs+sRbSCcqNQ9AMLBgvSsj/WH4G1VWo3G4NN45fAT
GfEGdaRi3BAQkhOFR1YhYr9RGupeIIkoqvkHqp1vSXiHlppecN1Sz6olJYPK
iMmxMFzBCf4cuLt/PJvIhPSyKNi3Y304Yzf7DxwD7At3aVidQhavL92sxsDU
RGXKT/Px+pTlDkbI9K5xiUHtIPM8pQwFTV9oG8+x4GjzwdwfrYgJT3WDrwKc
Oz28ehspXDFFdkX4YFIdnyMa2kmmVY9NdgCQO0Bc+EFQeqqj0kL6wwys1oKk
znHL57dhUG389udONcua4PO6J9JkLEw0PaLOhZtvP0YzKzNtdA6wAj7Ytlaa
UFZU2szdaKRZcpBjLN5ROfPEvYmYbuq+xtuKa/XA7zo7erNoa+/SF5noig/k
6SglhO7x6z0cL9TNgyfdQr175eQ1gs9AUuiCBxdd/amWDSKUZDFKR4o0nhNE
yTXVrcJb1VqOtaq2KoH1EP3DGfdIv35uogp6gF+Uw8XDYP8W4nCle8zsKeMB
+DbiT1kP55EG9x8nP7k16XyCDPvOSHBtlFdSRMqdHXxv2gjxuF86J9/gMzQo
V01acEgQRG2180w8FbiJPW0TiXD3pFR0qeWBci8VMPeU3THlcbK4iQE1z2TM
ynFpsxFLrU6wULJO3qErMASdt/KX57tBGRYblkx8Lar6L0dISbTkjpbJ3lWo
XawFnnAob8EyqgR8IcGCk+QbdpUBTxR1YAOO+YUAlUbndHN/LM4KLM2wELa7
8et9dz1qThQrYXUSxuOI58MarLt7z8fjLTphdvVrHMG/AtMqV/Y6ssGtQ9Va
b1EAcG9AJPO3xw8JvGqKxWLlfb6Yu41jru5bz4FNnD4taDd9k7fIntA6wPM2
DzsqjH2OVP1MCVCn2UUGs3ngyHs95cQKbNeJe/yt2nABxezY9iBM7Bz+vi2I
0ycO1G+JIJillCAMvpYOpNbPgPpIirogYVHe3BoUlAy+n4vYkc0t7rQNEvyr
eTxn0HzZ+NHaoB1OmM+EludaRW/IEfTQ5owC9Q6bkpoFK9cyb1y7hKk7YmuV
5jWKf2MuQ0n8kYUA+EGZswxt2UWsbHZlIAKpx7pw+CDv/E0tEpv7ERSBYe7o
0gXFAM95t0cg9Q0kN7bUeyALgj2erC7bBeMqgELosOju3phP7VAg0RfzRSnp
AlTnbxwSWPJFfAjcPXta9FVrcLjJ0uFhOXZe7QJyzvqKmEyTTRN5m2MbxArM
LjRsn/EXqgCvU2bcbeoxpzxAB+riC/Mj7Ja3t1XpN7UaJychlHibkWVc01nA
bmCwjrKUO4HsWf15+VmovM07t0I1A9qkQDDOC9Uul9Y+aBVYtW7+TE3f93fX
X9SHrUMMlNwTxNucqyFaJv3sfYfvS3Dx/FhCobLkDUFPAVNbzZBW4fGa96kI
VgBdI7TwVQHyetgE89zY69cMksi5GSwL91MVH6Qr6UnHeuv2XewcX80RDGZz
ToCQA8yiaslN/EjAk/SClUBAbJBd2oxAct3MKWCe1WLGSG/0W3NY0d6BNOIM
9iqrEfCxMxwRVGr5IOoN4Bp5iV0McGL2aJchXpo9nb1nByr/uCJQm+sqxin8
V8NuyBODGJiyYi/UX+Nfy/Tq0w3cTVMTjiQLs0alQQyXcSJGOVYUsORtUbO9
CNd7jx522k67/3I44Qf0w6XdvWQMfbdaQHqC+40N35vl58MCRV12Ac7/KIKQ
34052X8JvgSj94fl5e6+0yMISNKnCpJEfv2RWTGfM39nlzK/aaNGIM+Nj5hv
dc72Kmz9fC24+gpUP4L937aMwDHQDZznewRPN+hNH5l6hOzlVEVYl9fcTOD9
KKythArkCXU40WxSzmTSWRs8Mv/gSkYxlayujxtilR33lbzHBJzuPjald739
fwwhfQgMR8Gxt+2fnXqBWQ1vgFE4vM4Let2jXOBPF61XquaF5TU50eHVQngM
rjGTJzolPzjaXVUoWngQAncmxZZbYuhEbgq6AFVtTo4rlHprHX5ueTps23G8
tr9Tf7V+a3Xxq8X+cIkZndM9B5+CJV86swjV+xULVQNC+c8H2Eunfv8hpDsS
HQca6IRC5MNvPH8C6YMs3Agt4hbOoiup+65HQn9m0R4qOi1fRSk9n6M9SbPC
a3mIOStD3iaKIgqPy3cQ95Tx2nWbY1bvB85keMyrwyXY+7TmP25EFoE2mGho
O4nD6dW1ox3caajSmvR/OTFAsNiBIrqkSSoyAsf6+Kh3brqhu/Olccg2yum6
EQ6aW8EQh0T8AyMJonSM4iFJAdIZzTmZ/1ii/kbmees1LhTg1KvC6urbPm6g
LRaCriLIop1+lHMkwspZRYNG3IDOHR817aJzpjvgnZxMuNBq7xLPFW/2IJJH
xiOG/uUwDk6ZODp1g6tqJZtZnHaNbAGUuA92BeGJq1Dg+qZUS8zkkCrmKtDx
sDRV4l38xuEOWFfMu3aN7dfxYuckB1iTVWSRwBudOjC19aHcC2rKLZi1uiov
K0ZN6prIaoke/ONXltdmwukQkTOfvqXTu2Uc84uL0JrmXCQQ93LBsugx6hrO
6mMzl/E4d3dYY0uL+ot1P52zIJzosXfvGaocmJHzOs9hpM2VQINtOqlyYw3s
t073JwC1/JFhttyjhEiVn8xN1Z+BC7/Z1s3eAe/ShwYS//fqjN8MVaM8xOWs
XKZHXVUh33xt/rIr3axbH3kis9qQzZXy301i+Wl2uc7rlF4FCYtaJLgT4HbX
dSv/OBmNtA+NCOLdQ7EDse78JP3HP2ze5ybJ/cHCiWrTbYhFGzwp9OwK4/Zw
ttQyA5CWbPQ2yAtULKy7oDyUrw2wVQy4eXUXgWjPfEHId22uRMlzyeND6aqH
g7Fz9VXlrACQ8zbVeywjFoOSuYGhBgTCJnAc9HKzdJMkA/ntwSuwy9RUAsbv
k2SYFu3JdeP6W4QIUNxJFlOovCsIIYE9ZgPRL0OAdDq1I5/o2RM/K+YlJt9R
zl1s2poM0VvTr7w/vALw7dmjch+9Uhj+xIrkuJSoei+J8mWQZKUOytKZJcIE
3V91ttn3hPRibm8FMwN1WYBFGYdWxTGSLjwxL5JSXjZGA/Mx6H9aMiIuelVR
1tAvR1bC15CA70CSEH7EmgtjoA9Zfoxo60CyhkJWZ1XeGqTkNfddOg2/n1Z+
J8gJIeJcfQCDs0lKTdEymItXhJX+0Nd8B8JO0zADMHWsOkeg3zudsjZwFLMh
JlVuSrclZGBxfvtzrqSEP6/1dTrAumNyT9rPgF+KLyIZ3bdDCnYjxDaHdTR6
0JlsV/Vs8GbkfqJJ8Mx8Z6hfxvUk9ypuZQOT3F96/nVs9ZYy7CT/If/gdlJb
1JW7/P5iSF0F5XquDy9XxevrWncbQoZXIMskHpID+fZoHTYtu5mMGuSugSNk
salzwUnKW7z5GOfrRhCbtA4yVRzF4tekbH+2xmElkJ3bZHwr0poXaA1EFIi6
RxBmmZHIrr984Si2bZTwmpal9yIEDPGaJV/yl2auDI0Y3nIcRnE92wom7PId
L2mbfg7jMFlkGLUSC0TNqGWcQSjxn/2RT+zbz0C1TWVNF765bIQvP2BXjCFp
TwsxuhmGfH/+OgS0cRx6QU9bjgArFHDRpeH5o0iK6jRt9lR5N8nXUQ/QOf7e
o2l1W6zWPIPptlk7Dwz+kL2ZNAGG88EHZP68LD7VSkSOl+0aMU2Jk/w6A6Al
OsbPrC+1x3omeNnmkaijU7bnotWeOd2iNo+NEiSkSC5unCsxrvCy/7KmnxDp
36wg3Lsi177RqImmoXIi/yMEJ65XzGvy9ngC8LUQCiAsx1SY2MFuj7XOV4A6
LAqEGdo4RdbfsZ577gS3lfWuNy+ejVNdQQSw1BJSotjIRMW51UlAxOK0sPAr
trAZy7bddvrbZPxERQN6nPUqTmEcb3ruYWPP1A3HTKcSQ5T4B6EsxQ1um1I0
3CRLCqWRLFtPqH4kSe0WlEFYpeNBQWh1xCSIn1G9lWv99KY1Xjxd7nr25zLn
mruB0lw0AInZFnodQga/Gxmd39q/uDjkyFAHyypxqenRIrTvNfpP3dyngVE0
ejokp2s1GM3s535GhHLjL8t/dyVrbpV3hCg9Gbch8DTq0xbroJmJoedUCftg
IRPWl1CK5RebKnRHO6gJEnUkgmb1Yf1EF8K5m424MjPth3Iy1Q1rsYdulrBs
f/vpV42HCRYZS+Isms7EJQrswAW/JZAEf6xASJYwSAdMetoOmtc0qR2V7+uH
oDX+mFBUn6P09F6YKHPEOVCZ8MJ3GN3/9dlX2UyNZFAAhisHwxoAzQIL9ojE
M/E22dKGrnkO42SCYzkN1oMIK9QDVjci4sGsNm7xYYxfreokmIr9B5QiAKwa
oNgpvSiuCuVBKYeFyPzL/c1SVmWg7lC5TnvVwwU5se4pvM8QLW4nF1epr2Ec
rpQPDfOU7iMYFug1GCRm1BGM8HNLIvUm1vYD07py97ExWblBgOjNS/Mi7Eyp
3P03tzu1wehgO3ZrhoxipAfeF5ggN/PFZP20PgXbmLuQsDnZs2aAHOVFG74v
5CiD9X1wLHWHJTKajWiU7sut979fqZ4CjfcOdgAU3AD+ZY/CuMK+NrSAL1Fn
/fp+rX86pP0O8RHc61QcB7jgjgMa69xqGhP8iVOr1Fpn3WR4X5HLJit2akdp
Hy7k7AREjfmLiIOqLnqRG5EnVDZIbwJ4eaE14uV+fWxAUL9K3jdUpKBcy8b8
7EX72/EDFFSjp1dGjoyuy9CqEw/W+9OHfL47vYpMXfuLzRoozlaRW9EsXAR4
9JtZAIaehoQAm/OnUBYjQL07cqzpHCN+x55K43f2s2ix5oxpbJMo9HsUd6xk
bTmzE9Wdfa2B0w7AzX4/oefrVKrfUnxMzZN4ZJGO4sIqtl82jrAVxeD11tWU
qwcCjmh7031Ey8AClH9UW0dK54QhK4N+8cctUaFaytzL1yaTbofAw1A/LZXO
zNPaJFTVC0L+LLjZIrBDR91vtqVWDJ3HXykAT7tIGq4uM4gSzSoLe6KZYxn4
EnJ2ehk+RpmPJVpiAL7HepAKbNmXMwR2kXrIbbCToM2Pfd9191jfdwrQ7XFB
xHaHyv6ccYTSRW2lpYlxMYajed0kNMgueF/OVD2HVIgXDBDt0zLUf/YhvuLv
vgQ6BwsftOrZomCMroGQD6p/HKD6237FJLg1EI7k/Tice0m9ISLV8jqJ5xAd
PriWOLW7LI2K3JkqG+9m49tyhMlpyEewlHppTJIrcGJQOjYFipwtvnB1V7wl
Db/PTp3WA/GJbaCYiYAWJBuRo0+9ISHqt5USUH1aoGQMbDEz2XfCXQHp6tes
S4LajHM0FhnrgYlHyz3WAaJtsKAZ0H+rEI/NuyR/ms/wxJXV2mf1aCqtvOOK
EhkDeuw1a8sCj1gAePdeP5IRaTpDuT8ctBctY3LfbXSPR/ZZtpu7xGt3JL5B
vfBHedbyGdwGHRM2y68uzxMV0/1KfCD6nRXUEcTg7uQFlMQudSlrK0crd0Ma
ajixSo6jPUKAHpuhp8j2TskMAg1SQqz441Nk3kQy+0hRmHQKGGzNDta6leKs
h0UShI4kM8BZ9FmoFzB4A7PPor98pnRin7KyK5SOjpbkAe+Jo8Orw5NcOMbq
s31Qr7sEnFg1Bu96PhwsFh06hWUg3KMPWS8UvhMojU8o/zkFwdH+KrFcgDyU
RBSM8AV4XKdBPdC3lN/VatkOdGIXj/k91PXetkF7jQXTcEdCCdXXwyV+EsqU
g21kDJY3rR5q8qM07EJQGFNyP8qftTypYMIlWENvKY7yDaG3UnkFwFCWvrCt
QclqMdunvAwInAVf4DrmkOMP3hkdfAblDrQW7l3qvWobftnircuZ0LqG/lwc
hJeidhH34PYAW+DhXAkr9s8V7eA22So4lzST7CaubQK2X8m4CgiCPh3UaZv/
+W9boBOOxOV5TKKNX4rlJY0CdktDOnLgQ/uqtPGPcE/oufp4C+Mqkam7SiIr
uLA4BM/9HSAonqEUeQxUJ5u35pEDW4dcsCsu9citrTaq+GHsV4tH4Le0PQw6
7binQNMzesoVUcD1b5HHRKLLEXBRRRPpVqT6QI2fjMUw0iOp5Wml0JDpNo/S
QAhke5WHOR7SEww/JNvRNJMO8e0cLuH69nmEwO4yfFGb1kS1GwWUotyiN+35
fBgDuPAKd1D5LJS4b5eK5jb+/QIsyDPdg8lgTxUX2szVkcmoWvUebchIaVbf
FnyZLk54u4zGGHRGOVifTqL+dbn3KUl+hl+f5gomwUwqpjVngVwaH4HYX7yf
FsuZwSnmfTsqN3/cCKGmj4YzDp7BQfcFHm4JsQPnPWBLGjTPAP0JYqYJV6qN
ny7Kqn0aegMLJcggoz2Erj3MtFyjL4evyKT3Kfig0OKJVVivlwUXI/CWnM8a
ucDAvLpWJjKjxGCtHJr30vjsd1U75Vtz2Afdo17UC2UrVafy3DeYjnJdpaLY
UHTn9NOYlJvFUKOfYc5ZMcAW4V6hqPgeihkzzDFSfxOArCxdJfZziEqIhfVB
hiap7ExiLOZFbMjgAX6/e4wtfyA61lkvB6b6XLWJoCS4gOTlRFO1X8xoPS5g
GiISmDQbkgb9ueTyEmEd1BnrRMgvRRc0pvZ7xgozGpb0Av2aftsB446xeGZg
YGjrNee73/ZKv28mtBzWqszGaBeCD0oI3KGPK6S2D03kkZI31MdM6njtUPCg
436TrAVGUeRzniYrePpu+YlGX4PyIirfKVDmr9W4B4lPr1PRgEZ4HTcACXGZ
/MwnHgbGW+hx6ZYlA5pSeIUbeXXPDdpB7K3VEtW9aSvazgou2KfuLM3Btpem
AoGEQxBdGjVc7xRzKRK4bRcqdazGRURoYLcaMr/d4xcO+p/GDI4fr+ZKmbtN
CIHXCOvlA/L9Q1Vkw9XU/vg6A1DgZvJHGIBbswJhI2fvq7OdeAF9/Ex4iWzD
5ROU1kgVPfSeCgmB2i5mO8/IA1NsLm+YAlIkbaW9VRNlZpetSM3PXy90GcVe
BB8H3qJbE8JHNlVxN5OrK5IexW28Lksa0QpJqiI3SYlfZ3zRXiBEAI9lugKL
UC5c1rbGlhRMPSSfE3SvttVUr3zHm1CUCw25YiKoIeWSM8090OJ0KiybEQnI
xY95/09jdvT+3ru5pma/l9v3eHnV0gnBzwyn6YdQ3wQT3+J40HiaBf4TUHdU
du4P0EWYoWYaRs2tFZGIjHNEvpoGIgWr0YUN8D/vib974Tb/SA1EenzWHhTI
M/yRGsAv0psnlZA++IxV4P93l5AaUP1KyqgI/sZQtoV+ic2X/w2BM15WwYk+
qiATMgjsG3v3U8q8UtUHIBcxRuuMtzeE53hKjXOqL4TGcl3wEmsEY5QXuLRg
/LmGLoESSZnwtYkBtRMpudlXobKc7AZalBR7kA3oLFhgHiEo9EXYW0FJoymL
gqz8401EXmAzKjgukYqrw5d80//xREjjmXvcWB26WPNry/toEuqbLid7KBXN
Q2F7CF/QHc4OBtrO7Spns49OsALdmAVlrhTpCJ3o72kAfT76L1W2qWDKwc9M
DL55lE/eSnDrj2HPM/PhLZXTattbq7DvL3sC2CeU0m4FcS1pKQK+/iAcXjA1
M3POInPTkz46Uo8XfSB37ZwDkMa5zVn/HS9pLHuwuAW1Q5pAnZvta/rzFmW4
JKlQAqkD0uFhZcVvolA/bbGTice+LefozpCrVZHGgWcNnF9SJnrHSQj053ST
AqzYTrY0iNSVvD3E5BbLOG1rOpRptHProytHWurzcXICx+5ElFMFRtvUSSr1
DqBLm4byt2kumM/9Mn7e1Ew0hxv8AJHSyF30YQ2npn8+qu7mqahdBnkcg/V6
m/mc+IDPWhElJRKKmYzbLmjiIF3RkeKWqzT/c/P1myLBov/hF5VRvF92o1Ue
LOADIbpCicJ8a+28mR29K+3T9IB1ldjMsyVqhos=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KbwiNs+RESicQ2bzfXCvK/hI+b1ItVxDsrmCSNROzbcJzHfz2Sms1ItENuTGzrJJLGtBck5zUG/LCdUa+GJTGipDkM4FN8+6DsmAQWkZrEGTjdr0a3AN4EpBxWKas2q/cMheSUzYp6AETxScnZwa66CbwRnviXa4cZPPANps2H8FBwTL8MoUoG/cjRGtB+IVlFxpwT8e8qQuc62VoUtC1E/13JyWbAqf1g2L8muKg45M/NIrRrOsV/L+RaoBc1LKA+rpQ32gBF+RgWrOhAUZBGmtnK8skqqFoFeXzUsD05mMo6SIFN5hI19t0Divx6j9De3SDhsPvOwcb48Ud/uEDvBuqoGZg8kbnRo7dxgGgNNvp0njVegVT0MCW1KAr83sTSZmuQ90lDl4fCaBxkDPCmD7jV+AyB35fHIOO598RAH0Z4Mg3h8JonzXqjbCz1H12cVD6mVmaoDvkjDqrwWI3IpQLdcyWJRmJbmBW1AhXOS+Us63MuBHmPv0eJVNz5WpsWoone2kGcGrZm4FJUMSg/epVpQ6F33AwhJPg7HBLkeosAyekG9Cz4mwACvvhg/qA86lIpcfjyanyV2VeQV10OTPypW82inWZ8Y0ybyVh/jBt7C/4k7XgbQWxhB16iYaV5euzALhawpr7l1pc5LpyjdwCXUTWDePOYxYbk8RZ3m7k6rG6AoohidlOBgZzh7ORyzJ63YwmNFCMZ6k7DOPF3SHPImHRkIMICLr8amoORenziLHj1iHJAOQwUsg3RehAYqDwA6z3qVaesWkY069rL"
`endif