// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ejcfqR042641PAuo2MG08dCvi31xYMKDTNFvMu2OJucPnXb8qL8uRz2hLQd/
Y66cYzd22WQU55f29PyAe6l/7ejCqr+efvMWfWex+ngmytxIft/8Idi4RNV8
B1AJ5Fey4bfZK2OmFYWEX6r7N5RQjbpwMUk9wM+yiFryU7YQHdIr0Vch+WKp
NNMYcPFOux2BjHbDoptoa4rN7vngAlCa+yOBFCcnXdFkVgxcFbJMk/CuObYV
PQY9WaKhqxx+osyH1W5kZrE9Yyn2yLVuSu/K2GAqwqzEUbepeFz0QMtYc+UL
fhqTCa2cZwDJnUew9VOyUPtpyguxNHKtB/H8Z6/mKQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dZ2CtdY9GHgWXXZm/1n0dvEMdwR5hH8iXD7U0yFS6e5UHb8ubu0aZCQpDNB+
11yecUbi2ywfOd4UwbDSa236hy6upqqExZmqOB5Ko3tsS+kojnQclkOPd8yO
Gi78dV6p7a8E0ZsG6Yz8ZvMhh3EL9c250d+z/YrX7Y0KYo1lwmXxBgzqxAWd
1NKYqs/srVLkFCaf3dQd4k/779DVlOQR6TWohiLFeuMLHCXZ9Rb9wIBH7UIb
xoHEpyPqAwupFKkPD9E+YRgRAYnl+nwx6VBnZcLq+JTHO/8BEX7QpurRaBKN
XK/45uI0AGEtuR22dU5r9O55MT1w+oS2QTCrcHbrcA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VNLoMFSvEmLETLtWNrwhYGvs8XbozuVuG6nL6VvkXq4U4f1XVnDlNMEWzzuH
tnUQLKJ464Ve/FDGQKuvU1C2BpQ7b6+92MI2mxvZYBvZHRLok5SiBh7YvF5T
Dx7vMB+r3knd4RRmjOhvU3fC0s9zAsaA2EXBPCTjmtrbHolFmUNi9tDLEwrb
7tpcdSKnVREoQmh8xa3pzIPdTLYyC7HY3xQGYKVy7jPRgQ+eexs61SQlYEED
VXuVwFgE+wE6DoBKokKBnBwMRVzt2LXnPc+EcMi94NNzYt9y0q5KOdSx+3/s
jhN3hS0T6hJiPmcK7kvLE1zbVOr1s+sD81G5JY7LMg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MkrHjz70aEFQK0h0XScnR5CX4n7gzDsuIUlwgrupCMe35I79J6A4EFYNQ25h
jKoqDhWrR9VyPCbN7FosOdHPjTqTgoRLjOk7OaZpqM3M5fIikwE50B3UaFBI
JymaUDEp8AA9QI+0AbY5wF4F6+8//Yen3uoOM51Rd0mjSdQJjPBsjA8htUAC
REVn4eMOF0lLRor8kC+Bf1fCin+olfWKOUoHnRv8Q1qeIeRdCwJA7JsZ81xM
ksw6sJOMGdiIa/+1XzDjgmDZ2TmU7YcbhHW4ve+11bT4Cgfkb169hzMVfZjG
0rbRfxF4alCOc17KnGoCArlqNlXtMsU8sbbQGCy+Lw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kU8lw2mYLVmOClHRHYBrF8KuU3r7C3uLpyT9mAZxJaoyR/waC+5dFkpe5/Lc
XSjxYc2KLs3xbgHi3bV30Is10Tta9lCd7xgVPntk2ac//3ekn7quiPw7KX+s
AmHDUQTKoQA3Mb86+bKlz0zSZKx3/QbaVi+Lg5L3PTNcsv2x750=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
QiKvJkpRNNU46dD0cJs3tN/WiH39Tu+0cWNJRfQo7rszrTbM2Fj8D5FIp1ci
M5ITs1dJboIn1gqupSbn99ABlAEna7VfEge7pmh7NojIm3XynxWgs9MK+iOZ
3atnj3ln8XcH3MluCmWMZMeC6P1Sv+OtXhZNJS3M+QzbVWEqt/l4UoyjUBKN
jp5VrAmtgwMvVArabvKAK5PoDsRcEK0rLf3GU+giDSvsxC77yJTBpm3OFzkC
chQm4mLMqmcZE+M6bvZa7FE7dzCV9tCkLIilKuvukPIKiWlgBeLpLrk7lZto
Sp1tsP4PI7pD9FByBb7irfUeJoEGjnZAUzPP+QnXfTA8f6fonHxU5xaGapZI
pV558ZZDoYf8T9Y/C3bY0YuYwlFgJeDzYiTNcNlUXOcb/7sgbeJnX6P3Lvqi
h2Oj5dLAv2vN6ojISxqQjJXpQ4PuWmrDBaU61VTePBGmZ3tLVTAtQMKoCQ9M
7ZOocbCnYxuWI8c48t8n2S0EoCEKuMvu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kdG+7Rm6BWvWdM/QTTyLIHdAJtw0fR0ISZXyaDSWGJkQxIPwF1JvydB2gTmX
FBvxGswxjCxg1YroYTRY0xRruWEZzkxyYQGRDSUVk4lGdZ3Ao8BhVZ2Ghr1P
1OPnNtGhEmVbC0VTY6h0zalfJkP8vng6BcQFprvmE+QX6ivzjOk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EU3jYgcdmrt3fIvik5b6x5mJlItDQmtYmiVT4RcBrE8GNkI9KSvpULqIeiP0
nohgjg+5DthKdJ5UzNmtokFDyupaz8VmTck2pROTGUAKhj2vl3vMKAkJByBb
QGiQCIUODyWsqz2tyukF2/tQqetI7ioiAVhBgOh/am5Rt6/nxg4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7360)
`pragma protect data_block
gGtlnH4CpU2B1eYC92agBKD9DVWpin8ZljtkupvIOAjKb1IDv2l7rmDQ/hG9
WHqfMSVK4QFcAz8DjlsSUDDtA6zjTSFCRPwbGVSlJyEMUhIlKEvCjm2mHYSx
b5tZCziFh0yzw9DutizSG36TbbzxRXrFrIjeDOr3UKNbYHnl+FYGn5GVsHSj
k6VdemgfUfu/P4Je0+dDYDaaEafMrhd3ssp+rqJDdXa74uBtSj7Fuv6EO2Xu
Zk3ys59eZhHioDalaqKeI3ILqBb9Tc8OMaw3UMRLuPrbUyqoS+Ra/UE1f+3w
ULneNLdMRSnj5pYIXDlLOLB+Rp0DCYTokAI6mvG8mgT0LRbV6T8nnIflW3qc
sBUUorBpVCuvXISabAy1ydTy9KpXHnUtxFt+dIvZZGBydKGvGyRP/mgFinZW
NON5eiCLP9l5GffJzD/4fcmT0FYsqurCFgKzqkueW495H5ekl/uAr2Q0ToAG
lizzLGh9K4/+KELH+1OemTahXtCqdpZOCeUkiwBC6eIlx7wqcTVUogVkQqiL
y7QyfhsUQU5WyzEWPyMb1GxCVnWF8ZsVywWQKrJZ1qpQKxKMF/H6kwaci9nb
TVZmzYolwwaxHGvunSALiKSDoi7pz9BcU/g8TwU+vXIdwj/OEUzG50GGjvvW
m2Ifdw33quY3ei6HHlzfT7aydv2hVXhmakkxpQ4rAhxaCY/TgE9kGRxj9xyV
sWO3b896CFv+fkNurjv9Tf2/IXWrTzD7Oz9VkvHYlM6eLZhXQqWmufDFxpXi
g5Z2uCX1DXbvZD8NZsnwR2ovqvf9iXS1Qqyd/DIBlD2hpPCvwI+rHIj9CKR1
Brn/lOLwmUC9LnYFbbyJexWctz+oHQXILwm9NmlUlAiaUZajYazjOBeCIQTZ
mP0ftf9W5HQ1vyrbSrr20yjd9Mr0/QocP4CY/VKN53FPrlrRANeo5k4ueWlj
aAxMLT51E+PpdM8n+cd2911y7Ep8pY913Od8QjyZaGT+xoTf0b2nQ8OANX44
lqLRMqG+u2LWe0Va+AAg1rlSgllFQagfErwX6vxjsfvGulbGjokZAYnQi++3
n1cEfv3ZLs3lhh2Tezmz2ojpyDJyDJjp7IjPudw69EMxnn/cBKIgek2BeoN1
4nT662OuJ2tC8J/4aRpMGnpCvOJ5QQXDkZspHedoAxKUW+0o9YJJzpn5MRkr
s4wjm7NLl1nrjsT9xwJw85ojHYfx7Qi0f7QV+qNsPg1FRIDU/P9jovTxQRsZ
UaeJKjZ9Gjtt5N0vTr4UhB4f5IH01242qCqwlONJWci5ttkNwmlXd0gmi/KJ
Fpj6uijuslFkdU26SL+E8pCkZfLOJpSFGTsitH0JC4g+Zy72mq/576jC8Gff
jv/rtQUNNHQQrX6mg+ruux3GMY2hD3zvk5Z8gYBOMq8+8tMGD2On0VLOkV1f
mmlOfKV1rSkPTFpjM6MxPoo1Ic9hBGqYL2yYj6jNsi5+bYlsqVvp2xI777qJ
qQ9Mz/RTR8zpzzO4oE6ZxEewQH2/NJmCL+nlLTRSyWtjQiYfMMUCiC1xgAGx
EBgBX6U2CpMcBzQwoy9GelfDVhdzCLmIqkuQJN8Pnmz3FQw/1f38ACN6Add0
WBlNDYZIs9d/1QfjKNPrfhnGlTmayaMBPDIZOzOeFbJ8vtKnXJZRUsQfrHSv
X2TWQz05u7yZ92ldu6wRhl66IzypvKARqZn+GKVK7H1hAu3V8grQjhzMGfCc
4ZIb03kNgtYa+P6vA0OwxzZdPL4czbgf7nrMcpuEw+0HF9xEP0iNmKhgscfP
uX03unp998JJY3wr+smAtLZdrgbTKIBKkMC1wL1Fpa9geavHrx3oLC+kh8OK
6U9y8kDsaMScPV+IF4iMBy1T6BpUGh7lUByQa2tPh0i9+ihwdXFuNIisq/qm
QVXZRkI0UkaI2N2DqkkrruYD4d6v8d6PqIGVEAuesrTmGZOiAQ8rRPCw0Fxv
vttaDW2oS23ClBur7AZ+GhOphp8x0qVfQ20Z/kqs08i9YA2un5FhnSFIDuBt
jms4IGmxa1S2gamtSfru55D/rl7nSsvCQ7gp6N5Fg0eP/UYJTUYTjJFh7fvC
X5W6FVVJJz/zITXWBECeAvjgmWdF8fSMEmjAgavzF0JpD6NUrJYqOqibAkdr
XBAXPeHqpaUYhmRTDgvOaeALfd03RvlZoI4esgSuZXpOsldtcWIEbe0KC8ot
biOGehEz6GxLZ5uAUWh2rDQZ974lkP9Om7WZX4Osc8zUNWfuRIYH/PqzDcW9
IsjMd3OVH7JY0iZqNpDWvsigMlADkvqkf3o3SYd/Wr9drXSQFNUOBvllAQp4
P7X/PaIW3AUX7VnIRTkN/zGBz5FqkcweaSkM3Bn2oJYzKsYZp+Yhp1EY80/1
LvS0OiJO75LZacp8JpyL8TTyvNPy/A3SS956DDCInHkLWtZP+rYl6RIvDu+O
4lxi6/daNNK/GrKU9wMu5bsgVypa38B99NbDIyvI700ESbT0v3JNj1NsKfVk
I3idrEcts22hjcI2iqnd0g3S3sUUl0d3ah1cACJVBb03cAkEHe53tbAIcybZ
/LgWrbT4RpqXDJHsCCW3f1IYIJ5iQOZkuj15SExxq4igB3x8rphpSin1Cs7g
ACtkQ/vM1v1JedJnlk5yLIWa36PD65lBguoQuUx02gU2zydxVy1XXoM6gjk+
WoV694GbZq4F6SSBLpUeN/bTaJU4F6OFoYRDoTjESu6qgocDUxGRRUZRP7pv
wlHV19pWrkNcaGggTLKoLvBVuvR7iKniwZ63QNWXqfsrEUogIVXHpdY7XZSk
e0uQgrz6awq+1oTFCghhjqZAvsjWW62B66cubEFLTjArcsd/5bW1AxKeqaaw
7RviDP7lgbfDujU017qEf8ObnQSpOr+AVHkzlYkBdh+1O2+1CnbdAllwwcvq
zsmOY9SyaiUD7G0dM5e8ZInaXtGRVHwUH/0GqgUU2JJ63Xf1e4ji5x3VOLSW
OTxWE0qYnAcUqObd1gok/GhGbaEOmBQmsfTguMotHmx6vkFuryC3S94ojCHc
VDxec84eh1XkTAmtIvxlKVkC7pLGULiUBgP3pYn4Sy4n/rz5CZHzstYMkSvc
tZtGnV8UbKsFducyFRpREyt4vReEooV7gSvUneOX6H864TI7AgtUNqMWP8ms
bnXJ3R1Xry+r3YWJ7LxTYAqIIeEWf5ooN+aQxExdaAQztyKIHhc/vZOa3Egg
xq3I80KVKOlJ7dxkyUFk5XO5NWcHTbmjcLD2Z3f2sH3PZHqxa15c1zc/u/X+
6kQa6yabBJTIYYoqo0WCYAqD3ov349d58mhWSM+j2mBWwBx2OO7fNHLoEIhQ
+Gm+2P4pOQ66AU11tT/t4uSoj/pLS5cgDC97Lj2SCD9KNqjLn4c1/zNGauFR
TnmNnoEli1oivqKla14kLJk+AGStUIcxdTaQh6F9iyh1UHxuGrsm8UmbjaMr
vrNxOTAvErwcNNBMkKMK/g7gvd0VkPXhySyx412fGQIZhXd2v1sdmic81XJq
UAAcgexGoD6UlQYORKcvfoZtpYW4ky/md4kDfO6zI9TELG3/BUkBqbZyVAcC
Od4wnWUHnFO9i/oli2QanayCgz3vVAqQJFc2JtwAZlVL0cB2RupKhC2PQJe2
5U1npvdJtMqQN4RjasN3n94gjpADPoxOXg0HIApuW8bPpVTYPIRL6y/ej2bM
zMalpIFg3rV7ne7E2m2TJdfb7VTEheOaWRw5WZDo0bvwL6mDP1im58j73Kf8
xPKN6IkhTEaOFYcpbLUnoNqRuHQeg2Dmy7noMnjILHDsIegFQ7X6oDW0SIch
R2GjEral5DsFcNX5VQPZzWab/6MY7YgPrAWAt69+Z1uhvLxybggxwXrDDRGO
GEZhBt3pzueS/XhFSckZz9bvTI369VRMiF5rzZcu9lj/Yj8VC9LmaHFfY8ml
8NolJISWIEnQSfmN6qNMGknNEiyufiG1r/zUIoxwpxktan4YeyRkRoQtkF7H
gsWr6+7WXrcI+awCnn2f4Ih3Zbkc4vjAWM1x/s6OWLYaVRKFIeKe19djZXxE
LTVAv1E5SH4Il4SHlv7wh4bIo7h6PYW18L5zmmBdKFAzqjFALEdWInmhfzEX
svI4578geO/aW7Fb4++cMgEy/OZAe/ET+eMto8/2GuHgNHfhzPIi2P2vRzc8
6Mng5lHJvoIbrDGwFyAIleXGRskMR/5FLlBFu32HWnsMEGhehi2/xlfQOKc8
qx2rXwsju8FXGUm8+4L26g0DObB7IsndHaaInQbzr6RF1SzwGrW4Hg61wvC9
1zCxrahURTkqItUp7lmLvPdyUnrfGr1mk26RbDTDRJ85AAoPNrV9vmrDVnEb
YG+Yaw6iqvQyV39ynuaOnDlaYPSGKUlqab/v/SxLbfpLXqY3ypQtzalRiQhs
VaBKhx7fNJn9jJD5olnXIFnwueAeSz4jVMxac2WkMF8g59tybHmY2li0nGlJ
Ab1DVlm1MxURTZ5Nb88ZLvE0suGyALNjpy8f6TKMCUl17ppjSDRHzho1cdlf
kxiNRSK0HTI9uUfWFBX65GgndqtRKAlllyqdz+o6qCjIwWHuIXrU56Cuzqi0
xzzEYnjUvOSz9yFNIzoI/r5S+22/HGHEWmAStJ6PHTqESJOA3iijr8+TOHqw
11vI10f0nakQ/LIhULEIt5H1JkTKYTa904b5T47Z6igBtDlYsn98lg0vdc1c
rkydZuswXxwqxv41Q7MVvyHOai6Ndmp7GQLljwhLvDSAzADmrROIcUXgVf7R
8VVq6wzSJ7QVcoUScNW8sDaWb24Kw57z0YW29nKG8ZFexsElXbkYc/uwzZ+Z
1TNPqRxWEjeIiYjTYvhAEXORGKIMTS2W7lijyYYcvT239++OAS9r6oEjWGEA
02nj5ioJKq8HhWj2u/CFTDTkQ34mfC9beVnyAZOkbaeKNuY94zQ6C7vuJnMt
AfhrFJ54UOo2fKViBjwG5GIchsrXm9rUSC+39mTIYY2Sl2Bg9T5odNKTX323
GiAzAti2PpTaJh5JxYwQWCxkFwmz1FN3nMB/HhPdSOJb90VvakbnEFA1pbqi
CJAJPSr3Y5nzdLcZmfuSXdnYavYjg7tORRdoU3BCkXOvs+0hO8QNTWxE4aYZ
h2d4IjMWVmpv3ARNkgcdI5TJIduo69etwdjo0sWdWLUYqxAsXHdgFaNwyVCI
23xhMHSezrvCT0r6e6jzqs9q0x7ipxW+zE3Qkg3T1vrc6Wu6x6PwW1pLeoDV
izDcvyaWQ0t13DF1SvTy/QuU1NW+3+MAgcLt7wq/5g53/ZvjYZMRxdIiSuio
neBOtxR+sfhd5rYWkh4NNMhNdDk3onlXK8RrUNwLIr6UkegINBesMaoekA5G
Vw2biFvUlk67v6gTDtSJTqhKFvRFO+UPui6UhOtPBPFYBF2iAb41uljbaoYm
7gHdOWFWShz8hchdDc/iiIw3bXbrntIUk+6+IYfidrq4PbEgnHoW1qN+7DEO
d75jYRoLnU3JkMr5XgUjn99ttP9JU3TRZgJDguQF3mv1CwWcLeAT13jiRmgG
7x/z+FEEHTY4YPS566n6KkYLl22PADg4ZLCcd+lB0+Lxqt/njHhlFYEpZ/Id
S3G5RY6vOngL5nBEqlAx35VYyCU0OLa00ylbYcnGg85Ch9hy6LrlcaHCODRm
MYOqtPAO/CLgCBMVCUcT0dizQBr0qZ4pSFPDhb9T2klxHq77coVRrJ+NyQ2i
TT7qC5KEdqJsqlpnuEvh3KxMyiURedUMUXT9lAfANrJWnkfTt/9gYacl+ZLN
EanUBgPfyzL6lTnjzGXqp51pRHTkOOosrxwyEQZm9Jgw0ueW49E/5VnpT27b
YriqmWJ0zTAyzVNMbh9VYWBfghwZNbUJkKRRluaw4T9Ku5Tq2K7VKK4D6fOw
ZiCpxRssjjJz3reR/im+quFKViU+kRkYQMGa4uJ0qzHVonBpOdo19usLLIQJ
Kfdao1DRHq54Xf5VbqRyTe6DVCGrSZsNAg+TrlLnOoRuChY8Hz1P8i+eet1s
9mSskQFz8qnCn0xiE3h2sEIv5abxLBSnyddE7JcM71BDrbzM0F7YvycmM7GE
2fPVGbaU1BsCyabkrGFZhghObcqiqzT8cRsAYzqpJk7bRp0FBmvQ00WHlJRT
N2JzXOGJ96/XH9x6XJfoo6fnqGveMPywOPqc2R234Kn6qvRs2t33wUTkUixd
QC+YAjaET3tB6LWrXAN2r1qDawkX42HuYE7t8oez+gUO2UKvRIbuOHtWPC2f
YbNAQpTieiSQMLKmUuUA1AFOe1PAW+6cNXWUMBuJNTwBobU1SEZrGDq/o4Ic
hYRyJA1IZQjFIboPRELmmsafYpn1dn5lTG5Ug+TbpU+HwYAb+ggAvKUskMqA
m3z+YpAuIn56NXPF9qG42AA+h6UNxrwqUOVXEVhTFutf6Yx5Kgq6g2LRk8nP
f/6b5iyLwaPpYIBLKWC22vvWZL2ygbPbsagtV3mggbPeVcFKw20lGatunhNs
xtDvwu8ew6yLsUP5rSL7aLEqFOeBWAp2rLz8fd87P6nP12tjStYM79fck6tM
a8dfEGM6/869018X1PyaK2z+vbD+fswVqXA8RfsSj5sueZcvawnO/hByc91y
WTB10ZKXPhnxJsF+0jkZ7JhYRVw8yweIDReArNkmlI+ajeefYTdoSbSm2MGX
exHzR9p2J/tmaVzfwqIIiUxWwss6XwkmlJGggZ4+7iAyjkOnz24i/YH269X7
Vl8xBH4Uk27P4BDwtXRc0HvHtmEfrIBpFvoN+OJ+Xb6grktBX6PNUKqDTHpl
1DeK/usX2VQS6iCuewbrdFsn3FnpkxoJ3OV3znTnv9s0yfvM8KBbLdCzSEOL
8o1k00L1y6gO5UoazHRniizDmo+5UdWJCh55pgV9b2FFznmwYA3wciEklLcu
W3BO3rDka1Y3zYcAusfIULM6MHXiyD96XOtumCBpTbb1uuos2fLodr7jTM/3
Fth77RET4Kdj4K8YnQu6NwYkspSrKQH9uouEYDVSASUlRqKTfDtZMRzxAASd
wCuPTrIM9wEblsM2UMOVcFSQtCvWUk6q9U8cCxfD8OgKoZgmK62LnwV2xlrq
vd1IWMCmH7c5B7ce3TTLOQIo+u8zxvX207wU2jzaxB7KL1Wbp78g1BjUfcHQ
Nfifs/UZpG+TD87B3REkIQEnNOqjNjeaAe4JI4BM/gnF/4KDyw5r4nepmaJj
CGpAyi8OU70kqPrLqx3uO2p7OGHE+QqTY2tEkTX9xlWQ6zE1iyZQGVgNKqwT
Uc7lqBp90uZ46R+gT7z+LGsau4GjJWix8K+q4b0yS6gP2rJzwBYCH3LQiDFE
WRw3uLPyRHuDFfQOlPCz+Cn39GBCzL12h5+IdB+6/ytZr4kk0+WJhZRDXDFg
2NdGWnmKlcBikSX6uI/TX17VouCp/4CWcRIg6u34u9GHQ6hVJjO+eZQrIxhE
c/FuQBJTD+TBVlS+sh2xnXPiXCm2Fp7hOqZI+KjHwEqI9C90wyljeqi5HoDK
eEvwnzUnHf0YFcivD/6b8XHIbPDK8Cu4Di80Nus1boK97NDNnybqtxYWceEn
n3M7hWj2WzSbNRByN+EEL3f8A7MDxoPM0W6rC73GNIiWvVdnsWiqTpwn9D/b
Vy1O9hAFbm/bXZA5foyvsoumZ9hfjY1LB7kE1CP2OmUvbciYZlIti8K2fPBK
rCQNbahhVs467i3S1Z+lVAlk2DSLiWDDJjJhopeuO/seow1izygF+nhMcMtA
r18g267/DN3QqWOmCX7vYNOXeSf6q7/DbVNU7TLNWjcQh2/oHtbCj5oi3W2W
NfHOMKNk8Dp2JneJxgdIDjmHi5ZPQqjqe93UF5mMnj2npvf5NfHmF7/Upkyn
nEhh801ob3rfkeGVx+PnHho9so44nGJ+3PwaWmOS5/6etg5VewlwihpaUjIW
WYsP/oj+cXzYQA9McX13Caj9twEtxuVshCKSbOI837gSEBaL+Nr76KfeE6Iw
UQveSBWSNjIdXDjQJiZGT5vlJkupBna2Nge/BBL4qvuBru9m4Z4bGv/XAaYY
qd6JISXRrvujRPtgBXav9Ka7ddmrX+QLDYLYIpTv3vPhZI+r5fIDSdud9Z/6
4OyEBmrPx/VrkJwl607K3f5YKS7vgaTpTCLDZAeGFSLRz7WEWd+w9tS4UyyO
U+oqX+WSCdaZ/WR3r+fraugYy/kmdKpGyFo8ShVa76pE3vIKwgAcWiDzKgoX
2A7BxEiyOI5beCEU909bi8R+Rc721fZQUqMr1kxlW+GvIsoUGnazoKbzzXWT
KlqI1RQB+Hx0HNCGjgDfiXHAcXViBeZ/igbMZaEMNywLiBVpJb6oVR4QcUg0
FzTJXy5Tub9B2gtlQgrVksKNYMAi4VY+0Moy1ufRV+pMrYaRe59wNEyOi9/d
o/EILLuV9zZm91G6d5p+SCKFxfLUmOrtCW2lZ8MqAheNqHanb/8rE63nS/Wj
7ox4HplDXL+T+RyjIkZ4/8Wg3ntyWldFm3W87W57tEBH8dAEm0pSgWnCsRVp
j7/IjnkeuskQRtIizKOlUF+kt3jy8Uy+mJmlmrJlUQnZyMGhb7KksqZ4M7Wd
OcaKhvX5oUCVspBB/q5Y5f/Y2GNxgFUU+6d7rAHqTUxV0vT0NuVc10Li/fzR
s2rWW0nUnBYjOpQO0AiiGds9NfX+S/ipWYyctDKSWhugYACYtNyhAsZE4SdR
Njf8Uo+y8b/fhn/xPE9LwLCrywFB2Ml1ByuSW0WLgcVRY5Vk0rk7FMx2gT3n
P/jkagrLLSX03ekjzs80nChKSG3RfkUbt0vl5zeWoDIy+RsuqJOoUohh0jmq
7DBYkllDqhLZ/qiUL/AuiKPbDd0fVv2jxnkhMWdo/wS6gjxvAb4Z7mBKwgr8
X4ot0B0z2ZKlh5Rt9NOCeByvn4LG48gpc9k06IVBE0KnPB5RL/2W7FtHDE/x
fRRXqxW8I304yQDBgUJKHffjeHU7s3FCJTMKiqqf1a8iHRpw4nAgU+H0Zb2L
w4578AZyGaPaTbe7eo8LssJz/VE9Eb7VZhxt+UHbcIJzPiFCTGPshU24mdOJ
4jCN0lj2qNBmmkmivfEYGLKy3LDkcol9A2IpHzcuJH3zGgTaTan+8zBau4/r
CjWxoP2BLL5W+EB7r7oAH9tqAG0CUsCC8GNS/nn6XYghfMj2a5m5wxTN+w6n
N5IXE9zhfgzVvqiDQW6PXs0hCgw8FWaaRdodHeMNTpbUXN2PS/TeeX4z4iab
Ty5n0fEbcYvaO1gOyIhWIi1R4eRfy2Rmu6+ZcxImacoHekmLG+1s5V4kXRgb
Rb8VUPxcwFRJw+VxSZsXNaQqpr76CYwvLS6FRLsYEnOzN7j5THlrELUBK7+O
GfYu0FB7cgQ8UyaURgdYUaZvFLUGIFfuDIxbSQM+NlbFzXVF1hZURwTNZRCP
AoeXbxMrMCWjqlfnDZJ4jvXmSlb50Kys8CNM08gYW1e0NRV4DVG1PkrGK3P7
tk32Rq6siWbdu39i7w84wr9rDsYHeHwNOP2fCkvIhqfZ7b2qG8FjfD9j2u5E
9417zU6Mz6gZYD4QRcycSL8s5JEr5T3F8sKAxhVMHPV7TWWteNy+c1DP9IRN
uOsaooFfyisn313N8cGavrZWkl8/uVHm8D4Aa+k9ewkNBcNvk5GLeKBxlZaW
IZ3B+6IYHbRm3muuVWSWUDzvF4DlYNWMgFFgQKb3fNpMhjcRpmTzTzmmvpGa
UG+OeiheigoGbA8XSwv2SMTlRm/IrEi3Bw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1Ls+JDU1s5ArkODTcHjpEqztPkIbVN/Qes3lhqaE79khLlkF5I9oD4DhvFhT40bqWHM8oZeo28JYThN9lWQ1NSmBmfxMmOshPROviLKnzOynk1Tn1z3VVbbgUF+O2kPR/G6E9/wsP7ErTX4IpxGD8g0E+7EL6JudpTK/s2iURJuk0Yp468doWO/cVAK2t49yQR3ZDtQn757EK3KyWCOcYRskeGXTViHyAHQK0F/Rf+JK37yMXbjSnre+j1QR0i8abV/9BcJ3o21oCHLAoSngrk+IiY4pY9mIdQ7OE8O0DBXEFJrIke+5qCeeC0IC3E7ZiwOnQDRTBmCTtDLHZzNr10tHY7KBjqUEK/2xZCCQ66gtybCRuTZdimZQNYIiiGI0FVnN3bEfENJl/G3LSQF4tdHMqsxMOafOHjHgM8xPhNG9KYQJpstq/akKaI68xFYPWyRGTZHTsfgL+L8ghXb0iSA8v3k4ZYcg/LTFRUDkrSELX6gjtc/IkJ2pU7YNJV7nOjKGqWYuQ6gSNzmeyg1iUyZ3r/CCtZs1Z6e/UzFzwHKG5chJ1tq40KDPeL6/XUTCS87Ce74oaxjdkRIFdgYK9GpbpJDteLRIBZjHaHJqWjCqX0L86N4GA2epYTwhhJYWr7zbTE23Fqlok2ndiSuXN9kx4y3WLttWZqLfb9suLfRKttpBCcXfTA7RrWp/Fhmw0NhAWH3HkiTBnvXKFqmRsySsSM8/X8lo49b9gWoUOu6FI6H1+Juqe7r9o/U2lMj8DbMnV0UDSGedVnlVBr8vuri"
`endif