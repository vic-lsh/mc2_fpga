// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p7sHKiunB+AlpMt1Elxji228vFZ00q53QTJpVPVtD6fbB3Q0ceFnnzhitBxT
w4xGnGvyW+3XfBlodo+n8+hA2sEx7v1FNQVwVBlj5zyt/9nGhgGQAK6zHLrk
2xbCe4+dvjsLFeSG/gpOyft9Ft96QNzkgwi7lHdxZUxj64/3HQmvzF2DQurT
QT8F3S9FqrYPweVycukBOxBuXm1lQbdP0puZ1DEncsvdxPp1eT671+4pKXDv
tE205LjAQyC4xwgDSmFMeT0aKx0HwyfgL8a1uutnGHhBvVLyiD4LbOJUa9KT
NgTvyxLh0i4JUTPu6yFfxMrnsiiCLu9Cji8t9cYrew==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
amo0mg+u1ZkFP39IWuZfq4c/VcUnwq6XHNlAh4llen1pg7rZI20OnQvIpdK6
TyvvPDW9nJS+zMYAYtYV0LZb74fB00GCv9yJUfi7K+q8DAppeEDuZzEII4K3
hP42T2y51VKPWEWsZD2uRClFJcxwM7gHrxV+JOcLg74wkAxqYkTmDOppI8YL
bJoJQndmCKk5psdzJ2rAswJtVxRMsgHsZlpqCuEgP8Ilh8MYyAOI6YNUuiP0
m722Coj/xuas0tJk8fZPDmGPdI7oCQ+1xTMXBxrhL3BQI9j7WfxIzBV/zxmH
S3jDvwS0j7swoxrQIeaHTxE+uPUGlD90UJcc6sCWHg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rNLsgxFRvua84ir43m549CpLQJquj0MlQp3NRdeJb4+zUi2ni9qZE9FMsJEs
isOaEh4W6OW/PrzMeQCLX/yf1tsyeE0pMb8Rcez+HN0JzaUwHdZotq0UJf4e
H/0fPDqhj1d39sj68l+vqnF7m/3B6m7/JbmIm3ADJfR4Fr3hXn9ZZqmCFXHN
XrxyCg+OXO2rWsW20RDuk6Fml3mpXd0XbaiqWko2PNTVIGe6EZrIDBqcyjSH
+x89p26R2A2NnoZ7CZVC6Zbdr9jDuzKDBpEFBXHJRnZuNyVXMZRiGEE06zA/
sjAIBUk8iLaZchTF/w2XWPQ3z6MOybi/Yd3rydxNCg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WXZEaqNbyafoapoCzvcGHihntRIVPFd1fgPvQP7qI53lTyUYDVUtFSug03zK
gfPMFa+bTMwxr9hJYlqmKlAKlB+OHcsKAJGkkWfqbbJrxuOXA6dl8fl6m0t2
sdDlGNfMIAhF8gONrF3yEIF+E0KbqqK09afMmGENLcBYp3wSIoYobyrR/Z35
tMa2mJV/9kUs1rRwvz4puVQb3GLff/IAhYBSfdk1xO3n6eGrqWb9c2nj6RgQ
80HezqMPk4Vey5+clyvCtaCwz5W/lJ0UZdMOAfUpoQtFonqmKlyK6b2Rwrmt
mwQMu7ufEbOalN2YOdZZIYLkv+8xb6RaFGdQw0GujQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nKcRuyXp9oW/ssWO/4RXsI7azbe9HUBSse1u5GrFlah07UjH5VjBqV7Ww5Jp
kBYAo5N+VMBKb6Y9k6B0L18DulgnXpJI8z1NTIRM0wgw6UqCgwaVcVCgfljz
gaycn6HYtuxT5UtJtSsqV1wSb5+VMBvk5j2QOXh1zzO1Dt0PApg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HovCFpvNM7FvpB92JaFiIACXfVkmWdq97oANfzhg5d6oG4LUAbhvTmodmG03
6V9BSwH6CWlEi3II7AD5j00UKIJZnqtRHwFmvd/0zGyMcK+s9SGNdvYWKI9A
B5AQH8JUG6xfXF45T5Wp7odP4+4ZyY70dS8ttcVTgEM9jVy6+IrZ7W/pU6D6
IvAUvfzad9Haszr/qjSDGFW/kqJa/C4ryg06ZqgriXijIb4TO9L1vgvEjOea
Z8o0fqI0Cu7t1N6IV02ABLR0EAu98q1FkuQy8z4wtIblZTAdUV1eMiBM25Y/
cARU2n+ktWUozwTRc24TPEqWozPSqVilx4niz/etU4BnRmEhk8InFn5hLPak
It5irtdHH8kQFkN0GyQfWfgFLcxqkyvqj0a8mUWRITS8ZqyDkgqr5Y6FWZ8J
J73ye8o7xc9F82B65s3ouR0PalidvYCu3e6fpDTwRcQPcQxaQa26qUtrhkkK
2jasBDnaQ++onTuIsNFgraD3gYV3jYzV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LqC2KWTLPDBHtvNZkGMFlcG7F6C95dUR2OGYpSRJU8b7GYXh3iUs+6Ln4ELK
7OGPAAw6ec9UddV8HGXwDl5TZ96DWSK59/bTbiFi5ICiXXzc0gFgmgVc974m
dDUDDE2jQ1YSr1jIevIQ2BKPfrFC3wi/NZP90qvZpwA9pfcjqzE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WGgnvgvIhn27lSaFC/oWy4F3NmNoAYDJokXsibxX0w41UUUhTK+wKeH23viw
dxqJPUgFDvHTreFTztgZ4OSnJhVb9UgedfjCccTVN+nAn0BkEUWVU9eV7s2M
ZfwzcyVRXgBQbTZ/9RzyorLHHzUIc5b1EdlURJBs4ku9Tr5JMpc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 36736)
`pragma protect data_block
TTf67jhmR/5pfEGJEmVukPmcIHtyo9Cone7gWBmE5JBKcPvfkfkzTWIghdXV
scXqAlLX3pSLDcpw1Rblwhc6Jq8ZlEi/9OxSmiuOpvBHwFa8DZQ6DXhj2+PZ
qd3CaLH2A02q19Aakv8G025R1uLT0Ge9LYMRapxZhxrPkpD5fAd6rgo5ouCO
XNo45inE7zR4Qb0TKbg6hNoTifnX7/n0El2bYXTBq1xUzQYTkf5kYdUohduT
8gnb7twvVYIWiwzLmMMZb5AFxPMhu3uwk6JpPOt7X4ANGqh4DqjvHS46q+2m
q8SV8Ce1gqvEuWWK5s+ijcw5dNslkt6iqaffAStH7Mi5sAlKoAcfrMFRnfxD
hrT68tPqdan2xcNy+kz5d6qiXLjg/R8VD5pRvsrlpfUjmjxibmPx29XTv/YI
I13Rc8mZItY08kibjRCnREvKt6BhA4EovOMLVeFqGwTiEVqeI2ncThqM+J67
shhnmMzeETLzuyShtzPfI/kExeUnubyMz/5K2Gog5dvLQoPnstWaUEfvXM28
82er+21KetnGSWzuDGz8HspgGE1kcyJBR3Dri23l65vsvx4YAejI2D5ZZoiX
sls6GeNuG5b3yadrWjLhXzHA597UDLLq6ZG4E8vL0m0zq0/wAK4zBxe5atpb
gAly2ahncJuhE8Ns/04G/YYhw2FNCSAjdzEXIWzzw88ba4iwUO8MQodigsq0
ypE30DnK/L0mte8600m3/8ykNB1HsGWS6xH9GkW06nMWsFVk4DRXywh3JysX
Yl9aQiQ2t/CDhGn35hwB+wtYsxNN8sqmroFK/CO9yameLhK1Z6gYNwLjxfnx
ec02JBN9BKkTwUZ713NMQTVBTN+1zFoE/4QEPyfL8+DckLkElAdTjR0VYLja
7Nq/iQbZ2Lc7Yldkyh6j3yr+4qqNqaouNovCoMLVYhpUG4ZfkLIOEbVhfKTl
EwIIJ81amhUSyIHZdCtjUyzfzNhBUBZ2F6Y2R1Klek39SLXET6MeNMquy4sa
4hq6RVKX6dtuCU3ScWX7QLtq0iKsWfUh4H3zsbRWFmUAXKBv9AvtjuqAUVxs
QhhmBCzIfz+nkyQXluPlUh7ZZg8wkli48qKL8NqW1hzrj8+cAt5B+DxQRPhT
anIh8hjB8PWp0CD2uOSWRR2sUy9b7qJEl8rdYq++kYzMVQOI1ZwamoiraDlS
fL6KmxFMh+Rlx+xmxMiumKhRy/tPH67PAXstLIZ/53kRin/bOmsv5eT4Kvet
e9vQ3H92E+YYxCPqo1nCYgHE7HVLO8rCA4Wvkf/43HYrE5im+yeUw/Mlk8cA
f4OW3Q0XWcfavqzpdpponyZH6JAY5EFY6fyb6GqghHjEA9z0qJrH9XK6UGNO
GzbIn/iyQoQeevFVn5/VWuCsUWQt6GbXVUXFfzJlHrbruLy5aWdrQ5ujT3h4
lDIf6vZxxfvXWoJeU+Dfj7mNkDetXXEcvEngANeLULfrj+xlKvUBJRHiOGUI
641AmkhncPIFxSttgVzCCDrI4ixROg0e7zJ7L5beJkX+IXNnbFkvSYcSyiMm
sTPNbACEcTqGwnl7UZU25gMzWfa0dgrTi64GY1JBRMCuyLjzyuPr9pljvH8w
fxqMWxoqOdcNk966fDfxkVP1bFcFVnEe0HllUp+QM1qVy1d9g+ofgHjfJCAz
B9Igy4TzCA3N6PrEbdT8WW0qCMlor/Fy0IFQNwAEkjkCnn2cqcSq86HSM9QQ
GZ0Im6+DCnImM/RgLQbqbYR39ZkaSJxeIXyiycG8NtnB2Rf3mAlQ60AHmR6F
8yyotjHG041fTM+u0WSRB9OZqGPvq8C4l0H2DsncXvmPWKfKZw2H5nG7npVs
K9vyE31D4b+RdYYrFwLUuyCLDay4lzsva14OoNpXKIxieX9Rks63ksqFGp3c
nTRxe+cR61OES0ukLni2uoBcHlClYlkLAffFYAc+/LQODUeKzDoVLbzhnKZ7
8WBqqF9v/Eb/I1IONB3lzxWUqsCjLRje4wvCWJT2A7JSBFioQWTN418uvv8B
+VpgFEQ7VZlfq3rCvr+HatXKUheb/BdifHJGYzaRKk3JofEYN7A8njAJeylV
UPjKd3lbtOed9mXqF8KwxWeKb+jVPTkqIF22VoLHeoFyriJJiZkBB9dCGt3o
rN+SOLkJo8Xzi6E8mnymnW2HWoG9FyqtOKizx9eu/RJHBz9O5t5Uve2truWz
cR1HJ9vwXx5YWrsDvduKX+c2BIs5+z5MK1p1dtN1qHmaHCN5T3v7byltFoA0
N6d8719rayA5fpWaWrI4+Jmcu8QWcGuw0cicAi9+oEYnCLdrakb6csb4Zw7T
u72nMzRoJ0hNJHrPkBu63m719E251BX/TxfUTwy/AjwOcbYeKtPaW5AcPGQ/
uJR/iJPoLKS0Z8O+PqCSmTznOvAqYKWxlXoFGkbH1tZhb6kVHTntm6V73Bgk
vraiiHSJY0+ncjSSe2JGj1AkEOwC35HC6mhsgaH2OuTgNyP9Im7ne5lFJ1aD
ZPWuaiC0mzLwzGYsevs+VqHIks3vp/0I4BP+ImKJafkVcMhBnj135yy1qIJR
rLZ/WLNABsqGWFI0i4EWdyIob8VYcLtSigJIgOZYvIWRdtEPKMr2S8r9H/f4
EeLiLBjpmGr01OQ3Swurnl20E9qkaKSuhh653CbfShqnrycfASIJYvJlcIg8
xSlqE/CR6xfgkelPUYGW3BrK3hVRGJGcydNM+lF0uvpeqcsj66Y5WLxR12Xm
G5UgcbOrynn2sEjVvcODpJXdfYDxZkyh0DQ39mVpPiLUjTaJvVowbuKyaGw3
RKD59Hld1883u693SqHYFmMZR3R+r70C2JLHBbjhXSxxTf4gN3jeUyrNUIeN
aO3nrfaT8oBYr3H78LmD7aLU35XcFdpj3wW4WyGL//zIwILkuJZz20vbGQDZ
wX6f+0LRjr5MbruDyXL7ynU6D4FeyE+jAgwufsFhcPiWzXNjF2+XdDCc0hM9
2moywU5/vI3wgno+5bsWGgpyZ4elBmDrV0mn/AaeDLkAUWdB+KAEYhg2fhbQ
HU4ANbdk94zMfjSs3BXxeuO+qLp9OxMOTM/oGzVwOkwX9fYdHTViX80V1saq
ToZiicGsrne4aYhqYy74X9EVVXfU0L66Ys1A0OecLlgq345QpWXeRwLgldNj
5ANhGUOmu6p7llQ9ncEfrUHXZlPrLXPvTKn1pj7NnYDWy2Ecd2MAkPpZhfGl
y0n6sBUjd4b3nbKTJlHgcBlyQkEzLmA2o7dY1eE+3MG5TrdhiZSUbu0HbykZ
wLaXm7yOwK5ZN+4b6o+QJrseq+hFGPFVyuu6jdsdJiveDS5TBXN+SugvUKnR
ODusFr1PznPOVFoOEB20bP5K3i7LimnsecU2/FiCJHerrcZTjU0iwpu8wHiI
4v6IRzzpso4gfYDfnlZWY95Mjhb3RpqjX5GmOVkLGbXvwok9LnMNyEi/+Nph
n5x1TCayjEkHqfTsflwweE2SyVQtyIrKvFevWaoacLWCrt1zZCrdsPd14xOv
zJObCj/2ANVmOJ/zBO1YzmjQmlo21pTPWd7VUzdV7GtnrlG0yqBYlj6rPAHA
ZAhCtnPfSnlignr60CyGdhvlJwxEhtGOI+WL0fYswt4pymsfWn1XWg1nRvjd
/U5FqwwwDjJs8bycft17IzzRMi6L+72rZuuBY671n84w+l9OEgoDfNogr/nw
bOnW0M1qHd10XeaM2kdNIY0sqcIyqz1cI58vT5p3TgcX/F2A25P9yPmLJS9T
S1l6GgnVjJAFzqFaNMN5pdI4AA1QOfnfY307zI7CnAJRYaW546xZSb40p4eL
09bG39jYnLbtODZEsyNiUZ/LtzikSCOkeWnteU6A0k8KXwm+8SfA7QJ/8v3I
LqrvaO+jSJQ9qk6pVnrJ/dcCginXYhxtGwCLV/w6H/2BA07DwtFOZWDwG6tB
wUZnMWxJR0o3lshT6400aJXw0WiwvlKv1BjKJ4BOGIiBGYXZbbdFvCHur2gw
qRwsKFXQtcM3NGGFlTLgK5DyqfEiiHYYrxZtNAawmoqIiVi/UKwqdR60+cgN
0k+DmKt5I4WNRHYHT9w+A5giMtw1MowcSXQboFU58fvwTWOSj1U3RqMkyihw
miNLVs2pwKHMNbKtNUNkLHOjH15FlNkxoHj3NOO1OVRs38Mn4Co+FIEgyffu
RiTpE4jmkPH2XAEfKgNtdMCGUAuMNmxYfbLD28SdDH/AC6Y3fE4qnqVhtzEB
x/bjn0+MwsI3n0NjyTQfZWW787OYKhxeoRtGsU5v2RSm5P2nwXHpAAobHNrX
f3wiFJXFBxfbqQpqtQyn+IdmhwwAwJaonqowzgiQZ4y0hQgNiQzZICaSESkF
2V/M4s5NUMLAfD49PabhGnuO/N11axfty3CddjG/9T3V9Tbaksn28Q+AdkYC
D2mHZuaWKiyFc26ftdd/eE2QwLWHzDKqzNPf8i/8RAS/JM60gX1inpIp61DS
CEMJDPwD6cx0qwvnHHx+4jsGqbresCy9UTj1ZKP6HQzmbk9gQQND5Be/m1Oz
YDY1HLBhT5wrzyx4IB6xorz4UMBUc7/Z10zo7ZSePKSiywr2Ay3N2AmCPQUJ
U2rkJ5hQiPQGq26DNBOasgs1TiUzoC4ZAwaY/+68Bqp6EZxOYSaiW8XiRI5h
WWm1xYKCCeRqEsIKlTwlytVXA6hAD/4IEv43UtkMLgbvmTQoJBPJO0AT+C9/
3pEXQ5C0t4iVHtah6XskDt0fX1ePQozOP3lE2BeCPezhxtkDltwUmk9zQwlD
JMM9M06Qb8o2grVYi62IYxRDtgIpXqKG68hQdTzdu0B8xLQ7uQ88CKYkH/Q3
V5DBb41zKAv3PI2j6oAQNzbPkO4HZL6tzsZPMlh4dkMVZZUYjNVJcFSd5ZlD
2+7RHOw2fEc8MBRxb19EvtTgeI5x3uWGJQYdUPv4rI3qHUDqMklAjuPtga9L
offEzZ7leCnnOi+6hi5mWI44MnU4535O+ZGsr6qlexadojAz7S5Sj1NiIsxO
8nK7tx2FWELfIR0jiZitmDIC3SK6Wxpjo3R8Xt/32PASBIq6bHW4Tv3vDJ23
tultWFr6LD/QeTO4p0PrQ8Brh1T7wQWsz/Vrr1+V0cvZYU6dIkxRnJCymFoo
+MNioS3fJGzOci+sKvAppPk6OqetDnA3m+UbPLTaAgsCOo5fzgRLrmgNGISi
MIoyQDtnr67jQMowg7KZtkm1h9FMZ2p5ol+Hi7TXUXNEuhQnv+Wh7WLQwcBp
z18jadFJf4DdPngilgCBSjRAr49+XEuU+aQ3UrMD2VMaXp5fs2UbRYzKzbed
QY/miQ5Qf+27zjYniEEbkh8XIs8bHSK9XfXRaK9nxYOWyoa+vpJaXxoibrlT
999NEQHN4s+1vdi2mHgvbfjoOHU4470NgRDa5lGBpXV0AMZTnRGuD5vlGetQ
UAOKgT8GyUDbRJNQEs38Kh1QhbKBjkAuTe9ivujOtfd5pHPvENmmUwtmpt5v
Pkydd6iQ+jz622jdF5NUzy7L94rFNCT7q8VnD9VCSd3QKgQs5G6xPC0J6YyM
9A5bYXb0dRUc3F/MNJRyT2svU6+0LQPetjFdoiVrN/gA8IjSGo+XxGZkX9Nl
abjslqsdjXA6RfX5K3xuXlLpSv4EM/KbO8jp3OQtwuKQpJv0YFGqZNfOrxiI
GtFvwhp4XfLZbRZpq6EodN+benAEjfkMX6m2oI3T0mjUjU7Sc86DZ/FyfY9n
NxGvboeL/6fVyHkYRPy8HDKjsiAF3GGsXk12Qm3mAsA6VmaKxucpciwcAPur
AlnCGcC5tC5RS+Jkn3cY3AyQ9xJXO0CuHtqIF7WV8oNJDNH+CFuTJgD+FN9v
vi1V/P8U65ZndCFrctE6n23rg8Sw7r8dP/RyQxgERJHgryHH0v1cKDJInlwd
YJvpuHxdZeJRTZu+3IuaFF94ZspC3mwBYek2wrhy/fAnRt0AxtGfycfYdYvG
WYHzO0OH1gyQOZmfoAnnamX4eDu6jIk2BSrJthRshYBrQxP0lCwaX21rJwz/
I6C+eTAVpDbLlvwC4/ddWaBAWT9Fv3VV9hre1GQ+U77PVeqIkm4nFYxvooi2
kkSOATBOld5386E72g/FdE3vVM9t5bn9s2c5V9C5RpI5jErBgrcaKJPAJbnl
TK6RdOr4aa1eCtjEu8zS3gpuha/AarvXMt510pjY1ushjTBJgT6ytrDeyz74
m64xapO33LcUJh5Z5FGj+fF/ngcTVZ5fjo0Sn/sJzfSDFxVBqgSEU3GPm/Mx
uTuqYy/ZAweJy9mMzwIYpryacnrOZClz32Z1cuxwdN855ssTgwypvLvlSybU
aAh8e2XPXM4n7Mc2knoXqPChgifyRVFtneaRpDztzyvtjZkFtPP/kLHzGyaP
b3c/ZfpMYPZ/LS7qKVba2gZpJl3xpfFqec+nIS81TbSFP7qAvRRI5wN1xFxj
ZnkgEEa8YUy8Zpq502e7oUIPWG+68lLru8QUS+NsQ//kgAkozXgEVnMvXuxx
qrfuMlbXWu9ydCv0ptJIyIhNh9y1bzyzBEj7y4yD1fh9I9S2nb+tKnfc/4s+
mhdtq1d5N5S3OPwdUejESZbw6H4MCwbRR3bz681qXI9ZM6PgZvJJyiopcfOr
LFbDtnVIQwrTmlv6IQ/0/Wz1pMzd5oEiIOAP+W858h7PRYF/Q58Sj3mNfb3+
zvJnmVirSmMfXkKnM2RlLzk3vurDpiR5sYp7B9EMxQp6blR/E6Cxjylj/Klc
bBZwoO7ZOT+q6hUZFxm2ctO3a0O+m3PKpGYj77QHuwxPFyjkLuELdIGjGSg3
ZYbEOTi9rc2ftd9qst2IHihcnPFTMRHLnkKHJh7v10tb6O0u8nRgSwGYn+l3
F72EBd1IGB73FOhAFQvGPLpEF/pC/dcvtdYp/TzKC4iHY92MPyHg2EtgenSt
wKwM11T/ZIo7Be8/AJxCTrr6tikMTI90uhZB18WPTBQ4k3EJTRhro8xapJbc
8WRV65zDblxBzECEyy2naZhQmIFZ5pXAr6H4kxysvJyrHU/IyO+r9SO9Z+qh
G+WTLQ6c5eX6u2XcOu46v/JoPxqpJSIFwhmUzf5rWTfPSHHpLNg6QQwM0/1P
aUyrn9XbRj49htH0Y0jMgxPX8R5VVHapgR9fMZWR6FjpzvZ3AssaUpHrovj/
Ur3jHPc0X9z7ijvvbc6avHOSusFMxPbFg5DhLvqlhbd4st1UcueX13gWYVSX
USGewhY8u+tyKu3wPB7VsKwSif8SvLQ199Jt9aEIOvE8q2nPcKFa94VIyDDp
UcMV/VnwabMQdXWPh96gkZ912opnSCSwb2/FA1AQJM3c8bgixU4EQaHww1gP
BLhOdN2CdGu0sFvspbRj9exNjT+l7LFaWd9+4Fo8rT2aOyEJIsl/ZfgQSyKP
P9ZfECfFdZAJJAMCZvTtgLcOyEYpnNoo/FwrRp/6aeZKINJmDycCQTm/u5m7
tGhbSfElKf0gZ9VKi1QTsloZR22CIZsYs/8XaVnX6NIVx+A8uCfKgZ1hWVX1
unpHNSIy1zih4Tufvq2YYJSVL6rJZvUrvoFcK6oZrK6yheEmoRS+1xtWz/i3
AugDzAeuTAeWFODVhrrey5r1neggGxk6kM6HB3XV/3RDBbiu+TjsnP6ulMp7
xV5O4KtZESownhHgbe48HMM76UZxX2PNYVWT2+9Tv/2cYT2XX7vr/kVG5kQD
Ns6Qh+7BeSXtntCszv6UgdRvcLQ6jrwOJ8N9pbDZ87fjlxaOSMs8CtofhpKv
YUoTXmyf3CEHRIf+Aqs4wJ+ISkqp8uKFBwiwHkSJjwU+JwQqnavLop251V0J
KjCcFP8MXbqKpw2evidG7TJdchRbivniue/jo5wtfr2y6NMGgurWHcr4CYFd
xPiVIkatVzzmvghkUYtvAEyOMI4FVE40NcqivC77UHcdFpGZeiiHAPkRW+Sn
MoGAbXBzcLjFfMNeTCUOZhEL1o399PNJ2G8cfFmQ72diVeO2lP/y0Xes3Fs+
OagZNq2OkEqQSclvOuLMOMWOWFAYsLdPEtafO7YVU5Ruewnp8SVJ7IntwB9j
iAdAjMJ+5NINe9xTUh6OmmcFekE2HS8ALyjmsqzueXfoIQ9PUYzhL6/ojwXr
i7kWHpu64GgnE/JEfAVQpXLnCFxLUnGmog7AetqcGmxGUB8ZJvgEer0Dhcnb
2qz1d4YkS3Rbf+NcTt2zGMX7DhuICsb4zmWdx7gxI4z/rMAA+OQEWqqTtY9X
+eX+1hfJHkAO3orz/flr7yvpQS6NOccmuZ2RByi7nr5wlZCBNp9ArKAQhPfK
8IUnSsX97139uJ0a/we5RCu75i5HwQ/L4PIwR9+2XEeiDGDvh4+M03YGSmRn
oi7ptZhzMn3+5AbJyLrTK/nfTpPFUvnW0zOJliXB5Vp2Sl8UZAo0HkxnbOv+
DxsemOX7j+sikrJe636G7gpjreEQ5YIG74es+b0j0LMWDZbXiPi+cCpKq2fh
tCN3al5O6sJXp3zQnbVxjymfYFZmOGCUL+8AcUPb463PeLmrBAHaw3eTjFpc
NsrUnYx0K03R6ELwlqz0KD0Ny/psTQcH8ckoD7/EE7tGQak3owPmqJcvdqJy
pmQdyAqvOTBSaDw4BJdKU+VEgrSL3RlHoeCdUtgmT4b17a+o8I1a38qpx++k
mQ024qPPF7EOU5hgfslDgCy/8RXY6qdhA0Garb/C379D3SeE8D4X5t8IrqLE
S6e5NBg/1kEPPsMzqvJFvV9DN2L18gkcvBwOS/OUOU8pMwxvhVSuv39wO9Iz
GVK5ae5K0oAjpgrYthEaWZLeP8gWgBavspbNFuZVSxNvCk7cb/gyHRn5ANMf
B6rsGT07qEfdIa2re2Jk5+8TUzHKcYtnet5KJUExNUfP1YImW9ntcIiV7l12
g1xM36rxL5xr+kvRzSlecu6L1lZzhPVmB0uYv10vWvQx2IXhrFlAEURIzSPJ
M5zIhVTPUc8dQ4rkMRkN1RYuPdqyCNDQypMO1yvNX/2g2+YEJUAXitjLVEsI
w0XELt9NhIWKpU3xpHd/CvULY4pPZW7J7lBwiWw/Z5hcxs/EvpL5I4H9jIBf
BnlaaC1WEqJMpt0IM9iXf4Ad5Uw8N1Ixxo0UPV2DhEHJxIVlnTOwON5Z0gIM
PZujQ+Y877+vtMnFg0uV1+dgPgcoQklgNopfZVQQGwnMJkrvkontjyrf1105
zxtJ8urApNH5BcIJTsU6r4kPeHad1qothnjY+LplGi/tXBNiJxezDytrh4Ww
vcexHv/etKMfZ44r0ZPlb8jMK7qAoHoGKOr4Kn03h2DjUCqmwoJRI3x5wnRF
J84w/0a7CTVZuJT9OTSyOgZovvyMWwrVtJRgjmod/x7qGSGt9hvy/d+ZhDGf
0AuSICnWf1m6sAVkhyiv8/EnZ+ekeCmNUF1GLW2ueoFi9QRMxX4xAcGSOOy2
xu82vRS3c9cavSVtbFcLj1twR/80ot4hllExS1ZW0yI2IxZqR6h/vcDkAj4f
u+KZZKaA4pMZHuHBkZXbRhEtGWPOt/WrcI3gDF8bSmpj8kS+8I+MvXnROAYL
m5sfB/mrVAI2K1gvRmhr+4MjfjF4rHIEEJ+kkuKrskpugvplmix9dpbcgm5S
w4aao49hWAaY8qtWjzz7eg1KE8Jb3/MSq3AVkcM3IxwwhCIba7Q9+bwaflkI
quVLvTO/j/YFb9hGUDz/uM/jsTUpIHu7XYe7/pP9h8lawPX+BGULjyzHaS+I
8/AfJdpFVWxbMZN1ti1GEHYujKVJln3IennxvWAMd+RBzyRNuPFalxRonrXj
1rOL7UZfvp2I+iDk60zONOSD58Jl2iXVS0H9J2bFr1oxE48uT6Xbr/nLkrqU
jsZnLXaSa9Wwo61iyOyqklIkMg1f980GABIpZimHk88vegNZcZ9KXhqaXiGi
BI0ngVyznycwthplMik1YFt4ALrBcqLGrERjzZbIoMeoIhcPOx6LuODHSb/F
f6bLEQ5E7/kH5gcTF9k2FzCx7boRejUaPvugoI7wMFRMJ05mW68bzh0ZZnl+
ATA6Ba6b5TPpnj5u7fi/Bkj5r27a8f5efeDlaYTyZA3HErHcj4S+j4vnOcEZ
i4lvoH6qhoBUwiV9b3+RP46bM/YdpnExUumdcGLcRazcHCcHj0gF5hJRoMHX
erK/56Gi0UzEyh78oa3xioavG2uo2cCUwjQ/OczfS26dXGgNQkjQatTwFjy2
V6HXMXHrPR+fdOCdu5kkE7RMJTF9pYsHObLtRXKl3PqY7R9gL/h44p0yJTFV
nE9HxMZPDAYs8I2z2n48JjuUJfcGloZiN+4JhNnADz74SoVSyHZiM87q7Wm9
S2379XVBHaoPqBvdbFYSQaCQT0q+5iVwPUS4jErBheCLQDVgRnRkZEg+1K+F
spvRkgQeq5AzCawPWPUqwON2Wghyx7oKPrlnPgl/PHqYW+yCBz5Gq8qVrin3
fN9jIBoQCBdTDe1t1RJ+ZN4EDbvMX1gcVS4N1gOlW5aTdpdOIcd5rSPp+Nud
nM+v6AqXGj4bPSPrTRPYAafg695KTvburTAAK5XTq0AbuMuS2h/sj/OcIM2y
z4XXFsnHpO8T5ZeR7toHCG+gnkZDF4WJ/3PYKSfaVvF5cDSn6qdm+12RXNCw
YXaODpDnG0+X5so6fdVzEnqvwf5UuHR0uKnLVjtnQ/J/r97mNRjJE3S7ETmB
hhbQENMSghPt0USYrSecZF/ToOJ3NVJYSoPn5nyV1M7jco1/0Dux5DrfIYuD
dUatk4j4rd5lWjFaN35RqKfTpONjFJYMtBEetwIe3Q5CYq8WjREdfuI4whil
Ca+zUnIN/IHElzRtW4EUBwT2ByVRGI3HHNn09fHG85F0wE+SPqFmCKjP1fww
ljfZx9WtuSE9ffcSfZG3+k0X1KBvq0wOHiKD6O4JRCqhrBqoJgwHwT5ERvll
F0ttYoeXyFdotu2H2Z1KplIj7yVhHVHRO7YEdfgwYVDkZVkH6idGEqqNchto
nK97pSifvPt7lElRS6Qbmi+Jm/b0ogUODM2qCfGT52XCcZ5xkiGnx9UrSIUT
maOhnrXsPz1cKDiGuvK6v+vPmN4IAAUOQgjboePhtteQIWTsqJhXYWthuej4
KeaIRIPH4KZYT82U7iI5hFf9dURJ1JAu0lvK4EGepEjLdkckDxVFE0+C0+4j
ujpdQMt4qKUq4ZBrNqvZrz0+fW5fmMGX0Lw1Kpjf/RJi+9YOf1YntZgkb842
i0bUADUhkEVLDGlaOAuOZ2RJ9qjSCbfXr9myVPKJvzv5sdoCqUMtThIJdDXc
aghF3Xc1IYczDJRF/FFh/FV167E5MCUPnuXOQ6H4G/ZYwsGhM2e+vBm83HOz
/cyPUM7C7p7NWprqNWGfCbGp4ci/FMCCPMoWW5s5WHqU5jkZfVweDLxBw7KN
tjazKPtdrBcfFwEzn9A3Z/++elH4kSPuun9cC6XM/j8N7hXWoqd07bSKKoky
NFnycDZcat8qGECun3aAmjzM+Pqap0itQUDb+PVBSl9NoSKYbzM1FhbWxOyG
IGLDv9T6nINFTn+UD5M9BeB+wZK1WagmVsgEBdwIceAGVZWUYdG3q3H3pEur
4kpsHfqO1nkRMJWzI9LAHRCrq4r+Z8k69RLFXx+ZpFgAuk1/lSGgpkU+JBLb
5/blERzN5jd7KkWR04yXywVt2Smi4DQVimA0uQ08JjDtyOWdUa6uyIUtZfwS
rimz67x5toohHwic/40pPizrsIVkQsYGtmBb3ZI1TQj3xCPPyapsbfa0kaau
n5LCopE4/UvqWDS7Qf6WAfhvh4/+mbEAakZPtbiVHq3Z4Epoum1pba0tIFIm
lD2Cq4VnM+18AzuORiZNP5P9HDGOdMugBOr0zmEiINYbLiQW6u4eLh3Gdp/O
YVssP8ot9/LJhTTz8eBUB0VZzBzYsaxWez3idNz0lH0nd/U6yw5inX+UKYTr
rQCixWhqRB9trOeXN9mQ021y18Qq0UoK/9yJ5MnMUhsvKeqXV1Ypm//QBDmN
+8z5/s3AhJ9BS1uFWAKruVsrEtu0FDrZd1xUAhs4PLJldEzmjSmtvMmdvOMx
fd338KUx8sibRYW2a+sl0zEeARFzqBVd9eGJDrvrkxgyZAIEUjjRy+aXASdU
dLYZ1jnp2MjZKK0zHNRhSwk8RGGZxZu20z13C7xe7s9P0TCHnZ/sGKmQR3YA
SR4dUNZv13FxGuW9APZExz7C17vYEinKWlr7El1/ts/n9yFoCaslAz7xGVL/
t8heb/6ATSqTSPbFgNaHm21X24W7gGFPhjr9yMYxsqt8yusV0zQSCOcIzLJ5
GTWIVYc5vzik/TIyRk+yx8tFciZe7UQW7hqnHgnWNashRlF+Kd5UPUtyCOsb
T7eYsqe6wunpJo3D4iZNpW5fhAX1p0Y2wrkCDI6UUqiGZlGuwRvBsCFJsNDf
OUMH3JyNyHR9YsKnr6iVDq+h08SCw8ouGhKYThz5L1WI9qReiTGcDmYqcMBi
wNONeMGoigE2TdA9nzqQVfQNw3KnADeZcaZzsDAAA27QnFpK1qQUHvBBTIdZ
Ai0mMMa75uNnQ5NO93e5O42ZkH9rOFEV2VEHe7DbU095floT3Jon+mKcs7Ns
IPu/e2MnE1OI2myX50gOjULwZj7u1JnGQbYSQ9kOz9D9TkMxdsgrL85LeuLQ
oxKNQk0vOjsAxQj7RTfLWigvq6gE2scmyUPjLTirsBEYna/e1iq+REuwpcvC
Eocbp15xh5Lia4nfZO3826s6NM1yJPZeMrZdrb/KPcGkeAGvdYbIoDeGZ5ni
QpG7yOZerTVtZ1WJN4cuZTj77uaz0SnUd38JOU5mw7ELtf2TRkEJWk/Gz5S4
4Fjqew7lnNza3NkNnKerbpKjSUI6kCaNkM3DicdebUQ8zOr0MUcVOLWchTW5
iW8J1zhG0qsSONQt4A8cbmEhITVrBWrC3z43Gj4ooupl8sZochPls1xamhan
0B6znQxeVHCE2l1ySYGIXNkXSKASaIQJ46jQHTSn1e1RYWQ1ExPz1vqFmBOD
vFfXjXNR1p7NjUt5vGZd3huinbjOlJ02p+/GnA0uXT2SA2O7MzDSxdHkR6Uk
GRrlhS9ib4oRRD0Vw57VKFiFEtk5PHo34xdBwNQFa6LMTh/vX82fErNJoLYX
epnwvovlJK0Y8GGts1S+mLL66OsB9HawTG/z4RJrKuHZH+t1uWbtmTjq7HXs
nM5591Ud/LdWnX3ifAiJNo7TlnOr8cu7QQVex5o8CxZ88OcS6QAl/tfkKmZN
fLvofgOqErg1XYd9PyvI3oRuIdjeSDX24U9vh6b0KivFyccT0YfeRo6z86Hz
dq3KgOd/Rf86RtZJrcmNV3ml8ek+1l02VbYvVCz0fr5QkTylhtzWfD5IbCDG
A63kN1FTeblSGTqjhSCOZsiiCYb8bZegV0KN7j0ZT8ApzM7ctry1SWZ/B8Wi
FaCO2WVSKcLEiFAxnsseaCzoi8J3V1qNlxa6T79KNWorvsx/VqJlpbiyWNE8
y782bib9FygjBbu8lPfISV/NSUljUEaQ5tD97XOWYBovRiiO0ZOwpJS/GWyL
AfcWSgLkr7fM2b20H//DDCZdeOgTDgzco+OXhAN/WF2KwY9ggQ9hlQL90TFd
KYYSGm7bOnFxp5ciLDLqOipAQXVRPfHtbpWzJe10XBS720DKWkNvHwDweDBl
Ye/wZD1YexCPVDdxjf569CyAOnPz0PpU0L8VM4ibiGaRm4brHVH5bMOInLOu
+jX5aYtV1lltPFLoiExKglxlDm/AsY/2ksItq12q2mscfT1mp5mFHBbMLZOf
kxjpi42VPPy7CJdacYZRsgkv6oWyILiR2siKccO/2Vf+AG6j9jIb1gCaUUAY
jneOFWpMv71LMRl0oeDx9q+st/cATLxqoIFerhIAObnsIRfY6nyJthtSwdb8
cDnJMsWWXjlnhKLIIFO5z0K0CsrIGeQaqilyn9l+fVshn1L/Bnb/bZAndzBp
di76S3qx27F2IuhdX6txj44rOqTWgh8cGsc/q3NR0bqyWkn7khG8vf+qUMJw
G8OwVoDQuZneG1Q6zcc5Ihw51EVDSgMy/KKYJCRYZ3V+/ZyiZPSO9qbKiwEf
LrILbeVnW5FP6YjqeFrhSjHWi3qOTcYj59bh9Uq17Lvc6WA9tymjz5fQjFvt
/yXdDT5YdRk2m+kKFdLyQ/W2IY+dOKxYpOGK2NFykfeIb7zoGiThloAcPSvy
U0+mF8NV34+w80xJs00DUQ9TnHIyLEQFX+0u2jciIsOHigDso3SsQaYROVMR
MQJ6SChRsoEo6qezkTenJUraX7EP6hZF7Xjxndn0c8uGD8Oi8nuPu/eHY/9A
bpDyM99lFRBgFUFqfpuUU5/rfWMFZwSOPBUGaJ6KnFevD/rgp4Pur/gRqgXa
xVoLh3hdHX0epoQcFvRoxTH0IeylZJRBNDrOMk1Ia8+O7n5wLdGDAemPCkKy
JIZKKFhB7iPSxqMsBi1vdl/SMpiZ2CR4rosodOhlKgTEZy4r7CmxUHVnt8Qn
QY955JOWjW2c/LWujBjfTYOnE8sGHIh0IVO1tNMTk0duIM+oKP3hjMZnb6ca
qaXRFCR3zB3v2658TSUK0HNhAsHP6etch29h2BwA5oBtnrYla71ZvZmfpud7
kwbPty/6D5x/wG560wC838AjV1hujtCBWLnzGaeZzkW/SdrZb+A1PTKmPiJy
ysywCAYXBwXe2Jh7zONZNfmTWqjg4zgd3Ir8Mb/BP0Qskjyqc8GlEilps6XR
tbriwk3WNImCuIvtsKFonJCXEtWZN5Qs6z+YXsRT/0kDokUUZEZbmwnts3r3
A0ADKVd8KVq3VxZVqZWTYvU4pqFKQmsQGZq061CcejU3F3M7ZPGai1Z5r75f
8BCom3wmXz645AZezLMd+qAD14a1mKwfkRAIvUdVVwD/OvT7ngH1hBAUxDiq
ZyYo4FLfXDyO3QDu4+vvApgtYCNt7ZRGMETADPWV0LSpVMp6yThFSKTk4hK3
zf1D1s/0JhnA2z25DATrougr/i9e5JcPRjAWtBLI5cQO1BTLnTCJkqs19gkW
TpNtBHKyA69nc1bY4y2K++cTrQk4D4ScS6NjBtWTDeoacbWPefM3KiH+aOp3
HlkvU9KGn86Tqzr/ovbn4YUX2Po5Z7fZsy534jDnzhEGYArIihahJxMdnQCW
37IXXUYybVqXCByRRHBVEC/H/uxa2WRWeNorhLLzEa1mYytT9935R+eCzi6c
ngdmT4Unh1u3NVujqNzma0C+a+0SYR+4MJfMFFD1O9AtXtBjgnV5YnpFEzuX
wQwchAtHBc2RsiTjNExRqg5kCPGOAS+RNtuw1N2ETaDod5ruHCXO+AHTV4BH
cj3P30lV4mT96HuzXBRfozsToAOSeyecNuxAJzZyr8fQ6KfVxECTTiO+/bmk
l7ByMM8CSYSeSWzgW+VKRxEoi6iW98SKmRMCBj3P8nbc0RHEteRMD3Nn0ctW
ZnXd5q37Jcp6VDcxFiORD/uOh76T3A+ZrRwveFfI7hvt1wiMCkLfQLj6COPm
P5EJDr/wscRCgPIMt1e/PB46s6Dd5FVeM3F6s5k5KZkyXWp95HHr8OdfO8yg
WoH87c5dAMAuZXfZthqm/KgGTpDxllLijPFS5BVB5QsE/r3JrytPyKtGooRR
U6YfT+rthoVh5qk1S+KxLipLCI/0/ECX27Gho6IgPoZchfSc50XcwFeXvJcr
0IjP+6e4sGR5NKiFOcvCpW+RMgNoFHMG1Tc3bPSzdb6P1GmjmHu0nZ2G4OUD
P791fK4V+lEvXVwKddc7F5V6/v0SycMwIBXTT730EM1oo+aAQFge2T1a1HOT
qmStquH/URIPCP3OEBp41E8bfyfYqWey4/x44MF/YhsPjcvU9GQ7G3gKxSa2
oyVXewEvFoPGygRzeYjXdw8/TeO9qq7+jYFUlVPcPCjdDEwKQvgpKRlyK9+e
upRb37tmbxqnBSIvxjeB9fufkG6uK4X+nxcf6qvgOg2WkEzRcrpr9HtwmeKe
H+LCgsiRxJJNvBqXUb08ywk1pDA+D9WfnurI4RyPL5LCDVtrr/A1xhWSNJLo
v3hyzjFcfg4HIoana6k8Pd/H8ei3UoIkRVCKhWSWDsayk/f/rCoxWSaIT92u
aouxDUUjp5XNOofBKgl2u4Obnyshuh5fx4m/5JtRO4xCUKOYJLLzBGF+hfqr
wyRM8PBHwhuz/dAoO4vQbDQoyQqg8hOx6ZCABhQQQ4RV4aEzP+D4c//+rvky
t1fqEULUmLxsiTxDqQPaix8+10I4o0RD8Det7y4VI1jIcWg4H20g9z3WKEvF
fufh5aiVoUrrfAADyaRqesHY18rbHC+EZ/TUrSP+qVd4VPscGUBqChxjn0aq
OmI9dWIyp8aeDrPzv+049XBihpreBpDX/8Xk+8d+dEE8+RdfJOnjYGKXIKgW
dCmHqJHlgBCAXGRtSjN5s4GegQbPKNZjqqL793e01lSHnHNr/cqE4XVAFWg0
3sVorVghpMN/BzvrB6eo1gTKA7aE6KITtlcuR03vcUPoXxSozmmvS9i848Cm
zZsT3DtGWSLmXn+CJg3x4q1m5uMhgroniq/DAD5c1gUzusIEg8BngB+De9KL
traFlO8H6+7eWuONH2mEUGnnfCWV5ykbLj+bnAaQzoIym1zcWr/FosbDC0Ng
eOkJc0+RR7qZbi8W5d1mrymT2JEgGLwsTnhO1TPbDJzXBZVvhKvHCrEWzytP
Np4cbpkoG8iG4ZsOi/qFOxJa/I61L3Kvn5LNm094a+afunnBSJ/eFcn9NJKP
W8NA2hmiPGFnh3qk+a2gb5jihUM1bzOmTrS1R1PnqB3tdyv0Da+4NhZoSQy6
NWoWS3hy5hrM1Zc2Nz3PsDhw2JrGGbIERfmkY4r5P9iNDECVPImQ7+s4wUaZ
AHNNPLSYZu7z4yEC4PwX/WXVvSwH4t1FKNkFwGCUL+W50QCyuqp6fByY7b6K
lkuAdP+D7V/eq8MbLHRk8wf0RaEtgQ638+COYo/zO1M37w4h62/fwj7cOhEg
Lphr9yp6Q3zdEkBPXpf/w7ZzQhheVGyCNBaQHfQqQ4EyVGaYxZ2tga/lz2NT
gm/uvJ/zEDtXIuc9OnCbMHZSu2crAuEkyONZ85fh7VfZS2xcsH6xeVo1ixpe
wIOf/cEhTwfKBgmox5sndqU9Y4ogXJP3y1rMffaSn6cFUFdWtCwGcF/xpOHt
uar1ydDTMS4kCQFd9MZG8m6xUMf+I21cx2fByf6cZx9HTJPTSEfnf2mzBlzy
1oTRlzqVXF0Lz6PKUsh82Qx2S4ADLW4VC7Qc5i1fJduxNY1Cadu+V41oxbR6
VBBHKq/2t2KOh0x5qUln2Lr/rKlvuZ+ykry73R7PJDLGjjtIcvNe6WPb7P8Z
ipEBHd6nf5kfvRNXwPv9ouBCPEH33676nmaMyv3N0jsi9eZ9NDIL0AlgdHyN
neoOzxjyySigGWe7XwBkwZXtvvNSqHsJgwnqCzmJp/afHEQe3OVORj65w7o3
577GWxfEuhsWao8skDSGHX4LGgimsMEXDfjW7SiWEO9MYVSkjaDKglwh5kOa
UNugLI5f0KMIGHlwBxPuFKOIwCExTmMuaU/WAFVgmPFtsfNi44J0Ne6fGB/1
f48EeNM3HtBDYQQ/tZuNAtGiuyX0A8tL3QVbwYCOyhQLxYvEkM+YiJQZr6Q3
NHa8w4g8g4DGoBNxL5RkDBbn+2h6sciQeH6dNKaQhxne7bUobNUG+oI6WQbW
zM74p7a5Nd3RGUD+beCVpHzrRmPuZp3+hSMvv0hPzW/GleO51DLM/7dvLCT+
fwDbaDrfHIHoU44bw0GYRqqDnjjP5JuyWpIZ1kmqDU/Qg6xPLNQC1MZ9znRz
xTIzsgSaL2DxmJZytDfOD7WcaPgi5LfGDTc5ZPpYsvgY7FipVCVFcIohEz46
cHbReM0hCbUMYmRbIRKYSAxhnJd+Yc3c1UN9mN5v9z3+rY3f692yWKUXBBHu
6+hXlOs+UqXC9cqhMPylAFMb/SIe8908ZbZUx6Bj9AzxTbUewUJt8PhCUzyM
eiETSCm7162AbgS+SB4IG/vp5TDg+xYHfAsy3tYcNwsH7KSk2LE4nW9gJ7wx
xyhxX89cBQ98939mMFBQUzqxrtBeLNCDkuQxUN/ofAy2C/V+yZorS3V3o36g
OU5nSgAUmJ5MjGvkkPXH5NTstry4kzphCKzCcOJKjhzwF/K6VpKDTjT3f8L9
fylu08NuqL62karPQU9lE0AjaCwV/DcW0Rt0cnO5wUseNtBDx625TwLy0I3D
taHQCmJlPSIKuB4IwpRExSRyIyTtb/Z399XKBKA/g+GSUWrx6fF+XoG/bGeh
nDPUZ7CsuBEE7YB2E6HQHmQJgN761CaTbGWHSJz/D29mCsfa1MdoA+BjahQZ
4kOGTSZbNDw5DOKTI1jIOzRnKOwbiunXNk2N6jo0EZztJxu+8pR1Bl10sj53
1xZNOlRLRnU8sR93S9qruMc8VTfye7si0Kq2ebsJaSt5pTYKphXErQRsdiN7
KgV27Fa4jBHeQ0PFHLObXP3Qxn5T6DzEhfnip7AzKWSiY6JndSU+kXjXU91s
7gn16a/nkfConCytwKQPnQWCNwnJ42rkhbAIPS6lHt2j1dZWUmrMp6HujxAr
6ymUjD3VYFsOGfUYgK0Zj7Gu67gjvw/NQEhVo1v9axlLzRX4YAJ16A6jWCAR
MEi9+73UyqVwp6saQ5HrIfYXnGJH+CyH+rYFIX/QS6do9Yflja3cCcHrXHfN
3/rIX/eOrFPQ1xMSC0F+lDEP81VUBdimD7cK3nRPOlhihpXufWFp4AufVG0t
nRbmIoup0NKZKbDRIdb8TVtAnoWUGSHdYCFsNxjeCM5YD8m8kYwwT8JM5WUz
6IP4LWNG1IN1x8Vr5xZpFY3DqHqQLtF27x/duidSZY8cD9ImDoRrONfuAhh5
XYJPCG35dQw/ipqeYB/iEMRhG2o03YA3cjneGRRHybpOhowCue3c7ugc/FEd
84LaOxPoyTDE6H4t39rmkKMIrNUK1TE9tF4Yng3f4IcZordsFLRs/5lcP0KW
s2ehc1ItyiQ5cgvEhqX0beIU+KVSr4gOjDbx+ToaCZHS4WeKc/uyF5GfPJcZ
SuKiaKeDe6joR9Er+swhd+doOqu075/kdKTnsSO5me0udrfx6ABJD5EZ+2AO
RXOiOKqU9qiik3xBzpDB7QezZUtUc8xVOe71InwcApOYVzQEKeakDT6l9Odt
xZBxheN51z9UUiRO5IcVbr0siWi6yJfhF7AxJNVjs94O0HrfaBNthcsz5xTV
IBupH/QwF/nVQHje1bbhF+JiOsq21jhH3SMm9cR9RpBHup+y0v6mmk00Ax3D
dONW5+3IsL4suLZ1w5d9dK+/+SIseM4fDNtOdZrGcgKtaaSZ/sC0aF+byI7O
nT8x+DnlYZ7ruei60XFSP958AtQ+3sQ8MzOaBNlNqgVCMUipMBMu3aw2OTiq
9byHtQFUDAEYpMek7Rucmu9cqGPdkIOtEqN4xT4OqB9PkNHeb202k25LQNa5
BNYr13dXfvQSXJdVeDZ62HdqK2/Jhs0bIsYypXqeX9NnKT11RP8oL7XBYLsC
WPgtX7Ixk4nKFzFhgmb/VpGPwDHUh3GWs0p9Z8Co5bvyEwN8OVUTfGdHuTx9
/WDkrthSCQOi75BRHk3MqjGcz7mtja8agSs3H1YitFxcphaOLt7wVcOzGMgq
rkSoBxUoRyJxyYRpN+L/KfmJ8bcKLflBYG9w3RmEOsIRvfJqOSDaOJdThxS/
ZYVS6U3zAxsziMEA4+hzUGp6u0i4+3d6ZHU7p6lqklOTtAgJvnNAGoN0uLg7
qyu0MUNW2n6Ndz5QrUYhOijcmg2WcKNMkj9IXOpqBHfcv9RkhCdVUvBZvERK
EdLE2gHsoa41veFNheLpN3ZP8SSGnqMq0BFswj3HvPyHFKg1tzSFq4jN+mdT
nH3w9YVOIUVKTW4V9Xmc1fdmlXQB4kO2S80Wn+RmYz4yV9mAu60u2eJywtR0
qSSeMwBj99BWI0q4hIxNCEJdKgZXi/dG62m/ZIEAo7h2Zu/zjUn7m6eX83jr
gra3LMcfHYF/g30JOPG0JrYJzH7/Zx5+nCJzDt2DzyMNpyN7b9Kuu38KxSSN
xjJM7ZouOsf7PR85WBdKir9Wytjrc9WCtnrFvwxAT6puXmuKkpNFoBYoe0P7
nhGByjqVoEdjH3bkCCDaK/Yok/4K/pL2jVpDTyFBfnKJ2CWkKDVACMt4yzcv
Buexem25oZ17D4IKQiYNnIKsKAl0UxGSZjZv3FSrTtPtxEZih8VoM6qGUtRt
UhSAuvlbIQd2mGAKfhiir52rd48owGdy3imRT9SPduoAdLHtayJR6d2DKton
2MvJw8gjSU2Dpu5yFutbOvc7Auz3diANtQaV96zlORyKk2K1E0ZgQNZmI4Bd
QRRsZ9r/r4VQDtCs0PajwP+qnzzcaxGDrl8u/tNf+WxkaQi7MSa+gP294y+s
UWhKrQnCU/mNNGyWDBnUAjfJKYv2SoVzoKKj+lVApTN2S1lOkwriRLij927j
OPnYEez5DWMcK2YI7L8H5leJQtsbAgpxxAkb6g78yg6pFLqyScGLM5ECbNBE
GXsCCCyAacWjLK70ek4waNal12eNXbmtJIMPQfq+exk/esH1flMkZeAWybTg
tPnx6478PH9WZPGcbLTfqn9hvqMg7aEdRapC4I0WLFuZD+05h3iXCwYHFfy0
hZ8ZHSip1s54NHSuLnvS4Zkda5pZCHCFchriwEt95nPjZn0jgiEwGHBmmlyU
ZVxmFm/owwEmqn+VUi4hhTfe8Jf1YFv5r+EpkLLThsUANghX1Bnu+CD27jBD
dRS6Nmn4Zba1GrS9pbS4XPezwxEOT/l4AoswlAOJhEbZMUDul4B07B/I1UWz
QBjn5xdLBpC8fmMHF/NmXo+nHQ9KqgLNbHU23qDJ/6gYopNTt4T4q2LCpNtk
pX6V8IaxI1iCScyhYSZmCC/vs2LoCXoVMFnMw2N1gyF3g4KDWf0IkHfmvbcv
OZHcqxRVkkirGvvZrLc7fblyfKnMycanPCjJKhQ5YbTUXDPeV/zKuI49HUhJ
WCmqftiX8NFq7VVHFd3uCWwQ387sCMeM1H8NPkbSFE4Dk8K2vBUO78/If3UD
SvdCG42WWzN4WLRqRdnLv1JkiF8xYUuAMPAnLctxDkH7p0+11i1gO4g5Yyqy
5XRU0GhDf3Y2urtFFBsA0SN5BajViwivkQPsP6HBXzj9KXE1Y0Q/F9PynqrS
LTXDyupdf9d6wz1L7v82Lcgow6FI4zHCh9wsRTNsNwU8iUdJmyw+IFDbTVA5
tlrDMYaiqGFVdpgQGaWXULeApt9TJMd4ea0XMtpnsEJbu/lrBETmUUNsf+vg
4LmQYwhJSwtYrd16pVfZK0d8mNASjn+3KJAiaRPvYXNk2s6m2rYRkEDof53x
44yBTFn7uFfgj2G3R3UOQQw0Fm0EAJ8ACgohp9sV4EIIl3xnDYYaBF8mbLvG
3/7sB1IFrYy/yAJPmsXKTwWgejq1x04OoB53ma+Nb18XCE1FzV5HSDl+vko/
UMDyqOMXaCJOwbbgHC7XrMOYoM2JdRYFOauJCw+GxYb85uVNpJvHfByONes6
Uc2fceFKRq4WsmUnQ7sshty7Nx9A+DOh74Uloy+AEY5iSZjyv+VrA9bW9MI6
B+x80f/xSDRHxWJaRVvsGP74pBOiw5eGJz2Q0zFvOw3HAf+85M1qfR0YQDS7
/SBZWq3GdKZEFLdWwbr0V441bwn9Gzfe4SLTE+27SNeF7j0pPOrn3MnjkL/L
ycWHtpP+EO3w9cZiC0M0fP0piYlEfVyG3ietRsG5quku71yhnaLkMIcPSSlt
byu1T6q0M6rat7ujaE0ZKALqLDPEyHx0bskmKwjvDwULf7ocU9trsm2htUlx
LrWCCDiHt4PsRnmU17RBy3lX2PpDcdG9csIbRpe0vHKN+kD66yVrG4DwVU9+
b4x0Wb2qUS3TROQbyb1UsX4RGNXdymUxAKx2CTwVcko13n6PkDLCriFFWmC8
RMqxWDeMhou9T/zaffLzY5OjuV8iT2nY7Y/c1s6trXME31hgpMYwZACC+Z6L
bRzDGZ/ySB6x3f+DiRfTsdP1opuYLoHh7h+1jEeE0OG7hrodo5SdXrUFzRy3
ihCj3b1c6xs0i3I6IwjQ1naHgSRZdV6WFn/oZft4q3WPbkO1atMek1Z7iIZv
9kzhW2b92YfNitDG5QrX/Qb+I9xZbJYWRiboUlRheYg+v8P4D1Unqh+XtV/O
M5ixnrRB0lNg7n+9WfhV2IvpSC53xpLfyR7Uf+mnXE942fqCV9jxvVxNhUNz
p0L6yD9IRSUPURIhnQ7BREByTO7taXhPQD9ofUUMpKz28iee9Ds6euYuqtrs
dAG+v8VvGUnUZD9rpqJKfSNCLde5FIsqXXtBJ1fAhZ4/fTcR9GwzVGU+Ctv5
Bzts996HjMdEF1ji5+LeagG3nvTCNOxtdTn7EYd8WTOZ/ZKU/VOonDJZy4o1
90hn2SltyHdj/xGCYa0RtAcbF1WCSOkR16z6eVTTJCMuGjSmvppkfhkzpkdm
RZPLwUOs0lXsgpRas87zLZypd30vuL4XmMpDja2ynvDOOxZf0xcm/hZz4vTu
Ke+Gfz1DhDWVsBv9bvytIZpjnuPaFIwWjoGIk2rvV1xrA9S2vNOTflHmXFH/
6keJNCT96Ib1edaTN8AM6cgyyZmpTiNg6gLFv5kuerY+A+dwpIph4gYK7mrL
LhxDaJXd5JL501KAJa1SVUkQntj2S0X3dVHrCMxHQDdIYgtmEe1mvBiul6zK
eqpgCs7TZuKkJIiPV0YoxGnIt4WQzIDAvmCE6KCjIw3xk0oQ/APLVDzqAVaM
3ULMtM4uQO1txQt77VZ3CK52V+4DBmEC+WMcKu/hgSuo0yaf8LOXGwgzjENc
fJBhfXKHJ4vwOP/0dXfJY1lJdYz9GNlrzroMfwqJwrG55w6sW5n8B8b7VlRD
gA2APN9o7vmemZT2GzwkzOf0AMf66rf81NHLHekLCJMqpiTaG1d6zr9N+BF3
HKM4idBcL0TTlesiuAhMsM0xOLkHOWxVFPx0g/RngG2Fj8mIri9032iqa/HT
oPjQfpcoZB6tGRxk3RdAOAdO5oCaMRpnYgyljjKhC3UpMUUS9ct6aua+G7ft
5P7Ka6W8vkVqg/YGkDIj3AJZqxTOT2V1rPCBildC2klx5rVfEqFcychkVcxr
3kOAkp5ayMj8caKbnKlImZuGYoD3bkBMHvgn+dUWTIWo83Rq6SYYQQcTb6iN
vgI0tbHcYuwms43E1Ir+eZ2oZmGO+FZmJZzibTiIAy6pq1g4YPvQ/XkaNzzM
2S2fUJ+PMnVoPm69kmcmVi1hIRruWs+Db9DY7v7UldLkHESA2lEw598eNNhr
BZ7DPHFsAVCVxEYQv/3sWx09Iqabv+wtNIA0RG13kBdz/eiIm5yBAL8BOcxY
SY4IMKn1GSlVAdwHI0MNB5kw0ZrAqQlqyuf/KJMgJau8OQ3gRZX28d8CcWjP
4wSAbATXJIL5cdnI89QQ9DDx9aSUVMS+LJE22MCh805AY9/1Lx6/+O71gZLC
meGZAQ/IfefUR9ei9317SP426zoc8N4GarQTBsCmybbfBTbwIfw6iAPXzhbH
TBxwBJXNDRe/1eI0Rxn8FhnIlvhOuXRE1fVif6L2DEDdl7pQjrHkY691G7TR
gfx5P9usywjwdgGU8gOwzJ3Rjqok1aNhsd576ZuXnyRbyh57yQD8/hBXJZE+
R3vOeZL9i5fuP4cfAEaPIzw2qFuUugX+PQxR1eDMD+M2LXTAxHiaWJQZA5n6
pcBQUXy/Azb0qVz2wqC2Cc9wjTQ+5AJ5p2/tPkebHVAtFv7qDnVMc8TKCLkm
afhKwPjhexBik46fQtRVaWlGrZg29hzzDQI7eeHXR3TA0CtpAAPcU5gcDToa
FuAZaRjSOambe6tL+d1tpR2t62KRv0PC5Qm8FvdRJiSWJnK3H7Lpp3Lv/oFn
vbi2gmMsrcqT2CtzGqB3dqlTtoeIuxeJvQ8wWRm+hxmGbvrCVIEy2pdjcN8c
vtEAn8MAHQuZKZgmgDjDA101NbuA17yxvFjuDgH0/WRNPnBpXy9+Uc7xzFmf
hOvni+jpjsxqzttgVYvS8FKBI0c51+G4IxFsC8zxXQDoh70YcehsPAABSJTy
XDUWi+BdM0awO1ARcxQvPkgja6rXEcU3pis316otN01vVvKHGGcGQqey6xLj
UxljhE1XvGat3YcjZ0KAb6cOYb5rDtMvsO9g9/GttF8povFBVtg/wZy15X3h
2XLBNBegR6YstwBjwlzvyYteNMEGOGO3NRtOUulFBUF00v1VV9XkE7XaZG5e
vHsWOkdjPwfzdxUUICOcYKCXPXL4YMU11Y7IUqcKvDc0EBsU9pJ9TWA8dsqU
oBrqxKO/mJTf5/+5Trjkk/j/IoY30I2kNMQPWXhVz5brW3Rs+y/wmzQ0dYTZ
fPq+MNAK2we95jaSfhiWhdgApxwRZySgSxaEveCRupL62mPqOfjUUkcZM8QE
nMCzsoACX6R0olil7+1TrR7Oi0a8drcrCa8wB2NGN+siHFjPwMJ686agFtGH
fk0AaYeQ02nJc1piPEMQvE+JVqXQo5NKjBtVNa4KZFo9QxfUmmZ7DsK+Vxhh
q2DNfUQCW+QLhH6xn47kE7tzcK+jzW6H4VY8qn9iibtV31wJEkNEpNnkZ+4g
zqsZsnj5DqK7W+gSxJxAEsC+CemBGmXhHbdE8yAtfZtRFAe40K8rGtBrVYNj
fmG0ttUad0Iq/Jlfp3J+2iXeZEoQHJKicBV/08RWAHIkhxsDfns+c8Geka24
USfxCGNefEKtwZCwZdveqqa/YBLH9UuumKnhgLYChHuLewmhcvxDe4XQgb+0
oIlQjZEKBNj6JOqKJny65JiQdXqhusEGnqFs+muJrbP96bBECQdl+kvmfdTC
+dMbIc23pgV0365EYr7U2IQiPmYMDaYvzrsdq216W36ErpZhQ6qY0clvGAW3
z9nNAsS4GMSqfc9gvTOxu7Ho92Dyb91mWU4o3DmGoTvR1YADpAMlH4rj3ohE
JG56KwtxhPNU6Yw8V1xF5PHKP/uYBdw8sCX0OTGPXKP3pXtDfQCfDu/Jqp9R
gDxsANGys4SZz/zV3YyFAJsCG9A2u8bk7rtiHALh/C93st40Nfq39UwLDU0s
1TzRz/uvgZt1wGOLZbMjtTyj/1GzM+ehDEUt8M8QQ1pjkoiHRffM8MCmz7nO
Yjy38ztGx3KMtBUIN0YN8Odpu/EMmKK+5DGq9DOjyrleGEZp9xMQNg1YhHg/
/4SE4rCnT8SEDMkTK0nMbU//KMcNQRy6uk3OMQgUvUBXogwxxUDkEo48SQP0
uDCj66Fvzzz1VPN+BK35EzY22kEuz8q8yA4RJcnrwt42EaPV5s8Ao7J1vN+M
mS2H3yGYgJE5lmeXnNgTmJgzEzEckelsp0lefmNUtBipHHLeR3wZtz58heyl
3OKvAzUhCbpKLof5mvV7KcuiBt0p0AKVXW3Rk8weiYmqIYtPnKUOd8NBhuDJ
NoKWojNp8baTIE3hDuJlLfT402gZRZQUkb66Kmae5tx8ZBzklduTfZO8j7hs
yEYNER3VPcelUGNf39BF/KTSThRd9f4zgWBV2cbbRKL8Gc68SgRKYmH9P9IL
wgOapHt9CGNwMpwZyhHMHu6Lsg76gp1TmV4WLL47MDJ/MkIQh8gOwylQglbx
fZy6DAyh4YNpzflHveaGWzPnayFlFXumMDtHkLHJAq1B19fddyVKnF4YDL7j
/G2hAvMbpZpnaZWmb6k6zI+CslgzO8eDSSMVV3MpnwsgOxo8IATMBaegL3PI
o5UVH0LoSNUqCUCcejHZK24ks4Ygjj6wkjk3JvdBr0mrHXxfqGpNoEtlD3Vp
zCR/a/ei/iSGMYxQlI2KSNApRZ/eeyI3ITDffWtUn1UVxm164o1D0RWUw+6n
KfLPsi9qcQpc9nW7ivTiG0a4efn1mVNDR2Vw3BCYijyb23fkkBm2BxZeGRGm
8RdpjU8R0JhkhUEniYHMVnsUWSf0SWN4y+Ct9Sqg8jrgGIkK3aij9L6u0h91
RoV+EZTJulkZnARCgn+OtjNvdBbr9j7vVBTvB7XBCQkFvX5zvxxRaFiM4a5Z
4udRn4ZKHv5so1xhShWF9FIh2hK4LqaynjVixnB2T90ursuks1wwhe2REyDU
iV2TZE8PD3tN9KWVQ+LJ8WnrEA62vwW/m8nIgCkLUxmUk+GoeCw8aCpddVbb
MrGPjIvoKitiroPEew+qkKpKCrvlOFKFhkOi5uN1FynQIF6vXvs5B7/91llj
8tZ2N2eDi83H51hyfDhXwSsweQKbD12N+pTxbrmyhFjI9PeLjhNtcuViMjNa
kGyH+7vt9ATWHMlPd7sDzuvnbPMf8SmG8HIo8YD8k9zNnCCsTbbpPzXUrusi
VYizGGIfZcUE/e6p5X6SViPIbEH+H+XF3A2LyGHhg34C4W+74F7sjd4WrZ1U
97gj89VMbrlYKfCOBEJDI1zuOkzs8B6mUvf3Z77POnq00zVL2t/AV9+2Prvy
qRE5iwyIOUMkgHw86WtVR/yF9I2AZ8McU9r4pJPfN5EgAuA9H9srnHtOhp+X
TX/3sDK9ChKnyOAeezWDffBrYndCE6sQU1cxRVaDhUacweJrjfGHNTmGyrdR
C1u2DA09Ijo8k6rgyI+hcgL7dsDkRetgpeBrB0auBXDjgLK6XNlQpmLfkwE1
kdqWBl1op8lYJLdEXrs90JWNZnMROmc8kuew58AaTzifdSfmwe0DESyIfCJ1
+02z2OdfYiRV/nDADIOBr/KpfBJgK7VvvYwgVx7LE5b06I1gEt4tgqy97vD5
lzM/mbFQR5BqVJwL65IZMvdT/waAsaF4WEU3RMVPBbPVOtnV4NxGHcidd+zc
MZMphSG8BzSk9BXmNA5GGJSJhSVdZ35QkNjM+DB2IQ5YQ3jo/xdnCBanBS6L
amDpm6X6xKM660PZM80oFOFY3UXg36FX8QwbKFyJI/jVuZw/nxPB5+1+rmwZ
hj2HwSDDWT3sGuyWuyiRtdNG8eewf415Gd6s7czhnO/jgZe8sCTjVvXppe3B
Ns+jrmOiBqLEnMVHp5NMvMpgVDUQMyPjtRncWdpVcXQsBW0FINj7rvU0DS/w
N9c6wRkW+cn/mTixlS2z194q1yEarmWIw0FIXlk9wp6Baqp25UQohhozs0p5
qOTXwNqv7tlpva1zqc/Bw231m9tJyoJ0YLbQv2jtOCI9EzClEaLrNeh/1yR3
SXgH4cywb20WdR8cPugheY+5p4GSW9rNSaCkwcvEtW1vyuz6lmDWNnpv+Cqm
tezyNZV4fNrlUOlFfZ+gAWKwIbj7V5KMo6WYckkmaJpQmpuyJsNbbn1PCiac
Xi6ayq9HS6N5t3MPK7nLAOaksTZK8qYqAqrkb9NVuFW7yw7Wwc36ETEzG8Jv
B0tYXL9dPwHic3mSxy+A6u9xtPbUSXkFtcJo8S4PKrDijp7ckx80BRTAZc4i
ogVcnt/VzsGYFu7m4o9i6rDrfOGDbwByeEm1LyufGMHeTn2F0wslLXHC5vD7
aETX/i+AeknAEAugjz1lcMjfDv37gmT1PAWkA0MCmbBIdtjqK8q9M7lcRgti
4Af8i//JJNxdubODR6evVzelAZq/U6e6j3QPmn5Os3MuUnAMLSGRW437DEiR
aKJwIfqVHq+6pcTBxWH/MLYD0mtd76faBJC1+Tq0Mgn4kOiGs0VQVIMdKyLb
MQSheRnUrmD4QVec/f9Lq1UO4j0XI9PlGyuvjuhaSPYVoGmQLpzJkE8pKGUU
I9C6s4M+K2e+CX8JHxPlgqQwT6VFCjrUuzkJsYvISjZE4al/myyRMuDXp9dl
fVMaOgF6gRsv1yMi2a5375rBRvwrg+GZ81mHUy7GQL6VaKavPEqIdi/wnhj+
jZsuLZDMhExi6BmUdjg+B92pWkEtNJtAz1gqAK/Quf9vkvEApTG6dYoCbILT
ihp00yfIYrAbw3SPDs+gjQC4188a09ILWQAWOyM1XnWsHpmh3Jgxj/aq20Kh
W9aUGls9N/Q6BY4MmjpbOhRAR3F8e+iX/9DAN3LSx2/X0UzOGkKZoB+mhWZ5
eUEiXMv8OaxSXhec1stHaAthKlcg+wHPoKl6VLmWNirXIjWfC6FXMddjTs1j
dCMRCysFdvqbU2CHeL29oH3LcmFr2fM4Q14gZ6qdu8yHonvxwHNHxmk0P6Vn
SAgg5td8KRSyYzzROoks/NGTflbZXorFB+X7oFMY8WjchURAwM05AKPxVV+e
IFSIt28jQHRs6DQw8Cj65DmGhyGJJtjelo8L2niezoJqz5CtO1Lguafz0W2N
XmJD4oJ5FNrsr3ekteCdeJWgBDLmtANLA/DcpPbDA6IzSu19m5MMa6Tr9GgR
8irVbj14l0GCHrTRmwge+hH/hNYiOajPjFVpF8GlhPBW7UIkSGdvgGoa4lYc
zcJHwoziynFDiPZqyRMIrcS/fCAykbRz+Aje2XhTTfSQBPPS/3WkfAs8d4i+
TV9Jh4s7aFSYEwxAZ/NfApr97x+2bkbiADoBI/GPvwlSSIlbIF3GfykB7R3X
b2rx5p0VTM2MCdoz16lpKmKf6uZe2+1zzI7qxvJ9CzgVfj/v0i4F6oVkUXo3
nbCayv9T6MNSLj6ppR+BBE6DCj5334zX/FbDJ7jMOjDuEWD/qkKOW/k18WEa
m1sDHNVi50igrk//s/wMXxJME3jRxcdzy5GyH3JfFD10hjwWi0E7C9z+vDZ2
iNj0bHbb8RIdO8wzmVcxL78KSkrv2pJ3GhrdASJ8rAOcikeQp86IRExHARSR
8zsGrmPQ1VuT4O7Kn1v5shhPU6A5AoC6F64QWykiD3SeXjeTCKq9YngdlKEo
yCgp06ISuIWpVTBwM4lMh10sh+/UgR2VMBuuE1F4huucUsldy6FyGinliDhf
pDCjLhAdL27vT1BZRf08XL2PEa7uLtO7wcpQn6EvmmxiX0uaiXx9k71y+UMk
f7KKrRbsfpvWK3H7uxeWaARxGlqaTRLByvZ2tE6d2OQMwfXCNlhvsSyvb8/L
cXj4cLqrp6F6G5mG7oXcv32pXCjZZyFiw6xR2J7aRs2rry6PZxIlmfJEip91
H6eyje8ZhO0cN0dky7lS7rloT/rDjzyb1NIj0Y43OPS+m2JnFG1kulI6x1F2
FcRa+gXiuhB3WSkAPvwY1mRLA3HxJZLdF5hp+bnyiyioJFPbnZxyKwBZwbL1
+yDkM8mPYh9kzVyluncvCAgaW1NMToUK4fGohggZ4iKjLnrWfpZT1vD1wVPK
j+/uikdBMtfo03kyOEpzDeKceviBTxaioSTaZUO6kIBIEJwokUpp6xv2n5Z3
E6Q17lG9edIiRdaTpGeWUpUlz817IzC69axuaGVQDxvPPMTox3B0UYOBsXus
4ztaac81o8Qg73TmndW5uFWuxEJGoWKC4dPGk7gTqV64EppmVBTxjrGJw8gg
vhAFTpB4sM1vkTCgwY9CylJRjH9XQzlYX3HN7JVhz+StqGGrbIDiufFZsb53
KUQgDngRV957UA8BdaSs2z8GbnsLIzmaLAfOLU8JZ+tDM2e0tr30Q9P13cup
7OW6EVJkjYVQeCDPLH0sI3vuEFVmFYLPlAFggq7tayblF01ZOMW8mAvenz9c
tGBV6phvvCg+jQprLdfYePUcfi9dS9hnuhRab0zTS1ejWtKhxXkPUvOCIOqz
Faefw9wzJgSCbjSQg2F2C2i34xUb/GnY7LXvWFdeybad4YQ9umFFrcylyIjR
cOkKKHDrt6sGHBCot/bFoCPEKZnHhfqLOsAjTn8gyRKa3b04Dsao8jExV3ZQ
cMyPrdaxUb2Few97UOARbqIH6+/LuuY9ON+catRset+3jWCOQj7XxBU18Wuo
jiBE1RsUGfVMfaekoG13fafeXNsW9c+KE9jsHEsWmLnhF9O2Tvg40oXn+PDi
v88GjaoyJ6rtrhhoJtP36frQ504wk/BgCzVOzPT+gpEWB0MNtjyHdkNVODGn
Lh6DArBsEOgJQHINvrqrEv+f2kWCx/8auVExOJG8BB+G89eoiZ+UzXPhtgPB
1Z66ROhwOWbX6VB+hz/tCswwQTq3uac/+L8AqFt/P1Sm0S+PkH4NI8kg5414
njvEOY4QlyQg3FzB3zaq0ujp3Q8xz/EGKuoLXYyeIWD0mRGY+Cry1c059fCK
y5Az1dK1OIGQWtw3uIEhdQRzEhltAmsODPjC+S35ptyy+S6hFSMIR8x+NQ5U
sLOvP2+X3Ymp47YS+XOEOY6SRL0cA5JnZAZQbTgYnJNZYayA6w8UTByFN9RQ
o+PMSxXkNjYsoKvhndwNRDHj6TW3R7zQMItFC9V6pCUPIYkrFTaVQ2We/ByC
WqzhhNsB/7mCLE1/v1vHqy36bPCc1w2zGa5YzJF0EoLV/t9l9IARai/4yPAN
/fjZKTYy/Rmb/H2uKXlJe76IjdTN8xfUIOj5Dngu9WUf5gg+jpa82wJp45/F
AQl6JPfa5k9tUUEQuBY5DorB7cGPsd1sWOKVPLmeeu0hb01/LyBBXTGqNPJI
cs0QuipB/XVvm3SOG8W8Q21rSmLI6kAH+ryGn5NKylx77mGIXKQM/GYGmjrI
ibG8Y/bUHJH85sFRGoDB7dk00pNKw3RVKCbvHW06efcawMzLbybxZMYYDYb3
tsrJHkuzFKhggFV0UiGhOIsBvmwph5mUsBtWXiWwaehmHzHL7oXB+fuN3gsy
80mtim8oWDOPc+cB8ug5mEfnVPCru9ynK7WM8pUwP4cnY/jgC4Uyyqb00zD/
aDnDaH/CHWyPAmEwXrUC3b92VQXwhHHaF/Dqk9+qGLoMQCTf6xmqtp4JTZZc
ETtu3cPstKi/9KkWRYR5elCXPx8oe+3gvceFmmRTV4jEice4zN4fXT/uILFa
TL02cCrYO9n4uI7AxU4U3sMciRvkZInkGlmcf7xngfkJVvD9lBJBl8AZDIpX
EXfSlM0tErKmK4iOV7T/9rqIO7p/6YjFOo4CTIZlF6SIyvbMt7/6D4L/pjz1
ATMwJSB+0CgehlSzdpdtY+5H5HPNRFWMZ26TsTY4j3PcL2G5DfjEuAE6/9fO
QDhf6Jsg081bIm9anG308xwZIFYz1FT4qGCtyRLmfUALQoEhIknEvzsDMNqz
OJ1tSpWJ0Y4jFb9eZcZzhc4IqVnJwgRaD5JyzejIuadxrkVO4XkZ/iaiIa+/
RC8b2D6QkhMWaDPfRtAxVIZwi5A6UatyK1+5dacdetKgnOkzxHpZJ9hXNZiv
gvo63VqWGzdVOyuNcYe40NaNLesaMUAmzCFs9LXH/Kk9VCrs0X0IUdf8k8+x
eMOzyM7Y/HtHich2ar+LviPq57P6Cxvh5zQefJ2EHiKWmgQsxPjsY/cnX0t4
lnYzphA/XM/SMAHOQ5d1nUASgdiqW5I2G/Unk3LYTFKpe69yQOJ5mDI+Y/Z9
qMoUjo5y5S1VAiqiC+BITrW5Hv+T5ego6jeq0Wu1W+wuLgpKiRXHJRbChUKC
tUUt0DWw8eorpkDct/PGNHxktfAtL0U4+iVsyqOOZ/qIv6e7Q2AqCRmcgyWm
kkakfDJ32JMTGWaWhbvQrkjseFEusqRizGOI6y+zRvpx2yPsT6nzJs8fcK2m
mSKvoch8wCkYFu90R7nif14jfgb3rL9Oxsz+N+wL2Nt6HYmIDFPeB9GCB43p
tSOWbzMa6PLjLQLru+cWNwV7DVC9JA+0MucIB0xZYB0+421pvuKPhcyNvkSW
apoL6dLb3ZK0eRrZjj5qauKUuoyl5Ge1WcYGAirDMUYq1ezucqqP3uwHYfpN
fSVYQK9u+9pkMAGl2/Fxxgzav3tMY7xfsAeo0ON7vaW7B8mPSKC07pMND2n5
aleVflV0r3Q1yWN7d/kmYd9SMGLjMnOfGh0Geex1nSmWpE8w0UwiUqKchfZJ
k8B02pYEUMqJLJFdVEiovwmI3fPJs/g/tJ6BZyBs/8S6iXfbJ22BC9GCuoCr
e8m+UlHrQPTPqBOsTHZ2oW4yLG6Ls3M3KO3+93iq049F6cgyErNDxZMe89Sm
0jBBKZO8nsTcL/uj+BLOrlj2BiBBFZNvpaFI0uyBvJbZX/j+HnLehGqP60GB
CQw/40o+FC0GD5t4Nt7QNA+Jqb7L7X0W6qKyQ3a4BCqz5wTtSOvm09fZpXsv
eH4+4z/ZL+sPXbIzS3c3pLka6VZVt30PTVPklqZgfPGN+lv5q1p6q3fthu8t
373K7d0VT0Fjrl0xwFHhzyjOcjmS+bFuzFRiegzjz3mNFZxnpTvEmczjTERP
u+mmqOz7Klz841TDOnnrCpNgXS0kn+TtkNsSkgRvkAEaDGiV0JUXvno8CV7r
goQ/M90X2bIBJMsQrnVhT+78eDVuZVdIvKlVb20uXVynqb77wKvPxwuUgBJz
9PnLlA8tYF9thjXRkxQaW3l+XSPbkc72cRrXsTDlkhsrIX2DIatdAvuCIWfY
o6lp0nlO6jHi0V6mUH6JW96XzIrtDw2Ka9ozUhnCLNNoX+LHXU+5NP525qkY
2CylzXyKxI5hCbB+NYOJxjBf2zGL8k5zsjo396i0GMaRmshnESYD6vGrqRw7
gZmEjPhRfngQBnAdGxX+SKwkKPfbpYGzV8TUjux/0S12gzeC7xQ7vgGYb7P7
AGT4kmxcovv13Qa0z+mmoMQ+r9RaOWGZOA7thsFvHqR9kmLflIEHvv0L84MR
K8OoCpvleEelfL+fwzsHV0s6c7lgQxoZWbTVkz9rK1tD3/hl1VAAVkZQ5Wlc
WYN0sY2tVFiGPErqMKuZ8F7OJ9qq+FuYi8dHqI5NexWK6oTBX7o3MGzmctTF
KjDBnlpJ+HXvLOsM/6DfYG27fv62n8YayZLZwLur7GuV+PR4rCoF/0qQrBtL
d60+jHMz7sMvwLQB5NN32+WXS3eEKyGkjpgcWLDXOweBmXuRDe64pLkTQatN
NvLmgn/lyAbRM12uo5Plp5UeJO78gtvZM1/nz3XuATc2M0GpiesRW8YYd7YA
jcgbihcDW7bKmyzGgvBC4L+5lBV25Sk2C0QV6rDAgjdTJQ7Um8TyLmIhqd1z
q7rkACj6I3qSD2PJxWJt4GkCvMAdjQrHI+mOr+mofaHOFMDcheF1lHOwWlwh
VvQscLT6fVa97kpkoSNaYAu2F2vUSWz/i5J8mTf17gzhmfQp3zy/2Hr3eeMV
7fEtAGwHPl7rZCj/xqKJzimVh8zufmqtBwZiJNke9GTmKNdGEnKynVeTJrTr
Oe8fpKVE4ySRWbIanNOHJzNxKeJkJH3zsgLg6daAohGt+I6zhX9bDeKI+UHy
if5baBBLDHlj0Iqg+BrAkz9/VVkBqg1C0WxpumcoEbMh9A7hAFjFWTrVv8zw
XjIa67eB8QLSQywnkW0qYKrtSFkOFI50hbr8a7eBWv9TRI+L7Dtxhi51oKPo
7xsm3oXCXoFc0RDA78/tfWojBr2gzIAkvaavKsQdB9k8VAXL/zCatQJ7/IeG
Nxd+Cm6RZq8EPts/q8FLwlED3hUfYZTA8/2SuUPX8PLr4VDiYuHa0dK3BTwE
0iyIhzXpi45U9P7VlU+Qq6uqQ/4bltNwOiePWsTcZ8OEzDlI7PaOKI7Q/c8j
jPlvxo6i/3XJOMRADL2tzG4EXq5+WAGjTk9sSDAxKQXNaY4R8dVAOI5HqenB
cwFYtYwD+nakacTnKOKU481v7qV46fBVPlXgSnl+tt07m5f/Sz/EFYUwZrMQ
SxzWmEUldsCQmPBQTrVT/WkHXGN6ojJoYP0p9TWS0EvR1ktGX0xT8haNzS4S
QY+kqYs3lM+r/uPAYoMSPSpP1IrkjkmLFRioj5PhD2MhYjkKi5ezZzv/EUzZ
CrN+un3UmLOa3zWy0m/EBGbImtSUmzsahBCIlXBMd0NRRuvp/Sf9/YtBi4Hp
OuWsNGJhIvoC956iSvJ9NsrG1HYCreJ+Qf0rH3rGPM0ZgPSSm/6eO9NG289u
Oig3vjhc7dr33Y1E99LsDXtGltgoUQ0x5mfaVsFvvPvi7OphOJoGPxtnDRCh
STAYhNKwNN8BVakKXQv6i++VjFj7MXyvWtmWKMcgawWCxBIBIagCxcZQJfOK
M+rq7fzBohDhkOJQyPH/ckrg0+9vDx9So7qKkSWpZMeOEok3aic35nvPNW/k
jRCrnn6B8VH4bCxltigwXLFIddMV9xetH0HgwsFH61ltcnGw9k29wDNzXZRe
nnPt+aX0uy34XJBDBQMRihCOmaaZHq1XR/pTLSHAWDqRFKH7dfaE2uE9oZhP
0Qb8DtQD/Km2eJPHDm8PuG9UB5dZ883XsBotXOuCryHNEQxz8gZcoHE5/cRM
AmiAbsJiL6eQlKDPh9PXJ8cJ6v1JjZV6LLpJmiA85v5XVxr35aGmQl2kaUS7
VRmxgnYb1WkIvJ8SYipsdq5rMJuNr45bRxSDv616aQPlEkPEuOw6/aGIKnTN
btjlPzevZcpdVycikTRelsbMiJucxirmC1GIlwHTh/BCpJN/IejECjU8vZl9
iMvvPslzGtSPtcashmon5AenZjLO8Ximdgnhzf6a1CWZh6o+OWvu3u9a5/Da
toYJMPFHX2Ya0EXnWTwOnd5Wrk0pWmRauROgpkqFeYTlpAAKwavMJJSnts8N
uGQbFJQJ/Xx+ZdjX1Q3fXbXP0r1BDF3znm2Xb/Q9D6gUtCjSKWA/VRUP6K3P
FQPH0twPwPu8ZxX+BQdGXalONM5gAqjJRg9+/Pohx6d69HcdSEios8LTt3Ab
A6XnR+dRfmwBq9RBNYMM5wBZHypFjxSP5hW0ySsYtY1AZPWp25Kw/+olbIAK
Nw0/wjYRzxoFMR8X+c88d0ENomCx3VR/YHZuDLl7X/xiIto0eVn2SYnstqvG
xm7GKc81w5AE+n1s5fT5vnXdEv5N7JJGro/JlohlIordtuwFuD1UeuTe19v5
ylBUeIM1r5Rdfm2w5kUomN+FROB53CTRga4ex4ucUAj2C6eNfULN1T1Re/+g
nC+vBCvUR6AFsGUW5VhIBk0ObWRSxI7NafGPr/SsrbSVxZv/+hjW1qdtive4
dyIjBdIqrI81uALv28R0Vf333sRaDBLRyXJRYRrX/7YH+B/Xn1icPhvFbdjO
t7cZr/T51DOQxuu3/HTkvk++J8M4C6fucwb90578okWX0V70y26jJcOwHWTz
b4Hsf6yOUsAfTQIwBJO/RG3lVTnwT4Xvs0IVtkdht18Ajw1hQLCuZSliGXXe
v9lPqChBeNwxeo1WwIMiklr9w+/gIkIEmbmJSx/dv2sm0P6Q8KMzQfLa5X0K
eBRCIupUNo5E58yx522W6BQi0lBrXtWzDgsGNiSkaJGB2EUMSYd/092+4hSm
t3zTvtJrQz5xuv2n7aYFxhOVlatecBUa54L8lLzsqAcWCoth4ajCQGwd/eOz
R0nvz5HcA9WjtGDqoD1hzNAAWQaBvUs/1UfOsxgPO8XdSU3eJyAvlqB9cMhT
Zseiw3r0tvfhS2/r4/tRHDPn7LgrDok/Nf5AR8DPu3kNh2OiEfU+4zAXNNy5
01DFXwUMKpePGwX8zmfCYPw9I8VJEQgLiog5NpUbtv7tSgkLG/R1IDQxaAyw
xYZAXF3hR6x/PUdoZTk1DGf0aSntMMABv9T9pcD9StbOGNpC5SPeVuBaf/Mn
VL1GzLA+2w/0ZXioiaXzE2ayM9O9JBtcZcDELqRlFYl6g1haVBWgJcOCi4cH
8tURwhWPHBNyRr/cLXAlLTtd0VXETMq+jejLxHfXEDYnVj4HrB+U9jmLhdB4
7WAl0XsQp7p4PgT5etLNqJNg/60EKUPigh1lpEYLQxAHbgibhm/f0siIfsMU
NR7B3VD3p6ZNdrLEfcfoXXx5xKu4JOJq2paR+wZAWMSZT+vaWWgQX27GI/kc
mnA+IJKjqeaTpoAYlv4qzF2oXU6MXPPgfsPIoHi3a+cSIMURschow21KiD/A
G6dXJsqvBClFkCVL/cDijBT1MFH6de7TaNCVuT7Hy8dHITpH4m1UYO7ezwiu
fXNDGgygNcYAO4dq83odQEgv0Pjvuv/PBrWzl8koPQDBkzzaNi3xyMYk1f/O
2qxLyYKANhSlcC0Wmwr/7rgc0VXUdymQdC2//x5pqBTAfTMv9fNB9AbS6lit
D+sibvwoabeex2BldrDHZGOazNiSAlpn3yn5fVO8iQ+V7Eztscpf9UFUOmrK
jAHLmFflJ60hgLYTTQ7dHpXZR56ZDwv45VThedUMrdmMJ+ViUT+mNYCUpYnQ
T2y9EzKT98K11XLixyZTwLxjw8WadsmbINMU5t6ngUuPgciDTOS9dOorMOaX
N/XYM+MwMuPXeDC3MsZxGcJ0FEHvBMF25eTJODfVy+vkzq3uvLTS7FP4NLUs
3wi4EXk/DSldVL0iwYZQEkzE1q0IMh0zhAE8+z7JhEHvmToB+biQlqPq/yJc
IkSmEe3/d/rBhCt5fO4tEUTEvLQBKf6G5XaddRFDR+/w+5nPDr/4JKEP0L6z
uh8jv2WvoK4PE+FDve6x3RwfXcJF+kT86TtzBlTRqGGgV3vDqKTLiHtBbcV0
xeSgPwLwclkJBBRnUlHLCZ9yRGDTCVND/nMcOBieJrA+NezxGguADr/Iq3ps
L+3CQvduk+d421KTJsoDLXj98ocDj1GzGsvywaw+1iX0tqD1EF/9OHOX2TVQ
qNQu4UiPO1mWTC1JO0Ln/TiQ00H71LbhXzlolOTx/+14yppJbmfiIoEKjDGx
5crXZHGbygkJvJVLTQbOp20LDTVIXHxu87eHveNCpsAO37GeP6Vxa29t5P+m
OQluTO7l4b8flyUitd/ZHtVnQ25yKrPnQZhrNQ6LRd5YaO8c+gnO+bHrkL1x
KjldVaRP/4Kz639WfOt8ODk3v+xUtKlGbtH5+/itiSxlHlyQDuJKEe6qGyMb
nBbs6NJqvFX0ry8/fEY8HL8tbKmjW/wDlwvWI2mQVVFd7VB7sk3N88f6v4hk
pzeZEG5Nu7HDtO1VxDyaGwEO0F88CYXRy7SeF+VwjKM+XWv9KZMgTGbMSJ/e
b46bfUl92CiWo3UW2RcIADu1/tEX0+qhjxXNoZD6CSSYaIrmP+W58xAA+mtP
TUOouBtgVtgk+FqWD4vI6NcyD56QAw7UFjOvN8pii4VoNqGgiyL9c9nW1iCm
lpbGVMXkhWIzDbf9EXm2O6cUjPaNCpg3Y9qBiUm/8/Fptpw7JQhiQOEki5DM
URIheVDOY9VoQi6hWbZtJgjosr0PPRbH6EQzVqKS1oMoK2o9rltmOX/zxX65
R9tjUCFiXjQBVwezsypMcq34W6SsxUDS20lXAE90UscQODcG9pUTk3N8S12e
3Mk6bTie90o1s7P3X2yPbICp/lUdyytD8i3Y7QGtuIiGuqPh+wHY6UnbJTGj
skfXlbpw7/lEQ/rZ1+qWeGboL49+7rWyOW1USZ1FZPFuXJccNLEbVa+B+46Q
kiglJuvDl3luIuIgVg+hJc15+1C1eFe/IcLntwHOTqFr2EyRr5YnM5flCmBt
Hpdk+p+ZLjbgVY2WW7wClccagaoSYC73SWZYuPyOFOOCIyavhWa2AAY0NmhK
ugM/SZe1AAp+glb46/NV5jmj+55OZy7648YWMsuiM1XeeHABoPmD2eWZ0MyU
JdZYMgPVK3pGDDLNrkGleYTmlAQntJxjoGf/GzE4ycyDgna6fGuhqR+hxATu
+LAETU8CTCoSEfsw8t2GEVlIgNdjkaXd0yDRab1WdU2a3C1icwy8aa0U3Bap
7S5BKzJ/BDhA4jJmUCk7FP5mwFLct7j7J+PXzSldIHa1ZUdCC0RBexXGMSvN
9HdMwhmt6VF8wEuhnvZLqpmOei6CXiVRN1qjLP/OdSqXLv4/tTJ7zJN0kIKM
oH5eECFvuI+cn3VQKytBAVxJXE1CFKxP7hoIpECg25FzE/vncZavh7dO0uXf
qD2o5sc2t91ZOPSkufTfGxfAp1DKBA+6hkQS5bcrbzQcgAUbidXPHhtwh44P
67udHU1FvXuOMUgcxwPffRF0rHU6wxOS0ke7H+qrvgytphG7bWEBAm6ksXB7
Lg6vazEojljzMyLoX4FoR3grpNmJToesPLGfT4ZdKo8iHZTdQy91PGoUIGBp
PadEgINLltN3u4hO3PZrSNbcuyiGQbvrnuTDEOBBG00/Y5kn4youEzRALey5
pUpODl+g71A6ak8jJq/GjezGxXZ/JOgUnYJQGflrjGnIEMPkFAiZ9n7APi9o
raNjP4w3zYnkk4Bpfvkr7suo+uFcRc2etig64Kx3M3q2dT21vxrOKDJqbLJT
N2pXHWsacSIYULTXJKayd2uiflzLC+DMjfgZCtiBV0e2r3QL+BEs8a0m3UY5
HaCS6R6BeX9/zuw6NQUh584HgXp65FRmIV0owHdXwd/XnOADkTBmyDlkoL3a
XbbSO3xrQ3BBTMhy78hNXpa2dOnasbz8m5oXb6K3NLO3b4ruomJ+OMnGGcv+
//zbqFRwq6re3zsk34ZRntSPQIOMQsrgqCyeW42KeAAT+Ywda2ARiMHmz3cT
wKH6dr/IxEvo22bj8mQO7itULkkOiWgdCxKEOFpSdcY8nUjlQ+XABl6Shu37
2JlqKNm30AjBE7gu/Z/k3e1+B6sOEDgafNyTz24hBFDkdc+11VEm7xZM8jVc
cHYKrj+tfbF1o6epK0ekBxw5WMFTG8TT/4wRi2J0PAnSxQkMfdOQkL4LcD3P
i6J9Ruqz2L378siYVJ9Bi1nSyEL26K2oMJ2xSBNBGRvzR4KuUkOqbqChdFc5
iOGkQRA0nA4nbUXSK4kf1kjzJJihCTBVHX5JI0PULp39r5tQsQuKdfPMXZvd
tv3/7mEQM8tnHHIWBg6sKgLOFvDN+SGIn68hKpSKyPJpZZS9cOJ/HGX4vjJ5
cV5hn/BbGR0V70wc4p5NdQHUapsHqeq9il7aFyyD4I2HfgJCx8fzp9mtNjLR
SGWSXqnOuVQS0yoKXL4Ps2WLAQJH7qz1WVyyAo1Y9Z3271xv7b+z7PfVrxde
WsyWJmkeSbAzFYbcm8JnDM5Yoqp298WZyKbc1lg/8v/wxzs5NLKdviR4xbpY
OieGqeCfUpRrSoMPShviddnhERxRwtVJnsjxyQqcAHm94fmnfbvubE+GAcWU
VZZlZa9lEmiME6J2f8FQSCd3le+MWYWE1GT4uuYwBGtC5Qpt+8KOKVPPQ17D
nXvGAqOQ0qyyNrOhxWeBVSiNZRG14ESo8mXTg7IbNMkGxfRasBAhIszvbruw
4mROFLeBO/LD0fITDFw+jecJ0ucdSBTnjbqmtqiq5LiFsnO8+iC5qWR1G658
zMcPM5aRGH/R79hN2aINw1y71gF8oO3AWTJAwCm6PH2ryZq5F/WWo2EPJ67u
WkgqOAvEZCywnchu2yNjCV17IS0ZRXjNOzaLIl0fE5uH9cWOVcq+WfWoAtMP
jrpXxh0pAxwDr72pR4h7CTUrOkSb4y3d+PP2zwmoWWKmi8ChtzGO1iMW0tkR
G9fGe7FqN/6S0JHdvAXuSf/BTnzKtZus7XRNSHXuFnpoDUtIIyK/aGimP+od
/9zFYsYi/O00IOoxD/DRFMIq3y53sbadYGQNnE1qW+sIk6Rmwxj+9sMueNWF
HSGfxugHmd75fSLezRxcabx4XlLNSYDLk9efReDdcMnXLGT8T+3MUbyhnXMh
qIkGK2d71l9JnTEW3GTb/7y/plavpeaWSthBCPuQGQcpYCnV7cYFDNcGTMJO
GjdH/EqhLRIWGDLcbBz9Ay7FWZLrrscTx472s5hI7kxxBWNVBFysvPowPL4L
R7UHcALQzTYKL3NBMYjtjXENI9MOmwJ1uZeN90P0Bi23iBFTdFRdtPAkWgBE
w8Cc/4KvEpxftq3Pa2ctlDuQSv3orKjsuv94IDPusQxSTYJGu/fjjtV498M9
xCxsyH63jfO8cYIuwQUbZJ7ogwJqK5/3SD3mFp5xsTUR1fywA42nmldpX4KV
dZ0F55RW0k3QR27/ujHNepJ4RMozrRm16Sytg2Oq/iSXioyefudjaZ/BIZXD
uu5EuDBjxOpY1bEmVzl6XKxpVkAQd1tushBxexU5BkUj2vC6CykRA3F6Z6Qm
yommflkc3gsAeFG2ycHZO61L9CDn1+XmZ8Ze7FGnD8vX5anJlX8abkBy8Pbn
mBchxAQJuTatAN6XdNsb17jw1blB5e+MUVs8/4o1weJK88xOnehw+X3zYToW
33XhKXH1UX2dSNUAiNkf2eEsWN0+10AzM4DPRWdP59iGNNQNVWG00JpK2XoD
4RNkjMj2W2Ew9H2mXA9AvyI68VoQo0FtSqZUMUQfguN+MkdpziWy+AyEBTsU
/nAL8IrrJ4z6W5+389aA7RGstTNFPlNf0nzPHS2UIZKg7yGrx+0H6KcVHmOE
5doq5d2B+BKolVREOAFE4fmgk+f/j/r+J1A7kIkBltMZ+kyEpVlI2LVVpj67
A6VBr5OQ2bcTwN2lFiA6pCnNNfEXfiVu+3bzxIjMhD37UauwXhl5D1dH7gop
H6DwTADr3GWthz+hk3yqL8PeemKLE0wEMO6Flv4oSXuMzU+iQG2SLNAZUQCh
M/E57wWCIA4Q/MZ3b23nhep+OGgURMgRF6VPhbQXXxb9K2ehzlR6em91DTet
nXzI+rtPbaWj3+z1j22maoKxyCv3MTQJfrc3NkBYx/Mvebsfk30KdO4Hgv35
ACJC1oWyOFJV7bC8TNUBkMYsR0Ze46E6lK+MB85Nw8TPzdfw/J/ZHf4jmMM9
Vjnh2pkLqCfJmBkNNasXvvj84ea0p2GJOwdloyqLolEmUEPNv0YCqvuZQQoC
TDpH5E7MOpqx0F+daVN/VhLfJMfI/wilO6vmHGVmGZU8sSV6pS7gZ1t/Nx+1
2ucxmBCRzqa8XE5Zw05SVAsdzltzaOmFLKJFurSaXt0guaVymGANNaIlbQ3I
Cl6ptWnz74dYbk54th44AlsGNR6GNcZN9aa+ruAj8JR+VjS0hrJBNGRZp4mV
bU+EUJl69RTgs1qRAav5FjvhDqzX31lVjnuGRsd7layO/9tUwL2vzDG9md2I
ebmFOJiDNNK0L3MSJvliVAeoYHwyyXVnsQhGQ3tMx0kN4Svl3k29n3FRwIyN
gC45gevTsllD/8C+o7DG6+oMbo3qefDlBoP8yOvBqyAHmHx5Nf9A4jGzry6B
GfZ2PI3kX0vW0ZD/Te4QXsaIsVN2ZJahgFUyBnaTjjGV2FwQhS+xTClDlXAA
m3Q7EfYL6W+Wb3+hb1qObzdCxEX1mZrPF4+UmWTesk654BXQtGU90myDDZ1A
2q0jJE87yxP/NHLKNIUJhXNRTcjwQXrrBOEMWOh03fxWGiENjVmvbR+gtixO
S7YeuM9q6JwO0zzjd0b+vpKi+SjEAi0HRdJYyApmBYlPLmYtiBl3JFTId48i
5cuiQRm3RYyVAmXO8Ox0i3rRytHkWn+y0EXMGfBfwcc4I/s3vk0iy06O9Ocf
ReEy3iZTZnLpkkKgrEcbTlKZLhf+TMK5XPOlHuReiLdrt1Ktp8ej9AdIVKRr
Ie/3q3b4BFERunmmOy5pqEaM31M4e1pT06FOjgsidZcX+TwHEybcbTEH+2bj
P7FQlbsUT2aJFYTTJwd1/+rd8fQ+ujNB/t6h21V4WObLqztqikgLQrVqFt2N
txTSJlX+LPFuirY8Q2Utw2JZH4sJtaRJTKKcJc4zRKPih1j9AwUOcw50Dseo
FbruwCTcK9ZuLgO63f264WED57onMlidmr+7bynmLgpIvnb/MOd5Y50NBw7f
U0BKMteqNKUf9Ctvq5KeNJAzSSESp0hfsTjK2FOz/33i14PEk1K2OO3Zc6uL
hfNPY8PjolIr0vyb/ZuLp9UILWKwmr6YN5+TgDJ32HkhKmbie3yjF+yAPU6C
nn6EbyeKX8Q39PzHhMjnkl1jk+mQvwmndLMX5smKuXoZ6+og7VaG6ybbqBub
1p28YyRNsULA528A9oJMmp9nKEQ9h8RaO6hJFdBDdokZ+8vx+xAd6LY1d9ZV
W5VY2cMwn2dyBUf4OHUlYpzYCOxVJ8JFdmZpuiWwaMD+it4QWsO9TPg7a6eB
U73tvtKVfsQL9cWtfJ/03PZY54PJDlRE5PZ3YqAAATHy6kr9LnLAwbCERtWx
nw4QBku/D6KS21kIegGIFFH1ZFerBZHKNpSCDQNshACxw4HWtVaYKuhx86ip
aHioX86ngrAGUZAT4MKuSR+gKhkyF3q8M0o8wEDanLSKOW9TXzn6WS5Orak6
l+UtRxco1L0doXujdbZPuqbQKXsQhdSkME2W9UOibHKgUJ4m2n21x/10RXZX
FRy5VDVMpf3mZxFZy7MNnc1Y0DJY4PJ3rgMRvCNX0V06bwftLuwNAFgwuyD0
C3j3f9SQEwAAouYADbwUjIWTmx48oo6Q18D0UNnFOdHWGhzz1G0oJBQWhdXK
FHTGX960n1D5wIZ4s74P8xfr6tSBHMrrWPT6baVUn59rxHl0AHt9co53k6YI
6eB5GjQeYBZhWfXQ2iASccrc8UHOelzTuVKv1gBrDuiQ3wrxELA+ljiv0byK
Ssw6LLVVBOK2AZaFTFipaqO26Ua7FXzgfTnhCLAeGSUGf3AnD/wPuHyijzD8
xzDR1uS7zGyQ+/YNnXWY9Bjh/gDknucjyYLwwE59OPAgm6FWnVvesCqWiS7P
TInd4DDbyDuvkiBgLNV+kYclpUXyjhawGEd8oGRqcAW08jQaZjmmPFNKspta
wlgdmATYhyYuv25+E0z2Sv4Z2fJpJHJl+0fS14OoEvpXg/2kWu+ckxQM80Uf
r3xbMtIGAzIDsp6KslIsm+UVzUDB3gZd81D0wrpH84VZI6KUHWhScjtsXCkN
Pf/u2ORhR4CC60Vg6iRhxyPJ1pFHVLGOUSbuCGx3xnDhieCcscbszZwwvXFi
QlmiaC/TeGNww5wobkWUWRZ0OHU6vGQY9oIblvqBh/Wyzm0hQhoo2TNNnv/y
7KrAyvPwafKeyCoIRh9k1AIWAcormUalxzY4ow8KnJzXNZmoheQupOFmTXbj
XPo538UJsV1yDTRJ3DD6QZUBCyCznLwOSMkpbCrtOho1pb1mEOn8vgL+C7No
u1B+g00xyO1EgGEKbBxFwP9QTs6tGJqCxHaI2/GBzDZsFk7Cnh9DmQ7WRvaX
SsWz149X23wOiMVS75RIQmS1iVolDIHDVnCbkU3OEuRwo9QM59X6czTPLZLN
88Bi2pdFE/M6c7dWL2MrDKBWpM/3bRVpF8wd8YsJvnxtmk6F4U+okOs2lpka
4qp2bmbIurIJxkswbla31k5/LN7eS8ggquCDjoUkDCfNN34HwWK6gzHjRZp/
8ArC+BKjZgQvzBRsqNnM2DJGyXw1nf+jV142H7SoJmTUnPZLix6pRzlmBqL7
C6mzqil6K+7wcivAizJIHv4WtsIv07Z4hIfqb/0bO42QM1kPdDMrh9di/wYK
tyg8FyQRKhBYlMfibcggJnCgmIiYoQfHdV7KEX+jCz/l6bpSEIqknXHIwb6j
h5aIVRbXuZDMOGMypiqvYJzYRq7jgEkoLDdNl6nnP4S2dEL+voLtJsD9rg3+
fh8lwCMLPK8EyBG0p2N/4dzbTQ0wpiuGgiIJzVzpekDOqvFI8sifVy5pM+WX
3XXAqcZ841D4q3L2pgequaLyvGz08M5xBNtXkKO85+G3PWexUdINPCqncpMA
8rPiP0pYZaj6WJ8EyquOZwFjZyXuV/kneHsRqQyd49/EisGdkgrebN8m/HyA
it8pVrSn+eOmaKXxEhjcpUR6HCu+iY+/YpCLIyR4xDsbTP2Nti0UvBH5BHCS
FJzhoqCh6Lc7d+Dlz4qffLvj1RHuBIoy9SHkxNuLqH5pitde81VnVtnVHw3d
O2yyaScOUxBCneNVZKIl8YEsl5Mt39bHNoGMUgICYSQCsdg7IuFPs87tu735
Rsxtux1kVP7hvlFaAVdivxTKx6n1jhhrBFXrnm7FUj/bxOOI1wcQERBj7yNz
yjHewRu6Rdk7gGbyd0hBvr0hSoZW4z6rVGQUXB/7yZC9+5l9zkvI3demlrnl
kCw2p/bglbpntVTbgBhcTq/cawkzUrztZuo9q77EOrJ/L7KBN9GZv/hSAIOn
bGLT/mqDKHs/5pvvH/v0G13d+JcYZnQ9dgCA9QgGmSZKF+YKmGh2uWZTXjVZ
ZO32KRZULSmOa10Y73KZQk7iFC/qiW6yyBzLrscC1x3Gotaj/W38+J6uvgte
1e+A6kgZteiY5F4BGW//Ht4XmpGV1c9gpKwuJuGt3C+kXsOpWsAbvQI4ADJS
75s9NBC3HyhC3p4xi534WkK7VgN1OxQZfVe3qA6bLqQrd672ltB+bFrbxgCQ
NWLjBRk9x/Aqh489aNco8emzegboLTjh0iEcnQjGJmZssaZp5HFt2PEXY638
S5WSKpmdrCQwkfWymuMADWDvRRBK7PZ4yFgit2kh9hrLWcjut1PGgwC1cTyn
K0ntkXSNk8tyzizziGkjoupAku8+61Oqe9BHZXNy4yHpiOBaqTrDMauuXP7p
whdvOEZd9iTXRhekuAIOu6P1TPrRXEKenAAaqBZ4dA/rV53XFOFEvy4LNt4g
j117ASy3W4D5ntpP6WsRQTSJIQ1Wwdm1eMJuIfkOZSynx5tR+y2HmcPAXPjW
lZi5X52RSN01CoqMp6+SO6N+NeLZzxYdBh+o2F8oiJb3CPw+kG4q5SjaO5vH
eDk8oNKxUbzML6gKGyZRzlCUq4K4dACATjFBVmvkyl46/lVAPZRQy8M85To0
Ux772nYAA2yx/QnuF3/5VFDqPn5QGx45EY1YbGcWIxiNDVG0gmKnbebhvq1b
hmCndi0KYWCeV8xwReQ3cEfgOvxI8dHKUUb5FM0JscPun9TgnTu9qWML+SCH
4TdVw2z0Vcj7+tfWQwJV87jQixxxtT/KRfJO6FDXQfwSuCLMRJ3ExDrfNs1u
3lxm2+DmnOTJEQYNhJ2A9ElaQsH1yqeG/K35kKt3nWf5Z0XDRzdHJtgffngu
MsXpjmf2IbHSutsYlWJoNDvmnNvQ3EoYaTSrmqLw4Yi20ItGlg445XnHAQ6x
xXbqQVjnAAoN2R9kKnIoCfGTxAiY3s7c+oIABgNm28ZGZA4GWfWlPXDvXhKb
GHRnoBnjScyfkE4OwQZXwLdnZw1Ac1W0spE4rIz0Yg98ZAnMFaRdVsYlHslv
xmZ8KqgGSYXz618JIzEs0i8+pJEkGTVKW+SZjhYYw8fqefcqBPv7OrbgHkYI
NdhIbMQ5pMNq3AZ3uGDHsEaQHbvaTKO1kN3Z1VvKsdWCcZbXo9jpifk5C2l1
KKtTxS+jF8jnVGZtKAYS5jX8QKkk993qZ8DTON0SF3nP5kgpEgjEmpcEl3nU
Wdb5gbrYME2ISNZN6VtyTtgBZb9lTJ7kXYPoSK20RYr/ZlfOlfNF2Wc06hx8
+zTEa7ezyYIKAO/eAr1PwrlEL9YgWZw2ye+8kMWDmfB6LcjjGV4tcQetYQx2
t5GikU7UFOH9v0Tv0PQ3x5HbxcncLaWkI91jDIC81i0ZOJC5eeDdZYdcn6J/
e5TpEuOPb2aoWvVB/ELdVl98YCb5GvsYaJeLMBaGKuCOnYEEdP5jYVaYU36c
LjhtCoZzBIodV+JwAY9mNmc41GF6hX2qsxdgMaGgPaay2DQH/GE/aG1voNnY
C5rjJ4wUCa67DX7zCOHFdzfLUGMEWD9A02Gxv+G+nb1xK49xPmdAUoOENJrf
KYyvg7u4Pl+ECRhztXBha32WL8UxIRFttl8KCv0QiMouHmvM4NeRvC+esppk
9+QXgO09n+Rp8TEHMensOGcHXYJdQd6V1mafKbWYNcA1kDv6Ym2pEMGE5C9g
75DlNt88whWlc0v9HP7WbUKlNCg9YVOSK86JDxyz4aqc0r/ouUeM3HZrPtBH
WzhxdmAe7uWOSkU+wbOgpYEWOOiYLaBEzIOuVOoGcDR7eE6WhpCsLsmR1JGm
ZDy4sYuvdTKqtaCW5yxW57R9d4HxavvJ36JMJawQVKRNweIXLHBxaon8143r
em3eqDNx4GCR/98QfJtTRXhRB3KGCLxSFc8Oq2k96Znk8OADV4RqjhwF3E1d
pCji07l+nrTIFkWkwn4nwFeZ2+McZybcT1Pa6/OLG7F58cfG453xIGRCsFEl
NWMY/Psu4Y43PnbOcPyKsrpE5e0IgVwhNn9iuzTimzhZcVKZsGWYcZWm6p3K
D9EqrG51YuvnsnNX1XdLh0OskJCErVKxCBPFwdLkLu1BPp52a4X8NsJkaoHo
u6jRtwOMsk+BVx0IWhTNYyXvdtefnpirJrNB7N6kbxZ6jmoldyGMyzWSsCKL
p5p/vV+osaIGEw9+8Z6KsnbV399dQrry8SRpyVSiO2Zrk3LvOivegYGco/Eg
iiNwPUKVzp+lNIQBK3UcCj7PvZLrYyo9XcssZPtYS919bESWGK4p+1f3PN+7
rML2vFwAKj4RYkhY9DSaCRiuaATzq3W47UpyDYWgTTzKdZ+u2Es2VKnxvaKV
0H08fcvxrdcXfNrJB+8vkVkietKdxPOmNvIPxmc65ZnTYIDER4A7ZJMcrviR
jWqnHVuvCmkCM0j8wVBvapfLUH1ojSLJLELNxgcuY/37yIoYO89KKyMP1siZ
50xROBXd8Fm8xUCsxZQngUuESk+uNorKSecMJ58pPGZ+9wvMiU9TDWBYh8Sm
MVKCpr2AWzJanIGcrCFWMSbnOal7OOMt4KtSSZPGUE5HaqI/jlbUTN9srqPC
omah+bsU9YM7HSYpT3tIhAgtuAssFbQd1UQnax2QkrvrJMLckGt/QvsSxwYM
5RzoF4sjBEK5Wha/zt4FousMR7fwK9sHkcRDq5wR8vnNEp9v1IS4W8y9SOPq
W2/Ag3jkRA/GVoANi6SkiaPnM1hkZmPtPZtCxfnaNZE1NfioQH0+Y8byExgw
E6zT2AIp01OGLj3EyYbGHi710CnzXokt1ES6/NEIpp912BMriuz0cGLi+Bud
Bzs5WfIq7M1gigFEvvfa8p4PqYI/zh2O+Jy9PrgDLR9q8/l0jpzCxkBX97gi
9DyM7hFcrWd4h/DhztcaLc+mvoCWe6WG6SWxCm+Jcm1jTN3FrXxqTcHdZU18
Qu40+1Yke4Dge2DwkHvn1ESbyj8KpRsm0qJrkXvgLZx4yWbU4LNG8k2dlVj+
Uts8QEcD+RKAXF1yCeJZe4hMevQ9yaD7r+jyaEXz2ny6ZQiK0RkiEwn3cmTx
Kb8EE+2utUhF9cUEIk9uqeW6q/eKADu8q284laZiXhGoMgLF3Ibakl23HxmD
PUejKnKmx2vXY4tphNuInsUTSczXV3CTHGwjpcZcbaiAosy+kGuFGxIX5L6z
NaiIn2a7FxjV7VaTFezsuh5fw84hMSCSWvUPJmnAOP96HN2PglZk0PbD53Bo
znWNqcj5K460YFbc/6DjGXIgNdQ7YacfBP+uLp/8xjXkhWncwN5C5axDi5fY
syvqxjMR0On1ITDK8JFOQC9l+/fpP+yLjeDpfBdba0G7WJKz6tjFugIaYfbZ
9Ky+hxqK1Eh9wYXeSFQrFks23dzpB7BHp1tq7w49+LlFOsG20NGTtHGXwSLP
NbHLlbTulRFHjfb2gdd64aqy1lhBaTA4GcHh/Q4s80XZCQ8GBFDit6Hn7Lap
ytx/ner0IBSDEIyTKDqm1+SHaFCYjxcuVAdHWUrZplVAErrkXas5szTfPiC8
MJDB5UhK3j8WZN4wphekCWYyLVSbvWskfXMw64N1jhiQO5I9yvvtM72imZxH
VSfxiL+CV1d+31PkWY3/Emhy+DUZ1o8NP3WSopSxVGfbCAQvJ1VoeTzGzxRY
tkptTrRQog4WINQ8QMxImE1eJccs6mkny7hq5Lw69SqtBnbaipfdH6zAHbMx
/tTGmxK9/dBFRDmOWTRZLQV3OlCRZlOdFRYJfQ36BzoEj3K3Lls3DBm5qD2N
iGkqIaS5o/V3m2QjZLu8CgIL54giPC6rcISOxSA8xED7+pAfL/naNLYP86+R
nZlA0xYcE8yVCoWYpM2aU8bw2cQIuo1jKuYsOcSOhV4l8kztFq3nhwkR0sTI
SNK1LsSGaC47BWW2TxAilxyuLlWsgtYAHm7b08n7ALqQAMckDabmfx4VLn4Y
VfxGofs+Ia9Rv7UBUXzKpA1F/7YmPa7QXApFhRHADx97foZRN3kC+rWOqzfy
yde90GKrIdJTZrM/6qAsVvgeAj4C4A4w2hFGDKaIDdr2kVaUi+Vhp8a1O+YY
owaXCHR3ahqGZvPY4cxtkdxOnu2PDE5E++v1Xg/H3lXyHhpYXAdxapDY81Ep
+J9qTLhvnmNsPtiMtn6MZPCuvTVM4uE8ND+yYlZlXEYGb/wLFitpEKVUes8h
uAq527/pEPbSpwMkOrLIa7woryXVPXoDVns2HkHm22Sje2jtZ5jhOq6SoUfA
ietcFDF2JJwUEBgxx7yu/8B1RNCVE1yVLHIjbiuQ3IN44TkFveiYi9780ZCA
qSFz5WzMWOK9sB2mpLJ+XJAagyhjzzfTMC1r7VUFZEnmjnaPlJWUE+XbJc1Q
cU2IWRNZciG+07/IobXLSt/pBeqehYjUCENbaw2LmJG6gSnyZsGqgvjV97oN
0AlVkzAi5pd2TuT06B9yzkM33NoFCu0JkgZlLvqGPdylns35u8iimyrTC64U
yI0sLgF1djBWpRjTq6xXbMMrrl2mDFxR3c77V2HTJcD4OnOAC/4ZbwhLEZSH
MiCr6OGra+Bvucs8XFoi/WKDpf6YsiHeSlFhc90aMLzFRjtr0dzmHfEiLI3D
YlxCZP2lPboIxDgvau9WIw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EqdW+P+2Ur/+7GIdbys4p0hb0gojvnEkP05SXWK1uakCAc2wfWheLJjuD9ddmd/kDeEmp0uVDqj4mJ1A3aX1pSV1AYFgxr6I1Y1759ObhNTnuMJn5RO7vkse/4/paTVRNDZ8XIKeY5M9KLvKQz8RdbhKqh2tjAnuiXqFMHoBkBvXFUNyArdo8NRz7+bCzi2miiE5j66mwNmZIWLdWWcBSwfi9afKlbHEJNtCMUynX1UmG1QRwxFkIGhI8JyNcydpKKRMFHLelRsc/tyJVzsFprEdgXCaUbOtlvDuIQ48s24l5U8NCli4mzsz1hRU+i/xTVaytmLQXlj+GZtfJVNNXDD0tmjU12JbZo5VdtHLMUq20/JyhiSV/3JXASLzYKEGInz9L6/3LQukD4BrVPjkuuZ5IqFg91dynoOhBkBfPJM0YvZk+ffUDI2dGFHun+6WTZlEDUJeOFhoezFSBXGtXPnzbYcOW6X8T8OwppMWf1+dWu02WswgYiwn5ff7MpuuB6eZ6Xh6c1tq4qm349bfVOFA23MmuK9BrsShHsyzCjFt4VeUmEEvOB3Xsfd5EmQr2OKJX4tc6LKRXYgndTdXapsTccFncX38KEs5cTf0xWy53zJVe9/Wg5f7xSVKav+oMLWoDdP2xFHtpOuQfMm0XiMiEhnywxYkBcKGpRyGQVum2eLRmvMRTJsherlPWuHR/b25/6fUi0wHSqRnzGUEqS1bkw+xpY+NGBJSi7POIlQ+CSmn9WS/r17kjFnRi3ihE7ZBmZkrlCW4gk5/eoMfW34"
`endif