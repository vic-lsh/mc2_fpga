// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LvYLRvPahRMJiYujDXr1EHfdlEfYfdfWG/UI4QGJT6eh25rR3oDHQV2cDtOM
p6eB/J8nqXO/UDbQ4fNYcz2JqXihLBr/k6QqVT3xm4J5rKKkW+g5BwL/yIQk
098CXFVfe1iLclrWlu0RH8VsUlKnbJBpai7EHYzpNJe9geDDtdJ66tjKz5YR
5iTZPuSZKjJCRRExQKa5uao+TipHUPaz/whov3TaG+oHLJLB8aIM2K74FzXi
guexgyff8Nz26+4rOQ77AslHtOeOPbMq7B82geGj3BPJX6b4P1EBTddAjsmD
7HOZKaTb6mvEEuWBVSq09vWBkFiIAJXjRAjQ9khaLg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XzpKuxoNLNsxUSjfhVcLq7MO/u/0/oA+nOCDSR6YzZeKj2krRevjPcUPOchC
e+DanDVEby1Bk/Mvp4knEMh1KW5xVMPLCx4Mad1KM8yTj27FG8o51Ko/HlTM
Engo69Ru0bkKG84UhnCrsoQpDhdgFfL7jdDevTwFL6tvDshekLH2Rey1OWSG
DM2PjZZRwNguIsqcSWRFQdgx9J3zL10kdVglMUTJMQjGFGmw/cvm/mdJezod
LYwQW5zT3pkX7/UhxwZgb0OTFzbOne8blhAMM+fuGCMW0kqSvtTX7DFK1VpZ
oNIEpgOs9K8NVfbwPGqe7jqlg+hIHBf/VgwCIvDjNA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c42Y7CU/BOXuLCSL2aHkRK77r4P7vDBTOS9nDJHJC+Zm1+tfQSrVM1OWqvFb
8nbOOyLTn3+eU+tbyUQP6FWgwndMf/EdET1w3RE93yxSmHZYALj/mCXOMuMb
0NEsQhRCDxkrgPfW866xm4UoiNJeo759JEjvZeE5S/Nrf9IeFbrTXZqBv4fY
95G7hP+CG080OMn14X/sxAum1nDcM80cQQ0FJOyfEgaMtbzPutJdAKWb2gmg
MTrh4JcxM+zFAgYO8W5WcEkWSdUDnHgWeGjTf9qS2Z5+wOrz/667hrbqwjvR
KRjyUCqh3YnLvYnz2biIZ/69HSTKNZJ+p3+30aecXA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qS5cLN+V/K1kbcQ/1HP1cBwSv8/CMYY//tYVf+HrHPRuPcnB4o9Swf3wyMrr
My608TndWbK6Y/i0EIj+OoUKZa8mkczT2uQlGYYlyTXS2fXjEhHEACsJw248
jy8eGfR34EVELHEXL3L+yt7KYmQ5abXYsRorkb5VToqI/tD+KqgbmODegT5X
9zPF7Vf9Zw1xuvJh3J/dbHLLKMQWdPROP9BXMHOMi2WEtpt/6KQJczPo6qAy
RdJF7xF1onQnKipJO8CPxboVPKtTfzwhj6q1AoTSdWDIv+J+JEmUvMyXaaDl
48FTPnU4KtVeZ/e2PxRb1M62veVYnqfj/l40EWpclQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qIIF1MUqE3MbTznlXOFNB0T3kG5PGQxyg53Vpg3sgRQcgr8U78Yg4Avblk6v
7BKthZ24rqDA3zwomP+Ja552X47cbEj/ug7nodVheEdBbm/zsakkllBO2RUV
h6aj9u7hwIKCjo2uGIRsPD5tNzjWFMdA2qhAQmQ0YHeBKIsQqAw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Fmx+gM7WjecCsbsW0QGw5cYlc6d0BdCFPtCydbl8btVDRLPiELdS40lwFYA5
hxYpVFkW50RA72so3xBHm0uToh2Mhi7aa6qGYadKDGpvvv6xi0+er8mOumzV
IP+azqzeF3pWR64lrJ9MChMwLz1m5Qkr1JST7bYN+xsoFx2qBwcajY8sRNUU
bQR/7q8p6LXcJNBKd4SupJ98OJxb+cYMttDARtjZr+ELXof7l6Gsi7/iZl7z
JggQxerEqhoa3p+I6ROVkocfp7J3M+LYwu0SRsnSdZRlLooLQ1dXDPVYS5eY
xWR7/LsO0cPSf1EJ4B1z6SYEsqU3VDwh7i4S+MJj58GciTgXNXeTzOlUYLoy
GyBn/cs/x8EPMY/nEVOfEzPiWugm8/grbh40/f2DyrFj4Uj8OGIBeiQSbnvJ
PlG/r5LSkX0TqrUNcT9aK5cBfiafeMovAASW8ZP85kZ7NBznGE25wvjne9Es
ENBuR/U5H4xzVHBfBbY9ncf7OWFpOe3Y


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XNNvpSydjSzCdhJqlmZJJCpyNB3Qx2IhWo+zXgqttHZoGbMs+zyBWlnpvNJM
hmBkK/uhpCC9B69/AAE6aslEO891GKicIXchNtuiVJ8kJyNr5mLUbaqL8w0Y
VmzrdnazFhmqrjQbjxU5XqVV4Ww85hGTQooXsVmFZRjssMI2oy8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
S8GMjeyUXzz4bjfY8VDSQNGGs4ZUbHyG8ILyfd8EjoegHNCPO590irGsm52k
Uu+U3RYLlK0kwXVsgDR9+NzxszAUSgJgMHtl9UVOuzdSVvc0Pfcp184js655
YHO+PhI08bFrAzBBLeSQq1uOhm5FDOdm/y9Z48bwNA4k4pmGIyY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10352)
`pragma protect data_block
pv8tBJpGCWlpmwawDXI3ijG9zA1+xWxA4+MWLQE/NwTq44nGk9cio9ZoFHQQ
NGE6ppMDzs83oF2zHULcImKrQwAyuwOby6Qg8+ul7Qdxm2LeCRS3e1zZFJTV
whFOxeEGM2VJOFtofGkApuPFPcGVhZjXhEE9qmckmA/nOBb6pZwvXPJqgCw1
XCQWmYfeN+wzyG/cL5Op+qJ5UHnE0GuEt4s8bc/m+H7+teefuRdGzOWNwPdD
vBXG8+mJSNhkOFjuPVZrkXbBpW7NWSB2eACNdsRCGlRz6oQ517L6kju/g9fr
k7lqJzKy/XSKz/RaBdTuqh+NOF6simV035gxeIgb/Ve//Z63WFqtmEVfBjiq
7X4Y4QLBVW1iKjOu0jlvcvuJlInBfGdY8lGaC30gyA9knYDA+1QQgrmY5Qvr
reyir0fgQXjsQppof6Baup2LSclfzBqFM8xKEza9XDdIecEb7sMkIXWca55G
wrDLGvrjFzBzz+JBxx0Ofzt/zCoGAp9pAoekakNQC6cxzv4/EsmsEoti0PUB
FphA7Sz6uKeXXOoACfHOH4VW92X/VVuLoi9XHie3fi0ojbTxQ62c07femTzB
KDODjxP/F/wT6TUNPfgASvmQFip1BIohIpYW7nVJPvM6+XWVCEvJFyn9DhYC
+J13vNVEmE5abVYuv02gBaUHhEH1fUL3f7cLhbiVFsVRR1Cm7WPckZSS7uA4
1h6jmcGloE1/OeNyeoUpaObHr0whWPJ5aJeefhFPMhAPraN1XTNlXkcumP0r
8JMM4GREHECcYWI5ZodWYREIHa4/Al0V5rNsLOdvmE23pZx2oawL8v3bdAV2
1/xamgyOvmZWkEFJGGjHFShAdFxpKZSoNbd7lcAvyy3ib0iPY4698JVE4l6b
phyEUxoiwXFsvouvHL7TyorF17cFSgqBA4v9G+OlUVtV5CXQRbi2w7xfjrN4
sCTHQ0Tdv+JolcGbyVj5pp1QfUBbRJinW2YJA/C035YpiiazXX2L8Ax7upnx
vVUAV/50y4+SbHhBVMzM5zfGHCkU5YNORybf20HIawK+mivuxZjL+WZ43hpA
HrQwUZkvcjzYX6hpwrYh1kGTm3idlyZg9gifdS8Za4eXpkVqPhhwlwWHbfsP
YcgnGC0+umpo8xyHTCJMBxb/c1k4iZ9BZ95iIYuDBEP/EoLmwd49htSy3oZL
DPK6HCOhguuh1cxuaPIRDvNHvj+2B4nh7ReiRGE2LeB/dznDp3ojuPHe3xLs
SeWqCSnXjvXe6vX9U22FGELnjPCpYAQWSEjw5aXSyYgdbXshFexAY+BwHio1
eu1PYuePNdFmp7bA212yJOwcVAA6PCoPHyAaaUEIRhjiNnNHrIWEZ8Dd+LOf
NTsmbkqerMmtdmbP7DVM8u79qEpY7Ttw9dkOs0NI1zVDXVbZOlwSXUL6jBg2
oMyhBNiJC7SsvvFf9R8UZ8CVOuBCpd7jMPFCT+iD2bZomGmsR43p68VnI8Oo
Wjni2FnQEVyImnZfZsRkBf7cZrF4p6OHiN8X3Pcy2qxcKHzPBSS/twTZmnrP
PMuvfMBtfLmGWbVhAaimvjv/WLYa9ssNys2weIVdEM1wwiTo3mK5NL9I5O/x
cTpxrzi/5zRVQ2z92yjN4nMWftLZWlmi5He0d62iXkQJ04gz9B6GcHREUsNi
g2yE0bmPbZqFpG3FsfIidpvMESquDxz7n2tRvLZWDGEY6TqNM7WnY/5exZzO
KpBGRQ/rcJwmrY+VLwJe6fA3ennc1DBFpeIg0KZ9eEgKpsXDXoLdzzHlgCn7
lwI7g7gUL3H9O6TsgqjbEVcOUELKktMGf5ZK/flfA03WfRBx7kiwu6As+Jyb
QCDJxVFP9Gk0sggaeMTh/cw8oBRg2MBjXKw362RU9DC5ig5Xu+9nNInrupAW
Ly3CV2xZ048S+J4oPzW5HbOWSdeH6dAZ1+lCZ6y8ZGreIPXc/HEaYEEbumr8
DM+F+owEB860R3p674y+wigdR/h7CYvAq1PRP4wZzq4ntWh4sLpMSKEfXyxA
NKA+iTclaUNYrNpJqd/FX4kS5fXHjvVmWVv/8Zgm5rraKqJxDbIMrDyN9L93
0goJm1meP4TLWyMrlgLUGh0iFdrvHY0RTk2o2rWg77VOUG10TNUZqmfGM5Za
cTZOUXqmMGP72P3kdiRelGh8M2Tg02QveruAzWsS3jTMz0q1yHfDAJuKTjKp
2XqA1uR4J131ATQ+HTwJa8lsbz6n4VsRLUHukKaOTKp9ydcnEg61Rniq5x8a
xyqT0imG34D4curACrfMlJedHR7MG0ylswstriz6uOwpVrB9jHt0qSL64WTe
v6VXgsr41R0CtG3tHEArmFDbCOJac3JWu6N07CuNsHLaqlE+xNX1tC7hhkUv
I+BXzUff5h7Cl5oYybq4UN/xS0+XklvImH3FVA1JbbafiGs46cPiAxCtCABp
9DScAI/0wYpmjxCxbryELr4AQFX9nQXhL4ukzeeYkzxDEoZdk8ibK4KgdU06
BeHDIdnIx1mEWfTEhKKarXol4A8pCBHGaLyTtEQzoR6VMmFPH0b1V/D5TqHP
2w+NdScaxgEzFx8SDrPFQeRgkOjyXbBzdRau4CVFrke9U3pGXQjs50vBoa1Q
iL9svCqkgXPb/pOVEhN1tu476FD9RmJnpcuK6bVDipxYbJ5LXgWz7KHJi6Gx
Cu6Q/IJXkfwjsBNDyxTC3rbpCk0Mwp+ImNST46cmENcZE27Wn1SWFRcZT+nS
qag7RBNlwsEJj6DuS6EQVRGX7YRRBlNfJb0cw/LZ+UbyKrCtaVrwCJvgKG/q
lGMZtXMAvCSDwHavzQBH21X5zGLFVeMtdkE5BUZoYiErkztofP5yweFUthLY
hMcQQCgrYlbrAQVSVWyS2wNuRCL/iq3KmKaVW+gNNrgerBlE/zneeXQ6mfBN
IFOuYhcRH19h58PZ5eVw3+DoO7WhPVFaA37PQaANke+RQ1sSNmvphEzr9LSG
Bo2wMa7/pXWA4a0+QXwcGcO8VLG8cMTVgjir5R/GuIAy+Vga03YQ71Xi2ouO
usA07hQVoiP/jm2TULwSSebm1OuAwE9nbWzKLykQXIYY1YbdBoTfTRdipV4q
73HtCcmrJKTyurKTJm26L7nQAbRX6BFou6D2vhVU4FASHgnarWX4MDqiW97Z
JdQ23HAViDwWD9c1gqHelqKPgrS+sq96V1Z6wMxi7GaCdmx0VnJTUHFWdRoX
+sh6kjZ6M503HlN+u5lqQAmebka9DQAQwrhrA2RBWUD7hFHP4TVDXYZOmm1b
yHkzU4mCcmhuREDuMJnUmTsnUBG9Ka25A8yZZS7YagElPs/2lEkMBn7GdZ8h
/aWeXMeJLZo6nwEfyVTXBOZt12j1EqgasFwUWULBn7usWoFWsuJeMs9a9yhc
aGyq74gCnFvD6zoMRaoXlfb5jTGjk6woDJMFcjlc/KvXFWu+jYhv/3jSpLuv
Sv0skQDr2p6O50st2v1WAYLDobhdaxVuXWh8cIDQxFO8PNCdoZNR5keI2d3F
Qp8mUZ4o19X1t1QEvron/9PqZmGcU5/0WG+CZdZ9Jsf0KSYpmUuLDaphAOy7
knwFKlA20GWQzdgneOmRfQ03aGQ4r5LU3310c0fJipwZ0QzZI46q1GxuB8St
uOYFR1BXYKtjNI2WfL1KYWDjb/PFgH3WMqLCrXeNi1UJVpU5kNNx3vLUCoh/
KSNcL6402c7c6xQZkqPBvoGJw4oIEQlwbFXuJaqJeRvN+Fz79vZ5B9791AiS
bjWiP59OtvUphyWHQs889XimTLRqO/myqz9Y2EfqpaZEpgiMGiqEHkgwvbij
Fx+nmF8qoYxHdtI+0T5aY0QsXQvy38mO4mDvl/whmocDS+X3cwwaL5eJhM1H
Tn2FD7PjIRp8iHuxVaqPQf9eJDh/28qF40Yn4czeC2/xKPfSjp2eR1Ip+aUd
cxRcfBGwJvveAfoqOamqTHkY5jIMV3t+lSgGS7O5h/Y4OvhftANKGn3LhWWG
2ffbxfAr7XaW3RdWxGJcv2lTNqzpjUMa0k0RAxDxQ66YrvOzsERlA/ftJF6S
3hOkbttsV3e2ytdkSO58o2lZqRjDgxUGw6f7wqo1f1cJv3VnPhk9ZTfFE6aV
vJA2J28rRiND1VImAsFUZ0mNuYOapqJZqhLEMe5HlQcvGBdzOW9Oil3xcVHd
2HuXFsvEPCBciLp2OxXslI/53UfTCsoEnLzQRYoXI/tQ3dYZZl10AcXgCBFy
sGp+IX5cZ0C/XNgUxN4alwqYqU3ZbXSCRHcXQmD0aNVQh3UiB+ivZ48xoiQp
DrqNX0UdEVnHfxyAUj7qqJf/EkfFka2XqmDCTsxRQixTRFArlzLd+75kGgTn
pgr0KF1qVhMdv7fbISmCXZJ0TcW1JiV8I5oJ01fsvtbsxwGjMF0xX/nB08pt
KeEwYyo69JUGl12F9ymwhpEf0O5KwwkahNnocVWBSVERVgZK1UpVVqa6kR7l
eL5tvef7jwZd89BDpi6mSpptlPt6NLFF3YSL9ieC1vq8lLnHCYZgWuM8sVx6
o03f0ZzeqJEuYkcYeIju4FqxQ/N5+Ib5N/MWFGPjMnZOtfYBsw23GpKSLnzc
uLlogZDvKYzILigbeTPNcrgJf4Z6SO8/CkPLX6gIsffHkkUF/dINJI0dMeZ5
5QNElQrl6bfP2AgKnwLIh+kXWXnjT6Pl9yE1Qno6oBX10zKajRtUNa0yvkyg
KNGrwr/9LlqsOHgyVGBEV5LLODOckTlfvsxeBi4bWFd2xOgpxMCNOnp1C2Bu
TCF23HZymvO73TGo3qqYgZQixsT3tYFjVGsqszl7SgUxau9Z38AqfGNHXjEW
RLdyegnPUqz7O2kY4YiGaOxjarDTsg9QBRhBG1KYX038KrItmYJr3atn0nVv
2C2lt6BpQexstFvTdrJGpjaBAhiv+4ueFi7D/lVEeRXtZ4VO/0h9ZAHkhQOv
LJdfueEI/huXzqO1nvNwHbZgw+1gEufz/WrZmCUXVjoBu2241bCgd6OLRS0L
yRTr1Q8iI8RxtgXrYjNnwoanGhcUjPsT6aGl5wiA7psNxE1uxZR/bG4b7gDp
P8YuvCRRhOt4rm2NVsXrk2Zy5X9YgxU4UvoKij77atU8xlzNX4UvDrICgwIu
10JbWfikHk7+B5XluQ/mpmBwGAEe1z/mNEuDzXrz0nF8tjvsceNurxBu9B9U
jMxU5b6Sm97NhP6WBJMVznv/euvZtf9qlsUH3mmojdsPXO01rUYWX5xhge90
tJmT3C/jIHg/VELb1HKIOvCjE7dub4/ZgsFFNoIt2bpgEGtkfY2S5d/t3qrz
JXIoHmIQbI9EIu9X5gnojnDTqjo8wtTygCa3rdy0G4QfH+6WMDdv/DpVPiJF
QYnCtfuxnb1PDq2m7W6lKD6g/+SzeIKpCqFyFkFT/2YNjxoEN21WHE2Yd7RN
m7NxlrVhCfkgGpcL36CO4JiLobuY8tZzbIzgbDpbeiRiIzNEKSzlaTOhlgFF
1tMH/cIEJhweRChObLXP/pN4mgJ/RpQOCMBADbTpnmriO5C3doDv4ViMrn1P
H+qcd7A106Pqoow6arq7zJpyMuxjugkwKCAvlAJHBjm6Wc/HtipAT5mz4X64
YpxQ0N4YOHeKljsmyGcXTn2VRa0hBejGatmqYLIvKtXD3Pg9G6FM/WPraCMB
TU3m8I+E2AICEQJvHUsRDgYkbJ5UzrvtuOKplG2NJtofALgx8guEAApEhGF1
CbPDV3GBrAzH1LqNeBuVhzH2EscRTs3Bkzt72kFh9nIzG1/GIjgMyBSCJqEX
Ky/Pf2uyKhU+b01HasinkTZHVT6KVl9Kmnz58xYNlkQY17pVUG5WFqzc+vKW
Sqp12Aye91MN2RdeqGXtk3os2T9UoQwZhUfDeyVXInYszcgvhDXNZXJOM91m
uyuBDvbe9b+F+DC1XkZRCQm1KgqWGjkGkfMcLo0uy6YoglY7CxQKJzp6+A4O
PqjZEU3XcWVnOy9hoVn0DVAfGZjPt/cUvx5TqV8++ZyR4jaa+6PA3jtQx1PV
E5eQ17UJd0Kf+OSA0JD92zGuM/PjoH/fveCss5396rUeVohVKPkttV/kUfCw
7MLPHHeExccCzj1tUkInaGIoofelN5qTPIU1vrcQgcZp8s+OFwot/Fh4TVQ9
RPoKznrL2do69DUIy1/l+Vz8XciYSzIm+9EJVozI951n60vRLk9O+zNtfLGz
KvKi+zHsY1zYDN2z92cEuwIq5awIm2vSl+QvAyeSLf6yCqmXn+ScrlgJBSQ6
isMMJUL9TkTDFP2+eZ5jK1vwvvcQsCRcBKqKFeVuxnHu5W/ofAjzrmYB02ai
DPvwbnJ9sLw3jo6zlAQCtN25oWmTlUmf0+bsamT+NeSg0t97pJUrmBJtTwIB
hzpBboYHEYWDJtqu1g+TO6H5RV9ulnZ+d/kKdMIoXAwCbLCfDqb44jPl8R9L
ionTldwOvW/dOU7tQefjHAUnMOwvTyMkSeynjzZjH423ZbzhsMJqnaQtjhAz
V1/5A+c9g2jklwJKM7SQ0cIBG0owyFIN+bfJOtCkN0SURL7cu7kn3UUrdmVi
S0xlfKkoyLPZTh8vTZshJ1Kwc4+aVv+rqt6KFNosIAVhVbSWYhBgz1L8gdQg
q9wo7hirSS8y4yO/gD3cp2t1noPBQFQkeyYHesbLN8byFDKPAvQFXBFOyO4K
59Q2MIokS2H+RKspL0x97kstPrIOdBxt/pKWDg8czcDTF5hpwZSf4QWQ4MW8
kDX1TH4fJJrBmtptXLINiBAxNPvZJq/fUcalBsIhEvb5dDahgO/hudByAjaE
HMV5nctzAZbu0skMVeVix0pCjviQbExFckPxoZXh0T9grdw/P2XyGABTg9C6
yqTks6kDOP/wjVKeNXutYFafMBeijp5x2qUk6Tuf3qzlXe7CQJ9RAblzV07M
ROepiK0GRL94oIB7su0OIdJ2rvNfhIv/inKhZ+UcFB8CE8pXBovLfec3lurn
FiXiC725vaj3VESkRB4wvgzENMzz6T4rF6xYgohJgQa9IDQ8D+ZqxZpdvzRE
gCcL2gPHwCRHuCsPg45/H8tb4qCvHVhpaDC9TCklTa72C0iSoLap6TfJE9WI
4kogvNeHwVh8EMRfiAfou3rYSo8n68XnA0Tkd7kYTklJP3Nl6H+lk8rztZfV
pRP8tJubtURbKmv233VhoKk745dUpIVRxok3efRAeNdHBKjOnqmA9gFKODdy
BNh0K/hg5gi4vIXEgNXFDw+N711QkHVVRSM4Gtfy7Gipi/IEJILSs/99IXlN
ex0EU9y3fbw8ml82QELZ2P3zfl1jpGCWsLlhy+dVbq6HBabDIQLH8xgaESRJ
ZUYK4Ccb2nHHiOlb5pEp1otXN0PpGP24NOZEF+ndIiO6jloFVAF+OTeqO8F1
iRFfxnK42lU+73yW24w9LZrB+DPTUzSwVFoScYeF1mWzI57FgBOph89yfyVe
GZ1w7loTp5S/NHy/JkWFkN3irP0KjXGbet/wM8RTHl+I14cfj2VIbxSeNujE
oojmBzBmRRzovWaoOF6CZ5YhqqREKiJT4kmUJcK0Q0rxlq/hCWxCWapXnKgo
8Gp1a9wGzT0z5hkTY5X/qnaCyJE/a1+p+wr+eYBFdiEWdkrzHjfYdhN4W4Op
lNCNp+7UG5uqR0EWeG321ZOoISy9cW1EnBtPkyQdf0JPV2MwVYPspqk8rXP6
L3BhgbSZ81nJ+Sz0ZkMxVEAIAX+Zg0ZPW68Bcws7aUiktF8u4E3G7YJ1im2R
5+LlkFkrcgrcyXS/ghLFnyvDI5AZQZIyAnLMPBUE1r4GzOPggT1GRNCGBElr
2kArHt3LjdDKkz9krpMzobpcLTwv1aHqA4DpSiP7c35/R9oPOUpFQBlHZOqu
Bwc+LtNNCB3LwiV5W/IElY4fObFmmwfGt5I/R/wuq2rhse5S1LukXYugp1U9
UmYhIu71lFMc6EM5/tvqTIRsCliT/R7zwbQyxHNiOJV9wAtYCZk5aCx4Yz5o
ZGqSwmazImRyviERG9O1JsV7ov7PDwDque+zJO/GO+v2pPI6tCUA8eXvXXn7
3KnSyDnQ/1r2rognu3JPTUE2Ik69iMVWzdvwoqMZ79CS9e7d9DA5Zrl29TBL
5SHdwGjnoHPzBcdvPR/pv36pvakSChbvQwc8jEjI7N3GuZFbUfhFSxttLfS+
pQlhWjZmemP93YyvLQ+FKrTwBixIDRRGDu0geiQdjKS2B9bqmlytnXjev2iS
ao2Wz9DHz1CHMfXpc0+JheocIzftzaRsd5G6vQT1XHI4ESWB3IzkFc4MvMUZ
Ug5EaflUhlUOqXidF94K1VJsd/4y+OC12rI79/SR10/uwDrWQOdkw6jkfm1i
GmwuPR+YzqRcPg8LZ/RZcmmaDDZ/V+0Qf6VGMrxrT0FeIdGqqZexF1qsmL+s
rliY50gE9wP/b36Fiuxr7dMEZdxc7YPhZU3BKG+LKiMV2OfCkIVpHk7UrtX/
yVRO5SLctQ0HTKxUpZLKJ6pJr4MrD7EIMTu38n9xGFrHPJxAU9CwBF3vJK6j
gCBBGNojYChy13/fektJ4DyUnKM/o+35WwU29S67XMN2vcRH97EuySAOXMps
JrM0puY/svBFbzMUc6IASJLDCE2IckjAoiNqNtifFZ1Ur+pwyY3+WJvRDjUW
VMtbDu3VG2QQupA3Q4aeFVOy/9VM9v6ttQrSNAD3RLksNc8S1cl2s8Jtb6Wn
jWlqsMcpSuFd9FvB8gDIpr9RlG8hZ9CvKcWagHc6COmRiO7PxRIsmNDfiQle
dHrSWPlOwRGNguXFslUXcqY0WYEWNI2JK5U3xoDZK4yk9/3v9aq1lEaYCWYD
eagoaM7QC8fX2+QtEqluhrzFpwARTq6mjd4Fhr1jRSiG7dc17HQQ9KNL+Txn
VJT/NDD4LajUymwaTdFvH3edxfU82cGPfvRo2+UxbI/njDouLiPeeIHjzmdT
Wq2weh8Wj+V14/cJMDG42jEurYBpIwdiXfa7Difiu602wtZxNUIh6vvWQcHO
Z+zSO8EmQzZ7wHjWanueIm/A+JGAF4Udq35zWTsvTPn/iy3rchXttVkhJoqq
2sAWUG+YJI1BLPkL60MHPxISn4Sw5xb+JnYv9JpmHZy708zK6qQsHJnEvEsN
yoogP4rTUDIvpaVkH+qZuOce+R5YU2iOjLtQZs1nZmcJPf8Yni0tV/7Lt1Ih
bobUdWf4bf8yhCDINlcof2WEn8UOgN5Qvqk/qQwrd9sFY15QgkRwg52ud1Tv
mqzYBdiMFhTqCdm20PidtMh7IGdzzKTPWlVcwwcKcS9VJm5dg/E95I9dYahe
lilAu6jk2g7kMDGkMLPUcdYCzzmQks2YQMWMcMRqPW9350Bpq2Yh/yiw1dTt
R/0CyLDo9WinqoI7GKfdG3gCCFzsAvmvloujFndhh4PRT1Z8py/YFGCrqAx4
/zp6Ar0L83Nq2logJSpoIo4E/Q42N8/K+bAt3G0P0KAge5A02WY4jdivCy2D
5WqVgTSM2RMYsZuuZI5lQ6KxApEtfEE1KOyZSs32lyFK9YFVzmjx9D0ibJ+M
A9xVeWi8OZHa2lOiEYF3qJ0vp7BbeKkyNIukJxrVofgZZflTGuDt6QCGbMRI
W4eBcWHPawIgghFS+kS/IPJlyTG2L3uWz5/0vACo3J0Sr1woI6qAyrOkUyLs
K/Gj2gKLRYiwDWY3aEEIKpBrPd5z9ZsiPu8vSl+FSW3XvoXVTM4k4K5xWEKy
wsEEomwhSSI679K9nyBNqCojb2n+rghqNe3yj1WAn8v+UrjRA6fELrhHVRtr
z1qViqg4ej8D3ZXlrwi4JtIZJrb5yH3jJmiTjhtxzp/1Y4M4ETpH88PQN3nQ
mrPMXVcoXuHXbPnnZGbMuvuGNddCGVpRmGW37H+DioTRfW76ZreESw/lUktd
ntvCcV14sipsltC5i4xofutY9MBl//p0r25u/DzG0WUlCH2zOwUxpRPJWiot
EyGjGCeK0URxuhuiclYmRi7PbR9k6Z0hks+gsCcNvSw6Xo359u+Ol6gQ7uc3
bupLam/I2iqhFJecOuxZyR5dafjXGYwFHJmNzTEv9FcfWo4LwbN0cbYdUQ76
DUr6V5KYB1wAQuKkTpZhOJO1ns2dasDI+fHbFbD0xdJhABBL7RxDcn/dpjOz
yPRTcKg9pmeYn4gVkxlUKdO4AtZoDKt4Bhh3Kg6MYeU9YGBjoV6m7HjxB52C
RMHge4Y7Obp3B9VjP0r1X9rglhCqv6Nl/cPbd3LkX9kAELkF7Dr3HumM/0sS
Mc+Hj5qVSbWFrYBqiwXqJioQpVu2JHqdfjwSXWYc5Ug9zAHmxePAa7gJtYeV
m5l4NtbykQHwmlRdyMhvXOO8qwMwYLD8IZlTY8hNg9ytvhbImmy+eeqSbFJV
0gE+NMzdmPab0Lfxnisv892YOi2MCCtVV++ALDpBjsaHvvClKkbNRTBY4kRt
7IOCamTuClGurfo2sDYcAdZBStuMhPgENw0Mg8iVQ6ibz5kG4etqvMazWePq
75eUVBvlwhaLmeew3aXcG/+8GCbxUs2cvrhnpMO5vg2lsrvJWvHkZEZ26Ly7
p4NpYa+nYv/u5QaVS9BSDcRjWSbWB+0E2rxGuFeqP4IOwPBdEpaBnLFlw0wq
mV6I+IDsUDEBkWBobCvWw2wxm9eug47gjaKSTWsb5gXu4KjCLK9hKtZy9Lqa
QHb2dQ5Kb1+DzyQfcwV23hLdJ/NLB0BH3J8AsKg8L8g5zZnNHyR69ZaZv1fg
jG596/Z4wpHBpi+7//ccdIUTAzi2NDMtLKvWT1g1teGWC6Mr/TO5VD+XL3Ma
giq3t2kq6Dpqsgmb4sBXpKgjoDGvwrnmjBOJx3X9hh89Fachu+H5SWQCHNmI
8L0vju1jWNPA4j0zqNcWxVW52/uDMei9+VIpC03hSe4Dnabbb0264nRCThU8
JO3SRgvW5JKRl/z95ZlMu8rbaVv90EULeocb9q2etjtvfsebFwT26xJky5ud
bXb+AwT7jUcNv00loZtNIaGWP7ejdqL6S6CN3kF+xvAIluBZ3mZDIe3sXocL
qgyEg/ZBYeUXXkW4sW8CzOBidbLs5yW8XJdtn0tnVs2GbAA0aBim7GEYko4R
TF4Qjff2303AzFMSuyugiIlf0rSrPUtScJkI1lChhDST/pBJNUqJfItxSe89
kdFb2VKAi00XBsYg7UJrE4qlMowq7rtgYWw2pQhf0y0dZVj6th8lwz9fseFM
p8CyY6ofU1hsGuzonppkwa+k6Hiuw1xaHenr8yOh6nmZNnwrU6180tcJ+cRw
N+h1U67kPcPPfNw+RNRggaCmlykZIaO7QezkjYtTHISMhdsSBZ6BdywUp61T
5mrLW2l86MOTzMofG4gBwjbV6QZto4qaB6Z5iZVl/J75EwSpNsQg0INcdmpT
5AtXAqwM06G0BgSvoVAc1iDywWjkj8BFlAmNCQrVvd75B9p84Md5uW60N1HI
K/0/SG/OWSu8pVBBgNzCLk/FtB3hExArmqSF8Orp/O6S+IBVK69POKZSZB65
XQNmxhDWxm5K0DjPcHM+OLsT5UNEsJbKEphYha+SXWweY3dcTQ/bKjKvuets
18vImugSS1H6+mAoegtliKxN4BQmLF+PvrFDza40Xb7JbBjQhGwmWAG3OvU4
bktx5/D+qEheZf25NZdK/4OMiF5nXiIUUhPyL43Mak5c8g2+AgxfULasDNi/
9yuKPgSAhV7AF7CW8x80BA1jrIeMgIv79k/kxykmeFVRFahEFfKIbUAj3KZZ
QcymOJvi5IV7cBGcaex6snLjjrx0VAqGeZ1Lj0rmUhDY301ucYwhs6jQjGJ9
s4DD1YLrUJuuNNKg9N381l4vUbSNg09biAQVAshpjEk+OOgcf6smPjKe/GRI
J21CVOdguma4VV1Lk58qzGl+t0AePvgR3paljZ/1SM9pCpsd8GAyiP1HnLQ9
CJNnsZC6rvU6+nUOUAh21jfl2QzFMtZRAlYRyrQJocM0xKiwzkrvtdkDIXpi
ssNNWnx+Ybu2SBkSZgcIis0RNtuFKhnBmEdtfdPRf7ty62/aTv9VSF187WVQ
pEJCUIBWN4FQ5FOJA8wCwyYABXdTy4OphNX/BTr80uuTm083PZKJixHZr9BF
TkHQR9nbwwZVHrZABfZrc6OBn6KeqMfzrKim7GgpwtSiQdqLkjrvsFifFhI3
IJBnn/4Voy7hDOz7RfqXavQNVSPgRRfM50uYKIljWcUccL4jea/18I3RZ8Dq
r4EwMy+eoPOqP32chkS1koh2x0ITicgRQZlGn/3FQS3vziUOdfs3Lk+mT399
slp3+6TrsqP1eVZVHghI6sRLXJLbmS2OoG5ypDHxQbKLoI4Q1PAc3yyFnuC/
PadiQ5t0kRr9+SfGPlasK60vELuRIZlU/ZgFyqE0TgtY3bQ9B5sEKLJ1pF8p
6Tc22FOylpzoeGhf1oSat3D+7HUgGYwmfXoGuuWVkmG6AfAfxYAZ5P+X8etF
+na22VIF/SN5BOSVBKk9AY+Ipd+bENowDiu8Ji5RZfNbK2R6Y/zUrScr/41k
8H3C4s3a7dpZpauE2iYiHKX0dwXKOtzsjaA2QyDVeg7pQhBIK6gEtmfcrztb
AHBITFG34YrewpRlQJK2hc/dg256LgIK/rmtEdgqcau1pcnidtqZKrsjky07
OI5WEnOn4Qt8nkKVq7I+bjjpZRrNiMV9Xg5sJOi3q+IZI6gkRxTL2plXMefD
xczQAqYqz8URxlebtbgaMfezMtvFk6mCkid9nvBPiPTfIGlo2UCinPixeeNh
igOgWEjBjwfXQjaeWvvx3h3B0l8H6eEkJMBqhjhLnMpMI8Kgdazklcd2TIzE
2YdNKI6OS7TiSGhUrvdf3h7/DwOoNBM9es7TvuGJtMpVygpL9eo4SrbEeSom
e0JBxS+2l6N5yYNyxTUz/gHyW+NXvs5/PdptzIVqm/n4TI/yFBaDHdr2Eqzb
OmHgEpfiPyOMXRA9Ji6ojVdBQWZs++l+D2TK9uu2yiKHLrWGgrbcg04EjO7F
t4Fl7HrKzl3wWPFJuaXkVa6oSpJkFkd5hVUWTKm4ygQR3UIl22AZWEZJA2hE
ILKhD2UIMMUptXUXgSdyYirxCgD+KmMWGgQ2eWOngVyR76EtEoEycR/rP2a8
A5CVIBk2RzJ70oSFlgRi/GYVjd80M1/MSjJKL9erA4aBdNkQmaDP5qtFohn9
oUnZ+hf/hLPUaADHXEJeFmt6c8LkXt6H0HQII6pCK2V+d587QtQeJ+fHm4Pz
0Q056sEHYgZ12jI2VzOo/FdoJ+kwDNRPSunPNDSGKzaWnUF68PnBzZ+YqmDM
w2E/SssFwZXuGf+A790tT4FQoVt7bBTWkKi74juHoMlsmQQxUfBWYdEkN4NW
F5qrC6lIp6JB15bmcPmbXIFspFXJ0Ihg5C5YgwDPOZou3Qt2Zb8fy8qoCC//
FL/EL1qpIkp4+R/eb+1u2cNWhg4UayiecNK2sAGFnBfzEprBwwDADRkQfKEI
LPfqqzhc+5Bhn2xmGVXnB3UraNTBzev2/LTiiMU5XJM6ePZ0xtt2hqL6wL9O
UUhSt2PL+Jw8u7bTFPYn9XgxZbl9z+v+57UvtF9w8ZunuFfA7rAQd7pcHpWt
8xY0kBShFwEmf4MBm6w1YucQONI3Ju7q1UlhFqY441UNelFy7iIMH+10YG4e
aOE3te5xmuzpXd2oZK1ontzpfjV7vT7j5egKBztKJonKAQUcqM7Ls/WX3qCq
8ZI=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KkMNIwxRme6bqdrcY1NLXxQQjVQv5QmXRvttm4T5sHB6ryJiitEGYreRWaQqqjGrggxKINqxbBJwoUXJCvw7pRWdBlxXWbHflmEUctkZF6jp0maCntFxXWDMBogCctht9A//KzwlvhbE5SZ+wyJ3TBmPvOh4GatHHotFskJ2IiES4NsYLPqM9+jtx7gUfv+yr48GGqYJ1FjY2LBd8YePUreE+1vLdlHC5t7ivGS5PfEVJOG68JfUXXKX/+56Jpkj5akUanfAuQdC1IIZrqvTCNLtDPsBL/6H1C21B+Gd2BFKkv1DkMSg1swBozQvWS+tIp6cvDpcJzFWI0I2elH2jXbvF/24Ab80w6UFcQoNPHWYFLdhNDvLzYyKgEoRA+I3ZfEKh9BMn535+5wpkvJLl3LEe/neoR0IBBXSLH6IbPdtIDFYm5huYAtuEfsxg+dl85rK8Yl45Mvq39ji1TdWHwwSZl52N+nfVh+ojxiwPTI1Qv9cmIrCkRmXr3L6NbIhoMTfh/FQNV7UAxnq8xAjIb3gGLywilMePROtLU1az7Ma+7+E3U3V5Ylmrboasg80rRV62DGPH7N4cwvzQwdEJeBH+rdBHAzXjD3W+op3j7wJs3CbMI/0BnPnLzcmMd8u0F7LmZJJCLMK0DK29b2/cIs8ZpGsPw8X61bHgyUYt/dkK5mUW8c4161734NtKlI+6jsbHfyFSxehOr5WOzNw1e4WI/Q3bJl/DH4U0m2oTtoUvcTd7b4xPRiKDNFIHffR7n6lL2GBMClB3EIAg6idUp"
`endif