// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ayxqyaIDLgBeYWjeDmZLNVMwCSD8K+1guwmlwhYx5oADz5ipz+/cO/04tgd4
C9OXIpSKbRZyymCyUIHJdlBFYRLvExbfI6/LjGAOlXMGZr6jVdToPO0ByVUd
jOvSSlSDze/AcMgGLKZFqKudUUVt2YBDWcf+E2pgTl+LduAyddqdf0V8saiW
jnva7sRxgpejLkr8OjpL6OT7bmTf0ndi7HVlU6bDNILFuR1U1FTN5l058Xjk
s7zKDIoLuTlzTCynM/6Ja5ypFdGVqlYk6jcZeCwWgIZKHf+vAb1hJ/mrUyLw
LCZFIuvPoxhSykuGczYnHgeH4F1k34WsFXNYR+eOdg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SfdQ9AG76K1DPExw1GHLVHVuW/8nkUNYMwf6mfQ6lJvuogaJFPqGfLe8cBGi
kf5oZoM2DdJY5qXWic1fKK1xXV4HQlpP0I83jiHqwNtVIyZUs1uHdPsCRpME
0eLYwI0tY35HrsUyIpb992KKopjgGHvQ2+ax+NyEsni+tAo5AA8xdmFuGCS2
vyO5pZWyeHY+Yzd5TNqxWYHpKxlVXm/tgh45AGDxA1Flzi9nlY4Sl508OWrR
OvaNaaM0HED5F8adfsoASvrmAzQTvdfw59z/3c1r8rktS1HvuYzCF8x6F6Dl
nAHSeKwzv7mUFpQCmZXdWj4mEdCgdkwRyNvR82jX4Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LOyWgSdijJd73wp7MPKZ1PtEwfbWp420Gj8Bc0MOpf8/fveeQkJihbN/2/dU
jHgVty32A3Dwm+VybgDi+RpCofjawOhXnd69QkCPd1fqkwwBL6mZFKxsUI8B
DsKzM1sM+7bj0m5NOQIvkvrtImj/xm5zVndEUP++aaWUb8SSJutI2GW1pjUB
HhkXZFJA9mKomR3uzPbxNp+YunO/ia0jywGZFD8UHPJiXmJ4lHT4rsRrj83K
080I+PhG8bL5YoYrfPpMY4oFmEtuzhV7uVjG9K2aoWfdW29haaIe7T39riWO
LKEbHHRSGy/vYZ7SXLPGwPS1xy431Bueg05tH9jVWQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dVZW6eXICHuxnbX4toG3dZ85fNV9YR4xIuDRLJ99xQya1EPgErIY064Cn9Hb
vAeLKANd7jkqmYx36LOD02JMUlouPndvOTOrdEYzt/yui7qq4dPBpPShS9hC
DIML64mdyULqcjjC4F1gFQa15j8NfbMkRq05htUIXB4qM0pISzl9RGp4lQ8X
kpE5MeVU2FakaszzQ/Uh0D2kDEoA6YeC9a8xHIyrmGih/mb6j3MsRCDd7ySG
QqWLZzFX9TuTKABJgv2FuIClwdxeZGqE/u3QZVFzMF9dit6SCEpBfFJZdZKF
Zdj0Vd1KPkF2fVK6avyexpchd38fnQzyBBcPvDXXPw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NqvdEWqJaUPwA+OHmnP/XczT8hKq0uA5Q9B52yui3O1cnCqhtUvYKV+z33lq
5FBV/kBUnzW+rNsMD+fsjlnf+Isb6tZREqN6ft3eX7WZJDv3/yHSgk1Aqs2/
nevjdmL5d2+uaR5KOTesIclPmyrD9nUbsqtwfdrCdQV1dCxEPG4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PGLXD6klJt2wTgO0hy7fwBrDnw5IFUC/VtVKO7qXPpPOMnbcbt4o5sFwKwCM
3gSgJ3rmjV8WvkcExW5nLmVUrWAJyQt1RIb9UlTaJNVUZMA1T0FsNcJHgVKh
ywhpHbQGyihAhL/xq8064rHuVzbN+/r6xt1FJWXkIl6/FS7jCTt2vyuF6Aea
CQPV+zkEhdL0iA3Reb32AFaUtMrrv8T3GFQZCl+k8Gua7RaCJi4JdR8Ojey/
bW94/ls4naG17QgpEC8A2b3vzDQsAKBk4qTtnH3wd2Js7wlIpopmE0gEGOpL
neacd+17C6WES5Di3nOoua7r0DcPTUTSwsDcKcDCP1Yb2rnprzerQKNlWeZq
tiLhw9Y1GEnLT66WEFQATQUx5NpDJlWSTkN3hVkIR1wDAjex0J45aZI24ooR
eVfiiIA7QBpLKPDO9XM9LkDbFHtd3pMuPTSt7VZbmkRlLZPdi++0bQWy7hJS
F5NaRYvHh+KXSF9QXijXLnGdv1U0NLJU


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ChR51S1aSscrz1vR2y9uUz8gGX7pk52GTjtSLTm6xYv6j3LFMSZZ7GSAiVaq
y/FTdXF/mv3XwQxKSnFHQcLi/4nhwdP3POCAbVuViL+wC7qHCoV7Ohr1OM3w
gNs7hSATy6oS6SlfHanh0vqaEB8YQ29Vgo52sCJ90fNxWvTkrV8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XpVAN41rUJyeHcPhXKusfs4i7W9XB9FPKBxd8eksb/SRqAftxQGBNeFsHx9e
TMrmakEPGSY+txNg9G/Jws0TUpl2rWcLwaUoHQR8coZWDwWuLFqA8zqLNZ7q
mf6PJSOJ+TmEnlhg8T+g5MNcMzhRkV8P1Ik/ExramGL6aXpTHYQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7584)
`pragma protect data_block
Ym8HqBuksvXwxeQX4906326/l+pjlVac5C7mb74bBQTkR5HrSk7jgiO/8GAA
Ha9mOVQ1cN89hcZpUVG37dxkF0zCuW5jZmU7O82D1A4bF1Z46GBMtELiM2rD
NBnpbslFUo6Gqc9q9FLEIA32X1R5/gUoa4YG8QCKc2KakR804utsr91IIv2O
8zLiMZUpwb8R2hSWMgfMsWbR8dcCbWQHZoaoq6qlcdLsR4HExqj/+6ypBFos
6pn4D5d80bSQCf3muv0QOdi87oDKSBa1e6cWy8w9xdXlZp+mAK9v1cA6Tqj0
0qEtQKcAkptPJT/YcA5dit4Uly/ozsKrRJT8ERjLWQygANtws41FH7yg0XyN
gyFB7TkjlH1AcMjrw4YlBVCKobeLI4cfOHEp9wQy6yzhukdRZA+Hd4ULc/S8
xX3S7mbFOCFGPOXRxGcQ2FqZGLwHEdVAqnESd5kOvxixCTmtCQIexbMv8I8T
b4q7v8Rv+Uk2J76xlijxTobG9n7vSoWWuv1bBtsHstI0nSHAMZdcjOZ7NRfg
MxODIEP5r3Zh2wEdHHeXmQ2jzBZP7b8iyPzPHirmahaL2sPVlMHdXQB9ZJW1
KV+ZhoImq7ap4XDZ8czlRefnVxKrxlzJY8Rdzbk++2iuN/oQATcxM2E8yc3I
f88jhgMs0kejVcnvh1fpwvIt1EmDKEUATKaRFrRumStSdIH1JOAeoKdVHFIy
nrZ+ITQ4yW2TSw0OszbOEiCZ7yeflBpt+dF8eujIugcpVZ1hsJNw+0Y4oyO8
j5WOsQKO85auBxHto1+cLZ0Mwn6zMZ4dTsURzeZWKQIcFhLvWjkUi5v7agQl
HdGRwL6e0hv/v3xPtfNM9nHP3mVCW0hRCY0CudRBgsnAPnjFwC3hgi3mXuIp
tlGGydGQ9S1QK1I1ccIvbBNLyeSxqmdhqKHVbZTAvjE5fqlULokQkbvTi+6Q
AuwpV6EoFkWj38qTrc11cEuZmmOB7atRMPlx7CMg37Jrdkn34gcE8cjm3tnK
NmysCPYBTXoO8TAEWJwjpToJA4ny01zqACHjA5umjTiHhdBC7WxN/567huTm
tB2cEaTdgK86aewlTwwuX0VLkI1L+Q8aHSkOJNnErrCRY7k9jVkgwVhSLXIR
N7Bmg7LKDKnELYR3pNUPfO3ZO3yH3Qr5yBQSSJLw9pmmBwWthSq7ieyRqD0Y
8wDFcLU49S00TKE+3uMC4v578wvSxt4Bhmi8sOKSYYrKgtdLgLrh65Vuvich
5byns3S/2Z8S4kGrEjC/QMbZQfIuuS++OAZWYxJirS1gfjN3xweXbvJjg4KH
iRGRC0BlVHL2s22IAp2sa5iLsGqEfwKfu5jjHyregQIFJSMpcW/ts2sOiZsh
Twa7nxeMNzbsG4Zbf73owG66xfzrcp5GXWiBO5IKIysk/ZqVSE6OmBBxSmSC
ToADu4Pvqvy6S+pvnPpy8FbjUVUBN5ti7OVOJjjqnyYPlQZJYyLmdkByDv8n
LgpPaKBFgHh7V0oG5E1PDWjbE2ARJbRPf89YocACEsqDTz8ixML1c7jaw5DD
4NYcWYu4tBoJztT1R5ojopfO9wG9bCRrbqeiBz2+39Gfm3/7GaGpLvVEqSM6
A2HgCjPCQgPJUxVclQWS5Bedrnb6hBTiP65FAz8iNmFVzrZxw5fN6WcVXtHp
dn+l2+BieQklmtIQCD6nV/UCKByoHvvi0YvKt7vm9vkW2hwuDCxTJEkY3XYc
MuOZqQAwUA5AUPXPzpdXyS0alK26+0teu9ekEet8lLbU2YPMJRqgQae9KRtz
Z1t8kHkWXjmk9Awp4XY2c6tMsdm+1b0Bvxdt+GnOdQBK+YgbCkjSws0YNtTj
BVDwhfR8MBs6wkftitU5jsAvIb91QtFi1AQ3dOqFlnliSL4dMA6bMa4YrRN9
+ueECDIVozhprLO3pgx+DqlmPk3zKpesDY6JgAsXCHWyFvkZ7Gi8nxuEISk/
uMsQ9w91j1qZpnR5PMaE+5V+/AYvW1a1AF1gtBHOYuwQQbmuXUbrEScDn+co
Xp10YV2vQKtI9xQuij5uZCi8mFyk3quW22nuk9cbihSBCazhFoNSqjjyK8Oa
f8VJyKl+eL2A6MfccoUtSYcD/yuOePdzmFTpSgoXveh/y32Q5sJbn8zVwvX3
GM6YynuHfVFNAm5aYaqW4v5hgy8OAcw0NBZfr/cRe880ds0mbwYAg4/nkkK6
8D40L6qKpLp6iK7qWZ42Rag9NpWA/KBQTJND++AF+LZm7zdqqmcVdNlIpGUq
0Yv6joQR3w/ih7wt2XC7Pl7lfUyXFqfT9Tvmc6KRWdWAns9a48DaVyQspMCX
pyITCCWxI1wbmqs824jURqiSzBd6Qq/W7tvuOyZt4lJC3eLqMF2c9aXG8H7u
MAsONc6kBqOHtu3V8a4DdxdfUDLk6t4so41GlZuerVMTeHIh7FrtAA0QgbTK
7HQS+pTiiA6eJm7wvVEY+zob3OtDHzkYDdul3KCNYxkLQzb6VSD9cdCHP7rV
2MkyYvPDFs3CFJJXilw+AqFB4wBonpS0iaIlo1zEPXzgK6wbQNo6F6iJkkQx
t1v67j1TTYK4dOnXEf9Q4E1VEvkVxCCRsfcqO4VscIMSAqWdyD432RDXdOfL
FIGUbXVNrnFq9S6SvW1he9cqS21RUN0ao/F+s6/QbXmPFCoAh56XKJQRjlG+
hrsJP56P8xjN2+SQdsaJxkaHbI6FFvsrm5/LQOXvX9hAQgyVCCDhnKtkjgGa
PePGQ+wpftPRykJVXSi8JFfQf9vu6saGM2IHcLHUpPD1LOQeto09GFQ8ouUv
9jXADWfxQJjjbpp70IXhQyGNpMog6z3wZIvWERjJiPQ900qMyNi5IZAL7UFo
nmmvZfWZ6+hH8//lcJSl5kBNqyxVxspgIZ7AclTUVgGq8NGsZWrec64bMtIs
hKRwSVTLwdM2hFKwPuemw8WdeVwtIkooT3+tPoL2mfn7T1O7cjY/CBVB+q6g
1SajANVa5nT+i3GNzAqeRD//Z/lb9KoDI9U17k/uO9Zwy5Bpx+bWpZTLzVEC
cQUz+K0d0ZzDXcMgRDDNjCfMy60ny0HDb8+VnETDerwAIngoaJzvTiQadfjH
7VWiQzI0kCAYKpppGGhsSAXE6LLipcjMxvG5+EznJVO5gzAo/oCfF0E060/H
XcQnhWNfXAFcuAQgEAudk8yst8mxkvwEEE106YW8hxpmB6ITbN5hFL0aN+iB
6DG7O0m2ii8iitg8r6Pl0m8zK5umFj5qeiAYXN8hVMojH5nb6Nl20/8uTo+L
RH7NyvQTN7Nt1sMNr6ebxBk/Qk/PJeXfEcY15kmeVaWwHvy6A0fRk4fxy/8S
KHoZtAz6euv1UbW6BPuVcOgyzeZ0maJTAuUczDVBOjGTZaCmq6lkwg2bVDqb
xV3lExfyaBXywMSR+kR6fJaBEcgxf0r05HxzzeMj1Zp+UJppoUv6yO2GpYi0
uLouQ7qtRAKjGUnxmtBpvQU6Oiv2PJG+vWe9Z0BPWkCXL4J0NQ7UaUNTOpuE
sanNfZx7oX151z4LlOcY+pf9p6zO91BmSbqCbf5Q4hu7qYOWMSHnXC3MS7Pg
hymcHie2CTsKavEgu2UIHCetQhRDc+F09kwCkFcNK9FRxYn36fUPFtMg2YIc
G/tOot2ErI3FtkkziFHzWqQkJCNHGT0i7+SfKz3w8PLwYmGZQ7IWRuuBe8CQ
XYE2IS79acvgtnj61SjHQ2e+Z5jOZ5dNdHQKnIBNkPPJWQEQEVkdCeVlLJQO
88/jkgMCHq5aqakpWoximce34ohjO4h3ak7a8qVpG66aBTBDY0MVZjzC+tv0
sdf/BxBW/9ExtNb0vLciMscH7sW34EQ2G0PpUpV7AS8jr1FE6CFeToShRWB5
6RSVJQL+XoEmZxETtEktmoiDbdJuIBr9omS0RqHm7VQcUYtCpN0gtNITzMmC
d/2jU+8vS7UpUZpLXXXfczpGekR+JN08zFea0oQNGDWkGVauG/zJovPSx538
/UeGIobeWaqjq2gIdi9RutAAuqKVDN1qgBXyufxikzc0Pab6xg2TeZw+R1a6
xowRbGlkn+3VatFmukZs9hxaczg30f0TUbTW9m6zgT4Pxs1FiMMDFwVgfz5d
nYZdrme3Z8pPognmnbcdiS5IGFYRrmaBvnDD4umssxqF6yIMeDE6dJHhbzGy
YDofBmvJQJoxsCPtzxrZH8tS7MzAT4cYMjV8cnLlJiog0tGGQ4gHFDtIpqr5
QV7asySx0YviF9trKp36xHdOkG5DsyNEIkGNsMFIriJOIUyHOWW2SeEbOM7B
Xf/z6Tq9EtZblQk8qKWmjb+ilwQr2GMFFj4vBdKZ8HHPn8Mm62G7otxDIQyK
T+Q1o2HCrirgr7F6fAIggiCcqeHy5G1EproDLMaxL/X45CuJ0uLUZk3zquIv
bjvePtFNO/0D9RsvTaQ+BqVAV4ZcwLIHeZJmjVa2py8dfiQczDhLHzasGdks
7iIGDSGMU/o9R8NkZIPNDY4m61ycWJPsSOL77QKKTO/8DZtdFp+/yJ8JNxOe
saTxS37Z/jccDYrqOmwcSK1dia7khMhCDqnLaewHKpjZXprIieB/kT5z0dnP
+808E+1Pd6C4tdRAPKPOnlDIK+VqpzQcnSoWJRSfHkWW57HRCSn8LVCNcWGU
LRnKmP+HaIN3opH4VmfPcEPbqckiSKOdrueEcelu42JCmeQlKs3AkM3rIa1x
N6SN/kknv1LFLeYH71OzwHUlOgV6vOMhVzHmETB5XHhzUAZiHP7iS01xv0is
7QiFhFFYc1fxKQ98EJx7tHDqnor9lSL5bym3yN570cWXLNax7w59qB48vU70
1V2/U4pm72zr5dn1dfbda2PgiD4d56LV6UXKlaxbK9kRyygJ5S6xKuKz2iMC
wy5rMqKBqO0zqtzN+kpyoNLiCctkCKS/E6TVdZhVGpu98bXtkQ38plyCeaYG
3pJ3rJ3ka65AtYx1sPD5fVuykVeMIYtsgen2cswwJFViuJ2I95/lJbZIwSUU
/Ad66j1hmr5qokAuy7TWLZFlcKzUoFgk2vtfZ3gdhtVD4VJHp1MAkUYmU8xa
4z9oNDXSfvLFyhn6OKbFppZXvO1AwqppUs7bFpOY5PEZnPP2FFpUQXLSmkfL
DIu6BSv2EHRhs+cuTbc/a7tZE7IvPOsb7dV9ypKcynz/GDFV/sPf8m1ul/KS
Tn8mtLd3kSyjQhaMv0NSDAe2WG97ePDocIhQ4BSJwsnUdTh45sBNoZSM56Re
T/2OCoLBIbgaV9mZKIVvefOMhFYDyLG2a2ZtnuWV5lJpi70plO11CkXIEyaY
CXRjO2bcjWkneD1U2dz3cH0ubWC8i+my3aIvkPkiMJVbyqKiL8UdvvZZW9fG
rBV1aPf7d2GqzrbEczGl6Ya07Fm/qIuNnt48zrqygMfBhsR4/RywQYYPalak
a3F+wsBq+NHOS0cKySF1fdEvADtgCtrZJ5DUkudwBP4jEF4bv/ovzqKDsMm3
5HxK4JTAo9uIbI+/95az4Blo6TqM6cHKjZp2BczxV3GfYe82RkPpbBsrHtkC
81folHUoLOrqvP48wJ0z7SZb+zb8x6P2jehQ9Dmqz4HD9mk2OFMHK0A6ucVU
asuzdf+duhYFkFvbSwiUH1sIAxzXyCqMmYTA14jODgwB4H9x+jK2s/NYxkdl
CXzrw+NWfvXkD0fUcfxgzEg5Ekvcmnmax/pfO00McVygSGKHxfegp0220fV/
MMnKwb3F7WQw4Q0H5u/b4tDEKFc0xMJKGvILgJIW28xcXxd2vD2m5bG+Pbl+
QHKRfpGDNPOjkvkv1dM3YIPnVaTxnqqU0iovlPPRlTNUoPWuqbhaUz3DL9f0
MCQ4YHRG+O5JADihDf474lxuPE0Szbu6Xv+b+MMeZlz6wRQn4xxVLeQy+DrD
vgV6xz4Q3OZ9I56ZUa9Ug3q3SEnIl52uDtpVfkYI2tlj9dY/YoF9ZTzwATxV
kN3xIOkvBD6i/t4+WyjzWt40Le/Hrt/ZyD2MOlYYFZIcoKzfm9HJ+V+Yy/9k
BwT7qHkC8JWgjcnDKkfW7nYgeIOdEhjhwTlIBKfJmdEJ16yOj71IYtF1bcGd
u5eUsfD3UxsfrGMmGShrAeW8VPbWKIQWt6Cax2v0MivivJiFbasN+fLjytjs
B554G9sb6nAJ1rttDLlYCZsO16d88FYmfmxxtdgIpElqR8X2zdo6fks3AsB1
mpJuor8G2AA/PDjqcpKHYCq1hvw+2Z1Y75wwOpIVqKis62BL0qKWT6gMkgv2
wEwQ+eutEUaqP73VlddOw9pxhIXxDFBq5u2G/VE1axyja5cWAkC8x8QN/h1Y
0dhFtF9Uf+7GrxAHtFi2Ljsyv52LapUtclbJWXn0JqMm8rz/GXeFeO0LEhxe
hUIO3nyTUd8BuDUB8M23a9QKYQpn+sOf0zHhxtqd2tUog3b4RRqZsq6ZHLSs
rA2Rrtv/2nbQ2/2MmB7ckP2QqND34/D1yY5dEptE8HgseqopB//2496tsfzH
G0HaQHuuVIRqwJkPMSl0aOSweXj37O4Jo2RVxDBX2gA4yKL2A/aFnRd8ZS5y
m4To/lDYC7qGxyK8myZ6Mm2IRt/EIq0DrE4tvZqL5X0fLxUZz1mPgCqv8E/j
EC+b/JIjvT201KJe9bfXZyZ4estbY/vWN4+4x9t2Q9chgw/VTrD7WLEFSxZj
AcUc6voE2IKmGZbVS4qg016JNsFPfJ28AWf9M/C5LsRP6J7v9rFueUQclFiM
rD4TMySmmW1VsMajrxfaFfBgXByVVDLUcc3MmxwoQ5dkh9rxsllutob4/0Qm
bfL85jXfFY3XqzuRNNOhGR8Khr9u1jklCt6oD8m0mUUg+uOyqxMwTFrNcoXv
3Vd4oRPwHzJ8FvHodQa/okt3kEArb3WFI58xn/OUDk/7m7fRTJNhOVKlFSwr
ivyuE1irQEao2fQpXS8+LjsIlAn0Hs5PS71N9POvlBImfV/gQkdRY3eiJq/2
Dq/t4xW4uFWSzm0mLEj+30gkZhOKXMgXkvhMECgm6Lg85ipxHW4+PGqg286F
MG7QwS3ufaDI9ciSHtVgLpjX0KqN/ty8wq+IEsT/paAkiKtx0km5rtb3f4HE
P4wLjQeIc89vmbAnPGMmd4GMXTBfKi0wdQAfPmlLwjxGZ4y0KxTCZiiDMAKx
A21aybPQ32TMxIQsvN6Lt/khUtRNIc8Y8xY72VEYKZ7awfcUf+yazDNQWCKK
ViZmq+XSTRFdsqavPDr738o8dF13BDXAP5J8t/u43lCShGs13+WKVvb0j6g9
1dRKnSlb4n+0Wvh5A6ZA+TwXzItSd5qIMLmdSMOo+ru0lVSN8hmNCu3S266s
clt+u1dxjjkGlL74825L9glTN/xtD0bWezK0RgW2CMrosfG0cahgduvPqO14
5sQmRWHQTvSY6DC+1zEpznZwdU6Or6zi2ZIduWy/W67YuxEucrikTPqJfR50
eNif3lZMYrfX+AgnhdS7hPb29EuKHztdWx9bd8iPFuLaN1orGxSi9buh0+/2
hS/Gvr3JeBRZ76RGLizkltiAM5dDtxqOx69Dw6Rg5qrjbiNe0vUcrviLcdcs
NqsARcQdV9ot4/TbCztakhMgoox9WHbAmcQ+SAH0wWhLwAto+eDMl8x/ctu/
VjdWLNKhGvY0drd17uyukQPNBXQ1PENuHdk8GRzSFjk/UQVs4jUVHKAk82Fj
IUTQuhYohIm8J/Yl7uXZk95tqpDVbKiQWdxdy3e1pqVRJ8x1p3riwnO8kWqL
oAi4KRt2NaMO466Yjl0DkR1IRBtgD/vTplClxTIQr0ygF8S7/UsOsSuqbJ1E
vSH5G7VRkreBOII99tTb5PExcUotCWGxHHqKIeVPnvlp8AA+FckIHczyP4fL
W0eYUXVocjt9ZM1Rm30OftwdhUHIkgkHeOshzIc14+C8wfLG24eNDYhccaT/
D4HZcPmsZHoE+TqsZQOCE70GMdsX8GxbDzj7rOTeOlLJoQdsaSujUdGIr+i5
lK5o6rRNWcMaSF53y2B8/sVgOOyYQMF8+WgIWzHAATkSn5Y2/o24TuDgnMzl
qXtIEfIUPk3DQn5BY2bkPYevtgexMlxp+seq1ZbzA02W+JUxTB9g9IGhdt2b
xEpwBJkSJmnrNxN7vCToXwg0lyEefiQytTaG76v0/rB0ZoUUs8VNRTbPrxps
2WS+sM/E+592CK7z2pq9XTLoC7duH/8hMvlVb1uB5GB/9VIySeuZm0Lezg6d
jLsviie87wSf8zZDn3JShEm3THnDRiGkbbDlqetoxYq7jqVGZLXyJmUoE3KT
Ya8eex3vYqlBX8BXhiIWc4CboJAhiy6K7lfcOFAzDTOjNSWUulK1Ub0Xx5pY
t7m97yGR/o9F7I6naiudGEuAmuAqqV5lKulJlUuBhUZavuY9J2qVPqsCaMTd
tO2epKqFBEWI84ckJNJowqVoKb4UvrZL1b6Ymu1YE8mBvH5alIqaIq/Mnsq9
vqEsY7U1avXNcSOXkD56WprMVSvkCgn3bIbmhj02Yj+PqqOagpzcXV+yiuhF
3C+f4RjJsBOwLprkan6J4U9iO1PUiJCttVsPzkrMf9vYi0Z7W7acPc1KbZiZ
2qmjM17lcP+5fv2ck4XmeiOAea+3+DVtX4KAXnYJwUROQz+F69ECJ5/Gl6lD
DpEYW48BTDaX965PumykfYAXUv1sqTPFun9nSVN1ihD7UD6unDh1WQs3/dAj
aPTz68O68PhD213AdhGXFHx9cVLgzqvt+2nrLA+PmyH8Jv0o/PG0tLWIkD02
Q9nmELcquM9ctxRmdNuePN76MM8Ax2jWYBWlz6itahRIQeeTAF6FPpD5dQOg
NueS/iWkJ5pPDinWgVNIVR4xMU+mKPrgy8s++JSGZYCjhpls2a6uIhILfVRb
VNK3JYmgIgGpQHC5ENHXoo+MJ0Exn+YtwtzEgwnBVYeNOGON65tRxncexw8r
DC+1Ixn+dBgGCejbBEYTGf5SPqc4qMSZybcl3u7w51YJzu3bOOlYtnK8hued
VcoZPizgd2c1IXwmIa5vvtBC0t67PGtI7+NaZTIk457ms8qHlKxIyPsY/VVT
I60VGQrUNZSjy6FZBvU25Jz1HNV9W2gsSoa4nrf7Sn0yYJI2Jb9ZBA7A2aUn
VPxvUtNUkMwlc23w7NL9B5jdPps+URVtz0Bun/Tgucyb5lctsxaz4H3yiP3n
mufslCzqeUjPwTlp4ysLzKx/n0pYotpnG5gDeB5/Yk9+IBg3S5WvAlEv0XIh
06pFZAzi3dPZgGEinCspQJYfbq2O2xuOxf1rSJBdupGVTymAqOwugzp9Zzdk
3DOnZvDajud1SOUr3OMq3gkeq0Q3K2LW47/7DmuT879f8FuIk4AZ+iZUJCYu
r5LknRg2wnstFX+A8edcYlRtXuGfHZc2l5xq23KLBFix9heK/SBG2Vtcy7ci
Y+YE5bu73RWvwctJQ4NIHcfiwfTmR4TTRbPjAiuO2eWm6iu4mQ4tNCpTwp6w
hQvILzQ7JjlLUVlhtU6QOg4aoGlFHxHgYYOKyxBzZFn5OJl9GJ0SbmxTscaR
cPBSjb9ZHBRpi7y7MEDXubfmt2BI9fFHzV//VLaG7/1I4PbIMp+KPYxQjYDU
3Po2uCZSQ7uB7iOFsqylNMFS+9CwFIkr1m/nQgMxuLSNyeybCBy5Q1x+MXxl
/cbEWrTfu90tpK5QxNON2HHySFHXX8xAwUcD5BeKe6OgnT2jo1l8eDFsha0K
A3Lh77Se1i3RvbaTTH4zz0yjYwMz3y4/ihIlF0A5OxmahfpMzZ13+q2beQy6
TRr9Enm3i0ayX1tm/xi320W40MIHOat/xslyTcRmkZ0r3v/uzH4RiontFpKW
PehSQPp329DB/qhXA6RFY1H+QKCeddZRI5G6dkhuLdBgmtfEuS2XCBog+Ddk
LINe2/bbL5Jo3I3kVYFe4fIbgh+MANgQ6m3c7PwfpV96EGkLHn0v7jhkdmAe
Zz7Akig1XVrA3G3D3xYx5v8ZsUWJAT5ZWs6IGtoo3wA7f/7KVZnH+fc5p6KK
WtmL56yDTTmohzBccHDmuN9l3WZNg7yK

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KKOXqpQh45LpmLPAIwSQSCs0frxy9BjcdR+we8li+S4Zl/xd41uCCGDuD2j5dJOorXl6gafQyUnlFzTBAL1KX3/veMUYtWXgiyth74J7lZw+nMh6/1vmmlfoSarO0Wq/XZQmZaLH3h+m+E//AqYJMcjhbRim6gPaK2vKE3XTNiTcsr0nd9u4gmsbi/6TManGaw/7iBgjsMOBNs89ddF6wGqghox/f5H9ooC7evnuHgYdL8ADUv/7eA8bSa3CXA3Rw4v9/RUjSnUEdb+r/ZXR12wRO8WtJ0PEshzxy58bttOyblsChIYAlszCwm93kpEk/f/hDJCB2JC4OKcgoW+3jdxi/NB4ZdqCOI7DVMdvGltKC36x/sXjn8PnVEhRLagl2zmz4bASg7oJe8NbFvaKDeN/quylRtCM3PyHXm1GFoO4fRIpqc6WcUb6MdllzEq6ZIdp76GL0WjFeifB5SaUSntT5M1FMIYf1RmZqG0qV2Z4gRH+9m4Sem/90tCM5yT7/6Dn4jEGCKC97vvN/JZPT5m0Fk6kVmfaQwQM0CUJySQdS61yM+Klr6CzrnjytSV5CnKAiS5pYilWMheQ4yyTad7Xwu4HINbcRjdEFvRSHesMfOw2200pt9+2IHF7HW6FcZs1nQkJG/gFm2s7+Ez/WyAyRTCwj+3Hw1yy8+r2ASthkPb3Lzr8QDHL7zgZqev7CFxaHD+jsDwqIpUpWJZRdytappjRRAOFK1a8WVCkdE4oFczf49uJDbdSM9iL2PhhvzL3HY2VOCG0TuZy6qqd0K"
`endif