// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
t84O4zFcx/pYSoNzsMBB6PPZXGUaGRkAS4EVN0EaeOpqPELkud8LxrbDa3f6
BjxxahO84dTkJJB7IL4gT/HPU4TAdsyBKbA5krY7PtT/gCnNpVljEARl4nMa
MhDllh3AEf3/enZU4hwGNkUlRSbEgZ02oDfCKsras3f39NT4yU7qDObq6b/4
xxk2H4O8yw7nyWGb5X/cLBZDU/V5viBm6CA3d/LsHIiFC9IxkTS4UaIaK0mB
xqywR96khGOl2hb6xDX4A+VmJ3nmeYrzXTS2L6dVvCmVVKcb4IqkLKDfDO5Y
d8ApAiCr0BaeRksMSdLtgsIu09FDBBMq+YOsXgkdiw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kVkCznmWUfdXQ5wtw1iHHxEFrpfcgf53GctBZ0xXNSy8yIPmgsMq3f0su3uo
eGBeoe688s1VaxKRSf03ys9wq/vBHTUfC1AHu6Pb6ECXIKUegJmJ+RX2/R/i
TcKexJfqFKexx37DcnX4JZOyMDW7oBu3KNmNnyxfuknkxAa8Nmwesv9aEI6I
C4bG61V7ELQ+KKX2PzImvVd+HQsu/6B7VRiNiMBCk7VrTbkjkRccebw9mXDL
C97rfjvDXdDkx4GfnVIDRQUVhFPXPbNT8S42XOVA6/Z+Lij8fxyXC62aFDOK
rLZLq2/qQE69RZtXKN7SxmWFkoAxhZekqUq9xK7tYg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fow5tNWOlxJloF3DEAVpKLhD4XMrhzL28tNBkBkR7KRN3FxTDerg/lLKbcwe
/5dlSBlxv7nSzcSTrH2iIN52qRn1Bdomm9eExjUFzSju4lAnWWyLFkkTb5ne
M2cHu9ZqGTaMlyZI5tmLaSNnbQoyBALrSpB3KGOwXZNzRe5vTmInU8v4ABqB
SzxmcKq3ODNfhj1z9cDry1ANZqSaE7QpyungJP76hVBrQ0ERLN3zFLkV62Nh
uGLKunH1GQjeuuotevT/ERBuc2WlA2bbW2D080ynkcCXGx2t5Ore4x0KYMsy
szVuZZP1Rnst7gkjFwLS++OMLVzbSOOirzYS/HBwvA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nCu8JlI8zT3hLZ3goYolYNzhd9drZrYFpakam38vZpTLK8OcpaPlgLJxubj0
qCYCujBR5KEBRyP3yjpxH3QntQs4nvIdCDCtqzZ3KEuQGZVXXov5oRFkCh1e
bL6PWaRAyumBWRzu7gQfpdUBXEJXFP+O9zESzCjSFLjifoOEhx7oRSG/lqLZ
AT0I0Tz1bs/vQAMG0STbHXOywWRlXJb0E3P0a5s5dAb1fxVyTxPbJlAC1Gmq
3FERzd+RtbolUUgBXoC7YATZQ4odqAkex6W3O23slmFWkiOhO/fZcfeFzU3t
hfO1xUscQqtehYrLYivpATPK/l0weK6vndALJ4B4ew==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PugZPXiybRrOQy+6IhYCvKhwNjRZBxhwKA6MwRrEX0szJfWqg/pKQrMasEdk
t1ZA80SDo89B69YCJINCDw8ZqMBBO3Pys31BfdUg7oun4Aj4dBsNN2YFoiWs
X2L4dEk/ZKHDPBi4opgrnyoe9I9Ksm5nsPE+R92LQ6SlGuB9dg8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
eN+oLMJ6m/Z4Yqbpo2gu7bjc6hOF+Qi7K80jYaK1U4u/h/U/TrFAHMoOx2B4
jru4OX8OrU3um91iQ56tMAl/NpNI0eur54JtBC3wdWba5FOrgz0tSUiEHUH0
STIGzeT83DJgwvrOLggq5WuXTfSM6khOId6x2GzJ/yoHpF/tZfgjzGgQUbLO
DHzy1rDB1Ilaw6uUZJzpEF0RmBcxcHgdm+faJrdxm2gPKocFri04TNIjCMxT
bCJHBuhhvNbLGWKcBtmV/GHKmbDH7ECZgQj/be217Bp/rQX27oZq526aj1EJ
B2k8E8Un1O0QVAT8sdcpBgDJvq8gK/hSAw6455ZlyFZinYsiD8+GoMYiDapn
VF2GDMdF+gWJfG4oDtTh1MaMh8e7i6jh+mXDkYR3gF50R/v9/1urBeaI2Ox7
QPhyXZwDKP+WSgUi2hZeJPBGuUp6axULVraZIoccMVWoVgFgva+3JLVuX6XK
Sn4woPG0ZOzN9P8KZnJE9+zfIPBQP+LQ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cqFaOI/25t1BuhpLlSUx1moIlsU7rs2CECAxXcmzslqBvBGT4+34MGzCLwr1
jD/Qz+kOQAsBtHwwXANy47n43cPnowOE8OT3witvlr8a1tsG8zpyui/F31NU
cGPAH1OGFFv3kDE1L6Ly68uz7xn+mB8V4gDGSIym+lkCm9fGyl0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RbPOrD0OU7zvy52GlU0S5B++HqjVVT/rpe2a9HNsL0EpK85zEo+ydt+G2+re
IUJs5gaDt5DS4AsTf8tl2fBHztIuNXi3KPEFWWdr1nih+97H6gyHVD6/RBgj
CjcUbzCynvPD5+qIxZSee0dGxMWqfuxePxDGJsSAjhSSdsvAFLI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 321680)
`pragma protect data_block
GBlsGNCyagllHd1yL9S98SGNLXKmQpZrDxpIfoNuTvJ1PslqvJwVcyzJhn32
2s5H1aQlAQIeP0cgD3hQnzcu5ih2s1jSuEspQAI2wQ5Kl9AKZRcNRBvKoAHp
eJWJfuX5mZr+5P/OYNmMt6Bvd0TRh5CVfixkoUUgx0bL1qBZdtykI2dSlSHA
dQfXssZGpkYqxA3VeqVkvL+S1j/enArzWztlxIw1DzBAKfh7UYgFS2CkyO10
7kQ6Vik/3mcDbCHcofbI9GRox7Jdby2aqHrHWKQCx58J8JSU0WvT6NOc1rpU
g3IvRL6ABwAExPKDcLQCorOEKqlLVFcQAp7oibfj9gIHAA+AmQaNt3AY60V2
CoX+gbbBZstxEDEbptuh6PaE9T+KmMYtRR/Spz8QLAwxxQttWRgD0MPQPWC9
SRWXOawW1GFyaZL5JiDVtdT8B4cpIipqR9xwyV8HyD+wS969S1qF6OUwdGpD
ZpjMHQCChf1bixzIbQsFXMWxRLhvyz9vZw+uu6vXf8fZyWBMzghr7TVKU88k
xq1BeGmhDORTPGef4PwA9ItalbDmJYRe4iGhgALc9xytfski62oWbGWoKfb5
JwT0KPXl3GNIoRnts0B979+NFonEIsOeR20zqTSbNKQeGjKVVarkEafHM276
2ziCdQA3QGVpUM8yiJpL+qyxj1RlErctPxInA6FgmgSjTdWPYDUBfkXJgHBW
uvX1+vEZv2tpkY0L10G0GxAZ9xs518+ccGoQnvJHBag2sotiVag/A7H8fGEn
CbTF7g+k5DgoCTRKXiUopPPgUE+dnBUw2/cxessVHcsMqhO+aJun7xee0vCJ
A0SCKQNT04Mr8r/QXw/3F8Zwm5+0A3Sjf2vmSS7chdxN7MzdCs9GP3Do4r0R
MKwW2wNqYaQTHb2K7RzTlNVxGM7D3sFKzPGaCyPHF6eIZrOXIagZjrkkpGm7
jx+gyU85WAcVeciikS/enaKXjAhyG6EAP4QUBIvjDU/JM4KamzMZFEwyVu4r
C+Wv046pWa4C9P9nHjp7+Ep+WBgZqufCdrDV6kY3dKZxRa2kXO2YOcBhLjFq
3ExpxCiJYoyBKFGpFlW2Mm942WRWCI94TzCegrr591Yo8Tg5jxBiVDC778Em
ofcpgGaNooMonmHaDeX057r+2EX2SoC3dk3yOeqGdy1XjDMrAZtTsV+ZXHWF
Wk9T15DWZ93BlKE1CaWSotJWb3ijF5duqWfpSdogPnLKqp42Z7JSvdiMBYq6
eGShddrS3IWg9bBQ1tEH5csC86745Is4tziOfSruje+JXZt8E7RzdirXuMvO
uzNYKKeEN6LHjid17lLNYiD+9GbxPxoL2RJtovyxy9D6KaCjaSoX78pr6q3P
aluvpplX/CXJhE2o16/3dqmeaK+6r7TORnB9nZYGwgMocjJDJDlovEFln0sT
VBiWItNWuZj5a6LK+U2KS6fOiW4Y2G/4Kg8gm0O9dbGcXRCjDU1Mb6EXOnIf
VGvmWy+LtCRyA12y4H6L0Y4kOAuRtj6Zbx130nuNSr7MpzsFEdD3LyYpgCCb
BL63gYk/tvO6UHn6MO2IofLsCwk3wN6nnpQusFFrD99uFwF/A5IxJETr1nKR
9nZIe/dcwEaKM2n264xblcn3nwvWzasI3bk3kL4HXKmpS3PyZVEgcuPxE1Ho
+58po2QEox8EFZr20sx+RKKEGj6ru5wCllyo+eSXUhLeCJPa+sqO94EJielP
Ry9Zg6RTpyAhq/DMdoxSlRVKXTehvy0WuIYgVVUtV7EWgJYHtVBi+wuO6JjW
1L0PvcCNOBA68LNqQzxgZ3UrGkev1gnPvMOf0HQP5OLDSEdZAFWSWBBlCX7C
sGVXyNdsQctd1iP1/VchIh7gkRE62tTFOP3QN7pBOThzp4O7GFMrLnVhb/+l
A/omhUBhXmARPMGCcqkIn47F0iWa1z4PdJ0vs78Z9cJxmc5W67vjHsTd889O
k7ibhWinlsIePZxTyMMH1InYXW+FFKwNc6V9/7Lj0BUCTQSnLK6FY4PU2xeo
BCkO1WMjbSwvD8f7CyHvTtRD0BBSPV044yCDdt8QkUbBYiH04qGcv+Jk5MZG
Qg80rjpBs6I10BHffHBZD4LSt4I+NH0Lh1auNquF4hGlcbnA1qVtaL71CmLX
zwydrtQJ47UJOSVa/7EfRqk2EC6/pOMkjW7Fe++2wAEviu6M6pHXpTK6spCQ
3huLD4OBMxNJRRMOwM+3zShOxNbjIgDh7IYaCHiK9CsbaT0H+lW4gQxmJTqk
g6USnPjTZZOx/KjLrSwOoRk2VUPsunfZAt9+MDq7lCob/gl2T6NvjiP+Stk8
hIpk5Ozwo5vZiAvgnKNjbgLQdWS+SHgMnECBqLV18cpS333EA53El91BlZpR
MVvGxsePvOG5hYsASQlkJluMsO2weaz+HPS0jAOmWgdPAsy961asLBD2xhM4
9J+jTa28riEUGNlVhd9f39U/8JI95PdJoqB1jsQ2Yz7baxE1P2eF7Jyg544S
9J8EkiaZpi/qmHskCG1Mdy5aBmKZgPFa8w+ZwAjv7NHPJskuB7gccxtsVYTa
tg0eG2wJU/n+0BErw5WbFB1XUOqlqAmGIwNwkS0qTHyEJTI+VSsWAsmTmZmk
fRMhKM//iPiqYzFx5+mzsHUl+HHVLPsve0A8lCw02dW1G4G+WhRNe7M8dlTQ
dFSUEndt7yJ72/IO82YcrWboHvb976q8TVeCzIbiopI/BjZq24ysn+DGC0eV
5ZE9qwcs9lQyLNEe7VpApcciTJ/jQXNhMw0UdvrRTCGAFZ6y4z62KSdmerU/
VfUeOxf+sIpdoNmsB+w+mQuDuahpfUhTZzlsq9mrr8o0e48VaWtmCLFE4o6I
XG7iJbAIgU9w5YG8BCD3kKgAyuoXUCWp15LUmvnT/dcP1oCoYG1ZTRQbcxDF
HPkUUEwexhRfWCviZKS33Om9gsj/6MzT+MXkgvZtyUmgVp/rcLQ4jzLrRdg8
CP9i/kKzFTW6DixDvWAYkWtKWNs//VtGukPOEqXyA5FHPAw7Cs4xwkzCDVo9
O1p2RHf8GmbV+iL2Y4+4W5jf0qpEMFdfJEx916z9snETPTCB5npKQ6M38yjG
Xncv0oreDK8RvUgVAcq4eoi7BcdO4uhR8J57TJwEx8aBAbJG08Lgu9oDKY1E
rlUN+GURiPJ6qA02evqCygvuK8MvltqbZOsniwRVtkKMnnbZmUcphgS0ByNU
vnEdt3Da/CW35gW5TPDQKLoNDL9aad3/KeWP58f9gjKOYBV4Ktmd9gClZXUS
j7U/roHJ5wFhq45SPHDWLGyUZ8g3q7LMBaabi7CxOnAhCbtFwB7N4HoEDil2
UNTPEXXZkWJZs2r2EFoyH+LR09RWwGd3HWp+0z/+xTJ3feZkuInl6I6pJxmK
/BeKevJlY1mCh3sCQTCYvlNpuv8VmA9EI2X1cn8tcSEMTB1d558/MlNiQYVa
fOWOKscv1/dc367YSaOCH4HgSp7EwFUNIlagmWzAjqcXzngR6OEIrXyz5qng
A+Gs8cuSsaBMxUx6dVMFt+4wAA1RLFlY98+4SAP7AIEBG9u3zHKuCpkCYab2
YtHGDOJ9lwA4CpJ3BL/HupIMs/i3QUGWGjmtG9N+3rwINSFWQhTMkk3djRH9
u2CXmspzWe/PJL6wjfRWQaVGn0yM4hziQSO0KrHALTD/u32ei3UpIro/nVoT
nS9xnmYcY4DdsU7K1Ut84gIPNAILYcU08egrk3EjVi0Jfd4fBQ+EOuGaQ1lU
6AagO9PsWXe7AQDgPpqgf32kpqZP86Au5M32QdczAoNiC/pCRF6MKcAciP3T
V+4LHR8f4MIbef3DbPmU6V25pWmJse010ZwtlUZU9rxzaR7rPLhYDpkBoxHd
6rz6ueJVWo82xIx/5j6Q5SLGxA7fbCZhY4x/ns5UJoVBStJ65I5jVH6SQSXt
POqv5DQ/2lMaG0pPLFY04Hl2jnXLWwQtLiOKibnUOMnYg8UFiDrOtVuWUaSM
/LeAZdFn006hS+WCbUIRjVwlSqnqtJ0+Y/5SF1OFxMYgsRWMHA1oA3uVw+LV
JBHbGEbPpXEx7WcPBn8da3KSJx61taZMBmKRI2jLgL+olxf4rRC6g40pl56r
sdQ89qHACPJk2V45GVbNI9Jvk9x2JxFrmUrwhrlmviu1Xc5tU0H0ErC86Xc8
M2YqJ1Q2EtPz1pGmFarVMDCKsYGCF2STxrjxjGDvgYd+sSgmidSuGrapn4Ip
f25NZwhRlOiI9b3/d2Tu7SFPP7pE2zQATfsAbCUzHVxDxH4pNmkd6kZlsYk5
IOjWyNYY/owsw9scQgX3DnOQvS3h0sAGhKMnfwzIg/AMGgbji0HoGZgHV4Qi
nXejSxlQv24XIsmau1OAEsKcJEhyqDBWPbdTcLFK4urvQZgvanMhDaZqzvxa
hO83Yh/c5DebTmuZ8RS5wu/MDnu/DpcVDGZPwi5Ep8NXzvVDg/N6r5XDqkAu
wY5x28GjSgJ263RfV0tkaG+dLWfa4/R2mHHF11j5krgGnwvf6lCs87/c/ezO
Jn7GUzk4z9l7dzVn1+Y++aRdCQ9S21kCPMQ/YbBrJnSgX3CTwpPAtpmo2mbK
qug/0ZMNFT6gRFPdltKPjHfaWyNAChcM+NnDdESrc+7wCf52X+25u2wfdt/1
8PaT3If3btrWjWFOE3NcqWLXhOi15CNPPaiWlnFtnglo65BVtBKJQxC+HHgw
yR0vSE26VpAgJ9QHqhy3ZLnzGBrDm5yNOm1tNyW+AZcAWlXU6NLe1KrUQjzj
DZHM4gCiZWJrwFJeFc8ZkIc/Vx/Aw/KMBzQJXIuw8ffcwmozQxqikyBRGM/D
bESBzPzB5kCFoC6xcVBtCSLpl3CId4+6gnXvv/u2OAf4d0QIJFkFSixsYL9M
vVQRh8MkKihG7NOiZnpTmjAeDQ4v46bTBFnbxtszWGld8N5P9HXHUqA6813M
Nh2eWg+P+b1biZch4RuZ+yA7c5xKOtTwis8MY2iTO6TW1EfUrUdtC+8oLs3E
Htjt+3r/SkkgIdgFUPbvW7+Y7/kkk2xqfTvAKfnc7xa2l5AFfqfI1r4RJ7Gw
DQT3zU/bT3F7H200SYMH/TFQrHu9SlE+Wqt6ls/PqrdQQd4IuxjyW/2WuZgq
nCnmcFuAunuE9QNR/HPsWO6k8z4QCH49AUrwpUZyacHNvywexp6MOGi/F1pL
2eYzbLDTD4oqz1vNsmyg5WCWvXtABWkKwP8piBTgagM3rzdAlmiillbmm4Sc
kBgpNjmbfxy/jVaLYnxNz9Ecr50X83BheTCagf4bj5cY2ZGrVLAF9tAm7ngc
kc97okDOE2qCafFLplo6dj/Y+vyWHT7TkR3Q4KieehnjS/1Y4xYPqQQzZpnp
u2luDmrgBtNtHDRYUKCwmrjGq0EswK+IMSWKQarY2Sj9ItSGlXH7lB43ZDpG
wSOvqh96i27C1XCj116ErwKFGq7IutTIq4F5Ud7gAl4PYZztkRvdXiNpn3Dr
6rZHPe/IQHm0gutB3VpyR+/dUqk047DmDOzCbkrxi8jBfz67JGfgLxqQSsIQ
PROvRVPoVJ1Vw+q40dTPyUL0b+UDCJJNch2pqVi+3yFZt+K6tg/6djN3ugU4
TWwxeYKIYT/iHRJLXsZ+ju77yx+2SR8hHDIR4/8bTRKwOUYT3Bqd3dCRxoVJ
16w35sPjt+2hBQuawSp+C1+ecjNkA4vgCMMvFVETO1O7hlgrTJ2k0F17IRQh
6cNWSTW3EOtzTFkY0QlwQYGRZ5utpZhJO93pnm7GXRYPVeExxpWHroS+v3ra
ZXJ9RLHO0sPzL01G5HdKcgRWnLqOfNruwYqTBX/B1LTNLntK8p5mCYeMl4Nt
cID7bpm2oBqBfyHSvu7O9CzNvHXSOidCQio6EOY/9OTxi7w7Y+dFr1EHNXiO
n30taM1bgTis1sGfXef5Ty64W804cEIGaziflciSV/oEMuijxgGHtGR6/oVc
eXImxKD4X3D6oXWMulgOGEn0lg0IOngFlBcMhjwr6hZ6g1rEEpb8kS8j+GqM
qFO7sQPCwBdp1L5qMaHGRe8sDLOgHyBm7iT36XPidIKhfENEesDYEQE+1OVy
ojMvoXFG4b2SbxDCzPTcI4b1YBymkUP9R+NyxT4Km9iB6cnlhZIyeYDhsz8Q
OChYAPqQjpk5PkSRGyCOrEZq0KPS8lpTJYzC6AWyrwZxWb9rDVCIcw62MP01
gdusROd/DHka8OCvHJofLc/zcckRxwQeVvNZAZIx/IeLxQmRHiLC8YVNt/hA
cSOWsWrHEfTodzWcHZIruvfGBietsAM56y7oHmU7iJjlPYP4xfDtVlUTTvEh
z89xvjBMCUSZBFsXra/+vr0dq1YTjQBBukBXlG+7WIT6mnwldqeyU/0+sfSA
SCzIA0GTCQr0TGvOVMV//+UzVbVgEyGDXI2gQlDoED3V5bof7nRYPccZJ8z/
YciR3/vBZKA5eulrignv4joBZ1kfAutGcnGkxSXp0IWtGCAqeGg7s+NPhz6p
0FB8++eliISa06e7fXVHzhqXfiLrGJFANMN7Gchnse7esYbJ8O7qmArZ8C3j
AcVmUi/BXDZn33mqTvEJAuV99UxGsQGQQ/YCrQ0CobzIr8GfrUa1yQrZdZhr
C9lvM2Zn0l08OCwPxsJqkdWPIyDiuNHD86pLi5zDi+MgvgElWuFU6F+WR+Jf
lREpbr03ap1+DgrxEUoWmgUdSEwU90KgJfSl61xXLyjdeEHeYNKy4Ko26cNO
rRvr3AJtGqwXFALRbQz7VP0MHlTtW3IhwQFxXOQARagOcTKHIhoLLWy3GtqJ
X8j7zSBwMVM2FWx+ym2ykPo5bhkZ4qfAu15b85E/uCe0chK3Tx1L9Cqemu1A
mwCg4Jl+AsCdqGeS1uUiCVP+O8gyjDkhKxn7lV0E6c6y7etSETfYlua6x+iQ
HEYzTvMg0wtgdQsS+OuPmspdarc4NdLKZErRMIUDyGXieLOTU4KAyt0oly2Q
boYv6Z0yMDBUzs8bqMn3DQk1BP76mgqEnpqvXqG3sVe2LIhHuo8svkAmA47e
+Nl/FaakAkUgWird9A6et9R6r/UNRZiR4gFeGyc7rOCSZf4flK11Hca2Ue4f
DjLLurhvjMwyyiqqqAqk7jTNWkw7EC+3t2yGCrNP7XB0Y0ZgkiSTiIShC5Fg
xDEsI6oLaSsHPJKg+mrljGrNvnmeyAeWxUqPWLO677Kqe4LYsw/R2Pr8RXi9
bn3se2HrMI7qOm9JXbhYX3rUatFqT8qWE4OoEuhgQaL9ftu6EtUSIEXA0s6f
gOT9hU/CjAIwIdFN4f/oOxdni95yjZY4p7X9CWXEKu/zMqc0hKaG7rWCFHgD
HkONatLBxUL7xXCdNwVsKHhVt7pMMAvoKWLEUsNCOEigGGq3ScdE89eGp2Sm
xcbFnnVgpCvZ9GThxxe2pP6CaovjRGb+wFocg2KOa9krrtKa2VCDBrjrUDZS
qfxIVAFS/mm3eczHByre9X7v6YPEL4hJpG7gGANw1ir6BaoVyhdmld1hC4IB
vLl6g61nwLvEh1qZfuaFl4pkuZprxjPJKqoPiyKZRXcKOG4OMirxGW4Ifjju
JD8/R5WY5IC/Q37Zx/ZhyV13kivNIEinIxKSa+iHgVvn4gBoCACKQ7fjuCBU
WuNwsvf+LAS1cDuvPn6yF1j/Iuq2ZXCcVRs2xEaHkk3Bt/CO1zCUm9TDBD+u
Hu1V/25mZhvv0ppaKjp5wEuHUWp6Gc3SIIiYsSlHdIsgG7P4EnVVqfqEAby+
d/RSXVgGme7tel5bNtyQrGuhRShK4iRqupYWprGn4Cd1VZFPGp/bk0qVWqoI
GPZqweOWg0VRH79gm9va/TBntJXKSPCjUXkzJOb9MC7A+s78jZWh7y2Fo8+E
Ujy2eWeRVSxHf4oxPCljLMLtC5haNfEfYGvN3mvtAQNC9dWHYVKkqBgx+fom
rOATyAujfVGxQifz07uyzOrTZeYnnbrSVBL8DzSCFqu3jqi1I+rDrvPU3r91
goNqNl1VYoeFBMJ6vQtf/ADNyD3eKhUJ3Vmp+tt/9JOH+fgAAGJd72/YVoeW
gMK/2iSQ4Lt0TP7M+97pJCX8+vEX2YfJdZmsjiLRiNNjQ6h3nuATen7rXSI0
FFwtYnZG4PvKVifW1WDto+rlg0LYCZFRtP3IWDFyqIysJ/+mXZc/WC1xEHr0
oynSFWyoSere9vdcVemwCtCQipPm+GVS/OMyWLly1vaT2zBhkpCcEHY8ZbB3
NTG64ee3gP3vUljBRLPLd5ffDGjOkXv8Mt8VKkv7uTrYWmA81hAUde0r1QiZ
iGIqlMRo+RmFBlQJ3tNDwauJ7z78sbfSpqdA+1HhNsiXvxJ+9CAw2xg3jL0g
bPEO/Hv07aQasMiM/fAs3foIC502zgG6iOn4Mz9guXh7p6iDv8JHMTEs/3o6
+PHyvBBlgfXKmaxJOTEqO3lEg0Y+w9Z/Psh94X9Oy6oU2V+CYPlxRQrBJY7f
LC3VC00StxhRlUr4evzY7VhN6sevdBVzixkKkN3PtzzPVDC0lN1A0viyTKk+
Y8ucL3/CrBuDORK+XWMiP1Fd8ZeOmL/jW0VfVkpdGxIq8Hf5wa3kScAQh0gX
zSIAIHinWviOx2PGJPBO4XNHzcS+S1cHX3IaFoZOFtaXW1uy/IanJAtOSEUu
vLqujktj5fNBaVwHUka91D4/JXezJiyyzEUQUK1zCW8fi/WIvpAHRPQ6S8LM
hxjPDJwl6pn4wdbPm0vr62Wg8GGQeZbP3f0CBpTveNknUr7mv41gyQY1f4ca
2y8tW9DMFzj9G8iLyL6PHnugnxsD1bWiLmRqGKbEpABBTJa50d3FLkDD1DD7
L/e0ilQzFXAsT6CRmC8fqNdI2vYpMISJoP5G04gPhV6SkpFm5FqW4zXZBaNR
YaLvChyr/IOFjYjTVTgLtN70ui8/ZZN1XGS78VAYFPx3caaY8KrWdFECN0UW
5CsvSLoJWWRJkODhbUPT+6tivmMXSwKpmcLE6LUttKZ/8tIJF3bJ+Dtut392
16znjb7zekVyhmGfh0m9SMSti0C7stSdt9ENqRs6699gLiJOOF7H4C5tNGzl
+20IHU9zS8tMQvfaK8myh8rUXTGyxJH63MTEOmUqAq5b0A5NrgHARgRL03lL
tU6E8RMlQDBOs4ybi2GQSkwa/BL7H+G1zjQsCSimFJ7xX2dzQyjYuRiK2vAS
tz8TXdUOJfMyUneuCwdehhjOagRA11colQQMjMjYcOusXpgKkhZNWsyhMhzZ
UNRGHiogWN/0jtB3KwecXDLW7JwGUmV2mtiGR/WgWy0EoTEbHYK7FJ5azsSu
pQf0iPPSmV58/ZQCLZlvqaEbhBKncM4xIEYBuzo8JXYKVR0zdWVihOIfyVJd
Rqju38xaIrOIwxN8IZbdOYfr/Wg7BEht5rZHW262ehTUJ2+bq44J83fYB08n
6jPH0IcAkWm1XwVOgiR66Jbv+N0wD7cQQQqqxb39LNGV8sPX2SvG45abrW07
X+JppcTIoRqSTpWaIfWjhtX4Y9/HQ7ulhbyW0mIY9jryYuCwodgRr23F2iDa
NKBse8d4Fj21w9HF982XFGYecR5EbiiOW6R705MBALHkbga3xC1+0c6xEvR7
/jFm8Zb56TXem8XpAYu+0o4b+eCnABRw3cckWzWzONwzJio4OjAUMdLYRWno
mYyr5ZixrWYd5tB7TyaAMA5gSlf9CGY9W6WaGkaRDdAOy4VRiUcUaZS6kvNv
lRp5N14OQOQMSsJxErOMwxeyVm6yMTdk2SOqEEbzlG+uY5GLuzRkbEkJRyiF
CIYTTwBs8VMxAAEmvwE47hpwW4wH+Wn1V33WCaK6IJAqF4BKxyACM/T2jC6P
Cdy6vm5wVBE5RCDYrMeQC+XTMO2L4F6XtyiyB57/gpL3/FJ8q9QACxlJFLCd
1vHr4vtK3lRQRNkG32+x8I1oQd5zDrumtJ9c/dOGtFxylZrhzDLyMVzNC5hz
HSYfjFILVyvFJYf9Ujme5e9bUoQ1NVKN9kTph2yb9jTuhoJnH4KMNVUNbua7
sGz3jRYH/Ha0DsmWdP5PatPaUr9XHvEroXct2fAFw+vsTbzl3cbbtFdwvXd6
rmmkxTBhorbMeOB3KEhtnU2jAqzMlwRk9YlVBu/gdkU/jvxu2bRGtbMGMP2z
G0SiJMMXtcK9XfzQcfeosQPM26W4q7ihLtU4oPKuPKVKnAMVT+6yq1Qkn3qf
SY1FhxKX6xECMOKCl9Ai5mbStVeGSDZcpf7gvgla8TxARkcSf6q0ItuGkKHt
RUuAn9dacgx9iHLUrShutslQwhe1RIk6YD9/2xM5sc/E2wy2/u+gK1iQirPF
gwP9MvsKAfyL38j65lvtgBjXoL/OghmVHM405pOSWldMkTk6qnsr3kuVs5UE
7ISJSXUH/iL8aMi+A5l02aQqtf2kTGOkxd5Y4t7QrvaEFJBVwaXlVRq/Zu/u
ZPi2FGIykVkr6h8KLd0EGEkPCD0QOJz3bDXb9iglKgntg1eT6o2iOg0mLChH
B3uJC9lf2ZzE3ctVSsoczWq8GHhnG1djP2e2OqKOqWsQvI6qsnofaX6txTh2
Z8/Y0K2h5gI/p8dG+kTHifAXhqidw9FhNOcsb6cPYnkIibIfrNiHTfRLJKnK
nUkvMpiqiK1DGIE2LrJw7nmGWmz82gYq3GeVhHzpxsMkGfBbPWi+C7RQeOIs
O95toECks905gOTod1eD6x9ylUAQ4Kyo2P/nihzk+rpqXZpU92Du4RDNTqqV
qvKz9yMpLL3dliv0V/OBbTSha25uJNVnNeuo+CFObIj0fCBVuwNGNTd8AxSR
oQEj4Fd6mKD/CFleW5gWzFjdW8/Ib00ZU9sJx9q9LLiTxb84XCiZoFKLjdbV
AkMrc+3EbtT20TptcRhrAidbFSATle0R/zyAprlhSbHOVG1gucLIRKeKY99O
a+HM/C+k/v7vhK8Opzq/PvA9f6TBXv32vHEanyXvduX0oUBj8N8wR1V/1Qfc
OwqOmjtEOVgw8mQ/cId7sGUMSt7zIS5KfZAbpDYILIJzuk+7Uf8W1LvWG7Tj
X8/PeaZyB/N8uV1I1C3x57apufuodUl54oUOvTt+IPvfz1Y0UvCEV2cHjiHv
Mn4SFFIB4tmnD2AuHp4sZ0hvRu44w34ca7Me8VCiNUsNKCJf3kyYUfdPdLQN
+Tii5i7+M4L2wYD1zd2mZK2hN1tidiVNw6XdIAoYaD3xB5tw5B4iRR+fePFF
/WufxR59ijh3NgNLjtGnTuZ1TdHeUaR2sLHWSKH1X3gyNV09ZqIjcLgnCDCE
KS612GZs0DlzN8qwsweuDwkreJxjdSmloeKXBM+uYrjKcdEhzoQVqeLOivcd
osISJAk/zoPtldm565qDEaV4TKhkIdE/EA7DcEnPhO9lwFId6Xc8rsWRgE+X
MKBELQvGwXSpuYDVU+XZLhTORFkddJnAiHH2GF87U9eaZNMl+qNdkldz+O2X
GCUaV3ghVG6azeCM1RIhz5mMQQE8Nzsu5zzYXgPr6b2bnYSOznnDyMVBvVK8
n6Zbjr7+ac75KV52lW9cngmdVGE4Yz3aYkxQZQ4H+szP7V+Z/Ks+zkfX+pUM
SKkJqD7zrDHOQkDc17Q4mtXJvro91fPCBKM5cO4K6TZlcSnqJHMkIuRbOn9/
FDrH/sBRkfPye70ATpdWOUO2+gKTqG/Fp/bg7aY+OxMIg6WRCQdycn9gz4vf
B74+kwUP38wgRzU9GwFwCFmLz9bGlRu6+Y+uIIKOmzp/0+wklxFp5kVc/iOx
WrwmYNJtogqozlyXel33A2uWKY8TNeZUGL4RFY3mSAkjHX5tem2KzwbkzIje
VWoeS69ZVeHtz+Zn9lS3dMRskfLZ9m1GS1uOUii8O9wcEmXGqZrRMRLKQoZt
bTSoAio97vl/vWZpCL9D5xNAlGMX2JLAmyjcfVLoKtAnos292DIyhgkyDjCY
sIfSVjmlxwGQGNAYWbWglvey5vlyGbmM9zqaaIieVi01xOLhMaS8ZKXtPdo0
PA66mSpqiaDgRmAp3tdQHhluOhIOvptiu6gi8zLDLE+yZRfXGXCEqi0t/AsA
GQrX/tSoZ2bO3HgjsN+Iw+8gHBQ/sii1l+t+XfKmvyZBhBtFpkglXCAbFzyT
Fdtdnm0Ek9TLBy/NzJd+N9ZUM4wc0ZFkIWNMj/l8ZFTP3yPzCfSGhY/z4oT/
Am0KRKs+MDarPVELDwNDyQdcne2ezCj3WuUe7U9qyTlua2rsow/Uh+1qbaNP
nv0Wj6T1s+VYBZHLr8/2g+VLk4Tq3hrcg2yq3H4Mh568EhdKsuzGnFN0xSiD
9+h19S/M5+Cm4uR1kAGDAMkcVuOtl2J8pl+kAk/QR/lx89xcSfrBqfTuyRia
DGf2wz7sGyOdG+xlX5obkcB50ekeMZtLuHBeBQspCmLAaRL00dvqVfcJb9CC
KuKzMdtqX1S34vtjBFiPBAla0mpZrkqva4iBgDM0x0ScAWFTi+VNB7Y2MXAv
YW1FR46I4TntWM4e9W+/FDdtbf1DanXpj8HlL4Nbje0+yvZlCe+eRbvdGh5Z
Jruo4iPqzca/+JM8NotJ44iksh7IeKMN5q8u6/5IerlPaCuDdDIDax5cgCP+
KPQ4ylGlmTMQvk9eS6hkzbkeX9xHwpp4HkIosKimOCiAAOctriuHpwAPyxaJ
TNwiZpUDG1zcAjoBF/EUGisQ45fGhOsLW9cW8ETIYF3exRhyZnN1Y1YaoacV
di/AKQwGHVSeHaUMAMbrHB9hUMxc/krvzF1Iuxhn18yfI0DC5+KyUKvY9suQ
JpvE3/ThToqJVh5unDIHOfkV3GlNGx745cdnhHzD9oTDJ0Xx5zYB3K2QLllL
ZsLkhHpTgFXpSb1saTB93HtRWhMgNYmPATEc0woIK7I/GG9+vF2+Fq2EZgWV
nPc/aBSreqZMNEUMMGpW1y8JXdwe7orqjoDbL1cp1mtbooIfWs8b511jo6F4
5TpYAqjYqzpkZZkU2R1tvqVUiqWwJs2zhZBJ1ZlufVZJNGjOP2dU+vJU6x40
p/rUUAWoPQqaLk5x6rjECGWbbvhQJKR2gs12XEWo304dN8IzpVfjbATSpY/d
yxjxhmRL+VEZoJZHBmEhVhPnLlFkzWMwHamHnJVlyuFq+YgNkNOwarfF/XF/
fag8RR6BfA5lPB/rPvHryf+NVHgwYZbjNn62wv7gpNyKo62zsLd64VArguzz
Xd3/YncBv+Q1I1oiwClwFFpKnvLjBpRLJvgkhm1/D7lWd8LUTkdNVu5Vu1MS
3JHDRSetGDrAg4hQ3DMPD9lzuA+9BugVNPOYDQNewtiIj+yrK9b4c5LSOnqp
SmAsq6yTJUgOfjdQhFupFUvS6mT9sgJQlep83u9PW7g0qFFHA5wtUj6oUTgf
QQypkaEwSDPbCmwvPfKAShykCmLi99aw3FGBYuL2AlI876vJxDhhB8XuWSly
I2iyJUv2yLrE5PC9wyxFUdJAqNJDurcOuEb810KpPAFHfJE7zBjHiIGzLIwx
XTl0x07avlSygfjBduUTdQPePs09S1biStrjlAvKUzI8+B4pHAfBJMWK6PCs
OK2L+S5xCj0po46bBreqqaQjKRvp+jLC7j324FGTn3mbarylpgjvG/DfIWmm
91J7ukJqi2LaVz5AGdtXxA0d7nbfHM6nPxysAAhRh5SXXlOM2lIFvD5W54Xp
cbjE6XK1an+CqUYIIBevytPPPangl5HV1sOljmEDt2264/OpETtF8MeIlEg2
m/GpVwLKf64/Tv67kRqzpgFlOg8c7y7ChS+7sTNxGT5DaLvDntxIPYB+lHR9
dFyahTDToz7SxBlvDXN65eAi6xmHyquS6zQbU5xoCdlgefcJd7XXE6PpRuhs
lWSc7wkylSfDJ6bjIQqT1506HKYlDE3zzCTfd5IdhVvXwc5azNwWRK1M7b1W
uR5YcxGz7t/DM2PdXO9mXBYExx1ObaaruXaRYKBZUL3zfh2yr6RNDoP0kp5u
FYCrvly3K3qerv+ymKrWi9yS5NulwWvS5xXHDBZy5rvQTlGBrgSB4CmEUiVz
9yE+8KrCei2d5G6fAYurSj71OwXhm8nFMjVG4X14Sw9A+0RfR0aBrK7ypO/L
HjNLBd/MT8Val42sWvszwKs0mMGNGPawktmnkMy9tsC9L1TSzb0x8bupPCtp
uAtjv0AYcmD4Aj1CNLlmddnoRqNRupWqqAhQ47dutbgRQOgJYDEOMDbReWwz
UVs4bMpKR/kVoWuWk504A+/E/hUKnycuvifwxACBWx5rFOBoICM45LF9jopJ
TA1tYoZHhkCa9EtenzEPnOll9AlnPAGJIQdhP2gK0qBP+SU2g0qbN7qJuQiy
FB3p5ZWMCeNBcCojip1p+bfATBUYyB92Kfx+aSP2hnjQ6ZXL10IZQgc1UZVu
/MXH88cMXTo7MXmHQWg20E/Dr6B/KnfkDOjOw6sBmb3/7R7dLIFwIanXPhaa
ZoD8z46aio9pO/Kne+dP8wZjmaN6hl/QtQoNNKjhh5X9egNlI/LVQ00vsCM9
xRrNP2QJjMpd5TAzFW+R0vrf7zUec2wR/5qi85sh9TluAcwJmdJDfoCCRNpp
8AAt7VmFATaXRV5pgMo6NqFghPmljssR23jg+Hayxe2b9mgnh69FR84Qosw2
8bCcgIj9LQ0tS/nmpvKfwXhyt1RgU92X6jh3iS5NuI9zs+wXUB25io3GoS8R
fQoIhiYiWvhg9rj2eV3Y4bPmxnqyL/YHR7wwclbwmvDkzQSkGMUcpyABePi3
yhtNgz3PhWUTehkCTvM8pkc93kvHaZqgVYHmgXJLzLg73GtaPVJWCbM0hnJb
mH6ApyYf+NmocCPLqwIlPylKyWpE514ff+Up6Z7qMWnfsEWFT6Qe3hZNo7Zl
psZ5n3GF8ufaQ/mbdJzgzQgL/L5Up4lOWyQufWpm8u71x9kINbvtxKEC8lsA
JfrwUQRiJ/lWv3MYP7dp3j5frazJ3WAimnK+XfhcJrUz6A64b2D6h3OqnyiL
36YLxXTr4hXhNG8+WlzJpVYLkEmgZrfSWdgc/dnM1Ex26JJJQKYhLkbvx+Cg
nvfkzdMdmbliY58BCW281ZOG5P2eadhQcBeWdp8iPg5IZC/aZDW6SUHBJ3a7
peS8KK65AyDDpV0i+FLgEWO9Mp81jPkhFj1BOsV9TnbTXLdO+YPrTyjSbChr
+wwbZK2buAWspVr3uHf1j9wpw++WAMcmbqhvAqMB5fgQYmc1SM5QwedjBLA1
6KRb7c2QkqmcnYVMWHuIgdWeA1nrkJUeGVOCO0/z65PSWt0GQQnRhoVrhb3q
eG+baQyu1QclLTqQdpjGM5p/QG8IsSmpTIlkIKMS1AwubqEMIBdlGYeP64m8
y0AOqolETgMPXy60ny9Ca4jq6qUTaQ/Tcw9my53k+eX4VonNDBCQElh9zm1f
SHvauchqbXmJcL+IZwJDG9ynvSmIg1xnRnCGQ4AL+tHG1IC+vKOBUXaP50vX
i3xGym/9mlbmd24ufiJn5xuQGk5rZ5t0bncMkVn4UiMCiR3PJbhmCD7w7hoy
jNqToYhhh08qWNfTUwcUYFT3r37kN8+HycjU2/hnV+5T8M+gjm5hNRz/BXi/
qS8MHdhPOZG9CLo/BNpPoy02Wos8Cslkj1vKTQmwCqonXawIkdlZYvJNVDJ+
ZqK5al4kPVBQtc+LUL9znlng/bjMRkGgzBfBH1hY8iHeg2ydTzvnKXeXN1Rc
2AN3/P+UcMnnmIJoN2fkLfbJ9ymEoRVDPewSlVbSSGqzEDIFNRaHEopr1Mkw
dSozS2aIn1rEkXwOdZCFooAgqoNYO/HKL5jNFE08Xr/1zJDMFxUauL+ATrjr
ePyodBlF6AEd4C9t/oeRnh0wqEWDdGIGt5JawiRK2KOoEenQEQEWD1MthdIQ
wAdMRpSs8a+xIw2PIneQQ/xEp9TQ9qy4Db4lCn0EN8RkItTBu37BAJVqF+g6
TzWlVV60A4Y0WoUwciVcXC1U3yOZN6z7tIRXRUjG6gTcA46rPmlfFQfMnukL
3Udy973NBg2l/ek9uDhzbDYIqJwVdLmmOYISu5eAKJL4BUTxa/ulHnr8NEcE
bBZiywky/vYlPo57vEFVH2ukJcfQ+31FhzoRyoQFsFL9LfxK1PAA4uKuQdzL
dN5/UWuf0OsqWM5JdU2E0K7M/kidKtL52zYfTlvtW/er2ibQK/Fzc2gnTzBy
v1vRipy06YvHLT7Zr94wVZoPAYxo/iExhlmpltEJHRqFOgUMbForPZrBaxxC
X+uELWk2kTR3Tx7ZgfYA1MKDHlFUu9ipWW0CpWaylGAvJISVqTd/4pfaEmBo
XPbv7bBWlErWjXRAaNU94/b4VXKBkb460oKd86xZigLCV94SuNzQX8XB4FyS
7n6BqzkBZcsRkGEV6gRMGzgHJxhFJDaWQPu3UkI8cWAtu8Q5NRDEx+28icDb
u8XyO9M1i2PNzVnTVapdHEEj8Vj2H0BNLLjK2zHeEOIxco7oohPzJhICPNHM
JfSepLd0OG+A5vozIZvrWT3Qfc9QwxO7RZd/WqWO4zyHCCjrX2m/lzm2A9F1
WW7A7lHPJu9osbwPs0m0GbA2qTOxuLvrgtOMCMS1W2QxD636KpaJt5aRB4Bi
QQeGCP/wpRyqjSxkYsyvOrbGlEMshHzg8oW3EaVrnOSrX7vw97ifPvL3XO6D
xpBGNtOtPCEgQTpRdpMVSnIq8o9NiZvaqKnBHWgwtJao0ZQgrDxr8fEi/88w
ipz66U2l2hX2vsnskgsAfaMq0F+75x6/ha0Du7XstTQOaozPqvWxIWk0MWLg
Sp3MUUl2RBAkPFa1czHo76EAKMynnGI+1bzy0kl8m8Nz8yLOhCYaZeJBTK1j
+hAyrDKRE2DWFm6UUv1KFQ3pzoWzz/zCuKBqUIZgbEMy2o/aUlvhuk76xLQK
LQS88Ed8ce+NCj1DVYFGVxaj3uLfkFY7RHRbWJlYDp+S7k3rvrGmPje2nhg4
GITIXRDJ5/9AJ7lGdnVLyDFazBEko8lA4ovGHkHUG+KraNQeZviRW/o9CA1i
kgYcIYgMBpRlfN5ZOKBLO88VMH27RXznuMIY6ff6phzmesFwCwBB9K3591ek
OacUiZkncNBWZxmW+ELOFGMbmxBKZfeGKAkh7MWSY3GFqWDu/gtScZwJoAd+
BrPfpHnVdWSIVWPapEmkMp/Yaf38He2QGwD+1KL6rSznl5w+2RNJ1u/iH7uz
3hcedE+Uu4I1ZcLtk9rnvGPhMyrHtpTRsUSn6l+b+YjfgC8f3MCVe/HLZMjm
3k7XB+lGj+tC8r608yYMM6SHCb7UPlMFo/lb82g2bjxBBNzqm+thNRP7g+np
zTAklKhPUu9jdjBHFulD2mLzGv2x0x+egPDXOAu+fbEzmfElgKULX857ULs4
NGGkv8+Okv2tGo3R2CNyO7bfPmghUw0o1U77WQBzHUWWNZEkGUYHnmuW237O
3TcY7csn+QLt5OKTqXv5Qdb30W2xtKslGGfE6uEZxZvxB1BnPRylhl41wpHh
/rQRkDepd7D1FGM5L1ZG+FZgUIzmE3vCVNX1/TfrbcOMW58Nh03IWfwzt0yZ
Rv9ETX+7Uimhan2dvXjcHw4oEU2tFKoVrObP7CuqCp+n668gR/PbWXERhq8H
U90CpB+QymGr5JKN3YYQH6JrmEOpmx6CWnK1uwXUvMVop2HHwIsrJMsxcSCB
U8bB6un79YBCcR3X7YIFOouqMbBRwaH3V8u1hWVkmbmzaiFkAb3rVSDzRgGS
dTBmhHy87k96W/zmHowb2BjAQN0BsVHjBWDGoXxGzB8FO17ojM3gNX4JjDSp
zlDIg/OBQwHvK4Wsd6HZcb/PN24GKQCCmVzQU82efRXBGapdh5wooF53JRPS
fHQGkzQudF4BXUBPQRCm86wTibVMMcBFkmaSfhv9Smfdzi8IZaikm7eWbGe9
liH5j0lRgRAJ4Oo+HuvF25NHtnLzrIkCMawWl49WvXT4o1hySklY7RoeDmjs
+XY+hAam2K7f/Golb5N+BZtzW//SB/4UxcqayV6Ce0okxChyD20fq0dm0FJB
zMd33rdHDPR/mA+5IgNBREoNh9V5gPrn5Ann2LjBJKUr69w2IcfJV6tBw5Ow
dCZ9ps2KcLb0NveFT4gHH7FuD6lpeGZyGZHrf2viwPxQmuEz3Kf9RhU15Qlu
tziI2CYB1skhHLH4bD0ItPaTcsqHc2cxHgTWqvCz3Upk4c5CgzLmxyIfgvTJ
rsBUpyUTWqlfANgZZ2yA3+8XVjB53BURCwgpAtKWgfmY+0i+E9VcDsxPb1lX
RkDBSk09nTwObTwjp+3yj1lAwKUNRKNodjJtDa6qayoSlnoHOKcT/oWp/S9E
UuvEejAV5o5bIjKwhDGl3sqq5DdK/aLVzwvj+7qEEi9FWQUd4sdkDTwTsIV9
+gKJUOoowTdGtdZRtY+Etgl9mmV0WEC9HNQ2JlTPv3kdORgJ0tPsUtDwGK3l
BGR/IUorx1wpDWskrN5z0rAuJKCdj3RJrTR1gA9+sClU2xPmMwCFGyP9XYxD
rEmYCtXtG+p2lQpn0LvVeMIqren2RhjL8hlhMzL5TUvrxV089J5l2IA36ksU
SufKgqOGUsJd0+LjuSFaMtzxY8F84YDlU8IZca2YizIbLkH+SIhlP6xnDQVJ
Bhh6Z2e8NHCGgmXr+V0zU44MrGsnFsO/JlXaI5YVzUA/lWbpkVgxVqsTzRrl
GbjwYlxyp+SPeRswnsthCvIf48G0vrMRV8uQ/71X2jaQQkPv9MxOK6VHKvdL
FaA+eiLqQoJTE9IrUMfA/zjLtGhSWr2mcx/aGJ+MmJABDJhEy4ZeFLexmY1m
jqSWvbRHLJtXyV/0f8WJ3VroU3ZvwrXjUEg9VbnmVd3TooCotQ7knSPQThXl
tp6a/MEQ2kjUGyJmo6qlPNZ7GkcZCaC6YE6uSqKPm0IW7WNzCzbgeTJFr05m
fNLeS1fhNK9drZ2PecIaB4os7ygrfogefteJu6uPoi2RvTlhonOqGOeE1Hzd
zYUDfp5NcPOfhsL0cFpmSOxuE4UfM8DNuE6PchBoWuooPDoVYSqV8GZQGn/G
cXL57e2hsPHg1Uc9uQvEGbcTcfcojNke0ZEfC0l8qcIawlLXU1SElq5JJAby
2CJUiYd5fja//uY/UWWbs8rfiq7WPlde+3gTwpO8/IO4nMhTdQ5yYImlGDEC
y5h4IxBl6Sy4P1zivQsYdzJdSJ8IPXmAJkDvOPfWWzxP9iL9rPHXguQa5LNk
yAUfQ67jHiYBWVJ8YLGh8iYhz6m9rFlBylLmKK5pTi/88CSwF56Yv1rC4xuF
jByS1AhUEeSWXVNql5Nru/rsKgbNp51AgCWV/0lru9ZxecDOUZgQpT/9WzdU
TOZqU5A+v5ygVH+7wmeII5QL4n/CwILTfuLnct1mKWaFszEe/wFdJE1s/Lqt
FVVzP2JaLy5l4a3zhB5B4IduiTzr4M/sV24wNAGu4y5xjUxUfqYMoes0wjCS
lNT1HXSGpwIn4jtSUvBXdZfMrEnFxW+NTh4OpRg1jxR1K7lgGpfjFV4nGif8
/FkB3up87iF89eXULuyKWBMATTnJVWEBWfU7AJjQplwymaM9aEE0mKcMVkVP
sEurezGE/AgJvXjalgcecoahWyR2gQEncEwOHOTGX069+7TKyBBEG0ERKTwS
WswLDZJu2SxAYjpwEZo+cCopG8a2AID7eKF9ZstTRshtCaz/6fDx7iu4Qgk3
W/waHDD+6KI/2dPraYQ626EoJd+8LkaMru/cZq/sTHdJFqpRR9b/FwbChHoR
cDiWc8sxDAoPv3ejHQqS4E1LUGSs246RpEtrCkdo1X0a1qRPv1vPpiqIy/nA
hr+eBEudtaLvQuz4ZycnzSJX5JJkZEHAKxQUig4cI/dJfHk120kHUFLu71Vy
HvC3FgbPuI2BTxUGeyOw7rfSKY1+DnN9EZrRQrcQTHMSA4xJjmskFmfuREQq
thar9aly2ERXgE/r/Zs/TTRKxMIdyyDSeizo8Vbjau9EnU6JBPSygrPiMWPh
FMytoysLQzOnUoclOPGd12RM29hbaOZ5rDGKA4eECORULCe9fLsMzvRCDXvj
Z0Bd1s1l2uNF/w1TxevFBZDb4iBB6bFWYqpQu/wep8+hA5MLD0+f9TUzFfNN
JgCVm02vQAFFD/qoCDU24gL9DL+bJ5H9aP82BR4beVfDJ9n3d7mfg+MDrjdb
aI8z153pnTc5sZoWApGlF1+NbxX0R9sFTm+OOWg/fMpGb3n7seOcBk65556P
L+Chvofv3JxV7ph5lxPuwSDUf6aEqjZrjEhGO25xd+2pV0Y5k0+Q4doy+ae3
E4Dj+06EoIKSur1fGg38YTE0KM3MxxxwZrv6h4C4DR4tgYL4N+tz1/f/BV+S
w/DxpqPBpWDqaX+m68IxE8h/VIK4wtl08c0wIwAy3u5EwsdGiU3s59y8ebe0
uGtGqFMi09p2sG/42b1wemelChbwH8GQ0iy/f/OFR7wCUpOJCmEfAiEwVRZb
72/JBn2uPRFkwm1J/zXkhEhhdEKm+7qIxA59c7SU+ol2fT/5zXTyoLcAdxRA
no3oXYYoH/GkUPLRMzXL/n3RhH1p1fDkUHi2IS8Wrw+ECiwU31ZQHP2fqpVw
cYfNnTBiBFYRi+HyoPNWU78DKRJsFZ8AmvqccHbrzn3blVap5r92sguDoyC1
wX5zFm4xKzz2/UqwcoXY6mFYxpW3RsSDHu0eiEUmEWVo8ZDvoTMVBIWIQu6V
b0+E8mBRK6RLOlM8/AC1PDlbaAjL9LPS4IYpBrZWp2EFeqfEZL7deVgmp0ay
0tEr+59knZGychVG+6Yec7NHyxq+NKGh/lGdrdb6fOwTbupI+epPCFDZvgkI
9P5ZMHz03xnfBTEFe+Mbu8IVAEzsSbuWbkusqquExVb0Muqvvie8I/0U+Zkb
blo1Dlf/TM3Xi+amGPyXpy21V4B5+8AZYpKr+0A+ADbYQ2SKjl4fzjBsSmvB
DMGCUz3g2SxK66zcEb3HR77Zs4Mm33lfMV1OWIWVM41qyDQny0NF+QOACUQh
+KWbW6g2I6omwKk4L1Y00cdZss+CUlApCQCfkh5JOn7wgmQ6J2GSo/Wntltf
UqG6m3VoPuBgTScbpsGzR9mUoimM+o/XMFQGJ4PeWV10dFpVYb0fy4Tdkv43
/yekUYiBQEFb8toqTvkVBVO33FnbVgTJ9upfi3tScV03UJlEQVVZyen1JYvk
OUpN2ebqzMaCPaqsv+ndCzKOwDuja/RPiWTJH+S2LfSGJOJBfKLW/W1/nkXC
6K+lI6ZoWpLxPYGLF+G0I9NqdeceUoxOz0WpKUg9ywWBp4SW69lHRDpRedWA
mVnaBVGYqHyKn1IdTwSoilv9R+yHo1C2wf1W5v8J/Po3VdjieS874B0nm8Qn
gDhkApiplnxCexkDlYrG08MzffQEz9AC74HhSwhYuFFqRsihvijc/BSYen5F
niULgnu04cmFn+Fl6zeN8ZY22iNPvfPq2UvGFto1670iDWYlbKZdyO811POK
kBTS/HnC1F/E7doxtBTWVQgcUwJJtG/zOQEtY4vifuibJwg6YUreVPIyNt8h
xAsaUp9LtD8ji5YMc5E1NGs14M5tNW5Viv8s1wWbhW75KuVNJfQ8LsuuG7wS
lhduPBy2pcJxeJTufVCJJKm1owAsZvxz9WbImA5pSZ4mMxgxwKGz1rqddIG7
MHvPmTu6EHjdheuUDT/6jAfbs0zGiNPhM/BoAgSwKUfbjs6QVnY9lv4FeTYX
aoj6B8mnGI87vheHgKXGoAI4r7/Xc9Fi3bQZVWk6Y1OvTdpDuyAtL6zFrhvm
cfx9pgzP64TP2Enyc35daGWaNsKUJsO7hd2TiESyKbExNf4YNwX2CfSwzK8W
3nbuuEdMe85mGSVEoRTMDSiBgdxhktEMfq62v1WahkL/xVbGhDMCSHyYBOyi
YOCIFeG9FChqiyt3ffnxvmKk9gkBk6pIPU5R4A69Ypia3lqUdyot7hgM3voO
r1MNv/aln7eyv2fQt3tcOSbDDBSDbB0zgTYYuybZzIUIbUwlElLKfqi1O334
5tMGIqYbT19NKAOu5t/q2Z37ePgr51LxIiUq/usObOqeAVy9Cj25G+M+lqEN
78lVMmwUh2sjOZF3QPExvZ1vlu8Sxlxa/izhHm9fOsBzgJSpIYVPfNRbxAub
40Pu2//NOw39DTqCGYxZA39ltovB9UunwobHrvBfxvIjLikVAzAJ50yCgsr9
hfh0mgUxgqle9gRygxuN23s1Mv3EiMIvAQEY6vHwNAXtL2Fduwl9nw4IizN/
/ldWS+5t8DD9f4lwNwk85P3Hgm4Pp+S8PZioM6cORtiuXg/6OfKRJKSpV12Z
fqGfBLX2sC+Txuh8ySES8u/xtN5y3t+iFb/0I5/1pex3xesK1j+zvDXz5NIJ
2U8eIl2iD6rZPSeL1jM642tKLxsGBxrFeKPJayB41x2wYSq8FwvYQCCVEU8R
h7bGEDy9kTzswCod5n+u9E+AozcTSjsoNM7vc8IZDLr61QGwAR1KAlsqohrT
Fc9OuGf5j4j7D/mgevJHBPaXUtNc+zuU/ubsvhXMYBUsKHeN7xym4e1yd1Wg
+WOErnCWpH+2Yw0elrXyzRBtoA5D7T2pvSRgviwYLKOm8GeSHjg/0/Q8IdPg
Y9ZDr/Bc4JVpgCg+npiYBlD1D2q1GPXKoq6WXXAndprMNFrQf+WqL5q4OLST
uoEb59UyKXCjGC/72SHh7a8Y0NLCup7ZJGf/crWJKBtby008sDZpK9KnTjPa
PZP/yY4AvWAEdgJF5mARPMjKp+qB0GoknjtLPj0yrjmt345j0TsvyAnfPU13
PxefsTs7y/UPLNg9ZE36aFmtGtMJQ/0CX7SoTgelktFR6PlDFEaaRrIOvxPs
Oc5ZdiE6tgSeX680SqbI1kBgob4LVqAdH/RuCjkpavpeORn5HUjKAB7+LaKg
oa5Pg6O5rdkTiwMH2JrCVnZZNhJUfTeCg5gKsY4rD9ooriyGRye57QZFfgei
zL1bBM9qSQr0qkuWM994Y5qFPxVqsieXtSsPljozfGw0cyfeu9ZQFL9QOQMZ
zLIOzqyPu54nn88AHf1r2Nf9UnSsSasp28E+AeAPJcdFeaAQ8SFqposY0/8s
8BPwEVCe+PaK14V+4RabQh2kVdQq2rvUUHnM2duWfdqDv7fzsF9BI8j07Vqh
TVG3q3OFtG/bfWtHFB16nukth7fhpv+irWscJ4dbw7FtlDovOaVP0bYJUlVK
zd1MdKc5xMYnugkxXPE93eKxwK75hlLQnmqGOZxg7Kzw74xbncFcULgmzE+H
EOVDklzXXBZMBZl5utjobSpEtH/oo5Z/rVB7681q3yShq5/X0GaMAxehAv9T
ypWDjICmWyw+D2ecgXhnO1Mn5LtmOQwSRz8ztFW4yST4HOqGHGhabDdI6hWO
WfRkocY4ajIiZtgGDfWCw2nHqrGLB8bvp23tCrNWcbVc6RtLO5ADo8nZUhNO
VUhMLgCiNARFjIGe9F4EtmKSs58OgRVRF0RzRydpWG/hLty8kuVGQFqpRp/+
9a6ZCVb4kV5Qxpf8+ZFV7tcv3T+JEMH9gHECFM+IR15LQig/K/7bufHm8MRw
CddhPdAg85qEMsRTuKHmtRHTyLUQvwMJWlLSK142A5nexFZJyFxIfEArIsd+
pj/ocvr5uNpTK9kXyZrS9zS7uWsw4Ni270g/MtkKMqm5GUKxMsVcpqaNNO5X
RiR1bTGQMg45ZH2UkJFqjg1Fkk+CxlnEkGr/7Ge1/awfPzTxQH/e8VHY1pJY
uuQ8AUhFQ9viJZmluNaxLUpGNrCt+TsRv/xqCeaoC9dXk8EYBu1eozh1g+7Y
2liLXqQMO5RHWFFC7BGc4Lg5QKaQtHOUaz/qtZnJzICZXfifdps7YaaPN8Pt
SQPql4z5HTmqNBtaOEHzyBjxMEBckrVUFUmWzsCCz2d3Hnjt2y4gbCyyYcfF
AXVA7rtHi5k7k2wvwQMl8o37dX1CIv3zSMZKiK4+4Nqkourn6jsY0hEEmaT9
TgW+sU/JJn7eeBytVzb2XrC85i1fxKZm0mULpF4eAkzF+TjgtzDhnZcLo57j
jQ59cZMZxwh4N+PXFo9ApOtKWTn6OqL5gcSk6AdTOu3XJ2/jeBlVN+T6I3+I
B+xjSCTiK3op3glrwQDQdPS78wblbZYZxSi6Abrw4GmkrwxQiuv7QFi61LJT
9Jkk8c0v4JjmCVQxqcsc2A0LRBk98o0Z9uvPGWtnPKxAmEcIk6l718/u7ZKP
GBdSU+cbFqplzBgg3AJCOKt22uKgi/v7AdHuCwgB3oPNieheDiVQyTq2bH/I
8+yuW8PZOtGNyq3o4Mf4+bYYazaV+zSItm6++q+bZhBqYStCo1IXPViQF16y
Ggb8h15f5Tu5xsWgJPsNbaiJV8R/368ru9p7t3IQPk8qUsSkpUqkSzAXRZVV
f9fifV6E5zn1IdzIWI4ynJRaEyMbh+EoAAxtahAXxtyr+jJR8Q8f+rQ9YXnd
5nXPww0YL2rVPJ78QiJV4Qh9rBEFfUXHSB4hIVyB/KrNpYHSMQhLW+esQsll
DDZg8BB05/2DU3NKDJOSi0FqKk8Hohv6TpWKjkx73CD5Y79lEzFuNmQY+/WA
I2ojPtd8mO0HWsJ21tdz9LJDyW9x7YRbzj6En8SSqsAfJi3UGjT0gj5ogcSb
pHQlGPkx3ayUAE8E4mSQ/ZCiwvETk1O8FnTq5bmpI8JYl9qrhb3PXVpQoHdF
C/FformVs414h5LVzKI8hFiznfGqWcjbOMzeEdU/lolg6704fG9gBwyGHnzl
BHAOgLOpnUfxpfHABRcxw6ovoOCDv/nOxRTseLQJIlfCwaJ70ihXc34TDwSA
Li4V4O5994ufC4eEhdBF3FWqLauiT9QcICQmrr7AUb+ebCdxZjGbqZXIompa
rMLHAO9LeUboDU2gYHIyIthi1TR0FsNqFeLREBKTrLOvvGdi3btYKOoY+P8I
iUE1MFubmTjHY/qlZ1jkg6+643wOrBKTGjFE/w+vYEkY5l47jHP3lK/VO0Rz
BTZ9f4WybQlBN58EqSRAIrnPrl8BrcAmT9t1zcX8zlcZnEokUAyQ+FiB5dH6
KXeZo/L/rH1SN6CA8Suj8pm9Rb70GL4TK177AgzIycrx1Fr0JYy4bIpXVdWZ
bNUEgF38lo+UAH7S+5pKc26I4dbeC01d93cubXKPXFw84MXc+Y4j/jyoDbng
wlaErQYN6J57wHnfNNrSccbeHotE16KyBFvEy7opNJbYWCBkiqf9KsVTnJI5
7EAyPY6k0MqkzbzDJP1osG2N1jvT6I+K1pvRYTPCq/DvjuOEHWbbw5swtpvz
+GS1p+GYKYMDH1R463TBdlfD9w9fVS7Cp86RuYGxkp5E1cxjf1ane78qRitv
Rl6LkZJZYvDLU46n3hB24PMq+YIYobwEjsr2gdNaUPPsF2CwpDFcWpBtea/x
M3ewVKKt65KYntNybqTiQhCW8Xk0xSPaI6sV1vT4r3qXEEFoKBGkKO1dvRZp
CbHmBQ5WWYtH4XsOORQAniWChvbBJdQKVX76W1anznrBJCSduzBgkVB+2FKn
xI7Aoz3DeZpfssguy03zc8ses2SemDTZmzJ8aGt5UJgMW/lotcFmxr5stbeg
4Zmb44oYaMR7saDR6t0Lm2NNl4g3iG3WhniDttQQ5BzOvd8ZJZPtus4iYLFV
Flj/iPbpWyZNCF3VWzEB8fvvPdiYBBOVv8C1jldzOZlWUPxDrKQJFNduJ9Ec
LT6hlMBvL4LxeAZeO5SuUsMO6KQ6TOzhH1lj/f1+p9ryxfNTtnF07BgqV9sm
2ARYcpVDHgAtVGjKQ6s8AEghqSKghXKBxrQPSzzxANlBdBV1uPFGPSUpWOlr
Wle2Ucikpn7WO7Z2zx3DZGacVszILQLPSdouz1zmaOxk5t8lF5NP89y6ZtTo
3jBF4ciSl6GdAXqm3o/9SbmcCLVKO009uUu/snF40w5xnzRGP7Zvpq4fITzu
TYzfWwGgiCQJXw/HBjh/03z06yWJ1fwoWCOG9owntFFnHJYq0kaXS2MMN54k
jofY/MZBuXj0H3S8SuAYyjl6gzGU0LNls7tMa2TNf6IMAzVqS1GU16ci7mlU
QMWXLizTmIiKapjcTrC8CK2nb/XnUHDqJstW6PLSyyz6O2oYUosaLjAP2fqN
tOCx6bOx7TJDkoOiclvtsRcYx5azcW4qpF53HttY67bs2PptlwpyPIdiBhfc
Fqdg+hqeXR97iuQ0ho/LCs0ID1IWmc8+tFNVXYcOj9Uvnkqarya26TTrBgyI
n5Xt/bZpfNX64Yrs58PgOGv7wOD5QiksTFeLJsvhg+LyhZPeaTRBVmFNEEoO
S53Jr5WGV/UtZpcfM69miwdi/3RiLWZSdCsIKpXaFp3rIExEXm9Ed03yVWsJ
20r30scxBD3DyzxNiDZJyK4+9VCCIdkFBXspRJzOeJMKTh1Bw/r6St08/UoA
J+V2/k8vI3dhRpE3ZRl7XEc6EGFHND9+PSpOHJbraE9O5I37iyrhzTSB5/ir
+ZQpWBtKDwM/7kr6owO1lHq4+LapmE/scky50chD7WBmVLoHvc2osBdM8Be9
JmUNQc1/tjw+mYTYp05+YrXLPXHZ1m5Ky6TdOtf3zDip37BxsQMPoUbdnBCd
1U030OmG0qGSnhSYEmafVN7p90er/8ZZUTPFCygB/dW4QyjNL4TIWWF7qnLc
bfNNVsEH/RVEQsluGp5ZmuKMurYEHj93nNMcCJ9DRjS8uTyPKczrwPIazRab
Dil0qn6wtHu9wf4+Pgwz8yFTBcEQPm87PAEWhri+RlYzg+uVd741fxpTD1tG
f3Gjr88J+s5OSnJgqYUDsrKuy+VcW2OVyg3fwARjxnbRUmCQwdKxpAxCnUy+
QG3CfktnvszlVgCAYPHUL6MH3nnX6oAL6h8EtHinrBBM4ZmQ/9qIEFBl2bcL
KlfsR6DMIuU+ktBZ+Z1jhvcbpWUJGz4d6QZdcecjuNezQeDyAJYLXi3nLkfa
fYo6gjfGBb4BbdKAfV+p16hhhrd2c9XX399MXJKrzobsYZ06NxEDXUJaIiLB
HNJeU5Z8jkD8F+OWN0CtEHS1tVmBXohPIyBOiZlPgxEGf/BgORLfHAsRNhzo
IOl9aLXXaBHbitH4tja5SeGlCongbahVyb8ltlhMeoN8sBPwoMB7A/ikrpZ5
ENJxmBWA2t4HAvA4o5UKxrESSvJXAGIpod34Ehs6SNU7zX3h4pSXUz2hdP+m
o4WwncVks6atWsbcOfrD7e0rB5+ZXBe0fzFLX3nmU9jMoZoflskyiUKgDCxo
mczEY3rpk3BkfNKd/6ZVAuAuWmXI6Pgxhq/KJlCtNVG4w67q223f3ST5Ilqy
8HgZqbJEQ6j/NjiQqcyAxZildqd+D7DT41IbubCH7GdS9FlCLRdiZpKfh6sC
M9Ns8b3KgDetMyh2+GUOIVcxWw1BIo6QIN2Al/Vmae0oKUWLuWor57Lp6Wz4
yjsQa+Y79e9MLt9z1E0vTPJaYY0n0+V4E+DMlvWt3O+UR3ik9DTXkUIFlCik
VszIalJZgf0dy5P/gNAJk3k0RLgl2yhBMo93VzXwrg0zZpiNvnx1TxOYrx0h
ZXNm2ilriM8rdc1EVvqN/EitjqHGoxlmQ+PUVjNyjRnSaOZ/3FN5xgajQTKq
h7FRGD78O6kNANdthhwyQBLda/KXNMAfFtZIKZh2dEuf9QkxYlZq5ethprp0
WcbwmOLSPsJbeWv5sWKqnNZ1rQv4E/F42GNinzKmgM5qcU6S1trBLguul+nc
ZB4qR8o+nze5UITk12WQDOTh4eJUZv+IVe4d6kLL/iXEZfJmDQyMnMW4nEp+
tYFhDRsjFRT5mv0ROxBwo6zJH6vUDpEX4ZNJVZoJQOIOKKa8xYLIX7cVcKce
+344LAi1NH3RAuT5Z542C3qjmHx8obAqK90ve5iSelHQkmf3c8opM3RwVTBL
RUr2wgQrWcMOkRrdVof4j+H2JUCcDNi9bF++ttkkZw/ReP8lbsijXayrpCaR
CEErRfSi5ma2B/gIeZAzg50hmJDHy7T+TSoy3jorEI9K4oYCwSP7dUiieFc/
Chn4QhVjnza9Wo4zRzZUmcfzIR+k/1gu8W39H3Ksy/IWGvi7yjo+XvGXLFW2
JJzxiwlDyH9Y3lxwd9X/SvOblHQ/Bh1BOnumf182y0m/7XiY6ydL8BUilcc8
V56B/01wGZBzyId21w1u3mmr7Rz8qcniM35ZFWBY5Crj3fdYcSz9wN8jQ2Ya
MsL8nZq3gPLRjS2tJ9nOp6wXlaSx5V3Wti/GdTyCbnbNVXU9G9wj91Vx9AE1
0q7G3TmZFDaJO4IzkDov20p7c6j3EUyyRuPCnG4Ar3A5q9ZfY0RYu8Z4OIdX
Pvn8lSAU+NvYJAQV2BmmnXT33lvKlJT1nmaW9yS5XdgbA2go9aHGYcAoGC32
eUMb3B1auECrg7P7ExIki02r0nf+ItsfPksTRU/Wbd+Iy/UQ2di1J94OIkBi
PCqfNBjI+1Jhg2pXZT8wOu0xi5/LmABHPRDy0elSzQ5No/dFhJkUhAm1kEfI
O+FISDUGclFo76Vm3vKYadwy6PNvWe1WyUOmNLm1uMMgDzSBoBZ4ViA695tL
BUVv/plxSrA4BumPrbPPrKdFp5glB2bQeparNV4ziW9bTHb73DEp93DJePba
4FRfExO74LDOjV2RxUGnZt7zFxoeD4KL5gdaftnMEFFhcqswwsTw1jFDzxFs
CaiRmIFSWXroDtjKnM4bOkVuW6UCYtrhU3D4Driz9VcwmWDe371DqNEnZbHk
MpPzxJ54SEhv9de3np+mVVk0r8lxZGQfpT2EFWavPpTEmjJU99hUqk3hwEC/
hk6Y8ObhNeOgHUlksTOouw10f41Uzlge83h1Lql1zJ4ASjGWV6ERMDfA+FM4
Ua/Ud2Ml8EJ41VasglGUrR2ihbCT948an9blIiQzui/d260oBMclC9LnRR3d
7oR0UF3NLeDHTVFIr5NyTRn+DDuTeCmbjV6Qv3ueMEX9Jg/NvNs3131Xyt62
fm5y6Ogmvn+BRuhOOfAGjPK+YLFdUwhqvQ4NOJ54m68xLSr8uxF9eQDDa9Mv
EKjv0n97zufqwpZg/oXmN3ChnHZYM4jR2FnBDLKbsn5bc37GDD9nV98+hd8p
GGSyaSPCgX5wTubMLLYihkiWW6atZ7b/OfB3NVGJ2jFMaJx6Of2kwTXyNiPM
YK5qFgbSfsvSkC5Wq2vAWHUfEosiYyhLpy9L/AqE1pI/QLy0ixF+uK87ZA5K
78XuN377YqmfOqjsBpk437K2aukbOt00i2vnYJ11wpYsGVBymolgxI9GKVH2
NJx6sgGuUl+KruRWoqJRrVWCRmHO4AOjskc3Vp3RDMD9uJID1w/skKyD2Grs
V7UWIURLQ/iIU1ibrbmtpnvVi/45YgOIjRne3oPIe3ahxM1Fdb4+MeLBVUWP
q4j8/TmaXSLMqHhOnz+cifXGLbTVKU9JQZcGdTTueVy4TV+4lK0l0OxpQ+A+
0uqxZ7XMh4MgtVMIEktlxUE5Ug9hAwi5uNvihfUcla43LU4VR3hPnGWCPll7
lhatMqSIs8BWJ3oTWVmaN6rO8iwyqbcoNJnC8Iarn6/WKMBk6jf54Y4zvmLc
aQgfjofZiMVdHQL1CAUE09NkwvflOxTtbLNZ7gJ11t8vXMBJsfksKodrdz4G
fZmfpPG6lVZ9oF51VIntvvdCy3oxZhteY5z2/20TUoyT8S36BzOoJZo6T2xM
EqNoeqQY/pTXENzHglCqAqmtlROJxFBwPCE0mMK+wLYC6K1ODEgApptrvIjC
J5gzFVYRdZVBO4p041gv/sFg1Af1/yktm7Zdd/b+utUy0F1vquYIe0yB1XC2
bwzI5j57XNI7MHm2S8F5NwTdAYt5H3R4JsWqYbwtC/qeiP4Xz40PmzuGp6w9
7MoUMNn0mrSWrv0fa+2u/JJ9/76jD6VRu8zVMUYHLzRUWwtnqOtihTJfqgNF
zQih+cFw1LxXsbBHLTN6E5WH4zADV2m3pnzj3f2zkd42coaXuSFaIuvGM7OV
qS57w3G0J4IqqWfOiwRxrvIxOt/94Ajq4DF2V8YED2l+uMXDjHW9IP5gKe7n
hbI8Z33r+xU8PbSDtGmKdgrHqTzO1B8pQsIAa3vRyDbjtateOl3XJ9LC8r3D
ZQQsICxbBH09MyPJj9sCbLiPlFh9XxtOSNMO9Im049kAXEkl/rduyWqlVzes
PxNhWksZFQVGnerGw4n73TyQxYecvZLv27CRopssfTKvV38WZ+kLhL43WM6h
EZgkSJm7T2AMz9xYFULkwAXzZJ2oaq6ZpdicBIMvk9c2uCGGs7ouueQvvw1F
FjSjvZk7iDRWW2j00jsb109wdN/x88BjG+oXlVjigFkO8K4MNYMLLHQYmODG
qpiFIwrj6rVjOavZiM8F6C5lWqsMAl9QIYQwLT8VQEF5wRTbEuriHph/ntDk
Al1Z7TNA5ESvzlrv0YxZzcJ8/tZ5bPbIvSzJnQGctlq/4HFkytlSfB0XX+0F
IWmKiy6t1/usXxQ6e6JhGDrN6fip8kfvVRxO9z5Ocj9XuXcBu7fJYqQXVECk
O8Uj4FfzTRd18iXfm8fTUcyAJai5dSRFByCuz/i0zHuma3KkISq6wOyzfVvp
2PRjWS5B04RgsP06RAC9kkhn1yJ/clK9Ao30oqza2ewZtQ5fjYviFSo+3f8m
N2Iv3gm01yrEapR3eOZiS8oPvNIRGkXixBXCcp0Jkbhg95aHRrpmhmxWmrnc
9gcEUa/dXcds3awUvoPnoeHKFidUKLxayQZrc7aQGGX3Obu6KWacuebnC/H3
+b9gR46vhbt5btBoof47g0FAuTSAg5RembVF68EtA0sp4iP3lGqy4ommTbaV
ixIpQ0I4bxjbu22ejc01KAUofXxmAIpWzusdetxpjV/jN1Y1zYes/SIpZ5Rh
V9j/7n7tquMHUCDRq68BO2AUOacEtftaHx/pjV8MbSjo3C6BNJl8QM2faTyT
PRhMExVLAZh1vCLLvzQ/Qii2iq41+ywIRbOM6IRH2tBQmUn3F6XHyheOdqHi
qqlOgI72p/yClFz1xhbVIgFpZWQa9gG6HIbw4w28CC7MuA1BhwNTLQOo1v5o
IbBgNe1+8oCR1Mb2HtikN48orvRrks7T8M+XFsbx9mzaT6jHp9UZ8BdPcdSL
MBPlWmkVeqjzBvQW1Nx4HPcj1iWPLmXArDmTCLdHs5qy/dtVOO6aqQSbJOu1
towhjQW848oDR5n60OU+ArptCDmU8L4YTMP09Jgtsyj0yC7TPKJ2krgEESEn
bZMUV6MVw136P274rFbRSzcMNcSajQ84CG0Ci6qjLDOWm7DH6Bp+DF+eQ+2b
FdEAmdBlHs0+Dys0PtUMG6Bm4zca60gehrUVlq8it6kc00MuZYPFJk02oeu0
CVtW1+1S+HIz8KZUWiT9KsLnns0+QxOiYzUNLIIbqAUPBzt/ImYAru8SrDEi
qe6WWj575ddBGxT3yInie3EgIxyChXJv5eIz1SxTBw+1eRsJ0fUy+Z1HoHff
Bx/uGcQH7Qby0Unh8oUgiTSKw+zUHYoT+pFMnIK7vXPBamslz/doZufixQhQ
gzjsiWL+D/nlKFeDHCeYOt+7GDyK52Q0vcnFjVjBvBb7hHhWv3LPPAMY5fDR
Sa249lDs3z4ytOxqdgwZFKvwFmkGLu+VdhK9GPFtSIFvu2pcOyF6mzxsFUlm
OqzEc8Fq2hpXKIM98juMpAlZUUg4qDfugRbNsmgXxIgZLXYJh22bES/goymV
kupBdEXDEZ9GeVE6zFIfzlQf4cAZoyTdiX6e4ODZKcFMWuZvo/utjF7Hi1RZ
KFLakHvnF1esmV5+DFoGnfuBB1c5GYXK1SmP/T/SCkvI/NL71US80zASENvO
dVC2UWaBHMznhxm9sXLhU7H8DG580zkK0Bv6cI13BbI8CcX7KXEsAm/gyaP6
CIjPqD7iCwFpk1LXj3PWngqwv8GGoF9PqNOna2yjhavaz8gKCgZNh82sJFsE
2r0/F66EykcGwRQhi8tRqiGXHITuwrNmXn/nm+KUZJ5LSjjSAZ14Jsr5mbgT
BQ/v2vVQ+UXfNDOX1eAE5n/sI1xMTrLsI1QIxu1WIe8HhTzm7kbKCyfEt4yw
KGfTNf/ENEL3xds7Wvx1KTW9m9HSknVxv39gcgyveio/zA3IW8a+yzaqHvfI
eTCN9gpqLlIzG6kdIgjtierZvh8hURPL6FgxZrMPQ23x9aMj/iOE3gORVnhK
0XeJol0zip0uPTLnGDxYDbzSx1yIV/j+W+NTW2FNeN7udBA7V3VJwRimSnuW
R4gjOb4I7GxTHZjLBEcFQM0a6060P7YTOT78IvhCRLACCGAcy/FhQ+U/d2SM
9BMFtjAt8TPh1jwijqFbON2dij68oKtQiRYj9qovqxPsgpwlNMxpY0SlzAOt
BgOSbukhLwc88ogq64g4hhL9+/8Rk1RsELpfRs06WGKYyHVe10BBXlY8JRRG
yuSOc06a4YGqCGw8AODgg37mbcT+Cmq17/XDxhGYi5n1MeYrwDoImQlkRjqn
7f8xNRcD7FXr2g5zJgYL+IQEzpQBCYA71N0d7aCdFQc3dujgX+x9r20ZkJ24
PymRkABTcQllOO4tjTgHW/WZ167cXjh2FNFxO0lu5FPZBER56BMrtYpRQ0uz
1yRBCgYi/CVw7oJshlrP3wIv0Jw/1cNYUw98u5US5sf6jmjZEvkC9j2Joy4y
6HBAOmQvVBkOSQxTJktEK9vTht1kYZqjeRLlXfHIwEehAbvdVf3l24RoVCTI
tH9/sJLqc8gYcj/CgND6hZOVbYo1HsN4zFqMUSHAHwoPM74BZC9972b3/PDW
mSpoJSsKeNXe3pAVoJ1yI3VZEiphoMHgJP9xrsn9t8g5H4P6q7F3EG0eEijj
AP9RA3L4QGk7mulSDb8NRZfTTugiEN6IbMnG206LdDA+5DEo7CTWEc4MiTAH
bMp8nFtxL8WevG46XmQgyeaNpmT+ZeDm4MWI5Uer/VsalXADaRv4oYxi3GGK
i6m7JzPamaQd3wFO6SYQyxsiAi0k+6HW93BBJrgsCaRKaeZcv1Cyx6OMQtsi
kUWDhhw/F8PeTnqAi7lVV1nWxEhusvMY5fqH1BqUCzIMfq/dlXMLII3z1EBo
FH86aKsVe6I1bzkhfLUyLaCWQqCBLtdqeDWW/YrR1+l4MzUEYIMuqHYG7ia5
DYmfUwTeP2BjO2KnysYt5SXkvaYG6EqQZSBq3C73AVThrcfdKE0WyjwY0vYj
NigS0OdtGBlCBjw8loUC42xbxW0VakNUSNTGPtoZeO5p7PzJAqw1o96MBMrk
Fxsuv2ksaeNop/dHjzDy4wypn6B/gEQXchoRc5uNFz7cukus3KQ7HOaGZFHD
ZvPCXlZxQQmpQG16rq3Ld7ZtpLfBMzq0gGhHB/xlNPUaAPE/xyQNKoZnRDkt
3prTdRPTaxi515P7jIFPTLGmVpbT1IB9wfSfIoZvIHCZ1OzS2R3DOcZKqNpa
KA2uqM30HrsTt3Zfn5Ncmb9xuaD//zSh5v2c+EI1QTR/OSfHJjAOZyFetOrt
t2u072D2O23cMA4qTc4PGTpRmslN5CIUhgp2x5j9Mb3cQOG0ktOWjufvwYDr
IjP4hPFlQNWxvLHLr3njGXzZN3cpzZIMEsHUqBLtkL+pAqcUmLzMMY9MGA91
8AE/+x/r+P80OePD3FFvWkw1kkdeCjhg8mD2JD9BUGxToA1SM28EAArqeyy8
puOmO6TkBTt/rcYEBRfsVsivWObpqkt4vWaoSt0qnYEYXCAx2Sp3WhZl52ZK
vlA6rkmn720NlR4M9f268wpMgibGDAj3bkTT0x8F1bYT8irfSeS/jB/zRZQ4
kzo2hreO95S6p1phNsnUEFf7USpTLzLgUFbgiUwnBvl12ojgBXlSkX/WW6gb
lB5OxnR5kQELTC5DtD8anW4xTnhE1xi/2cUVfba1cUYauk4OGyZlo0pNmT2C
1Y4cQx0URKSI2fNbpE5SRoy6ICkNH2AgWrDrd9JBUL+B9xJIogRgzIjwPaWj
WgJpNyshsHRA/QmKNrJdmP+pfqlCt6hY9b+AttaKTdIJaT6IIcyUJMsx9bnc
q3Bbk4/5vR88v6qLyexABseqTih/033Ls5dpRG+BZwde2ZRVfgpk8jZV3Xqh
5h2qbw8ov3eFZ4WXE/gGlrnj2QSLPDrOqW+22R2CR9Ld3qUk2TcMj9SmfjxM
SdPj/dwpYNxe6AZopBSp1hGin12spykETDVZGmps+8igrK199qEWkxC+c5wi
IehJ+UEJmGIe3yO9++ncLTDhUG6UEpQh6BzMFPfT5W9Jj+uwWPLG7JGVpy30
FdOUf9waAug1wptM6sPskrBYo2ErER4eMoGbdGpES7zx7P64LzfcMU22J6RW
I1/gldEQyhRLjY3UTQDSJeg75XTI/vhwPlV6LmcAHcu8FXMnw9VCzzpjivFK
dVSzc1fQBbb7Mw/fjxdiim+CTFCle+54la4GNd+3LYUuVu5cy9Ta/Rv9vq0K
AtnUeRTbkxo7jWYVP1D+w9u7vjM5n0ooduffGSBgb9KW0GwNPa9fgEOSimoL
WdbJ8ge6E18QembLEr/6wGYRVva5MiPlk5HNeAQQkULBxC8mop5gbTCTG9my
1fQd69k9a5upiARkCbLkGOXAWAhlvhZVWpJDj2xdevSzlL0kNHMeFhZfNKPv
kXVd5S1T6zedCQk8KnTKCb0E0tl7GD0NIO1/LuxxUfKKQjGuNK0iZ43FSl1O
ZRDsa7WF2qgVePtQODny17CGHJFFWMvzdsQVEPXubK31NLwxMrNT0zG7rV1r
E3pxdZWW3p5gP7hGQmGk6cfGWGzm1y6lUSfp4OQL75mIjLsLau+67uH5Jmmk
tNOuPnU3Ox2fYhmDxJ2Ylh8ZauTFZLX83It4aGjrrpFjdXLTHWBy55ZrDv97
NwZcsZ7EaEF6WA9QPa+m12lzckucEvoPipi9YJgIAOz5TVGTgjMPPQVYikNt
S0wu0BLSP0X5E9fkR3o/JyB4zQ1hTDJoZ4M5c/vd2dQyt5MEjygDLoT+qpz4
QCRRwr11zZrb7BctnKmwDaniuwSPzCpMJrng3OxOwCIOvws5kj46pBXmI6nZ
wu1xrLEK2qlEifSuDs6D4wTYcCPtZ/2Ee6KepEkSOtDd2IoqF0sMebmxAk1U
mesosTvAmHpuNMbLF/8mrM5DuxXss/+s38gt4/riaDJNIfOQyevLc29//+vD
kEbMaum58d4Dwvzg0HoTiglYcfAsNPVLpAr9FeYBHJZNZ9Xz+sAWxK41kTQW
zk5pY8bAwE42sqY1pfCDVC/wcXo0IehDatso/y9lVBwWz3uJzFZlSR3wupt0
Wk7q2OGHAwwm9B6qaia/Y/qORq3JjJmlr6hBcyNR+OTe9BdDNkN3xuuShAWH
ubMiy18ybUsiByNBViqhYpKnvdu7Uwr134tGqlW5+LHHuKMQNPLuKe/pDXsS
z7sBTrCQXtOZsrsixgF64hJJxI/zIgkOvesiwaNVrBFXnvTHEavrhCEhq7u4
hQhUQK1yCcQO/cJD3d9Ric1Vp+b8BynCnzu0x+wg5KIcKETu18qUDeBsUxre
BsKy3XXluNrPqLC6f/VJ1X/ClpjUb5vG5t4OmicPtZXYJiokhGSGDALxPcIp
D697SenRXp0REtoji5SvNW+F2cAuO/cc47UbsIFzAjxo1+avwKoNK/FVTUA2
FIUb0XlztQD4qq8EgKORxo4vA2bB6cawXTwi+Jl5p1hBT5OeTcvhWiEG5gso
LhLWN5GrgZmH8QhPPgx/jPM3c0qXP6pmZt7EC6br0Oh0THLHXVVRPu1k+/SC
Xbwi62pU6qCU+JUpkzu8ljkmJeRl2Oadi4bJ2UeAp6xjG7+jWropKXwwLGxg
DMYLEsJWvlnWFatWr+kkeJiwL60BAEJ+9oCnr6DpqKIjcS8IOjb2EWNB8ccA
isoK5YvojZWC1CVt7EQkjw9WolJ1ChYaN4NbeAFGkNQVZHK4PpSLnrist+1C
XQDvq53hKr9eYCAQT1dOdY7OMV6VBLml4gQt0EtyrJIERzOSaUgWUDBIJDeV
M/s/ixsHE0J6ISw3EweKs0UhJ1OvXBHygcQGtkWOZMuPKrB3QjU9YAe1X/pY
2/tHrBUbins8b7KDmwDm8S4LvDovsYi6JT7O0hPsXWxrU2otxAMK5hGmaZh1
9v9WpQbkYASHzUEztiYXohiCKuau2+tmHV+v//n/RRVbS7zq5jjSy8LftaJk
TTwImKImAdJEXK4gPzYdIg4XFFBKx0nUkvMsblr2bYBsi4RmNWblZnua1Vw5
d7sSOL9Q6XMXhrjhMvZod2rysWila3cAFnOVLQWWNBlkoCPetdY55KzvsCG5
iT8in/ntwGwBmexafE+v1VIoawN8x1H+OPG4pMHjk3HC38qHoX488FaPiVct
5QY3n+wbA4zMUO7/F3+FC/5dy4ZUWYGPVYyzJ337FwfbuCpKtWVgOOlnwTF6
dc9X5q2IJg3VouTepSDleL+q8kv8ofPJrgIgea/3/c4+yEA+ht5D0s/xL+21
EZBCfklEMmEw6t7osNKflglEKbwYaUtFhOPXuMm334PGFmbKC/U8MzKdqv+R
thniXpdqszXl8VA4dPuPo4niYDTXRYTR0ZvwnwvkFaEsBTUFBSwvkN4RTzhk
z1Frt+8ObWA8HnwJRtTojgUU/3XevzYv97IbiJ+yFa5BfisQk1VPwVpOX2Jc
XjfLM9KELGuS/19tL20QDPiLjtyTSZAkVPnyUFmN0I9qZxPl2Atbftfwg5q3
qTVAK6H2PLZlx6/WCofU9B2Q6pccL366EdEGjJ5AovN9GsJ5hr4JO9O11Txh
68iEJ42MahG2kwIOag1h1CibUSJit2vQIadcUrjfLUwA8fmJD+ETNOlZZ8MY
egLaI0k1XLrrFR6BiPxQLowoEaE//UcFdTR8fFdhw3pFBn//kLUMdbFGaFuU
6g4Lk1jm4yo6wiUcP9q933WkenmghxE2u9Eud3Q94uWBCpxKcmUV82CLvnM5
rfB1BX04pbFZAEHkuqi1JiK6V4DBo8Z6er3HpH62+af4cd/2uChviWcHD9d6
AiuzJ/sYJDICLivEGVlS+f4qLJjDUSVKUgv5IgS31FC8qEOouNz5P+jBpBj+
zRLJTbhHPz6uBMp3oqqoHWPKyKDFQuzfmUFzOHHXwBmHgzBwI5gjS5C4TAQG
IVtLjSq8YW76VDPNcRvDIwuSf0EgI0Gq/SP/kUfXFvmc/9T/amu/fl78NItq
sfJJr6vP1xvwFi+TcEZTJ/I8IT14WVHbsRR+Vh4I6Q5Mfir29qxqp671A8wD
Vzq3IWVMKbNuFzm1roVYLKdoStEQ/UaH3SqTpHEEqGm7SdIdfAqyPyeiSrfw
3fje+dMZuWWEAUYeiyJ7TMybdNF+I+WAu+OzhwsbO6rwsqWs6J39Uj7tcx76
daeRMxziHmLwGFZjxcN4PYIDThvG1OIr7njYGmDyrUOQEqRfQXb/9c7lyHQ2
+fgKjSLtr6HppK2c58u/xQHl3WThaWrrbvLDepeh9ssXNYJJkOz3TlV2gG0Z
yBOvRRdBw8n8vbyAr88X7fJRj1jpqqIgRMMHGACPln7E9U1IuysXF+r5oaHE
CKqc+BgVV/1jTG4S8q2Ad2lnbl3JssV4qWMCzwxqn7x3EBebCZfaM/M0uzpK
Zf/XvdeBAn0VT5SLYZb7LX8N/VMWzTEYcAqqmMn5yUZXVAx8OomNiU1S2YHk
wQDk6B6vcblpADjTfZ5JFCrf9AkeWJJwPtK0pud2QmCsZQM9yVOV/M5uUHcQ
hFrjpYTYR5wghbSvA/ROoNPP+yqflqca8LSKRNlY5ku9iCVFSRCIglp3IqjL
PLrLdVa9W1BWMLJiBoVAupwNwy5PtUKZCoBnC8ZOsCPppX7ld41tKUmvoev+
UlfZRypUeyUU07tgN5oIXAwJ4Q7n8d/Fv/bvJjjSA0VZzP/BxyucJVQPfO5z
O4BZEeeO5mcDLfl3v1jQhD1a7a8Sg3Wylrk/32gZcW1192RX+tZ92GoAjcl4
3cCLaEsGc1Z4kIkC0ZJ0cMOGGbEzpp1ruXvSupaS8xeh1Zwrqqpk4eLyogCA
/HdZYy4oOUjDXjFe72dMNBm2ZeSfyi3Txy5fomeZa0bDtKW9WJYtJ5uea3zL
l/OfqLW5l+AXzQILnyMr/rhYLlfvIi5HSKHpVSg2COGKmVfgURZxUv2RRB/f
Y7nJma6M0d10vrb9qsW6h3Ubv0YDO/gIfPMvHsAUYWhgyXDhdBlg0yTJvWbt
FrCw5Qa9mHV9XtK53zXeqnjcGgglsWNWhbscc05G7BFRK/0PI9ibOqK1UT13
MU8emgJ8Ubthau35SB5lWkA5HyoB1upwTWU0KjXW6+F6c4bBMMTaX8jNqjC1
xxTE6rGOK1iXRLenropduz+/27t1+Fk4Tj3oVqpqXKm9+DtPpkNFUmSbCvir
q9evw3nKQUZseuFWBucvu+yDWnZp82e8hbrDI/asdLjTjiSF40UBlDCqRM5y
d/o4ZLcnF+llobDAcyx+Wm9x70Iwx1NAi9qUiX35kpkOnFhIUIbn1hiIKgC2
KrNhdtbNPUnh/BfsnJBwSNGcziUqe/hiF+Zho+VJoW34/2dsGVPb/m49pJPX
lNGwsJa0le/Hx9yP466LnDy8cDI+Md+85p4JmSxgv1rdFFDqUdX0jgbi2kwI
VMXVyyKqN2wynpbilTQrPkmMq1dHGnQBCLdtFkTlRgPXxZJEvJgPy9zEUcPD
K6l19SX+JyKgpQCwTB6m3Reg1CXvcc31Rc1cWDCY+0Z6MUxDZNvYIr5BSS4w
EZ/kKIVk/zJtuxVswf9AL4XwMYgZ3czqk1QdPDtVbLb2+O+ifjheATP1+ydW
dBF1OYpqS86INYwZeYzS8xg1tqBBbwIxE/0peEnFnjso/3EAYotIWWsHmTdQ
hB0BYwiAXDQ22L6hOD7sjnxrcYT9DxlHKEwmWA0GpkG23K/0qu5f0BhUIsbo
zymyRmNI0HcUgFUoAhqu3ph0cjQaul+wCcFoE2XMlJTcDb0pAZfXXwDtWrg+
YG1XzVelmi72vrenqlUytGtwLjdSJud2U/Z5giiHY5IaAOYRTUNuB5m1jn2c
wg1xv1Zi8DPJPyWyneBPvpvlEZzt9T5QYmRETGNEUoSqgKsZhR8ZHHAOl6ND
vQTl+5xREvc2HbhR8FrLJ7fK1nbsGvGZKgF00OO82yiI/Fv/Mmj3eRzMSE3q
yC/AguTgR8K6X7h7by9/g17XHhp3sDhpK8kjseIM9e8424i5fuVN+KAf/Q1/
BNmR6ufsatNo0a+zfzub79bADg0XQGSh+uCga7L4NoukZ4x3pR/yfs/bQyHa
LOhSQElFQ0qvwYhBsjiNZCIeAnJOF5A6ypcor0ndxwJtt9FT8UIb9MSjYtm1
EnADCe3p+R1sg/OD+2CPVhyL5LER2Arl7AIqHmCjwOwbPH2zH49tX/5RIrs6
9OFoIGzpvyj/DpSrSjGr7JB5GBkjXkuTJTeqb7mxmEtLLa40ENS2Xli0RWzy
6wNqLGz1OnQ0gz0o50zwfD9bZV9TGDXcA+V0+ekyj4OND9W97ynCsP81SDZR
DEE3svVZnPfrYV0g39lmrIQL1E1rFZd9puuX2w1gpcRfNogxMqwz08M6tu3x
/8mDiP+DKK48amcWvluS+bZ1U4ZmR4PGg6YFq3azDxaE/40YK8EYaR3qZ9uq
Anp+crmfD648SlmZaqo4j9MQMq6bjk4BuZeZvQk3Ni/2FEXw4FNTIYArW5pE
eyvGaTQbJshDK82pmfiLl0eeYQqA+Oi2DkpQzWhC4dk4vTIaJix8QgYpXVbs
cOsGAYPOvipAJfAX8HkLp1L9IqBQwREiMcIIAXNnpkPSYMrk+R/UupHSKtbF
SA8ZNYWeKyxvYvZxJsS7Nf3uNmqViizsQFPhYnt473yEayAFjk+2G3pBo6f1
7+BXD/P1yWNB2KZ+lnF9c0CzSfL/77OjqxS4MVFsQ6k23gWPkzYgpUd2FM30
0iHexQeSfAy9ecf+oBiouC0C8627s9yCJ2gk1IAgNW/hCpnqsn5U74PCUHi/
/6810MwAhtQ16daoKz0DeUfHI4SANXGqxsyxwiADe8Y6UsK9UKcVfKcS9kgA
RYJKbMaUv0uO++7Cz/+SJFbOfSOVh0oPEaY/eN08CR6f07g/lArjosDF44ME
UnrinxXq/qORQVDP8nTVDka1ZfkAzm7EVrp8Nnzq37ZSkN7Cu5uO8OSipR0Y
2OBq+lyzj9LXq3LE2nh7fQa6uQKjlyt4kYn2pL7Ymg0FbQfYVH/sjYytOZyS
cjT0bD14bXaaPvtBSgcVYS+EH6funb4/ay9eobLLXTG7I1Lyi2Hj7LWcwQVd
7Rt8W++BXUiRNhZ30Bd7R4R4044oPpNK1FG0FV9ibyGNk5zGdDO4q98R30Xf
CGvZU4B8sfyuFoOFlsk2oQa0ii/IKQahZq5WTyqppSw2Nyb7voWwcpY06ykS
VoofldsPse/xXWEmoTmKUC8lmnLgalhZAJCZr/QuPea2G96idRTg9M+UaA/A
k4zVgKANAcArySAEC8YqyUL8pmy3F+KT2kn+3ACjoAh6+x6kinSneHbB1K6r
sYiGdQS1WuxbX5OUMlVYGoPenIqMOgOYNJw0c9xc9CU5rZqsxepqJG7FPPEs
dLcen3iOB3eVxcEDFm+Rv2MT0SGboRt5Dtw3Yt3N95erv2U5CFWL1W9nm6Qr
RTcYCUqxaQsRLEWKRrUBwfHZLuOvY3ZStR+myfj9wTLouYoZpYQkjdMZqXYu
a/X4tiUz4ukTCenbcdzWxIKoQcG6qSSrH84jhxzvGV6bNuJbmOKgHow1U+L+
Pjim4Q4tjf1I5wBJnMgPhMSXdyuXQTqekSn65hvwIzqZGlHxBnzNMLT8AmpF
NIVRmb8uiEAiCLdhXIMI8QgTnULDxBMhI8kxNaaFNzZSqMO4TwNT3KjuIIaZ
+cdCD9baqMJkITCfzcb8fq/4YCc1SLXrQvkrrogPA1VxM5GhiOesQmjmeYLx
11XvJS2HCg9Ay6+hzm540aw+0PXH7AiYvgrGIW61ql0S0HcrmV9LJjhQdOTH
7aTSFZEEvmJDr/Zc3uU4OCVICjkCwpktPlmPQy8jkdwgS2eZ5pYLxpM03fKS
ifur4EtVuOFHpO42KGIimywaNI7ahpzqKr3W6qmL5OXsBD6Q3YH4w7PN8Nt5
mlLq857bI/YHJxf+Kz1K22sbbXp0+sBV/XVr+milRi7CgHHEE1uWkT+/lF5+
uz6FZj1MNA9dnRVb1bM0itpEzAaFZdlybPqZJuuBkoDoI8HL+cO6asVpto3I
a5okX+S4q2Ohj/+ffH8xb39REJDDz/hTFdJJMTl9FkjqiFCyWzWOTDHzSmPK
5hNJojFG0LkBIuDLGTyWgFiicYHq6t0yn6E3uO6Vsqn/dMIV+kc09OE5HN0L
aBXDqTN/8FHMbTQrVWF8qd5K+xA0+OnzyGUMPH68ncdqRBhV4fc8Sw24UeGQ
I3BkOyAbscYi4Nlspok9ul75MIYChLrKv7CsuE++7201L6bMDZaxbTHdqedU
RUpsHaA0kQ1n2Z9jNZf8ZRfm88tvR8QidWmlQwhygRo76mafnbmoxkSBTPxF
TtNMyiTZscrLfDNmEmjNTrRd6/2ItydCz+9CInyXz6qb/G+3BodvTUVbIqvv
AdGOU0lx4RKD6mGVom/u6hYsluYoO9sDLY7dKWCX+k5clrucUFtVFQKGBpKW
96bnRtdjuio3YD2PA6MidHIgJ1QxoDSp0FgLzpdZsERAxjoQpY59Lha0eFmy
9vyLx4y2vzj+Km5TLZCeTRhqEHQ/GWTG/Z7c6Ivy5glqpRWoHq9O7LDNxyf9
vU997y0RdX+oTePPoi1M8L4rbuEfkuxSvKCkVi0dg8xM7p04LM2Tge2YL04L
c02naUZt0f9BfuSrtNVvTDfK9gKMxhbqOgCZOy6EGzRu05JXqzyVQrZLtjwn
T1NP7DMPuMa3aTqI9rbKvxx6UtarxMGcsyFloYX5YrrDjYtHLjbOjFgV6kg1
HdnLPhkyzZ+sVA1Z+ymQP+gnNS9UlwPwGfMR7IFcs0O+n6OUNImdfbY6VgAc
cTQb4PZtr7OhMI4zdjzTgkGcXrg65X8IWFJvJKII02Ei84XO3JTQfvdBcqNx
zu5hDcFQ7ka0H+attIyc0vF4/6wLepE+V3YCM6gRWImz7Eddxk3KUGqFYf+F
xz0rsv7VvpKxBkkueMwtKmywlLHUv3dDLImIG25xJMr9ItK8guV8chquoJ8+
orhAXXhwwyTT50Wmtux3hGj0xtAOI2AbR/adt1QRwc0Y4QngebIp2OzLuq5x
KcdAuHn3IOslpTrzd4XNI3N2WXOlofpokXNeF2rZAcIoF14Y6IP3oRlFLsFu
z1Wft7J+iP4YCk3Q9XKrH6bDU7sOzHjlTSIWehsi+5kNYghVYfg2RKtwU897
ZaVKpA1QK+/wEdJft4eueW+czZovPs8T26d2s3CkTzxLwSXEiZ7kH0IuvoBc
x7DXM1JJXjegwoJDb1QOH0Ptap9d8dK7JSgyKo2wjRPKkwBdKK2ky0beJFYV
c3GQbTzCgLqumfbL0rHz0m/EolZW56xs9JSNg+2e1sZ7Ym3w/oC2TuNzcZji
6BVXwWuobBUlabV29WvrKDqgb365S7upICg+eqbvNkDv2c0gux6RiCfAxbTE
xjJv1vldsNpvlEl233zI+TqZ5VF513GCcTolbIU0aZMoEkqgY62wQ4oAtp4m
npJpfIzcf0rKHeE5HjVtNWpM/fkPBMl1pPup0rCDXXrKBS2eYwDmL0g8RB3V
kaIC8SYwfmUTcqGNNHxUpUa2h3yGdzA4LaWPiHaVrunZgc4wqhgXOc8aytd5
BFlt6pmZQu30C9PXAlSo1nRC9RYhUtm3A7Gp+Dkv8qVtpwIlrfjm4tBQmoce
TkY7zc4Zh8erUBP9T583Hsp7uyvhqZi3j/6pmAwPZ4NOyIrAbgkCot2F3IVQ
LloS1muNOmbuAxVy5G1+U68vBPeXeCDlk5MXh5VRaPHYEZs2mp82znJPsdco
nE+ii2CHIT32bAaImuUoKKPBAnuH7SKU7zWkxAH/5EpYfsHXb33OSwyfPO2B
0SoHzmw4krjfl7tpv+PUxs+C50MwhKZO6qs9bS+azUjB8xT98FURhX40iRiR
IQGNtRgmArEImJR91uQthCmuMQrn926fw0jv6glyP3rgKoTmav50KFtQQqQO
U/Jn/eYZhxIKtH4OiO757HTw7lg0QIcTUWl2JCH2tSf3DaFBHAYVZg8i3sXt
JrOI8b3CcX2b/+Jlqja6s0MFh/g12ZU0PG/DAcAQkHZLLkz5J/eoVzoqfNq8
CRtjfcjRx5zNpajHYCfEQsLlyDyZk3Tbd37PwoLDjpjWORPPthE/cyHCYGg/
yJ0cEmtS6bp8zdsn6ERaqlzBBLplaI6PobJQyiqmLoIkeBX9S7Jrwg8564+U
Gmsro5mYUE22msadS81StFEViHjOVF/ZoIVranYSKn0tpb3pUCXwCeX9NVmC
Hp11bs13ki5+G8Dx9sXLyhwSyc5xkeh6A2DyxSSkNzPlvTlWMagUpb4DwTx/
An5Wk7tdXjAJyB54oYDCUmjnIhMaxPvTxwDvHvuxcG42SaPG3P3k44HXQMWe
kK5bpaRUuUUNWDNSnt4FS7TdSeo+xhPaE792vMcJB+fXopop42ToCr17zdG1
RDB3BdlpnJIbmG1tJg2twJsKT1mHvWTd/ZU5HZ98EjCcU/ivzODDY7j4c9IN
7cD5K9rHHizqNlAr0OZUeUfNiLUe6TAjc38lUWgRRTRLgUHo9XFVLJhhO6nD
wd/+aewB3jC6USqOtSjeCfo5/7s9hS9/DkhZMhG4k5pM1w9bXvOfpOaZz5mI
IY4OQBbFBurRvGP0mDwG8OQ4NauVhT4mFx8oaFE3AdIyFT8CJgDwXWiz0RWB
ZCDQ00O3YoCHgisyq1ljX6koYB3xGsJi8UGVy90CX7UrEXXK/LYfVLNAIB6e
elCK2NBh3TnlNw7xopSIG4uYUuQQAsVl0WYTlaVIQgLT7RTE1SqjDb+7DCy5
TqxzdKsAX/5Bf6C2ZTyglRbFRxH+Tm7Cl7dXMuvZEoJfpezST8SQMPMloYOE
deFs85VmI0GH29kpUM7uaREhb7uFRsTVqTPUpHGC9T8yhdwW09FdcTd5B9nF
R7gxLMEuX+nR7VzY0KQ5XmxX6UsfXRmkBSycWObbAcMKoP8ky7ezSz9vISBc
sdzbasDG8JaVmCIwB59ThWovRNv53iSfq3exJreL2YEOXExAuTZ2lAPjn9bj
nHZBJBnjwKY8U28/KYF03iMiiPeHUhbyXL4bTY8qSSuU2vu+P70lx6GDjLCL
PiifRkZLoTWrS/DA4Vru55runHG+xLzcqWdlU5fRoVY4yD5kugFTmyIOilHc
Ntj60F4C3WWb21U7wKzZGvmOhfdastMOeb5zJmj+aoqgWIpvKZmKrTEO1SRJ
55OCQhFahZOredKdQQpiN3GNDUcfxaoe5tW243SyTEwfb+VBgZwptzIEdRtM
/cjpmq32J2bhaEXheqyN3a8wTer6J3dRvSml1kLN3BxhHtw1Bua72AirJ3rK
eILu3d2wrJBXnjdf+OeIlN4RTu0gQzuA0ePvVXlHMhT6PT75XDWAcSxHyb1s
Qli4/xpj8O5SwSVfkiuCud2WHFtUkIUoGEfIK1gugjEmyVweNynnBVAJ4GGW
BIdp7ccACA4J/wKkIndHGs8/12hPz3XnnwNoHR0aQcabTgZFJkhBQYBJfvzV
PS7Tu9hb2LcOtbWp/2hjOBilhrHKhjRmpdcq8hwoWOxqIUA5Gv+4fq6aGBkY
NVuhC8U3uYpq8FtI4yo0KPadwtpo/uzB9kpwZGwWRE3lQ66894vtqqK6KDnG
ZRt7mh8vet12+ZWYJ+BEkglNe8U5X0fEndG3/jhpxovwMyDRw3qZuWRALWgG
aiy9OpNJtSz9VLGw3E4NFu/7AqllpMJB4aaF/Vk7O1QYvpaGlx48U28sUiF1
GwMDD3KZwmoINUK5arOvf8hmqzHnFs0cJcHAX4PKmY0lXGImIJQOzQ3ev5V1
wYogkPSQbe4LGm1GCliacc2JmhETFLqPr668WCXIEfFX1a2YwLEGZJ0K+Auu
M6bIqO+957NNdI7xj1Rk+89rY1mWmZ43uyBB7U7WqxkWQuApwNFyaI2z0r7Z
rRQ1xqvQT8uHYSlP69YumJ1eYfBE7nAS1WTiMNMMOqLnzVV4w0+6DEahuUfc
aOogo5RKJkOqF2Vwf2Uq5ZkhTmPfEVPd91EzJrhjP0qdJxmaeE6TSzsQIdUk
zJWTXgASdfSVhENmIXB45jsQwbbETanTepYpbqqivnoSomdcOGMo0tWxa0FH
JUdALDo/P4cz+GU0aocK2ZVuHw0B6narp4ckH3DMae/EX6UO9um+Q2Yu9mhC
lJ8WK/JlbEnZIo93ke2R78hON+7xyMlvH2IFh6vX2fvyHDNMLQEJhtM0NmaT
lykqvGZH+1tnuQBr+zvXV6E1HI7OD7Bvr+HnVsERizoU1F3j6SHw/k96mB+E
xUa6PWEkYsKBQiVI8Wf3UF/Basv5e6kLsVirzHsw9jFR16xxFPyaGvXRVIks
+mpNpuNl2A5Am1fcjwwOAO2mN0si3/gQbm4vjBzkRMPD8ZbKmAkYtiOJFCLS
74X4ssI3kp6ByPNWSzIjxmT1nDxcPaRs3s8WJUReEbbFM52NA95x4Sgbja8y
tYmBYdQALcbn82XW0hAtHX2JTZLddIbFwTCgEKcyS6hEKb64kY5Ei9BkQsUQ
WcshFxTNgCwRHhjxvW9QVyb0e5yWJkyzVMTM//GgyMBKjKvgcKrJ2+ZhnlTY
KfESAiVE1Ky1zI2lys2ny9z11BbhJ8CsQk1kWoOlgbdvjy9Hr1JDCquv+YBF
qRbNqwEMIT6Or/BfDqUp4iAJ6K5l00OmbxSYt/m8iRXpybjpADfJBhBc3OeS
ylOD9J4Ngp/IbJJn0jywgym2ekEvSpG0TQ7GIRWkZGtLKf/kfCtRQ8/nA3kn
xVpuRT7lCCpxdQZm8smz0oSa24p3uAB4D7BQCIOPOJvS159PI9rkFYmije5B
HLsa7NZloD3q4L/OjA9uxuFz35geZ8ehs8GIl7J3OH5WUswXtz3pAgp5x2aa
/gR9rtNwBt6xD612Mg0Rvfj+O0/7JN2JTFTw5d1AIjl0ZIMvoLwdhOCdYgcv
eW2acSCN4wWtHkiTqiXU8xBPy6wag+rT19ItgPr2GvxYgiD8xfnXhuinPsTI
KdjSYrxg30GBqJKbUVUyI98Mz7JRQBU3HY4OrPbQ2u7LXH/5M5M65Cg8YqWf
SUOgXFOD4PdN45YzTWt7EHTltIBHOi1h1bEN76rGjL0CiVc+A8Ci2xfBs1cZ
xlmYU2d1jDVPv2qYxyEkl/Bfdo6haPU3TB+eVycY+ifpPsWwHfS6SzhLyZdD
ORqpqVDjtWipZwIw09+x81So34nfCeAFTtlEsQYWunjbhgdTCUSGuEDUOLq6
o5nQ/bHdAhFUJDxbgdiUPKvZTSpeZY9Ic+CtAmUDhHeZkGpZwnXzowYeOTyX
5ypq0hqxYSG7pMT0nCn8wHskSkPzSXLbrTaE5pKekpmihiCBQe9QXWbMr4fI
8h8e5U97m2KvgJZ+sxERYZZNu/sozUjOSJP3i4AU9kaKQ+5DBpM1wNZRP83d
qXgoNOkxg12xYhW3O17BzAJYWclcZLYIqL6IllUt/pwS+p6/oyC7sZU1a/gO
LPZ2WpzXgwRy+XrBykyoH++vdhEhlsBCDnMfP1NhLmD5D5bC5uwaiEJwRS7e
6+xayL3XztDuihfsePX/0g4oEi16HDDfPHejWXBvUKL+XJ6uqKct8uxQMB18
hxqLw4jQ9yBygQ0Y2DjLLd/qA4vTIFoBfYT+1MsDzvVyAQ3PAiANM3b+tyFg
aWB2SRbxAtxNlvFKs5njrBWWFK/dOlmFaNwT7ANYWVbIm+iy3jKAIFySpC3/
Vqvmi8CocLMRXbNBwFTXnIguXtsUAHC/QlWZjb4IsVYn1/xSGE4hFPf9LJF1
RoJTO5CcdjcR2kE1WB4VUA5OZgMBS7lVobWePDQ+v+CuZD/RthKBwd4ROjNi
U4Dtu9Rhfe+GiDlQ8s7cellUhKKEu3gKeGTdVzv9m7irqMYObFTmDfDEZXrM
BGh7g62pBzPoNyVaw8BlCw0P/Rtsa4nOa8OgaOslVrBBBEhGXq1cSmF7mM01
6D/SZ5m3xv5g4w/HUJg0UczASMKcd42v5u75L/MaQ2J319R3SEl4w9HnxcK+
KPj0GLdRekW9UJP1ZvHN6n2sMFnW6czBBSNJEvwN4Am4vIe5hjmsg2zRmFXn
InfVJoTZ7DL9PiRrZVeu1DohphUL3SOojH1qeNkfzHZfPAOLGYPS21uN5/3c
8k/2f7KlyTfOJ71bEXEypA/UvUdWFquItW5FBkNhA0sxem6ZQcxekr9rkKzH
bsAHX4G2hjmcpPnFkUNr1NqPH8rJFFO8+As0aeDNmt1n2Bd4M9lU9ybI7MAt
nrzvhmE6aoJpTZtcJ05PvzJjBnhq0JOxrT5ChL758uoKYv4aM+3QsUQLVAY2
vo3EuvgBNNQHr27pYSF6aLF4/1ApNVGTpRTD1WMFAiGucvLobJaCwovudjL5
U6X25p+/CfL+wwhsXWS7dGOZYn3/xVas4U/b75USxseQQV6Ld2w9q+5jk82A
kd5KT1N2fpIvNtwBicMft4XarHSEy/PXFaDMjlgrx09l+A5Hr7zBIPWJIjSV
sPq8ryPur1dJb9VCWgk8asW8ZWRIXf2xtKF66ps5KoL5WGpCDTGsNv2JgkL+
moBrdgDr8uHMAL7SLEhNCi0ZaOU2J0Lnr4A0J4M0bru7OEJ45xgVddK7kkxZ
ELT3FuobLc+/3ftKc8SIXVNiGXv/V1Id3t2emEvQ1lBRF08+qL3+Sv9yY64C
gx1NhvocJkQBapyaNYlVzmsGzkXXG8RlyC30DdArsv08Ebyn0BcLkd92LBQr
q25EoBcvw9sBnX79MhKRj/TfwNI9d+6aGI9KynYvC5zbNNdFfDa7yUbKgBdR
rm1HfLH0nQGfpD0mCuUgWM7cdLN0mLfj1NsrwJecy7vCZauLwCyEc7vROGEK
ClCLwobMw/Xk42eSDv9wPqT9BB0Gez67NUji9wQ8XVwhZncp5rCBMSf8v8rg
1c0AfTQj1/X91h1fYipjG4dvRtR5EwpMf/G8J/bDaC+1exmqDsYJHtlvnbKK
q/0GX/0knCv9vaemJOza+coaXQGLTW+vrCBgD8fOX6akVbrJw7MvUp3PA7ai
PWVLfOlK3CH/Ghs++eD64nwDM/ysWhzisZzXLlgftOeq2Rpy18yO/gnSxR+B
AETFv58YnKvwS/AfskZ4CqOnCrMPG92JAgQOKQPTK22ULXbP/hbEq98+PSAN
LwSrsSOgjCOeqQk1kz4mPDWCufqTvbsfDaXfkt+0zKWpOqRt+TvDjBDCjWcY
lsZZ+MNLwAfSlWZknb73eqQhSxzaF7/QEKNZlmCIpmwG0XGuOMyLEfXe7HdL
mNNltOJHdVLLbyxVx1ls8leLhRlVrL9/sAaUxETiRfCLqxUKhdVCSUSseKTy
xc3MAHiovceiQvsW6d50qxK/4tdXcVmaWG3zDFSYyqfltmlf9nv81XtXPfqs
5GcA0Wqw21DaNk9KQf8RjO0HtKyXse3Ho7rThRKm2qBTDYW1B/dI28BTxAUe
/frCP6U+JqaoE5Uw2zAIw62TcvaQ10RzMhwsInDwabbRAdcJPW7xjH8healF
VSLw350+dsG66WZpDUT1G0DdGcVKIfnQJ3TFvPBCFXGUd2bs6I5ykm6D7Ot3
UVcNqcUVxcYuOf8IhntVS9sHc89VSmw9bWEipR6R5cYjjG1isVXiq7rgntDS
n8fDtmVrp/r4u6kcXKLXmeVRXofzGRvhk4yc/SqRdmmyFtYj8h2mSmSy0jsN
ttE+dbv/S11By9cLYpOYslvz1fuOAmeNWA6itXEuSKVOFStNnm4GrZXxbgtu
Hi2EipmLGSRtg4nEb8n18VXKvWStP4V+1FoICQBvTKkNNUXU8AaUCTzfyVQQ
p07QzNdZbWVKOCpe6C9crEbFBbm98jkr2x1NbeI4YqNVwd47p7tCsfNBhhJX
9IvpdZYDkwTYKos0uo0yVhdpg2Pnbxzeh8VDUlULVGOtOgCIi9cie9t4l0nl
c3nlCoMPmNlXmDOy7aQKnX190Bd8r1xHX5BOL5npXsntbllXahFMBkeXMQT9
QuBFmA5DJmxcSLUhHQm6ytw6C/5ahQLx7UYAtGnRUKV1pGYqt1gUKMWxGotE
1TGpdsxVyoOoHrIayCurrt5fOOwKxFrMMUow4kZ8ReZ5YBlP+VJ/MIrCRoll
xzjDfagBDvwNx/zZXVbGJOO6nCMQILEvI6izviOLzqANtYKIwpCNgBmFiq7c
Q1xlE4H3EWmXU/MHTj1KrCPGYevnJfYDc9zcLbwM+DuBoPS4jjuwXIwt5ueH
uIPPnf+fqftAjpBeY1U5sml1CfIE2ncthCqp4CpDYZiBP61/8ib2XF+0z7ef
Dbzfv033HVS66RSrFA4kMAkm7o58GKuWWtYBzChcsqo7U6/zGSxTcnkHJCZ1
ehbdq9qTAmrZrcCc4DL6d3CeqVvFqCK6/3JPJJlMxDQyZnmyjv6cF9xD+eF1
xbFKasz7pJpI8Nh6GN+TscNWWbijjwOA/mXkEkvl8m3VOieibotMe+Z+u/Fv
Nl0GeCsKcwp115Lzyf9vjMoyLVGGawDppP0Y00qhy/6OZJqtlGHGPdgzgqQJ
8IET6II7l05Liu0bZDQ56wgJzVdBiT6PYRjCbxbrOtQFYVAEcMp+Jk/3K6/D
mnjFSRPEwWFm/9lE62Ejw6HSGIys1MQ7Iot3VHz8B/1O/s1PQDVoqOg5//sq
0qnTNAeFMkPtDf+Ft9/fty2AvTas0Va+vWrc13EoxJAEDgFfakNBhbtfqAHE
qG4DWxqhyygaT2dYLt3zVE7PVSqSTOaIJinf/mLkexCfT09NIWSi1Ma4H2Sl
zXEdeYjTudVY05YLFvaADnt8HZx48zUrA/QxrVpw6FF6WXNJ0tv10ey19gnA
45Fj3pH2YTAp7S538oNy41NZb2uW5L0Sn7RFxN360TQ6oi5hLED3k8iSi1yj
+/VDEMO2F1E3lB2PFzQ9w6Lr+bNRBwyilbaDKkwtLasq5aJTsF/c1D08xVzC
zmrZmYw83hoqUwJqEaPW+3yb1gFnIP2lC2056ABsK9mOZTGDekuFy2CRqibH
tjlidYekN3LBbiLisuAURnGTihXVYvTO2seXpiDi9WNW8jconOEv9IpYjabG
4ZOcydkD7cfe30PfUMRDStadsvLPLLfbpQxFZuQIiLIoR+MWKC/UI+WriYlF
FrMcXRdVvGcxz8vHxDaSUztAzFKaR3OH2g057uUnjnhdYe6Dl81bNF9Cooom
kuVTbgMms8DTJcsd1bMnIBjx25a5J+Wlk257xA3KSzoaEnONl1XDzKIElHvR
+GVoKeK5+CBlKbsLAPaZ09Jn8P18bX3AdKWee9k7ZW2DNC7TvJePqVrdDpz6
lAH7s3sQakJCFancGrfNKZyue+t4lff9Y368l5moL+LaT5RtkZQu5dSG4TLB
GQYJDdjBTKPypcLH+i4f17CuvyhMDKLjY5zNF/L3N7jUl13lkgfQwB8g2OmK
/FVIdNOUqWzysXppsvQdpZry3xiXBsqb3iJz5SYf08+1Qhqj8O+BwVW9btkv
cD8A1ETM+H5sloBF9QPE/mZ5ZBBMe+SjulPigBVKFzcuBR7roknQo1jnc/ur
DbjFzsL4SUDmyhA6o36SoAWj0PPxfdZet8kSgaNoARfXP9gmew0Ey7eP9hiv
hlApLigx9WMVjYEVAM2ToJ+sRRPdMV3nPw6YHoCJUpnPEygXNK3vb1b91+LU
poEzxYpPPSid1voQaaCkELi+p3tNAE67+Vnl0uAsnLiR2qzlX0jDwOAxPRYW
wa9HF6y3wwlQfZAGcj/IpjQwhpfEyD0OWacpa/uQk3sqIwRoYowx2LbBiVGn
2KWVsOexEabBWLXTxdB1vb/EMTGu7KkDLP0iCSj0BkFHkTVChcMIcv8wdn2n
o5fhlsv/GsEnXgjKPhi5njWBca9j9GSvmDa5I8bZ9MsjCqM0rS5cO0p8g0/c
GQ6LQ+qtvOVSzgtehaD0oXiL7KgClvQmrMrsTMjsGVsMv+xE70TFTxlMBrZC
VT/ulLXJCP4b2CBYMqTNlN6MZpHVqMeHLzR3jRAL5G2lQQza9n46ts7msUFZ
LwI8+rar3LpOk6fOpxvXsu4cTA9W7ipomH1BU5YBGQT5OnvDY3tX8+KE7p89
ULw0JeI8wjhU0A24uaYvq40lIHLP7DJ3z3HH7EJSPNxuXsL26MuOBeTDTYR6
4NZB2KeYaXQHqoO0ydSjmE3Z8JPE7Ghxdi6MLO0zzmCy5ionBg4aWbteSoIq
yykJHwbuV2bXoNIHTZPP7YKnepFtxFjaZs7yYhckAq6UULY3eb5ryqlQH28M
vnyU3sQgAK3ncxIBF8DVafdwydto5CjDsuXSlrdDCj1b0934wcLaJenfOC+I
AyhtNefzltUY0Q90OJ1HkCMPUyZa9Rqm8vze7A0u0PvMgFuKraYQR648ZVzW
3WB2ShSvFTNZIoxt3wZjljCSHE+Jgov9v5SJwPvm0HoZr4TRlwmnLfkg4+84
S1skR/qLHRqzj9+fXKDjHg/MXTqFw97kKkCL6Q9yjA2QJBWpmqgwtcbX7Bjo
XUJA7JPyMS//WAsQV1G019UjYN+A86MRqKXhFSaaqodoxtd7imrAlcl+8vIG
y45gokjHa/AZsA9pn4+AtdBQCgytfPlDCmMtfSfFqOBc532f9neorE5kkJJI
iImXsdoAPgXu36NB9zNQ0dNcod+vL1FzIqbCYxRcxeKAcxLwcdXXv8uP6mP8
qT7PhtNSeCYFmkI9HdsJmFNCigNZ9/m0cBqZMCU73GoqQmB0qHxmlnMy2Kj5
k++aRFgqDbWIREqS+Kl/OmrlwPUiJV3IlN/YBgDqyDnW0uun59n0i+lYZkE0
sY24gYulFsk9efKEWIqGOwtMu7kuYz60wbXaMiKympLvxavtxKad4A+EAfJq
09mjugWasWX8A2nKxEuKyGOq0sTWU7DgRQeI7BldtUe7tToa6c8OkVPsl/jh
S89CreX/nInX1wn19ukdptHlUxkIPZOeqZhGnKFH5BVeJZaarBjHCAVAJ6su
Ws8neTDi/6+w9rYpwgrlQBcKvNIYpi4ILxnnOaO9187o9qd/MUHz7bceadWI
A3xP4Ws/aSSr1ZRXvPS6QzfOiKVXYgc/RqqkxND8XPgC9PQUIpAEnurHJP3y
MqHhQbYO7BNBxbWldvC5bT+xFhpNFNizygiU3SRcqya9IUSVgq03veMfbtWz
KEOWBIv9VZN/ALTjITccGUeqr2jBkgTE2SirAnsLEsEyuwMhTqwA16yppa8X
nxBCbj+JexPuhfaRpcV1JVWXJQ02mAky5hPk+3IOtVtm14cz8lqZEYWQIeve
ZPwkrwGgx+8zel2ZU2dzrnYkKkBtuzPABo26qGLY1rCv0JcjTDZkxAtSL9Y4
3fCaTTsnRKWVM/S4g6qOKnmmV8F1JItH0SkeuEJs1KRukjhkB6/+UdHhKjA5
0dIPgybQ1NPHZGyrpaBCKzTIOBNhXRmdJozBncvbSk+E408Y8UucM+N6g59P
hp+ni2w03ufu83Wjjnj9/GJq8UTXiTmZQAmK/xkCe+FR6F+h/rKn9+1wrIjV
I/GGAbST6C+QOmcbZT8sA6cXrg56axop5EOUMC2WAz9gt8aPd+z6K59TTKOf
MqJKyXn4sPQBkhwm55keUE0Lj3ZFWfeQEw4CKUf0Ls0BbTxxwyDfk24O8YhO
sWHDVwuEpt5hSo97i0Tzko5+4n0Xp8vGgmODkFgCnyoDtoE3fSBNtE6+pMjL
JYWIB0EG8PyjxBmqlFjhnTRt9C1BmJ9gEPlvFLN6Q6Y17Hjc2il/nFf3Er1j
8F8msiYC6OVMnouc5pLKRUm2SogrBXXHkqPbMVYx7It/cWYtJk6YbfVYT9V+
PyB8SOz7BYqJrwCmw8Ibo+erPZG0LTD+7RqwPlnPBxzpoi0ZC/a/TSG4rNz7
njCzSEXXlnTfPZ4FLTGD7IOuLapGRlD48NJqYBpcjlkT4soNqgniQFqEqIUv
Mjl/B4HY0uvePdKzj1ZbKqqTUPrPSz4hmpMRZKr7HjeBahDx1Wqv6rFhVuxP
4dw8YmVKTclvK9W3zsz3vYbiXuStIN7Yt0P7spJsgSuaOXv4ovi+olc9hOO0
VwRwcuR+UWKErpD8xbc1WAZrHiYrTk/NGEucWOByNhX3spYne/O39Ka0C0GK
VxtyRcyo/j1kMmQ5xLWMJFqpBf5rTGz/UohvRhsKr59rmK0wfkSefK7Nwsap
z9YltWtHMLV/EQX8EeQluV57AW/kUpovKErZDoT0/P4I3HF/DtqjduJwqIeM
pESsdOVbwlGOkORl2tyZkjTtsZICOg9O4e8Z0Y30vltzgq/tSgX9kP5nUnYI
LUYlX5ccB9ld2ntVouDnqhCCrQeKCmeUirnJXka9ggeLwTZTazsuDXxv5Hfi
HVThQRFrhZ2yMU0NsIfd3IxbLR6+1XGSOLF9z9VD8Rogza34pPfDiI8HxKao
+4s9rv2cPX4TI8vDtrYfQd8in2WJszPt9IvbCUz93zUeUFqLfsETzCV7vjDS
ckAD/Eq5C6QMaGvzWYpZZFM7RtRkET15sToA7GKM/CnMmH7qHM8QYSDcqhw4
Ua5UhcBkx56IuVEYqiJyCxbBs0L6VScYN8MzeTjgWnUp4NVOB8qQ7GuW5T4s
/tnw77Hr9u4oLHvrCeuFXMNjsK9+6qlKTWT+QGTUWXXLE24O4dFDhn3XUFb8
BMlaBYvo3PNyAok8N8jMeW858VgFIkaVazJVZjPxLJ5g/hBYYbhgKh2GLigi
MxqwQi8mV5BuwIir5u7QaB8v4R2QR3JosGMSdZ9kkninkOL4XeQZBt9z7yI/
LygfL/1VyCl81rj0g4zbY17u8uOpuhPYeUbBFt/mwwZhZyw9XQTasXDolzzZ
mbH/yRd2vUULNx/tRQbSQdj10/MJnujq+Kwzu18v+SeU13uVKH9qXOoVffIb
p60VE++YkrZAsUN59mOrcs0wNJXkBT9ZCFHF3EtktxYxpAuexdl6Pp5wi29x
3wE9zpkE3ta3T1vf/yx4cCfN9O+sPxHZGMd+On/d/dmAn6927A80Bb1Qy63/
z2G3xh/a3DLvNgrCHlAXYsn0qTYH1J7q/gQi6rSTo/R08xLbBrbstoCp7K3X
byv0Pl4YmOwuHhqq+r6q83eW2IqfMkRpQdZfT2+QDUd6MNz7+kckcucdv707
eY7a0YmFW8nDwzmYQOhlr7qh8K5mjqYyoPVw+UA2hd7FWhJoDcPdEBZokzPq
bVDo+18n9iNOTriEIqT3tFMSmzfsNV6k5W563WiC7uknWhfwpD4YlSbBaGVT
ZW0Dcpk+iatDZmCSO2Vl3mSszaGng1WcHrMJOUqJAc3xlMnn69O3H/bccYF8
tO+0bN1naZsCE16RPQdMi0fJBdiJotA6hp5bNla0dVd3xKG9w1KNPMD2lGK8
y3kf20Nnp3qcBwXZTOFRJKTZ+rHlBpLErR6/sbee+t4AKrgzH3ABNXQbjwRF
33mg9EH9JVUt9ZhhXkjwzHtZt5UiYrdmrO5dDSsmHd9G6NrbTiObhLUzyjcO
9FmeuKGwVjkYMgeECvxPjwDulRHyLqwHtTMC654QuEYEXDDwb7JYkwSMDZde
0Mpuem8xZ3fP4Ub+U9hx4xQ/FLDAIyLpv06dqAdfMCs4giv6L/rUcxj72aRG
dOBeiD47A9Xay3URJ1ldSYT9x/fXDK45g3DRkYgyXgat0LAEkrsWPPdkUAwg
KG8rta+Lg471pK5ntOdNoSc7JKqvLBTCkZMD049RdycU4TD6wkiwutyjnIVJ
xMP7R+P8MWwgdpfnYxgJdzIsvrHS59MCjXko5GES9y8d+WlxNh0KukjKPu+w
Q4xZBY5N9wZfmKBgjSYbt+3TsKJuHfYpRzyMCkIWCaB8FfSY6FiOm4Sy44Wo
Fr7+ZoE7NK6JR1zptFW+wrnGUy8som3t/xBWaRSoAcAIWSzyt8BjHXfozbLm
3HgmxXbBF7qC7c3NyCRPMuJtG9S7vfGEraBJVCrCdWMt9ZhWkn2ed2oHIAhw
A1ngvczpbTkcKeTwyhNI6ZC5oQDccWT0JbKvI9v1Fzb8RoVjLmilx/8XPmd7
TMLS6lGwSkDFZu8Snnj1ShvkvxCiF7xmNg7/KxYsjsIVRGWf7X2j3awMYXwv
/KDCTtZqKo06924JZvGPW93HON9npNSYQQ01JbSciJSzUUJDO8Vep2VuyGoB
pAgwdzc3KxvSRE1er+aCqhfAGJ9Uqu6rFk896MKAEEB+TvArVhAB2YN4zj+u
ZKw2yjBDwL1FF0lp0kscKhkZVVuWWjyK8Sr7JulyW/szRvj/gWEYRVdtpnMV
pkVlM92erC58fmcjVG38U2JP0hlegytKKY8e9u/zKPnFJwBW4voiCKLMSfk3
aP+/BejVgcpozOvuM1tTs05tdxDBnHUC6uXdry6ETd+rpe6SF/iZQOaCpYAp
4ZjrfDn6VrGVaR8BfWhwqASAxbm/NStfAO3X7rEH3iVsqrS0RotfPGBOk2PI
4QaMjXBZyGn/ShXu6gfHbIhih9H7H2YaOKkTGjKe9P0LmGQoBVPG0DQrUoh8
fL5/kY2n2yDAwzyUAT21WWvcdCi0wutqbGUhAq3BbUC339d06xSsk6viOa9m
IgYdI/0bsi0hvEN4fmHM//W0suWc51GNur6uA+a4NdylOgZ7RRq+wW/xBgW/
7E/ub3mzSZBLO4YBAOTk6cK8PtmRDQbioI95n/6Otnj8cQGlu8ZW5sEvdcBc
rJhHhxSMkgOfKEzob4aXCMFry0o6QH2QX75qe80aVJyqqsj/uwlxGn1keEPB
U6tGEyzkK33dru/hpM/qGmanNw3/1LH4gl026PBOXWAnNk+7F0Am+8dxjVjC
xDOFRc62Dj2P0pEoic8MgEkYSKr+HNK+7JdiIWrzaIotB8ryCi2gAKIy5PKW
yPQRtN5HBH9S5FaRtdt2A6ORobaMufq613j59Kuh8PqDmTWtuflj7hYPLtnq
+T75gwP10CKXjX42tK2ph8Im/R6Oe4OrCqfv8pFpc2u4w1CRv4dAioXPUEW5
XdZItEWDHm+segHvqssZvfgj/mRwYNjFIWR5NESFevwyJCPE3QbrDaidBXeM
HAzABVEODtU5wLNeijqOX/KyAGTI/Uogwf8rKhWnKJvQdxq8knhzSwPZhDcU
/q99B7COdcVVIlbrsz+KcHFHpIUlic3L6fGo283L2n7eUkHW2vSdllHPe4ql
MJ4JLGPvR7oQCro8cG2E4RAJhweMQYXIRM7pEgfKmXamkceCaDDF88NZjtea
yIcqdPJyJ3sV0UlUbaRXDohvbu1ozza3imBVqLWshzLZaNbTHzIvPulUXJBV
lptW6QzhKZrIsudPkELR5rjBPG64gAlw7Kd6uYKgHhWKnInu1BA9RryHALpo
Zj1h0ELbPVdUNoq7On3EjswMgenum9ErIX3i2LOd++e+pM6yZ+Opok5pgOEX
t/QHj+B0WRxn5bWYxsYKMubCZTW1vp7i05x7kQlSxZHcOCK4Wsq4yX7ScGzc
5XzefFevVkiiB00CWp0fqv8L8cyCT8iO2p7jhwQRItOkHekzBCEtdEv2fzpy
d7CStTtls7cuWkXj+UTOIi4qMtGDXcuLkMNMpEZBo3PLcNVizkq55uJK0lbw
WRyVohL/BWmU8H8SGMqxdRI/D4dBQQ6NJRCI3/h5cvobB/Q2WlmBzQIDf5Li
IxkfI8jsvC3nKVp3oDQny2KvpjfL1svNelAASnSsYjmmt659G2sLWK/j+EiG
ZmzZdpMrqJO4uEBB4R2l6AgFOcrFOdh+rxHqET257h4KFTgxJKLTP3OVuSVd
d64I5bNRKKDU4v16PW3PJ5y5snWxVCxIfqLU8IMhv0fTVLXIfGA1ljYW1BK2
DllVOH+ny055Ntaohb6CAmeXpviUlkRN/vwJcJusuJP6B2AncthvP35IdxnE
2lgiQHsLBFUfce8KVZbJiwMefApQpEkumW9OKrMerCsZDIKl5lQO52WKMFdu
hUlW1qJ89b19NjnW4nbVVB6BpobIknmdirDuM2M03CSDLplu/WeQ3T9fmTXq
j01RV0p3sFKyFoaMuvyoUNAFEGauNv6363m5DKxTzuIHtPt3WdwJM2KMtsTH
6bKS6tpI75nTsfj9jHpl1G0npVq7sKIaGoLdGzhDgn2XcGZ4ndPQwDsPioz6
5CAhAarGCJffvkRzC8oLtBI61z8TVQ5HtGRiAhJQD7kVPq3EGSAfq81k6QPG
p+vBtUF4r0UgQFqj97qF/9jxJg47qaaHRrsc6T9fqX2jNvIpHxFyMobqBTjM
xaG/KOr0UIl0Vshtbmdb3IFruzch5NlBk+Wkga2W1U/dj27q5FBVQw5snE3i
eY+hMdojSie/STlrdNIxBZL++tTIwXcj18tUxtJQ+KFfpfYK9TefFEx37Lf+
ORMENONVf4wpJziRHTei5SzrS5b8l/iCmtmIa2WGlNYVOUSLVd6xgo0ay/WJ
71cTljinqX41+ypoTes1o2iJcA6mPIB6RVBxPBTTfqKIFdtjYgTeTO79yzkF
wuSqK+VAqaY0qisRVNCFwSh6qZlvZkAXPnJJxQBA1HFBFiAKFpf8ExFNicny
RnI8D+5iD9SrjnFGrNneXOK5HScBuWPdiZrewGEdkUEhRULpUf0DdqGRa8se
1SrJTROz4ke931t+qGVsv7HAOOHsIGNHgDpMNzp7frBEACkDPaRruS8XgJYt
AQfedsfo05/gGoKtGmcT1lF2l4Bf4l6717BK9gpB9V6mrhNbISlIpgsGVltf
iZ7Kd+lbc7VLa0SxIC4LwLj2gd1jmTMXfqtFWYf4n8ZMoje1fxHIGQItShEg
xjlOIgofFgkvJiDMR3wjD8GMOHDWyp9WlzeOhjJqCloJswmpKVmy6c6QZ9tC
pki8nMyYLwGS1/bst2CdBk1197Ay7byFMPYOm6cLEVc4WAxPhVR6ixRvLLha
hlikCmyE7QMMcS5gUhPshIjlHx9YRMfX+ytvIF9ODnXmnnPsHB2QtYk26KPO
kP8jEAx1Ql4uWCqZlex/F7jbRx1kf6sTRQT8Ix5iTX9iqUxVH20Ain2/uMG1
RodJJ2zAy4jVhA4vZbO84QmvjC0yS0Qoyk7GWMJHhxdqjMvBMU0/M4zppSpp
XAQuLaIw3VRD6mxjqpIdpPY1Y7RDn0VO6xSRXWpVZ+BzroXDbNrdnScaazKd
nllTSQLVDY0/P2DtGueYKk/ylluHSVwX/LWV8pRsJ4pKvd0K2ryHSoSrfXwZ
N9CC67ydIVxlGobaZqZaXlG4RJuJOwI3o5qGKDHGnGSyK9bcJLhXq+gwK+ur
RuQlLoCAAyhPKIPesah3pmTmgzkp6pIsWlYnJ+84d2E7OY1ET2eQShZriz8F
Wz0kEi+pPh/5vML1+FTlYcSlXgXtia5XIV6DLKjMXvBixBGk0moF7pPNbJRa
TWjODaTw74F28Wu2bg/rGmzFRRDp/f/ZqKBYAUj6Rr2+5pNtpAAro4EdR8Q2
iXe8EfzY49zmIx+7DqGUXIp4eeNMZ6Du7YDaNRcbmz6KYsEimzd18PEtPH+m
4JJzTaHYMaP2HZaKknnTRQEqMwMhUypMPIcFLgQ45ukZQNLrz0dqAF3RJNX+
ClLno27H1X4JkSWW9JiqCltBycFfCQ0qbAV44kaY+NdbnXHx5Q3t2xISzYW4
uUcs8zsOy7S76im7HdR+eKqWeekhjZ2BNlekzZO9N3InPixOyYH9tYAPncdc
g/HBtVkUuTWSWhP7LmOF9ckO8XoWkB+0Wh1g2W/D9Epl9glJ4A71lDVQSCJ3
xWHnw0bwZT5E9fi9nRaTkpC2rm5ABxbLagMPrbslWouB6MRJ+9boYXb4HGcL
KGLw29lvSV2pSjHxr5DhJ/XYQsJkNh183AsdUDyI61fyK5n8wpD4VwzWlrfF
ufuQLRS9qytPw8qnlK32wCDHN1MJogslHudOgwFDppJLQE5KMQk0ABPv2HKW
MIOVFMPqF5j3RO8S1D86VM1qMOvuH1r5SuH6DrSvo8xHxf+t1iTxaJQPp9be
W/mMkSv5HzXcyLBTgPzVheAk9Fn/ws2TnsknVZbU2UVLeUwHOajH9jowD/9Y
q+hqHp1PLPuPd8pwFVmZW8VmHBv57pxJgXS5jMSlMNh9DkmXWMLyFQyMEWzN
p1C6t8Owz1nsvI/LgM/7acJE7SrN81J5ZT4DtnKXfThZBjYJH28pT/L4RwSX
P01isLWuS/kbHOAWVOdWRkyye+kNZdcjyWfViFuZEwrhHdPAGTchzqEwkn6R
CfiASSrB84L7y/Qnnq14bFrc+YblXePXN01iV/ZC+IEvbeJtJiJQV3yyMlXh
/kYQfBixTDYyn+FA2Be++EINkS23bbuDFiAiXPyh6xsczWGn0AWciw/DPYVe
/HIk+6Ma1OjElHjCa4FFth6B3aBTP84H/GbYl2PKbjYQvUXVBP0WlM5hmgbi
AjaDGlZOSKT6+qqk7oWiPedDf+BYZ8GXgdYITuBpmz44xewWjAVsZ35M/s7Y
wjTXRhnoUyZndbmb8SPu0jCfnwj3GX2A4KJwqq4TKKwcqCOv4Vruxbna2xS9
mghqcSgDs71DwP3m6Li/IGfnYWEWkfxPEDs6vm32eYM+upBVt4xtQKhHyLqT
jDGToU+MkeeC0XRe7iUMWs97HPE1mtT5Cr0jM75jqcBUN6fNVx8/4yDVz+lc
OUflKHL8nWHGP9oAwBPqEaj60rmJufJ7r9llRCnsnNi8dz6XR1MPRK8giemg
32QHvBDjODq8xKqrQgHRdYdMiQ+pvq3thVKuTep+kOz6mtuX86o5Pm4BKOjZ
Bf4PON7w1aA/9L+F8quSgcxE2i/1QhMofUuSvLkLm24gQd+wBdZBwM0mW/Mq
tccAmaql7CjKpKITjoTneWw+TVNkZHmzzIEUg18RGvmYWfVeQZBHfYeOg0iU
JHJT+m55WCviLS0o1IW2CP0gU1BVc0q1SqqM4Tu6apvVA8e0PHQArAR2YwyS
+DTT8MHkuQYBZ9Sa9aSqKd4gEX90SA1xxBlry8MBIsyiVwKiwh6sucWziPWL
SL6jQE3WQVbRJdwfQ/2kGNA9uul1ZDaD7vlIu0sHVlXqUS4b6rajH94iJEdG
tmUcdSljGfEVvDqmFPrX8ZNSbbvOIKroqHB6iI+sV1qAiG6mQ+xgvgvVvGut
1PSE7hd61ldGaZQmnno7U41pud1XL0ZjZXEsjsEkr0YqnqiUUr9DkEZv+oyS
BnfX99fXNSjYQiSF3ufRtrLMBubZA7Gx2FApplgiAiYM3xk7+klispn0J5Oh
862u/ln0zoiIAxED4H07B93CBntm1ZfRyFNmSUjqIOVroIzqTNcqO6OcVkna
JKEDEmUj83bweBUu/daPhrsjnsg7dHB7u5aIfljjtv37y7LFBXBHsjfb7V7Q
NB/CizIGDeK+vcIZI5U9jk7RGLlW7Mk3RAu4EiCeKNjnMmy5AhyZu4BtK0ni
2LG/Fnn9RejSTzIuctcLqALXOYrB6Bk0saCHlEMW8rBWJbcTMrGPsoDMGd4h
1oKMNCH0YSHjd+/klrgeogVVlrvNo70aahyo009JF+7uI6b+1vLp8lgmUiO2
xV5bMz5/KjZNGD/FuxWHdeShR3uDOYXE5HvHZxfPKWq+1P8yRTlFxF1Ww14c
h4cqxAaymg9fJMEPkhmOmj798s7+UyVLkHA5yUBXDgqyc+7hpFaKmAorRkaZ
AcQwvUbPWRWGIMbRQwoDjlvhCdZDV9eufVNXZas35k7QFDf8z0WYRPLv1xqo
fB8x3n4MbvzcTDphxUx5U/E9iaH8IBpraaK0ElK2jsEGvinMCjZFH1OhTx54
e+0m+fvihQlPe30MSvaRQcP2b3tDwO2ej9V4yGMc+Zb7S7fLS3PaEiL6+J8u
fFfjkifdbeafLCxYs5VSIA4T0LBLKJzKO/Vfc4GBi0SBr7SKLb6zPSVMrajs
0BfgKsATeb8Yl9nq6t4cQA9Betm/AnhuKzvR8SI5/p2V5Gjq3d9nZiXRfpA4
0iFoUIbMCdvbbQYzW/iRH9Zo0iuhLVRp1hRm+rUcSvKHbnPQvCIaN2uKq4fw
KN0r5niw28F+B4WyWUXvm2BbP411pjSlCJ1h+7GKmJBpKNl32kYUhC/4h2Tu
7HNU0IC3mlCPDFW0EYz3CpY+k4ltsRt3IdVsX6A27E1gXi2wNDAyz7AC0JbA
ls1huPaxFMyAxOcilH5O7oIFKboYDPgbD0GvNYG5tXvwLWW1j8MURvgIXQt2
lYYnPbMHbn2+fqQGnyw5EpWaMU5VCfoGe1WvN5nNaPWP76Jwr7U+91U0F3mo
U6gM7HQKSev6Esu9g+5x8pp/pNNKmm1CGYLiSUlRDHok2MtY9ybQA0epSajF
iavikKGa+coLO8M+rIlh9sdpwnXHTr34ZMdCxtY660huMuJ64NAQupjUxhm7
TGgkU9N3MlH5AgOyb7q4sf3Z+cduffs8phxLxWViuQFixamqeuiL/6laqSrJ
P1dPZUTuGO8+AcoSXNILRnjOPdMYK8Txyz2aaw8WTQmFCn91vQRaVd/J8wdR
rvfvop53qPqmBM1ioeaeqZD90mspHyXV6jpV54QNbnB5XfJYXDGtz/R0vAmT
VN2lDUJIWwdUUwiG5tEX+rLSruKZN+X9A6KLXqE7tKieLLRCEn/iBF6qkdmW
4fITjB7uw+B8+lL7ZDXc8Wd+MQET5vsAxvGAgeB5d0HTzPknttKJTFFFDwKL
Ck3F93YyKM2wA0UEEz9FaSN/pi5G0dQERrCZ99+MD3KvzPxOGE00t/jb1nsO
UJ7Ycak6wley5iwGoSKAYAVIFUpYhWXdNVRfuIdyJ+B6XhRxrpxYbLibs07t
j1CkSnPZXlLvpAbh1KHdHt64HS5WJTlH1qcXD5/tE3UwP6FgMxwOdXb5phsY
tBQNZfRUiKGkLcqPP3PZKhDkGTnic9aGdjlw0q71HPmKMEVifQMjloiDa7VV
SiEF7929Z8hWajf6s/Eo93Fr2KgCyVxX8hRXuQb8A8PINC/DH0Dv9X99kaLa
QAvpbDAx2J9L8827H5/dXlmw4d1WuVHLOjmvBC+9NkM6DmnrWqgHjKS4E2u7
5M7kX9KPCe1wAyn0zHW8Awu62ZVnjH+lLDzL45p4Hr9WvJ5levituBGM9Kkt
kPjuWpUSjLN2xcn3dk4a+x0xps57sCkN3TSMWYRP5ImIMYVAyAh+jwWh6518
Jg1Vt6+07ip9iq3QFgwxMqFnXWFdkWF7YbfoMTtbKPMx3oJtOIwae+XDG7lZ
3ynvpr6V+Mjq9aSO8g9rNeFJJeAZ13M8fS/BTwWWYhAnkVhzR4om/hX7EMnW
9C2JZRpZMWlfkfvOUZUZibsvHXD3tJ11Y+nNtrRoM1a9zUXzzzODDxb8R0I4
5qTYdg1XzlxE9MMTWRe/1G4nXtO7+APuDYZkOjvfqrl6R1S2JYUez61TEPwI
juvhRIS3EkdcTi382r1Z/62NxAyWmOFDWoBIrrg6NGR0Vdh1tKemDF+veMTs
cffcQHvAph1ZWQJUwZMvSuPPgys0RH1dWHlYeYXPfNYs5ka5iYMRFL0jMQSZ
GnZ9zWH5yuqmL3VPsVyvb8IGJjIlbVswiwon9oIbPdSvontPKRSfr7+3xOO+
w/kQ0d44d23SaVq1zSJLuc3S6PdYMs1mybLevzSvW3igQ58yASsda27evvtG
yHDNO396NTBHsmqg5S3HHk9Sf8D9APw+uTBmQ9wGy7e5T0fG+XkStEqTPn2s
UMO6FPxL5J+PFfvyYYoGaxPkJ0Qvo2J8HrlSm8kjd7T7tK1GfF8tXhUoQy7V
nLQLLfWUyxP10u/MAOG70T+bO2h0tGK9iuQRZ6gw8SS2ht/PxwVWI0S5v2JZ
Rd3z2Xg/57lyedEO8AhhwKv9UthmPN+v+VWCSJ8He7/qzHIXR7TTgRd89U1r
x7fbT7xMg5lpH6qrsgeXksQwraRxJ+CE8+rq7LBooS6+RsKMeHRw086GHHZM
YFWACC45g9fUDE2vCKTydvqQfnXVdpDwafwGG6hd3pViS/IFKBQqLbkyph40
11aOyiIb6eH2+Vg8FnC1CH9T9AlgLafEzmTTmkG2EL7fVZVJO1REH5HUD0NX
lkAsb+CuAZLUwPBE9Z9JjMKsrlDdMq7FlxugcH5bQTf4o9DWY97cM5/5jX+n
oL2Ndm0e6pn0Tq5kDvbB22h8BL5UakeHxm0Vxuz+M1H2GV7Aa6qOBlmQE1Wb
4hLiOlZGLzksrge+2wMedIKj3QmPiUO9s6kqH4UR8OgF0JybWzVmTOdfaWJ7
dEA2SubIfWn+FPCmNdY6SUym42s6LYMBKD+kY+3aB91ZQBcDMaYlm++1jwBO
maTXDvyWtEAIVc/YecasHh2ctkAQRX3lBxeg15gbclMHL8/Dw7b0g45fZdef
VkY1c8KCWz1Ch83Kmn4+R/APCOByV4GiBHD2ZC0JqfFof1Iw9qEH5SDN7amZ
NJpHGmdiMZdi9YbdLyxrcfjl+7VRMG/x2Yzp+/Vz9DX7Sj3yAXl+ZMzSVh6x
CJb/4PD1Ns5vlKFLrjeURhGJZoEcFYoXTjOrfze2f5M46jna5a/ik5eqwd83
ri3Q+IcbyCpVid3wIyumIK4CVDs1fkjnpOV+jWpoKTTPBdckI+V/n0z88NPp
MVlVJ09jrepQ7CpjKejaDXT0XVOkhBvLm213EOMWW3HIBXO8BPoQrQ+zmkzq
4ju3arlbuINBiXdCbmQHWACQBdheIKEHa75ZdqmhltMRJjjP4OFWWHDfU34I
QvwEoQBa135Uw0csvQc6z/Xkl57ucNR720TvVzY6kGvuxbfJ4Hbz5rbbbALO
n4DrMyxs1s6hLQB6uiHpskbGkdx0F4mMm1HYevDybz4km1e9GFTgwazbAwww
g4uPILi81NlFFkMlJGhT7SZ3WHag/5LKurNi1rI4G/TAJ2TFt5jKUaz39Xe8
MFz4w7pQEvEZRoa0idU9cCWWoYEA+fwvJxyrnlKeqWo3h3avr70jCVnhrLgZ
79MVOoLTtNdcq4nLRXGpD7xUno28Je1SCpDAzSLX6O1dnlj44MYV2TnbhCam
pbORrLODkjQ6OgmlSqM3a1bstXO/eapqgVCkzM47BV1Qt9jtwWo9uGl3aeo7
p4jRc1bkcV28aI31zzP7ri5t2hn+BabZaYLCTm808wF1E4IPPjfG13gqytIX
CHsAulLN44MzOxdSXBeyd7iRlxTGhal0dYeXtGNJcYOmhpiSKkul1DsXK/2i
GGvimVLNAT/g6EyELDNc4KVDQLWNlejyGX9sCknpn8izmh+R9qE37tgT+20/
Hm2VIxt3svWoxWxunwNZYrvRLb1fUsyX5F4HAi3ODpcVfWb6FWe9HDQDs96/
SwwIuBdUBC7a4lUNq1bIu5c4Y4yl65sFsMp+OXZ5wUrBG1mI8SPyQ9wT842h
D04anHeCHsxdMzebc5AlrjBxQ+BzJbXNUYwBKHJQUJ8Q9FxZ3Ahw4SEWZZBI
wxpleH0cn0Xx3WTqJpjrhnKMd/LYpyj5v88xykliVsNy7Oh+pZxs1tLVV2v5
qgYj6Py9AI6nPDL8v4Y7ihjSOUQuq7asWRjyA305eyOMojhqfYbawBMV0A5h
Ql7yCqCQRDTU8k54ulqb5UtMewSop9//uWX+PhyA5h97rOIQFEBEYEPo3STq
p/c2L1R/mmFktJfN3JSzOeafh1WK9iQMzj5dn0ewTw+yZ8ucPL3WEce6+D87
yBByHL3CUb+IDHXsHizwxBWM2mUDTjpN8Q0kNaMonHWZhlTmd5Fg/yJBFF3j
B5FH83teT8pSY7oGX7zPp2KoDriDJ/z4f/cH7JdHvg8QnhHxQL5izAl06wkB
g3hITXqOp0oPuQnqj6olhfqBdQBV2fqxohWH/Euy6dDpUT+mVc1qlWH/QTRR
Ttz54JIqHQ5NVcx4yCZ/J/yIoIHmkxl392Vcs217rvMqjvvvtvz62VzVLx1a
Og7WMpwa/vYFvcu9fcH0zdad2e6oDpXRMOjNLoKyaowwWbVevE+o3fNMlS5o
f2QU+V9GsHsCRsVVlhb+V8sA2WdA1XmE4CMIYTvxueGvJJlD4xloSob4CZf0
KmIv8UXsJ4PCV6N0xjjB8bbH9zKKmnlYmcjEvPnE2qVOZTErLWvKxJrIrqJ6
z0z9/ludj5GsPTNuvWSne3xD041409cra+RCCpOIRFAg7WYkeVYAA+MKVrxT
5PmylFTJwO6DHcNJwdH5L085eKQYPENZNJ0vd5UuLJoAxkC7J9w3RkAMBW8w
48tC3gDg9TwYGfTZOmE4oqRR/XtaeNfg1jxPFZqf8maEvXUJBb0H+YeCnQD7
Lj0anhvMmoAmCPNXZzBGg0dc9qWpBXECTvRffO94U8EKT7Dq4i6pH40wvelw
95esaFaweXx4QEh+Z9u9G69hIbgsXnfqTDN7zkh8SIRG6G8FogdVfo2YjH6U
ylngPzD8cfWCodSETXEQ42GxgBeH2XyUcJ1EWdYYr90faPC7TSLRlVhEI5E3
4VBXZYCNCWF0yo2vZw/dfCKP1reuJ5wZ2yqkE+HTObdrHY4vNvQ0FwwJ1+ie
NIdfBU6ByDr13ruboC+DHcLmlCIy10iRsitdBChVzNs2hS2pVrnN1Iq4rb7a
AJZpGSsfSrpBNQ26LRx7OK10pHBLt7qpJfU4C+9A8auhbRt+33ydanQhxAam
5vxTY7CyD+39hCJdsrC0kf5qTUxD9TOEJIazSfA5aWqUzNAOhwPO9tAiQ11j
5yj82F9Ge3WMF/5vbxvkFm6CfcNBQ2KbjYo4CDkq9hSeN/LkLCqSUzcKW/vA
t4cBK7rkNtgEKwmDhqx6Ea764jda5HBAnrqN+vBNTv82ZbbNiU8fS+sALbJ8
AgN1raltUqMa9fi/x8p2Q0ricwn5q0jyk++G+efItJKV+zSSoezcUcQP4oO3
lSK4FAV9xo8w35QlOIw93GYw9gMYSIjSYvePfIpgBXcoknfJYmcbH7KK2Mio
VGRQi+dxXP67GpSLbDfJ1jywDORcEffK5eaxGUkphs815gtIydtmBkkeJv5d
lx/klOLXo4ic6p0L+RHpv8/vN49cLpFb/OttY989xL21yW5JKXRfZ9aQ0VRI
kr1DF2T4tmEQoiOcbqBzYfMnHOV+ml/RQEUWtukm5jAh+cqPhbdYXesTdQfB
8Nn8w2RCnorHllMHbvaJn3b5shfpOklU0gjg3+5LjqnBYxyflbWK3SzMT+ck
TN3XUVdDL9nc+/3hM91f/wkB3Add81Tncu5GrGzHewq69HF3dHPdaERAsDtY
+3+/MYuN7qBcPbQf0f3sVSCxhiY12bl7d2WJ50xtGg/RiR3B1Wi48n3aGY8h
RISMZaIuhNVcy/kVtCOcl6EGaKb5OwCbuFxVznrO1RXUX7lCL+qnAhn7Y5ha
oFDR1z0PhpDS2t5pmU04uZuWp2B/lNKbUrhOgMCA4f3hZP2Kkn0Dybb6Kfg1
/QIg2S1aZrqqo7hdnZ8f759ej289h7rKS4d7UZA5uTAV1azKMtBRdhj2JCJ1
Cq+d4pwk6hYRWv3SQuZhDh924GOEyMffyxuGqtkKRjpzNgS/OWGx6FlCfq+C
ml7uj+6MFSUXV2WHfMHKn3v1GPtZP1jJAfOoIvcCm/tlkcRPCKV9WWBl3c5e
tP3d0uKO2Vm4UH3tmYJqOHxHxq3iLrbzfGQ3rgngEYINlQdJMwcUXvIQeA+U
u2ZcB/YIbI1ieysEUHe7/249ki9qqvmxitoclszRXIQaO9Is5V1EWQG9Y2MS
4WE6HVfpZJvZ1qygPQ9aDatU+df1FZe43uJaAl2PLUBm+GAH0zRzYzwWFnPN
xSCEFe9Irw+9BbpKVey3QJb6OtplB6rFaevHe5kDauiiOKo30d46ecGtEl8b
rgBUo0YYpqO9BwfLIEBDDsaamP+9lQRH3IG5r3jP9wxPIN7VpZIfPSAYZb5k
L9lbGAtvN8VJ3btNJBUx/o/CSMhZbqkPrLZtTqcghm410lFWmQW1icF9QTtb
2NDArJvPKM4h12htZfdK/p/Wsd/g6ZR8PfncPDnTvolwZTAkRC8FThm4pJCD
tXkeK1UnXtqdWBe8Z65uNXaTltKe9FJ2I+0cW2OZIvIW750Gc7LkVC42cpm6
o5gkoBT2xTLwf4m+t41/iEfioSLii+RL9vkX1JQ4ZLrCmcWcMLxukMuy7V26
22q/56DZkCVP/UfHuM6TgPE224++NZCSUj+x9eAzwH3UpdUxEQdPo87Aicr/
ILjGM3dDE5FyerIu39nfzzDjDWMT6aHZrCE6lK1mvIdLL/hlmPM8+cAWzIBd
A09ACGxocnH1CVWDXhoXECgarbIq6SMpNXYMoYpzf5kJnDg5EDDqV1NAQVUR
1lWGPd62/TkXGBV92uxncGGaIXcIwfihk2x3bNZ8lp0VB5rp8oY6OaWMqpKG
hXc8mRCEJx0FfMjjjcuk9o64M3cn7lLmuQMJbJ7GquF2U4Si09FCEe3jdrPd
ErQG5Uw4BAgyzZCpaxkdMeqwSqGzLzC2Pul47b1I9dx3hyqKrXPQWaQKq8xh
8Apyccj3aqHh4pafliHnfzyWCAehRF2hrE6YBeLKXQY6xp0btxtCmQp49DWU
3jw4sHrVZulfhlD3QBSminejRwHQhk+TRfftQwh3QwZ7mmLPvsq5dGKFTyJr
EXxlU66V0V7cE0vhpQz49HOcmgWqkAA2E95fK39tmm4yDLuOEDI1ukqriuZ/
qrhcia/vm9BPN6mEy+m6GQ8h2vZYxUyEsQYpGwftbE3Wl1MfUGdbxG2MJcIo
T2E84s2TxxptfM9C38C/0pA1eDlIILpvGd8NbOvkYCYS2IzXQwuggVR0ZVBV
V+iY7539II8ZU5iZnQG92IwYHqWE7X6vopMFz7eg8/I2dQuxBvnwnbsqTK3U
Cda6dzAPiDsfxBR7qlpkc0PT3Cz87ceY+D+CbPRV6BUwEUQc79tpdo3NEe2y
VUtslXYTpOUqsNkIvy37VUN+gmPReWqk0kGq8ro+oQSeKGPD8oNskx7EaxNs
diVo8kcJDjB7Y97VjIkOIP/aa4rN7Szz8pmnCqy2/MuFDSFQCX4mY+HEqmqd
NzKAQZ9adkflB1UAbe+5LV5vghUGeF6nj+UKq3J9vXP9jrg3QSPIkbf9wxrU
ojwCqJ67RryfXFfi3TUP8C+Rcbt9dDH41FTKc2JdkG14MlxW6224de5VTzuS
1A2qe1K9S43EVNwM/zPDVwzzd0xIj4+Wld12uK2H+KQTI4Dij+27XfnR7LYu
QPN7xDJJZ3P7n0YuU7hCS45TUKEyG699rB13ye/ocuC14zifthGxusOfy9yS
TNNgrZmXBi6eIwD1oAO6/UaQmmjgzNEifLaAP4Uz61GnxMERj2QyW4BIsrJQ
dmQ5HlnpdxFZ9FU8lgCw4bhJJiA9x/kbaTg2B6Prk0u8jIbYleSd3lhPPDhL
HeWVvCKt0081QnDFLxuAXn0fcX1maf7+z+pDL4RNUZrWVeaKCkx+BknRLuVy
O2HsPW5/A18y4nEY9s0PkE1f84wZ5yqQKRHDt2iTSp0tcTb/lEhD19B3rXqf
fuSOkR1IRh2ue51ttqk+ikJaAXMUkIFHaE3UH6aFY2z/9YBkNRKhBdXi50o8
nQDty4qNF4WWF+UzTU2EeGhV15CMmdBKpvlFHRBMP/ocN9f4mNXLhZQ8el26
jlsEH/1x+o8gA/dnlwTPrfaJwWGPT6tvnhZYWV2dLaWzrfr705/YAx6CDs70
9z41mNY/RQjKVVG5V/lpVMfO5rtOPk0i9RaqfkLbVxNd77TlPqD1vNXOS90d
XCMvpG7/Mh+OU8OpcxjQVkr2cbVjVxt/QOlcsPt44ejbXBztlqLxBzVhggyN
xOaLg2NCNbq9cNHvAIOXJ5/P4jEpMJ31knVgJZMLEnqMnonh6k11imOvxJvN
G9cEo25Zw9Zv4lbbciLmIGW3L7amYAVvkbLmz1SQI/sXzZ0IPN/8QPMAoFhd
OASLkBVb0MWYgkWxvxq8WWcjKG59AlIdvGrFj+oH3fXhFWxRd7e3xrfTlHF2
LuQcRqcKO1dswKFxP88RvLY7yozqLIhWTlap7XQPkKW5T5VjYGEZtKIO/mhj
rjd0s+07ePd3dy/Z8cebiMsQTalPWhC/RsxWBwJOPpdZG9N2kEkmIJ5shrkq
1BFVF/UQ2SKwhQzBHeD5cBo1GwKBdPVSqVeM0JPtOiuUeJZNz2/8nyIhYsHz
YNsNgoUzzGDdRlJLffZCh/nNS89X4QVg3oimj9Mq35RCw6emgJECL/QpTBjG
aMJeJFy+tx1Lyj5OuZQ+ldKfBy70RGO4q5bdy8eEC38gerrk8bi6i95gLp5H
lmCt2r3F68SxI6/OusuG8tCpcCpX/cEh5AAslxOUpgFLZnT5Pw0bvHkNX9t5
7JiQFLJXAZA9NJ1m5NeZfqWq9jTKG8ntNIRt4C03XL8y+b2SoWPO2LtG68u6
SXYf3K2mOlJoz0rmOwLasXw8Svr2aMkSMIZ2BCE9KzSpDxvlP+uuOvsCL66t
rWaFin6/XI5pIHqZKvUihAxYmjOuBQWE+V4zSDpBq1EgYjo+bBd8pcG+z71l
YFqzs8me/6TcH3I7dqMvOjrPkts4cWmmtU7GkQL4FCzgv2FHfvnENzNImuEN
X/YQaRm7dh0bvkNhE09AreWcMuBMkKlvvyTRbp+iRbQ1z8QsH/KGzBySvHUu
pTpyEWGflP4OJKqa/z73FKd80A5+Em6sadrvykmhdfdvjZ0yHVEUSEQS6whO
Pgy1JRwU9vHJ/PkUQN3/yC9enOkLJXr4TRmfi1jfa3ri7Mxs6AW5zUwCThxU
LDL/bqny8PCxryQIG2xMZFFcpk3eTHQPpZyg/57krSgz+7oXzCL+VXQ1r9Gh
pzW51+2VoZy63ZsosieDIbjrDoNA5MreXk2Vo4IMCo6X0LOwVkmkC4Eofl/l
+V3kYzy5wC2MIXuaSmcoqm4iiwDLe9Aau8gdNK8McgeQX2s9IGlIpPxpiTZc
tXZPBouvj6sfjDiqB/PsWyu6IxiNAf1juMbMRH7pdDV/jrOsn6xxXxFCY2V3
q7nDFu74f1FfrndTQnqCMLp1cihQi2p5bb7AvPekGkGVJ/5fobEIxmeEx89u
GReMGA2Ezq2VM7q3zPbgz2+Cn1lUGaMQ2UdGT07S6JP8DMi1mG8RPbLprDmA
KX4RvtW6j/SMPyswVfEKQPhVhkDZDcJl/h6CeZTUangt00kG4ncvfBGFHRSv
i7BpEyyiASTnyE9vCNGeaFhVJY6P4bD4k83t8m7xdlcurAEfsOnUJcrcVN1m
pbYuxBJBbo+7xXVVOMa42qqMnMBZbX6lTbbu4b3/roojq+cVFN1NNCQNB6yz
BjF9eTUsEgKVET//bfaN/LPgOjZYHFjmmGQeEapc2nvsJIjhiQUugkkw2x+q
j8M7lrSmHXNT3gT8W1p5MJjWrhTvAkkOG4BajKu1YYoFdUkHp6Apk9DQwXMf
7mpku+LDGbmGnqX3EH4G6xN05MLBYprKAy8Yu41yvE0CK5zLyC6gtWWoJfq1
jT5ZrxaAAh6MENo2RVFhs9hjnGZx2H3OvA0dYRP6igCw1sGv2LvQyWeadI12
DPauDnRt4Xr0+lvQwrdOML57XxZaDXxLszJ9voD11zI3mR2toLavRVB1IRwE
mEYFqfG2LMtRRkC7PcTu+ZAjR6nU41x+GucCYKUvVD6aKABj2oaIujhcBu7G
jG/dPmvt1Eidk2kAqKWsUq8vLXg32xWIAXzdc27eciQ4XZOgBbzSXtj+awmQ
/w6P3dokU5pfcXKvSUhwpl1pNoZsK19Vxafp4pkMNIP0HziZSD6WruBQt9d1
xqTxI0aplhYusHGE8m8CvwGy9gxOYLlLgVmGZdUMPC7D1XK+E6F5fKihAfFa
6niFVWgeTzr/9tpeVvsGOZRSp6kvGSo74m2Kssfh5F6JhhtXqrvuLLtwwy4P
KBGr87dqMcuzZHCBGi9Xh89eN2q0/7WhdGAoJCc8pPLuSlc+gMSNyr9pWsCz
AYWU0q12TEcueXdv4fJBNGu6SM7erSIlF9T/tYLWSlF9/qaXyzzp0GgjaWec
89pkN0Yi4MNyMdEpy9Seu8P2TxJWnyVVkEfX2VCC00CeQWbzYpskJc5TpZ1y
U3ViJPicjGMFF+DRnCBeiLuSfG+Y/k62cC30tEXHK/pMtpu0HvwYTAiSPd0w
VCZfwVRrOZr2jW6QrUd+asmhcXk7FpgMOJRTaD3vz8em5PLLS+iYvT5+TZLD
xe98ifATOa4nIAg+Ya9ZFYzOv3IaXc8BpTf26w11ALENnKCA6Kkqj/UL7+uS
ZfwwUmcBZgJddYhNDGJQ/yXrmNAFOVC5XBXXcHwOG33hPY1hj1WdaQPHPont
o5cmiIY4CCgT/aW2B1MGgKb46mbkcUXaaO19hVqldunluDVh64KHd5upr0EE
DW5259DlUD6fCnwyQClsw/etIt9g/mmNZE1dS8taN5To/0xxye7dweGLWENq
Jp3CTJvMQO360eg+mMgzOHXh2l79TtHQmZvPwBK6s31h8exqPsnFiVkH7B0q
QCrhctEKr0U0qVEkrW7kIvlNfUnDHUOlJtaADb4mjda5mzSKAufz6O5hs+06
EGW9ko8FmTtDClZryrF7u88evfD6GZ+cKNMYCHvCRWbPcFoqfJIkNBp57fIg
BjsxWsYVSJe2BEgf60RCQrxQlHTw0jbuoa2zlrqZ9yk7zoVtCPy7bjpPFqsU
d1v+qZwJIddfxnhbjno+ZLNhCYAe/MAShqHwc4kC0KqAOp95XbRfyv1gXHWj
hQ+6A1tTqkSqEsrVUPhnEBzxpIKAwPH8sJ2VOXsmVrAbAXhoap+nrJzwBCZN
kvIX1ct9CUcYpSqZFFRijsoTqoEXwHweH1FXh0svY7IlLoBh4v1zOUt4nPJ3
WEkJTXJ5ua6oSl2bMgM7+F6uZjZYnw49f/6zDZsuscBiXNQUsl2YDYIFpcn3
LrTNAuPHl45DZU+tM+4RinwNQDnAfaUT8YKunqEH3Us3HDGHAsxqt2igvSmx
YGYSDup71s3AmY/FiamMld3yhoC50YgwsnrWtuBuf0dendR59/r5H3If5kkD
EUoGPAdZljF2JYFkel8nFbvKTaxEQBbxiTlYvrDe7LHlX6d/sknj5o5fVBH7
wyy+bTJwzcdRHM1dGQwPTnExm1a7pgxbA+8t5BHUAFLZHIHuX4DYvNs4fQmi
W87/3QuH7nlmNTeVov+ZTPOwJRstc3DsdjKgfIaekwcLnFf16SwHrWrzivzp
aN/H4qKKDfcum8B56xE9WatsuTQq92hD2tgTURl2zR0erCcP0ItoBfEIQknQ
6qjXEMzupB/rP8TkiYdebsldveJZeDciCztGDiRQVF3ZRtPke91vu+KHo5CN
Lqg/HCK+og9tOY41+pyA7dDG/muX8cVuffit6PKzEfaKTfI4dqq6H5yk0LSi
Tf/t1pjKPx7Kbl7mxIQhZAq1ablZXLKZ/TwevJqYnJiyAbz4CI7XJOjyNkat
2b1TvhlIpMRHbBtTzk2ZWcIFa8NZmyaWydN0c8PT5Lwgf+CYwisOUJGZ6uAu
jjotMSpUiKUV21PUhKXLvaWUYZj3hd/i/3mXpC6Mgfit64d0gAjI2tmYXJ+g
532KHMnx7hvyaQg8ZXWsJynWpIsa+KGM7RgmkHs5qHhuFhMsIhlaaOhvZ/j6
IMtX/3wLZCQqMi3cL4SCIBzPIZkVE+svsRWBdBaqy/w/I58j5zcyo21sG/tK
y7RDf0yX19WDBNks57PkNLRzhi3ZxWSDDkh9wYXe0lO0xvy/oyCnMz8V1c0l
y/QrWpIJIkVa+42mIs8ahbCMgZY8iz18hPmgRojF9ejyieeapFw29XPADYWR
NiK3B3C5bkZfDBheOs4DOQwgFTOgPKvUZPlNJzS4EwupZnfUBup0CkziEGRh
pL3jMdu/36m5KlK3nPA28G0Zhhiw3M5tj0S8MCD92HnmUt4EHiDsvhb6a8ZT
IS28KvaqKqaMsbiXXiAfHlZGmtPPAZI7CK93LPqMVC/RSGTOWiGWQY1mISw9
VEK2OKmImx2mxSkfV8ppmK7yGUwJQ6CcooOBBOpXn9NLVGDu+aPCS1EJDniq
7Ln6Qujt8Cazxx6Sd9CZk4qjozM/H6EbM7WR8MzOk4krN2EjURXpTd0PEsY1
r+st3DJjUV5Td4+dOsg6UwJ0dkF2a2/lLdzn2wSmD+wCBidY1wdKrWOySAEn
IpWG2OrBN8v9frFna4b2QZLOlfSl8HeIYDc584wMLQqb+h//ceTWCOrQ36YO
b+E0HXqooGvJGDUZKmt2N3LQi9Bpw622x2ROH5oh5i93a1t5+uYMBsiF3lBD
RWQG1Yftmn7o9gw8UxohQTpg1SjBzcVN0E1Rdn+nitan5NatB2U/F0j09/RQ
pLe1BLCtB8Bn3Q3wZkCXzVSQ5zXx2VNiCORKBRTO75GXZLyIPXe5rYsjkuCF
F6aYqMepgGSav16/0mTSaa2+NgHIjvYxsTwecE/RyQroSKvbs4IEXIEzUw3w
eyZy95R8+MBJlIDBnAzJCKAiOTzogGP3wAa1E9Em08U+lEOs4aukKeO6Bk5s
nkIHlK45Fh9/7xDxfnu5oMc13fE4YOzUN/Qwo+nCXCQO3MNgTk0CSuULoD+w
36n4Ixe7/hjYPrHHPMe3lv/95zxSLf/DG8+ZTEOjzQ+zv1Ml/YODOn12qzNh
URXgz6lgdKdXNTiRzeqWVzXaIwzp7nypic/4jy4yFb4WDBCf4WAnMj2eorou
NSIbFHip69AC524/uuYvGaO9DzHfbZ4m1aQlwvpf9rGlJz7QC8hniUXgk8Is
bqlePOBjx82YHdknJXiOtu53vMlU4CqrWl0TSuQbgYiTrNATNj8FWtkk9aOB
FadfcVfxS1uzK6PeZSH5LK9JSHVOXYovCApX2+52vcqQ+A2XwX8MgHTPfF32
dD9iYYaR/7+yMEtwXG8R3w+/4N2VFr9aFvnfLVILMSPQYi1Kxj9dnBQq4LZq
xLHLIbjlkZnLNT4yH530JeOWOru/T1mmE4Uzi1udsmPa687ItAhpQA64pcm+
nAsOwj6zHCmOdefuRMHBx3S9XbTsKAeGM3vloS1TL6mPWXGDk/MgLcez/Wou
cJQfE5ZlPxq4rPq8ywvczCWBmSiIokbHk9i3knmcJg6xe4+EAEZwdh2N9BpX
0Ebw42UItiWO3+sXUpIEaHp//OOe4ukIdpf/nqqKdXXw0PnvDpFPB8tqLHPE
BTGQmjkVKh9vluSRU0Cn6SKKRAHE74x4wcPenoMr5lvg03TqZyXI3Y9XmhtA
+ND0nDW0bjVgKZoezq7GyXPuqFvS4hv78MiXZDSM5wa15GCfc2HInvK+/oR2
e3IISQXdOjCy6oeycSX3NrT4dm4LUF96Un4FyziPDZmaSLZg+t1NoXifohQ4
oIjIPyBLQvdWy0Qcy4FyVf2o+LQHBXGqSXOqQcNyaMXVi7ri31KjerwbdxOw
zyd/Hm1+Ehn7gN1CV+HwaITFqOcLGx1VCuVxrRtSuFd2R53MWhA1t94SUdnd
3PBm9oxcmgK6FaJw8hzbFBuDHxWNlHeDR1xhAcSCAsSu9coxhsKYOI4txLJq
+lRC9ABxFoD+BEX1ydAdBnfH5n6YzYt4Xu/kQEv1dT3vSIaZVTCupDYh7zS/
1CX4FyVTyyCqiTZijCV+YQZ7JmBr9a8WCDHr4MeKGzBZ7zn27N9oR7RoHmxw
wDrECY1rMLw7J7epz27XDqZWR9DCnwmKGQMYH2ocTLIr2Jls8NdsmomMCK4v
0k6hTHyRrvhHEEoeyOSkbWiKSyTOwoVumi92JKWe5yzw/PiDlBeFokXhIlIb
rP5b9CdWNq6kp8d310896WXUDuC0Lp4bHg/1kCHAQHyMG1LIale1Y/HUJc+r
hhXVnq92l+UzJFjEFLbvqzwnG5t1lUd01m56LQOQ8sfm0O/QbENrK3sOS5QP
+E4XZ23Dpxw2eyMhn5SgMIScHX7Glvq/CAR+MKdiLozlsg1aNJtFn2om+bo4
7FppyiE6u91HFMU8hAKEy+6m6pX7AusPsYRMnusEuZUk4shgkavqhfjFEz17
guhW88MjnKu0E9uksyvJFe7vBeWLJAwgvoQLLw5P6anF5pD5PXcXH4kYGfer
QOT3AagNwF0k5+NIkqUPbON9zMjhNn0DYMsWVvChYD+FxJgQCGlQ5JsE4OjY
ZZeJdpZgxLpShnQuRUNmSDyeLCQdNc+5wHojQxkDRqk8Og+x1L73IT0eCNOe
P1pTa2LR1U7DZIuedqZ74s1fQC8LHX1VKR4VhWZ55gIUxQrik6quNsOVm42o
6RHEjq+sCvVEqQA7+i3Pe0YLy1vzshP4EM/ijWducXX8HOBXrqI2hOUa9UUN
P5CEp5K0I0T6N+GhKJgVLtAMGFYR3XuTjvxPcK7xN/xO/QvJ9bwuePbm+KEH
9wy8QiYTj22N1Kz6jZ6FXwbgQDIsq/BlZkuzjvOe7OQ28YHjuoIOuK+95wQH
c7TshxxvoZpCh4vfYLuYxiJOxIu8FSuDxcjmyeIwKieneVYTeIdGlr1V+o1l
jcjPJXCRhk6xNWMp6mE7QywgyM3+ipDJmNe1zJkWjqr7s19GOKECGQx4Tjms
nk94jn2X5XLHfm3q5hxHNIvj1+VQ9djyWxO1j2zaCa+3idWLlVf3QqQTm4W5
V0a05igqo6fuXwvTArgV2ps672BhJ9Y7dFBjRfTdV0sRguj70ysBAr3S5XWm
T5PU26O1N+QxJjxMz6/o/xxTyVJxgjZxmDyNQJ8V4B2A5JF+K7k20YS7uaoO
7iIfiFJNTI+ygJaWPBupYEh1XnkIjeKuOlQjcojxSlQ+s/B0szNPi+yisAeN
yQt3IkviLWzoqveyTm2zoDTcF22T9zXYDs2c24qONSSShlJUn2UQk8highCk
7HsvN4lpDuI8Pla9K/GraeNboXXcrKwzzPA4tDgDs+nrlUTU0imiJoNRFqfW
zLg6CKGgHLrHoieEPE1IP9QRHhsRq01AIwww7WQVKTynTSw6NWaFnfFWsxuz
jvLobf6JX3ViDZOPJkEyWBYV5h4CGaxb774uJOHmX14cK4fEPRGazcGF2VdG
o2kXhTjvZKpYJSg6TtITXVaydr1S090NXoyHKix1Ye0+shzgZfsc8sYw4gJ1
gLOzR8nKnQ3RHpcVyISu0kez4+AjX4uoRC7DsJMXn5RgTVtYQPFVLr3Lqlma
iDotG9qDP2f2fYmeL91JwKqA/yOOhS4T0BGOnxRq+WnRGuzy2PUJgRuZXEmW
E1YHpDKAJ7WMPOjc15a2UvDF1yi9DL3sJTwyp8kGWgI/VjouNdquIhGXmKjr
0RLw2hQ895pq0pQ1cXzREOM1uROKvL36x/SUv89QYxoFzW/10nS4gl9zNKQ8
tPgdTYPxYXIjYfZjSNTNhGLR+ZdbvUo9rnDHgjS5FHwzRaexASgRUB4nz+er
QCXPlYZqoe+/YIjbXvEmg0FZSiznXEENoZM7HuTDNTFYFFvyR1140QusknoX
lZvceU2ScLGvc7PyCOCRBgm3UerCZiablVV/5yS1VuSHthhTdsHgFOq6UKIl
YRp6eQwPPsbSAGQ+X4FgJ/XXioH4SZCSm97A7xXxZZGf4DBkQFYua9Gm9TCt
oedR8V//lGBPfLSqsdd+Akt9QE0bC+LUEyQyRjOTgiVmE02n4q5b2iWZAaM4
plmWIPPtkHPhDf2CU3EIgm5b4+Xpd2sDgwuPIIVm4jTM1QjHArl5SRLzrbeV
B4/jTQQcAdqyNswRNzLaE0AvaZ76AGZ0o3cuscklBWDxDWZXkz8bPzYX5uUb
WOT4lsr72weDQWPXKzxyzN/vPaa1ImJg+43xbVKbq6tUiktcMbBfI3aTmJEN
fkIVSUN9cZzqVJQMC+mdBwNIA0Fp34O7I9EW+MKNS4UA7JIO9q5R8R2s0h79
kjYFpASx3+miE57IXdlNL+mO7S0SZHh63f/dUeNlHBPob3T3LVSwyR9lSNMp
VmEBOfiDgjDuWIZAaZItm+K0mBRcmmcmVS0FPluHSLS7EWPGAgkVLjKGvu+N
aUkghNkzs/sPKcUsIZDyxrqvRKj7uX0sWc/erQJMe8D2lI6CACnZGCdunwpo
P9TasRKnbdolZur4og1NzYPM/KwNPO+fB/GSdzCpHL3sSdSdY7YDPpH64pFJ
Eax5GFOhAYUt/GqFJ+A1qJ3Bpw65yenbL2AQxNPydBHWVr7/I1cGE6aoZeGg
bB0SVqZ42mjvII1ZqXQLg1IZ7mpiEf15XCnWNK40WyZg2x72AwBtNzxlyn7g
c9QvbJHfeN1Cb8Yr4sK2oFKdFS/TZbeGdathz1QKMIwTQcHiuQABAYq8iVRz
TFq8F87FjxxDM8q7E9QlHnWDNv3h9y4Lsp388MHgg/Uu0/SUmwZxhjPkwyd8
Gv6qEXI2gIidtli9EUdM1VVdEiM+u2nHmmhvbhp/IjVNPutMVSUuzJjIsIMx
8GTEcTQ8amPO1Yyc9tzWZkGM+UoHixM2a2dZIpAP2TKmxq3ipXEWdr3wQXSt
wea9joMLc4jrZlOhjkCYqkbpv6izY67ceStP1j+owA/yTQFZ+oQZWdAp6swH
y77LNX+u9eeLozffV8fysadm031U3ldqM0X5mkjsLoIpSWb/02BdsfoROxMV
zjBFNoir5ZVEJbj4EEhXV72RejfdbrUBAJWGM1HCc/QFIaRgKYhYm1BmvLmF
LPR8mhzSlxgRnH8B0XHFvqvcltAaymp9zGqHqV2nS9CMahT+ZuB6j0HeSWFM
Zyun8uTF1qpwXNGavxpcg/XcifaeOvRlwON5eOaKt2uey6/g2n3fPjZtvaxM
E/G4LeraDF4+d7xQTN6mBFnSuPII1BvPF0Wt+4Q8zpakUWx4FyxzCtXtdHOT
SwUwZ1rchpZYzdtj9SaWtrb2rqlCVshr7TYyAme6wuOxN9bwcP69qqqdWLVH
GFY0xcOf1sftMZGjKBxTvzL86oP1Y7SlkRi+LJcHgWcIExMKxase8MFghruK
PJYmOEX6CRjaC8FazBYLk2CU855p0vgSQ/IaIcr7P+lxBIx09p83RzLIwlHu
ddakAJVnaWcSl/NxwPpY/hdDajtMJAkP7iy2wYB0gjnPf6yGkYB6EF1O1I0p
nNJMBijGCqwIpER76e+CQ8QtOtApWi1H5LweWrM/unOSziBbxm9ehXi7TbY2
DAbshbxI9KH9zHBUA256vY0tgsEmHSiuo1h5K/eQlXrMrP6Cz6KpaPT09Nn/
4jdqiv7AvwtHmfWTvK6I4nMD5cMpmLuJOqgzTzYwts8dPdvDOCquSuEAUDvI
XxkkYAm2h/gjRnycG+0w3sCzX3ri5RNNK1lBowuy3d4cvVkE6odcWgEQTH9A
pTBsJbybqjzdbjSYRzcSj8dgBqrpRGn9mFyn5qqnlvnYswmUk+jTxUkmUn5D
mX2UDsF8lZ29mYdf2zF8WTgFThrwqbU4OLFXqud5o3F9IdppJn4lkUS7as1w
s2BB22bHu6joDclGT0eOD9UxEUamsWZQuIRvmYoYXbM8g1C/mhl8DWn9MFCP
352UymcHDWpHVEfwlCCm0mYmc2pxah/nUnGf9xMIlLlJxJ/uY0S3/t+E+TmS
TB7WAdnUl2JSachl0Df01ROzkNT+o9ymzbcC/CbCNQMfr1BSLhVglaoWu0fP
oDRBruwiybt2x+ip0lEdJfKZuZWfhRzvjeZiJ9P06R02dRC13W21LQ1ao3vh
bxnsVgIlvABasVhg88ZbDeNxtiq7pap6ilFJFoKJQ96KGsU2iH9mjRphZ39N
+bRkySa9QQBGYPu/ZIcyf8SpyMeRV9bZ0rh66kCa7ujTUG7n3JZhxuuCQtTB
38OcHEH8/un07vhNwtfIkp3bP1rx4m4MpXkmH5nljrEmKE9JDeDsxqBMCYUd
bBOde0UjvSJDy0rxocqDfGEgb/5bZ6lcrt9ptVw7CAEDtWctKWTIWgSZN0Sd
8BdCbHqsAnHmWt0NbAETFjWtqnfk2pRXPcqS38I5nqfMOp7T/EydNR/tDUVg
9+WCgXqc0XhSCF1iL8v51ClDFMw7WbIkIg2Z9YOFzA83vidyQ162dX06/zb9
fAXK2yqlV8NH3U946beTe4fNY8nwPaMQW6Ki31NSE36FCMiWWU7+4FxL5+2f
996yIbxcuuO9iH+BAwVmUCAEocZWoG5QlAZFWIlV9gIDaQ9UmWoGIhH7/98j
Xr/i3RdLs+drLizuFRMkBofIddQadnGH3e9gUo+l7evs9bk522ZhnELklNax
AVQt49gwS+Y0H0tHsKgEJ0v2SmUtUCmz1WVJmCCd7e3FiiJxhsefvsemCMkI
UkKII506n4QEa3vudtBovKrbo+g1jRPMWbJulIo1awaOdl9o+xjTXQowC5nO
KmuxEeF3zUQ/CqGXY6J9eoJtIdc1vDFgCFSLa0swhZLdHDdKABT4AAadwqGp
FvDxqEFN2MvBhgZas1Vv1W4aiFesWZcZkqyi964KKZmm4aBhcEnhvkYm/jvK
nRacX8+nOtT5Rvb6U0LUMmFW2Mkw9d11xfks8jm692XfnsTNWE52fbNOTJ3I
xBNFt2Xx6ff/+Wy5sWNKG4HdqkNt5QxS4acDwlq+kByAyXdRBXlTnubN2W13
uNwHdJmrt9kooGtaTshJoIy1KJupQ3bP32N/giwuDJfHlURhq9MqYU5beTVj
+tDcG4BqB3wk6CXBRlb9nAeFqk1A8fuWUkCQ2PiyFxTiYhQaZrfze2OjUm07
hL/i/Iqj709aLBFaT5loLhc2SXMn+7rXbetI2OTsy/K4LG4mx7UbFvJaxKiN
uLfVtEBQs2tbZZgDA8VHF+0HoTHBJM5vkqHZqEdFcNs0OdcO7iwwRt34cevY
sKyJ7FKZDAzDBsGh7J840kLBU8JDk9LmqB9uTRrrUKumLYC3KqibCn/oLJwK
PZIlfxQQ6y84WkLLUeSRTQT1cIx1QDgVFlVYd2rnode08Kefr1/u8Pwu2jvT
HChOJSICX1Y4PdsGns4pJR45momGybEK72m8/xK5rePtCqRYj0pEJhnhcLzm
yz0r1w3MXpykAKjdUjWuD6MlCsOviEjqQhaTtodEYlP+QMCxmz0DsWmvU9R2
XVN6To3NtzKOnqcZ4SzN2ssqyag955bIAMGYnfx0+OIBDIqUIQbf0nYYVMF/
Pexn1MQB9tLdkhnTx/ExWPziIFAldyp7wrA4AZFY59X7JBNh4a2c1rQdIUFX
JpbfO0TL5wJlLAxfvO9pgh4CVr1LwDcmUHXizrqG2fk+7jZ2KMDzP/CKWZlf
ihTsmgAoPer6t3HmjzYIYSVfwVWhSlWGShMy4Fuc4TvZbM6skd7PMs1eul8N
zVJGthkWJFwFCePAIt5I4bp7uUZX/Hid0IM94LmH00RbDU1sJ1QjRo7Iy8DB
x3eIrlYu/h8JuzG/1oesvhjuNYBH6VK9lTsE0uTohAHCCK10esXEMmOKo1LW
3Jt3iygzUxPhqsTihYNXLZRr4G7LtHjmlJCv5BJ1Ot+JjeDgXFuR1T6yYdYD
O3UhKv3t1QxWMpPn3F/NyWRhnxvKeHHNj7fEOWZFJclsLHTUrHWpGENAuJOv
HLnH+932oAaHyFQ2h1NLfFfcjqtqCS2eUW1PYzJsMXa+o6oFDBn0vdDwRmQM
B258KdpvGF38+qkbwu1PN6QNS7iC6KHDVixldwGaVq+PW4ulFztL1omwzeZk
Scts/lZ77i7AvnN/3/RSsqJ2VP5nI5yD7Ak+P+rLtW/2eUHeLfKx+JwgucP0
GsrSIWh1TyAT4gZkeKWjMtazEh5kBTAxd2/EDTmIxu8w9PkT1GZAEkN3lL2E
6ZPlr0K4DxzXGgEz8D8XFCLQMW0STGxwtQ3UAzjJspmHahdWIZgsA2olRE4G
jAqgMAcq0mQ+A8ZaxQtfolMW4Neu2NhCDeXdpT9Xx++vR9R5Z4JC1NhGmsLA
yHpKmNopIzC3P1SIPKf7NmjjHrzdHtPavHtnLKUJgK40tMC087J3YfxETkAC
3jRt129d1C6pmR4AOv9tQ+rihUM1mdChYg5c7n3bb1S6JjmbqgTLxAyv/16J
IjHD0SB63RQGMwDNqr8Ey1wE9oJJCMp+UR+qwVglD3wU/5uZzKX2Fm4Lunm3
fN6R57S0AG+rbu+B52dgtw8WNSDecDJAuplNwtKlhXE1jG8a6Z+ND2WWmPw7
F5S8DHfFBWUP7ipJogFGFna3gfpiMUAyWpWfHpXJxSptjR8j6JsCHV4HA+qr
180tWDjSE8JPuokl8ih0N0HLMKAZmLeegmqvuFuzI+TeciaHpsgEymQxJwCG
4P7jaMldBgezQm4o+HH1J2fWTnsaAutbq1C6GasrkibhljH6SwEVIV7tjt6s
HR4Bkfwg9RcrH+PFH0J8NpiVo3FPOVBO12ZB0mYr3LCxYQDYYuWIWB2by3UY
tXCZCnRUFIePXJyZD5RrIP2SFTuDQTGFJDELHCEa3LnBym9jAHFaZR2QYcld
4HJZH3baJAZBBwK/XxUaJMSxe/ANP9acVhD6aMN4hqSsmnjXAIUiuEl1t+hA
BLBpyKBY7clxOJfxl30s4Zfn3I9x6SjmyFqJsrNvGbpXrVehpjOYyr7Db+Qx
414mzWEzmq5Lnxl0uDuOBRCVoMuP4a88wx2OSG33zdmYPVt3E3cLbzSzL0Uh
CM/1TPdv4nCFhpn5jbEt153u9Jx1uOFOOYM1ZJpQ54jm3G+9JQT3sjynpWnA
goEj+khxkgHz1Rm4O4zBMVyUN0/X9tXgMV/1Z2PI5bzOESDmtIU/Kv2yDvLZ
O+6MBSJ5Z3t1w8htqVenPaBB1NHtvs79bcLn3lFe3b9owA3WwmDjqx0Axul+
WhkVv1GN7T6fGpuzKLafkEfIkjTkYshf0wHPeMuzJQlqtDeuhpYfffg62IkY
pmTYuSwaOtkf0FMAV/4vlGZfOSF/9v5RYgaEAMOjuAn4z9XDP36iA+G6O0+4
NqbCQPIslMSRcJtSGoha7L4ldIKE+fV1tm6JwbX1dywEprVo1VtqxWlWabTg
cdW9JxzZImZIt+jvSgnHcbOoHuU6E/kCD9L4uC+6yhCbYu2o7xzODVSZbBTa
psk511qC3pew5AaBGflXOeTxWy8pWdZESksNDe8p9v3hsNFEg7wTXdTa6eEl
rhF5YeVlizrX86lX2ib9wnDfJx0+qVwWVG4xjbVUshKHuE7EOkY7+E8d2Icn
CPqiDG0B715WepboUx52/M76U6ZPy5TC5KVES7Zpy3F1NzPgsyU8GnkOqUuM
gi51xHmXQDs16l63OavsTjjEkQFTY9+0l43vu04X9Ev62Bc+xCQDU5S5xvMb
pArgL2xHM3avkk8uNXqbFHSAZunnVpXYjq+qOsa45VIAKeH0pNZD8Yoni+/J
zbnbbI6xffMO1utdp0TFl+Rr7mqefnH0/L3OC7QHZoe4xw+u+arNoTJftv9g
LdnglY3e0Ba6DBXgktX09auqp2Aysy/M0obavNFceLKynxBEgdWJfo7ZFwLh
G4TQKEIY/99ZOT3kvwa6N7oui1gPaKh3Mi8CFSKmlVk9JdXS0wEbu3K0bouZ
6QGXghbxXqM4vO3HLtvlUXmtcl3bRuVUXOtDBSgEjFY3/EXmdPAHXT8FYYSm
M9aweO8AUPlJCeM1rMAYf9w59KZkKSA2AX5RplmUXuNWpdOUqjdPPgvhVzvV
4vcVvUUwFs+hHC0VYQJE7R6qZqHe9lfVxW5jcRLsTO8LL4OYVLWXFKn3yaoO
YjRjd+s4r1PMVtViQdEuMxoM6nn0//ccsItojSmB4NoZuqJzkXIInXQvnSte
EXEN12s5zpMDm9p2KtYsnBuQcngj4hEdDCZ+/iOuCQaEm/BgpVVaKEmIxkk5
6C4CHyIMkl641++5RwCd9cdAih2Pnq+L7MN1YIZnzCBvApsGYJhbbHfWfs2z
jyN5NfS0oYVKkL1NSS7EJcPORcxK15dT+eAhhlbFrHKmY1D5eUgkGGSffSLC
IRZDHM6ukRrQmRmdOAlno/FZ3rymt+NNjqKzPo/R/swY5lF4W8yvxKizLQlE
X2mV1Inoco8esEjL4qhZ1aAfcAuuqeSJQugBZrp78sMBdHYrW/Nv0flkWjCQ
O++bhWuJytAT38hV3VuQRAAR75VMHRDLOvRozrdMo7JSizmBYWlioQTsCUeU
bEaYuNFBhSwovlUVcjVAazX92kTs50h62nwm+3x6z2Gotn4MnjzFd7O3UU4S
TOt0nFrgGA2nw035uPWHLy8ENSRGTPlpQl/eVPnQmh4/qAmL8UGVACvd0xMJ
mreLWJe+FR+EXqrvfAY2ZppLIIx0/KawBWYczIrANKqv5RbKB5gaVWUbZwJ8
kRUKfrd9VscM1Pb11TsZy/aGXcZiYgrFSV5ECYstG3C2euBd77xdXQJUJGaZ
MJp/479iFOCmHolVeuPVwKuaLEjEYABmfg/28HClZAowHgnMtkrEp9bjqZeF
cTkL0mYUtXqwu6R6zOs6w5w6pGPW1OEp4vrBU0JuXYMjQTArsrtoHYa33b28
VanqCwtEaPccb7tA1+W+Uds5KqnqQVTilX8YVS/83k8zIEIpSp1po9H44o4a
iLy88u3SeRChtAkfg9T1lIqpjvAZNvraPHZ2PrmLtdY5vytMslOAIf96FtLp
L+incs9z/vPqh05YO7lYIBdBcWCQ+bz60JGPWvsdW8+zEbF6rW8smjjlV4zb
oHDxlO6+rfSeAyWu4CXA6bNVgIlW8T0BInJLhS6yPdBZODzCHbAX6v2o5C61
m5pwC7khJQpPHnh4+JjznBxWM3jo6Hh6K40Rbnnzg9eT7WJUremAC75agtVA
qOayvHVpIN5N6jPMmLosKpKkJx7TkAU2l4YkvJFxJTFAqPxYPHFf0OLCRH+O
u7s1acbbNhegl9K+RG0AI+kR2esui4P5G+s7zD9PjIBWv+fD8YG2E3HPw7vj
p3JJZ4A72Pu4f+HT76kb2Rk6LtBxkrZHi/6jxA2gGRGFbSNNHr0pMG/F5xQB
B3OSXEDwtCLRo7iGY2sD6Veh/QoszSNua7Jm7mD9VfK3RI5WE1TtNlBKlaai
NidYMlK79fBFea+mILurF1/ontYYgu5ADw98azcjSxHxn/nSx5ntjALMCZcP
KNtKk+S1q6aE/5JcuaMYwXvKvqee0H+FXvf+qAMzhWmliz0vbMnvzNeJF1pa
sm/HLlu15u9vJfOM10e2afyMQE5nN9KCFIZc+ipFYy4ekgXhxkb0RkcSkzT1
jZjMpChsh8s09RlkFVlyyyHhflQcQAT/fi3JpHwKnVG12iI/l5yrDj+G0Gyo
luWosVRqSfw/j2kNj4CcMxV3f9i6VoCL1Imo2AzBPhXNbEJ70L+ocP3QHKEu
cX8rCm5PIENSttRoMxl+9R4uHrRV4738w7dEfi9h+IwqP4K/f5iZTcMZi7gI
Ln2FaUnbWdQo9JKVILWUTt4T53vzw9FUmRl+yrCSWJLPUSMM8BG+C7t1gyFP
14zxBNIkPZG0yx5YV2sZmjsGMpSX14MySVDOJ5uFhG48Y6+9xGxY71RsceDz
/+nXUiIEb8Xx3kZZq2A4bu2SdKG1gAj74I0JsaVAWZriCjD9j1y3MaIBNsos
PKnm7eHOIAAkuAIcF7wtny9dJJP7+P7LaUtewXcZDS3A4i7w3vR79iF3ubgZ
tmoJqzHg7TGWfNOfUfcRHrmV7bjVtbDZjD38x/3jslQwK+PdSH3/+VZJrSiP
AhDL45s+ofa4V78i24s6vd1SHq9oEOASHhYzfS3dXwoNxdu1vURtGbjHwOzA
50SVVV7vpPhzCT/JJ7LRJDGhnAh8ANy/bBJY55EJtCEDpxM/MeMDCAtV2pnb
rBMJCrkzK05hBCLOcXXX6mGx1Nbhggz1Eh+VXdiHqF1hupDIVd4waj+vwbNA
yb+LJFVkUf0cL5dTTlqsodQCyEUjaQDzPdIboNRoHqZFosS/nQyDmeJfesPI
OyaRawDIJRJiVzw/I8P6K4QryKRJDKhOvwqLh8HGnruP+sHZtOVOL3pGkPYB
+BdozXfW0RiOff8X+4uZ82idSucFT/kEnO1WAFgs2eia/mWNVaaf627eDPxl
G2CePAOlDDD/09KfrqlggIWLvVp/JSbltkM6tn9Y451leloaW3F4m2ygWjP1
0mi6Y1vGogkk7j4RvQzKHsjAFEvVtjkiULR9+ISFTWrZk7KUTdKwSCHQtrrU
gwzWX9vYMVPVDXONHT9mbYgNei45mHHY67Z17bmm30yvx4vVNdg8HF+tzdPx
V/C+JetVbb4qsDLoJSNM5apRrhvpGFz9e37OkQU0E7nbMrZ6msPxp1GJsall
C2bvhZkWWya59Q8grs2ZLC8SwfOLa3iN/GIeKon2osal4/Ln8SK7qP6Y/KB/
HcgZN5D+MXsef4VuuQbRRCaS0m16RbYYL3gBenJ/boKm6P0NgJgWyv5h6199
LyWRRWTVHuCsraS11lgvTLqhjMW412lg8HmH4O925Yia5kuu5rc4aHfNk8t+
27qToUMIwop+WGCmEoUIYi6VSd/O2V0tDAvtHq/c6/wZsh2evT4gMe/kIXrK
OBHrxDGWPTNUzl3iXyN44HDdY2cwA7SGNhp1K79uJ78zNwxwP6GEvN7I3LzN
6AnUNy1lNCp4x1qXaYE12vM3nRIudvdIdoW+7uWTzp+mWjoFcmGUj0wfVDWd
WUUqhWsDCTfh4T6NoWZL4uUUrcomG9XW8cFSerdlzfKdJSIaWhIM0tRlTRE1
eeLObKHGOyaaPlXxcKg3Yngx5yn2MuQPoS3iaK/VZ3Vm/nmrptcw7NCid1Sd
MN2U/l0YAGsis6Yvwqm+wC5H0qeR7BL2P+iGhiQIpvsTkVuUm4DpvQz5HLyz
/aD8xHf4BN5dJ8VeeIOipKCuw7qc80h5MIbbdq41WeWP/qgDFfzk7XJlXvJG
UKiX7YKg01HXvJZU/L8u8fZYF9ne2i7lRz4jV/BCeNI9VM//giq7+EV8Ims0
Fdxmw58E5uMkivkh/jHIK/K4YsO2jYKMlG3MsoOM4aEPVp4ECQgH/LGObNn/
mxftdDdX1vZD0hNRGiF6OdNy+SeFmV+YyHg5Ry5eTW5eLizT2EL9vrJJ22Nv
b6jcerWXCMZ/PQ53RFRxgoh6dSdE42DV3c1n53M2dux9RebMx4mEM/1XxEKy
fRyZRZLOeDjDlE01I+7mtPqOUiaKxV5qclT8tYAWnNN5BRTdVSXBgDtnnTd0
nsV0VZUVOUY2uSTK+vkcFXB4f/lW174Dhp6TAWEjD1EucE4QIp5cAh4/+nx6
GSNaK9kpK6r4WNUsPDshjUanP9GhMZVyNij4HOnlbfZH0trHgnVBJNIHv1hR
Gv+UpKnmrFA7oPUN9AFqCKg12Vs80wkoisW5fJO0K8gnV5MOsEym4pCNwzjc
gXfAJCRxDBsGJ8sptEex+gSEmmbc7agw6uQINAf4Q6v6O0ph0o4CvPtn+6K5
iTJNpGWgFbUQW8Km5YlT5GzBWGjw2M1QpQJKHdQMfgCIjNBl/J3o5/NA5sdK
mJ2D77Zn2Pql12TAyfYGu/ZgEtdyCOZyvdSZ0gRljPOpkhu6fcVtmpye6S4l
uei2q13lLUjypaeIhi3tTc4hyjByHTAyHtyqG+JalIGSXHRzL8bGK/NzDzFw
qz3ncIemd0T/EnMIbrgNCGiTuSE+S0cTRCOB4mkeEi6F5A3GlwDlNKKLmM+m
eVj2qPQ8at8fj4KW5bPfYlkz0i14lmWVIMpAPnsviqjjDjQNwYthWr8FQpsN
QlyuPAb1HVKcIseGbxfxFZA/7GTb1K7wDnCFNpQAiQGZ5cRpnQQSa0Lq+zQj
/4furQdhRgO0gr7fPFo2aHapwDCjIXAokMbc9ZCkoy2KWKApJPlL1XX30LrE
cyVS9HPeub1D1QNO64/ALasVrKoVZckwDXVNqvZzbmDzFAaBn9Oh+XFzpVj+
HEwtOzjwk63ptxxl83tkNx2w3c0nlJ5YcLruQEYBJq3pc9RGKZ/DNcbM1IoG
EqcHS0fNS/KhCZ4TPlj5ZXjvL8Ye563e5Zr8b2Vt/BOtuOVtyTT4kIhHL9d7
gREOuK47M9OxTStMhH4JQbmu6Ke3rIlXkIz39cQw/aFF5LxYul4BC84P9Y8S
cHcSfa/BIr0N4D4e+TH9fgNrinijYUZ5xJm8gLEz7b32nNkkNHUlFlIHmCLU
zqIZJJgk+WEZu6lalsOy1pMRnCmFFovlTDAy0bKEU8Wso/Ao0OXmjGj0Kbq/
x2x6T0o3q7RrGKCy/GYgTrQUmdZAW9ATUELXheuf5vy2qTPYIitGjelf0dyn
hogin3qvjZaUyII2H8BowiWE+xbOvUP+YA6BTCl/sI/OR2VOrt7Kr4Hi0Gti
1jOr0kyXl1cOXzh4iCVyoS5gGRpMRlu7yUf4ZYmhukLGRUX6WxR1ugOw6kOK
G/ggO/RurU+WutD+LYjhgh23DKxIN/+uYxequtRzHATxofta/W5SJCjuVgDm
me+CRMJHqRog0iRnuoYT338Rzu6Xe+02JZDPgfhEt+iV370jNsm6toxXObnq
cv8cf5H9RCr9ls1Yy3Ti0ffIBVMOx8OyNkkJ7Beqm3C2Vy39klU4g8cqWPiR
W6vN+ZXGBfmsx+jLOlk3JPQ4/wVngFY1WjVwO6P8zU2auQKLkXOcFPo+Qw6m
nIonUgr9SCwO2o+jSP5EK2v0OCqOKDqqnusxkhawRj0Uk4rfCW/U9cd6AYwS
MHw3+J6EUMAx3KkihWg4uSPXmXr/MCxlbsFRn1Z3hGXxRJTEE3pLlXHb3ij2
PMQSU8V55nIO7Hbt1CrAVBEdiL8nY08NFW0tjzu2UzVuD6acMosGVc55ty3c
sR0HQwVpldEmTZpWRksyAOEq7PmjKGXBS1pvPiXmGUKPc24oAAeSdnbNcHim
5T6VNENRRDz+uEXtnY7DDs8Tt3zxl9LzY+Ad7k3qbFO2ZYngs8PRRHHLkEZ+
CCskS1Vm7W+I7TnZj3nF6JiZnjp1VVaExs1sv8euIGGZqNPZYZQ+Dn1zA8z2
bKO8GcgCtP3Hx4tqch9Q8AVfEG798JQ+p6I1Frd5MqRxVu2GKPmMmqcHyFEp
8Va4qss+NSDavWTYtRcFZ8bqpmB1g3OjB53t8osNAIA3BtuC52Oy09vtc70q
mSm8jKc+s5v/HyttDw/piDEGb1XIqcP5CvzMA5oJaFImSYukSbfXa1ggEcZr
UZVVSKmA/MdhJwbA1lByMGmBsV4xj9np5RB2i1C/E70kF85iKwQLiqVl1nwW
hD5LYZ/pCJs2w7liK/CK0QHtMd7iibeqrWmAgFpOQfDxADWH+5NQcXb+9sP1
Mn3/sFnV+3DmcCX5SGHH1lxacDmrP0qo0weq9P4dxaMgQOG3NS2QP0sB94vI
S0V6g0ko0GXXQ6skWoxy8mIkJymDKWM0P5esOUbk5V8z7khWYx3WWeapL0RE
TdL7Et8EZtKhMICGBQOdlpnsPydpP2cXUVz64UJsFyWCXeZ+gHoc2TNJcP3r
ywQryWTYiPmmXJE+S8pPDdPk+HSni7wS9O9gMmcd0jv185bvF/2ibXJ8ayR2
AhH0qu9lmxij+G9oCy3Bp0KhVB0OxAx+H9b9gp2ZWiqjrZeD7PhGWrhABsx/
zUvTAHmW8mox4jB5FWUbQIFA03it7xgbGKfPaOQuR1xwOd2sGCcJlVWl9TcI
nGdGtPLKHr4ilkokxfDxKes6WN+PkhBNYsPuQenjztYyoqbDrARml1XKBQlv
WgaM10sBwJJx0TOilNwd3ea6LGyoml2wzUrbp7p0s/QNSOc12tOiStCPk2PH
6lMTWBmPbqR2otge/ITrx2Gh5jGnDO0RHCAt7NixT4oj5UtpZ23CxtI5oLx7
lomx1bIdlkNSfgbjRXrsobTyRLFnw/mlumI18lc+C9E1V7vDCyv9sgCeJQNa
BU17tMW8KX88jbHa4Cbse0+QA7lq3OFNpmPhkHrX6t4MGFcMG8EWn6d8yX9F
dZ0hrbYEXqm9Dw07wCdynzM9usvTPeu5tdjTzxSWN7AraeqHjoIKWOQOhlW3
8Ife2/puHlhb0jsAKgO2dAClyfAaGb4d5oEv2pCZA03oTl5tasXSmGg7s+ze
olWn7mGtg6VfboOII2jVxFZSTNHrSz2xE1DfqFEtkhA2NHZRDUz/5DGoVLbE
vR16EhYWBZ/Hvh7G5fnNy9Ppth0vGvmuRVhn6uwEP9EoCMVy15M10whPSMGY
K6I+SC4hGQqM92zsHWjc/gvuL0wGMstqL3vWSgPwnYoGVyyxIqX30AdBG7Go
vj+pQe+1i8flbQRJJtHgdBSxH83gLlVwOJ3OKrXCwCR6GgItbFIC2oZJhuqH
eNWDHfFUd++XuTgrBxWWBnXKQauqJo7U6JryjP6jcHaI9Y8yrBOB7VBOQ1Cv
AUSWfhoKRtIBoNd2TFhfKmQ8cAKIonqMauqfSv7fbjUmSCfdbxI2I4Cv8TiE
YvDArVhbLU4SxF0VL7hZCyL9Tt0tZ5wKGRjEFex1KrSm/K7cP92+GWVOe/Vb
iw/cBCkMF87Uvff7lf6GJ/Kx8Zfn9iEBraLAaQ5s0aMht3nRkHcFidyii8Rm
ZAiN2ZR/bXuWjUoCNHo+eBPcog2LaCrieauZ/d+YR2KpF9TbAPdHbfg+vlO5
AoTaQpvHDKl6LHuTJVHYNvZzarnOhA1KAZwCbdL2zKPIE3phnMQSVkz2elf+
+XZyQu0Hq2rBz3CFmadsmgxHdMAs7HBOlStwCzmhjQ+mNOz9mVThcQUNKtvS
5N0EMS7VKvZ+F1H8sa9hGYoBpjqHbTzOPfno2+LfT+5O6KLYCZBqM67Fu7HJ
CiKizOTV7yy+rKuwVMs1A3CEZ3WHC8NUtyMOKixkKuxxWcpMgU2TM8XIZkhU
a6sgY4B83W3X4xU8KS1jbO+aYno3AXaqsU7WwNx+nAD2UzRegma0aLxwT8mw
FHYXnYWYoVWswL7iZKCHsnoNuAqrsVAZlKRZqgAGjcOsFbPs29U9rUJLplhq
TyPcT67TCa2t264TQZtvuLJspJU1AQvhbsmfKd3Xbw/8u5jvemxmY0mdMCnB
wqSyu9AZUbT39Ttk8nxYsTbSZCbD4BPe8h07gc0Kfgk41OV0U6g9hnAPi+pb
3+tqVEUCCXYyfve++rSlaUxGzfIeh8LlPncb7ZBnYSLHX6+Sl+WK4YhQR1Cc
21KH53ueHdZKuUt9jxF2xN6I26nq5GXP74Ai2OGSyPXTTLwvRpwpP8azhIGM
hrzCN5OVLXhbRz9ubc73Py+2iccVu9sSKTgcEfnk70KwHQu9ss3dtBks0wB/
osLA5+H+wACo7Csk153VF2FKsSnPqCfZ54LldYWiswfZkd005qHppUOiK684
+UDY+xuMUjkj3xWKOZwhczSaTe3ENz/X1s8VfluT0ZE1N0eSTbqWWvDmYKA2
A1pbOo39OCxrDvJWH2O/kFpz38X1aCJgBnT4IR5ZxBnyRZksFNY9HE/4YU6N
EIuFFhz7+6gb7b3Lqe37vjsPFurUB8pAVqBuf4UVKUisHMzOQu7aCR6eIfym
roFG2PsYELI4pB6i5soOqjDfo26gUArUDN7cqa6JqnYW76VK0jmJdjIbZxB2
dcxQwZVi2xaBh+2kedI9q1F8aVJwTqLJhqVbLuGJS/7xPVZxCIREMAcq7FsB
trkRcU2FZsdm/oYbNosuccoV14nLJxovZpmdG1bSJT/cbSBngnr/PgkgIuEq
cbudzfF16Ztb+wXLUG5fDmKUIoBNqbCesOXqMc7SCWNsczgbrlRkNihHw1dO
aw/jqrMk1ELfwpmiKSOWxgoKLJ8fcY2y9+U9OFMUAA2bpRdvrzJ9Y9vHXnbC
Co8O7VSQ/aJZmsIOIsdkSk0bCr4S7kxp/bTT6MlFRBJYoAIWKhLmc/XcOIap
5gXE5UXu/EYq6mA9qcWOXmj33dN6VQUVsBSsj05c78zEplbwfT85Q/1BS5zl
i/PGXitJ3Q+5RVb8Sp2OfyH81TOMj9pJN4BGkRGpHs+frieV0D/jD1BydYUx
JCj1hINpxk1MAMoMTw+YRZXLa2hhrWUdd7vbpJuIlBnYClou+Z7SycWC8rgR
Xojae3BN8GY0NLVcPKo+et/XV56Qbnk87xxYePQxjEHOkC375Ga8uBp1OloX
f9MfM+rbsMbWo6NZ0R95yK1nRiDC4qG0IVCqdTP6TUD9jIIUgJUlURaf6Pvn
teLOAfR2MUwj7JGJQJSx6H4VHGOzH5VrFvNfs28dz8+C9hNMMho9zIUrSocP
dyGqiYF1vkQ/2+hmqi9DVQ4ZDo7nJ3tvhAzJRvYmnZB643guQvOamYybX0XS
gtFwhBU2PpvIKOwe92E0umSI0DV1hOgNeEq3JCNoRbaDhJMPtWKOkX1SsDfq
rQuzDUkvwS5ux1TcHU69LTRwXspPJAP12wjVcOQSN353M34k/VQJnYQwNiwv
xh0m2XImsnVxMGjaktSMbudDhqgYzRd1ujiNp5e2/L7YVfm9sAflz2fuEwYJ
01v58mVo6vLpxht59/F6VqCE3Dfl2GXCazN3+K03eped8TCVx1sOkENIcrdj
83LAXGYmC1j2NryCv905CzBztaOsTCDtFF8Up4WMUx63gkazOWS3JryKfwEE
YFsAQWvf3JLNuS69SO/RXycEyyz4H/ObJD0ahpVrkPnsfF+k5UwJjrCoA19g
vL9REPsZMIX03Za+zJVNc8Fxv7y/Gv98m05vCT3taJtchVCF69waX/i5PZre
9hC39MeEd/wMRMtYIxdIrM4lxJI1/DZCOSKJGdh/XOwNveoLOTNVl+PA0MX7
LlUE7b7Dq3k9vwdummCLTncMY842yLM7+AecUFltq6Yl3LNHPkLqwnQFse6m
p+zvpFw6DNehh/2vlFgQ4QNIr6/V7QFYs2yox/2ieO4j+Sgm7gJBxIenmWED
C9cGHPIxbUMUyLwfNB5F2+zk0mcHcTA0QGDXCjD/kkmfkblf1gmuP1LSEk6/
uw0ZlaBDP3ZBlHwMkwZ9Dexceb698ifIudsrnV3q4HwhyO05mJ1x7At/FBOL
EQYOLeJEmqM0PcnPQMkCWC0lD44g1I/lL13dkBPu0PYiIxxNmMfnA7p1h2/Y
EkncT6fxv13Kh6EHpG3D4iRovOfiasdkduJm+br/sO169rgK7ZogBiG+HA7v
lSo167WlLhu9KC9F//unCCutH6ZWK6zc8OM2l31heEnc2H3CMNkG9iPUPtwp
qGlqT0aTmav1RbXZYc3aXuJRMQ94Wz0fiYWyMOvXgM91lRcfTsE56kE2C3uA
mzlHDwiSYOVVE7PyGlRktAHtTFMWgmTxvAmfp+s54SR3o6DfW6RlWbozOCFO
zoqk21y6FrQLQz1rdPwd5O4H5obK5HIA0+/REPu8BFz7rnyNJeXE/oW83AmD
6U48qrVMjD2uoapUaehyTje3BYfyezowIO2hqIz432Gf/EVlJqmK0BAZLa57
mjCicHFT+W0mMf5gJ3oXokfOUIIXJdv1Np8OFUe2keNnLM+wJOuspREMv2Hn
7VAK4+16j9yLtBQIDYDSqeEuUAv6NvOwpHmvdZ4wZVrh3aE2wHfEIv7pgx78
mOXz1sFOGCP4I8+GfdvdkRAdkQK6PU/0H4uzg9Tt42/37CQd/bgWpF4APcS4
0xPFQ+XYBV7XIBmICSzQ17H6XzaAWyYf9nEtAAxb8FqXHXOq1h/7ZfUpYrJl
ziexsU5BSbaMmTaNzJ1isA7IEvLdWrVBrV1Vx0yGQrnioYg7nsexHYpG2+rZ
VdL3dDvGp3xA0/V1Vz+OgQFphPN8eoKnxn+n+kR1u2PA7XRDCamXhIgUKx/l
e7pweRHv2Ut6tI8gr+QYekhCD55g8SEAPu1IHg87HffYwc8oZCcwDqeeh3jx
yBbQnyb6dfCapHPBBk6dgwAMpYcYiUXpn8ZZtWC3YQkb8pgfP7P9kcBiUCZM
dxn57iHEC5q9hLJIQ5Od7/UhYKxAlfvdmrzmvPB/ulDrSWkDVYTIQcMWQUh0
h3orvApPtpp06Fgu3ArRYyNYXlmLmimoj2xFewwSm7VUo/HEp+Z4VXKvdBB4
QOEVkY+fct1DP2mk5IZnx9WtleZTgPew7TE+NyGq9UtToZSzF143L3kkWgWZ
M1H+v/wfZLds4vxd6IHKaBjTDAIHvhHTAY7IyENbnrrkVr8xaHRK2BE3N6Bq
GplTaneIu7yjxGyGooE2yD2W3mLY1C4JkjTJ9x9LRuyAM2+5lQEF0IztSKcy
vcc+JNf6oXxwNhzmNwGtL1k3pOtMAZdd9sPq2kVMl9ActllyD/uNYrEW4U0O
2qgShcL4UJtcanuOpqKP2l9F3f07MZK/wpmvSMYzSDgH1vYYQCrKpi4/JW1E
HcaAwjkLySQwir7xtcU6zxJ6FN+37bBLckyC8XQQQJzSk/sK7jypWUJMInIU
lVViKHYLbaw4w+0ol5ukFXEoRV0GSvShoQfKXwDcqHLU1mXK4BTZ4Oa0T/zN
CG4rnn36gWq/iuBrGK7CxmjOCgtzOx6bSglNY8/RZ6+9urmlGdBiC0+D4vCU
zfFOpjLGcDQfqJZCc2gEpSt1y0AhjSSqgL3N1e33j/TOaNDd4O9XJMGrGpMA
zLXlkdA/kF9GXyloEncgMqdniiLu2OzcQFCvyE0Wn+rJnXf+/zPyqdPrICME
2hv7zQMTnY0GOQf987jnjzDqEj+G7/QWrhCyNhAV9ydTtIAdmf5cqhlnuDzX
g8NsZbm3K//NxP4Jdt0p6OJyG9ItuFDh+/C5cYDzsdBK4mLxd1N8ZilSUUrf
uL3euJ5T1ALfEaEXe6p4SzZmgf0Emcfs/vS8oBpn9WmMC5D2NpcsmZcBNDe6
gGAjG6WPC9D1AG5OZGX+MNphl3czHCV91VFPaEqCkM9qQeoo/w529FXDSRfw
fGiigrtoW6TgKcPtOqKNLvf+4YjPX27qtMgaFFEpXmcGwP7OtlXdE5cApDIW
yv0rwgzmTp1xp5V5vVIPXOFaVYVOfZlHQKKygHEGMfepj3CWaeNcHcWmbZmV
XYyCeoMbTsPPMPvMbGlJbJDDDoY/Xs6rNCk7AAx+itVOVfmaEQbrvnGU01pe
JbRBlWbvSeBrVra7Nd9QCGEm6kJu56VKafZ/WANpsvi8IhQFHA81U9gplVfG
DXTA/Zrh/rUs86YOeQ4M8TosOk3lUm9kilrJ+3AHfCE6jbQhz1vdDIhQk7ya
kWZF5TL66v1JPMHGvJGcqKT0HeBj0wVRqBIluizQq8XiQNexIJ1rhonVq0Pb
MvYHm16cxZJs6DuSu6m49d2Fk10mcp+rBQEGF+XGI4pxtan2Jdb5dduElru0
uEHlYmLM150p6G9w+F5on3InbAlQjwm89tv66a419zq7j6GRGak5VQ1Bqkqk
nlG1oBj3VCJcrBko+iOCobzhRfd3pfiiNb7W3wExgdXBM3/IpR3H1XtzsWmZ
JdKMrUDMu8sSHP3hqWOOtH9JdhpfIbODKDnLLRhwakhYbwSL8t2qtGX4ot68
0LlaumuUG5PfkRMk+TnvcdsCZc1/sXqvahM4TCo90tWxDiZQ/nD8Btwix3sk
w5dSVIgOXHwqBZqB4Z6gB3A/5XYhyR2vpSrZVdQEt0sRWC3UQ7VBlazoyN4j
+ZrZL146ZvF3fLdarJpmVu2HO+Sq82dEtCx/cMaDIprwRphGZ62f3hqTzLAO
1iBADdRCKeIClCXO3MqMV0ZlbGW7x4cC23LPcvNAnv9LhInjWF8zPhv+Me9q
SmeaklNejnmmNpbRAsvd/WEqKT4rFiCtbSlhvEXtq9L0hEDZtzWxSvDaJMUb
5qBeqcAwvFzvOW1dRPPJM+hNgtVZXX5gTaQxgLSiaRRp7jG9k9B9HJDmoHEV
5UeD+pJrfP3TIQ3X+qZFmdqXKKAz9f3PfUhyY5x0FYI110/NumhHbdK6aDJR
jMhvdMuhJi8Gi5L23+UQNFvw5kjJVMCb7bQDogObPtp0gptJp++baK+6SfZm
xwrKn7crVNXn0VYSq8yFQ++QWypN7SeCdMamoJI7BH+t1Y3ZiLwON492vmk5
nQL4iG6v0aD/8OwdgOYB8HoFcrwhNDEIg7miAdJxrhcWZ77qOsVu7zLFstCR
qastSZZ11pGbpz9t++ddQcWzOsTArHWyUxvaWKzG/uRTTAin718MwFl4KtSW
PbnASE4CxOhrj1rysvAfc2sRdsNT4Qc82U3+kyfaCo+BJb7i1a+Y9wPx46m1
DwYVfyisEK6xcC69eVl3hfHPbMidiwfQGmEPnH7L6Vq//EyUBmHqDpbsi9eb
jjoL4JmDiRW3JQTD+atm231jcfpCs/h+VfnffQbQux68RWy7o0iWffQ9NnP7
+wuv/e51ilhEtRmsHL0Jc+TcKLnosFExgMEMvFtSrm1mUwE2r6w6IjnFnaDL
oTzometcCzGAApYCFNIqoczw7ZC/gf1TqZZ1pH+nBYow6m/4Jmu/2+d4mkUH
+EhvnOtw8J6NdE+DfObxGW9xyVrv2ZIYjyYhmDa8mgbtuhntf3tJ/jJGe7Sz
L2RgJN3l3dLu3///O/UjV7Qp2t4sH9cMKYbzUtdQ8fW6mruWVatYqpvjcYoJ
KUbbLMUStg7D1+01KQMecNvd4XwIWhdtqMM3hsWOyX4D6DgV/raA1zzCyfd+
u4qdpxPNPZwW9t6JEgKs9pUa1798OHGWWonaZEkYp0JPRJ4acE1sEbHU1wnM
yWr6rJuL0yTCsLtOaDQ1BVZsKSOEEg4MklR38tD/KDGSMgfU58m9cjHE27yM
zCWFWrWRbq5oto2HhMOEq2MD2TfEv6pWf3zd4jYqN2V4TsPisBN/kGlVRqy6
AMt/M9mDRol8HDVXpLMe+OmYlIqFrHWAV9KpOoQH69RFNMGHAGs0qXZzRHaD
PIkQ5v813UBzZoJaBMF/TW3jPCCc3fcS6qhaYCo9LumIlCpQDhCUkDT1QE2/
ImU3dSV9uksOJS3hQRBf3hlfFPlzvt7epyUXP+10fNtfVGXM1D+pcW04w+Jg
baIxLABBA1/C9eu0rdJ3o4mD3PktUCV+etcXV+iyi21GH6waDaoOEd6/IaEK
1WS0YWD4bUrhMFod9OGiJzc9H9oe0oCHqZcesQS3m+/tMkXkWnQUDOU87tKu
bG5VUG9J+SN2DMxBoPnO26KFXBCNPwcOFsF2jMViGdtr6v2un/OPU0J5M8VB
w4guHGNfbCr65ODORH7TGnjod5Uhw3C37Cns3cnm4vug0mVIcMOgjWFdTNjW
rG8pBOEaV35XlSMYfAwkeQGuf9dcUx6hTHKpqLHWz7vsBClfLE35+sJMjIdM
WbV7O0aaOBjAw1ZAoJ1FxK2sbNWu4JMh3UIncqAhLv3SnNqkmJ2HrpQvxIvP
a3u+jtb9o3nL0cO5xGH4xxlYn3wUcnY78T11O1XmOAdYPfdzb2rY2cmMFhgj
eKDUupnU8Y33xU+h9iSRld31R4sr92cGbeneYGqYOGLEQI+Mh28jCargAG7T
KV1g7z5VOd47oOPejs5xuGBtrWbrnVrL/okW71kkyzn4Qrbqk1pfhR4ZBjV8
ASQAMlWghZMQP3d8tf2M7lDXBfm3YOEKFMNHaqL6panZQTN1CdnzpDok1R9i
iRynbXbqvzYdGrQyfeyWWFT6+EqReMCfi1w0eKRXOHRXDbQIO94ty2UBh6BO
r5534huUGk8HW/z00uBnV6h4QOlcOQIYwM/CdqUS5xF/csmrOZxw+l4jRlEL
n4FzDspzNXYF7tQx67OxMSJoa5fOp2ZvXA2rscycq5Kzd0wxS5g89mxg9Upk
TtczpjCS9w6k/J3LIZkD8y5pg70a+Su0hAvIvPuaamhj8JngOzgwsqDk40EG
xVhiO1WlVuk3lJZWdswae7iT6ljzFWdFSo0CoMPFAQvCF2QloN0ROn0ES3x4
pmbalUbe3LfBqKZ2tTj3fCR0WWPm3KF1Z75bqciuoXdJWHUt6kSgtdwWHGpz
qR1W7tNBlc8xExhZiqeaGqdncoCNDj8iRHzxYwJYt6FaCUQYJ1JRN2iEnSlL
nEEMUTHe+Yp4n32cttZfdQ+qu8cIB1QrMMScJxRJxbdyMwqP8JvSvHu6hWnY
op6wYPw10qMmCHeoYwwCNPRTuW+dMFruO1MxILZwtzNT5PGqEY+0iXyuo8Da
6f091t93Bqe1thRBDpbskF7cvvwx6ZYYUY0A5Ov2vXY4EqopxHHHDdCoy19S
pjy/DRYc5ri7i/VsYDvAqMkQZW+bJm3wah2MuXhWY5kdlDKCMY1usYaYtb2V
FVlo9HGnG8o6aPKtsDJDuf5sdxqrNVEtvkqhzS1x+WQFmHFmBiSUY+bxZh5C
+gqkNI9diZ789iaIJq+zorX5U8Bhrf5RV1DR15h8H1rLift+g/Mcp1IONcpP
cRT16vt3xLAdIPv9NWqMtTcBOJTtTlb0GrEabXHtPWB6tx+krP6woluaGwoQ
w4d+HkZIWjI81gBJn/rq5DNGF4ieQokUJKIuaIxsKmHfzxn5WYMvRcEJ77Id
RmCNZgRmMb5u5/uDaNGk5HAyR/EXqo7pW00FW6uKTpA/6Igvi7uTZ3GFX2Ok
ixdSvspQ2TKDli2bhz/X4oZ9OiyLe1j8e2AkxpWMW+bINUmI+8R5reu/dklC
t7miODDodLtH3LgQyeqOnBJAkwh9DAOa1ZmaMIEkrGE+MJ2fFiTN4hP5Y6wk
tGRnSQDfRfkjHBSkFUnuIumr5TFGfuSuipE7WsFKteg/vZ8wQs5tmU/eCuFR
LeSQZFUdhSmtsS2P7rLfaUmmxHeQvRaguJ9rr0wTKQ+gII/+zPefCMRXZtv4
hGHIbFlJvyBL1zp+mcsIS5fou+81k9K1RplnXu/D4b9SlaMYagTIWLu8DECZ
lN/O7GbvheI4J24oE9EVGmrEX1hj/9PMCY1Njz50wzq8pjJFZ8nTVs5dsagP
Z3pzin9FrlV927nmldYb9aZ3rUkveHfnpDaL/xzCIjAPJv7xb9nNm36vXIbM
a7mivli6R5oTNMoQdWLB1O30RtOv2Nkvq7dnK2qgmUkl6IocDqjLV9LH3rnC
v2bBrUMZB5mA2kK4xW+j5jK9/dVn34VOI336DcamgTJfxQhBDv+GcmCn7jl1
GunU0q5RSgVvSlU5v/2ksMlVaso4FXvQf6uXPEgEUwlA+n8j/BvH6OxJrsYE
jVpGGjbA6gMcHwhq+k4wCyChtVAV3uRzGb+s0laugrsM2p7cuJGTW6/3aTwh
W2zVsN7pAYqfHw8DkDr8ZeMShrNBU3amKP3K9sVlJqkTp4ztFnzLMe79+WLq
EnT4PIUWsmCe7etBmVQ7D5NFpXAMAuSmG7/ub8wPTxjD3ogNy0Zx7eKn5E6P
RCrL2Qovb+/8VC3LqWJ4co9MbV9ec5RC2nj7R4vYGF40OQVC+ePWtBQ/mUNm
TYCK2n0eaw3zwBylmqwmpIyQtxrw1Zg7U52+5WgOqsfSYUgpidbwEXGhVU7f
ABxnd2/TUNgGq8HUDjyHlGRqSYnmY+iIfsyM0+mxqvH/Wk1n29u8ffuM1+AE
YhID216cRTG0ag+EjhsUrTgheaopGrpNSuBvUjSuVbzwcZhxiRGPMYTG4XuB
VjvFwtI62FpgxssC4KhrUUIPIuqorJN69qgfK2ATaq1rG8U9PAuPIwReAyix
dsHusF2WQ9ybdSfI+i8bRvqe1fAuLAV8d8cn4d/ELckNshNnIHTyvofV+WlW
iF2/1UdQv3w/d2RZFqChdBM9lmO9MzYMqVJxOoBYIsTnNd3H2mtDkaFoWsgO
v+djn69eQ7mJITNKlJ78t/oMnlSufmxZ4ivtsZWRzTUm/0ZTXGsRvHiSJUIc
MgrDbMd6w0xBLdm4GFm8MzfgWcLj0y/6o2CoZd3O4ruDiNnoqDQwQkJcPM+g
7gSmptT9PLr1GBY9WY5SY9ZlmXi+2XtyLOK9HRVXeC65ncOtDFGUbVszkDqj
u/FPxITOpvp5/2zW978hkOn9b2lV4zK/U4b1BcTFCC8MiYibI2tkb7CO67yw
bBbXZHSRoAJMUBgjAmSABSuE507Ljyl+jiMwA+wo6pxQf6g5DzMZZWmKZQNY
TojfGYme2WaDQttEFHqeKxkMUsAUPx3t0DF5MIBWLm3ys+iiGXijaDIPZbQ/
vD/YHlvOjs0pho8K2WV+Js4tZxPBsp8LYVJIIMWf5tXMOoMJ+N5U0bzMagXN
jJeXl1ANXJjj9gvW0odbnMF0cWqqksEdRarHWFQviZsV/pE33TLVceWav4z6
tHbc1NbZBq3m+9W4VfMuOJe0cuTHij9HhbqqMYNiKcKUilFOnLFWPV5gH1kZ
zSWMtOtKLYTMjdoUbI5rgTNYzFub/o4/Gpt+5Ne+/itivJEnZWQ0YdRvF5+U
w/ylRfuYpDqfKV4nz0MWhTOG9fjsGXLLdZYL0brzUZwtiT9QQhwQJR4CUmg8
2HKzbt9Pr8yTA+02riNgcxrPDjDxFHpG4iWPz3Wpnd172T33stgTos1hiInZ
OCRUZOOk2ToLq6XA1NTZJy2dvt5eQW9taHhGDT8ZYPiv8k/nTOaI7Iznk9ge
yWbDAeo3i73O6k16VSO15G0fM+v+kmMFBjoRwLYw6GgZ5A61qoIyXwKzx0es
+0hWSU/2UmnYQg3YdSlI2zUDomr46GBhRAPESqzUTA3eaMYFdG4nz6cSA2kd
wWpDGl5jIdjf7yOc5w89JRRrHsujsiO8kAo0MvsCq91NUJzkrg9thu+UVB3t
9PdTwW/fTntb3RgKb1fmRSC66PJmdqZ6pHO31d+8API5MuqtdwC7AdgI+6Ln
/q9rCPhznW2WsMZJ9RR3q90fbUkBn3ZerSygdJlECi0OdSpMcCYgat5vPoKo
tlPp9T8K6AcR7GEFqsw7RjD6oHzBqGlfx6Yjfv4l+4YH4spFb+2uXysVxCTy
J54LovnC1LEmYj88nFQBK5veJSvxj7dUPAKAyezqA5hBKcOgTTeb4lhXsiCU
xBmgannJDlRvkAbJSMe7PHiarnIZOeUmhF7yQYN3gdrzOGbUw5PQ4Xlub/i0
3eenCp9KuWxnfDfOktMAriIcDYMfr9FkqZ5+47IQ8QCbZKi/dAkFFES6Qes9
k/ceF97WUer30zsWWy1bzEYqkcjEmnGFkstqUamME+gjCJuZdF4mfABByUjR
38jbpLzhoVcXHsylyRzj5nz6Y8hsO2cNv/Z56gknGoXYTL3BYrg+UNAeEzpJ
Ei+BpDvwfDU7UySTZoXzUR1cyeSEegfSDLkjesl/lfQbbJmq98LrLKg2tMB6
eyvUai6FXWHRMvoI64jcYfJ1C8VDRbgRXSmHrgMEgjIHJvXO/E8MbM+Y5Y7k
xUC6P3RL1/IGlA9G98JX14dM7MzkYiLF/hwjO5MOCEwVI/a5tMNXaiogUfZO
La0O8TtCnlhIERXQv9zRgXpymA5vHa8R8IZZSuJBmfmnY1YzuhkO2E65bWt/
1C6788ZDSDJwtSAOzJqmM8fYDw4mJup9Xeg4QLWC5fgLuYTiCB5JsACeS4gq
Lfqq3ayFIozCmrNf7riOZCHAZ9GVYmdtlPuv4uiWpKgzf/xt8M5fjsZQtU0Y
XEkVxgTgOVT7i/O4+ys3JuVDqGnkPcqUbRAkASXtSwJbI0BTFU+wqzNsNXkj
5qUQcCPy121k0duXbebOkL2k5ZxKHmK6GNEPMr8sy7bNaxIZ7ccZayL5WI+F
GR/U3C0NGnf0cXPlx/+1/XsBEziO+0qGiVWFSeaLED6nS8UsJe7vgYJ5HCFa
xSHsh8q7AQsAc7lxLBeCWmjWWVLTM6/rlN/JaLNur3AFuzrPpV6Ay//g4TSG
1tSAQWc1Uv2FTHLA67ebqMch7yzedsDvtsKWGL/qmoIl5LAFTkxsIP8imzUD
M8g1qlBVm19CaiXETXAyPhkHz++S9vUd+S+FxuoupE4HhnCPS9hw8DPrEdJ7
0UvACM81b0S5cFIGmpPSq1n/KITpukCc11LdxtqOcsctGsACCvRceE0MySne
BtGFFAYFVjKc1sutLxTMW3oVT/gWgIaBZyZ1YVSWuuohkZMzjTSORJv5FevV
qdhN6lT43xZie6uPLi+VA+UtfvSZEbkqwYfijyyY92Jz+mxbHduOX7cBZmBk
tMozV/wtPv48LTJbYD78X0yzjS5tQkhY5Mi9NQxIKNMo+1ejLrv1JGysY5cB
uAIKCS7n8uN10Ezv/cK1GlfPdql5wpCxmwJOU3hF1IMAaGkIAPViLj703G/l
gKRx0RARYGtvV/YK8AdeNPv3NI8YKrBPIy9e1w872mcC2vgrmES7YhwyHab4
dsHmGbe4aBzfeyT60Gd1Sd7oRjwrkoDn/znGesqpp82Vom/G1ploOBzE7IZ4
31MRBqwvXBUHZaZO/pHb1dTLOP4VlZUww0d7x20X9miQIApVbDIgrBWclg/x
Sf0pziXaP5ejIH5e/fFGF/FCI2PIyJZKxEHD3IrrsnHWCpNsckjxQRJe491R
Gkfiuja+8nGUiubHNUNTQa9/x3Nf3rxYbF7qYdXuTr7VgBUSUYzXv+1A8fU0
CdqI+HZiKq7zA2dmgxbACfU5AuuOEOIEesxxAjAomgK9CB04EOvce2bap3t4
btGt3OC1T/ugtqZzRYKH43kxBsPZJt1h8JJ/NukDMQc051JfFXwatBi4KFE2
3nokl3M7tsWx+C778smrWyJqcMrFUFkvJ4aAP15aI3gk1FpFa+04lsmGfOI2
HdVmi5aolVVGqFC2FSJ2dyqEY2Q6qHo4choKqJsGFfAER9vFQ6vW60p5WoQK
tzAfOujbnxPioU6nitXs5oYFMb+ufwpsSaTUO/3hMbueoRUZkMRnnIqj1uI0
ibZ5jYVr3nHGhZaCmqSLnmLWhCbxpQGXHdpL4vYi1COZwGZf+GknVVPfdYCC
ocb5MFanpfea/v5/H1/RzouQYoi8zDZO+CzWCxJOjsP0QK3zx11VjWWf0OxZ
KLzfc10ldEuSh9lGVwKEpaK7ur4SzzaZpvGW7sXo76bTEIdHrsHJDsv/12I0
0UkdpPWPxd9GUpo9ePwWw/uA1emEltgfyfCWkBPnBEuaw8N42FH5OQkTGbOz
tn4Kb1P9yV28kx7A34ITf95atTQCaI/9FgUlaL8a5+RS+3hPCpVD4Jvc6Htu
AXotbRbpxPHJAKAx8/bA+lWQnJEKj3Lz8TyHufNrQ2YO/Y13Ryh9ngsQ7pZB
p1b1QeCQcsKwsSk1qCmhf012N1lACt51FWkYoMsn7AYin5T61Qw1avF2c9rb
JIr/Cf9CIgVJXbHrN8CbaykK+VvZohtfScK78/5s7+7gMukV6CKzFED7vlWf
oAPmlGrKMRxuI9SWRZbbmY2ycDjecJP23GIwWn+L3DGC5tRgLpWChzyjF6wi
Zm9g+gWHiwZBcvT/knIkRcOn1eImKgePYGm4sI8KCVsjzTRzL2oYW0gw8G9c
j9hI8+Y17AlRUGhaprtAYBE6e2N7/miyrbBddwHjp+nprWsOH64wWSf69XvY
ssm6H1sI7h3vId2q9P2CqhhluXZMGdhvdh2chCb8Wgh4zAKJWPBcn+KlcrLp
Rti/uVWoMmj4XDBCUTULeXeMQpgDBEX0/JH79thjYxEXZE80oEGw3nZLsx2n
UYJeTZq0YsRvLXoBdSkEQ4MesuKUEb1NIEsjU0D8+nGm5jmECCxix947k7m7
5yfndLn64+SE0UU9TRVXf4/PpU0Vx5WRKqK3lpF22VsRSb1Qt2DXvuZ6Ujrj
KPmV/gJtSrrSAU6DXswqZGlq5MoMl9yDCLcNG61syk8G7JtUf2YPV1LxsZ0G
7EktaARr7bLHMsmwNOLfOpz8Gg8RghKsGSrZDPypD7aD67H63PzaTC3L5EuL
xa7tIHbYTcSnZ3mAN7TtNdW/7e6BHW8TDtFkG3ZNrn3oGh1XTtiDosLlh7qy
+upvUkeVbwezYU91eUwsz6OT7J+QzVP+EjOj/Lucaxp0PLwondxKjRpvKFA6
v24AtAfcGslOYPwr96b/GYjcU2k3lX9Ab1mKXTTiAOP+Toou8cZfWSRypspS
1b8ZWxsFQc9CutHA2UmWA0caFYb4OtRWzRm3kRBzDk/ES6yv/U5i61n/D1rw
CeHQczgQPOtDd9oSNkdTuw5L6+4wp9ZRcQPy9UOarvz7pF6ZwXCjrAF8YIh7
NaDSuFiGdEZRJUZtNDgJsZMOkILfhCIlMJk9FFGKKXdp3wHqfWMhz+9qjWtA
scfqTkufdiVKOMq6MJKK66nTUMcTOGstS6rQ1IzLTOx9gyxL+tfQwfQIsHJV
CrhrIRkdSq8++Ws4/FWJtTaYSH4Pp4w27r+QSxrifntGuXaP9YAW/x1NqfKF
+1aUs473i1LUuxedvFoeSa71ZtTeDmwaySX8A7s6d8tDqL6j3g+26rey6qgL
rAxrqV6QKJj3Nzlk/knRydgFXRuJdaKYHgnkk4eQN2Wx1jVNQtbElr5zicoG
d4XPHaNumPXcCupV+s64QdqauXja6T5AczD19yLDat/U6jLn0JWc3gLVQJdi
YJmw6kIkzVVOSBin9ACtx9ECef27gYPCcvOvGWQG9Z59JXlaLgOK43KwfhQf
cZ0Mc5lXDV0gmDSZm4s99CzvEa1EjaLFxc476q8DLAfdyVUHA95KkF95JkeM
dJye1tDFB8FevDjvUGlQSpH6IPJht7WSZFTGmUY/Q7FIU3xeH94b950rApj4
0DHeKyLFPITyquucViMxE3TRrroBi3a57Da0k7pi+RKYfGjSjSaU/ws5VgCS
m3aMKEASBHFtl01sLAme0GJRqozVRr5g8Nk8o4PCPh+4wWsgmEX1Vtxu3RFt
NosxjyoaABautxRF3sjc7YLUBq6PJ5j44DN0f3huwewaOe9tv1TvoecRrww2
IZNLCN6Y/ShRHXLjbhwoWL6Mxc560JGewiAOYrs4Ffc03hfIE30biQnEm78R
wjLeq24ZvFeH0O2bv+8k3feCZpUhEcKcyiC+2YsG7obhti1roYabIiy0JHOo
L0BjdKCTybAopQFyJ3fgorwjsTnLTMfR/I+xUSCZYmtdzKj6gxG9cfBy+VvM
ZbQc8CxULTiOiUp+pUGuL4x20EIfPfrWqLttA6EhzejfFA0vTBM5/tItu1Uj
DiqfhZhXdspW8jSsY9ZYwu0LKKKEdnhCZCI+jq9vKPSAC1Pc7AwTTXXGh+WI
9ZDhd299Fx6L04W7wNde4+uaPGSueTr33jSGE1XKkP+dHFIl7TQoDJu8E//U
ElC+NWL4T4ix91VQOqsxOYCOCRpz5AZjclAqWvq2FHKIdPN/Az43h9dlPoDF
E90dTYnT4Z4FAiD2q1NcfydMVtBYItSqplWTOglMFGgecoo27RkUUR9wjHuK
E6lJ/6NixcXnej8LkBsYJZ9cW0z8nCOVIc3RUYOt2v3O9WYLXIYmETU+dE6k
xTqg7q3Qe97CZqFU6e04BTF/CJQw0sXLlNSVPwxYtGC5l1HY9aExgQnPUA5T
x9G3Nye9CkSHrl9xD3jOXK+XAdoe82ybbc2/gzsxymALAnAEFNfJJSPGsuc4
vQxv7Yi6jrmzShB7TQCGPmrPsFeqk7qG0Ed8OPCi9oneiDG/TtYSWoJWWIzE
BH0X7ODrhncTOKwPjamtvQPaYj+aUd9DKbqgGbipVbY4w6nFuSH9jVk/99e0
MRhouyYkWWNHGorKEbLPdaflqKO5aJH4mDbpjJh1nnlG1RSZpkUgdx/TFCkW
nZYBgdfM1ziP2Gni3s68vL9oMiZhDd7XAv3/g8tONDyRvtZZ11ogvBABtdQt
R6ZFNHQfC8kppRv2QVF6fjkFLzwKQ5OyiVWJwvXDcXpYOyWz7Wa0zt58KouA
jrzAo1KkUK4uvH+iXQwtYelPWnYafkulcnN/Vr+FF+gnyEXgGSTmnb2gRnaK
LKMDHC1Ijqf8tQR7LGAv3nUSEbqpyvijr2jnD8Gt/4adPLIi2bHVNls9F+8f
huOw92PQrTQfLzG5lY9pxeMOExZNkrYcdF5JzIpx/GJvRvvC4HdsQ4GziBCG
Y0BcOCd/NK/K0HDGOUpQy1Y7B+1z4QAWaQoUDeL4XLzfehOYQmmffbNbpIzl
c2lI3JDp97h3+N+e0Eyht02L1X71WZlr4tEIPT2t02BOfYPX1HP2nrl6M9XN
vJfWcN6TPd6Q001VLIHNln1mjlWUi+JeO7iH0yUNsvpxWRa14RUZ7gRxlEBh
r7k5QGzcENiUPNWmuM605TZuuyEp/CzkfKRkiqdtNCrRIqdFR4P1cOp4RuIJ
dCqtTFnqqt3fc1nAnJUQ0itttXivxsUneooB6cg4Kq1HnYKIRmFIijV8YMfu
4aShWV95yMPjcMkMn+4+/CxZe0YVjgBSC2c1vllFlVu20ebvvKWB69zyh5qJ
1uwxENm8zKAAbhKeRqtq7vxfNOMRMnMMXA44W1HXL5T9IqNHBFKcKKs+wk/T
b0zh5PVfdusCRWbOFN0D2iC+8GMZp2n0baVBX2j2vTI5vRo1+YnqFKOZWa7d
unF+i6Fg1VMMEdQY5lUT6BpqxXe0jNsuPELohOf/CDkerv9TzzYIoPSU793A
m5zwMILfBncTXdw7d7rOiXVxRoTewysksKQpw4tPx/+SLIpKRZIa3l4Gt/HZ
qtnb+SkG6GCGBc5WGJebd1+w1gK7YL1QR71IJE5FsoimNlRjrKDtC6V+7P9x
DMSHrxh5vY7srFMjsQobtb1oOtW66TeuUNqi6HRokjAMSVh29pHvgHFafN10
5tcf9SWxw3z0SE2bLEC4a4TgHm4J+NakAAXBTPsM6n3wCwKza8js5BErEvnn
Tt7eDA5YBByx8IP1Q9JHT2hmvFIULnrznYvll/zrnhmV5H37LtUcxvzM0xv/
ArkE3u8Le452pDyQOzM20Cy+zj7kksWoL8SAYPj56Vd5eKNjo9jR0mFnE1jy
7sGeiwhBLmtVYTYhEmauk/kjuyZsVCqW6ivs81Y+9jS3pIbZ2cHYD4de+3Af
KIWtdKOGikZLgGXowDTay5khDPkZemNJvAVMcOs65I7pXKGRwQ4KkPcaUKtT
yRex+FgxwCLcOqDAk5D2fc25QnNJrEvxA+maFaWzwtuKztnZ8OGGVtOq+UNl
9ziGsGbY9hRG7TBncqHKzrWRzq8gqvPgV8WFCqhRpJmYffz37unapSR7zKuo
3Blq9rkijeZ8n3W4pfrdtUTAi6gqDyHFXT/aJQV36l5o2azSU/ESnYOJcPHh
8uIFOmUkl+ddJ8lhCvxC+Eu4zIE4UaXycimYysKT9W/6MWDAde861pWeB4tg
sl/q6/G5p1R1e+cE+af05TYjJkrhJu9Ti5UucatBSdPSdUZI7IAc5ZMJW6vl
duxKPnfhQmMK62MQAFXutCaY17f2c3PUhHWRa9/VvZ4UimGyytnztFcq1drm
mShsLolm/2G3k/+nBS02W6COJsqTK3bsuOC0zAT7N+9uCglhXm3yxOLDH6iy
AzY2uGJmxPRaonw9hvrycGkJtHj7FnXwJO5z9e7lbtckt1uEvqy/ZM4fLQGv
re5tNgc8Dk8/eYMgjHYJMqXeJIqa6VXmmVVF3KGeSzAtIduPUbWOzXIl2B1k
nddRnAXlG9gURPgHHvWafKoWMpT0POXF28vXfj0o097ICecMITuoPACe9I6e
N7HU7TUzrw3ciKo/mKr3U2Whw+KswMiugBQasyuXoywkbIyYWzwXT6hBr7UV
pJathNYLQjoab9VVo+rS6188ox/D989V+73tDGJRCXfWVSF/5imtyjgMfEzi
bg1aWp7gQ9cfjIwbjeHeA6Pg1u2nlT1WiljR2cmffw98snjtWPho1GwjArLH
hoVT58iHfpQf0NBWpLvJ61i72cJ/ip6AZzEP6kMLBtrCrQhLy19xqwgxW3eN
z3b6S2hDH11+pwFe2+lqqzAlTqlpcIE2/54LE/N+hjzTrNyIRIsH5I7m3nwN
ZeJKIvrrA/Df3g/+LrlZxqPkot2L1EsV0N/gTH/dCo/SNugqEgfEUGjXnIAS
B4wl1cRaOonsxBq0wiD1F8+wRO7fi92cMzB3fuTrQgJE0I/5zU18B0QcfFqJ
mddGxHLxCB5PNopadNUksl+/JWZ1hI1OVFZXt0EGOKY6BoisRPuWexdsTJtO
Up0BCKSZZzPK6eAMs04J6ljNtOAR1fVFtZJXbv+GzXDaMRskr7Uee8Dl5UJh
+pUsVSbvmgRA67r1o0/xCYt2sfGDMq3yPf8kFnfAXwjF/vBX8zp/nPvCZ5cs
UVx3Ke3CrsQzCZQLLkNmYHvIM4a1JQAc5dGZ8hWRuGyTg1rXHYxSdvzIaVR/
TBep99yJfkopRzNCg/HIobv/NGILQ1Wo1VOye7jftufM/2AM3lPgkWPWt6UR
RLU1MPcqziVPtpQQEOSbScEHD0RP7GP2cyF6IuWFILO+VRa3KyLBBNABspSI
sSqE55qEyOBbP7ct1Rylim87PRMZIFIIgRgpBMjdScsVHdS6tPUMULAFmv8m
5C8m/wh6S32niROnl+6pjoSXvqnWt9fWLc3SfONH+RtmpB+VfSrfZ2xX+0y+
MPYLfkvHbv7YH7bKStD1UGOIwvBOy+dGOaYDP1aRx4qqBEC1Y6pzMw1iCcfy
CVOWCT7VfTVdzT8AIzfcIM8UPBOqOvgwU99k1ptmjlN52vrBvdjuWvBY7/M/
o2A9o8aLKxT2y826JfkgH2MRQNnSQR4zvFZ4PCjDiHKScOWXwB7Dl/8DGlZk
9KIIfoH0InISE56l3DUfivwVV7WcP824PnsGeMkgVGqdhRp7R1k6BHS9Wzi+
NjAxG+Qvi3JE+S8rWca4Bs5txzNWrQU+ddVHdVsJPDcBNL5uyHkFAiBYAUCw
WGZsM7cAZJgJ9SqHhvnSvcMCDN97fSfcpp6/NhFOU73FlalNb7QMYeOh0NbI
f0ui0HivSDM9raP24l1usPR+Mo7cAEC0cl9nNB2DZhTnBNi9HFEAwVSUqeP5
8lAZGXaR7oQ12iSyeU/IY+wntaMvE59lnfbmIaTzISGWB0Loqm588hL0kqmD
WSN7tSaTwH2sHz3Xiq20+UJ20VkcEYZGAM4Td412kL//6tYQc+JVDDqUT7vO
Z7M063IVwSWbFmtmzaJSUbfK/HRlq/kGoEnnELOIF7J8ozl8cA9JBTuRh8+H
gen4GC+cbRKUbfKB7rqBSXIh8UWLZQ7geAV0cJtLaT/RPnFzUuB3iKUT0Mqp
OygMZxsWYD/jAa3Xv8eDqqp1UxvsorhZ0t4ZKj/apa6dh785FHoQSy0e2gij
UcBF71A1x+7TdPI/7mb8448OluH7/e01N6eYkJOoMeRQBREYI5QpyiG5h5JW
T8UHRdbRONADgsoWXL7/1j2OtXKmZsMAUHVd9dqnL3fCr3iQcK1lw3ELG0HL
t0B1/WxKFbC6MpRDqzQKpsCQwdOIaN/JeCQQl7ofouWSLc15qRgrhtFKw9RX
JRrEFyzxWVpIFClgsSEvMC9YGCbpaL5Oti/xKcRix6cnk5bVCZdqEo7yM0An
mvma04cum09E9F/74bbHoIsendFTm20xMtZ/RtYTHyAeJXXboCziNys4hgqF
4ZueTDWrmwqImdvpcQcIsn1E76AlUsrpU/CJvGbvF8mTt8DpLLO1hweKMoCj
tL1RlXvZNE1DHihFdMd1er7Ah0LTiQqF1lhvyg/XfyCzwu18/fGm0CAHf0Pg
ZVXFqDRD5cRQsgh8+EnrHNiyfc/OYv6FkcBHOylBVjCFmbl5QCh0HlHJWC+J
JNORGSwxbU0rGH0Ghf2iFSWCht6Bte2gij4ysuhBrznuSKNxZCjWIiSDIQy7
kmrxEc6paePweqBUt0/2vrA0L356s1Nacev2fdG95rGlZrcLHti4hH+EeQot
pon/btban1hc3KfqVjma0BzvuL+1wlo0Ox5KvYnrM55zaxc1pem/tJ/OdOUO
UYYlTnmKfgXqLsKdzzaWq1YWYMkWZix1sCMwmgOd8s8SE55EDlit4EbJl9Gv
fjSoN4Ti6cRbEaHXYnzPdm9qRpb8M5ia5XhiaVLN3AkRxSQm8ffTUlAu18mR
yPOwJjZKdRyYWLn8m+bn0yZoZnyBDlWCzinAr1PmQjdEsmFkFzL19spR09Tk
VhvaZPuW8p+xL2+NFaExLei0IAAO3qc5eKBY/7Y4hWh0urdBLJg0iog/JD6R
C0iT7xOh6ReVXxjkL7BYFhvbI6bpMTLhmCxJC3xPi3Ailp0iRiXfBgrWmGFs
LLd5GgcywtoiRbO5w4R66mWG56EDGI7ekCafiIfXO/kqeAYJj24MO5OAhVE0
1RKIJn9NoJmmcvxth4UiDZkOHwsffvHHkvVrfXnt+Ss2ee4rO2ykNzqWoBPF
Vc4x2nF/aHOgUpduJyUPWq53zYQVmHaBvnY38MncEExcjwkadJNzDahsUdJL
VeOSR2e6sfwvTaOuTZha2+HHW2PEH/T4VydE2I1dO22x1Jp/ImAfaUxIXGpP
+bHDqeX9yuc/2ZPbur2cNwNVoVHTrk75aO7s953End9mnI82jneJrTGmmUZE
zyqeXZmi/KAJYUcaDNVWMNHGGI+PYn3AXzJ8OtmKbsQ8IqGLohvAHitt272m
5BFRNs+SDbrwxHs3F+9VEofk8UX296uZ/PeENKYq1+Y2yXgg4x+PTylwBfLF
CI2pJZkKrF3UgqQWZIAjrj+nVtZhHdnB3DXqRAVWxOMk+SvF0xoRZgdexp9H
E9dCchLY1TSY6+eqhBMSSeGKXjPt9y+HNJP0R6qa/MmpplJrwvQVkl/7UXds
HDje5Jr4ciPk7xjFAD1ssuu2dRAGtH5/XmHVIEgLKp1C9gt9qd1fd5wPs4F/
JytYiO7aTSP8JrPRANmwtIYmyGLJbWeNs9deu9VM/1NLRCAMLWkqKDMKu43O
NaO/iqQNl9I0WKvNjNkiKtE899I/q54KjirPxbuOuN5BiAOxB7QHAtAM5QIk
D+FjQ5gQsZAZKg3IEtGFdT1ECg64RvXNcnX/KaatziB7FTZS3ix2omTqqoNG
DhQQxKvSypFRoknZDLzzn/b+edNGfwkfUmrkFmhEVTiYibL8v41hY36Z7OYV
QezRwSf7YsEyP1UXcf5YgR0NNq5M4XRht68iv1UHqMZEkoj/yH/eEKk1TD2T
bolu9HKB7ZUussPZTdI3lBGIi8eCkpsD9FbI+Y488NgU0hnw4ntAxFE0pxMV
3rcwCpfuoTo0Ukos3B08oeIz7tV7d8bbll/Xsc4pBgLnDnLntzl+SgbZHYNy
ZZ71gYhY6L6KkIsdgBISJlITIzlWFK7RTG6OX+tuf0s8qNBbGnbdMVW127yZ
Wa0c8QHqNQFO/hH7PuuEc1KTTo45ScOewucbVLBs7qqq6uVausgo+1JKOUmY
AN0gAhkK0luD67s/Y12mWSEIXlzL8abBCkeABicnImuSFsqt2GK8fV29QSvN
LwZ7rwsR0hVuvPv1pEdazp3BoxpPw5rS7+NEBWkbs8vy8PmtHWZwXPw7SOLU
EcOh+abuG0EuDdapFIaQoy7N9ti+M6dZBpRwWA9SslcaUgdHhhOLm1KsXbCG
/Z0LVLGxK6dYXCnwKG+o+8dwCaxks5viVeF0MJ8Ey2akYsvo20fRiGM5D19Q
cBNqrCB7uE26Lk/jdSv3huf8yiapCNIzesBQaxF0pMaFEJ33gAfXNXcNr6q4
RWCG7ySpeFRc/IBvSxuDmEJrVP5wZVofDQjv/YrXWwFPhmLOxSy/vg16bMxn
TwQ5QiZgvrXs9AyqwPNkoKnr95EzDPSCOyU0Mu+ubpB1V4rb9fxsTawahaM5
X+6f3NG8auRkjtrdKa7XKGKR8WwX+MoPVV83j4KndjauFMs+EnwFqflHvg/B
hi4SjpB6L035bxVygomdHc/uMh/ltC+0XLbDKYJemyi3XU/rJYt8aMqRwgWL
+20oX7xfKNI9xhWlu9btre2/dRIKPTHiVk3hdX4De4/fqt5L1tyapeGSKcXe
hYvavE/LX151Jv6cuC8x99hA9tvHPGToc4/30jw3hGhlB1WNarA5OWtbXwtz
vzal2s1TYKJQg4qLlmOU1h1Y60q0V9q6dOnvxyX0qxxIlkhgNqYSKFlYKA8J
BXtyrGPa+BXGDX2niIV9jhEzuHG0/OHMr+u3hU8d2dDuKXqqObB7NmzEsidH
pBeXrrn6z4Tuv3neY0NIjni5SqFzHIXsSrPTYGi73B9KGDC0kxX1GOXlrBdF
9kl5BtNMCvA1MOOCYcsmKHJ++kaelOrmBmfax+d4opRTerfmLV3O/9KpuB5j
OmLcvmLvVU7kqXDCHPSSmClb/lL0rO1Mu0jEXCui1rz2VYxZIBPAIB0WHV6p
9NWUuefZo0j/nFEYAqFzHbCGVZ+MCX2iJQ8ZOdEBNmcAGupgnXWXgymcqW3i
UC69Iw8znaWxvEgUzDH2qZvhuI4SoH6uIeoK0ZNuZ+ZwQZI/jGq+xFXLkudG
05zG6BdLn8kLnLUBWr9cDif8/NLCJaymtYBILz5wHgSKjKl1GDf7AC3JSWjx
P/pBFD66jIlJHA95ylwnlXv3xUA3nSn5ugl9cnS9KuZXSgmJMZZ5ImLUgDS6
QEGqQK+fxnX1sdrKwCOg97uU9ngBx8laGr1jBoFjYldMBocvVNnecvKtGVrz
OYZSblfmNehNUyvBZ+xut21hYLOCHm1ZlCmKJFoY/to7Va1BaOJxenyVH912
1ENr4WB2TEeyCvgG6yhSjJPBjs5HYuKaZWPGzTlYyiCVPvULvjNE2XWQ4kD1
50gSqeJfjJcSryhHnUU3prcUdF5p3yymOaKaTGiOPf32EMfAyZkK89wTow1s
DHVQPRNPf9CEMY4DOS4d9Qe1PJisUblsgv7Sx3awK1trYyULSjgD9AMzifBN
swza/t2eCxYUiCkOFOZsRf80KnCC6XmzlZk+CtWvKuhLJJ04zf5eayqapbhC
wcjsbLEGx8qe8NNwS4/Rq8D4cFZdpFdvKPSO7xXu0xqWteZwAK9rrg/cqJJy
s0zYAZgTD0OOGz8e2kL1Y+USnkr4pGEGahY0FwqAlEzjens1WJd63gEebVvO
lKP9iCLexWx3SU4quSdfyPcI3ZIdxvKQKnku3SNosNXuukIBx0cDMFX5wFdv
TKGu03FQkyDcYOhi7iPeyx3TK+KBWwrtMQogKauswVT1kFIIiDmyGDOjuOPg
KdkMRYze4T5BKasN6xx4kq7JBIDHF90N039AvmtL8A/+5dk0LEswrVFY8QgP
odKicET7SmHD/WXSEyuDsCEJkgUnVWJYtxRTa2KnNBfI/JPtPnrXVH43rzZk
v2OfgFBNkPzitBsANSMQxsSUXE0ZUWfpnVeAzCIqipcDIZUQ2h18zhDfi8nV
OZSAqQOq64lKO0MTGnYmEQ1etq3xfDvGUEWJRUFBnO8X89crfPCIav9nLRvX
+GReK1/Fauc1Cm/ZmRegBnM3u4gEclWCj8U4gsgzWulxAZsMYKQMdFKO/2QN
NZXqR+QQvreBYeYF0Ph+bzU8VUs45qsaTGMCSStxLC5ANQWhRmd6m6uRxCCf
p9QWQuMamclYz5zL3O8TdaFrqlw2uVWHCt0gPRSKk4MARSbUPZVIF71DzSHZ
CW/U6AugptAMky0RGP+SR1Iy7FjYCissZ4zCoLxA1oCY54sSaHvH/BKKcIFl
F5han/tFPdOQ+9plz5D62wGyp/RCfwE2qL91mkMyOinLN68lqJQfqZ1gwfBb
lFrFX17aDRQxYTUl+5nI4h8QVgMZMLlu+eyUUEGmyNBCC5llkByaHpXQWR9v
uGEESjwveq1mnArCxxePLaDPdXcHqIeMAnVdDSSqUGXUL3fMzn1ik0rzn1qm
BDdWGXOCU6M7YTZzyoP6yV5Q4c3RgVkp315NZ/Emc7liSO90tRXwnRYEmufI
rjVsOrLHPpJDpMIRYC/R1zaHx+cU9DJ47F7okmLZR5By+NOnA00RuDpBDcN5
t+frz2u6vTLcX6K81aoBgS2OmeR5eyGL0NB4rByc8mfhiv0oHIGjQpbvI+Yt
IPA/eD7Wjm3PH5r8bc0F1CUqTUESQN3xqh/XrlGEfNYN6AJ4OqkSt54oTfe/
CYwDsbTloMLlsG7cf6KtshyAyxzUXpiCKhGGT5wvk8uVQl5tNOFfTT/N3qNo
VHUaJv8M1kax3ZSVaA5NG5Lrdf9NeuTfcdicQ2mGJT8ShCW3j5BdhPPVUJmb
mRjNQXWTP1uhHyst92oWWxlSyUese961WtREuQHh9OsBN6yPKSWFqTy/1c/d
kDpnZ+m40fZ+aKWqUCPnB260qBEXNembDkrtpy44blbVBwZIfoFJyCHF8dNG
RwZIkv5aesHekP3/dgnZtc5r9DizfgMlUYJqk0z2CX5A0oCV5ENMlK8XzXWs
klXCNs/rmjUyuOVZcxCLQZggYy1oWBHheVm0KNuy+gGaOiSCXgU4SSuBTgzO
vU2nicekVQFjZcFYxa+fnQB9dzVDx0PMPWc/rhV/21l5WXkPq5cHw0pk8GdH
cjxR/4tYzDjhkg2aISf+h7eXwP/epobL7V+pimxdukp1BWuXsj05y0Mf1djq
9CIywrV4XcvMNVw2nqnzKU/Fw0/l4LhHOCCGKFSrjfbKIWDdH4dmya/vo/Tj
uiltuaZLkQvi8pC9doTT5zYSfIdQIKXxT8SSg+ViiswnAc+IpSfllUfDpIF4
8qFDUaHboBYvtRT2+JX6iNcNO/otCF5A/jTV9ZV5K7h4vNiQhOYo+SCjlyNY
sHY156i7zrqZxZuGRCJqZ5EPxmp/5yXNeUD34dUZdHr4CQWYT2yWqdPMLM07
W7m1bYTrRZhbIsGrTjAJfxM8cC2pHldEEpis7f23k5bNb/HQh59ptpFngNfz
LeVr8BEYhTftLD3JDNKHaZSNkzBQrJ5k9GLwbJXNJ8HBpfcLH1SxNXQf2nkX
RsTP5U9Og8MxslIhCzMUsbvGowFdmE6GD3e0V5/XrbbnAJJja/IdxaFvzHhm
IZrAGkB36i/emm2+saRJBf09n7Lu6QDqXzVYsMSYERPmoso4aT6SLjeOrGDP
5Xsa6Ehznr3lCkTN4VV1wkXUsucGv8D9mlk9nlnbajeJcJ5rELPqzjI++OEj
UFOHaCPt9UwkPS9EscFPhAXjGdjDrUO2pXIJW1V16Ro8Qca4AfEtY+JBNqEf
EitCelhxfzTQDYR7uObncT4389zN2thdW1O1b031j2htB2kluAsujtvY5O/k
ufd8uhogO5UhOaZ0qjfFH1t8yfLAxtweQHJeNuhoNemJl2t/D5rxI7jnsgoG
6Yh7KzQegRt/flQkDOmRmN+MYMJ19xhtkDc5JdDZkGTM9FAKNDL6HPGMXsed
KqPXugPa+XoR/nlVu2xK/vUViPPARQuzzsrMYInsdyGPB9ym7c9UmnSCV+2n
9IOi6YwddbteBUlVBeNyO4hy0qn8QUBcdwtjNPJN/L+DfCiEPDT/HRZDgYOK
RavPdA8/Yxv2IuCL+Wh/Tr6ySEn3Hr1I4RZKrM1mP1WaH1WVRrlqyqfH15FB
8BLNelxlxCkm4mJhR2WeedDnHUxeR2LPzBDm4EcqUhUQrMjYBZuD/TbqI7tP
Afgc8yMj3FsXb6eO15IZ5Ah9dTBCBaf9AmexLkM1zQekQZ0AP/8+sTl0g7ed
/W9GjIWwiNe4O+k3Em4/Nubsg7XX335kxjF/3yXKG+3n7z1S98dEN7wT1QFx
do3c2ublhoQ2z5l32fKfp3BQ5fFwB94emXDoIFcoSai2kdr54rz9cpkVldU9
tfUYUwY/R3zr8oKQeo3AXdKWgj2YT9gRNPPk9Y7T2zyGVE6RSiRFESs6ZJO9
OMmzREyRjFPFVhuJjvxn0BmpArs3W/7+M8zhiEwS7kKzTpGZzHoHcU2OuPwY
X/fyCYldlA/JpJMXo+Kjl8YyGfCPJEKPgpKRUSPCLerjbWE9qaqwHWhfobsF
YVe/GavGFzzkSoRHhhxIaCiZjzzr0XRlnhTgBCMbDpwI7mZMEFJeKiL+aJ9h
UI6ljH28AiAecmEU31/Ed1FRJooCgMiaECNrKMZ6n8BueitWdWqenFVyRIUu
SgLjJ47dSMr39iRkxGF6JFoX2Q8U9Gp+sOlEXMYX2Pnj7O9Nse92JV7YzxVJ
Oujx8uL4Gb9JHprhbQVvRyZGZHmXu5Pbb2Mch60j/e4c63/GjCTqIvkQbamm
VKI2av2Clh2ueBqTmxtNUzmO12sZ9Q+ylrN4+t9DtOP9jALS+kEsktXjgBEv
yc058FXr0p2bOEokqungEIGRJ3R4lgk+GGyH+VTA5BklGpu4a+x+d2FnUh3R
ZGwratciFu2PUr+YzM2cLhuS3uPUFGdJwhi5JBAekLBOg02Rlxfk+YcBMqrt
lyDQZoirwtGij19YAl+UquhBR1fRgsRdo31c7SyNa/9zzeIlVjCbI3bMn4N1
LJETxuj3gE3DiVSSeD3bP+3QMLF0nXrKHTCKrq0KNxHw/4BMZRP+6w39w7yg
Ij1UjlC0N4PCKcdmmxcjgx/3N2ujY0jW4Z02N/ZE7UnaR/kUhCYvUDDMw2K6
aLgc9oXAyPCAxwhGih9hfpARP1hMMUS44MNNaAaweOvwF3WWzQvAsAp99/a+
vww/4xt0IOkaw2n7cU/1DzVSsJ/XOHRkVGDIhC1VgOl503Yz073KCgBsyt2P
9eXgE0OY3Ve7Ty0rlKBlrMR12mSw+ziAUSuDuOqo3Cox/OHUaPKfjbkkuHsM
C7RcM2EvS1Kz9/X9X+Skysz9sR1cFQYJVTX0PlOB4aNCc5ukaakQzH21J9+x
EE935PnOxFdVcomzFWcmQ2laExIvx2LeZ9+WjGNrOMxqgT8NvO8cCDqF0VrN
En1b2n+AM2Qx6zJybtiD1uI8k8qf1gtGNYzs/Qs6Mf0ELDqWPBs8Szte+xr5
kJQ8XxVjU38y9MCtJyv+mOzKXHqmMicTVQ7EaeQ7ZfuzWNwNlsh2Q90dNPtE
HV9nIg2miwAiaX0YNnnJ+chDEIjDsepfipDqzC/dqK1zqG7px00KUzZz2obU
dxKt8B3rU9MzsXTJFyGbmMb+mQXmKSQkz7TfUo8IHlvn7P4sn3YEFae0MANZ
mk9fxvy73OHytNPHEDM7jfwY4G1BCP+Fqt1VpkB3B1HvtL6QvZAqpDb7Z+kA
Y6nwgOL+azBoQvvCslbFLt0zXMap0pXqcqmMinwP65huJs2UdUDV3uj/+11y
LLCivIJNKicyhLYG0H1YNF0Pv9v3aKwoUT6rSEBfhEaSQjyFleKJhrVI1OnE
KaVnvfCMtkWjtnWcneRQwRaDFqsTBG/Xm59md1g5hVr0W0tJnY59XSDZh3Py
PAVYZVK59y468ddu0EuBGxmJfPRfutmyJUFBdaO6i1qco7z0bXerF9pA8bf4
L57jdEQ0JZ0dNJSzSyinl+oxMgNXSaq7aiuFLi/k6+kUniDTfHLnfn1n7+s9
pUDl1v3s/xnE+8I0TPMW/7MfdX5RzHx9pAnLWbYCxhU7ePfcCIrhGvTLqVPU
kgE5Nq6EoOp9lofPOKP71QGnssoQhpdevoARmimrGLYwBG7vUSQ0r7aLaXx1
H9LD9V+uO0O7UIP7BzfC4ApBogr3ChApI4HxkjsvbjiUZEox9jZtelBd0VCm
LNZPT/h3HEo6hp8x4l+Xn444izraLVtq1oESturOxSoffn8OwCsrxg3vpfjO
aa22DIBxIUuojxoGAXypfZmZZvVg6OeHS7W0C0KkeFt0tYZ3uiPwEt0J71be
xsfy6Mewd8q3I0ykPDSxBO4cAhM1exnZey70sqsZ/loh/Cx37t4B6AM0tMIo
rz6dU8IBNBgYFj7fLud0RKCee+dBMJnt5/rr4zOIUz/Kf89oGQlxwDKuWwld
OAO8vJym0Covkbn5iIEEtU+CJGC/8QwzPIyT2Ribwd6a1a7AlX/qrnV8WmZe
37EoMdPqM62RwCu4QUlwq8SurR6g75ORurLS2eug4SllA10pd3fo7+y0XPL9
VJZKKwMKXYxyDDbReX+blqaGc8k4X8sovhCXHEd+TU9sY+WU/dHPQOK5MpsM
z40CC2C/D9cy/zKL5No5/0uvmgJJw3qSEZ/q9VkuJcWRl59+AYff5zcGCYvF
OsELfAMOXiN+lvZc+/iX7574TEYlUbW6/oaKpoMERSQSyKZ73pOm+mBIpAIG
Xu3T69qYn/P4dDEbduOyNMYmE4joEfqdUP+E5TSQUf6we9FQqJCGSz4VU4kE
4c3wKJFn/6BfcSckd4Kcoyemis3li+G1RssfEuSZE0xdmlPy67fiQUM+rI/W
PeWGJv4xHhPnEYQy/6tRqIYjpab7t1aFW8izdCXhprpEz2ZdreFXhkK7tVro
uOgQ0tdanMN4U1HSwfbaRJJQIZ6UghbvtJZ6cr2H6M+xzd1mWbBzn5lNSDhx
9TG4v1Ep8q99g3nVPWs5ItF6Y7/uBzGVrHBNUopB5qDNjLIp3fc28f3H0/uZ
A9tZCHnMUWdMd31Fo0lDhPMmvttAS/+Vr+FBiRq9E1EENaf3Smf0V0uzR95l
mFsbMa91TWiKYAlPm65qcdCrQemKlLECR5i+3UcNpv5ipHQBsiu21mx7ajKa
t44ETMtsioijGIw5aw02vxZiAiCe26uyxYzNAevLkk05EtGKvW5PnGg0LerZ
ZBNyHDNcu6B4rj7kIX6O4HNIEWHDRKbsRd85ZIdSNJCV1TD+fulwdtU7KfrB
Qe4iyM8O+k1PTXfXuoowN76Vikcvn533UWv5NDe/p/Eg+ZZHsFwmPUA+HKMx
DrfO10uKhDDhjfAwfVE0ib9ykHTwtNVQ8qmz7S76qOIonWpWq2d4N8us8drz
DcSr/DhOxd9ow3y9gcm4Obx2SYCRwIB0gZG7nv4QXs/BpqdNndEmL+mImqZa
lIGJYQK7EqLbQg+p46wc+D6cy9y1m/Q55HWCdm55zf0T2qaTyZ+QZ5gjdg7j
wcEipOqkUAcLYJKPBP0Bm08qKoSuEipgDCRfbf+mxhwbWBfg6IHSGgawfb/d
idehD6NIpeZvTv5l9kK1YeFcYf/pzJAAXSCI9cr81r5Dg/hovmX8FBqqcHF9
hOoxpa8qQcVdxg9p2PB1GCuHC4i7luJ3ImNsRVhoj8c65x0eFPWcbiqUz3JL
lWddfO33kYQ0TrH1gmcP7uMl2Zg2i0rA4D0jjWXsFntRltTJUKH0lkH6GqTu
ivEEg2s5GvQyb6zzMcmJglP/qPcQG+7gOuLT6wU+f+J3Y54MQZGDIWTHk46G
f3cuPp3yjkofdFJSDUWWB5WYRRWpWsMBnsJZhgjh1X7VGFeol1pSJQ+ItaDo
/Zac3AfUHbgGXRW+RX0WulRuVFlAwJbyKWTYB3r6VyjpY8h9P9PWRaYG7bMF
+Zz3ZwnHn9u0VcGDAxs8JnDbngdxivzXKOyCmoo13IDOpJnltcFslM/W7T0M
ajTXPfmGmgihlNp4Ou7f2I0U3Oq/snDjJT2fubM8DjqSmw5C0ntjnRL677qT
8UmkRK60W9Ahoad4neLK1bWshPTmDpM1EWqj983Ancm7DSiLQvijYAK2eDfK
YgafAlCaLSUgzc1BpX1VxUC0N3C3pQFNwBcd6YWJgwzHP9Q3r8BhVkcV1p94
T8PFMynYABT7mQY4Cy8DPHUv0HbVeRUE5gplbndXEHteV4Kv9olm0d696kVL
iEWRhqGS9jhTQsM31nBGRmnprhF7uR+jY4LYy+7/khSKQCCAJYiwkcVEf/Sw
tqGs67VEWjSd8HE1+EsFvmnwmtG9wWj4wEAzW1gjMtvrOgi1ZXog9oqBZLde
7ynKaoONo+aaccdCYBaL2rtIER+wXF6A+jYxSTcP8v2Qw2bXcUlZgbP24hyz
r6uiyfObgUIYWfCimiE1o3xEdMjTZJ4KtSqr/jel/DyIKL+lXHsLkzndbl7o
dnpNgwZglUDP2EdxZhUBZonlOP3poyh1/u+qUTglEXGGXprXf5OCA45ze7Hf
77BOCewUokkIp7XRG63QBu9LSP9I0Eltf0lzglrq4MhdG2H+tJEpZvklfK4y
KP8OJ3JbNv9G7gpAHcyGZ/DSK1GaDbZimLAysdrfRlznFOKT5pqMhATNfcRo
wW2ebAb2LMrb+PInvuwXeDKeIISjbPgH89u3+hZtWP26BCauzmbvo3aY27H7
AWVailXioznoXO2m+0fDH7WrQzjqsNx0tMIb9dYGEE0EEEToTLu80TiLPJ4t
sAOzONdFxz5U9/pK1oQJuZtUSdLJAYlPVJ4G8udlbu/iulG10Uw0h+Kyzheo
dd3sfrY07JX/Ko2/2VEYKAQ2wv07E7NAORSsuYJaL4j0tujPixzt++/1Hbnq
zpa5e4AlcdfKljAesjtwYbjFwafBi/qycA3meNx6aqfQQWTsJUmpy5KLrX/h
6urffoCemFpwzFQrCmgVWe4OXw7SwTr71sQvQXLGrkVqckd0qtDeQfbw+iGx
uXwmUXQApMC1Ruh5NcLpwwqSos5LfepMxFgNhXi6wleY3iB5ONm2gfza2y3X
jNpYMpKtxN3bCPT3zIE5OzjuHvQw7Z9fdb03V+MnFgj8ASN0vsdL0tfrUeUq
eESAy049z3rWd7DNzRPGVhTVhbRGsmX8CqN+s9Nbm+zuC8sHxBufSwbUYuK7
En+2Ta+AxwdDatOFfIE7nd1EsolOk7Ouy1IHIjeZrgttXM9j64Ht++wrQyHQ
ctJMcQyWy8XhqOD6c09IQIHkLhYMepZmtJIvIsMz+7j8uctb7jEW4xPDNmU2
ugyBwvmemQLQs1TaoJpYu8AOREyfGtjUZfhNi8d+EGdml+NYkY44qSp4vfQ1
W9BtDntYZM9ZqnNBBImE3EzlvGnVN3LoagE6jIfzzs/3EDMX4B+Tg/LkF7nR
36gTSBHr/Pf3hUcA4uwLtpYwAp8SUKChBH+NflvSReRk6eYb9/lsUDYlriZu
Il60AFJ8TwNPdPp9Mc0fECE3mposHxfB+xlZnEj1vuRJCXlPDsTit9hfprCr
BAyVtiyBHSAkLmvu5PYNPNMT26ub5AM1Bs+U3g/md3rfzitGwt2wZvDm83pE
f3ubK3Rj4TxHc9yJOP3pLAw7H7MJ5DPh1n75Sfln5jYwBk4jPBx9UpxhEWWn
lYJ6Sz4Fb2wFCaKwBEMsff8tJ73Oweb/n4f9fe5re5+8noZ/F+cXo/VcSNg0
0abD7IqYN+LbxsZDIUD1YQcXNPfjAOcu9yCaTqMM1Ee91dUdo53ZkOBMK9kB
p9QWbTBa1ceAbExJF3QQ/T+VdASirds5zzFlG/RtDXcCGsBBMXrmmVnm9w98
h++zKwM7rqp8Ex11ekMg6YMvN2hd9ZsYmbe+2OJ8GwVRnMu/QQB2bSxthxGN
MI6LZ1x8DaAw7Yjk1xYkL0tx2028igjS/Jd6hi0XQZuz5T2vK8CQD3eOk5Ey
GAsq7yS7a94BdEfh01qV9S2hFuqwcF5v9bcYSLAMjgRVNGVU3SjN13NMpwYR
sMF/e/PlcwL7ph3MdS0iwW1B4mv+VAivNLaGgeKFokX18yXsdJ/wKBHOaK1A
2l6hYDlzaO/Pn/poiBgXzQKTd2Y8pKbB9JrSnNctvXI07iVa0HT7cfkTOh8m
hkoFNjI0DtjRYvMlcI1T7m8bOadjvKXqauwbZoYHdkWIaOfyIt0uCcDYbBzd
nFSrGSIN66a8K6oqqy3Cxkzc9aEc8g5MTtcc3W3m5UdUlGrndXMjMeQPjr+K
H2slVeSURbur3tMN4ubncXpc+nho+3Nueae1XsZ+j9R6UKh/efpSvCHVri49
IiZLVOgdcBB/Q+hdVN9OEhfvy2095Jnk5k0Mg6Cx3Co4DSRjLLaomLwz4INS
H1BlmsQTlfE9mRRYzsApHpmgNjjIHJSgcmaRnC7xOh0DI3mnsVRiKCw1jTNr
EProFqD4do0BBU+heADg+dzoqIDvSm2X7jnv4oLhPJ8oYyhZAYFiH1M1SX6G
ytszZEDGU90qiWaZNh8XWtpT9Cl1DvEoaMK4+0X5RpzGIu6ScceqHn+gdOHM
/j2D+8iCyEWpekN047Bfu1vmCN8vb4Tf6xLs4CLKY9dZ/KYOtgerguE5Us6u
b4azMURqLbMo4XhpshF+78L81HqF07jyetbAYVLUIDSWETWYRyDTCv4CnzXs
P/mz8OVYt93/4xr2b/pnkYKw9pDA0P4MWWr+8dE6S4swo2a/xGAPAdadLiL8
VCBWHe+vYLCjCMRHPMmdSB2BIGelk0H9Wr7ZKVHHmWogvVbdg0FTf5Bys9OL
J9CNcnQqOWVPyKqLgf9w329m/71ww3I7JRP7d8tFY4c48RkeWVhhqS8OalfT
4vv4mcTHXGcuSc4TrEOuaUWZv5ocnEGJloRAzBrEujoL0sTt7t3Un3Fn42An
S5g7/W8PBWolQaRaFQWqzq7cwvhzLWUyvq6vuv6iNUQeilwTMe7h8IVmkfAQ
hbMW3Cb7CwSknuJYm57mX1ubRwN2gF+LP/fvazisGA8e88VIUn5bEXFbVYfk
Mb4E62fIDdht+dDYsfEQZEX36p7+GyQYajQ8klyG1UcyZgvX/r5C+Gkx+VKu
4hLQAJJ+IRR98qd4U94X7NdPvQDmXN5Hn9NSqSEGAXWfXItWTujAssbq8I47
EN/vnoTKqJB9EkDAmF8XADSemlOdAr9quzu3jmQfsEGuvJ8SJlS6HBKo983K
CrcSkz+Qmx1dOoOfU4HtsrBGm/9YsE4Bro8k7Dz7F+gO1Ts8lJeuThqAWRiy
PBo/CAWakL+X6dc+5R6i9Q5lHG6h/kQ3SJ9tiqISCkTdbQ16/Iuo/XF93U4k
4FPSX/JWKMLIhPX9+io5/VDVR7TByRjiVY12XsTgYA6jqGMuL+oMxaYg4QBv
+eGC2jb/OO3oIikAixD7UXl2uphqCvB8WsuhOvTg1Y8PB8SP8r95OSEIbBES
DmIx1ZGu4OpjA0yMPkRD8FOWqpIlCWhRG6VyKfpW4RO5Uju9UHnDJEAAk4zM
WShE+aW5RPjZueiKI7gcGM7iKlvhzh4pJQE/iI4yoEmbaKfaoql0Ajw66d10
kN5U4F6i4x+ePaybRaonaMEFpr8YsfgjvnuNN/qZxY848u2Dyk+lT2wgqAea
jtYm7eS0NODTsGy9xwOqsxL0tQNzE1aXj/sSH8nDmKckfhTAIp0QCZMTgdSm
qieDS19qFs3oRYhQeqH9x9oA7gF7Qt/gxz35jht7Bmk7s/Q8Y+DY2Mdn5UlV
db1rM6xVDqIAexKCGeOMjdjkv0L5XW2JfkjZefKNS6CvVj6rJchHrL4kZhfh
FoHb84C+tHHWEDUJX2Kgl2uAc+BJZf/mIhjLgBGOEz4KRRp3KtIFEUMKdkN8
OM05RT9D5RVFgI3k7swdouCgpgcDrl3zpzVJ+o0vpxRBthgx0tqfUXauwH+J
+HK1dOG67eSTyNF3xPf+42s/o8h8E6MmkZqdiagjb1Nt9hiaRNE95vzNagwU
B7vj8q+Rhnrl4449Jj28zVRZChdlRrdt8cfDgP6RVsYiH4VU1vFzUJ/niMH5
82vYrTltV2RDLWoz9kXOxpnyI+q6XEfwtwpGW4od+Ie8HQ+93M9NuVmwhqMf
NYmVbg3Jit5FPhLrYZrAr8iYJ0JFeZDuceRKVMy/5Co+0R09O5a5EiqCsqTp
EHAuo2YZ2dHtmDspybgxAs437VPeSEzr1IK7XG0ju+c5QVS/wadluBCZSH2N
UUxiBcGD6JFVQP1zenBUh+Ut2X1+R4WfbjUCc29NTTYoEoxrT3wAO+fbYJMY
9OKG9Vqalh9B35qd1NG8nQUYy9e8yrQRlILS1kytnNYtm4ga0PHcNxBpR0p/
DFMRBL1BP9nCxcGkp9sUc8XgnB0/rEOcxFJeqianff+rdQItjOJ15/W2qFEG
OYAHrdYXynWW3meU3kUfaBb/4dBxQoEPUERRAkmSTGb0CLXuyFO9Yaj5BitR
8MVTVY0oP3cL5Snz9EKgLY+FIdocccUcYs7G389m/B48AuZ5SDPowoyMFMHN
xAD2IRUYZZFdk0Y71jSzTcEXqMlluTsudIyQl3KnhGlLh8KViY+kS1tW+8kO
s+OgqTnZEIZ4RLJBzU6OBUKT81s57mYpRu/FRRPWiX7ZmiRRG36uRBDQNNIl
DfZBwDJwy3fvHLRxUtN9gTDw+ajlO2V8bEhYuNh1KH1RUABTcEyKpX/WxdVs
Ghsx7QE3D69h8SDKGP5tk+C11KsscYitDzpG9bY077fOKf+5uejgrxJbJYaT
V+og9TXy4p6CZ/GByf2a+ZiINsQ2StXwX09wCTPWrZ+whW5rVtDrwVMM3IMj
nl/DTxAIyd8U99XNkfshKVLoFcoj88RQW8kV+RmUhTnvsddssCvsPqT4Xi7s
DmGdpVR4kYoNY4sm+tAsLG8+/mC8yZGpKU2uZ4dhajPdJyYbRIz382Gz9xLc
i1kxtRh0Z8t0Y9iUM3mGK2IGfLIOhEWkv1VcPm7nDjnd8XmrdSelRxgiVJDS
DNheelsfjlXwKLUZmO/c4UA45NeB0qriDtpDXZOV7tcvOjqS6JDa26PTD8TT
fkk14fC1ch6nqrxRnssMDQwc1hrIg6THfMg6hS7Kb8S/+ggxBe4w2nn/P8Za
2jHezB4JIxKqNr99TDXJY6j0A3dQypO9iMUZwXweJdW69WcYv3kn56ioLZWT
puI1sVjbX767CPVviA0NzU+c2HpwQFhdbSeJKZkncuRMUlZ91wjRcj7uXye2
4EfQTWdHuSzwrmx5dLXeWP3z+EFc5X8A7w4OakXHAM9yip++AJpJxjgA5c2s
B/j8zzKpWoXnOAq88ScL9l9mZkOPCvgwmVe1dx0DzuJr5HnTVGV5XybQIgnT
GwII3OebxiFdiYLuzeO+XG+9itnDt3RQp2/gkZ+IHUcC2raM3BOICnpQxPVv
uL1BTocPEKLMjKoBILcZF28YTcqDN268RXZ3DDTqAPdzrq677YuZmahwhMSv
sPc2mmNDiRsU3lgFNa/QCjnN91mk+ahLbrwYyNdzj2rfwK4zAVbLPsUHA/sB
dMpoUIFgsHApC5qJLW6YmxXUD0AE7upOJHbZCQYGaK+pzWN1hHubkOrAdung
z4h1+WYjrUhFkJXIOlfd11vmT22NX+ZKwekBRVxZ/kxXzF5q5PbZRr+rnkh/
63CimoL6bP0NIaK1Bv8dsFDlTLooe/F0DIXB3nHcLzfpLwoUDXhJggbPHP+g
mpaf+61tXPdaQcqwPT3BHfXfieo9B3p2NcSIqfVoZIcz0UWqiTBXmwBakAPW
tbQGRphvYXNYOcAoNaRAMDPtlK44Y/JN1OnHuK0eDuTumZcCfUnza9Qp5Ser
m56mj4UiohZlef3h7wJY+6qSETcyKUD6QVjVZ0p1q3+sj2VoLmVIpK0jRPR7
D1JHvFrfTL73VyNV+8jgkn3JTt7J9Dh5j2gGeTn4EKO5Q5QwEacfw2rG10wD
YHLOPeQD4/INDUNURb7vc0Xyqnq2mpgbYhiGDBxtVjRXTFeP5CMzfXfc6Npm
dnn74rLG0iWmTuMjW0+kJUMXkz45kyCjSdT3aTZvUSPxgJsdoe5muel9N5Ck
+/kaGvd8W1aL6wEg3vx9BfGv/n1KUbTymA2vgGlIvW1HYxW474gWJH7PSRsL
U2btrNra4F1gmOhL3+XZO8MazLHmKDC4v+LZo0YP8e7NxzY8vGFUWpJY9JFZ
xUMkYjC9EmjJnGcEP1aQG148EUn/k9d5lvFwpAJswGETEMZJtuKC/5E6T5VA
brO4zq/O/s06b/pHZKQzur+sLSukqkpbqUEP1s+dJrhjmW+vOnHP9skJ/Zxw
Z8MtrKRv78mybfA52OfR9nJC/C5JuG9Ef5gIsq9aA3uuvY3TbBXLCiVIgHrE
6j6BG3pKoUGHDwLSLT/LfNbaDrkqLCcno3moixRrJ0CxLA0Ykd0Sv7dctHQR
ey10hCwfHaC6u/tWfrgMuRguGQ+ZEAb/czydv0Ly1gm49U2Sts+bNpBsTpl5
g/NZiAdeuAHU40jAnsawpQG+isi3zBM9fpBFRmIVqh8Ju725vzJCi/epXu7W
U1L6d6jm5Za4ppQ10cv8qcjwlQ3nSrlrk5tByOkoZlYL14ijXOa53H3jxu0t
jBGiSDFnU41Gq4ZSNl2Jm9ez75prCbfZZzNeSW7u2AVCt88Nfh2DF4tNcapm
3kv0hr59ucI6GGEGI0LCECAj5eD5QAAY3uVQIWmMTPZne/1Qa8KqV+svSubB
gTgnaOyoas/TAAak1rjiY3hWvnM3tYvJXUTuYGPbjeMTTIkQQVz73SUAtQp/
3Cv1q+yr8GXQdTnud3FhMoTWgobXlYvQJQsmPr6xRBUbvMf5JFraByFtMBrY
pzqmd4GHsyfXeqFWDnFm+6YJtxbmHDmzg/I/N14vdZdPhG6ldcLFc+rR8hak
uARC8OYYk32qdTG/DqsSgzYwbcQ591deXP/+foB9isPtlU7BGmTZ+WDw76sf
ypD5xV0E+CdlsQVFDYoVBuQrxSCupn2xoF91Jd/RmGcnvdc7J1wrv+rQfX6L
+BWSUgYEh2R2KfuilwfIjq+YtpuUxz8kndAUir/4j/J0kQjkZTC+a9cJDcg6
uaoAHYqIR853wfCRSBetRXBiWso84HmnH7YEY3uea0Xc3wsUrHRPqg3XgHEj
rA35uGABbBxz0yUc1W8bB+sorGJCEYsJcf7YznSuqwkFZs6bbYeSJAO3QFb/
MukkpHuwTNoIfBFb/+7MRh9n2ezXLMG7Me2TQ9q+6aeNQDYBReFaCbBuPwCy
c/e0MVknzoXHTar5JjNmoSIx2gV0nfAz+kH9TLe8+BC2AEIOXPYsqEfy4PfP
yEFxSsyMAfWPQ8bHjHTkAU0sJWhiQ7jBra/fTt481ERrqmpi3+HY9U8SlUqs
FWqboR0Sg1l+0sPJceRQPw7zg2nauqFLw3PpUQBz4Y56i7Esq3/KE38hqrDs
0XvJtx8z+lU8q6ZO1gVpqmHsyyiSk+4pUqjSAi4RIObsJX7vXQZpgfOXWEXx
qHkk53kTH6rBsYjB6VBbypHaRh5cCpg0Gj8MZK8aKQ7MQJRTKtc2+2XARkoZ
6oNT2YksC8LF88Dx2BbwLYzfmGEPl+uUaWYL2DAaPIZ1bbUh65I55sfAc+07
mciRnNsqtGbdC8ep17b5pI/oMmw9XaRzTewMt+/Dgh1Zh6fqjCOAGJaZMmt4
zXoMwYOJ36WC2NLx8mRTUQUsj8I50y82uU0FCIAXAHRF5bm2NzJ23zW3V9UN
4sH1e41vni8gVUg08nlagPO66T/g7MfnwTkM9y4jG2Hu9TJixmqDO3mEtBMT
zNT0Nfk52ubiDISkmDubx8jaCMSzA4ukowLUrSqIUhpVfcBRnweDTZax6b4j
wc4qynxqHceNnyJRQVIkjkhSfbiGwGA+kLHD8P5wyrQNhrOUUXNDNEXheQ/W
jFhxJ7dA8Yhq7QYaAmTmqqOpYlwtbQgOdeOSsW89sGb3E0oX2Gwhr8Ut6Msw
fLCMVGb5X5VCZSGPJ2dtgbIxADL75XVrvveJLmlxJHnJ1+uAO7vQ3j6oYdQd
CLj6mVrbxID7BBxLcNg0rA2vLqkbyOpAzA9WTQpAgt4K+j1BRo2JnGcl6mT2
jY68Ts44ad/dLvFOD5w3HUppB7Xo3taQ1QWXCmSCCE4PYc5k57jh8IA69D6T
640XTizDVLchDOEewVhYLPbtOySj62g02NPqZgyPtJxHxe7jXR15O6DGJ8S3
82wY76Zwx7Fyhi67j8znHR+f8n5lLCo1+EuCK8Ux4Hw8ucVnkkW9YoZv0al/
KyMPI9F+SoxTK6bLoCMwzStqJ+V7MwXBWI6Iaia+7hyhR2jjLeuqmwVjQTF9
hZE88S5xlxWnKoHtTPwaJtzzJWxL8PmKXD2rD1DCKrYAIX97CISv30mM/6p9
0PYETFBIwkXPk70CYJbl26B45j1qTlck+JC+FOzQsHsnBzx4Fr/zACAarfYC
x42b8UjjyZZ+Ry92BP3OrI+R6m8KVtNB2FOWQC+s8G2vcpLMkKhiUclbcWLd
tEN2I3Gxhiwhdrqbm5Hpt2xvBZDyN1aCOHNoxgHsdcl35OoIep5hiNgUoNUX
8nvvobjB0wBbtOfe/UXXaTlvT3QqsaHWQRRK7uSbqAIAK9AB3dhX+vHWJEob
3cmVQ7OabLLkAgIziB9NcQnmGq0QADryyfgWLTQWxThdeczhqJ+xUheFZEed
91YhB8xIIQzEd/HadbU5fys9MdnvKiZMY9gpGchC+4gkYBdr4Eux/r0if1g7
lE1jZB9JJVXWTralgKGTbjInGNy4pEZpltZqU6elVTMOMRre+3LJ5lafglCV
HAABzNAhLS2dCtcnVBGFRbhBeoIZ1dWJnGd/TqeUsBOCJwKLi6KVdtnQNAfQ
GIyAWyHqP37+Rjv+0Gi+v+C6jg9HEawfUZFMa6aszKcAdLwgx+9T4H3ejGW6
wKshqUZnUkFke5uOfjHmGMymNLVuix/n3E9XlANBuOlNPtAAU298vFRtlVoY
0jG+X35mZHu0WD76jemQzok8dvXajf70Ys+MlJ3PaFg45YRgK/trE6/k+m/q
kU2KVaQ+Esar9qQ12OnLyKF5mumf7L3acW+Pxt3FuKSm7p4m1jQ+8t6qzszL
4Hn6F9sk3fw8LBcu1hEJNwWJ7Rzy4XlrlAKyAO8CynnV4QjdUowsTEis0Zt1
9hlqHSUMTtBxeFZxxyap6gj9lAA0CYkHYDuK0Ojvn0SLQkFNEHCPVV6YIPpj
TOG9cGl5TqU7zoxewOwczbbD0v5ADeNWLB4HU/v7W3a2dwOPfcR06RlD4LMw
esWLS7UBQpNgK4hXI9bfzXnNYok6rFQIC0wyVk59E/icJ01Hp8vEh4cJC+ID
ob6CzmMQGVgbjdJMrf5YDaF1Fq9GRxtq7lBuyW4Nf8ViLprmRVVnbpdST4d+
mchbhiUrs7zrk2OSo8E9p8IW/7yMcAv+eTNnrA97WHgdNwJcpKEXxcPbNUlm
41CcOLS+hkrv5rcmYe+vwd3vC+JJNGcxL8haW6tpPdfLRyRi4L0HfIVyb7mo
ydgJj4Jq1yCAN0mi4aeEd5U2IvUIMho+jOws/zZMRM89w2RsW5iU9AXf3Uzi
CazDDAK//0PJM9sqJvhZMV/VUYAMLD/S/kcS3Nv1czj9ONopvl7wibVXDGPB
OypxK1Sh5v83ah/l6KOqyiYLjrRZVNuPdPidBGcdLM4aZViVvqFdJS3dsIcc
3VZe3lhXH/jVcLXcbmamdLaA/t2SXrmppQWwZRsQfZxRDyr8ANdGMsPFOU+7
jerymFTv2Pg/MbFftwJaZVSlq5rpZXMky1+Me8TvUEDwJO4wIODePJuRetiX
2SBmEG0gwmPSptmUbZPCyGDompz56wWPhNoE6dDrAzGF6a2ut6QV0jmomtRn
lHYAntT8jjksXaVFR0ugxL1sPINLz3Ca9KSYwsttNriCBKDmU8+ypWS/tI/O
6KRAaQxXdfQ+IIlcRgxAfJJf/HKuaHwMfCK76R8VmBjITcdX3YjA4SlU/F7E
WaqtHRAagggUt2ISHDO8H/tV5AeiJ2w3geOef077A5qEv0ZmkfXOwfG0hX3I
zPtr3nz7yEVRLmq4JnXsx1v7HylrSeNIkHVHklfHmBz3lmVcxfO+HwTasUBg
29M5EcqJ9iR8a5d7S1KJ1UFwGoDApNCsx3Ufk1SjFyDSLCEdXQJpXg9Zr7ce
2QAxtAKZZ47gAXseJeNhOJhH4cZ53XoQeoEqIlHAMwuAvIeB7NPnAxSDbO/Y
8/b7mpZfp2UYSkO6zjflYfUUtvqyS8OITCn9F/AAv72pNOrYWMZQf6VJzQje
MmzO8shvFEUer3hfaZc+ZSUaq+lpp96LYFr+EsjnTidRDpvw9ewi7O7VuhWt
hzJc0NhqhxzDI0Zm0VhWzY9KXbILKT1AIHCCoJuU44uAlV2ur2PrwXUOIdiH
y6CH1W12gpMoRynHsQU5NbR1VsHH12paZR17D4O/R5gEci6Y/2un8hnw37FD
C2ZTNiridj+W+FlNeQXFEQP01j0N/HbUpUFO7KYKX8wW1Q6MXaDoBOlmNnIY
/qYpASH+h/7E34HlUVk37TPx0mKRTpEMjFhUj8/ISDramlBwKV8AhLT3iQp6
1Z1uEPd+VvNyfgHbnz0YjdtICNHMyLaNCT1/tcUoxcffDqX4TUc4nL0Vap+r
RIpy9Ph4mzVOYDRMH3NMehjO5jtBp3VtBVDzHgRFeZt3gtAxBcTgO5+67Yod
kU6yQ3e3LDuOTJc9LBikmWoe/2rlHU3xnDoHZaCtJObA5iWqxe8WQLZtw78M
jnZ+kjZ0FrmfSEa4LFfKKWAs59u81qkSTqFm8hTgmx/PfVbWzBQjIYvQRhG6
UBwO7klO/d+KTZ3hiq/oNE5W7diWRmoJKM+tSxSdYpIpHvVEeHPC84bnBGFF
2MYfUKxpZKGt0h3iYwvPEPgnX2fawepWN+DV4m/Rq3SKZMhwlbqyKLRTtcsC
ZW+b2rKfHt1N1/tLW3wxvlOLrYCk3hiipYucWSanB0xFU0IGBTsgpbxhXtTC
fDy6n+mrUHkKdKhZlyf1zI0iSZEzeGQiakekbxTdpjQPdORFoL9Ty9TNujuc
kiJe7+rAfIfQ1NRb2od6N+cBxjeu3q9CRH/oUpfKn6wyrCTwrWFzwpu0UQrB
1kxu0zaUrpGCC3OzLRDpun9CZk8OkHZFMiY86Yab8Z4IVNjBfsfBgYShv1/U
RFXgTMVI8K0VB9Y+EGbGGoSnc/4bu7wITTeCvVMG0nfFA+9bFaYPIDySulWG
6JnpyvQ7tpus58qxac2bVUMUrfrSsbfxSkB4jA7R12enGJieSMxZJhWlrJXc
Wvt+ZYzFcA17KzP8Zph0/vssEjp7cnbPOmfmazwkTHHuHVI53hUMoB3tCR1o
mJ4TqBodw1+vqxLGpqETuX0iHw7eq/zKoyIq4+CuPOOIqQLCtuNi6+UvWE5r
1NRyYIycTLHypX9bw98/aeBXGquFgf07QCtXGFfFACHfvvJCWnTX8kwL6UCW
7sNeIRPEra2wim1i7Wc8Jnpal0k3jzRADa8nDgN50O70TRdgC1VJLLrIfReV
x7mK3mYrAK0+T4tBknWuETUlrli/WOlIpqvreiocDlTksaFwXZXK0mwt/iib
QG9FTpVaQGgsovhVObGqpTYXQXOLQqMmjzr4KjzgJhXjVWktDC0rIJXHCJ71
KLSMCS9Jz43ReyzUZQxIJbGsy/1iHQAHRoFmZmb+0kVQPOdHjosEJAQy9/LK
FY7QCy7V6hmeHd8so1U4H2ZNVQHo9qDaBRBWRlpjrrwg3/OUNKOINvqQQE7r
zGsEmoVipeGXTJCBp/5GiG8eebwfZbga3zEqmOJolxuDqDJCm4NSOb+I3ygM
pHwBFL2jvMwuY//I+1YYVH7ZO8VGRKTF/NGvWrSG0bGouUhx7UQjaBZcCgM/
9xX+S7VTvDE7Z+0aYaXd5V6CcCNQ/j67Vqc18DxlfQawdFaQHzqPd197hXpj
qSTz93u/lc1V4xn5wb82l9tb/bKBbY004/TG3n8cmZYf99myD9MGs51gv5bK
qGvIUhgu8VAvCLjKVNjjMUeE1hKbWY+f0rksPv++qZuU2czmQsl628m3fmvL
RchA/S5wHdEweWziyyPOXAbhysVDrGEmLPRDeuJRjHqFXj0iSGHQ3eJPIPio
TirSxrl4zdGyVAegbl6MWfl5mx8Rz+7XWxulpgJoeC/amH9Yy0P7AIYK8pMD
mSgD95ablgjgubAlIlmwkyLBGbuXgFPAgkFoWwtyvXET1gi/rVpGmXjWoEQW
U3MYrHAuhkxlXkKjCXnakEAcK54M3GkcnzU8gfNlRAUNFr7pHpdMEFQNbmzK
GHD5VjAIsV4/KuVK1nMD37qon3S87fBiOHBjOYoZ0HuEbEi+9+rtKmWEHhec
ewQMsS5JzKmamIip4O26XIhcNxaHiTjocLHBlM+fc3gvfnmQONmvt5XgNjLs
TSuilgJDTBRlg7I4U92s2GbhO9OGbR4tMQE8kBwHc/4WQi1URPoGz3FfcpxT
w0D9Wfs+Dw6/f2p6ukzNTxHhAx6haHdN6ln5TQCZ1zLvnMuXslQdWcSkTmE6
qOJEGwazd4M/ZeXBRyb4G/5LdUT4NR843NxxPcKNMpCFEf4Ya+a/igQEg8la
SmrzGBqcaYMD86inU+ltaqxuwZWHpIUnuSvF9dyVbiv84IVH+gD2pJw/Izb1
i8Ko3v6x0Sci7KZAiBvMUw1D04/S56IhZfMFYOea6iJm57Q3L4WqdLfht2xP
/g/qqe53mvVM1HswZzbA79JTgmTLx2IE8sJsYM1Ma/Ef6xZFLe+yQtS5Qnat
BmA/cqxw3puFdrj79Q9PREQdNLiUZMxot78JRUfCQFsLhGNCtBFtfmoCPim8
jtew6F3taOg2RnhXm9ZXNadp+gave83QKKhYPB25mK2gcyu9xJ57ZPWbo6hE
pSWHRl6p0FkezLt9oizLn2K81bhy/dcEF2cCTQkdqy8dQuKhQIoNYkeAT1aL
n5Wfe6LC+rsT1QeX+gk9Gr2W35C54SoIxE66dK3otGhdjBmuHgyxJfHtJmnZ
VA7ScOey/LzaAyE2qOxR34FchEf3weosfc0jvHBhWkOYo2fInfF7n2gzCrqL
1KbOknSbqO5r6wAlxsJbuqe1QLLQsgXHzCz2wy9Hnv3mgEZAhiEFDctIJWZM
EZMHrtTQi2CR24J9IKxHFS2lCn2Urk049mNqSqpnsFvMDDRxgCnTI8WrWz8E
tHgLpVk8weEea3i1wppL2h6h7TYSr4ZbN/J3hgjD5aJIyxTao/10oHIttCvo
hOm+GfnW/BO4xMcEa09iEWYcl90jIcM6jlu21JaHlCbwvtO9S6hwIwwiDwKI
7jQu90IISCDPGSw1c6vXp/1+K61It7NdllebPYmGZ+a1VqggEJi9sow+Y1G5
yXkMpONHTHaPtWJlkbe31zt/CJpJF2cgqMOkWRkC9Tfk3tGmc8J4ptjENP5C
MCSNOEIgNLgfsezp8tr1oNywtrvwU70lxLsCndo/NfTBzXkTKAZYAclbMyRk
WM+NF2jAnH02aq570c5vRCSCyp0CyksuULjZPejx2bLRmSmpNSeWvNSm3sX9
zzFa4Xj45QvQCZ5g5UXDkBQXX13Y8sKNXBzeARZtiM3dyp+03llYLxyg1lPq
WqJqL4j+mSh7gFUTxzpbknKt15uRZ72mg5ym8CEXoUqwsP1CJVTxG9+5p5Q3
f2XxbK3PVkoqlRcDF/IcNbtpBe1Q/CroNlAdlEaBS+6EfFP+DIMz3308DOVJ
LoEWq/dc7PLWMXNBq+xG6ffjD38517l7tohy9vjIRqnL5n4/4YR5v/hg5u15
Hapz0b5xk9YgFEjn8ZlolXlJ4nRVruiw9Elyx3qBgjaSxn1ZYI+yHTWoVuZ/
+jZLW2Hk88mJcpzXLqVYF6n7borbUjyin0S65hRdNnfYGOrJqOveTpbLJLYm
7tdgGIuXAbuf1ekGIFnwqxOhmF3SnbVrl6PsLRAp1V08yL/AkW07ZSWJIN2K
VpQoJCHhqnSHPTCslVSYyQx+UVRviNzYvu9SNMppYxhMGNLKfHSry14dZf9w
AfXUSL1E/DAl9a7blLefcsX137bDWxDVjtJXLueP8isvEMOX9uayBTF2JoDm
byO4G16hoplu6HIJde4TOVd/BNElCMf46ol9q9I2ZuvABVlfKOARq2zr5grm
xIBuKk6FCw77IvAyTEiq8adTBRm95oep+OFG7jrw0qZa1d5PYekIlGAkmEHI
S1RfYw6ed2bV+0/D1j9yEUe+Obvml0iXaM3N58GByzgLGoMGIqTWhsoC7YXh
Tp8I9s/FsDkzGGpWA0v9zcYWLsHv2I1JeXXWxAvbIV25R4ieyFKwTBteYCQL
2n99S5RB9SgWf29YCPuTynaOwJe6Aq/47CH26hQk1SAmIR4xwAuqHh+6sUl0
F7zULdUyDCUviC8lpp34ZMhV5pFBxlWpuZjFPkR9rTdST9B7hDj8G0tcR7n4
HuRF1VkpyIkN5oeQP1Xz6mLUn1kFkeUd7lQhlecHs8i6eI8fQmOau6zQI5ku
1/89gLo/SLDYf0dwBzEdxhybVGNAK9+AXRj/hAsd/f7xe46mBfYP10MJ1zwa
Cr/h3iFGcqPyi3Gep2ZovQvsGKqP1l/2loIei3AZPV+bMAawgiTXVQYkQTO6
444QsVMqb6aib7Wqhm2lqG6P/Wrajby9TS5XHAPDiYAjs3bmomOlWNAXFfc+
+jugFgXW8wRvbwvghtcygA/UgLgKxL4SwNuzstn9kTO529reTKKCm6rsUtLY
bCORxtdq5SMHmClXJNaJYEYSarcIsC5zUwMMw3x+eocEVV5sr4NOX7FBELau
1FGSVtCvD9cFKScmNm0tACOE2TW/BnNhH6wZ2pxyKP55AD8YuxwJwSLLtyk1
AXIiTzx7R/LPK2D9O722wtb1gBGQM731ieQzZUOGc/ETi67K08A5vnC6YJOP
TiGk/4DZitc2QGNwFq55rzcnDinzgHqEeKE56vb8jtwfdmnk2BWBxA7YLGAM
PTTyh0kqInbsMACqUVw6o6u4ZOUSLuEQ+LT5flbKEmx0MXWWVJS9ccKDb0L2
wDsZxdd+jm3G5PooXdxsHhi+CDTgdXaMmKAbPtp6Uddjd3+BwLv3g4aQK/aq
Q4RmncSjsESVR74cOdAe2Q4vRXKnSgCDWT1dlCYkN3W8m8y7pT9J5c1EoCj8
MRLOgNca/VdXxIBIKH7uSE7jHeoGaK/ylV7T31HGMJdvgmPTiK9T/pvmrt+w
7PiYlZ/n0EZyL3nq7ssG//WA+jZHIOGzN7gH8QGT7w6LCehE3iiYarSHx28i
inYT0Tlcdff9wfk2MCHEQILtLU3HS0QHpaATdyVZOXxq2ZMMyiyEs58KeAhq
DEcNGcsVZYZP1A1xHZzhjZ8iEkJjMZ4QSkzDsp23YT3tE6OnLFfYrB88G26Y
BobFGHNGPqrieY4mGcvSZvhVfWp0oCse3RFJ+fcmTnI1wDqDq/Ta7XSU86Yj
BjgYCL1TR0mkrKywzPZNLrKOITgt8fzvUxAaj9M1tZaRrceEq75RgzBr54gJ
o/WnA4u5H4ZFzt4qShu9uXalTI9kLHmPyNI/6GuftFUXWhTUsOHt0kQ8I635
L4yO29/X/BgTRyV4TO67stOBxcAv4Gb/dT4+YNKMgmXeubcviwSN/XsLTpup
OqSyJaaDOZo4RlFqVGdYUYaaieojdrpi2CCUMzKmMsrR2joa/Z5LEEpONDL6
mH92y2tm6Tq3N6rpc7YnVq5oBp+6F4hoZIkAUtVRKHQtUW2QKl2hrGk0xqWA
dsxn1dOHWaoJ3i6DEvayRdI9dzkyM8cEceXm3sir4wJd6mqOR0IjEWqA1r7y
VKNwlV3Rlq4jDUIGzJ3MEWuMqvGl91FQCEN9n4lqMaxWaoy7IKYfqJQpnq+M
7vDaGK4uisK2AJxZk3R1a2oqQX4wgeUX8upzTnV16VPajYdX+DMrwlyTt71b
KiG6jzi3iwBWdUSpuhnkPO9qgtsvnh+rfDLchJMu6usAUACgJZoMXAybSjGT
I6rmzVqJc5dcuQK76kGwjvctQNb650SznZhHSsJtM6ru6Mh7lwQUt2PDPhbI
XaJRXJMsqjb94JDkLkcvBFNzakabvpWav+GH7GlkEqMMtD/2C4aq9xcGagkq
p+/yauUsNZXCDtcej/HK7XdcJz1asYV51i+WcgaqwjPHg3j7njZVcWpCWN0k
KOTI+YfMtj4+rJTe7jS/K62NzDDfMCrXADD+XaMVDoDdN5hRLtsiLoXPyOm1
A2rXuDhMUdvpEQ7MyMgrL1PJ9FM6W4YXs9RNT/V+aiCcUrZWi3R6uGBX3w6h
XFH22vA6NCJJ5ofeM+6JInwYiqVMTQNDoEckX5bk3MSqlwew7UQnK/NgYbMQ
LtVn5y1FhmquDQNbUcNXYIYgAyiqiD0Iq5N8/Rd88OWjE7XwKkzX4SMyrjsO
u3J5/w/G5OoOchBn0physYIMJh/a+lhcDbUibgbLwUINP46lM0jgZOpGYWFu
/x99xTucAxzeN4Ak7oQC52YUsGO/ldQBhW1Bp39QEvLTQOB4T+g1aHnAUMZl
9wASnjNwH11n6WK+VnmU/3k5svh47JxYyI0BdAZ+v/MTDDa6EDXUod0iWCnE
nzI5CMKSFi6H26Zfgt/e0fU72TK4E+UQ+ryGCrCC7E9VnfssViTN+EAcWa5Q
tikPUuIp9XY/R9xWqqn8wM2Fr1+tSBIi4kHb4k0siknQKyJbOUb86xdiFL3F
Q93wKKiJ7Vdnn4OUjUpMvEpBEmXBJsvXBO/7t/4fg3pNbnjYME5x2AxEuuHU
qH46pP9vtyqLJSRUATLLWE865At4EXiJKNu4r1lSHA0gRAP8zU66ng8lgh0L
qvv+F78dcINyIKfY/l0CVXfxMDA/WkAbHrAiRQZxmJstZ24yvM04nXmif36V
Nil5r5uXt15YAKKci5kMgmAc90XglUo3GVRajl4n8anzCPC4fUt0nQoXkwQM
K7e4w+Ux4JOQi+SmfU8fsm9+uKos+sLi7lKE4uzjUI9Ga+owVBK+RpSNmEDH
Oh/Uh3W/v/SGo29fUqgVES50wGvilsqRI3tvHf03EzazLuLNu5UKi3YX8T7B
9KVGrqysQL5RwkVR/8xciiWF62GgvcsGfVXLWu6jWk6rne8EmQvq3DRb08o2
Oe0oIKfFizg7fPAsLAkiKTESYCbcfg9gjd+6tMEuTFThh7V3LONz+U1RqBom
076/7/B+1UYCbrwa4El24TR3JRQXDfs42n5q9adc41QHYiMEKMzpmhd8hx85
rbxAJS7F7WS6sYspkC/Z+n9m4EWWkEF5oWODpZyuiExCq/YadpXfwlOOqeez
2EPDfTOXVup4096ziG5xYb5BUUnr3XrVZC4w7K5X/MIr8yjXvDIRclh6miYj
mqFwajMWEnyG6EwhL6q3eolxs8+rzBmYy9Uyadvpx1jhEMrqv13X5gdXckdL
0QJ11k/JZPeZTQPQrwE91WUQuqe4HCLu7NziBJZlqWUVAukFrriNlGXDUwSm
xqHzyvcdfBYEwSg8S3DBHUnTTjZBJDR0a2KKedIaq297HgF7EjaKXb1K1Yve
JAst4c2p5W+Au+V9M+CQDrzzTlxv9TQqEB85tDXpF9hYH34Hif0yTiYJ+3Fo
Bm+KQcvuef8sUGfEAk/ZPTc8BnzrzYRSAHBdx4H8h+iKUK3DanUBmgqm71Kh
JSQPc72m+aqNx2shyw6wagsOAH5pSAn8L7Q+VUDsNnlgl6u/ApSAbncyJeuX
ez6CKUZFuaoBFzCirOdS6xcwHAfoS4AJCD0J+dbAYDKCQCfPU3QH4fTQ64y0
dY1cwW1hZKTdCRZWAUI28wOSM98HPsWBLfXIwsK/wFXofbBRXMPe6MCmZ4MK
QU9RUGoT1/4qd5ZcduTQKun5aoklEz0GD9FMfd3m3IWwEAlh2eSpU41g6EMn
jv8hpcneiSpCSMstHKfZjRcuS1ExsobZsOlrDvY0h/9Jv3ey6ZahWPxBlcyc
plwmTvGFXthNR4lij8j7OZaEbZwsTXZO4bo4PUmf2+DMtR4WQlMWe2uoUQKv
aHv4sL5H9aYZZEy/AuuZWZ+YHofyEkGSpQgsjy8/Cd7IM5xvVpHcPqU5od9n
fIwiTiO75pUs2wk5CHzXTz9qLo7fFuyw1Oj9kzop+WqGgRTk6QCAE06yUtDm
o5kkJhgFicSzVPiz2tbDLxmWveI31zp98qk+zuTGVXQjTUwKA4juxTNliVrT
JB1qbkJs2i+ZkGn1GK/8+n2/Mx7yZYVko1CCSbnH49feW5uTFYJ/pG51it8P
yngRCQUl8UIn48RDHUJX9vUvCTGVUGVHJnA2RDFhS//FClzsZ8mZ9Xo1+Dhe
ENfnmlOsnCzdozaRFXiO77w2QgFnKsWL00DbMGXflytFf2INnIZnFQWZHtPS
4CRxxnXK7luIOyMK/bqXqtUGsVtuEUsrwtwH6uH08wa4otL0se6yhuO/OQc6
3Og6Egpb4cy4e9OXBfJ6extLW6KXCEKDTssFIBnoth28f8pZU4lSaoG51ETf
WHhNWk4UEXE705LaDmcucGYyFeFn4FE41bpH7NcTh3ctmngsH2xcbwpdnVAd
3ozXufmN97zIjOy/Nbmbaxm2cnFM4cS+gtN+ksznp7RwpVcEiCj0f9gElzRw
zWdgbeaaYLkj9rcHLx+2om8rHhe652go7qjqIy3ywF35XMExD62GzgqGMobP
3NsdHX+Olcne+QnC9AsRxG/+iT9y2k3ociiCM2PQariLIPYLnYVWIkRvIATF
D/ssBEQEjzAvNMVZmPzyPHrtHKqwjYbcLiraR/Fi7KZYr7HH9Cni2Z3bODvj
cOveW4ah3vl9N64RyrRSyZ0EELZ/jaAttKTKFHGkq1SI5gTGkirqBEAgX4Tk
8LJvE5IDbRxBBOrjT5OqVZ91LNZaLUHQsofft9Xb9YvH+s9qReaX7VujJ8hv
GqiBMYJ/zlZA1tIyq7jT7mbZGhPXwH0bWh9+sc2NYGdrXLy/BADgfYbEwho4
rzysi4GxDZkKXuw9dyNQiHjlFVxD4gxa6pkD6Hzcgq6ycd8w72OY6t9oxmrU
aLEZNffqYMeDDc8yu6gwRgxiOd0aItwqsS4sSxTGihu/uRkAsO0wmEVXwlhf
BhQ4Gn2+cLB5dFT8qUqdbNHknfy3wuZR893yQ5nXRqFLAdBJs8TMp62OGqnN
X6OovrI7+IRtBFFKZTcPLFKFTdYyoNg1zG2vFmeMop9LiI1oUe6Y7YLoKK2d
j4CItmRAfClwwgxIYPCjfEqKbztcQjs0uqZKYRiIIXgbLEpuH6UZjWCenjxP
5NB+KwySfwZFxdoaYNlVussKdNu5qdsCg3ODTlvKNMZ3w7IoWnhN+8bOoiSI
5z0g0HOMJkpcDNc/oIfRnR6uT6461KSRt5oKEMayFYGFa8xjtMkCqS7Evbey
+XVYSdUz03VJSVzJlKEuQEGI/KKoH4ilVFmRWHhqyHSJ/JdfoK6DFrWk41DR
hvgfKWEWWRosLl7hOQLI5LzWyToAA9kgHMbEm2FFEKvr/cyDOZv6hFzaStwa
9d5UJbKLPBfVPgzHHncwAJFWLh2dYd1P7299kkSG8FCPB5IvYzPd1V9MBNK/
I7rYQofDmsqO5l4GdZpgRFh7Pi50U3wNy5bzaasby/TEPb6bSTal7unlenBJ
FUvzipZ3ndYNlMGJL02z2f9IFsUQfawY7hs7ILoJO0ylGf9A7gfudMSUNZvS
vLb730V94j6YYYqwpYAC9/opXpHs+ZRGMirxgDCJ4lOTLtVxw8s2ATZuSM2U
J3S6qQW45v5HQx8rpReMnhl+daMxEbgyvkq5OSSNGnbGOnkI4lkdFCG0hihm
k2x/9XPjSFcJm8PeaZlomJyPEne7K/1u6zUE1wQ6OPatHASiAtslkGovhQmY
TFiMmCbYWXGyBMJI67y8puAiaRhp5LnHa9vC3HHbWsLvSBob4DSTxWOVC5tX
y7pwabac3zfyrZrUhwb2zwtfKy76TZ5FftAU7PPK6/N65rud4Nkw5FVgab9n
GNWpNEyO+pCdA2Lo/W3mZEWlkPyUtj/4arLvqlySRr2/Zk/6FALX+yMI1+3L
oohr2C5OfzG1s2nLxLGtef51mJQMr9RDTJu8X48Vi8SPYtJ7fivgkm1DjOyQ
z4Ih0ltr7PTr5b4G8ovA/jdT6C+mGR4emSQsLPVnld9kKgkn2zWiulN/e5g0
t/vqyns5mFOPC8v7BHV8UqAmrx7/8rgwhU30dqH6sbNIsK60Jq5YCVL0tIg3
l3HoV4IW3nrt4vxPawBVgxIv6+8Lq+jPLG4dIgMmPADony0LdAH2DLjEQDvm
irNswxCHpZuxnFRIwxejESPpoYdFHgc25iNA0q6OXhVC2stbQjWMGz2uP6Ne
Cb8oSWP+M0yjtybSq5i2kE9ShTQcqSTAADWnAhtBy7nvwvC9Xl51iqHZ59JB
MlhGFAbmyEvYn12YS0TCDPaOd5qwR1ZkcAf+ikzbCs97mq9RnXc8oeVfkMCY
4UOo4G0gj0Hblx0sFtNd4wtxZUD9e/5IJRFJCyzbvtDl5hNFXCE9HgsX0HMw
fZ5Emuxj8XwF9vMnowuiGuLJylDNXeOJJnsYgeaanuTa0Ra0+mvcfi89dGGM
++HA8QYsKFiZ4E2SbPZRgwkuTM7g4veG/ik9MpH6EpeHJd3pm33YuuU4YEHx
InedaSKlaJ3J8cROHV/9PsUJZUkWgNZQk8mZisKIdYblNz/jYz4X1+fb/NEz
hA7HJe+PVZoLxi0UubRC4FdXUCaA7xq3QEC0YPEb3WHG+G/ktYCL8zWK6NgN
nwh31KeYXCxMxhQX7IguJRTEh016CBhT3UIF6gG0Xuo2B6aPMMUHybDJD/70
aqjOsOr74rj8QYiXs4PlUVXkoxw+GuZnsg7e29QgnBZA3E/HhvCohNhzbcei
V5o7T23lZDvwg+mwbLmCSJHX4loLZeiA21OrxdLgXohv6rDrZOzF6mtIyNNE
2yyo5JIgN/DgyKVUKsR+owb0QPwmD4rjVRLYKjIi07UOFSZFtL+JsyWV+acn
5scbQbLCd/MMQ5MncBq+mA8bmwkQJ8oB3BS2ybRyXZJmGhmCCBnPvODs3sxe
s3BkxVULGSG7qaK11+nGyv0SdMpErQIG6gRdwc5QIPsH86HSgMEt1hBEDBEH
gAYnGa2Bdodn6gSDi1TwSFIZPIS6ChvcctK0e06fg0NrczvyBAu/rEC1lBuA
qZOEiYEBdH49ArjOKrx4MgzF7TZGGr1NXxom2JFxCawWNqGDROxeaZ+R4dpB
2XgHls3T/YZdfMAQ2zE6InRPxjIlnfhDd9kZCR28lPpqB7xGJm7TDgti6cJM
UjkP/Y6icDHd3Z8EqIT2mDAaIar5l99JnhGzUjERjs45Ag6vdCh5MZRIWWu+
JePI5kcxRpATE+Mtj+or74iKpMbGEOxmf8EfzkAejdMmIiX9z2G3YmKlwwzQ
O0LOU0ARvdPQ7s9neHt0p1iQxFQJGQedzAqf7mqvb68KafC/uBmxfGefsl/T
GeJU9Pb2/Wd3eJvEq5F+VJnrfoYaSimrn+CDQiIiYoDtH3cza+vForeymZld
RUfJVfOU5XrWRTJXwEdi1HF5TWCmhzLtxPiQixlGUX08F7ZBdhBGZ+7jdKkY
k/clTAK/uhsqY78JoTfyZp2yL2V8c6rQZ0RYUC4f93t2h61A5WddzmA6KylL
3l383UJLllu4kBg5OWE3HWLCOJZySz+CirXqpWuUrT8YOUDS+/AwzGoIqap5
hX9AdJfidbJDHHhAP2enkm3gqsFlhNPA22KAElnPmJc+j1WBwoEbMJvRF5qt
FAkIfSCdY51kKtkWrWHGT1+TAsGkMVP/4gpU66W4eHC78RuzoYVSFzYSIfsu
9f6+p6U16mHH9rsJNuQ+Z7IDPF07e6UVL9HBJ9FRoogrL6OsJygdH/cFMbZ2
upCuuP3SJeGdofvA96YGreUBybpOCJna3OhlKA6Q662rgh5lH9uwUBuguH9P
Un31x7joxgVy2w5MsfcpuQkrSHBRQpr006Xmer7dmty+VUJTqShk1Z0Yutqd
NO6GKzZRuTaUAYHZL2W+uadBLlCuzOyn/9/ilB/RRMfqtW8oQKc+22keinSU
JAs959TJqHkSvVj7nzCkZz1p8+LJpAOJijgCGcjhCYjPk7zdiXbI5kefezPD
1tIZoBPZ3YTihJRe5jvrJKBnV0F1r9wxZnVHc3xkoO/0Ts0U23HzwFGkP2JE
h4UK0OVAg41CcJuQkVoKjGLy/PJH2wp+yh9JVQZYd5VWKIkJ609pbz1U4qGf
Urhd8yy6XvVZHKzUuSUSBB7LwQlPzYkargjLY3c5e2Aw7sXqTr2Px2Y6aPiA
I4VRFxNiCpiYXZCUot2BtuFv0sLmIHQV8b6bsL4xVi42S9UFeWDxeWXmX4WF
In/ZX+IaSBCHighcX0i92pde8+FhApKSbwfiG8JDRIuTkk8TLafOsP834Lox
r1kUgwcRKXK0dK7OuWS7nAp6iU2ouTK9usz1Hvpev2jg21ymZc9r6voRp0na
tA9TnSZzX7wzm1B0LhR/cozUJVmAK6/X+aCn971PHHaxsQR7RfDiQorFsznZ
BULpN1UuxlaRpopUk46dBjEDqK0R85pGr+7NucjmvD9WNY7xz+qDeQvJU9i9
uRTqyBXlT/hdnoDSpoJcPaZahdhjhIl1xrc0t8+xi1MH2fYdMwSjdcWE76Rz
2y3qOjyuKk50VBvk3FvrQjU3v3SfTQvH3+XP9xU2QPOSaShQBiz9l/DEg5I6
FSYEJOzgX8VsL4XOjuwQLk+gB2j10lH8JKXWJrq07UaUWpnOMXuGRW+g3+hk
xWyqzI5AYpGFTrEmvaIWgzV+1307Oge4B5T05GsPsmjdTSQ/cx19bLVeCIlH
0KC6R7dVQjKqXJm5PiIS6rL06SWySQO62Vt/PcprLEFTF4YAfbEtYCllE19e
T0fmVUUy1YsTNo6X5WmtVGmiqrW2/if0jCZ3I/Oh2Uq69chrDSBGb0KQgk+j
tO5H2TOk2a7oZJNROsyJoub2dAkB3Ie2smRor6Q7poMVsJlElBTNI60CsPz9
6aATw/eh45Qvqa144gKTx15hsInMjPK5MrxdopX+MFkSdLUlF9+vR08bhsFL
Yn9tGfyAt5KUAnna3Mv4NWo1KOEgMJ1o8pGLy6pF4SOm8YObijqL7sIGnhIk
hwbmof0GFPoLZxhoLNpjVu90lciwXGsQOYKN9aHkD4iaj6YIUAbgQnrtSx/Z
Jf3KG4ksa7leXWWK+1GfQ5Y7w/VGjn3t75WXLc/6ErDwatICQqBTmyLva3l7
j2fAsCrvC84PGRqWzv8MifA+JIbNFjOA/raeQ4AM7s6OHYZgD4wYC4kX4PUA
znAxZzMrC8bRryLEIBLcA3jE6d92lZtahPCrnVf7M+UJZJAIU/s63Qylb9el
VyCrXSZYTCoMQRfw2pNzuQvFDGl2Ry/8LkDWmYfPUQPdefUD2wVDrgDIvOhb
OrmqLEjv0Lfd0VTqKBwzAdjileBd41VncVa4thGHXD5LK0w1B7BvNGMyoE/i
BLjcGW3ffGGcZ1Z3lO0v/RYvShxvleA7NZ+2QuYW8RVB0MbnIQc35YdVB+yE
P6CDy8pznvCm/FqWo9pNry8m8zlD67tp1/6wFOTQv+b1qiaMEnLe41lc7a2h
WYTP4TWF0vZMHM93e3ZqEliSe0XhNjAySlRH3S5GvfQ6LJFD0FoyG6zQ2njr
QRU2tojf46/lHrcCm7lGg7XJ53f5odXXNq41oQ0XSWQzUi3HSv0XIVNJTj/0
RBnP+7Bz87xkf6vBrzaTwHIQBqIrNPGC8B6K68aUtXwfbo9397EdZ2Mn4ZtE
chFvadIOA5xGxdMMBQ9+rnhjPEOycBWgTTpTF+d8mVm20NtDpBsn0QD1j2bX
PxSK3/3y1wZ3+UtbJRqg/GY0hr+5xQgxCRu6EJR/ol8nzRatfUSnH01wR9O/
1cEP+XjqrqiRxaWeG/4yzc1F7073DWf4t67pRXnCxAJ93xeKD6aps9JNAavm
PK+Vvr4qr6CdMZfXY+te9QgLfGLFqnPVsQ1Mr4la/qddi/sVaY/1x1orH1zs
VK3wvd71Qv53C4mm7X9VJUPvVXJo/1tzh7RiIJPTDlin0igVV/N42tqRBdDd
j7+ck+Iszpmx0QUZsIkxy9R/+wEimSaiekQH9P2DCvzI+4LoAwv52Q8jz12M
kn8hQvebNsFw5LPJUhfeYiNgIMqkoRVzaDQjnL/A9RvaVayD4qba/NH/eHaS
xDCAeJM8AYNZfCGsyeYkZLfxGShrYmbmhiU3qpk5Nzlay72X8zhfiuildQYp
EMipYu7bLgyeb+DqcoKJ/+bkZyWDys8zPoMdIwWINE2aWFoapnZqJAfuoSCa
tWSaYAo9eFVHkpQi8mv1YhEa7vJaqfWH/D/GydX8Qbhwd+bSva2GD82S8cS7
1dbAZcQvOiR1gjnwcPrk5AKZZnORF5qhrGXxN9LwhoMyy35vsZJQqlqS/u5W
NcyZty8NwT6sLzRYyE3dkMuHc57z5PU6mE2yMvPggSo6h5HLEEzzREXF43TG
yw7VQmVoGtBH2qTFJaHEQZNdEeQoaQAuHzfkDE3w7TbvgEv0nfXduJ9ApcEP
nbC831Nt97Dbn/4i21SoZW2AAYCoGi1vFpML13i5jbSaY00dZlSdu6YRVQ5W
dfn6xESyx8MjPUBP3DrnuxCp6QwuR1iFNFO/qNXJzFdedIEAyPN+3hQc9Pue
HBGX895NxYG4ofuqDyO/FlQRfpHxzTCg1XPbMIcWPh5XjwH/k8JHgFqbnOPh
OeI5pO5790aYknQfGvho+RLtCtPigEMr4H6K4xFlABXJdl2FWcfvx+bODqdw
WYSkUpgpOK5seMFJzxTnYlVW1ggZQMezZW9aLKfc7iYCCCofvfsss7allcSI
j2M/eI1yzZR/mg3hCpSZ9n/+mmibXmdZAD/IuGoo7SDcyAeypga3tC1QgLts
/ogQBDAGKL7FpWMdRhqHTyz0/YjDao5wa2yAQboP8XPVAgQpQiRgDUBrwaa3
9Oe039vyNV1AQXJshsc+2HEiud3L/cI11mCcdyJlpqPFzFSbGm3ETnwLV9wc
J+CFww0TtOcD1GjraLEdYVriZQiJPjwfwPdSg+tVzBKElXEIIA54D8JJ8vKM
qpRjIXmjCMSxkGiHF6ASh6Jj7IWUx82Cmk4nh0PODrd16LOVPey2wKJQgU9H
4uVNJxlsHA2O8X3TYGmZ4CoHw2zlgVsp7XZuLTTVXf0u3e0QUNLZ1L5IBwgz
UdS6bViWhjNPKxW2lR2FU+xz1RKusp2P/4prTnH0oDeGirnGflVZzaj5B395
tMelRSniLgB0vzElx83+JqtA6g5Nhxd6ZW+swZz5setd1JyBWVL8DR+yDvLg
C9K37m0Y5cFyNX9QapxMKjk3D/EtfuosNXNJSl2ryjm10fO9xQvZP+VyzBRD
DsifwBvvvZGj+8mPgOSXLb4gQdvsDh8AYv7DH6JESBXsEYBYAfTJxG3wcxp2
m9fiQLtpZ37LpOgDEYSR/mJ4NOA32AbOq2IqSVSktHOXc4B/wbttp3s6797U
iY12hDTRjYt9alKA+6521p7j25J9vULJVOleRCywcm4h7OOa5PLaqSgrQaRL
xqFG2oE71SSCxDGb+zSchSINJjvuH0AmNAtOx19kTv7suz2dUfH1TEhBRSFo
3BVU5YmJkaYvPSpPs1J25MCyYWYzkbfFHc1Fv4NvJjfEOijXqGGlodtLk5Bq
2yqT9iNCUXPAO9rWr8VzTAqaiL3wo5Lwmx7lJIqbB8vFxU8P9Js3pznfzmbq
/Wqc+rcWyuWHLoqG7sxzkMymt4Xq3bj57nX8jwAABJ9E8jXy2f8ghyz/nRvv
j+XwBxtFpfNBdT3ywpib4z5HvpuSKxBp2bwA3/etW4GkkccRYhCdO4QDUiky
guM8rLdZIrCZJxQk9AFSePY5DuI9CLzIi0ELZ8+P/zncun4AW6NEdYpEZYKm
6uqKEzk5KtaIRLUUtkXcP6lM9DYCfvJ3k6Xj+3qZcZrxLprTNWViXYn1d3os
0FX4c/pJTxaC+l30LUriVal6g8xrYxBBiTK2Nx9dHJMMJpJDojSx2XbQB166
wqZhh4o10pYNWGSTi4lKoCz3vfc8m31TdwJMap3YtWwGgowKfIkGfU0Bs7UQ
g43y86S3PTepm6PFYk8sWVlt7xCYlIgnpzkjPH2VdHxmnxntKWdc4mYkGEW+
gzs5wooA5C2Z73C9aNSLgPd9hh/JhZ+mfybBF9ygQjk6o+nVHFwDZkhIAGsA
ZhihXVSsd2VJJ1BUGIxPjfc48fxsw4HEpdxuYJtzyxBscBgdcnkfL5uvpNfx
Pe4XfYdwBDHKLBt74WhV1zIM+3u1gkFV/294NPaBNtA3xVfAOhqp/wDtGfqI
TY/aVtMF+x/NyZ9p9QlpN29Y4JaARqrpOZE1/eVONm/GlQJQYRrFtuj3fkL5
+vYJZ9lmpUPUUwnv/d8UvA/DIdN6JYAHvTOHCqyQM4im79jsSYPVIPw+SOgc
dCX18AGrsH0Sbv/Nt8rNLxkgCzJYHBN0mlz9Qm4XKYfHkmiKBPaIdY3fFHiA
N8eKv7zU/s+nlm9z2jCDhUZdddtpVElfiXxXBeM2Fg0h1K6eUJVh+6j27Vg5
1TE6KpRWkQZsQ6Ns2pmcgpKzHov1FLQCMTG4cy7UfhIkbkJrX8gb0O15BLqu
snhxm+fhCE83Wff4tOWBOaHjAdkg+b4WMETZ6wXhyk3lnK6KfXu8N1A627ch
n7OfYX8FL9li/NU8z/rTzE9BpaCFlS1oBHuznv5UvYGpLhTJLpjJNvFjrM46
uP3TdORf62xK9SN7CHbyKmLs3ai1gqjhF8SM9O36eAfvKArVGWFA9l/egh8L
NuhC0uo6bFEl+DUuubs9tNswQyY63rb6G9dh1V4YDfpcdi6f66LcMXQ0O7nD
ugDOl79jEXqjw0DteOMUS3K/PTD0EJFFUGf3SEWFPnBQsDWuXowi059Hn2qK
yP4iWWegiq1Bi3EepucVfgx0up3CxKGDpqoCvYNbxKor10ERBy+Xe+3KWg65
N2jQM/WWvqOGbvKsoV4b5Z15Aeqipprgyc2O900idbPocvxkDjmPAkxvijI7
Uk7DCXoSKzf/BIgmbwbSMsMQoLCUObsQMqW+3GjMZxyMK3AAiWwjMrr94qUs
3xfMzsJCxUL31S+krXd0Xfu4fTtpVnsXE7O+L/0wiKKiQBkL198lNEG15eWn
i3GNN1N7b2KFG3ZXO46RJmsWw1Pmss49BE8CyNTmdjxefKDgv2B3Lsr6DuR7
yx/n93x1XoWU6dG/TwROZ110V8G9xU8u0WmkQNFlF9Xm5enD0+38pUtSOWCg
GbUudq7nXkfcZheViz2sfotNoNzn4C5U5T0q1ROWVWFLLYuAAEtWlqFx7V80
vC2ulR3ypu3u0V4+7tcf0GrOiba2bwyxZUNLf0tK1Np9RXURM3Dgu8W467Ww
FFpuWf/yMdUDItfJXFLbukuoEtgPwSIkQkvpwU2mdnMlbRMx+E5jFNnfImOL
bZBKpz1xTDyZ0i/FuHcZM16ftFzRO1Pk3CewxlTr/geyAmf2EmwZNz8KD0Kd
j4T6/oxGa6bIyVVxxJG2xlCPG84WnbdfOzoF6HjGC08Y9GvtmYrgDZNNA6fL
qsoE91lr4jab9PVNfIrBg8cAKd3o+ErQ950xmUOjtdViI/CTjRYRVQ0r46DB
waHX+PGwrs6Ysn2Lo0ihZ4Vz5Fx0IvM7kGyJUwF3V7I5t5txi8LeJZKmOCsq
ByMeCD+Ul7Y4cqBNwgYYSs0eYJyqPGG3LgiHAbzc0UeVG69+MTI9jOaziEHJ
Y0MsGmhNta3+20UD6o5cfAXKDkqS3VdRO+92IkHjhK1U0ieniX5AsB0OZsYt
V+4N2aAeG5LEgG0fY1S8dzHl0RPWevz94y58O7sUHhREaqCuR/xCKcvN6Qgj
pQFrhwI2D2/2IrwRjGtUr/zUJYgJRYhODsIQkn50BXSBnUufrE1D0b4BF1I7
M+An6sU7BKGuSlu0Jl5iIhRV2Ufmh5L49BIipex4gDkO72qW19niK8ivzaH5
dFNohsEZzIvTTqMzS/JYhgk4SBqW/PnNUwHAyv1vCLYK7dIad/VF6LLiIYmf
v9AjVLLekjkDxwBvFq1DXF8Lpe9oOBZi1n7PyWWwUlPX7soiv60HlHj32c2n
AcOcRAGaCdpUHRku1hBi7q3GpkRiZ/Wc5Sn6FDzpwOzH2ZNAKEfCnqJwdg0b
mia3X72dj1z80w75mIsiOiFaelq0/mU0dZhB2daM+WGMnCmucx8LheOzL7Ji
6UFe32LQMOv+4s78qbof1Sb0nq91quSJhkTydfaBZvuZgusdx5VG5gKFNeF0
9gbOppAclBSb3PWmHE24MKfXnouOc6ro3gKw8ze/MfYs9/KA1iHOcwyra0vK
EPUoQ0MpPM2BBRglt7/iwE4yJCXx6Q2EVlS6+5W/cYcIhB6fVm422FI6a6A/
BlPJdpE1s5SmUnjFbQXDJev0g+6CdqKFo2u1DwyFpG9hilDO831Igy8DFn9k
N18PMggA0cel7DxQmjZafH6C6QlImmOD+jAWv9e11b2/yUH99CEy2CB05p6R
i3fnMVR0ZtrPJCjpfcXl2Ps/5JClZpRAc+PIldoOmMyNN4jda+YSnb+Mnujg
J+c12OkU0CJJs7wEG0iZ1BDgKN2BK+2RpA5u0i86+TruYmONSN8CjAY9z7+J
xUK3Uk2GO8++vN54pKahh0d8TB+aTQ4Mk4J/HArC5Nbq2BFlsnDxYOA/Rn1s
fmqZXj6foiN+rDOWcYBbGCCmZglBrmx1CrBQ7d7cVHlbDATJKcEFybb1TSLc
XqsaILs3A63+kePVtqVp5/jdkkKU3++87ZnuYk8cqaS0zFdHFYOeRzjHsFhc
QSShATaswr/7o2JXxhZ8/h/N2QV8Uu/w9idS/uvgqHhRB5bm2ErsDjXaDZRm
jXqImv3Wb36UbMeqcvYHIn582SA6Bzl6KfRtwXVKbiBjxL67nDT0s30Ja5T+
F9DOnGqKLFE44XLOK4krl4rWQqrfaCaLyBkju1QU+8wFxbrMdtmXfWCknC3t
eFs5+nI+/gd0g7FE+3Sq+HkO27A+un39Kolx1I72XbY9jclGyXduqp+2/oPM
sVEmBbik8hncTOTrhXKwa8SdFENnN/4TnCoWHS2qABPaqiNvVyCNNON+KITG
aDiKBiP8quzs7zI2K+SgoMeERE+gt5L0L6sIqEjlWNpP0WYtx3P8uaSNwAed
lkmk/u30NNoKw3/ts07i3z3HOxgrzLWGEM0/EY2VY8wFv+2m10vi6ylQ76Ed
kjLiINYMMtkUuW/vpU2POXezjlp1L6xJIPmtFxSa43PkIGI9SRJ5sCc05JIO
LXe2Ed+CTH+bxpjwBYVT5Vgg58FWHKm6SI4Mpmj/lSbW9rMfYY0UpXuyGtHM
oJHh6pC5q5qNcIvAyvaY/5fCy/6aD1I1z58r+QnbTpju8dBOPhB2n5PKR1OJ
au/NXC7onuocAI0if5mrJkF5qMep9VnkNP0RvZIid3wC8I2Owqm9Bm8sdbzo
Xt7DtM3GuY9eQ2lcmEPqGP0mR9+PYYNokPH0M8iBguX+tmdf1deN1BXuFS/G
wK74jkEJGKwiq1KaFGiv5IaXqqW6Y2C4ZB6DrCAEdTtvD5bLYre8d8Y/g7IR
wHUl1uiv6VO/ufM2Cb3AT7e7LMt6DPVPUNlwGAiSv6dTyoBMcO/QQclE7s94
8qp7Dq/zl9D4IORlIOtLcONv2UT/Q8grcxMeo5ORz9HaOQY3Dma42+IPjLbU
6H7SSXfzSXiM7eDvFUocc+3fwZDppW6+GPv6Gwp/d0RCxOCGRuw2m48lcsCM
UT59KfAoHxfJVqFdX+Vk827GZoE6366UpPBMHZ60hlhm1KmafiRUJomb2vE6
+XlX9hAP4nN80hm1OwQ9NJnru9OzvzXpPunY7XYHNr0YC/gFczZYRh3Rb2YR
7sS+UaGqMfIs1EtkcDF92P/wZg5R2K4V5/bWsuO7X40ztCX9drsoJxjFewEE
7YUg5cyo+N6L5DHVO4O7api1fxGauyBsAgQ6pVNouNthECWyrvB+UFKfh1WY
zUpG4xsVhRKVDW1Noskgp/CYyZbLtzToTJPbTDr/BnAA/+mOhgqsHSIyFa+t
jnV+3iPxbOO/M7YKWxJyFC70QZy7mGWQLFOAWgAdbkgh11AiB4qazByhIf7o
5uQDWSxieAIt506wbE/U7wyVV79hj+AqiLFvRTmzLNVjwboyFsV7aXw8Tlcm
rq8kJ8ldskNhbbD4HP/Wcaajmjitn2G3JqiE6yNbbq2kifnqyk46MZvmg1tC
sVR00W0HIpdcrSTg1GdSt6SoU91SQmRNq+oL0J0c04O+u4YioTuomTfvEoIw
/WrNG5wzBDdXFNQSFd4L2p+nSOysG0f6kzqMmJDNDj3f0sfndm8GU/thIU3C
4q2sPKYdw73c8iTMKhy6Tyb6KFTf19gtvg7sW7lC4hC7/Sh//sn4ZQqVOrLI
cZHHmyRLwIpLEO+G70dyr49jZ+imAkEQficKjxlX91PW97BJ5DR3VLPBRBAx
3t+2Eg6/ff8xHlsvTevEI3PAucWIVUGFXZdHJLCCbmUrZ9ItaneSs4GfUr4O
fyyCIGBhdc4rf886x1y0qe7dUWbeCMn2mFFJvL0+2eVCr+FX6S5DHckOo9Id
PNvvwooACpRB9kTj7WSH8OsIGVHKVf415OGNg0B5cXhTERH+JzufBBh0URg4
FjoDC7zbieFtO26hcG4PxVL1nVFLrANXY6vzxfrlNM6o6cxwd5IaSTY5HVH8
ZIu4yVHuKXKWSrjl+EWOqwShNswhHctsJWJiVjT1sbFJMLvmIBUMVTh01xca
sZYgCJqUt4+IcN47916z1eJR4jMi6szCNXyRIDfG0bJA+yw+49g83QwGvGJE
2Uq/Uje2tB6qk/Y68iPqHDhYPWKunbX4gnrRyExFqDAoF+0M5N5mtY1/nnDd
q5D6n1KwD5dkhNBn5w4E8hWKjki1Q55MqbYeY5Zmj7oTEWcgGeQRl4HOILtb
85xQSAP5XpGkkGXdVF0uPe6+0r8s8YfY6hL2vGVE7qLfWL8Mi9MUfrthb5W5
pDQoqTw+/1w1YBiJzUpiKPpSsFZQifWKGT1o/Q/YVxjqIEvgAosEfdHbI7sz
fOH8j1FgchhZQbMESQNTB/Ns6KBOTMv7xqKEWfYkP7kgq2yVQkIX+eBL4CA3
FiKS1RDFOTicCHiqnBwl1meNBU9Tte2rNhv/Alxt0rsMNEBsrVXp5YowP0OI
WQxev1Itzg60RFvztdmZ1KRGnwzTiQENxscol5ptb/9WzyUhCuM4AYa08ieb
B5JRRXYS/G65TTUHHzMsnZk9TJchx8uG2SuHBNMJ0FbZHQvJ+Sxw7qTzTrSs
KaCuBeQfR577SkgZHrJb0FwNUfGFB500r3RvaE+Pm0gUKvBgVi9uU9L3zo6C
x/RyRQaYxhxlNhlGI3sDjJLvM+DrZ3zuD9hcw6qEXoSH4cTXxQpjdagJOU8I
f8gXr4f3Rkf93GeJpDGzA2d+W3VsOoSEWQBCng3iMmQjY2pNp82GZwtliVD1
HUPQTt4e4ReiGp/LEVAIyAZ+KKp9H5wOBaLIeY1wVN8IsU678yHK7p3z0oL5
cMMvvnWXC+RiiGJyes9Y04SKDDarEtvl8E+q6BNVtTJfUyOyshgTQtsj6ySN
qyH1UkeEVY8LwFh1hbtIFXnhe4HeQPqkT++8uJJW1Z5hL7rMoZEcecZcKA2A
t7+3sXNcQveyg9c1g2PX9t/O3u8jf1JLbMZpGYp1/M06r2VcyCqxbxXS45+t
DwmZ5dyO8ANYk8oHeEnLsteSuf+Z6zzPjPt6i4J3LhnbrinhqtSvWoOCFrfC
bOvq+72S/PxljLmt1uQRLuv+1lk1dJv5bZ6iXA+X1I1uXqMviNt33NDhXCkJ
7dNggmM+9KbaMZ90d7fOw1GFgk8D1/vvC78QmMTJ73+6I+EFiHfqL0LgJh+h
YtDMAhet2w4+24SUSgQ7Z2QQqpsHM3cj7xHQbL316ia2kRxbI0daul0iHXm/
si74t3QHrkXyT7bi3WTnL5qdVo/kT3bAcOk7E4H5CGb4FxLxXDCL8rMxiX+n
U6Fl4YuOktDlQvO9g6XdnJQKGjmXr7JchwAl4eZmLVbJTuT5MJk1bNMVb/ey
a20QtZICXW5Hu19Xte3Zyr/EtFGL/30Jpf4y2He6kR6yvVqT0VQYMORW26AZ
bhL5WMSlhDi85jInVF2c9cy6jKUK9wA1kO7tXrnZ3ftyhKuXkrLxo1wq+iag
soLffHCZzgh3enamRUUA8Lvr0tHrJ8lUfj5dWAo9SrciYfIogO9RjeQQv2os
7WMnK5LWhqVAev6QR9AqyavtBr4/4EuxYIRj8L99CRb0dOq/X2eV29gJAMpU
StVF6COXqPV6TublWx2TnMq6jC/ry1yUWCeKkAIrQf1Tb+ewAXYfT9YDxrfY
lGkXZcx0dilQMAtR7Mfj1DTgVXSZtAUtKHc375ezXNvRw9uhy/9oQEz8CGuH
xLFtaGGlnRQu3LpM7m9O6dl87VQ49pTbq2U/DkwsMUGVRguv98TuUgIYyqAz
NglqJSltt1kDuecG9KwmT8mannGz8CqJu/d+e2dC4/Yq8Nv2mk5MnoVV348L
pzZ59uplpjnQvfjyqxKVD+CmFtfm9kFzwSxfWWBGH22isSh/MfD4EI/f1cGo
1qxzFT7r9O4OJgMFLAKcuGpX7ab7kce/XbmQXRNw/I1FOP4upx/r86E10mdW
bJceFBuqb27HM/8+OVLdACWmM3NHDtW+RwoLZZs/9fVOTAOtsQaM3e221NNJ
lvfAl/rw0KaC68VO2hxiKd50j+psh6HLAxT2shh1rU80ygMgXu+0OgBTXPAc
1ASzpBTKnz5Q8M2unlcX4BSC3EWmoJyBdw2CQ6ny/Uv9a8bJFe2AtwcmZtkH
V4n0lmjKF6JBfHEhUTDP7tlpqIA5WiotVh1Q9qQfFGM+kx+DYxEvRjKESqF3
68pgylgkOyMlwJzwBY3mnRYuMlOS4LjnWH7s7i9MoTVpookyJDsOM/Xla6Ta
ya1pV726jLcmeHJ+ZqbLgCYPFQy/PTzrPOh1xscwoKc7KcsMeiiFsaDNm667
pNt9OAfX9L2Wu5tQzl0rudO2aauRa8FbE92oFmjBw65MbIBmN73C1b5cAH3S
C4bIXOXFtf9/urhtd1emHhMcVCmlVdYB4kATHnjx4ule39O3LwA3r/mzI4cX
j08IDIexQ9SGdTgtKXIMHhU44eN3kDFy9CgptX9qeMjSNTcq7wg4afoK/MrC
03tIYxS+9jo6nutO0dSkADpJ3G5bWhGu7J8poMVdytJQKT3KAyPs0ptSEV2b
si7Z02xB3GKsy+VKiOQA7fgsmBiwlXDZxrtRE02nazAuAR1oisFS5QX0Xf72
cRyG4FdTREyG1dThq+4FBIyriQTCMRbaylKUzWPxMhr4N/dVqrwr/gc5BLyu
u7fbBOS9WglLgQKjJcVMczztpSD9UlEApGdnrs9gRsFw2i5Gthe/arkQZcSZ
0OXR073QNn8Ukd/M+v2rdqYa5ApthM4h2VQLvgZGfi3OSmxgbdEqTRi24he2
p5nhC6f8qCLRcYPkqRglLKJbCaEU4qiqODxp3ZC5bQD1tNTCgKaZCu3EMWyY
jgNXd86d5yik5azm3iAOmG9KH/L2grTnuDjen6IWYUd87nUVWcfajtAtG2+Q
AGLHVZo3ok5SmRcABYHsU+/xkZCkq3+fbA4GSJKeLH+cwlHxzM8694FOTIaf
m8fdX+IM39jRjFetEpOaU63KjAVhMaJoOzCpluqE6Oslk+3uWtDmdNtocMTj
csooYx6WwNR1zVaXmlySEeXJKqewc61CLK0PcA9aDW31nYG1EjqUBGxKL4Ll
rQp+R+tILV8bP0MonNRUzs3oDYFgSAlf3cc34I/lP4rW7xmLVZ3ayXFH5qYk
PhOWKZG8wNACEFCZqhrjQLvEhs1xzyAYlRbqmeFU1w7fwroRVnZ2sFHh6GKF
2OMHx2bau0yFfvImLBtYPA6K0YhPlkQlC1yWWU8mawT31A2d8iT1osyBQvlb
AlNWWvxhVEs7BP2Jz8FN+Eg+PO0y2eCJNXSWORnclGw+Bx6/nx2tF/pKsAIf
b3dfYUhCwLq9qyK7JExFOMbqWqjcsGRznkDan7qEfqp+tqSf8XB0GCknnkMv
yAvMuSm6xAH9qMKWOGWnAdM1qwp63kLe6KxwKW1UV8T7vVU6fAtQo0nFliKB
/lXLmw4AsGx5YUkfI37iMGXJE0H+FcvwVHxdlYaQQ4xeU6IGWglH18GO3CRY
kyxaKKcqAtBiNGg/lp3HWleff8qlunVMyMeOvOOPiH4By5r0J3WXq49mteHO
EzXhOLPslNC3V74AjvrnHICGJXvPU7qCl9qQRgm19sSNhSozICcM1M92X6WD
AsdGWEk8thfvdlDYJFV+Vpp3FHguSR0041PZeOc10nI+m7vaziyJ4fkYo5ly
+qQ8+Xxl8VS3QSp3Ev06vwVBw4F2jqRCyK86hTMrQLR9SpzxaY4cZeojq99+
w24ZzlvdC7vhlCsq15A5Jh81zjLufhcaoZa0Rfu55ClrsVLzbvv2TAQGt04h
gVOvRbtJtp5JPWxbV6XM9X9Qx9nj3q5BZdzHdp+U1gIlFwEWIuSOyEv7AonD
Gz0Xp+YHiJDUBFjhkfjNC7RoOfHda7Y7WisFQtfJybtqorLzq9MkXoofkQ5p
sW4OILuG5/bn0oyKUWtR96gS7c4PZBx+6cTyyvaE8gaU7rFDc+apMHGahwTq
hpFAKsipGUw8iOq3ZqLMIG45W8ZsOWCNItJNgnefuUNvJi1/quK6FbzljiFG
sIXZjHBIxGOtcUrVTU3WMg7dDlhb9tDwDQj61AobeFbKBTaMo+eX3W7n9Gvw
92huwK1PWRBD/COZTLoe00v0JGQIoYHbgxc3G0VYlIkmjFLs7o8gJ0b222B6
kgrhVeFnH0I7fCM/dEs+rCUb36QZB36EVBabcLY3aRDhMJ9IClWZPJnUGk2t
wERNWvjjAkHm90CE9qCp5W255IZyeHOxRW/JK6kh88Sut8nSHLyFOrpXMagt
+uD9AbvdK5U07LqYKpl4Bt0d9csv1Uet8spOk7PpMFeur1X8qCjolvTsCUUK
OsoWytghRqYm9NpIUEQvg72wmDNaI2SUVY0uXYpsqDDw0SUwLCQmsZfSkG+c
6qMTs6JukoAaDPFFPcnbgxBWSs5kxmHx0UL8SLmW+SYavsIp0fJS0ZAHdVJH
KEZn7ZkErjhpyft6T6kP7tPUU/2/rUeMuyj2qf49Ri0ncMNM98wdcMQGyTrP
nuQMKnFTScm/jiIXyYfN+A09lBDEopvlZ77zwJD51OBKIUz0/BKse5eSxKEp
jTYJSNxW6sTUBkm9O1sRJgosdeoSBTpa2iyrIX0lJgKNTlJOMJ3tML4Y64I1
CjGla/OBcm/1K8Qu1JERgooucVTjlSvmUmlhv6Ny8VDMGWMkn2fOBAl/5y1g
792n1kR6JTML3ragbO6VnYAp00MErAPN4/b5C4aTV3bcpk0pXsmtNlClOtF6
aByDKKBaHNCxeJZ/6ucEwhy93e4k10coAGETkuHQNRsvmSi+e2Mq+bxCd74V
smpiUVgmn7XXq3h2iXv29WMDTsysoO+FIYmbtXAMDfip0iL4AN85HXSMYwWS
exGatI//oeIPZUxZMF9ClZ6OYH1CvCkBDuL7MvBVj36MfSY69jo9pdxf4YRu
v0yvmKoJDnguh/CfnD4DNh9tEDtv8is54K9NTzVCqf9iuueqveLMlJEJa6em
oMt/axO3KV6/5znsWDG+5Rzcu695spl8caQMazbpRwtWx8dsJG3oaNZ2nweO
j3ZwZEtHy6kSKD53a7plH5xHM5PmtMpVDYAtcOAPXlMF9tQn5rmrKyq76p5c
vslXAOlC+iexUDOTG5PJB2pBvrRJUPDe0fbq9OEv6Ls9f8IvyhaMR1heoZYP
Ge96Hrb3kyxtMLZiCz7USvWas8t/ogdGfpQzeZxxQ/s0l9X6pUfIN5Wna+Qx
MrnLrdo8LgW/2GF9tlMug6Em5A85DFtQFcdFaurARUNLDDqjxWJ9vKCA2xc4
wpVBixa6w1j024qZJbMXHLQgQWyxPSl3KMnaQkjEtnFoE2epgEjqSpjFoD2Z
j/XRTirmoMFYdhYA63h9UwFZ1cPB1l0PsZEyiiDj5d8nxsyQUK7xBLqNq0DR
HQqtVuDRWalfmf+D0HUjtOFYfP/uoZv5G1bhUjNxG7R6YYDVOBTu21yA2zIL
vDdxIJPlvEfCDgkEjdaF8r/NRzklm5MgEYv/4MVunCaqIw+4SE79TyvvLqwl
uFlAgso3SQ3kaAO1Xzd40tXSpAp+B7bOnOiQTOfrKBr8VVtC95+TudiNaPhP
ou/+iryfA4VQ9Fc8ogiRLvmOudMTXwHZHeArK4WRKe0NP7RDufCkwu0SXBZ0
PgBNNBkXmME6ggX/G2agD8aPmQDCkHCiimkFmtPWMRDBsL7LMjIaHuN6/F6T
/GofyCeK2pzJdaEKMPPd/eGfU764neoS2lq7V+nwVOzlPk09HBac8qtZeqiQ
PtxGBbJfTtUmGtQx3FPftaJ5CfgqZoc5hxsAIO7iVYqdaCjSCTn5cFrwEIom
Sy6d7HnCYzv0GksLcTMHKQwoGAqwDVq9A9EBonTjwAcNHoAU2AOvm4NVdAmJ
Be48wApImxZVnh6RZnR9pFoLGjmx8hxo/fwC3xBefptAEeMB8Y9Y3m8M76uE
ER19SNvZDm99Is1N8GB34UL8MBhkcSYExr5Lzog+vd6Wc5vmNzV5LYm8DJiM
wF30YES/5pkf4JGrl0NXOlubqGO/dJB/GZb+rF0CYENdg1BxCY+YhrPjSDtA
X7rWCSUXM/bG77Yc3TtvzquEAYmBPFW6k16vGXIdiFndbSuW+QHvl+tx8bRr
aAZguRla6nQKrUzA3T34Pov4VqFBzCJnfK5pTYZe4atA9hkg6A12bQnkyE/E
4xhy6SvlZxOBLSnstFfn03sTD0nNuBq0Nw8AZMTXAy7LS2SlTDoRmpFlbguW
A3FTLiGn8HgxItX0TcwyMbcfh4Uzs8faYuFgWYTvSGPnA8Fg+6XfUYp8Ct1P
EfFfPWDgsTpSwCDYW09tJ0LTYgiEFyRDm6J8/mQyqmuKyMrBV7vQyY02QvIr
DWILZ6im6DxOzKcYZyoiyx00r7X1qELpdCZ7gx9C9ROpwRY/8QgJtDhg97t+
gA6q1XEHh/H2pzChMhx2rEzUJpOlQ+J/k2uOLrgFDEoM0ymceYTyqT6UY3OD
vMrncc3liVaGOXaMDeDJ7Fxh2BuZayn+vZsShEFTJ+yxZ7ILyqw/J42i1m7A
FVES1dlEM3uIxuZ8OaXMaMC/1ZKVjbVN3DEZTt9tT7HV1acKaRksvI+Lyy2N
nFzQX2Et96ZAhuZm7fXTKxjjxX5H+vC3fM2ZuhL7D/3moA093c2HlEM/fRde
eU4JoPmkOOXe1/WtMdO11E+9aL7X0ptII+PUhHFWlfHf40RfH/w0t7alUXy5
NT6361D0nAwK5YOeFFlZej9k85WaiGkx6QVsP7A4JxPqrPzEJbHq5Rvt5H2c
Iz6IwaWMaILeaL5i3EQfXf1HUYdTpLO/kq/+fchzSzwjwXdHW9u9BVxca+fQ
rjia7ZlHuPHG5zsIB1NL2qx4Z3NV3/AGfflj7LGem8bqs9yg7ikVBBU9xSpX
QOCQjUj3jTNO8yKdJ7zrAJHUrSjvPI/QT3EbpuDCaTl29rFZCYHt/LegcHdv
GC+7GrhTo2y5dLJpz+wFBn/Szofwuw6+oziO3vlk/5dcAtvMMaoUjRPlmrJr
/VtB+v/MmWYjCkh0O3GA78BqKVs61m94wQLi+6jkVNgOy0U5fItxEJmf84rm
rLA/5RQUDohUE7bQMIE9lJolHOndwJZAd65zFYe8R91e/d3J4tsMJUvGonk/
5Mj7VYjc+vzHyazAc8f2ZNbILYHOF+52XbqSJBJTSmU+nDM9O6IhmTOrelTk
lfDjdnJiQowBtRfCs0E2U2TPugX2IX0YsBYfuBBSg3f08sVobPFk8TLpTtsg
Vk1a7GsthaNlc9hD+R49O1FWSN9NCm1AYfX1Ql+G5PziRyLEGTjEDEElCCDn
29+2JSxG9WpBOhXyj52mv+qDPUHK1oub+lH/2aQfsWgaKQYHFCqh1CwnK0An
E/MFvMq/5FxULsvxw2zGVXg8qZt6Iyt506uTVTt24KkHavWF3Lb/QgHMerZl
yoVb/LwMLs6GE2sN5NMHc1iSYItmNdUrIdkwDPiCQZ3j4mcuChs4RBPtfTb0
oITZz2NVSyT6+lEI+yf8D8/CXyj/DqAQ4a+dc1mTKRjfkVjuRX5vMNzrxFR5
a0hdtaBDlu+knW9BGHeU0myZvQ4mtBOrxP7Mm6+kZvOOxIrn82AiNbwu5mRO
7kNOafvd8z1/SX2oKWpqfDkRCRqaM3dLLrQIWdERCgX48X3W7MKJWQHG6MXm
HK3LZRMPpAoi5QCWvb8O/Dp39dRU0XfGbtwnsAxCArfD6VQE7v0On4ZT6jPb
108Tin+Jx2+9Q25sYnqDSAyNuFTQq63YBFb2qLcrWaN1zWAS2oUXJXmxfC9E
jDNZUkrJTJZQEbk1ck++UBfzZswMIzkAW5IRbTXYKzhwRphYFyJN2OQjEUO9
J37+7nZ8F2vPQFaDIzPXoPci7u7JwBlo0meseKHuuqgqhhvz3FGb9KQ7ojFE
U+uBDZvEEcP5JgpmT6mKMbo9t82TgteaU66nBkz8hc53e459/cMbIaKUduzm
hOqOq/5Ce2sbJ5geTdYXcsKIYFJcg3PsUyilVLBMPUHHpp9iGza5e30KISnG
OOhJPai9lIy+qxKfv1ToLzyiK9sq46H64EwJbotK3Xl8lovsgtRs4X0DjJwB
Jw9+/7guktSuCc67dOmzNGiYK2jN/SD2IXWivKYR3bXLknAUeOoukHVlQbye
0MACi2x2xJfDvUTcKT5gCbdz4Im8mtNPwclbOkLc8sxu9Cs4CDwh9EFM5OxQ
Lg67Gfg/yrn+Dg8KMUIGsA79goDdJw58f4nJytkGp/2s07+nT9aFhica/y6a
eFOcFwra9v/oL9aSNnnl1fvL2nVzBxwLGMMOvuRhswf/esAmg6n/iz+dHGsy
8ig6eFVQIxf58C5sZ6vUx6DS8Pn1Ek6iBoV3glQBi24wiRe4i78KqQto5Cm3
Hn+w2vW2+gcXNzeNQdbcbVYO66vU25xLXsmOOSGUxNuMo+Z3mN/Yvb9bCNwn
5mQUW25UgLLiAdnnC4x0LGThAvppMcWUqxB/YEMKb7Ij9c073lsy5/ON8wCC
Psf0YA1Uxz+ypvoeZ0GbKpoNqbr5j8ijDC2Gy9utS4N6FVtWoziIU12Qg/Gz
rwCfd8dM/fk7v2rgy3e4YUSwz7EPPt7QLGAn5LbUTydW9GPP5ott4JKVA6sx
vg5+E4//1bmOzb7dVme0BPpArwWjn0UYmpegbCB5ECsen4ybwfEe/LQHzYFx
z+CrzxJboHPNxFMFZIC6OurgjwrbnLODJDCpk1WLdOuZ4O2/QULp3O1HGRJG
E4fOg2Wjs+XvBZannJv/Niwdl4s1Mb1kMCamZYnpJflmX2NWWRS1HIpDlfEF
1koSDGBJLWxf+ujjguQXo0p4a1lmFQZbTaAlo/Wzs26VKvW1ay2qxlVzkqgP
2sQ7RDA0fkLrpw8MSQPwjYz/oXUJdTB3eAiHZnAkRGkfcyFNrOPZIaMLEZ03
LcWbp1yXmiHZH3Xf56GL1L6fBINWvvKjImcNHmZ8ZDaxL3y4FLExViueQTyq
0JfVnc2s9aWkBJAU6MuopOqQpiAYYjl0HPwfoIlZ8epFzQRbxydGOGGn9NYh
bQ4AvPl8A5JFb/J6nPhJMZIeXb5pJOnHv4mKlwPukoXX1LXG2Vo1R2q5jbdU
r0D3oSrQ5A3ex0/NpNpqqln1n4BXK3FA2Yj3PWFsydCx2MlxdChymP2zwnEt
re6kzJXuYevQN7aZalsEy1xQ4vAYaH4NjjQuI33grxFLiB0d4uDIDmSYc7AY
6IFkm6ZxqpzN7ckes0GQoTUjVa1JbahexVgeUKkjkMKE4AlJbfnjpiJiozH7
xiziVWj7369OpFonn38CH6Fn0YVfK6nNVSLfJc5IVIuAjrHyOCAbBiYXQAEm
faj982NsQHFwvx03gzNpXJ+gJhwyKYug0L965ZAONcg97u/W/eGSYSFoqjBz
ZngLmYt8E6HbziIZaBh4AAt1Uwjxag+dmWipvU1MmQRVsmxGxtpEwTOVZaNl
xGPJtb6sP2UT7xzFBzSnY/JSw4gajfSpZCiGlQmrOU4h7z/HFUTRPg27AT2Z
JtP+ManN6mvqun3GsuDBo5uDfg21GOP7vuHGDGlwidTH+Mds5ryosunovYEq
+CORT8iKvFNCaEDCQcBoxH/UTQUt3xIOjnlVfQIYG50oukNu46Ca9iyVzqus
MdQ28BHPsibvJKGZ7GXcI/q9Iu5HOvbBe7w7Ilu+7enlsyeLFFb3faGP0HPi
ThlfRSdqbw5Q1Lg08L75OzEq/4y29VtOvzcqv/kE13fUv4iTvIzLXvfmWUdk
e9n+vABfgXnERfeKxtOJQJZ51Ai14/+2gc5X9qO4Ka3ZF0baoFpuloPdqDJx
b3EB8TnrHOz56Xh2uClpNUw5fRy2ThNqHhtd/KYSO5J1riTqynV/GEKrxmU8
A82YEGpPVH16Fh650naJ2YvWh/y24EOKxAC0/goJpGfcvMod9lMEaXx2Q8GO
Ont0Wm9h5LcMBRefq9PgEGXUr+zzmKIfBkycnnp1kpUwaePUfGab9f05G+hw
BoevdUEE4HB+Lij69ZrO99efzAwoBQWW4X+EihkIPQ5OWruyND2v1NKbJ7u5
qZLfS+dENH17j/mzxX0LzImQ3ZNlxzEfbsASjBfGBwhrkGefHg14uiF/GxGW
kbX6BAO2Ff1nfLQE8EllpUDl/pUlYGW3Cr7HOvAYTj0RylFL9tj4NMDQ8ldM
8MX0TNXOAs+viacyhFE17BmfvKXX6muhbRIIchVGB5VTKKevxYR6trExJ8Gz
NvzWWNlQDBawaKoRoUCWqpvlXM1NgRpNrum9J1GU0t4NMt4T1f3LEUkHTY6F
d7rUfChFS1Nix2RGqfTJk5nDvmyP4M1PKv0v93ntWQCfq5rwxS5z+kiiZtm+
s0kAG9zAGmKdo2e3pOC5EaVurtd9yxVsKZuvEiZL6MB1OwCdLSjFhQ7qsMJE
XLl/yH/P2KsiLTUaXu3u7eJ6NzCFyy38LcA3C7Dxy7ZdJMSX/QFFJH3M03iC
EyBzSneROwsEoyTLcAPKNbKlp+ReFnpkLXpl2E9B0YLGFJAg0a/A6Fb8vBIQ
LNXwQL56v6LFceTnEQzGop+j63fKx9LsIDvmZljUnUogLuyL1jZEDM6JN5lM
4a4YI3soNmq61whbl1/YNQ0HjfhZVnmLRU5e2riWpvPU+wHCV+kmmoTrg124
6HXgroLkJMW7hTiT913Mj6PA8V4eq/MNJJ7mdIMV7rZ2lmeAdh6my/M5N0bi
CjsMxL11rFTjX9sjCJlhhpiIRp++bKp5O9k+bHfjQDBe7pQn4ZUUn3z7ve9B
NDd+y4Ew7egwNUOqYEBCi1EjQu0YHTb8w/L9Zgu2zusbmfngLSghuFhNuSs+
zupa4sxXt/QWHSK1+U9a3R0/wvyV87gVFjhk9QQcmdxM7IDgVhho9Dt5Sv76
rH8RtwzsIlB4famwr8cpv87UdhYT8yR67sqczn76X1EpoaNek85RFCoYTfKe
yeuAf5lEYQfSdC+6n/KvjALgnp1/GP+21FNHd0woZFKARGPMN+WasPMWajaD
ziYVeZVdLBPCvAIMbh2T9xd6hw7n126OV/pGHETiey2YNAaELZXVfjw17oni
RSYsSDGD80d0Br5PVJiml7VTwzrfKpihzG/V4SGfI7KHHisSPJLVjSAUSWk2
PoDDp3YkL35g2In90bz2RyxkfA29GNsf4ExPHM7peL1VPBSoVZl8qRMlekha
O+BFOJmGy9k3qfPyeaQrq5ANygS+9D0M0b4vVLmstL4xbjBdmOxRYk+fmvq1
pNbqj+tCARxjUEPYNx1CAFKvS3hHlQrzzzfCDgPWlYxfCJx5zIXmsc0a6qOH
gMum+Em0aj9XfYuWDGpeZ89l6BJ2Fs88QBg4vC7mBt8BR5+PpSYayCII3JI1
vIrPnCVXPsdWfWyHJ1EvcV+CPkC39v5X5wMWGOwRsDRTl3P7im8xgwvsqos6
qAUOUXBqM/fxu0G52eiNuMogkUJmoV1t38Ne/amXYyZlY1Mfw970w7OnKDU8
ROKc3e/thRm3rF01my08s+LFrN2F8S2tSLWQDNNHAfH7kS6NMndE50rhg0P0
iVcaG1U8XSoYy68ssBD5Im/AFvKbVczeKRCq3iX5eTIMoirzwdXIZLA9NrGt
kXnXNPcWqZX4lq83Lbq4oX/YM56dhsf6MEG+rlYUJI6cmIfsYE2YYFQ1vvkc
kufmClUVPvzTAMUXvw5jug3n0Dv05YMADn9eSeWQYr5US3Y0y3dxp1BU/CiQ
eZBBeu6AdqDofRAYXSCI2mKhBAt9NdidAM4QSApuOnjHY7FCyULnrWSTIkdI
8Yh9Lben7HHeEB9DtmM233t/61oTWEywsqJqSNWu86euuK84+3Za5Pxi1b0U
xorsbMo5iqNgIAB4qd7K2B/d4n0zIempwk8wQR20UawLJ3ehzitV6SBE9X7J
/WMWoQ98M36667cGEcjbLs6RLxSLNvhwV/fi0E0vioVbWOf/5l/8Hebt1sVU
M1jgmcomu8T/ipK+beA2DEvQxJ7PXLoJI8xk6oiP1FQrExzJEzgtLYk+g5GB
11dW75miZC3QTNxqRgmktmiBPg/xKYJk6AsP4z7wm6scG6i+7KAmSYF3+wQ9
2emNbhsK5reHHGgt7saSDRbrIzzq28/DDuQfPW2nSSPD1KKGRwcHqjP4elAr
Y5gS3z85jRtNP/tgLBGZ+r/z+Dj86QlQ4c9qj4Tkksk14W7k81GFdyApsU18
TMmBKz+d0LqMg1wAJglKK9ORN+RgXYuPHEg6ISBlg07dBqR+Vpcwe++Oh7Ui
sTm2FJvKfAf0x1SAmOFrJu2itpRLlaMkxGM3820oxZ3A6IiwNpt2/0A3+Euo
4kF+5NBstqbQnR38F4GAaAgiaIIC4XIQpMlb6J8p+k9Qcg4QDxjI7FBF3edl
fLsXN9GKZVsdabEPtKYTHIzTw1qXS8VDe+Q0dBhZ11z+iD9WzVj73xHPNoDG
jHj5aG76Aoj5Z4cgYjI9jExGTHUzlaK29Z3sKyEUZXGxUTx1sDdCGE9fmjyN
18Z+vX3vU6O+FlTv64xN3eZafq8Z9sungj6OXJhWCtxdDiYob/TogCVvky1O
E8tmSJTYaG9AVfctIZ6nQNi2Hy1j23PPXaPFXMCodW05/t8JvAddu+kv7J5/
JyqfPAJRvyUIpB5/6KJN1QPWn2aea5s9qc/n44lzrSFsx+IqwnLj3w5PBYNV
Aj3vGLcv2CrLOwdMFY2mYk++dnfEm2uaB1l+Zp3Vy2jUg16R4aRo95XH2rVA
m8bnSw0LpYu5wlutxSasf3BTQ7vf9GrBByY1/8aT0U/rafAyWcvrFlCjFiA5
5Wlu390wmq0bqUqrGw9/mgJabBffyI9ojRizABLd6dDdBw45Qx3a8rzn24ug
0/XjJlUmmh43NZ9rEy5MRW2eUZlOll6hFnyhGQHIuLE8KaUJuVXX9Q5W8b6s
XdFdVjTr4FB7xNyP9Nd3/yB19k4IFbIbo42mN066UIW+mdIWIqHagoANzBPx
4Tp6PSxYnH0UTQ6pmjmo0gXNPa3XEI5uRaOWZCt9tqyznQPe0ryK4/jZ1gfV
CAr2/m7QOQtBP4oaSuyklFS2+ZQD1jBfUb/fIPfpjwonZGBjcqjHGZcOkXq1
XKbk0D5QU4Glr0rQvq8VMgAsiBnKuABScfVsHIisTJfbDLRH8n927NpUV0n0
InnQk7uZNuwdollFqIUvXbtN6p/AX8Wtl83SGsGGCy6Xhk9zd7YylS4LHhmP
ZA6CtRt82wxUgLyrdKAxAPV6vXeMRP0ZwHNAd8Mf8zrVl0nZf5Ymv388256W
qGKzYjWlcdVKfP7EDUhYvc9TcAProEDYWDGiEEJcyHmEXX/oJSL89fzH6es8
R+1wU6y5O8HvchdK9MkSBaTu/Ta+Uq7N/i3rUMhqzkC20WfJlZ7vXEP1VW6U
MyoZ8OB7x8pxzNV4Nz1l/4bGUnhq0oiCvokVrqDWC7BhhkXfgXpMVyhhxmTF
Zpo1hMU/w68OLyUHyXZlP6aZvkoz+zYsMz1XhMRzGcOWdkprmujbe+CPgN3E
dPLqCONGlmnjN6fiuOOG+lrthkdvEP22Lr3gxw+4S6rN2ALCmvIVMk307V3O
vrQ1bmuseyYimavg/6xyvsHwn9QRACP00Fvp0vaxJWBe2UOeIo9EUj3SiJi/
KjbPrcDzISMavDk5W42W+5fEC1DoY8vntVTAnAa2jMwV0mehz72pcnllCI8X
VmyNIjdaHiBRhc7zE7yN4Te7AZMZDano3vu/l4kuxRNrNGB69DepcmpbxYnq
oiTEjRhLBHLhlmFhqHMyRFiWrGPKQxBkfTPqPckn+MxuHtU2KXBWWR6nQa+G
YqQN/t5F66Use0dnD8Jua8qRNb2PavyKwaZlPvdDr2iT3AI60585KKkuz8Jz
QgfSttD0H69p6907l70KjUQHo1iMkkLPWg1ZtNJLasFP2azL03NGrq6LCkzh
2wAd0qie+v74RojV16d7902SScMHjtLx77T0Yon/HY2d8XWFkkLn/xa8Ijw/
+z+9J5dGLmPr+x9mveU9Ozx8VozAIPGSEOe/TNlYxEnYaatnXJXfU4LCqL+B
EvYv8AoygDgWxNTMP+drG3jFfSrJmEUH4YjTvLj08yrcZ2W6ID3BaRxwLmSb
14HfJ2NZrDtgtGpHQYAxBw2btfWGn/JRBKzS+zG1oEPlIXiX7tQRXob+uuw1
bx9wyItu5waDSibFCJqBNz1+tck+xZScEQznuHOgdpUInJ1HLtt7Q4j2LuOZ
OwaeMwA9tbQySMZzDQGf/++uCE2ZoFSfAuWzYGiTcriV8cvxHZ2bQrMf0ogG
sPYx6bfgs6DHQ26F8yrGJU5+bAJvQclvOPCReh5qbBOldqvGPFG4xPbGTwpt
mr+7XceSl/lIbCnkkBLBbJ9cpcvj4poaDhJxUp2EyUL/SaOBoHKrRZF3LP32
e5C9rlG4jM0pLSYVcqzFUFA6KN7T5J5WCYsMU6Mdt/5dYoYC3owoHnKIFH5Z
fLDnGyRjCoD7OAYhX+vICctXVfTxoH1rh39t82IzJt+u2UCbovPzBE6JXOvo
pdAhPKzbsWyjT7J5U2h2NuZiJZcnZmOfjoTjDxEDkloboby+ZQUpUShWjfAQ
Nrfd9ZJsYHMv37BxxwJ47D7o8nGqCNSVMRoTdy8GiJkJL4AAOq1Y5/YQIqnQ
QpLgqrFH6w/yx72KNmxl4E9pN3CiGsXSWGyS4TwrCLjkZp7LR4Q5xJl31fAh
oAGb988YSh+zALLjRcCIAAB1AQQSHbBpD6ppEZCOl4KRD/IXrh5JgTj7MJw1
zfAF+qGOwicCpmgScBbkR8qBdn/lbUiNhkDySJWIU2AigwI1Tm9if60FI6Ez
+xO9ghMrWiUxxUrWY2HawaA4v/Q7U86t9oo0q4kaRLk2oEMU1efJZ0IG58qB
aB4YKrp/AVEFB37ouvsNTr2c1zgeSiAQJgGdIpxba6bdpjX8JUMJzBN1W4CI
EjCVuBvKf/UdVYqnpH249/IgMUrk/M/6Pkwzu88aMPwhCNKE4zByQHq3zfau
OTsAUQJlpKYYc52L5y5bB4rjkiRewdsfmgdOGTotcfXjxry6EzeD6JyRhe6K
404lkrGhgclUYZWpntCzXtt8hDrV0/jE+umce8k3bhyN8T9/f3NU3Tk22IKG
+wh/97L8Ihc3LLk+Q07Esy7taqn4RTZmYLMG5fE471khPoNmV+WZIvMrQgRn
6S+/QNAC9nZrZPd3hZVdX60SV+hsVL5bSUON6WxC+MWfXvPpv+zSl7/Lphaq
6wxDZhbzw0RH/MQY8Q60X3HcRscAdHBUVfOv35KVMYai1URR/9LMdeXhKhlZ
eTpWRoARC3pZ3CQWS7s0kSBTM9o6M9oMehZWFcd396Sn+cK+GTQOKYkTPqS5
II336WIJBpyaQua8Yi3scYtGpb0CHyI8VOqCyJeKvmc+hSDGi/4lpxzG+Zw9
1O3BZlOxrrVRCAbiAd2Sai0OMCp2JVEQkxz6TrbG9h21jE0w6lkWrEC/P4j7
bTD3zDI6J4LUrj1dK8TC+YhhXuLUcsG1k38wiedoWPmm2d3sHJ4h3i92xNDi
gw+9l8CScSLPuj82Q8JSSxJTUfteKp0n4wI7VeZYMQd3ejKT6QzycCzDLrhE
bGa6NR+7xNRTAQ666o50ReUjJAiXFepyOpybjAzNvfRnO0zPN7dijXk5dic9
/g7/thapj9nwpwyMnwlnKXkkCC58tgwHsR2GZ73LIvElb5TF0Tr7OzDqXvbK
GHgrMpIz8J2e8pesKETQLrPwNluO1hjsfl/wnxwl/vy0dQREzm9xlytDPlF7
3E4cvuvas6Bz9rco3mkuHHUd3wEhxiOYvyCOVcfYJ/PUFCLM3YV67eOqevcf
T0PxKybzX2rq95/SuDft74lQHrpHwZurnMhKDj5rUM3ASGCxD274xLAt6vS6
KQAe+SIeTtf05JuGZh1uSF75QzSmUzlIyVd+UyrIWQ+nZEhGUxzqVhX+dPyQ
Yhmc9co6Le7FI9HEOa9HR1V/ke6wUGV112tkG8xu9z6D5MXDlo8YC1gSUe8C
6XB1GXhVPotVwUJdutPIFV6AEu4kt5ubwp/yTSPlur4SrRVBmC7G+ot1JR31
iakP8EQvvlO9CPrtUW4pkz1UZuaiZVJK17U1CNoFmPewfLwCfZMKsAsFjr6z
WYVw1+dJixhR3JV3+m9hm8WvPDXsG7/dlkNHtjPwU0XHV20zSAh/5dDcbHD0
vjY+hS3Lk46WLrSPcBG5QMI73JGUqs35+jUa/wHBSEUdgYtYil5y/RJhMgOX
GfawaQzRP3QYqO6KBuThOlRx+7nexRX2vWuiuX+eZAY6CEgtc/cafOaJ8diX
Fd1OeDotUwcZNtpM7avn0Lz5FB1JyTWYl+r6+idLobzXf4F3Cwx+VcGznq7V
NJQiGEsqA31IR+LhkfS4pX6Odv7ytq9IIXgz4MHmDjw30mQb+aYApghdA+gi
4Mtl3P6gY3GYRXPRdoslKJ+iU0OqlBxpxsBeUwoC0jg7E+Lh6btN6EpftY6L
0Aa5o2a5GMwoSecsoBFoCgkEq+On4a7uzqtEKPhSflMYlqlTMCk8jWpfU+eh
1k/uaTGZMlE+r3r+jCHgwSBl7CVhYSpA8V/BaJ2wyJEeD1/nnsNRwkeKiWL6
AW6YLKzvlEOlvo1Rti7QWD9TN8FeRDifL7a4JYC5gpcq1izIwhTwKLiSfdMM
U84x1w6MoTb5Mei5G8+G5qz93LMSz+b11lU34mlaLWrrD43QFdahgDaE5vc9
cGN2GXxMxnZYrMxH7hYRvftngoVV4ek83h4FzPqt/4QRy9UsHnJl4Kqg6JK3
57T2SF0XqsP3gzLLbvu7XToNVs/f047Wv48MCA6NlwBIvo6oGYlGZDqg+15/
aIoTpo3cHVbBrjDvEpaY3E6n9cdaUJTldjg5+CoXLFGGRx6OdsSDLkRRtVpa
h1k94KLa+hLW7wJIOwIeWiE1mgYPxDMsAnViSnQP0ZoKYIt1nx0Ga0gCtOfI
kYruD34AutIx/Z9cTIuDx7BhfEPhMyRRxKkYI04VMaMuziJkfdnFBaN8dMaP
rC/n+JXs46x3n+Zzq8dLQnIrRafkVrp1VhcExwpW/8a/fLEPEHFIhsK/HFPI
UqrkA+7dFS5Cbv1wmcAZsiJyLb4Tj+lup84ZWuZleV0SuiW25kcBMgxUFE3p
V9BDaEyaoX4tNdAfAdYA1AcdB4eahw/gJcGNoHqSngbsdhnB1HrdXJGhXTwx
w3Z0ZAsFhTO1wM+1nechMWrjBXECEOc8eG7V5HpFsBNMLYV5H++ex1hqofFS
hMMYDrRPMl+cY/3ALtIwjq/1d8I/rps7+m1fEmCvtDtzWk2f9Kwg4i/x+1XW
28WYDZd4Q2GHGgoyWmkUfHNJ6U4J0ZcipmqyffWy/YriP2RwXfFQdk2zS3Ve
MeK+k4vD/mAUcr8mub/c0tDWEwmZAjLJyHYYIXEjX5IjuZjkgFTSWfH00zHM
UiltzFjTDOBMT6618e4AHk/pdfaVnthFtWVUgQh7MIrPnDsLIUPYfNvEFrtq
s3WOkDKOQZG50ceMKWH6c1xU192ZA3Ou1SZ6qWmucBc6b8NQIG6b9JkbYIg/
4c1aHDkM0X352pspOpIUPNUH4NjkH8MXOgyxkKYKhD7PfAOV9YxT4fcb035H
P3/i+qTYzTMb9fK2RZkjfiVD9sq91aX5LiZa0UhrwEIqOhJNoYTdO+mUAROt
AZexyc0KFFN92miJsBOU7oxettSmgWIJzx1k4NKRE1PClE0L5umI2vhRX2p9
mJJSkqSjDNeKIFSOYCjM+L74vhznJjpmpHfwO5fGufgTbbVN02KQ0xXYYlRv
AnrTHAQ71eMUaUbfTlgw4rp6Gb6OtGawg6N5gUp5LaRIaXJ0XHRFsihA/NWE
BwWvPZDKrXK44uGdmKrsfmqtC1ABDqOc47WxuWHubrkBL4lSSKjXEbczo2pQ
0K51FE6bGgGb/bMy5nm2x1EcomgGFvTNjRTOzcqwXv3dy7naqR1MDRUnkkgG
ZASbxWKEh2LxZiur7m5JdCbh9My2LjEkzgZFe5KRaGONLLBIIdg9B4GIxdW7
CGpiVdLiKYm3XA9Mta7aA0UQ0e7kT2GHtuk67XS82nIFapf7Ug7cW13x4EuA
7mc+Qutt9bIpXlpJVKZfWm9jYGbxYJ4aMFkysp7u/JQ+t0DcywJD8Z8xnpq7
9JOtkyMoNoiiOeGMYQDrpW9WHrhBnqNZ9tThvxPpAoTlivhrdRKzXUwMjEMK
AVGDzOWJOkLiI1KH6SQRRIki8ALTxyv2KGR6rtKJo2Ci9jx6cCgsCBZQENmI
jyCXSdTOKX2t4z2d1Q50dUAkmmwd/+FefGlYNa83CwLdZddmEATYg1xL5m+r
Ha6Grkz9jyDyl9LA93IO9A8WdRoTvGTqlql0hQRynBVzwU5tF4DUa9CWfcOj
OvvrA0QDV1d8nbhWhc474SdhW4h+baTl3BOzHPoY5Ke9NKsr3TwPFnFvQxy0
qTCci2qZHM8wfMEm979fW1iPCg1b1+H5JaJ7AGqtmMEJ+HcvjKuszfmwOf24
Rvhsg+oLGoPhVVWC4KhcyleARJ14k3La9cejiGA+auLKYCO5uxOleL5zn5p+
olp96QFbaZjmKaImI6s8qu8avikntQYKwl2Rd7l+hN82z2ASvYZXP6vkd/HO
g0+pnPnYWenzJEOq19Of72p9T+rJIUMfyNrdu09QzbSABmwY2LQbpY6kotH3
BcV5LLB+W58RYRsCZ3mVmaH5jSwi8GsVWntpvW1XSefp0YlzlnZF83/QU+sv
xkDz7GsZXsE81C5afKeDF7NTZpBQYqOoiErLbluPBojyqeoY3L3waDgE+Ulm
sF6/3jig5YjcefuaUnJJYCBcAfbkL4j719JeeYo2g6BG8XDxAfj9DlVIQaHx
H/NlN8ck2ODu4iQdglqIdo3PtktM/SotyviQp4kfZ1JqFXyXLabaLpHgMWmc
CdCvi+6Fv5dgh7qQG7mIzkXFQxfHVhzJeuA/hpKRjZWYDFj2k7KKZt7oLvqK
XRTLLAv9gydl2avNmSWU/qnzvO/pDFeIpcs5BEFp8kdbxK96v8tWNM4Bvr0H
qtTdpb6leRmncyRHaaHVns4DhC1vos/dgOSn2qL2cezdIr0q8E6a4pIwuyB5
f5T+7TIo5270AEX+mb/QaSvUOPjXDLa9GdYZojwb73ACpLW3sAxYgBuLOnZL
s85qSrZys4Vo4mJHper7BgQwhnEgVPyUvVC6xYBfnjEkoIJaSjGI/mzUqLrh
kMhhrcafFayrv6iDxBh2cHIu0h3FruLu1DdRBXLLMPhgtxryCV4hpAVMfIVF
4dzABCAzHk/iqc/F/ugfAvjdDiEtolYEfeR8PCZ6C/wWONBFtq5lGc/R5OOO
RI2ClFZroJU3u77jaDp6PH0SPJuaboLSRqd+l7VMp3toHhaS39YPj2xjZvqB
eqVVrCv9i7IigEr/VWZC43/WtdgtmeVkxsyiaglNsyOY+dC0YFk7aRP+U5wP
IUt5KpQt460LBS8DT0kn5jEF47WjqU3XSLYI0RdzFObLlXvWEznGhLQG5zuK
B9zQ8dbdewg5Gt0jqdYfraLLXKqb0WqXyWvQZ4VrISz8COEVVmJIlXx2a9aH
skpUprp9aM8w9PZrGnGhPhACE9hOiXvkUQdBzySIagq3wsmqzmUFdXaNhqf4
fJq5965BcVXFLvmE98YVAUQUQnW1CapjjFsSCuP9FW46nKh8RgQRWaWNMqk4
f7lKZbzW0LTvlvibDFGipHMcNfkiHTg0T8dIauQuBt4HIZwlclUf2nn7ktKP
MnCuFjOSrFfd/sBXvVguBLnw8lHh6YC0YAeSgWtICbW3mTPwdpyTpMdC9B2r
tUNN5n6sW4PcTRB1/KT3t6WffGYGVWwD7JNffGCLGddT3F6E+mJXMGMwnzn/
8vfNvD3aRaFrv2IJwwp2udJceJNN5PIncMDdvie6ky1D32yHlRZcUrnU+EOu
PM80WQVeWu7XXZrzkslDD8u+KRV9aKvyr7rpwtN3G9etsJXHid6cLnYFWmb+
LIf7U+qtBIWeT9JRVhzvNusVSyp7qqB6oTyQtQd2wmj6D58f9hkYkhhJraym
q4Cs6KdHXM0q+U6USyPVvzpbpe/Pb/gjBpvtD27rAViWLTOgflDE0ThtNTbz
ilZ41YjVaYFF5Qn7NG7lzK92b8JUDruqlLPsFKTl4G/qXWLQBbptLuzubeSM
oCTR+4b0PwvCuHqLuAZ0ynxnSKp4l4RtwPKvg3g2NB1eO+VG3Rr7wVD33S33
Ab2c7va855B/b1vQTDLdMcPy+FiV3WDeOSJVnE/RGy+v8HWU81Ul07A+7b9s
IE5XJH1if+sHwKxGVvQ02/gHnStOyyZWrIgu4ihROZujNNW/YTDuMt4eogX4
0apkXPacmxqS0+pAAG7PuJpMvWyhHTN4mTh71QmNbE1IiCvUUj528Q8EDGlU
rgkHVRLZmO1++bEFMGspJre4Z9aC9D+xGv4so4GIJ+bSKqBgH+0s+9UcDvJ7
kWwGN3pshiLvUOQ5zu+92R6TmkCTpSQfBhKyFrQN/b1DEYrlByIJye6+F0EU
zeifR31XiQUIdgi3aiVtZK3TIB7C+Z4Es+69ovh1VY2RugNewYCkK1Smkfst
yUfwbPYNsGkIDbEWpkWzuf4Bw7UFSQi7FpzW27uJCdGhJ2x/gntNNfZ5C8Dy
UYNMCl/AI53B+3VzFjP4b4a+CccPIv9oC3A45SPOmV1lWRju6LguQVk7//Zx
dGnb9gq0gzkm1k2RIlUYfsWH3Ae3hO9B94g3d8DHWs0UioYqr2AAOAxS6PoD
/V8y3f3MhQKMp9LZJnHgtkjWh8uAbNP1fBvNI3JZHdX10ohJeOdyWU7r38qk
e9eZ6misoTnB4/jR92CM7NO1Yqsmv5VYuwqcUV2RqlSGidvgfIXXi7dGEdN6
3Hl7AW1E1haAZxsy9vWfMxM64EHzJK9w4QH1BWdPwT0nAnMVVsTl46KzXHna
MqHfKmAxal+1CX7AOV9lfsmJ0y7cfsqheLobZSvQ5LZuaq5yzbjty/t/kocK
6YNwM0nigL0q81Z6Ed3LajKTJ6U+WiTPxcyTPuTgllEEihYGyo14701mzcUj
F8aO/UHguAcqi1er3tif2WoW93vtMi40FikiCz1MrzrCwjxHjbPdqQJRSp0Y
gj3yR1y8IFdjR1K7idFQNg+K34soe1ntyncBnYhruWpawgKDxG2oIsbTmbKF
XNxle7r9N2rZcoTTHq6xs8otVO9bbXkBeIMa3/mQMwF9hGQoJf1nG7XVT8FX
rbrDMZ4qsPOhAwf/A1MnmD/PRgdytz0QYGyBuBGkEa9Xeg4xEhaoVsk209Qe
LvTWJyro8myC2V/BZJhLfQ/T7XN7ogqQVxtL+PXzcUVPBTIHnGWkhG2/ldnE
WaeHSJlOgRX46q4F5Mtrz1soLFUYuwQDUJ2NNL5llTE3PKnMbkwWz/EuOigV
J2LOgFhP15QjCYNp54x7ZywfIztGsbLYeRTYVoNzLu2RfMSevPGsPoA9U45w
JAHnSJ+6G3uY409x5ymGR0tlPVWtA9y3G9WSrbNY05jVbJRNBr/TZXQD9Axv
pvsM/w1vkyojtK2TQoWS9Gu8vQEqJYeyFLIGoiN/5uo70w8IyMDmOVZs5ohF
JuUbxHgOBFVodoCGiSPKeFWTSqxiFp2/5fwCLrbZqLWUg8CiJtaXW5/bA7es
KCFZ+RIrHMtAGyEHErF83bWlc2Q5sl7gBaR3gyhpnXtw4Cf5s121oIxZ2lMS
/cvd73876EZdUOUFtWxu6iVF3KoceC80rjhRykiP/4iIOW9lOI9lz5uvBRxh
MGj6uR4X/LjbOJaMokeZnp9B+Y2OE7853NrsOZsG16fRuNlaBIyWWDIl5EtE
4uIfk8qqUsfgLry5Nl94duaUq636K3wuCZJi1twxGcbz85n4i1Z8yLxDfmrf
ie37FbIt6VPYLWj7Qd0WCUQUt0BmvE6tVvkoNh6XhxoPJhnEB9K5SWUtv8Pe
nDF6Vm8kRfi3+vbSFFaYxKQ2ao+s57rCzc7a7cdOJOSNl3xqvxxpXJEfZykq
ptPU2iUVx/DbTgg15QY2e8YGeXc2M6fsvUHhDu3LmsIgEV3nNR9hebsTXy2L
e0oIWpsgrm25C3SoK6a/WV1Coz43YvB74s+3MrmwHXZsztGTG0/3Lm/TFnh6
YrSeoultAfZREwrrtmxjWImk/0eui/lFQuwMEMCKxwLwi+dXAoBD8laQwbif
pV5w3DEUvjilbrw7trsFeZgcUkZKxir9+eHT8UqRZIqjoRmpgtlUlhezKtCM
nLTdXkckv0ZMBhcKpFChcXwrnHOXlHHaD40QpIgjbBqAfITsdhE7C3WGco6J
2ZrsRCPH0GRtEqZCDgKv8ofRJF3J/Ybhd9QNMwdjAqCNFHqdDL+Y3Xd1x5Ti
ilsuCXs5BBZrtb8Xj5GVqCjd6Gozl9qPlZuwXk9ARfRYQJNE/jjbEDj+rSmZ
zLbZNXoN9sIduyyCuzrAo15QZtxy6LMiTszNsfEqHdpVdmtqo1D7YgIADup2
qtr8NuT4TIP/N1csOzHxGw+gXV7Y58QYe0wj7RyAmWTEdtnisS5XWCfIpaCC
cFG36UonRn/n/NhtU9aJyBdQs6Yc9q7OH/f/Cjk++qtooRAXjyRr5GDRLv2i
ri9sCFwq0GLrj3thLZenkNUGByR8ESMEnbT5Oo1wMmiiHcmv5zzkF/epVsq6
Eg0jJpLwZt6vMZDSuc8b4pCLE0AiWGEbJmTxEXlFiVDo6CUoY90L6ycBfTfM
ZyXOPy58RQAKr09q38gO8K/+jlfAJegXwxv0C7wvB8vYliDv6fgF6eEREzRt
UsXa0FOKKwOYz6/BOdLJwc7PoPt6QM2dSklfLCBaw9/P0+F9lPuK81SmCkBH
wuSx3VKxhWszuBaTwvgNSMWPWIrzJTS/CDZiHz9teSkcuQ1TfG9JWpjnpe/F
kq9Qr2yrzmJ8VtwwGvZo+0yaBbxr5o7YvFWXraaS1oon9l4xPfqH1/Felw/8
k9AC0wdMI7WHxi04vju2SmPcSejue+Q/jc7nvwW8jgbITqW+dfiL9ed42aVg
Tni+GaUhmAvNcBLj7Xopo/cGPlEMaKmCoClObH3h9SFkB8588dWryjQpSV6+
1pCYrqx9Q7BCzcmJ1WwCnIJC7pmLhmhNFVktGtWBEBqHr6GGFSnYngWkfmZt
KMmhPCO37anWljRaHopvjYNFHM5FcA6Z0mCQhOuWmyyquOL4FT0mlaBJesYl
SKFCagRfmiBIZEhmHB1mdE1Qc3YlT6gIDw0XotkcaIUTURGke5xQElJuxd/l
7BHHAgxkW/V+ivN3CV/edlwYOFgu+STZ1v+mGNFVl+z0Icmoql8/9R5GrrXJ
apVsErERcRKiscP13OsUqPKvY6KhgGdnG1Vas036IYevzOMz49md2ORL4f+c
IUK+/Ao4plM9fpP49Jy5YvlmopZtsY5IvPid0Owlebaux3P6T4qOVgGbTGnT
7oO2ZZM37Gv8BaInMwCnWX5GNiFDo3YJacw3GlfuE51uvO9KP0GONWxBvR3A
C9cCvzjufWRBIL/pYtWYMKdFeK5pAWWBtAwt9onsYd9sBGMmxYBvTpO9aMR1
BvCb6NLJXP6g/X8fKcQGiaxgp4DX69ttrHIGgpT3+ERz6Q0kj1sJUsFiI+SA
xrtIg6vMT4GO7N5tMJ2D7lavOAEhgdkaj05R9jD/uIs7K+54YSrEBdEW/UTt
RB45UKWgzHgGvILgF4yBpbz58SVOYZTIwxw3gEPeo1E5D6DwRL/uH00X/He4
wInaTTrRf3fA6FgBj+qwQs8T1/K5BdVjOEPCdCQnsmz6GDD2d5CLRvCzK8NJ
P97vg4AB5o1OUuNJkPUV4bM0MVjnlg5/Q8d/5rI7RxqyPN3saMIRTZtmulS8
6EmMYQ2ED3gKBJEzwouRyN3lZ4dTBKzifoIlKzcGxmNxfuDQUU8RhQPb8Vsm
PGHC5bdNBEGj0tRYp87P51e0Mb1epy2uk5dB8o6phiqPhwRTwgPxGu/SpTd1
yE67vqqJhJ93ZDm6YBbPfIDy4RGVh66cSLm+XutV9teKivk2laDyFHSVJWoU
889l28DyRrjwujD3Xm9NTRlyatlN/KnNz2+4Gwtul0onOqxI21whpzIso6/n
9yDmSx5ZdLIjbGvRTKusCoro4bNbP5D1FJe6u64JiHS1TBlaIbVbo6f8Z2Cg
Y27o7DIPGo5JaWqZmUxtewSWWxLCoZedj2jWiXL3DQtVQWOSVZAVaaqDf3al
WaMAi++R7aP2dAxnkiTSjjO1mf86fAR1E+i18YoHpCdQlrbaKfyO4mDVm7WU
WOGrQmU8FiZFnODzkCSpgRxceywI1e+bAbqRYkJ7kfEmObKTE+hAFEZyK9S1
+UxVz+pp78mWd116iuPCv2GJIGE1oCTLKkH/3gXi4QGqgt/eSgK8JdBA8Hvn
bZud4VnNRtRog8LgJJ6g6EhOs+LFWr6P3aRWN/a0qtWHGkGmmX4HgoQ2Ij7u
BmevKTFGxTnBi6w7ZH3oahH8EO6VtRgw/qjfoa3NNX+7lGP1NxFHth/YtyCC
eBoynoQY08vPQRwODmMahAcfkjXHJZvhw/gFbu/pFZzAwYvN7trm50cTr+f5
7pzGjXS5D24moVqEKpqYPiMVz5Wm1EsSaA4bGOVEXNXNdvAQvTvF2hL5KZaE
FG6XFDxXeuGtt4sS4N1FYyq/ULxEx8QLNPGH8R3sxvlo+IqJ8UABreteIHAq
KYFnNoiTvmHvOAG/aqWt0LCD2tjs4TSsbDs5MiR93znSH90p8jAoX8Nyf4tv
9YxY+S7so2feo0hB/tBNFIp3ophrc6l3jy6Mrc1gejjA7NEA4zR5FUP1iMB1
MsZwDmJ/oF/yXJqUmLel9BCiHevyFpmC8WjbF/KXPFT3432XOJosc6+Snk+z
qZ4yOYXFvh7CqwQ7q1/8aOKV3UsBWoTnInbjAa6QBoCfBohZgXeP3zx1LTic
1Aine+JQL7/cPm65xvisZWTlbUFLS007mCFt3aqE8Qwqu8Y6I/AxJfBnSGx/
xf/iXSuwUj0L70hDF0RHxh4P49th/NUyC8spcxXuWGeYMtKmeuOGg5B3F0Hc
40GMOjRXubWqK0Z+4XEKWKBMoognHAU4hrENx6RQzyK5L+xHQ/EGZU1/AeEy
VjbE8E4cHSfay7THhAiy0CCw8ul2Mz90yHFkBaiM96FZF3fZKyFlUCKi9K3M
ze9PndUII48Vx2Hc0/DyMN5EQQ8MSUo07g/EzlhAJkVvBYfW2KoGuRrbf1nl
ev4zAYYWwyEra5ZsEvDjL9c6I+C9+KYYmX6Ttlv/da7LUcj/BBJP/mYCnOo0
xKT3qf5UX7HA/YpzaDTV7P+iagbzDiiYpKwdUeDazjFvFtHp7RANyjfabXPa
mDQxwkrrhUSr62hsUSUBTl94fnVwvgjjkS9crM7JlC9fC8IaAqt97jADakas
Q5UYHCcmvR2NDalGG0bn4LbqMvGwsjd0SpCjEKxaLVgwng75Cv+wRf8H8D8O
kP7NMsY4JcLz+wat2/rAPixRK1pgvvVFDywwXv0PC9rCGSXtAxCkc3ztHBXr
z4UoxD/MvIv1NlMuozDuYnviGm48IPvyKnKtlRvkPtuXsREVB2WXaooPJK4d
T5jOVp9jqvcENuLuW6tVDwYBAVs9TPn13HsoR6OjXVDSYrkMRn9qsMuXErKP
r9fb58eMh2/7O9LkafEdUA+vikwoVCb41g8fX8w7/h+yVU+rpdDIGYtGXI82
7lp/rQQpM2gciGU5Qgu9sDqmezGUtJjVAU+Q+DauUH9aqwuPi4C/IeDHbPPG
iIsY0bDraH8mmtOrQi0xwRoLwaU+zStTHll+DOQ/sjOoR+xVfcYe4UUHvYik
Mez7NDhTicbZjlFmiIxRhgcdpZ5uiCM2ykuQ4HS/9+tOAZQV+ZJCHmC0xA16
SGljWYaXEzRnasW7W0F60p6pXzuEHvAZjux297Ku9iNL0wfoVCQ1B71QEwCt
xBEebkMEscvyW6pUPWpd7udz0Pjr3m5InveL4Nijs9wr4r0F2CUpi3u+PbtK
vauxgHG8DEYmGxq4mFpYI77IyXlEvGMJQJh+MjboO2HodG2rD8Uz+KVPGfiL
orN8mFCdda110qcpr+4WOqmGkGamHTuE3zyBa3qTROJiYLWETMKCgrqkB07X
8ID9WUKYiUr8prt7qdGTn/6x3ZRHo021q5yjePE3GVjhXy4agRRluuyM6FL2
qTrRBynbumwZlo0jUiSeBQXfLmi7WXnr1STnZY2ugMqL8w2cRdya/ESCaTTI
XMq+0CCDLAwtFbtOH/Brna1YTK0DgYDJ5zXMpShDHc4mi0dJXyTno4aIkE16
LPCxpt4c894jhkQAQEgxBosp415wOWL2D5j6vD0LsJo2ZQKo6acdXEmbcHeT
ytT78/saTJ6+sYiLODFVm/HWbwNhWcKrEoJ8emuk5fnSA1/yVvqVRHI8mG8+
R6wYisxlK3FG7q55Tz5AI6QU/1esAOqy02vMKRpVQiQxL7fpzhiukjmf4RE0
1zPJzJHsluJXYdok+gzaiVSrIVYQvSMbg24xC7wCCqgcAhxWPX6U6HpyhjF0
qnYqNLxkPBN2dFUoUizP540xfqeN5olcDrqTWruQLnaGy+MJN1Y6E7839OQ1
07HTV0ymrK3tdADIc/Nq/9uRbzvbxl7tYtGNj/pxjUZ75ARWN2pobTnDf5RV
koCVnKoXzl0t/NliL1EIutktEYCfwGr3WC6MQ/MzOydW5uTLGIYZAr4yCTFp
bv09gadef+nxOr2AwnIBorQv2Rj9n0JQEonAFkL6VXjvR5pOYIOv7zv8AjQt
ItxTfHXwoKD/4t0vDbcDnQr0dE5/Ey1BQSmo67FUwzFC+y5BSRhMD3kAWBl7
KIrOPK4tfBhtug0xGHib2B9PlnkkYPyN518YixpVqDf3XDg9wH3Qj5pm89f9
iwU/QaFKMMT915ZQCT/ETHomTWbtY1BvN/L0XWwLuffxWAzSQ+7mAn5RQ/kx
kPt5MIvEwvLnyCPhiaxkJgxllyJYz8ICekA5/kCUzHXDoVhmtTj9hAFKo8cu
SfDwrC5VMpYc60Cn4fNVrQC2P261NmMjkxZVAW+wN3ggJdFZRJooLtF0NP9E
hjWUF6FTNQUgJHGRhY7rZ3YOAxUy36Mm9nDDAHGiUFi9e9gfU4mhpQAfbJxL
2WEOxYHAWiJ5kUwUVxgOYAWl5SFD/iSq3OD1SW014pbQBfcLYIE569SQ52Yj
jSLz0MvYuJAcynoompX0zppA8m1pJbBC/6O8Giw/+z3sXlWVJN8uA0WY7ydW
z4qXrjNJXJBwTbsJFpgOVniuk5fKDIGXSMLJHQ8pv/Ih+7283nU7S55GL1sb
lksekeWVPlcx2/xfKFO4AtmdJgttxINB4xoOSHoKmCA71ewCSolIb7OPJXLJ
mqL1iRK78gyeGq14J6Hsg8q/5ZHQ27lkbwR8Dkh53h44ijnHHj+igV5o+ZX1
0S66PiSvgU5sOpBWWuJLh+6SNwt9WpfDS39QMRWnUDqpOZ/HZJkgWZgvyU9j
yFcGcBI11Tw2Bl4PFaoWeOOLMw5ArhhL5kxmnfDLg7Jri3HgYSREkwIhOSJB
TmoHz0BJlOXLCzKUMtgYpi5cUiZrlaxBD1w4sZVNN6mbPdVZ4bT0G+op6Gxs
fWcsZnvmYsTaYnqfWMgf5nXBOcBPC2Q8r51ECNfwVGqsfB6Vgmce0s4TgVQl
gvKPn5mgI6V6I7ErdIiFfFgPaUhVy5CdxDLM5j4rGUEcRtTe2+Sj7vpUSRhk
xhur2pyd4i39aihj+/TxJsEwCD0fJPhogiKBx9LUMIHz3Un/SDADDrU9Tqke
e2M/98Xhwyx3mvIBEaFwXnu5jJO4EOKv3ZuFcHJQQW9Nt5LPS4JgUwZUydG5
mYInTkavEJ42V5eP8AARURm5lgkzqHsavRUIDBejXleg5PPSph+Wnsr2ai4P
pftL2jz2yjgOnd1QHrUJEAJY9pk3jlR85QYlTzz0D0DtS9cE9s8/TiC2iA7l
ywvE/j/g/DEJUiay2jaG2/sLqUETXBoR92FbP6kPUJCBdUCxJvpvpYcrzsNZ
m/dTIJfQDHI2CSa59Yxg0KS0mdE7ksBxFdXrKT2fD4TJA26cfUg071AyorAb
uDNNZz6HCyMcstwmY84MLT8UZpQPqTph3BewZ9HH7l6DgM1PxKhCQAd8MVCQ
HuGbqfN3uSJM9xxb20jUXl2RVY2yd5Ua23FAr4cr7bQOyJA6V9+BQdJ26mpb
h5Ao0Zha35UKBb9y3PKYYt/OEEnAm0or+9Z9tGBWeDmEpqLYhKmLMUZP3HOj
UZ3wRPEjQ8C0GcHD7PEfffiKDX4A2IzajVEJLfTRe20g3plF27h3XSSEJyy9
DF8GixcAreMFSTv32ev+x5Ud+riLyovgxR2ed/tDdHR5a8J8oQbRhRMVts6n
Y0yNORRRIxVBEplJf0V16eW5P7ToOkqrrgsUf+DM1odqPCG8VWoLGLM7H4wh
oGH0LSjqZPvr5SUX7VOZZURxz3Bghm54jDK3GFzKuGlHnDxsTlVACFloK2PH
KV9z6zqun5JIXWl5ypdYbADcZtwhUSJr9H4hNH8gPAm3Ou5XY6xuXmuec0ZW
FYRUgBMdKufu/2rRPY7LBX5MLMdCMyp3hqLZDi5wPOXFn30icFT314U3yMqj
SAH+04X6eU2qH6QJNzPhrczkT1wGmwOB+NHuQCcQX01547gg/4Agfc4iLbXv
kxnEDgA7vTHKIDHPHMdadQP3fctl9ZafF2k9P3k725SpWZRHa4Az0SBvG/vT
vnpvTlRI+bmN5Ywk33t+9vpIcNcd19IP9V4LKijeL6Ol7+/yo90eOkVlulUF
0PbtDdQnWLNeAtKb62lIuTdX1xcBDjbgDn3oFhrN9D8qjwEd+Dzk8GeS32N9
CwIII96HviV0YjRLCNysZ0gtFsD8XDtxR6YQJlvU5IZEab1N9BDhCJpJUjRd
G1IJ1EJQ+Ci1nY7GBRRKT+C/yJXucb/z4VkHx6yNjJ1WyEWUo1k1hneoRkgS
DvlRyKBSX0whVQxIt5dI186GGzjpv/+gm7EA1EOBkHwXUj69+Ht/UETQAM5F
s9IOdPOEL1AvUTZfki0JALVrNpCWkvghqwKeUP1i7p3FkK2mawsEIUCIuJMU
fxyvNutAuwMZxacusW3I+qNJz9i1fdgHRKi0hVmuCvpZOzvi79uj/RTtKPPy
POgXWy7wvdGMLpoGFC5BtLQiEMlvwL801O5U2p6TZhpBJYOuEU9GTy7MSz18
tI95HHLzYZxJavjne7cRSVTwNe7hJpIAf+/a8Hlpe327oYF11je84vN+e04l
N7PBF+z4znOhFBJ89BzcGlP2WPTuuyiI9BF3CzD2gNkergT678/RDiUP9DZp
lDqlUbDLWC1emeeMOf2BUzdgIumJWXZ7xS9hr4XzDhvlBcxlBRwVIXUtKLvp
f1Rw5WlrZY6Qwg3f24gb4xnuWtUDYizQmo6miMv0T898ugDspzYPSD0FF7QA
TwQTNCC9pUnitMJkKlNC4BPlfzBIeBCpjJ284ZVwABgsDCr/uFsboIqX+YaZ
X/9NHMo/lNPnDDwJChXrxL38J4OL3/HdytbCFwO17UjiypqaswAsi/xyXOxM
7Woc5ioeDh3OUNmdqqAeOFNRQlwRZ43pRDwfG0rlwayNNp9AfeCEdZp3ZLix
zHq+gX7X6jtH5GjZo0C8QYM6TSHAh1qfF70fZu3ISEMVHpkavDXogW0WXGL9
mwVmSvOXA7kqm8UAPZLAxxBb3vMD2F4/fLxCn3tFdmi0zlGb6V18IPu5btbK
PQlyL8rH0A90C9nzEZzp47IwZq3jTJrZ0IzJIsvSJ3AsCMmLO/WgV5kHbF3/
tSpMQeSegqWwFfA1Jpvg83OU4ZKaFbUb7ft9ZiDm0HGK8zJoLZNGDhelbdun
FrBV5/fhYkToYYpTyaaKyF/fvTNZnVG+gOBPrGSA3gWXQRJaaTsI8oadvRho
1QjEFqf1Ck41Zc36o/cBDHS4lzh/J/Rh06FExmx/VP157T+wR+QqdhoUdQ4j
Yiq8kHQAYY58RqoXoEk4JfchofDXitKItmv4xQjnDrvcWlg7zcbXZBkygdzS
y6WqTDYy5AZ5e/XbzgXy4jibDn1SKddR3YDp7C419HVNEElRRLwygNWB1xbE
UTSnFmZ2/LqWvL55uU5EFXtbVgH0tjNS8EF0Wrk50ym9uSZBfeQWhLvklkf+
J9TnNfdEEee88+vNWW9PnNoktM4Oe0D3kziw5o398GLjas8B6em39A4KrgK0
lCR1E5MuuA1GyE/277LWFQ0j0bnF9zvMNPfF9PtU8JmmmYmAUaQt7KDYxvA8
rb+OJ0rQ9VC5zKnJD6znlm7jyN9FpU/VNLbpK4sVCrqBS7o+Q1/WT2GvV09M
nfjk21owm/Zp1DiP3Yo9IFD6Jiqe9MiqsLBKEPsV/7ekfGfQ08hLLBqLxaeS
5jUT5/tliAu19zUsly3e3v/g6+MNM5zF9FkFCbyf0IEy/3V3sfaNFUI8RmGc
K+h0eafD8De2YnEZ+CWFzmeUR3gzxdTf7/9kshhtooBCoi+Hrblyv3gKLCpM
ONAc0/o54svWJChHDD5p5d6pbCkGBr9TP4LuK64hNS52U87zuHZWpcvYJ21F
C7HgwV99pxIJC4AtGCNWc1sppublM9HqU4Iz7oA2OAKkVWmIVpYEiSs7frUh
BD5gi8O9BDrq3fizn6gw1qQ040TnAeuB7Ogph+Sgp2SZ0CpRDiuf8ytQnWzI
GTUqemVRxVhGlnu9ivkf+udUGer8fpoC4TLbkqv5ODH81XUHG8jBXwmGtSId
dtSpuhhjvi3MUpUPdXNVEU0xvnUfrGgyT/i0iIAJcw65GikpvQWPdSbkiYBo
9mOhuJukXndPOw4ljThfz932SO3hFdKTcyvdgGPlghm/gxwcxlH9+mKuFYbm
NkMHY8h01fuy9KkoaNJpUSV9nwBiYLEic2Efy5aoHL9qAFl7d3jRF11SAaL+
APSDTpfIM2fv6ml+TDVP9VrGNgpzjbZnlBc2PZ2axFyZ3i6rwpMoAkMKabpU
VhP50AWK7hPr/7+IzOu/F1t8UTmyePUB4PyD0CdWTMaQC4Mo/9BaT+oxXuGK
J4lMgp1L/BTJOc67hDIu0dmSyW2xe4lso4DSosIg9hd4Yqvg7mMHruTM8M7c
uVS+W5rY8fMHqfqnN0VDEhh4O6ZYqI4vSjMCyiCD7GCMJjXNcgKk20WQ16ff
NRchsGwOWChz1iZnNXdPL6mDhek9bTOHljtcy52e7CJ+YPMIXPcSvQqlngEf
6bpdjk03exLG5eSBJS74anY6vb/yJoXD+N7zoEAUWzVPsFZqqVyoB3LCCvEw
e9CxVUJLez4L+q3wCTsnmoJHweF6CoxuR+vJrxOPzts7MBZPuEtZIAc5pUWu
rXQHwYqNLq19uaaUwlhI9jz84DqWdKnjkkWbjQc3wRnZHPEevaeT496811l4
8aTNjgDR6hvabUTZZ/m9CkfFsc0G4GuHjvEsuEU3zG29oIo5GACM6gQWDvvz
Jp5nNUO7JA6peXkNP4WArk1LMP6ypB5v83hEqYZ1meMq36W12ci00Q/eCux/
2M+0qVwFEMB+CFHgIS4x1UGaV69nzxqmiQksWyIX7dwp+hMSXaSPQbzBxAEd
8b+bE1hOl/dFEoN/M7TrUI3ZXRmnuYcUiebTYSq76Q4muaxiVgdv+m8qjSWQ
mtU5DvacBXUXYISs2JCqrVIg6Gp6dEgYmqzCc3Dm3l7JWgeQtuPUqkwtIeG5
fypmn82c8R/d/yANuSzdd6vtKppP2wO5eOvrwp0zTbUyx0awsMMZlV6wywpr
wO1CQWfUDNYphHDWeSkbZyG+MWHMEnfZm8hFWTnPw/MPruW/N7m7lGhQ+BSw
DpusD5BBajKG76BRuYYt8e/ZoZwNcqBB0RPbO1oj0YGMyeTCw0s+LWjo9Pk6
kjbJPJgQ9evSYosP4X06jae/zgC7Oel+OvRzpM888McKLWYY40gT6P7AeM8Y
ex0NQEUWTdmHIpcyrbu144ir841gc3KQ3KayxZn/kcMRnaT66Pn84xfnzRIC
l5nT3ZZMUKyoO8kl40t24l85OWJZq+rfhZDWepVL15WO0E5L6jKmE8/zsucW
gbvGtAGFE1bXxMmVj2lmGDF3lM4Igf2t91HgM6k0BaOqCXru21FHjxrFtes7
H7WQGLNMpauEGS2LGE0UGuLrfRUXBsA8iN/qRG6q9u4W0LP2d/BI4guGhfpm
WpAvhPOAgyFK1gU9m5TxSYiIjaKP50scsC6ctGThql6FyQWF6RCFSCT6J1rt
UToOpU69hIlbV21j/pnu1SIBdUoeHuGOpzn+cMEcTe3NrvYy37I1LCO5CiKN
f/JwA5rR3XFdIMFS6IEJPaIRD4fGO+ExdORhxuG3W/ib4s4IKVG0QxVipZ7S
bbKgGQzC1EtJP6nxfggKUuymaLNRP5S17qzDblNPbFf3z4yqa04imy9ndPet
W4RI/rh3GjG4ezYSowqygYvxYKCjeXu0eOK58nMNtVHV/rwt/Fhrre+7bObR
bIu8H8Lc0lqBYNW4BCjiKDN2rPRiRgvWigg4LP4kF8Qde6TdCbhmosUlvF7+
Z958kes2TRiTa+5RjUhiJoYLXFoJ7r1rasnOpSxNd35LWgeEidJk1vWniSBQ
gAiSiWe5nWLoPt8flR27INmUDzOMLsytoAGAO10h3g8+Y79diRDLqAgVXRpe
w+vltFpGBYwuFnHwMIZKFLVMr70KDhS0zgg2gK1mj1tDBNZVnqBOt7tlaa0L
7DXECQOI8dZEhYUz65vZ/gc8AOcHijJhEOWgiEKtofUZN741xRZ+q3V73qoC
FeIyC/IVmjwV908BYDYqi2zDfeOdLNUC5eaDkO0MYCYx3jo8L8sk1FFM+2C6
pGqSPZT+8gwUZLvh0P4w8mthJlNf2XZ4W6q7YmYQzSlKiNXDTHbe6j4TQl2D
kUNSlNx2tW5WQMdhUKYfd+G/aZp6TZYaP2THn12VP7mDg2cUfcKbaGLK/inG
sGif9N5dTcKjuwLURaVYBoL8uHsvTg9/Gy66gXoM8qTZe96NZFeA2Cy84L6U
Ixczu5rBCviaGK8AWHh7TP3AEvYTxwpkspFHFsvhBJNq7y4u/StCY27iHWHk
aUG8fyIuETeyyLyTAx4AlHhvbVux9up6n0+roeRqnsDWgBBeS6Us/Pkhohv5
fozAX2g9ZQljOB3WMbn85JK4wmPGM4lNArWVJsbzTW3wFwTRTpNUTVX47PxZ
Q5vF8t4zVeHLKFeADUxv58tD5RE9T/hmhe+X3J0ipD9TbuZaDtsPWwU3864b
QdCI/u7YwcWSIqpAWH6A77/Y8UQ9cTUQAomYWQaHQe6gAzw1CW1wy9JD/CX4
EqpSlBUR4jLQ5QunGtY9hPanlgsEuTLz5At3jIxPd1n1oOvhCtXFohXoV2zm
VFxk+UIsoPWuH2VWGQ1wDa/HtoOg3++VJ/XBX3gqLtBOiF6HK9SuX/51qoDo
07wFZB0CNngLF7ESAPeMeMKGPEepwVBReElpySYDqyI4HSoXKNu5sxMvZAqS
dkE7fEc8KNLLoBJ2lqRPS8IMSg0Dg3nmULvyKxDDu89U8g8oPl9ROxIID0AF
iUmDcqI3407GCxQ5kedrGMoQt3UoOjznn8J6HL3X0oiXjmAPCWV58ju7D1ZS
ToJUvVBo0+Wv1SVYnFnXLGNlTxPIzVdGPk4CWmrZehegsfqn1bTuQcRArPV2
IMDf+dNZDC26zbj00sQXl93O0lNDcqmi0np7RI4zdN8V0guuwbeNGG1DTZf5
hLyModz7LvGNAA6/5lOz2EcngSx0g/sgBkQEdAJPrk62+ONo2bDnDRc6mmxy
qizovDZZ+iqIK+RcsIzWIa7+ia26P/ZlnGyPpgW1fiB9LlDq01tD/xqWu30x
1KZ5pKbQeVmaSzfRTU3e1xjRo4nowzxYCv6FQATmPlAY9G3S8Qn1VPTI496w
S7N6vaa2eZ2PZPMhYTLhgahqp/ldLjXC14qT4G28fJlN/ARDVelbbkMso3Lw
M46tlFXTrWfcUQiScXo/STbix6kCkMVqB/f1wKmg8tkpZDsHtTGg/6MdDU4R
K0jg9sIwdf0kwBBL3cq4zuUfFfx2QtrnJERu4LMHzc+MPSgLu71QAFsXyvsW
L4WTN4ad02OvyvnBGrE9HWEMhIjyBumLBZ+zVhWzYKorOLS6SCP7LRk7wp/y
+GDCDc9eLjwS2RZ1yXCdeSb3N4hjbWZAzTL23Ux2mQT8qfBZuFGl8NmAc9Ic
vJmKGYLosu4t6zmRbZhPxdnIYaJUBupUXF90WZPk3clI5Vwz3/cDJOZKfIxz
wgQr9nmrHIFab17diqcauvDEq2lctTcztRvwOkaufQzp4sD6GYR8FyODFiZG
fZBZIrfbB/Py4ZPn0fX/ZSvuLWhSFfoek/VeQBddY+L/Lh556utEEqVmd4lV
JXQvbDfuXB5O/ykmKru1v91uIVzwZcazBbUtsAACORxpsaZnfIH9C7t6KOe7
E0nf3eiIzV+AYnSTFnnUtngBrXoDTR31ae/OQ9wIprKxGev74goU4Xir9kh+
39zLEIl31r2aPsSxe/4vtTqjOSWgBJ6tlQnmnPaxljWQTa3J5O5tymNCf4GY
cACyLvaCq+PHmRQ4/xbA95vavNbNuewwcIqUlxOkvQme/BlJdPSJAxVY+7wi
e9hcsm3qxPUz4gH7GUF1nTVg421gph/ZsXpgRia0ITJSgU3HJ3giTy9VtNFp
aIB83w7pssGgk2rxHdD9WoG/HuI7uJPAYgmE+DNbhnoAaPgPycGvVSOv8Pcm
j+xfNgPILZ9oBFrqwbkJG41pRKeDJ81et1qz/efj3g9q2wH6EpfOJudK8KBC
IoLTdLnuC/Z9J3z26E9gEbCuFfiEA56RO5Jy53He7moSXniE87nk7gvaVg7L
g5uTmHMRTpMMBkvm86jAJWVp6rMPjHPKQLqNjRXuHPgoH2PDS7KC8NgT6CoX
KM8+vGxJYToKlMfboY3EXQ1STN244IzOTCXkvfLqp1ucPARCGI65yKLH6jPx
q8RlH10OqzmelC/G3VZkQGII8p78OlINXBQnMrzJd22I57EpvbfoJF7C6SFq
UGxjXbNXF1xpUagcdZSoEf1TUmF8R36AwZTfZ1u50IjqKdQ0fgbSU4ow3+kk
uxREANribQiMynjgpxSLXbxaly2VlAAxr1MHpGqz4DXbfiajLKKdNvAFjukg
YGmm6ExxW2RliAiJ/7RlVhlefFSpgeBapU7Pm7omdkMlI4qyWyPrRS8nYj0X
FeYGioxeXhXfAH+CTifpUKvYfvz2DuY1gzJdnSfBypxtw1aSSBOjmcNA8mXU
wj4ax20lm0qUn9SvVmESrZVCrb1uZukIsfkQEJmk0e0YGaTjtSlck9Mqg95G
4l7HI43MH3vJ6SqZLTKkbgyZ6BsxBF6gmQHND9rryfcMcuI2ZnY9Qmj/ax00
DVtuFP+bxXBsDtdK5XJKIh4tedFisqDJ/LwIkFH12whneXXm27Ce+DxKZVrS
IQ927oYUw1A+z3nn6Fhohz4GJMaJCQLOogeiHI9HaQDjPbxsVFlR8gXNQtmK
14BktUtqW4DiLw1xPe8MFGSImPnXynSjeA5sZyycUIdBgpBzJ7KY3LtZe36h
Dc3rbX/RWwjxOQh76iNmOdEcXqQhTzotUrgFATHwXVBeWUP7kAegygnIum+E
wPzG1X7n82QQkBs61h/wxbcmhxIdi/sXayLN6q6MEQfJ6PKznwOj1R5jifxL
E8o5Ed12Aol0Le2q0e4zxOaZgVfWyMUzDGRA/R6ST8TI2eleSn0l6o8GYc8m
3CAV2rkzhpxZG/02Omfie0ANoot8VTLu05Ych3mUBKmsRUEEBu2xUVxHNyRo
QQIYwhoYvg5vr/6ANToZQMNEVYku/X8VyTUrSyADE7NbZyCangBZqhJ+JTJi
y+zZPkucGlI0vSfx0E4FV3ztFPYkzvW4nRD6Cp6aT8FrdJNhSGsQSYwP/Cct
TkcqbR4ZfEhUWAg14xbIYQd3im/F73hHIrB4PEGtIp9BJuo04M+oyWOkjZVb
FF0oTd4ar27Auk+VTdivel5OpHkkPn6QCW+fFManh7FCRgoCNJ5UxMNqF/eO
ryM5rlMdQG3WgfOSKSpiYK7MXBzKufUKEsf11CUzH3YSzAZjyiRGwKvvovFi
QMOE9Z7I3vsArEB+RGgoFf+kqqavACi1xQExU3GE4yIqRVmVq3sRVPnHfe3p
rG9dt1P6FVPh23vFmjvfDWFnffRl3cFBzxoJKT7YHFTTW9YGPATG7seko+av
VoFFIDhOSMAN09FLTbchDZDGy5kFQIdG3Fm8DlXPzAUn9nThD1TsT6MCZfd3
3Y3IHqagxK0crYe07lTKdY5Y7Eqol8e4KXHqp7EBSMe65yerBLTqug/uMu0w
Q+eIP0ZmkTQ2ZLYCH0gtQlnMk+c61pmTTn2XQeik+NnJU5Uey3n3lcOOYXAX
jresdYd18HrU3T7GES2i0Pb2DncnMrO+oNNcLTgNUvAe8LXV6bJhIlRHeX4O
1UHZOL5MmNO++nM56u6PUtuCS21VMTij7k7TStkUZCROoy786/DX4A/A9cDZ
+3YAaaofWEHQL1dRR741MotZfT9UGjVUgpmRF05Td+Mv+U3MvAQv84ssAiRD
h2+SN3AfW1HGaLs+mKOqCyg1KmDk5YXUw6jdXrM6wbbzJqOLn6jDrIT6WDUo
fhtDmkzgR4MfGh/jUnua+nlLJfLtkmwTPKRwCETEv1VFXfbF36UjClDjixz1
kkL5T5PGnpyTP/KBdgoNOb1I1GCLPTyOTV6oGrsIQJ66k8kHxmFNjziHNLo/
HlyhtVzCrjzRNgD8FIK/ziqDPUqRZoZMvlgJjtben79xoOe91tDKQ9QAMTP9
NLK5eCVhh/7E9r6/ICZPntovdU9brDM459oS3MN37GUB+y0z++qe4QXpB9DF
76wawqu72g4kes282Jfwtuy2ZgclWaa7f07JCRaIPsoAH0zic9ukvfhMgQBU
4wjtmzSMHywQ5NBH4VkWymOHIXzcmnVGhlxPg0m6tpXnAOi7OvLCbTVPq4NL
NJ2AtvNIofzIKUMCfQIklUJLs1wmgNAz0XxgrzKl/Drrmcwft1iLq+g5KA46
BPsjvU5V7WOM8ieA3hRBEuUzgeOkcH3jo8ujJD1V926OCT7DxKl+x5cIKF7e
5Bc3BiX3RPYS1EVF3Lpt63kOyDyl7/QBy4t/vdCoAdrZ+9rG3OssgKQVWTxY
BlpFD9ee1Jnic3WbrMu9xQSYjUsuzUjxy06irHO9fULYD8d6VCFbMubRdIBL
NvWK0ZIhGm2vsTgo8X0RqGwt4DXov38xATCI6TYISld8i5w/2aYhQ+Ff+gA3
FPtvQKo5FQt6ZGXmhpfilBwgxdw00ZjQodgjag4nOdXQbgv2Ic75p4XQCZSJ
ee/cUheb0eAg+k8I0+01VbIfKP97rlv9cpNt0Iu7Ww/kSnpma/N171jxZ1fa
4sqp5UJQAyU0v/ybAPYtlG9tTSf/mo9lQxVdfr7qjzK0a9dLkJ1loRDfPUrP
TcvMJs3wQH+XvjCzrDBg+E3Sz1MQZPzwPi07EtI/i8Xu5SebIMN2xhDFudmT
FPNNg152wL1B3IejCxwwa/v2oSEdSueYnz6WMtL9e4+ryciOK8sCLMnCldcy
olE6m0UTYw1UM7u+Vat6S8kMBgvgIa+c1T5b6YUzH/z0gMEQVIo8wIkonprn
h3dnDlwe+ALmksoULKy252pyC4BKty4Q6eil0cWvaZm66cR89aX1iCxSxAtI
ioPyrrwBkHa3ukWqBakQpe4G9YYlAlpexs2/0IZza8G/G+Zxea3snFIG03ml
jVGr3PEcrqIgE3T39UbPvObpG53WNevoM+ZspJixtGF2jIibeqvSg1FlNpVx
5M38UXdBcZ0pnXGYca5UREem90KdJVScReUKoHJ/ohRfBLUkBAKwkI+KZaww
4/UKV00TwMgQLwr1nc7s1iEk3ywPiiG+LvRo8YoeQoYvKbpy+aloydGRL2J3
JD39vpD8nG/pcNBQnqeTJhw1kx475AQzqeafT2eeUP2MGB49VuMEiDmpHXAd
LtEIL5HEl0GtmtxCkNOgd0rEOfReiNYSji094BJdIxlHu3ENndEC229vTOPy
pNrLISbO/iC6Tf7BWCJ3YQcwk7237SWrt/FaxaMdg5PSyd9Om6WBHix6qCnI
eJytIQ94GiBN3Jv2uZWZNdtb2MbzCK8PdvCSKqD0TXSbpdZwCHF/dkiG1dzj
8/5/jO0MKgPLDwoavuIq9WtaH4Dt8msr7YZqv3PPeeO5Bl38SWyBKnjZfk0D
ysqQpIhRPjzfmVxfHUf/72Rnjw1ABLx2AuMJuXFghSLPxpv0ANZiFeHGFDmL
ttzS4hpOh1pgYGde5G3x6Dd51yq+JCZP7Jr5AZc9gshJDRdSuMLZMwikhpWM
KKPWu2cWR1GOsg21ZjI5k3EXaSF01UaaS7+5cuqQLtj6h+TmTXFTEIaDSo0q
s6uuAhuDCVLeRTq2Jz9uRBByqqmgB0U1Qzyt/f95uDpbo891f4iE0O1lhOLk
tEKyMTOv5yBJmiCLU0GevUtuAKZgXaGwezKr5OkrmBEgyMNutGoled/lf8Gb
jAkg1yPCelLj+tKFgyid9QuMRPBR/bYMrM11HLkqRg7DYaFttAW/vJP6bu1A
zLPUW5bH72J635UTx+8A/pkgC5mnAvQj0rEHtjtvufqIt1AyqiqPioICCbom
RlhXwhYyj/scVU94dSDlYI7PAUuYTJ5pHM5jM+K4bRRFrM20XgOF+7QolaBs
BUQc8OJmxYce85sKIuMdRQBtouUpjjSyBpK4i6AbopyS1wk1BGgqUsf34O5q
GhM6mhteuPjyaxlC7tF+LTPmoLfhfOZLJCOKiIbaOdVL/u3lU5e+HQ+9ZtGs
Fi+/YkIKuJpfX0xXub4w97tWo6UPXZpVOOaFrwjVcJ9uFQzXNVXo3T5rDM8X
2aNATSDBqy0jBE71ePVJYQ4wLLry9cKdqKMJEbPESaDFW/e+Q+jGqF1ZYz+2
bXClwnY76wrdIBUdZbb4pTAnZ3Tz1PGriXlIcfsxf0aKWBMzdK6RIneits7b
V2iwIHYlZOyTyDJvR2LhtnPyqzLU9M9/3ss8YLPTW+UCBtWmAS6z1ll8KhqR
IE3M5EyoUSbTSm3rWr2IiU8gTsr5clXhQbq57up0mIknrizeG/afOlgw3eg7
7kAnHqQLAd0KOBnpFGGPhN8AL42CvCFiHVTOLxynOPi6mZeEtvpKOt8e9Yuv
k14iQNoiaKiAL6+DvX6KNjmjLb+TBEPUFN6cb8Fu0Lh4wWzTlqFlcHyYn9F7
F4MhJ+pEGP6Nn48IHLIwH8QfKqAE3x6f0M4OlwID9U9wrn+chaCUw/K9FGxx
OqZPcySZgyno4H4iOEuvAd4qP7LQG6eKgXqPfSa7oG1M7+f0POhppc++NE5J
FA8Pj+1ZYR7EwnS9wqPu2uYw8N7MQIyyITHjjnBL7hdauM48TO/xUEHIYM5k
dpPThIBWoSVcGC7OSqC1ACAnOBRRv58jowysEq70IysR6isdMim9B36N0mE9
Z9D/QdqgOlyMfDek+OMirb/1+QN5SWHjzjyYnSkQ0ITEjxAztKbT9rFv3ay4
GzSMNY/zhAJoyY8siWXwthdD19VMR7RBPeNfX1T75ifOy4aWj91aCwr965U6
Eoj05iteFCoE0w8/PwhrTr7CePytoxUVVK/aNpQV3JaMHrGN2HAg7UEUy9GF
3rHBI/YsLUafMnFxYAiS2R8X9uycRxat+zPEsI2+y+m4rSXqHD9Q3jWDcGPr
Zp5TqbG+xHIsbIdRaYTer0Q4sRCGwbR6N0mY4HF+WDIKqfkg2ruEIgmOCp6x
p4kjK4onbu32VkJ5SaKLtcNG4cyV0RH3sDAtQvobvrb0OhTEFbAAvpW/kcWL
nD1rzTDmu1qEPnxHTAFnKuV6uXtqeKv4ggVJEr69CeFBlg/glmOt13L8IMMY
x5JpLiH9E7htPYOFI0hgolLwpKM6xglVOfPSqBDD2gkCSYtQnlh4gUQ6SCC+
HggXT+clSqoAn4KRN0m+vdMEbfnNQIrSl+oW/6PKSsK+B9ZrgqtslRfof4fQ
dmeOMhsWQX1D81c3zzpD88z6JaTZMYnM9rDwILtuSaUL7aTtBk0vi1kq2aSN
UEdezpjeWV80c4dCEMwsOPnemBC2MZHSJDfwONiKnS2Le4iCBgz9t2HpTELU
x2kgqSN9pD+/RaOWACb8Fg/+wzKys5q5JUeqDsCGw9ta5Ox+ychRXdkeP7Wn
PmukDLXD/qWuxM0jqKfnUwGMj0FM7/agVRAngapHuwNOm1rDBu21d51R7ZWv
tSEkZpwS0XcLUr0I0ItVRPaHGrBBPNYAFcqi9w9s09svB9fbSBT633h6xXFb
oIYNgdeNDWDIPyebDbD74gsqCo024SllBJyGq2ECzS50Xv6cKZ0RS9d6df+G
P3i4oByQE7iY1RbZQnTx+mfqUrbD80dRW9ztkYnSVyaCgGlv72na1ya08Lt4
3FHiTOdszweB8fmFfcwUhmXRew43N+AACiHd8aWiF7NF6gRBz2i5dKd/WzZ8
u3WrZUv+tzM9zwlxM3y8JmJLwBw4fJDnrtGpME1FsRA/wBAM1mN1G6nSm5dM
X6Ey16HeE75VVYEiix9WVGOLEC4BuGfWKEsbgu0dsnaYU4dkgwHjn52nRDnH
ifbH8wR2Fa57uVCC+LoMZpoUkJ33q+zIvMTwLAmXV4gfn4L+SB3OvoH4igJh
whaRwNJJAlI1uZthGk9/VTx/xWI6qLT3MJcAeurPJFVm9NW6BnjwfPaNbIir
lNLl9w9iGtCbAfzV8yG2YSTJ2S1NR0vwIEdzFtWaOAW5GKrAUJmAFFuR1SXV
170hsY3YBd/+KhwjxsuUP0fJtUJ3SSRc2Z6xmdYRfuFpE5dJtERhZ7P0rK/u
nYSycfeBtWtGqpejc9lvAYuy+MOraT87t2cmuuKCEIp5MfNZtOdCg0NrExTQ
4Z8vu6DhoF+S3iP1KC/u/JIOvuh5iz2lGf5y/06YpYd2hgY6WCWynd4yBw+s
kM/WhC2yE5qD5lKvlhTZcg/qXpJffhktm40Kfzh1WLiCuG0caHTHEiueNMQx
J9SPcxqz58hsKpK11pKAKNiuVXQr4dkmT6TZ2pnvA9M7wOsUQhM0l1X0z92Z
dZKdynfccQ2eivkMrI90I7OcPALI03pkdgS6OGdKbeabtKGQm0VU07PKlCx2
jLmvgInqhDWjDf1gSVS7s+uSVDlV+N2dWpzTPFnxZ7+J+JtOP5h5auq2FIrB
wG5zZAESzVU/nVkypY0eGBi9rfk0whX4w30ELl98MSNYqnzcj9CwCDFoLP0T
xMF4r7GVRxq2TPfhVYoaU+8+Ap1AkAvXCdBj1KPgeXHVnO9wit1D6Xu2iZbI
TCJfyAF/SW2Aem95xylLFgjGs4LolSo3DU7NjmGl+67WMdZKiLiD3JLRzlVO
Xed2LXfADKlXrZr6K0lRwt92qIq0Ij2OI8+RcL1SbGZsOEPhyNo/kmhU8Tja
84Vtlmz1uUEU4LmHfjPjVOpKGykwmNDZcIMKPzKcWsFz05zgxuuXNuiJ/Cfe
AYcGrP4YuA9utcELfEK7wXLkOtpCNuZq1l5LmBCBuJ0KTmp+PgoC/rhzj643
Y/fvYAIovv/xuc6giEzrhuZt5PY2IFvUTIPOfPjkapLkgY/q5BJdTEe7Ve++
sotCW8N/Vh1Kj+IFLXWOzzotCJ15ZgRB42pd0ohnab99tQ4BKq37Vq3SNtZS
UwKRiHTp1s4lny0i3SnM6T15nUKiGKXFvlKHaGkd9XMEQXpU2G7pIM7bhlBY
Uszfrn+sXKEgwfQq04mwHQdUT3eGTemZpAdk6jZOip3amSzpSKr7SsGT9wSm
lp9wbJDLl0ZLwXX9fAtrTAazGe4ugq088akV5BDGtVobgAu14deyx0/9Stc7
8HO+OVrVL+fimV2uFnMqSdVx7+gQ2+dj+a0TXHcOPEgAO9qHDRPeBgBrCfYy
duGeR+tKVeqp3MFzcf91vLMR6JgC5Kp4XnqfRE/hoN2pZXefJyubUyNB6c6f
jm0Bc6VG4VjNBg6AGgighL9Zo5S8tkISvDw+poT0SmUJD0jGQR6p21G8/KyN
xjiNC5RlqkTEMc5U/O1uBtTHg8KcXNFZ/69tBtTAL1u8PZeYtEpXk7PXaZsU
SlZg3x1KXoC/oP/WdeWWvWJqd8p2bNx6EdqMM1ZRNztKXc1hX4f7cuXuQp5u
pYhze84zczRtL+k4zJUdwzYmHr0jJEvymhpwkW1VllvGMp5PM3opHchMAhVE
kU7e5av4wmbv+4VjKUVJUTQgd9N7UcF5TipQpII+12rTpQAKIYRnvHZSVLNm
DkgNr/W0pF41nLBFNfIpWqH+yTsIIAEIXrechCAmcqzerZYM98rouYd0fhkk
R2CbYT49Vw17be+LldvlBUd90BoMOwVsNWAsBFGSIJkEGZFSGjkFEaQHF8eV
Zpg+uMIONF1AWhjvm6wpWRTFiz4N4PEX2xlgYBLDp6zhMWlEDUyWi9zOVt5e
5RYZW941UPyIoMsy3mFWmgJwHC47XtO0KUhuLMlQgxVEcelBHfEW4Wk29c9e
Zn6n+Iy154rLoM4saPxZHgdcGE9OWer3uKiWssEAIQ8WZEcVB5OiIserDUL3
pFj8cJdqKrD95vBeZc0AQQInY9QHa7z28EwdtR+KFK9jMOjmwO9lMDJxSE1m
TGnO2Vsk+opQEAEBHLIJB9IvpU/48fh662mxopRstd7E6nhRvzSsYTJNfqvY
3ZvHVmhQ3w7mQoHkm0XKncMcqOzAvhin23S0jmOcCCJkV9SogLWUWxy250L8
RH+0zRZGvpq9V2ja3Dl9m5KQOuQofjXJ131gwwL2c7yuO6Zt9PdYqLjFILR8
A3MfPhMWaJ0Hcgj59PJpUnCvmNgunjforXgHHhFOK1VtaANOLSAahty4FDJS
yHphEBUVbxUaoEWXVC4qWstYC4sUtqTa5UmeS8w40/ATtXsgxXncL4tIioAD
HkNKdzNuk6dmL3AJK35ue79TDhCtzNv+I9/nNmcDBDgaTlqQVMa0NS5OnBSI
ID3SAOlzbUG3/A6oLh+Tf8KlhNQmu4HrDMZOhAqyihVrogstYRxSS2PGaXn4
ABFS1L5IucKTLPVI2DR7D+BLXVhNjfsJ/BHGzqKuz9ou9IvDAEoOO1sapY+f
uaaWgZmOIWe4rLddmwQqz60bbVVz4Z6Q+804F+ga+Ug76vztOFEoIkuEh0lY
2AhNBo1Zcnwtk1OHzEkX/nwVsJ87sXmHkFtyNu7d1XOU+NF4m92aVYnRRrGU
YXdpeSmT+gYu4tga+p2QWuJVH2vK79lsSfAUnC55LntuLSqk9uRZhNd+eeBz
jnOz1yZ1zQSKC7Lb9Z+9a4xz2jX3f7ezlVtoii9/z3ckmy3Gn81l1ER7MwAL
lY12GdwPAYeaHo/5ku6WaKyYTEqrK/5Fx1wcH4X2RU90px18DwjUagrrsfVG
TINdffLGBkUa6JwKxDgp9rR6/c9kg6giTw5TD1VNNvTW5e7UmJ8l+oSFc1h3
R0YWYX1r8rscPoyH/zH4B7+RSKS7JegXdxF389inwIiCU/YyQ+0ivVttQnLS
EFBVMLBJ4EVWiYu5IghkRgr0mv5wE10YgICw5lm+Br0+QgsqjRwDY6PVbtv6
9WR9VSYgKazPfufaViudmLyt+J4p1cDDmEux+4QyxW04iAv4uGmxOxgWUBKo
aAV18BB+BofztMwAswtN69JypOFBoG0BDLNovSulxRmR/RhPBLp0RX8YI05p
Gz3RRt+SQdBCmCs+nan5//M4qaWi+N2ShFhEA3iTXhuj9dhEOlwvMziDDI8z
TgtutML4T0wRpNd9R8MQg8dzs35O7E+3rQxCApbvEVcZTQq3x9VDKFwhxWGF
ROtJkjCB1wVlalGttbjVI5SwTtGP1P1fm1EwpMkKRViUtBmFTFRKca7ZwGZ2
Bq3+08zeeS89exlIA8RBJyksr8+VSmhbKK5m3I/Yul++T46fV14c9Mku8vJp
W17rkb+TB+JT7sVxYROWHoxpa/jfCzHaGI+Xpu2kGlLZDDtTF42iP0AOehUr
qL/v/z3V4kU5h91qv5C6sgqje8zZGWnreN3ft9bjtAUAXuxN1TQSOw4S6Rbp
GISPn9x3jYeF84HSDWZHubG8TdhNNbYcYQvuahpzlOknU2Yov9jEEbWsrxxx
NXBqQjTkPKE78f4wQ7bj85LqZ1J4cgghDO0suSebSgbSjsBQOrAVNHklgIWT
JD+10z4U5t4tiH9dL9IfmV/aAsrYu9P4oA/lkiXDx6ylBbRVPiBD+YKVsCWy
rrNnd7EcHPvFha18s3wYr3nH0IyCXWSy/LZmFigjSuGW/63R/kNxFzzlbm49
UEpsqFJFisSzUDoPeEPcHDUUiOi0bd9W7vyiIKcxUACgdu32ZfnyslP0bHan
lv2TTvDMeXx8y4RvaKjuYVpb1wPBzKUvly3SXq95SfWwpPC+LEdhlPvxPEEk
BkzdI5IS+579iTOSwaRL/cx9U4m/RUua33FpXwULPEFFy83aZzeCtnNJElRW
1Qs2LLhm2uH8RAgn+DrzDwodZDLtD2attrZ7QwnQ/coAE5YqoYxI0YWVBevv
5Qj9NZh6fUECWhn+Hnk/fotVy5QwIwf3aXuSqKxmEcE5egaXizIvkKlNSnY+
HMqpnqdaqit7xG8D4A/PG7QBfbK2SLpb+965K2y/SFiwNFuvk15q/PKyP4Od
iPI5UeezpUKUSjp4WpNGxnXURIC5VPlZ3u0sg9rrbrJfbUPhAVXIk/QZ1KKj
9MMReYf6U1O1LykHVn5RYOxOiC7COg5hJp5pPHR6igpOtZ77KNlFAimTli47
Pe7C2vfKBa7k2IVBBtbiGqS8Pk/r8KjhDLNv4llIUUAf+LZ+ma/IRpnydeZb
h07xRaHIIAqBiD1zxI6YKKgtOgNXtTZBDQZM+LSpH7YTNGZRD446tEZmrxp+
lufoUPownOrqf8E1s6rkuReU7s2g6F9V9cKD1R++4qPiutW/tMLjNiR7LTCY
rYjxrAjzIlaeHVLY4tGAFeYIF3zJSzv7Uj5TrfV3F3f7NivxBSL4N7EMawL5
8FY+IHle4AKCHBZBt6zN7fBfVBW6YbuOsYER4vQ1OvdQkPXwQ1feL8MgRbVl
tzTB2HT/wHzMj32gNfusrahZGpxf15LI+DxYhHWjbLIF/9ytIAUunnuSdUB8
Mvl56/p1UXgyfrfiLqv8YusV5MqzYiELWes252EK/zlc+jpEeHXBeLquir9V
9xxNZY2QNtEDH4f/KuxISit3DMwRrb1b3NDD4PD+41N8lUIlRhIc10A0XIRw
swdiXnJyeiUs3vnETgsHvJp8Ql7dvRHM158+DY0Mm02yzDl7pFWRcrMkTiNU
Dx5yB6rCSHW0jWeIyoV39SWWyF253jT3ysC2Clbv6L4KU3eomB0G+PQi52hC
+1eRtRE5YZra7sRBirY9PDit7eTVp6s+x6z/ROaosTPoc7fwhhioDrp47/Wj
RZ1w4rAm2vS/KECVjd5oFbDTGcE14PmwJxN6SDdXm43SXwx0EjyNytYOKljw
J06bPxL1+FwJKRey3MWVzODRgjOajlq0bMtd7Qgms7mmdFaAYC7IAMkhO4DT
lD2iHLEEYgadp1rK19ijsVYyRc1LPd72sKQ7lu/WeF9ODZ8GXYRBs6Z0jg20
iAecrykfTOFNks/heNUHtT7vYXO4eca2JUzF3dZAkVrRCzPF49/gAKbsB/Tm
ehj4khsT09jufy/6OjCCs5w/0HKORaZ4wo077zHVgyD4DuP6o4REniGjPEcY
kzJlQn0gD9FC5DBWwohPk51M7R+8WXo7RTFS/wcxJeIzUSEjyyJDK8Y6a12W
npAz6CQu5eejXfcUwxL3KVlTTOGwWBqo8iAsZhbC4QPQtkBbyaAGqGWEIK1B
mOhPzMlAqIk19U22zWnwr8aWa3BSYiWhQUw6GJdbqsrxu/ekZdA8oHwFVrkQ
aiTFT+Wf2u/WLCFXBsLwQXntIttji8PVhue1u8QUr3pVeR71R68mgeNTc03b
IZcnCjnE5pBhJWG8+mIeoTpmfuLImYDpnGeQa0QQFm1i2VzLUJsfqTTxmMn7
ILixDEBoGifLQ1oh8r3eh2EK4tsM1ZVa8bMJf2zN7FlSHW0PTvrulg0BlRBl
ksAwaBC6HFH8sKqBdTO0geKRyi4MwyahgioIzQEMY/LFjg8eetxukrQhKKcp
LSqU6xYv1d+4JfT4ruDJY0YIIfpPyM1Ck0EWAqqTmDxB7d/fBF8+7BGMioYP
4YtqZMYrpwC9505sGyhmcztTSLXY4gid//2ujlsIDfhupGpGkZAfOzDniSoR
k506jVUyS5Z6GyItV89nYkn0vX6pS9QWUsgQ1kgjzR57Y/odY68kmA+I81/B
noTLr5/zH6SHwX8a7iTwehl/GRxzweiEum49yh+LdK9xv6mc6v6WQhKLnspT
2GYi1gF4wnsiuTWS8yYeZiBdkV9YZq9uTzncq1vvJiUIrLiNdZyRBOd8i4Yl
brKUVkhnUhUaUZ1Xn86JuOYQGOTIrCIVUjVPCJXRq3xkqcxf/cyWmmog1/Zb
6Aw9LDcwcd8GKzLqSquCf52rwWpOpb2DBi52u2CET0lhOrNxvm+vfqKE0foX
jAGeKKYt+kXuUkVxB/I6z6qEexjLl5AmiO4ElkIZRF/XiwQL1xwjkdJrX4z4
+xZ9Bgj8Kd5jRfs9NOjrjHsbMhMJPN7VIFd/sDGd1ycefBN17uJJN9BX6P5j
OLXR60DT2AL/CP0v2hBmgPAV73WgH/NutEx7cuVXxqYmzz2kY0TrvsPOFOeT
CEZvkUtNofML6jk4ABpQIQv3tAE9VsdslqVqgqwieas7Ruc5JLi+N2zc1Cg/
GPRrLDIghqJaiaFTId70aXXnMadGgx9toCFQ8n9mCIMgCYRJOfyvOfSIXB9+
CP+VGbcjzfXBdWrsfm8tpFIdCUDxUTibdDh1XuJ1urEay4K6MFMnYLNmciQL
0yBsglQ6IEVG+eU1PtPTNZ4/miPCl8awtksD8Fkgryz9fIuZyf08OkERDiHu
qRzDql9MQQ0W9g3SZTmxczgoEYqQQNgRc4WK0uDyRaZI4RA0vujDzx4q4b3R
HMDMDPP0V480LjXNoiPgzpP8jE8W34gRE3mevQ1IMwm6v05ukfMFdwT4D2C6
ryjRI+N3b6lmEFglkpee09OvqZJ/gJ3Xdpd+4iDpAw64lZJ5E6QpDmjaUTdv
4Lhqml3ftIvNpDIf7ob0i937Wi2lfvxekWMfadmEcxGJXbZR+Sz7KRSyYjFa
E/0nxlL4K6vMDC22PxZoC4Ql4aSUwKL8b+BcIBPBi49nY25+hvSlK7yeCtAv
e6AUVkweaU2PaPs2rAlP6zZA8wlR3SFdxnzRDA1VMzK56fFpUHJ9jwvUa+IS
FqxZxpzERPfJO1eEZVQ2jaBMug7T/R5MqAY6yLUciZBBVhDa9o9rUjTrUEu/
oxUnQpzDnCGROGtqcU1o29KzQoI9/060AZzfWexHX7iADrqh7NtYWVzeigAg
43P9jVPxauULUE1pF/RTS6Qp8ShmgIOqHNCMP3UqGFfO95U6L+xuvViedDK5
+ipq689ZJudxKA2zcDqF/xqDHdmm+IcFwIQuImPXBlsUJluCg24qlIHw1QQY
C0ljrZd6EaGtgURhp/OqnGFbIthY2bqU3D80IoGO5Ng2dGiGDbOA4n5OeTaa
/C167yAeV6LGQ/I5UkzlKw6Mk9kxPHvXqB8wRZD2wxsGuLv2gs0Qx7We4wBS
mU1woJh8oJOPehfNayU6qYa2ke339h8BU00aHYbKEn2TEqjHpOfwPAtxxfnB
mxUGQ7IdChffxsmL0Y1YzIfOzKwm6yWCKTi21VMmkkWWJ1JL+FqlyxlMePju
CZjzWZVFVwJG8eH6i26wnaq1h3DB9CuZQwWlzZtqtC3VYC0y/zJAnvyK1AtF
2seVTTGBM0HcGm3DP5yPpp97m15hay+hmC2EL0jnnUsK4JtSQjc2paRFwLlm
BP6QFM9QcwP11muVdPEMm8uAm5mugN4pDIedfMHhSDvYcZZZXq14wfdNxGrT
2d6jct+fWvjkcXrAQs0v2LlvY3nNiqGkh0qrCmM/Y4MahU/QA7L1d+k1Byh7
x43DgM9hP+8v/tFs7D6kxxmtLTiWtqn96TUdhy8uswvbJAXJTQTN8WJ9x7F/
Oj9nr0pg6UZeU2kydGBkI3OPTADvmnUH61UgFd3Xh8hNYaRLovaCwsQKWYwp
t5cwBBqQkTYH9GrRL1xXHAxkXIUW33QAOeOSJB7TtvMRh33GF08eMJk/ecLQ
11nW4QOC4dFwntNwIExURbfyuBvWKGp+ELph4JmlO8jaH+5tUrTe7l6VuSeE
AIzNryZfEg6nqv8p65jxw/kRbVMtHSXoTM+mFITqze0XcST+NU3u1UpE6DlX
9zbUaKRjMUM5kGFKP5Oak5LllYhp8RSmAZFG2LfB850zMmgkU1LdxFvhpMRS
W6DIo/lzix8y7OwbdRJfI8viWQM8+6Veqd1GnsYo1LHj0CJc9SYduB4cVplf
NNPox4pLzCxYCiheKMwS8GWnzaroZNdVz5fzNfbpvYihEfWkMStHwKuZ2MQf
UZlUit64cRkbocQYO6svVhFbj6syEGbR+6VGdgkDL1/98x8nrhnU36jnUty5
7dAInwBjnCXvbB5+3gavV673jEtk0HrzHhhMW2Jwom1xUXLPkIeuFhJovxX+
5pQLk6HZbDPGY0ZSqrspp7FCkqWhbn4YHeTvnrMrvX9KifMRKQ9pQBijWtA4
iQyRApwnI6ZpHjKQsYLMcDbsFPFdI1O10ejXpiYGfldZ/nhS1BmeC1guWT95
ILObKXiUU8N9Fy7vES6E2RXEUh0rtzXAjLDsL3gNkQNchCmvOe0knZ8xpui+
4ZCixtXQn6I0PzK9/IUUyJappaeyGUNaMIbln1fRA8DJTYqgr/85THe1GZZx
MpMrb6xan5hgxfiO+Xge7fYLCa7zwP+UZKqCSHLBk69HSeJZ07/bErW73ZU8
kAKcz7W4RSXl0bMNUBF3pL7tBObT/QyCcqq2gJ3WFShQ7wuOz+GrvjEDtXJ1
UXzW0zsO7oyGPSmANf+RqPkLEFKArRz/dMgSglnyErDdXp6FgcURsZLFA6Ls
KOY+zvskbXbvIWpUznX1ySXpj+IF0xG82d1M5D8M19n9+YanFFeEQ7VKggxi
TMmc44UuuD0F5x92dXgqbXYL4DdxsbFq3y1i6V5PsboTydanvMt9RWYdCN5Z
Wvh+dQF3Cze3SP8b367N37Erva3DVswR2hShia+JQiHxBV5/e5Kx2AufHLi0
5iv0hjGDUeUDrr5cJq9JbGOJhxmqjIip5kBSdkuf6mPeCYio6JE8NSCk3Esl
v+NRx+nbjlMBAmF3KYHhupXOXlHAlBod749ujg84AtRg0zWvBlqiAezB4lfi
TfGwVzsTDJr7PtjNJPbIj7U2fL5Zpw6aVTZNJx/gH2/LM6nCxzH32OUHNsRV
HwOrld4RiHcxX4iWpSGlcZeF+GIwNsjprtL7zHwKRVpBPwjzklo/T+jHKHxk
0LpCDKBleynlxutZfeA1Kotw6LcmsEEvW/Trf9V/OM33VAPT048vmuyV0FKD
WQZ4bzeDWnvu53rbXW1GjZC+lIBF/rP/FEMv/QdcR31xIyenQxahsi53bVB/
Aydl3283KyzZF5ap7dABb/BcdrEGeakrLy+MorzieqKlK8toxVxAvEfSip4w
4mYSAVGH9SJ3hbFX/V9S0qEKIai7dn4wGKfwdJUXVpWS0AqlDLW3XkSl+lqx
OZDtPtsxEjOIjy97JIu015z7e1+iw+8Ccm27nf7hANanyz4UO61I79HTovhq
HRNQc1iydyV1qZ0U4Ymbwdn2KTT6b1P9BcwSi3UmmmOnKgzqEQRwBQCfWRhM
7xlAGMEXzOwGrDqrz5OdrKVPuGb5oOv8+RPWOYzgTAM/4vfJiWpI0cfYqUMR
63PAhciS1ku8/ws/tiL2Nf+O51kIs2JpMBPKRInwAov9ArEYYzGIXPUvAscx
tBaRR7RBPkzXrFzZIzvC4rD1V7PzCTsAYVPSlugOC2YUyJpmQoV1YoLK1tqJ
F3I4QQSypAxaqr2PtoEfa5+DvQmVYspP8DIaeZiH6stqZqALmQjI/pmmL2Q/
YYvyIAI4JSjU0IanI94y18np+O3AATLmwVR3k6lc75HMvzsvr2oRg4UMUFyB
1CZGsfAHGhi4O9jnNTlkw4KTSp08M4wVRArszK2s4+i/4CcCcVzrOE/KPYYR
T0O866U5fw6ZGHwXnEhx6HDAHUBZz4MxyfjX9SNPKnJYLuhZ4iWQMuY6YYfy
unV5F8F/+SDtN5RJlYTk1Lu9TpBJszCmwTBzh4gQnADIe+1Kl2M8l9mQmfc3
lVlE1xEjpeuBAcj/DeVBaDL0i9wpfJfSFKTNZRFqziBuxtJOayNRrWto7wWX
54Y+X+Nxq1i9XJES+Xfa+AeQu9+IBUT/jVmSt39lQuTVHiacJlEv08vsMQZp
Z9Bjmbt+5kqKH5K2mzJ4owugF052s0s+Ga6lxCM7Naz/QKciNiyobKYTS7H0
mOI9ltSIkItLUMp7uZyqr2s0O4zaxxt+mtZ48uHQMVcWS39sCI5rSpWUXmld
YS8pRtk3+i9RlbVFH4Obwny+DhCzld0a8sQ+MEahZ2pmnB9ogQdG6LV3G0u3
QiwdRV9P2o/aH2rQyz5eyKCkBue7GDZQHBx6pnR8EaM04W1qMuKx9fqEqKUi
ABKR/e5AJyxrt7T9Vnp0eT/Jh2pj2M0mYrKN7jSyQxSQQLHeFbPrepjaB3sZ
oSbdLz4xgzG63mfd8nMhOkaulCiZxTQYJpFJYmJ3QFSWVWPeNbweUHpsZrcv
XF4/GHs9hRr95EcHzu+e5FR5Yzmf1PPePpRROxVClhw9jyLLpxHNecrQuOmY
AlhkcKJklK8wHAsJVrmJ8VOuBFwPpjKa7ucsqLRLGw0MfvjDxqUzEdH/+778
PqpUu3wsT3urALz6qql388OjXVfWk7qSkzkG/BpLRt6oIRk8+nrDGfT/Yq54
p1HnOQkL5NGeLnAcVSSXKelRr6VivDG/OR5FFcpNghrzkMaAkX4/rdvYif5p
cFA4Q681HbOUlyq2k6Pppqs8aa9LMdDQGRwm0vqJ/pWSRY03OaOM8zIAvX2C
b+e/z2IiJu6ENNuhE9r0ZEmPBWw2zJ9066hMtogh2Pk+4HQMkQkMf2PkhdBo
uHtJkMS6y/6qOxsiXN9/Jg3ioJu3LZktvWZZhMquqFu0oeARbc6pEGQF3M5L
+nwXD+YOtNmhRSiQBTRG1nFsEhAVb4SGdcVI8JQBDGlsV+AS9m6rmnGs003M
/aUEcGqWLYVUCFDzWIfee4ikQBlKQDrGerwMMdbsFQbbZq+HTwKb7AhanItq
F/nN4eZAAvUvLqYxhAN+WQUd4HiEKWZIrmoXsofLdImzc9Lp+YKzEUuZ50MV
Acq/A5F2Llz3FtljttMv+YprHXFK8CN70PiWYiDCJDbE3PZEoRVYQmb2aJg3
daeO52UT9J5UxcmNQqDmCIU1VcMmi6llY5xbWJ/xpjJbu1PI6BeyncycjoMb
2JUpKVUGyNDvIiTvnkwFqetfNgRtaWNZlts6cE7iY1Ean1x/JEvOOCli5oK7
gdyjqqj8qPr0s8G20p+E19k/0Cs2xFUuzOOK1san2UhFCfbUqClPdewHaR9f
znzwHcDwGtJwB1ejKQRIwFC7KGqa8iqH0fZzRZRdgB/L99kQ4MebultZKFWu
XFpinyVZ9U1WjZ3ytaEF0GhDY0TJu8QT78o8wHBHBALOzJ2b2Ao67EVO18Nm
JbMjGHcdKP1LolHbS6tIf3Q7tEdEzcRLBeD+6LIA7xAUcr4FwZEA8h8nehdy
exVgesA7xIc488pfRGAmpPgJDnMONFsd4Cleak04gNZa9PrANea2VsG2pO0M
HzClDIZtmuAepCN3MJA0d43vOq8f7tSKl4vxA/Qjs60R6xUfSu6YK0mTFtOB
aoPHE/bN7ccBNeSSv6nY27pj1nNCs0FQdDLR0e//iJs/O20XOa3Yl/W2HhsL
dkoUwJ18DqYWpdY4WtrFcZDmQgNEexdkjG5sQs4/Qk3Ehbl3jMJ+PVNwYlkV
2oPqiD5Fq4/SQLkmV4P/fRwglEZbcQidFcGRU8eMG+dYNfENya5FDtSFRjwC
XCCiS5KM8k8A4a/+8orwqlk/bQ62Pk3fwHk5vCWnPBc5EXo2qB79tjZQuVG/
lozFSGZk2jwljkKo9lrigDtb4uHdQGA76BlJKPOPEuCrheEQGYOFFIAGCDjU
Q3pUXVzawH/F9DUGcBHBj0iNBYaxHvpDal64Ig1fPHTl8GSF57/Xe2hZ7YL0
2hyt+p3dTw/vF/+L9jWmmXX6OrGqxQ429UbEIIS7a/nD6bt2j/3LW2YrLrnD
b9yiOfbpYO7r1+FuFcT6rx1tyxvHXBSRHLFrGiUbRFpVNeV0Hje/GdJjJNCa
BQlE+lipUlL+w+Y2efehBwcufoG79H3jz80G1kxzh2jwCtVUQe4oj6XcQpGI
5PG0+GIm6BjU0G7b70uxxW7HenMSiusrZeBNsJxDseHP4qXEDXWTcwCfgD/L
uAvQAFNFp8B/lgRnZvSjavMULq4n99NeLPdmnokwcP07VNren3IEdmTtS83m
myMqDk153WiwdKDViVmjXZYC9BsVZ97LGoiqXBZ6epMi9nKOXjW48R6r+9vP
ACoU6ZzFtR5cjmdt1c52i2TPcTxoHLVHydO2E/L2Ryvvx4y2ZIPjPnda6uId
PYkB4b8Lgo8oEbew/7vxa549oO2x7J6YlahbGCgpHmRWVgNoPyQubqbQ2uBo
HjzUaMh9Yizq5COKdJDBciqGNyjCX50ZJZoNXtRlyg1CzfMSH8ujO77EjEai
6wjY28Vn0Gj7HJR/GLmdynR8kdawEdNB6UrPJUSD0Q+no/q3E1NHxHG2Z7kq
7bv/L/gVH1apGNJbV8lKmfv4HziExb1iJPOM6eQhvOHv7y0f8zBZGSn5y8V0
1iB46gMZYikRJRVSOQXOS+JSWD+zumr7+19VQbFXVvwXMQ+l9v503MwZveFS
56a1OijKGzpAQ6iZL20OWFPbQ5d/sJ4GbfAEeEUyTZPFATi/WcqiWC8Faj0Z
hrGIocRLW4hjycYzusfhjJiCZYKTa+Vau+z84+mV+EFZ0baP86eaEvlZP+iW
nYIFMfMSEd530J10pvx2TRSscwZlsuRinhgrtGczS9aN9apE5iO0oEil5rwX
yR+xkGj88KK7rhBypkiguTqdqgPov/oFKqajWdW003RQRX0zRabSS58wBV3H
0ICnlm5BfoiToIRyJUlPBvc3OWHVvuL7mcXpOMT1wxdgXSoVCL3lXlBU00zF
oQIPH3P8YoYCREFe43/SlHtDdmEqye/r3hbKxxgCU2ZuI+mctWf2+7tHwOkB
1tKlKwp6u6uf4kqDp6de0LIVb5wgt25xMwIHG4IfnFtbwJnJvoxelzUJOx+7
etcVMCSy9BJbtVFqe4ErJijUsnLJ7DDT/3dzkfPtCNZ14x9w7kLNk0lLZxRn
8wpuIAtBou9zmQuwwK9vR0yEz+GXA4PuRL9mYs/bOeo4FkkRthpZcCKs8Mrz
5e7WXn2x7czMJLaX3BdUNfgc5+tFEQNYOuhPOP6CrwYOuXFrWNpMrN9WQmaq
2QXk7Rx38VHUV5n32Y+XKQlkLhwT8fW86MnU/i0hSHnREoqfRyzjUs35R5QK
DcSbQIvKo9IJ04TBorpYZLgDiSjHi8Pj0P0LEXKGQbUulPQpFcfT7NdcPM/t
fQxd9ET2Cq05WTSYNc1J4522Nd1FAgH2RA9WBE4UCEox9OwKNI9BOierCcUe
K6ej9Iyo4r2cTfLRIhnz7UlHtwCJrGczYM53Z48Xx84ShetlwMZBsTpXBBLL
ke3Ka7dsTt5dghM/zobm8iBfCJ9I4/InwO1miN82VtpED1VGil/zV5iCISTq
yFdlKnx/SLa+4qXtx43uqxuETVxq4Si+ELNmTRXLTuBOlLogsocGG6/XVUOo
58gAo/aNTwjrPfdIEs346tepDWEDOktoGogSrU+JNj111a9ccrrZClwoqN/Z
4w696efixc5rRk3cWB2vi/fN1qp/jYtLz6bPLHXoeby9m5rw5P28qBsH62Sa
GJ353WYKG9bgmPDjqUWVO3i4Dq6eTAYRnFEeK/JxZb1oH+woaysnWTyIzlp9
3chrqFrt5WhKNm6yU1Dletg+yckz8vVFW38NkPTW01H9LmfyHm0036iBG1vL
iRc/J5xqF0WEihDi8mrCduAOmvfKyFHFwENuGDbji+lqYzvmPcuoPzjjnJxc
25leJD/EAEY4yqqsTcrg9g1nfew4RzZCLMJjBAIFWiGWz+bzY/OEqIrvV6k8
8RK2m/r7NjZZCH7WosyT0LK1R5QligsUReFFmCd9luXxqXok3PKxyM4Je8uo
HwW/7A9Z25xCN2uFnK1xv7vmdWzkn+3otvVqeNbWmYLUYV6yuSqJL7AT5lyT
wmGcl9T/noo3l+Ab7M2uc70KOQFypkY2bIpCKA/30elWMExFVWdKGqFV4JFR
U0XX8JenhiZO7L2bX6Qnp+0OnVOUn81FKLOEBGvZS3Nu903uS7FoYOZ3HjeK
D2r0Gjekx0MzBrlkzdpRJmleyfVzXzEhj/cWidxngzhgFrjzLJ4kfjt+XQNd
+FIodvvG99R8RflT/jrjwpaIrBu++lvNs75QnfqLHkjaSwd+n6elRalodrGS
37SHhhc3pqgCS2MT/3PDvwqh8u4O1Ck/Ps9B0lxzwod2WPqmDM3MDoMikXjC
btEW6Fa5xctTWFVfwfbXxeXg+NjkJs8i0Sgp0yoZ+JsvTs4D8NgHKidbMLn0
MfZ68S61qBciRwc/7t2qmUTsOa+8Mi4clnFlh6NrML5I1nPVSwZ08t8wox4v
YTpbhMQjXxIOEsrsghTK6G82k3tyr+TDRhw15d4sXk+lGrNStRjL/DPu9NQT
F8e+OD6PBBkWOUNxTrHkmqa2fGixCahKE4niSCggjpz6HsIlbG9lvz7fEo3h
9PbYtOUXpULqyOxNwilE9y21AVbxBX7B6HSYNSco/JAbkZG3OJ7BAvlGgwgE
BjzPYIwFZfZehzR0XKTsWW65m+yOo224Z+oHadAWNtMrRv6QPsHouKnicB3g
MNdFahyxgQ8faIysjKkqRmgMXFEKQNQbFk3CKLbvAnfAYBzFcoM/IGTLUzgJ
DbW/WdnBrUhGecSdMA7MxN2ZG8lT3cfSnH5pHVJXt9Znmn+x3PeBlW+d0eik
R/qOqTptRdYDJ39fwb3KqQBfkZlZ4L9tXjy9B3qAKzhu9k7H8mB3pE+vATKM
+wOL4Hn9qwEmBpeD9sYVclZSgM2gBauJrHV99P3pIz791KfNSf3h1UEgEHOv
BiOWjTFy+EKMHbgV9+1lZ/pZoyov7hJYkb+IJUWI5/unpyet3O6X8jJgLTR0
jeQSYOSWrT6RMSbrkaSDPK4+afqSP8cnLnP7ZOpGqcd4ekybM7NPRJpMVv7E
HmmfU+rXBuN0ln6XECo5IXmtODo9IO1e5cH3VXghnG6hT7ciQXB8EKbMo66J
+wL18BsUtl6/kKe4sxOLC9zWslg4zhdIEHQcf7kbHLPu3JDgc0RmIyLgOs3D
6jPjlVVEXGgLThfC2AfXg41r9qpEL4HXzhdVX+U8cNo3PlHQY8vJjndx1JCI
Q3NzyX9pI8cjAobJSeJlVhgdSDqS0+Z+u7fCO95X59qIivsHltTOaXhmWt2f
Uu5hKNCyUM1FrLk/v5p3/BcDIHP/Kn8/XgUeml/m/ZGZhcnrGoRuQi2lt/pi
2pro18t9fq/8Ubsm1gCdQFN9Ayf+eZ0EtreS2oc3BidE9bt0f/yQJIGRspnL
HVmYOdB3bxURS5E5h/3Oe9zYJyiaIxr3fRQn8b2HIvtM9xQw644vzuXrhY84
eioj8AG7dTar2zzFfq9meYcTWn09FzwB9KaZQ33MCweVu1VYJ/GuopNuTdMW
L4Luah3VGC2UUeWW+zQQHpTLU9QZ68rLRd2sTpydo8GNMWvP34igzIHCNne9
bs4VADh3G8VnEWeZ6gHqrqrdq7BbkCpyeK9PwcRp1e5i3Nn5qJkkWWvxLrYX
WWbMS5bC9Y/NQwYcPi3Gmq8mA9hnraJ8Bl+u53yqJ7sbyXhTCYTw6lDfkLvb
/0+ziEBa8af0tKAZDZ+8DPQHu60UvW7xZbI/OH5SedA01f308lI/RU+HCEIZ
hqGmF5zIFVl0L8MwB6M338TYRtdtS97hfYc7XewyghJOwh9DKWHZBJMfdF1r
a6TL4gYIy+LArBpgauNQrwSPcVDHRxPpFfI5tlkquMtJ1wb7OP+9KWbq/r1S
7tsFAx6QMITfNBALA/39vpTIWTkY7a4rN/tNy4g6l2qQk53vL6mINNARXEID
1h3pp5eza1tIOiBM4MYaVhQyauNc2+ILim3wKX3M0IIPf3/BkoNdpl0CkrZr
tSU7VUXGKqz8vR1ZJVUEjVBkm5wrgIWkVGtpd4wtwzN+tD5+LiLP9VchAc9z
NrSMuH+SxCU1LLI22PPGGw43MCJddb6sfuugXzoB1QJ09ZlnCqraqlvo1hQb
FCIyVYbb3IhahjXoPU+Z2+zbOTWH+L48OrQKZt/7p5MpriwMXNQhzdxwAsoT
mvS+sVJo3ow289d8JZ99FajuHeYfbtKYlA+C2ZNzWkXLbrhrQZfTuHLpRKLJ
rSavF222f+SWLm4VSC2TEh9OO55Pxh9dHIlp5swxPUcz5G+yi+txoYRvxYVK
PahlMkCwoW1tx0IfQGF9l+VUgNDTibtEU80BI/KwTu/I39m6zILcSBjFHlXx
T0RzSF8GkZh0gCFqQzqSUy2ULeQpZxbJI4ekSxRnFLCF3mFc6YMS0vxxrbNh
+PcGxdH1NF4TZB12SRXRxVdrZ0EN3kp7G4xc/MzSu13AUAwCAluEWmzzBA0H
ZWeJbGwWuDb5o0QHKMmlVctKXW1jcAtRidJwNwKhZABIfkWjgmxalbAxzH40
ZPOlAS56cbjU041Iv+xApGZLmYcYZeLm/Y7VCniNObLzaErDtIugOAGEnYEZ
mC5hQmfx9rf5E34C8zhWF4NBGn4KDUbjSo+k7RItzq/atrhpkuyIY51tVyyQ
HOpYoivbOdB5TQuo3sGrVE30+6yBRRwjMzp+gRTmHO00lLpZxefIwhf5EczL
N298wGRba/csYK9MleDaAtuFqAuF1Rhh+IUzXhjVQLfFpRWqxbXO/qtuVdQn
RbuGjD3rjfW2dPLdWcQ/ClH+SWDi9LZqeUd4jeWoF6OO1c1fAt8kPXwKGfBL
3Z+a9BWHtE72O5PsFozOXFcTc0DOBQ+yv7sU7NbzzNJLGnZ0EhGCk93tl8d1
qtBUYvOCPLncm9cgSAalmDLjlWYlnQYlNl2en3n7MXpsD+vhIVlqXnVFr5E8
iqR+6sZQ6q1min1DGLUhovWl0ue64sW5r3x1iefoJxyjUaEkcvHqIIcUvi6V
bf46iRZYqmPuduuRgQ9BRXsR9Kp4R52li/0IjWLFmHIBTOmke2UyvcwzRNF4
N9t3BrJjK07YAjU/xMMN36nYVv+LrYYaUIRHCrUTL/wlD6h4gXSOlgGUhfRJ
7Kd95yPbYZzoz34kK6aVtf/yKYI51VYjN6kcXtuG/F0hMVPDMvqz03XNpcoX
9NjBUGhL1SfETSd/ga6H4IYCS3f8Q63gEWr7e49hmcvEY5qpzmtPFGtlCRUz
TgybCKhwLeOyTmBK7rnHk3TFzHeUhQQi4XmLOET4BKV49lKVeWHZ9CTK44z0
B0U/f5+0qZy19CNAOj40cK7QqhgihbxFcNSy68OLIZlNSssaqAAyrUgPR5zg
8X4FOgXOgJUMgpF+xe2Qfb0q7VSnPXDh+MwKqc6S1MwdE2HNmOoWjwIrVL57
xFfVk8Be+pDIvcfrGBKbajCiHPZW8hIJUuBgiEjhO59G0mULTgemxAo6jnnI
vgxBTKy58bMlhqzJORezvwxLXJcAwn4XewWpCe1yZejnuoqhNdScRnxcxouT
0WqdJt0hZ6DZvEMkJHbQ28yXcFwTe/pLL4eBpIrq3rh5er3u7gMQUPlU92Wn
qPIH1VP/xjveI6aZA603ES2VWbQa1XJJavDFh7UOz6mpjfl0R9fNxa1oiViD
G7Rb4by+5rgX/x8ER+Nn9PdgQnaWamQkIZwWr58VNyAeG4fDg9/du+rzslu4
ApvZfWZYW7kHXTs9l3DMqScWLJB7p2jvetE2QZeRktRXI18DJtlQGXdUBR5v
D24bXJ43lq/MEXufZgUaT8eH8N09GInGBf0g9nMb1tCjoYkouQVCmMzLK3V+
C9zUqqaCxXdUxPMn6so/F+qHK15oO8JGE5BQOpdc+oN0xTb6Gz/RBWn+tcgC
ev7Ca11D1Rnmpg17QtD00/P/aP4yr1grcpZVGVdnMTfxNDIN6iWrvmACQXgk
TXPiswSEw3kW3AS24A/PDoDptN8Z8YUeOZ8/qGJ4VE0YmtBhXQbJ0Unxb9ZL
0PyFgmv8bfZG3hEMeB9xMojfYv0DxhBfm4cMLN6xGwgusfY32UEVlzIGFlxm
4rNM3FK1ODgVuCDJvn+78KUx/YX2u+tyDLPqPrE+dgOFLkT3tyAqbm0lyqei
gRrDPHSRgyjNa6RSnOjhlmDF7SA7BtZ5HyDZc+Ll6s+xuUc8rJgBwUPWWLlR
sOf8M0Bl2dTK8ZgOE1TgjTqMXbims7bHpoWjDKLP1gvz7gq5k/SQn/D6+E3W
26xQ1QzTDsPoulOoK2p4EtSj+swHu8PAVc2ikhdJ4QH4nNLyL1ApP7c0T/nC
sm7DHwFGR31j4nwTVlmGAOsssCww+9fwD7H9vbGsfKSDv9QHWPJCnmxXCGkH
ePhgQ0PKeLt66bBY1DcuVEzqxcTLs8Ge8UX4H1mUvK8oUe3J+SR4FYKbgp/b
93piJJYvpJviNBQO8+vt4TLFjSCgZAyt0HlvYmRNQl92ua8CZ5AR4QarIt3D
p9OXU15s+3MRoi5t9mgV3qQP7n5KrQ2fZ8DwibRSgheONyxMnTSJdxYMmYyc
JtRC/HZ+wmY1MaFOaucasarlktyy3ZXgvnR7Y4unUQiP84c6o2mHyRQKoj9p
2vEyz/zkiBiWMM5OBbQFFlN3QXdYrFEjnMtkc+1h9M296v20Z/MEFHi9s74n
xqqB71QJay6MqQNxychWiTNwrsgUXxUkaAHX9YqSpYur6KwKjJ3IYnPq4OZQ
ZiF0uuslp8uAtFotUxrf2BgR/jNgmO6Q7uUrqM0OSoKTYtn2sAeSxTq0sYxG
LSLY98lx1aa7rUM5miVYFZ1Id93uLZ2J3DVLueo5Uv+Pi35ACh1QZnUlXCQr
m6CB5cVzHv0YEZOHqWa0mtJYn4J8c1+qDF4xgowQTHkqWfeaZTyEnjIhU5U9
FGI5e+SswJQsqGuPaDedRNKyyLFPCfTODtjwNZ97UxqVWgzDdXquaLMCrsbC
LVCjWl0wY7NzDlcok3g4N//b5yhX5CmQzKsT4TGtVM14yqKxd2f2o1bzrsPG
xfrVb0mP2L8OXH/L6r6L6YphZ42suFX6KDW8ut/sAdcLbR/MrCiYzD3JInXz
7R9eOguEBdFD5spPZDFxSh2C9vquAv9fGT1gZU4ggRCxKc21NyR54TaA/n4s
hnAnXBx9n4sB2IG+hlmZJhyWkGEA3i2qIjvNBF8nhjSse7VN+f8195ui4ERu
Jj2I9MrxmLFZlASnA3aFGxDO/NaxXdigOXrbD826ic3zJFdR5VMejRsG/U5S
nFwweRKZugLDRXTa1kkIK3pHqNJX2O0TF91/9hkzaLKZM4+C2qVDcdXYJyM/
FPBW1YUPA3RCpRR23kYVtvchlyNirkFHCXjUDi8XZ99QHhWiJZwUPJtOdCeJ
QOI7XbqpJ67C0wbqgPiVdkTl6++3Nu1GwhwrDvt2QWTNHTTBgux4l17RRrl5
tpR3FXmbUswwjI/m06galz2sq+EqekrYI4A6wP2mcN8bocO9qckEsyWuQJ92
KM1BEjKMGRs6t9g262H/+ikPFdVwh7pRvOc5kexNLtTKqI46VdZCa31Mu5Nk
VcK5OW2dAmkOJV3KPE3dsSg9xBcCcLhNWrdMEP/672c/DXvtKdTIhErBdflm
2R1z3TMogAdeeo90nx0LwRacu3lvh7+1PPR0N+L7jCZJq47OZiGKEeHbMEHy
NwK+TVoSuTh2RHb0txqyxPNov4WPRvf+miOIM6/ACCnCeMIY6uIKMOJvUQAs
v+5MAky9+TsoNRjYSmy7o/ua1DU+tRxjmlywQ13fBVpev59w3oodWmckIFOe
1GNLeWKp1P1dip6CzAThzyiHSoRVl+RIbVYM8VU62EAt6rwqpyA56Kj2cJfF
Sca14yRs/k86aas+LhZLWZzukMlVckw9pejE4DroBUdyJfTy/AvLJ1BJZSHV
DMBoXYMTJIQCiQZW33cPqwZu7WFWMjheC1Or1MewFK10z59iyRU87wzI88AS
wRU5ixJsTm9GgTW/rxd176iXZfkkUJ6qqGDex6N+UXvkGRWIcSEMu0gXFBD/
Fs0pCPh16ZockirUtxjoQJlabebqE5d3nepIagbYC1I5xt2czYVM15Xaw52n
sp/G0agl3oaU2Mi5RnXJ1PtU1G+yOKk9QEU+EhkAptNvxV/rf+nHWxHf6DpL
Pk52N27mxgC4AhrZ2mI0ljW7Y8HHxRKrhJj9je2DcE0jcnp8zxwH8LRr9OQ/
Sygz2qP4m3MdG1/yTavgOnnffij5G3D3N2HMOUoYzfKGPEPviw3ZMAPuEB4C
wlmdZzXY91d572hpa+e8l6VsGuUhO4+TOKBp5apf00V734CIi6e2EY+lre/t
+6D3TD9xiCNwYTysvPXefFMI/jFXlBy5avXTBFwznQi8G5FhoEpoN92OfLnV
e0lLpAqCPzTNEoCaaFtXnDhf0Il9444swK4YuJm8vWX+vZNC4eqWHUHpUZ5z
IwjWXD1MpbHxxXySJFN4q7RaXpinrj335r8XmemnC6UbHwxLbLEtrCjgaDUQ
k+Xhti3QZfg8F6kOsZBacHvV6PSHIoNWlz7GIR0wfan0FdsuAoFSc0f3ZtSc
Fmisnecjk3SzjnII6bqXOG6+GjySo4JIY3oJJr5kgA5eyJWGO5kwjqUG/occ
xeXeY1Jz/kGI7+hwOr6BK1iZj7963H2ipnWDVxnDD5E175bODQVWFS1p70oi
2tnXz1pItpaD0PCEu53w3Ftgh43YhR8bMkZV2xD0rQqq76dw5+Me4/DUbxxX
ECvNkpfPvn8sb6C956XdB7FxJjaeraSyudraWBeKn1nxJgvp2DUyCmMs3Xx4
64oFrnSmThEXbltw7xMIYm9x7bROOS2uuImJ8+Bt5o7o7Ot0WgOAaXM+JjDW
lFEcogKjwN+F6Zd27TZfSsteMYnyPPH32ibCZv4dZ3V0DBeIZjUXH83GZToE
QVm0Sxma2vlZc9PDgItD/3nr0oV2qOuUHeKQDC9ekqyuXaDNmNgA8SVHKR+0
4kd1Df8aSbavnMFZaYoq1fOlwhcWbcX1Q7mvBk4zHC3ppM8saTHdKcJ4L4Oa
rx45TQOE38UUJbJ0bPH9tFIQO+z7aDz4/5O1sIpQULC9KzloRvSW5QoNqzXT
TnWNon5r/+QGKnc4euduBkd18LSTSo6Fk7GyT51WNvF5BLJSwVBg1Ji3RSK5
v95ZQqXOdFttmbkj2u2exSzXOMXFP0W7Ef31yo00TDWgKtMQSIEB9x0QzzrO
DJtHJGN298Gi0Q9wrVKIrVhkoOKo3eO4ZW2s6pi+k8hD1aPwrUwwYJFgmFuv
17nUZrKGU93FOVLLER5PQjcF/TBboaOCsGqT/C7nUnDIZcC+Eb0HAE7DLrcB
kUaUQIvPLpIEeVDdDme8cPAMuwwwgAAHL+bjunCfC3Sye1/idkzeHLjWlctn
53W+NZtUUhBad446cQGN1e6suNrEjs6bSPMHRzy+ReqlRqALF2HhSD65z9fH
Mg/m2gTdSUd+pPpb6Qt8fsz5w16Y8cDEZsEiLcxqH3QEoevMQ/wKxuTjMI1h
nx1eJOmq5AdOkgVxHjlDNpnCUQb8M2sXLkmLxzy6v6F2wAnBVy0Quhs9pLaV
Lwyg8rdtyoyOGGra6xQACBAQ2YPE55ugadR3dIS44zLs2Mil0gkdsvzohzYF
HPwHLSuFmuODGYDL8E3E/Xd3YEx5D6Qc1MvkzxtkJIq1YUQgKONS4jaj+1r9
wCrvFVYAyjUP0bfKTliaucqcVei/6KZvHL+ghoqoWRUNC+cNguxmKhIEj8ns
Hv1mwyor7DRvxjHlLh4sRLM+zmZE5NRH7cQnTnBtHsmPSZjlZtNrXICsTlE/
AJnepGF55fzDIfEa5MH2aDnNcPn5XSvdlo1jfGidHDNV/VvUczZuRddccznh
BPNemsBUMyTUlge2re1QoQqX2pGlUTHDvQv/NbLtgCJTTgUjz18dFmsNxjMf
/AOx1j8tR4S9E8Gzy/wHluuxK6KRUYzcCvfLNbvi0HrfR2Nron4MOIq0tr+c
o0Hd93Vt8/TAsJRMqmBAUXbcHT7Esh99jd2IytuTkXW060qRLKSa5KYrmnGs
fX5VxOqtarfzxbGPtvWRXHv306LhzE5UxI/2k9cPfYE2HiYJ86tZJKDbZR7S
XpZqRJqzK6cAcQerCypkVJgCW3prdCqJ1xAQz0ahyalzRwFnkHjW6FbrNb4D
YC0EcM1u5MIxqi0oDGUmamkcpzYXWNU3T6TMszig+sMcnKiNyudlTHL60GhP
jl3A8hxQC2SKz0q7nnFYqRNRHBRoPYjGl8dFmreb0igfWoNk0+wCM3R9OQDl
yu96ewRoF5gyg6374cHVh1e9Tysdvsy/87XtAy/exLFvKNKFFWEn4r3h4gU3
iiU1Ppq6pEcpghfQGNYubfEd8zduTHeWfBwXWSP2YTiXzqKCuPyPesbiHLyj
9fvOS/nZ0ycMZ4v0E8o1j09PQCeOELA7hHL6gq6irKa12kwp4PAQYSwtcSjM
c62tpdhVt1deBsbfB80Ay6z6bcwZ5riEps7Tig195kJNLTqEcMT/1ogqJIYS
A11/zGpoBuqFKUm0L3gWrKletFum7Ae9TWHROpVJw4ohI4zC6lhgllgicUfV
lOiulR2EWuwcrU+i47DPYf/MsIEiQMosr3BlOZWuzAN4priDmTfiVtsodCgF
+f+46/pOYULKcdL9Tr60gZyZ9qsxDieQYozMX6sLDoblIcoensBMch3hyC5M
zaB9iczS9CxObECdySrbQxwpUkEdiuiYEFRhXJpBY/CeMJhCz+ZAuvgSvMBH
3uv5iYz6R1M8OrDc4DIbFoMojZmAOIPdSiDQ5KKGwmDItFK5eFWKQ84rIIxV
TcbJRjPQZPl13BJrrkRRhD3W9jEcb1pqGGfEvWRBOhDzYQ9VyKETRCRuYPhD
O3NYd8QPaVpCow44UpXXBgKTQDZchuyYyxWEVnWMsS5Fdi5yrjaIHBnMRF1A
NKHuV0U81kFCeIF3lQeUTLRIWlKvJi6xeo8/QcFPtp5t1WFh9F5JeRUksHij
sEAC8dwfzkhcqNBf2ZpGyV3PIBl4oMvnI48UocXsFIEGuV2WxNlv9k1iAVZX
VdUZ2IFcGQvZFo2MIRYymzwafxmdESKlY1KxECTy4bMKpaFyT13M49fiw6bh
8pvHK7b8pYjhOfiq4+Gyg+av7p7BtOe5j2M9YqSL7aVH1eVf0lTeE4y9aw9V
ZEFylHzgE7cnz6her4TfReRJoiDwLsl93gsv8V/lVfXhY0y6chN8QU7iTKlA
NYXPsIql84EB7/pVQkV0IbQakACOageUMJPXvHPqC4bnqh3eLHlSiEdNnwbk
nycGGZyQRDEZ0rM295+zIA07kRG9XXGkLwoTIAsSFvP/u0xwa2MZjVdxIABc
7rEOwNIjIyGj5PFgdcQBhXngFyGdGAOC+Npy02dFngCseWcYYnhXJLm5eZKZ
DGzXt7V9Ldc/Ihultprbge3D+2zQswxnC5auGHkfMtACpmeiSncYQpji6WoU
TcfyfIeQYHUGg4nKK9/4ZXfj2K5wOJ5Vql475Tza4/ACInKVGyENbMJwG/n0
nXlx1WMUyGDbViq2pgaJOrHEwBkHAfPnIP+lBuV6ELIiLbz0YUBIXDWwxQxT
BI8GqBcE674SfU+KjI1fnaRrzJRNg8JDLlPO1pNcH7gWPUyIo1c1LQT8ZFbK
aCO4z7jFVhknew5VPeoh10jyF3L/giNxLxRthAR2zyxFTjfl4gMlMnucoK+M
L1remRgYJb7lSUrJbt/FAf/5ExrP6v/LF6K5DJ5vicR0qB0pnaIi8vAY624t
CDOCo005YtB5Y8ok+XoP14EegSrs6uSa2OeaNwMYdnTtKlbfHbrijuqKRmeC
l8K759msCxi3txPbE1n5sw9TjEZy2xgPKUQ45yjBJw9OdiQHUHnXb5orItLf
p9U+/l+0mgwzzFVHxRWTBOyRZzG2BwiiOSnqBh4r/CTDxrqS6ZfXRIwm6cFD
zlDfTBBpX9wGhucCAKFNYOypnOnSuIm4Z8nh2YLWfAWVFSzbflfzWEr2R0fq
lwXsH7hXnhZQYoIYv+dzko/KsSYtlGk3PICvoBVT1kld4etDv66ppFXcLn1+
Yn9u4+wTiaZ6g0DIuFRCeUe3yCPj4jd9wMLex3UpJh+bYH+Y9GUX6qrPNMTS
vopbPkWZy8ty8H2dRdz09Nz5LwE3SiBJj0I1/LpM3KY1wguZ3NH1A4SDNi5b
rsq3REDvTtmXMLTjsCh5eQXUirsgftiVWl2FheoMBcHPcr1LJgw2c3NMqGeR
f+zbPjK38PLoPOiGSYdm23C0AfHnflBplZ6D3lv52J/zNDVWxkoL/SXWS2dU
yx2ngRvNuOz6127UnfUUpaVnZLgBfA9A43yJIRajBeC4IbxXlETUXwW5xb66
ZN2lxWnEl1pcWL9reNT2V5LxUgUtgpyDu6rzWmF9WMziHbasdUC+FVunQTUg
9UqDmjMcFheJwA9JmGNkjAlb7F0KiZrMco71q2q660ozMV8QDj1UjanhyPWV
nbGBQwOZ7coCdKaieMNV/L/MlQ03+1F5t/4DxZeCQx98m6YmgS93C8z5xH1M
+l6BM4WcBA9ITVK8Ok5qfZ40J05yL7FLBInHYCBN/Uk+weYU/oL9Ne4CXX2g
681+L/nBtz+jNj4/k+Zp6pnB3K3Z3e2FBZQtw/gIDQl1+m+GE+37Ru74ckVC
Y6C1b3+vqrZxhdcOiIgPsajPpnZInRPtn+xovvouyuxEpzAPwMtIGnmyWFyB
tPoy7+WxS3TiUp13FdssLSHY7ApaIVO9APZMhfSfvfFXf/6c36jNj5qLHlAN
kTbIgkW7J+9Gnh/m6Vvp4ooHjKeHHiXqA/oNwlqZe70TeViirkT9rtUtuWRl
e0S/QX5v6fzmajBvA8XpYfdWKYb0zNd9LdqT58ZDdKKWGUFKSeLN/BOQZ7U5
nbm/zgRWqmJWyRA+vjB3GTa3emKiFoLKPl8KY4HWwSvIBfp5qAgbkqfw/rgy
eDk1YQpI4eo8PWcQ+U+AMBkEzpZQVa0uKmpRZZzPwimA6vJMAYNMg5nTPPgL
wx/V75VcmmBtj4tw42SwD/cyPFwOsOiNpenXvmLlqhkIBIHTlekaD2nwVI6V
7W/rphG3/oyZ5vu6Dz+NnnC5bvexjUukzCM+ZXOum73tn3A/LjooPXnrw7Ll
9+jfmxB4Ltq48Bhiy8uy+m2YYjexyPOS2Thft7imBbkDaBgm2sMTdjlVTUI5
gYb44bMVN3zD90IZLuEBBbTybVrmyONNExT3Zx858OxuMah3/JGJImXK346A
AyaDfWNgeQE6TUZlYj3aUv7wB+niG8bwP2px+r8opDZc5ZZDLLEJBpZMaC7X
is5cLl+S4/xdU/ogM5K/sd7bj8DqSwqgH2EDPIs5fRSXVPMe8H8NfS+ez6NA
4h+QzomisrCrwVo8UtEIPdypApmJFdwkpkwGkcq81x5cjOkDCgRrWRmidotq
xZ7zLsPcd0uZTK54+eB7jho61O5sDW4vY3VrDllQKYKxM/CI53DZ+3m9ZrPY
dgOWrIBIs2p7Q00rxC8/t4UbmqV6JUi/4nKkU87/zPwu9KhXqOuzF9fmG8/o
+vuF/nXXbDjJVoM+CkLDTymvA0q1W6/HS7V8jhiZ3OdmEmCrC/at525qBwdm
hksEfxeEcKKeSIxR5TzzqpbRiAt31m6fvynzHD8GU50O1olcPHifdC9m0GQt
4aZVs4RPhQoUxgoXbdekIntVraACuHMjoSiqWhvIG90hsmu/ZARQ79/7ount
D+MgpWJAoQWx5Gq8S2rPgVRZfia1ZNIamNMZgA4i9rwuBbWuUGYm1htwUOoY
YydW9g7Mcdk4GFTSCQMrwxRIQ3F3M06gRT1y5OOuvekv2Xl8rWtMJMA+2/vv
V946Vo/3t2P/zhB8IbXRM43qq5njnihsRVkRdGXHDtwjw+Bhhr4eu7e4Sq+G
oQvlnGRj5yaogTVeLzlDIw+rnuKoSaaOnn3jIQHh6izPkLd7sIt7ww/qWoQU
TttbR8JZ6wulqJJwMXnQwFN2539dXsOrGtki00Lvv7IF3iCgH5A1pTkEtCmu
iIzDbu8lh9MMBPWtbvt5zyyctoAZMnIXE5mc6WAeBEam5ByUiarkWATPNExB
4mU+G7WtYB3uUkKogDIiU/a7xyEhy5iR6oMocEeq9lg87+O9zVxCvlrM2Clt
QUJy+X4OX10hzkYHlOCo52srIcPllXPt05WM0SkFL2zN88kknrp+s0anvzoK
6WMyGNvZCeSWbQEntIaV/BK7wy4I+8ZCxuAyuIASoA27HcUnB7lFrXQZ93FK
WNcY2CNYIYxOfyqn3YnyE7bDvdf61PdvQA4MBZSYU2bsHxoZHUaXM4o8w7F9
SualSRvLPA8irAV2mQm4tq3NMHoRF7hCrxFzFZ956RfYDHEQuhNmVwj6LIts
k7NZpdcs7qZZ+Xrk6QSFDonO9BMsvqABbkABm/1QExPW89zv4L/B1mKIjjuF
W2D07BGEWjgDbzHsjy2baq3CHvgGSHtcQ54VS8ErG3cfl+0ryhgjSZiZ5Lyv
y46HJOviqnrDHBz4TDzNxvmuc5b7Zs5zjQF/UdxbgIilnfrV0jhwnpRXK6Eb
DlUN/bqG0ulfY434HBD7e7H0YseMGYMi4npJm0VyX14YUkVfvtqTm9hVzCMT
xnB05CnA7V63mgFQvH9ZSxWn9a4VU2vi+ae+BovOXyJp7R5HBZILYtPeN5ph
44xu8HlkXE7WvxFzwUrkKSFwOBcWmHWUlqv2whkc6EQSXjiMtoc1YFDczTin
8s9eN0x+N+WXvNxphXHHh1HgABcmnpgfNfyjUqMZbL+ziUUU5Lk7VMOYV8A3
mEWGUjAAHPWnD8ZxGo9BpT4fREEhRp0kkqh3OYeD8YHK8VPxGjBvD3SSoZsm
ZhATj/BLaHHg87ukRGPDOemrezlkgbGcJUyxOVa2Dg7JG0l948GtFk2Rs/Mn
sVo2oPaFtS/nH7M8XyY7UwzAkpDFgatVvdz8LEAAMIdCmIM2VT9jruB3KzIm
0U43SnXB6d16ijs7CI8TfjtJ8hF0pVpY3lsLl9d2yjDh+ngxNV6ywPe1Ec4g
8WgCJ/27Rt2M6wwdnoWRwdT9L3PUMA8jgRug07lTY0nWc5huwEY4FcWJL8jx
BaJRzpfXx/AzaF87PP2TUnUhqqoE+NuGYdM+ogHmsb2xQO4pv2zh2p9HsG77
t9CfvyRmKTKpOLcqBiaV5Xu/5TVzwFYlQE8LLoSOVXBFYnHxHbKkKwggAW8z
szx9ANddy4L7mSN4p3K6YkBjEvsb1pINKZ+mOx90xodr71eiFLORSUyS3WRT
hZuvDnyPVp4PnCkHqjWOwU4Wve4RhuHSw/uZUG29dn7OQyYqrEJ80mhfImWh
amlYOSn57nhV3m9NofcS2csd9uFHQV7Nd8ZT27ABHItkeMuC7+h9PBf/h5Ey
QTCTUmzMN4Do0BQWUDJhMIiHmpHzKv3CwZJlUPlxkah8I9AekidmOyWYCMUP
Xss8n7hkT2s2eMYfv/rXjZxH6+WUt+lg/9KQ+fG/zOfn1xrZCqC/jnz+OFXU
jTLhTh0IjKvIVzycoR159Rf6o8AHuJdpQeXzFQb+XrtfqpYEfcC/JJ7k8n/u
4zMtVjOaWF8Fy7KQQ/+hxsBPZmypkDpE7YDVLR0f+j/67ZVElxywDRT0zP98
o1Hzom9arYzPZeBoPmksq1oEGnec6MH4T+XagTlS/eEDrOTRGLpHNGhQZfT9
5R6hw3y4fFZmSSKAL7GARrTi0KOdiX1pXUTl6utcquu+mqn5HSW4po6uAIrw
XAznz2RFAFWUtTAAXycEUx6OxxTqAkOxNueGo+Of16r3QaInWnzEmA1JmFQl
gNU3YyLWEVotOSsT/hUpS0HP4enE4sTMMyb8kf1f+PuQyKAGzAnOYA4DJ9RA
PmVXWhuQAh2USCF5brH/U0LL0X8xCnKHSGu0JbHgDH3WBLjayGlhwGhqzY6J
yTXu/s9tTgmYDD4WTMEyTZo+TBr/Q2oTkqo2tDqfcj9daV8/3BaZ5g2PdSX5
HPTufn9MYX99RyYelJRSoBKYbp0ilWA3ukCLsTiE7ZX2eZeH+TctMa7qmRD7
DeLxHgj4Wy2SsZwDFtxFYj7qQQskBAcENzcqSK8FB6qJgvQnitv8tEyhxu9j
GDDow4VOfRNcMQj36ruVpP5bgkueu1z5S7pwT5vAvOxVOUTzY5Y+USKIPxPj
MDD13sf1Nn7Efg/1hhU65JCgiSWZV2/NImQvTu2ExZTALkYxLaoG/VNQt+bP
Vx3MUiNutj7HC17u+lFc0bvNsT+ig4DduYvOvRic4FmgoJRvko9e6LwMwPl2
f9khI/pAf1Ih0KMBMeOq9qe41jf60WhHWZfgBKVZtwKYfYPmtYl8lEncax8N
X0vgZum0uXFlRPhE9FxaD5/SX5/K0CYLiSmr2RkLwK9u6sBVG6DEbGRUF1A6
W4ypS0QKcjLI0Dv08CoXWvxIwab+pA9BPAAlqah+NwUa1pWkUOqIw9eEJ0n4
ZxZlhrH92PYtF/ZIVdC83PYOolVAFTUZqzdAkGc9Hd+3cZ26yzCVtAR3AsaA
qE8CAtY9wmmVB75C4sUYYnRFsxEgY5Yy8VSablfQtmnDPYqQFu517V0Y8YK5
yRj8qyt7e+GxT0nDDuwz6v+d5jEpUrdDIu7l2WCu7/NYlhBsgwAg8Q0SVxVC
xRFiE1n3ZQmIhim+FDhm72WtKXNjrRG9FMUAsEXEiYjO1aZ1p2kwz5LJe/Uy
UMwQHeSmx5HXGx+VihbK7q0YfgZGPI1ZCO5SOIwA5z2q480pf+uT49gmYub2
0ptO00yU/lfF6ZwYWbKSJ797XVHiqie6hsJ5uVHUs7fePRMYH/nS1wuDBAuf
yrLTkKxCNG9fLv9LKHMAx7Wk5jvkXYoEDlWI+fjbKAzQXh+Q/qjKAxlnIc4k
eLzwNHAO9cxr7QNAymOIbCbs19wWnMgUwUwi20l+w3h1/ecjFWc2IZTZcJzC
EdQNkjGr4yjXnOH9vZsm2adR/HJjmst7/X7DPHYN0du2NXeyP1zo0dWUXrAP
2z7moXOyYXsq6dwDOE1qBwbmSJ93KTqc3f6RfjeqRaUvsHRGdYax7iPbh8RU
dmE7ikvdBXiRMF/UzAqEl5LF2/huwxMjmJzh31cmP1MDNqC+Fb4U8xgBVu/L
JJYbW0XsTQWCkaLJgnJidMXxqKOf1OlC2ezizebGm20qG5ZNUdzPIsW5RJBb
8ou8ep8hD0Ue887STF+dz11APNkoBYkZMCXCTgwc30SIGEMC64EJ/gPZ00z4
lFJLvaiYlXfF4O9kr/VV8iWdJkIWnISyUJLLIqEy+ZRLcGAp24yNppRqH8KR
rK6CWeogd2Xztnf2EDI9pH7Xo5Ypzy3mbWn9HHz96mMQXnqpS+a2yPKFTf9r
oTLsU6z0R+m04CXQ+of6S0RMkSANMH5xl9bmVUCSXdzJLh1y5HTnyUpfwQTe
xpG5QgrovDMZC58VGvV0cpEYaHTNBY0PKtUCgz0ixKaBITRTAvCBg35IzRsq
Ym2OY05JI9lxcDjxoqP2EMQYT27ssjLvS+59bl8fTPTT7J/oS/SHmP/jXavG
IRvSJ7szhVe82eys8W6Tf2wM1ej3XT9OjGMEDoZiee8j1aPtJCmL3drwdB7u
waJbZEhpOKYHbJbvdaYWZPOqtheLlWdXt3jwPCWf9D1hf+QP/TSLeB2Nvu1I
+C/JfBiWvT1JtwnU2GnDtDzirCUwREQvHNXG3cnvVQm21pk5bqWZQl1S0s7J
RJmqSwsgAzW6SYmgGYyi3jD4HYSWagq475PjTVTX7CodYMIADJ0UBB3XE9aQ
11Im4JoezlGBuvp+Dwxn1LA3Rx4WqedON1fWFNbZb4wvOrh8WFFQSS9cCAJM
/O+/xQQvbUEvlseclNGbaOxxVkOzQNPKmZ6euVhmLrkBSYC+ez+Pj6TaWXiG
w/gZql5NzJp2jGBEVU8vWA3XfzJzj+PvngxvEBQA5n8VOSKUeW8EU7NggReC
TGgo0BDJMBw8h0qOkH5Fm1AXqMxXY1q21Ywwsw9kPMT8u3wH6hMhcDk2a8Sz
Gfd+1oSjohcSeX6Qj4iruxWb/+EZrR/KAhRJqk5kuvIFKYEgQ6njCC1smEzs
B8De4nBTP1OtK9/iWXXrOwWa4jnbCLNexRfLduA0RK1Rc4JIjOw1ZjO+Nn1d
W6s4xCquk8zcJpKKz9U09Z/eTGxgWvNIiWc39Go1CSUbA15bS9Mg6fVVyYKg
wZfsgXGcdjRzWtD4+Cwrrjo5S/xBIUnf8CSRzlnepLHS+NrSixasj+V+345u
chCrKIZcnAinLgbUg4ylBrahTGJColkgKydsZPV2Nnyb8+DrNH+1ew3TuX/3
yaKItaKrhewNfLa+sCbsRVP/sYvm06xcqperoswFXDYG7JpilitR9d8gY8Xm
iq4jULLUO5xr6GiCshGgfqSBHByGarXs290u/+mBlZHuskcwfYOybS05f4Z8
iQnyMwU44Omj3NR0kLz4sE+UC7tfe5zUxNwHSfc58PqQubNxIDx1ev0pJAiC
zGxKk2Y+dZb/KP4b36x942uwDpP1P3iixK/DpmKvD8wfA/u0bzO2ceyUeHKo
7RJ4ePb/wys+VuLlGbj+hIRhakgPiZ8v4kKWgJ3qqN9QNTDPShToWs6R+2kU
T1pjXmHcAS5zP/J+6l93E3vrBsqO2QCNQgQGGnoiN9Sm/YIHwMzpCXoKWtl6
MqBMZV6tlgl5eYP8dH6aABubp/rZqDifGgaIu/xmPazjNAjIU58o8gvdlJo9
BAuYEJK/aZtQoWUaPxskotDxydQr3MwKjmgaI2TyP6H9/RqS/+35R6VbgB7X
VOnxGnK9UcjRpCe6swh0YcsiAE1tRO9m94eBwuivVeXJIOAOaapjaShvzT8A
Ya62VtfPHTyJ58Q34MulPEiO+MecyWxjlggEQebUp1VdfQao2sE7e0Vf2aDS
nkz6q8KcV4aMPXfGFPkVi+SbUZ7ZhlU7dKo0ejjmZn9Krru4ee+5fcMzmsHJ
nYX9GByyRJxG24oTbb4f9MIuPJVKwJ2NY4OM7LRKCMjdApR4A9cnGJg6SSx4
o4DwevRKpxMQqWgGQcJtG3bx0OsUBwDaHup4Ym2WmSzbXznK0HSVFlymOaPy
xiVqfqQ+rpKso7aEQzOj80kt6wjvIfJ6yj2f2obBWk2TllV9sJ0Bw5GhridY
YA/fDtM0spemgJaBaSlvY6iWYnRXh0/eIRo/9nI34Se6d1/B0pJaD3oA4j7I
4Ji17x4y4qs0g2VYUdaxCRPjgSiAaevBJY0kn4GEmTX44MTPxGvkEQDT3f7g
04hdJyuGiP3ICN9ySaBjoqfozpZ2Ir2cB4szwGyPixrLqV+KqNA+Z7NC9BYP
rJ7WGw0Wl7bPJPbcSm3hC0jwj/yyyh/dX9dYqw0GX2le0/pGTBPllCGmwiWv
P8h5cmvkXnF0jF3IPhhlxtlwMwmkUXJUlCT/BF7478DUxkzW7Ov2Jj5nG6Kb
WRGVf8AtR39gURc2fraLltc6RwX+KF+CPpM1bgwa6wiyW3n0doo5EmrKUFP/
uUQE6YKo1nuZt7L8n3zlmpEvYj6547kb/YcRKAvPNcTtwWdAllGnpypQSPw4
Qp9oLRFNXdQvTU3+Y0AmsdDMNbVQoCu6T36xOSk6nJSucMhv/v6ZqPBWzXqt
gq7HceNtyShcyikrlUbgxllO6g7XFI3D2M4aMfAf3jSkJhPXbkrSSs1dFxsn
nFrzlWBJfu7SCqCRGMCKWwyppc17ardncPjjk2WplgoTcpmLr/Brccdyl0n9
M4nVJk2yBPJ1BVWGkpmH/nZN6u9dozbfz104TnVD/nLgDkxLvvPgrxbOv2dj
vcgLjZgM/ndvOnSEfejJatMxVXrEGhm/vo1Tb7oPf3RxIKK5KGEimT3UqEq9
g4gAlvyfUxnaUBieMjW9tvedA7mJXbPF3WInYLkLKd3noYu2rUK6i1MngYrm
Cc4z5Ze8OASr+7NJP3rN51n+Xq5+P+NoEklGXiMYdjahfK1pFpocllrP8Rci
MaNyTkEGIWrCnL9luIuKs8bSYuZmO7vz1lE/aGH9FPziSUKFiNK3dCEW0AER
n/KTUitiKYSqNGcIQlnjd5S+xXVyoKAwbfkqHLjFKoBwnTYJL0dVrweTCa2H
qOuoIjqVJ55ZBHQCBkV2n0L5a4qIvoTHBWpK5y/ZSxz1DNri/6aRWz3PUGzq
vvXOEMDE/B8vENZY4uShSSlVDnZA7RnkbhicqIIfwJDdZHVgOf0dBKCJznwK
oLfuT9VCvK9p29K06EcVsKPIHOnxdrvNNANeXXnI3A1JrMkh3sRzjQXJ5PXD
D4zAN4moMf1JgzdSxLfGGoH9SKm+FWFZgLt8rAq4cD6VuJwyG8q7Q7op5SWu
dZkzg9evPAyRfK5P0GdptQLhz4Z6IZtBEp8muWDj0ukve5eNllVdd1LX9Kdg
U07HDCe66av8z1ogO1rVgDAUv1TTleiAvN90p+Ui2PHKfa1r4yn0+vaumMn9
CTwzN2CMORwtlKyRJ8egC97YmlEFLhqTm/OjX9KnRjiT9Yn67Y0NVlVVZnZD
FumQAZBPSc0qqe2s98QSm0T3a/aB9eBYf3OtRGIOzhUUg/Z7VPdvLexVAORS
Hq9xuS5TNaldazXSMbLXvQ/SzXLRhAs6ER435Fe+Nv5dnCdLqXf5740kRCie
BlhidhBgFAQ7dzOOf6kUxI+ij4gPDc95wPovzjifoSg+B6p5pgylVNPK07un
2eCXG+Mtbr42fGzF4jKTEAFmEcg9wd4bV2QjdhYp37Gh/5UWly5azo02mKcc
LsMeOUQAINPZ/gpm+pV0SmY8b8E2yyG68SZxeSOoJX2dZQYx5+X4iKQ2bsiY
cd7cXiMT0h3KNXjSB3c7zj+FhKk9jI87RGtZNMxu218fE8gRcZDLdu13CM0e
YTBJeKNM+rhNHqlbTSj7B2xN9R0Mu/FzUN12eWiuFjFJZOFgOL5jIsNFEEg0
fVwA+MihjYNZRHgH2Zdrc2KyC9550VxCecaseRo24N2EDiuKA0ydPQp+FIQP
xoAjae4GYuQDYJiz2MlW974YyFgx+LOLHbGNp0EKWVx8HIb0LDOhQgeJtSSH
stzxzYa0qXwDDTZ0tzk9l5WUg8oIWmyjwDPGSPF8D58ZHuohxWW9nSFbGpYd
+yg4ApwvswGiQ7KHOtOuT7901CZZXSI7Kvcz74kGI7iTccP4dnQHRWyRk9lQ
0kjUAGHh4L94SmpBxrpMSZvPIk+JK24/AT0SBOX6xiskhZYrR/3gnFPNo32x
beQyeUwQ29a3VKZaK2zlvyF0DRR2ykWMpdfzIGYVINpy8dDYjZT2wR7vssCz
8pAafKDXULi4aJjgDT+u5rpYaEHG6UV0+mYgzr02f3IfdaWz9gMxAhb26cNi
gEsHuOFx1ngfscBoH/fzqwLsf0nLm+ejE5BpP5rkNJaCzdvfS+6WmXGWj2dn
Dhj7MbqFdIVdsZAlAuK3cZvRzah2look70zEeWH1d2UXBB55n+FiaPPcbxpD
Yu0fLyLrBj1iEK1ClNaA2ytFIWn5GulD5yfDoE5YzR0YMomH6FF9/54bmlo1
QPaV2STg0nOoJyfsJRyxp87NrCSfmTmRlmato66KiBAltspBhAzWXGm88675
jVG04B2WAcO7a1F9Oo1/fo5PNKxhDW3gYhu2WAQQ4KOIgZz+QQOPJxB/HcJa
jFK9zpXfXYCGQIYyMDZeHEIcfkVoLBzlqZ4OM7kq2K/oGzZ4J4mnFn6c6Dno
JAmWTL46LH2rc7bawT76TG213lhRbJqjmnrcPr9uwIBjaHQhHHL6DSlwVqjH
qOV0SQ9Tiqqv7mplk4w4em8OeTh43noGJdl1R2QbYHzqlA1Wke2RlEgavhTw
1tZH3t/gvknPPC9sOlTACwcA6o5TMtvw4nO0G/mIvqz9nfIfcX4FKoYhqu7S
OTjA4/hvfeEI8L1txL3ngMZg7/VkOACuUIRDT3o0s118Fjc3FcKHXVt2LcPp
7YlcpWqsDtX+YABptWgsA24J45yZ2KjzxicNzyDfqXELg2ULPspzYxmxTwg/
d3klFSHjZLiqWTwlprM8olzt6gUjCOrdae1CzSPsEqrMRZ6oxFxokW9Sm8oK
LQcLT3H9eoTxuFhnPRJJc/d58L4tOYF8HJpWgE80hHYOxvvAdC6lbLCuWWqw
PfUsgbxVnmlApcXPd52t7gHxnPjTlavWcWs624/6X7VW4myYw/5aMF4gJcJg
Am1aBNEgpbJASxx+aftl1d8BegiidUbIeGGpsAwNWQoiWDDTtpm+FxB+NJhB
hcCEAGSqgGapC4xGqgIVduIPP23ucQM01PZup7hdJQ4fC0DxXsEoaUimauIZ
Yc1+tw3eka+4jWUTZ4tKCUT08lTVPXoac1EPjq0NJeSR1rfImI459W+w0z5l
emayZDpx38ua+anBLZ0SJ9lyxV28hqcVomTSI2NlHIt8zwc2OOXSdWk3znFW
6wf2orY83IMOx79mGdztnwlC/OMHYgEYZ27l7vqdENxY486YChuG69mlbF5x
dQHNwa9IzmF3HrceQdbvBWZAl5FqcuzjjIovomNE+avrddUu2YSMlpkiIofG
zGgggOaZgk8zCdf1KD/WHQvQrSYgs2nZ6Kbj1sOAfbRTChkFQR2k671JdDCl
lz3tstxBEbU9bWDFI/2FEHp9d49GUFZ/T+WZcn70lk8x6xdeIE+UvlIXSSYr
nghr7ID+HTFSzyyzz/tNMtJiC8VpvcuhQbg+zuNH7/S8iLGflSlFQ6TFMKVn
+sOA9DMwhesXs2MzVT45KG8+I1LEkRZ0H8pVByFjt8uF3d3j7sl3IeS6S4tY
82jY/6FYcetDHeOojXOtAB4DCJd9KhkLDZAQailYuecr0G+7enLyQOlpz7Z4
PE4oEaMC4mPfBBv5NFZrOdqC5XKClm3pipWSSPwULJ1TbfQNag5kAJAIyDIP
Liu8eWSEuadZs4L4Z6VRi1ordBEz+8j6ymdr2jKEUyl3TTXmdI2l7Cny5ANN
Tu3Y2SGWJuFp+SLVLBJe6MyIpcnPCtCyEXFKXLKh1VysaJT2QIkqf/7L+pHU
oISvF2nFEHK3PiafkVQGM/C3byu9qolTQhUICrGGIh1LN7lVeGKiw+C5msYe
5mPQMjCdei1v0AIEtAwXx5O8ecSUEQBaQXeB6IvPgh8+fBvWBDDCHicZjwD9
QLJKZOXPfnBxYm/lhM48WicjfpXJwWZApCbh0GCHaYEx4IOOl8m5ZoBTBOPw
RrVc8//6diV7CqOM3zpnOC5D0m5veGE1YR8YnJVwmMJBq8G43G4Hu2SWcmvB
qIl34xPAcrqwxbcGfDhy/mjsilQnR8Y9E30uHreYduwpgimzD86UkrBb5anf
zEmNBq2FrI4TF9ctpmf0E12XVRvLF5StGeiBs1w4ggoKrG2zHpwGTzMl8y4U
VYHf8/xxeRvvp6XOGAZcwR0SbCIuNIv+A6OpXvpYs7ou51b3VHwHnW5a4uxb
O/9JRsyEBUJTo6uVCt1tvRXEkC/g6qKDU3bnfI0vvKVzLcewED36+leEMZSL
nSYktXjV1wf1hXK3RpDA5cFPjCPVBTaLrIXU/jimzHuk+eXxPTLJm5DqElXg
M748OIol05fBlvxA9MysEK2D15IS3FtZv3zLWuNmKMXrm+KLHEfy3BXluHsa
jvt7G5f+zZrZEIPkREXjiEAHtXTHLnP6O9ozX+pOCA+q3Dx8jUOy/KZrV5l0
ocJtxpOYIZ5NE8bIXiPwSRiGgx3ck4rWft8NReuefTCcVMRoOm/spyOyBlrp
vncRGC3NPJF0DqO0n8s2KYAs3o00hMIiK2XiitvbFCb8Yx/pYGngfOXSgvy7
i6zEz5nyTXZnFf20PQxhcY5fY7O3aLbBhyYOmRFuKi6PD8giqlg1iQijKaae
If3yHmFStFboYCE1Zu9VLzol91gvK3m5SN477tdzBONAY5Nu2gwxoumNZ+xJ
piPkLU4JiD2q1pSO4YL9M3qQQgLeJmff13CyuNX+BCZPAu7bwv9w+ICVE9He
6EXasPTCUEastd/YV2WNyqb0TTFrBijOL27sFBjXhlaQZJr9mibN8hV3kfqG
QbVoF6RrJY7/0IUR/Z7aywwHs7Ehs8oWciwsdkP6yfl+WMcVB5C/9iMNjXzg
DJftEMTDYF5XmuvUxucVqXNUZfmvs8D7idWKLjycH9fEoGtgvDjs3huc6SzP
EtUtpQoWkOMHMmi/Ypah24TQE4/o/CMSQ7huB3jjGTHvqkkTfRK4k55Ajco7
9f2qlcUkJsC/1aOVOweJcjP+dY8CAhL8xYfU1rkiCF9lWDabh/cY0j2BRSLp
i5lhM2jc3+ufDokk3L4OLHZiJnwttY1UIsUUOJbzdXZOGkO+YGdsdl4GbTtj
w3fJiMjdsAhxSjw2JdUbe7+nlVe6k5iBR2z6nUS39X5Xv2qLJurW2AExstAo
J5NGEMjfa947sN9OExfICd9hRbKhov+azHLzwmFf58JXnHkH9ImUAUhLsnH2
qj79oU0AtzPYnSHHVL8cnCusd3Lv2E6ZHC2+sNUm1vRTjLP4kAZT83u4gr6v
caeneJltRt0D292Q92cc53NYJ77mnusfxXZ1EgH7HAEsi8tFghAANXJQL6r0
dSP7Kt3lWKW7T9o7tFelfszv8z4VLousFwAdNY4Y2ZH4wLa/wLtQ17wcLbpM
Cuc39Jj+XaXuT91vAsaw+ms+MgJQzKwiX3iI6m5sxGTfLcxFaR8unssZEg/G
ONOW/qox09oJvMfCakeS/ASAW9avZPD0RNdp6bcXqr3sOuzLy5x2To/Nq3Li
2zCi0Dg5DSSCk7TZkaKzoakP5svfP5OBsWXwYfl0oVU+bfrAR45Hd+PSddb+
AUvQaCmGPpVYDonnvCtwZ9I+WllERdK3LJZpxkLhawPDp+NIHBgy5fShETpP
FIJ7QFMPw1W1Do5Pb/OBg0ixtp7p3V1Ng90c5sAEUHq7csaTO1XmrWXk724H
OcsXlg6kqVEZhTVSvOoNNELajVE4NU7/sVQYdRkCAF4TLy8a3HqDJD4KngiG
wTWWfMTPEIHux77KNhHIXSn1v/4kBDHYpWAoueNEzIewTQIolYeKHbPnqbPA
Xgp62QQLx1xZsTwzM0Xqr1MSD9IWziEb7ExGzCIyGReTnLDUD7m2gxnJZx7z
8x9IM/V1ICxLUMJYzEUOJNfnKL6d0dL3XC1MLayzSZ1+i84LenVxHRXxq1TY
HRyEvedkSrmI3jVj30+Nsgjq35OsgC3VEcZC2c8geuOT3PTo0XPEpsL4KLus
DJ7FGgVEieGtvUCjBb8PTR/dqFG9rmQOGSYo1m+jC5JlbPmutzirbIgm+JHl
myV+NT9SkLJ4Cf2+yHCgk0l8H5V5fflfe9+hEC4ZwKbmI73K1ua3EOKy8b8J
J3DvWGoLxEa9zeOxfdOrymwp51pAxJKq5Wqf8+YRyDQErgRauHc133IeTmIi
4BMcO5V9RFbJS+uBrS+T1tcusY9PjnFI4ZS6yOFpGWNk1GZksfns+//0PQX4
hnHSlIizi7BReKObmKFFFqhLXWpd3RIEdwb7DzRAWQ+kuXT69SsPER1Cni94
5sr/nJWj6Q+mczHLZpnxleAjf36OSQo0O24/c8al+sZUx0DAcHDlSxyn4A+6
pszK3td55TG9JJTw5AnfkFSIHvitQ98irbNTWKtzqHR7/da1+DoLZH2VLBBZ
agIU5yln058KtrMgz4QF0WMDPmtlrgOhjaQ0fBhrV7c4rAhoYrEhm8Kye2+1
9YksN/OQSEaVU2EzROEaIP3bgVLBA+j7WS4ex/e60A4BCvUfd4MzHGxS4WRl
5slVmKjaZUni9NeKuUrG3QqPNhhcVUUXRXnypOaUU9m1gSfgy6ubKseu82cz
zk7EAidnehHu7tG99wfYyEKe2/d8gMl/qI406mqiMQy20otewoTgZKEOGECW
Ayz+Sq6YT0EWRq+XpO9zgo1L+s1XpK91ZVDuK4LlOqTr6ur2pNm9EdXjhZ90
YzpBVnX+IoYoa6eK26rfNjrhLxjlnQhHybVMQHBw/sWoTGxBFEaIBEekPzxl
8Dwf+mpClFoJr36ii89owP+Bvaf5w3HV5LL0rRgrVaqkiBshdu0M6hnL0608
KO5zsPYwVGiZivIavVNkmO+uUVu1a0iYmcYwUo12xxbfEOBQ5+gUXNkaDdYW
xVy0GNTgbS2dhkK/sFHYfh1MYR2DenQGg9ruTlQLvnq02boCuI7k6eZBWpcp
NEV4vF1Y2BPPt+BZCeR/5MJxg+2CJ94Dwt8axD+a0QIgF14tdg9PbXL5kdAI
hEO7vuXYE0oSLMwJp2Gn0i5idzBGG5AMZO6UYowxZdP+SvvUJe9ZvciQdxRW
2Y9oS3DWtpqXGkOU9F5BjbWgRD/4ZIXlIrbuFDZ+3isK8z0tjWcaNiZJRbE0
jibAQ84UprolxHC192wONEeBq0HM8HYEGp4UD+mhPMyXSJ/PeyzfOaFTHXdU
B4MJYEDeV4Z7E11RurL5uHTSa2Ti0ORhz63wewWLcNjOPA6P7R5/Rpcr36R3
hDafwTAMvpXzxLxn8aKMc2TUpjlYJMV/IIM/vMNFibkB94o5Zt9iIxmWjplD
xQkVr3PEYoG4H9TUknAfagTk0b3p2n8ytsuNGatlwQc0bbnpULKHWkERY4Pc
a3xuRzOm82tuHqXaMXVOzUAKjLIudgf4AXGOv4xOJWRvqkUmSs051HJC4fzE
/TdIeJsaWPdECj9eyuzV3RVcvRKLLBNlLrna1iCABnKOac+rUN6p0cULE7cG
/EiaRjGYE7HQ2yEPCa/NvDGfejSmTgljG0LUxV3A9ORoW+IH0+JqxLKh60nD
SlrdU15EUvB8cQyP/ukezyH7R5oQMIUmoExhFk50kPtpoA6Bmjt1SuvktfHK
5PYANMdjjv7SsUt89BUeXrnX5WUHpNe0LD1wvBkqXU2LEoINeJpshAfGvcnd
XPrHRPBU2iZNM3DLm34S+TJEJiVNDo6ID2mQqegZc4rc33wEmpw8T67YnUi3
/jBBKpi9e/gMgdaA8Jj5jOuPAKfkvXVxOVWLGUlOSvRUJ1YhlcPha2x0ZQ2L
dr5IvK/rcxrFe8PcbQ2MTmfeUSD8G2xJHSaFOPOXuenJrw3wEA3XqFn3eKq3
NUvkC0rAy8mYIWc7AYXWD49iSBVy2MrxEPCKmKiE8XqkDFiKQqtuHcChw0nD
VWbxUXVhhKgw4B9tVIt1zMvfdL3Fou6cl8+LB28/a74X3b4++f0ZD7ugLDfz
x/3KPXTNn96fi0GTdxJiT7hzdNgGBCKZ3Gm4LYAFII+K7c1vIgLORnO5Yg6l
V1h3V3CivmcWb+kGuBjB6hLGMsGwkWeLgA771exaLVteH79ENNtIYI9cEzMJ
DWLReWm75vZgeabIXHmNy5bcuiHwfeixhOtarSjoRhMFqnBDocGO9xlwyiTN
az4EIGrYLy6y58snj61/Swf30GjAt05TlX0hXj9nBKywHHbNqaweu3h/eFYg
A8f81sJud/VggG9lPSPT92iTdztRwq0T868Q04jDmhdnuRDq/vIin0KWdWb+
0WJEctbh9XMqQtHQCqpwkRWA3cN8fCHXPvWSez4gypFrv/eo8s4hbN+q59QY
Oix/+L5nEbblV41uYdDj4mn4rEB2fxemgLfUfDIybg00Or7xm+MR/QykzwDo
ePRYWduTL58dUC95Q1VVelbLiZPbSCw9Ujv7iRmDsmveUPISM10mquXlKzin
3e8gADnKXadGhyJ0bkXBhAtS7fXbjnkXosGeL/jeYYNx1ogYCDxZmDUOjtzc
DEuwdFNtgiSKEyINLEvRyB+UTnpyYHuuBNURXAMBaDWgLnYwyH13LEU+fg/N
+FjfZoJ0ZYY6Z7s5Hgv2HsBXtnm2s2zPitg5stozmcL8nE0O1PusYxa+LlCk
ouTfIVeAiZm4JxKHNVJ+CTrRxSsG6dL+FP7mEfa48cjuFCUuclLifBEGyJZj
mW06ythDzqeZY0OEY+9ZQGcuEtF+riB6qLNS/RkWnLOfj9IplLWai9J4IvJ4
+Rjxo/R4sY887KIGcPCxfapDEkEcnjDANUlnrwSrxuG+WhwFi2bD8kCZkZ6U
VVcSKcF6cQBUBmt88tSP5tatNe7DyemHIRggO3OGLx0o3O+rxyk0G//7ID6O
L4CwIHulv0CgJ9OAsbHDHnKwTXnwg4OnL1zW8zP/Xv6KESo0Mn8rTttyOOwt
mrRFQH/iwYRrbRfZ3XYxWcANzzNG1AazmKmO/vd9fIYnPoWaPjgfNtiXNv67
JewRCSNd2dtmgRNLDFwP5rnoMDK+gyyMRCec/mM3n+Sncwz08ZEMqrHYeakN
Ha2nIppgL7p9xKiS7Y8tCiIClfaOi/baT9g8vCxVwrTKufLcCK4A06F6JMDu
1IUXu6F9UwlXtFMO08PgGH9kx0Kh21K6ij+SVvK0JeTMTgvuL2rcdsTseggg
dg2qz/yTpYQrCKpx1LmtqzUSw4bYt9ZFHRzeamiXB95YWIt4ibMSfzHtELut
LSG8qpyL7YaEvdXFlLlVYOS35Rz7g4iD/ZMki9dQUH1hcNV96yLkcHzuS4Un
TPbK/hU+i/sNpg8CzQspL5zw4iJD7F8s2b91h3fBt8UGiMQYlhGt2k4aLICf
i+oAMPfaD+Mqwmv1bud1U8OrgnyLlZPqHxmO1DSeT6ZIVIC+bLQ3XeRDpB7h
u2ZsrYGkbultQkSjSyngI7IBce5AZDgSsJ5Bi7X5Xz227ecy+beqNjA8cPRX
hG3dahWFjRtjen4931uVloaE/DW1a8m2B10ThjGNInNRr5+w/94Rke2c2WNA
WQ2MHLHeDYzoJDBASHhd2CFHu/BhMpSt5MS6hFysLT6t1nWnC5u+bLMEIqTj
KwnU7CLLdZAkgTXoc0N65xmn//5U2fQVPfkdrkWg+VCGwAinb29TIdjCULtN
SAMo0+DhJB/lDmzv4ayZx3VPl5ZLDy3pahbBMokIxDKdHQyUufQ/2OeGLAsJ
2/0wHUW9uv9LyginfXoE1fVjqWR4s9Fd5XScIlemLjsMSZQn0xyIfw0Asqvn
lIba9OYnFPaKUsdVxBVe9Fh8TZ14TxCMyu0l3zQl4aiv+9wxq6XSJh+vmje0
HGHClX09+SYhGmY+CxqCh+LMGgMI75el6Oteqr/qcAomD4HUqYDJh9yoXnA/
9JERPNwAuA0WCNWooWSWgcBjFAMB+sGkXFBJEkWXun4yjDwK/VEMeksqEeBh
zzvjseiSzEU08Q1hKFK0HYWIkWDrdkNk1NBnMsDAueYCMPpaEWwKbHw20+As
6d/WbOnziRAT51DTS4jV0G+pIaXW1PI8HIVvvyi67AWQNRnlEFZ98LOj9AyG
/KHqW24rVnF+yoy3RrHGhrzmsMythG0bNhDWRR3WnqCP0WEigQ7LU0KnCYYA
eEXDHbzEfSqw+dnUpDIBLg05b7tmabZ4ywLtVMO/nWFov0ZhvO1qMGSTpfrj
vM5TWqsqNbgMrsGL3bLm3J+XkkX9B5TlkzlLb+0TxHMahYVy17l9WUgBblmz
mEKUCtn6z/5z5uQsbM7+BJdvfgvsmcUzAlpifNurs2MdocLXqX6PdPx5id9S
uG48AeLBpGXTd2KL4RmyRt2o3cDy5WJ/Y+dJJ3PPT8RefvxPXM+K0kw/wilC
iBpebcS1VS2Wmq68MQImwUv4orhcDub3qy7cnRlwuTP97cP9uYVekIdUtK3u
paiFN/0Fx67tdQ+u3iVpMJvNGFJeCqpF2IpEe3ZKfPcM4IGRSXDQYxLpITaB
L/OqfisDXMZfAuSE9BxjMOHgWeKqD+txESUeubhZl378mnCUatDKZa2M5Mkl
Zi8xxUgcLsg/E21dRtpgj6+ThCoN8DV+pNb+V1A6NqfWwjSmS/NVw/5usHL8
9aYlOZLVLSrMSjq5eUw7it/SiI9lF74V2snXWU1pf3P17mWDBJzYw+fFvIZm
1SN3g9+QwcXs2UVf7d7kY6osOcRsJiK/AA9+GK6m75Y19zymbzfn8nplywxN
A5sPucd7d6vzERkoJTppU0tzKao+K08mksPJ1tAWvJKznZbajkuiIrOWA07x
FUg84vJp3FZVOL4idFi+vIGMni5khDbiGbNfmkzMjy1FZyZQDMI6l7r+YNKT
4QXuC6n7RKGJ9QsjREYbrWoAJATNLfgNz+GlSWwCvU30x6u7Wfbcb0kr3qLE
RAecrels+M6AQ922vdJ51eekDvhJ92l6n61RByDbBMr7nkf1pFLu2gZnueQv
R98UJmsF3KRe0ydUSe/BnxjW6TjEhLVI7ukBqZhoQHZjvHnV+oafpwaG1R1G
Vzaxn9Y6ZPmZWnhS3OLZW54MWkFBLO9ZBWfYrOBi5iQjJwsqXxRUQ4OMs1q1
GP/PQ+P81S25HHUvEuoK2eye8bthMbVbFSvuw+R4bSa9yswcksZvrpY7si/N
fB/N5E3H+pYRgkJaEYQsxq0rSso/hl9YtZ8PuiMB3PBCOcn+tN2F37Luxcv3
BVL5q7DJxMpxf3N+sLK+dTFpRj3WI7kW7ozCm0zKfgpfCgAyX+J+17YbSLFu
mOFnB7tDRuKUT8I71h9tzIEnLaD1I6mJEKECmYlDJjr4zh1t4IggvdlCnBDI
vYQhnEN6eg8hqPr+4Qo0UxOyQ/pqjJ+UaPMnW5HBiPKHWyE7ffBX7D1Dg8yI
hmjV/1WPQfhb53ihtTlFiTDe8OKMjm7vN0oPpdUEX23Gj7IEXjaUGXUWvMpq
7A4hbfqyisorNvBCxkNhMKm25GiN5plYEK1AAaPFOfTHBalDBeotQv2VgZum
Yp4LnQ6z/d26te/fXkWldufgw2ZT7UnRXaTZBs35dU1ZNd/JHKatp/Ft6jrY
PfY0+hCQLp/HTc4q246qjfyJFmzSJqY7GXxy6+mb2PxDZIKrGo7eT7axNjC/
9rJVWE14XnJmots3SbprOlWOHknL1yP8H6PwaizmbLdZsRwLeNbEohLKYTeb
Ea+b8Ge9n/TjscGtkyDkeSnJ/+dGne4hbiPUojv2kWz6yWJD0Rwu55juBoiV
7AkBtY/ZZV6U7fXE0mezjLmQw3y+QZ4xa539OYY474xFmFnF/gMBmW7qgEZ5
XJvtoipVmQCZOyl6PV6JVLXRfEUcXvHwJ39T+3nSl7AEAdD0kovSo78R/vAL
k32XSaHSQxJeNfEAOOypA7eOVLrY5wfNyfw+TxuEsuIz03oNgRp2CBOYgbPZ
sWYOa60JSAhRnOJK2hDUH7fqfEd4SV5AkAn1PsCoPAiBSP68V1QYWpnmOB+G
iBLWEFSTFE8rbTTmzIB8Lv8VuyHb386AWw8YC9YsfEpEuBImEPL9uLDnughZ
5pnepjGuw0hdHLIyHhcXolBo4QXweMhw/1ObIY6tnl+GCfg0HMcnrvOpR/cS
9acDGopDJdMdZB62+EUSjQfqLOeWMhIyeonqBZb40IYVrXShrtZqCgsLOzH8
eZawHV6GxAteGrLIL32E7UDc+borr6PXisQoDtHzJggC4drd7QZ9mdVVNUzD
EPKRvKKaGNUWnWbiT4MPe4EmB4KqGJxBx9S9/P8NYchGsRVFpLSLJYVxVEGU
Itw45F37MI3fzZa3ugzRkP8dSOYvitxGFqk5G7/BXj3JNfF0Sr9hIFWBlbqX
LYhnZ+N3s0Qn9fHQ5Xx9P91fSmEd6flb3UW1DkwiJswgH8Ub86pWBHHEBbIJ
FAW1O+op6ZFMvvXyLu6ru73UZXaFyKfrhWCgt1lbSKTgazSRH1Nfwyge4MNh
FdLWM3DN9sqP5EGf0iY9eAsnJ3wJGUq5piuGDXXa5Hrn6cQoobCt+rnP+5HU
QRu+8UXZcdIk4WJZ+PPzJgVDO6XuwJ6b8O4pnGLgBiVZ/w4HICVQf6LQXd2x
0pT+IWW5kCS/LEY3/w3oi/hB5t8dMwF4qvdHl4FGrlWEp1Cyo041C/prn/OD
QBF6/nXvvD0KhecSCj833Yqu9p8DfhUmZlampwPBwnT7dsRl8v1sB81BkEGW
r+VUQOeGmBt/xfV7gFkbP0aTcTAdD3NwFw9UpEadhMq/fJXj/C9thtG1kTUP
eBX7VEI0mfS0N57m/jxqDw2MxOnPEFQYorZo2ESpmlGv7+3zI+sjt/afaK2L
MxY68t4AgfG3hGJQhaxisiHxXT+oVEoo/YHQcCju/TY5Mjgaap6706VAnjsJ
iqLL4nO9HeLW2W+FcPDrUrEIxEVMdJG80ef6ljaAJcM0w1SZ0YwaIjMwOYVL
2x0+opO5Lrn4r4jXiuN+D3gKwXdLftYmnXx6CZ1rKvbSZ7ssKgn8+IUsG8se
4mTmfxE33+ucW01y5/T6D0FftYPKljY3qfN8M1tbkukhupBFXczqRtWJLtbA
298mbxfOCyLXSYube9qiyxixKMdweMoLJSmU3J1tOQu3bJdld5ZuG/h1YD3o
fnxERhDSSAFBu1YnGwacSciQGq/pVN69QXaxtSULQa49aXnr3VYWPwqEti6+
2BjmwGGfFV5fWxWKHMSFLl7B8xZm7dPRMSvwyLBpYy0wd48oVxdtNEBIQYNC
/BEHx6e8zb2yssgDcNeuFVjCr79NiWGhgujs5rH0oXmja4QV804UC4xXY6Me
Piw5ftcPsciiDRePr/4oGhECOxSJtfxOpUWySsBoAJEDVJz8ttvLsKrnPLqK
iaxLRMNdJH0/cFoV1hzNEX8IbFHyHgrlXZM/YQhXRubx7ryXwMZnqlfsTahV
p1mjSn+o6YIMJql0MYsJi2aBr9FeD3qxf/KktnmDjPIqZlRskPNpfBy1235V
PUD/En2Ttea7yeqrVg0PzoEgaQAPHDWyiZDCriHlRa8xdJy1a4aJjWv+wc7L
hOR81bMzA7Dcx6WX97hRY/1sVGvGEpjeIlOrkr9dpXfzIYKO2aXYjqRPprzN
7Wm48XxKbbEVGDEzY1AVjmNE53E6VkZuRa6irt9CRtsPfRY6FeZrMLIPUZdG
/5TdiHepMI6vArXCT8nGCHPPGFGEUgZktjiSlyLJYxPsYyKBHB7YjueR4q+D
048SN5jCRxTFFEg4UeYMw5P39phdgZ26HnGzwxIOCg9bswv6fdKSgX20uV+g
gWrnEW+G7ObughGYIA2e6KfpGH92/fDRmfqfM4qxXCBM8D9G7aUyEKPkhL3S
sA77sPEGGoxtQEDIMOjxbJ8rJplvl9Nwudb3sSelZ0/6P9iS6S0oDiIOvJBG
Oavi48X/tZUtKz84dqKF1bWku7MjGAePpU6pHJsTu0EBA2cA7bCW4NBCbcWG
+eG+JaqJVGVA7clm3faEFkVcB0NTK77ZjWyPX998ZeMD2gCtrRL57p07HPbU
evPyyTZV3sdLlzRNOQcf35j+s4f8lC9UkAR3qMtb5OPytqRd/t20xUPPtKQE
79Kzhkof9J12mVPwJEW2vX0ZgWTbz0GkdnK+X0IBtJ1jostxhN9dDGLOnQ/8
4iH9IDeF4wGmw0ulTslvLByQrTX4mqTXCbpXL2QWkF0P5oy97JVAzQNWxxU+
xLJ2XNchyXyYYcEVP8abnZ2gYZqBy06OXLam0QYFgYAIRJApreYKWpzx1pYQ
z+K3PCjRVmyxXu3EH172aQYZ8u8QYn00Bj8OLOanhALufsLmv7NacsdX4BCh
fgpVVPYcbBI/lRFPuN5BQs/e18JCRbGPOkWNdACyvevaFV0yHVmK4wZ93UkL
wKgmeZ53ZSYrXhsTM/9X2HjOxgDhZ8Yuc3GxdOLDLXeYKvfHKHA84q4v5zam
bowaHptSTgXCIIjFn9Cewzyp1n9rO+REQt/3FwVzITQXUWKPJFYnrNuuU4U0
obzt5M9BeBZbQaarKgAldL9zmt3GLpMXanz2sAosq6+Exnqe09bJ4CcqQIfb
7Kqqh5Rn/47UySnByb2/hGg29zAqiQmX4EAL9FejwzW2brW2LFIWm/i90Z+/
I8iEfk5OpFyriIJW1nz7pdfyuy/i+806G87vmsj29jt59ag+2sKEKww5+oKO
J2P8pxDSzxcGfhUICfJjmZ3jlyjZ+fCfCHGrL+qgsKhxHdiJujxk850/OBXk
UaQXd012izDiHgeGFYMxv/Cx8pxAOglkqKGsbCvXa1ZXggCNJaCLoTO9XMd9
jTlDoT6Kc+CnOdnPelYE5pFb3IKm/d98PEIXVufeG4HpzLY0VXNFbFAKAG1f
cSctFoT7aoVzubJdh0fTKYvSx9htvvYcajvOFbt/Lndu2PsoOO1qtx9locVn
OOrom4TXXhPA7Jf8TjhUEHmxwjhd3CX4MRVkgsjTWwWC5+YUwZ6OhyKgTzq3
09iZPnY3DxoCSyVgBXTXKPhBuzCJ4/04Qnuds00ZEJNASMljp+b4hOIbr37l
ASDEZpEfSlApMt6iZktOM1FMOkAuvPfKUF48B/tr5wL7CEtGHwHyrAeAMsvv
EmS199hCBUhffaYa7kzbChOkSrGns4BcFRwXD2q9jr52sHp3h9TGZ9vnrrsM
benoUQqTB2IWipsELHcuCqJL59g4gwIsg/glSsm7BV2Y/S10CIO9rNt40l0S
PctzyWOaghLp6uaqwbw982nr3CCyPJfq4OfIlaHzfelfWE9A2hA9fRhPeHFz
rrTi/Eq9gJtkveu8kb0kVyL951zVZfgp7F1Frf7lbglwXH6lGR5clJdeNhys
kyN8rOv0+9pvGSW1JvEyyFQw4ZTrxjnWPAGeUL/SoLwXFGXWqw3mYIrchvoj
qunicJqJNHHf/aGrCzh9u5aghk7J+5npar+uZVHJlQCMySrdShc5ixdFjF/+
MHPQ5l1e88E+uHWC2t7Qt4mQ+rjvOcS9bBzlATYGb0B8fMYbYIRUO9WHH4bq
Plv60F/Am3BMoPMD7pNJG3vwQftxcRt/Ip3Ad1Op1QLkictVM7I0lSbN1FB4
G7lf4KLvk4cdWSOpOg8SobpufDbJJdS8gfj0NRjpFm8T8tQQXiptYYtbeY1R
kDOi3Cr3w4jBZ8xdftAHUeD2eEC6CL4Iscz7GtV1pPVHRijn2M/L8AMN05uz
8bX1vlKuTG1V17HGKc33V2AfRR+RCMWrQDRBdttADHtnww5OThkB03vJ0ywU
Bpr1TrV1AG8naYAdLlwr01/4Juol2E6pVJvwo32i7yFn0YpcjvRM84RzuSkK
mCRoMzbHYdCNtQgIYXCCSi6EgGz80HS6f7ZtZwAFC7k0/+ltNdf1vVtOh3RC
9LlpIjiHLFarddWHYQm4h6ZlfAgfdJqN4feeng7Z8M+r3vvqrUQteKP9o4Es
IqdxjUQytSu56jT4pkDZC7DOXvP9uhc6sPYMzHM/emw57P6KQuPTxH65gWHU
gk9T7oZPJT5qyZ+h8IZ5bWiXncJc/tKBbEVxwhRAFi5zzedfEnYUkoeRTqcI
UZtH1zZif+0NiFb4Cdy9HlerNbIDalUajY0lybkTy3p+56bWV4uyvB2pOpMi
Dy3CZ9vwbWy3bCrr9nFcMUxDHy5O/wMLCozcFF56NYbLI9yoGtRgo50VNKog
ca/gHB+XRr5FOV4feD4ZAKYiWG81qUC915JRc2ifUdlSovkaixvrJMX8DZG9
MgPg6tO9hKtE6ux2jVIzkHg5tBkSitMwNdlrP+zOiT1kgzX0cJEKBIKzmDgh
Xvs0WZB5oi1Ztw140goczvwTcq9VBV+vKt7QRPQETJoy+j0OtR1xgiGtnObW
MGb3DWoDTn8N3MBAed7VjB8oZeSVCSsUnuF0QgKw+md/J0wI9DN60DggbkCU
sqK94fy0gE4diwpP+/XwZL+RYY/ykuJTv5Qx1hqWwKn9bh9ayPhNA7XsMm+i
Qn/x5caRL3r3/sXS/Ai2Xv69z4BqF3F+RDhdQtOQDllViX+YtxDAMG6pJOWD
F7JUCJlVbXj+OvlpdtETbgaGKwpjqA626frEWhUp4Z3upbbO9Vbf0sdOsBcS
wFN6gc2GuP3ozZv70GGdTbxnI4bwROR4xmKqKeWaPsEhucg6I8YJ4OmSxIDt
ii15rQWaM4jwY+AYEEyk7OjvroJUz1AhF195tEScJgRTZNAlzE7GIBC71BqC
jmGt3SoOkPNZjOC16nEnLBvLUIaKFMta9XEzd/UvKgLEHh0cIzZV1fvpBuD+
erY0C6Z7/ZKLykGzVXg2eMlYUuOAKzeolD9H9isVNqKQ0rimeC4Q66WK0ASm
cMf0/djZyj+GAE4bwDJbRgsubZ/oqG7Lt2lzaTxR0ubTT5EqLDCB9/cxslD1
kQuBfQozAoM6xeoKPxkE/MbqFlWGcG5PpHTghGfcjIXqag4T8hREX5Bgm7Y3
hZOxLE9tZbL/QTRrr2/RTtGLVqFbDvKnsSqnoJaM9O8MxKeKenY45oPfTYCS
a/No+e/OuX+SWBZlBVcvR7dvCWSHEwiAmzt6Xo+LN5h8w9ujrGafnCyZ7OaI
2cRSKnaGsgDfqL05qG+bb5nlBZbGypph/ogttjjLsGrhxQg7oAFdSO4/+Qu/
g5u5dii2octDVn14RWzSmj/ooiQyPUs9XrXTeVVzR9lK9n5iAbLMiaoeT89G
RnDtTGDfNglZIiz4Qr7dLNxqGD00R42uK/eHY1n+AVpNIeA19za8UXm+4X6v
DLMvu4MFmOfRq5yNDnsfBZsvE4Qu0KijnbFTTle6eIgcCI9EE+BOu2MjrNRf
BwNfJAZRYLb+zNkdTInghY4BOroniHdMp1vnZ/YHoSqMTbLujYEUTiOgHR2s
64AvKjkw9JH6Jp3T7/yNgi/3ZoYg+NJzmoR3Ri8yL6nHmhA+pfovU2XmJeSj
e49tZXZ1EhYyimhTU2Yp2w3+aqLqZpFEN2hq8mPzmFHxuwxh7Bmfl5QTzG1P
FR0JJm9WoPsD0nOexhaRe27PiCKZxf9LwKPavyBOJBeNT4DaRqguVDXagXXz
XDaXwXj+NWxmN3ZIoY8SaKGo0Wi6B5xdzSv9q/4SQrGbVgZHrFEmcK7qUQmp
za3Z0dpJKNNQJ6yTL7MMyJOc6R7RMsVICNc8sgNRRIIMc+K/FrOlQfSQmg+y
UY7GAD0Hz4iA1nyhVHq3ceCyePyfxGxAP7bHzI6g/kL1xXzxRlfA6V+MNTB5
3azR1c6oWDASmMd+FHx2L8MPDl1gLQj8t2IxpuwBBjZzVtbtgQD4XKsUzrru
+GI4XvKGyoPOREwrLaQW5tSXD0wVPm6u0DBuNTGAfV6bD9IuBoaVE6r4apRV
LmQDzD9nukuvWalC9JhKir8uZq0yQLuA/4miZ4E8f+KWk0q/q2IE4QS5vCUw
1A9VeGsZIWcVhYd7FjmP/rzGmEAV5qmbzpixMHpLQH+2RgHx3LFrT+xGh6ri
BC3WaSdZEl0UQcyATiElaEptRLzBfrlrwpzPDoabfA/qVU79W4HLb3GaEOLm
i8VwbpffxR6CT0R/hA1CBHw/3rGMk8wWewDnPhRu+XjXOYq1a3sYkWopGeVe
60uzbqivAzB5sz1MK3VDfTEy9qvLDcU8fr1LUnX6BwWezyz+JxYxX+Y+y+Jo
xOziWfzOrsAsRrnLzyeVxv3oxRsv5Cx6+7lZmjCsmFTTnbQ0p7jftFTWHX+4
D26zK5WRG7nm5T4qNcUS5m7ljyP91u3NcGMZluznBrBpVYcx3sJLnFUysDK6
868rn9EDPUXmOX0OKqG3WBK6q7d7MCgrP6f91afd3sG7RpaF4EGyC4t7eqo3
t5FOHItlxe3pyiDROjavLGeGUUuMI9NyTgXIRJyzuEkyy7Erg7HE03VdALQ3
ZDeKsxA7pH+mY6oZH1wdjgiu4GUxY+K6Hymi92ld5l2luFacYbgG949CbUqt
s2Gyal4nGgRKjTxasQxO4W1xtrBU/X+LKzOqfiE9x+Bkv0tCKZ07aHlDQM85
RwluiAhGuEVXvlPiIw4QZwEPqXjyq3UiArCWH0VG31hwgk5priUulhUyftyM
Q0Y1yu4beVCiuzY4/8HbVC3HbVDp7gsKLgh3AzMNcmkWqrxaLXapjvNhI/JL
A29eMSh3p/3vVNZQHc35opPPFaIKjb2ay1RcNAl5fTKs7DxMBr6YOsfvdJM/
fcOn4kHdgP/LeSBeRka5q/oEj1D+pFOH6aAKCSVlKwaCnPkZ3VHtRckiw6kq
4OBfdgirPUUXnhg1vRCbwNIcbmKc7N7qgMQ9AXa50wflRQR5fpIFzcLBTeZW
uRaqjVQPpYXNnrcYLpDEkUaM71UZtJ5PPNJAL8jf3MLXrqDkB0aeG9NFiGFJ
d+yYyptpRA5TB9Po8MGoaW6lRfNtmnEP9W6vUk/BTkkiF3McF0sQiA61RkeD
+EOiwBLemdGKTJfZkOL+BACGnRAGtv4tXkGxBdwGPD/xRarEPV1eLfM5mQmm
9OccfyCkUfgFSO1wtqDhA+7I/FblwjYcmrn370VDWQzaJt+5qVMaPb5Y4txU
DmWWuHsJEfXcdDrsFag8BkC2IufjfFjYsCO2cB5M5C/rFGp18xWvPB+ndeui
G/kQA0zy4l7tj+qhc5BjTXWwapp1T9BundV63K+j/SA3JH6QSbi36CkuT7lu
LG/dY2D8KgpeDhN0tNt9iYMs8hlGkqcU9BpnOCilBpp9UddXnNXDOQMZHFJm
uMi+9Rz9EXglowCq8K2Llk7yHpLRzvfkQJTGlp0wVnRiFWzKe8IcsoQzCgGe
UoQtuhGhdPGYlDl2vXg44SsmLU5J9BkMVpT/ij7JJ1FlrpBkCwt+JZYIcOVc
q3gjV7RoyL/yYam3Cbo0Ns63NzSlVI/7NCglX/kO83JT/sdqTEei/PunNrKg
3QGSRmy04JzVemM4ByHVbMLcx3nIm6aUsRAnuPZGwl0buVHXkQXQ2GPCFSrG
gCTZ3B3tHcZ3F32rWVDHmmM84XK+rmxly+wUbP/e6yus1Kmka54UH6m+vvSn
0xZvDGI+H6Wr0KVedW/dGYT9rB7B2pGAfzHmOTkLqEMnwhogNtXnzSgOHocU
7pTk2LdNUWSj+VLS04d3ZhZz96w3d2D/rFmy4ohw1g9/D4/yZYTdnw54mK5S
3sMbJVV38n4GKV10kzULO9Zz10jogEuiqpZHoPHgimTvXyxRS6psOKY/29Cw
6CWmszT2IaC3XOnMpMw3c35Bq+5iQc5oaWr3JkyrW2XXu8acMRgJfvbkLBc0
EL6wsrk1KsyBW9hBb6B8aPHU/2nraHDorsnY269hFYcBGwpNTIJEzI8WX7yo
EH+RhVGg/XByNhttVubxmauRRY1vGAKL4KT3gkrjNprTCLXU1d5u5f8MkJ8y
NljfI+koAU1GCevMqVYBEKoz+DF3DJpfiaY6Vxd+Id6q8XuYbC4RztBKmmhy
6tVZiG3Cl2V24Oq6OIHU7enPFjOD1wwfJWU2SxFU8yQSnf/CGBONOa+MzpHD
E63QkH6xdvzl0sQSm1wYKpzP1GwYKlrA8k/2aEhW4HfS3KFh8Ef2vuIV4EFG
RrV+9Z9a8mRN1U+oem6LJW2YUR0SDdrZDjYAO4fhx4sxYXHYWnux5rRSrRxt
FNMfc2ewmJ6DOGXtZkJIrzWir4CuLrqskbydLuJ2FfLP5/m967SsULurrQnj
JpxIZCfaJ8Y7VATs5fNyJ916rEadlEcxpUpsY/ssIRU26s5sQ4nHWQyPJpQQ
SU9ixZKUyGhxlmrXdiYFyLhpBIvvOGygWsdhTGT8NRUjmYYjmKQpw3uFn0M6
/vGGg5F6zVmDubGnJTCU1HeuA9fHa2JCuNMGzFGIO+WYTcrU1tbGtIR4G/1w
loIjGvybbnTtDFD1GWDidBrTjHDW7WQnmOUUMfv9gAgEEfvSIzJ6YovNBCSX
Qu7CdXwYYBgK6uGGfqscuS/h7asWFvLST3BTcJhFWjTAVkCNUOiJmLUNt56U
OLoGIzWVA5MP0Bsz+9DWrfpI3kxO6TYTHanfthsbG3lWSSoC9c0np/PggGFF
ElKzJiizZHUrOvFKwW1n5QmTmEB/HodiIixL61NXp+IpE3S7zzM7UiiuQRHD
oa45EXtzQz9vKaoSeC/UDO61AW1acD5PRFKxM9QqnwLKVpZ/PnPxLJCSvAtq
KwatwPJCrqRIC1jUO3mdftjjavgXANFD4f9wQOTzcmiTKODspMOhP4ElqYJ+
zb3JF7QeDsAOFAgLHtTfhMpMsPg/1CGj9kyKnwnym0o54L/Fg3tFXi+eHxJc
kzNEkQrIXDPHZLGXQNvTImbber+UgJaRJZ+sau4A+3QxBbrYE9MoTsd+HZW4
0eJIiBOAbkIim7caaVcKbKndTwWrkZb0tVifkrqjK2ucBppFjDVgyLVHLmrn
TNuip5+5XUcr+vI+tcGfX+m/zuRcCCrTOgZoFDCGKT2/RgcSPYHVhTLofk2k
USKGU2ctjN0/hjyyORq5WMAgAAD0GEaF1c8Gow/cThV7gDqSUE9js/W5YDYZ
Jl/4m8Olq+yI4NCHfNhdYeNnaq0R1dpiFvpwIZ6sS0ih/snvIRh8Vg6i52Wy
lOcAxiQ7n14WBXyMvWQ2Zi0RvzJbv1xZl4m3E5CAXT1LaalfWwsyyJsl2Os7
ogruceO1QSNzA/DCn6ipJI33XA2NMSNA0gGTQWRl82QXZ8S3WfIfMo94UN2h
Z+0qHWzp1M1ndCIeB3nqZgFmbgBBBuQZalGHr8bBwxB459YvY7ID5s4PqoTK
xov7J5sfqZnx6fFBCFawgvkAJ68seDT5D1FvQKFTZedKLPeTkH1shYuu+0Xx
kcAYsegIndRecARlnSD48N8ZcIBg5RmrZGf6QOWwq1AQnRxIA4km7eJchnnv
3LVLw29mOeFLtMarTVYd8yMdPX/EJaF+L1WCjvIzm5FyDMYsppn06zThp00w
mf0LgETIKYUHYxbEnnYfxOfdVFWq6S8g2GQ46tygMrmpnyDk5bMSRAJCFqQg
cU+UpOCmFsMuxWwCDHSJ4Jjoa4ccYc5Vk8jxEfRt6rp4dOUSsqPQJ8ymvDyN
SeU5LClxA4C9kLksGZ0jgsgFAbr5CcNCSRsIa6khvKWchqqhyS+fr5i3Ajwq
t72C4CcKdo1PRkKXXNcbcnMutgmf38VyyeqiAGRp7ULtjy6YOzPyi6HVH52D
dzublwFykZyGpCON/D1ZVuBqsEcZvWCEGkpZkpZ/hkuYntiO4em1GNZ/SbCr
2bmRy1ybB2mugCm4ObI4fIRSgNioX0Uv0wmml6e7601ut8xscM0wHTgXwzeM
41k+/SMOLZj56905p8YJ63nPULxKXmbGJ8FlpTF7WnvjoXW+bMcVXmR0YqPB
f+mjkNDTOfQPp7U53S0u1k4JRT+qiIfkHRRD689ofq/Feb4VDCeyzA8smg8w
/qPbpW6bNqgKBn93sMbh7JJAmfCNcKdwCO41DJl5hPH+z5XvUPOssLHvnQm4
3mabfNFFDVwaHIg+4aYB9+zqJBDtbMEIPKDnadsP2Opg73tVuv2gJ/NNuP+f
j6POsvcGj7dSF7t/wXtsBL+JQcVdaLECz0c58FSVmFL3Q83oT9GSqsaS2XpT
S3YZtivPelxJbre8b33EHwLOHfHM1oWhk1OD7Mu/lO0u+Fu0Hi0crkCN0NC9
odLT4XdZ8snhUaH1/l2X5vSKuvdKSou2NdCkSR/w84+n6z3pOfgCf9/UlrqD
3hnkidaCJRf07fGkIdGfe9+8gchhuRwLBdTTTMZTfyREiuBPWD/rrW3J0ts8
fb3+fwvqE4voK9k59X9Xg9XdjnU1/IxOoxo6U7CAOGm8Dy+wg/LzeZy6FLpZ
VVw755gtBARWFikysCivGZJGD+Qu07IVrnamSh0Un1BSjtbHgwNKasvGHOIY
LV3j1isRZ6cxChkBgm3dd+wmjUJZ5ewnlLo2dypxAREF+uLhsJfhZFxfaBjg
b5b+X7G7XtGYJeQqVpvNpsfBFnq+RiiByq2chBfskePPdgn2W601bcmwQj1e
ms4TgdTpZqJxYHX0XYj3jwYfz69OxZ7iqHAw5I3EaGnNaIJWRYb8fiFW1Guy
+wN/JFov/11Tffb7HVnDQqxAzubhdkIQZeilb+ZFGSRn8zGX17Fbdr7luA5X
5/TmYU80bDQdhWna9cx6iGzCQNsBuc44eAVoPUXLO3Xtbbl1utn93oNl22AE
wkApnpD1B3+JPVmEt3H9xhIibOxT1BUWyTxEanT78PyRfIBSX83GkFrC4j8N
uQ87GwOzohyJIvUrMWedjKVjQhqyxrnQLEsdR628SM7b/aUWDJfQ9MA+n2gZ
AiUDgZEhcxK6e7GxycyTE2CoEmx/74D8NS5Y8TfnRNH4fmAAazQvp4vgXJJH
W/fY4g1kzHge/jdgmXC4ywmSnjp5Sn1Y1+jVSyMeVu6heanc3KRDOUuuBtN4
5OTvv+ivEE8N/1owkHgnMoBrvzCUnw/kcvhVhcmFIQQrlnjRjR2R9mvC4/ou
qwJ3RAPu3RL3jxqm75LlHGaTzV05CKCi+n1EBhAuVyG5piqWn+nDeJ45Ut3o
g/KZzYHa/qsnZs25FZ9qvKpZ3oCTnR8BLRGGAJGOYqPvmcM+OH2JR9PVIWS4
TxeWCyNc0kxqC8rZpz17PPaQSyI48ch9BwvLC8Wv9QNgTfBnWHwoC8PujOE+
2EKNB0eA2DW3j98RUCw3kuhhpSFXislibKjPwivtY4nxLbr1oq7UlbqT6jMj
OIjwY8i44EYz7o2ht2gotKCesNwzD/+4mrWQjDmO+0VNXMu4CwCIo/q4W3/C
m92T/vG2D7m/G/TFnXvwjhLdf0rGgukVq4Ny64tsPw9vNuuyPZ4FJmbUAsoK
W1GDQwd7xglvQpuh9j1ht9csLh6s3Z9aXEXh6uUkAhyYXQC3cdvNVKErlFqj
JI72vC6wqnFqDBROU4bkcseut4PcD4Yc6inligKtehoI+iwsVT25L8QZgU4/
+N/g17uo3HwxKKTEpNc3+a+qeEIYWHTXyLJFLXibDwVWuSwzJqsonT4c89hF
pEGAwLEDJJoZD5QC+Mei9MksH0S3rTlG30ezRu0WgyZ8Xewmb0Fbz74oxTTv
f7fXSKLJlcMutAN9TKO34tsRVrNpBtwY2DefwCYenLLwElxUg90juNx2C6vZ
XOJbgb5DSvwKUu6BODqJ7JhIp6eWzD0//NwqhI+z/uoAnycMWboA843MOQJZ
/eEQnjvFh8N4rpoir98gISIm+1hB5BicCqy0f0RBosv8OfgizMBqnBasz2cH
HKqVl8QCGBo0CNP8xN8YXv6M3XF6wnJVCZBa8HKIsaOdlPcVgndZlAwnv/xq
CLjqBomqHH9ICaXcB3yv+eYeRPQDylrNIuowk8a7q2dG4HCfH8O/EisMIlrn
xfeVcZiYvQ4qgZGTgRB3eu1ZABUeqWQXzAkeVLPt99R2h9wR4NdN8w95JeCS
4MHOPHMyumDOo4D0m2UMmV93/qL+d1RI+/mTMkgt5N4PfzYiWjgVnjtG8by4
1q6FwbJL49OmYHowfy1faWG1EiD+tlNUovLfGBZM/IXajhWSOY9C3jMM1arm
Ij/5t9nNmYkvLUjc80e+fE3pimOiGIw4auCA5AubY1q3YlEKRhvdVt1vgG7C
WKDQrhqYfeH9iXmRhuIYnbGcDQgWW0yottM3QTlFfIzWZ1/XdcJyAaaQswzp
mvzECpcD3HDosnOspY2IeiiCvaxUapUeUb7P/T961mbfKjXvlePRW5FVow3O
Vyi9b0GrB8L9+ezMP5ZSDSrb+EnzE5smlvHAFEfU764r3v6PaLCsSx7FKopE
NjH6NOx8N2b514p8KC6vAUoiCOnRlMb90KMd4bRfbw3jJ7yOPATvLCisqY3f
ZQ1nOz4ekeANzGHxwN10c6b5n3vdI6n0DysGBNGawGh5siSaGfCOm1zM/L4A
/lGiWlP/ahdOhNw+nZJhVzUg2VaQ1QfjTyXQlKLCxJmJjCY3QmcUbxbIWhOT
Gj/dphWDXNlqt/60HevrSb4p+1OcPq/+tsUcN32980zR6am2AUI+/Lkeuy/H
kgWyGpVODHer8wvAibPYbs9Ovi+cvWTzV/TYGUptu8xF9HkHDmTcfSe8Ozf8
midtJSRlcAbBfuwDiNfs+t8IcjJcm19QLEjIN+gOfwMRpdb6KecKAFIE2J2T
l5DXWyy8dUWCkCdYcMrgHfhWk4yRgQZEWuHvyGZ9xid7H0N6YeWwUMpQXtJq
fvYLSJ7va/8lLXM//tMDkp1YFxmbTrN9Decr1jaKOJZSsUP/Pd8Wc/S6UQPd
nyfBa8g0sPAV9rlnamsoUP6eIvfan+iDSFMQa0hfLgfzeCe3hy0Pwzghopdq
9YPyNz+kEwH2U6O5gYO50WdCnDbc+Vlb4BZhPkSJLy9nSFnrA2jM5zOpVsW2
ESvM2lcM7sEdAAXP2zGGkwLbUHyAeitSQLgaEF/aqr/1uJHR3A17kcM47v9j
nfewG8zH6LYZYsXKAtjkrrXE4FtPY14scYbNV6FlKhVu5j1E9390PsvlHLpB
fciPMkNe+uU2kYSAVelOQJ4Eyzl+mgEFedDuC3NLp7/3WzzIIK/TzQOUxo9N
H+FK00gT6ERKs6mxMB22Up0MCfj6wm5ZU6/GOkm0+bgTVV3Fs2xgLy0ZVMO2
RrytO7t15z4OqGZFzXpuy+bhdd6f5MN950a3juJVjUlDzVx5OUmXqVL4p92o
EYgAGSVhaSKTnGOXTmf8jLm3lt89Q43G/rTF26usxghSu3w/Gfx3bw7OR28z
Sv/lWl85JK10s0l72Q/2WKb3lAQmdFJHm6fXO24lp90KDXPoM6HJ7gwhkTmg
TOBmHxmnR3SO4bxn1JFSUmAB/4u2T5SkKUeDkxn/SWVc3AoKKCzTqqtJHL8W
Lg+WNooqK/3JjWWToYRdil9eITEJVwXBTAVg8RMGEYaqvTgVWmWL6mMvtJgC
PHtHGQxlwduw0zmG78FkbYQoLHqggAk/JMDNIj5XGy/6dAzDqdf6PLF8s1wn
LNKVQF+bmIceq4d/FWv8Isff1qZOoiChK9+Ibb+/0JRYQvcD4VBDofJZa+il
JCmqvEa4TclFLOvyKT1nTMhWDukciQJNthhSo16eCYJtPrjRdmlHOQTkNnMd
cG2Xoi4XfOBLEkGRBN66Cz6k3oatYLhuuKSZk18LGeCByd+zOZJU5XYhNW1y
1+ufeJMH3THBnbSAC1rJAYaJaoq6JAr9o0FG7WKvyFmejf4CzWjM+9YaqHd0
y2wxQTQLY9qY2oJ/wLyailOBchqM1SHmkN4k+B5CWaSBjD3Zx15iwiWQ70cj
Mh5D8uAnc2bRxbfDI1sS1//VHv8Y4R63bn9fAlPsC3o6fH0Gqanu1I1HqMoB
ionuf9CpW0I7wdYjDDLRSnJy4wqOoVyIVA1xUn8UrKQLd5wFTXhwCrucFatm
6pJIBiXx7VhYE2oyVn8DLpK8Li2PX3G6GD32NnDkVlyUqwOP0wUemN4lbTYi
HScF4RSfkfItJBgpyZp89xjkP/+v0X2S5BukyY6WbVEHSrsv8oheZ2uQ7wm5
y/HnMRJpUl6Vxl/z/MCw/jWf/GgHi3C/oe7AkmpRf3mEuHXfuRtXduEPpGu3
3Rob2/F+tOobmDVGZhrp8jO7UlTs2MVfvf7xoH0hzwjIYqa0oa/LWiEnqAH1
KtSRr93FlOGeoTis6DSv/RQVkiW6YBQwPcyorOR14iM3TayA5dMjSPFgfeif
+d0Wb8TYALGZfl2tDxRVnKwKI1PWVyhebtdFne15XpmXPmmvI6udAVPSJjqE
sdLOiR4XPW5ClKH6VR/Zd6BHJdKIVfTxDxb6wydQZHsx1s0hAdhaNdUzLOpc
L+yCYcp91RkjSlt9GlMzyuGvqWjr7AaPd4Fdoo/u3QEZU0m3VRauFbqKu/Hb
er9DgCglfoYk01NP157d9r6RCT3V3cXyUBPRxDFW7vZN2urn5uVPfG8Thrz2
ltcT0Dgc1vjMBEgHLLzMcTvJU7G4z4KuL+jYqav1vQtUdJWx2HmDURuh3EVd
E/5o8UYL+RgRrOaZJbERe63xHs58ojNJi/uX4OCqn3GNsra27AbfEdsOKq1B
JYTMYcWPoc2SIUTqlzcgdXhzi8J09SzHFMYjhabboFRYmIK0veBa9ubEQEtc
Lg6yW5B8TOCcylwBszsO6Sov9rcuwR1GbLGQ2vtopwchIyFvG1JkwWSKW3SV
EU8oqumcukwyoQQlONXeQP3/j6UfaoAjk5vKTcvqc10TO82mh3Gcbx13ia33
5BFbVyXYZVYhEE+pePPMSEkHeWFB1b3sTG/YKz80TAhlG3HEIqpmKUgVlQGr
1WtwkjaVFNkrLnmIv8ZiBvWZnpexKSSJdaOo+WbfyoDwYiOQu+1Bg6iuztAo
dtzbp03JKKsi7kh6H9UQa5d/ofhy13fyaOWqzQP5bwrO3tXq6+CY9UPjXnCg
nOxqVKTX7toK32YBGXfiiGr38PGQIZ4fQDi+x+kv3bIYKP/CBNs1m3uGKPbn
I4qrD4/+aZ4zLrC46tBWmj+8FSa7sevVbe4z13prLigbGfTrNtpQftmAUUlB
JgDCQVv/C7+Amk/bTDvF3YWU9SIcc8+H2pKGCiJEK3SUQ8vAfRASiVOjuPVd
h7dGkm2+5KhuVgk/cMpBzJxoT2EYbQooFWuMkF2rT/aJ9SYzj5n7WU7KSmBh
AWko+1m+dKQ7ZA9V+tH0emBuEO+rXjq6fEmNsOz7RgY9ei3apVgqn+YGj6I4
qIIwlqSljzM+eO8OFvqUZMS6015Tg6ngaJW2ToJJZn/bOQasgNcm5DlS1vHO
H3b9Ez1/AOkag468D+9DWnlC7Y2dnITxwlZltsjqVpl5U3oT9ivUPfNEd3cu
TpRH7Xn25YTTPSMgW9PudxrUcqUSn9MiCzfNhxgpjIjGlFtfzYjhnl0KNECD
H08tsEtGARAznmr3M/gAnvMiF2S5yAIuVinU6lqG8RwZn5iAa3DCo0k7mFMa
j5HeZbvusMpx0kA8T2xoov7sWXyYhXkLsP8gTMy+WAo3XZCRnsXhzPZtNCzV
GNL1g533EbaSOrKt7xnNHOyN4+GE//eoSNajV2oCd6MWQIr6sDAkGpt2Cd5Y
DOCI5H2b0mvfJwWKKRP6Lp1sFQuHMlhmuPGO51X5ajSnS5Dv3S9TSO9u4C8v
FjmdlmNdkCmxM1AAhkvGeV9hiLdPrGBvax/UZQZtLvnj5X94EhyqBKIutBLq
Af2fsXYg4SxvnKrFNTBvNd67OKpbc54LoZ0OvN0Ve0S5WjmGoPuTo1w8gqm3
uROTgPyCA+sQkVR+l66IxHRlF0Fy1NsW/EpdbCeWFSwH4DN48nDx719pPiAy
fz3qNKtzS6HZryD0YTA8HoAQLSzcXUWE3VStQBk7pR1XtFc9hFDiFZU31gCB
68kaSsWpB4Lw3aDg6HjDJwOMpdBbe67rG2fybYqBRQ1RhpyHZMgnigXiFuB3
5tns+iJj1veIJ4lIy/94z3ttIPebNcm/NJFKTV3XyH3me1dX+4UudIW8SNIJ
s0WMR8f25U+dQijvAqslwU0zJBzJDn22JlKn9RTsVQslVfIHUE4avz450C2Y
pAC63ZfLGGb2ac8i9MUBgoDkn02sel2vCUtl0SdVcs8jIJyYPLJzbWOYc9JK
iWild8LroF4omuuSvHB0hgTQp6S0fTLJKixywUM8tgnm3qLvpGeh76f3g4YZ
Tj1xsLrF5jHlym/7+MyYO9NY2fAedYSvpk2mtnpzADcHUJKTAoUg1xGwqi90
m3lf5kMk11+LsJKeREwLUCtBB4XwJ5Wf+uZ/WEdAqCgvZ5U5bwZCFUNfzFcT
n3EvuR5Pzqsq53uTaOXEObgRJkRziTGKAAUE2d5II9GCCrHXdCy0XP9beU1S
qjubcsrEFREFGY/XR+p30n7v3VZ+8VtluD2JvnMgr/pv/VwTFanupZqpoIde
C9LHUXOQw/6NxfIz5Q1zhZm+fIPW1Hu4PsmNWKQyEqUCX8GjfDycF7eQqlQK
rXI5+czjfZJqLRGO07GQyTe+fT3jvSoPG+N944cPI4+rvGpeddFSFVYLGIcV
QgBszKwiIMwc9ibavc6DpaySAh7hYWBGaKi/iv1JMNPHmi67djG0mfOzl1CI
TwjM8mbCIsBEj/kKx5YAiBXDxb/OOkoo0FKK3/g1e6PPmkgeZcCKrwILDqvu
Ab6+NKmoKcjrpsrR8awNMt2Dqu1tFK1elgTcEQMacCZGG1okF7ZeGfR9o5CK
qRXuhXWbQ4qu+EimWh7Edyx957GiV1OQVKlSBc7RJWW6my7gDTRD0h9CV4cW
HFnjPyDwebBj5NLMsliK04aQ0xmTKzcS2tZnVEOo96Bgy7gvsw0pfNsaKPl5
LLE8GcVU6rIb7no+Zu9jbfbAVQkxc/+6ZsGIV0IrEfu90lEmYNN8QNPsCT8D
SO028SgGHDMAN4sLmzxGiNyLC5CougpmIy6rrgXOonVQ2Do84y/V+kf/h90w
KrfPQSz2lEd76cVmAAQnoLqssYYZNrU7NX3ifSlKNMsEZt2btz+bV/4s7JAg
n/fUS78BGLjSqPQUpqIV12pB+RbKE7TTcBhjbgsmnfxvyJDM/AEeGIyqVF/W
QSTkRqN9hO+YcYTM6IWVfXF6BJbQJ2iSLW80HaXJishtCK8E++1YSkSs7Jgm
AhjdItXRqjOikBB5TGBby4ZKAXob6Qefeg2vjnMy6/ZLbD6z0GKGPjHsspKG
4OPWkqNFaMQOAGoOBJ1pBt4eESqStifs9UKDNR7Uqr2JjjOtx8kPnkhJKVuH
KfbZrOuiY6lyPQCFuQSs3jt4RxQiZEEh5SYQBtDbSPgJzOONLkagOdnDQeCn
DR/fU4W2qEXPP9Vfyrthk59pS8U4D2VIAC+Q5SbDBI+w7BAgd2M8S9X5qPjf
Zv0Gm/E3suuu3Qrs1OlTI57gMxrV3XidbNwoHGN3h9E5au7lTv1RC468IU4k
cEuiwrn9Y9g5HywEVjnKkHbHriCnIaJkMis8gT1Ttbrtc7SC9AQ4jxwOJxHA
04fabHYGBdGjQpoSwPV5cRka4eD1D/+QjxdJd0WkftmoTKQPSnyVjRXNV4QL
aHpVd3v6OD8iVjylHjIsxOKHEWl4z2C/79UJbDc7Ln0oCtc8HMsyLIinJ4/C
XeM8mK58gxqeIN67dUUlTMMkxS4IfGL8Qx2xma0FS/s9gWk0OSzL0O2FRoo7
oSzwGfllYwkFQMCQieVs0H1TLjc2iJG69kJF+7thBfQ2XETcxqImlrySdh26
Ui6zqx2f4twgNS77i7TKuNEZVtQ+Ic4x9kPfVi3O47a7JJioLFkA1Rc6b+63
aSSHcHpzkXB1EJQwRjcaaVd03YzmSpcyQMp1BFUYgi7XZUg1tOpRCddmroxc
P0aDT7d/kdFI260cSZ979SK/k7USWrz8+hFjPsd35z1ujYCrdr5yPzFlWt8I
zXEYX2SDu1lyApjtGUw9SCe0RftNesNYLJu0CkBZrmaITQ3X9M8N8t1R8T84
Xabtt83l0RUOogPN4kGi6Z7L4GWBotaf+rTWmeteytsGfDmBkZk5UNnSaVSI
KxD1Pg8woJ6icCu71qs1H3Uh+g4MQJPeZ739N5TC6sbcrD6DdZQgoDe3Db1h
pfFPaXT28los8MuU3Ba9HC751wfHzdJndJVunhPnhtlrGjJ0Qs67Kb21Qxe8
XAGT4n0OG0YWQ9osxrx0in0Wl+8sRGFGxFFZplksdgrLkEnL40Ok4VFlZ4bM
wrPGbxGyb0OMvhLEColx6lxuMBXpnkC0eD/P7ySl7FLuSay57+/QpxO273es
ZA3a0kwoPWefKdBrUaX2rhhd5jXU7Zy67EOaacpR5BNTSe6/+7dUs4cafegb
He2lOV4auoOsUa7NqTTYW9nEx/n1a80iVDDLezStN8GkguK5IT/d4T2fRRAC
dEgD80n13x6yFFvR000WbCshDf9JF87c87KeYDlT988CSs2flvchbZrQly5x
6IGO+Gt+aUsZGjGdtSMOmQjX97jRsx9hk4G8DToFs2iW7Z/QISoc6jGX3qOD
w+b4Q3oCd62T+EBd0QQLsrGOhEwimDRkkZnQBn88um9831Mf/ZoGLAl9INwK
Ck3ml6y1Q0e9JalIjw0s7hWpfE2BnHGJoVVY4ULLaElCHqpl5r3nAPdhNVkB
Vd3tknT8Kt45VNtGI17W50nQ9jMA5p/w7Pv9FR1zcKJa9t2JBuybr8AIabDs
PkfHwccgLx6MTJ8YBZpgRuq7RpYRkSi1xEJXr+gV4v9UWUw4XE8+a45SAVn4
NnXY1QL2VPbftI4wePZDvxzUC7aVnuIgalYZ1MLy8m/0qDYCQwhYRlLldqSu
C7qE5QFIDWtVZShfB/g0nRXXXD5X5K3EVkqi+JfDMQmVTj3cLl2gDvjBSbTm
UVe2BI0xxVRcv7/MK4AWY1b+B+o7PFq56Ni+comNgVsyrVtEv84OKqOsJCA+
TzRoYzlrHjnYJU+Ekb+A322b+t7ah5X9b5/vyGfLC6OsPQw/lh23aFo0vSH0
SuWkoD5rbXFIWM+QIn4ctGB3lYDfLbxfe5zQ8/EFzjw7H28e3ghE9212nIh/
7LDlSsPK6EHsvu78Olb+B3SwipjC9XAvnGbglXkaKkVdIUXORcYGKlACuMWM
aZvaEHHKgu8d1G6ztamJe0CVOW8NIubt8gj8anypRiDES/9+I5PFk/ZejMn8
uNXbbmvu75J6mKEKX9LP4sSK4JdtI8B0TDb4MTuvRkgi3hGBhPHBnnQcFoMW
ae3ZdMU8mwADRQzs04UKy5L5Udf1lppaUckmUS9IelcD3XUpvChygbpf8BNV
G9gLMlygd80W8c/joXkT1TMUKjV6cn0QuQZwwpd0CdWFCdUseG4Lhu11FlM+
cIqX7kLakCx6fQUwhUzCPn7k+Wo7Z3M0Y0NPDoieO5sSQo/ckRGAcojhkEdZ
K1uv1Dpf3oCNDosWm49d4qz/xxn0TT7tF8E/5LhPBR4kxVBgjzwwfsuOzxr3
MDSFBjkQPUY9Wacm1GnsQDhizIWsbFxqrEjwdkQxlH7h6/BYm+THWu6nkwby
ImW6RAw/dJ/VmHr2gLnsqtStfo5swPB9TshI9dCdHOWSdF883mF2HkSzwZs+
B5Vtu72qAKrkbRuIuLs/DEOuw5XP5BqLenPRiy3RLzTBv+Ujm9HO8NxDue+Q
mqEaASE2JjXiG0DewzS3ddMuPS6+B9liX12sqXvPYZI1oCEcdsb2DR81Pzj8
N6b0zRcud9Gjss28L1JamhZl1I/POVMfJ9dhgC6NrcSRRJZsNgMgrIUQ0Axm
jkE7Q8+yjcNduQn3iuhk2esYPRkE3eUEAaBuOf8lpuZ9R8jlVaz7bmJ3PGnJ
IIN8bMy4RLjrn0mLZ/IHr/3rULoPcsEod5jEf8XoRoXvbUTAQVgcnlN4dGcH
Rfew9FS/Y6+2qdseT7+L0lnknpWVvyJBQuIJFmpR5oY8siMKcl7QJilNr0r4
YZc2OwGfds/A3MPrLY/pgOIqKyUyNeWguFEEL2YxS/2rfkmaG1m24x1JcYdc
L5Vf2c/pPTBNjagxMgdy7SCZ3UsG11J1y3phvta0l30ERdYx3ShZSFxLe0/w
QwBHntNRLwGr0gA9LFSMRfLW8tfx/gYf//H3RbDsvqhiS1V0KroSU3KeLUpz
kBRzA8c580GFpXHW1U0KS5i+q65IJFRYxFaS8x2lsHaD7HjLF4FzPNicTOGF
9CluLJbLAgKE6w59/X4EPThO6UCZuOV6DkJWbItzUjOa8Xq8D8idJ1kH9i3j
ROrsxd18JrA3EeBIB5TfQHMXVdp6936tTG6ooxBnHYMN3dkGwqOu4OXqTcXF
K3pwrf8dAJnIxaLn5jeSELDuCoHPjyB+5PzPP0HhIaWd0NVNmliokk08Dhhv
eEjjKDBjioYiQmx5zbMOHMDaYOgsMv/1U0lJnEhALT243I5y4b9XpJZtdw66
P66xpCrG7qBbrhcak7f0M9/fEycaJjzUPgyJ7YA3ZYyAFtB+mbHD5rmo3RmR
ZHPGJXecrIZlO2A54fFsNTDy1NnV+bRqdgywuoUgpcFFsFl8JpbZT5Z/ogXZ
UIkYyYpK/GpO9Nn7vhwq9z0gwjG4Mw4IYS9sbIo5sIAHTpHbRgz1Q9Uw5Y4b
peS10qJ1dBkcJFwPBF9WVDee8C4f963ABjuafKdvfa1bubqh+D3o0ceszccw
W5OayP1qGzJ7s5rDKHicHllpp4+LsCWjsj2JJj/D5aM86Q6heETetkwQw/R2
X6SbMsjkGWgOhtonOwhgdV4H7UJStEBz4TTotVZFOtHmKiiI/M9YsNLB+Hge
uRj3oUlQ07rWISDm0/aMXHC7+9r4RHJqUhlLJSHsNH78pAwNCJxWwJmYAYkk
zMPuPLTQwFutSHefZM3zB6+KuK2a8AAcFPkDZQxJOPH8/LI0LOUjsBrXZJv4
X5AyzVKCyB81cKW+9iRK/znGWqCfuqR5QiON1gRWFI6PKKqh+k9rj8dhahDb
/4KcTUF4opctNCWlfF2MVob54TWnqw9FMH6pDJlt0Vd6tU9Y+ohqRJDPY786
l4DerJYTnVERT8JhIndQOXtSnGqh0wpyAjQOaDsw1+8MtzMqNrDR9GCwocSM
6TH+eZpI4vaaNTRNvpdNll9xqx7OXW7ddcEzIFHMx3PIbfn8VzsU2v2TgqYj
fcOFmP1fcggaEdtPHd8KCSMS9wKSFX1MMMYSm8Apne23noCZt4xtsnIX70vZ
OuU8cHc04Z9kA9PXToRyho7gDR8OJ7BmWC+YyhIIJ1Z3aDv90rKBV0gqE2q8
ltaf7sxTXqKWhrKcJkqe+xpsrf9ezbGj5s+cR/XCZHZ2ET/semcBxThg1s8e
A7cOkG2ipOQnzFPEnCK/wADkLimN9Pe/5f5gidffb8UC8y30dmOu2nS7zBSK
aKdVE8c57BvZs7rLG7E+L7mHUYZ2QF+Eyf4iAX2J1x9Ay4judqKTcEIevlBq
glYq+yYiUPwASKgdRzkk+ObyrFgOheavb5syMHn83Mo+BdWE5m8cX1PHIPpj
Mud2faNC3uq6h8UuYHUuOaC7lDjh51JvF889HVtAOLNhvsjQLJIiFTPHFH05
cH5E+l/az/2sizaqCQCIej3VVMbd+A6K3HxbX0LEha4QAmfK1GgBM57JRpFh
STufrWevvpzGlmdYvD1qb1ySehZCpz7dq4Snx0p8GjKYirQ8HOvcmUjkRc5T
gfBD1ivRE0bnQBety/vUD0Ga4ROj45w9dKVVrYNi6OIC7oEF8amserbgOX/J
Q4inAwDAgGktlfXeUYBmb8VBJGq8xai2E2UR4LXFCye33nRxq7rE5mRpVB9f
iF11J7fm9PdSaAoG8B6R+wxFulwlHrWaGFW8DzzkAgWar55AihzlW78kkena
4F3/VA3ISdD/D4jgHjydr7F3n7qjetNxmB1TlZkI3kvHRIozuadITCrKbX41
BjkE1XIkdgCoWbygQNp3iDeqs1RSNvXnCKPjED0/D9h/9ypCW4QP2zc4BIcX
kKAchHwqe26RL3Sm7hdL4GijDXC4BVkQ1oQP7ZMkOUozsUvNHmbioDkVpt0m
+s87EOXJXnw8Vi3vq5qo+6eOK51065QR4pFK/zh4mUkC8vHCFfHB9CovmDaJ
lXf5ZmtxJjOM1y7M2ypFRw8F5p7I8pfEkMC5JHnNDohudsjF+ERmOaw2V7V0
fGL6AGnczVj+FCp9PRh6vDLEvPhAwk73e63t4Jgc91cTFdzugq2iInkBEJtl
zpYXxycxHRC66NBw/1reKqS98V0mkn6MbvacOiVXN1+jOSQiWWtZhkhktzg7
qkSBDVqOojpzshXAq2q7SDjDc40sQ+9+QSUVjrsE4+gC8m+LpAqYLfgin/Y0
UybKB33JHcl8338MTsnhqhUzkSUiw1vZimDDO6pv3Lv3zL0aELXOZB5LWEPB
UMG7/UYbcJReoal6L5fGqa3G/JZyyOVKVmU1f0hcJU2V8qvO0S20qOZ8lwV7
xQUJ42l37rhmLo+fD0tQAu1RH1tVYQRdQTMUjxWakU5vrWHLen/ZzBacK1VN
+KPVbKTxqJnjnPBmsZylnyWWFC8rzWChNEQ3eZaW0qDRO/44+bMGAXUCiyky
INtuTWx2+L/l5S1WduaEGIj/0oaJm3w7lmDgrTWSxr2swucHaHky/S9FWOtw
y051Pa3saoJLhCT7fv7MoeGqr71wINm5nCV4G4O06+itbk7ySyRthwcXlIkD
7mr3a0Bqd9qOr7W/f0KC0+VQRFmKx1wzmr0QUa9SBLkRiwhAA59azOvE7Puo
/QQ9tOKbCxAy9QhP1J1PdTLVo34aRxDQw4JhP2NuOX2anBjLdSXscK7K/rnT
VWFN2ax2wFMDeE8bI2yWLsyjpjbuGRSkUVQ06A+0H39QRFITWAFhh3lLMm5q
yuiXqwEdb6c6iw1F2U7MT6CfHYILPUhWxKiFJ6tzSanX5kB0AOfW8S5o9s7n
dwE/t33zAR9v6R+0w1ZiaKMdf77LLHLZBSsqEkq0hZnk69C37YKllEd/wvpI
u/DkMiPKNQZNGUc2FHTqoSpxTR1aYFhrUankTkVHjZypdZY1CMciBfhu+oyv
smDT3iFCcDAyCyZZSkfW9NWjNboYLPzOP1Fx1vjCyVVjYo0Q84PQy3cWqgcP
y8Dla3dkY5yLjYVT9uScpgmu4WoRLOLEsEA+cw4OSFQXIdYeBMGzYN7DmsFt
MHU9fP71/j3GCY+lvA+tagh4MPhkubXvQYKfORMRpnSoETvrcgo+HV9JUGlq
H17bVCqTSUqrayAsDmaakmTJRApog3Kw9n8iRifyD0uzXIlnPUhXwwcG1Ma8
CCx4mbKmWaFBRH7Zrc2bl3sxMuY+chihbqF+FqOou5MiQgISfK6tDbdzQvGX
otdN/+kh5A57Fs4zNpq4clybNRBdhh/34qSf8CEJth3cR3iwYSIP33OzQzbG
uLBdK9NYyV2AqN0rHjcoqbHKLKoLeKTY57UVBiux01eHvXkYS9i4Pfe3K/NR
aTUYu5HK5Mv1lrRdIo5BGWLMhUF0SiFJJ7pFi0pxjuQKvNXO4TpSIDwl9sh/
iwDyWqeJefcMGat1W5RFM0LArfZzm6dDClHYhiAel6OC0mt23KtusBOibJbT
2sHvUZy3Zfplk6NtpbGeRentdN193ZuFcRGT5rod+N2Ajhz5O5qerbsNaSEu
MrgACX0gkE+dYQpECzDqk94QAWf53qkHNIUopzK6kdwuyEvYYoZ8MIn7ADBN
kLZE+tKZng6jRCT+34sqv9Ofo+QqIM4oUrjG80DqQhV9fztM3ddZ8lIhZWbF
R7nZgbWnY5V2f8HY3H26YFdZ6SbfPd8LLFC2EoQnaGE7wSrMH3n/SmIyex8T
hLaXfXuCjCXgyJ5VHIHxn/NexgE+qiT4VHINdC9sDuaH95Xe8F5tTwpS4YFZ
rlasurT938nlYp0rWm//+hIFcNy2OdpVcns77TdfKgvyFnakPLEKtgAwB5Sm
55jyD2fqQNhuwuW/K+ENXiwJi84oxISnXus6fRZH9zOIAXiEAbt9cT3OFtq9
szXgTaOoAHzAc5ig7smoKsVSGi6uMF1KpPFfR9bXkC4zBbEIeRJSpCEOp+1s
8XCLPA5CJ0yX1kTrqBrqJxnf+jnu01GyOAMrR8YrqnHSkZB5H7x5TdK3UtJF
SgUOu8APgnzsJS/kIh2HIES9TICAuy/lWcQfJyplLYSOg0MTcX4MWk6aHbD0
TgMRK/qPo3gANlcqLx1iNbB8uMwM4QyLcdKXFGg405zsztOnLXRHLb8KXdnQ
jC9hUqcxJsaBGQibE0f+E6CSHxDPK0Dv/nfX47ao4MGarSi3tsYGb15MdttI
6Z7gjw1aHeaIdHPLoAUkjLRTC6Q/AFwnfPCQffEJgdVpLlW6NRvH5V7YYCZw
BeSTc4IxfqOU2yH4dvMkjds5WMFp5LeZpUAH1u7elqAnIM2YqD/kkTRUknul
h0d2HUgqEdivZfSabxn5OoFTTbCXM/Gtm+jd7amVrcxsfC3amJQfuChmSfOu
mD6Dtmc9hfuDTgS0mNNhMWUdFlVSIpGoPtupHp86f95TtMCHZ7Xb0s6xsJVs
DCUIwwKtcmwf3ULgGm8fh+sStYBLbV1eSPuoJU122dsVtpHr29xSh/yhRSzg
jb9pMndbsIv1ZTaRoI1J0JzaAbJjcvKvtsdVYNMw0ojgqwToL6yJ909/bbFV
PUe4K4+1SuiLgiTOFEaHWi8wkwMLv0CGjpAV+o7P3+/gVQ57ZF2QZ0dxEEbl
VEoiU/7D2GhULhWQnoz5fdUv4DB6TF5sV3Yv805IOarbW2AME6ux38P0m2Lc
5mW/m24Et2n/iwWIHLtISrWSVY9p99l9pvY78N6zfr/CbcotFnDVJRbYy12+
u20gGyWrkMAToysvLYBetCvUBcx6kTUBxPgM4qvczRq31jp4XbDLKxOkWsR6
BtdWZblw8Q01o9uihiHvrKOixCaWd6pgTf4cw3zAYco8O5mYELhlt9VeMOOB
2uV3L2lxglee6bR53WDc1BXAq3vsJwu4YlNlPWPYk8JWs4ukJBl4Z9Qc+bqA
wk9s3irjRXxkTVjkC6HAUCR92MUHqM40rOmL64LpDxRSETBvUjMm9oWQMIYU
cWzPAJEWzRuQLcra4nkkOlu06VYaMhxyiSUAaY1szkYlKHDtjx8jenz3u7BN
VA1xEYUF2Mye9rux/hAyf0gsvKvrVaJm+HF2UZFhGgvCLEDrUL/B/ua7qv6y
mtZC0vUM09Uiucm7pCoUyp8ZWaTziOcVN3Q8SPfk+CdUiUMsnyNVwfhCmFWv
4Hi4fkfWd8ZGdcmI3IvnU7AZaEIwIA0J6HyI+0zkE3DdAh5Lzrl+um0lP3fq
18HpUESFh+Nl1ETucmBVMuLG6wxDxAmp57ah7Jqo97Q2RdQL9RLG8spsu3al
RuRu9a5QvT7T57FsvVx8S0UMOgZulHEtP7yjcu3My0ucjyG5z8u6eNNWDfUQ
CU4dR26X+p6hg+9jQXIS5BCyS3vv4oL2VC9F8+TXbHmUhM+oIPzNFieJQBHq
jIUo3iQkluxWgNDhIMAcd3ClhNIGg7HcZAmkk5VudQ/2q8sbI5m/2tc5mABq
slVPbLuU9JyGm57ZXGO8gI6/9JwSX//GkajmREEb0Mr1guiOyaI2R5hFkaaq
vUS2/E5SLHqTmrnTIw57ANGB0isEjSeWTxffR6fnPSTLoGkqyGQHcg0AoZeR
kJUxJBMZOKKGm9vdkm4HQ24uxOxgpmLFmvOQaH0JP3K2xLq4TF8eu5X23z77
1ZTLyz/H23V2hX+Xg3TE0koaaatZ27K6vCvivHMSOjRWqOis4hPPs4w5jul0
07WupL7u4merP4fsoe9K4yZ8zqvXZJ/ijdNeicKBuphrkW/qYhUEeec1izqh
Oiliw9xZkgPsTC4sHe5czduHtbgw488WWWsE3Kl3ApOCRRdvYy0ZgW+yyJIb
yRSDyYrGXbDZesvEhDhGF4jT3KuLoFMoVw5uiMQDMjhaV+ChUsFUDwfCu275
RjWZtGAE+AUT3IlfAVXAJ+6e1/r2ni0/8tUTyuMjo0PSpI92vu0rKyP1EZp5
YzvY1AqY9mx+ofTwnjI5nXpuegWzW8nB2tuKpaXEybVv54ugoSaamD1D1sHU
8C4znDWFiD68CT00Jh4xzOSJu1pu9CwkTAAQILiJEOpPfoqiKmpmDf48J+RR
pR3G0C8Q9jqkl94G2+81JyTxYlMOt9RrTy5d1Ai7tFbprCO9hE6BUPgdjp0n
PxvXCK8d+oF+dnrnRxbM+lODvD02sPU2Aq80OsDmM+8qg/7pKobPDvYSIRg9
dF3VtuuhJdYItGZwNOefgzt/kVKuspKsSvDyY5tcslZc8BTkNTV2zysLKkdO
455Sk9GBQ//o3WB9iT4o0EeO1EJGIyiQsKbo0ZByh3Vz9HEi3qcihmc/NNnc
MW4F5Id4RLXLrbC7FQKKOmxU/6FFO4593+BKZkzTApifv3HGyLiLv9KF165O
52yvvI5bzcHcHajfend0xSpWGrxcTYKdMl2A379H9gvXN5Vosc3ulOe4yTUt
LOt0KYkHLTZEbNRu24jwDChFgi/UNs5DgBg4xwWiw8uZMXmlCJ9OVK6iWO0T
K8i0Oe6VHTISVUhDUac2BduR42KM9xioIFwnEOhsXUj3P67R2Ieg1fNwhA2N
zDH5Wzy0yRFDZOsSwMznWur/HAiua2I30p0oRMddo/R89FOoOmRNR4w3RrI9
rUAK1/71dg3wd7IgtpOH1g8z/ey2k6nVAERwsu0Y9VsuSg5H/pgyJaoTsxNY
S3PYG7VMx3jBbcHoopxVppy+iiWSN+rQJzhVzah72t4XLTVMkogsJpIPxkL/
eGUI6vMwiLwEU4H6Um341FAR3Rgt5s+5TBueTjyC8uNY4SvEeKHaF2XP4h2t
yr05BijHAcyjFZwMyhVpyjNXv+PHEV/RZ84YFCbUzFtTxKyTWKfdseIsZizj
/Avd20vvBgta/GLUo33oq/7pQZ9n8g6vrVTCWK1ffDe1DslWOjSMi6mXec3z
PqJajEKL+s4oN+sG0GBSraBOwl+W4iMBtrrX9MbGE95aLnnGb0L0ptEAMbIC
Zg2YcFc1ygS1KN1C5/telU05LtcxEt8kgZeI7sxwClLH8WxgfSIEZPsdKA/w
/xW04eAQYaZyv4QnN05RjCAjLO5cMN/WOMqBvZzXyLXRHzRvGTd5Pg+ccPHR
lreJb6AToAPb89MrYR1NvMmlHf+WGoGlSvJxENwWRw47wToH7Ng8XXthqLhh
00hdb6UU8xsNfHT9xSrkENaavn67L+GwjMmGqFDA4HPU+jW8wg4JWu4FS+Bp
NbPFTF390aZCa8Fs+9J0OBuikCcRmVxTp7G+p9RDW73YHCOQaAAHpkP7srRE
Rqw/Z9UYUN76VMurw9Uru2DXUEPr6AvOXMSHmf+gsWHugeNp5WspmcIRGr6c
VRgOXbmhoaaK1NdjE5WMR0ZYMDQjRPVHqo4zoDE9pXgL9bUSiPbEWbkIOT/e
CQa48HeMrfhnZU7l0YdhQqfU4DKviyjQV2AA6Z2cCg3zwxZJ7Rf+drCvTZ52
TbEtPdp9rk5rexQj8K3Egw/FXQapp3toq4d89j4ioMNf+AhWrmEgRGU3lqPs
mDEAUdYE2eJT6yCP/PkvwNWgMOBNTqlz9FiXRYRJy0Imz0qGlfTW8zSHV0/a
w/RlX+DeV/hfiildd5LJLfEjsA0d42CiKhBGrqik5K9OST23lyuKw4jv/Z3O
vSHIVsrwoTbi+nc/4l8esD5B5k3JI6WoL8VG6BfMqQO+/3+sTP0NYAjfASbT
dX41Y3ZX3BxviS9HmxunNfGDyAe7cg5TnLenJOkdHTYXyyUzYgaS1nKWaEqn
Kc9BLndJa4mBlgva16Xnygeu+w/nt3S849On9D+Kf/LZhiuUPJud8nvPpUDz
VeWA24Lj7WTJ0UJSlznMAyhL3rFUZZ1gGQUXLui4/UlhOoNAkdG/uokYZdZp
GBEWBssk2WivBh8PNd4sDYmI+5scq3wHGOmbxBWR44WFk75Vcnziifd4usx0
iucD0JOPfZc6vdqfLINBqtFFCPDe7SJcS15y1P8szHlOkebSfaTaNSAdQpyl
5JoQkHX9No6zHbl5Nr4H6T5mB1J8OkYxv2dQURZahhDckTiLPiuBFlmxOynV
zpF6oyUL1ECWFX8bHr3yjnbd5lowHJfzmyK3y8yZhVQvY1HUaTNQUn/GP3O4
zTuvR4d94RD8qQLs77fR7Zn0M5BrEAem1LYkIAPFW1VzQ/p/CVj5S9EY4aMk
SjuGfV0mTyH/AiBGI6kkj3QahxAcsp5+D2aXjE8l6a+zsWrr39MGQc38xQ8F
BIo/HXslyj7U9O1/UK0oSqUuwxbEQbdBXe2GyXiLTclnUpCV4StAxYQjHC4Q
EStNn9zT92Yzh1Vx0Bh1F9wesRbXYoKTXNFmKxoXi6KCkMTJPIo7Gi/Mpn8I
g3/q30AGXInDSrCFJ7WgHszTsx5OUr9jdHZFWc2BGPtvWv4IWO4GGnRCmlTU
DdBEE051sDswmZ9oeHmwyB/cv8/pqen803zlDfEmbqbRn9aW76lKO5JUNxyy
oAIYNzHG0Ipdosup+YIwfjTPhBomX5lihajbaesMO61gJvLcojQd8nKvVp4Y
Linbti1WxvWlBnS2r9TEEzRo6SKm8pWiDILthnIJyI3NcIU+aoksVR5MEjfp
Qga8YoE7M1ExXPv6UWzl9UFBcf/Am2uYgTWlpbNTGj7LGB4t7iqFoZ+4awHp
0GTbh3gGsRZ0GpsoD016pDnPxomqcwM8oqSBgOswVJHcQ/o3Dh0mtGF11T98
hNgSyunlWlDQtwOgS20nsGoRZrx0oKV8dHm5kH8aFv+pMDv91SVrh/m0FDwT
BnNeNvtmdhBYukQ3RIp7lLUzrVyQHmqLDyIxzRTOMk8/k5dWFcB2LUGOdv1G
88/vuDUW3T9909PNytBhtUL9QrMgwTqC6eMLqBB08lrZbbCdH46K9cJPPE7d
FcgP6Fh63Tep7BN8v1mhXMiW4sbeQ8TEGDmBliipj9yUQF8n19Ztx1Opiqzp
4s8Z1tG65Js4pAW7fkwgwUfh98c6YNfVt1+73cYxjFCNejFqDVQlWXTZjstP
usM6QZvEflcIpru+0App5bcUq73yh9s8fI7RYONMBV9aM5XHyT/uWl15rSSN
LwBDdQQPZaqjrCRZ8+CQc7nqJNFBT59OUN/e4uXpX1T7q+rIxjb35iKIrIxk
vwYfodUHDHMfWWaHNHtsHVIqMkoF9oXfQze2Vli3UAvDw8IrNCruWrba8Qbr
YDZqn2M4BmPi2+0s1eUc3djTsKkaTiVprSA4hZl45TqvFTTE2tqEj/oj0zNr
kRsUw0qZh42ZOW5V9KvJBh0zx7PUMryO0v4ThroI3nCQqBXQoOhFylr+AsR8
Uge35+3JV5uoJkuvvkaw/Ckw3JG9e7QDr1bMmwBDh8DBttTKBBzp9JaWkQwM
yzeIgCBp0AiZiMOc9fbrXIrRH74No08VrE+tiX/UJvczZrxhlwC8Gs/xAZBb
WXX2SxkR0QVg99XAGinZifoEKt3gEOsL7Cp79EvIQcviFDiN+ArcB8rQ0n+p
hEExDayFJWurFHHoQLzHxLAeM2JjALm3OJ937U49ojfc4bSAaXhm8GnE+It2
Ed3uurpz8QfJROvO0Wfg2OUiKJsiKfHB5U1RDblyUQCeVyrs7eCrlkVzSAAR
wsVh07fdEP9RrAfyPPORtHmViJJM+YChlVy0BFjM8yYbyqCnS9KEc4mE5MDe
vuRlwfDp578eRemQMmZQ9oVk0n9a1pHw2ZmZ5XPcNMJ7WuBdPlMvv14E/0eW
q+cM24cFdj8HbBF3wEmWVF/ggFCyt3qmVD7HFbKPmwOMAdw0LhbhyHV4Efxl
2dUQJfGVVKSBmAmRmZ0Y2CDhAgXEJbLDTkGuV2xatElYhEFDpiQf+DB3GGfV
pysqXdbEN5q6goXmhqRHPm/NtRQvDNopRDtRuJFkvkxER2M5qRoCOLBsYgHq
RVxPH+3xhfdwK8O2Se2v1a5uyQcWIChEyck4JaPLTF3x2tKBv1kFkzAO4noR
0OHCPx1Vm6SmMPA8VO+v+0/Mw2aZCtyU1XY0SfHRs3nhRZ5KfUQw5mIqgcNF
Jybn/yMeHJjDJoDmwt2ObGvPTFoSrdNee0xzdZMh4uDh8iUhOv/6HQpJ8Y7h
7Eu1CTKkd3bjzj6jDszZDuy3mENvE7jsN5o02Q3QE8hQsniehIJduMlJ0+jy
dJ0unfgwT9RGe8WsQh44/OtOpKq46UlwoeoMaIv4Wq2OfvQaLgF6viHRSHOf
IGz4Qp/LznXSgy5VsJYbNmhhJ88zReJDOVSQ39sSkZ6DuBuF01L/oWYLvm4y
lrG2jjoVBwwsJPau3G7s95kgTpEy/Qt3a/wMOytTsI5qyAiq159mm5FzacWb
conZuhSb0awoJnhVOBneVVx641MjdtwpQpTeCzhZ5mxMLPhD4dCc5hpz27VJ
N9bsyIbs48rp7kEPZcF1E3dORFSk1Vgus9GGv0ZaoKwQGJ4Pxf4e1A2tWhT1
gTby2Jh66f/q3LEW1QFYUhhBrNEYimNfMRqH7ZqLDgxJX2b+62JMMYAsJsHz
M7n8y6KF6UMrxuavaWVjsgk/RFKIK5hhxa7CYljQkolQbAuh+C/rt5OOpoTZ
FVGFUtWzgg3mkf7VVxpJwe5HrvhNxKUkoSFh3kprrLQ2iCYh19EBHAmQkW7I
bJDTOZg3sCq1bNcjfietOPpCZpjhAEQrNLHuj1/JG1GkmCBfEFg0urro891D
sqcWRk7ZNmI4uflktc2J5n1rCsi2mN+T1TJ6Y63iFqN2U8dcOEapijVm6ADr
R+kw3WQ+R0twOk9QbNSsRJj42zLpPi3AKgxUC+ZL1pyN3Tl6uWm8miErW/kX
MlXQEn/Ny0k2CZOj+dPRFPXrSkUOxMS+qIe3Cuh9flWQ8ARC8vFPXYnf7ALu
Scug/0rp2+DqZ0yaDD6tObBOK1fvNZfjYpwrgSM4SrPGc8ur1rUZY4kZ6d65
rNPJbbnPrQ5JbyUtSTqTX8SNp/i1RJzNHNHhxRoV07EP+nS6i8yLGgXTxtj8
kWrnq0kQJ82kkNTO6O5iTTaYSvOnrlaOSzkNDWunD0aTf0T80MBykAyLvm8l
QlGF9xwgSiwNhz2i1P4VCqkSoqDOTis4vMx8VPoouitOj9pp3q12b31myPyJ
rRqEGwGsffXZZ9k+Phw/CEJoNPhAihWI+8lvH2h++0nOPAmiRpsw0K2HYVPy
pcwkzQVS/3ANaOZh6D6835PccrT6M33aitD+XA4Fvt/JiD9Mj7nl2f5amXGE
DPatKEGsWFUtQod8z10PRTkhwI/GkTTMrZIhOC+JwWFeDWlF6g1aof+ysacd
iyZ1S9T6Uxm9Xsvo12oweXJsotiR/Xl+bBMTuwQ1cqHd329XmWPf4wwQHnF8
dx1z29xuIjh12jRgx3v8FDgp3zaiVXE3Bmoxoh1pW38m/kTBIvE7x9uxy4kx
U9xWkWC5KHnCTW+/uy2g2gueqlYWitTvR32HnhTRT9jJGx1zteZdJocVKFJO
nxLg2hxln62izpPXENe24wqep3QaPIV3rbnM0LMYee+bWat4d0AjkOt2HTUY
bQbMy8EepUpN9ZA6G+oNtVbbM1ZECCiKPbJ3H88zgH+6GbAZtSSjmfn/Xy3N
+OpwcCyw39JmN6iS0ibyaZbHzBuPEGbHsNkno/kt8ou+uw6+Pgkfry4gUkr+
iMAmQSa0/yl6+yPBRNP8Rud8BY+Df/QL8EZZDEP0foP3C3Lt1KfhiaufvPuo
AQ5E17NExN+IixZER+plN7vJGLRZeJ9HDWuEDwwFxC60nCU3bxM0VDB8S5MJ
ym5/x35YUwJt4gF+5H/JyQFl0UDXiYwjJEocC4THnbXcYWXP0jf0rKuLa34B
E3r3xW2tyeqgU1tPkcqv+kO6BN0WKbgSYBeBseLbZXN6ECSR1lHuH1zaOzIv
D1Opj0f4+ciNmAXmcgHCuiCjNLgT6v5BeVfVlqNKTmAp1C8sjiupqPNGhIfN
snID3F4qo6nugLVHLzLBc4PhUEItSwq/RdvZuqFD/MGKsQ8/P25w/ZesrfzW
ChPmLPkRaL5Wo5eP4jabeLkdSs974oTPq+nED7TZLCmIE+VAxUoDDZiB6rMF
AVbXAjO0JPowze1OtIzft+FywYaXpvTpw048UKCpZxobdTDoy12hIAIy2EsN
zmpzHCzu8QOxMKt6KmzQJ9YV8ADGQAZ/1WniqqK+8CehowbHgyXg0vlZvuIm
UYPwfZqnYzNeUbSqNDx3GYTZQHTrRukmQhtigwkTPfhVmqVmNy3+vlFrjos8
0t+6nzCSc51+wgdkkEU05oDEhIfNgd3/Td8TPRRIvojdJimEM0kePhJR/7YM
A89Iki6v17mpQIU4loDqkJymXENnP2Ox6kkIIl0hbM6jHUMKjSvyAHhfgz4i
lh57KcD4h6zuQgccnhKDBvz2R0/b0elVAcwjApKxu48n4XFkNbAJBNSbO7Ri
YIfEO/lzHo96Syclv8VuKlPCgFgonyna6C90I7pdG067yL5A01tQ9XLr86u4
SpeY5Q9nmMGN1TpGhgwkijWsBYdiqIySU9UgWb7NWSx3SMvVaKMiYkwFkhrl
2R82AQtAgHBIt+rwvmMOfVzckAf5VoQQc2KZuTXiObIB5YiKp92z40tXf3Vt
PTqzMrITS+AzETMbSG25ESqWAbwS2Za92Sj57Rs9cpbSsB75b24VT5q7f+Pq
W9ST2indX9U8TitbJx8yK8jQcY2j6Mf8A/YKCXK22CkS4P/Mgbt7NOZbQKrh
Omuur01vs+YyGLtLeqkMckoT3Q4a1N2Wdl4W7D1QbKkEqIPC26W88WtvAqjs
+AoXQ8yu8t6ru4hubrtFHOa8oAwCga7psv24gyNEFaEoyWOhKs/W+YU6riVv
BuEgGvg7fEsLOE07YNYjSdlqy9BVbGrDH2dzkINuRE/4RwTOdoo7bWD2CmfB
VmMlj89ll6VaruYjVMB/FPzhVTVqMB8r6tdgSqSO6poQjPivov4YOCj5xKax
y/P5XXWKbNl6s2sUgiRmhqMSgWfPP9QyVcs9I961u0lm8P7OhPMgoKIc+t0E
zjYxry6GE7pUvDmk/e0s4NKIjAnLZxkF+zFeLRxkDFnRXdhLYvM5VIgJTGuN
tToUaerP9yY2+6WYSOLCW6vMvx3wSHWV8lwgfUAfiENx4+ru/JqzXdcaBZqf
wyVCKgNxag2pcrFxYkO+oPzt9O9/iPJUf0O6EV8lUP1i350JZIj+jAYNP73c
rv5AFlrcG2xsIWj5/8jZwAJKJPbbUVm9zTs2NUTvSxbM96jyw2TiVJU1d2ep
PC3yPohJ9Iwgqx8OErb4AZW/14fRrKSb1jwIgZH+ABAkvECCe4VLibV5sNGx
3z5IN/Xjf6sIwnw8NhKYrigZLcx11T0KUGEKkPHAYpHB8A6PlyupmcFe8mle
lgfjcuHTSVQY3BOmoa9YFgOGbnleo87jF/1V2RocAcCV8TsGkuzqurR4m1rK
4EhNCJ4kcpqVEk063+PXaDCOTXuoTgQYiRZKhIWbeDW7r+ezD9F1fL9MEOyY
r/JOPIo7jLCKqxGICbfgD9wKjxK0KwoIHJlYsHyxPhNoL4rK9JWUrx3GR3WC
Q7WhSPtQ4Pn5w8RL0J5LI9mUg4/3f97bL3B4PsRBJu3qrEOuOKL3tRPkkqUl
vHdwHobfEwjsGU5vZBbxcumaE0oCS1EJWZ689W9sRK7VcfNB8hvDHYvTOBXf
Rbl8C+2Q38NGRmok1imRy1DQh+NRGZAW7Kkk3b3ILqTDf34ACYuXev1Kvyko
HMdTJL6yc9wk1PnAzLzVtLPl0OhNaFxviePx2Z4F9pNifwuSauZuKv2gqT3h
k0ISAJ4Db/Bs5RaqKDaolUDFd4RXlGjRzs6zTgSgc1MCHEZIIbTrb+lp8v1n
3SrvTmzmQTpiDPJ5837g6V5PejV7oWLCRaae5wDujcwVBviLwektIS91awij
pcZ7sVvSuMOmwttxXfiwsoSHmVWms3Fdwh9gfCOyEk0KZWUCOki1YNrYHZ4/
8DvhcFSxXCcX9b04Ot+7My2lxAKDrXAYXF++bRcLzGmFPlY+qF7xEG6PKQN7
prha7lSv0m7L+LsgxRkgT5WYj/QcaeSJPNNrfUOBY3jvTLFbfux/vr5u5zpf
hv22inIlE6OLpN9wIccqQ1RR4a7agXleTyZNI+ImkRTANemxGq3GRSlT9O5A
28aA0PqNnaayuoRhRfTYl3x29+2ol6d5tAWdL3GZP+Ji80xsrFaLoZ5TwGM3
Q6JkW1xX3CHs5WD/40GZ/w6FmPQ5eCgn3fefblhDawiprOXZlmulNG8+SWFU
fFfQvE3plJdLIPUGLExpy7wdTby2/k2dcNBEWBTJ9+04haQte3VF7+cariEH
Bgf1xKecpz/MDSf1B6IRl6M1cEh50Gg3Noz24L8Bv2TCOhidmv5Ep018P2Ws
TO1bIADJVXF04KsuS1DpCFlefHappb9UltSRBHZWeLPJKlj2dMVs0Udo4SNc
dl1xmOd2rgkqWNYQOJ92oZE25uzoRcFKkLbBi1bLCn5fF2tWr+mwJeLUTPgl
jcjJt9pDKpOmB4FROqF51AumZ78FBOiXL1FymWh7+1yONmMdiZ0TnBPh0hn1
KUQnTBB2gfCCSCnkN2jxHgM8jvBwm4Q7FasFG6Og8jylRbR+c5VCeC2jUegb
UT37DyHyNiApBG+lzyWGe0whHH9UcgYBiXtjdxAB1TiEEtaHD+LrclDy3xcl
XyqJzWu4E4FpSTBDuLGKimhYvfXAbZIQKTLWjgG+nRyz6dhCkVqIKOyc4zUC
40e5DDZPwgLcBr+EgOVQiJ60jX4hyIw7/6jyc3c1+Afnq64LH34B+H3OEgRu
sle+CgNTk7nNZ2AcZdKvgobHlQE6qhv32RH+P+vbCd2uETv/qn5DGDH87vDv
x7pdUPL2Iw/3mdl9OFnHO1h9NOq9wtfy7Q47OH2Cp/L4PnhuzB4O2QqqmqzE
1osQf5dOYJsTtpBaywyvwTx6F6OmbLXp5ByXjlW7SnwttDoMoxoLxMXUKr/W
uoNOj9/LDECGnx2K3A4o9XRrfHHMvte9aSicgjog95G4jSczJKnkQIv2fuKW
Shf98hLmou3xJYCppcZdnK+6P/unDYHSWrhIpgsHDYwEx9REQi8yMWFJtuO+
QsCdtWwgAVW8raa+Wcmi3zwgY3ZM+jsZCE8XjUXQM3UNxAjR1DQ/LMpnV5Aj
BuKdQad+rqaRFb5ZGOezNr7nhDRRWzYG1x0oElm9CXrkcX99jNyOwJ9aHsUB
yVmekjNF3Lmcrw1X2idgSgBm+SYOBXJU2A6b/YUWdfIz+BylOqOLSBiM3hFq
fEz8hp0GZumzalwrzWNx0YXNT9RVeqXdyVDzOsB/uLWvNT7u2nyMNynYtz92
JUdm5yNSYtersEee5d9ufrTjQiEBajWkNAFq6kinSKF5fpPboPdON9wlyOyA
Kq44Ez8SaXEAE/TGQOJaDZrkiI1/+zoHddcCjDkwE2T9uaEwYi26MIAf0ucF
xG+ntYZHjZiy6Hn+I47RT48KeGqew2k/aul+oEzKYmpVgqjbVUMiFsVw/P1D
1vqwxjIaJqxh/WlHNXECWt6b+q7mTXYEWk2lGeA1uNuFwxKSev21l4u9qBvu
psHF3MtwpZXYoF+Eyr6/a5s3kqK+D31NmtQGHKQSUKeGnVoh34QhnQhabecl
t9W2g5TfGz2rO7gGytmVYjeewz/PBwhHrRod3P8XyVdlSRJXllFXLx3npkZB
8l2bNk2vkQScVac7S0AsvpLT9hcLOXPrO9FSnbItiH1Dtaqbr6epIOXNYAZT
iLhNouCC9eyCBeiuqPyvFa1gjNwms9nNGCSJ0tZLht+C3jvHNxL53Awnld7f
5CwGTb4hDtRExFJElwSzqA8okA7KoJGNLujK2ZZuRI/C58CZyQsrb+hq16w3
Nrmb6bwJBfrLKHpgVs1PFwir6SqXb3f8RBvMpneE2O6rdNFNalK1HdrR6BBq
lPdsoDmYR7zTXyj2fd4PBnStky5BUWT7urvVkpZ5L3nyDeLRLqtpAP4UaeqM
z6aqG558HHea6b9tdH8aH12jozAJTrL+WALpUkM0miZ+IsmWDr3PxqJk4FUQ
rdAkzdtme5LAHoqfzWBIP2YJKV7CtexWFpgRS3lvbPK2+yfr5/8jkszBR2Jq
qKJiOpHneI7xJ05sSzM+s8LRIJJ9UZEYdJfsKaRhrjKx2a0caZCGYob8T1TD
if1NdbcjI2qqSDE2QjMKyqtSzvTDR2Z/Wv6aEUrOeaC2lrxWnkvIxq23gJn6
IqG46XUL1VPYJRtesdmmnVk0UYKD2AXbF9Rn5X/rfTZ/AQV0RKUaMxyXyF6j
v65ki+UAFJma55rkUIu/uAkufW6LcK/p3iznnCPtRqQhuudlUEqh17/5TxYP
nA0n511A8lsLSv1dvbvdnOXcI+IGzmSb5Hq9LaYYY7CDM4LPzviyNTLTZT3z
NJvHsfPqtZpoToRkAogOXfjxeAj1sXaQI4PVrp/O4oVZVlu3k7f/9ZhSJdAi
aEEYtXDLChCxyXpRerIsP09mw0duEWKhm6ZyhoyabQAHMkNqzB92s0eKVJ6T
Fi2Vsyu52vqj8vUggORI68Pi8DZXg6YEUNzw1YhpUWwz4TCJObR8haQoIos2
t0uMG/pKPSCZ3P2aU2IyZvyjUP+2AEmdc+6/ypfUyPHiTicISe2hOwF0U+KY
m5l/5TNbfdpngtS2hMOAIGW7Up2+PO7AYXOhGEZn6+R7rN1iKE7FBlsM9zQ8
UrRnjmIHSoJqwhRkDcola9tSQPItQ58Mi7HD2Hkzxpxk1w5PUhZi8Yu7nofr
dkaG98C0PIn110b1o2yORa3LYSgceHq+jTbfpxNnxjH8y/LhBRldAuMTHrvZ
I/DqM42iJJY3ho+jKVWg5e5IHIzyt4ND6TPqBCCuW1PxIngAbOe9vbBpdGK2
+4jLwqnLxFGNQ4ss3PkGJMpd0wRm/Qx5OvJl9iDJ+kwscsM+wAeQjDNJ4DCk
N8PnAgQPXeuVuQaytHLw4maAj36PK5jGx+p4UuTjLRdSnAL9vjwpr9U6Z64c
283BDUVxagdgvaYH6Go5SSwye0df/Myj+u7+9G13wV72gbX2e6HTXN8zzGkU
RPdMrJCWBrBP344bphiR35p0KM+CFLTImUvfqj97E8eg1rBvJYP18okCVFZS
c5HAZPTzQB+mHtwYUeEHwOIl2HDPZ88JaVoju9v4g3eO8I9PIheh4Kz6+siO
VOi2OSqKkTJdXePa3mMws1mMeRfJ7MKzd/ZAUWZnbfB7ftAyGYc4yfUpwL7w
lGge49tD0erOwyB/5tbINIZz415FkWRsZ6FvjLSgU8MadYxeq64h713GtMFY
RQ5F//peSv87UQl7+hE2u1cAoD/gdS76YCDG4ZsYZ94S277qwUSSrNVWwv3q
XvmS+pD9am11ims8VCfww/bJLWiX1OkQLD9mrvLExTuVMDWFYfOrLdwZUMxp
DL49LLmmAL3NFNxfbHNn2Y2ZVSigT91IHVrIYeOb9RFj0+s9e6UTObgAarNe
KspD2vODBWCXOE2lokB96q9rXB82qjFO0YZvdrGxPxoqBaVWn/lhDtgDr2Lf
SjXXKu2fwgA/yDWil/d+cHXs6IcFVVuyWx8M5nh36UTXLNaMizilbBGQpCAR
Hi9DdcNj6v1F3KUIbeWGvh5GhKIyX6Lvityu+TXkgghy6oIsyCNnwKb7qOuA
CedEKgrWVmIwJWDBXJre9NpyH4DVJb3TEV9K56zLdF3z46iuNwd3FAKpMMHY
uelefn7+CkALx1W233cBwqtYuAtQ+wwRYFOIUOEabnDlUzLFC/mUH0oDYXrk
KRJnCSljnAmIt+i4fry/FkgeknDnZxHeiyCYazmfr/og+ux73wwGj6olB45q
mwHuFfVbDvYDTfEiT3aoGDMAUOh/fXDAmLD3npI5xa86j6gCYqyVTP/htcaX
lws7hXd92fQRy74o1RbM3f+KjbeaHkJQWF2JGnmyvpNzPgv3/SeLuIXSqyFh
Y0bHgTxHkE86fP35+zr8D6VXS++lxN/ZWBWyx25MJa48NvJVh3pLLZZ32JCL
5Pb0ZMLtUI2EsdwfiIY6+xz5UN9WAqPayFoML0OBLDdO1E28kz8/rgu+sjKT
6WigHHkwi4woPlYmLevtqxkwMUNudgFV5dC5fA35GNgzq4UzP6xX0xX9qGrm
b6Og40bgx6C3PXScpl2Or6U76oClVNFvFmA1ZGqRJGdmu1Vlrrcg/vQFEcF2
pk8wYaWbwhwlRLdgeU93AfX/LUwhfchyHAVXzgb7LcVbjQFxkcYj2Dm2Xf7R
LabxNPOluYyhY4nvD7WavqJRms3i5GsVkZ+TeiFA87yTI8Ki5PIZ+lnQkidd
HfUczr+qGDbfVnLSx1UCgxVQSBxnaRs91RXFlC4FmES9u9w0HbvMl45wpbCG
HbSMihbnwXsTZBilGSGNC57scfnM0tHYLWAuuogZAFtQQj07vPlhEb3XyDk6
ljbAY8MSBnjCO0f3aVewWI9HvcwXVBqaiwicoidoojhmZxa3BnMZ1wF+HYTb
EP/xzDOGDboCpec2AaJhbBQK/4DZtv8mWr/uf7mqnykY4S2YthB5HuW2WTRv
2Jae6L/4fEBpYjJDgxuySVAwa08+1q3fLFggcqzcv0qC9XZMnhi4FDKzPTGJ
rzWiZfvjiw5U3lDZXfytT3GRZcQGIh0vSgCsVnjSklTYNS5sCmKLdmttiULY
nooytmn+dkGRKMx7TYmeAiXlykYuzxxYlIhvvdB0XxYK4C+t/D6SYFvOhLzb
nQHW1kSVXXIx0PjA2qwe0z46zeYdkJPn2oN8AftycN8QdJdJC64/7/41+GQh
GPfiIAIEeyzTamVrtqAn3ezNz/LgeSkZHweMj6i8PhaTUwqrp2W3K49hohr/
Auyx3CkTYwRc+v/9xvwH01xnKznov1D5pZB/JdXMk7XIyDVzFfa63MwiYINc
g2NWo4ehEe1VOimXnS6dqEwr7AlyF3vM2a7KQHsZSxi8JBUfhUsK37+Fc8Sj
nsds3P0yaYhLS+/I3MAXUGHsZ7umc1SJYMT/8TnkGGytG5Go6QeouozUJ7Da
fphNrVw3X09U9uGIFsf3gtKCe73SZfYYuMefSQHAgtP/r9/ZESoFlBKpnVqc
owLC8qSZd/O0wpvCCtE2WhOipOsjT6t1FTYl26O3zSxrEHzHrGrJ4NCHdSt+
iB25s1E4bobLNXgzAijzBDWWnwQT11odMdI4Omf9ofN0aqOXaI6kyl4vNBhP
KXbq9JukzdB1t9GNhrhX5G8+hglqpjjP2qgZRbzOAvqjNAC7PNqbLYzQlv2l
KbihUtjbeJLuBnwQPyVfgAdF0EQv1F1h/fAA5T6kTnn+319vXPcI+gh3AXpS
olzNzsVxjeFp8ERssm6WtF8RAAh+p+uAPvqDl81lLROE/yzc843cbpvasXJj
iFQSJDrXb6E28+BEMLng78cYJd5yVXDvjRWsWPNE5DxhN+lyEpozloAfcPsH
P9aKA+SMEQSGmN0u4XIKeux4I9GgtlcOGS7JpARqz4/Srh9OvUg2N79ShCq5
NwiTougj6e5nBCWEJUPPmlFCjJBNHGcmJfgivvHgyKaQOeZQAg3YGt8wp27m
WJPPWTDpfCbpLkEWTHV6kx535laQL2ei0WhxN6Vrnocpo8u3U6HZYzDDqmVf
VZM+Y+ieJbd0Tq8PhDWLBB4PWGQ5qxmOSblQJ3Ptqg0o/yoAqXpWO6sd6D1/
yVCesAWnVnpVe0m+rgglRJRstk+8d0dq04Bctg5otx95wOP9zul3QVMV+3SS
gOSNqUs70worTSgZW19qP563bDfniHD9Ki6juFGPwdUcnh/lUA5ygg1e18wf
5kdYecP/r/b+IvAVfVs+olKzRJnVCYRyhjnPN/IaKfiAlC1tw1djTA636Eai
xDhdJfQ2l3dEeLn4H2q3dfPTmugqp5L/pHDAu1UqcmvNwrIRtCCYB6fXTOAL
hCuihSvkJvUmlejQMEC5qAWIVGHUuQozo4NfzhktmTCg59+afj8OlANP9E/s
mbr3nPST8h4Z1Zfd73DkZdsCUociQpmIfNsdxlTxDRa2znS+/09xtAv3pXri
xMlfKknuQJ7xu8enLP0h+UfbAbLvMLQVv1KZ5p/PcNe4Sk3p7OkMZU8hGXjA
Y9t1VTJPPiUDpDQupJhvcVACPttTrCuCJWFsBZLfSaOzqpNWSk7hOTGCh2IB
OgGs0C3yhJkPRaB4JhH00wWplTfrlRGdCldMJ+kp20qXR5fLjyceJqdjRptT
TvG5x+ZmzIr2wc5mL+iefU0rAB8HUcTtE3lTaPxEVIC2hIKADQ3f/Qfi3c79
twivNRKHGqi4J0JyhAMGr7AIJs8LvfCpddKPczitOQ1kwKfX/LDV6LoODP86
RFDp/gdaANBFrMrT/sWdMZo4HDMr1TNsRq+JO0k0En4C7KueI39jDr5ODfV9
0ysE/VRoe2vokY9YfIyJDCpNyWphnD1uIkhnHlhfaEGXbdMaNV528dKRMy6J
d0ELr+QLZ40V9U/C4NvtBz8MelM1UykIRkM89X5aqUIyNP1gw2XUyFceRftb
2f4EXxlukkyt4qnx9Gzf9AeZlTcXjY5nRWjiEUCQNooZ9MqnCkxVjV/qGldH
ULZUBCvaLHfvjLKZKmgEm+oMaZgIri+mXbhhNIEFbue3Uk+WkC8F5OVhoe8G
fM7rGgbB6TNkCNJmK4nC2wR0Dv2mlUjLWvaPlUIwTl4Ftwdp44Ob7UTNLJYW
jCL3BJNYaqTGjCyphIJ+YHeqoftMx+qQff7it8SbEhU11jOyPErLvaoTtsKZ
dGgLFgATjST2FRHJp0gv4gEHrQQYi7NDEWp7FaOlpO3NEKgVFm/z53usl8rL
mJPk50yNPZQPry8QwqUqdq2W9dfSsUO75YMqcFBN4OL8fsNvRQEQRYpm6Y5y
4RQWKg2GH5YvGaAXDdWmxsD+bXF1HJW8zE0RRiD6R3qm1OLCf+73hKdIby4T
dMpHj1lyj0WdbttDxTA/4TkWAClg2BNY0LPLDdwGjOSlVmfN6xQvyikbxNBo
vMUlDwTcw5Iik9RTu8fMxDgDOuPj2ptyC/bW9gegvDPVZY503wOnBx1oAeyh
u9S6CY5XN1jdVbvXXx5qwmxM/9NI6pPsxCpPexdjdZYgABpW6WZjV0/SZy1i
042ZdASu5ML7Lm/IKHdzNZoD/8mzjKV1oJGWVrYqH5Rhj0BvLIITjcZfZZk/
yRgkEhPJALeGO7r1HVQtVQLku+zeps5vg60Q1jQeWNYIh1OY6363Fw157zZ9
Ik+TOrGS8dWby5n+CGADh4RACh2oybgSvk7dL6hSc7vE1/qqXq+/TeXQhv1U
KFPtEySPsBl1xNLFtpwnaoYricnpENv0WlHb4QZ2XhBxePtaT5fofKWEbIYY
D7dXtXxMKlXUkRQXdBacmp4/lIXa7zJBb3jmWm93XyHOW/0e84RzdTWn9emz
EaViBsJfi8XfR32i+S92puTFbQX9XYROzZ9iA7gMElCkINLME+aOx6EABZjx
KXZ1/4iWp4WLBuJyWgxKK0ZL+cDK+sTDCubxMUsKCKvI0z+7D9u3Po19IG31
fQjOfbU7TdN7hdp+1AahT7fGMWjztow6gk44AK6qhzOyrMeBTn0YRhPvp/qQ
dGBmmYJzM6NWjYnx1KX1EWh4J+Cmk+iIM8XSOubblP1vGQi92ypRWdHVvw9k
MlCkEGlUI4+azfhfNDclg2/iFzci3YBle/jZCl8hZSvSxam2r+8rJgc2tVRX
G4uHHK5ZMVeNmfbUyyZL4KGnotcgVQxCKIoFoOEN/D+XuhDKHAkRC+0s6g94
MRo2zaYuSzLvF8nCWOTCxlU0aAV5HrgpVm3Fi3yg0gf0SKkEjzh0dnkSwcDW
rLi4bKc9GQ1yJdvw2cmyjJIgSDoNU9KvKIsPbrlUIwmExeWdf2tRw+zyDDDb
corsS93RW72iBGCOHDB38r54Wvz/3/I+oKC2Vgmhv17goTPIVgQwt2mijbrb
WiqOHJ6TpceETOVQHpkZKwr8YMn+WOZ2YW4P7un3UpUntXFcU7WjBGsc3/1/
WvZQz5YbXNGYFDdXI7UhCrMXwwAn70JrxZuu93TncI8dFruCdN8O/Wn3wqfh
hCMk8zgcLTh1DIeZbxveqa5lw0xkIxCxdOK6MLU2BE42OHMDhKiU1q9/PIFi
R9nz3yCltC7kr4kjCwSme8d1sk/SJlIyTk/407Sg/e1osf7vfejwt3JRLiXd
mCUV/e8qcscs82RkuiEMGZCC8JaeqcKigvDIK1LtxXl0gw9mieFZao5CPKMj
GKWoxsN3X/CnzjByMWoSVJasMGMRJE4tZYIeFpGinIzkcZPej4xPdSjjrBkO
GnXJGGBIhN5tFQ/KmVNdhKbhFv04sp65jJVuBRH/Z2ElPtbBTYFEM7Yuncc1
RVU0QOX7CHiGVEPzJJ/oqk4cLvGMwtgB63FMcWUi8pyH/qVkiIKzcYGrWHjW
7woGPYhK5NdNBuwMLOzgJXD/bLr8XW0pC+VzcHZvKhdITBafgcKjoWoM+nL1
lzhXMgvqVCA8NHdOzFszDDhoOyocTOOICxLrMmOHwOgcnvHRJA035CDrK1WS
pAKhGW7mipv19hwUUiPPYwvJXd8J0Gg6Hflhyzso/e0u/qNUEj4HvJItU3AV
g150bi/JaG70HrU72y0Yjxdn3ClHDGCQBq5X3nF5/sfw9decsba6WXP3vTVw
T0sI/kdyp++GrpHy1OEh/FPZ8k80UybRLtHH3WwBdsPncIXKvwa/YWzNMvZx
iL9ecrBrkkfSndyf79oTjaCajK58BpA2WGbzubxn73C6YNhGVtKmaIG9J+rT
S5Yp3clujT/+heblKhSLUWIYXG9InyifVWqfYV5e4qg+5O/Dk2Jdz8V6xSSb
1H0lGwVWWAMFk/iAIRIBaoTpMkVYg3oMp592qjpvnNtyT/0ATMz42F59p4b0
WPxbkHIybl0iz1dLXZ2kgaiSSB8Bnoex19sit0JOaiw++rWo6DKuNufhiBr5
522XtuWjiSe/Mz+PDTNRKtvPXxOCxv/vHVhg7SMB/ajTwD2OXQPhRd7R4BFr
BiU4zoPIEaGZIkKtmh7rD+ybwLWE6LszA0/dLjgLD6Adhg3Z5u4o2YKd2Exa
AlxYnQUr8+zR9WXXqZ/NRRLfb5Y0FtzNcUrRcyMNpvwWodzg4Ajer2Dambb5
Sx5ZTPiUogLY8mB8yBLWvR4eRLD07txWsGAD/pITzxm4ENNgNFSdlGk/y1So
juFt9HfK2+Eapsq9r4oj38TdmB6VmIBQb8jCsXlj5s9RdPFdpt2UtNztQfr6
o0+XIlAfxfInt4PPVacMrdNKnPZFO00cl8LHRBFyEoe1gvuO8ie1fLbFAcqJ
c4/kdm4Y2mersVYnkWnG8wN0UHNIwWEj760moCqrqlQOPXYq+FF9b+sZXxxF
YXeEyPLWwqm0Fom5RKy4Rt6OJM9tZGVSUPojoV3+GRo8193JoVsYSh1Gflv/
vwIr8wSKdcu/RspgKuWhsKLeHHwrA1LYD/I7K8sK1Mhk3tmuC9Vg20stvw43
qzSDiP1xPvdKRglFuhffEuk3gSyhUBUjbkGNiE8in4Eydx3v0FaOQUgctz4N
M4StZMp9F2fl8Orvw8hzHfqRHtfzFNxFt+ojbthvUOF7tZRyzbj1T6vIEfwa
VgnVNgwWSk3vqyyEsD2eyBgE9Ruw5NLNe8syB7fYMezdK8dUlK0UZfvHWXHG
2ee0O9qtdKSHcnXU0wzo3S7iH96VYWPvWy2+2IjWrckxkKwH5BEAVwoE44B/
0PaMa8bk2230q3yeSI9f7LPuziz+lUqeMVy3pugmjRm6HVILZicDBm5ij8sz
HnUyHVha9+S977NL7YWbjozZyWBXv9rvzVn8AYb9x5n3NBrBqSOwNUtC6Xsp
bXiienehgV3jmFMg+rEb9uyQwbRz1pBGdNYW6Q1Eihb6C2onLk3FBr+dyxS8
8fShgH2EJ7OrgeKrJzPeDO/vcbHqqz6oTiC5X095NvT89T77I2izKDLZ8WW/
wTEzEKQCc8lMFQk/pqH7StCNSYwQUAmuN6cclDVa8xcKV0/CZLFOsmK6HXTe
iJagpnQRMF9NFiQvRi3z80kbMxk2NpM/ZkXcru1+PkTPCS/9FqF4BJUuV8+s
KhhYKvzw1S9LkKwfj+FReV4EVq5n7IZtSxMEIQUeYHHI5hKlaaUz9R+0RPcT
qxUlM/PW4YzF7JL/f7jo/LxDaNZGXVcTNJD/9YK0EfI+Ntcz8pqjFVULQEpV
a2QtmsId17xVv8mHsMqhPeJEsBmB3HE5S/6wncmRlAbKCfT+agR1FbYwGAt1
UONCyDUYQiaTaMMP0WHhts5a40rhxuanmo1cKng98e5MyuHpid7mXDBvXfcz
Y+YeoyPozUFy0N3ycXnX/vnRtznzULFHq0l0heEAxKzWjmvo9+Y2AzT4omdI
MGM+bvqWE+ndQ7YFTreMhtMOdnEm4XcnJJECz3iKAWaQbBEmmVbZeY+Qn7wS
Z+lFwElYvqhCO7iY9QfnhlUfKfm2h5gJxOgqqESqCRJDbJRr/P4vieMcyKo+
hbzqr5iH94BS1Gy4+5e24uHaACkRzINwY4r9jYnJS8ERMpQZ/xqO7VopFHgr
0WuOPT1qJXnQVjTTveLnj5VPjLwEuAcrUTt/6e3QNsNKQprHmsukXKn+yJBy
cLI9m2868WWvlSA/3qjeNNY5kFJfC+SnBqQTe0gZz5Ng5y0+YHkTvCRpJHeb
IQ7RzFlr4jW415j/5wV4vcuWhHeNa+32xpnB1lLuRgi9eUajrimKMYNTxXop
O6GEDxG7eAuYs5wvtvIBa6+EfBwa9CS8hiPM/M+55h81MR7Jn4DtoT82M0Hs
qhqkg9HhCxnADOqVUvnuwxX5M+aLoJBLUz9UHf6RzluWQFI2VyW8M381rZc4
FJf52HhVPjoE9gUhTRdWbbYIFPGFGXGLYXCicW1x/dHxpXhe01oGtm43UX+3
/cxuW8iCeaHhgKi+L0GTChUgsKnLdGcGWhAft+lKS+j3jkXxmvoL25nv3w1f
A1+JXZXxcmsGcEbBopWfsXPPHDsRQQpgtTiK1QLj9/d1LaHVk0tlbvudcIXk
BZ9D+KG6XYoiH/IpUYfmI/lwCi2Sn52cR/vyoqkFyIrUtVM68wPUOFAzOJzJ
zLiDQMr3jKTAWkRtF6DUNYJFiqT8RvXTRAj/PHyi/YpGlTWOVagqXs4ggHpV
6E3jGD74/YQH9SVYNfR+99jkSPoJ18YJevz+V6FGxmbyxDzk533iAG4gXOBW
tfnRyzu74JsQmI0Sc7NIE+ZqJkfybBqG8OCD/S+1/9WpO5TVbBvOvmpeRKjW
QGOrpU5tjFjnOG6c8H/RXd9JO9u4DY55Ed/d4UmedBSpPZHBCPQsZt7IXYp8
fm92UnTdbxd9jZBZUyRXuETJ9O5JaNuVo7GBqMsvQjEBjHZx50e4ayf0nFxI
WENrJVP1WU2NpgZpgASeMxFLHOBsY5s8MVjYLBNBUu5zacYOGtPO7JoO8Rkt
S2LvAzn2pERFFuwU0BMT3o0WkcprGGfKRzCyMxPb2AoyVBixaviOssYGhI/a
8nVBxCBBha1r70BaTq4CDLZtW0lv4TYnzqKo8f6fGJx0PvKM/shEhI/v6RjP
icCyFMgWK6qp4P1Ja3ZH0+I7FyBLNmHgUvWH3DzzdFwaZOR6gTi3lfrELCcH
a/Gsp4E3PvdmhIpVJVU6p6w3086fsKnlJNObpkDMXswUwL+r8migzeZK/gIO
6FYTdeH7Jlkl9LoGjDZJsoSRQjobJBA1Fur7v4B21oJq/utLm05i87nWMurG
5ukQ3eAeYc2Hp2tc3H+vCf0GBVwjFpkJu7RzKo4FxRXCVI0SKerK2k8km0Qs
/OcCDB4a50D7Ef59jGJe1ImdjrYksrLLlBaTw3XdVKaqNCTCG0fQkfa1viFN
4kKHoLIpj4vnHr7WJdaRmi6GSSZLjDvY/bCMBtd6rkjQu7wdFzvWOZBuCTUQ
QKALryskfOCVRBfY/K1YUMzowuKNmzoNGAHcX+j8a2cFKFWVPkzPekzlJ1wv
nVCLNXOk7bWRB0kWrBFyI6TZwzlXrR/wZwvLBymNaChJZysoBtYwQgxD5R3A
GYNHuRJ9VdIF5wMLwro1AxBucQeGeBNJHB20NautVr1J5Z2a3yeS+n16/jbk
tpn//Z4lpF23nKOHnU46NxFo2sM+3aRNN9Fwnb3dcDtY+OnqqEgIHHmJswar
KE7vYvPngjjsja5eOvlEyszvOs9FSs898nT+bHXSymmGiSCrlxSJkvRAkrqa
lLQQL6lB8N/13wkB0JFO6nUvmI3R0gb/wu624BM2uTy2qUndSTZoNBTpCcl8
PL3fd6aWQs0RlrULLRqnVCU4AciZ+U3W5hzylW2eA9phseIlmyZMbJM3rR/y
t2oQFgb90uRPw3eQhuWnHTycRT32QymHwXhsiFfic1a4zrJYkxem3VNVRKis
nJvXWo4oCM1YU1rr1k89Lpnp6YFJ+323+ueGc6fwiTcjXnf+zTHP8tXaY+mU
JEf6JMAofiYlmnJRvSC7ZlIC8hL9ispk4rCsH1oyWw6f12MkTbnlJ19NkdcN
AQBuH1v5ZIsEWkKSn+b6BX0eIP1uDpwVXZ/0Dj58eDNnyldaZqH4gYaiIQS6
Nu1IJ71to3VFliE/qeGIG6MN7pTiCZRzhfUpsmCbRih95tG3H4QJ/qAii2ip
eEqoh+Ank5ohIwaSWbWZjlsVdXnKzjag3dxes6AR2kQNV1zFdE+Cu2g0ROWg
TI+62UcsAhEwobrBFEir+kZyNDHZTZbPLD9aPqPEEw4NZPjZGzODKf+NA5LF
ZIXTLy9OGkUj7viIhQTSsyUWoBh0wWOqKhIXLuDJCABi0ObRD+xTSU+44zT6
9DWGh314AM7ZtkzKEUwk/Zi1ts623M2qS/UpX8/8NyR7v/B/9xmQ7U1oh3bI
MbJUJOlj3uI+3rWRYIvpAnd2kV/vrt4SuxlFofv6R8QnQhVYGSgrBB00DImm
1wO0FB0NAzzyPJ+SBMgycB1jVu+sEKmCgpnl6pzGyLMm029G/+FVOhPWfOAp
SLuswqx0ftmyxwexzkq4ujfpXMEiwmAgKT2fuCSqSachDtIYlPOY+zVn9dXB
+VS/tAptQl31FDzpW3PBwo7LVcTQfcsGEJMFpl+/LizXTKWBkcY4cJYci5xx
4jKmw4nod841nS6CTMHvpXmc7eVLh/7uqu1AGvQG0W5AvVj2efUVSflMEM2O
KB0FsubuQsqgN3VkTWl9Bh00Z2uKVibBd9pU7nPrvfM0OcvQkfV9bHjyYTSe
AKiMCdP0l3YP0GRxm2Ox19yC2StHk9Mkl3eghHov63d042nS3vRF9hU7XG77
PTT0z3R6s6Derh5jBuOfZkD12oDBk+6de/GXulDqRBVIuHp8P4LjbxuMnJ4t
AZZ8E8dkM/tqsESUhQADzWS7V+wH87ms5ahASK0HrrvOg0GgamKISW3VW6hH
7LscU/ErJLimSEGmVhQUPAM7w5GNWarGiDvZhx0dw2nEBRR2YFkYGuhQO0F/
Yd9GkRRvRGDPHl45ZKlAFYM5I5PPttHc2ttxlEXg9v4wNCU6GpelZz5uf4lV
veQBRJ31vk9F7lO1W0HlP5kIDiPI6Jqa+vjbmm91TqxFKmqNL1VT7aeNRTfP
4R4aQrJs/frMg3Y+H5bngZ+76Qhss2ic/MhbaDMYx4cqrvBgPMPNgSPCH1rG
bZIy6opTNdbUqswmE6jv4FDZjgcBoxf/HWl7T9K8QaKFxuoXEVjfY2cEWVlf
KDTY1WjFJhFRm4dNU6PtEL3C412YQsQy/AOo45ed/JpHbx68O18/MfmQmw9h
pp4QKd0Rjg04xPxB8jqXYWQnhimNY4EuXKddHQGTx6V2WRf8xTuUVjmnoJ1j
NZsA8z8GvpoQcZA+IojUb0Dn3CWkU2hS6tEI/jHefxgwAGzLl7L0w3/q9QnN
oy/icBZuPCG1/c4tdFxGjwCorK/rx2ZfqqbmaFIHblGpV2gqCBIaELd6i7Nd
KBPQPp+pmjB5rwipLquZsHQTfR2T3Gnv0+JGOoL6wSWSdV5A/AOhdo8KJtL6
zgNptqGYUS0pQItOtuVFyQkKdZQ17d6igTxGR3JzCMGidMcuSpfBq3zystsu
Fd+YWehm/Dx40NMuNidLMeuk7LVv0bDBmPTcB7N6oLIGnR5FAJguhPjZ7dR7
qiWsHfEl3NVpYOpGKhZDgNrFO9TSfZMZ4efmiLs4ONJerDLOLVMN/Jis7S9D
vec2CVJHrN/0mbg8i8GJ+jTXE0T1jzloM+CdpAV74X2ZVnLOhu1LwH9KX8C7
6pbTodt1LpV20ZXufKQY9i19rVbkHZQBYC+cP/zCq5NK6uijEYBUmWVp+Pyq
hswjz1iwPSxKBko+wzVS37fkGYxvhO3LcLMD00FYF8v/M1hAb1x2zTP0naea
cyFV5oiHYFti/2M5xMcmqkpzjYqCrSb6cFS79olABDsKo9Dpm3OmcxeV0uIr
lJgfbjVryxugSIDYwHXVZGtjkJNqxDTarW2Zw1FONrF7o6mVuLMEvKqrXN0m
vLfAxqAIB6J6N+g9XNyPXBncUGKU2ALtCwaX1oQCmKfMJFdMOt1f4XgKxsPS
waAHArHwOoZEVzEeNuD+bdP+ev1y/G7BANDlUE/TyXhXwd/MLNr5rBDgcpxr
BmKrTs76icqvbqeEWA1npcwdYNJA3OUs+FNoJLQCWOBNA/6au9Ol87GeJMnx
wS6fEPsnioPksrtMd0rrxFXYkM04yGXn8/8ZedC0HV8cTik0oWQUWydQWvvK
PXfGYKcIMWtiWT0y1xlGnPl+swJujPqmLP4RqgDmCJdSkNJg5wAkGJDswV1k
OqyvOuiC423aldn4fSqOF4vEKPIDIu6kxcIWimy4VVGtmVmqlU6xLZRKUgHR
WmteYF5oj9OQJO2/dHGzNckz6DUOxAqgKlu7iTsg2F8WmGiJ4l3AyhA9Sjw8
SfG27rZyEBW59GdCL8r1sKZdLYJGAyu2uYKqVcl8qAC4nru3WkL1hPz7/7jo
rAvUYwlIdyMhlAKzJ1zSrRaEmeH6W4VKlPkVwSFjDDEcAzge8yTTDVoeOXoF
Ncko2+fxff1Ee4gBXC3X83CKHjzvUjVlXOOCVMyYlIWYIENFg+kGfFXXd1A0
cKayuWHXUi9SRJ/637tOsghiuwIDmUuJ2NvQ/zEjRoEOzDX3m9318GD9xPIk
8sjIPjxFH+fhPNdteA7zcufeNhGlMMELrnlPMsszFc6BW8puO2r7JcOnPBWG
TPMV0iAnysofruM4p9jq/DN1We1NofVTH+YFhanb8N++RIa3o816A85LeX7z
Ei+GPCe+e/+2bRa+Z97vyW5AMA9O0Y4M8rOYC1M1gE83q4l/1LARLK7vr02Q
bcOxoG2u/bHIr+dbtQOD5l1Ekc6FWY+A4bJjl8ihyzTeiMLlyKOICP76Ldye
QyDLpmRbq/RQR5Zlwkl2+KyyE8mhoWZHgn/4VD2w2awKly+0+y9pbWiKd0N2
5QEDD/+J6LrJrQStzQe2nnWlAMOPJeNtbCw3AACnPa/5aoP/8D7lD6rVBY5R
/etmDFkRGPI6ol+jyAxguGwAaUvdcNohA/8tgI2bUmgj1zcIL8hHmJ7tkA9w
t9iQXyOkovXmwBCTt6R7tLKV3WcI0NQEfN9LhEZa9Ylg5PRobAg//p3kKeXc
iQq0X2vi4ILOgJJUBIeJ0Sq/yxNYadPOAjTINmIBaU3U0mghWqtsk/9AS8b6
3CrDg/O814lazb4DIZAvPvqgMZdfFv4uif7lbjCLacIrRK+u4b8VOpMWnh1u
nNYPalJclDwN0Ll4XSpWMVHnEe8LFATj9idDvevMTCAyvWEsV+XFJ/Q36bD6
O2XJkJCSUH0Wp1MRNfLjLBrqh97aUEVWRf5dkVUnDsVKjlWYuyaecdi3FDys
+vEG8nuA/V5mN1DYZihmBzakMqPJea2u0ZerT8uALTZ/c7h+OfVNmCAC9mV2
muqJwSH5xl0ERS891+BoSWp3pGIfti3qkeAPV/JCbxLV/gfas/n4KPhz8wej
C+7knp7v83++q/muTBCdvrz0ppmsnpH5UlyMLH1VldiLbaBvil4SlS0k65Dv
LCJ4USXbnHeJoaRt2phOjucZMACKcE4CPge+UtXEUw9Qucobxv6r1eQEmzMf
KSy58oCDOoI7YpRtzUXTlkDv1NiYp4adJLxz6icrX06e+7yE1+KTyBvuaLig
9HZC6pxoT8l1gbv+9uJyuXUqEKwtm7QaQZWRGouI8EJZsIkj0D1+Dj4+h0aU
CqYba3LgJ7N3Q7g/ZaKAUiP1bnOCVeVF3+lLz+thjbyOpzDQFYzD0VLSFWm8
AfMXCAruF3agpHSWse1v7tXk51H6zZLA59nF7GKpfX23LkxXPfi1PyzrNOgv
CargVeW/osOU6GS1givyRsrTKTUS/Bu0vvmC1GVd2hQFeZzRSmfHhdYSaT+R
ry8sw3iwXWbk/VX47/5Az7EWA7Gfk9nohB9TfYPfnN8XziEmXTGTvbBZOjk6
OS3foEwVyC1vmjLY1MQcmODqoXzngOdoJj4V15HSUFDKJjExs1Gyhebjq4SI
Ui83SChVwlK5LxVOVE8uybW9XayYBgoWps1tjoVSoLyGmhFXxQMS4bpZ7nYW
fLdSCwVpCJt0clvdJ9aw82zPIYe1/UmQqf0/GXaMQVUDmlhgQ4l/NWCm1s/G
ZavqHl2X6QhyIlVcEZopjjTVmVXB7eFIJbZTCNHYp2f/gP8x+2Ucw68ySCWb
ZYuarP6hetOwRuCn+uEKHD1aA5FHDt2LG4CkyTURZJYcf8Xf4HMpN0k2Q6rl
xldrgcvoUOx0bEXghbekWeiHzP62MuampItakRo5Gf6k9WqTaQ6UPTnQtep9
Ki3gwfu8wuwCz/h0n/jSW+PcaTK3qp0J6S6Fy3xgl1vZdpm8QR9z5LOnn4rz
/ugcVvC9XGKBne/RW8hM8RyqQT1+6/SeJKTTAZdvlskxuQ18pCFieL1jUaZB
lX9/J+ujaV2SZRdybCWG2SZ6jbZ7wyXljoJ8SwT5vPZC0m59X6wEhJ9mbZVY
YzO+ttjAZDTtHxrIfX2HTpJ0+hxPbIYnO8v2o6tx0eECofVzfuIQXoFspgTC
vlFz+ZsV0PzEz7bZcnRGdxuIM2/Nv6oVTffDIZEXwrUu92YB066H7Fjuaey6
xplPxyqSbfFy+GtdgBHGz0rQtM1plmka3oetAivxYZE5fSqj+9+aOBKyUJkk
tH/UFdJ2gk6rmfq0IwVYCVvI3O7ZEMuzHJGsHMVATZYBVJga5K/xRBABGGbX
Fea6Hz9jRbKcAxHTEhzTIl0rJtGyS5wHOMWhvOMfgb/CgkNclQNsLqNU53Yn
J1g6fp5NgGgFWXMGfj/fwlF+FNgFPD/CUeG4awC46WNtuE6X+YF6Lpd0E7Nu
9Rhd6F06Srw9B6M5d39n8UA+PruN6w8uIFUoK9GACIopJ25qf7tSgYjy6Hsu
oTvR2kcHE6fuEWh81zma0B7jEij4iHvJPnK9mQNHW1397jQbtA/fo57opq3V
/aT3I02xRAxxEBXpu79cdLH7Hf0XhmqW/YgXHElJUEgn3XYTumSGuN5yoBuW
mvX5tyoWATDe46shFAXwPJSRHB/pKpfMwX4c0lAGNJUTpOjOG1uQ7kL9HUu1
BKkYnV7h+H/064ncX5iYdawLdQa9pXndRRgad3mbigNMp2G5uqXekU9+OryA
dwz2V3fjGD1Iq2UTuAjzvrpiidQfnbANGwuvP/FjUONEdw7NOURG95W6H/c0
41dswhwexyDhVqpPtOsprQqTJslxCABVWtcGojGRYTg4v9XRYbgjbDgcp9d1
s0MdO26mRU3Rg4O3X6TERocr9coO+pIp4zU/lfIW154a3mihlsLbfGx6s+pY
V6uwBbyOyYMPwrSWEMwLWCkvOdy8hKyMwHvBrOTBnYTLCDG0TeyM26vCkJYc
6Nw8TMplmTsVIL8v1VoPHoxlPl53G030yM+ozObtvUl0lNEB26bnMwWR4XyQ
ppMC+EJ4D3MHvmPQCglU19H8kzGLJYoGKrpmg97SMu2ZOF1VnPKINKHdFe+c
IWMLDRz8BEXTREXUxCB4XiAtcpzuzGGVOSYsEXWsfK+k/bj1MnLZ0UhSc9/R
l5SFWbUimZDP/3xjh4h6gOgsgItjyDQLAxMS/wqdp6ExGfczcfzgC3exFvSn
VIlRplBmqf/xlM8RCwXL+HhPFQDiqVfxKSk3UaCGrZDljIRT/zSU0Pqyfk+N
hPhvcgPleXTo+q9IILiPsxIhPaVJg9Kb82yzPBjCZD+/LNAbFvQNx7RMfhpN
JNlW6R0FBVlWHXhI2Mfd+H7XFvwor4/H3o+rRYpBbhP8JL2Xh98DLZ3ruf+l
nLFHscWqJpw6ZGaCbGT4lOra8KBuImGrEPtbm68jte2B+MlIQsexCXjzbUj+
ihzb+PUwOwHadXYKV8f8hjGAiNUMhAeeKz9nfabHMwhrAZgucsPa1kX7raRv
Ik/LGdSIG89rrPwxYZwTIMOOZbXkCAqN08n7hHqOk0bxcEERn9SIE16NiHUx
FjL+If7/RdFKT2Bfy9s8hSc8abk84d6uFySatC6xvu8PMPi8bU/H5NFtH927
b/jwkqTG6EP8rK/dT3vry1FZ96D+CdpXGGk7nPANz7Mgkv8HTj/eM/YCEo+w
Y68ad5G3SJl6P10trTFtmGeZnGLi3FBSljkvzOqHeN5OXrfHmfXxB9oHSFns
jGz5yBi77qkT90UVW5Moh6mEOKVlA1ITgAXtxkN+NkEdWKTiPtNUn/F/VQzB
mMtgW7Up2Tq6KlFPGoUV+dVnJaiG59J5An6v4TnIsAMKs4TRd98tN2ZnB0Ye
2QXJa+hhOZ9TneJh/yPpFyVtIajdJU12589CFtjz91jgMF1vtTdwjuvp4h1r
qtY43ExiYqCTVwVcx5qjF4sEJ1tgS3JOlW+lDB6O9KrAA6RmzEXRPNflpyKW
96GoBLqdw76fjiip6jom3PUdhMAjjWSdcnIPz2uPQ5hi5wJiZyb1vy7Dq0H8
/3A5rRdc7I4c3PaB7uZQXVQXP0tiYAK5Id3fqb3MYL+BgbliIznPy8e0J7rr
iYV8vzXmEIUJuWGYrWm3eu+vAgkMXOvUSzkOfXU2DIh+linnueeOt3tE0Ab/
8YPIkW1DzCm3IiabrcdKQZmDU8nj1j36e60+mol99ltrCz/uivFB0McxYhjE
XtZnlM3GAxTGYx8VdyciLsXMgZ3b0PaKRPEtAaoOdWNIlWthp9HxO/dxmrN/
whWHTM1uWXcdoo2wytIAy32tsW+NDQr2yoIiTM+DstErnbgwGAftR5yFlAZx
UwNRXecoKIVG5xDKhBPjJedkaThSeIsOs1wJLvNGhyXEIabU6C6PEtL7PJxB
r3sdABNu9Nx4gwpmByFWSsPdntEKBcb7TJcuycjf7yBLtgwARNwlS7HEJSUy
WivjHy3CIoU651t+owLx3dvKwjNFlFNXAzzHaTOeAA8O4bFkVAZ0UGN8X+Gt
q5DEgG4GQJOJaxAqsc/5MHI37czDB/UBEGpINToJBKF4szwKom/9hyR0nXVe
AqGrmgFxywbn/4Pei+odLnM/KcSwxfy5IQp4s4VbBMInzvB1mAvRle3ETlI8
ff2cBsUgwLF7ya2kKBIQIfqMEXuP9riGPaMIIj5milW3+HEWUcsYHYSa43dL
1v3ftUo3bMRcZzdtupeRne9xJbnaZZwwe6I+ahbaRYgkyFwttk+Fr3Vp1J2U
Q6HYXlGh2lvIDeVDOWz9t+vdVQoUnn6kpSCb4K7ABH9W+S4WOLp+oOhAUjFd
/w7av4Asap5thQQYzs7vPvrTYPGc0QsBKOXLTCdS1Nm0TA8BRD/92uAK59Km
phcb2wN3L7w5ardePWCXKpb3jLXivqON1KRMzuZNAIxRQAi844MmgoaAlrQ6
IWLSVxtcXBReq2GNQ2TD2WIn4rtnUk+NDZUOMiHJ1xnIO/dqaIOk2UrbdEFg
XQStkrmkhfGfpLG2ecXu7Fn33BuGX04iT6U4ViXniWEonKtO4lWgYd5m+xt9
bQMKuxzj4ThgdtiHP9X/Q2LVtxddce4Imye+MsYK3G9GpN9/LgruH3ClfCoL
zDHLNIyYGelHp9daXRfdesVIiT7c8GghTQCqszVoZ66ltqljTEmwmWmHfY5i
FgXoAd8pA5ALlj4VkV3f8oVjSNpXAp5RVjP4OYasieiITCP5hOk+2S47MG72
a5RN2tRIr1HNRfe1M+It7xq58GRdi5cyg3No8tzsGiIF5Ddi/M8ypfIrA/2R
fzVc7b/bAabj67comWc4AiD5gkwo4VGx2NusoMhiuNjE0aiTOQH8honViIPW
accvxaKGL5eKaPThnpVLopv9CTHOs2ZYKPql3WZXnXRpCrL1Z6eB4B7jQUce
HgzaoSot6cnD6Mv871+6OhEsCnHHQ2eN+eCHCZFTu8/RjVZebpVj3iRzBwXO
kb9sW1zUb26FBiVTsa8qH5rpJOjvEAyY0bvlDFTYzPwI+Xm4ZKho8Fvp33nj
b3bDLhWiMp+KWLb4eJm7z/MQ7mEMWzlIJ3VqIFF1id4dh7uRqXjoe/dsazs3
DSfI71DKO40AIUSOMNtKe91F0Y3yH1TcXoNVOzXzITiEbAhGxVrVkf3YBMI6
reJIugDfR4AYpr8JxrydXaFHuldkC4ThEK+Gv+qYmRckP7qFTrcYcxo8MiJP
X0/GeLCvro/esPy6FjAJUYjH8QCgfQSe3P/V6Tz4M2WamM/NLFOSIamynNvu
8t6ZIheNwggeA8sSsXNXniT2HDkiIogbuaF4/huYEzb2zl5K5Z8DRNta2sw3
0mjpa6aq38U8ukXG5ZqL7DaKD4EDbTMfzG/LgIuaMixvTTCVE2opvxfHnX5W
Rb5I8eJuabXC+5MeX5QLPwtxecFknPv5ssAV8YApZ4YqIs5K7dhlz7W/8uxm
BvoDSG0pMgDyAXvC7Y6zv1KYuUcCQ99XMfGi8ssUAW8HNTHrpqPiPttNOrZY
vQ/ImIBv2QzMuHkVgTAH8yg8qxeJXcT/8Rsj8glXaKQnukujzs2onwki85lT
8PwMKtv3/wWgTaL6EPYuRYD7ICE85gAixlEwJsz2s9CaG6Di7QNYdiGXmovy
AzBc4FAUsQMI5LzVvhtTWyS1HHpS/3U4h7dH+Eb904WCg6zG8PStIqp2HNm5
tU0X/QxNH5jFyOuRMdYIZlFTQ/pAPG/iZbVmcnr/uz/oaosBuWf828I7UpEz
+c3mxw+ZrXD6TizzEiVQ8u+s/yDuIVe2iwdpLOIROu7IO+SwqiH+yGvfrYRV
QSV4+I6H3ebVLgmbs753/a8LUGZWxB6ZVOUtvTwFpVsGhreiZCy6N7Qnkfyl
TkCfL3AfLQRujUlkEwEAMxh+Ln814urqwK4Qbj3XrZi6+f5JgpyH/3sAlmGL
VG3SFmOPk0O7rLt7Ht6aPie6lX7bfnW3qUzWBQA27msRlnkgZVYptPDEAxQD
E6/LZvHL97veO0DBHOLJEq/QxtfrCTEzMjzSknlfsOQPJmrpFDgaywIEE5Aa
V13wy+Kitei0XU0HYn5FaE0DB9zobTzWOe6C8sLQeTCgAwBBSvKXpQLhBNRn
PwUVbn8mBw0c7xMb76WpYhzzb3NTDSkM3EQIUlpvd0O48uWcdAWob6Xo4awh
5/DHMFUUtYKqOhRIjYJ0lLP6ajHJvT3+cuLl9SzK4HyyOfAPLyk3PxTafN1a
OxmzY01gfduNBT6eJui/6X1TI7N9LTUkPL4PBIdI0k+X5+Xm1QSSxx2vjKPg
pLFFG56LvHrCqS5H6cawpZqi07n6eh4I3rea2ne7cZ7ZBk3sXGwqEy1X9JFj
QWQWBptYPfhw1KJMfwfnpg3zV9+fMdeRH8qbhFiMHmxioMpbKjF/XOipMHuH
gjX/bj5Djsi7aH9R+9i9xZsPSC1OY6QHaJNqkVvHMCzRXgu28NagiV7HFj2m
CyjzQVly/Q2M/ZZTL5OjnSLZuGdOayZ3SPOHHMv+jw2WEmOukrG2OJKF+oGd
zPUi6eMfbEjjlA5OvfRKaoXVRs8PPnB4fKzg6i3kuwG5S5LTTdQwbb+ax92X
VCw3AO8kD8xBOc8SQXTnobdUJkS1I0714IGdJCQOelozuSzUWId0zFTKP379
PXG6olxdYjcvJeBuekwAf0sediQhTKRrzioLBU4IopNfeslP0VHm8P15f/lZ
s8UFtqa+nugot+4kMQGg9cXT9xUR0ADD37lmajpWd9RPDK1VUVMx7itQu7qP
Wz0QIDjAudNhSfIlZvcF1MZ2BcCCryRWkeNgNwGMpNxKD8/4Q1s8qEyb0eeC
A+4LwgpJhDJntMh3Cmz1EhU0ci7V9zajg1bFtjRKF862r8NqpHG5ZuTPf7Ze
9ZIU1V0D88UdNEeqzyewC8DyTf44KkL9cPDNEkpGEZs42GMvFyToUVzZ5FRq
Aj2AFyxhMXihJFvSGphtWxfpRo612FXyMd5vxZG3Cc4uziUERRqBeER+LMd2
IYQwYmTFNtqc1MFTEmZjPa4k/Kl5YNoPKCel275Oxrrjp+BgBMNw9hOpu82i
ZqyAiB86RDtNXMao8ZsHq2eFUDY2AB+kCR6CKmbwXwpjw2L8tDJhEyR0wado
Rd9gEe3wJ9cIAidmuScGABu1BAlSo20TlUuwM5/B8eiM5QSexFhOeW0YQWd7
Jpx73prvzKya/oyf4MWwW5/h8sUpaOw+EYEoeEVRzvg2QUX7mo4o6tBh257y
qz/3OnhTu5G7JJH0NJptrRg0x0S043pHx9iqLymvPf4JX9gzjFJAdQBduf8g
dGbz9hryOPV/uhNoWpUpsNzNN41dLs3z36h5YntJT9o/8szi8zWppZ+rL3iY
Q94tiPRnTU9evDYofzI4BgCow1BxXfPkFArvdKksM/9tMCVqbEodW/E33qpT
kv8IibdgFc1UgrRxYaZctxVsjA6usWD30BTStbwkZhopnytgfp0ZVxpZ94ac
8ESmQOPWhl4nXvYmki3a4lyBZt0KK71JTJqC5DcFd4l1aX8Mbo49rfaPwEcH
5PI4e/zOfozogl9egsdX27rBSYoIcxg+78M65HnbBot7jh0xDyBM72n8UXyh
1zqLxyNPcH4VhX4rwNigdnQk9SKbI39gDx40lTvcX6421yQn7Axh0/iK9uHf
GgLRQ3dFRp42ucx9OVn70VJfF67sErLFSEUidd/AH/7IUq4OUktsoNQohOi0
ZhGravzr8tBpyhz50FSloRgjpP7XyueXPMUlv6ynPj5T12GhQ664twrUDTF2
RIQiEXH/UEn47TMmEV5CK+wmNDY6qdP1uMghtPt8oAnE8Qbw73/qpyglyrEY
FRS0MhSmF+uXWFV4lrPLvg9uLjoA1WMvk78T1VQMTYlInhCaFldTFwiajwYL
ERwpMa5CIRNYIwivV1NwNueH7jG2M4aX6/yRuJiRtNWsXMGO7ow7ZorzVFHm
73Evifw/0l7M9dil8sqXUj90auXrVuVh/L6G5aJcdDbhEJ6M6KIZYFk22VD0
Ez37JV8f1WSClhGeYjaYNVX0t8icQ0gof0JXNO0A8sfEGpJOV/J9Rdvr36MD
LY761D6K789ei9WLyfAwA7Z1iIXU8hcvx9gp+GRFt4/y6jV1gf4B27Ih6A7V
jij9igmC0+Bqu0MPrBulOGOg0Dp/u/ZQLGMluydlq6kqrMddcaFinRwmHmoG
7oizjTXkY4N3UoysQA1Yv4fBllWiwblwBQPNw8VpcW8alR8QXp3MF8kJOaac
1wotACYbG79XfmJNHDwC5KNsxlrZRsVXJwr1zDTAlmgmf7iURFc3E2szTZC2
SQ6b0IXfRJKoRDFQqsj6/8wV1XFk/3aWz3GBXMUB7qy/kWLX6Lx7Myf3x6wr
xGWgqyirhvRg9b2BUqxXYElg0Angc4vhr6S34MgmqDVuqfmHn5EW6gpXNT3V
LOH8auHEtbrrDwLaqhOXok5gLcJsz3uOXUuNBaScWmsLpwt17PFk2JwvlBac
HdeEjaNf6vGhThqgCziSNBT/0DrSe7ZBpf7mP5zMxvys/T0vF/imlQsnBVwo
B5GRXY/rAB1X08/kTifTPZoCKqQklzmbvoVY036AnB8JCpTt1KzCpN2NR7eR
JkddYyzqWYDxs+/GiWYDaYVQgF/9sTDgY/SVnA/Nj+RPhJoShvjIz23ZsVyK
CqGWNmheJoknGpJKVMvfNnvXJ193Uq3qgLl+mpQOOLt0cwWiOTBjBb0itPEA
KbrtdrCclMdPCz7pguR//HtMYZClBjm+e7Z+0CvHCNbuZbOnScKCr5/uteIr
vypq4mjEpqsln2Y6y7oIfBmYc3vFWtJwPunCbnKgKSVMOnYO65Dg47lnckGf
fDIKHf9yXZsDWIVHepypPmfnWbvYxJBCMZH8xNPDuJyl4PffvjRw9EPByMtN
wPpGDg6g6XVatCZm+FO75a9aQg5rtRcVMkWRYgUI8UKA2xQbucpIzG5ozleI
lC1jyIVld6f7a9KYOlgOxMQ23FYEizQTafBM548CwxXMjiz0clfsV1vuqnYU
L3hNMm9vIXM2XFyTbKkhnDcMEce2gqnSMrUUW5TuT+yV9jHQNyh/H8pmJBmQ
jF51D/U7iuOROYmsV2t2y/F9oKIh4v60Sx2P50s51MheoxrV4tuvzHtLctKK
7/N4L6YBa+WEnEZ5Q4ushrTg1mh/a/krO7cpDzmmvPMIKMaCehgja/o6W5uR
wAAUHaL2mmZxw7IIUgohJWu73VlpzZk9ZGz+q4YZB3KYNsG4HRjUNETc2i2b
CVnvyzLS5z8Y7hNeZ57iA5XLwT+7VJnaCaSU2JnWeyRmoaD2viEKCFpl7zCH
zMuu7Cg3RvKCGV5GWB6RbVqnUpQrwYiGhuigpeyWf/pgGUEmtNvNCdFZrfF9
/7okilF/vnbJCjsk0xx20qibkMMtJy8XIhI6MuWAHVBHxSccmhsdgOy+u2Qt
S5zgWoXYFPX1/rZjzhmpkSVZx9Jz3WxdCTTZYYMZPPf51D70gwQ4bvW1PwRj
Uj+TbBKPoQIdnEvR571IcvAxC7XJR68dgGMNzxTPuio5Q3gNDlLnCGyL33V8
+OZ6qEborv8aKlBtcDr7d2tWoio7n9q1BikU0uhwBjJer+EaTNBdtgtnoHaf
ED7psYHx++qPDdrITdM2cb33/yfqrlbEB2524fqgChqqFUScOhUCdznqx0oJ
mSVgTLGhqxgVP1mK0WrR8a8YlBblXnT2j20mdhi0MEvyFVX+mO63wNwvXe0l
5rN4nDnkfMzrc4l7S3ZaP0VOSdDWufacnvqFOGeercs/UDsbs0aHyWmLStyu
uAue+2OtP62nNwj8goZngvX3R1j8oVCPfttbeFF57d1f1yac09cliOqwbpYT
CHO/V7dWjk0PVihNsRC4h5Zo2K4f+1i7B+n//wrDY8tf9m2fbZdpRBS+KnJm
yTrP1z6Ol1PGbE+JDt6PROEGzGCBfOeneQNiD4waYnfe0JVWfnfwzFaum3AW
udEfRp0eZPq6Dp53j6MoeCgD3yGlng/lh3CpCRuBnDjLtkv/jmsc0/Qjrwr+
tC/UsosWoGsjPc6a8EI8XvxnmczuVQFiqphz5yB3B5RRaaxTT5bQVjSDPCrt
XjLFm9KiIxq7RvqO3VmeMwMGZpBxmHZ+Nn44UZgM6VfT8vpbUDXYYpp8bzI8
+QnEiQiz1CJ7c0WDh0N2TgpswbB23CW89TOFroRxcU8J7+Rgqp9XBYeSNn6x
KQMdz1AI2DLtBPPBVyYhWK+t1QTmYyxpXrg2knDoDadkSexhcn4A/WzxyMqK
UjqJy+QdLaFeGwLhZJktwOLvA3PL5P+mvYEAXs6w7tyfu5xZ/QbZmRWL9v+f
fx1bmAbjlg/AB3bLerXUVGIhl8FoTqmrSt0dHYBef+ANXIzGJrKF/5eohcUQ
on87wM5gmgWPY33x0Jt9gWCRosIgQeMDoEOpwdIituXEG7PRsxEkJAXfLyFR
hiDLbK2euCIilUBIphmTc50U/puLuYGtDenRqMJND1+PKE3RaKY2BTX8v9Du
a619EMLWJKRYMfl8bLEGGoVUZLRMc5F8GBZfTQQ8ps0q8kHrNLvcZBvCs6Jb
FhwNY1d+ronOcUlsbo1JCjG33k/EfK72XiCyq7whzzOuGWdNykZN+m8H7Yn4
Rm5QvdLLWXXJOBcSPXqhYZuV4ufRszmyJ44IpbodlIYq4iB4RABiypmGadmv
uH/1EBTi0HeODnQMa7jjYguoHpRJEhl9YHfayg/cf4sQc79ArO3PjkLTpnvP
cFuHnho/LFDCqfBjngRYr/fBcT4oeoxSO16w7SDD9H2Faii42ad8nSgSymfY
3gbJtAOqs4M+T+Ji13uceed8fb9bbYknVHEssrh+lFJ65xlaZANAgDOfc2nG
DnruBPHCyUB7z2Kr9l/P7mI7wRz8/TP7TGciJlsavHESGsOO7qtcPiXbJQco
92kQ6W8frKx7WluqECbc+UdWzBTKBNP9T/oF3ehgu+ydK+LrzTLca9O7i39q
RDEWcdvMmf9RKJjfVnnNfuM6Rdj4m9AFaibyo2MFXY7Y27S2CrZ68ZZJbV0u
RlysV1S6FoOTVd157ZRtqFvC4Q/yc366jfdZ565WUL1p0WEmPIvFSSLeVqlI
F2JjxMJd/6jOWLJipyNUA8vvjKXUJE1gKEZn6jwA/QFe1YvdKu9eEPe9z+yU
zl9q0vC/gitOaw8vweds+ArOxFxUjswdwn+zqr9R3NtrWOs/i+jl9buBelqa
zp+DYXOwfNrKRSwmwOWoqenB332DEk0Xl43VwB+hjBCUo/Dsrhrm1a3JKJeO
3HiRM8Ebbe1JAKZSQg4qXlfDOGarmAkmwQQh7sF4euhm//2R2rCfQ303TSvm
MMfclsxPBSsEZDeFZtk1zACglnM3PDkn/+SLrqOC/MWc4TCfJjI1oipkErXD
qW4ZlfUoPmW7whGXC2KMK+hnmTFe/PU/yTkh0wkvHxfi4g0aWqNLvzwsijg7
HDlovQsc7qGYV5AmM2b3bnzankUiiCuj5vlV2DuZbHsLY6wVs8KJAYvfFJS3
UDNhPYJOk/7GkKOQb65p3vsYqm3gF+BFpWh7BaKXg6puJ8g3QoH8yNPhYB43
WHCQ27D8w6FyB/M17zzyjeHLL2DkoCLb5vqvqFz8Wol32hHyRqhc2rcVP8be
zMGesjsDuDX+2/LNjlkyiOokVzrS1u6EXei5KMqIe/oCB9JrAYGvkHBG+Re9
o0sO31QcMhyKpHHlBfdfKdeMzDUMdepFHdfZTKANAntm+yQaMJteZ3Bzmz6N
gX9+EDEn7n/J6P4mLKc+e6s4nHfN5Lh6KxdY5oLcscuXdsxc3x2hNqdicPgK
GrjFXfBlFgYVdZvEARmZmh8EeFwaP941bAd9r2sxiBwDUnJ+tNOAYhjeo/Bd
hAQ+9bQXVKcvIYZAKnXpy6xEqmEaUmuUV3MbB4R/a8JrJ33WvtDbC6sCfXVZ
fPI/KZJ1Ps9d4UFkzfmpPFuQltUhGd2JnStG6SZmsVQRmBsQ+ujiDmAH28rh
tmvSC6cyD7cWq8/634t2nhqOmzy2TREESGYsn0ES7BR6d+kN9lmx/QH8BgUO
4+UFd8NgfnHamAiUdVv6FNk+4brVvfANtLy8nnd1N4YWN13Y+JquikeEE4dj
LvBAZDyuP/XkhHnhkPaoZ8A7p00p/+ysd0BgH7uwOCRU9IYFgedd0pgRc+c1
4nF0Zi144d7gLSz/Vx5dy0ASyHZLgpMARPNmehqJZM+MbgFMzD3OliXgIIF5
W6l8Hah7WMXtAVbpwv/vvmtJp4lDFP9fopaIb/IFgttrrxdAwErSiephZlq3
593xztdSENCo41aoU4DDh7/u56gpWCClRqiqhDFoBXo0Q00+fOlpEG4aZCPg
sQWfJrOB6GYp7HVQjIv743gawI1lF829514OocF0VRtt+o/DtA2pfvT2XUUs
D66hw9lkEdOphy8yotJoh+WkzVrHyhdadC/TugqYWImbT3CBe8FW79OKHOEy
81FxzOjcGZjKrm1jFty19v48dy+vx8O5s6VK6FmbFOoncmdi3p6a1GMnhiQe
IKIpefgNIHIlXceqAnbm1j2zD9bFW5Fw6n57/2BNLEHPZPpu71epvhR9EWT6
vmFcIlyxj624zvakjNFetgq8prJxDoPKD821H9adrZ8catsrBgWjEwpkkPMU
UGjWchd9A1RO8BC5eWxx/PTBQaudIzka9CEb9gfpIEPn4Duom/Fp07KfsfOF
K01+ah9oQU2QUWpwUeR5/X+0IupSJNY5LQprUEtzzhhUs9JjJK8yiqtx85WZ
utKjZSkTqWgqkirmDNTEQH5nqXmCUlslFuexCEzyaXPeiaN9Iq0JUqJ+AGn1
Xwo2n/Ddi3rmJKsAgtUECgymxJFcQexydrKGAoweKJRGRHnn2NnnQB0USXy4
S0mqbDALmiyWgDgRgzLMwycnrF+5oKZIcNz7l5ZCtrrPQkbyHer5eFAb/W7r
aOYNPeknVhKBDmLJcT/veNRcn728u9Rf5y00LcdY7KJ1dLHqeAidLk8ZsnPH
VLc9NwDs5p52KeeMkFZcDLb0Jb6rwzS9//YgGOH1VVg1NJ0iKLoanOasIyOl
WGmVR1DsSlPdKGrJBbxEUbkFsRqGIBAvH3/QQIY5V+4fkfpBu2zVeeTA9J35
QtFVIWz+lHJ7d9mY+2xfNI7ri9UHeglbYHd13jhaPk/+ZKCfQ0VsjyWkY/uX
pgWovDhsIfs4oSNNJpMd76gT381+4NTTAiQGUiOfnWiGzSrEkMgneD8kNBjI
HYconN6Ph9b2Fxp4fy9TfxcWv1AEOu4pA+R3bHIgK7Wk0hdUgxlJNQiX0Ppt
dRyQ0JjktupyA6UTvJZz6/vnl+wZLTdKOT7N7yUcGDfTrd8PUKSSkNNcQTfc
1FjrXX7nWColCY3LgVZ29UNVPcN4fvX6cW6YRO3jhaLAc+FKNZrtgSF2NcA1
BCMG1hw3h+yekDln8hwB4VV4d7vrg5W5LNbJbCD6fobMTAPkZ0WnmZtGgu+p
mYKyoifDLtPeFgilw36vWuR4Wu4ZVrlKrQuAsOzWdkqPYUiF2FUOyiFSxymG
TEA8Iihr/hh4SDZplQpkvSODn0P2B56HdCsQIOtardp8RWydP0y3pu76v7Mo
AY6+uurJRFGiikPBFB2YDbDZ8dwj+wM36nfsdjJ6c7LKQlQL1QgtaglU9bA6
AIu+LaKXvfDbcjKdyGDpqBfn2glZkk/Hzk1Ph0uFyd0VqSpIu0LQ02U+K0SQ
jXccnTTBMPKh8hDALmiF8TUPUt9xh/WVqQqDGcf7oj2joLBT8QbRFN4jqoFG
dmuCzm3i8GYhmYJmZyECNjz7NdlNTI+2PrBGieE5xcoyo4r8gLrcUx3+NWLY
AG4xHbvUsDy+1jrYWl/Ga5/rggLlVV0nPjHqkUORYDZ38zbQU4LAiWAZZqsR
au+7iTQr5w5/2jzMCJVOqgLEu+Vc+x2RiatwnVkuvE76zQRj1twca8tLhCbt
+N9ujC1IpvRthSGivYcyVpq4MDpFk0UxySYCAybpHPYE5o7LYdj3g5w+bziX
Iuukmu+nI39pEgs1Wen433rgN5rDyKkMpehjW6lsHBNzQRSXJTfXVPsojGuL
9S+fuDiKVuP361n1lxt5mj1ShIN6FdUw13D/ywPA4QcL3xsDie+j4yvLXqFX
NUpVfKhpbIv20OsCXMDqWaVZgXjtdqtpewPVPQzf7pwRtrw6v2HaIbL9RX3s
f7T94ZgD2nl1mj2bjmtY7QfGuIwjVe5nV+SIJ+5gfJmH8mOSEUbYTZ1JZEs7
Bz5Rck7kOpfXjbzLcUG5wwyXxLjtapr0oc5tD40BaGakUUTV3SN4q/thB/Cf
RDSv6nPv7lXxt+JqutIu3aY4bRROjvwVLELJEBA3QFE94shulOIK7Gczfzas
t6kPiPlHCmBUtxH62nADJz+lgDfccDVygCFT0hXVohjC5A+OOLWdhDb+bRF1
WYQlyOhoLUXs9BKRQGas26aUmhaDUt6bZZ4e/iKHevOYQ9nx/hAl/3A6iS+M
TB1LJ7y276VFnlc0yU7OW0fYzy6GSDcfAouBcB/q/3J4Mbt112TQCmpY2FSS
iLBQ2w3h2vedn949l3Lp52WfqavbGexL//Qx1um86Jnupuaj+30iABvKcXOX
IjLNFn52B9byvh1sbaSD5HEpjhXeJUbZH4UFbkiOvhfGxBhydhIAXNqutClW
pfCyuDbeWLi+diCKCiX1uqXndWaLzq3sz7gFv+/YPkJm87vOpx+mkE5tA+Hi
vO1kT2ZrWVF3qpMt4w5nAjfeAA6PMH1/zW/zkJ4zXne8bsluK/y1kxYmk1X/
ESIO877FLU4tQFI3a1AlW6VAV6W+4dtZnRqMuGgat+HFbVra/un+l9xbj5/U
KD56u493qQzwWgmqWesHOKYrCy6BWjPUeyp9Re3rhUSQt3qPkZaGZdLyia6I
B3xYLZRVodQJ4PiuLMj8aqJphCuXGclkOwwVWphukn4DA54koWCYh5RI/wQ8
BKC5jICeBwJSNny/Wy9FnuFdvU94OTTGbfiuNvYl/nlPcnfrTp7eAEVvewEh
cHpTPBwcgkwsKA0PD6fRMhy44HOtMnaLY3gnGR0Mx4vOFXoBZTcEwGDxpEwR
6jReAmFMX7UslqJUz++mEjKjkvlKrnRbRBSl0KGJwG+tdCzVC/Gc2LYi1x/b
0eq39gcpfUqXcmWrzJvTt7GjlUj0gKHXMMyFpg7mo/c7yUY2tisH1tXLfarV
1WX4+G5zoqLb3TklXedivkiBVp7NiafntMLbxMeyp78exE8kM4wNcHqGO0/R
6UNa3u0PSjK3nJirLwGbBz7zhwg2Ttw84OINNim4zH8yW4sEcXssFSFffmvh
EFZTviku0GuBBWcRhL+aPxI4/N8/hqkfee5AFxkSszbm5IzMO8bINEE161Lz
JspFwsUjvsWZI0UZqz9D+CIv5/Pv1+TA5uQ2CJXNM/LsfRMXLoerTUU+fivM
jOYWAcGpTCjZUor7g+GdZs9YHVPUFUlUveOg9r876q5pBpFRD4DMSDht7zR9
abHfdRtvyTPs+o22vKNvuzAmM5ZLKHkgAhUV6oZqL7Q4IboOD4rlUsDcqwss
lQ7ce1mPAdHkib3TnwB5gwU/xzwG9Pc7FF3w2bF0tHj76yByGD7inUxZnwxC
oVt3ieASEzbNTSStnxBlv59GtCzec6hT7LbTIZF1GmbrWbK7lUveYlgEkumX
ZIUl0zuJJu5ou1/mlBWnQPO28Sdq1vegqnECA+dDQvlNM/AjFqvOKGMwVjqz
zQqa0pd+r1MFUHt/tI8H7ZgwIT2AyCJdO8XITdmcA951F6zINSJdTLqt+vCn
m6kQHqJ41AAVfvPHfQ8Cb2fC3jG5WZCPNd0dyAXl+afVZys3m1UgzU5vK0wv
PU5Mkv5uXvPYCzKOdLeBWZCMl/ugd+Q1PgXK/GdP9nz2D84eF6XFMfWHpNYz
nmHP63BsZb6p4hoSK1Ji+iWULTqSscxe7DHo/5WqvnZTToKxp/c/U8rYJXfn
toAwjPCLUreZV9P33o58SyI7LH/NR4AF7WoftBNkdLh4qfs4G4RdvfBROVGF
NXrfsbU+TNZyYzofJiFALIwcyy3aDF6fpKadalz+X95cfH7SO0puFf2j+sW8
xTfKKMi4WUwBrrMyrlINZRp3VCSDE0yzBfny0HVv8K5MLumvA2mLDLQBaIU6
rdd4fcuMxkUs8xxOUTbUqVwfinl97aCDecYOIzj36+jI+hMxvoEKqQqyTult
QHlI5xEGztjqGnkAiLl0NQT+9F5F9Bta3QannwJGBF6lgw7Gsx5cJU90f6J/
53xCc/uAc9NRoQP2v2UHtfuDnrtJaFbArcyzYPN7EQNqZA+iJtUDg5HlcreF
YEEszBMdDrsBH4p4TG7P5GIuTZG9N4FtNpKrlCQ9Weqmcu8bAOrSf0QugpLk
Xe3uF3fDutvVZJAmcff6BAWkytQd2KQ31jmodmqwIEFgun/uBBJ+0GGr8rFV
ocME1WDFhmKPpIbTvT8TAVH9aIEEeDKOzkVVTI8jSuqB9l5FItXI3XVXLmxW
86dv/UyMtcGoyf8EOC5MIKL1DpQzcEIz9LcVWY9LLESuWgv7DPPCUdS+c2l4
FYbXoWak6a827rgxlCOydmML1mD4xeyiAfxJ1TXpkxw9lnxt1+RIARdx7X8u
7ktW1Fa+LUWLeszUp65/ArxBmY4SrFMzadJCUqHx6SE2ezA+YVIqZeS8b8yT
i6USoYmA2EboOXnGbBdBoNYi+qjk1mX53YgklRBxutH3K27PVNR+uHangp9F
Y674O+i6FjnvRqsxP2I5Wog/it3EnMa73IUAaXZCJEq1kLUWcQ3FPCxMsi+i
9B3PKDB77PCkOtyxOVL+CKVcpMLJgkJTqukHplPMY9CFFiI52WW3tGKgqz8+
+0cKgTiYLhvUFTWVEwzkJw8mu+I/FLo7n6Tp7bat7lsA/fv241731DWbliTq
7DYqukiiEsHLWaL4lP2pblC9yzxq7pmqroIpn7tTRG1tUyhvnV7Sb13r6jnt
C+dI4GAlSMbkbZedXW1Qw3I4pnI23NTHJ0kM3Wfo8W61buy7l6E6ZgWoz43W
uAGBG7kQp1QT2Aot/Gj7Ah+YtfoXS83LIAZIQJef3vqocZrPrO/pW03ADtam
lSjbMC0aj8RKPAh5zrkiiXWYbAzsdv6SMuFDYedKhZrkNgCbCxayR3OjgTht
op2q4bu7IEMnGJDhQlCSr2FlIGubuLyxdJn5BGD+TBlwhjss0NFxqOcbABz7
bUCRyqP779mfo4+K9lsZB4r+RNPG0uSyBvU08F2cMtn17IZHjAV4m1niZz/h
dec5nP57bt0EtbXTgFcO+RMIe5kf3SXUV21BdS8Tfol17Kf+pRD+7xEOnX8c
l+F/6Xh5VdYwvvYCKaE/bENt789HSlgdJHlGzvlg5UmAgYyB+utWViq/nP0D
Dr1UUdgPdaExlceMhNVqh+4Sz49XShge5nVCkJaAzV8Za+X7wfTcHBPUCUsP
zbjfiXj+FtoLSjlqmkWWZ5K1Hu2BiAe/y+4xwPxFJw2JEI8LhWl5/w/0jhYN
PxbmZZJvH+4IgtPxf8Fz9ARB5ZDSwYJxFYzGcCfMKatXLyURR7NdXip/Obrp
uRNEZLjyqCgvjNmNVpaaqrb64p7tTw3AZU9zkSzpoEFTVMbr5WDqlgVAb/ON
FMss4TpT7DIzQ7oBmZ5bkclPsXcLZ2+uo/X/8AB75FxoVhH44g6ayRBUlt1+
H4TaW/nYA4ePE4MphiLnRKfHByxu0599oU8rHugIm7CRFiYKO0/YyLBJRbal
nbKKmxB/i0Vh7jd+akriQ1igkRRWeoHOKjvPdVuIrqhD1ceZqJgl+mPlyTVS
fBvQTWr+U9pwNQttX77xjc6/3r4AZSA5Y/XB0rYq15J1FneQKAs6KJxcnL4n
/1oADqBohSSFkTGnsnhzR6A62Nyv7erVaY054Tg+wSAPjo9G1+eRlaYvV1Kj
76YzVq/uypRbD8FeAwlb+d3hW+7ZZjpkZ9Al0ysZpBzH4yBtJarVD7a6vh1/
/HnJv4jNI1FqJO9UIMis/zrg1fAGbw29D7X0k3vLWVaYTWNgPPhwaXP54FUi
j/hIPHve+6ws9SDEjFEBBEDgBGgDnBSLnVAIXlHXv0SN4dI/HaIR4bKaDBl0
69bZdW4H9WFBjY66gVQb1WpxrXzuJLcTLe0RuD2ECaIOpS9XM8BAWdaOtoFE
GjiYJl5vxeTi+YOOWn+f/IfJZwB1ZdWmqaH2zctUmnC1Wj/Rk0ZB68aP6sK8
GVzdHjOXuItrFs1QG/1v0uUgF8QwfGOFiEvYUbXmumDzsJKIu86n2rNYnCDd
WEZo9uWg8RbbSgbaC7BCSLHNiWSRD/TcNKjRYx90YqQUmzVtH9FWq4n9NItw
YVJ2kCXtWrgCIZ3f93NgqoYfksCb8Ht509zDJ5MA6CPF7vFVv7A1Qh6sdi5i
ZWnKZKTozPRQWf4e6lOa01JJqNfuYkXAA5qtMCpLRn3UgIOFXnahYaa1Qxuf
+9Xbz2GQD+MyoWiDRdTGt9UBpOR2r2LF/IAHcmhTZaru5I1yxd5muq0jP+Bm
z4LyktBId5GscTYpx7Ye7s1wMWLs+RAfvz/VUIOYJFu4xeH6vLBxJTa77c+1
kQ4tLTxxEAbYOepsHvvCoxlOGkqQylEoCWbHfnrMkLFmhSbiHswg88eP39j4
u8u6NsSXlmwxLxs92jLnXJUwtW3d4DLNRxPNdryoaYxrhYSa2UhgtPBjKfOe
MzZvxqLB3HxO7CBveEeeqede0tUUohiQlmlJmSkBbiyWE3XCwS0w1wh7tv/J
zDw5QFKWJCOJR6c3pQuHnq91sd6qsG6+eubHRAHPE6r8gWHPGjxg1iYeJl/j
y5DpbKUmEd5cqtpOuC7GhDzJ+sMB162P0K+vTWH8lKpBpILp36yInFDOksKM
AQYTjI5Skf6mx0J0To1fdezqNrkObpeSS3+lgds4Vq8YrEDdBgV2MfjWZxYR
F6u9KFMUpVFoYNj8/NreaD/XGSVg6fZ6NMHIis0+O6LrdLHSK7lSUEQnGGsj
aHS6kh2z5qZ0/cBEa56SzXN92WPRMdvaPfRo7tXAmNmSxVcth73PIClROT2V
85tqaMvrUlWQvR9wOArbG3N7Q7TbffSwMm4vB8DGNL5NbAaS0+ju5ODvEWGs
fTiH+5zS66Aum2ZipZ7OkxBBd0vTdlRMeVqK5XjSxceVQZOsj/g7EmY03hCG
gMHE6TgHZErcS6SnWmAJgvqgfgrwQu1jnfI0evP3RsTNp3hX833eBQMSlbi/
DhMpIHsR8ZxAHM3arT9rLbjrOhEPELph8Boos8FldOIsdUaMfdYZ++CYFieA
IwhQf5JZ+KywMPxB4vKWpKH3Fr3Qgkvd6Q5NT4tuFkVYEWX96wJpUpHnf5Wb
e6e1e7Cty8NUAj/AYnXVK0MowuKM+7nint/wZDLg59ozyUBqwv8ExEeZhn4M
FEMLzd7GYN+ZFRVuWYEI7LiXFkLjAKNcsBEZdmyL1d0xRV6LFIB7e0t4MsUv
nmERfqnKyKrZZ9+jkXrj8Xnqw5fgpPf5iwTR2N1QszBodBsqPnGDLnqjFGIi
u5/l+eMBChgZ+097A1OqSPc3jxgNUiglgSbohX9GMAHCCoJ2sAaQvkm8tt3W
77MMJtuH8lTZp//WtiOcIBZ1JrohsUZnBJBv+wuqek9GUQDrqxb7HBwmgkMB
jTnz6I9Yld0L/cP7hv6KgQLyHc6wvC0J6DP/Rwk8vgxywDGz7AUATkVV6QFQ
2pGPjb+tTixCCd7W4z6gVm0BPUBDepnx9wuuTGuwgC3raWuvaSqNi09VbV1v
Kv51DlX6AFNYRuiHrl4bs8EyMyBAezoq0/GmEnOipabHt3gIRyMLl1mzjmoi
QdXrW/Bt75uFLdhlsnXnad/kzB2U3zsctbbW1rJ4sn/cJpmWOQdd2WzGjQrs
DS7fe8KiBA7HwJI9J9rm48L6I8cDH8l9LTdIoxGdIMaVeE8nZqCpHSvHjf+d
v6RiBMTDIFgkrCygW5DbkEqCMUwEk12tWD/9CM4Eb5rOYl+59hUiqlLpQdOC
svg/7wBTE9XswmbCwGQ3kC+1qld/93RRBUgSco2cehWZfxYQ9yqyJHbAjNno
xAyAsd0OBSgVi1ccG5JlnwNLemcH0SgwUyoLfEyGMgrYjXgLUlL1IKx6I9yH
6TvGE8vVgPed5K7VyZJ7hn0bPBV7c6f+l2Na03DuD3RTWJWLefUWX5Qkuf//
KOoNr9UQ0ZG3zfsECD+YfxkwgZINzxehtjaXPFYdWbXP2kfo6eoXQsHpEXWH
iUWlNrvBazUM4bQ2WQ8Q7mQGYdu7urUCgLYJAZMRf6YLBeMiKMlYZXwKPCaZ
xdCs8gg/NqFuHrlUnD0OwHJzLLjSeoArvNVdzWtxnea6uzHa9sTXmfjyiWgK
dl8uu2USRt51EOgSJDz+SkhFKp5pDffWK5DsPSWvtjOnOTHrbr+z55f45iGp
emCxnKftzbdMd/e+uj5QT7XxBixlh5AqKieLEFkfSFx+xjBEMV2rIt6JzkVZ
ky6khL7rp72zV23FigsTWcERxZ7ktmUXZRbh4CQQYnUGLvFyZYPKibmtvYCO
zd2Dj9+jSBFdWTxwwoidB5aXZC3Qu7SOMTr9skxeLHjpE9knrO0hQVjpL2WE
6afAWkXamAo/RdBsNHqi0mxaXkNTisUTs0QJN878gkoh4HVsO2Z+OvQN5Psl
5/X8uwk9kvwQSvk12yNpivcu6CkzjtpibhhpIdj9gtzzin4+ELN6oy2fRh0g
Z/vUP9mD0zO1G4NWQ5A6PAcW473ESCZPn+HtIWXsWLy3fcOaFE02Hk0JKjk8
e9bjGteRW3k+DOrwnDFHRapQPbH+rf/z+DRfrV9tnoGcOjCqNTOMbyd4VVW/
UbHs/CVZgnkYRmgMDjpm+/CJRaYjrUkjoWUKANpn+HCJjl44ddPuAvNuTEDr
5o4zS4vk0dc1NAAmuKZ4WEAsZaehNMp3tP7h57vqFDZWB1wryod0yk3oqGDC
w4Nm/fTmgCYkzcQy9SMK+2My3sA5pCXChY5qPYXz5pQb/9FkuRifFHmm6ccK
OsWUfMVgvMikJlGB/STlhjhFhBEZfjGjvsIsr2aA43flhaP0Ylu3oMIgDu8h
F2nViLwLphUqvKn6IWedgBLqbzqqYUGynbLLBNejwbu3ofb+AtvzGejEOXyb
74udq9K6iY2OzPN5chuSoyC28dWfGNRb2ZNYoUW0r1D+vQB2vHgFHD/QZ3cg
gh1pMdvxfTYS8siPZOAveRggEH7WZEv5zW48cCISI6xnit3nehCNCGgA6Qh1
W0drrK5FgASbApYRBJQAHsCBizHJPOVVySj5RrVDPOYMaqi/LNjchLmCg6kR
Sh0HdYyZESKwhxuHEboJXJRiWhNd54f2o5bKZALmWxx7kGh6xSZ6PrnSGTf7
rYzfCgHR5jym4fGhO6PjH4hikuOn2qXos1ctoXcyX1rmydL5q7rESKZlr/oB
70B+S+LMsWzZFTLJiVNrB9V8DHZgSW13pTU3+UnbD5skW0s563sOifh2wG5W
njN44Jkfa/aClS91bn6jtSQmlwZGQQDyDUhbQ3hWVs2WgunFXpPvhfYFl32F
fXWDSTty+GJwgRMyJ/StLvVtE6ILXxe+PDygXfVL3otS2kJ8yhf5bwQdjixt
vpB3cF1/RWa7jdLnupJHug/eU8wDVDfZBi0M78oQnokAVBkfxe52+A9UKG+G
kZCRbQavLiBtPG+kVmq33roG7Uk2F5gdE3wVAUhwpe56FbSfuqPCjwWEfRqX
bz53hF5cAv77bf4z+xauqgNb86g1UDbbhfrTr2Pcx/8/ywpz6fjnA6h9ucdj
x+EnGI+tAwjg/9cNPMX+3pd1b+qpjMPw+0BGHFmTKziHTZoe8pXanP2qD40B
4xGtDl3kDmKATGWmUzxJetLi8PUsPEvG58NbMVrBhX84Zdk/czPKbWdOoItC
NTqRsD8Y6Ecq7gpbf2wYvSq1EBSnCCcuTFsLHgg+nqp2MPW/9REZMXZD3cdX
X+EpHDWtVWdfGwE1fdu7l5ssGQ3kxgfNGUJOum6Gg6EJvTNrx30kxMqAztXk
GVsod3P4g4Ub/o17IGjnA1e3gTWB8D5tzwIbU66elQSPdiGPRyskfQ6rjq/a
zCc2M5eKYTvfidwqCclUC+QSGnEg6xjlo5/3vpYd9lM9nDm0pqiixkHgLUUe
xHEz2JL3ElYAgkHD5plgDedUlt0/9ZP/KDmGMedYwZL/1pAOTY5Ns0+CqHjf
6kpb3izK1q4a0rjmHeUr0AHnRbQ0dWyaE8SjvDGPqv8dIYj7aDaVcBkqg4GS
OSg/krMr3URc49NJN3sgNALKUtOI87UL2e31UhbS+8jA/19RVs2N/8yVzb+9
U6xdcX1Lre12BBE4jtTPmbOYaLcWZMuz/UCUXRoCHxEF2PTTENSHolrwlq8f
nsc0ieVyvcuFF+9yATJYN4ia3n3NuH6xso3+PRREJWYqws3RncDbDsTO7VGB
V3scYxpZVohbDcco4Td5wmkmFtSh3Qb0M9nmH7SpKjjCEDV7shlJZMvbjK6b
knFf1aV2R6qj8Di2vTjau7JgFs2+nUMpFr0cPg6LrOMgW3FSCBbmSzbNovQE
ILEBQkaPkIKFol4FJ0qbAoek3a6RHlnBstpFX691TBnHn38h3XfJuKWGcgTP
1FXca0/Qpvr0eDlLO3dLA2p36aS4irmrJoicjwzJPifORgY9EXsrqIgVz22f
wKs3P+8Ajt6iIZNTKmeXg8T9qnGyztVQgfkYY7Y4qtYQeuYXeboAk/yKvYFH
9bJvTJWPQnuyhK27pvtqJZm95yhtauTd4/IF9TUGWksIN9nX4blR3JJG9PaH
HQXyg/SGLQ4OPeQbHCfLNlijAzHT/nPoJ/puvEbsUzG7rpuwrsH6Z78G3ML7
RWstVjWW+EJ3UJYmR4M6QW8M/EeSpPutzkTPe1KCjL4Dzs5aakVWQ8vOOuzU
b7aZGjsz34iQAqsPYSSzizPrCCr87i82NApKVgNZJVRvw3QvrmWxVwAU9yZ3
hYAYsOEw8TjmoIjRXFRoMb8JR6JB7C3xyiPih9YbxJ5oFZ1L3f23cuex9ugk
L/Mw+KJdEEGCAmtRDEa4eb9S5G0QJLWSxbGt/einV0bMcOSfYFb82RrIsHXS
KZ4htfHMveY8QsveZVJrZkuM81n3zmQGdXH7EmWMn4/hmBk5tfAcnbvrpa1h
XKz6fMfDOE0PqxN62Zc2FlwbK2R+JGd+5IQNt/07fxA6gfXRSF2YfdNZVk5z
qhibV1uD6//XrZCcNF0ABvgK2e0j8oHzV02EYCT8cyoY7ZnlRLdxvrRHt3kZ
OIdEKWG4QMbXtR5E9m++tw9MIh+uh8xIHI6QkQUVBZlePEttYT1jdtIip+o4
qiA1hWFW2KZk3WE2W87FW9+aILn8rx4X90ZcskpRZcDgmc5aclDUDPZbbEn8
1IoOiWbMexIMKRuCkLL6KWvrkl+wt92zmkjJFnpZ89xwTVDIMsUsyi32OG6g
yACDYNY0BZvtgwFCKdq7M4QkQdtWXSo0UFRLnIdPqY3cIJQ4budenTeJH+3C
gUt3s7MfX+PPof0rdbVcHq9WyuDyDVkSvL7c9s2ho56M6TlNG8cyrHt6NmI2
ThhflEe1K9LEm/fKJOxSczJg6cHvku1/uk2yukN/dl7b1xnM4MeIc0NQM9Xk
ziwLvWVYeCgv3ruYMyNcMLAvMNbeMa6I33KvlWDPk20kdAf6ECHKNdPaGa3p
sCNjSMQkhD+tfwQY6/QddIF2dPrb+28ud6l7TaP438ZCtC9CmyIA+Ng07OwM
OqRRXobyrTWnf2nDoyXjkVunBcCn8AV/8UzCjBwNnYqffMvNbfR4P9R7bKC2
DkZZ55ukwmoI+1SLE+65jvRYD5TaYY4x74OWhUZ78z//3rykS6DL+T5UcoQ7
K/fzOI74SbmU4EohxFkwqgF6ZMS/UlCAYtDLdVQfkRXlfsKpU9j3NiTe6RDj
VDzrsLJJrB08rspsR5IxvtMmtWUVLnpan7S6ePBZIDc2eoDt2/Gdxjp6BE+A
Ei1dBCBwQE8sGrrEANWw+Q7eE6vklap0eJ5SwVBwaIqHpVAM8b64+ESqycCP
aenwh9CKZ12+IH3ln8WhIIbxX9slGu5idG6TYcBb4oaN7jlA3aJbPAoIgGSK
Xkq9bnDNehhPq3lhNMoYoTQbzs7ItqDUcmeb8W2RHt7n4cOgpFjehXHZ6HzZ
/ckUwBOSqbCAqZhZH87YG+gZZCoJGJJyIIZEU9XqRXGwx8m99Xiy9ippFt1P
tiYAK4MP3bJrD1lj+mDK2tvF6Gb1Sx9GFt5kXvDi8F0WdN4XGF6nwyCi/N4W
2cyIeImdn5eeN/l863odhiuAbcu2NB6vH0z8X1iqvR8CMDJSdNW4hEaQDqIx
rYZsSIIwpLwg0qzoI97LnCu6NaYEugnNOb3DGwUwHJMHZmV8TclMbUkmCdJ5
fKnDS/adtmu+9smtAEOUhYzVQ0b5Ty8RBgSkBv4RvUvTMeKZUUEISTaLFl5o
naGVU9RFvUCyE96U0YgKI4LHE0Zs8dr7PLMf5PjS8Tktudbf7Tn7+ND8JgA0
qC7z39beWdhEyQwPhf01Xe0m2NnUnO4Z48P6o3Z+nEJWMJ2pIFQTjuwj3Q2X
kCf8635X4ur99Wxsp2Zh7kMr8qLeBFirXuzhKEjzVoj2f0urMKyexdRyR+iH
FyZrV0vj3/iQ55snAdimgzG53/iaIRNszeHqgysOJ6Sy1m0m608oRJraiigm
uGySi8V1jh1rdIz/EW0Mf8UYXnhwzc4N5fokhrEBaasA/M2GpiFXqZExw6DL
woEu78PDVZDAK7y9S1fF/oF3j85zh381HbbslJz4nY75GVH8UnuH9inhOAs4
Ia998eYGG+a9JgA+RtL6qmr0ZA9eFuYciz+zlFUBbrjyocv1W8Plwmfb1vYt
J3XmuP0+2uw4cSXnladAODLqBvMkbmEZ09rhe2si8w0fytSMfaNWduHm67E3
XWH93JJWI8feBiJ5VnV0p37y/TH2T80RpsT3RTeZnSWkDjINlq6nt0pOQWJZ
5ahN7Q8vYR8n9MvGnZI0ZWAOGpgCRgGaO2xpgsTKBoU+oBy5ZMiTGSdh5Pd5
Xvdmitv+ArhC8XWJLtfQ7MNTVahsbwYJoI1db4iu/sPrJr0yFghzWFyCuPri
O9/wMuySyES4atJLuyhAOGz36UGptcL0eglDBDwNaV5hhOXfux3IYDCt9aMa
4zfkmmRHWToF2zzbGZYSGh7yTqzmLRdin/3AaQvsW+xeaFXBKVHFemTm/THr
MA7PD98TZabF/zAPk2apLbempSIiZH+akrXiT8kxkTWacboiArvY/yxyTNUN
q+eUZ0PF/Vx/PBVPunIHlQAiCWmmrCKXERNo3iqmbU0sbOnUjKosa9PKFH2R
eiYk/rg7EAb3VaZnV4VYJKw5HQR1+DwAIEtEbQniwzqaz3RsVSWRsBXlmEkk
taR/770Sjxgq2whwFC5GsqfhYZLCftoMnMTWqjpJV8AmYw1QC11VGzKXmlRL
fyDZn5i2vUbzq3q4KKpfLvDPT1PJ3dwSAUC3+5RtCg+9zDcw5mYCQd2bhfny
leTfaha+Dd7IOXu0QVVbAzbNJJhV+AlVUmDM1Th51fzKiF2LaRpXrMkX0Ct6
Wh1vR7SKgrjAdrFvRiT5xYgoJ1dTMsk3rSIsFSafCttUjRTQG6UI0XL3Jt7n
dW/CdgY0rk0shkAnZncLP0K6evCwHrhL0J6xlEWm4M6y6JsQ8AQ3REZ0RvB7
7ZXA2La3uuvrets+OHgKJd0WM3T3Jp1wswQ1a68qggAsAcuy8RODgTeaf4aU
lbs90mB6H6j/pKNis+OpJTn80fDPkcigUoG/HIAcgPz1Fjh/IBK/EhOqoAA/
eItl5JvsYfFZfmmgJoXlrcelIjJyo9FbaZJIgaA3/O0lD2X7GukoU5LeAIbM
7IC7Kmdxy4+IuSRCvYrD+fDAUtP0vrmMxL6cTYeXPD3fGe+A6HaBngBYD7Zy
+hmnCcyb2RC4Ar+XxuOur01l2ToeCtV34WeV0qtXm3g/mXrrtF1dCSl97o7O
h9pDrq/ZpB/e0czqxdEEoxoPSS6Q8/2YhrNqHWfOOG9SOoB+GCkEslqt/y80
kkQafUFbSk4TIbmhz6a3lICmcOpeOY6SD8QFd1ZJ3xABog2zU2igavNbmbBZ
2oxL2qdvhbeRxuEA1siMWDl89clzCsSAson5LKoDT7FgTecq8W2CHBq7Gdh8
/UhFR5ZCduStNrAbjw2R/tHwYm/uVh9ZX5nt8y4U5MlNJTCVg4x2ncYBxsF+
Bkk7cZenGNW228hRXkjiqKzBZxXvNwY28Ocly7/PC83GQ1CuutUtikB2IPrs
p8Tob5YvvYuZLGUdTWNgyYZts4Uw5X6Oh65qA0wouuyQ/yrQm+8TD79t9Nhr
F1s76V4u9jgFgJgRqeyTluaRlqjv6Ouubc3AjF2+v4XjBXEGg7e+qgcNFM0U
a5x3bCl8H6tUyOCQ1/UFiYuWBf0sX13UF4SrHtBAXsgfTTKxKYPTI+Isqdjj
xAYwezY3zdbhvarLtDhv1R8bTWPuB7Q4WCm1WDODqipbSstOmafoXxSwD3u0
cDrFnR5JbBQfamSeP+Rk2lruktqP/LBAIpGjYGiwn/BmhV9Gi7u1B+b+J6+O
nS7Oit+3Qg84fJrEtHV1juccgzoBU8Za9OOmqNpFgPQ1qiL4VDF3P9N38zlp
LgqjVAqyjMi/ijaame/7PRfG49e3fCFKR164hj3/aR8e2yxxt82xQ/IyWqpT
ThA9Sni39N03qWG+/tU8QfGaQllD54yjZPqaRenU/eWIgKMA+wf8ujU1qe6j
iYFC0o/VKNpOmaB+Lod/QfwoIVv7hmAsOHnMw7dHy147ud5lNRXuccmw6YQw
YccCJmf0CEmu1AVT2hlHZJnBd6DYFYE99tgkhaN99zON2EPMC7u3CMc45wVx
tfLgSfq8uOKqzGbhj62V1ubgG1digWUKrlWlL3/tSuRZPer/1DxWc/qXJ07S
DT30qydwDMz2n5g/3Grn5MUJHXvunyhJyi+9UeEzdrOifD/VyoGBy4gypqL2
fAE6n/27/ujCjhTgivfykBcs+ZBgfFOMYisjfOlBbgbHICBSFGvhx/Qze8jW
PzUeFhqw5knGKVmTpuG7MaNs4NhQucU4LrpnN71woYlEYzrFuCXKrW8arTnV
jshNSG5iwwLzg5qG29AYxjFefDXCOZmWwIOz+mTwswgD14mKYUZu6mkm6S+B
/M0lzPvyqcHGz32ZEwzgDAWkRs/fJU4OZC9JOzPa0WhtIiTDEnrF1/nqGBOA
uaDfQcnkFriuB636FPTdeJIiIzM5w2RlWiCeIqjZnXG77WijpOhHdTyfQ/N8
WRV+54SFUkylBizTvazjkcUC5ShWVwCyAGq3eo+j39D8vgE5pYRgALppOpm+
i4W51kPFm27RRmwiPdw9EbuOp62mClO4gATdVhzJefKc+/fPAKuMw08LZdNO
QEIDlHNB2JuJJ5OPFl5hNvnYbAMYg+AhbWl1q9zXVQN1e41WrwmW4JHI5nl7
zzOeKBT9ltFgiENOU+TksMyq9bAnT1fTG9unDsFNAt1QIeOvJju65ycdsAfd
qSY0DQ9NRYRaqvf8kK7TeMfXcm3zq4nZ/HxI1HVmcv29LcBWvqiLca8kyF9x
PN5CXgmRc/gsdFaZkFb6XgSTEEmYqtxtf+nE4541PdAm9nqzYdYhonCk5TvE
hl1ygm6oqCIGEkdIPPRRUifUvcalJrVps/Qt+RNSPAaPnm8JNs54GfWD3ZP5
pvUMjg7yXBrddT3qSFkBPUfSLxTMNSpMIrXfNiZzoWv4SrFyeIuqU0Ik6INH
DRbpkg11j4lvwHe0Jl63HgSffrBojKeYyppnvcTcoqkVahvlskRCHbui9SYU
hfxwUp1olDNY64+yklIeFCkQzp4gdV9cZgGs/y6VFSWNVhFU2sQYX+xNGD17
eczKGYtjcZJTa5JhENPDaxB7QvABs9JANzvZsyL/zgOrjwHzThO3poN2Z4j2
5s5aGw4ZI7f6YfUxE/qtEMbAr9QKb+LSU6JVsKNRp3HOms84kyX6ldwRZPxR
lfPLqRoE7eWZZ6BgeGHIedddqkmt4tsUPHmFWAWNIae+M2Bz5NaBvutI8BO3
qWn03Buzx0vlb8OEJm227H7XMD26RKj60ewRF7Yph08CTRoIDNMbRS6Q7HrM
A6OOoVQ6jH0RBXej0Xhs3da3H8+hClN4szqKjpaWBxHr7S/hSndUOBnUe1b6
QHYBKdfaCK9BRm38e/+fHulGmvv/XBHIFgbc0SSGZNwI7iABtRzj9GJ3NvT2
pTEII7g0BoWxG15/1pNlKJNQ5o8WtBkZXOB0DFB/PsxGyce6RYaBQ/IuZDDv
CsXNFxQYuKy6Nmj66Q/oA+mty3klPn7eGtjREUEGzFgdhj1vf+7HooNJNOqp
rV5+oVSDsV+qlcCcK4tt/BL0N+uagNSo/tSPGOgruxb/kGWNUQ0N3SALL61y
m3ZgMIpGYRrxJ0riOYmonqZLuDUY87shRsaU9QDECIYOx9UKgGVWrl1gMMwN
PArqCNnKH8V3RFrV5qcK0vlnyQlWe+/CglWgUQwExnx94RZ+zALJ7bEkQwMR
V8O6XDrqTAe068BsvcF36iuL0Ocz6rPY7Z7eISb6kuWABZrt45iDR0KZDSyD
NNKxMZ3ha0K1bXMCP8raRs+8cXvfsuH+qFbil1W0iSqu39QEedfB2mDXpycN
B+YHIm+6jk42iipHYcQNPE3wkuRQrK5h1FHxFlR/NPO7nfm7/cfPGBfVW8Zc
uCa5HD6SWozja4cifFGZvy2QO6ZYXGZA/wDIf2yUEHqjJe1N8Vs+eVP1lj9W
6TYPXRSFztApjEyzt1r1W0OqJXsqc+S5MMou0haLtSQwn0NuWt8ZCs9KDIA9
3d/6MAfqCTuoF/bLwkmpVsCloAAGMowAoZxhXvxE2jC+JLurpqxA0iOOsrXj
Pmcd6tmB2STa558ay9yWEXYhdi2hntrPg//n9znAVufV9YsQhfddVHbqtd3I
G7M0gsmYqDFEkwCJ3iKmaiesriAg8zeLAw8QWT/g7nmBkgh9joxIEPKzgxS2
jbif7+tcZxJPgjqT7CDiXXrI5G7h0Xwis+sC84hYpG6xM4K55QGPignmeMBA
ovLUtlwEPsOQd/7u/681GTfnewgfcEM0XG1HiPQAiHFlnhr3PuDCAOfeB8Pi
lqOm0AKv01Eg6mSX3BJ5MkP5DlIpsfEyS978ZCokQbIyLr86qXJjm26mIn9i
bsd8yoGlu7qIiMQlnmZDagSrxseDRBfGzqAHm5eZCO6TXTYqp628BFS9mBO6
HKN7qkoAgtn2VwBFZLjptRnVSMqBPSXBWtnuLaKm7un673QBDlxImoCx271Y
EsrMM7ZS8hMAzxBcZVCahlTiKAgNswUY4TfBHDalcuFIB7MjPGggaMtuafIK
EcE8joWL7KZ4Pdj7ng9NrJQdca2lyK0PwDPNoFQ8GId2mbxaEqIV/bFirGI1
5nU4X1cPuboPj2FHMVmNSxzxLcrWun0oakXWeaI4HzsXbGAZc+TKfaBkCeXC
66rW/j2sooFAR9bmdNrvYAaLMFZjYabf/p+ZJNK2TZrUkEr4Vha+ZoV+/NiT
A8DTNF6qqyw9CbgdTui7IOypPxg7wey84vVv8AzHYfr+iAPjy07YPlcLPrzZ
WrlB70CA7aTBgCB5Fd+LZ0xotL8PTgqnMEBeVcKAYnKVBr/CbZrow6LpyVnt
iODsYvo7lwut0CV2w0WWxgLgxqbSGOSeAGiqnHqT1Db4YWITXtduec4vFGOj
DCOD0ZXdO35/T8vhP9Hzz8Wf7x42SzU3IJRP5lV4j8HXNCbakIoH/KRUm0S9
WlFqe3a0wqBUUKK2EMARk5aXd3PySxUJpy4RuWCNkwwQYZb1TJgSLR+0AkbM
GJ8nxsBgBBbbG7weEIslcWsbXDnl/ctk0rp9SKUWyT5BWs7mFObHmT+XabWe
h1SiC9ZjaE39RSaUZXEkLHAuhmp1miM9LkZ2+HDjdjCnILh5Md5vbiT1Nk2c
eToPXsSF6ASNzzHGR7GS6zXVsMuHkxq3dbkAgfdOi6miJ8QuYmIteUpvidRY
noeSI+MpzmXTwChj3+zBvFB/+jnygCni3hhumEuzkKwIhR/quHoWWyrxA1lL
U+wylH32PHiPBbwFSbvr+8+hrz5UEH9lbhaVwjyALRdjmImyAh9bIBgQXTBo
j7U5lMIkXAk/fxbot3Tg07ex8lN0MNybBkK57HvxJ5TJdd/lG/kx+HzkYRri
2S4I6K4CiNZwx5wZMGZDWq2DbBTI3YMKG43Istk+yAiGVXF5ji3BNqJmz4wq
kmRF+njShzuiWqQkzCcY4tJNdvRuAaCE/yf/6KiYtyG/RpF4+amHylHEuE64
PsAb85KC/MEDrzBGpGmAk9ZWjyopy5+beNDZt8j7f0VcKjQD4LJnTZfP5KER
mW3Xy3aiDrMfmOF1JBl8552f86OyG6NfEMhgvyjP5hbyqdnuBZVCHzTTJsT+
4lAd2WK5BdBL5CAJx5GASFsyi6L/eLHNeD97fL0tshAETsAZV3SmRKalZ8XV
EDK4Yuz+fOaWXNQVPUJRAbXxJm+w0c/hSoIYuWBvn65f2xZ6snTzlsKPFXgM
Geu9wgnIZSpQGu1s4g8yXcV0SvuqRb+LzCq3693uGbpr7nTw7uRIRXlOgeZ7
ar0yFKYZxczknDadiHGVZoaIMM+yCQG3BtyHiF8F3rtYwxStvp0HYQxRqF+D
wcWUnGfR7jtT1pXENaQgfDLs4buX4nRQp3sBr9HgmPqJYUaS8X/+yx1TyZyw
+iGK+6U40kgmdoc70RhnP7/ImroKJzqPz3xIRXFSql2LchmrnTHmE3IOM9cR
AZgRi2xheLnk1u7X4lM21fhyKUL/rdZauxsnEeS+V4gkqQxxCuOTQutn3nvc
dHvZDLCBA0HTM6wYIs7jaecLwKglu1KwGK2B2+ZdgNRxOZnfJXAGR7mdL1Fr
0WiKyjyOZ24gyO9aKH4soygNErPpuGy2Ar3iDkYE6eRnKkC7Xvl3UPzNp6FV
XIouXtbB+ZhOp8/7Iy5ZLUwmepwn9Z84VV3CS30tHZKI88O1Qf2ENhUucy3z
duXrP6zz6/PChsCrw7bJ9bxQCcyOWzCVcTYmlgO4zPTX0CN6EjiWVlWBghzj
73iCrxGNZEipU7raL0IYDAQGsYrAFF4LP0xpn65hAnhyAMmB896kGuJuZb8L
CUIkW42MswSsN4JuAv9ua1BbIALm6zThvcIyZw6YKocPiOfyugwEkVIh8ng8
8sdAIzFkG2++zRaFTWTEBcc3kpYClm1SRNdXqjAFLpR/aDk7n6lMAewNh7iG
FXbXCvXS8dTGaz48EyNaar3s26FyZENZjZAghsNVrK1Ngn+ELCp0Mu/1EdOy
UZJZIHL0IQ2/n8kHsN3jkF2+PQMZgRAL/MZre1apYjt06mJ1k1VGXBaTKetp
t5WWhUscRxf0ho/usvApVkfC4V8WCHgSxuWGPOPwFR7nQiFobbxZA5MZbI51
NB74kitkEcWzDxP1Xot0DBMB5LufbTh+AaLulNg3fRyXpxMp6Vmo3q3am/Ii
3ry5ePutpGvf1S4LdQB5CKYbo+KBl+i2Swhiz7cMDj9B8c9hnrpw2Mj+iVOM
Br/BSBJNRtEzsjRf7k5lHXtsrLUlWhrHQlc7KDHOg/is0XqQlioMk+Czm3zm
jGjBqqvDZw+WpUK/cxC2oa9hlQFbqlZbrBuBhINvgrCGO+asO1Ryxs2Fo3Qo
GQdzPKPbSy0K+rxaY+eU6lVUw/u1qDkCdy+8uMufxqtqiiRnMu07jbh5uXzL
rkLvAGX0vSn4uKg54zczVPQpITL5QYjO2xC2NSl5i2Op81jWs7B3wD3bbhZF
JGi39+MwwNwhvFwCMB7X2W3ie4vFSAAFz2gXnp6c3qlIneKgvg+pd/mgFYcX
80Q5K/KRon43xBKAKV4Nvpw2ZfyWUsjdtcnIQnTJSbiZkomEgYpKgPZjTj98
U9kXhJWB48JcidlcxIhpKjF5WTZjez6d/ln7gQ0hLpOtytuZkXi6RlyuMnco
CHrtxnYk/FvWG6L/4djjHFh14g7aOls4wB08Hyz0sZCWGFbIDZ0IkC/XBzUv
2gRseMlLU0lZazpmDTOqfUZW/IP3mW74Mq37pI9BYkTfMg5yhnckSPMic/Xb
v0yYBcQZ9lCDPB/3udgVL7cJFZ2M4r9r6OqF6AnbwcegPv0rb5m2n1kfBdje
FYMtGeANdObwCtiucfLsm5KxnveEWXmeUaqdKqmHqIs2Wv31uS6FpLrJllMM
hChe+rk8dLm8mZAYhKkh8XGJ8D115A6Ww7wcj0zDxPwtQbCnhdzh+zcJJCFB
Crryr4jtlbMt64gjdvntyJm6FRVyqjAXXXh7JRm61OulCxcbxq068neEqCPR
/b7POnNmv2XgcimTyeyuy9ipxwTrlMTybAOvy6fh707OAiio32g+5Di/hnJD
IGiU35h8RajpGggcN/I+S9pWOdHpRqTFs42DkdjHMlNW4zNzr6UtM5+wvxpX
NaoU7YQFWVotb8fEjhPm94/5tljMHawDLBFrlGs+A6BB+8dozo315vBx2N0F
YKei//WeMUDV+/I1Z2LH5Z3NwirO9vVZfrfBBUfKx0XSqdQslamxZhepEg8h
Ax9KKig87BzybDmHZLRDYodxvIk8KyHhAXme82TnzL62Ifu6izZED0FUtxwT
iZusa12ED0ayytMyXnmLn55t7GTEhyj/d6Wo2gypN4vAzUJnpBarNT+iR2mz
y4x1oNCwNJ/uB1IcE5XMGto5rRNQJIYPY9a2pZIS4MZrA9+7s/gov47M+73m
vRPSUCNmA9v5Rcdpz/fB+j/P0Lm6VCYMwHRLhY0aZrD9+3x7pgqRhLqw449M
bGsD5Bc7FQVu4xa4vRbvVxAXogFQIrZTnaFDkHSXEF7yUsKxneyiWsxLr7p6
2oPJpuNl4ksj0D7zpUyH2tSUuy0ZQfie42jyalx5r1w7Y5csW9/y43iVKVKH
Qmk7EHv3N1JpjsyyV25uzGRkzXnuSEAMsNzZBYgdU1WpQbJPZDHTSWUxbHRP
YagDKM/JVATKVM34sNRIVZrch0UMpqNc/L6ySuMNbt76JnrL/Iesu7HWyQLx
gjw4nSaRakQlgeg281kYeJmbxihQx0ktwJ8pwWQTrJ9PYm/pF82kcM1TLX9U
FGgzcCWZ+N7UJiphURUSSsa7miJaWNgiEfEcbMR73cRsgsKyJScbxyU4kEpv
7NW1h836/zSaBtqvaFLGjvYAKU1Y1sq6Q8ck/mcd0UZIpKids1HGeGjOp6pP
uo3WdX0pag5xoyrothxMqs2CnqmlwEpYnPvXZi3yaGtx3/LvKJA6CI5EQ6k7
n9fzuWZgJoZk5x8P8PjrcesOGHcpPzE06AIPaBW/6PCzNkZBG9VjF3dtWB6f
00ouw5eCrmO/pEDai0ELb5c5VOyV2S3XtCkSkT6pkp+WlNx5IGGkndSQTIWY
3oeg18+eSiJRtQ6nwhIyy5xFaytXp1hse6Xrj7cHq6hL0VmNQtI/DR+cNphG
evkaNVQAS7fARrJG1DVvtiv3uUevu4evF7NeeIqDVDBvQfwLty2DGIZucaqK
5pYm90u9rdvKCun6aSObQb19sdOtqluJJiBHw46AcMY61SVfGtN+epyAyX2T
nSQy/PLSIrcyiMVtmE0Tb64nof8JMxGtj0VXpAeXcTqp+6lzdK/OuF19mGgw
tlzSKgEBc6+aJwwG9L3Xsc3+9bt6g5fc1EKOxUMUrZpx0bAHzkcpOA4lZELh
Lfw5wcomrOHIG84oOWAPcVbksF26VuKxio/QOQDLn35IyXLnSY7w6iXSl8la
K0pQ02Wh2iXwSKeJOB29Ya1WFjIWS6awJy0sAqG+3qXsnvroAJIJdQR2FEkX
7TGCMKYIgUUbnFbDs7Nv9/BaA5CQ+hgFrueGRX0Wo6oNfUAu/JDHmh0fCTEq
umdrBQgxA+BfAk5HMpmQBpAywDlp33oO2US+iRaEziRHzuX5tdW6JDqRyxut
c74fGioKQjtU8GBF9vdcc48daMNw6LjMpXuPQpflsStSAYlI6OV/W7Y54Vh3
gwjHbgHO76NbtBHk3QbK/SIjzWtyYbz8za/K4l6ANHIOn7SpXXGD0BISN9te
AYCzZQUpO5JXq1x5Gov3n92ud6IuqDzp81c3ovjimO3p07XTBMuTHFBY45zY
sxNEOpk54vtpaqVniVMBhM70HXjZ1YGoMpFmKK8GCcF5YQcvAlcf16zrGEJW
UbJ7JB7uq7mJRu/hjoMxBa5CJZHaNN7N2FiL72Irgr1Qwmm6k1vXUN/pjQby
ZEyH1kXTTrJvw12AW1IYIJVu8Eb8JaxaAdNFMRUDzuXtdArFwFLV9YqJWNC6
QliMUUupfHws7sgMlT1y52ww/0DP8fLuRjG9VlJJAmf1SC60gwc6LpnGjPvj
NjwZ+OiIW9xeCpdN7r1KeKmTdGdhBvbIA/2ktBw/XtCJ2ZiDB/bi/ONW0Mtf
n2BuinGnVheRUtZGETSCDHaV4aozGDhAdh8sveDmdSpTAwOeZTC3N35DPJ4E
ziC0MsOTVWCgKvYTJ9C+FcTsL3f1G2l5Q2eEzkfl4VKeZ10nULqooLJfwPAn
pYFj+fTCZKFvq67kJgZfRG7Sy+mfjqdyCJUxITkAg0tIv36X9ZRBRHVljs1F
RTWlcwttyuWhq8l5DKb+pGDfA8ltOWkAr68zsHj9Vg02Vi+h0achYt86sXeC
AQjCadIq5r1kxAz54JOOKjERRXIcZnfXF+7I26urxUYMQPUZvT/m6iNW7q68
vPwovrql72zRuxdEVRv1YjC+NBc+0ATJ2ImkX9ebR1bgP3rlkAzhfJ6kTzKa
PPiiqezaXUnN3Ju3KobNbPGwvK0rUsW1iKjLBjoqW77bpFJXg6Y7N9itfe6v
39ewtQJUSNPaJK8k0B+IKBGQljDsubh7nKNqeHPwu4xoGagfPn37n/vcuk+5
kcKItuwqcws5S995qHactabrvWT/8GxnoCpndwuJgqylBW7HiFccHTTI3qBZ
205ye6xS2DviiOLPnx70eT0TMn/v0Ol/mpEBPg6H506q1KdFshMLcP+4Namv
Pd7e3MDRzKOmGrTNm6vBFtq0vp/HovApVq0dEyWzaYw5B4++20zm9iAe1Q1n
GxFYcF4V8Wf1hy/kGxvj1Om+TLJedrk7TzYU/ve0uAr4jAie66h+CXuU9LAY
DJ2hnBVspjvqB/28zM9LLlwHk10vp3ARFMHFj25NTJZ1clmhIvlLMYWsMjqq
H+5COa7sSMQpHagF66ipIwMHX2aixj9pu/2amM/mEmmKxlqmM4ke6HTWqkCQ
44CVLmXICRWHWF2YdV9fZxF9hI8ffQyY/qcgfv3NYGtaPhe6/SvUbbghpiAd
6LE/NsRNdZfspQ7kVdDm7a4A4vcHR8p7bpuLwltlVjUsLIUYN3g0ds/ZypkH
FaLwAENm0H5NieO6zn4Se9QA7QO4FILxUTsvekozJZjRlPeboTqrC1C2RbzN
TyDXmf5Aks+c5ceHg82aojMdn/7LNGXkYLl0gfMPHN7WAygwCtSMecRuchz/
QlSCyOV5e+vPBxFXfp11190zJClKUF2SpeafN865w4UC/fKCH356art3YhCN
eSTqGpfjNAHp2Ldk6AJMZMWxvg6Ejbb1RIKxUGNaFp0e9FaoA5AogDOAcgs3
aFxNvww5u4vVbhDPb7sCHQKpSUgpTCqjJICENSPSWsbSWMie1ker2jMAnNCU
Iu5VndtMgG3GMEr2B1Zqxcn5Fys/MfwaJqMNd8+NuOl9RHFweWDntnJxov2M
XfQjPqrKTWPvwSiXBwQDcT9KvuK+SeUjFhgZ9EVdDrVMi8+jp1PxxImlLEr5
YTqbiKhsloweWxDIV+J07i98qzLFT4DRSYZdtRuioYOdjbfwFMcwTOsDc609
miyPFRLuyXQzv7wiMHm9HAsYs3VI2PhuX/dL+wuAzl7ctB2wIcPnfy2m8ORF
bOVevbP1gKtY0eTyeG0E5tDpQn2XdZle+XdPTWrgtcdWbNCBBeshsT9MzOMN
x0NJn7b622+QF6ozw5wlkqz00unPQZcu8IayYTua6x8m/2rEu6kmcjH1/8O1
EojKf8UJF79K55Oh0yLT2FxKWti6WJu+ZUD8SAEYD6qjITACQQHTUgBZA5ZQ
8JTYyjuolWlwIsZzvEtY8ZjVXv0uacSo3iLnshMRHfw8ndGDv/9ArV/jFdFz
7k/8TCxnhY449UF07S1jbDGm3Z/M6c21jPt3zQhv3HSHeH9W9PL92xFOU4qo
+dmvUvW9om++eOeAgRpy0mu1VXP51WpgbEyFzVBU+4ht4K4vsTiAE30NPuAj
IZS9DAtXyHhLFrTiwo/hOMV0hPxbDT+8OLgzcU0EaIgc3dpe7Quu27woecp+
f/DiLS4wet1utSue+v9BzTrxMwde39zn5rK+miwROSxEMkpVweH+gKg6IR2U
qHN93na6RZJzRfmK0zQXxwoFiJ47eO2xoToiHE3Bp7Y/JdJJgFJ/v2AxWFHM
1JxuabXtDe5yifsKKrbGa+qg29sqqwkqXnNzxFKfVjeZ0iI7p1NF3DrKHPOf
k2KgwB4SV0EQrWCJwOocZAgwzftAzhWk7QXXlaKsGaqStQ1tmW4N0PKhGmYa
nYCHrqw5G5hKVIVsvUoO+sC6wiqKfs7KB4VzGZrsKc2QeUcMRC5odkz5Gd/B
jrgRrI7hjsUkEoYRqxCUNmU3fWVzxNN1uK1TGefElJnsG49ijrb89GgnKRky
MZl2zHaKBHAqF5TZMpeOp6w1cALs1+XJxmJot5jMQ6laexZEZbI7DG+xFzEd
8BgR3Xf/bulQm78tGJcZp4bNWoYRrhd+OWT/Fl1odS8zBs/mnf88EM91w6aK
0SxG70Y1Noi36qhKYlB9FIR1ozO1i9d0JtXOHE865D2jd4gqNSXZVNxiP/Uo
3AjqnFuymC6B2nKgkAlDmj4/IvPQkWXT2la168K98ED792uxg1bpHmJ2TJsW
2SZcfWErw8l/CujlOVjreBirFq8o1J35Sg7zbY7gzbVV/LXp8FFEYFzgQX9p
jzF3mfihaIBhiFv7WO1fVC6pvP+/BZUTGiqqc9woqyZmBKtPwp97nMx8qHX4
jiT2qTgKVpEUZ7weMUtnYa7oufXwfVDVyTovgM//sz3UO01x9tVi3bzg9BWb
ArltZJDC1ebeVei8DHX51F2sftKdzKp9CFO6x5jZ0oiLV1LFIW0qPiL75X/V
YGhwS8tQlbtOf0fhQOLA63zW4SkdaZfU3pjzTYwl9KB69VBqhkXf1uwYrM0K
S+GZVdf6Oi95QvoNz9HpuESf+tvoXLDnR+/J3hUic9KZYM+v2iXtKh8fAok7
VpYiyB1e2V9StC5CSMPmEyuQ09aSNoCDojDcPR2vSnP68xDO1mYvjByh7VwF
ZwO0F0uxbS7r8f2pbUFsw5Zd+doQtDA4oXz81FySm8WNYDfPpYqCLMpntIA0
wRxh+0oeO9RLTiF9veHPrAdc31V3CIjeQfHFqOuKp7p55Kyk6TZSkrWk7nrQ
Xmq2luxdrgT0HVnFxkRy5/ZrCgAgd2VdNxck0LGF4bdtVVcjqyJyBI3gP6xi
yztC7B4zp0QnXrC1Dl6tPMnwQuNZE6Ax1wAaSdwTRmiXt0ZqUHW3qCHJijhH
89eCFhZE6KnDFsSZdkvX4d1r64rHjNfGc59qH1pQs7xsfs4QCbSmjyfs0AFU
ap168In4sIVIuNyuE1NqxGdIrKrjt/HWtcOh2w6c/aTn/Za7EhzKcmJWcfQH
VgKmfJBREYaOORo5QtHClKvZUw+fllGj2MUB4hhgTDlCLlvoKOHBwrIiFqIG
HOycXOzGru255LtzXrB3IJQlKr6WN+2ltNpXkie2n3G7ZutKuAq8jjC6ydd3
j5rM2+GrLj/tbEGVBJWRy2fNMhiXR60AqCjzpiPnGUU4cYiuFJ/4rnaSmtcb
SUEfK3qdoYAPLIAhR//imYu+6KD4Is/F6WTUv2VtL8zPGiu8cQIe8/rrs65w
ZpPvX4zQ2VgXB4YI3t25BINPRQaX9Iuklfgr8dTSwf0LpMhU/ck9ctNpmt87
dff8ppuT4rKWwc2TkVxcPS9T+w/cqjV20JlrXD4LrC2wYxxrR4rWibfXvb8O
yYgI+xLYQ8V9+PZAOh8uHXPnOJ3YslF/EmKVGjjYcZ/xLMu8acsAr5NPjrUB
Cox+OJw0SaUKm4h5OasDPaTA9FBD0uo5/f0mcGbpYvETUmZzJA0/Qb4bi9EV
ktC6fyqFK6MrHV1NW40omkorhGDhUIsEWGV8ZKPbluJMJY+vcyvRD0AlbZik
I9NB4j806rF5Quayte+j5DW0KzEPbrFx1LP/njXREmJKQNw/o4z6oO/G1dgu
UDzabH2kCMB+MrNXrf79BG1Bo25Fo2ypWht73ej6mRyi9sHC88Ly6ACAxhTc
Lz/AjecmeSL1hnADFxsNdUKtZct93X8MghWZbeIJ7vSuVZEWfs9CEQiW4uWh
vh6vjguL8CnOdigXMMHbtx67HRHx9U67K1Q2yQ66JEDmcO6si6XWWgx/QTSB
C1GoXChvXEdQehrc5sVkxsDzL1/W5z3vBDB0V+LnK85DRNJQTMWwsiSFSw1y
VgkOt0fiHX23wiDGI6HkrO71jVDqljNOG/M7CJS6VmqZKapOILg9wnCdAR8a
KO2yPfylDkkOoepGNQwOzvlrBlPuUh4TiHm5h3aktydMZEhi1ZeA8s+BtVS8
lDdM3HM5TvJsJFQuSLvbUNPNRLztFbmoadYBtowcMWzUj+wt/nmKhtgUCu43
BCkCLfClgCU7i0HA3qU6X1j3i+TVLE1myfF8fLLLNwRN9mArga94b+tiGFqy
UJOOTYJRIpLH6Ez9EKTo0xGE8rp8HWyixrknZ2cRxXne5irFgjR5aitE5MPw
oiaMjhyms9S40rjkQLFXBP8QiIiO3u1zXoRNgP2b+RF1zlMN/gSdfQdupR19
+3r2UtrNUCWsPyylgZkrPDNZfIzYsG4Me4hV2F7avMypG3W5v7b96NmA7g8T
UoH3LSFajBe5niRdhN4Ovm2NfNSlpqJTKzJhAIKpmBwOOUOrjnw9iHWiHoHE
0T7SMzXFQn9gu12WmGvtKbamelsTwy6tlXXsgs0f6VTui29w3X506blhVArD
/ST4Nh5Ds6leaGrr1kM/iFO9sQAWsX5uMDareg8Gf9Q7RZz2mRlGPX3IOEAZ
9vBwCyfUIAU/a7JHX2NIwk7jLvq16Tsu1o3E5foD0D7naGMX/2uSUJ9nhM2g
jJJU6Clj1hEPyOoRYKofupNNn4vFyLq5Q/O7xZlu9uaJqO7PJlNa8XrWi/kb
iihVl/W9U+eAlO+lKeV49j80B28zKodby5COzsMbi3kfkwAJ085VAfQAjTMn
PA7E7T6LqoYTdIkK4vINEywBGCOiB51T79R8mnA7j8Qi5MBHq5vBa+b5hr6y
Xs7m192B88X2BFz0JOT5GiEBeeWc2KNT3TAINNYMx4wlsDwT/nvFQ2+/odD1
xOuxBTKbjDsX1ddZEAualsk2zaqGwOgACM4nZFzFfv503L0cu0+VD3UVhZIN
M+AHsejxd/tpmvi19uB1uRH/7G2X9PTUXQriin1nQdOeuBuWXWG+2j9RPvyp
IX+PnQyFT/nz2dbcOS6CwZhTjvP3Jgk0z6kk+NgEBVp//FIn8aVXtUaHbokQ
aUPHC5z2TygRK+KycNiIKG5NW5v822D5PY9hOrwOEJ2t+wBOz2Hc7ljEk7IT
y2vUFXr4UDMUXTEKwRtzMaX5SKjmsOIXrGoZIHDUJRUf3Mwaa49STnxCslMQ
siFAAIdwNr9nhleRuYwJTDEpIyZKzgJI/wL8D8zrIxqqHnxMA9thtrBcfem5
x0GpK4jEFcRJ9KuqCEpkVewxhx2L9PxLUNUPMcGhBvMNFDW8rZywZY8sG1A4
L5cQ6pTjyH6Zfllv/USNcY4WJVfYB+ufhbClhOlPvaY/KXTAD20ugwjbFeEE
yUnHrDEvXX6TscFNjB25SLQ1gacOnYC77lgFWIQEdbxxjnFsRy+FN1vT9EAn
hQh+ouq39FHufrrZfqt+Dj9xEKwCQWvxUxUe3jWA+u9f1qVHGDCbuz6F3KRz
Y89QdU36x/nZ1ujxVdFskwl09N53AvUPmwKL+Nnm2+ZBKPR7BkICa6G4ic/W
K8Xe39Fa7bzSxHPm7Ul0VUrnpIsSy0fpPHF6AodftU66o0qee0JIkz5ItSCs
jZ0ujBNznrPWtqi7xl/7HrQ4AoMhX7dnAfEynC7/jD+J967mOIOwR5V6LehD
ANGLxoxcjI/lbSFV6aHK5Ok3+r13ra2uk70ggd44QSzwYUNfF2/CJ+BgFp/5
G4oqaYFSDi+PaZlOFIhq23froZf+RMH+Kc1w1z+6R/Z0iF7y2NvNc3p/6k3U
UM3HoVgYXOchKZDV1mkrcN+QZFlixBuoBey7mTyyOTO0HygtYtveVhGInVID
Fbffmr82C1cI62vM6NbENw8ZBq1NnPSQVwTkmzFA0bbCvkDQf0Kgn4q0GIKc
yVDaH+V+bpaTH6dNHWljjEeu1ogTCkLQgkTxhdXcGY74HRbbl9N8hoR8Hp9G
B3GSwnDJjbqlSejZSuJLOKc1xcELqjUc5LVmXmSWclXr4LHaX8QQHLYFnBW9
xFCOrp9eA12sLi76t4oKx+Oy+rb61A5StudCMU3VX2n6ehfppgKhi6hINLvJ
NDQLJROjrbeYMwWbeDkit4CerDRsewdcs4kvtaDirliIcoT4b9LcZl06lkTD
/9oZN2qyxgPjAd9HbIUQYFL4vYZpWtFYEUD9EzFA1ELHjNKUxUnH012quFNx
RHOCJIaJp1jds7Y/uWMoDGWkEXKoTjAa8Rg4XKa39DSe/4dz0Xb+n/QbuT6n
4P+qDEtQuOccHuHlZiWUgXNEP2PobVm09CrFlr+wLaBKfrfja6KyajG/aZhO
riueMGdeL5uxGTqZ3nvzBN9SRAUPfcUo622nOw2CjlkmX+ijre+gOeTGCjTD
UjXi2kdu88zpWK9nj/iyZ4xMix9RrK/3i2MtsXCgnjINn0OEux6Vsrb9Znyf
0BQqyDtKGmARGdMITJsXIkSoJGrwcsS2ehzJVjrreOT0niwySH5LFldeOkEF
hNkGxwMKgwvZLjfJoWjdkA5Uw75EcBDXaFlM3oHwILUECI+FU4oLwXOjoLp3
DMaCUWSo+Qg6mJ2+vmoHPAJ/nI2HHgoK4hZtxBks0VLg9+M/TbweS+Nulw80
youMeuAg6tfE/M7NKpc4Pkk76xfiGY0D5ggSfgIY4ggRBTfHtAKa6tnKZZ4M
fik7mSAw4KSzUOu3D2FodyafS4uNS7oinjHdxzahJ+FBFMpNaOK26mezASsR
wBtEr8W060ytbOTKy4MNBM7B7e7wM1+/qzxUsXxKOXy2igvYmidAEeFNVeAZ
cV1LQSdkwTeKWxJbNrM8DypDux1wBmXS3ORYhdhO6dL81tndFXtAUZV8XUTa
VeHjzWtE85VdEi0nzXaDU+EkijPwlDnn3Rh1YlVAF7XMqfMFGkl9K+bsfWYK
aaQMKUNkr5b6oYQ3HHrAJz5oh7+mYsNIpUgTbnf5E+DZ5zKmgfgSafi00XEQ
PeFV0Jj0ZVlfcwnctCnM6GTSgo5+fZGWIA2Q7+J4p6myeADI5rCf3m8P8vHr
Z0bhOTrbcUUdFcmU+2AhtnCpWoveE60mZsXrVXWerg0NW1GLiYU1zHBj33u3
mj7ETxtJZfYe6OLzvsBukUQyVG+XdXJyraHGSfOmNvWQx0Ro22muZIiqzsH8
6/5lAS3GKT5Vm6D3zM7iAe58bYHiSr/xbOrkM2CXAv83Uwa93Q5/lMI6iJSn
aucrJwxjGCY6sO4nZsniWBzx5Yt64DqU0Y+jIe5lFUG/ypDT4JgSEJynjP7g
qoKpC9v1RAj7ZhPBvdkfoBfi0qttcLm9kNFedwI/nOnDJgRilQ69R1Aset7K
TJsyGajV+6GafeFDGAuKKNHxSz8Ru26WIRl5cfyoHvP5oJWbWzV8c3P9t3gn
ccdz8RN6oSlOMlCTUxCmm3QOMF2IR/BpqftamX/lOvQ2MBw2AkvJ5fjaY5Y8
jIt7pN9ZPHgBG+qOAQZx0tEQRrUNvP5u5sxu97z0W6ptTxJKH9olGCeOvAxt
HXgmR9VNrSqAQS13Fy5FkSPE8mYbqXnQgFNOQCWJuwBxcx1j+g+5tlHjRe+Z
yN/MfhWBxi1LVt2S1+IVedyx6s/koAczafN1V92oqaEfSFyyb31VgwsMWNCp
uZItOUH1wJLWcnOL7d18iFW9D6+qFjm+/CSGAzUzKLwqY2hSWYQYifHpJhx5
ooU2pV9ThGq54+CragrZyLIAs/dWzdmBKwkXgCPs2PozXVLlI0o9hnT8Buvf
PKAxnVGcQ1IxS4gaP/MMmzNjqRGr0b847KDkX7loE/CxsgwgXLtV0sZKKzTH
wh62HlS8tP3aJw6g9Bm9qKy7FYuVGMfMnhQNoeszgAR2Y+ScufJccwzbZW7l
yOebeh9fgHKuLNVbZjOODnNlajyCQrRMYQxHRnx5DKyStRmN1NPMIvwut0Cd
ahtEaoCRqir9hFoN4EQD6Z2vMUr8mSOgblgxXjuVmf6dQ7oqhR/KxdJZKl+x
dXskSpX/TqPA5ioF70gHhvt3/dl99aDo2jFnwkLzi1QXr++vIcl7vQPTyawS
jj7mLGQAbc5cbHYZLa9KN6vAutzjxIR2df9mf5X/Jl2IaMcCve7KcXAqMt1X
o6ToTief9AJrk4yuorDbZ4LZGMzYSnxGLdn4qhV+KsIYGigFd/j7W5oinZzh
U6Gh4O/gi30NMwWz+HRjpgWHN7k5mMUcL1CRh+ghlE0Ho09XLPQgM0J9tAVm
GZDK34RzC9K1zCjjuKMiMcODkVWn/+RR5keWiGRFd7G4slssk4ltG6wC7gE4
mIroe/tRoOtNfo+GW0peq1O9+YA5TVbScYUDRhsTzoyPxq8lNu1Z6iStL1tm
Uef1cLNTm5ROEvI/YzRRBsVyR9LsQFtg5EaP3NZ69SMtHvUiBsyA7wEMUOLl
KtcjZ6wpi70f/CTKo02KLRXXulTAkbt83SeOuiLNcvd26khqlp6ULbx1Foem
+M8oy4MyTyXVfP7jhQELyz4Mnbz/T7RpkFPq93ZZ10nmuQk4NcDAG5YUqUKj
wK5FNlWvlpCsU6BIk1sKvIvSBPf8MQ36BtRvnufFaEIwG7PmzC5zCH0kUfmY
si9egyBYuQjKHfGBQlV8oqJL94YkPG+ceL5htjlBa9qnFQbA+kHgNCzgcrtb
Lp9Kwj7HuKE4RvNiCiqgBscQ8X9JLyMSi7/2e6yKkAh8UCkCPd0Si3At51DS
GFIvQWWV7k3zCOHhmGlIIEPsymy6EXLK1UlcnK9EPMEJOpbAKteRNSUDMOYE
5OmKuycH0EA5RlV1VcgGNYOeNY2eJq1NlNlyUUZUoaXDOa8MZ3RjfmQcbLMn
1w/sa1u4SDrrU28gr0gkDO9a72FUycZ2A4GCOZU1HhCWWqRYXrD/FvauFybd
NENf3udnVMr0u+vSmEK3O5/XHWeW6JQOLp6Yxl8COCZee7rrcRVWwhlhWM+L
UaPefs7cfhviCdUCQTWNdlZEBCSjW4JZM2H0CTn/FZ4AEjjoM/j68EtfY3Xz
i3zR+TkroUbPZbJ16oLvWoFqP9yUeAxpNG4wxb1eJwBsUVzUjTRhNngGKPjd
2QvZw705RU4lyd0gzLJA8FAlOJq54MVj6yCFPPHTrGb5T18Z6pLy6Xn5Tsch
WVRsYxdaLWtR55ivKY/ISw66b6Z0cofOhJSg9SdcW5mXOR5tpLJsJvHuiWzu
dNL/gmnzy7jZLHkr7xG3PtX76/YNYex5koMgquM9lKyfod/xzNI/VqlTgH8Y
6TYHX7NnaqsNrLcPxx+V3iAiRbTy+KL3DuwjY1Hg+aCrNLr7sJSIvgnSWfTO
OZADZJKLV3DW9Sk+sjv+jVR6gpq9YyflEfwXxPlmpP2DT+JJRc7qCj66a0yK
qz5/kuJcu4ZB+23y9at+VI6EAMCFrex4rSjUtjYgY+BRK8wvrDbvbah05D25
R9fFbcgEhaf+jDYc88NnJcxnqaLiUUygMK9lAon8jp1/k/+HGgNc82POfNZT
79oBoGPI2TZXPT2poh72nbX4qLcC/GoRYqewR29g1iXxejWqA517CNJJWThY
5wMdvuintsn1nnPGNMALZlCnbxirH9iXSQ22MfXY9oEPDqRMHw1Z/Q/djFEb
xep7IHGYHcQCqyODtjjwlbA2ZwumRLMUQu+W3C/ScFs4hTrj2a2p0Ev2q8wV
xI57ymTCEBMs+OJHEgUl/TJSIf7kkU2Z9w2Y5c0bsv45gaw8+f9izSA4V9fY
XPLVlk6+lMkz2dFtbbiVCf0EZf0yN+Abt57pQ/tKblv0k8c+f4PDptPDR0G9
7QsPRC4r5T3+UcP9T3zifGKa/M4USCwsrxqam3pjpaFeVKGjCJ6dvx8pOLxR
rSOKxnNnZ/8CCqEB7BVq80RjaBaLlBjyNRroesKxO2liLVFszNRQwuRYhoqV
d9YIXR6HMM8H7AtGOpQgbl6rEEmlk7imZ5lpDX2Yvetu/pdHb72NXUxKQxjQ
8Oxr3/tGFOBgDiScJ9mwsRIc+yH23vg7JbGsrt5gLENf2Iu+cMAezvWoVoGz
EEi/YeOwqLJjR8xul5Y/WxwJPm8T7ie/HteItzuZV/zK+OQUgTW6ihopmS1j
dMDEq+P4XlW2DGQIcvoIS3j999dIRzeBi/ndJNpd0mvNSgK7QL7lrnmZ2pDv
LuziAUSmaX56hCdb1Y31LotZpA5EzRoZ7ORnIXUWqS+0J3PS1f2b+lTJjVU1
jHvTJcCu8tQ5Vit+sQT9WzD/CdWJf0CcWLh3iCLEUXDPAeeMXvcnDZXPrMdK
ZsOy8GwN4agiLhjWHPqvXS8lX2BGtKNeeaINdce3bEjWEYOeTYbptgN/kKsU
hTi6hq5Xl64X9uH4s+HIC2JIBE58hSQ++6KbHN32yRMaKSU43Jv0HHwl0LzX
KCUiGB1xeZlfIPKIe9v0UM1hlpHMlzt1TH3ruMIpHmhG6Kzg0BGyU2bKgkTU
LqyA8EuCBpDOIPeogaNF3NN3qR8fjytZdR5284E4v2XLmRilE6YRt5XCPMDD
uSi7Fny2nhAMOHfT7b7DKJT+9R1Op0joCxOe7+FISa1mRKHhmFWuOGBTaYoB
lt4dEM6rojuiJ7STOz2k8H2+aHsV5Eqhfr+C3V8TQ7s3E0jna0WuF19Fesyx
+i6n3sxlBDYYXTq78fR53U+eHoAigKeg4+/wvqciesvPa74PFMxdasUh4sEG
c9aWwObHl18k+UhG4FLfw3DE5MLvS+T7H6C0PKXG9tPRcB2AiiLk8/O4GlKo
lnxA0A1nEM0/bDTiaYjTs3YZ+XDqbupmh+FQfOkq8+4chSqJgt8a648IzJDU
NbO63ooVP26je6i26/MyvLQLqVbiTqHc6YO1hPMit7kRidRk5nawkhT6DlOF
aaH3pXsnfy8sPCP2qS1aB5/eIBC0EGt/eMp56LLAPI89bqeGFvxTCAWqS39e
Ze9RYpJSQ8rKrziMyvLUOI7wB5hTAgUIXMSlQm5QTj42VtudDnU/fEmN7pYm
mHsK5mbHzdexNtCgw5MlQlbFQSflv3Hb3UDNBX6pv1oTxJj0zKM1bC+si1ls
4pTeXgv3UfWVJugMtKuYhHQFmEHKrIIke+xYiaekfLXnGhZnl3UAxT8tqZp1
UQTo68KNC6bN7E0KGEDqeB/d584oMjyo7vvQiIuY173n3Jnop+xnNQ7tZ2jG
VEyBS7qcvRUKwVm7XZK+/g1bcw+x+Ig71sn4I8RGmdHQEMMQ/s+ZTLC20u8T
tbj62W6SjIxTX48gHAgg9qeqOyYKDBAHxyzMlLT6GR/qhgszPMyMqALv75Dv
Y6yVEhdx9H0IJlSGapt5Q44PfyN+m4tby28tG5k90JQkmDbzb/vol7VlIL3J
8Lfwl4oyq6WtA12s4Kc9grMWwRt/gsidp4GPUQJkMPjcpK/EY4vqs1sdX6SS
1hnIWTh7pw487ASi0Xl6QaMtH0tXTVCt2LR5p7KtDWazGj9aM2rrXuYwlWGH
zjLEJTnJzKA1WxngImJClluYEDTwMevqmWenw4csLScpxUdQPZBuIke9wWw3
gQp2vG7X9Tsq6mchjBo4AL3WlK71/Fg04ZeVRul7KvcfJ6wSk0xj6D8vIhOH
P2Lo3kVHvld9W0KWZA47gVTnSVxKvA+zM+M3f0p5UoRRb1t8Bjo0xrDlfCiH
PhsO/UefI2qtPb+mRELtDjyM8vkfMi3si6y0IBgoVBWGdrv9OSs1O/qZvVlB
iEoHY2c2Mm0pI1aqJZNbxPMn3rzfED5j4tQ0bLJemUFWKNB6RGDKZHgDX4th
mM8BHyIOUCjSDxpB88U8OWyXCl4t8o8NAIwsOCMVsO3EIBgMAThI07YKYuXU
oxpVeWJUVjwzsiTe0vi1iRyiev3ZuT2ZBYSQZFhT8vwOTm3AZ/HH051fZuQM
bxbt8hwrmjBNtgPU+cOBuvn5gEaZth78OEJvNohidMjStGh+3v1NXxXMKzv9
HUlgxi0yxGaTPYfQQr7M5Ggzck07VPGDIJ/rqP2SABcy+qmmCwxB4Dhm12u/
PT3OsPheht1Oa7TV+v3C67BqR5dspp6qRBkMmTF3s38rfxIHNsz5rzkfHmTw
xs5tZA4QemKz1LpSvHkOOSzv9q/pHje799qTDG3k0aGwbz1N6jbWmuI9L29H
sEotyt0igiX5dOH24C7Vp/JjO5X5rfMY+UdTaykztIIiLYNWOcwlzk01EBNX
HwqHllsiCI0xI8jh1FoNTtQ8sX2NAfboUKHla7c+WGJ4n/RW0eruEia6I2Kl
O1v1O8XcmP28aZ3VXn4G1L1XNAKey5f7uErwHtZl0JrSF/DNcugT48y8G+53
6A2i+hfIVBcDeOFBOUrwF8VtxTKqQ1SJT+yTCj2frRZOae+rmI7nLjh75d8n
5QKfEc6cgDgXfM7cLXLixaXVEpEHd4csRuhsrG6eM3HaT0E5OceeY+A5jneA
Afwvg54jRn5FRF2bdJ6UPm+E4mrBCBzLGMJd90yRC6h1udKXZBK7mdnCTzuD
2sVTtsfIenJJz1EUNmRtr/pJQ0cI0qaljE+ITu++EbGLXwNka+Oxf8f1HMve
Ftq8eOzM8pUL0T+jQsyTKS+uHDTopjr0BPzrcc3IOy3/MIiE8lxy6FXS7zjP
58rt3Qau4S40Gt0xNhq1R/9DxJ8s9jbxvAwePYhGNuTqmz1IKNvnm78RzxDT
SLUTXv6ZmwB8qLgmZsj21M846tE+GbmIk6veiGfXIqVfnPC2pkAVV8fdS1es
3VgoGECzYgtSoXtFOCriX+R2UVDNIDPQJqfxrDQeQa7qMjlMOfoeuKl04FFQ
rx53JJ3r7Rau/vwnrnB7e/tQplyZt+aLBGfAFDsqEg+EjlR9cw0S89i3+M4P
BbmOIfd5GEGlFI2hkk+yNBj+iFmUTivLsJFQjXXXxUIrn1COlZu0C9Hj8RCx
NYRoQogEDvImfMEs+1IWeZLL6hCGn03lnkHCYRDFBcKU0lbO52m0+gJSfmNF
ULoWGVhKbKoIwsXSm7Fx9QQMc64+j7i7CE+obVDiKvW6x7mZnKL6p4EZjvPc
qFm+tXfgrpCsw7gqiKYqF7zh1lxUWdXI0cH7uS1xMgxTYOzsYjPQfzml9yga
9D8VbiNznWS9FJR0DrfLexyGjqWvL34LKHyaMFfs6jXcd4Rf2zctIqNew3J+
KF8fOHt/s/h2RPyjDxKsjtzeswGWTQrWP8u1aoftJQKLZD9WBtrJ482sq6zu
gWAbujDJp7hJW7SY2Nv11qYa5ss0vRbY2PekWDeavO0Uo98ELeUnji6RC7ze
gD4TP+s0Ot0nnzr2/zrFh58P3rWoy1p9Afw2+ZMxTfnKJjY/tD7MD2PGt8o3
UfGhtWcms/k+y8nzl+3k6hYE+YKGASusWuZqKEWObTvG/4bQ5I+e0YS0w2Qq
3PpAU9qAJ6yycwDu4olWu+bvqH7M+eWe/sx92SSrfpB7KTy7F0UqGgNQaiar
2h/Maj8FS0EUGVTOV7xpZcU8d4LQAkwBnDG7pkkwQYZkhwddhlP+GoUTjnUw
Hu7caK08ACl/UO46DOa9kVjt9CbYLV2eZRwfAoDgsS+af9dqdvbPZ+hA8bOH
abHXbzpai9/3bXz7M/eUV4Mk/QZYOKOtiw64NWNTTOCa8AnTiR1wcCpqC2vp
2ybKLdLkQcuBCMpe5mcgfKxdtHfnYWYOdR+B9HyGtseOCg2tYP2BV1byekQX
MpyvgR2NvencEzB1oQockqZcs6MtAabSMEhnDu5PujpqmYyLEY9xqe93bvhi
vjnpafhT4vlPa3fJ7b+t2oJhP0P6PJkcd1/GxOIMoOBIaUYaojkKRqTrZn2R
wnNeP/QK4N21MpDYEx+caIdzRcL1rSCBTLr0DJYbXcRv//SGuQ/NAgW6xm+k
TU9kQrER3AFZAf2Z+Px7PbTmbGHi2gzBzgusxus1SGc7J+QRdgrSi/DBLcpG
E+QAJqLKV4A3LjSvkpT+WF2Fap0KWzgigo7iiU7Igq/pI4i0xZFzvlThLUPt
AS8C+cwIuHKf+bxqSVSjFSEniummOsq+PUfVqNFy4dYp+23AJ8ZdZF5T52Lz
E89H/NQk1DBxCQEURSZEWCk1y9q8kdw49bKyDDivH+wecNTco21z4FIBr0Bp
+yy3K7C9cDhTvSZum7nwfno+kRquY8AH4LkFzgyUwLbxldnHswyna2imlSRF
BX0x98h84TmiTtl98D+6kXSkUa2sbvob12toP0A6hzbHp/I96jykAoR8tgdY
N1wVxs3Psk+mLqJkzfgSPhaREfjTXsPLWzYDJOk+pRXrgT0cfUOtjlrpO+Kq
m6V1Nze22nwHAcOZnz7vG0uAGisv64NEykmh8U9QLx9Mla+4p5Uzxh8x02uW
YjxOLFhFYXiBA+0pRrHcFkLHaxKpBf0zuV0Xy0jsZrOpa+Qjfz92dGCJiAVD
KkVkt1E1KazypwG0I3Mzkext6l1gGB74PuYJhv4aGHCxjHtbWKn9qit95Dq4
KRsSKRBQ6SWN7jL4b3xMHHefWuH+pBb/AE35twReKdqcZ2/HFfP40ZCxzEMZ
GMYo6M2XJmW9ofTLcyyRygPPaKk5/gXiDp5e5QdOkQ/stf7F0/lLWUoFUFdx
MaKNVRhid/u5Z1ij40jungBeDEgB6mcP02veu4grwRZzpxl2fhIaXpFHVW5R
cIiTh9Cl0ArmHmkQ/2iIgj2vtQHiMN8ztrfezbvSoCc4Zmx7WgWC01hsx3sK
Gw3BZtyal8rgwfopQFA78yZ09gkvuMXkiLrXjuFoiuVC0sRgGbCqd9DQAAFa
m4fwgv1AGpPQiQOMFmFHh6sf3ovAZk3z6QVxPnekH0/jNgV82MEMCatqRMcL
Kx4AbMGZwpo9UVl0YKtUjrde1Vjz28fiQ8v9x8iMBzo2KqsiTu3EsQ9URZSq
7ujQBnst09lqaexRGyEfCxPoRIMgGnVABAaMa/f44UkDFQsDXk2Gqanlkz6W
7CazKacwf4EfYBU8nTa8PRj8kNUIniYnrSWX+Z06yDW6evbNUgAjQOXswx6c
wTTCpAGR3NsZWgPf+alAKWZk0Sa6oN3cfIqG+deQJQectDyPzMc3wry53Ie5
wvx7BeQ6er1QVSf0hnE9dJ6m8TQ2ZZeGL9HJyQhnuP+mB+9kYepNv9riZ61x
em7uYiGHSMjyDHIeC+ehWgo+yxI0Pct7ERRMmLGSR8AmunW24538ZTcZ6bPM
zpu9AA7v5FYupa6FjVJm1QwXZO2gp66nWlIQBeQjWatSKOoj/8XWRqL7a9lL
jair6XXoqujdj5ZjnKPCyu1eUiL/YkcA2KFcUJ6S7iejdp35lYoWHIChA9ae
M41SuXC6Rv9QH7FdRUrbwxzRn+IjMM78k50/YshNv01MzYanL2xHCpPYS/EF
c3IZ/Zphlepqap8AOF3kWqdyuK7GCK3tWVoVkKFYKY4vufPyA7p6mhhK26eN
WCNL9+7opzPY0mBMsFteIFkswJk99x2tg9D8EG2E18Y6stskE9yqrHUgkkqm
zy8CnSM1/teGpEbK1RjOdrDwFFTa73Sy8BJLxURbRhqFv3qEh3KEdN4PyDCJ
QpLbBnhKeNSFN1bJtEO5q8Nv0HUI69P9WJrctBrX5EVLJGVa4pu3okB3aVfX
HJVG0YC86lVUhqZuNpuPGV0e3cbxVPW79T9oCBu2SG42Cx1SmCmB+GYq8GF0
VFkQifKGZsUGZ/XQQeGcr/JBQ3c4ZxQH8UuTH+y0+nQitYGRsL4B6SRZzRqw
xAT3zc+uCOF5W9gLq5PuvrootS1sV466dqJyAmgNQAX7ECcONDgovMx03Jbe
tcwBPrNHmVpbj7vno5vA+kA0e/maPx23Ng2mbLSTVDp9wm+m91m/trHPxspF
20wMhthytgJY4jep1MAijB0/zhKOgxhrU3uAl9sYSMIdL/jOwYt90oNoEWI7
9e1nEq5/bMHnMmRTBHrUTx2WSM2DfToRk+I2/D0KgKfo0WBlnmpZiOk7t2fr
oJXfZqCnlr/3+nONfpK3sCNGOa1BrD2hR3bTWfzfLGcsVSO4nuzeMD1iOZY7
FCxT3kIf880jKBwhg3N5N61omSsJlme9N4Lidvr1jioRB7lYtKhOO5dMVz1l
ndZ0AIU/9ls3fUE8nLA//MRxxgaz6jOufjUur1Io+UsjiG0BU71DReMYJYSM
bUm5o2xlLoOiSC6Xt+Z8FuNBbhlXFF1aNZ11cC1uMzInrx83kueqDJ3Fn5dF
bVch0F0b86VEr0MgKEBJWI3XLJJwImUlhXUMZlituHw8yMlWtf4S5qLBtJH6
eKOKzyHiakWM5tIeH808oBZDt3jChkeafLTDPnHBb7wEcEMOUQsdbInn4GNb
FJ2M3FlEpeaKbCDDS3+dxV72J2mo2eDmn2AsOpRHbfOxnNzZM7marQvTOEEo
8sITzDQehgxclT+WfE9JXpDEeFcsyhRilHAx2dxpmhuuqPjXbjRR20Mfwo1U
ymOwKhAdyRTHUMHGlwcRSMXCfylFtEOmuth5xil6ON7yv9wneJfWhK8vFKnS
rMJGZT/47w740kU46O9aCqOWNWCulmlKxV2N4e/qvswmjW3q6+TGSHn0/uuu
fKCvV+Qgf19S1A50PSKjXSN+bL5b4D7J2warrjMaWMv0Y/l57hw+ML0/FuDB
ayEvTqkWze73hMF879TGBBDcr8VVD6fzj2lTp2hQvAwTtH1qxyOy9tMw8BK5
N0JXiJoCvDg3sT4JlC+KPfV31AOqarKdjvZ74j4i3DfhlLbRaUSq16/x6+vV
9SpJ5hMJ6Mx+nmnSuv6v/2beQityThM7zw1orutQvGriYGu70XujK/HOEL6X
nb12agVQ0InGBjZhW+wbwKIgOKQA2CKgp3hIIUx1gQZqg6PaEUpYYzpSvDKD
rvQ75tgJPmXns2MUPXNoRYmnv7KmYpD9VcQelV8m9wbar0LqqNSC88gXrYEo
igiSuS1FBhrOti11aCetHynSVEmirEfZeMLpoeIVlk04k5Y13IMYeySWmkbG
QVXPTYbiOatRQv4BnqWU05c6KhKo2Cj3eBhxb50mBG3ELajx/zeDje33+Vc7
WKp0stvZiVq024ITs4BJeap7slL0/krtbvY9AvP2zgr76EalNtqTbVdjUNKn
BjjwOin2hCG4guqo9a3i80I9zhEHBn+FqvYYPlauW/vFjMtttbG4MgO7DvhH
BD/TRfKx3GXOeUscs1J7+YXjprGRJQtY+qfPJhQRHlHKroJIQiEJu6BgQPph
593nranqzfx7bVIEd0BSvtElb92Kf3qD0tx5Al1RX8FwxapIRxUl9qkCv5H7
vbjY2gUfhhkh1Uq/cPYGoPnRZUaT4Fq2hJhwEuKnCOoQrX7gKzLEyQj1Ru20
OkzfQlzVjbnIsZ1BwBeN6js+i+BM80mpKCGPL+e7Rh4RuGE85nzyPHotDSSg
B/5zq2Zkhjl0PntVU4fod+D9rqc+Yop4OxFMhPEPcKEeZCfFJjCltbt6TxUd
3yb9EItuxo9RzVuf4kJZjDKeqUPtW9w/cXD5WKE9bKp/zqPB6CyueFIJ4sh4
rvYujmP3EsJ/OYYRDeoq7zLHkkk39HOODmUS4tWYGyUnrIX5tW1u21fWLrHd
6LxQdsrNWzv5YqlCk3YkccUe70KFz2uWo2kWBYcYa6NsYvAm76sc39aKERgY
lnX3ka4CF2lz7wL0vQWr3qPWjblkJnumJlfd/pTPehN7is2zvMOlSyCGgme0
a3XCeJJD3OcDt8gS9s9vRVEoJYpMFTcszV0kTKc9VJD3AMdA6RlXyonqphS9
klaJj631W1E9Apf+K7auBa64RaPRAv2elVVe7MNSbmhIeIBbHNaPyQqNsLXl
dFVRGEq2V8QCAZmBM3UBl0GcjnQCCyh1G+kOxWQax9zQOOGGOEcOjQgndPbB
zJ1Du6+PXh0wp0CqfHh0orqIMlhyWkW3cyY9m2BoEEKqrIpYWN2idBWw0epV
foVGrWCHtZmRmHhPhOu/W6h2ZVjOMYeqAqCw5eIigBq1vKEVeBC9iHkQd7wP
XH7DuBw+7DdgcUqpqw50QG7Be2ffN0TkXGOX92vlAfB22IDQP7OnpRs0Shxv
DmgTmTwPMFCu9asVZQdG294LytHr3i+SWY+QSfBYVnOsEF+m5uTpM4g8MZTy
4qvzbuiq8nbxuyAaC5EybLWPCR70e/OmUyqWwQKA2Osgv790g5ldmMHt9Y1u
lJn2NsG61+8gAu9tHWODia63LtAV0RaUIubINIpaAE6OAFDZy5wmWtGrFrrY
UkASOiAvknj4LMNza47URCMf8PYrjZv4D7dLfKRuWQp6SSb/e2PcDcSqUHOY
e7U9K/qqvHGI/eLik+0PGYwq1PtA4oFIsqwhy/7nRiitECNLXLc2C6BrjUEE
942tfRPYmPzXNmlfqbhRpuu89WiKk9Gi3t1ptW/gUnx74OGLlhb+CfCdvbIe
GlQL7RW4Ng19zXHw20b5R1a4ahvdOYwmmpffes3BjcbeB+Pct/CezQyCy3MV
Yy0DB2JcTOtDXpxokFvwadP22vmB0wrlD7LgGurU8CHYJmGpbQVJH/H6MVTm
FCdznwiP2K//fT4FPV2/RGuVdrJPE6dHozn6n2p+Xwj7/tCEVwLpYrDyMCTG
1OHhVGxMne9OzKvStu0bovCy/ntbTR0AFpyyRGZPmWRdJ6WMOBhlGhroBEwG
Y7+MXL15fBzsdHqqSGMANCXWLe3twb/pjRpvmz1f0l7wKXmExjRn7srENbNn
yxyxeYhWwbAGvRRmZzzgZlyNhZoge0XMz0QhdausR1YNKujCLnMgScKdfjh1
MBVkudyZGyOieYIxEkRQQfpacldTYAdgvSE99HBSr/OSrrjCRD5dBKgaBGkp
dzUzliPapiidcuPyaZ5Gn0x31v+mWw2+9z7hf2pcByRgerCLuJ6A3kk3zzpr
xqp5xbNYrNJfVsBgzGCP9XhAggTFKXt/kUfEDTGAJuLQCPJu/k7ggBlAbKyL
KVdjezPkmvawvexzehAfRWpGQ0ZtvxuX45b6ErLpZtNdltvAl+Urf1kLbQje
zgMsEn2hXvb84S72gV5X06Nus2MYqtBhyy7MaukQx7kbyclBgtPUa6AFqBIo
N/sa4MjsEQX1vNX8thIVnU4UP6GknefEtCGYcYPXr5xQdRObLqY/0HDDRbG0
WVzPOprpt/luyzjT7MWmu+yf4iAoxq1bSBKVmRwK0UUlydIcQqzZA/oArOPi
0opQHSRZbAZwtEpaoBqEmXb3k4taljnqBX7KWBOoFInon6OGCl7Qlc8ylkxK
YGKxPckx4CdRUYmn1hDTETIpcG0JwSRCJ/ke1wnTLZwYIjQpLJPM+mQcIAXY
Q0WMkmJOncOxhN0Xa7S9ZcC0JW64QLXDIb3IAIAkr3Wisy6SDQ0JdGYZDHF8
IHsYR9ZCECRIWizogmDjm0Eldo9qUiIB0QyCv4YpQSs7fa6nIyEGFuym5wvf
5jrQjGD6A7YezcmCXdcuzQYgxBsj3XE2iab4SwyANrLw1v4jw0WlAik3nTT8
I+FiqLC37GSZb4bi2qzxxb9MdWkvzwJXLgojX2yTlMQ61cXpL6yiVpnDnhTP
SJfOLQcAfnmJKzcRKKJ9uSxTlQ2KD3K/9wnTlhA6leq8o1hmFeEKW5LoEJco
JHj7mtQ3F/trRslzE2ws6t49K6shgJK6b5E7x+pLvzbWAvBiPkEE1whtalqb
kFrOJ/Zq0aNCXsBATOv2/B7G+CCGZyfrvXdR/gf8VFjdzWrGbRFvqXePo+hr
gnDb70utPgmlbbRH1xj5YMmZCLK7X4C4qNCSPvBtN1IPnhJDrTyNoTVPOX50
TPp2tg97jIwRX3UUqlMaItjTBMfx+i65mkbGoyqSQADnsxR40CmDPyKz283p
Q1wBpWgNBfMvWp42loAzvmd505t3NF5AmG2paFZD0/GO0+qw2babfH3STQq7
ZH6FD8RZ35/YfwyAcYkC9lsQNwu1a43Th4EXZ5GY6czcNwPRhASUUhhrsRyF
xVCugPUjq9ejTZdlethVD8N90O5fV5Uqb/az4tzXph5a3w/ruLp0s0IZ79r4
6aXp06hmKUbLqw1Pq8DN4+eDkD9qFDJ+MEcaB9qY/WaUApSGVTvdBp1IaofH
e26qvc4iSkq0Zuxjtync7h5Jyt7pjkyaQvRVmGsOArTeMtNmbfFdgH7AICJo
EbFFn7CTBsXa3XFDaaBosWehAk/Km0uaTVasXJ2h+gI3i5Shkd+/lJKqrAm7
FjMkmjUEeBHiH7wj2ZAANC3H2e68zW9ULjppTQ+aPZwpSTMih+SbTOgTxXLI
NnYc0QNpPGB9Zhcor9cu9C25ZhiwibGcXPG2HNyqcjf7J5XgLIeQNkVrkAaf
PR7n3oel6URhJQBsXOm1IVEv8pp09f4HgxaPUyZF0nPzdE2d7fxc5Npp+XPw
DBMVdDMD21rGtAnsu4zZu2tnE/PJPy3J+hFp6ZAfzKhC+dKyKsYw9NtNlJOz
rsPNBn7N+CpaqACLxYEihDhw1cUxr0rn6DmoU8cEkM0zennELN+T2P2Fd7KY
VeXEOkym/Wt7C8XgX5B6N7HXQ6LyJPdRfF0jqQxoAia6rZfGSPznZmRwjQ6/
5haPwq9P4LGtm2VqL4X1jHYINxxXqNpnfttMqcmFs96GCXyMAebJCcvgni4d
whx+VmOHilkeBFVv2dZ/de3PAMIHUlpD7/iXAFRqgviXu2dwCeGNrIGXsX7W
Kqkr8lJQDs/eKB2MS2lMu+3e03stgx20AjJIpHLeLJzOBLGVYZEwXiK5LcGO
/PWKRFCDwRDYt5E81T4io6+ElL0f//Ogj4Bi8G7uVJOnCFpx0E6+7sBnyqq0
az6YSd80WFXzYRF4HSa17gSUs9FRdBWhgAA5kOLCRWf/R+yPsjKhsKUxalkF
/GDyRmB3Sk/FJswCkjwMK9ycxlzMgbTioKnV4PmB5DbDnfvxCHVkNjkxN9jQ
LtBuGeifb4pMT9GN0p08vSL+bXjKreWaByX4RmTALiyr0N19MPmUxV6EfURi
PZXcka3V6j2iCzkeVyL/6Aj+ZFWIYzYeyJ8sskquXYXiD9hwpDIpOzaiAD7p
j5Va29i//GpB7iiJnOpaWh72Znh8JpxQ1cldts+HbiOuNQ7dUEtW+NYv+rCG
0FUW04IpuSMpJLsRZLEo9anmBYiKMhrCwnEZqRyteH5I9uC+gf2G2O/RFBPu
uBBUTXTBwZ4WtcmvN5o8tINnITd+2kYP+1JNZyfTNL4aI05+R0GO81lrR6Gg
YpPlyXIzbHIVI24DGk57q9NX52ySuvDqfBJeiE01ZYMiSB0r+wlj8aC9Y2MK
RHMjHMGCx6LexTjaFEW3EmtliDmoNUVQpcKmhPEjoTNU6ZpBaS2ukggb6qMh
5p6bSYU4EGk1vCH210Ow20RTZ+brLEY9znMyIk8JabiPG4RDxNaSL93Avi7D
YLvcySeL/XpKpqYDURv/pG4rxT/00q7SYweXVybtm1Lbr3XXnPSplQk712p4
NlQqWgiGuVHkcd6PFSuNzGkAojYX8JW21wa5dcuTAwYTqK8RiXGZZ5xOY3CV
oDhFTnl95g2rGaqcslmKx8jpCqOv70kvBkEoFL3MKLjCRvWwqQGpmafpjxyL
tL+4eSuh+zkMvO14BqPb2vw8HYX7XaZ5S2SqPCjSW+xGioqWw5E4hEyU3oXO
ixSVqWio6Q1bVXPRrs8vgWWxhFsBuOhoaG+YXLH3jy4vZJb7vEx/j1nAFOed
ycBZjyhjAYjDIrgtBuCN7f7sv4vHr5mK3Zpio9mcFI43LEcHk75DgkfDI5pJ
HGOkPMM9Um4mTZVh5QHzKZwL3kC4ylJwOy80hXAL1oe07naOuRJW1m7oQtqn
Y6oPyiOvvUZHJz6MN7b4JfDK1NKCVyGyDoppZHCObWNorNhZR2qHp17kj46B
8iN2wbPsSPwK8CpdfqHH7wgESA+5BZ7w+FN1erBTLDBpN2CUmrlrcmo+zQbJ
tbQ2cMy/uyuSigC64ERwupdseosPgSsuk5QjVV7rHHofdNtjCkqstllnUVej
tyBmn+VpLz1J9JBAd3/gidZ+K/yy+OjzQInBRS4Ek9KcwtEbVLUNqTpZvmjo
M5n8pBsWEzUd24zqhEI94hkgocKvWzZyZ2PsBJDTUuU/Hnp+8dd09roKRC1z
QFaf9apJpPJYGdD9P6Uq0OMJCqG0qDD9V3dV1em0pZZe0qoymXVkKF00jSmz
to/o4urTYavGDc6LT3DCktj1CL+vQIDrScf2SRYJlncSxzVZbMfYBSq2NPAs
Zj5nsdvM4GF+30Dab8pJIXomhW9JacGGedHyu24ABqXXsVxxPhchtGGwErgA
TOSOi7iRZXHfCQ9p04VzFZjQH57hCWU9pkihVyaK9EMQwu5gJkAol2O+8Sfy
8S5Djua3sxpwVa7P6XMlQGSXK9pYjRvxP6zkkt3b5J0YOIAdFoM5ExAhgnuM
vDus49omHcJ90B65WHV+WKT+lOFq459kfdXqi8mD1mrzo+3eDQ3bBDKJsWOd
mNg/FcNd44qStTK23OgU8eMMEz7pwLDbWkvroOzX2JyzNxg+8zvpsoNxuxSS
T784YIWBmW5Qo00HW8XbU+wGq9WgtEO4m/Axn/l/EFziWK2xi7Zq6z/7o7HF
3IP1j1F6Zv8UK3y4SL+9eZKoMD4KBVlck6VoifPPd5byFeQ1eS/b8B2u7y4Z
lLQvdAa4Acx8cutMUrk+J/191qYSqQXg8XAMKN1+PmNBot2ZEOIYkSnV9Vo4
42D8HQB+7YSmVOmA9zRPbkwM1yU2Hy+9XFVn/werC6/r8lfY9FzEj+8d6Wnn
h+yi8Uw6wDOnUeA5YpY92fsDsQB3JElVDiFTBWKpSqm71gc/BQOtSbYyMcyS
0KFiswwOZ1vy2a/2sN30r6e/OgczAepgn0fklvi+RZf1i1fXdIKnJZt4UNRU
FOoVTC4O3dldYKhO5uxzZQsynzjDBI4M+tafnzycskv3BTac3oPpxYGE3U39
XGSCkk7Vf8DDBLts/HFtaU0UVSC8F0mWuyhqE458WZgME1zHtRd6ncOwokKt
OIzC5uX0sGSGDAJDc1kKcx7QIr2r3DXRnNYvVJM58rAKtSsMln5ktYig5Smo
yH7DA9O/LTno/SnaKEzRMQiFYxktDz6hCkh3M5zYI0e6c6eUfqiMW1tfmLo5
+e5GyxgP0w1I/Fggbl03vZj9f8E8l/9Crcax12Hq5F+DIqNV5eeCe6sxlLrG
ck+xgHwfMp2D/hrtGLrklZlu/xApcv4U8sLjcp+jzeKc6QGQH8EC2weWdmJl
hdD7uhqgsXoFBkuXJbRN/hoOeq8hMGsTI3BZjy9GHLDjxXOmgBU6+4AgB6sG
6+YpMlXCsjBgoaxSn94oE1XSUIhLW00DADIoRbm7bmtTT7FtTEG/2huyjZhq
Qsphv87yGbcE5GqkOkbT47Xy0Xm2UTskk1j2T2HoL3OYdcpSXKrQCSDbiUZP
Rgt07BgPBbRxWQvu+F/UJKun+Xs//fGotESbymeib2i/+fQI2pT1pCfISLYx
qCXzkrt5kbbGfMpI50gq+b3neIvYqUeTRLd+veyreO6UA8ffsZdXD8ck/ypl
w6aoSU574qrQWh922X6uTYkwV3Ndaac9nzslrJWWHXdRb/jkaKpdKqEcqpz6
jBfxVYTHEuQh3uylWgttIJNiyYQ0+6D3Vf7P+KK7SAmaR8ODtS4WKqqpZLPR
RJUf4BlwXr6b4iZYpOzWRzuyPqbBBJWeBA1MvNXPp8o6GnNOuGQ2iDr+jHla
5xiOCc+hu8bElV7L/aF5zE7M+DSvFajFXQuMh55ze57L0EEOfeRximVXemuq
CBAMc31ch2DmoCXC9B4VdIX+82wG7oC9EBIfP+CaNZR7lrnlmvdFT45H1vMH
fjy+2zHxQoIdEfs+Zy/HymTKYQTbF+Lp9Hp03jVZRHE5oz7DTx8KdGkvcbmE
4NT/bRjh1yDV1AQ3ddFXEjmp4qBEh5baGenBwdZUaFAgiD86aHO3eJw2fx5f
CFlHc4MOGh7XVRMvqkLDRXpIOriQIrHHuv+xAxdDQ/nBsy72SQGVelmemOSy
Kxwrea725N9/Qpc9SKjm3RBwhFvnh4TSjXsQaI78wVhynQtYqW/zaD+BmMYF
Xe9oCuU2eKGqDnCgD5ylYo7qO78si0tCT/Px4zH1TMzIR+0MyNB8AGysRQPI
k6Xta2LwkMvfslS7UsVJ558+od2UNsRfgbkC3OyWb1E+Pr98SZ9c9qgFbEQW
QWiofSCdZ7A1/9dHx0zXkgTn8Bq4rf9VYQ2N4ABWyFeyA0IcCUqmShJmLAAs
tzVYdmM0iOs8nMOj9ftb+g+qUy2BTYP9ZQQYrKhjcZKU+0NTJs2SBsBaBVXE
g6MolWuiL80NpO/dUWVlHmpJGGpDHfqPsCJR9EnjxwclE5UcL3Xb9dZ7426+
0sp8jAoc4PlnPusU8+Ey1cj6HAXNxFhEI/7H/g0mTMWYPnqwEznqU0+5Mcsd
YbPzam1ePFH6cIEBfJzm6XtFdrujrvxyEDYgojp5Sy1orKdrfLVE8YN3Phb3
P1emz+cYjyP2gFM7snUfcDD9yEMoqjEBKV9TVsk62SllPahRUDtTkTGl4jjU
mMViZxgV0s2KYwIY86sgN+Rz2VMWK89BSw1ySO5qxKzQKXxKQLLJCjuGhvFt
Aoslm8o0CaIjXz3tCRmAbuqSsuCREtJcKQQBIDrpdf1bRL0nJUejhSsBvUfp
UkdyEwmOHQq6SWEhrAOmy6THQn3r7/TCJJ+oOUErnrmzzGZ7Re1F867K/H/J
AxgSaqY+OwL4UbNfNwQLZj7PMm1ZTxI8frwpLJ8oS9BI2bQx4kL0GidhXSqQ
GkWWjtqujTp9eFhv3qGawKOQ1uwNp2/xlVe2KMBC9gWDbGGqHvAzKTmfaMBv
WnTcV1u8K+UV0uyaaRctc2/exgt9qGdUdogHs4KtWw255CvxiYNdU8AR/ANM
EOUOPK0eXGnTdKkILJlmZRgRE1pVV6VX8NVjo6PrcgRfUIghl8SKVllgkjgL
vdEXjUyvgDsUSUy4sxA89ijkxHeH4F1EEUfKabhURbJSUMXq1VTdturzbVmL
2lTnLBNSuDyTwkT6HxtUQjMkG7CkwvnFT1OP1JeVbevDqWy/WqZKyfJh7yNc
/L1ANfgOY2OzCxvty3MFWX09kcQMIsa+h9De7r15ZtS39ssd9HKoRwc1aNjP
ZijtDJojFBcrvCG2nUkpz8oovO8Vbj1dxl6hcZITubeqSUS6EZhfj9eVA5o7
r/OxgC4AcMF3UGCLrGlDTnMGJLb2M8nxOIlXpY6Ki7mCgVJjj1h51s9YA7Xn
S71CRV97Fvt2iPSTk1yxdCc0k++IVxMMk9qN37HKk4HfeKKF2+MsWYTRhAzO
+uWvt9xtPqM2Yulemxahd0lmcOAv038xe32yoRIrTp3o8jgiCOK+x5mvPycO
0hbSrCPpYQ5o64ojidd7FtvymikbQhKpaA8TEqKTjDPj5iLe18MHA9iuuHJa
4NnxkNMklnH/oAZgUwfyJf2zWijYSXGw1obWz9SWXrsXWN+6r37A4bHoAh59
cz8Me7JY0nSpS/dEblqMndpwQwalbsn1FKOqQ2ASwDYWjb5rr1HoAiYJwATb
RYwmsOi1P2+jmc3Z3jdi02q/YSN4K3dEcvNQ+jK/s1SoguNGMSfTgHsRTVtc
qE3vjIclSh/I20rvY04Xju5JbiOjPd7RWSWOT0WmwW8aDww+DqSXaUwm6gJI
bYaUvn33TXtLNCYVF1w4UasU/jwRopWihOvnD52vWZdj3/8vLzzpm2z7taCe
bc8UVTacW1j46UtFUNHz3KvMABwblHfy+OniUerk0kyQAbX5m0nVQE9jrNww
TWFVo7LHDdpcNKibulik2u5lD+ClgY2g+2QQ5AMhbpEM14jVbRJP89VgPDhW
G26TMD5rxf2nJy4Zz7HJ6V+qXyvHO53L5MIC9UDls5u+ohN5utZxPyFilDEI
IdssYRWkmTj7foFKqGJV2WBOKOmzulPVc207qAEpVZLrl4amgjlwx1H8eEi9
9QZkBx7cXKBXkNHl16NRBx21rpUP/L7TG2AGsAvm8HkBu/0YOIZIHDx4GomG
kgft4oSV6MAx0IFwCsS3ksJd/44CzHXU+CRFf+kfNAlmYwxdhlAvZQm0jiDu
bfkKHdpapz7AjIVpC/F5HzyzErHfeOurO6olCqE8RQqYKscmeO2lMsS1pOIy
FVcbuxj5Nj/IfWLKgzOFQLRcxlEnJxMrPRhGvNgi0jxAXEz5O28GaZ5J31k/
j8K1T9Yx78IzlYeI4Fgj6JV0PQUxeHaihnr2Udm2ZywI3ewc3dIxT3pyZlKL
XdbQ0cyWX4nr8qUY+jK3V5a8BbN2VOmcrPFdZ20/aNmilwi2F8nBg3dferfh
fKVWtSLGUH5Q11nZKVFWPxgfbHHSP2VnEiruGMcI76dJ9ovIDkz3qQ8aHxOQ
kyVSNa/2B4igHTfctw5YWfbHEU9gu2IXNHU6WW8ppbmpfhZ+zKEHbZB7aYPI
jGuoK7Z3MAl+TyTnNz6NrUElFRxGtbJN8zfRn+mCAfh3baYwH28OAd4in3yX
a6pZFJkUegPUbrSkvwUc1ilVSSTJekWHqQoEVhgg9rLALr5jMnZeUfOCMcpc
V/CYSx7KgDo4Da2P6AFZUhzohGx44BDnt5ZPdjVzA41cLUzQ4WAv8pUsMnjl
Msu9vxDmEjwFPOtln+4E5ERt7xrXsxJnogTu61jd6GwAIzVR+RDdFSwN/37t
cx2qerbT/CVgS4ENyWgi54eWC5cUGhobvf92HBzPKYkmuqP3qVtYZt9RaJlN
Q8fA9grj5Q3sdtxsQGYtWPRmZ2+rlnaAiufF7swfD7/8+uNDWwzzxSt9/+/N
w5hbcNE1ZBNiYeQpFb9WxSRQ2ne/xlE9nUdHjXl499MdS/Kd36dJQxAkjQ3N
tA1t9tapG6PKPVBMPHu4++Owg8RCQk+Itvp+jfC/J2Une63p66nlHzhjE2P7
0Cp/baxk9nriYIWu8qR5S7UVQGp6IAngQ/tXfFXfYEPNx8Fb/JdDMOIiWEA8
5KYek/GTc6cw46YF1uq1k0Fp+JlCxltwtEksteBIqezF2brn84LlCDOquczt
YJ3kPr5P+WWJEq5jLk/Gxrf8uQtOER46IP72vx7/FvZR0/aq0NKpv42Ik06L
BwgEbio/33hQYpL22pCUkg+8Yu53BVpRBnLjcOWk6vM8QNdjltLNYIuKEKNY
+NXvKhiiDgOcZ+1OV+3hMdk7W45JW12M64sCRiipKQLnS7aF6RcTYTZrYxU6
LAjMi2DOrPcP8NaxsHyOSRfdhHRrHA6n3JLSrkzszDlrOqT7I8JTOEIkXDlO
tBx0GAPgHv+pfaRf5h+ASR/HvHWHOV6JRWovr0KaJNfLdyqLvy0ke00ldh7a
pdaoMpTQvkW6J7pOh3YGfga4ib+KNQM7kaKsSscTUfIsoDAtMUa6nVwC5RUB
8iaq1+on1TpvwPQlQ/RN8VyZxsJelPLRnrqPfYlhVa+/BJy71s6U525Qeu2z
fqoJD5oSIpiG55cEnMEWX35PI/BhxOTKKPfpk6G95NRHQ0I/W/WM9kvOE8Wp
+2max5bwLRCbxl7whylMkMMUlCMV3HJjM9O/Zwf8mmkv2IEjmFGuKKb4d+tu
hXRJ20yPhMUes/sdCjhXIDuacwlkn2oZK8yr/I3BjMEnQjEoQU0LMon3q3HM
gMnNI13C4tsb95RtVDNATubtJb64ZhJVnSnJlvbHAS7xMQcW74mVtBFMSE8E
S7VrRiygyKObLoGr9wzaKgLIsOVRDsteh4FkgA/rFdqirjU4MIIOH2p10/gp
vh4PmWr5Sxcz9pWuUb96tykbcnXrCmGxaijhSxULjJHgUOmR26C5HPyMv1XZ
iCX8ff0B8mOmjPQYCbvI/53aoe7m6exxNUISX5rD4YdzWTBYbzR61Ea+Fe1m
QwUFhs1AEmjDfVAvPVQa/wWqt47xaBTqFmEZqpYydjpxhMzbcJNoa7pPN75m
bvKbJjKnucsHJKAw6gnuLaYP6lvilchWXsdQhx4DA5GO/rt5wFU6luKiPdOo
yJ3Ph6eNKYeIcnqWDswLJ/PS02Tltvow0ktIAhqeyrmOnzGDWAJvi5ko9ebO
1Sx/K4bYUEZAVUIH5xXyfzppMaYFiD+jfakGaZ3D9W8NWavtEFhsARWPedc9
oUfScT9QJLT/xqxsrLpkTMPAbi0EB8GNL9Tgic6PWAevprh7RnYod4uepC3G
ScPMwCHogxQPczEnMEWq/Ku7JJ9uhbioqjJcUIu3RDzAABxBqtKJLj+J+Ws5
8Q8acDeCvkdexWnOQgFp25F6aaS5ybkRMEZdwgAtlHJiPBvu4nCBzpaadkEK
3YViDmi8x5TnarOb4p1/XIScDiImP7hj0SiCgKRIo/xxzH9w3rdt/Pan4zMZ
ViQRSzBBQKsAEzBmDZZx54zc9eI9ebq7NEaHWT+EDTlsKbdzbmUIhNqGXTAp
e2YgkIxsXLNiRIevN7kUqIu58q4JTvpK4a9KCz0aGbpVw6hEeSDwxesvoO/f
ueJZyUgbfnSmIzjhultLQhuEmGxQMqO8vMdBiiWKVNoWZg8AV2epIrGFkwjf
J9tqfxygOpb3Sgd24B85vrzaovwkrrq5w560sl1XUmvIddNxp9p5V9bDmA9P
Vu/k3O+BnxD+ZHVZxU0G1kIQ5xxf06minGpryIjnzBYgN2da5GWodAjFeT7a
6/mybs/RiItAP6dnrNbiSYKxTHXb2X3ESEa/cQn3rmKTELUGKb7d6YUeuYap
GDxuS3Me9QkOOfGOGR7qp7TWoJEmnxpHozDNjJwowVUEYU0As0DNbIbF1MBt
aneA3NYgOLV6XdK+fxjy9/Pgsh8VGxcl2+K6kbZWnE3PrOKuESVoo6cuD89e
fjutGLFrMWdTkV/SaLzQYgwIvar+PufctEzitAMazJaGp0OihPKraFGKWCs0
KBoLrJ2rOqPh+8P9Y0UEWhjF5/PLzQoxHyUjl6KMZs+mo9rIwQMBEw33ByHm
POCrd3KBPEO0DVZ+a5L1KjfJ/OyTgDYe+MzgA8kIyzDNWDWcJadMufmddAbn
Y2fse6nsmBkry0AOe5oOfKJlRb92ChhXbV3PTsiUmZzpg2fwLSXndP63xR8v
NRoKSJ6GKVQWvHP3L1H/hOZQJcI+aadSKkPPbcAvQ1hwiY7tIhp0bNtFaTV8
oHnRnblc3sy/rLdRgjHq2umz4img5GPKPojdWzSIrfLXYrf2TH9u2HQVzUAG
9xEGsg8VYc7qRc5daCvn8GmwtVp2+PkfX6EASAW0DtQaMrRiKsaQgYiXOsyr
3WTa9NFgnyqGr0wEwlW8sl+qCZHggV/YqZSRhx9Bfa9ZsuzTrBvrvxFOrcYU
I+ERcFLLtIq4j0/VoEq7JV8AgJo6pTLSXj7AYGRdyJK0MG+VVZbnwLsG+RuJ
x/PnfGqLzU+7yGmgMTim6S3HB7yZReQWr8W/4Yyz9bjSBc41val1YDmvgG1a
bfQMuZJntC3PkAfNI0UqeEyGsBN4Kber7CXcqK/lJFhSpcU4EbKqL6njRzLJ
zCSBovVyZJCmCSacOms1XEnlchZp9jNb1GoKavpOk43A7lXZOtuPqoF5oyL/
FFKeWPSiJ5UH/Xu9/vqz5fo+sP5UiwjetRXPmTwgxOSOkLY3n6ubQfyVpKRI
QyG4XFABc+hTVBwsxEVcurZO/BAvtOgqbm8b6w2eSqLN1B21LGeiMVj4a5bu
2mq3hPn/0lPmJb45DGcnc/6SGLVywMA0yWoqyamg6wAvbNO59/cKwsrX5WQg
D/gc1Q2EgDavqLIXR8PVGuypKsNnRvXoVUPjAaOToHz92FbSwJrqgQWFUHe+
5o1eYD2kATWcj/CrnA2peGGILAwLy++PDnY5v8AaDVXHjShJkyZT7tN4viIT
inkGxPu249lZzFdkYU6xso7TrbCRBmZmmEQDaIGWtoRO56qpQ4jYPHVYaWJF
rTmD2ERgTLX/aBRW/H4sMIN4XPe2Jge1JoQ9zS6gHQCKd0Oh9Zdy7VWwEDi3
4G4+9rCupqPrszN+7DiS9+foT3VDuQBcZtbwCjtUpiL9pGWt47LHJ381A8GP
Juxc3cJbLgSfhjYJRBzLNxcc1y6vAZ2DB5RuSJ9EnPUnfRvyiXr1B3NKqVXD
hTIljf/Hvk4acWHgJMLbYeTOdJaKI6ZxIm8O4qLtaqSyv1goncMHVfmOukB8
RtoHujcnz4IPagVDLC277Bqx5CGdMAeloqSdSiem/Yij3jljS89zwMOwZruG
5H/9kt4dqMpy0ZLpKtLRdWh045yrW6TjsilVD+KzlhikGoqxwVpQk0WgCnTb
v/+76DpqZpImrdSWbr+UTrQRz92ioDI7Xm5qHSpw5Uia6zOW5dOhEkzPKkOS
8IVqS5laPSMb5TQE4LeKOg9FCtbeVZKk9ltLss7ZtUCzUs3sXmZiV+eYFMHl
EzxXOrV5FKI/FwHE+RSSdjT3f4nmbIBCGW8srZ5z4k6dntF3DLUqdVdmYsxY
GGvcAqc+jwKufy23Ygrh5xpODrNB8oMcQF8qh5cHvqICuNVH4yaPXCnCMf5a
C4xVFH94vUL0Jj+VWbcRqwDtQ8kdK8+AIDW6fWy+etvFa1IIvdlqftGgNGIc
Huf1zy0G9YH/KaIyD+J5XcAu6wokuD8nB5WSb6zsuKrYm/yS2LkT7iLseMvx
LwadKjqdk/S/GDmAsCp+wTL/h48pDsFbhi4HB7qLnIFGSTYR808JAHPHgoQv
fDk3KEjjhY66EHk1u/h7y3p3x7LdXPaKPbQ/spNLrv/aSvbulXGTZeLWzrfY
T3H5XuocSS4ItfB82h6cj6KthuBUTQMqKkvF9Yzcww3YjNqR+l2SiWFFjxvd
lwBBU7Mx0jd1KiTe3l0NB3VqMcQv8jUCZPC8wL6PMzH7E6TMPQLx/HunjK2A
coXKmnA99z9IrWO1fQcuCMGEyvF987r+a1hX45HPVDkZ4Sr8CCCgl7F+stOb
okxmcpG5g1Bdvzbq88SnJBJRwu5+w3Dm89B8/BjokOWuHDmwMATY0+2NHT3u
ckyNmxa76T0C/Dyar15AaMAdeA09dJDl2OtlU/nrvD4gkM687IjbnK7B805E
hgzUZe4YqCX6aUguj4lapubNQut8/zlKguIK2QDlA11KKjKTuCqH7M0XtGLV
PavdWEpKr5VncOx7AiF8pVi7/htpE6XV1TD3m2VI6fYRDZHQaQBvq9093Gl/
w2yPpBvrKD3ialGfG6SImngxuUT838ptcxx22p7fWP+s8dB8B4k9aJVUHTyx
xHHZ+/2hRVMZTN7WAERD9ublTikKMymblgduy21y6Tuv0tJ18CbOzYWz5KSb
i9FpS8nQOCIk/TJftw/1FBPGZlgS5AGSTfnZuSe0aGSVr3ZLtY+PjJ5HL3um
/Ec/qt68jsYknAf6CztsRsLop8t3Bk2sISupP4XVWsPpLGrhIvsljO7r9ffT
cc+McyRtqrh5deBxRhaS83Lf38nNSyH0BtBF9BilPBLZOh+j1J8CHL8AYv6v
TRZ/24c4sTZdiCiXs1H32q+lpo+QuCgNCl9DFRag0J4bjCzXS0eA6h/JmIW1
6O2fI4QlvDaTDfUfmykkf+NBBHEkixSqTcI7AhkPr+JGNS7IN0P3rE4WkjV7
K/VNGA7I4z85ssKx8WbSPpWSkVhs07lUfAKhNID598SaC6arG4yOlxkHdJU9
3h6OQU3B9OVoj9Ef9xHGAttWj9cMFtvjVdtFjVRENql9LDGzaHgcEDeCjbWD
Xmm3EkNrMs8NLDrg5HnutOZj//45+kXhCJT7FCfZfw2om3+AqNbi/PGWFS3a
umlrDEWNf6jfIxsGgmjYhySLiSMwD5VkW9IpEUTD9LQ5goO4n7NdNtVgK+ux
3uoVIVToIFOlyPYMus+4Mg08BrCBB42jbARQl1BF+QLKA/+4hfRqtpspP1TE
+WB2hMc5ogZO6Ik/Xq9nFsYMa3RTJb2PV1aMjdSqsbS56tbBSSnQn9wlstJe
fcrFf+Wp0ZDwe/CzhvMXsAMHpX3yDNLnt+aClcKxcJAbmndrV2Kzi+NJAg5a
EqFcczv+dVqa6v5QCT7YFKfgZL1vvL1k/tWNEKt0p+wYSTkjX8Urhp4d/f/x
CDBCpsJTX2DaQWTfyXArNPq45SP7TZCjRp0Pc4UvKeAS9Bvwg79QXMwQRaOI
ZwA+NLEtABANp590JCo9qS9B5r3iT5BIB4Q+o9ITfS6FDZgo2VdXo8MK/tsA
CUDMxbcpJs2MrYeayFEjhXcKIreay/fOL18DRlugOhXKWqjStVphdj6QTPEC
8udE/WGYQYVnhK+B3smWsBHg26DxHAKMjXOtL0W8OzJElXIXqMddn/EweKz/
02k9GQB6CWvJoGn69vMGjJ0o3q8OOmwOhB9flki8rR3UudhvA4xRaBREb9ff
uWwMbu+zUsqOuqbfqnv9wMF/ZV8bieFZ8wokGl8rh/qrzEtRHW5HroA385RB
WQAjAatFsEvm8HWCf8MCW4G7OMvbK/+Oyz+lth3dEWeyZLlRgM3xT0rzFl1q
QgCiu+9aP9nrabD8e9yymeolEp/tXuVpEpPXr6Uhm9lLFqr5nlRTG1R/L9LN
g/gtJBGGtJ1+5ZqzVdML1h4G6EAN7lsqZQmGh5p0YccWsKa5fRvwBKPaqiwQ
EKCdrrgW0kuMu5pbZgiFnYrsMEpfz0XrHXrMOQzDDuF/tRoya0B8xJSLqc3a
9xXRGASoCsxWkv28wsaKfKdxZ6C1HGCzWc53IjgkpHS9pc5QFDOAGvJlC1om
YZr8s38zbQ2OHDGoaWBcROXTWTLx6827AmORwZCBIr+6tLekeEwWenI+Kp40
kN2EGK27+mMfISra6a9P1rSnduJG+kJsOLaJRvep5ta7v6doE4a6PO16rC8B
sVmTjulnYuarjXxC8k1WR1vnmR2yVkxxqx98cqx81CK9vSZX4IR29XDZTrpO
VTQhGduYy04C0c7cu/surckQJP3ESFqkRgKsDXdH5pFz/i1eL90zEF0F4e8I
hKGrdYItf8pgpi4XaN7Ber18gKcMjT6Ngx83B9MckuArjwhWamIuEpkMtYsl
BVNqATUIhOpV7PglKzGvCHwsEXgFCMF+LERwj9J9AgDxHqZoMTD6NfHCJyro
HNZcc5H6SyigMLU1GM+Ex0v65gMw6GGyeQzC8xe6ZM44GeQsEgAGdM793Bgw
r2VNtlIUoFKRJmJc+81trcdni5u2m+gG1/vDQGCdNZN+cRmlqaydc2H/Cnkm
nJhKO0v1iM1jQfXZejK+RL27tzyBNFqHwGSBV6FKOeBM6vAg8ZhVv45MGXnM
Hga+i9ezkhxoohWzJPdnB4KEHQQwO07PM9afnRlAuYJQNoTj0AMQ6xr9/TMj
h6WCr+Oomx+uBPr1FPsLkwoetlXkEok4AMEgRDPwbJUzeCTTIP7xSUP8aqRV
2PBTIrWNBLHrCGNp9hrigk8gzwLlyVXYY7+Rr+AAP9DLLyyrQ3DsweqUfMG3
k0B4sPP51/e61PWvdi7el/u9Y1oFIpXN8vn8sGTqXahcXMypp57MSW+4siXD
Ze9MUpqoIU0rATSCYMFZgnRLLea+AQdgGp/emlItCb4R4FJnUqOhgbhIrzgO
sS6L25EXXRtl0Ee4Slw0MAoQMYcbJ/UVO5Vg55i1u7cHWM89Fv1e/voBZu8U
czqYq7Fus/LYYES7r1n6uXNfDJmty7wogSmMq6y42DB/1UzUe3wHIVTXl+1B
+rfVuVPb0NUKq3bgA77r7D5HQ1hE8zoJ8UqPKD5K8pz6bNGIchgf7pUw1K2u
7C0wKney4nlcOdsGzN1T/Cy1HCdqfCfUKQsgXNBHyM7u5zApwhVs5fQCQ8y3
qIuD2QRiRWQJTlNgYHmeOVrdNjToO8Oy+bLu7cUd/EsYoi9Izua0TALfhjuj
/PQfp1zwdAtxOLVW9mi0lPrAMppvX0aTrYCid7bE2Mu6vDiC+ms2/m7eUQcz
nlA0iAqsVeSQ5IpcfiQkUhfCwbwJ0Rp4elcfizrNp7WkUW+77xnz2mVx26nc
KUVqgr5VtbitAVeSMdrhu2Ls2YxWQVphSMuozfbb7WBzU1K+hOVRSFMEw4tS
G/sqMAbTSS7cVkRB9z0pRJf35q2pCA5CGUIcUcPnGJEJ4yHmz2u8lCl9QZAR
vse2lNIYg9RUyNcrgAtYMYRwK158hQXB3MBa+eYe9Zk3uMBEv0Snz1UWo75S
EYW67N34dqz1UPtWkLGEcNrZZX6SC20M8pADwXcPR5PFvk9imEq79PKpsnkA
gxUc7VaiyTyz8/mzF8eyZw831++i3vcgi5vXBaM2/mZQTDON5WGflOYrroqf
DXF+I0rBqrGv9LWMEkM0lifc/sPHJAD9CpN1cOsarG9waSzokOWMw1VFg9Qe
Fq63qk2+T9JS66rjHSrTXVyN3iSdNc8okzPKSf61H9BByDfNjHbhr8OCipIE
5ikDOnc2JMFwp2t1/cARhPG4IMOY3ht6WkNj2OY0PRewpE3M6a5tpaaGL90b
3VGFQeKsazESDSTc/O1l15140SUkrD4udCT3gaH29BtWdU3gzF8xAN3SWTny
pkxSabDJ34LazInmLXDi+zGzgX5kX1UC7qj/f3Z6TohgZyD8V61fgqJd67J/
AfbNK3hVwv7YqfAXQvhUtLgnAZ8j1F4RBmJPK3j6dVbVBXhiRr+YYys1BgD+
uWMGJS8JIfRCQhNnm9HUwKdmFgfVPCVw15g04bfLYLPxI34uPanVEcIKmQSe
ly7tHfdqC8RgWDZkB5HQ9cstj/dtmLe+21W0JYxPUYPQtUdhTMM6l/dnDQ47
u4qWANmr1QnbHuGMgowZNOOwCbE7ggJma0YUGocfIWrlMR7rb1FUhLIvdz8Z
KlhGf2Z0cLoCN4mZKAxf584f4r6+pBf94a+lOnY73CYXuEoJwghqjvof/S9A
xmsp3GIdhV2yAz0TOerfokqfTaKO57VRfo9OGTw+rGASnBY8HTwmUbn9VHQQ
CYLS162LeOpWjBnRs+CwNdN895whxzs8K91oaF3z+GIBS3OSNO1O4ZO4vYxS
Gxaj9CleKx8sC0PCazk/9NosMVi8E+qw7b0toULsZbrYJQbymDAf5K2DhEFt
n9ahWX9V8gmsQ2ufQBEly3+ZWXJ1EURy4tTlf2QR5DWcasN4DW9nK5KfHLgt
H7coULJSrTRW8zsqGzmQtCnIp5gfR2mbDiQU2rWRcyOA4QbqmmYQM7Sy8FOk
siGH2xUo+/kVdePLeY2ZY0zNk8AR2hupnWiss7JV6VA8OovVS+UbmZkjuPNQ
rSusw0LcB01JH15DgGF382OD3QydiQrkC/ogPZGETlL47gMzSi4DUGQwJOcG
CrRHn/J+aNTYU+WqkX/MkBOoo5vHlu6S8kJ+Zlr7PPoydaRZQHIsXIAyzslG
g4xCrQNQ0D1WadMrwPiSQKMcqFBfj39ubNHOLyG2yVXKpzcMTnU94NQTCH5C
DShOnnwbABbQYjg4yiGA8ptkFyN8feSBq22SJJk+LC/MhOq9Vtcv7rYQit38
bcUPziu20Kn4DNgrRuaRF9Yvl7mzXqeIgKm1YxnRpJnrAujF6CDOV7FVrBGd
rwQDs9u7vX4Jce57MJJtMAYCYGFvzz2uPBxn3gV1NyMYega8gTs8Om54cxMF
NrzE22Ai/TRYZTZ5JYTYfKqT8d711IZUPaC1Uli+QA0Ug78ns085Pk3FDT40
zLZy5fy0lUDzvThBc8AEWVz3aA3pDVYuEzFaeSpcTlqIABLF7AmaWdDMWtAT
tgj/ItZbnCBKzCiEq7wNx/pNFgUQg4CNXvY/+6YvW6utXdwO3FBCXBsl9gFP
0/YpSbhtk+2MQu2em9mdpizn7/GfwkghmDY0TQGt/1JpYeXuk3TkmF4o2riI
p1tkTS9kQDIBGNFSw9YL0mmbaAccP1hA2MW9yO4q8ABOclmDA8W4WnPzBidC
ciNybg0RlE04S+osIS4STa5XAQS/7OhHNhq1PCJ0cuFfDxMu4V2Tl3Iq1NTe
5X0uQn5tkZJehvuGuCE3PutrX/A/Tqfl3x/sEtlZVQV+VWHHPilJiKdG+yRJ
YGsb6/WwzJ+jFi5LoT9f8HxUv74HYp/wzy7YOhsfknxKSh6iAACsEECXR/lx
sdbi5gn+ADeyTVyySdFEYZarJaJlwt0U/b5TaOO60Jr6Vu0XbzEpzYwx48gK
b5+JoqHvBsElaXTCpp8RhCgWSgMdUvmR2nCMN1QcK9yBuc44H+BLWbnrRwpk
6lRBaG3N/afhTNCsuEkUVLYPMpoABWMtI7LZQE8FTz/8gqudbTOE1YUlbL5D
FXXQHBP9cbbPZ+3dXCss8FbEF5iCLxXhrYTwQciVrAIkunIhOgZgpJMtkjbJ
8Tlfm84wQxgk4USHh90In8EDUsccZPlA3BDcG5UP+smfgTTexnTa7h8qR0GR
MRpJ4WAiBcEhRIXLobNBgQHFWE31chwkFQXjIQxHX3+N1DQB/a+iVjU8GD9Y
XTptr6bfqpYY7yfcdY4u0z9NQmDNTkM+N40eQ22KOQ5EDTCQkLm9giVY8nrZ
aAfD0M4EyXbVyT/2Elo0EHcOsLBfESoYcEWQqr5TXkTdA4V2vtR44BZ6mUIU
hlEZ9Zz2QSMhG3PuiSyvonzmnwix0e3gkvfJpZibDDsN2A+/pbLNq5Fekcub
oL1aoDYOg6Y+Z4ZtVNbGYCTX3QHdl2g4cV3UiFUBv+ZbKynCQkA0bdrpNXth
u40kl2DWi6dsnSYxoY0FCTdvjc7UqjbELSHD2QeXIkdrYWGFNNTL7dps87s9
/VxPRxKGwZZFid3Kn50CrhB4UOTy6+2CkogbMQkatlUnrmpr5UWaNiil08MR
nP3Qo13og1sKILSyBdxqeYz+2l/C7XfdmOmSYG2xOAWAio7soQFGxDivausz
0PLtWciKKY4qZydqHbNptKzUn442lae20GesgbqSYYSrwcOV0pYpkVcSU81C
IWJcA+pKxNNgMec+JF5x/Qpe8VuewQJzTJQIOkqmEKc5mQmgokd514Kt4x6s
29j4uDLPvopGBeSIOe9/4MoFj96A+7H4cB0yE6+o8sJ3ir/WG+TuMiY9rBwd
cbgKxSbCuDo4Z/BMiF7FEgiT/Pdo7NtlLZxhuCONMFRR6k/P/3msSkz9dO5d
gPjY6H5ggX7hXi20IgPrehlWavdlLDJk9pIEYkI2j0P+wvFF8TpwjYqcBlq+
EYkxu34pcZmYWdfihmBq02pgsJ/kmaPAT50jK7HO/iaLdOUZczdGy1L3KUPz
gbf+8LSVnuHUgZxHb8XcbwXRreANC4XkMcNMXEuF6KX4SG02Y9LHW5nsazvH
5OnvSdy/iWla6LtumSy7FWUFBLU/xnxEJS4MJZp7IRTsATRA8bQ+fwEiVUNj
s6Mio6drm65MuQig1SWlWEOaDAkfqo2u2qefnlNGfMybApjhwjmuOfnNmzIG
pAffmNleuxSXDMnUNEWhiUapXm02idO9NtykDccMyBlJtupPnkPq9Nx5sjCz
PMHbCw4wYaAmU/glh3r2S7v5YYdQ2C+fXBpkUhLPnik7AbU+srqbEhZNQlj7
JKj7RqD5msaBM44UJpbSuOS8Z4l6TZJ86f+hBYFJCNzYTzBqnth0W/WFXdPQ
J1Zcf+wYFgDajtSWqlk9UkmTpOTd7gxpF2GIEYnefZuW65ZVktD/1uwX+zMf
fyFu3kNDojZ6Qugqt8HzeEw7M+ipfUXiogwRbWTBdPyGVx4yM72bx0pXXRF0
N9S+ZkzCEWeMfe6PIFKuE3XrBgWwY5QF4sqJfA5fiAa42wuVzN4VkiThJjah
sg4W74pMbjsnpxdniSLzFAHIOg0g6uQQfZxQpYkt1ZWRcl+zQc3BrNEKLgId
a0IaEDt2V7BuezIgEB3ssuj+UVIz7xNLvdDmk/0CZcmUhGR7VdHuzklpSXqU
UZgjwkIWg4SdR4rvS4rDEyY5St2qFLUvPtuNsYPY5IqdWjxqggckT5q81ZfF
Sxcs31An9BN6eJ0hbi7ohKpJpAt0p4+Zw3/0rZWh1kuXpsrDWeL/j6rpXdXZ
I4xjR6soxMvR3DKuE/wf90Hl4+Otu75dxuYgrr14tiXm6yF/QtiuAKdtq+MM
bYOekOI/TmuYABdkye4e816lA3G/XQdea4GIF7ue1iHnF3GQ1MeijChXWVhM
wZUKC77e8MgPIaQZ4MS5UFSN+wDFdDYoHS1tsqkvMgUyxq1Mcw4pMN5y9m/4
tRHHT2c4pMOgo+gWt7VlbFVMPmvZLn1PKWBABLUNs7oq/6JO9pmgyaWCXDrj
gdn0V+xLh3e0bGRvReJNHk0vJMfjPzBkuP5ZBNqN5cwJ5/0Y/outRwX1Jmfm
S/LM4wQ7hWw7mTSi6HkMNK3c3v7m6z6TUFWH326QCTzCducXXCUSZpUe9WK2
YbYBYZxGOWvcCAjomtCARpob0DZBpOM6nPEqi427iVKEFvuwHWUxomsMFQq8
MriL9eWMzbsN4qMnRTEHm0Zrvz9qAT5XK8pjC34XUsVecFxo3dqwJ7hiUf4l
gKiaW4sYduHMm+xpOnsT6k+CU5OuwwyzjxK86WNvDSTCfsUzN00BqgUGK6uI
GfIRXISZAHBJbJcCp0i7fWYBOVcLZQ7oS7HuZ7Qsqu90zTkPIV/UvveouLpn
nv2ZBndaKWgyHq6QLsx0BRRyILR6B1VPm1eNubWRXBQrMJf1SsLWwmyL+liM
h2+lgZcTxrlnxJNYiepwYQSDlUB01zQflWyYGkZ6CAmiA22oZQWC5+yaD6Qd
ZCHkZIY5QvaXOftTTE/7sFgDFsoWeV5q4po/FkqL8TgIsPqj0ufTUALzgkR8
W5226z6GoJaceeVYM2x99ap6FwlMQR1swzecGIGolWLoU6rUmVGk9HcoJlrm
xmE8qCEjRijtWA1JES2SbCN5sZ0SWzHKPiajECSYDvNqRK2S2w2BXSGVkmzi
6Lhk2q+hN0S2CnXqolzgpEEWB1MlBuSp6qIav0WBdx8BoyypKtOW7Nd5HQcB
JvUVWLQMREWY5isHHBvSpG5LmlaggDinrWTSF6fQr+QDMVlY+UfR+X1kIbvt
jJzWtPvgPngMKDC2KcRgGN4mGrIwwtAhq0AExOs120ZbY0vN1WbULGZg19DA
kLGQqz1PvbbKP7PwNXCwnHmkdKJoXFGYXIB4QWHFRAIwDbILtqwNG36aQIjv
SqyMpivRdyS+kwwErYF+Yw4vxG2YqBWbyUAps8eqvpVipSPz8MrMsns9uryE
LPyScBMtWIJEtlqykHazezYNHO1gQh+OT6usGij8n0QVwO7SMarcwAE2g2WE
VfuRMkazgEauYkvBP3yMA+xpaE5lXmO6wdKCrLMeTjhFaJfIQuNk/2mp5vxO
sYHtfofODyRnN1GY+oQsjcsD8Jz8AaackR0+jNh//iTgm/aHPeMby4QWudtS
s5JRtkZJ9F83/5Djot3qhhcFWgjscKwPZlsdWMwBQCL33ukWHwACRRWKFTVa
fDAcw7ToTm5zGBZZKRHIAaXqta+laZEEKdS/lT6qofOcpscVDaZ7B29k3rU4
SNZ2iTSUvCMPpUIA0i/B3t6KnrB+P5iJywtsTCPIsodV6AZBYCeon6LaBEwX
CMRYh7dP2j7aMPb/OoXkDEPW7bgEOotNiTCwzOzRscBC69D7N0Y7PF/0eVvA
EpKayVQZKNdeTg0bZhrm19l4EgAZcHZqQnZ/ZDRdLLHmkNbJpSozriBPF8DX
WExXlgW94oVukXoVl0mwxuVnEkdJxDDJLxljb2auVe3xVoFltFlv3X9kk+tq
Sd7JpPlXoGGmBLkWT4SM+1O1ZOOtRgbOF8o/r5a8NeDCRCo4ekz445NgoOTu
G9XcR7YMn6GLXWA3O4VetcGxfFQGphTnBshOQ0MF5LTd1azZSxrTLtqmtO+c
ZTX3c89vuclIV4oAMNesTnqcy9HrNGp9xMT0cWSnluozzuxVnaIbd/kVhDfZ
0JcBRv8HqbF8Ew4x0XNTINlUVh5UC2Z2S3Y+MdHkZ//znwRiIh/E5CZyFoGh
/fTs90l/mIQEuOa4FkALf78ei3wW+YEuCX1zjY7t3pYutgC+WvXuJ1oAF8zm
YA/WbmwY+YWn9Qg+ttbGIx5NqDDyIu0KzVgo/JPff305/OZ8pSwGgaIRBN07
Np7hFwZFqVEEQ35opeyXyO+AMDQFNVdh/h2pHklAr/IV8Y/TMCF+j9z0IByD
WxorIjfJSv+hH9//jV3nF9pXVnW/NRvqXpjzvlBD/j7/d5XyHVObbbfYLsam
7ACYbu/OM4DaY+Uk2kIznQ4+r+vjmW/UvdZgrfJgpNJPTe+FQP0D6jke1q4o
JwVmJ5XnFq6+PcKuReMQ8+uDbgGu9iC/Tgl7KP5KPuM6iXsb6C8bFFavMHoL
tsFKZ2h76GuGY2xBVFxO4KP9HuFstSIv8GnGq6lzWJa1fWZdpLcZgw+/WZ7q
bf2agum2e+viGP/hhsWQR/y1WBPpWNXldUHutHroXHSsmsSW2NnoGUeZV0rm
dVBCRpj+PTx5P4l3XqnmhR16imszBKB2q4yekgE4oebn1lItheVHAfeNzYBS
xk0vHDvnYgPuizaEkoJKCJJHcK3/m7nAy9Zgw+08nD2ct4OSy2nXKCWAlfez
n2E0xkJVLEOOYkTTlyliXe+0krMRm15qZl00MdyTKsftPHr41ylTOvtsI6Xy
1n/t4KAI3NHcTxWVxESS6/kh0MxnkcvuPN2YwkxkZwxPa/SUtUAgPj5iWOIL
cgITkGGBNuDLieiz+TvpXLllYlPYkpQ4p5ArM8rmt2ckSvOdQolWq0U94Wcw
krDfWp4Y+z3yPrSkVHfV10Og3qIgdp9qAdh1s55aEPyg9bmE5SMw5Rjf9EPX
o4Iodd3KQfC9VZ64Pd0zwJRBi9Z2gh05+Yxeo7T3Vj3xESx0JTDGPgXmGJEd
N7V+e8QRNrZ1ciaCGDl4MGCf3S12XO28LqA6Ns7Knvh+KAvNbayxTJ3G17/3
sePu/x0rggGSZiJ6eFnEds9vgy2mDKUgYt+cvylQRrnjmF2IginpavZkP6uZ
hbZaJiQ+dpo77Y5jcheiWdKeFG3PMEyGxWLzAJ6ZbK02LzhTGivHvOBeRfDT
4WBSyWOOisAZfLBT4uoeMIWNvKgQILSBP7jUagsjIy9blrKxpYeqjs3gea+m
BscNkSojHM253tfV/BLRwtPfC62ULeYK2Nk7XU2fKM3ECQdYM6i3tMJFuDNH
8Gd0cQPUxuLky9uAUpULyQDJjGRL1W2xsLeQ4XfgTRyt/J9ThlBqZgcdS9FZ
GYvGXHhD1jLzKvdQCrMO5jom1Bz5k8jV9zs3/JnkQ1UzQQE2COYZnOq0V+Ov
NzM732/ggD1abzyu65MakG8iCsVZSb3cjuyAbqlvube1s+e8QnoKZGOMrbEc
/uK+rzE61vZbYvbqFf+Mt6Xws5vXHaU1nNs7y1E3vKJZysNLhqPak4GW9wJ9
X+anebPXl/OfCMS5gBVD2BXX33a4T8y/N9BjBF9XLwb/8u7rBFVoAJ94nYaz
2ENAg0+qPlXhuc8iKbohweapaUfcP2RkW4iLicvtQaJZyvEOm/f5g3/RnDxQ
S/Px9LWt48QL1alJ6DnmBoF4Lps1MwOYVPRVF6WPkE/d66J0M2D/jKii6C54
Biw/7OliR5wPF/qB7E/v1HJ+P0IJ/NATbbKJj0NPA1/SNLE1ShTU6LHQ9ioT
3bdJFqyS739yhzqJGFYC043PkURWFscTSIVa1i/T1sU2Nt5wNKs9pvdZZzLr
8ghkbI9C/0HuhyqqPo2Zz8CvjhDbCjPBVMEPmdVzpPO2GIjSkKgZYmFDfXmd
NSzKEAzbXLPn2PCy+JFWrsToa1OzsxhYYhSA0jcb6yenQ2co7X8GEk3NpMWM
5RGp4hxtsS7Qg5MBc7Tlrz6prwTi6ynV0xbBsi+ed69hqRAhUn0fqXGF7Bm4
W+aL/MV1OkUVSVXDqIyxGtDyFykoZ85e/ZtXhqYPwOs0mDWYIem7TPmzbdY7
vXV8j2A45ydgdeSLfEdOz0AQ5rTrjLTCkpGJ6Uurs8grZ25wxLYztmJBZ8BZ
TAQdj6Cv4ezWBvXT12GY7M1zB049H6pAIEkpa6qh/ZWYS0hZtYmuryaEKSsJ
+oWtBbJnkj6KsngVnNxq1JvOH54UbSb8Zi42fujsm+pjT1j2AdhHzelFx8Rf
/BYgn27vn4I3v9RTRg0X17p3fj7xRQZxr1ITwISuW234io6Wr2b93Xr2RLBy
Vs+eB5snUMVoPSkif6cdzoZtAmiWAvEjiQdffl1GaeHOiV3TiWot/lvrbNpd
h2pIDR2uJiYyQx2UJxsYh/Zc1dzXGk5QAf45Oerm/sNljOgr3DUuvUlY3jsk
nQPq38DmjNY6ZLmYYBybcZMbcEoVt5xVXnBMBpJtG1Crpy8iINKtOiSrx4ds
Nop9QMkf79jxPywfPN31gT1k5HJaHCrSy3BJEtteZTx3QA42Cmq+RaJ8xS3/
H7X0YnSxgVLljBP+8gbcybWPsJp9Y7Se3GaJaKheBRC7ASVezoMEr7sXC8MC
rGXj4kdXE35+5aCfnJmVSS0RCdB7wR9llb0SzMJ+V70mXhA4n7N7QE8+6d/D
HdYGudcSZIgJBF149cKYmOWtmuGvorjGdzJV3cxc9v6Man+DD+fOhiX4IGic
bD5a/43z6a9arH9eeCBnFzz7zB2HKRd/USd0npYQdBgoHGSsT4WIzjqiZSkX
mLCrI+gMNou6K9Gge2TLc2uEFleX+xTi/5YmhIv4eS78U0RXeIO3a8myU8Pb
MJTKuOIIIAgvlA7RlxYVDnAZzXVhzYHx32HlO6Gkud0uUyJNgpDTQvQXLLaS
yZdLFRaEnWUYPZhQqnLop4VtYGv8i48N852UN4zqQwefsT0W4P0n/Mr8oC54
MStYEH+Kc0WcfW4/PXnGKLf99n9q7qzHV/dsKUdV0PCcjOESeFdkjkYeWi/l
yIEYjUr0IkPeEkq/4Q3DUGo57sL8uYA6yLmBJQwhuY50u0E3a3LQ+IHFq+2c
bAhYekTuZC0H0ydrFKq+kY0HFgH+mBFd9ewROsfW5rQI4tY79/4Ziim4ss7o
lIc8mX+mC5RNAJ9F1oGhFBF3eE4ZXP+Etwx4vFY5qOaY+Fj9a/rTl8qeP09m
4XtY7Q6zWwYeFxyqFqE4OXI8vMM6x+qGXfdQI/YXOhSRVrfj1LMsXiIPnAcg
ynK80sD5JQoLOpkrmekSDUFo4Nu2PVSmXynEKA+P85ECVzaIaMWuC6mdSDkC
5znhNpcAr96vbADmyHznZxAdpuS+AFAW2pq2iXRJgaJK9ShMsZ1JLSiUELL2
5PbEtkyAFUoQ4YmovF1MZaLYRsplItzaU5pOS0Qjg4ESed42c/3Haj9UHhXW
pmbL6zadha2KNvwOaugsfIf/ussJ6bUoJiVZS8RdISlNXP9qILY8f3Ep9XKz
wnkT/dSHJWHqVs7f9v09P3RHK2/v6ia7TsGeyZ/BejYp8oiTrUM7wOzFvCiM
oGEKgdCNA1zL/qH64o5CmFPqzjcsIIJluqgJ20o/Ok6CCx+Fye+7PW9PSUIh
+/cZ3pmTgGDQfjACWxk9VRJwgkSUI0xs6hJKSJxo+gsYb5aMr98/TeIH/2Kv
djbeF+TMDX9eHFiOp1ISaL91V8Uo04clnEja0vd+lpgo94IM1yDZdwHHXPGU
8SgV9/t7iWkRb/MvIvm4gJqs6nAbRF1dv14mKxnvLRBt3GYzDIVEIHjsIQXA
CfQ5gRstzhv0D8zYDzAl8jjCaR4r2SILcB20qRZHFFITdyvY5v3kiZI2uvDn
nFaF5WBjBIwnQt7hjtk7Ro7GdN3y03LcApKiLEPAWFwe4utt/hM8y2dLxEuP
H2nXGTDMXHv3y46MPMh0dvUipFPL3t97LNOQUOdjBF/FflsV40kqGfM+OFkh
oakB47xMZDzXsWvTJfHvPEu4xX7DlTJOm4b7/BUD0EYs4nahkGIJanacAbGn
xgSuQwuYMLuyUVLTmurk38r99+qNLvzLtPXAosNURQ9E2ci1lg3JlsSkOMHE
tuqQ5U3qajLrt4h9vJ6D2TF1QDAJfF2DYkqKfCFsSPtNX4gAJscWDeJ+Gm3B
49IMdb2eDeXnUSsMR/sgqpMAIBb2vd3Y2eTR4PYo0wk0xrn5JWHrUtCD2LZD
Rvt5Gx8P5+IW/BsJ+SubCz4EaN5oYTmCsxh+zXJ1aDFUUgs+jO8ArH+Hf0Cp
6W9ebgeoFKg/COh3HPVcQSJ8uQsNCVrOWMqi5vTp0av/5WwMBMu+ktwBAF+1
KVzukjdSDwCnlzUNeclYl4J7S5p5meobBUbfoyMXl4CfaPf/8xXDAGtn3NE8
CMl5InqUcgkcFOLGQ3OYtAYT2gm/MYsBGOjpR5Bd0kMSVwy85E0uq/q6Qhaj
O5Y/uQl1VvhWMzkR31x/8MRq8vrkMnfEyuN4qwStnfkHykfIbD4t3ErftKaL
KllBg1ToHyJzg28wW3xHC7xG3Qi4lcB7TFhp4qXHlexeKJe7uy3/liSbCQ/R
uJ9c+BiQTxSIbe6X9kuIMXqBfIp+DI8lI/A1JnIHPh1HLBEPgFyqZsUySCe9
qh57lvFj3ApEg+u16DGks6wALDxXG5pRLqHwWpLt7QRzpWZ+FJOpVEBgJmhv
5Lu9UUMuLssCA3hkzPBH+p1Dhu/iyKPdJ+rD4OrJkjZuYVLmU3aA3RsY+3+H
c8+pcZq9q6Q9KsetGIh7BagzfPN6T1/q8WhCZYutZhTBdS3MjwZ803r9MHc+
zm5SNGiyw5DpDdDNoRbdC5MrT3Uq21CFwjeR70PLgWnklSm6LTKqit/DeSgB
a3Bf3skQNA5EzySjcqvEEso6p6AERMyaaJ+As2PuHoXRD3fISODnJ0MPk9Jt
6zcf7wKyZpsOJ+UgZuJxQ47m6aQVm4g26hHTOZ3mwmFWrpdhCKkPeltciplt
z2fMl2PhisuROtK7+X2OpDqD5iSy4hyFOs+f5gJynB9ZhVgmr30bu3bdH90x
Gv/QOJOUKiXqdwkT7d3ZRTJQfjmAA5pWyA1Ch+Oxp4/o+TOp3zn7Ef6tmzbb
B2pbPem0YTf3s55AaiO7wTCOA2pmZQp7KyLxZQYelLQB13+JwJAbmZ/dW29F
YTfzTWfzi76qfABvTKnWg7iF0EOxR+Dht7/Ki0iEwafZ4Xai0XTkmmyDO0xk
vcD4boJZBIbKwpsvS7PnPWPw88jfIKaPyPLRwep9m4HV2bAhCCrN3iOQzvAu
lId3qKazrQnqvwdD2xqQQyRaBiuRRyxBB4qTy0Qu0IwJjsWNNsRycVjih4Jj
+s9C5UPUDbkH1RR7es22YlFmmaoeJdafXtnLwGTY7ZmeIXmg9qKRtFNkNvJ3
oVcCl1VvPu220i44c57WnUl23LgVwZurxqLvKuKm0TDbUF4FZ8QkWVnsxjWP
7zOscsMPLJRYwsMVCEgCvv19CZgWmgr1XPqbnV4ynR93XQRBKmtKBrwU2Bei
mOlwuEzVpxxRibpqkLAZOo1CBRLuWa7eOq6aah3j8zbhxo4g10ND9uHs97Co
WOLe46dDcfnY2YoJynShlz1DITAlPJs0N46pttjmxFss3oSW3GBdYRuWrjcA
JZzHpBAhNyG1ImU1ybsR0d61RFY8if6zlfcJc+I3MALm43cDUlO4om8ZoS2e
wiKwnn6+tjKBVGMMkYO487s414H1y2IMjuWXPrE3GkCUSi4lI8iyRPtM1Kj+
RArRRg/G4HOxyipWQT2T+2XPKmln/cf6Xk+TaOdjd+LY1NNINJOkFuEu5ZXr
a0/CzxMc8xbxm3gMpAZphdIPr/0/lXhbH6t1I+rgAZ5MknT4O5upgJuY2iWJ
N3LE46rbpNkr9CqMs/QGmlRb/2fKTDJ09Al88ZemAtdFXvqFQtG4vlPP1oW/
7jSegtt98qzjHoG7wejrcv45xCvEzU0F2h9SQHl0MDiT1awJA/MJel+FFFis
MZ27VQrCgb06AKWm/LNe8vfsK9XcfGW13c48aIz3YBjqsloeVEQwOVej5QuG
XGQHjH4H6CrFLzWepOZB2+e5zQksCWm5yg7TWQUOBUKEVeEojGP1ZFvcAXss
M2Jt/93SntbhdR1gwDRVmtI40vVmQ6oH9rgw3B3u8vz+w+BkcBq/sJWP08tA
qeF5E549eLcNNb/bmEnJxbtpUrdJwP0Er6ZgDkSOq4hS4GJNhpej/wfsqZ7c
WDFaBkMo/QdS1o46Vagp45rRk9pv6HEmF9NY1bF6Bzg80E5vHLwNOqXwqySX
/C/cHVd5ywbqFXXbbozdmlsVZgajyNTHSu7kR9KAF/7N8d8tCoWhYOYRB64r
amqpNJs8kGKchZyMe+Vyc8BL1T4q7xCAaq0RkyrMRGCb3R3v72U1M0IC9AqF
wTKQh0dTLvm4nknAGzHwLUZvOFO9oKYj/gG77/zbaZEYIWO7qed4rizTfYhg
rEOvIVzIoHkADt4f98UkSW+D9vGX4g5FW+Fx5G/DVuW0574VydpnkL8rCmaB
+pofHIeqHgWrGe3oM7VPkKZqJm/GP+pgyQyxWebj207QBBu43WbW9gN6wZwz
X1j8hzimB3BzmwnYozKyBpIeoSLaCuoolhxzKQ/o60Rpb96KTf5zXb0b2KOj
z84Kkbd3d4NQ4uAVAFXzukYio84aDpqQL9JGAFODgqizt1hLjjhCj9lfjM/b
lFAfo+NvaYqTXdRm2HfGVK03dpDTXsAVBYt33Sq5upVAp1HF+W2dZOd7OKLg
F2Un0o7PxD1wc8fLc9QQEJk5lT8B8P1YOeOU7qGFEKk5CaKjPgDle2A+XF7A
kWjOgaoikHRQTSIRb3SRFR5bwWPlrm8J2z6vGB7JXx67NnPkM5rl7moYRVQn
zS0e0aHC36os2CrrPJXFC2XsXhVGrRpRXuh8mHHXbDA3h1QZu/wOD9Slp/2S
oSDzh+hvcCRXETVAPmXdP8vKqkgXoWe06eqYTv6bwFmeY0HvxPhdgplWd4w0
gTuXfaKzwhZojCB7BDlkYCKWaYOXLD141+lhJJFRrr5KgcyA1bFhheE/Rzg4
uEEmDBaN6e9od7yRReGqwK8rZd3oC35FwiBBtZTe3C1iJG8vqD8o+GIc3Pfk
3ZetT6NsXcZlnxMZbuw7zzUckJ2YlQldpJ5jNY59KffHchZvcJ6nuwzZuK/B
LNUfY3FmlBT9iKTYkF6jpTCu/N/DaXebMO0DpqnGEd5n+8MT8+6ellS5avtl
Jrp4pefGX/sVj8ZfGf4RbT2WEYKbgw9O0W25XjEnnU4V4dygzOyN33oH86xT
LJs9LCbUMdwMd2FKe2CudOuuVk7lVOQ3+k+5V2n9mI0dHZDqm7oTP+M1HHey
kf7vAGundiDRSNXcojMovnoOW/WIEe4GPGYYmsIQ3NclNPQX5ihso+RS5Qn2
mD7/1f6U1P6QejCqiyytqsH1xAdvBL1Gz+Yx+5coSIaSvBLRYcyAVqy5rJWt
P8tdxbuNsNGp3YXeuiXK+JHOxXVClgToJ04OJQ2mw3yjTZyRnWLSIhJFQVn0
RkZeF+AdeQFq6o4DwVIwE6DlVhnWXtdhJcKC2vm44vZ7CwSVwL3m9hh0s9I+
/o7weNb5INhcnQKv3xntuP7U+5YqOMGlmuf9i+AG0VCpByIr8iRrUINfzwT/
UMWmdfeG72yuYeMw+wSa1qDIe5cx1bwUrPhTzCvTjPiGAgzrZwe+bPZU2CX4
Hdv6SSIERKOUaLU1H6oXX0OQ4CtU2331LgZnaqkLLjfScIm60VeM8qNBZZJS
sIXVwxGHS16aZwLbAPjTuSfHcBh86QqnZcdbBzHZ/hJJpGorJrJusqpZXxqW
1uW8c/+Gr5sJhr5rnqRCKs3QJDhIIvbfD7qvkKBeAfBGB9od2jr9xYaLhtTN
BTKJqRm7km5xu9DUm1fAMCVvTuz/iSpSbGkgmprpUcs1D1+yPRYq1i4BHUsk
S1VI80jY8PQIJIGlBJa93Mfj6Wl/v30nairFDHmEtkg8aiMMA/GaGWKNelqR
DoU3riAN9EuvAipXr3hyigVhNvn3+aQrHgDOAoC3dmgbZoa6TuRvfN6eGn3l
JS+SQKG8z/Xh8KSaClpW6LrWt/F7ljmjvM+QIHfWrhreFK7FG6ZDUXk/kq3d
TnoXBfSKKeGVLih3/dQaz+f7Bk2snBIh5aEJtUcAlS8Gxa5tbpX05da5YR60
RbFUL5Hyh7UzBm8i+z2EM+s5lGm2DwmqtbvgX34tm/VbDrdc5ay82R6PBzm2
BqIgtxaUvEVlALFqBUYzMnoKqsq0PuMIkWLBx/p4Fm5WYzQk4TLf1zj1QCGL
grv3miWRNztHTYfrmXVB5N7RTUliYUJsMmjmME+5r3XLbAmuh2CaLlp6cu+Y
vhv2gkknDkqLaDQxCet8OTSRFFxEQXiqhcAJrOrWEQG0V6DheOPhjDgoFkmU
LBcYYI6qYIYg84/f1a8emlJdMEElQMZ0c21BwBg18EsPKJmHMKH0Tzz1QTee
o5ithkg7zDm/tRBr6oVOpSXWdtFq2kebtLTgc7PPYSFibG1W9DwkcMQx8EEg
57B/a088YPQqZN+9rOV3kPMUwPmZWtBQVBZZKT5U/kJL0wrhbVQdJ0Y8jZB+
+fgfX6ionQZ9Ubw3uvwo2+craSlSvV99fHaDtUjYsLnBFQeWJH6DNNVekuru
0Ae/BubI86pxt5AcCxFq+TjFpfRMCnmE7P1a/FpH6DCHMkcHx05Yp2NGM8zF
uWFM0tNIHcL+swgrHpCOmOsjcfDBg6upKyBWki2Y9ZQaSppVW37h4R1Lf7GA
aHiPVhTp95umlBIRmZJmfv8hCHEdLVHOtELa0PugJ5HNtWhNbOs2nJ6P+lP2
24zNwLQ4vOCrhRAnzWg3R0l/tUuEYFELf4/5CX8Ev++nO16vzzAc8XvY6QSs
Li+ogvwl5x/xSIKkSHYuoyQns7wt6MjL2C+jZ0QJaXnMDbLevApznRIR9C9b
3rg10/cMCsvedy67JPVlyhaIvDiZO3VJ3SR7W6mioCQKh3UyyRs99xxI4Jr8
8LjQsyfWo7INCnl2GCLuA8lexatw9xd+0wtz3K7twpnuK5e56W0Lldkw5pq5
VRKpz659ciO0m3c9VrWRJRUAMepvF5Ngf1KoFCFU+CcwbzLaHgeJz8JDsqel
VZFgFQsjM3H8/xpqGqLldUmHbRIFmQpzBg1QKvDya1CaZGS6puUGukTuO3Cy
5cWxgTi9NzhGW3XaRA4xn2Q0liDoufQbltG6RSTzvlNBqSKpbhhOD6yiedrR
qQ5B6rKzvJxJc9dEFQ3tBhyop70M4WITngwtyWPMWUhv1SWOSs3ak9kRlz59
TLFzTX3/SCNmINl/idKANGgcfwAwZytDh/9cP97/STjRX9VxP+DRl30Hsv+/
MEcwcxV05QH0i01uP7qbgp/IsYpKBChpmjvo9hh65S6wWVKbt34vlTjjGI2T
D82XODRXEUo7RaogQbtZDqtYbaHICYtIyi9BAjC1g0pwbn7SjvD+f4VxgV1k
al5X156Z0slNdGrQUwPUcbBcfESb9Juyp9rg0SIKX4IEioVvEiC7fY3bfBZl
18+SbNU2f0ObdAg8LmEhRU8WyMmikPznVBREYw/dtIkVTBtntU7BQc8O2Kbc
5L1TT6paNaF9vInsLfny+GbQOE40RyCguZxyl+KRT8I8Cz+LcmTVLJnicGNG
1xEB/Inai60Fo/+reX+hiucxfbz80HXY17+SmLQaRR4HENuklX2VqMoUVXQu
bWYJmOmGh7ty4C2S2pKjp+sOXomtRQ1rhVNeDnx2iizsI0mv1bmaw+oSb7Qz
Tqthku40e930Y+e8BGavkLBJpLLF4A2o610FD/BlD16dvOTltnXKbDKbDUhD
UMzrT8eNwpLysv87Lu3p2XThQ08Ijx/hyYAaYH0F4j2aQ8fxFzjPVyfbRecg
og7VnVj/akS+XzxFLwOavdVY0HBsF/KECGIr9tT+ccZPPrqBflNJCZu0tUlK
Q5KHs7svX2xKlnfycuNzs7skfe+qpuNS47SwGuOKz7HozND8LLyLrDXJONuL
psB+VXFvpHXtwKZS+BdeIdiyZ0a9kSBgonIZlGArDOpb9mbXF8nvOuyy64Vp
iQMXNbY/iyY9swO5FgFF4hLP/6njrgu6M3uL+hnGWE/Dh181sWYZ4ex3wvwt
N6wLYe4+LeuvWHfsQVBoAnc2/rZ4+R1tYmKsiqxk1FTajFTXlXFrhb7xIuSr
bZigR6neMI+4kxiwcCeYB5Z4e02FMluRQzfF4V8T9LfqTeAHh+yvhWScO7o5
3R49F24A4x2GHqFq1RkNKCfLp4xB7v9XHz57eYdMkRiGbPzBmf9lGBKUY/Q4
5QWYmk8Jw8Cq4DoN41c57QYZo5kzfoBfleb2ZarTAUUPJoZJSLLolVMbdBgG
ICvlWFbEbg6MOHxwmP4E2lZCbQMTaPjBVCQ9M6ZsHf5OruBA84UBFFuI1AFs
LPBDDZPrdWBGIyl37V2EoxtlKOkJD3N3JLs8dTb2g+GKLYcJ5CfNVXYwd+/s
WWaPaAivyqGIZ9Q2tw+cmoiqnx1nvobEu201aRh+DXiLT9smchje1iRBYJBO
jos2rk5GZr7seGVigPW7T8fOzJ/jxDiKe2E1zzSbYy5TAqPa5PFjJztC/Npq
fKWErHi1pDCn0R8w6KSFyIADdZ9cd95IgaDpzjd1xWpAAfX317gmu71Spf6i
ESwQS/x1VYd+UQYAfIvSu2BoGQV2Xmpzp4yQv0uoQrNjLOvoBqXJUtM3zbiw
8ynQNA0l+hZKG/ImXhqH99GR+zJ52yf+68cxtVvZ+PJROn1oMzP9HI0NfoWh
a0eYrWqRTGKryE4p49UaRnq56BBlro1JhbuGRi+06kWbbGsOsWNf+ntHBrMN
GVLfV9NSn7dsMZCthMfdRHP0sl368yJ6iOPY35wliESWZkzV0Kva9rHxLIy/
agY7Sa8W1/ETOPYl5tKcHMgRxTqUza5hPYut2EQJBZQ0o4tsjZFuZeOcK57G
FTno4xgrnRwqGwWumy6K9NhJvUYclagBj9JT55+L/gUx7wQbqFh6HGbq2Vgx
kY7N2ZFryk4yDDM3X/dhZCsqglLRUKCOlqTni2Mv9QKlNP3bhI4t3q8ynWBX
kbHsn2zBU7gNr2c7YjUQVWmpXkveB2uiU8i7HJbDiJej+4Le3cMk2LHeQvOt
xZaGWOHUo6sqiV5GwK7ofzg8e+m17S1ucuFogjD9prylE1xfGWukhKf2b1dw
CKcLDn9fuZjXCgiRJLixyg8LbiRF+5dLodjrzoWp1s8wq4DVcCEK3Xqs5Kml
t05XZ4QVDd/26UYBEAZupmEYVTL+PCQXkm0FmveT5NgptKdl2/r3A4PjIYsq
qkLNRQNKjkwtjOvsyUVRFdr9wsbtt6qhAD+hxL3jqCcKigX7oPR3Fb+zPLiL
AXA2nfShutYMDTQLgRIQ8/Lf3nodgMN1XyZg0Y6N9u/NN0wWV3pEh2dAbNRJ
xYym7fd4E/5ZDPD4kSTcEjulnaKcV/xQf245N9e82uPO3dKVxKmHYPa2/jew
i/5MTyDHh7ATsmv3JuVNdeOX2XJ0pzRle+K4Zj1eQsDTAcSOYslsoXB8URC9
Oo8Fi48v2IiveyfBvAhta69Mq9Sw9BiZm7rnUh9FjUwWc1+SQ7lalLLOs6Gh
rpqHPJ7tFJOWsW3YOU/AE9w0YCKqsK7W/trChmJfxpOROkrt9PosNEjA+fG6
6QtSawlOGpHYjk8R0Q10Eg6bUS8FPOLQ1a9jgg9tY5YQ68NjY9k0bRTNpy0r
ybDk37RrVu/UlTTKBt49k+2bJIZdcdchMSfUMOTYYbGxBhOh9hD7JX3d3cbX
uW/y8my7vakM9yUkbdoCHGBoTeWIo7CM4px7QCdBrClW2bZZ1W6l8RR6LQfI
Orf7pLBjjX1fD6Hv1SbgMiCcU20/L/e551DHRM/Byph6OEhX3QeElw1Gms7s
qwgG1FQS+5/AFbp+658fGx7vJubvHIIseS3Y7yqh1Ew+4itrpv9iYkCzX9mn
bVHDynFPN/L3qhNXMIn1dEr2OCu7p3M5+0nNPu8bvrWaTvS/OnGiuX9Sj6mD
2t4SdcH2hsoTx2Eon9ZuWmoPZLeS2t9UYkrMSXbODD0JFEod+E6H4RNUSAD1
NXnsIPq3YsSk6le3Iimepcb8nyk/KpvBp1COeNOMLzj4BS42PT7dt25Gx4Ho
Tk5/W5/cpqUkFzAQFaMWCpUSIQYtEo0ql8L5yDi7n3PUGZVSU7i3pA3D8Le4
XEP/1WGC2f3+VZlP1Thftf3G++0Zng/JYnTYoWWh6QMdxxxFO1b96vOzcong
iZ6UF440jT3Egf9nRKcuqTYXh0tR1GIdAwed7s+9t217KatEJOpb8pLNr5YZ
UZ5uu6La/WD+Ijw2zGXGjrcNyixh5I0myXM+PaE2XPkFUmDRfJILPb7IckHc
QMx43OfUSTR86fuFyC7AM43RMu6+WqRZfxiO8QX5HufOmrLxnUBjSbwvSbx5
EDu3CZb3lJccbI9JPTGDY4XgOeV5zAPoXtAay64iARf2QFTJgoAL5KXjgWEf
OlcRqV5PVGT1cVyZGB58TLGNqQJZQvAhPHPhv01z6LhDt82s86GD3oIeSuqe
3B1qKFSsjTqSJpCxlu6eOfMnB9LRea6uUUPX4uU2MFQxWcjENKOKaFLB53ZJ
C0806pcZIfdkxth2W+IiiplHpsHMi+dupUqdwS9McBIz7+9YIQJC0IPfsGE2
rZuYbjZIzt4Kk+lRd9TW/CmnWtg+DZiJ6tGPxf9yAqrg6hz3/RaiyJv2HTkT
0JdzCAP2eWNhsMFli7oK50lqKOtKv1TT663B+i6E7Zuw9f6Lvu+zB/dypN6v
NTvk7pR8ORt+46Qqj3CxW5R57hjDA/UG0CtGw0RIaqBNQyDuRaXuHgCiLYC4
FUiVBgrPwqS+tE3tkXSqYH6YDHiGddX3wggmZb5ikMlDKc9j34HM4EUxFwb2
kFHjcPdEaEMnZ2yltdPo/6+AfKW5id9rQ8eV2QGuB0MpvXEdp8AKJQS6kFgh
AwISaiHfcF6NRxniWYG9e/+MqGk+5/BTrvtHSRwhAcit2lWBvZigmpdFuMEP
XQD18KSYh+wTYn+TxSGCpF0vdDZ+rk5v7bCsz7yFc1be+3tYuLSzhHQ3eg74
HvlfXTYpUPrksuZoLXkOlCjOhuPUXK+kBiQPO+yMieQhvdWfTzp33Ll0EH5s
QRt0OnauKRD+IHOIfPR7kxyu1GG8S0KRGZFFiChCTCRAOiDP1KcwXRFiodbs
K1qXVebxHozsB7Het7b578ayKpns4Wu8LLFSJKfeiMbH/hUZec7Ir+21iCAq
4V605ZILM+ePeq6oWhtP97/e3sH/2nw2+KncsiGzu+0ANOEX74efsWFakjMc
w/myR7ivJjHhEiY4SaLcpfd2PdVSQTbbeEfTuDn4DhPuuyKRgvdyEoA/Whj/
44hSDPJfjy5GW2pPjmnx5y/S5oaKsAGdOQf8G40fFUyTekVoNAhqrdoAU0lF
OkQybJZaWmtx8pA0+YfvmCyz8uWosb+/qLPHpvN0CUHdsPQ8k4I9Ms3Znbsf
rzWN8C/P7NfURJV80CoPcqVDsyTnWrkGM3L1jKsqBR0zSDyGSkAa5vbzOU8u
ESxhCqMuLH4kaZJpjiu1RAZBZNs6NBg1Sr9LdQXtuv5jaO0dwgaW6d56hlpj
jKNJO4UHdPyYqyG3jq/211AvedCQ7rH+Aimu+isGWo8/sHFeMaI4iICZ1dvr
xhmBDihgyeAt9SWEg6kXkUnDdPmylYbIVME+Cpv95vOJAbhTbvDyH6kInI9d
+ozEooJGwJ0DLQHlsi4xdHdK6f4CzEQc6fP6drENWhZXNl4H28n6YOyBjk6T
/aatf4ecf86FzDL4DbNogzkPDAqcORC59q00qTphrPVl3lu6gpC+A0Lc0CwS
jMkQiltNZdU1nCFIt5P7tvdfrgdkKno1YQfNmHUYaRLjnBfcGMdyipghlliA
byKN7dfyVvxhSU7BGAC6akUrM53Hv2HYnVTC9l2IVDkm7TYSJvoNWLp2Blrj
r8keUFYR4PSi5c18bZAv3gNXeHRoWmzYT/I4T+/vMNagK3YHAFlIKo5kLcoh
43nlHTcmFaEVmxLI4WJbYZsB5uCbwmV1bTsoz/Kt2yh7umzzttbNoOXWVGcu
RDgcyenmW/jLbDijuM9YxEMLAqhsGxM8yukDBKA+xT5Gvqu46Cg4OtckjG46
SmKzfge9f/dOJ9vhfvLOekkMGI6Clr2EJVPYtQUXEXSn+FqtBZK2hQVjAd54
5JGxJUcECYAOdlvJtCwTDhkYY44O9rClZE/a2VOe31L691TWtpsmycm4WL1x
97zR0y5knHJmZtxwdX/e8zlg1xh/IHhO3ZOO08QOjcSbXWrLNZJas3FAMUro
m+5TfqsP83/tahyknxIZQ9JpK/9Esmm8We8vt60ajNcQoZKPZLTvMPNFBaaH
63lH0jolYz87C6sFYxsGiBOPZk7wyhgWVE1/4T0jbR+Uair5omBh8CribBwQ
X4rjSWNuvozC4/XzvnSwoq3BtIY4aR7JMoNkdP7EkjK7MWjfAkbQz4RdS4pp
4yrYV0ukkwckghwIh+oJT8HITgRvbUf+RxRDFokITV6PjF505AccNlxvFhWL
x0QVgz2mci/wv1pE8vmnyCfbD8plQvb6GCuCUy8s6XcxbbhgoGPbPt7Q3425
aFi4Sw66c2flhje13EI7e9BlIMoxauy4e4HD3kQgCqK5mvgptP6NysQ/rXUY
cmzNVmh4WP2hD7qgPT9E07cLWr5IlJ4if19hw3/jbakIUhw1AvgD+xp/gQws
ZZMi0/wNXCb95Zp7QlTb3V8GhysByngRAJbTzuTW+bnA8bPkigdsDsBj7/vA
9b75s4koKhKI+PG0VkPiwfyr92rZgGnCVO5E0HMpjM4aXzoT+2MUOMWcUCj4
eSWy/nDmPxL/6FoOD+5nS7cqKB6rg2UzvJfoMNrA3U4bjFswLxJC28wgLCZg
BrvTQPJWOcefTOz2s0VXT4+5SSGdVAuL1B/IfpQKdVW2sVNXQRpa2qHTFox0
zxIRk4G8Ik+7Fuja6Mq6A5gzYf6bkvHg9f6gs6GPvg9h/fAukUvtaeB6B10b
9yWkWAPuTBLvfCe6uzO+/Iwato1pB0AtSnECauPQrWZPySAEDDLbapjRkBry
NDyhzPx1vsNDR2ad47uc9TB3d4rDcRkzEnoMcm6hcFy7EGsitA5FoUe/heVz
bNMhK5RAeWpT8aEB4yCplvvUvoFBIdxIXgOlgn+YuOLNjrmV1cgYogUZtzUp
tqZRpf8I+neQumJNSbYO3UTqffk8JQ/caCB66NHApLTTUaXQL4bPh85FLkuF
A+g7ERaTZR/sMwTYj/XnaZQ+4oVHxS2/cdNCV+9XxfRIav7jO+q3ItaUAik6
f73Yt+MA/6W+0npJZh1NVzaqZt0zWl11Y3DCa2Si+bSHGj1UEGzPdS2/fYkG
B9YJxl1eJ7JrIs8jofGBihkz4zRNPV7KHvAVbyc37fgp19E9PZRZgTouQihv
/2JbihjG9dOkpGx3s86LQkBQ7yoZBgKqyK5kq1iM8QY6hgFpqJxSdjaSBdFo
tEQPRB3PYjLFRAlL5WQhXhGYs/d9k2A6jEqbNd05FOqP/mlvpDNiB4y83EMG
yNtx9xZuYuR9Regr6Kv8/dZEIR0e17We2kvN/N50q1dkHT+8cxgNpR1Mgq+k
m0SzxuyNSU1q5UsuAv8aWrezQLPz8W8+YwppvD71nDCU/uvUFwFGjMmfa4Xy
tBZp6FSstLdGCxmzHxHmqGkfuO2lyDGZ1r6UvWg+EDx99dyEo5Q718xNiw76
jf7j8mAOEX8xsTFUOxT1StsR58pRnf9XHg5f+lFiCg7wMcIzHAAaIcdimJH8
PVb7IF6+5gPgYYsLtr+aFQPLpghXj5fU8j/g8wCFDmScZvkp/S4WMQdKr3Ju
Dz0/90JgpXSAO56NnELX32dmWbEK8ho70QXS0V45udfpUMhvGLT+Fb4ZH9Fd
TbiSHdcN/Y2gFKKneJono5tV8Bu3Rq1dOFaGMjlbFCZxTsASGPzz0n9d8hWl
AyZePUvEkJJqY0/AhzS0LDD60nikhKh//FmkFSJRGwJA/EF1uNVMfhTnPNtz
RcWFzvWiCf0xUUxl75ZW3xFuWTmHlvLjqZnoBaXTKioUwUN39MN5PjUP27Vq
Nv2eviWmFOpEUcTuaHZHZbigHp7SQVljDUKYxu93hdOikchm1iLjLFWDPfAa
9dlLa9vF7l3T1fE+ixmuzKNBbirULc6/NvbE72PCjjRgwww/s8evp7pidkNE
oic1QK0+sqrSzxPYjgIDMb82fXnZkAnA9E5bY1p+A6SNAeCelNUdslIi4MB/
skTh4vXVFkV1IqZyad5cC6sR8txYqbR2OXMTXD8Y7YwHYL6wsvzQ0g2Q9Tiq
P/tD4rxB9hlpxQSNvAHQt/NunrtoF5jdMjSDgxuQxzaD+tIQkQEWAo79ssFv
NUMshVt4Bg7tPdOuA7EGYwQQkWrcLCjOaPbDd0OfHanbG8UY85rrjSNO7gFq
9IIrHZ9vWQn4gja+kNEQR47l12gfRIov2U2X3zIEoF56eOBqVUuYzFJD6dNg
nXdwglag8Emdvu4+CG7AFMSDPRnYYc3PM+M7/NIB3aarglOFIJlw3KywxVV0
EHyeYA6DIIyrh2zSWQZPBeBYc2zWcNxM9oFMP02K/sXRPHomedq3sr19SA/A
biaRRb/WJ29zSATT3g9tRRMR1Ln9kXt6JVUp53/LwrwU51QLux/j1zEfZrdx
8lpxKVLjnSDI3bduyMWeUO6MiW3tdSJixQhJP+wyMHGnUsyqc79/IoJtlFam
cnUGSEyJra5vZrTDzMbuXZbjcYhMXw87Av+qjTjk6ApdY1JtjS7lCPA7cFiQ
HrKDd5ProWEsJIjl/JdB6Wafxxtf7OEaKlmfFfoQa0FdMvNF/B0EQ1h2X4M2
1P/mHvSEdtpUOnLvNlP8i2X/kuaEJdnyMk6/mDaTHYBU1SQrK+dSRvnBoVkn
qJlBrtiH5xyqtM0VXwIpj22UgG0gGvuDH0e5UQEdLFtWDnjzMxB5kXVRCuU4
sctmahY1AWx01zNledXRTbv4QnVWjdE4SY0Ib8LUX2xH7yL+0qj4xU7o3lFI
UN0U4Mj99nn0MDP8OhauhJ4Jzhzg4H2ZHHKc8Gzqlmgaqb5ydMz/GPW4Itvc
N5xzJMyWsaRjqnuXF+DxY/ZUV2Djz6H1WRP/txWsEzxXTJxldNEyMuvWr1MG
FDFLWq4UgP5sPF2kLgwLsA1kk7yoI4XWN762wKHjmIydDYf1eock9dUO3bMQ
GwZLg30gMN4jcInX5JT42klDFiQPVg9xeBjW0gFVOQKTiOMr7FjiiENyv9vd
QmpZijgyNvWSaschgq1dYfFQPlq45Vhed/MFKT3trtjrCqqZID2WptMUl7tN
7WOOiMuVw1Q511MBFSfTynUn7MJuqeQd3g9uLQTBrkbzmJuCH+KM/+mgmx4z
rNZwt7TH+42R0+t7FQ01cuS8RqN3+xHsX8ffz+4eGNrkVyNb8SY44W2ul/Ak
o99cwLViUPB/5sxCeIQwreCxa2+VPHrbYTjhe5FBNY7h3RJSiTrPL4Kgv3XO
UwxciZl9nYlUg4yT2ZL96M+kKzF9W5Ibfwi7xRGj9og9ggQNXeJEnNmC126F
hC0hvmcSRtCMV7PY1qVj/PDjOdS2g1m1e3BqiA3JfoBar9oFoN6JRhWMtXXv
R6Q4tLjf4ZVaWF3KCefXzWI7Va5NI5f0Y/VG+U2ysLI4I3Bl4JMFmejoE88S
7M0dRFtAXM8F4CKnKsVpp8q2pCSUTye7kXKFPgI6AnWwJj/KxKkqve8q2mv/
u3j0uzMMvcjIUy2fAc59BL6not318BqRVnvVTMA8rh7k4Scl3d51nmoCJUyK
f2Nn1y2xMrbGIKmrvtHlS23S0cM4tGJwhXVDXh7NzXWVb8SlkOxgSCq6Rbyv
pdVoYPLLjR92qvlFCOkg4JkeImoKg1D8i6OC1ewm+xOmLYAn2fwo0wgff29C
DlErrTzRN2NWSgXhGZRKBbWgWMfuvFpiHDJuwa3g/XUwMVzVgKpOHYjUuP+c
AWHAyn5tjNu6rqQSd05/0BLVGYMz6dDtICzY1NxvNZXfjoj2bDxMDq0wScUG
GX9hw5Y1UmTQiKGa6u6u46jddJRZ4ovHiiTbRna9zW5ljiatWx1MPKG9WBzu
lHjMDt/AGUXO4LJRM2uFzlclnpzLlvRrf5GZNOQoMil9fU3de0cKmOVcIPLk
h60lLP8OzecUXrllOKCzQP2r1WsAMcObfpThrxc0WAUt3eRTp0UYQVnxK8t4
8cskaOjxw4h9bP8yEHffA9zAr1RE36Ymn4HjkHT2bJ4jT5VbxJka0dRbFlf4
aFUHSFk3rLTrxgO6UZSnJSB8VEOeeqdy40402jzWFYRrzwahJo0O5SeIykdt
2GBGaUrXdEdh4WxcF1PILdSTLUNrKdXMcR5q9OgjDdCfCzQEyEkcDU8+DH1U
jxwrtpVLNfMDkt4B+9wWzsfhsqu0Aa+Wl66RO3/8WaWEdZiQy6+84kA2RLE0
VL4otUaZiRr5HRfbMQux0TtqS6Gn7IAkGagpDklJvikllg0CeUcl/RTrUH7R
Ed8otQ7ww65HGzoH4ZvqQdT9+ozMZ2BohAwo5i10oeQxCL+0ph/BDj0KkMor
Z9+dVM4rLhUtl697cDWbbly+l04jBWkxsDyG9R8p8INpK9JbooIBwQeKxIGc
sGi2cFJH4mNfDTTS/2i3YoIC6i81ml0AM5TU47vWHC03kpGMvKZ5NvMVXSwR
WgtjhHyoRPuPgHyRaGZ8ymUKtuHhhfuEUKFGPHLfvjz6RsTxgCYG779VSMvm
CSGx737IOzIpN1eARXvhgFHZjf6AsfFxctwU8Sje/l7BvhwQtVFPruTws0p6
eX+8BUedRTiihFvXv2wR7BeDoWIkyz5vUJ7ejIikFff8VXYTB3igh9PF4sUs
fNB1MIJ+idDYlCMQmz5GPctoHAOaURWvOGJFk+NCY/Two0PUXxb5vnf/v/om
eb6INZnb/JdSjEhT1w37lB6yxR5z+y3AGB8QeRwyREk90w3NpRpvAHTd70Ep
1ypSuLvzqmrYNETDI7ulRL7+0mc4XJShE/5wAh8bEOuoI9atj2dqJxO8upkg
uvM7r8pEWhrULwcLyBBRQUXQ+89qiG2yH/3eYPBnzp++T5jg7SAzvW7c4BW4
kr70h5t9s0qR/nCaEbCoHSQL7tNUretY6MiAQyZV1xrPVXIkqBkjR/z6fU7l
vxsDKBj88qeOMc8xLRRiD0YNmb52cl+Qpq9qDNaqz42NH87m8GzqkEHbHTQs
AP2WlOZBPI6AxmUGag2Hcr1aEIPqitvV5KIq9bIax4UQOyOCPdTJ6k5tvdhn
UZwg+/PSk87XV+WxFAOip+UMHBJeGy7RlF6/yjIYUNuc4pGqn3+fb5aXsPbf
3mKeYGAlK+q8xFlS8HqnLnPb0PijqM+1vdcvPXOENg9qvOB2id+bEEAuUdo5
rezc/9sow8lPtHolNWfscNgX4uCMJ4wErYhjnFRYyD1ot2W8uqkMZ10iq6YN
/RzHP9VUerKqc/afb/xSZ0jzwix/5JSsCUn5V/oD/J8YoWAn6nnLEkCksICd
D1t05XV+c6cn78wjEnkzYqXUr7O4HeP4TOID3IlQNiji8cY1ly1qZ9Rd+8sQ
RdLnSK00ky8U0KuRT6HJIGBDlzN45FKq5l95mnFmv79Dqem9ot8gO8Q9Pgb3
0mwAEvlgzenovEGEpCBhZ7ch8PuYw6KxosudV0lYjlggWOWN72VsR90UVZ7d
bcn1ZBq+hbfHOoZO6Ojk2Nbpdj6F/u3FFgr5t8tITmCfaAddi7QIf6Aj2TyQ
aIrvsG48q+9rO4NcbqDwPoQ0Yaz/wGPo3AKZ9HX6dts284xmao9sLiQ8ncuY
ikek4/Sp+7wNXEiUUF9Uegk+Z9x3JdKcg75FaeyPzF146TUzaX25w3VZrSJg
Fku1Zejl6ydjYw5GEroJeuSxPIqeXkIT/RhY3LLhiYEOqZ8OsVRp0HyHEbVh
w74UuWdKBS0DnpRwe3Ts2zo69pLw4HKnCh27rP/ZabHILIJPo9lW9l7oUEwp
OG1vQ9l8EPwepMyCR7InEz8/MtO/ImpA/Mc/r5OnSWV1ZDBfKpn7aRgVzYHr
dTFQH72gh3175Xiic7UEE1CqcGTMYTdqOuHltcebu2SaCG6Ns6Q3YyQhuMzR
TWyoyNLEzRdI8u3N1r6nTD0ECsiI9+khTVYaThEY+z4UUNVIZCriVXEJaoJz
y/PdtBkc21HA8wcNvKu1kVLk2aLMacehF92bqWHZdEcLZGFah+q7xy+2+ovy
LmA13gv6iHko+V/qPkXNcKY5lnstZU2iiQ7oJm4lfGa1ellDnOloa0Xn3r1C
vzID+G7tVbBpMql3b7xlCtIwOSEY+MLVK9tRIO8vkCjX1UOt1gI15AUteBOQ
9rRxwaHo5pMy9vFdf7CLrEYLTI5ETLxBovgy6Ktly/an3Q172dNNEuGo/1xO
wpuXs7ALZaNXSkAnquI4CMG/12o2KjeQPx2uGd34w9Jzg84HTa1HqeIbKf8Q
jnsRcvoW8ZSzuWxkS/VeCe73oPQh+kKLJclRD7h4A0ITzoYgwClFLIcAuqpv
TVNMWnDRkeE3reyr0bXvAPmkXvjSl2WUG26KFv7oDH/R/v9B18JxfMz7iml2
4iqRqQ14GtGEeF0kFsiHv9ZT9nRWt+08Wuyu45GF0RK9c3Yh4X7VcGuDE/W3
Xhias39bsstzVaVziDeEzr163h/64DUHgw7U8l7A6B6Yira750v5QBVTv486
eSiQ6ZiobuN2TsJidaaHpNJ2KNmrZEimYiB6yB4YdqkwEi7nFPdmT2QQEVZi
GxQGJ16945L7cWWRv1/UjmIYuEgpSImpSpaXJl9wReem+GQwVHkMHjygqMZk
liWjarsDiJ+CugVCe6AHPJJ/Xfz/vmZK+/dR6s5VeT3AFNUZAgforVqjPXwS
7pFL/5+n+AnGjNKMij9YU2d6qeUMmpESG+36mbPF/jRtbSxwDnzNKOEoqvAh
d9nRCZ7NOeHvtzVTo8d6OCrmAdLbF5DfYViqlK1eHgFfNnZHb5OMjN1KwABm
ZWVb3Cc/nPaWlIm4Q/0wusW82N5pBnk+7umkhskqfoDa+AQ6egfraAUhyxVs
UrcXo0f1VYraoYql2lVqSJClJKFZZWHRmeaIfWxcW/RrTBd+9WeatwE7lje3
9TmJ3hrP9wHWRApXY3zwl3BU5Lims19lAvqrEV+z600Mk+CC6hO43U9nfnnI
sPPLAb93HCC5qLBV1wh+cWWvcJOjp8QhBUrJ+DqOJHScx51J4Ihj0B4ta/HV
rU/BR55SW5wDh88GD5NLV4M+tGXoDEjq1LFGQGN/mTyR7pKXCYf5fxgoXFeL
tU7tYAgjhkvqqrsWHGAWLImBCwQaJFPL+zpT6hj+6jkzonhsG6Lf0KHD1pEg
Gi84ISgh+OJTyeZxO8zUMHpn6sEIFbkQaLoCqFFi6UWfLkZoJGExqetof9BW
tb+AKIt3hBsJyugwC3U4dDzIHRuLTv5zGLEioMT9DgRJrD6XRPPGaGk+0O6Q
ruZxkNHfakCtr8RSEipT+j8LET6DlSrIFcE24sd+uezm5ymtNybLYLTcVuUW
vtzY2qVPNf00DnH3HvdUy7VA1z4PVlSX+FqySA7aBNMes3YF2Da+zPU9PK2Z
iRdf83jKd54+zqBzw4p/tT+WN5ITofgZduLZe8sUQyg2fDiImN6j4hexvQgM
5am5iQXfvSBj4UwME6kbgyBwwKfjG7P8GFhhJSsfaK0RvlZBzUyxwJqTGjV8
XsaeU2IYkS6MCuOd74nhRFJLkdgyNJYOUvzKFnZOB0xiPjsrug5B0es8wdFm
YJ5beg/Qy/rNyNgIzToCOzlxLg/2Nruu0GKEyqlEGyOvuZfvB7iAMWiId+Bs
uGmsXPRoCaCAn1nsBsPzYGl2b1LKuwcoabDXq14ZWm4YkIo+F6CD4QNs0Met
17aqXix8EisJoPNTX1PsJVfb7IlIfv2YTBHXzJl5vwipCN0rlbLVGP1MuMg5
Miqn15az8YEf8DLfkWkqPC+yVjBCd/bTUKtgkttswHJ8CJd5VeV+CKpjS2H4
rh9B+7txE2ee/FY4hpssD8iw/eW0ACivwQUYd/SK86qcSKXp8Dc/SQf7mL5x
Pks8ybX32WjrSP2EqLSppWznwFpf4HpI2tbE+xMcwJ7DWByRPP7TMFovmzQc
oyUAs/7+i155kgtsQw+S/tGoAlhGIrJTnKaeEzfMnzzmRJl8hWAibY2WCSU5
KZx+PkFdCzSgrYx2PafCYaL6scnuXwW3C1lY8uwDtowF8AsMFpjhhrvJoYLI
cd9MTcvd1oW2I2fpTTX3okEcSQZMU0N6Ta7/CJKxa5nkyjIPBoTYYnWVE+f2
LvJrVBgNOUUK0fZWpgzJ8mRCVRSAjl271BQmkMKZ0uCyadxn00QihtCaQiXm
Po0uEvU0W2ovTYww0LRnxYLCP9So/p/YMzGx26WLygldqL/RxdPII0PomwAZ
UBSW8ReMyDH0ZGm0Jwk2rJiSFS1ZpfvD360itzcrOeCmVpvEXePDnodnvArX
J0R1k0MoAFp1fVRhZxlrumYz0zRReq0m19fOQDytoAQED+7mBupr7o8H5B0U
/kAjGiKLyA60zHx7p1VZ6Vn8bMprY3vGo/jMBQP5qotF5l8DHCqcPLQAiBpP
ahZHMGZYINWBvvxcnguKpQIwFJ0Ry4B+JM049dFRHlgBVByPo7+YZkZYCg6O
3OIYrre97V37ZaXbhmpxsJLKuklCv7xkkOriyOksrTBZ8LwG8FsXpo1dPmdQ
kkDlXPfEfHQxLMbI5wYDB7whGiuY7+7cU2mAqHzhXNCZ5GwBOpxekb7l0Nb2
5Eq9IObSeW1u94fn3n8P8Ggu5jIQ+gAqcln698mWdsd4VDBf0nOmW8eHV+Kn
ZjOS/en0fZ0F+bmAdfZ1dz9n3HsEqlYxOcrNEk3+/ws09XPZ1OngmaQGKoyD
sVXxSDtQhZuorWa/TIqBUkerhI6RIoqzFvAr0svkteUROyOD8xDwLanYofgR
GQrZqufXxC14m8fKE1h4lnEKq/QySdLDyn5IwL75aed/SxWrT+/79Mmu28eM
wsc9bZ3r0Wzz5Zk7epw5zvka+j8Fhz3gtbkLI6qjDefpNL5tT/Z/q7U59/jL
z3IYWjFNUTt39m+lp6vfXoqFftm5w9ca01xZIuXW93MusEday4J2tONWIIAB
WHOTEgZh7kFUQQ64Ieb7rmN8NG3lXnhvEK+A0LCYgDG52ns6M078qImt7wWV
akXszRwNvr+6GERo8neqm6cLl9j+4Bhz16jsPCy7bQNJZLa3+ECyYmFN1Vz3
MW4ecut8xKwTj5XQ0cZRNzxdRXGYIo2Z79BCdL785s/TfIhEDH9aVhhlDzL+
Hoe7HgtqsTF622HOkFa4w4vLk367EEn3UW5CeLKa1sRu7qhjomnI6phaKZtZ
u3qiTqulOrN2WgpmKi1jPw7omAPMfeTieU8Mo6Bh4fnInWW/4V/Qak7NIo/D
meGvItTIryYmKVsvxfqBBQd62imMtsCrzaNUml7+yYcRaI/NyfSA3aks5/64
x2OVeeAL69wxenHszPAANSaTAMr7dY/7DWjuk6/RauTGHCoWYSrahCj2jBb4
+qbhUj0q9VxobKBhQNVCTWXwwtGzEmhLwkYyAPy6I5gGirM7Xke1hVAYIcXF
5bQdD/tYLV7GGhgFpAENXA1MmpOXgacxbSvtiD7avZ/h6d+s/hYuN7LB05lA
CksoTm77w1UAIbnCorMmSDkPCTq0d1xUzb/TqwK8BpCz7ypbgXralY/bY7po
3wLJaP/a0CX/KgByOBfbl5LuK4PupiPPQRomTcXY2TxDPR3cbSujoS3eNU9e
ByFHt5P5oTpbI55zNKnrVagW4tRPScjcs5M8oSRa4Rhf0zx5XrRlYoNGjB1v
+eWFddzyk5E/RzYk6VcuemHoRm0bQY43ssZpg0YeqbaK5eI5s3jia+JBYNDZ
lP/jWutTPJGR4tFf41XWZORX3pjDdOvJuXMhfxSdkGxgbCJ4RyLD+nRMj5HA
OSOhYrCQoeJEytIFUlKsxdEsJK2RYCXZ5hPMsP2+xvJQa9aaXD1131zHjQQu
al97irv1MSwYzCuRQIPFANMttRun2ypB8R0/oheO8e7FRDy8gECPTp9+s3bt
YiZ32N+Akk8rb3aCU8m4nEy72/fNCFL8OMHwEp7cvpUnpmiszWirSs1Fqi2V
/GGSp7VBrdGY0JwyFlA9NPV6MbjhHyhnBDCWvRWHLmtWYnGEJJH7E2GtnC8h
vAVmoqx0cpQvObsJ59iA3f5TEy66NUF8htGtQdb4BJOVja4QVJZZom0mmvke
ds9HOhHzWiBG4UY3K0bQkOnC0p/jcJ2tyC+1UFuK4dK+yjM7r73bnUIOVfGy
T9A+wLIy2sCQ8qM/taEpRGgP+8+419zNUEPTs53JIlbNOg7bsyKetQYacwlX
IM/4Def2FCMpdzvH6tuPZtfBFnGBddcUSo8C0FGTI9OzORar1+iMuSLfkXED
ayKBHFyqprsH/c+OSNB5Np5fDPu8/Kwhbi+cyVA96OXKVGQwgRTvomSvIuMy
XsXwarFoZRVIxmFqsXRT0J9fa0CIsnP2pEODWUMWlZksaGDGbVf/nD3oaW+3
9LwR/vYl1zrE56TelyBN0Iv6CfwlydvHrt8VWa+zwqLIPLpuAwcmIw67+9kN
NKkEusUZpn9nNS2VGcF3935Jqf7oxNyEBlFZ5QUuKcXkSd6x7us8rBc7nonH
RXbxsgB1mf/S/bEcMh57h6cTR1luKDUqK+UQQTEYiCzc5zfFYwkBcZGb0Mi3
FxdEYIRNFwIKCd6ThPony5DliZLZPcscI0JuJF/DMY0gvzrmuba9ZLl+Uolz
vlnns5e7FNz2m30j9Ld8iP3Lb/NLXKItGTNqzZh+o+CKEn9EqLiTHtIc+Kf+
qngwy1iNsmjMjHiISCXdfQ6VQvhREVIkum/P1IueghoWnYw+E3fGhqDnkTUz
9eafNgpwh4PXFuDpBC2/msvrfAFu1XEVGgsm1qeG0IoWVJkrgRTJdusx2qMm
ATQLACL4s4Qmaxg6TRmKL4gkh+YpPSxrYm4fo89fjauNyPg/hYcWk60w8tpu
U+xiv44q1EUtJmCfBiL12jEBe6wAUU1GmuMk/g/rY231Aelc258BlztVOGND
a83vxsnW0JCz1tTl+3Gfmw41/LhezQcIwSH3h6A2Mt8Bl3s0PA5xUTWeAZnB
bJDrX2axdRQNgnq2gt9+s1ZuE6te54nl89cil79AqJyv8GqMlm72bNyZOXZj
2lB4IZm/Uw8QhbZ1iGAHLQszNXWtu1flPDqyJx09oynzr2WSOcZe8oLUEx2p
jc2rTTl42+M6M1xK6vopNyGloFtdxHCaR5bsNZmVa2Q1Uf1rZRNL95nzlBDZ
NoYkSb4UN0Lr/bYHJ5chUqHHBBl0lVxKldU4vknhcFSAodnimiCQvK0UBE3Y
29bx5BLN4Q758rXKeAZKkaLCsB8IS4HJcmhFGHynAp9jw14BjAn/fhOMW4tJ
zk3S+RaaAtKk/hIBgSIswiJ1uzJ4AnL/eg9LAM3P+VYCL6N6aV/VXnw9Qfi6
9wx4P0ikOfO16HZ0RfLUFis/lMl/zdcejITbM3wB1xhfCsRvfTLYxq9OjLym
KsA3G/JyHmzJ7/7fqH8sjzuFJCkhVfCHtEGNd2dz7hSnBVLET0cqbGlj6ChI
8k0iJaTjYB9bEGqzyK+wF0h2cRfzgFFAu5zfA4tk4iQPowFhL/SERVsQ5MxS
LSh3/xzoMg0qxJjxNOxcQunbQnUeMBRzwzqSUwPQMXQEFOvTug94lzo4S9cD
5pSGieymaJEYfqtk4FpfrBHWpPTEUBcGsO80lMzLwIXdlX7XD/XigIqi6ik6
bmi540PiXJzhvjYuaPJHf1HYn37AyvJbItXYrfM71Z/UywoufUqU+iFkW3EP
kcUS3RgO2xjJ4O0S/xznoZ4c9vnOnDWhhLKyg/A84a9SVKb2WM96hPqOLzSa
QgrmnAtvjjGpzs3e2PcU++2Gi4Miu39yO0ELq2/TXY53CKJq4X2QooCs6GTS
2Hh9P7W1NfsZ34DoYlv9MliDQSEzzaRLdvtS2Iy/bhZlweW3vHwc1drGYDM1
UgERszEoSOP0VEh5s0F0mLVAR1EXnDIO34YSA8Dser5TccwSkGPhu9eb4dD0
5Qe1lbW89VyGZjfQBOydlK6pYxdsL7HjuxxK7Pjej77GmYkKxAsS2ToYvlpY
xvGrAtD/UK8qoQIJD0uU3Vr7tBsZqfqqEeiacXbC9SRa28sm5ua77dbk6V0W
bsVJ+WEDTuI9i9jKjP8/246PWMdUFS6dlnsy+IpCLzUuVuJzsk5A6iCCHRdm
jrYlR7GmRx2C/kUIkoUAleIfS1HiXSbjee0wx0mu6ePwbVYp+Qub2uRRIdHE
q8/fo+CzuAmT01gZUyC4Hq+ydDihB7yqSerKh6IYnbsv11am/HJCJ9+cribN
MRRC5lYP+ZiOFs/JgaR9NbWUfnW9Aa+vD75afP1eZBQPl2uxhKXW1dkadN3/
O1uCx/Tw/GXo/0BOugIqZj7H2vuzh9k+FgsKbvOUm1QdnPP+9BDpRCDISgjZ
opYejyh5OsOh1jCVEGZ3+xTYga7UPoPAZwC1KRwsmmfP86ybntvjT4EWAQeM
UNe4Z0jDCDabeqjbmfSqZrdmWq2PZnBjB8QrpqWoEBxOwegMcHSYQ9xn13AB
L49nco3QRudOMy+KcH98wwJrM3l4lTqH6UPVFQU1V5hW1OKrKP/E2GDdeiuW
0zbucF0t7GcJTW7tpVhppGKlI7aBaXEMVWip5jVwyq/Sai/Q2WwDkkdN01YC
D0blO32Br7f2FrG3XcRPe2VOVSlO8vii7SAeG/z9eNnk2EdvMWpaYym8MmPm
bG/cnsZypZwQezF10XnVw+uY1lA+fQ0ycCgLxVZyI6P1c9tTUs4RbhyTNKf/
PL1aCXqTvffxuVJv5SZW3MUEyaqOspGVgKFXc11BsPp+f8MfN3Ia6AyFW12v
W961i/7OdIbMzymBNCUYKdypwLcVU8MP0u63wh5qz2IpZ+uUcUay8YlYx3hT
phjbxjVXOTy5YwubyYkqBUgO84rhGDCySBkg+ynwlByGnDEB5AdTfET6kIDp
SUyQMAWphQ7q7KSUPYqoAjp8p3ScBtJLbEIljO9fFWuDO46v9fufOQaP+wE1
2wobeYlj2ghsDhAH2BZ70KXjyVVDqtFiAI0ynU4dXI5cun+CpMIiazDc/sfc
gaUQM4eWI6GVRb1RFkcOCC3+MUZzGBn+iQrG+nMgoFI3HOlTTecgxFlruyzI
ByL3Eq3c2bMYufEtbKjqIVyUwVpgyEj7fsFBAYiX1trNnUh6iJhortSZgcya
2gue+QLaNr6WTwPu1uitoGJmh3xP1Vdq77PpPRM5KXdvYsFxQa3HMtRcsnWg
rRsMb7FvrX+eu63XuusjvcyqWtIZ/vMrRKSQsxhYMLuDgKGuIajphKQ5UlQk
5qqvBi750GJK0AtSluiIhCjVITJiwBCM3ZPNu+ETWt/Moz5e5kUDWrS51vFV
atPKi0TJ4GO1GKIK2S7LqIG8SEoUWA78eERKkHF25pW3chJr1N/JF9SsnAGE
fHc+xiPzjUqltlO3eBbETqNQu7n8tTgbR4Qa5s6nzSjrmj0R+ish8KQpry9r
Ng2FQtD07dEXIVlc/m8K4pS63198goCTNofILYEu2IIwyAbZGWwWrdtuE0tj
vG4xjxPWZH4nGP2E7nCcKZNLOZN79r2ZA/qcr6lAGznrBaCls2FDhpqoaXNa
cpVQU9EDDuzVgH0yMq6yWKTxunLZ1g2a7NlJRDQ1lPVYhiQ1R75nIPn0dQeW
ZL8NExviR+VwWE9wAyPKDvkUO0YAEloKG6RXkGmjEHHHj3r8BbQSKDWMBKyo
cfbBO33st62OHGnzuKFUJqwVIEF0q80SiPZ152y4PwLwypUVv9zuhn0SEjYD
PfCPcDK5Y/P4LJqJusFpEmpzn3OxD/ad398/qR1heKEaUJD9ikGg5Mk7lTba
QjHikTorMoHks4r1dGVPWyHWTnPExhHlIhadWaS+25gYeLaW15q/0r0Ph97J
hOo8PtDa56of0F6h7rswrb7aHlOJneXWKlMIrrIyIitD0cYDKYyzuD1lwkL/
L1fYQapdzM1aNgTWN8cGkEsG94QzzG7RM4/oQ7rZA4FBUtPsR+bnEmxmBahN
g37y4mGDjLS2s+jwmXO+5DRVI8APs6BfXpn0EycmHQvjR8g3xvnCQulqOlDT
vg4D+bILx/kJ6j/nZA/b7pY4SIU+vFRrYstMPSH4b3AzSPl2LIWrXdCSxJC1
x0Vk27sJz+htStRqqiOGjfB5KPk+cp5kFDy1xusXkGk9RV0PSuY6X+b6TH3Y
CUwR0jLWI+CEpBkMST3V+Y7fuChI5IrojH03ZnTCsejtM6Qvg1ZYUhDzMPsq
hKLbzlhkhLIRyLqLEQM+vl3/nz2WFW8baXcDMGwX6Belk0QzH8eJ9C5O4eJp
TrBnSc1FkAHgxJ+w9KddCD3KzfJbEM0JhYbN6Y7xi9tq+c/FBMjqfl5wExmd
ZgEEApww1ZXnSMFbNimiaeaSJiWDL4D2/NybWimR3iYygIa8T4aS57TQ60Hg
Agitsw9Xw8P1y23wu1o4oMkHiGnQdym80gr3uQxo7OZ0+eOvbamavYHsisFK
wTT8SY/Cw4dn+HZOWv46n6movsUAjcmL/NF2usbtVpBle/19uINp1K+bD5Y8
Nzgk0/njj05Adtk0D7Ny3aC2TL8UnIOqKo8s1GHzkbszgQBmgpA8eDLMreOO
lCAxNkOy5A4dOrp0+kZYTCV0LZpwOJqKHhsTywedVHnBVeDQRZAjvGLjMyBc
AX17QpeF5i01UKItgLbwAbx8F2y2/ChZYnlkn/6daPupF4/8sj9cLQE5+JNk
UlPcMAqetYDvTJdnMRXZSe5LaQ5oQEUs7Nb9uNVOlD5Ks15JaB00yWTcNYWS
plkfZTNcCfadnx3c4lrZIQKnzK6u+qhzd2Bn+q6vwcUQumq6EBAJMaAH0bc+
Oc00X03R0VQn4nu8T7cEL+uPzWHd9m792Cw1gmwcPm4UhVrxKzIlM3UKeWua
qtHZ6hzQw2FOFl9gWGBJXaIkDkq2t6r9oWjNyaYC/tS4VYy2UPLzjUdm+l44
b4W0seBBBYLOFWNCObpnOaZ9e5y49//DOrj/AtMWNwovQGQ+wGTY4SPLiHJZ
Aefw9RCiUOBW1jAIGwPXaoGvVUo2385uQXcBeQuTqX2kzslQM6seRD+Q61g3
qB7d3+FhPCgOzVt3GqjuLYyYYQZ2eh4ETfRpzBSu5PGx+tG69kd1VIHqmSJQ
20+qLKiNLRIMXCh6vnCCcTX++44lIiQdixggZj0a5NUzLvFiNdVcpnNjGNbb
k0yfUIerD4t1I5gV51xtGhMsWHZBHYyuMpBW7vCU2WhlwJSS4SrauGy8M/l3
ZSRklMG6aNXCdXkgZg+5nPf/Oa9pwXJjj1VS3f4PObDlSgyL2K8B7WtLyF3g
wHw0w2qP7eWBpq8D2hs7s/RWCxDvpndhrhluF/n+mmgYck1s49X8Rymuok0S
2oxWrJ9FyDciQXgor7xq0BdOgFd6gC8skNMJZYKbYbpbo3TZ0YPOhppSm5is
2OLf/aNsOjFededQw0Jn476VYtiBQ6XYFiFjgP3dxuDngr1SSznYOodHb1iK
Rml3Ek5KEKRpvyRyJ5nKb2RPY+PAp9CABo5r+PTI2fq4NsgWCvfiVBt+4f8K
XFltq4McrsesiFRDcB3j3E8F4Kyk9SS1ruca3zzAwqF4EMFVJvkSL/bLW7NM
b+euK99meoHeKZBK99P12v4qVdCQDudXbokyStpJYO03AMGGRMWQXM/D8dJP
Tdls1QpCyQU7RPAJkQ3GWEA6DbSIvmNGEcwfkORTBPZXFxB5zgniUJAC/vdQ
GXumeLLzwnLUKfuO1632YmR7cx/USf/TPRq0no+h5imtKNuFqa6s3uKR3O2H
NVwWBIgUmjQoJNcm+Ogv26yNO6iuhimUYRtGLSKSkIcjEi9yV6BsttU7AkQA
DxeILH3rhrwOC0FR5lts9E7iKE+jQ7+VDzL4pLHcIAd3MbnqA/7ZLyCS+QG5
56+nMshX812VJcgh63Y3dXses0J5ugakKLrSC1QVe1ebrcgjJFmjYMs7a3G4
bNaX9t+LBrELkkWnVgcPTY17hSlXiiRnVclFDrH2bqNPisQyGqRChe245mMx
QJHjB8GM2ls93mTap0nLKpYM4jXV/HjpDkx75WoGEbWfhpU0wUxIS8GIYPyM
HwNojaulpCculL+saQhG0NN/5aE0wZpPS/2whvHuIQxwOY5tOlxC2m3lIjZw
ShBngPixSZYVWIh+oZJdZ3IEfiOck7XlGlEvZ/Jkp/akGZrpx6GnqVJ40ILH
FNdWEw1erwT89PvWrtwRoY8gXTIYXRshgUTY/byJWFyO6BwdNMtKvSdgluFs
BktRK6+4st72uUa1anRrmdrpYRlUmsL0RS9FvTKOTWwN8hfaOO4AzHyE8KCH
57Vfeursit78Baorusue2f/F90wkOUGKXTvJN23SCKReLYzGbCLlBcbWXXce
XRsAbK54ifVAFrBj0774pMNGtTZKuanDE/564sSYNAu42+o35UEpVKlbAPjs
pJ3rJyD7EUxdD0m6HaTzrX9JS4RtiBz+kV0+nezhjGEPsijhXkxwK5a+qTSI
9iBDSPmj3ZAB4WF3FndUtpyAys+TGy3ezq4sOoQlpUhJunzP2AxLZ8nla0MG
u6X9LpRSI+TVCi7duzxyDVK0wWNFcQJ+upNFgduQ7s/ZojhVc07+HFlvkWqz
2QwFR4HfEU8+ktJUUCla83xLTF1Y7c71IHUJ808wZuP9vFFZwgHpTOCi3oCS
DbIgZh4Tu8GE5XKMGCrCEX0SoA1WxAjMXw2kKgOX9q2z1OMkjsdjbO1qZ2or
L1orpbXFfG6q6M0I3NU9YGjdjjiqHqQXEWz2UIJDp537ivm6MJPO56BgSSOJ
vnOlhqigu4Zt0TOvo4Behy4EhQcROU+/oa8y+iO1nIsSV21YIHL3gkywdZge
oWAbUHC9GGRL0EGRcwZE5SS+zEh2Xm5mcyOTNFt3PesUsNvGPQYhqL//OpfY
97XeT+sEXYULo7xpPalwxRgcQWVa6ClDXg8g0Waiw1eDgfFY68xL6eIButtt
CbGWkNVrrEjs/yCGMJJoEFV0axtgRoe43wyiPYDZfZTdEYm2TVWTUge/zB0E
SxVUbrdC2Cb9RDTORQm91UvWpp9yMvnWQR9Prz9mBZLjDtbgQn2+JAmnaw04
iTHadtZ0/9PlzOOcW32Yto9uO+doaTdlssN9pZ5mo/1CU/WIPHxZDg43PwTd
8JJqO2UalvXPszoMWpzHjonDBYjEGVr05EdyExJLnjNYN2PKFGyNIlc53a3L
dQy0KkhVSiOCFYzhi61GA1WOSTzv3OHGvRn1IgzEcyvDGW3WeQF94nGYwChB
4Us35o1S+TOt1PU4BNxSqh9UNGmZWPOR4nRyO0uJVg3tqMsjHR+L5JH0kjTE
XtsmZkguwMo5xv9GFHiV0hUVd/Beu+ikfKXlvLYasxrTshlw2fOZFIdiX75p
4MiLMl5pwB38iy879/+wVRVJhPtZubaTXa0lP1NGIZCDeU4/dBgf4v2k5Ko1
WHPnHvtY4NLBeFlcEeuu3sBdtKVIwdfr3ATlw3loBuM/26UFi7J3MFaArXdd
NxZxqMVEk6uENbLlUn5SpBTXifJ4NlELjK8Q3lRKJoRY2hPlRq/0FFm70W+i
MwI3FSs0RUtRwH8qYxS+o+tQr9LRvnLJdPFlRRIY435VihjZCrdjMLN7Gpmx
EvKb+cBheHg+kv+BdyDmZzjdrxe/oOt2cr2Dt7IuiZMbCTZ2/f6rwmKrkQ5T
A8h/Oq0O/lnoHiSz3EoZ9I/QSLhwOf05wVVseNXT93g7BpW7+DXvBUrhg/Ap
c0UPF/EN7tCWJNUeIRM2c8ey9kfUVclZSo/vdY8ZXh9McCVNgAjzt3SKT+zr
RmKxbGPcGXdnk1ioaLQeB6UUQMieXnJxcmS2jwxzoSXQ8rhLXSkv9JLe2pXz
l6gAk1RcknrgZ90kR70oYTikRrgwioEAfQA1fm1s2fTJCYTv18pJ9aFIccab
e3UbNdgiM8Uli9qfaAISVZHSRiN5Oapww8gUdfc5QmIXqod4LxlPvEsBfCf5
gmj9j5YD2TJABO7zGR4JHgx9AQffKpe+sB+aME4v9mSVuK9ujXVXyYkF2gB6
GxzqU+fzDbnPRmF2J5moWgj72iVNt+lw7rANrEnmqIjlypfpy+lgWhUZPz23
8kc39AcojCM+9VnhP3oC90pecqVF3fwvwQ9kuTYCNMpDMmVIh5T7iH+upM7Y
KD4Pl/GynuD7FekrdIvhXDX23E3as4qbbo89GkQxPyNB+Ggz0YNx6V3g03Gv
vbb38lrjmBkbEgTTknJ7z21rRlE+GNAIifFEkedIqioYO0cpml78Pg2HOGwn
OQO5g07Jd/i+R2Z0k1HmjO0yOamUcfuipSI4TcUGfuX2StsMyO/2WHkQk1zq
DCSyvO0SgcYCGQRGHbFbyF0PfyPvof6+YLPtVYFeVLkBbgOT/hAcePi0Yuno
0NJDEnmM6wUjEF5crxN5JwvcAeTPw/qhjD6oIu665ATAnz/2ofkmx3qAQz+d
Ng+qyF7Tnom14iqQZzcvRFF+Vz74Z9ZsLNidMZtQ17eXTmM5AJjDgdoNjAmC
SK/jgBc6eDsrR0ae0RVAUKgWlmPuYeqWGQJHE/qgVbKHrzjpQ8APneC78arF
BuzdDybKfhUA2lJdzbu8Qaf2qhYoojlov8dEXtzERyPwSAxogvemo04QkRth
Kh/hoU4eofkQU6aY37YHjLBHqg1BcKc0nfUm/qCwPYntkkAla9CIlhyIYVYo
pn8SDF/ZoYIt/5CPMUUz7fPp6N8AI3qlx+EhaGp/M+SncakEslXbSqptudcg
ARkEktM+iGihai4MXhOT1qfXHin426lGLFqna80QgJ3bIyGkjQqzTboW5+IC
KyMlNueRZ4PaUPI5HpoWp3+gBf8rplDTvpw6l1BsWjc+62Z4m0jupSX0/iwe
eDqlH6f3c/jMncSnv+xn7XlRGvqZah4jPn3ubuuXsWoodc9KHyvxt/W/0oyk
zDjpKYyUMmPnrexIyKq/TJ4nB6R5ryvMZuv7tF/YR0fy0LqBGmM4VOQJMEk5
NNcHMYNX9jGzU8w2NOk2rIXzRCI4A4fpBRVzM+3qxY2khSzBTfFH5S9CmcZX
RQjLuj6rrN0YWEY3llKJp4ztPuJ5558cKsZvaYRD9EksmUbCLSQeX6Bk+a6H
E1/qopWwDOzt5GjStWbWsQqgj4MmWM4kha9TYenZY7tyBgTK8WMHWYVxsODK
DSsSA4dvIUx6rA9mF7LPNBVscxRVW0EKriNgUxJ/K134dFcLzDvpjiYfzm1e
7k02llydWZLX2tFqEjcxL8qm72mBQLqaAXQ+SOYZ8NmRGE2thBgqRKV2J1X4
XZQl7DEmKvzJObxw5Q8x9km4pDi6WQytgSmVhn5LONsraLplD17ssPnSEUPo
tvO2uDoQO8M7d2a9M/A8n/HQwfFvdHnRmDZevldekquOqkw8obibeck5UlF1
5ZDZACs6OxPUiovqWAfcsZteiLspYBQ78V6h465+/hqhFBjUt29UD6TjhduM
spE/j6KG2OBXe5z8eA+Zcr1s7kftQ0eKnB0CXW5AYdJsPvykMpm1VruzOeix
9fy2XPdWj4KA5U8BtAFJIP+9UnM2P+E7/mJQR8fgZz+4unJ161/rPw2OWObM
0sMWrEq9gA8/+b6pHEgEuyFsAdwwhaKldsU5/qwkwLXhKeDzHk6suCHCeFHC
90lWT7iKZKZi/bmTz8/KxYdoDqysZQkk/L2mMA3nftLgEW/mn2f4czX11cPf
zsou7HyWDUmpJ1BJ3SGv2ESMQaRa7+V+DXsvyXzheEnCOkYrMgDL/aML/07e
XmtA/nZLDX+L81k8+Pe4njG4W35ZPWc0a6FlPwTAgX/KuYhZwmYg/vR7R1wj
/KK0Z/3TN2BOHBpE0A3HcbXk6irN0/GTL9is4dPVZyJCX/EUKJw9K5okfpnP
UDKzPT59OagYxeTBHsmJZq0NzOuBGNcuAZgzrwS17oSoqiW7TE0rUk4TOR+K
is2JlRJ4aY2aHdrOHrX8W2JtgIInwrUGBgSviiwVT24AWPJ8hzBBSYtlHnej
5rpmBDwqWGZeFAMoAy2ze/2lTKwXX7ZsSh0gdxv/zGei5pqzKAF1Hwl1KIGe
qCU5tNrd9U6GSNVjHWAWsw30F7Gd/eDs3AujDaP08kX/6n1k/4PbH4+03Hfd
wWRNbi1qCElOmULr80TT4Oytg4ll8eQxuXjac9t+re8BDfxLfxQzB80Mb4Vv
8j9aar1TLp1JJRy5sT4r7mXUZHLj8BfzsHz2jrO65+dolkZ5ZgbAy4nk47EP
ZSu+oCUF3GyhaJa+mGFBFbsmv5zEOtwGhaxWQVOD0dPPFQWejtYOZkubB3HL
PQk96UVBmkxTp3D7s773B7DO5phPvzjZaap2nXBqCmeaJAcQnwQH0ks1CvpV
tqRsYabjyuHU0KIZIP6AHwhklDoFKeBTjKvCOosZAhUvetNSxXzBCzDr4uY7
YpVlz5R8VKm0wtb/DnLB8bs9o5qaWaAOpdvj41c8vAFwCBiGv/Ac279nXNcW
YCpwyXc8ZdcU4iTi0m+FRl7i6Bz0WjPtnHdnr91om7yXpwSQaqJ7Wm4diRPW
CgIOlAbuYUjKlLJdsPvcNzegQdm70uZXiyhsWpNC/k0dR9Y7eOcf2TNDFBJw
6TThf4+BR22PW2hlQ4SQXUTsvODyJBkLNoPk5Rl724f530MW02Ps+9i+nFoB
O1R4TvG+VrLCapoLLkYwUBP7rnHnlp18KVT77dw1o6p1qG+u+cMK29767m9w
6PvueNrZZFD3qdvv//vE570veCGwAYJP/feAFJAA7HFDTpVjfQI84er4Trij
jFWTV+Dg0pdREbqgJaY6/gkLGmU+urxZcuoGFssEvmH3MV6mo+oEsKkSRZg8
zIoT75VXE0fFoxqqlTNrJtaePPguRbVQoIWTSoG0exONuP2sYZfzBNvpZD+4
jJvd7XomJm1+NHw7KwLXrup5gmEQM4ij6hVAqXHXnVhPwaseVrxaDbGSgJkP
nfHjAculqCD/YuFo+xBQl2JP2iA6NvNHIehM71wgzt0YXo5mpQyyc4gEidBw
JJgvOdGu1Ti28AjX5AafUBsB5eZb3lca9IlqSztvCMJaLBs3cmK5PzOBy8Bt
Pa8gXEvv13XOhm4InkObmHO964TneUt3yz8DOd5uvQ51z3egaEIQZFWBKx5q
PQryijDCCBnSi1ccmQrk8oLZG/m4F8vjc74+aF3sqcwb6eRiL0quegJ67koE
EWrvXIo9G56nGFpZh7BEcAY5X/yDbZ+5ffF7DnNf1aI1/10DP+kDuZV8BU+O
NPDQ6Ger2EwCbJdaWaUHjor8CX4YppK6MxPu0W3Bd3yhi/+MSiK9NHyld8Tm
amoy+FuzhQG03HBPtfYPciclmoWQHmbZQj389Wu6ZM6L/a4mTJKjaDXd6Fsv
+b+G0rqsGVV6Wv57lANxRAd4MF4ppQyrQhRPUgVxleE2PJE8Y3EhF6shKzoc
g45StF0+GBUq/P6pkZVzNxQAdFXWz1dhVmoT23AtVUSkzZVvElQH5ghRUvzI
O908PCpKvKLEoMxHkiOpAvqacan4MsnDCu5W04I9NPjlaBHv5/WlLx6+r5uu
Vc66G2sSzfewykTNzFDAiRpkewir1aLedwEu65QyI0Fr1rzxxFxGh82nyKP9
G1Mci9xDUAKRGkvL18JjLMCaG9rXUqsa0Se+VChaXYgNh6+SmEIINlIjrL3C
9IH2i5kD69b3ZOjLHHevaLDP6J/xHfjQob7Nv3FSnPaj/1D+sLCC+1UhrEKD
BiKXTu6GBWOWND3ZnTc6SaR2T05iegJJkQRNZoRxklsGPtzvzrWuGRG1Rkuk
M7nlMPS3G75IgtkCgHTwH5Zh0yb7dJFfvhajM5qHAOs7Gb1kNTFhDcLdjKsy
pcixYf/zafnh6cWY8E7FZydvU1bNaOxZmeV3yWdP/0fM6MuYkGswpZ4y/ljv
hzoUzCOxbRb3dPkPy9eAcXNX6nsz9DyUFN6PNR6TRgaBjoDOFuhr0ep/EeZW
kf9spYQH0mcePcyXANjzF/pdxrK0sC4lEWCQveM5EXk1Dcd48bIHlFrAwx55
GRxkUWRpcwd3q6NjF3MF+ihLU7edizOjMG2ZkfUrqs43mmIvH4FvBKc2KdYm
QhN74fyN6MJ2YkHO9D2SldBcR5d8Wim8LgCau6unaqEej7B2ID2SvR6Lj0i0
xCAuvWE3eWmv8FKDnbJ+1qXMscyRLsu+YCUX5E1hpk6sWWvvb3T6eeGjoI7q
jXn69nU9B+SjxDE4s6Qi8w7STcp0VUHE6EjjIASSGm4NQp5dfBj/KM8NO/nW
PtzjOeE5rA6cZhsC/898kZOwrTpJnN+aRtkeT2ayXYl3BB1GkQ7HYrefPrJG
p+Mlwb98QmWNgHcTIUVFa2ZP2GAZ1qybRlrsoQlYEd1Cln7bmoNbP2S16FCl
eAwWBB0VUtEAy3+OmnY27tAvLkTNJdEJx/yEfmjYNnM6KJZ23j+s/OTdm9bm
FWwINN57+Wqmmdu7gQOx8nF0YDut3tIZjC5BRJvDUkN5C6jEt1NWN8ty5KNX
keaDPXKN3Hm7zxwsubBR+Ge1Xf10jFVsVuhbrEuuv3veP6oDYBu4ZsnoTYJ/
gnpQI3uZK/Qp+WCMwIfbNunuNowcJ1I01utn8lluzsw0IHShpgAAAn2211Xc
4SEkTHW3gOwb2u7og499FcCIL4PFGIMxEkJGHOORRKBDWk/5AyQO/AgGyvkP
ggpd8SOX1D+6xkSpBQFUxA3wL55Wb1YFJJBH9B6vGpttKmzpRnnetpVybweW
rETTJrrsHOEl/5WDAyH0Z7oOdhwjVdYx+11isnPiD0l2eYhhjckTLgMe+WEq
GbUFgHq+cRY5x/g8j8TbUUx9GYQ56xhhh34Xcu/kY3bcvFRudzsvS7/j8DVu
WxEAhkf3jiC6HrooctcLjvC5xgdVIWPdr99tgNA0XwXCDRsy0q6kdzZLd329
KNyarn0BEJktSgXT9xypZ7o7yvg1ffRx5I12eI93FNOe3B0PR108EKnoxYbP
sX8+ivFtvYIfw7M3xoYN499O8CEiFUvzEnEV9TEF5l6fhpCXlKBl3m1pxcwn
cVRn7yzwSQE2eCar6STnGG3FVOYzSJr16QR2WyzQ/RPw9nrunoD+6K1fv/YR
OzZtqr4i+3Uh53ZM2kW2usLhOyr2QRDgM3maMA55tyUROu1P59C7DqnKLTzQ
b2gMp35nKb3VS8a65a7iueoLp5qeJ28PVSWCL3ilTTxAyQPhKFvLkkQGlEM2
66juXOvepU0Pe9xmoGgGRvf4YOQ6KuRJkjUbHsje/3SNG40wM8YgRO41i8i7
H5TAVaH+bc29WOt4/fR7rNzKwyzjZ7effYAkNvf1on4OxA3S+Ju+rqCVlYht
ZGITwVi+BEqMHEIMgVfPuVfX7+B9GszqCPJSjzexBINfryIXfbsMQbO71tOB
VAoN/0aG6nt/G2PAcZgXw04OA5RJBc8NzOalQ5WmLGmsDKZvLkQOvd6adkeP
04je33tIQ77yewL8EeWba25sbkwXzrkdZoMdtyZLL/5ZWnE4f5yLf/br9Tvh
OcTmMAK3vzR24KZ6R4MLl6hCGCRVvudkuZP1nFJJx+h2SHwT31oqVhGu2jOk
TlPoATsTjCNuImIEO92jKo8kMVhZk9miSJAWxmVft8680RoX5Xz7ChQHdAcV
6UCU/aEqRUtUerkpSopqHC+/Am03usPgNi/y37mYD/pVxeng/WGXkCjMjOwp
BQnVHfrXzUd3KMcksfZn/JGC21bkIEAeodJrpwoSdtlR7SSGb4ZqdE0JkeYS
lf90/ijISR4ltdG6u8SbQUwgzM932Z/vIUExe5uZSgexc+1hxZIl3M7Le8/i
2V2PQ0i5qF0JQqfB5CZIhKvYYb3L1mU1bQM79Y1eF/zFXLJYiOTG8XubprQ9
TBGsQdrER8CJ91D1uv1IA3h0NnlQJrSxv8VC6CbWvyZcQcqxe5iqcDnWSwIJ
+r+XA1sTNtvDwTFwRnxICQpBaMtli1sDRR5y2ytkm/Nns0KuM2RpGqGeFAH5
KsAtMfuX53Z977E1hUeEi6/KjHjh1ObVqynjz9yjqDFkQHdsFV5OSmmmddon
HWPIQrlIlxW9I7l+tFjDYDXnMXgv3lN8tUGl/GiYeUvZDPELedaoRg9LuSgv
XaznPgf6QQJ+EXCfp90I25IdkZLiv8Q8iO55+EhZEveEWvaJLa/8pXMx6bnC
di/qchyS7yOXG07HtGIq1iirFyLrvwpDa95w271hq98JXZlgu2jlt5knEmu+
iyzrxJSEH63Q3A0GfOCyF3XkKIMMqh+VpaZXJzoJe57EUVl6BiygdmVIUeOn
KRj5vug1cAP95hJwvYImUjqTivYot1qOVJwfTd+XBFST3kE4OFwWGzgBmgiS
iTzo2E0D9fidI+Xxt9s0BsaW1mDTSkI+i0koGkucFxqZpm5txJH5AjdA1Q5u
XS/VJw7t8fAj1/bpheV05nfBF1lOVecSyocfuhZRtqc9LvDoy5ZfBLsEMK7a
xQleG42THjPNDEIFEgdILqCFSc3nXD+GGN66stSgrjRyPfiOLND+CbK0yn8b
EgOR1o9IMxTD/GfwwUw4VTYhNUdyg5DltU4IZEfFTzjiS45Z6vS3YXv4JCUA
lVfEyrJMvsnXk3fvgrc32qb6sJ55cBuVwoASq/peXVTXfHVzTgsdKggnX0Am
7AKzb8n7BVLeefdPMVUq7gaumON+lnYPsutcuiwifhKqmZ6oD0yvShDgiru5
+JtWKyr1EQaQviKYJnU+JIksV7OIWP87erNPDyCWwYKmHXWgtIlKJcUZMqn9
sP7AvuYSkXdbpqDbTT9L5PnjPPpuV43gdzWJMBpFmVNmG5XYjTlUOYIMh5MN
XiwSoBtL2SeZ/VLml/RXcdxmMKIrhICyV/eOKgjedVlWq387wYRhiYGNLWTb
iWc/gAkIB+AZxayTGoKhve7/yrJU8+KJbKdEWk44xe7t/nNGj0sOA1t+nThd
2dl/k5vCqHB01qpi8XZkfkLGjAj3rd+GoDW/S/kToRQa15Yk744bmKE4MJE5
5q+UpYbD9lRPe84JXybDEcoXlyrTQT2pFIQr7lO9v8z49BCq4Ojljn9aoXho
LG1OJUMwn5PbjuhNBF+IZhT2XV17a9iNIy+DNkwL31DGzh1LPoixmEQGqJ6d
8YVGV9Fd2Bpz7aY++9r65L6qoVRvsT9mlVkIysWMIsYUzZUVvpED4MlnjdRx
0xFf342mmoxvYfhdNbdr+b3e4VPgl5Rk9LVq7usUB63nRBJZnKORb0xGlywq
e/h9snFnCW3bv9dg1r6fqqYyu93KkJ1pEMJgFEidQwDYzPCq/anSr7xCIN3S
+QxtSEapSz5Rc8Y3QG6jCYzRQaaKsFOOxuLdEnf3eNZmsFRds7VX50E+TBMg
6P1GR+jn0aiUADRbZU5F5VB5ZbBvNrPXR9yqL5+JMkUmtTARG7BPHgTBsD7l
JDs0DLXLEOY2PVsqlIGNCu8A5GqYkb0xIc02/57db7OzGxdid5fFICGaUejq
gObxQyL2ehHv6NQsgntzZ18HZ59UrS8/akp0oXTfd4tSIc5NHAnXQtZ+qIv5
5Wnmp96FbxFQTM8XbtnPeLdqSj2uAMy8MDjUlgUIjp+t3Oq/3CFbi/X3hQdF
8MIdMrJfh9DhsDom291sGVoI0fbjJm542WkBJXd4IRVGfCDSozzgIE6gI0eK
LhZsDng0pyL9SnOvYKN+KAj0aTc3qVM4RGbrYXDX8BEe2aq8WwMUQaqCek+5
qPO3ZdgtZDJRaQ6WojYaxvkiafefer8bWukohOZJPvUm7BpbDKYJdd7YCx25
/JHlyeSWTbmfpqHtbUSfVljHtsTXFOD5q9NUpy8YKONFLt4XNbhMOvixJ9ar
22k2Enal+u/CnEH3FkrYxglssssJKOoLMlE4rQpt1NUMLqMzPtFIVmxk3TJQ
6V7ZfflH37f+P75JHjmQA9sRN7RXMfgptB6Eo35vtA8x4KVsNEXYfNT4mcyq
jgoiHD4uCQmIbKdEa/uX+9uaq80TMm7JSX9aLTapsHGxJc1l2F/qhHr4hIeO
6nWNhR+WC85l0+649SPqyr4Pq/mx2Rylp0PEvadKLFxHiSMYnWOo6d769lDA
249fVB5qmQKqCNQUxio7ZrI/azFeUxFka8wGYf48c2gL/lJJc0pK10uFV5f7
SRDrRUxhSY1b8Pygi/gOJLBy5553JIojqhEUyOuLNrleTGqF9kI6Oh/+0xOU
L576YwC09suZ7e18Jg58kEdmMB81g56zVxem1XrNQDISVngi+Y4BUJQ5n4v0
oD5pbsOnRvYb9Coyid6p2FyHXlOKyEcaqirrr5BZR6pGUKS/mA/PH5wMPcpp
RzWgwmq8aq3K6d0UJH9z3I9otly2BTjBDfvKSv5KczqE0da49FC8kvOpedQV
a8vWAr5Yid2YohsDmp5T1eGUrDoN3EbuBiBt57D2w5nWGT7UJt28zRx5ePgd
uEu6Db0MxtlTlGyh5jk/PXVPOCaXwRxGbSijHjgN1FevJ4GX2BPKPRJhbyqm
/iUG1+zzHTiweaD4xpoEVaMSoQ11Wh6WmEQ/0T7HdQc+wakRcrot9MtSxXc1
r1uESEE8hb+AZTSug5ycoYZIkCRH3UiGh8mQcQ5SDVGBUqJpwxkN1qRpJYEv
w2/4g2MJ2N+k2sPP/0UPK/ni1hm92smOZE3m9rLfcYM+CmOOlSOS3OYgybIr
xBVYkB19ArFTEUVYLHVxFcWcI76aS0ke0fM1uoNhgtZ6zd0ajbETJ80VS0TD
zRv4SIqZ9yELCVlYinDbCugbTaG3aAJXufkTIEe/gbLW13Y8EuOxUEVxwYHd
crWLTSFPQLV8oylGH5hZW5rKeqoii5kFdCG9eAE9XwHGnrkHU+MixrlFomb/
yeF52YwHDpDNK80mlhG7s66+/YOy0gBAXLE84QRjoAm6TNkRjhS3WASb3NxQ
ZLpICaGZRi0cUPpePm1VtoPAhASVKYryiYSKFTgUwKpU7oekaNrP15yJNM7b
tf1vhDcTspW6+aoDJ7x04yislgNvwAFCRp5dtpA1KTTf8PnXZqMfNbgd3NkV
YYp6yGPTWs5758v2WhrHapYDZH/Ify55y9dnbE9RSG1zAIdI/dDCYRzVqJOF
W2TNRxHFnQKSGbcyh7AYDN6y5U8jTSPFaJQeMEE/W070IBmgpF6vKIV18tTb
tbQGQImkwgEt2bJZNyt2cj9UNcsJcSknL6VsrLZ9sguTmge1LWaYQsgEeRtJ
qprnn+r7RMdZVU+3+togMqDNVI9DYX8EIGDFHpKYF88dNqVLluHTBC8m0cRq
0iNn9sq0pgOngQgh8fIvqgqdLrhKTBuqnG4i1ZlTrYQJ0TKh30dXPvhWpEf4
qyWP3lmf0C4uMXFhgtE4q3lRuDEADjG+YeJtHVdV9OvDNuhE+24f/v3rcE7z
v8je6lUO0KSEBoxX9oDeREOGkuJ+eGbI3hzmHfR7HUCzSKrC08ZIa4G0zkC3
PplFlBDh/ty1FLCfRe3ey0L/JuqUtu/ksiVeeYW8AXZnBvxbQOKkbQBCwLuL
RF9BYz3eTLc0OqPrQjjgy8Qn2LjgRw0l2UiXoK5juGQYJ1y5LjCF5BxeyDMR
psHNq9oMkbeK9QAjtLDKgPqV1RJQ08deifsMV92FSvbjpWA1d9oMeWoGWxuH
5pM9SnqJF39370uU5tmkB/niLd29z3Hu3CSeLJAt4b1Mtk79SSVxdCtIvR2c
ti1wzAN4pmT+JV52XQV5EcXDnO3eDgfeztfn9XWMbHNVuL3a7PrAV18EElZ/
o65MGM6NJhghC97DhThxftIQxm+LzM1f+xJNbQkcatRwxXnnQvh2ePZGidX8
F0qNCINSJx01Vl93wrFDaG6D9JE1/TL+5Sgm2aIKMp5z2wOWSV7DwzAHxNwm
rj4fmBL8BaGcBg6qvFPyj68efjIq1yAISgVyzygRwxMgAzFFNMd6iX8OBwnC
b7hedCQ6iZmgfXvcClJHN8nlniA9tqfzCrGpqhXviQE4vcjv/PlXi6sdR5qd
+ZuTK/iOWkhpmuaHTDvji5OhbtNCZHNFIApg7q9xNRpwiXoODNZ1FSSRkrAY
gl+BjWHjAP6nONkpsJK/p5Utzj4iqBNkUTE3ukCBeeU5pJbGHd3hsIULipLE
j4KIB2nk7BU69/fo56WY19b97/P8gF6Dgc2zJpMy8PdnWoTkGTff7a2tHST5
RunXNJaziwazPq6n1kdWsBfXEn7+aRWLTqH9nexZlcBkmuRCXfqpeynEj23s
1H40PPcwW4K57tPf7qHcRZku1IL50gqF601o4JW0Ma1E+wylHqVOAjyWWKCE
FmlsxH//QP1E5gm8YHDgteWIRE+wsYpiQiAJwRg9DgKrHgeRQvKzk6Ugp7jT
6FbvNGXZ873za/ZPD6lMS78s8JzLHxWts+3prZXSuS9zI+EKXRvMY6TIOz5N
yK5KVc4Ye3y/tceG94M2qjGuaJzQep+n/NkEA3Cy/QMXr0nVKaQ6ojb1XfmB
61rUn9TrkCgp2/eQ+aDJoOcWuZhgwE7fZoZp1dYFQnM9KtdUBDv9OIaxK7eI
CuIA/+kE9xDXHvLVpUXIKYMDHV221zr5Mx35TMcvKQZHRbyhiuOmwXu3J2kd
VT12UDRc/qC6SUl0Fj2R4iUT26IF7gYsyTIT0h+h/cSThc3ZJzoheM4/sxtb
4zKDBKzpDYqhoyHZFuaF4GrGXpnVOFhKWkykzPvu+WfFTMU6EEHbEZ9ae0pv
ixgXrnRxIYLp5ABudUWTs8MYlH7bwnUAAcOHwxyuzlOsEeA34O6TlG8pA/1/
nzs5XcL1Fz1gfVe8UTTZcmYudkCLfe+t/LQmNxRXvSGeUXKXtTrxXGLcEOfM
UgDdgTZMuoiZbeXc7t/9sDFSx+yADk8GQ3tDhd8a8g+xxUQEbH5XhpVOiIrF
gr/VJhKxhKKWwku4oPTeZ/03CLheIcI1SjIFxSCjfo97nAjr5XhcydACdeKn
8e8xX0SHMEvNwsfOBmogD0Estfe09ymD0av8IsMuqMqs8lIqYs0MpUyPd7rL
W5at4TKtZYSsY4w/vyjNZHxqdZB4pc7zZdD2h5vbaRmWXNCCJ6/Yv4oAGxdG
PK+eBKmuEGBt/rKKLhgMqmqhNbBMmBCrrq6SapjDT2sTX9Q4sFRHMDMW1li6
1iL79DJuZD/UqUKbPQP1uqxJNY8VdPVtQ4Cs/70t21LDV78Sm3vQ/LQnU2rE
LhNk9Y8gJQNaIORpTm/w8EtoJwHmt/fT/sawBxjiSWkGfAAK2yaR0megVcPr
pWuzq4iH0MmwfI75vltjnK889f37ZAZaJZx9PGKzMUiztrAquj1O5Jf/NUNh
dVaIJNhg9unVJ2WsepNSdy8MUp+IQKCD9sDCXYAwnb32Sysknx2ebCuKho3N
a6e7cnBmmazxHplgM0MEiWmdsw2XICA+ht8rfwbb7ObPg3N9dVH3fmS6pZiq
JHZFsWaoc1dpE2t2U0l7+CTU37xS1i0OBWPok8B/JLphLzbHi3L+yegNrcCw
rFHKPNdsz1qaIfPMPP1U3a1KdiaSWHSkWx/ypN96BIrv5hbyodWUgUVrEoNG
pKoRGA0S7LllAlOjFlVK/RT7UDiBmgEn+naOczqA9IU/+PT+iZmksDTxV+3g
+rEa3mazuu2eJepBa2u45znEH18G9tGQOVo8XEAcZrBDKrcdXcSofzf4PrGK
T81SH9M0fEg+ua/lpyQq/IGn/3NfLsCbPxcTFWrYd/kXyMyLyB1Xn0RXMKh9
wXzDDaYZ0xRBclGB0qXNC3l0otZ5vcf2fbmUGs3SJ4gYjrW5AHE0zh3dJEBt
DBDOmzNuSNKuGWfe+H67GB0afd/YacKBFMjl+Jcbc0yRrmxY3tKsAxkeVxHR
OftTHcAbHQmx2pBQ1nzwg3tkRlwA46b+/7hJe7pud5cJMFv92a0/YqriSTDj
dJEKCGIUKIKm3naGKFDERWLUJPID5KU8niyEku3lFvIM3kJ4Es46Q6YZLS5p
PZu8IyPEgmqb3A3wS38bdevKOmnwi1ffwUa6QlUrG0ivBBJirUhvrvb6aIqx
TespEM4NsZpom8sJslS2PX0nCXk/r0CPQw0v/VpBcCEr7++G+tWvrx3kp80N
x1gDhxMSkUqmWucR3dlD/ixTjKwSAdQaTPxinjcpPfHcuWnC35htWhxOMOFX
c5UwHl3SAzwudk1m6Z2Ibe1gUfs7q4RBzZuyiSQEohGSj79VFNyEfbGrkWaO
p73irEtI9ZG516zWbznUhWIhhVksZMijhUuHXEJk18u8wwPbCcffV/EUwkCa
jB/9m7Z5OAGGBnWY+GkKyR9Q+FMCK77JWPTXppKCFX0XuCHxf7NvC8NbZj9K
AEgWvWWjVQKI6TSbZ1Qpq0wqlRLD2+w3yBgptpscwFABlYgeUICumWzkZcSV
mQwY0fVmakB/oNlKaIOBZKZU77u3ei6LYvUYUpW6yo22He6BXnhCAr9gVI7B
v9fxG/gl+fVw0Z/Djbt0IEm7l9LcDRCqJdRFc8vAv+iowsDMxtbdveP9I3pi
RvkmVZHP0J/jgOnADGzXM7sL1YCk4tTH0n1wg37rFHDSvBAp2Nq98c8p7DNL
S6bwktg0GvY7/qCSi08qqGDo+EjinoANhJx6rzq2rZ7x1EOpLexZLaiv+SGM
z53Itt/RWhLvwWrxBeyKuCnDUuJHqJv/5hO8kvMaUiG8ce0Cxepua21H+53g
3qwLTsWOwSKjOCJVnBpjcKtvuQMl7BbUsatY45qvpSB8RijEo8NYVcfABcC0
67P5JPiGG6WLBdsayKxWl/yCWSWBnsomJCIaGpgHHDx/BANThufdsvAz6Oqj
IfUmwgpANKwF+3n1Se/OWMnBEvgJyxObYnvcoSvdsxxhqEcPxP2nunmAvQ9B
OZcQcPIk2naP7Vv8cMF7re63FNUV3RfEAQxeJUSg5xndKz2FaeKuyEonOhPq
zneKQK7oFRqTxL3HVLHU8aPZqxfqoDbZCq7xzwfwaue97j0kJUnPGO86Zsir
qvM/OrG7PKD9PsqjI8RsytLZn8rMnBK9fsM6jKeank272Ip7kf0jX3k2ZNq8
9gKGGktFgmZVWWcv6ErHS8GLRMkZ7rWkrTtL6zytyG31BOKQ7qZ+dRW0bY9H
6FQ9QkxUsg6MYZ7H9AmRO3gyiVqoL4cCpM0PKBUaB5sT/Kt0zmWyIfw2i4xd
7ccVDaNXAhv7CDedvV8KEvHGutIbAtXJgI3Axt6eVUCljQ0jzgjjd5QuVsLf
lg6VHg4808Kc9CdbiW4T43FReUxWDJ9BXtACqNcT3yw0iVLoemG1BQPW98vh
63HkmwYTIok47KkXsL+UZjje8xGi0W665JHMljtER63CMOs3BAVekxSJ8KvB
52oISByu6YHxIBh3fUR2776xJe0Gvr48dnkc0TZHZl02BHnNOrh6PKaqCDUe
tz8LdivoIADwju8MO3LRFdjmbt0duYbz1B9XRRUXvu9ri800Y7U/nPYmuFeX
NFg36f9ymHOZw0k7u+Ez0ocPi7zL757szj4TE1VmqcMAMzZc0ywrHTxCGxjy
JhnzXAjA0wOShQZO4i0E3bZSTPMLIsc2MrkX66bp9P/UzC+y6eWwYW23iD1g
u1pYUr0YzHzVUfOCiEjDtrxzP7iHbqgwnes7jV+M5GlBxEd+KCaZBQI9zXCN
a2pRZMokbDfNJRWFt0cCxh1tYJfx2Gk/VeDimU1wnO5W2nBFLkQoYGrRka+K
IM+zjSatJ72qS7+wwlYvqa6o8boMq7s2YdCBGdDkiiCvJD6S4mpOBtE19ubA
p92xnGvsFApWWcewBr8WCQZN750xmUVELZY0KqU7MvXZg0edrQi+PGseCPRl
qzm7LWL16wl7HHHQL55bhUAQfr8Mf0zUsfHgyOT3KxJJSGFgJe83gLCSCX3b
mmUJj54D8YZuz3q4TJUJZ2Xfz4zr9EHilHGpCC00Wih1HFS6lvvWwM3CUB0Q
ls2d2Lslf4x3fhKfSLXBXOeU3XwsUEta/4jEKeY35JE1JvmWseXiYyxzw38W
RgGdYJI+9ozZkioDX9jkEE7B2y7NnZcjoIE+OYxj4hnpZIFFvf6zPInS3Tss
K+vZ7KJKu4DEWeehZ7lT/LWUG2vcDOjrgqyCk+leDXBeJrsDNkYyAyLtaeri
RyoNIXJj7aomZsrb5GIPCjQfP0PuL+zZvSgun2Eh0s1rh2QTGcYoQpUw7hRT
H5JSh1eKrlfTJMn+B1FUpXAbFchBBb7LWZ8CUXsyMJtRnDFEFmvz/KgwrXwK
KM/b50JaQLUkU/2Imuv4pdNRwgla0fpAoDZBQdgaJvyGEbxlXn8Mh3iNqp2G
Te0j7JAWHxge6oo7PHej/iCBCjnmAemzdPYsNQtLiWsTgtseJUeAB1N0XUSs
+ePPacwNk5aV6LMlL+fF/sz1scs3N3PFo43B4F9N3bZaIFU6NmZtDVxG2Pv8
Jldd04f3q02pyW1QkL/LvYp7c2UWiK1LH4s0BXVf9nhI7JZuZe7hKQmn+td+
8rTYImo9jFAjeWjri1Hd4i0Z5Roqqx7KPteBGC4gTL7sXrYS1vXL3YAfi9Rj
4J5+iQ9Y4Gti8uwRnERlfOBFZz7HTRvwG0rI3rGciB8waMPAVUeXTarwgjLB
+7mHIiIa+QuXH5H/yiF4mBIRVHTI1+7amTWiC/lLD+Y6Nat0mfrg0kEMUabQ
f9l9extjmzDZhgtJdgr5JnLIvtmzsMOObPkdtQjCKx85lX6Pq0KdawSI2Arx
mkfPkH2MSNrH0chHBPIHet/HM4Kem8xzCOURSjee/Q7U8L5C67VNNllmH9Ja
wYOJdSVZoM0lDQoZCqk2h29uRlMhe8Pf7k51hSJ/abivHqM1W1aLPvc2nrOL
sRa18LwCK4o0Opyk1PcblEaRN8hOTKDtL6HzWyJlHRxBqtG0GrUWCmrceoZJ
5AYd16WUSG0DFM5BfBgAT/bejx8le3p68Lv1HH5eNeBvybXq5ohd+xOJ+ukP
QoDyzd8xbkRIttWp8UfFA+OFCBT1KTVJBf+L59cqRPLuGlg4LSQj5iPOpfm1
agO6F+7BFeIvIknjAFzwcnLgM/d6SOdzyygxomTQVcuhybDlNJBB9/oPnaRo
5uecsmz/OQhkbu7Yj+jOfesOyBkALaffS/CA1cFd6wbYsydhzi99ftOuEZFF
WXlIpWKo/nj4ddeY3g2nA0xxPuk2tAhHBezhLYbsMqg+2ik8jtdn+9h0OC04
Sb4ycYcztjSDCN72yaFzEll8q0Q6ILYuX90W7ZSTv9VLJeaPXMGsyuFxulEx
EUDXF4gNI5UFZDmnHzxgZLC2fRyOWZs0gBTcY1SQgcyRQc4fsuyUfXX4ogd8
DqdCvog7wcDtNqIpNC/vmKrdUof7kcYlWp2O2QIJ419uJLKOn/caSlXuUuMx
4dR+fxtr0hCYc1D1BkhNEHC9LDIXP33mAWo05kwGi+XE8+KEXRK849seVEdR
69qIHBLEfB7SvaCjNXeBsl4V+q6xdov9aolRk+F8irHp0zsMAq4AS4ZmdoUx
aYtUoXLU2i05Xtld3XEKoFytftuSJ+Kvp/fAuZtFwbgeDbUo0mTgUKCrO5zW
Fn6i5ZHLOWGbfSUi1XJiDFcVNO67Rg7o3oR25AwrHbp8KgEdDkHS13JN4dQE
CDO9rOOWVVXB/8HhoEI9YTn6J/c6qUdDmj8E5CX0dw7OycPevvXH7jPe7s1G
W9o27EBC9iXcNbpvKWeMOzkYhEizTPdORh5tdrmQ8v4xZb8Et2xTTtBybXeX
w1Pd8NMXqwnxRJC2WlIlnTWDa34uwey4lcSdlOn+ZxCrQBvbHJED8JOzicoD
KuOHAggtoUvP/RKmrtUqhZ9rHqmxshSVrjsVc/DWW0czUP+Ec2Na7qXP4xUn
qKrdoALriMiedjCn09QTgVz5cHPjO0ZtxMYUSzAgaZFc1IinZm96SbEuxuur
WvM+qYl56olXG91OWxF1nUWIlCQXAB616PeW6mLt6E1fljK7C1LlZyA4m15S
UGh455Xo29mAwuFgQ3y/w1KqABWTN+d/AenYWr3o/BTV2xWttCp2YlCXhB6e
z6xMoUr1+sJQWeaxvujaXZ82f2KKDfU4SBQW4gb7ZWC6zyyZ/000hBEjFkEJ
CtI8R1sDSieF8k1qxV5iju8IP0aYrSsJ1UgkPEBUtOukzcnDIeXBqkCbrp9Y
wUzFYp8wquiWemVJIYBJkPhTnEKoBWV4I40N9OE7teyemY9QiYoNhTVvsC4j
QyM9fAbBTdDp4AG9sVIzTDLZjzA5CypB/Eu/pIpnayHeDqBJJ+CjSdKH9iAD
80lxRDSNoT1bJjA9qk9NU0E3pA1Vasjsy7BWr7Ag/C8G4fdLsSFaVZNfjKCg
Akti+KChzd/qaNvSPo/rP7N6ef+FsqmWi8EDngTCa7WBHEy+DSf974CoMSID
KjtNxhrwwe/sOIus5X90g7zKNEHtzVeFxMb1r8WtGd0x12UkZkfsA2HZWSOI
ZibDSS11l6719+x68CAwv4RngNqYtc0rujlU8+4G5wJdVehDdTJixV0Z+mcZ
OwZ1m3LPkJRU8aqoTWTnAq4CmUHRYC5OrjovlGP9px2o1wmSQgggmhb/XEdl
l+k2D6xxl67qZ/7s7Z9lGc0VZFxk2vUqp3WsG8mPb+4SqsD+gnf0glItiBN5
hkSLNBX3Tbidzzqu04je6501U2QPC9lsIkP+4UmvQTe/kn6Mge3+Linl7iV3
oMrb4ikqEuwS4UvX6P4sO0/lsVkf0FVJgZX4vYU3dt/DowZmHZ0lbnf9uVWQ
oRXxmSlUT3JCQ/uty7nJaHkLbgvhYRMcM+YMJf8HtYp59hwo6OxUkXqFbFxV
isGI/s0cowBC22+mWCwNG72SSw4Ty4fKPEnrLoQUW85h1oGb1h06kPFVfSth
Mv/+NwZekRbKtSC3jUNt5StrK3Nz8Nzay3VYhlyv72NsgO8Xa+3Uu5SHyEBF
6u40gbTRs/2P6phOznr1sLKvYKy8q2+pHjJkofOfXJmsYuRQ5n75hBJcGmlm
7YMLiDJlAJD0SGgzmthyArQ3UYVmGlTmqiJnkl9ZbZuLup/0jG3H7nX4qxKB
O07HryjcB9YJPRg4WSpGyLYEN9G7SqmF2JREB+4agbcN898jjX93MHXxuOOx
ePtQzarJ1zUjn4ynGFk/s49Cwq/V0M+6SOlSS6fg7/tzuK7B38VJ4xKrl4rd
td+GwKMaWDaavJI2W1Zvm7FCoz7IRl/NgYXRMptUeuemehLcz5+A86OW7yEG
STKUNwk3+cenxVDlAD/aF7lSxGIHQoEaHjs94nwfVVI1tRksBEwggy5v9kBP
hMOCMrSe9CuOiAYO2VW72euGnhrf3KCkp24yyfVaCtS99P27GIZaPjHc7ht6
Gq8k1WqL1TyCYzgESheEtLEV82IXe11FzudC5MOHrcFSza0lwemUUa8ZdVfj
wDgnPmb7MLaxqZqqfTHJv+X/m7r32OjRRDk2Bm6ToyBEznYzde9XrJ437uk5
VW7ftka1I4Fn7fcnOi/PwsN//j0y9mSWJlqN2aJVHe2mUpSRyqwDGS81hwLr
ZTKBt2blwGpLbfjfwM7/qGhHL+6ckVRGSaYy6xL+RWP+E+a+dIGRmtUFSFct
kSHNlbk/7MbwlW07JRHr0NPSXpXG4ylT3wvhi3ZSm+y0Lgf8pM5ToHdincbT
7WCpA9voHK3gcvIgme4mivY+mrCLQyxCiFd9HWe+DtxNODolS1/03p/fnLv+
OAaR8Hlj3vE9tA57wkGKVqwKUfMa1KLdDpic68txJYVkM0nHnN3lK2NNIWyS
ZcEE9Us9N7O6uKcMZ/3ZLDJGglFb+qGzBtlyFnjlzSUoYmFtZ1oyZCsp7cJf
YZEY99bnfLbBKgA/oValTJKIgyfd43SPI9pysJZqsG38OtqlAvta+st05JSs
kNj5sxVDbPuqgF/NTcSzEfYnfkssvwbHVNC2Enc8ELRaYwF2PeUR8kdbnXkz
ecENYr35DrBtk8ZW4PICyOCZPEeMzLy3UwWFgT9HZ1lcQF58xd+ilcfnuc+j
8Yt8dSEhqDGnZMaRmGw3hw9OjkAQM8QkCcLTF9diunIG6X0rg0H9003TANGa
nDEgMOK2e0O1dH3OyySLL/Km25G/pVhuFRZ+qKgSqyRMhq8YOsWGKigXFBeg
HZrR8jVUZIu/ohQ6w0NHdh/U1XPS3uVLnnYDLce7JNNJwOE4RWYPyCSHNZim
juAH8NCO2aZsoX9R8/4SwRPZGRxGp1G9Bv8+iRe+YBeIS3x6NTggvt00dOR/
rTsCxsxcAGDh4OYgqtAcPlOqafeCtgbYypTsUN3HhHtn03U1/Sye20LSfH5F
V6bcElt+PpyI4OyBAuKm0yTEe/wO/Zd8ehqEMjd2LbrbuYQfkq69m3RlgmVZ
M8nBRPqQvTCKsLi4BUOHCY+yQW6/NVrrQXM3FDvihvLxBXRphLKVnT64Yv3E
TD+7JOEJj5F5Lvk9DjGCCbvkdI1b5tN2PdWCrQQbOXX/0huUTOb3Myp6tY6q
C0aTkaH8AyC3C/KdOenN4j1PbQiHNFJPytHIEyitgpG51ZI4VYIRymPDpIWU
IlJriT3FpO4DrBcT2hRRtOf/hzGWZu7hBvvbXDRmkY2iYQqUgbrsUTyy57B9
I4voXBS4Ckwy7+Z5APrbWgl2li6nGNYTtBmt7kbdMj+UWtCwBah+dArWFiTK
sS7f/VYq20EJkd1Sn5P6geHo+6VitIAjgAuVfxpLrBXcWjZ7GEDipipWuOte
AmXK7XiOqhztTOZl2Ty8Y92TGSFFnFB/PfAlulrW9YKWR57M++/1RzqOfjmR
j5X+MgQRssu0VnGI9yFnyhKKAHQD977aVxyXY04v+1IutBAveWPBfAC8SUpH
+WP2elZFPHyE2PhCcyWrGpBcjpGcEbMeJgrW4Q49J744cxTaZrS/IC4u97wk
avK6M5B8ZIU0s9Ln+1e8XlBcHHs5QrAeKq9YXCfXikJVMdXHjxyO2AgiYysb
GPPrxu0piIwLo986R09kLgI1RFZfheNIyVivQcir6DSZZaYwAuTo9WtyeNra
O/poutGXkxXR6D6NC5s0b7zg/UBXTB9BYKyPt47jEzJVpmJZjKzKD/5mQ0Gr
m/c2p28VFzqnWcLLt+8uUvGe45rHTGjsllzyQYAle9cqiAuImGZLsr9dAg6a
HYxifnnVWZDfWt7Zly+dSznPu4+scnMSzy6Aaes2DPSXIfbNoGh1APvbCWfv
SR/L0RE0/PQp55l8JFiUF+OX1HEa8751Xk4aFYWiQ7rXFG+16LvpALHlWMJ+
huCVNt0s8+2MqRgm1sJkve0eeoDeXWfFHMcT6u85csBw/OJcujZVu7M8+r0W
DH+HuOPwD+6j7V+MAKEbzeTfgCKIRlrduz9X6w3I0IdZ4cOB6iLC/SvOJlsh
Oidn2R5Yg/qaFv1A1euml9WApVGDNCRTPeVBTHYxDbynlItPrYSIEu6z+nH1
45q2K98czdRWJnnEm9opyCW5mCIO13xsMeAUU0LbjHbldGmi0XbTpA5uKAff
4RgQFo5BXGvbNZFgoJIRTVIlQ7Js4I7vHzQ9b/Eu8EIkj3JxhLU6blbKIo0p
E6prp2/dLjgrK/MzhpgdSoU6qcn33ZtHC623lPNlOo15MPBG/XV+KBR58EaU
oY2KtsJXfk3UPQNauDY8OKOj1rZJ9PlWOSKdMLc2XL3P3ScjomYVtVf4S31a
fkg7+YFESA6BGeM7BrZa3rH+imLBxsvE9Qq2z3mCIwz/Qml+FNw3HjGsgIdR
PvbEKKgLJLM+uS7EUK0gU/9IOvW8jjdGqVoMakbZ+ibRpmygracjiXQ/pEyI
fp5dYWRcZGFtMIhNquN/blc3s8jHWMBdFEg3U5p7SSGkzemcUGbrcbe9WVgn
BqsNESQMst5sxG3diJeyHljm++SBKDB8bAqJ70VRs/sHkmxQy27osC4aeWoU
ymswZdAzs/FWr4ReEAlF/ORpDyNegBS0PQDhmLl0SzyyWKATioHTqUR06lii
Wyv7PZqmRrn4Sfj0/BvHN8YHJzkqendZz9AJrC6gPo9ytZsP21IDe7qEHLO1
WYOYefbgO6M4ThDX6Q/XsrWRwaO7Ux9SdUY5b+mZBaJFiLcAFGkT+Wl56uB8
kbake3iC/u+to6j/T0r2kC9i0yaUWY15PWrtOVt8bdKhyj2IA9H3skSd31jA
rx6gfULMyXsLLYNipOIvdaWR0+yA4b5wh421uY+1piq51DipdtONChj/z6qA
ShA2ThWT0g6yiVyqM8UqUT0BMZ6t0ijdVKAs4V0xZduJ0donHLehx+W5gO0A
nTYa7age/dDhwH/RkX5lD4EnH7QGShnnIgENae+VHRCb5MRIiMpnjxE+ZxJB
hYXVCtr77dPb5mNr4OVutMLYaHs7z80bG7q3i/oyvHb2AKvug+I2HBmvgNJ5
8dNgKllOTJ20rHAAdOw6m/qPzgw/tsBvGbsWmFyh2Jsk1Q+WPWbz4HQsCVYH
1IOqHpNAJnqmBPzSr1l/EV7S+asdLNl5jMz8Ym9vwOx2i4SmZ6/ex/fx4DxN
Y0V0BV1W0xzyHc1IZrMC1XlFjR/q6EcerChGSsnYK08filUrSG+8uBmSKhaD
vaELfuoFCSbvaQhTmSEvJXc7iC3WeoJ68w8iHOmy+mCYIx5tenpJ4r2PPYjW
XOAi/2OAf+P3E9Di8bGXsQazBhuTkW6sgpzBTjodxT/dSIYOxGX9Bc6+X2/P
frPF3ixzBz4TR7ERKN0k6VRaP7B4HLvmPqgT0HF2sAlVqOnIKBGOjXK5M8bf
odWvk0D/vXpH473jNdCjuY571yHS8X2z0jIjlX52Abhorbn23M36rBr4XCup
WXwkFyVOooKirwJ+fMnNoI/OC+62gW0miGvUj4BsCQnvimoeKSvmMT/Q68vD
lsQsu1iriHISGicFKxw08RBS8uBfngJGE6boX44i9bx8teJkJolVa12dCE8Q
eQF1RwYBW6KmbfLOKKkvNu7uN2QRwMWJPrw75j9dtEmSoXawpuEpTQMjPqA6
xcuHVjWxoSwkBXtc+cYg0ZX+ZA4Sng2DYkVCO8pP2a8FX5O25nWaI+MTD8IK
PYtd0vWqoEZUC8N49AWswzp7h6mGLUzZYnEjwk7jyGo2dv60pFo68RrIC6vk
KT5BoU8ECSSPzVj5iuUNEpkUypxOn3KD+5wC+YeXrwHmxZl7SEmRo0RaaGDZ
gOM4IHxw+sr+ZMeYxFrOhaPb4ERwUTa/vpfshlqwwJSnFbPPj9hAaGU6JozV
sAceUwDFXFhaek074KW/rv9+F211PMV8fT0GUShyBS4wgCO1d/CODiLDRV4c
AmpgrECneiynukPWKlCsj0W+Iq9SH5XrtKG3vSPbXlH5yQNu3wBbZCBl2CM3
IzFc6Af7UQpSDO8vw9tXIRO+QV7AwPPAuiyz5c8j0MGPYTKyJy4G+KhIkT44
+uU5mir44Bxb0s6ipKFCsyswX48WK1JD/10CPkiALbPDSuKpLD0Db0gHjuCL
LdmibfcgSfjlQ/GYhhSiOP53BVVrw6cizGf6ZPUfHnldnzVIkI6Z1ok22WPB
6La2M8ZnjmlgWU+n5MFbF2wi0TDMGQERw5Nl2MJbt5i0Z/pKff6ASy2po9Vy
A6qeugu6k94iWM5UdNrTGzxUyGtOjOaUuFNYS4AFHv6SzBRQcdRtQf5iEzpf
6ubvFNW2fLvNCES9D7PVCKrRbZCT4hlumlQ2B5B5nPWRzB/QsaOKYWNXSyOB
VQotwKMfoOzJl7uWA3UZZNttt4XwuHGJLlp93nbYpbynCPQrC3YRKo4wnZGf
iQn3hvp0xP76zY0nn4pPxAAeSy+cQud2XKsEiz5fIczt8d0D49phzV6jt9we
IqW/qNf0FYII1cQfMpOOQ5EQUE7CnXcVKfoirrMLwVszzJUuv0z2IHb1+G1o
wxPuyxTayLpGxooZaqYjzBCaAvuiz+5NwaqU9jkXIyLLtYC1LIU/lfHxILpk
CWPtKfCOK+dbL6CPbGofi/tMK8igIizOys38ylv+9ryuukki2K0IyZsKtILW
vZ73NAETk7e06JVciPHAKUxWjvAwq2cPLliALuwTURbCdeeZoIKEqXXGbc4U
UIbhdJ3K6GCl44p7wlADCHdnzDtn15YPsYdVxeO9Adw8AlxL6EnlcOeONBjs
HLZpfu5asCXuceIwGje+ODprT+E5PvZ1QD9UqM/5xFAS1W327+kodFjW7o6l
bq4JQIO1m6Xg/H0d8KEIzWFAN+NKe2hDFZv26Q0eVD89RoG+cP2Cx8MduGdk
2qeXvZ8z30xkp5RdiSxcPDQBLWJWQuAIKmzZd5zaNpHRQVVrmpcWcLpceWD3
hnP/M9CzSpWhjBOCVMnlB3dmpXhUX7S2vLJ3I702Ul8+l6JmZlCLaeI1Qh46
111OHkO2P/8bHcWnKfvrdeaPsFttVM2t77EdRL1wnbK5MnHME2AyT0SJFnIr
0oFGmpUEU/zd7HXcEGgQo2+5BAPSuHf+ZMpjrYkh2aLOM6EoWv6bM81qkAHz
cz0iuDU7FbeNKxYUtPKfsfTo7L2cWFFUmONqug7QSopSaRdiMtMwG+WuWWNd
1KaExRmMqaDogJIq4CWwNlbh9yyUyQmBf+jJIwMNtmLeNe+p4ArKV1W1xEir
AJ62CoEEUSLa+oyJAWL5BqBmf1402VvijgNpa0LwAGmo/bdvcwTmgcjWKrtt
EtwNl4LDlZ1894yxTXPk5IF7V/emRY3NKHUuUTeLtdcPFe08GHIWmP/vY7Dm
xEjxLshj7vSqX80+z3HqDF7Ek6OZEc3ZXXWjWC8bJfMo+gqjtas3QwbAW0vp
1yQrc6VH0VSUIlys5SAhyhph8AR3nrIiOslNT8omc+0fxRFOQjab3pCoCjOJ
nhlH5uQv4Q1wj5ZbGVA+rzHWwTvH1DA6XbkCIY2Bz0ARUyaeTjNQ1plIedlP
kT83i1bG4uKcukp5ES6sDlCP5zyS4/+hoQN2RqQMg+lyWh4/a7ZSLaQJoKQP
O8MaeZSnHzCoxHPz7q3gI/IEgSWLF5cO7DPwFfhS24YpWwwiP87zZXPNw0Lo
K6EPBCua3J/8G2G2nvnPnBanc/sWgrWWXmY7bSrbHNZJibxapPv7m2CJ3GRN
uihqSjzcS5dLbqOtW9ufaRo+XOYN3XNOmQ6z2orhtn7JULqCH/jW8yJV5f5E
sJAR2IeuPu3onl/EJ7IoX+oQ7wFIGZU2Djr3SxtWwdpsZsm9/Ta7cIX+wE+4
ovQPFMXWbllKCdVM21xcWW+rXFPHDzSH8QCY0d3I4JhsyRDRG8wu241qHj1F
MJ5jkiwmGGzk7tifXq2Ha6Ee7tbiyMdqZZ0hLiU0FOC1NRJsaiOQopYQmvT2
6YEHObRDITFjdgWwGQwl19Q71tcc5izkaj4HcLNGaxhY5OpjD0dqL0gNdA3H
qXTSdYPfNyrP4Yxpur4tUv3IUAsUd8BtDRU8SLBlbtMIUgAHBbmYDsuHHTFQ
OZLqWFvnSxCagTiqFOtY1MCuR9XaK6Oawd+5gzQCN+z692MV6VoeqkF8OSEC
rEuPoUaPKG6WKge8UIwAlTyLIMVnqA7wvhhM4zR7vhQ9BYRDSY3CQZ+PHWym
fhUR5we9k9a/48okhh+/jb46HSChZiUu8Jg8Ccq+9S2aDWEaF/ZHugytmlRe
XqBusBy+1lYIg9CsHWISwW4Anvn7Wgdo/EO6h5tIwkvpJIl/23OztgQF6jEj
TyZZuaNdJz3wQvkbBdYdN2qU5NMq++O+YFXJ4RjhpW1cWWrw1s71yJaAOPTg
uM54dtNmzQAmoXJ+Nb96nclp8BV+P/jWFUPtvRt+pshXx70WRq7MKOajgP+c
RoGlP04fwqs4B9YQ2KEmFtd8wUyKxs/pnK3uxl5pHB4EZnglSvzf05dmKje1
qA2ZQs9+z2mNy/O/DD1OgJKMiQxaD4RAHPZ5bRVlh+3IEU0pTTRaXZv4J0M0
q6xKbkLSjH4DUFWOkUUVEat/1JE9XJPEOOBsckIYJeCUWyX+QEpkJ+rGmsdA
68WeUfIO/rgmzXDr2N/MGFisSnOvUj2BiKGmfjLaqCL3wwGHzqkNrU3cTyIS
AKcMMK0eYK6vsqbm0KnpwPicj4FtP1gsSa6JsIIWRgWodS9otUPZrsUN0TxD
MFwlhPJeMXVQHCuW5UV5iJdRuyo2MkcNERY6zaQWnYY7UO3MxoZQsHkhGP7P
t1tdFWwu9U5s/mq1v37GRwALZkuRAYy4HMVQ8yUk5qPWmNC+qXv8fFToicbi
JEMkQiTrwRYJiGgDj8M4Wc3nAGZr6skmXdLDCQuh7YeeTAqr5vponbysoYcV
wRipykECX4j/CWzuU37jDdnSTMzkp5bDSwflnjr9bDLdhr5YkTiB3ElRlGJu
HnslcLtl+MJ8wMdf3NLSk/sA7bsUBWeLaz8y/wUp5/0l8zzybfGEYgX2nrIR
LDhwgJ/3OTYwo5PmP1LwpLcyV17eCp+/ebyQfeTnYiNCfIfCvQTeEKVtLd39
3ARayCQsfjtXK6P9jtYA3M8SEA5dd3af86AG7T9nuFjjV8BCDw/0RYkecHvY
ifnGyv7AhVPn/yElc6xkWwFY5vCK1WNSyQMrUyKWY/KUi9Sg0Ipz/Huf/pg5
nuC57rbdy6SGi8xQ8RwfCB08tuQo3/JE+kVi1Bfq8BxC2Pip3pscEtTZ1LA3
7EZufQZcVfHyIB1kgXGIv1MireuBN5ZckApngtYFxNXAHwcmd73TK8waWTaE
V7obzWUsoluWPl8BKAkpVHF4I2pwz0+CPf5x90/TDHr74Uq0T01LjQzWqUU8
qLfMgT5Pz03E4o5yM0v1Id3pYmCfFb0XKCGx0Mmi6QtPeLo/nHSQkcP4Z9lN
VVxnHTNnFvvQj6BZHyD2dKVAFIjBDW1EGWAHJi1UVO6Ipk0rAG5FlPubVAc9
oPtrR4BWixyxCpRZB+IutPWZo0JEorkAjigc2UvEaFWds028QEIGDJgMPEGk
h+kWpE/yQvuoXw+j+lUJScIOSQvHl4AFbJKjC5LnlcLq4ooYW8ioDOBjkF7h
VYK0lm0zKqb0rsScQOVNfxHfIWU5iNc3rT0SiUtPnH/495T4vek4Pszxq44i
ItKsTpfcl2Ff4qjWcB0j63+wUXVtB2KdJd+zgc9+jXDGvrEiPNJbqk4Q+GLV
68/yXTPp0WDlNwABtmR6uqUxtxUoc5uZFXRT7gkt9DYzLZs7R9Ef2Sse0BTH
TJgKosWpN/bwswsABFjKLnPizqN4ipDjMOuEq/QgVavVsxP/qypwh+wfGaNe
hBNsZzQspeE3nu7+SYh10lk6P7p4Nw38ctrXQkGVjtNvPQu650I+1yTDvzv0
MrfyOA5nToXm6qScsLVyvDirgelsWY/VgMxUUz4ph1m0H1OWphmGaTPw5e3h
WaYbPgYrFQZwoqApuQ+3/Kngblu9zmC5kNd3+OLjZY6BZpstmgM0bZGLpMl/
19k4kI9Oha7LzZYkwLjSmWeKkUJihnCLqZnzqwHYcTqn+aGzyvIcd8ifuqZw
SukAQpsY12/i6Kzud/ZV7e0BY5ppoxN3csbAUATAMXDD//2IfiBvMTkRkIiM
uZx4FeHZKERufN2z40BrNzXLglrHiv+Bu7LHqMX4QaSrid0rID+ycMTjQuR7
TySCkJcOvFNDXIm8jEDnBFXRxV+yaXcnWdn7/uN2x7rIcIqggHB51tL6j9jM
gtu8RTM2bq3TJH6qmjZaYumubrV4stpKaG9rNtFB971+UFm+stOqSygazeQ/
bOkpTZrRLdHskPljR+fawt+qFz4qQP7CHYkJB/kanYC3HNqNB/WcbuVhwI7o
mN5vp2u//8o9TDEGMHTjfszPKWXt9heKUC9nv7TrNm+kq5BjIdDeBTegyp00
lLWwVmUV75Wa/kVA7rY5msv+XVg+qHtQ1SbuSOOyorU6Mik2t4lXpjpDYTto
51L7+OZt+2jU+FVk5CACtMeArinjiWWTOlQHq/+PyrNtzFDQV0c+T/c3CQdu
Q0viZoV2Chmyx42TdkxaOwslnj4UzG4N2XZ+Lk16n8/6Zc1ndDEdPocFDKtz
g4U699ALQ1P46a2VsG09Ex12M/eFPVpzDlKstvIeugyDyHiE4t//DwwoqE0e
g4HmgS9ynJ4LZ3YKBgDqHsD1vpFeZFDDwjFZYFVJppmNqnGjz0BYvZWxA8DF
HCiDE+fvrYVLZx0ftLSFdivB9BGwfmNmVYuSV5EcRP9O/FyBzQlnHq6JuhPi
hCQm+dAgn+WyKLeihcjP+eJAGEp+V96AdghCyHzuHWE1ApIrIJTsYSt8q5E8
DDpvKL/YUs/aoK2gQt0ALvyDOj1y6YPyaXLdQQjdZnvSptR7jzqmbcwmT5jc
hxBk7HUTdu9UePqggEDVfPgSzSpp/5lMMj/l/cnPFrjrKaT0mEnabDjwkPM9
ojd6Xv/WC3A4/yqWUO/lIqCW89tOSVRAVJk8k8dWT1n0viT643BK4Ig/dJKG
InF5B0UaACZUzzcR6vbBk1Q/B0N7lSy6Sta9Khz6Y2c6FL8jozzx4yFHpQE7
VB59ZsZIuhzBxB9aT4HeHrh7qP9At9rMh+H+s9mxu25Y3liteQs5VPnCgALU
zwhamSRYWrdCodHYVvw2SOHJV1w2s+izKYmDOtUuWcp5qv0LM1YkGfxSHAOu
jVkGepMymI1CDv7ROr9gWl/EFFwwJ7aN8ohj1twxjHnJ0NTnIvhSNUC/+Qg+
XtOQ+B+1273damlyRj99y+UAYz77S45qWzbIq+qOJJLTM3NkE2CT13K65Lsf
t+pEwEmCpiBM993WUNPcTQsrofJm1dZtB/UDMeTqIerhTp4vpZWv9+ZMnFXV
eFa0RvfqQcip2kgPRgrndjJWRwgE6SG9Cpmc74ZzK8O8ZfZJWouAyeC8wfQd
36MtFeU1CmXVJs7ZP2TNCiCvZyr3MjCiWSUt1cm7pT1KfPHRevtK/LWAjvBX
xUDuDt2xntZPgW2pg/FZAcoOc9jGxSmcF5s8k8Ecl8Bxkc5vZFBlTXruKdXs
Z/qMy5tXvkb9QItUlcgFau11SXOQRXFh2086jYl1OCFP0jAjN2iTCU0lpTZ/
9A9wInK5lLU4YsW88/pN1HOeDtJuFgNLZ25QHsJPbrDzhwAG5KI7exGa0Xg6
fsRT/V/mopVFoWmdLYJ8X7N7XBi0d5/IgLcKJ1ZHB0r16JbDnEv9J2S4Ph27
HlmkTNr3hMpI/FPLbT0VEybvgySYV4rpAHioJI5m/E69ojPa1xyUlkE8r0eE
gWcnwzxfRlvasxO4w3FzAMbDbN9YZbbMFgarskpXyhiWgpKEvYcP8hXMk5m7
slrqg/2u9l+V97jRX5gtca+vObVPgGbe8VEsFoqkCg6drCh3GtGtUjD4MiHw
7pfxIfzLkxH6Byb0RzR+dvyPdhECKESlXrUDkmHZEft1LOx5x009+raWc3kC
y2AmCJJSpf0Ri7n7gn8P6QOmxGxAZKdDadecz9uXnAZUnP51zFGemjrCvqv6
H8eFlRhzCifTmEGW/np8sDWEotf3bkduNwug6VPFipL51ScbomtKS2Bt8NE+
S/B9+fu+lAauRMMWDumukdzKb1nyXKzstyL34S4S0C7+7nn+B7eSr6u5iibJ
T1Me5XX9tFHD9L9VIqylcmiJOsDNMzwyrxI7SP6YSNCZmSptnXc4ng+e1IzY
FhHSRq2Y9SMVXG8QPZBOwdyZY49Ut0Sa0KtX+H+PhSvIsWh6TY4HVMaTs56G
DTxdZ4dsnePYx6yMnGGOvAn32OopJ2Hm93fZZ0ExD7vIN0qlgfnbjNnB9EvL
yowQ3sHPOMc2bG2PwPTSLzGDyAv2H5gtmZCdOOQnBjFK+5aPXuw6FSsjBL+s
VGhwtdOJ2sQMXqyoaOhpn0EIwmECK1pPWvhGEBc1yTYADLot8d18RZrza0da
3tqD3qBVp3FluKMqVE1352DZYLuEKZBai4q21YwakA9I0QscwI9QgDKdUjRZ
PGQlXJPw/K+k4bW+v/gceMzcyIh/AU71be6GBTXvmzhJ8yQX04Ur6n7cVGAh
JAMvocXHnlG0/bjVsxU/5/BwPPJVQ1zP//hIaY2+DLxrAEKKMOEVf/q7JcnQ
MYPqTF9O3Im2Wkn5Ak3COvImEtP/c9T1RRtT9VjP6Tv8cl+bEDQeMEGGwBnN
pfNM3/7uV8R/suTWvWdZDz7vbdAYj1sdM09UnFCswUCQiMFI+PO3jnwne8ti
ySj8bOPQEWkP2HkpccJK7mWoEgKGrjblsAUCpwAmfOyTvhmeF6C9L9jcVaRh
IFI7XVjEEcCu8eWAsrxx+dlu9qpRksoEIbqInf7TNWSTH/VoSmNDlqiSlrUR
wKbCFbQ2HM/4NA+p9bnRSqafvv3MXJwubxxHdiFBZ3WM3VuryJXTnePMUh9A
/6SvIYvaunnu1Q3LdcLv/8Rt/MuEtbGSp4v3MSfBc4uVZ++i3HXuK7W9wE3a
GrE/7XDynEEht55RkldpJobC5z2FzHJydYVeJoGj35/0cHGfC7vUcBcsK+yl
eDvYWYpmILmbj65VH8Dwl7CnpvCypG2FD0Hly541nE2V8KlBRjr/DOFSgote
dA5sfVp3unrvy5wapJLquO85rz8ZVlaSJw8V43OtXS3aFwPlCYZZSMZFAK2u
VQRdWS1RVYSeT5DeQBvbznkWfdTfafLdKz9XwBLdxcATFBJ6GszsVlZnhdX3
SLdwxGL1cMoTPNgprKWwiYTMoo5oE4xJYHQ+yTsCCoNgZ9kv65BTz6xS+JFJ
+CF+b9n8slYM6uU6CifjlQYzobEbeF4IBRVUCQzZGEaAvNB3OikG0kAEU88j
uBTnKECq+hKH4jutCfoWRRSsQzsHv4cZkYijwYTG58ljcnwz9weVzHQlE43N
tcyJs7RFer1wNXUOQqw4ytkUYaBn3CzXbwCJbFhG5HCWRzhr0Xpul1Yar84z
AfJ2MmL+y9HNJJHl4AV2u5iU30/UgNJue37zAX2I+jUDpMiy5S3UO9vmi7If
WDRweeny9S5o7JP39qeiW7GmOvI0Z4KdtRsMWpoCW5zZzI5IJ9zhgjfda4AR
r9zAmRuREkDDVO88iJE+kaZc9hrhUqD1S65toepQinS3dxm1PjN5tQKOYozH
PHQARNFkig8dPUltxWryvAMBcfNHTR8P9R+HuHN0+YnZ0w3x8crIHsuRdseP
ajl8xefSNSwzpwdtlFq7GQr524wa7lciy9Or1TffWED8jsk+NGSCJ5ScGr3f
Rmu0z5BA4Ud12wBD87pw6LwsL/SQi8EMlYfyxgp7JiOpUZ/NE3MzEQH344y5
HwsI98itcn1PZTGpbp8iBS2MxUaUOpPxDO3A7dijwkDRm8Xm779GmEv0NgOs
kFBXsUJACxmoIKbhytsKgoCj3MipA/xFr3JsP1f1xCSLVpL4DOfedfDd0lcc
vhBuu0ZvAtDHfasnrMR2iy+tjY9knuCaQ1xiifHZPlvvnkC1HBXcW+IE+Vgj
YxHd7v+6YgDOeh1Jw8oGPO6PcHzpU8H8s+XfVFDgBUSwZM3F+rKAQ4Jk4g9o
gA/2+P5TNdauejsO2l0TQ8gn6EmiVee7FQlVeKwpFCTMNazsDwqh3VIDH3Lw
T8p/Fqtg04ikepUxt/DXU8ZVUgZHA8/U4rFyWzqOqKoc0eewPy5mlzW8nAv8
sYYPou/BketFgPJy9g3sVDJHu1pvjB9lxVrL6yQb6E8ysVcFkjDLYmCHXbTi
uI9CM5C3ykWaadhUME1TxIu1+Lf54GNCeursARmm4/Td5vjlDyueqTXT4f1z
7IjCOwL+s84BLV8ui3cnAma0YEJ9eyMxAb9uxUnkNHI2eqjslDAnF/DoF6Ag
CEt16W37riKIYyAEkXMuTxLX9PViMEyyNqptM7iS5Y++JX5CPF2OXdy1Zu//
szSvVW06lC7HxAhGW6k1RLbzVHtt/FuxjN2jgSCagPyZmY8u2dwAh5IDExUj
1xlMROmOxR0+qt8o+Dv9H9HjE0XFIxi0w/19GII/9zFbnb1bjxyFmcJ7DZk3
Gfs7Cxql6sxdTlaAz7fYlqbCDZhOlk6VwB1NPxDMdMKyEEHRyXyj+T+QRUdP
YJ3RBE/zEMhMl/1qW2m5bxrbuuRw1CM3wKViimeq3yFfvJF9r2mSPW2IZgoV
iYdZAyfch9ve7hvAqyfvXnq9O7ak8VPcK3ZVRvxTiu1erWVmGdB40y7p0Z/8
sMH2MJlFAyDDWOT+nzGXOZ2bECf2yitfGlLRn0TWnXUIJN4YOfa+pvmHUh/W
ppv773XAnTq9s9SXzMyuUqndrFuRZC/yIz2eYVN0EWEd7eOFlae54wT8XziQ
cb1SDDQSOUnTW6rEqJit1AT9U9+6SxudA9eDYIU51/ODYybeZSN3iagAkDOC
23GDIcfS0pVndg5nO41SThjD+H2XI8Xe6tCERvdYZchTwNWQk/iRrITzPGin
GI77Gb+ZsyTHa6+dpcF2+kFgvcY5xrKTMeATKaT+LPAIv82vF+MAFMjHaNoV
2jPbgHA3xcTNvjpRT74qHIXL/P9+Ln2wrTk5e8WsdPtaQLi80EgW6uTCzaQk
DEozo+uRwt18l5xloqeifGumG4m0flGanQ1hR4EBvmMZd9+dI2q4MQVjKo1v
TQ5UFiOfoQqoxtcqJcD7+q8OBT2bulXDIhii8aKp3RWfYyQoNtVIgcnCvyV/
tVCjzKPybzJb9vzpAC03ZNez+oX3OhMP/vlGpvt1yJc8l/7zAvugyg7UDMK9
d9CdWkxM9F0ie1+cdglz5Dc/8ST8QPQB/NJyWEEXPdQFaKDXhDTTNSBlCUnU
lrzN8YfTTW7jrwG23UM6o+G6K3fES2hjHRUj68apwP+lSwD0/pDjgEub3EY0
lO+pD+qzZPcAkA7zNfVB4pzR+414W9naMdyHX7fGW8fKiucLwp5rp2bPT977
ns2j+43KL43QTzfCj810FbpVGBG4DOxh4fV9aBRpHe4o56AiwHlL2fbJCOLy
IKOkJOXH7Uig5xs7haM/zZaf8PWv9YHLF9voKE3fF1YgaORre74ziukERb3m
0AccE7qnOBhmEFBdWz1IORh+CICwFopvq1Wrrohnp62zS6rGVkTqO+29eIXH
evYfS7zI99+dP6y8IzaLP4U5wfnyuqGOebNOmauU+crMp4SnMULMpB6FR7vR
g8Z7nwc2nACdgG4RBWBM7TjB7NcwKYsPHZkcMDBIue42lwQ61A0gmytShZ10
akd85PbV60NPk8u5ixJk2ZwPAD+oKGEkSEJpeKjeMwVez5+6fzuZ50oiU1ZM
Xz226mBqvIrJ8bfRTi0EmRdFkd5i04qCjaBfBuqr3UQ/BsqR6oXFCmeBFPPz
Wet1trTF9Dp6M49E/ir+o1/sRp8amD7OaUyzlxohEFySVcACxEagyrHVANG1
UyFxjE2YbPPn+b5q6Tv5i7jfFz6hovGteDPwn8fqFAzED6CQMDqmGZilZJ1u
1eR/opt5nwLGAUoVIqARlowum8PaLK+CpIsxlvSiYteXdKFKYnpMeH3QffSV
NuoXQbM7wrx7bxlQUiCpzr3wrkOCS8kSIjlyqLN5kj10zLZqGYYRxdN3xQQH
nhr9DXHSI907pt8S71Iee6oJJhwFgDWXKAasLXWwZXM09ihTk07ZUFTJONFR
edwQoD2QBI44CvGbr+rbuyJrlDotHrcnF+9jxW1vF05IQITZLV6n2QLNjO7+
ntnO/NCU90hC6hdLS6ZEU2oIKSKhgectprrHwsZ3fiJVYl6FIe+A+DSh0/CB
QQSSzDYAQkOMvOK4gxebyYc+wknia3R/dKBMa4LrVdiNBeE9cVhdr92aQ9LQ
bH2kf3jTObwzsJ/LLvKuaMcR0xkr3YcF0F/Sly8UFZ4EruuBZKt97Gnjg1xG
AZRo0POxTjtIPp70THRdPKF+xWuOFb58rS48CUPTGi8ISMuO1EIZaTiZLghR
LTQTQssrCWGruu04PftsB1CFVvNNQmR+TxYvzQv3SnTqomkqnuNrbHb0JjG/
kDihRAIgH0ZPA/rsMg9MZ1YA/76xWkhMKLQbz4iGPGfxXLlD+RYkJ3tjcdRj
YBZPtGuOO+sH0QrusxT2C4nsUSjfJdtCFU7SanXT876oAU5A8LU5Bha5BYM4
vTLYGZ85UoA5koov6T/F1avcL+rVrYJfVh00VmSvxdwE8w1AUQMFFTXoBPmO
x+n0FshNX88ms8yPNfP+U0t7RyzPe1yHjH2PpI2tTVV1zGMFmWbfYj+DcWxb
5G3HMLd2tV+puidsrwFykjcUi5ZRSaXrs/AR+6Tai6qAf7S44UFncWxfS4yD
LYbl8PuM5wTqq+KI2AxFNItYLNHyq1weCXirZAW9SXnAm+5Mdx1SP56CeH8X
0C6NI7EILWOoNUYJc+8hq9l8a2L8Ad5tngWBJpncV/1iRQTCjstiv3kNqYTQ
B0F0TLtaXcR0rFL+VBoj8IsRDo+yCLct8hfL4UjZEq10amRPzUw8rpRjC9Zh
XWelTBtpiU7YZZXd41rrXNyBYbbkXpXIhIW8Cr5HT1G5LD/Hb5aYwRkBIH5m
7Ucg9am02gkJVBaT13aVvGFmLLF4bApAiwqFjvQT8FY6ab+FL2Xg/yWa7EcE
ylB+V3B7vN3YJH/5ZbKZY0aokjBTSNWBm3yG6xbD3z0M6tY58c7soLzHrtrT
8rpR5WP1b4ytiLODdLYrnWjHbd5eeC9I9w6fgUejj6dV/HTJibNc5tup+n2p
yZYwVAaQ/uDdoRHIMTXHn9ap2KyPD+WrehQptkTg0JAzbKru0/9EWdPxuxQg
d9/ikIa4g1xmRYbAVymnrNK7ZV1vu2OP04LpHFlThtbt5Pqv6/zSBG7r9uCw
8b3y0N+U/olJwKFAAEOSixNOSgtSL21joKlqrl/1iou8hKSJy9yvPs5T9uQ/
Hdi9JBgpIy8W5poFWgbon7/c+k3elZu46ZgseYcWnGyP3PB8ehgoJIk8LFnV
t3Yq69+1QCjs1ziH09NSag3f4tXKO89pWbttr3IgY2Qiv/AUmwIygkoEcpsf
d0QyQsKyPoZ1Is6CALc/e9SbEgOxl2ThXM/oGhFknc2FVA6376ub53M7I1Pg
NOObgFSqunY7cTlG4v6UfjBn2yXYdsFBA2r4dnW+NPCLNR3AEFdgU3zeJW76
mIGV1dQSl0xgvP1AHBqzYmiFKyUAcy+snoJkLJgiTbqTN9mZJ9X/YCAptAp0
waCQIAQYZHfVSeRYpN8afD1z9KnbfLjWjjRpFLidQ1w9/sEX8PtLExhg3pkp
ji3GcsD0NPDfRFcPiEWaaryUhlQ5XAjREgp365Fw3fM0rBuNmUp7v82j/QjI
NlIn4H0qWYGRkwHdyVumzStI9Faq35OvtN3hfUA7sg1eP6qF4OlvISH3xzNz
BDQepa1YrFOKkUYkf2sI3mnXwYaIvuJ6WGL5Bz9FxMm7MMfk6NHJIVHriqd+
WS4izgeRIliOHjcX/LlHbuCuY0ejwN03hwwwYuKgY317ctl/MjUJe6t0umLO
MD4Kn3MfPYuZyMydOzyr0/THbrtBecSMnjQzxIlyP/PWfgQ7sxW+kJDkL24D
bAvzZur2jIxkm0HxFGacYQnn1OPFP1Fq3byJkLxzIj3m+jCuy+NVLUpPzLyH
aEjMhoSYVIhsho3DO2qtHhTArResyLO00TKGC8VVulJFALB51ktLSFEwz2Qz
rPtgiKI5kvInAXrIhsgK5oA1n9F996OQ7dPGEwYTNcrW2vu2Zmk6TTgpLeUR
QVdiD/X/BH7aHRvV47aDujLyL1232e/0s6yZOJY4FtXC2rCp1MdRSY+ArDMD
jU8qv+Crp6OBFp7FD70T7+yPOWd0wSYczIGV3QS/o23iGpAx1eyT2h79Beh1
ppjofuI33r2ngi+W3kfE9/mislAHQS4iduUvtU2IkkyjvA6ogaEuVtlVHjTa
T+kkjP5dgF+jAX59/HveOotj6D+R/fmp+I372NVPrTi+jOloPtdimLmcv9io
C4vOhiRdKSQslyVoersItNPoJSm/w2kXvTK673Un46CMLJuoqnz4Ivfgoap/
nTT7RGLDR9D9vUJbba6Exd7OSrijKKy44Y3y0RZaFpAuu/kdUUKknQdlQdOg
3OazVCjx6L9q5cKKQKY5QGAQkLREP+qfgsp7tIg0XtimwuKFWOj2gBZsmwjF
bMlMMZJYysztk1ITTkDjATj6x+//r5Dw/4JenuWyXs27uz+t8b5LRGkDOJxO
esJZ/CLWzMH6hDXqnvPoOKEbxc1QFWiSTzwK8AxtYOSRC0DaYIgq748ZcwqE
H1u7Dju2Z+LNgCG/rQe3WoqRTb1cGzaOiCiOKpKs7fYM9NyQ5TZi3jQFCdX3
locIwOCzGJo9b5bitOU4jrKqu5b/u8H8+pgm2ItKINIGMOzF5rVj9LESqyuP
X1LdNH9EOcvYwQ4sV6HB3Ts0ZG8OeXnCGW8jFbdCs33N6QOqgNq8GnHXeXz1
URZUk+9eBBgyfkiceqaCIZlEsjymYtVJPzVVSRQbO5E6tVHF8hn2r9LYqvon
zb+X5UKWZVhAMAWUms3sZTjMcuXvZVk6HMjjZ5JT4xc6b2TcStnZBkqz+X1V
u9Y+dGjdZ5/kIuO78gOMqJCTPdahPTeaZGcnQwIrLjb7oT9CXy6IJGerQAR1
Fx10BPtoPdC5lSP79+Y81o4JI6hGACiAaUampN7XQXkIv4iR7KZ5E98SVKBS
5KlaTLIQAyTp4fKhbom5fSNJ+zH1W38UwcmTYCQsNeBAPrJf9yR0gaujiYTj
5elAbFZNU7ywpP8CHmbLH+6+MHp+/7/Z1irNC1M9IVPqt421MxJwLjDO8Y3R
v9LLv/koir90+Yv5DeghKwF5E2lVfF5OrM3orERpPciC2tcEy0SPSUq4ZeD5
cfyN3qXB05Ig4G9jUyY1ZMpWgPMSVB6LlJSH9CzVb9TnCahkkww4iv6jr5/H
keP225O5AATL8joMY2TO7e5a8GfZe9K8lBwWzaytwPFhbtHc0UmsAiDvyDu8
joO0VGv5gIOnzJOwIMQ8HMVg403X/o3ngumb2vlSiYICzHwmFHwz1tTgSsMI
RqR1rjv6AP5VjI4jbCvlMzyxA//L4z5omHweTbF2+yy+DTp2F2frahW+GH+9
YkSoshIxFbO2jlHildMgxid8NYPixJovfD2c3T+UVqEQX94CZW2QUEpn9FJV
crcbMxXXxT2/O3DRUOPX25GzxKeRB1RIEawk75G2Oeki5leR+u2po/wJ1Jqa
DOd/b0tAUTTeu9SV48TuK2azE3nF5WWH6NdoWl2ei+kbjGJBBLEQcWXOTQJ2
ASD1iVafedpdqCujfg7xpHDBWi9RQLGJza68KEZ5hKwgHCv0SccGmrv4O+2H
ovtlfdjML/JJyj2rEFbiLnUkuJWVtuFS+MJAHK/DaZRZLx6XwH91G8OnR3Sl
W7nuz+5GDK5d11tr2hOXbi4j+KCi2UpW+W1Wi26bdBKPqsDy8nHxw/vIl/pU
M/zT1v4f/gNNwQW+tKu4z4Eq0yu6Jtu2OVypZbq/2hx9DPNmA91RFMT2Vn6a
gqoxYFYCOHuUdVoOKaKHZqCfGG17QWAqIG420g2bs98quqH5NHkSHBMy24+a
WgVlnPT26B2DHwHvUzI2Veevb9FyJDRoiIbycyZteS3KMUsgSTMw4kCSbSIJ
l3FI/HMkINPmJsE3iV1OjECuFAkP4rGhlxM+zPdjPONm4Kd9Ef6IvsDHU/iE
E2M33F/RrpURn+oAjkQbAfOMx8i7PS1qGXz80Q4u4n3n+mL00oNNV41410bz
I/liVz4zCzLzachWv0zCx73hyBRzMbx8Bn/B4WrD41lMPGepscsESQJ7QYwA
RJ9g5f8DGsnVcz2s5ojoTNvlT/PjraokU2CSa17Klk++JI8v28qu5YPrBdEK
edD2fRF1nIrJhiGhA4Vz0caUOoVpaqQkQ3Qw2hup8PRpu+lezFwds/oiX8UM
v7emVk40WpeaCT6f++6Wrd1wgTyaNdc+zkWNGNElkQXJ0cNbmVof8kFnZ7UP
ukecjMR1a4uVuDjAB6SFccLaaMYafyeCrbMu4GEKuOowJc3fu8XoAWvVk0Y7
eM8p1t3HDUkaddKZWoL2M8hkvCr1/qEBncnm0WMxZRtSSmcv48xl3BF99Eiq
fVK8Jjx8FbWInLH0cuxgI6sr5Yd9g6r8mAFua8Xwj7tUVhygpdaVgM0iBnun
F/OCOhgnFwTud3K31g+dX7CyGnyDHiXPlxvJqF4679mDCvsSCJQ/0KNwGG/1
f2fKIr1fMGCXeu3E54j03FOr3pCY+fKa5FU8WSjqQjjS4Xb9wLSP9EbAu+3L
1V8yH898gjdnXbFokVCKTWysV4Sz0lYr53ucqnKMZWHJe9PzDYk8AYgLMW8a
a69YIvHPmpRx9hNPGrcW5BMe6yOjYqKsOqhQl8bk5PZgxVaBQDxzJ/CkedK7
bihg/+9DmcJflNPOKPHytFQ3Xvk9J51EvhHxQqBqSfsey/UdS9YIgDibV3/8
WiKXAXtSuKbLQyMBKIYWP4WCo4myM7n9HixDCZj93SGz3D9IQIHJZWVW8eF1
ygSN7JyvdAnlns8asLdeiuK0WUbl8EpD5Fq3SSpsCz1KO4cimA38W3AbaFKo
PrUlC341VyH82ASH+G8p6iK+6brclCNv1SB0dT1f7yqAEhniOSGmxqOMe73z
586oskBEeTkcC9XHwtiPCbXquDAf8hmhfey3LLXawkLowmgKFShOMMfuP1c5
Ek55+BmhuL7no52f7MBTYbdk1tqUpZxjXDSzFJImI86DHBkwYqDeEnXhZBK3
HU2f3J6DdIQpYaZy8a0WYzyoQ88bOtrguIpPTGFBeLwljdyMLkFgSTrDOpTx
8u3dNeeCLZn65WnB1X1D1kyu7ZTIBzOULOdXOs7N5RVO8uN+lShL30wlLuhE
RlmYt6CFzKtTDJ+7dshRu5HFttRWBWr8mxyG/j76P+K1yV1WbvzjGLLbXZk5
ANX7Nozquxsm68+RPpuvA8nBvC6mcbLBLnaCVGUehf7MdzjPPqaAsjFnM+lN
MyM8G5fb9m3eRFsomBPeJSI0AvprxAJF3lVbFrg4o5kzaYkAxzs5olDao/EG
VGfXsXc6ATEQzq8Co4cw3CtgBkw47owDbzvKtN+/mxFefhT3fWpeRyNdU+WA
UxnxnUWMtEzSWp0zw/Y6WFXedIAvLDO1EQLrn1usMg+ehRNN/6LI+Byr/0Y5
5SL1BMAY27NaXC31OxerSweHHd0MtxZv5e13PlYt28bFW5A4J10RMCgvInY4
IjygSCqOmd3vaKk0x2rQqTIeEV8zLKfTlrRMCx6lpLSJk4Azw9tiEAUOvz+4
VrfvWTQgtvVJANWF7Lfmm4USY3k=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KLhwMiudeU5Ct/Swbt+xbzn7Z9fslQsyz7LqAzuBnNrol3mzBEhTD7DtYKT6kbmXRQEUx4oHPgQLavKZ1yRy1osPOnh3nRp990b4zkKrM44omuylMkZX0NifvTOvTRApJnw8JcZ7iH4jiToqzkE052y9EXvWRzopP4E7ze/2u1RxGhx0uG+OxB4zuzoUKOka4oxCl7JVyT4I6M3hmtIjOIIrxaE8q4ohuPhYJ8sRvXf80Ag2hDOIS9oEhbkTbeusJVK9OR7EFtsbHuDK+EM02yT4vdrCMNNNUiZtie4KB0oTCyUyzhdOeAK6mAIt/2YzHrS6mRlkJ1XqSnABbiuYOrIucHiRj94ZeHw3/pXFjosnTC8fGXO57QV56p+wuXCUQQKA9bLDnFABFJQAjeSB/g4feTR95Nh2bV9UQLj1zuVa7dE8w8zdEoEnm00BSdnRZtJAeBPB6Rh2tx7fDouTykYufxYElOqfwOHew0UD0vpO6XMc5sp+FQ7TJ7baqeElBvS9D0NZ4Nsi55CazAZZHMomBkEs11z1hHE+O1VdEUvQkXkSmP73XCq7ULj/xfJAbXhie8Mz50LP3CMziMmQmNTppW+Sz50C1YS4xxZRVrtVATCRL2LgIAvTv4HCpwo/jA/7fTICNb17lStuzlTHx89sTAkMZ2qzEBSJwYvXBLJVq2ZdBIOZz5Ur8jvT+HBCPOXZzo7HI/0gLKr6roqUJAjPZUhtAgj5/2+70SCRxKu2Mb1+D+7xNXuCgklFERF+TKFfPqwThSoBhjxck5X9Iv"
`endif