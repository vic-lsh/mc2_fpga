// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Gm55qQiQWB4FuoaTAPKC4jR/UhoSePm4Wb3TC7cdosz4whWEvoD78e/4X8DK
T1VwExqOYde93U6chEtmLdMxsOnxU9Kbq1dxxLdu4OeiUNlLCWS0BQOwX3nf
0k4jZQy6vNt/4rgcgVMty8bGHAcANiL47gLfuE+zJwU83VzU5eI+CBCaIG8e
rCa+jFoeLWoPy4fRR6mtOBIL9XWGO2o0TqI0lZP873m7VV/gZfsDAXATuecQ
plMf1a2EIxBCPPSskjZ3b3Vlcsw0GScM3W1Tgb6gGHLUwYB8/hvg+kL9dp+Z
ZWY1ObXLJ+mMMpENYxyt/syqmazfwnlbzWEwsj2Lpg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RSZiUwp5aTzKJXLKUh1HMVpfjQTYFozhBgpYV+NdF4GQmNwjt475pkUMVJX4
uW6jxw2tNqawjgNOCeQULGwkZdMQ9MN7cmYAY5AxLT3JtjiDTev0cwILs/PE
cGAox8Ui0OmAAy9d0Ji+Z1yqDou8Xl3psqSfrDbZT5BtohBu1I/PV53EvuEd
lDvIfg1KsiDMZ5xEdPI9ZlPzjF80Dm/9vFKf6KIjRwN+W8Mxq42BrcNyYpNz
sDrWf/CrI0phNLkrw+uIMPvHxFU2iOL+/SUd2waG1Rpb4cW2Lc2r4htT6tdl
deWcjitjvPJFT7UCwYDPafPPHW6fsudMvwvR+Vv3IA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cWMDHebjAdVf80AXOLu1d5KdOqTUJPdK0Rq+AMO+0qC95mNTLPi/2OAEHkwi
lQDz+NrSEyRJBmLVLt960E2k7bx8bvHYBMSpeiAFxuhKzDW5oRD7fnwlvDsx
Z2kO+QhhY7mcS02/gfd8ydA4P2Mu7LUITedmDehxNF7LaY1LqxmrUCTnIejV
AlPJBN95qPcwwfK8zxKUS+rfY5WoADVkwAsTZ1zc/PhhZd/4hO+dgNxQsMTn
6/9vAVrTMG3tMLGoqgsJ2EWQ5LQPP9Enc7pMkwGt/preTcphM70fxxzw6QSP
Bh+dEsI/cTyAxsPHxYaf668ExgWBc4cpijXOfZp7ig==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gNHxatQxZtOM5+DS5KbaljREX4fDLZ8toujJALklLaEY8SeOCQ7fZaN51At7
/XxwHXa+pQVRO4VgwS+cfw7TurIuLxidDcNCXALd1N1sr4IG8BKqsMPVEgit
iF406qs4Jn6CkWBrK/5xQakp4BOZWBY5fBL1y+edz9DgEySWk+CzcrnQ6se6
gr0qz0uDUK6eeY6r9cGGMT3sgfoLNvJI0HklRycTq9OjJeFdPo8Yd1ItPKUk
SV/X4P7+au3D8q6OMAFN7hHUiUQyeJys1WtI5wCffC86jOUf23/6xuoUvINt
J8AZphxh/J1uEYTkwUFbw8cX/I5VFykfhVPLmD2dXA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ThTiRjuAFV0aW/cg4jSrn7g+8j9D92LbJiw+O1mu2CM84p/IO3QxPoUM5XDb
xHsyWh4dJBDykWLxufDZTidzV8i9u97Mfqebhe4IC2faQ+p1uMzfZAgLyg8D
Bkuk7GiAmYL/1+Bl5pfmsptNNO2kpbDsElXwHguRZokLNP4WM0I=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DMvGs6fNmxcizS40Jb+fmYEmN1oFfD9910hVBHfIOaBnGDfMaTLr+XZzzty7
qfAZXWlQid+yQd9dz6ay98Qw0k7gOBNB2Hs1X+XkNk+GhB40GyninmjFp0rM
YFK+6MKGaDckDnyCaXzCWldunqZHj/EjxAjwz9ErYixEzO7HMOEZ2Lfx1R7i
WkCnOHc6fiBFdTH1ltIl/b08S7CEnuyjkt+Nu6JgqN6ICVP5lzwT7lZznSjm
yeARR7RL0lt9Be/fLUwOeX8LqdMbqrnO9doUqP+2kHE+4imWbchxjRHsUxpF
XkSkfYu41UJ02aneanYLCoXSWwHcEAqiN+W4Wrzgdj7GduFA/gX4ueF/0gSJ
fx/LWDKYDmC6iq+beCPituqTVH/9+e7YFYwsbNQeCgzlVrVD2JdWBQHa+blr
oYEgrwN2NvBtOCwtV7EZF5qvBX3HAzbKJYCIq/hbEc7JMIYzleR7+4RIBWcU
VarMWpx6AJVmxW39LTZOSFdYp80Cv/y1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NcUWcNzskKoxIfCVHgvSJb0yZ1L4vA3lkXtkYUdJ3z1dtlFW4W2VZxOYi/z0
0hk3YuecLtjFHlnudLjOVyCbVSBXRjEayBj9B3V83PK0bXhPkmW+/W5lcaDd
VFLNkBEa40yq2W9SqbzZemk/hLwzifMfTjEjinExLwu5zSK02nY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nB2LTn0Fx4ZdWN0+Gq+vRkCNRZVGtQfK0SuA5/goCWt7nayfO3VcyC5fxZPv
mneTnI/gMHDkexmTNF8uyOM/0lDIIkXmmqynFNl+EsO1AVJrI8sDnBJC6eO9
SLBKpa1SNWm1YTddvyvigCbd3Rm3Hcy9CdEWaQMJ+yVcaUGpj9I=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1024)
`pragma protect data_block
//bWkfrV7D2+A8YxuQSfUOgCK96zwvfqcK9kQa2vmKzBq9DZsgTls/M+gM+j
czPA1GT6zI28MRrKagtzhSqYvHZI789SE35+c51TEjD9V+zmsQ5DvknepW2A
nHWl0Xjpq85GasLoAoepwbUphyjdCPp1aaaZ7gsKW9UstnkZ8zF4J2PdMEHW
ligDqcs3uyFgzBj1fYQKcb0EgWw6d3XXRUXyGYcb1/xWJ+1cpP7mBn8uqITc
PiQiMSqdnYubnFTwoC5jnkAA5RUE5aBv8Ias7Mp/2kO27bzEV+EF7D0Zj7N7
08hJ7zRn4Za+fTqZHlLG/u9l7Kqn0YMpJOt67voIrxr4PPTSU35BMZArQCfS
Ug/fTY51e03p2Bh6UWn0Mfs76dgN43jztQf/NmDyVSbnUpuwIb24/uUkg+Uu
skOcDg4Bh6AbB4nFyqcBpR+lEEeQ93F6cL6/HGNJ0Wl9DoDFEdDcHDT2+ATi
QPz5bV2Okvn+wVkNDioGEcQ3JHhekftf/m0GnVQQKPf9A+H+AsctK53gmgqS
PvG2IH0RVscg2P3B3ENUbGUQ890UHLcj6tJz4mxOQWgpOqNv/7ZAkhwmDffb
gJ9HMf/QYGeK4brKCgDkGmQBmv8K6P9iGYVZKGg/sFCWqUlhXijq9VNUlryc
9UMVP9Kcs/3RoseFS990HLS4J/1D6X2p3BziMgBF80rrqLxjj25mj+bhsINv
fMSAgs5I02xjQCSJYpZnsyciuIqD7IO71ZzGyS0vRkLa1Bg9pjIO0ap84hRY
1/x+6UIWnKMOoy6Ad5sH32NkIUL9Oj2k1ADsVwAWCWdMXObB3Loy3ith3HA1
9BIUzS8KPVHfcOTuHMZjezFVGaZf+o2Xi0iFYgrq3N/ZBUEgbB1+vRl8nXZk
WcO809CJtlwEQluNKJc92wzUxvfKkauJQ/EQCyVGRpyUFyFbPeHRQb4HF5Ol
+ZMHAlggLlbr3YyTbTiteSDYCNPocVlc/qohIGQtUUvmFkMF/KdbZRyy40Jy
QCbPDFjLRwIC5mCgGC1zPYwfbf9pB0VPzZIKJlAwDVDCbb0aSZzTGrMgNv0L
fv4XidNLxMM77zVIirl9XDG3kJ2uF0U7vv257SMzDoWoQuphlMJMJAFdEFvW
VuB7cWkd4lFNXiNzjfzqk6AeHMyUNcq/YK1Ow6V5hQcaWO3BibtznkyKprke
i69FI0EBD2tNe6sJuE7yXnglfJbyvoTqRFePNATTtpTU/jTTRrSM9R0tKYl1
Uud51i96Lv0HXPJTllePaNfmCcL935CtNyz2CmmobXxt0l+s4yMF+rJauHte
D7RbE3fPjt6y/jGtn3frNdZPVXatRMyMFa4GJe9g+1sw9Q==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqf6YK72nUsP6as2wrB/gzP0PoqrilrxBL9km3l7sg/oi3E9uYIysd9B8fMjpYN5pOys+dvwSVWtcp5NgXS18+WeJGIdsDcfRT5LaRv+hY08q7PDl83OS2h0BtuyN+bRHcZmUowBUYxiJjBv1GaKxk2+HLT+txbpt0Hko8PyUXs/GvPJ/qGxu6MKKTtZcU4LX6UKlGf/afB3D9YYzKRZImnKTtjH0k7g62G2BeIQ9AhKHQtPingKaMXsZ23Vjeh8CfpHRIHcp0Rv1vjSVd0cHxojjw/+euujqjmkQEfEASUC05zkd9sJQJ+dkF8NGVay4fDIaTFp7TxfGi5N5maAaVnPWoM/eNRB9+iiUdjesvFRPsxecv6HlZgguvf68XoqHJ9zMMDlcPJBIK3i++Uq1jCtS34GS5AnVVvwSiyFQnyQ8IwsBSKGsgyPu6hCwX+vmn9IjbVEWyR6n7GvFl88Ua8CWYfc6VAuEWzXhGRA67xOnY/LeGAi/nYuvH9mAFR0RmEISUcnl3RyB8vhef3/4U9V+vcpjAUVuApRChG8tY0Tmn79hRGAC2wN6n4C3D9JRA2NBGi7cQZzy5II+KSB2BdaKmOF6ySBxeHhkf1naZ3gSTI3VE8PifFjfZLcrQTLqvIBmFts4z+5gxYSfxtntpDIR85/kCBke0HY5gjJBTHBgljbmcnFB5qh6a/DZyNam4DndNE4+w+d3ZbFtCTOwoKg0COqX7w+bqCxSd2e9l1dORJkLQILA1Y4CVGNJyINcPjg+u3gYM/jyeFEXYE6fHoM"
`endif