// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YBze+Koz1jP6caZGjAQBz7KcRO7CWG70GZbHHx1jAdFAz8fWvJ2lo0X1oPzs
eQj57nmeP7ZE667M1BZwltAa868G9hrQBFZRm0O1Mo5loutP8FBE+nNcLdIU
C9xgryhXE74mSqoOQZKbDZCkWVY00mesYrbJPDjXkPiDJoo1HvoK1N96Gj0L
Cb0OnRxHNadpCdB9o3vR3wNcl75L07ZiaPOmikl2ER2a9XO7nKT2stjydTZd
9L4j/RYyRqKmfc1ZbeTa/qnYJ5wGb97CqnXzQSL7G/2lCWDMKJdv7Ak7PpTw
xnd8Fs73P/LS1kW+pdT+0arHAM9HXm+ShF3I0Qs8hQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jy7cOIrj9ml9Dcv+CTtyfxf4tpwnFZ5eIXupiV8S2q1Zwy/erJG7SyrTupZ+
aiCn0FHTHdrC2wPZPdY2w271SuYrRgImkESzEaZEK/XXi1KDuokmy5BvnsQO
G+Lc7yDaCsBr36QB8JSskjFztWuPl34QF/hcpvPhxz0qpu/f0M95mYziu7l0
7dVJ4xr5VtHkn5ZKjIm921JggoiGfNoACqL27RGX8dThc2DcqiMUru/TH5dj
abdUOXsDMeRjPeVY9/QN85nfNC3VVhvhNYzghgL0N3zTDJU4Y8Te7Q0JN7US
vXAnuA56kVcoXD1kporApUifqDhkGj7XQVISVlWcvA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ilNfl7JnSGGE1C5wLm3OJ306llYu/0jWSy6AK3VZJoHvIQdpdxAq9wM1eAjm
wGl7ZODqqO+xKeYxm+hIq1Br6ThTCaCj5uWzdd4w96pLNo0i78rri0wH20ZA
Q5Wrm4mL3G4UiETAI+UStnkS8eN+mH9mJ3meJYCGHs7sK5xhFc37D7oK+1kp
87UCZAD1wtBre4XHWwUSAv+zFbwvdZkZRTERKa2gODsBoh4Zvvzqr357G4rV
Abnf0dxS2dCQ6+PS/pmjMwAt3yT9AWvXV2bQqrRlLNbVbzgCLeEFw8OO+Gej
wpB4yRkwJBEN3bkI232Xiedj2neaJgxfOesw5OIqWg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OwZpqh+eiiUWFpH9OHbGOkKdRxI/1E6YUhV3kX9LOfduNlOvZoWxBhzeg2eK
6IX94RGpkcHrpkISsNPhCgUUsUIYIFXO4LW6fIgW102cb/jumpSDsk20ZdVh
+VlfEXQfIOai1iXvyyUVzUwCjd402Zp25MbdhT3+f6RwRNGoS7rJZCxwdxAW
OAqR9zmr9N04WN9sIfbMmdHmPOEpMLKrAJA47sPVB/WeeVJVtrOYsLiOHCWI
OMZr4+H9sbpJy4KfGxA2PlMNUGiYVGMQfvtC4FkyfP9IIHUVkevsWebRZb+A
hj748bVUFocKGWReaUeenDfgBajWzfdcrY4DWR95vQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DwA48Wd83B7faW4qA1PuxYakbJ+xYWFvdr22ekvh/pXX1DIevUvY8xc4C60I
jPMCUh2AfvFrjHA+jtlMV3YARzloXp26aV8evZ097Gc+0El3QesfOkq8eXFA
WqQuoFBvzfH18zPAK0WEhXSkFqtMqPYHSb8yfkB5flEyVc7RPOQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
G/I43rzcR97VerN/cBwjKuhqfWJKd4Fu+01xj968PSTZ5lF2LjtZsE1HppR7
h2KVqJf4MzhM8anzp+g92ZfKwpIvgqOa/70TKpYU4+/3bBO3qQm3uDqbLeuF
zWNcP0es8CJpd/ZBtq3+tD/c0Zjz2ITHiwkd4u9XvGo5ZxNVJrC0QAnBOjMa
qKTJktWfcogwmFU/pT3PiMPmMj/V0rcM/VlPPAU5a5KrT4Xc/Oe7Q7jWcKlY
cqlx3XKkdpyZkf6oYnRFoiwYVD3Uj6SDKyj+QhE9kT/h/pLXYea7eZ2p2UCp
7qCjrTaQwF6MuIob/qrah1kqM9O42OvIybki/p0ZxkZZz5wD5Mjl2JrqwLMy
+nHU1dmbpl3wMhGESJP99WvMpETtX19JQI0zUd5GFtQMM0LOy0a612il6gIY
kxQa1vxF7QdcGgg8W5iG4ldsgLbD54qXg+PGFU2IBZOMy3igmKyMayDzqA5c
WLzEDA7Cnvb6u3gHNCotuJWVWaAIj97R


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K/+FigicErnkSJSMT1NVC5oy3pQyBbXI0tsfRatLqDPHRuEv7+MS8NBZYgbt
vy+F4h9sdAWk8/Dm/b9w/6VrKihLGU44H4e6kpN7nVxYz6OO462ZANQpTZev
iQkdBcqsea4oEc6Lah7IDE9b0vH+upCUDO+uuCAOqI6evvJa8QI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
guy3+koizwEzcTAarAHyaOg3A0BEZUHz/aUahxVm7HCj2tJo8EiGWT5V2YZ8
UYxVEZTEFFmo3sv4uaLtSGwJcr3Z/vNU9+XkPNpPgZvxCfwXQx2VRA75DmTF
npR51zm7Estni0SlB9//i/5RqFkv9+etL93c54R1nU7qhuRVwG0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8496)
`pragma protect data_block
Fux2W4Z5r6MNTzYOqCao/5h7VyQxM/yWn2759RsxYep1ARwaQNvQtivWOPh2
Mbiu85rljpOTVX5Rj6951y8AUyDbh5+X9AQKqxeQp2f2OM85yx0hmR1reYyM
5tC6FMZUbchD/rX7Op45pbfFv2rySvNR1BBtI8TDNsKKmh0XAdfyNyZTWmyq
zwwcNt9tMGzNqg+XyEN8uUDjZzpbsH4/bf02/BNpbF8SNQPDijKyzXESEkxe
06A27y9eGAxB0FCfxDuoL4Ky5n9uXoRXa+PrnZGwOzOsMhb5uC3GHj/w/Dx6
o4bxVaWapzmSqyS2dgrPaWkV2LyrfTT8j+3sMlla2uLhzdzGHLEXDYvSfMk2
2QXxTeug19r8N5w7Dur/9KDPS3OH3Qx3fpEWJCa5UF6kvIVHh7sa0AidzlFR
z2FBr3G0OaxtH2b1s2XWRjsrMBZZdSAAlO4y9JGqIBCZyREZ+6iD9Imz/EXT
nVC89zaS/tbyPfai9qVLErTUQejKRleicqrEWNt7LYeXYHDJ2jFqR5f6DSdJ
dSmx9kuCt62yY8i5Tcs+ERagqJmF01rnu/3MB2KA+ni1naQlPTlbGaq9Mt04
lYk0RrnBKzygkH898QOKP9prP082GLpr3zMcCIxV6rq8+MoepwOczqtG7FVl
dMyt5rSBSht8jJRzqnR89HJ3NEQQYdAIZ9NKIoKsoMA9wuk2jUOjfC//sn4C
HTHz+zCdLZkBFMxxXTdd/hd50knImYYMxFRSWG5UE6EMh2Sbm0RmFWPhlDim
hz8Srg6fhdl/CfCphv51EgW3Pa2rRrWCgtjPyeFGQVVQop3lkNpa9RJsE7eu
sK2BKeeHOQbXNiJ193V3ZgYTi6+AelBduwXYAlBQ4Qa9lBGaK2vv134HsJ12
txtQrc8VfDFx6uxBs0kqPuedb7Y/ADzlgGQBwCyBQTGjy8Tpii+0kF1uFYcm
NqWG8Lq6OBCYfECwqpGgIic4D4khiIHhn3tIX1d5yIOu+kWLOvaOkQO5LGBz
Y/kSl4GUYLSkbOoxrvaRzkp1cxfgGXRNr/afywONQWH8oqLROck7eJrABxpI
PHYQXXGrkd0Chs9kLRp6lqkHFJFhQghpvKdv2rmAUBQFaoTC3eTbXGRX/Yvw
+W/3G2jVnnpjY1KFwOPJ029OAMAWvA7n8OhOSLQUFsLfdEstDLVIkQqAuD0G
2W94z79kQ9ArYPzSVyMaR7aZoOyKqCYWmFNSMR2n8lQxDIA9HOUverPJ/FVR
A7IeosVGSHcgRjww8s9Ay+DgIVfJB2GJ3dR7on9KnrPhSO5+HP3TICs/5azZ
06diSU7ZNZUDGXimCzuWe9gJA6mWU4yMAwMG4kqAGekL/ZX5B10TWXb9p/W0
VmiWjwGRZAZFFvGBKN/9I1UvsirqZTXLyPueJbrHsA0ztRQ+SKo5ruzY2o1k
cdeeRPBrzfTQdKLpZedDzNqxE3jy8jR8CAGvM1qed4fogiektKQnbhnW6xXM
tHUZpJ8SirI0b9ui3t+oGbPZ+uFMh4s6AJmPmBeMv0EKOfo194dPVCJxiwUs
C1cA+xw8SQSXg8RYM2e3MGAcBaz5V04JqXZtItiEE2kuCyh9IH2/NN2P7woT
9897sMFdjaXtei2vSW7viE7MzTM1oJo/V0beAfTzamDgj9JqyWW4bUydF2jL
/RSuXATVUXxjQnI3s6mLXpkPVXbJINXeu7AjyPIDwD+rwjyZDvUZW8tMzZP6
3xHzbz7IwECeMFNXXvqUgnhD4rQnqpUbBg8iUmY1Fg8z0jcHRkznGRkwAIWq
Jgj+1IiOWzWFZpKEelMkCvfjeig45qMGWQfszahliz7QQxyPyQT+PkOi6lUT
+FYrZs+LP+zy4w5VRN4RjzbvsLv9XzXWuTz2IkHRNJwNMsiel6OFEtryJzub
BVs1kGOe760e6oO51u4CP4quZLafuB4wQsUfoL7PiS7jsnxwEOyI9v+bPnDd
Pccp5mvKnZhfdfC574caRFdV9+wwgk/4MTjAcquMXMLYSvTSZbkwhhxzQudh
6u3Pj4E13s2yUODpox6rt+CKXUMVIQLeFHczDSk4mGGriT7M+4o7xgU9WzY3
QXErcHI5G1i8PmtOKMDb42Sef7JzDp3sNStXysI+u4R+rkYTN9WVJS8F9Mvz
7bpVLeE4pYrsnLFtor0EZ/lkJP52uUUxZ0vq2BUHVPRG7rSudOnGyeS5y5LT
VVNF1cSoH4xlwpluMqF3NrWSkokPdo9AGqvQUcdf8ff/MO9y14e3/yNWW2p5
f8r7cOlAgQRP0hifqIf3t/p2ozfRCNUgQyZW9H+ipTGfLv4AzPykofQUf2PI
0S6EHN49+kIRyduk6jcqLFodi4rPtFNDxo1WFrZmm/VWs7nzS2OozLHNlCTj
eMMVTeVZlCpv8mppJm2MyzPkcHFEdUEKDohxX5TBHk4T/58gwuDzEcfukfEP
LuLSxEEtuPeHvIboCK1cZIq3Lav6OH8hNkQiekiJm8OX6hop3H+J0AtC+2H0
uiuVb4n6JGmlgxjCUnXedrYPdP8YLxUnNhm6Ya6sPIFO1+gCWdi2jV+K3oU7
OLc4DyeyDRRBIuPTwCN59HWpWO+yjFjz9EyI7ib5g1OVJvgSleVuGFJEG2w7
QgLROZWRL6gB9ZMHo2B5es2iCqm0IbOFObriwfwKzNxT6b1qYSn4AgKck5GY
UwbPtFnkjFnB0x51QS2DHADKNVz5sdc5K5H0jLT1NktIBRwe2WgzNraASq3p
osEn84nPSfqGF+ud8jakccmRhdGN5HqEA5ZzjjQd+CgB7FVB++YCRhhGDN+7
kZmRXnyBtkctq9mlpGie9D1HQ4z9LlMW1ZzC2Dl0hJOPLYXcX8DHkpUgOr8t
05ONuIgPdNAugkf8/nYHiYxGLAMKJODQ3f1ovgOcnvQAqw2PlcJAlNg2yVok
WK+Dj7rt9YmpoEtT9Wtb+xAx25uYl5yIC4yDLS6/Kod75y3EeIE0nM0b7rCd
y22O6SiyJ9MBcdLf1q7RlF5SMukOBEr0ibVm+7FQH5Gsq00sSy0lLQ0gNZP+
syDcuuI0ulA5XYBN5/7VZrwo1lO+7xLCg2ljfmsPOc+vYsQviQY8gYQ8mv70
tb3G1Hl1jDR9351jBdyBek0XaP9deTYQEQCocvnZysu+xW4GMTiyS/vziMkq
EgE0+F5g9xV63O2gHGnpkoRHdt+QanveQQZkkMGMJNFrZktarxvQ+grGoVLt
5g+hjsAMdxaZ8hNXyW2UrlZg/pNtscvJ0ZDC4qjax8hRpqDL2Gwof1weQ+Sy
cPjdMcFTo4iHy4hIvjeMWJGjYsdflfhUYX3rQJT5/REgwpxwYlBlvsxw3w1j
jJqTU/Ub+Z7QuPu42YAvB5ylKFRXszqKxD4g0QxQW66zf4OWZh2KQnmIpqHV
kW8pyexlvrcy8ZHjAWAkc8rOvJyDD6aewXNQUZ0rPbSy+l1HlOmOWyj5dhDW
d5/WgD51qssya1sQWe6G0B2kC5HeKszAU0f/WxmQO86X1oevyci/gJW/eJ8u
vVQBI9tnbSMsQZqYj3RCCLxY/onmDSlAVF/2JdckU5LVFdAjkFfjdi4rfyDS
ehHL+LtiPv97miKw8asuyYY1N8kwRiXEKHR3wMKplQWZpuB6K410fZ51KOKV
QhluzGXxILLI0BBnfuj9aDWIH78aVLycBMDDM6h8EGsbDRKYF2xXDV2fW0HE
/cbqw1+XRhrLRmSNg7NS1c20XqG3+t6cc+Co4a4U2Rx5fhrkuAGLo+7BbWso
t0hjM3ZPjTts3KhtZgp55mkzOwyO6neGBimebUb/al596245GkzHsR4gWPV8
YyCR7vc8troPUXPXoDyxg+qqWeAMxA6iJv0gHS+e30lxGFh+Y35ZeYEi1FRk
t9CNjLtXKHJRKsww1FREb6IlgMZFg1EARrftbTvG3NObm9MtLWzE87Kxgc60
JEjGW0xDSMN1X0AipfX/DSvr0RL1F8QJRfRt42ZT2ly7koBevaNuA35JZarA
+3Uylt9Sx/v8Mb3vVQ1LzmRjAcRilnMtipVom3zvU0Ng+oOd+Elbpu2v1070
KXgnaZd5sNLLN28FCDOf/M6HAgz/dwZ+Nt6isytYCi2apcL+BP+RLzTQ/zJq
3V+E4J3QpxFvNTI2SNaaQ7cyYTL40xFEOGpLmabWIJSsmgl9XsYb3pNxySGI
G7zhumSzvzCC2s9HLhF7uNBxpsevcrziUqC8YQ0n4VubwizQemPJxuJaDaX/
Y2XCIZF/tScBdVWgv1xzkCzS56LTDGFg5snz1gGtgFyNDUHeG2pC17lL1dAq
vb8Xh1RFgkLdy8/ZW9DRwlo3WJpPsHpn1gwIO+XGwGkZT6AP1BlUpA9bcVqF
Noo3aSDtx2vFCjcp7woue4o63z5venL1PwxDGdf6DfY1ZViPnLi0XRvJ6jqY
hv+Fl0Z8R6Z2whmDK+V7cdK2sPvia3cVW9NtjLtnQDe/ZzvNeqEGiYNlMb9o
7NOGHriXG4yJl8Qefuv/EPO8JStHl6iKULolezcewIN4KUS7pKCuHV+AQIGZ
OB92hRXuiX/hXljMXbFHmPPViOmmEUarz7bV+7br1vdlPgqmunt7v1kNgXts
npI+tOFIibgtt0e0fEFSvabwuJOj1xWIfgOVNHOcXX8snMWRYDqIK2oqakPz
lXyWNrtrE+SldisOBhcoxDfQJt7WQZVo0RI0osbIi56GKseiyrjmmpRpEDhn
oYh1gqX9S7TysXgUHTZbenevyFAiRVSahsyVDFRq8uJkfUf9dYtqkzCwbbgE
4FkknBlU6pMgQBQtkYjUbwfi4IrHLi+lbnyVrY4KCRr6DJiFHdktD7Lrq6+K
baZdz6yiK776UA9Y3sgaE5rOIws04xnbPZqq9H7Ph78/xbYZCaavBHuHEP5P
NNLYj9puaCCijNrq5CNFc4o/5rqe+QXg9+YxvW75EiJI4MB+uePA2PSNrsrv
GDOQs+PoARGyuXZW0Ghh8fh8C8Jd+qt+rQvOdzxAp8RSIP0RniCpxmt6QdXr
vyBssV8t+8yhR6BB+/TLRkC6FdayMvRp11StDUuH/C0fEg+ltMZqnLMOjHaU
YJqXti99vReCz7rk9271lg8RY16laAkkYiYy+NvRgl6l0+7VhG5D95BaIlEg
GZAsaP5c3kcyuRdDYxnAlF4I4ry6ZTsNIgNCmWUHBH1ekRHVfMZSXQaKjEoF
iDINlMzR/CzSU/JzMaxyYbk3kSm9YnNXfC3piZaycxwvHpdtThPsGnP8DL/s
f+f2hjQ0vxCAElCgqacsIlhBDL4Bv+5FzWvJfjhqjy0N81UxCeKMPcrpo1QE
bv6crRJV3X6Y68JHePa89YkLI5gAGjTrbs1aRSnhM983hyiNqzjdaJ9sUbmV
t1Ke/IWxS9kDZdvDpPGMFCtE1srKdLfEl2kjbqalldc3Qdcj4A9toAt6HuRZ
oyc87uZHNIxb/xrSlNByk4/3apO5Eyqb0HqQ8ITOSl7+w4mzAJc2Ff+Q1HSa
ZxJzfir8zdjd4ePgaGCqyDHBt1aqctyGz8zzSg3SLbNJQFvbEBSNI0+GwnUe
5DLiAQEolezgVsz/03BgSYK4qyzt54S6r9svZ7tNFlJeynfEwb3VtK3yhk0u
9/vSnntXQsT69XqRhQ1IRC1+2BaxT5DKswwyRsEP2MDYi8I3dOgyxGtIQWmB
6AgnSwKxWciqV+sPSfucQYbQxnlKQOcfryBeRPeVzsOuv/lv9V6z6e9L3VMV
vhn2K7c/kPsPrboMKoVwkNjIcW+UpYwONkp3Jz/czyawawBlxaXEWe+3KcBW
4AEWxqbwFGrYYxqUAxNn6pUKxlLxImcNiCx1sg/b8f7ccAMM8E/LoO8Y0Svk
SvBoX4qRxddHjMBgWfVZYhhZGKW5ywOxKm3GXQDhbMTq5jbety19wEEphINa
42z1GjjAnDvCl5QC9cLAZPZhCFBwKxXBgTqyP5y1B7Z5vp9W9JyNydAOTLxD
x0tGfYS0lk3PIGMu+nitCKFHYHEfuYLFC4QIiwfIiAvxV0xL//xr3BYVGo2w
sp04C11iqlf+gDpyd1MbPOMcV08jWxyHu1v1b2TrG+F+8fI7BlP9shWxP0qC
2daUzI+K6Vue/fbmINNjIZIV0xaX01kSZSB0bLN+eX9YxewIFueTmjXYaiI5
fvcXtBnDR7ZK/zyxzAQVmd3KUQW87D5EVV5sCwQZwtc71fTwN/PglpjSoS+R
rP5f+hjFEttgqMfmoLz5nOm7qRmsQ/8s7VJeI9jkydYHCbY242ronYy9l79+
vMBqVEUtuFMkfD9L9ykLsnC/6Io1bPijClxe1/l4/4O/GLcc2ewqywIXX61B
Z5lkXW9oQtsFb4B8Me4VOKkYoKjU8uwCBs+/WxEPw6MEI+yBgLLPqAoV9AIU
rVLhRb8JpRttF9z8YHvVX4MoychY9HG4FOvNoxrMouklNNbFExbyqh/ce1Wj
t12lToKgCtVRSNsJoT1W/n6cR/ufd+a0Sc7rD1uyH25cEuD2iCdD9UZaTRa2
Z3/Ob5uQz/XZJ1eiip1SbvlOTLCTjViamgi2pCbejfZHPMq8qxmz8MhAQwSP
3xfOvaQsOrugcI6WPf9h80ZXD1a3FUMtay9eK/99BE8Xx1kLOUTnkLDdCd2O
8fz7rw363R0WFax2+8s6OAQJvQYqHhdl3rpmdT9N9ZGS+UJh2s3mVzLLagrK
CvcH6PiLWJImoVobfROMEf/MevCT0My9gCGOGhPgdELnXQ+HtS2su5PXewkz
Xe811aK0gFp+cvsN7g2SF4MlhivkDrNS8kq2HFZjF0dzbS+/vXo1mChpGeRk
mFZNjw03NkObv4gVC59rvuu5/KwQDBkCY5PEJhVVODA7qite1joA7TXW8dMt
TFNxxC343ao86ONmCT5Zz6rnasV7LL/vDdjWBj2l1tDluU39HIhqPalunNbK
IohdzX+0+Oy3GYdUTuG6Ku9ZWlUI44Sft3bOoBwvd8BBLEoqFnv248bmTVl0
w9xlqmlnb5ISYyraasegqiHOKt1uAoiansWiDMwOp3oo5RO76L+agG7Cwexf
FEfJRj0h5ssOs7XHtN2yGqQP7SJJk3XsMtn/yCbUD3ztUaK+9JO0n5ARH5yv
SSRJRgfYX4+8yUmZFytkqJKare57cX/LLauEr/ZAwJV8Lh+lEFHfHftLESw8
Au4R/4S1/vTdKa09V0v/veOlvCfbW44vd1s0Hw7UqN24Xyg4GoQpJKjyQI9w
5SQct/7JN8zf5M2uBKvKxa1ysQwD1znDa5VDQTf23nftWlFdGLImquKBygOn
0GP7m80KPFMqxEMRZy8qRr3kIqOofmdq3PhE/xfVqhqmcj+rxyUs0d5F3KGO
zqyq4C9vtOXgjcTfrAxhqtukEU/W0u897zU59u8rUhLO9VHaV/coWpLzKBwN
qumS4izFMN4dYFKvSJMmmvw3f2TB8hgEG/E/6Dib1OcKeB5VJd77CH2YjkaN
0Y7mkb+HatzTdzhqBfIO/VTU+GT/mWw2w/TNa9W4vxO3EqngUTwNDAI2GKSz
v6pROfRPwt54HoZoH0z8VPeduW/n8QHshVM2fKXcebUnUhSZ5sxYdGcfZ9RB
jUNO7M+5eqXGTEiH92WGsfbitsIFksaMa9br5EhCJRnwvYRcDgNrlkC2lRbh
9MDDbcWB4Nylym6HS/T/rfcZGJsB9dFLjwDLFIAt+4d39fZw47IqUGJjvZRx
XZ0tgcS0SS9G+iu6WI6x7VeKsfeGFIT+G5Ti4Mr3MZbP3tmZOYFbNnoZDZOr
Du+ovWqmaHH/yvuxNNqAcXQAK8sWmhIwe9It2prlIdh6OFkaav3X9lHMoCDE
qp5Qoib0zp8Kwm7hxotah0W817ywIRAjDortGBqtynBeGsBxpQXdwzLqBTAt
2HW5sGbJ5NAWbPKo9oFUQuF1n5qcZgNJdsiNhVq+ibjaa+rTrTcFXiunXdRA
ZFx2zYdR2aQUZjI3xmYina02rPvSCzH4HJMjZWj57sgVjCDzudLjUbrOoWA6
/cjZNFaqGVp97G9pld8DtXMyA9JhIoMHwx2aUYzB8pn4I37Sj1oiNXZKgnp2
iD+HLjDxK7O8teROC2Ez1aequFMSTaquvFwGrW2XyPbb/0R4ZI+9ne/vY0ES
/G7YPb4O7Jv6zoPAqLfIIEciDnuXbkdM3KhVL+vA9hHWlGOF1JOMl1GwpL/o
XaDNcHwRFFkLWtyMcRModkFlsFl2OHdPBUzhq1qFo9C6tU8vfyuZXb1hO8w0
194G5eZ4GWnT/FWAqmTij2BV3lu7C8u70yoIs3y3z7jRveY+2AyLTWEfv/0e
sBuGjUvkQan3SwCr/DE8SghuGieb8QMMltSqslrbjhSt6OePfeAm3t/0nUlz
yiXHGP0+FdPnizJgQS7EBE7VQ+f+TdlK1CQfNKHEn5Whg9jGB1fOmz4ihsc0
kjLezFPrSc9GhhKQnjg3I+DiJwm+zdljgI+EaitMt47baD2Tdu7I5qGjki58
WDojUaKwVdFB2lnywTjEpD7/sjxmqKJSxL14ydZK0UuNR6S6nnsanIXK7zOM
GZ+AeRh768VLLHXtRCgU9/SiMJPcetcuxqzU/wDdTV4R8oHIUAWS+uBypUL8
GQI65yBUSRevZ3ipGwnCvxunUJvrz2rrB9u1SR+q61LWIK8VFegg5xyqvu+q
jvxDDJOrPfL6w658QVuyoT6TfeSdRfGCQ6MjjY0mSpoXo6Ur+OUJWZBx7eR4
KbCqoXcmEYKqfHS+8l+VpFVvgHARFW4aXrcFrKvpdCzaNcNbNpLdPNZAK6QI
T/DL9+JGtyo16xUZFXt0OV73Lhj0o3DS5D8FH2MtU9QORR5E0+IiLUd6SfNM
gOTRUWM/FnYgkOs1xdMUp6M2bTtO8D7FbJj2c1kDLQgPWQVFk6Trv3IGoxRF
RPAoUI0TLmG+ZAsNUz30Jf0L3wyqdAEns36fSVQpcrIys6UTjuifIwpIk2XX
V+v6INd2ng1NrEQX50ji7cKXDUjwJsa1OxufvSop1JTJat3wxtB2OXJwlzth
IkyBHIzwnWYI/F4i93Ke4tq7ChKusZyOSpId5jjg2sj5g8It4XS2y9knTL52
ELTaxxrWi+HNvFnMAoQiSh3Pjx4V9FXx4Dko9HFG0n+7Radu6979PVqQfmxS
iU+b00m2xd0H2kRx/k1K05BlDbJd5oR4R2MgmnejSqdOHaS9WAJXCcO+KPjM
upwzpEI9cJfqKtRzXEMlNVmEvLBkzNRmzYUz6LqOHsxhCqt6pJudmRngmIot
y2z4zyGmVuOmIcJxEZut3/hG8oLamjNOIF03AjdSHNPkjBXJPj83bRpkwPTX
L0SKmqm7UyipVEuE2AO+4DK8mrD9zJalINfcmTWpAk7fA+zIr7Xv4qI3oB6S
0r+cr9bVYG8oLj5QNGg4PMHMQcc2IqGPFNvq8/Og6Gus5QrWF5qy7yiAeg1v
gzYeG3pKI1KakCc6gYpNTkGhzP03r7nobgmWe493UaBBkw8h6aI6yqBKDknL
2KoOEcHgweI88YcfwLJWKyluksbipgFrY9mFxwM37+IBKEkkNO6BIkKOb3cK
0BK5xnh/7atv+D5I6F5ZqJtx2WI65MWEfBYO145ip3nkTEVTovpWWz5cR8wc
CyypnNqvwQmY1Rf3NGiTiUtzLGf5fxXnTEE7PTvQfgaePWl+Gu5hTuBHU9u+
gJYQVhH2+SiIP5YoFdSs9PzpHut7bFdXOHDaeEWOJX/+64DdXwQWKbKisjnc
V8y4rbZVnkaNMr7Jjcj9UPJIh+pfWjh5zbqq8ZYO6EH0zeTtw2SJzUw41HmN
/jwi2CJVz87QihDk2LByLRYQ1e/yY4eCZoab4ZjCFiS7tXgw+xCR1VbRZ6KE
npFnEZjJowOYwlBzKspO9dppWH+YvBIB+fA8hcKE5EZ7ZdcngV7zyABlD9lx
vnj1o2SyuGxA1e1JluaGlCNZSXdTJEoPqS4aZdojHHxpSRbgnr6Q9nf5Iyv9
J1yafgiXJffAKpZf7zfYdSaTrp+00efKrj639CkWZG5VlS+QN0LJArvTa4AV
fp8wXlTtNsbly+oxjqFgW06LjTHFC9eLlDkSbZhtsAf4pK+SmQMMw+hT8oFA
lXuluUrrn6UYe7EiZ7RQDEVEofTv+x2v4dujia5tt/Pq13zPkdvgUHgIToNP
LLYVy9VyZGE5LyF20XSH0uZsp4odgW9/gf3z5IwAGEIKqwOFqYUEXSzMZoQC
P8MnXmcx09matq9xkUuFGtWYoatcAG6+D7+RzjCFIaVjIfD40iCvqZ+yBGaL
ByS98AR+hBgb4a0zillHpBQhsrJIccfnDBd+yw2nyQ4OzdraHtQ8cAcjEleC
ZSSuaf9KKskrLUX7vda38JBf3KxXoDYOm2znSpZ+tOOhXISnautUGvTOdjPw
gVPlSStpvVcOA8XAKM8NvUughJkJSNC70yxHIfSTZ5h540TD3+84eYnQDFmJ
BAAfyuU6uTHdjReXG6a4A7FBPDGyGCPG9MVXvW7VczlWepRQf5eEZu3GhbyG
VdePzeybR//JdT+Ma2GGt2fXlXVQHzI6MKu8ihyCoQE7ezWG9XvbUkx9i74T
Rp7I1W1rYk7gLWqHfVpO9lC+dSrzAXORzpAxQlGvFRPx8PgMYJJ02/J4Yq1z
prk26VoJm1HXwZnUd3YmSYvZ/VGYArUMfT5SV8gyVTRiqPAcYvQzgV2RVuFn
LIUKNPdg/eQOMOEUA3aWGt4OgiWWS/QvNVHOm+qwT4jxuk8U6grTqmNvQBEf
3ZZnF44f/Zfh5YZnb0a9CsIat5XS1Sk0WyoCBn4iVXHkLH9cR1hviZa/EbHw
XkUkoEFOBoCKBsQ/hjXAkYIYJva/X9i+7X5LAr3WJceWDUd+Ny7NZ0xofUlh
3bc8MRdyqY/MZDiMEC7Y83S5thp8TkZoT+yr80WsvWhflNkAER60ae2lUs6U
tzARHyAT/6Z1nzTrBUg6TqThwXK/K3SU9SV/qceKqk1Pw6/QVpi2SJtZUatO
MXbJpTQQggzxfONqJ6Zm606burY6Xyg3XWBNqPLW8f4tTL8GyS8XJKI2NdVw
fk9d28vBIcvpb7OKIyX7xiC8dRMV63GUFYj9WqCnidGpHBZiig3jpTSDmQ1R
JDTRFB7b4k+hxZQJgTFEHPfp4GoR3MO/MtdkTa9AIl/P0oxJZUqf3larPNqa
nFASgiDJav/Q9cKs82SpMvco+lczT0xpUHJ56WyCqq8jnuQ2xF8PzsehZOGi
SmiQWy29+eDmBvpZIYzCvWW+13HqqfXInl0gDkG0kkNWH1oO

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wi2ZErOZWZn8z6E1IHo5+bOcIGFFv9StacQZVReoiDJGtM3bfMQQ6JOh4A1u28ZN/6nHa3OtRm7noFWHhbSvONLJcABd3Y4YiaAPXH0BQQ7ByE8a4aFdadyZfxxk/uWEB2/Yp3OSkYZN2aU/8OurYoIxdTOWI6K9emjYe7Wili9A0kzoy+vT6/HDTw4OLzMFKcgJLaDa+4cOsNHtPqu4Kp/lPlLE7oRIaufyVqAHmj8bjUtFh0MCFuKPnp+tEdWvMmUmJgCKJLP5FzU+nsi0CnDwxpzy42C4Njqhp04OCpgHOPRKBAc1pofOUsoXpmWU+/3F+OP1GdlzBx1YfxcYMC0/DaVEteZesan6HMhaXAkGv1KZHjjLwiKO0Xj1HL3dh+nPogU+zIm6PDsf17D2qFeh727cOgqjstbi6mHsYy2tFOlu362gdOUuwK7aMkTekoiYj4qE6+1KKz/KwNjv3/P3aK1W7TJDStVsH28uF9wctdD088Im5MaiWAiwcdyl1VJ4f2RmkRCoceW4MZKEhgDUKl/jvS5CsbQ4no4mnY3vIHNqBoFytSRPdmJvtcdREB7ymDS22UkSs3F8fR5IM3zFn0oyMDi0mmfjF2Y5ogEZ9s66VBrtRGtBEmsiY6qAdsVvM3JTzaL8W7pS1nEOLCMX2hn0usXzs/erjs8JK2q8t0SKKwde2/h2N+ttHYjQwMDl51r4q5qGe05br4umZMQhVcanEtAxGVGD2qWKFH51dfZoUhtDepLu+s+V9Vg6VkZqK3+gQxELyxn7WGOORMl"
`endif