// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dM7a/Q8MpoJ0cngFD6WjMruyjPg1vyUzZeSXMIMWhn2r9hNi+WsGsgpz0fs0
QbAueG3u4YSCnUoCJ9VY9GHGVGvvWyjs7r3EExPzacoBenngrABBsMs4ocwt
XYdZ3y1I5TeKr2DCdUv/p/gxdHE1e18bjzNmvM5g1znijv42PgYIiJeX5WXn
OCWt+pqaDez8V8aze6GBoOtu6+gkOWeLWnJgi4veNCkEpizUf96XeLVCZQ0M
HgBuMbJqzF3T0Eh76UQxUXNnFmBOJQXeqB5lYQZe1H6OX7RtT8icRbgKF5dx
sQ2GzAQ9mtHPrPJbu1xQ2tpg3sJpdDdE9FLWNaZF/w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m/Ov8laEfZi/Akd0vhBHokhnT2LspLrWWT4/lqTyqqDLTNKyjlSPwrIa+YUR
jP1id5hqVS5LJIWFQoYubXiEZIJF0Ipb8zK3wUIw2RtAdFQa/lkIpFydPc28
8qPY0dtJcU28nmEyQU8r7TtqP7IDOQLwgbCvqs1epYwqbdOUlGCf2HhmwjqH
Ra+lKgWZGGFfpvGq3/Bd4cQSg7uzBNd8pJnuUBoEXzxnJMGdWDX8fNz9IADV
OTQwmcyPCJQ/L8UppvOixgXurj6XfIJPYfcr/lHX+xmejhLxendTtW/E6UC9
FOFe8AHTaY8aoqhtyP5sg/iC1+75uqKOEkSG9pxEww==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZqgetLrlBNeuN3M6A8TxJByf87Ng/sXW76xqkTxp3KlyOLqIVdBCCmTXMYx8
Z2tjzzQEv4ArFrjbNWCF+U3GTmYpLhzLMtTOpW3f2fua6AB5wOxF0U0ZezJ4
IOUjwluFXUCv9XWFTwT3y9g1Hi1KSIhqV29wXRqdz+4pIPJvf1ymVJG6SIjO
dmQ48m6iNtn9nJRegHarHoFsqTWRlHuE7TEOpC3LGjTx/koYU54WztbKEV+Q
aPAuBq5pFcTPdujWhd/E9QtiWRCBzMsqNpkzy/BD0oc+sO/YHRhLtWKgoFqn
xxzRlnnAP4fUJDLKcg+lXtYYYqR0h2fwXsWJxRQEMA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AUt21ZN90m/L01vvH4N2b/3we5xBRwhLpaeoG6s+vbLWM8D7rqrdh5x2xke+
irNwXJeLAPmHUeiig3UTI3YZSYQwroLn+Dq4fNdo+mNlpvfw2cTHk0yOJ0BI
HRpZLvRje7kKivYUUzUVxhlXbn7bMVmomotYrcOQWIdXo86aZXaPby/rICLW
zaIBkA9Lty1s48fr/0BEMyJmFa9dbSMHdwpEP6fj2c0+XzNP6ZJrfVq4i/nQ
O5jMDFswSfddy145E/oMBNULmxqtFWitnQB+gTQ3EfUvY8Z8A2BLsWq3Zi+P
mZBtfkcZJ0XW8n21hNu9+YZuLzNSOBmCX03F4bunxA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qmehz0Xw88tXMY7FOPx/DxxMiJsLYJ9tRk05BkhRsY67LWDLMqlXkSo3OUgk
zpAFHJlfD25ILl4xYlI96g7NKDMdsR4eAFNcmly7BGycgNghAB1sTRK4oAX1
WlYpbrlYA+9xSBfKVyZVg7TXtwRFPr5iiWht6toiT0Y9dJgkZno=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pTZbzxUXkmERUCdCfD9PALAjIZZGTSVEnI0/90DGv3JXkoEJ/tMXcQF9vpBR
iabU6FbgbkbuaKcZVqg53+X6NA2khcm29uhxjf4OwPUnc2/0KHpD8uiA/3bx
KK5Hu5Oe+F9JwBQzExOA4dQdfCLcT34bfZTUQ5+5u/odt+zyJ0myEoNhDK1y
Z4GDG0myFEJlD4juhqySE7IqHgOX80ex47gTbrVIarY1JkVvBqeQY4+73i5S
fVYRgh6ymoXe2X0SYiKtY1a6lGup697waogm0CX+SMvSgaIbhSxraltz20dq
y78gaERA/bR2tRZKrBiUskPJmhuvuhtyt6XwmvNoF96TRmfH4yxSHPB69dse
xMRDndH/td7cpu04sfR+Knl1V7KiGsfXKI1CDE/wS+WhfuFUogcssQ52nOvN
eL3qlxxGkdi7cv0+wYYtpNToNAUniWGjG/x/8q4K2RUx+274quyYRv9heMrz
WjAX5LwIsR4/J7N42OBS0Xub/bIvvPqr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jp68/GXJtUuYz+mewyCVhPWU7GhBk4+Z2RHQH0poWXk/iO1Tk4RgJnNpeTS+
MQ3jsMsZ2pDF0SDFDQX/32/14VcVClwOZZJ+vKYQf6nLxDd6gZZ/pJ2PhkIf
ov/1O5s/CtDqTOnYVseRfMorePlzTCs4X0nR5xBkFzCHpe2J4b8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iNeIPqnGSy5HneeUWQXh1jJU0ccNfFXYQR1C5Rytt25qmDrCgoSlalnK6mWy
eOylTBzT2SZ3MIoJuqxKjlkX22bWqer/mi/Jl+DBlCFwAfurERJGOXd4z0Zj
FZb6AYIctH62ClBff/b1Vo7aHpJaWV2TiPP2m5tmnlP18/CGgOw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21936)
`pragma protect data_block
+dO3TdbP6oG7qwgg3xreHrPbcpxQoi9HP3qSM4LP/RQbsQtEL5oHBQNH8A5R
cL7woOIj8ZttHpn28yRYjCIWLW+6/vPpEmYIc8XJNKQPyW+vsTeKP0HeVrLQ
MSMDW7i6vePIN050Jc69y5m38dEIVrRX2P2Ry5tyD4lA+yIA57SsaD96VzXT
990MxCqOO4Sto3QaI92KdZrzej3KZkRVejSEhEifmxNng+Z+/1KWCBFwBBDq
MDoHPEMdvm7LMf9GEM7+/0jGKEFuDWIBpEGE3jikEuPtK9llMDAyVwcPW7wk
k6LzMiK0ZWHiC/UOggJT3wN7stulRhUVSOuBqHF/vVcOe4komFe9f/0GHFuY
QPWzfrHMSv5FuzXcXhdpCUwHG2f1ysy8E/4KRa6uUVkQwaeDIbT8aAbtT6pS
erlRCVOQCIMixk46MDvA7g/IRqYqLEa9MiEoGaz2NHikjQwMC9Y9zINXAIgH
pJwTzd6Meb2Bd0j0P3cTZzC2fCDU8wsHv/RE/aghPe2QkYNtkcxbhsli0MB3
VWYxivqQOwi6rYCV2fqgTVxAqesRA6C2ovWw17cvQYyk/cyvB5956Kj953mM
ShZLC7vGMD+9L2CzXFxOI/pAlcZIhQSYPwFA2y+6ZRtWXNz/2LFvugacjqS+
dr5N4ecnFvh8NKKLDQlmYq3UtUAuSe91u8B+1odQ2edJJNdTjJgZwUpmrcXk
CRfNBUwv1vS38lcSNz+VQvGuN/9hhiEJx56BM0ehfCRvsUl3LNTUHsEHgZVR
9ew+u3b0V4R8uIByKD9UtkPvWdLIq6DAUFI4as9gTozWWHAq9OEKMR9CRKnx
2j2pfidvg+gUv8VIFwIL/MPCR1qXNIhRAs1enYffhemTthanJ4x7AYkKN/x3
nybiTGJrdYcW2B61QFZypHhI25jLsgnhC7k1zullDbdIm3M61UXwa2wU8NIs
N8eBFsefX3hD2gdkaGOxsJ9AJBY6h0GYb99NegM+wQig4x6NwYRdr/O/5Tql
gsVGpuoM4IbgLDAvhfOzxyYovvGGieX2G3zsocUAXpy1q7z7vAhJ1TNrQFAt
1/LFSKBBTYwMbhX8VS5jf9PlyokAQ4jXT7hj856dxRZzPRf5aOXUW0Nielcc
FH8VEfQIzGyuYkNpFiAFggq9X2VrKk8HDkDyNIO1xzvzjd1L0OBmncFizJRI
pIpPGulcBLmEQpDqFS5njOLAzHpg4MuQ+NHKPkHx3l8jpFuCefq2vnSqi7bC
4pCOhMWn3aGu7phTmpEeLz5lIMdRnY1Go2zJyP+1c96j4G9W/t7CPDd0mLLY
KJlxthmmwDTeIyFX7ns8U7ubjtozxgWq2Rugl6rdO2EbNaM4F+srWL7KThmt
aNSU8jW9E2KF7TQ7fk0thEEsw9Iqxb44+qnX1jNes68+CIHO2YVksF5yrVcW
na6rtmfH+tZmWD20ugqobSKYhiuFPpPWVo5Mj3PRz8AlQG/BoNQaWU/w+i3G
h/uVTvk1SKdVVIXXZRFRW/7XHnSAcex+Ik5dodSKER0tj0d8GHEL1YMM10b1
zO1VKeSRsgmR/OegBtS5vOVKEdRrIJnyMDBV9IXajXBgRlqllBaDrCdKIJkQ
oouH85s2Q29Wq9eeGUc3ClMyYhGlj+Q+ORpZ6eCxzQK/3H1HzlWxJaZktlBA
lg+j2u9yRC+idCHma4QEKVjxokk08g1DKXxvDq/DdvrVuVdmi1GZq+RxpyF+
dIPv+gBYp6i4MTkZavwALcGwoyTJC9wH4PdxSqy6V9Ia/LAOmhcfQegSq1Bj
JORzvYn+F/beTDV2ZERvCecIaQGarUQFX7eLDX+4wu4pft/qkHR39781qNDr
bKLqBZAAEdJRElvPv+hDbWhpXV71U/e/SX6XoLDZUDV1zZoemsOdXNzpZshm
Ktd5VDSg9xtq/cKy0hiI8APRfi9Gg4XQ5Oj5EmO3O2sa+J/1tw3TlnpxfTfj
MwJhKR0QVUHmc68CwO3r4dUP1wW41ivBCtNrsSaXhb5vSsA5+Pi6aybuqY7t
+vmNWKFg8L9RhHKKsIUiXxtIMAhdyfhGtPBobcp3hId7TH2nvspyNRQlJfHs
8h3VMp5Tgpsztu279eUpJwejRyLKx0+jcDUvsj6mJva1DClmxNWYBwCBMC6U
jP7wdi3PAicjkm6LG29Z4MefNykD17y58AdTiaab38a/kEutIpyq9aKKqO8Y
vmV5ivlTQu0BUpPmnrQz9r0q03xzpZbAKM1r4SFp3p6tmZgWg8ISXjd6vpY2
zB0FiAsJTKsVlyXnMIqTb3/4/q44ab38WzCOLLOaRb7dgR+koRKszxbQxWMV
HW98YLsj+eLeDV6jV8psOPvNZFNPmWHC4N2ak6vFLcLXBrD75cS9c9sckkqO
sOoxX3xOQYNs3b8Jk0RDd/ArxSV9AeV8AqEMp9aDtuQPIftET10PYViZX3f5
Bsi5UsGNosCRoXBqCJ0Zf2bG/TXFybb3rPM4j9+e6BREZLosR3bD6jGKoRoy
msxXb0oaUd75dtj2Z1hRjp5xBor+0s/i+EQi2bGiDMELhcfKPKG6/zd3L4pc
IMK9OdpNQ+Fr2YlmbY8/DrG3t/8YiwHDb6aoL0aO9Z1Yf10wyv1ZW4O7tGb5
M6Idu0vW5VUK2W8OxtekC/trxvx0RnBwRm20vXricMPBdZHYVK1n3r+VnfUP
A2PqbM5bf4uVsoy51u/x++oyhiNBDwCiQ1vuIUxICzmK2TbYLP1uKx65UT7e
Imz3xbavsFCUnzJHsyEVLNec70BG16+F5BuFrjYnvtz122J7uminS73m+JEs
vISnjwRDbirNnRyskZvMCQ5PvXtdWXkUev1OvqGNGxt6vSfMRDjRVDhBbMYc
SSX5DyqcF4+onJbMBq7e4VjurNJ4UAJAE3rysSIxcohaAhZuryIOWzWx2dTz
9H7oPMWPSmUZlyUcRSFyzGxfYZzB3jGSGKjsPQNxMf178Uh6tS9tnVvtwsj1
l+S3UuVNBx37vsgLr1cSsS5ZL+HcN0Qh7HRVDIHJ65twBuLHROY0FwOeRxVr
Iukjx85cizNFOd9CiRRZQlfK7OOh9XIh3nUSU28o+VVSX3cY6cw1zXm4kKwA
nAkjbNQ388GPcpCGwfIYkBjEhB3NbsbBF4DWDUsRORnFDl0QdmS8i/yVCRVF
SW6ebJI2LsXBpM2yvPSkt7LXUV0N0Je6QqAyF1nXthuI07w6lYdLlnq5+xiH
SSFM4CBarV+D0Dl/bm5k5myFRN8s+AVqeJ9mGMsq0UWnIxX0J5E+DqsNrshO
kW58OZl5eoGh2NHs1s7lCb7cjFEbcfPj6ZZ+01VvGs4bT+E4Igl1xpMDXfYt
Z//VybJDOhzKEx3GczAREd/TM1qLK/+EfVk1hcNkYeImg4VYZ9yuPy3vlEsj
TKSnBV+kJohOu/pjNXzDBRVK1sHc0QHKhfpDBpUisCEq8Q3nkmuiYS39LCBW
ed7dMtT83HVPKqPiga4K5cRPo5QJo7OdMNAOzqXLn4CLDA0CQNV7VHyqoIgL
/a/27w1q737YLcx1lTJ2c+AuCxauq3MNxKcatfSdTMEfOlDh8GtyO9PfXecl
ZfG3wfWXn3BWeqUctcgTMNMIHKL84aQYI8c4vnT3xCPLGXCbOOsjqmvYPP92
0z9GRyhwr+VtUU5J7ixKRt6qIwtfc9NqIhnSzqmr6mHqfzhh67G/msEQC918
6ND8aYAfIObA2Kbb2J0Eux9o8YhetrqcG+oDAvtn2IFpx6IkW5eC5IQOEukU
pn3dyMqZVK/1sO9PC7yfpMHcmw4L09518P0W6/061Gl0Ai/hbxXXmGFXSwZi
phFDgSlZHq1Bta/4d+xCCLM2eQf+L+y8NqtY7FGDrCnRLFE2LlrBnzduQSSE
9RxVTOGnpw8Ozu+G83e8I1zrqXoUQyykFwBtJdU8Y+TmtHrioEg7nV2EHA8M
FDDQQ6pmcXs0RQrcJlH87AVCFF4The2hrk1KHh1BDGnUi3ywajQHNCI0N7o2
P7VYWo9nVkhxiKa54u9xIIAtP1r4zkVa4rqSstM9tTgPjSjaLnLbxC03UJk3
c+7HXkgXx5G9XJfBwN0AyiM6XBZijQm6a9iUyYJ29HEQUAD3tO4W+FgL3C0W
gS6bmrAtUCxOQttaNn2AzQdapjTAAyNf6jiti1B/ArBrnYbVAwbYbWIPnFiT
+c41j1yZUlLzcBCkRDtX5Edc6CVPHvhog5XZchWTIHAKjlhIoZQ5GLhiLZFT
kzD1xIUaJGSE0BTo7XLdI/3W5bLsk2nsoaH9Gmo3mncu4iF5B++mpcc/h+eP
0EQ01qXSYwqFlrVXcmb7m7jxRZyS39EYqVFTTEQSVqwbUZHJ/xxEihOFkx8C
Ifylvz8mOKi/HfeIZgpn5oCf/jhvAE9oB+H+/CTDG79PYasAZ3kV3K3t2JxR
06Jh1n2ApdC7b1zDj+O+jhE870Z52EbL79XjV98wPpou9dFhJUKPkh7Ma13q
rf2/VI4bnJVLstLSJjbsPd6/zvKeynZQBxNdMLrv+0A5PEch9+tKJqd7BWRq
Snoco8NIVT4K+Q85G5/EyVH2uQI/hekUkm8pWPfIIWqp9qvcS9c+HjhUsGQM
85Bdno7UO2jBgIlKPR/H0mOxsQGaj8WkOJ4w96hznJLzpJk/+sJEZVWlGj/v
CAPKNB2M9JEbCQA+a8uZJSdLsTbN9oGe9uh7dy8VOc9JypwvUcBlMv3F0/f8
cuhqKBLxRTyXZxkh3opJdFxJ0AdBrSWp4VurcP41HTLFXB1o9FKYgI9dlaKF
gkAc9o7STRW2H3zE/JPvFMnOYfKYUn/bQvdS/mGyuDRRKOyivi6gt5p6d5Q1
WXg0RP5og3iaCXjv8YF4NHl/WVm3YDLAw7gLiUycGhVhglv4T7YRHcXvhhFB
E9CQB867fcgvK20I116ESfHRN0bqoa9XkOSMHZSUFOx9YzZrq6EfzkF6xqQm
QLD5ru//jcDv0amY9Pk3uJWTSNC7IQU8QZZduRz+3mSYAME9kgVo2mfvJ9qn
8bAEqDvzS82FBpVRxo7+d80Zo63jGofNg+y8DDW1GrOSpr4zJrMU5uolUzVW
FpICAEjU7Qm4xeF7W07XnmhEuA2TDHfzyNxngGrW60lA+PvLWvEQFPmon6SU
VKGgwnMcNqdvl7zYLxkwEJfyGDTJczkp9NHlwXPeTAPi60Ujz3p/BO3QR2K5
fC40vtw//jtU2mZB7UZmzhaCFJobaM+B6Hbk6aiSv1rosDoFUq7VK8895ZFu
Crt/nwozQmViPmLZc1+XfTmxDHrRSrqfHVMiP2SCAKUCWWY5kbp/0jIQ+01N
k8lVgCL0Lik5RtGe5eN3FnDvIEqAtGVSHRmZb/GC9rWfObvIazJNRmP/ziDE
7Sx7Ln2LM86dHmhCGKnEJwZZ9PKAWiauEPjVQDghIOCOoSuVkW9iA0Gh71tq
GLrxZHafu+LcXV7A3zllVZVJfSTP9kvlCkE4ts7UP7mEnO1wqpMXypyqTgNG
ak3atPnePo5JMSTwxhJnakFPTXrVEM88l45ka7dk0FP1+UjuYc4ChAOYxkwA
estRC2V6296cdEGIPd5v66JU7w485rvDlvJp/B+ZlyfIup7JSX1TbH/UIIfA
tnBx+HFSVDobUjPSwbsdgdHvnGkJCykxgOiC6SVDos86xGcqMjRxnYMk6D+y
JbsZwGXdP+B6cVt4Z4C455Tq7VXSUTv8JNwE9tD297EWyTpWKhEUnTOSPF5H
fTpaXGVnS5d1yfu97VhpZChUILYmu84x5o+2GdcMGSRCombJ4qmRj89tdPlo
XyQ1sRgOOfo5uGC0EJO5gSPnfo8tT3A4RaJ60PJ7zeD+kaH547dyBrVIpf7R
AzKQr1S5YCf5F5ZLLQKMxUBboOvvFlKGXshPvYKI4uRfgVUk00NBCpV9wkqP
efa27S8PIdkR72p7tXYtUFs9/FWi9IY539kt4S9zAOGVBXMjw/ctY0hFGvd/
NLiP/mfz3yY8alfKuRS8mnnHKbghKPJE+LFBy3eu01XP/jyCEw2EnWiFWTM/
D9kU9AVKfqm1QrnUexQafR1QBt+hElyFRRRfdaMDSs+2zfJzUUOZ/yFvftUo
9FsyybHj68oRoWl+o7huKmSuN2A0AGSfrhltENi1PMeYwEYaU9TLqXff1JU6
AmeN/iT4yT8N/cX+yUlIi9rRUVA2tK/iT1ObWD+A4oVo7FVN+FneLkcPby4r
uEAJpG3EwKHRm/n7j6Ul1MRCC+fGHBcD/VYDE0FW36f3uH2w2YobVG9aZvYu
kz7JvA1LfSukldWNVpAstYFcEsWmDeYQr8QWHH7vEfxCkzn1lv7xIfy/4/ep
y202LpiBlir50XOf5Hba9nsn4QLn+PGWq4ahz489Z1vMVixIOg+lko8Hj1JH
Vptctl11HeqpzVkK3NqswCkFP43u0nqorM139ADZGkMVtRjqwCoKqK8jX2+b
BtWiDamd+F5MZpkPBbvwh+sd5v6Supi6L0TslGBN6jlnA9Cw5eQDteVOic6L
2d9oPB1wi+dXsVBQgpBEpyJgAhIE5PCj961cU4bIoL/nblYV3JkbW49xXEts
KN4VIsOWabokTPVPvjJGyLX0mv/qxGwxHJ9ibouMLRbttRhEzdCQ85bGUROJ
XBM0KGMhEv6AzbOHCNghLG8u/IDXCxlZUNla30vVs7rsbhC3GLxOh+VVl+HR
yC10+cpjgw1agIsXk4OW8wXMVN+fchdjMcWIZHuLDnoHjTNgWJCForJD7BAH
cjR8z3k53TOFMtNApLxK6ttK3i9bTocuGYmPWX9dky+pL6HtRpumRjZ1gCDJ
j7a4J6l5hbE+U/6BeZCSIvn5YKuWnYmntayAZnKK7Q2NuyKOJex3QD6JtLnu
yX5OQtM/Q4g0oR1DUjGTCf68klkiN394T+fSVVuvXmvSztCAkk277VmossT6
3AxxtUGplG6lgnn5mPCn0DT3LNiR/MGBXUsql1XkexOgII2KT9KWWOgXdk7B
xPsyirNYi22wWtxshjbhwSUO0AB3cBUSWwP952tX96JE45GEN3dZeC1acBNL
wSmtnpLmFPJnQ4I8t9GxD+Mnh8ZXACGs3uUC0YbK1WyMOdb+hSKSJ5inucfk
BDlB0fIJnfc7fp7O5VL4i3BTBIMGasNSq5HRU4tYCu+t8jbFlcjCfCItwD1C
uZxkuxhdZnsafpTLmr2iODjcXiKIpvBcshOdVB3qGhIWYR0mO+W4B/zBfV4r
OpHvWMpClPyFp4qHixinwec9moHeHklxRNRRCSFjdPatF3+1qbqS3PYKTEjw
ET8gngB5FWdK4ADYZ8Otqal9xIX2kgGOaNwtt4wX/mDcSK87tmWKiOsuKPOM
mXKX9KC5Ud1Kv1RRUJQQydftKNQ/8IZ2bZFl37Lis20I7ViQqXc3xIoFfx9J
i0ZIY8NKkprLx+4prZF9/Kj0j9ksPWgNAfhN+VN6UC/uDZZgJfZ5EGqb1znx
MOkYfyayNdFYbAYc7qeAzd2RKYayN62LRaX4uMzCMG9PwZjy0cKYa2sLhw5S
w/SdG4a1qyS7sLGSWECOFOUaedxPmO/WR0acaoLvrIqh9RIb5UY8QJuk9hOX
fFnyy6+z1FehYn8ceN8mFimh7iZkl2LqAJdjjjw8q33ehbYnLCrrmUZoYPRS
T6gHXniUT0Xg8gr6o4PvuwgPn/nQyDCsi9KP5ikZf/fjVZQmzZgGN3NsoQcM
OOYrrVbAXhvud1qYv7MSYOZ+o89jPK2A/JoOYFSGUs4Tz8+nl8ASBF2xIY+A
yGBIuP/QbK5nC3gxJAkYJVaBxv/H41qeCgaUQKFtsB3WuLWxxK7MUiY/9Xiz
O1XvcFHTdktrXUumVIH/Nx7pyiBMXLhIFw955KtD7gkElx4tZntXdIGvVERf
F4Xkm/bdWyP4hAIptmyAEv09/iyVE17E6maGPT35dEWLhxRwKbdk4I+IIept
9vHfn9wRNl1PJUuaKOwdubfCBQJ5v7JDs08e1M+CEtjVp6RzenapnfNZ91Q2
Nd/kEkVj0FyyGXU5Udc/7ZvtBkL1JzYycgM7ZmVSrRX1J6NXEpvdW0pEQNb7
rkgLgx36QK4L8tacQsxp17eYrEG+ICUQMH0/S5Xts1jpbBh9L9xG0j3HBgHK
xMjXGVVtB3Q9+AqhBAwMqH7aDorEKn2MmWec3rWiiPlC+qGUPbIq29BtkFQI
7B4nW+5XpiQ+tIg9J5K5MyLzp9GPyF5Mva1Cz6R/Sns2kMQ54ES37RMdKdEj
DpbEHNZULsulZUoVZVf71xIpSrU/+WZXcRVoOLGHfpMhWcG8gYpwa7BwcNdc
3QKm/iRllJCoE8VVjbiyNCxknS8ezO++pJG7XwH7jvluL3TMke9Q6T/IroF5
2GX/KpiBwu9rs6TJFJnD8XN3Kf1FryObb8Yr1gSSSy6m13eZR8YhTnP6Y+Br
+F7XUSCYTglQwKVmJCcQ4DzQEakG1pZ7hY29BfkFzUwqzUF8s9qSBz3KJPqC
Yzc0seae6NkA7TChnMUJJpWzwCWegtpT4xxpguYtYCvRDnflhaXFIpowFrvO
nFHYxMC5dyUiID3WWdg2anDU5la3iQh+X+41j+PVvJ4Gett4MaSu8RIUSQdO
e4noPVSFnHiPrSoNaR4W2/5llJRHBvZZJSRkf3inG0S6zBCS0SDaDA9APgX1
45biOqsmCmHsvTkzbZv/LAXxELXrZZ9cGBiAk1DucaWDvNXYTJeGfpTX/fEC
eoZqLboUIdUwLWlhUUSU1KPyeo2Z23+daQ2/PvfFUmcrPjDbfIpgv+qhpLih
S8lOozBu+vNUeLgeGMSiXZWYrDO1QZ8nOZ2eqLle8s2UsXbZCJ4QPXhUbQYl
JrxprMK23Vrr0EfstLJ81iJnAoHiH2wA41bN+Pwb2MXAA4AxGlJQP9K4oOcZ
O4+VdD4p8/zO2+DsmJ+W6s3QDrZYOq4y6BhJ8CtxDJ2sD2xaVSQSJzWJxSpV
ww1lqDD/1GTOyFYNc5jVPfiW9q9xYXFaBIAQiTVH0v75M8R+6DtszkWyqBvl
jH4POvHhjG90LzhbSDwtGMNdWc1Noa9aOAR4a7WIFqvK0JsugIu+qDLfZ5bp
WdSWp4cmID4wB1py5v/cwYw4811jVhuCk5zuCFNYQTOm2qTF19xPXBHhA0WM
9t9GXtzzVO+bM9k12JrNInm/znFVfs2DaKmkVAm8X4ydgEW/+b1UFU0yzmpb
S/NPfvLlmHw43xlDXqkldCcW2CSVTJF+CYlLeVo6Zrjcs9xOfO/+A98MPHAw
hOcAFVplBwC6OOFg/yBHZlK43+16mCS1Lq8EBhiGPFH5s2HGJ2TIFfl76Ov6
JqORpjQebfi8lXNBy5pr0y4o/NaTgYdUbyCUJEkRRR3120yr+ExYBk1mSKT+
sMKXV9e8pWSj5P5jNiDNGBJURpaPww8MRxWXOhFU7611y3rWeCzIrEFC1Mwa
ZHI4xxHTctv1u3A7OS/Q97ru4Viw2jw0PPQvFqzwnrsVeVrGlCdZqYZRdj1o
DfHMh52UsrE/2eGMI6QEwp9sDdM5T/h15AHkdBgRAF2OenfRfa/elUvLWZ5F
+a9CEWMDwFmDcAOBGZr1+fsDlWzZoEVI2voMUfxIUlOMZS2nd4e/6saCPDCB
914/lD72OMp/9RcnN1kIC7jsU4OVovCdN07/uEyoYF5E6E0aAaw5hFiHqK3p
3nAx+UUn0s99olFrm7f65zs/dTRAI6W62twiWFboMnnP5AC1jEkO7yMAp+wt
sR+JH7QiW4MTW9ROr9bnRVLm82gYY74T8DjU62jE1FdJgvzK0dDCrLlI04/y
fpCSvflThpSDiiXn35yhmbj82VGj5bivIFBT5SbS6LVFH0nBoe6x/T5Jszpg
ZadhOM+BmjtZ8vEs16F5L1a299mnxnVLorUOyQB0gfmICo5wYVE08XjeUoU+
faeNON9a5thuImmG/JkOT+WQHJwmoZGyyBKgUHVh/AbhQgtZQIPiWEgwi5vj
qgyk4YRQ36+eIrfxSPnNyBgKQYz0+wdZDWFxSfscIJzO5W9zMpLktI82aUCn
KYNhZpfdb6Cmy3UdTzCXyFpgkUUkQULO0jYwtfc5xqswbfQNazkWEflZjdf9
zURr8fG5Z29bf9QzX90jLCZfvlGkFTGbRleBaC6VtUGxfydrIZKkE8Twm6Ml
MDQ/C20Pg3Ja1RfgkgrF0V4n2uWiIxkrzsGAmvmneGD1uwo/H6cnNG+rfGNK
woQYGg2iclUofM0kThtrYr0Kf/PisJy24FoppBoFo17SKx/pcMAQ5zpNerNi
G5TEspfM/TpQoitj4Ku0tJIWa6ue/Sh0dOC6SmvLtYPSTZc+BI1+Hjm2VPAA
yHGVIkLvbic/HwQgygsAA8mUQjMD5tkucbizaVr6QXo3bPcxbkuiMrT0N8yo
3V1GghKzCdVNgP9vzbzH9PpleSBSKC2mLxPLud2t/npwZoZ6KdlUqILRzBsT
0h24/1P6XuscJgkLsyPDfs1xjo7sd3Vim9y61beUZXlPeGnT+gNJkprm6eQT
h6eZ3IFG0bBqkHL1tYM6xp2pgnJuxH7pe/KUK2wkseHaLFy7thYgycRzk1B6
mAAcPvN9ykon8mTkQamEDaPvuXokJ6UW0iDv6/vmZ2xMNKKuGqn/R6m86T+i
7feGnC1LRPGD+kQXCeg0GuxwvUp1Y2LoH/w53R7NzH8SWisfszg6gm3cnMkd
ZeDJXy6sr/mKYcBWWoQ5Tuz6iL/vcftEkRJNbboY+1/gkkZfzKgmsTnpyAZY
dZhoPFsZGoz6GSeEVLO1zxykwMG4r6u7gfpS5j07kf5+pm9eo4LXbuwO4O2F
k8/sF6ELx2ripqk6cvkctkCY+WTURfjZAboj62uJAzXLt1B4JtG1vPJYWi6Q
dAae+zEP+nqPR2YDXSm/YIv5AmlcA6h7Ip55wBSTDejYKM2tBsl+qbi66VCU
oUKmm1wBbu0aoT+5tgWqLKsYPDnZDcmg+hlquHYiM/8EC0v6EOdEk91ykDQQ
c5Y5pNslSsS/mdH/9n2BSux5EEIiG1JxqYc9bLj1WaDDudjx6W60tid3pT0+
ie1X94pjLPC9W32EStpzg3J+4RStDqhuAXmhNxvEv077gM24N2trH5LBFp46
pfZFOoNVu4X4rIygvaSMTppIpyxJ5Huov3aiLrhUmzMepxyuqO6U6o6tUCt5
1bqSgbIWGilMHY25LxngLNgcSlkXLw+9umJ1Aaqr85+Gc1/L5t/Dl+EFhkmc
FJ4+7AIoUlcNuCdASKx946BMtgLPQz1RAG1tjQSXZLjhdVK4adamHqw5diTn
Om4UOAfme5oUohXb6nwFNxDPKyM5lQaDI4JkAWP6DVFWWyFUmriaz4ZP+ZGW
dWNpP/mVromR35ZU2D3ZPrdy7gN+/t/llZPhokPZ/hP48UsI7Rvk36uUgYW7
m722M7Sv/DruXrxSvsw1yOnchRxEogtK9VGsAFOlozGXr5XaVtqVKxT0VsPk
3wVD8m9VaA9c2M0VuvzqkqEX32M6p/GPIk6gIObpIM3k2ykA/AWbGvUB+9+g
fdcKMAOj1qkRLNPketxFYptpCx6BDU0EQ2y1284cT6bhNltY0m+BM/LoN+yu
qusHUCSk9jEFe5Nrbtz6TKOZ2lQMEit0TXGo+rnmJtGPiDko/wVLeOb7GvcZ
KlMHUa1XBFBUj+4hkSE6QH2dOaoDn4nNvSmUypS/wPYNLpUh4mtYwPL/BIpc
s6UQiRkD5dqSR5S/gu4xenkTMQ4A8UbqkKQn8ixotLHZxS7SOTJiO0YzCtLB
LhuF7V0qLGhNGSuNZofLLHMn3f1l5pmRCehQEpsocTcfOO+0qn+sN/JL5Hmq
lgpXieceAxu/DeFFKE/qai332bmDQtkVM+N+Wpp87bGOVwxonV/KiIBx/UkV
bMiZXti0s3NtmE6EsPzhLNQgL4cKQFzYFFYz3/Zq29gqb0CDe1cPGH31mQaQ
yfLHmjhbRHltCcdtBKn5eE7KoKjJSXCb+xUZOXqp3VpcfwpFSq5DENU9Ho9y
RygpPoTKBp+qnaqcf+/Hna0+5RF06PDbfgZKQtWwyxiNhFYzDvh+unEgl+Pa
ivye84RxAG5IOZLHNrwVX6oSUap5H3c6rznNUYB0pOFEH0GM6bVopAqu2g3S
qIdZKKeh3XSjTTwvv3veD9Kxnere8FmET9wBPswziaAGWvU5uj0lRPv9UAO9
8vVteWqTl4nyHSZl46OKYpAkEAll50TQ0wmP86Fo0l77/QgMiUJbkar1x95k
CVXYh+pAWMoAP47mbuhxwwwSxjE+as2zPqwxRGImYv1BFtZSTK18tHTyacCG
gDdzdLlhX3F9bZBMk6t+MpDJlGbDkSyiZG9PFUvAeUWuKJOWXSADSCU240As
skPJARvjtwV9V9waqQxqeBaZfhj0jCv43Fj4bWfN/TcCZz9XSYv4aBlTKH0M
7YTGAsHQXfD4MUWes5R+EU4cdZGbo0IoKyMHwHqGFvLT32rxIHwGgmb8ixMJ
lU+s/6ZDQh6s6CZTRof+h4v/UjPqIkNEtfeqxdUOcrr0AtrxaGgazxDrQyth
5vuiGFIDFMkphNEkmkJU0RL2ikUGfdP0q6C4wYerfOMcuX4mYU1DyNtqVkw6
s/0nzxf6B1QuIqDc2zxkyE/UzrOMpvsnMEhmIXUc2If3buC+kOiJytx1ynuY
uBTEzQmxF8qOMpZJa6oRGaYdNO69D1AH0gVYW2UH3Wz9ziARnuCPQY9/6skh
AmeXXgbtQiQelR7Ee9Z7J9C5faTL9pbIUi5tXgjjTO2/Vo7Fx2Gun7ZHzPwr
uTkTXpA+uxhl+4NxPszecG13ynHox3qWfXy8LfAHAtZRde66sfJGBl0UzWwk
WA933VOthjkx6asQ0f2qqjuQcxnQkEfkbw/lJ1suv5wJX4zvUYzoOR6HaLX/
L/eNaSfYaEo92ReSQfjOBjIPe1AzJGVhUAghm6Dgiaqe31VU3ikI7AKMB/Nf
KHKmxiA98qBWBg1hkTLizMDOrafOc6kLlbgRGQz1+tIrmEzibaNY31eWar9Z
Z+AoOk7hUzkSiWxUZWCQkl9JHldWjsOzHEswAn+bAFoteSl6TslZrPuHDpF0
nQqje2kyrw/xYTToXHoAabrmvKJJCUtgvEXTESZf2ZUUqZYVjrBBw5btRBa0
b4KFnuFa/lrbgoEVJcZe7xKUqInFTrTMXMgbN+aSzB41LkP233tN0avNoSrK
MnrWEgRsAxWlENJ/B38QPA/TsOC+UDJ8kjVMF34vl5bQVOw1JsPTBQkrlK5D
B9sEfWy0ELkgxASSYYKmUQAvWO/6qjuKC67b6sKeqRnGA6ke+xoLKTn2xJxA
Kh9Nu5SPCrGcu6iIYhVlvlcRLUOa0aRLDDxZVYx2gaFNuTbjB2CRuwYaOP6x
J8e1jYVLU4EWSFQvP8NMQ2d9I8dC9uqUAjgdWavauqpiMOIcj17b3cgKh7/E
n45BtVo5nUEItCTaLSR3ARNNj/CE84r1k54wcECzyiYhuDX9YKyEahgDKzZu
oLz/HQzSBi3R7N4MfpHUdcik7kQPs8l/97qM5PUGPLOY9rEt8OQOQQoRFJra
ufS4rHx/pSCnBLmMUiaXn3HRzQdvlGO7wIbiloGm1bWK6BTbfO37R/bXbfwk
Xa8OGSlKMd7v7TqQe7oIFQCqBdxu9UvLY2s8sk70BZ4clMXudJmhs68TmJCO
xi+h+8RnVeLGJYHZX7JSKbCddpFrQUD4TfSJpc2O9KrdbDc0LxX4pf30Ry0s
a1oL8hCGLoF+Yns1q3jIba65g3k3yGExPxPg90hd41M9XdaXZ4XPRqvdMRBc
t4Qi8VnDiahl4r8CkINW6qKpq28bAGrQiTNRJfzDqHFrUEY5b4of/Biaz9pc
NhpX2YMUN7dTBqSaEiII0ffwpdSg/czvMRu2an6smMlHxfpxWFWuc1Dia1Jz
lzdqMSt2GRHd4QzRvBSayFUsRPs/wY3tw5sm7N+yxATAyNMRLorYJ8e8H/y6
H0v9N9imisNDyIY6GENydLcgDJzV2XDi8Wv1mb6KKvooJQ02MLV+GlXueMGF
9lYiAefrOgREcQKK1CjR2A/wPqIkZSqrmX/TBrunfnYthqj5uXryDUSYXYcS
Wk6MCam4YgVFmkQ0IA0y6bQl1wbi5bM/E6aKVSi5jmC719HQUdsFvQh6w9D3
oQq/eLBmkl49JzCoaKM52lJNJd7fhksR9bGtJhbVoiubwwg/Pv2aTxx84ut7
d5zcsVB6Xq77Dnv2HUcEL1wdP0t3kHjyUMdw7r+r1W+HHTV9OMhipwuLZN6j
EQ5AMMLgbFGZ0HwUkJXx6XfeHtZvCrfidSqkgh3lsqEXh0rheGXFXTDMwPRe
bjyoEXrbKX5A//j4pg6B5RZUBzb3GM5Jc3cUYoG1pbUTsecDEYkfN0VzZi+j
R4sefMaA9pmCJCc+pHhKi2+CeKZfuAIOzr4DrZ1f0mwH5fD3qHHxpxos4iqf
Q+dq3DMl5gg/gbl6UprtIvUqo3Ce+xl7tInDKk13+gA+rfRL70i3gqedfuNT
tSi82QWK3WIxdP2n70ammTgrk+237IbyYk1sAYBXT+SMvIhy8Ib/dms6UG2u
3viDf162a1IoSPCusUcfcZMG73LsiMZWbBovUppkvYpj8UNow6dDp7jA1x7o
CpWPfHXpl+IGbnshJyI+oUm0g6ZETFoNH0IXVZIx3iykh8o1MwxbbyhttvMV
tFxye9l5NOVfiPs1rmkCxpBkWHxzKTVYo/4or4pGQmF8/ztK8KsFEvEHBKJw
H7xSufg2IeHVt8GKieh/0+0iTpv8W7KXI3YuRSxwke3t0Njq+SydXtqaLyxp
H6ZBntjYakrGIpO8FbpXXmH5DHJXcw1pTI1aAi+l3iSnpSzfatBoLImHTLts
oOYqQCgFZsw5zoiXHpheCmslAgMcSpD+RYRVV4HHmCESe03uCULd0g3nndTu
Z/8+Q2UPN8H6CVDKwOXSRQYWh1j9u9uKtOnMQmiAoFILioJrvK8G/II0+XIr
sYUkavT5thAwqweDtF4j8BzVdA+dupDLQHjhl9DgNcXYSOixjkEdmZ5P5fUQ
OZmqQ9z4Rp9X9HxslhjetMpGBQtAYMHw6pDSYhfP/anz+Qqz0wG52r1x5Rck
E3cB/S4Gryv68Cji0FIoQ1Gc+kL9/EC15vHEZOXFlsv/ApHE8HVZwWmanLWn
cNJN7iq0UwO2yI80n6bqWZpQG9wjVsdQd/96zkoZY80NKwv1SxMiAk3PpDzN
pPZSZ3lp6oItuoq+AWtzHWSWVKcaK98UtrWdJUc6klG1wmqVmOjTC0iKnjAU
uCH/ERcDdV/Bx9o+zOn5JZlAJ0kdmtphi3A8hnnewc7ebmkL6BpI1GmVqHTS
WOTz8qYYhFJ0Kjlbm/Wdh5cqHTnXaEoJ7TKFAanVlGZQ6XpHt/iWWSY+N/uz
FiTsRYf7z2cPOEijoFd/6v5AqVVzjouVk9BgEHm7oXV6JGY7L5bvV5f+waER
qQ6O2S/MaHHWyxYTs5RrjBGLpmyGbC+3ls+07M4G8XCgU7/5Qb7d/yXCCGIH
4Ht7Mb6Ol2gLbKWVINOMsV1CUW1YD/fbyDm0HnFCCOi6sBodo+VaMYyM8Y8O
81Pc6UqcxvtGPh+II9sPHWMloNpSCYrGNGJscf765EFXbJdLyPQ1s0cmOSZO
BN1QrbAc5SqjYWnxeB4Lyhdkn8r7WwUq5pDUXxrpccGptZ/bvrvzIKbNEaRs
vCbxsvq2hGmfi1KSWYjA0fjZ0WScQUF3Hp4drOveCG8MzLIqjbtAIT7oQ5RC
vUfmC9uub7ojRyATBZ9Q+L5MTxNy/QqYss/noOl0fS/0nOC5nBDgx2LtxWqU
gbnwHBJ1FPNJB5AjFulbxRojN/RRBOFqcmnJw4VTw1on7nD2E4OdwiqrwxzR
zNrfXvEMPCKnD9YBnBoaDAgx95gLKgEZuuwkdvt9yjDrbnjZ5dQO8Xmjb3/n
ZiOTuNnwDIqNVT/nl1TYsqW+uFVvvZ/ZVJnPkFFSFqXXI3oYQJBDZIHhXWKx
oZ7nNU+vz/ZQT++5/PUB3n4/n4SzHc7aeKJti+G2es0ShRlA6X0wEDOES+UP
ChpmMtRBWKTOVGIQnv1LSaucVmQdLUk2KM5881j8Kufel/ME/Gzfa1iXjsjX
u88tME7hFfS3Qkskw7vKEX40PvFWizjzNWHjg6Pw/LBbv/GuOY09mWKii7PQ
RB5i1fPJurVeuDjX5dFOK8xFo0p3MhIMTikOKCm9LKKjXnOne1H+VZNIEfgD
CpkVWscr+LyNPSB8b8VaiHnutbshf7AVdyHMwc9Jpkx27K/IvlVUjgdPhlkP
8QTq+7eCc0K9Ihw7yu/2FIhcnk8p5aWWtZjhtf8Lb2DVJ6/kKPQOM3fROdTw
m94lb/+oMmjX8mwahGIivSt5tTuK6nTgli6UWwFlzJOTHyZq6KG3f1v914Dt
z8L5uWvdrAnH0ZFGybEmhdtnBZwLi8jFvhmR07xTEOmvPmHShf8TOJheAtWb
UfJ82v4V+9Z61AkqZbo9D4pL0dJTsuWSliuGNeqZcIymX/5HtL6tR/w1vygl
eiVgcmNX+VoQ0mDS2ze4iwON9WkBWy701OHzrvfeww2/xgCMC94WjgYQwoCY
uT7i0tcKOujnHo0JJE/bASyuIStTnqKreO/JOGtXw07sPwlJlPNz2yeq/oXo
HTrsJAwie+UTdkERwrN3qkHwJO7cS+USeT1G463uTMxICwh6zlsd9lSArZe2
mM/HQtbEDzBSqM3abvdjofnbGyGsH8EtuxenKbmJKorOjhW1jkgaojuUUq/i
TeCsourAgEeeO2z6omigu8UrlacnMwDAo3Ws1qq9XSKe5MwXQG/Zzy6CNwR1
o6gRd3Q6aFSXwDkt+ffnvGMhN4+ZzvdHMpZdweDQBNhSFvf8fBEbeCW5tiZ8
oDvqDpozIdESpdt8zw0LTRemOrhnM8adceg29GXXgyaEuxymWaZ/Q+kPqp2C
9CtGFcTs9aQYOjMh10IJq5NwY45WhGTzuf8pwlV3a9Z8lzdqdG0N01UAmXUV
nQ/ItPlSKxpDbWcgOMPdjlXuzVL0EJDfjHK+DZlwHsqR0dh0qqZOoWL5+Kf+
T5Dwi/8jkHb1ei3FQOXY9yFhZkren/YnJTx3enTqZjyLcsjXxfHtK784c7yo
jngEq5rozt+h/OfZjwnej/ORHHGWs/x5ICy5ukdrm3Lr6Av//7yLAHfJYDnE
nyB2/TvKGd6EX6ftIKr4siaVlXY5hmFaEjF2ldYlJwn+ZZao3RsV5588hmGA
KhlEXOvRUAAR5BmCYgQ/9OvEqC6x+G/6B75uB7gv2dGvCdbvdrgbp5yaDrid
kBqSRgV+oAuusj6k81/X6CRYLWe6lX8P2ms6k7t4a6kNMpV8qLgeh+9z2sC/
oWE+HvEfzx+fDjKQTBTew1ql2LdMx0eykR9t2y+PNg7Zezc+ZvDvDOnxxmAr
TR+iYQ8yNQdYaA4jRdj2ik2gT3z1lHy1W34ihdUv0TcP/ACDo8PA3CQLsMXW
lgvSf1Y+eua+bBLK3Sj8liX61EXIiLyYJvcQvjNbff8+OmVmFhlDEPPJWywS
oFh7mIISl8iT8gEpvUB0EKHCVShwef+WyFDxuZCkPuK+Lc3Wng4Y7sjrPTLB
du1VfqqsGMCnOyQhoLDJ6EUBC1EWE7QGO9QE7gZePjbUGlBNoXiVaVbgN27v
ZMnEhtldVlACDX8Fo4iimcw9lmaORu0ZawpTb7uAd7qkVwwVrtyYI8eRh8SF
xPA/Sqr9ZkPAI72iD4CBtssagEHBH4LBIbnQEwPbPFZQkvnC0Lx0bpl/2gGr
OW11wtjJMpQ+Yv3flpakhgHEbM4VvwWhlBX+opJ5hZ1jUH5Im7nPCBAD4/zr
+MR9UaPNM+oqHiGBWJQT3e8hW7gBCRDMWVGDJcRB44Dz2/NHv1IEO9Rpzf7j
6itQeQ3mAVEAzUcyHkIPXKt22eiJ0BJQ/SPHfJQ4Yp5lSyJPM/Fw3dN63BiS
5OBkRJR+/JoGIpsJOKaJg09/ew7P5kaR0aO1x2ml9pnm/FK3nVByPb4L/RIe
GH0uTD5z7GaO3AqWOWyptGRTfNt/DnTKC7P44FGsxdfqc44iheq9O+L48tQX
uPqv19kRzLgyHbi3l+/bqTC9fU9oMXiRsJKnHDaBOkpjWXE2fJnDbNf/Cb30
sowwcdUYl+ENcZJ447PJ77Z00Ng3hLW93CI3Rd9LKo/vuxlqBg2gNCp1W87U
6iee/KSd5iyLDsimpyfnNAEvmA6lF1H8gVc64bmx1LpwyXGTcdqpXTzGzo4K
cIsSZ3MIlEESEfyYhPGi4ONMbSR+IyUH9S9hBtZWlksTjOgn2qDnevgFIQA8
GhSxyVZQVCJ8hLFDg6JYEpYQhNNtdImJULDOX91Mju48h+/QYryRQtW0qjsT
nDtMSMgNXqkGvl9BZkkGu5PaKrK//Syu2dvJRL3zxc10VepmIyOya7AeELXa
bG15CxYY4nDoeRVJDJn99hyqnkUzXNgaMvL7yj1qECMXnFl4tYtjIMYvSD2M
byjnzGjwdj8HJPKzRpGQ/dONZalKBkQVYyzMqee5DhASnSV851sVZVf/F4Nq
47TDjPzZgtc5oIuheJZJMD3NLLd7xxkJ3th5yTr4iceyirVdzXfM1tm/Ua2f
vFqeYnTiNdKivqDwzKV5RStI7U/biUUl8EyB/hr+gGuqF5NIdf0xO+qIHx0R
jYwL4MiUE+elkYUx+f3whL+nKGPEsZoYciWX38G+Qp8xiiBDcVOP/burxuCg
gkzF9A9YT6lRh0gt3RZPAUk/NJ2UQ4tlPjhJbgytfaFV/lR/kLZ0kOc1O7XM
3Bb/m6VoP9Z3hPPuoLSc1ls8w7h2LwjUCRQH9HUb9MMLcFtBK4FFmSbAjPY8
D4PA70gDhVRzEohJdYY4MOOqtAshP5A9EjtMBIxCHJnwYxN6qcy2NNTs/uos
JUEdTPZx3URCxPFZAL1L0lLz8i+PFKknrdQJN/Lgb73AZ9DZ8xPzrhNYIw9R
Yy3ouVDUyvAUGGCG5ORj1wJw/kuzH8bp2ggT7sM8HdpzitxwgGPmnkKqdswU
XCb6w4MCVy7qssy/RDg119pRRvzGNM5hYwP3C21EwLbvkOJxixNcDrCnbLDA
wznL/6FT7ZSgCgOhWLi6urDZEwGLFPSwqnygi0+Fy7rqY9ev3a74w0FnB7A0
xyLG/9m/qteRui5HUYr5oMM1wQz5tQhb2MStb8S2mai1UdbfmhNiHxRo+SWv
EA9EO2LkylY8HHZst0LYQCzoHHE9hWnoqM+3o8Bvn9hFQY8HWQcO1gFPar2X
EI37J8s0O3rbO8C606kXUFXC2ZJvGrycnpff6x0WtGoeEZYCKLBDdlT9r6KP
BXxn4BRSyCmUrHYnnD68m/7jLpYCUNkyIggMc6qRaB4ME4O0SAPzuNe+3x3n
QfRNKX5t5F3UiUy8b1Rfsd4E5XYzdxDATr3FIssh5wn48PDuvnVSaqoUJXC3
kiII5Vd7P8N7PVOqWKi43DGWA9len7eLFpo80EkpHNJR9DfhzHabTUxsAW2j
eoRceuArRg4oocrfJsmAKl395CJfuRaBScvMJr2eoKTMK4HklwBKoTiD71KI
opd4iY4Yb5Pk5fqF8qSCWXEXdG5GXnAb03HtR/li9EyE3c7NdgJsXrNlVSuI
4pyDfOMUHK/1SM4zTuztgxTIxvK5HORwLUg+jYRhAvTsg6TTqsgBqSm14vqf
yrXyenR/AmNTci0aADU3R9rhDWjAQtUy062oJidhsP3/gpZ2LkVQ0cGsqEWY
oLv7TvW48ULzV0risJcHTIhHnTfHc9/MxKq0a9tG5s2lLPqBUhKHkC/Eaz2U
xTNfXcJluXUs+PwuTF2w6PzFyUsevXODovWf5yHB4HZpgtbbzdyzmzMGy8XB
1zhWR/Ria/m9TKWbEWHT1ZPLrZMG6/MbmBYoQPdxJlFW0qrORHbm8aHU+Cy2
b1fhtxu3qD8EOH7FtUsYZvsVB7bpH83OvSPzlEKjhifj/oHBPfYD4rWfJq+B
wpCI/PfZ9M1BtWMvv8hHSU5RkaJC33l625cUeqGY2/lrji/VFuk3q+1cT9zR
P3O/JsqDQp2WKOxSw4tsBNEHAD9Dg+qcNifk1WAkrYqT/YtgPYfXHlqj5MtF
BxYLglpY+mZa3rSvHURy14dDMVcn7Wst0cHwaNomvAAWNYKBJMGHgd8CX+HH
t8BohPbTYKtgzAXyKSvWIvFyNtgguVSPovdXfp63JxRBF+t9D7lFMKSIejqW
L4WohhYtD7UK/H2Odt1x7Y3I4JoH71mjxe3Df6aofJKi7KB7QhoTrLHVJ2ky
fnHaFhRaPJjCTAYxm9fJvl2O3krcVwYNnLwwEEKkKwArCYJI17Ue8enaTb3c
EXJeb9ufyjx5+Fh6G7awbE7yAab5kA/vlm+Tak/xEfFoHoZ/Mm8YdKrHEBYR
Q+ucj3t0qIXHXf8GXs8TmuMXqlVQgQC5LrZxXBmvGC7K+uGkN3XkCzblB019
/ynPy2AASjXolFMQEaO78LS3R9bVbS2yiVGxH/7j4YzfYK44XeYC7A5AyYGq
hdbt4QYx+nhI5gsxD4n62X/gRbQgWdT3a1cxTjAvJJ88h5JijqqbClqiG3sr
TL+ka79q0q2YL642m6VLsVfDhgfY2J5eH899KUn2M6F7bLhqtIa/y3jkyHZ4
s+ZHSETQzx7a7a0xmEFEYVgYIz6nnxSQN5+uKYrzgRjXBb4jlw/xP3KvhIdu
HO0d2nVHEupPyBEw7RLCUFbI33gYKqUYvAXpaBepoIdBNU3j0NXXnDSwFSCC
7dOqPvc1IsXa06oMMMfpTS5Iy5GMdDY/Dl8/DpBsdVOYNWiVXUTWLU+dIG5g
kpNnuG3TdQ0zfrcWprU/jm/E/qT6Tbdc5R/ve/d7Aqrp88HIEjqhj9EKTrQa
9rB0mIVhCdK5QblUQ/hayi9PNwkkBz1HIjXAk5nv1+NGM44xPE0HMfvz0H1B
cg9xqwz2XbM+OUEHqJfFtSEuD9OM5K/AMR979dBS8mJBGSTwMCshvt3/wU0o
6bqeH2fN9CwYOpB5rQ6HYYglQ+Rh+LkyKg7ONbdR62tg9Lb5JkH2T15kFWqV
nu1/WqOmgNR02oj6OAZMySIv+3lLzxeoGkQP++C/wu2+w6bs5NO/ByD+9T8t
9Vt7xJLMv/GCbnLWHMeclZRuYDJ7Hql9gVuCL4UOxmnf6u+BWiUJsFHY7MwV
vl1oMp1/LUdFSLXuhVud282I8nxKgyFr95z2D+M3s3FfxBd5T9HH+dODH8mq
HPacBjH0wsdHQe4/lNUYu37nRXmHF4mKPqxhLcgf7RY6p/Tpv6iP+UIQ3Inq
KnI85YLLj4BD52a9UJDBLGu8MY+2Tr/yb3Q7szfarX5uMUJKKLTYdJEx+Qgn
vtyovZBtpDTpou2qg7y37BoJR7yKFRdOHO1LJNhQHkD8hdQKSJkvTTuSMi0y
fWjZJk1gDOe6Ygwo4Jc4Abuy0NuKimhfOi3qMdf0k9mDd4NyxqWAowRmLked
mKNEKMeqMil7b9orvbOH6gSVOu/lQkOc+z5403iQSf7wJSrx04d/iPcOMyMa
r1yvm9C8qEou0FKxaupVhTfXTJFh4bCdaUv7+qQh5h5TRs/GuE60sFmx38K7
4K7arhrqLjOMvyyXw646Aoiv/P4qLpHWit1R3pi2UHXzeD3rpecSXhj9lII4
yKaUzIuPdStsom5w46eAkOjTfWFyNUhtKHUfCmNhvp9j4hpJAkUFWv/eBuDN
jvsrGrIa1ka2Z+6yiy45vH4GgcyEKWi0ifLO+G2rne/4j+E53/F9oliR6VaT
CpoKMgvUe4LfaSix7EWEiX3e6orsnB+6MFX7/KL12KC7GT+TpsLqM4ayK+68
vHjYuqx8L5Q0cSVnkE/T7UgWqx/P2LFKhMUwC9Olj6FCz5vQdABKEpH8HcJv
K2yejitkRzCzmmNtMPoCkU88T7CpTcK2uHedMzmci8FGC22DIiGsJxKyxV0S
DkwVw1a8C2Zap2pmb/uXQOI8of5QljqPClkcZ/30aU3Ihi+Fh7Z0PK5FfAlj
sqSTEFX3pZ3neKMP0+H13MdPVbVcavWfQYzj4our/1OAfsRVp5QCGrYRZy5K
+lBun+KXPOQqK8xIc/HAN8WMdT1CdOuIMV77Yz/lq/epooMVUw6GOexRvuQ7
n8yYO1eKii0WnA4s/tWUhJwJp0sZ+YevhcxUj6H5soko50yosu9PpLJrgowI
KYmWzbiqtEbtVM9SrPsfbUuMgZm8gDYjoQznENQWdE/Typn6VnuqAAkonGN1
BlSwnCJjEL36HOJSgKXM4om+kGNLAioAhQ+2Dqpi1OnOMeRRYz5mykzzeab1
H1fYitMDBn60M8iAKPFP+y/QViXRJ3mX/nUSZ7rzu4KsAjRXv/k2GcfAgv9Q
buy6iwwU4HHXkuFnbGNvyhhzNZLhiHC8IRF9UYHBrhu+VlNn6wXFT/cWboEM
EtOasCPxmCOq6/A1REJ2KwZ69AKxyuUisN7SeJfODQ9quzOb2IZSubKhH0hF
C+WcJztKUW+W/5ATGQcuXrcN28zHR8yPosCpY/ESyVad8eRQMFZ+aSwZ/b0w
wQYRpfESPC2gkd95TCG1uMfzxNCYgVq7kh6PULmKKuQkMD0XVXbe+Lvi6t5x
g80AI5HIK0RoiMuk8P7c4n3aBuyZ696obdvtb/eFN4+3zpLP2SpodiOENQr4
mQ4iT4l+a3HBZ4e31Af0d7gh7zdwFxYtPx7L1zetqzcRyamYAZs8DXZUDi56
+2EkxiONBotpACx0tebvwqd7ru3pepniB0fdvhe+iiBf9yQx9oKA+wlGaQHy
Wi1wHucLnuoDHTFfHxZkh3ZReb/HICY6nNVtSQ5ieerFzKuyCsEOFtPMkpiT
qHslvvFNJOgvumZu1cFz/BgOAUWfbUL2K7cKZ/wc+79nDVzpl2jlOG5WyVTU
CoIInCOT7ljU4cWxwEkx+KytUoSZIztaJNk3viSKZr21PM2DxLE3ENcFe6ya
us0NvL222JEv3jd5QqrWcqirzi48LAuP3M5NYWN/gSfVNSTu1GXuHN6TukYY
j4uYkeyMWmnWActFJbTAAbfRh0vthVM/OPmmT8tQm+C0wqXGVgx0nu06ogjQ
45naQ9kVvGaKqPx9tiVD4XKlBb75sR+Ih8/Gc5eI5KKGEeLFGLvdjkNphZNh
q34P6FMsAlZVL0Q6AwPDsApGWKpBFI43eEk7afqxDdULFqk0UGpr/BIlTkU/
7qu0kkar/vozV36+SAUGMI1WVr/0BHILf5thEU8Hvib0/I9NPcTQoxF99BEx
51gvCNFRz8uIOeQ14OSsvy7KKzX/pKBq9hRhTQDJpfrX8dsK8KYSHYgZYd/2
iAoXmP4Ccje9UFqLKt2NpJ+MTUk4vWNyHnu1kWa2Ku3Gxbe2Zn33mlPBknwU
o36VeCk44b5kqyL+nbVt/0HjIplkNRBd5V3aBSMmTNLCgNqiHf64KP7yiDf5
zwhjXAxuReh8xmcXljdf/FAzyI5e1onCgvEcIHcrhG0/BAIMEKQbNhwf3NYl
XdNU3yqSfxBsC+/74qV/utEjBix4ldxLqSaAIMHpkVhtR2ldbHuKpwYRv9u/
Iy0V0htAJwMkZqjMHm/6OOEDY6qINBcGli1FujIE1oakrKtXM2T1U7woMNZa
YSsqjJAm27ZWkUu4B+CFmEPttw+EY8fUgzBUTCLFnfnPtFG6oClnbC9Hg8Ie
IZPltp3vtobeT7TaWVcJCO7HzImY7/aLmNEyqScKUjxwhu0bxAeb27YIiePK
O09qFjGtJIqgA5NdF/cGAnV2dZTtZ2nrifx4lnMEDM+eV/KqNV5bv0V9L4vc
r3bLToVKvKTpd1W3a9WzQd5DH1lWL+sqJnrX7ySqDCmZf3nLQOXRP98VFN/m
bJiSSkxY5sf7r7JRCgmfR6dOcI8jc6ZSoswm3vvk6UudlN577tvU0hGqmfF3
bZ0aoOT0bmZKIGLEVPWgVWo9Uto494Tl0J5GaTLVjxycPGBRzRmMiZroGdDG
8jYvpb+7V7eHYkqBaMIgejZTpBNaCHrvdpopoYeu1d8CaUxhWv9DW13AVRjb
Us8gMfPbosFwPzPGVFADB6D6Xj9MLTYuS0d2ECOl9Y4KZmutPGl9AwIqoSns
+7uROF1EPXFZ8ia6Tjo7Jto5depp4yqD7q+fg5DkkDmKbT94rCYih3F81IbO
INzrcoZe735ZTqkIhQDfdMv+2UDuhnKxlXapOhxeD90hIOul7pCg59ssjHG6
N5NT6Xq5q26nlB46uPaoDOkK/grNMrKK7lcYn46ULQFQ2ZtheKdrX6v5de07
ofhjsMSktS4HaeXT5wcVHxidAs1qAakf4q/UfNc24ohHFXLj4WFUpduNovDV
CMUr4G7g25t5iuIGWmuNwj0shiAN1gO5+Q+oXhdPrZqOqVG6hqrB2m2uQBtA
EnCh2WrciZuU7APJx5A2qgaqcD6Xbc5yxbVHztg6SDybmie1JdNchbP+OPd4
auG+zQ1O/rjhCjBMH0UhjoHbQWHQHLy5ChBzyTJF8/L5Le1zUw9Ost/dJJxM
lokhh+dfqZDjdfNmyXGk9z8Q/ZSAuwsSvvrp/yWCDsOYLeFr262bgRpva9NA
YXJUP7Fb1I8PSZaC5WJ95g/v2fFtVSCvg7QiA4oALiUA2LHZeEQR8i+9KXFH
fDDe1AAIvTuvH3AQBg604JOE7i1ikOpHuGEY7UU6GWHeCWbjn1JADpFRRtos
kXCoWo+PJPdPrEwfIqtIIo5TiD1RUPEwdc8H+oBp1x18cONTg+Ye6dubQ3Y3
PUQAI5eu13032n16ddUBy/g0a7Lk5c0PmSXOocQcHCiopWa7Wo+VfJl3sFUH
Q+u+c59pnaZyqZU3/KrZKOLh+qPsv0pstFRZxVKNJL4LflBa9FfTJ/RxnaP0
YyuT43jl6OGRaJN1pE0IzadsGj48RkOSD13sioIaqlSZrMOGYcacKpxOmxAh
oyDiurkeLjT3eASSPrssRjxqNvSW+8qTUpZoh3OCE6O42cSJFoJkAsz8gv/z
aWw92z2jYskdlEJtbVNTfOsXKU9yLEBXpz79V2SK7lkZGYCvJrGiNpi1oTzk
Gn5t2oMpMLIBkhy+y3Pd4QX4NWmcNgNfyVvASf0aIhYz1m15CUXZCc38iDVL
OF5LZOJ/jdphjFM8FMGuJ11qYxLeTuVSDl2VdEeaErG9KsdfJlsHPHF3EUK+
sopkSn22ah3dgzuTD2s61aS+MDQTOh+yOnUaSBLGFeHhKy9qaIpuLErpbCd/
hmz+HShdEJnI9LsL10WsZubrizgVbWuJn0G6QIvsWso1b0UYlcg0mjEgbnIo
f9B5trHnBGSKoFPAK+rhqJunnLhhliRvmopls6DhT7/oWgeEmIsnZiE8WIDp
tRTI5+nfc8KybHIU0zs0sYCDCXdRqC/gfSvb/p9xZyVoXuArY+Ot0y+uSum8
SSVTO2W0662VqESvhz7f+B+Tm9+U/DXy+uIxlJIP7TNKw1gnLKtj9CFR5Xs0
esBiB5vi0T82jURJzj8ggWF2bE12Q/cjEcxuqUPkyU4QPPzfMsiq1oS5bTkS
wd0oohdy0Xz6ZNM88hrhOA68e2wOy7RC7fPvpORXWN+ujlUAhQWjiumC1wt1
mEGeqyqiIJw0T1icjS0W+nh/7SoeaXAHEazSverQQsGh9DXlCwppuJ3Go3/f
77NR48SW5xiiN5vcgvx8wXoKM72wvd4g2uJtrOKjNq470PQjU9vKFAqw1OGT
D9jG+9hx6tZPF8gILRweerSv/TsXrJMi/UtTZtkziS8bSoBHt9oDH2pBPyoB
NrCjjb8z5XR1s5OZoX3KMrYPuB8xxNLVrqqWfCs/lAFa1oG2IfmNngtsGoep
tfft60zSKx/z7FWMLiOgXmCEeQBEheZ+KA82/rrncn2n5FisuaCRbG4QVR6V
lBNyFbRrYeGsCbCdYAr1z3XFhU5qWlh/S0TSq1KdjqPuZGfYBzzSe4/q/nG1
91qAwQ2CDqbpCXLLFGa+CINvQjeDjNS4/IrC1cHpTFdJq8A/870a/vMBfOal
+FTf6oVUotM9KRh7IUTPVO8cl9kv0P6GeYBcW0VNl5A532vstxTQ0Keg2Zb4
Zqn3dsXYyXpXTeM0XB/YJIiUDmT0oe1rMRQ4dAPvmHK44dwFOdX3tfH9ZmHT
Xj5hyJe6tW3YjcEJuIFaJ6cytTu29dqLxkDYqcQihEzLE/ysca8dEpmyIVVo
FdYqAW1LcU4E1OwuXxNFsrJIwJDaHl+n86YaL1nAbgcz7nBOV2jEcSDwwq5D
/mYwqhUiXDnh8IrrcD2b2z/vURp6Pvv2w9TXVdJRFoxfzbOI/PCcYuBU+PSx
HQ4d8nfhh1Cy5yryTtvlUjtremo4EGAX1X6Z2E2Ksplz8cZI7LputYIlYqTz
IBM059jZT8SPHt8oP6I/5+Y4CfQxugEEBFOBvMWkRRKxh3W9xzf7g8tsSy6/
ZAZ1mQoJPgGpTTMA5+vrxeNywRs5pR9GQKLgo3Xta9M018WOyRJCoPgIkufA
hnOQVAsotVlXe1FQrjl0cVm0KNJG7NUoA2DD9648/oZwBDBk7njHlATqRYva
ZKxlZD8T4o3K2BeRTY3pRYkOgfRQ2JDJsLYRJpzu5qaWhAAZT7ZbX8HalnIJ
gbZPJdBAC7E3PjDdqNvidbsA8+c3bbpql4yETUn1HKDKWabFOoYd+JkhbvLs
8njfUm6KbQdeMamNCeLQwM18VqUGzHrGbQkoUZkqSc2xjpavmXDipDChBWCo
5luB3gBFhaSXpdHhkmVrrZY9hg1TnrICL1v3HSsQ9VQ5Ymd2gmuVf99Ct9Lc
Fdsfgx68Hbrl8mZKhozLt20kXy4U1avNJ93/6iSktMCLby8q0ijJE9w1R6dC
ANZgnCdlLTZeuer1+0TCinj1so2UeJ7wJrmVF0OTSNT5j3zYfk+T/PFz7z3g
NlPjZkg3AevpJocDJCZY+FlpaOi+OvlC2aPMYqA4D6GE8zbaX4vCXP32q1H1
ZjLNQy3Cflxws62RxCDUfltbp4vnbVnyEBPaEKeApUANONtjFH7xNXbTLWnm
CMCkFbvV37gPFbLpMX9ffGAzaAPbcjStOEIl/dnKOMjS4Uw5R+OYGLIND7wq
AB4U5GXgVb5yGzDIWpY3zFfiEvyMb3HDOvKupEARsxhRapNcy5tx+I7VynIX
aWaOXKIUDA51n9LVORWdkwVUtx3KY6r0SWP/anX8QGPaeZdRebkub6B2uKsQ
pukoG0C9w+nT5vsm/+DVU17M+IcmYQHxbJMVvNCFrfxUur8YRLzetpgJdYwo
D4B3yJHObRu16AyP94iaTpKjED+tRrioGJ1NurD/36fmi75OVafOR5qd0Pjy
eFfNctOmT9voFGUgdi5yQ39tD7Ol8sFcKnisNqv67DHOYWbpbNcc4IdbzHYg
9HjSvH5I2MUsJm0joZV9D0NgLs7wwRgAO5bamGI6anLF32JfmOMj54eXBSMS
babto37uR2GCMtG/ljLIBTUMCc4sHx/E7c8qaRlxcaFtzZl1a7lV+htxPFMs
z1DJgiH7PFLydNYcvTtDWoWly8lH61DAyDz0iOaqMdlbIxvzdwYvr07RCHHw
t5lp0NQlLdcuHB1FOckwJ5RsoQrD4VraVAhwIZIjWV9iJDkqjbfrjzxC2QYo
RxdKd84k78LBY7NnUKSzZo0zsqzfkHObAi/k3ianQv8JAxqk5etgbU7TVRfQ
yq2HReYY4Hf4GeYbPGSaL8zDpQZHHvbE8Lh3nPYPg8tPoAuDJ+1/n0Uu9RaF
AR67+Sig9ey3AcglBUWEjt1WILyZ6AD11gsRm6xyydzneWnFKzzTJY/3SoJY
D29qSAq3fLBmoZ5nhk/wmmL9zCf+FAxyolnVpvJBGtSnJ9KnaGWzpDg9NWfY
D2i8cZDbZ9tKw4naDFA1s3hY/EGoDZ8UZLVdBWlj3+l+eWh4ESJrCb3S02n1
z97odo29jSdCQVpg1rPBtyMp7E6XVPeDSJXwqVbAv4IVO80doiD98rD+f0c7
iB9HJQA9m33WTRkknkDuutVOl74c2N4B0Ksdgmc5zQH2pWfJI5ayCUKoZu72
bL2HWuTVaZa+qCpzcOcVGTeNLcK8N5k31ytXDkUMygH3OP3dHqOzY7tuMSzU
fo7Y6VrCMPwX8I3ZQXvE10qP5nZAWwv8NASA7bE8A5CXaQO7o4Bmj1p5MfoS
Ptrh/bE8X6jhHk4ayWll8AOPVojlyjVIFL7LYYyXvKINVBHOYILKtZHLccQX
/OlnH88qR+hYvMh8mrZmJ9cj7gh5MQd/hSn3lm8ikEwWghSs7t4TWHwEtBry
gvACz27Gj70+TmhBmdH/i0Gw/jFMGf6YvKELyN9NpnW/bZeS36PZC3S/YTLf
FdmwNdNV9JEmZU+bgt2rQJlUds5xEu02Epjvzsb6cpJ/vyVhJkP7sfRsdIdg
JyxKK+dW6A5bDhpkb/412XrMMW9Ztr4FQe2bluwah0SGFLY08eMznh9aQkyu
8XD3Xbrm1fBYwMNHocvwtklmxRyBFgUE2GtzLFR1VVXzh+WHzIZbGzSlJ1XE
83Qu2quUzk6VBGcEDCHbkNnYG/WOxjSfEt+URwju3kLhDdM3QwSlU28nc6Z3
ZeOGJA1LOPgOzsImUdBmntTl6CgXgbV5HrKqEGC2kimlbm9ZUQKAyroAuWBx
VSpMBxmDr28pfCe74Zaw/orKYhE35zmzJxhW7lNKVrkUVf1FPrljVL8rdu/l
1QgBjW+Q9iSey58Y+F2WJIWCswMcOxViJ+DgAwZHdvxYUbhcBBNKGvGYtFvH
gsvcmVayFKxfvV+kGN4RMUU3vhe6y5+4HEvBS6KjeGFsSkRhGv+kSmnbRHSk
I3HswBkk1Z2FONr3mGU2juXVxxW3eJ9Mr4QmoCmeLvQkQnsbw41drRf2CtqL
7wdKJnIC24lurE2MMEUMYw8iK0KB5rUvqSO7lLwteTEGPI6FA9Axr6eTAU2P
b7AeEk7PT9wiw2N2wneflPik317Qh2nSrb0jptDBo5wtnqOg4AaOlMlE4VSl
xKxyhKuUBTaOgHuJhCLofNDH36YTm7XOPSjOZBtx+/H/7X13pogPrMRHBG5A
RxOQetgGSiU8eSxd4QTOn3tMoJM1

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyJIa61nlj5VL5/fMYSIhw+TxmFnk2pysjE/Xo9pJ1g7Hs2bcUgPRY0Yy8IuHxuw7en74shQX6dDx0vo6VG4I15SUUOOkRUu7dCoT3WwocCPe5kBlr/1TyDGvJgcQAHDlq8w0368EcP4gRDSKCHuohrlZHlNk9NfCsAHav/WowtL+ryJyYzytCzpzBfNr+Y63NqKqm+xgdqRMjrIezyRRJyEj91Fe77G1WvJWGSBksFQOSP5hMYS1oujxGoZjiqw9HRs5GjYRHmPno088AERlD775BbpomvfT7E5kWghQsgZWmvrlViFilI+/fKF8e9NirbKWwHX/WiariIh0TwNNBD60uthgw5LtK2mqq8m+1hjy4PPJH+HL3COUZE46BYY9MsbaNwFLTQ0hgpnFifbtdmW0fnsxf8nwsZxXOdZ9eMNb/Ea+j9/TAqs9jjOr8PIpeSjdMl+HSmXFBuM6aDrk/dF/T7fFK1yA0IkWbLbae8wp8YISaHVhWwyasq8pyyELFDxhB50tbMKbwLoovQq4c71Ky5RXmrNiyk7vkuOhXLRBBqEXgFaYf7EPrC/7Jqwy9EJueYUzoe1YvVzLc0h4hDxZTU2SUPP+6S6ylCImlyF23W6mlJ+uwJSevaczZER/pFPq8kRGINMJwU56ZX2xMy4WoISVWB9J2PBMLIuFTXnHlvwBUwO/g0VKCE1vQh1Iah86XeIqZTjuv4JeUYPF3hRV6RCBps3Jz5hjw4nHL3PsiX3mtAycQaXDSehMz5u5RFspeBlxxuZqLMzU2RHlY/T"
`endif