// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ExSmrsT2j2W9EJvM0sBnw/BHosjDE0s7USXk75VXt0el+ttBQ2fGKEBsMVPN
HfvXYSET5d9uErcxNc11V2s3p8vSCH3gHTUk67K7j4sbTxuAw2AxTZudGZa+
L4ESXOQDi/QaWvnAqfGOzNhxP9PPb1kBrKQ5zgweAgu44jV8kAn2CxDGVQgU
8qE42U9MD53U39n70P+XyAMZXJZDkRo33FCIHmPI8a0BCdpiAk+PjvZgKNWl
yGMnqmPovgnI4BYPb7O+rDsayv7JKmJGKD3Hq8RTTmjddxPU6zufBB202g5Q
K1aegZG8JZMgW6/mnGSt7+WW5JDynTVgLS4oVy8N0Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d4APlDnHlm4eOcb4fa/7S/2pkTG1p51sM9/GBi8YEywEENoo2TMCaGX74bh7
u3moxsCub1gtiyOmg8i3mnIG3WB/SLnu/9Z5WN8gIe/IK3LzWqRtkF4mFOkN
0Y0SvtYrg5l5pmzWYLHs9V0PDFzSK1eJWzRukp5bqwv+3jnGzb6ey5FMgkTT
ij4s4UUZ1wmARArHTmspmNETpu4mGVqllZn8XOeAtstE+n59TIp5ySz6roDw
ejO5fKcu4iwzKrifOybUpHlfyFMIYkH7jq1gBevCHVWi4eNoDExFjWGItqp7
Ak9FaIZab/GyozJ5bxPiAr9pvYzlWv8AIzKGc8HQyw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PbDqea9pCWu6Tgigwn6jD3aAgJ9pyjKpbwOxyhm5l6DaRhdS8Rz2eHJ2PZUD
0idRcxXIloAbrAW1Dy2plXY3pWA2blCVb+l8YSujAPJRCe5W/dcmPr8bDouY
s8OXsexOyQ0IfLFdfpogY/TvcCAydyMMRanOQUgeIWns6jReQbtBTKFBC5qT
yV1e1b8tGnhH/s3nTGtn5Nl6ZvLljFfuV9xycEW/q85ZK2feFnCLmkYPPAC5
ScYm50idaHuR6bkDl1dk/AuNv8weSEWFtK5ZAOwsuvjcNVfnMa+E6NrOPC8K
eAxNLsAVySoYnZgJUu8f1bMWYbw9fKiiXGPbUwgODg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gj2IB2gD+T4xnAsv4JP4++O7856dB3kanC4Y/cbnPLKNapqIgn5379fXRTvP
KRwgG1mrqIBQdhcxqurdrkLjrWGE4Cs8+p9auA1FSmckZGEIYqf7RKkIH1TS
d7d8FQWcD72b8mWcS9eE19IAACC6kD7rEFtyHQzc9jf+Jpstfkt81LNR/kIj
YeU4M+i7Dh+YQ5/K27xMbXgKrXZ7dKdLxfVhW9YevdwwVzyjeqG9MHvSW+XP
dDNra1w3jCSpau1FuAHCXZh4eG25hX0kAoWBP3L+nBpW49nSSt089GgjMMRW
lhaKaSMfzg9eLWYnC+nMhRaIU4/1EZnPjfporTDN2A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SOAIq7EESn9yvCi76HHPwbqqtnDincXwYyMqVvbQlklnAkWnocnzw9h2mKWz
P3bawGiSNa9sF97IGZfcP22heZznSduCPvBhWOvUrEHq/JyigOtdmbeWRZir
ibUiOr7agMKTUfK74BVXujpSYakHhChsEKYys+QW86Jqdg8oZiQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Qmbbwa6EGb5ibSUoLyxsaagSemxO0q3Q7ctOBp/u5ROZw1wKIEA6/O80YbB0
yY0r2xmyhgOL+uTAqqJotZerSvcQfAxcFlNpVKShzRBJKzTBtQR381eUSBES
szmsywBr8rhs9nxoI6DwevR7ny8/xoiU3b/e3CxCtibxAxasvE0nsN1lWyR0
yX0QbC+KysSNQbuAsSz8ttaYYXxAQLRtfVnSjDfSF06BN39/ihNRNbPA1OTH
uwOy9141AbdgHEvZii2jQnWAnIpCsQXwkoDHTbsZRyXykyvWSOjkjrQNeCzw
J4JUSV2jhXZ1j9jZFbAApGZKm/MvcW6ei7PS7IHwBFnK9mDM2SlzTvIE5lsT
s7bj+GDARVUEEt59/N/cYHZHr21YgfeASbmZoPv52ryseh+2vavXpdRjmOQ9
5R6BKUScHZQk8eXE68K1pT+sESLq2P8frCjztTbHLltFcDqk2HvYg46y/LZk
RMG+BhDra5xMWQicZxQiJS++FrZ0JRN/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lkOZgMideWlHEATE+aN1wYhZLg8ilQ94MT5DQigqYTJ/bJ/l2FiVeKIB+K+4
VIMmnuiN/K5sMQSW29oi5CnbaWxo+ggI0HhIhUgvdjKyAG4cNADs/PD3Nj9C
1Lro2nS5JzHlsY2H1mAco7MsvYVtML130h5ZOiF6TTAazUMGxV4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sbOjtNh7z6P0PsJCOtLLGrG9+aHsG2O5AbP4VR+qCKoU7qX5QCqU5dtC/bUR
evL+RhzQI34m/2//eXO4FVi74ynLJHMBxYTrrmolmQ9A5a4ZAeUMdij3FLOi
V2TfZVFATDxa4D6Iyxyhq1r8K+/PnLxREtSePFg4KZbLeI120sQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 58528)
`pragma protect data_block
7841eSP/cE2+3/V4GvKkN0IoQgbRH9l2Zu37qAGgLQgJdSAxK4kOVriC8/zj
FzMAVRoC8FzirPuXXLf8nHWwGVXoeWrBm2a4vx9GUaCt9KZ+EqlJEw+bk5LS
jbuF74lPDsGy+qP4fiBNQ4shIA3+PaM2WxL62nPTM/bwftGUHtAZ/JZTMdca
GwhQVWqR7YMRoxnCU6oziQgKPg27wpW15YSs+FKbSCLMJxuh9xWh6oDY3qAb
9QaHj1baV2ufYhLIxabn+jgCokFGbUCyj/OABsj1Vfc+h3xqEbPKOooiaRZQ
Hwp7+Ijmi2/IaCL9VBuh75IS5yZsGJTFgrTu7HYRUK9U+r6XM8d/8WPDTqDr
WMW5mnqSIGmR2GzyfadafcwtNkqOT8ZEoZV0S7mcIz6M4dgJN1yZpD7CUdgp
3dfb/NH71ruIPrkgx5mj41Tqe3Dsp22qJTvpnl9I1l9zVSDXUlc1QZ6ZYSfT
UtSdl0Oi5ZwWqtmvUGf3k5QxU4oD9ITvNA7uCcFX/6kfndze2NSRT6VjyXcA
CdzlmPk5PPOJjTgE0xLoOlJSLN6IpMi1FM6wge6pQN5XR1XFSmc/x46Sef/b
FiIUTN1dQpl/oKBzfrUD5L9brwl0wEriCslwk5d25vxsLBKvwtKmOEl9nEPc
f/HkDA51X2RQn/bybqlrTUySFzZYxq0Vhe8scNq6bfbnMR2424gqPgpZ/AAH
Zo0GGpxXb38GFKn3/dJ7htTBmNS9zjZFFAt/zCooBAn/+cE2chDx8UDZ/WDo
Xc1Ut2/YhFm/ZWQcRH3f8MOoLhUjIMRRSlTY0xpIAMOui2xTyej70gUiETAN
k61SWZilbTLCw97PZt5m659kt2p28FqSGcVuu1bRQ6xKFMcn8pzks7pKaoR/
Vt5VAPTPDL2uvpfv6ErfrAb0CGLa69+2Us79NGxTh+rTkuWaWpZ3FNuE9goA
zOAnAo+IPYrvHVVIzCoEhRG2BXTYwBZNuIFDHX+jdZtbMo29jUawkcceIMah
/ovMTlfnHCcpcSkf8UYJD/Z/L6i/38mztZcCEvWuSE9+vvNl5zdmvuGPg0+m
5Y4g7XDTfOkdRX5HjwSKJkzAvhszfdPQy7qZH+z2EImzm6rDSmTpWhzCFcEl
O+PDkw5crQdoIIBSskhtD17mv3/xHw1I8z5yD4Nse3oNBAq0MjklCyp5JQEr
PSEuBDPo3/F61wiXerdgGrD65CscRLsBJLIHW1bjCH3mXON50fI+ClDSYNA7
T9NDxj17m8wfFosUehyEoqN8cX1+NWG+fqVi9FbYBI8CXkacW9TOFYkMoNjT
gX431lHL9EaX6ydcLVf0AMkIIljPSZjlqAHwKSbhe4pPN3JJTwqEfFIyzH7p
bGNFBY1KnFqwEpVcSwwvkQkXMCPmL8282QqYlnP1+lRRubEn5vjeQ2vHGtvK
/lXVjSux9EAEtlTUjImh8jnaXCjCnTjKm9OfNR0x+0nXedfn9M2xWqco66DE
ih/cYn7zQlbSkQhiRHadRdyupJz3t4O6zSxr55fprI2cF5xnwk+Zx27XuZTG
lEH9m8EUiOS070uOysd1TBGSlIgQPO9q5Es/Pi58ESiIKPJ3kpIGaGZwG3Ks
Rb88xmlF3wMH6we0nLLE2Z1G6nigrOkGPEvBIaEONFyMeJRXPCUeXuyInbgI
Z0dk8E60R2nw7M5fzo07lmGhl5r9r1NPLbtGHBIulTEiOcC6WtIFJLLc3+TO
SMtWcphxoYeJ6QEgnmwzPZAaP4z2qmXGn/Cg++SMXMNb2SGq8Sy5J7TZp9w/
xJx+SOLe1w7zQj95Y/GqDnCO+xiZEZ/jtkuj6010DXcztSIr1HkQJFzIJORt
TpIAiVM/cpyxbeMhmWL7GtPGlM71VKX1zTZPaW6y4nv0qdVBJRq1PueUZbly
lqhCDRtx4w4wWD9sx073No71DwfQ2U+FgIvmHXS3BIGt2AZ2zXGhkPEQPkFi
tzcNawHXBfg8IugHDJdzbzxLMMsU6Abps9R0SsWpEqpfGGyZhzhyuCWXAgOb
H2LA1NYpEUpk4wpbt9seSa7POngPj2Lcm1EnKsGWd7RGR1nldMlnQXZYTfyC
BlXLaggNnaDIdt/vyTI1FFxcaQUUTt9NxGKVG0yJsBIJ6VwFgbiGj5zrTPsU
h9zDIqTzMVtWb+KHpz7vQmJ7Yzag8rL/yCfynGUJ2NMfinZQq1yjNCr3s9tv
mUHOTay72SowIG4Jss2qTGEkIeFr/28J2V3UZjvqK2NT3fHCZp4EWsAoxvZT
AO6xlt6gsQnz4jkSKjh4NlOJ4R5iVeADAjK3hb0KtD3RtstGzViDBQkkToXr
9VBJe/EIQlLJ9lawTdvIkGrMVqgKit1Mfs3wccN5Y+NYSU895VbuXFPXNFEU
f+YDuyy42r5rb5U54n4yP52P/jcG4yIm0nT5QY0q+OGQTC4nrUg5ecWREq8K
DsXBUxmTfrEfW75l9YqhNGk5+v1hwbe3wXgaQufFVwGajF63LjDH7aSbFQ23
k4xXhee4tFAoDw04GGDLMVU3M6gWT+9HcWxMWndRJyyNhlil9EPSQSHne3DB
9AM6Z858ZoSGxo4hLk2g2tJBaJke1+UoyUD1pb1Zj/jMUXMg+UuZSz1h6xrW
2gqhU4WCgQfmiLZCJg3zA5AMoscADQOqNGi7uPWLB7YcRVYbGZWaU9CiXHJn
FSgymwP1b+z0CAlUavKvAIrevWh3x242JHmdkIX7cCod15U0Sef9UaMcIY85
jRKP4pZBMIEBuxqR6l4fNlK85s+t7G/Vja9cv0GsHsCGW13lxMG4ZN8+VL2B
hkWsINT0OKZzvz1trXuCVa0Kqok7FJLjCItD1avncTv3ks1aQ5vHmIIP53n7
kMmYZUYsDOTkT8WJ5/mvKP/9QcjEF2lSfMrIb0Y5l5bEBEYSzqm8FkYAOuks
ihQCGjwuHkrIc2MwdWRtbF8mcXXKXY8vPmMO/DZBOY8ZfGVCbAj2R+2XUL7+
Nqro1HGUSOMigCUDIjDfTS63yoOC7eAEIPz7LOSq9ecVGpGJAToLVQzLN/mG
Tvgfhn1q4TgVAFpAJSWkG/3tvR6L2rA4x6XrSgqfIk0+B0Ar7lL6/L2Vl7Pg
bZ4sOeokn4tEx81Ae+PynaTII6CRcZak42hzCt951hGR0MTjORBAkJPdm2Ke
GiHloYylrLtop5rAzgeqGBH1i0/N8CSgILR+PJVzmqbj5V7Rj+B8PGXEQL67
YAf+Sa9EWLrV2BdUl4zQzilA4pvbXrguwUehBk3dttE7g+1UpJ37DTLJ9py4
i2qJWSF7uEhYgGRL6AfRtHGpQgw5FEY/WzjECgQ1vn81VG715PtneCwYYnSR
WX2gD9LFnNwIufsTXyi65J+Gqj9tg8th65KC+1O14N5FbVoPcEWHJ2/f9nIh
tgYfONjwwbcQkAuTkpfniucWmPP2vbyJXYYCFaVUc1iOWfcxhF0Bvj2vVhTr
EvCe6gx4uhy3+qzPtAEIK148QNh94UlFfhIUA9U0BAcWxtxgjhGXaY54/tV2
+pSWhkdIfvEZ4ydz6301adADIGWvo7Zr69T8F4SaHLFm8o/iRZ1p825ec1Jw
QQweALLxMlrpGEwW5F5XfweGvNmuYXC1OIO9J62aEDvxaILxAWw5BVE2KU47
ymERx4u9rrKVQPM0IJj5ndU9CPqiMtSUaLOjTeToa3y+SZbJONDF7WtGjlSI
RmrrI2WduSWPWR9lfgwq2TILm9yMrqH5WJzPIiLyoSenKSYIMaAs+xTtCsei
ZgxJ1anA8B35SuEk0dLdOhyFhjs1SWIeFQhpTSQL0r3XmrcU5yIWKLBxB9aH
cb7JNrDgDRbMrL5AHYMX4n9xjzNg4ryLCqZQyhwhBJbzAZpY8ouBci++3J10
ljfl4YRV/cMaQPSAlaBjqrGqCCuuTEg+gi34yGvOHxggrP6hJQApRikEKkPG
6ghEv39g7nVAS72RmqKb7WVeTZSA0eeCKPslQReUdI0xkP0dpiAF1lI67oy6
YvpgnZYRe/3USG8pmT8Izt57URNqaof/f66jHMR2Vfv+EfvXk8umUpaOXe1U
Ry1Ceb2ii17UrBMe4ntzSU1aLWvTc5/DoWdAO4fDrq92qdcW0zL8YBXReQ+F
aNTOKAevyUqXn68o7F9SJX4M4yGWnBzGhhgYvq9SHpaK+xDvO+Y5A0+xc8o2
qzZjtU3qCptzrgoqhKD+GQnOkDHbjTQxJxgYKOMkHgPtRWvrMuYIMof9W6z1
I5PZ+/0M8bireqqf0Jv9I6L2T2B12sfk2/H1kSb8OZ7eZwAjB8NsZWepX8sy
lyiniC5btXO6d+tSeT7UjJokyq6VhP6BNw4kq/JRw+j22tkOSBho6/Ch8XrI
UUX/RLOR/kW8W13UOK5J3bAVTpCI7nelfo2zn8c2KFnB1n3MeY1n8BY2J66p
TKzTNgcKqTe730kgXe32rtVIzeoyipmlPauoWEo0aOLwvVPmrEZn1THuZt4h
gC/XCVoTwXc7giOlnEI/ekQ9VpbNBbAfYI/7aNe1dHxtaq20iBmfjW6TLC/y
7XxkbYhlbc5rMCnJIDDdngxi+i4XOBnc7mUZYmu1LJsR1nTuruquCyGwoX9Q
91jRgCghfkkbgPC6efBi072XOBTNe53fp8ayFRay3ecThjQZ72umh/vhcmXi
cQDhHtjChgLlbxzhg9T2ejNJBXmhIe346ag0rN1d+hMCmJ66z50cwMZv/vlM
yXzlvb4vnTa3o4sP4djTw+jlWme4RK2wCTg39Oy3n7vkov8vVkyHPjaZIVA2
/frZYi3WF0r9Nt6PVqkTo6e70xS/fAW21QInjUxS5xQiPO85fg3PCRpQc2Dx
4ljaIJxkdfjphm3mYnxOA7cMqmNVipFEFAv1bYSv61t3yNN7D1QKtJrBGT1g
xaBXbCMKJ3MITQ0uQwJMpUK0L34gg8X0KP3qlE84+CcuCnfaSOgqXfANVK3h
a0WjPqwSulk8GiS7a0zh0ucQPwFkd2jEdbNIKCS0G0m8ustpUcu/jaNUo38r
0u94ug+lBNAkLN2J+8fOaqdBbsuGfX+2PBzUt9R4n0fOoTfKGDDFhgUNCnrU
3fUjk5XrbOQneoeZDxDvACi3c20NI/wVdcc7Ge5pqkCTOfasuCENM/mKmNZb
nCgrthO1mOnCwYEjffbRoOc/vkR/mbL6jACFw5K2+ECA9y0vimAOkMmUX331
7NPhqqF4NOk4wOJtQ/ds7pF5Zk9iDf/2jQT7WgyXbxxTE43NRWRGnyL/FROu
rjalJdEAbkD5wTCTywq4DGWF/pyjACcW490mPag0Uk1zt9U2ohNcfqfJAgUZ
ZJyC9it1yCY3H5Hd3wEsK0Ut7z9wb1KdU5loG1OfAT8hsHp+xXZQ3q0e8CEP
lepGDPS+D1/gmAOK4DA2dlRrVLqwOxYkqB/oyYhi9dvjymEReUacHDA/plN9
2OLDAyQBt1JRyGsE7FFouZj8iHeguT1U3wBR+xVItavuq8UQp3ifDH47OSbm
nS3YPQKaizeYl0MIS/Ty/rUs6iAZo/nMw9O4Eg5IdFfLbmJpVkLpijPtxQqf
b0/bV7BUl3UgsX+t6jUExVC1q8ZJp2LriBaRtlgiY+B/rrOIzgM9hk3jKrqk
ntWHAtb1suI3OapdEErD2jJGdoo2/x86Kjor9z8zwe+6MMbY26wlxWGlJb7W
FMTxj5TyBm4zRrRAUZIejBPI7WYKaU/mOiJld6nxBvmYEXvn9uiyFYnp+cQw
gxV0O94pg6lgTGnxa72Y5D3FgwBQZKzaW17UroebSra4PIfX4QryBOuZkTgm
ueZUfavXa+fwaWYRzkokxGOHxtxqylWn2sLMODs62zCuRY58ii+FHmShOV7S
InaVlO+MtBHKw/RfqaYsEkHVEpjQK/cgKM0Nlp81ZkbXIx/32BFPC8kLRPBc
bzRkUMadTq/cwWr1Eqlidw5WLzyCXEcWp2PdV81BXaRsIznweJZ4cJHBTXCr
LHUT7DMQQRYFcuGHi1zgFaPb7lM6UuqPbmSPVg5Ve/LcHT8UdeokZTnFZMCD
m6Q8FGkYfbsZQGpIaPPBc2ny2E6TwDNlcEG8OwzPQ6wXqwnW9lvNfW0uz1Rm
j0KhyukrNYQbb6/lR7bmQMWkoThIASPmV4qSaE/AJPefdGPN9rGQm4dmg9nV
utkvPaqz4u2+FR0tpaJzacjQxSZPupVH5ugBBFvyaEtnSBBQaZTqInsjkAKH
zyC3EUGnlAXVcas2zcvcHInbGnBGpHpDyHA1M4kivBmbNkx0ODmpt/qOj4Q6
wWfnBVJnzBuQ9v/Y5zToiSpjYv9xY37rP75g0YXQ4FHB1M1WTXaW75iWQn3D
ZL3A48TCuJlurnaJFPir7L64iCy03dPpUiFXnrn3llttp91gzRKNjLEs77SB
sJb5hnccBVCbYVbTBcMjqDBqn7xX+JgfLcUqYCRlS4/EngDWnlXHEp48A4bM
52w143pQ2LIiWz7r28dAk81gdXMzxTJtJu2GywgGBj1QfBvaAoelUBPpBse6
GLYEjxsrNN50H33BxEk0mtaTZTNKzLwRcpUiZXO16t4QA/SiM8Q5SWoB/gNC
uaCRjCRLeSHbZa27zPclQ4rtBMj0iIh5c2AlAdh4LKYuiSrPfXUaNTgu5fj/
9FeIoYQx7oJc5X0GzRBkYq4eGbRGai0WFJo8e7DFC0xGnkoZGPo2u1RsM1tL
YPnyDtIcDaN+ao5Zww++PeXi8V4Y1RbuZQpKBpAiG4p35ubPqTaxDetS7cxY
0ZxBp8sZUvbGW6iQihdZY2HbNCk7/AbKilUTULMfITNmQFutd5NPw81KZb+r
18smDJOR2mydKoh3zhRmKXIo51gVBS8KJCZw+4nxQvK7sJtwL77z2DhyRVCE
aszJfKw4JqQkTRc8OmCwSzBHFxcy01GsHxGz2YIz7jWRzGZQWqGAA9J+nOGc
t5IsdqP7gC6dr6yQ99OFADfL02B18Sx+aLXVD8ZaU8RrzF1TXAAWfal3SJ95
+7c7fAm06ugg/heNlA51pkt7eaU4BbaWLcizwVGdy1HCLCfChfWwCz+J8xnC
kTU71dCEAOj9QqAohXXkb5e4Fkcd6S69Okool89MHMp1zocR1k8sogpesDH6
755cOzPml8Qm8kEdBoUtKqjVrIEVO2zshB/EBRj783P3xeBK/QZ+UL4rMH/p
Bul7GK6wsGW33VccP6jF4EkgNvOZntpGT96uirQRD8b5zjWK98xx2exb5Bns
rbCzi32Fj+hjQGL5ZQapHfw/nn49q3mjtuig9XlpZTB+VfRVdHF+lCJLFGPL
+oM1rZySkMiqbQc2cgLTyNbD7xvgiBHOPK1GkC88LXygTMeKFvq1PvTWflzr
yidYf1mFE86g22t9h8zVqSlEMB+XanVCzcHpEhXXuuljLh4um7ao8cP8FQwI
S5+s/m7u3VgQtRp5c/UbM5nFYom3pSEvjYL9IIdICDgRsFqrJV0cEiNJdCnC
u3N4pj9joYnF4raQk75VphQZOO9kwjufuXJwlVJprdCy+ZyyEKC6A3ZLrnQs
dSnR6gJdHakwG1X6MTO7JWisciZ7roncLtB69efYNPsM285QGyfI+dBPEvPg
WJnlKxog3YGy9FIR+QxdbLJWMm0mgbL3aMHY8OIS8i4FAkU7d5d4owylq4Dj
XHrbq+Fgq13lcbTlGiJfEmaQ3/ytskDsqaHQWS/60AuytE9AtJwYDoru5I0D
coY5h4e8mi85XJFzoFSR0AHDMYS3eVWqOIjA7ID3IRFfYueQAgB/1egyyZeZ
nxDJIy1OH50p/mH1qdjT537KMgi4v9yP46D9k/+Jr1g2RZvhiwx/lKmvl01R
TbQN2ZiFVa7+cQgr+73La4Zrnl29kcXAQyE6Ovcwg0EqzAfGFbbbeYb2KSX5
O4eqRDYlTwuSCatU/Rz6sQHOmbjavSMBYUDnJyVGJ50VlXR9Cq7AiC8a8DGt
Wh1KxkFK9INZM/djAgDMzWeQpXGIZKTtK7lwNfKXo7ryd82DmU8WCTIvpDFj
2uyuGPyAF5FYsPF2BpDQ4lyMkdc1pcSjj5T9ZTSIEni4TmeJp6P1rNCV4LZC
joEjBR4S72lbKVctLrKeXf4Nldu8Ia8CaDOdpFGo0RUZL8EE4dEErfjjl0o8
MZJSs4hCLAXZUd75F6HFaYNTq1L62Zdbq0xwEthsOkYlRzG1zyw00rtWtQeM
6JVj4VQeknwoTor66yiBZ5+y0VzIIFSuK9ihKf1j+pWNh3EDfeVBj1ZOFa1c
IyrSkxCQYVT6Hg6IEFBIjEhLz+TdrwPiHZ3yd598QbNmqlk2cUsUObdbyPlN
gCTzvtXEnveaDPwygecFqrxbzXWE0gu9JyeY3g7IA3XTWD7ZOQgN3df+TrL4
F8kyDqPtNSnvw+k2zYXn2fQkukSTuqxayykqSuVGAAmSGEiHhS/NCOfzIn1j
Qhoqe5T42pppD0dK8qAhKI+bdHFNuKHZH+OzKF2ZA6MaNrRj7i7F99jiqNmq
pkqVmetVzXhg7a2C51BE24pmy4Rhdd3uqaXJppiFgni8e/QepNACkhFGXko9
OEuk5HRvC+dyTK6fCThc8SmZ22cD56ZL+vj2Mnqu/73/pKf0Gm1aF5rLRj0j
k26ozHu7N95btVYEeownCzfhoe6mV6dS9VB88D2rZmr8dCeamj+piOgAtROC
4r9UWGwWb8LQRl6sICGjqVQrBrIB5bMCH6MYCRN0BSubYa0Od44EC2JB0C3j
e69rNAij1qoTxldQt8fuPKP5+BgDQy679qrKKlVQB4Oq25CEyw86iAhW7LeW
93FICil4LgiXY9z+LovI7ulPfTjgBTswZYJr5RR0sG7ZWBwE3Qt69t9YlQTm
fSd+ZHksz+KUILSqvAPvNFKd43M+L6f+H0yBSN8cLiAW+JVqwHfBBER9n6ZH
8F7iFI9Xpt5RkadamOGOb0GUD4cFnuZXZZdZYRyz+pIbTF1uLd8Ia29s2WHB
k7/1uiFeDPx4H4z+rt0hqnxJtqoeH+D0AjD6Yah3KWOZ3U/VdmT/XAguq3/x
g58yvOWPPnaI9SdsVfZ1j3UP03PHvdM6A8oIENOGKJ8xQ6CraPiUCJ7Zi7Hc
FzxSWxViJzyG2oiqxuvmNdek7V7AyvPkZV1Ggh4hFm24QKF2AllDwYrQVZz2
5nvz5HwSsfrZPkmnNduB4vxjMpbHzS4Dp2g9ybhrI6ALBi5kVR3rayHfUKzb
Xs9fPl/ARG9q7LKtVBM8Ssdcf8rKcVOh0xo/+TihrzvSTQYruRWKl1m+0lGC
cWBTbF3nAb0/6gzb/SzK39ZcKyARo4Svcq7NPE7RqMrgcNuS60wKNMlkqtsW
cq0csGSOc65oX7PomtEdD1IpRyseVSbqZFd7EQtcmnOnfl7D9cRWNafzSNOL
901OWXTa5w73Czi6MrsVmCh+LvqjiVgP7tsDObpxUcgJGtkQZEA/OBA76x6i
9y7HWrLd6OeRryU+a/eEwLd4eyT3NCcWS9LrW1dXOnT+6fCKPoNUpG9r+sA6
jz3ZH3wAnHQDmU2YBtAPQSdtj2CtPxsjk1ZY8TZGCrdcT4Z909ALElbTw6sp
jBEasqJ9MDdNVRqvWEwR5iIV31wpKsB8vaFp76LwCn5JtXuo7bC3q1Gvm1a7
ccHi1nOBY/IcUUuMFQ1mED6KJRoUqxorkiKX9Sqd6kqwxZpNhQhanLzupHx7
lyyIujaE6zeGdQhyOjykP/ziAkfpNYPnE+D1pIwT5I2gz8dBPvNoQ1OOCGfC
ROePaVZrlXk4ffbj2LmE05JgxsYXl5He0Z/YcsZjGBgwx6dBB/Lar7SR3gO0
1jj65ZqeoDdC6sD6tAvKv5A/tZ1xjqcnEEtK6EKrbc5glbaAKhf4IdMbR1v3
fvrx4WNVfcZ6krMkCzu22GGfLRiQHrM+yfhLXrk1CQrPiYNTQHqHo3Pdx/U6
zLtBbV+yuFBxbL/Yaz912UNt3m0S/qyGkuvRdwYCqj8i1sDnZ0NWtZXSppRZ
qw++YLbx2VejO41CJT7B0Btpj7JqDbX6sMlArw9cA8WThYnPApFBV0GRlqho
jaHdmG3gclGJiNd1Rt+B2UsdWIYebjLu9t2pQNDRqS1q0cnc507fVTTmVqi3
mv527NBjXzSi1TK+vGbEKQuj3hyR00dS2uMIkmfbVfWcaRCiXOxO0WIoi+SF
vQbwDeEflnURM9sPjM7TBfbu3tKrz4vC4CCr++gon/1LhZX0MQHOi2IGNBKf
Dy3uS/gOIRtB25YKBSz5q/jtjVIhDHn9Wb5vpUacuIqEZTpaD04Z1w9kylcw
NiWWrr44ndsYAEKq2HVGEg+kuoZ1R0SJWXvEjaS03+uaY/pRLtrXl84kV+8m
AHmS3IOngI1tGsz3Eus8aK9d5gTOKvSnXHys9T9i+s7IVY9srLM0PRlK9SwK
vx1zp0VFq1Wwt99qrBugsH95yMIBuyJTlBlbbXvv6cdl3kRaxZu4o6Dy6Su+
mqKgPqrwdMpo+b0/frVeBDn0ed9WwPYJViEBRuVskOVQiK3Bhn6r1j6xqE4g
OUf2NeyuAv/dogbLn8dn6DhfJdDkku/RKf/gkBJ8A6zl3k21NoxjoKFrT084
Z8Xqez0whJFsk+JGomRObGuBoLEve9AZERy3ubSPhO/ETvIi+1wbbNlcd6oJ
+xDK7l5YHmeTAd/i7ncAgKJVHeiET2yfJcbHYq3Q8TElXjvL9CgC8wkRWe64
g0Ljl0U3E55NzCsrzWdCTyOICHgIGXG02q8ERuIuzR8CnWWM2x+uPUuEVjn3
OmUns87+4URSMG2yXQWNyOp3jnpDQWEr4xBdMRA4+74GF2k4yAs0qJMW0iwx
mSYLvo+93k6Wbu/25sFhGXZf+YU5Hv+1L4qsVaWuL+7dP4Xz4RLYgAMT6DmF
CqmF9lut/IVCgdmYC3tkC+2d9RvX4QFsv0zmIv4wLwfMwbOozaMLZ/vvdr2S
K32fCoId/HPFecSNTnXbDiTkhOecovzLGrY27pf3CzE2xVrQm+N3B3X6vxbm
e7NN3476NnRJrPnAoYfvOYTPSqvs1C53va7/2jUDgp+SQFeFCu7Wt4XqdZBl
b09uA3RiGSKUgesd1ejGnhzmipoMzbUChIUXeUiHBbfd8AkaO6hPt5II+HUB
LZQa+jR/XsTn/XCPBUFsdf4VlKsFNqF306iKviwPEEBAvH8N8SNBqu7v3/vy
9bsZ73roFa4fTkdvz9oLBDsTdlx9VXajYqKopzJqIQauPK8DoxGzquJ1wK5f
Vk6PPPZPZ5Fl2Zex8SSDZ6mwv+CPeapRYdZg/Z0xsYflCFE65TqkrndetnHd
4npA5V/OS1yoK2onlvZ+RwnBnGwben9/ZJXw1tQNYpBxYB3ZcySN/Vjw+RVt
qhYdPqdq6pv0MYG5c5ZWSvMYVeaZSOphw0CVpekdBOXPP2YqDC7D455GVtU9
wU6OTVyvzUNa+zxT+VpImc2bWzAqr2VjyX2oMis0nCf9mP1aecCjnpmeVICO
nfxuwadQYA9n12dPEbS73mfYzhUAwlQXp39u+9ifxz9jf/Vm9UaBjOGT9vWm
yqt248jg+jyFZNFkUqm4S/t8B6JB9mq37tY3QMYfMrcvWKiSeGglRl7SgHXl
VuCrxmNIpV/1AOk7dpHnMKvcV4kcJMLMxE3WyqESlmFJaD1IH5s282yigzFB
MhW9Nb5qnE5nHY/7p0bZAATx4KH4CKXcJUddcxyXP+gSsxanVNP67lpXLEsv
zQSK7rz1+LSs1rAqcPawufIkbV1lVYCb4QeZ9qDIvLxVvh2WlLgzEGFHhmdR
2C0MJBB7agYw7wMK/9agxc+ZaBi7aBTgKpO36drCb0UgLVzDRvBjN6tiFBXv
Slv8Ahy1BICTsetXEiNmfRKR55RulZ9dNmGihkn4tl/Y0YEp3pYs9C13B+Ja
hTxk8TMunQA80ayN+hX/mM1yVfRmXkEbFCffVeEGqj4cxZ4TFdf+pZctj3kr
gwmaZG/YJ+OgIF57H7ykQNMIIqlJ04Xozt5tzTpM+E41ZERSLGhhKUcnHTsw
RHq0saxnDDiolidvLz9gvm6pObgHf5Z6/AWtMkrCOs7eOZxRT4de4k9zzkFI
OY597aQsS5+ohtY8Rw9Ruz0jjT5U6ziYtYityet1Bf45FwjhEMlJLwZ0W+6w
4Z0Mreb896GJ4mlhZTMqoD1QywYlZsEka6MltR9EddpdqZi0TgM+WnWAtBjj
DLYB1PyucPU/JeQIx5XcY56ZEkCDTvR9svuctfd0vCSGl3wPmlz1HSIraSeQ
FvVUzxTm9G/D+5zfpYJfcxX+DwgY0I0v6B2+NeHa+LyI7EaxEAjBglRBcJAD
WAsZDRnBdM4d+frac8gyINOS0ywJil8mWMgtTsdKBmowhoOpJewXih8Gls0y
U9/P31VTAIdKr3Tmjk16UQtkrtWFbeZ9/8iQqNvSoyISxZutcuuCVS8BOk8w
NSj/2sKrahXUC8QfdalfEkCkmdSXhJh0febS+l+ifkW7XxyEC4mjHXK7wXZJ
LAbOChY7zj7ypImGeVC+46dI3BlIf2/oC4WQPGd3Hw1o3dPLz+sosbHzWfdM
9uMoQwBn21MuO7NRPh8XuApMog113bPfjWMIq1kKu4zp+tgXjB101mBBMPrT
0f4R5rhK9WZ/YE7LmaOepH6LEWECh5ZPE51UM3xA/MuKmo4iXYDViT2eOuDt
raAVWxHamA4PFY3Mn3njul9/MiG/Jnux8Aw/JYc3GazUYo/xaR1jbYWLGIXE
ukT341DStaxcFvozrYZILq0IP/NLTWLph9egWfSa1D1UnPfmtT5mH5UjjHX5
NNzMimJ4UDHRjnaZqTLbQazwPbp/n8iEcul5HeDTduLEPSpQr0TsHcpX3Xp6
yT2FNfPvtm3i5L6B1JzQLoCgc+cvC3dSzwIbUVWZA101AA3zB4FufCT1pRzX
Me6dtZFvvwqrC4FSr3TSX7LJ0NSubEvJG9K6GpktPtW1f+Ix8H5AVGGZpChx
HD9HSjPD5yfR+fTiU2uULTUr8kx/YmfvG7kXKD7kk0yvfp/oUqcmvkLObuYZ
6gM+eID/X7i+nanIRVbYNyuxecVugWIlII+7erZ6p63Y8LIfsVVNbYALW5sJ
RU2wlSiNh/m8nZ8HVyJhloj4E0sUGJRfxUvkg43IRYuh98PwfjVYtGd01OEW
yegk0MfBh9tDETthZtybO/5S9Ds4NFiDB+zYRfwIGJgF8uRiHg9jhYfKVWn+
N+qSLkPR1gw+CSro9LZoVClOXMuQmYY7KLIuU4+jud03lsw6MiK0VU9R/aBG
jxt+Ri+LMymE25cr+H9POfZooCnjAB8whgJxS94922+Jy88cFU6uQCWDGL61
NvTuSTm/j3EcKfs2p5XoEIj5PqIlkhR6I8wW38hUiTRiLtP6Q7/DB5/GePXI
QyHBLBFwygCvkqHwGmKqVX7fqrSFIFlzfYEGTjmEHD0Pj+mESLEA4SYJggz0
1DAXTaeK7AcsvP71Uaw+d2LVi1j62WsU+BPyNswDLeTn2WC+MIzCly+bhXPB
xuMVrsdyq5z7X/ODfYcRV7XZdK3P22df8lx6mdoxeTHcx6wwaob6TvIDUCh3
XABD5sJK2+hVQp92+nIUrRqUiH22ORK7G5GuKcsrLKVc1yLz+noAcOteB/Y9
QWG3mK7l2rJvgYxMeAWfsdIn9VyMlms/rP8W1bDQvcEScYq519t7yfn7PJ2o
4VLJOF3y0ppZWicT2G6BzHKL+r2KymU0WB7Es8wJGAOjt7Pttrop7m1a4qrq
3YAc+SQdTpyslDE5fVi1PsKMqlIh+HkOnJvStJ8FR/cb7qnX5pUY7xvWVxJ6
ce7jMA9Stk8GbuW/ISDzmKMfDkEpeitbxRfPbT7vsaquySrgUWZyIIlN3NqZ
0vR48DDuQYv/RVqEH6Ii2G9PZFl0nwGXKOoSR9Pi5n/VSAujONAUtnXrrTk2
q3hPGvVaevXeSC9MNH7mPM0p4WAtD3cFicZRtNY52ft9wWrqYQ3x+juJbv9V
cfBk/Qjra2lDbqzUaXGyquO0WZg8Qxq1beebz/Yj5e5FzQDiU5G4rpfpzmqM
t6raOrGz7exqX1sKXwnODr6xWtF+yPTM4yPKBfu39hoB5kER7th095Qb8JWF
cOIHAPG4mcQ/iVtyVIX1f8DVOZC12vclqnSBRJFfn7PDfJE22VsFJ01kLjDH
MWhlgw53UqXKh/YredS/h7UUQiZAxx6pphqi+2D/v/R2iXuR+XJQ/SdRpZcm
gAXogggNs+tiCfg386uvXrejUKeopAXuKuCS/Y2e0LAP2RogF7x1ed1aRFXn
9nrgPiCOW18HLkrXXMRcNdlRQrkSKZCXaWUTBzdRroCsQYofeInry6qEZ68Y
Uj4MUHJ4ECn20gYC9xtNo+xBXshwkfFLxuUizCSRFjsLS28HhWVZ8NahKoRV
kCJ9qtekjhNIx3oevWT/8AbGk+Omann3QBEnvMlYwpTR+Mk0X4pnsSHWiEG5
vOQdfnxaMNFcOVYkRA5J6UY5sBKnYl4KuWJ6/ZitvD/ksvEpjT5Hu9UFO8oW
jgtgB2H6gEvoztJ68M/ih2DF4JcoAvtwnCXla2FYhvKJR2n7SF2YO3zbRHbf
cUY1OLTM4b/lVi9fOj01Yz4uPupXf25hdsvl6xf+OU3jQJtiQxoJqR6/hiLz
oooallNnm7PFS+uCBsczeHZDZq6oAm6zpTBNniEbfoqlMox4JlliUx9uLAr4
JQKhYB8ZXbrw08Uw8mWmddITBHfxNcba1oRTgDVRRvMOfUCodQPoSz78CvSK
yo7J6tYcZDuXxytEr2krRX8e4UheAhewEtFKaeLHYxvS+LpR/F4kwBh4U5xK
ivNkfc5rinxvEbP1llwPLZywk0Z/uF6AH1IqyYf4p6fsds7kJRjJxSqBP1JZ
SYzDwo2eAK6Ud1hNHiYCtgamRouviG7UI8RuxngBcCJRBjez9yNh6/eIbYoA
9pLsJ1VAlSGID1+JqNTaweZAchtCcNuOcEbK2GGJ4sqDGtcVBvObd1Bbadzn
YU3BXPZt5E5UniSpPTmRCHOcdHQq7dl2BWG1y6KOJobZDHRIvVaOr/zWwhD9
vuj40qH/2AaT/BLh/pzHPk4BDevD+fEsAzQC0Yl+TQc96COl44SBbPIjfJB1
T/fWZU8zvUyQR5Xc0FyvKT9h287BfZdr66rgexSbkPdm94vgDHV8Zjbsizq0
O7ioClZ8IXkgUNyGZ8DOMl1NwXTa+eYUU0t4dc3RCwRttgEV4lywBfIBpbmn
MIi8xiK9/x31EasHcvmYTl2yV22iIt8mGIaunwSAcQBwj+HhkCbq05e6WkfN
6RZh2tsD063ho+fWg+aCOgwH7IhiYxn+vuQLZJI0IJ5dZ18RYJHFari5vACx
16f2irJMcyYXYBl/Q/OpZI7u0xdnG6mu/f/+efIdgGB2XYMx0ivy8ssfpAZv
liORgxNXc5JGCraFhips3GVspbm8XPzYWoe1DhKGPY8eyCfvVFD1aqb+kJGQ
8QrX3HICwOFwIFS0Lqak0dq2iHRGSa6NxsifklEhZS1k7SABRn05WUpsDIj5
joZj1gnzcP2jBkwhe8J2+BnUb9Vp+v3jI+QP3pkV7DrlqMmLW3oT6sq/qLlR
t/owa5U6s5d0K70jNjiqc/XAhW6KhgSsp27n0CE1YA6kK9YokfxTYoeWVfEo
gojWJcbP0I/feDEnQ5Du6CsfJhvti7dh9jprIssMm3tJRBzkOXraUT3KhoNH
/fVcZp6M54ldax858X2QZ5+x0ZDrv4WNxDU4sjLobWXhJDm3aoomgDPvlnpF
DFgwqMmiPzhoifVtkLUkluxD7oXgeh9ta+yaLuIYZNR/LzEQJu71KxDVCr0d
381MyD6RzmjAUb1a9hyYF+hpMkyWCVQUi7NA1vGXWPZEaOqtbxU09iJmBc7g
lct1C6cA8d67kBVJY9cIY9+zO+DqIS8lZidXihaHuoB8jKTlfe51rVrmt+KF
UHh5Y/pNjrFbxmdf0SVN0VHvDUuSqjMem/sgJ8XvMW9kNn+7LaMMBgoVkh8m
7RUBRg2WSvB8FsEB9CRtOyw7YS8muxjl0hXbILtP/T3NuGWB4Bk1S29IQYCA
Vc383zrQGH2Zvzb7N/igxmXUEE5bcKGC4QtvH8MxzDey5vpl1WyacHgJ7iA2
gL3/2RPL7Gi0ElVpKQclytcyVA9VNsW2Prj8Fhz2DxjlWun39NO4jzrtrJvs
duFnolqbzeiAw2Zevx5OczlDGGa2+Wre4gFf+w5FJMhpZQjH0EvBUcQLM0cO
nWuGSdYSIX6Fzt+JcR3OyJKuWAfrwxj290s9K0S585JDv/TWTsn5EeluQM+2
of3oiAVvK3cdx76VlKjNHL9Ju1HL/GGvnXAeJVQdl4oF0HgggMt4c7PvZ8Hx
8qprXRNcUdzJ9I92MiWLby36TjuJQFKq4qnAiveakUDfi50OhFm8RSaY+HKf
lXuQ7xIkc/MhHIxvwjdtR+Rsu48ypurILPYb4wzu7dvlXc+I8vniX5+eggsp
P4+ho0dAQ8WSVoD9szzh4F08Ka9pOxsgwXcttPC0EGarDkxJyPCatL25t19U
PIc2kQ/mHiQ1MSrTBvcbmzuQfOusHc7THuLoqb2ghiE0quk5lW2cwPquNqMA
fH8jJSLFxwhkg+pNfvxMqlMInIOeVCILegrqIwz5ssDt9oONVvfBP3G7+pvz
HGipTF4eAkSxh9ph5VjTb35k2bsQU+nxOD1zYIO0MB8ozyVi+QF8P9S+zRv6
l8wyfOVd/NBAYV9WA00LsUU5JHNjI/LXqGA393hHq8ndoacItrlqsGG4dY3r
Cl/1nQPXwc/+I8sxjHTFuUaFvVRY/I2qfgEWpsGlnn42UaJ2P1sienTA5CwC
yMcVcqTOj7sknDprNPFQgDFuIAs1J/OlfUHWgR9t3DdphsRuzVze7OkU/eBU
P8nUL4ZCJJGF3muT9i455d7/1wzrFW8+fH79CFIfFJX+EzVLScjVb8CW0E7n
c2pRtyKIY674VfIMaoZFgx2BqELozJts+TAtwEY2V3ajTt/dTvOxshql6Hug
ZgsPvpVDjBZv4N8hG6goPUYrqDKoNbwLk3f0Z8fniW9U8jRYksjOY+ZKMbU4
tyEoBKrGf8AjyRq6JNvMJe3IiNzrRafX4+vbRVvNc2QHtSg87qPwgS13p0Sf
QAjJVNT1wvYKxsA+UW/WW0n2+B0K6NXYAMKxq0VUhSDI6hMY4ZQWqzUg8Mz5
6uFAB32zgQ9dJr+os4MVMUkXMpAcCeJjP8K6exhMQKj0fyw0zN5ss3+4BDUB
GqQGhmKIKBNLb4DigQO7WSJhvsHKLNznmpqlv+XCWtOY1Kiv8KsakNBRR3re
v2JpobddFuCn6/QxBllFqsLh12RtpF6nmNBAkAtMeszIfHs5qfZZgcQVYy0Y
RLCMRqQ3mNPv8/cPNg+sM3d4sxw13qRu6VINS9BYohjh5DwCKz/+60y2w1K3
Gz8ZB0oiU8t0khmkD1cRpy/yir99dppds1C/+pugmiz8fnZ0ihinoSC539VV
cxb18/LG25Oneh0u+PfHkiekOQPyMc/H1vlGQA5peuJNaVWrgGnZb9Xi2RpR
W19U/imIdpE+MASt0OQgGHJcankX15qeW1dNCDtMLiJU2vmQ3xtVp+XXaZaW
EV6oYyRk1YykOxQSvwP0ZUo9MdG6qk/eKIIwNWZoE9pHfMNtch9g2McOL4r4
Uq5c6Us4bXMjEVKMq7+N2I03iAN6/ePks89u+2ZPb/IBgbW4JtEeDk5H47ik
d8mUUfSN1paJPSFayuep5ehtMESy5oq8MSzSD4eomYM9SXM5ykz4SSVWagjw
ouExMOlKP+NWaov3MMi/4MgE/vvsI57/iV74mFcpfd08bAJN9DJRCHNh2IUa
uWTmc2akUH3gM6dRZ9EJt9hlJbEujl0v6oN6pv5kJ1zgTxil6m9JDq4Nn3H1
yGDPCRiB7+wp2TaRQfjnsxlVdrkPcoNUdm1mgS73X+WTwNDNQg0rTPij62Tp
4cTE5aoc+ri/SNqhyJ65tPOxmTE3GKd8RsubwZVdQ/NVAa++2lbPhLvFPpRq
1ApDIBYV5HyXyri8s7CL+Xr07hckObMFWeERhXCc1Vd6EEUbR2BwrqxrkEkN
aaAc3pRPqMeNj5L9meO5G/TZdci09G3rBE2A3k4K4PBoQm9EqblYZS9SXZa8
72rV5eU0u1mks6exXA9pf0zD+/HB8zNmpRf8yz9+SDnXhOlDla2eGodZrPdO
2FIdKX6lyWEyaJucBodTAkg8ZRQxykVI+djjOGA0bu5fK/OQCTco4eE5WDof
s7OuqaeV0pCtT0v6wkl+3zyX4zBUTcyS+cvjJ+/AxS3KdoZkn311Mh21fgi7
MpSJegoeknNgdADfayKu9ggjJM5UJpMlkaMefnYKZ+MVPZo+dVhg8hcMKVaB
xJgvcce4LSzpy6GtrUxdCU82tXXa0yW1oc+K0DWI7kv3B4amFQAMk+447BaC
ufKYbeHky6y3xMXNASf6rMLQpieL7uvxP3FX/VMFZj4X/ftzTK+hTvlAyTQS
HlxHC3Hy4fAeDBK+1WEcTCQ5Y+/ClOrYjycDD+57HtkBby1zk6QFrIknn3GH
OLZH5dLTqPf6xPK/+Q3ybwZFKM5VmOVlWPrIbcLKCS+Nx2pkQDF8tdZrCv8l
GWFw5cWNmr/S3nNac4p7NQGuIDaC4rw7K2fGqUFNwGbMjEX1uFeveieNBuSW
9qEuuA7PDk1ny+gZwq8lLNtrjdVAO2rJgBCfuevTgSOmJ5K/UF26lD8IfbzR
5ktILnXsAbq2JkbYB36LVZXYKQTsZ3UC/UX0RWO9ZT4JIlov9RCJmrFN6Igb
uG/vzqNt3FS3SrHnbVq7j5unDIx2yUOaxeXJTyN1OH4iK4MQjGQ1GTY2BV+K
7DqrZNQHerQB835GJQ9MbtPz0Leb48ibQ6suS3TVjVju0U2qjsyj7dI1/3Pg
DMmxRV0inDmsSO5DqZMrd0QAkDKcvFFrSJtsy4cizorp/PH0E2v57WqQHKTq
mEMLzZeZE4nvJntP8Z8FBerIBBCc2BYnQEtcgpQzZb5jWCRKV0IGKmBpWEyA
ASZrCN+fLenCWAX3mDArZuJxOxZ0ipnIWTjTnKWCf3et3CBGQI6LYqPyaF2f
J7JdRBdCNZGzKpPK98kgGzIzeS6FXAKE/WPpTmO1C67VGNkv0MIjnA/W1oS1
56fLBOecMj2kE9d12mM5J8R9+RXHQJyuzZa37uTWItZqWtV9JitmTJD6cN6+
K4KIOoK1Q4zNdwfOf7kK57LQwQHPfn3U6n6as0fWSRtiF3VWtzhd6Mj0pN1f
FP9U/HVuloNcCdoK6Q+Sz19SnmI/LXjZmk51GwR/Co+5G7pO3fRRij8zvrzk
vEARVAYz+/EreFg6hOkT5bJWS6iUxtmUo6qDftBbhUZ3aAvbubp+khlQlYXD
jGlvCZEWzW4qkajSbTyGF5UzmY6HqLKFE6hNFMWfn9tEHGSbb41a9XhQjvPJ
RkzM39f7BqyPc2zVxmylj0whMl6Hcup+E+2D+XqffDNMMSR3mGXOf8AmrBXR
CenOqOU5YO3oimvZFMUPKhvMVqSwX8IbjJaYyEdp3KGLh2KsO+u2+bwzVDfY
halc2NopZOVsTQ1yKcCVfTYSx1XKFiFlpcOjPHm6LktMxz2S9aVc54hmiR0B
w6GIQPy8jpVgOIM+eHqYg2H1gK+hdVHbeYhsZUbLcoOipgpp4b13FhErga8/
RvMiWHvhOo/vFEMBPDtmONTea1Xy8IT6TxmgHjwiBGqNdaidWxoLuSoOrzA7
QgLduKUFlE4V597c6sNd0nkSLu2YwveM2qjziVPuy5UpSNa+b1li6CpXIrMT
KVLIFzlUefnB8tbYRWwtgxYHERxbUtGd2wHT3iN77kzrbErgFi1zMI+qgbUU
GBfV3i/DyZtJrdPE+kbY9Nf4RGqfEXHJu+R5yYYIA7kPz+LmIRt4vaZCGGzO
FPvtdzg9mSPgYuC7hJ+YzEfQKqHUWWPP5F/0cwArbEdxvtlSXWempfPsZAe3
jMu/Mf0+l1pP9AKE0QeqPZb5nyiTyKdJPfk9kbgb6VA/+2ykdGOLtfYFWPGh
bGIQUPyQkXjishT0uXbFpDySHa0+0JHg21uaUr5xU64kJaqEHE9wNJIgVUuE
9E3janroQAaFBPoMHR6fqqWscyzU/pXYN2ff9yujp9+tueoL6Jb4feExjAgW
Ilp++f76lt6MNmkylFEIt7D5BdLYxsTfvOlUc5TUMeTjWIJIgwGFEpvOS7Ol
ySAXBQ9gEa9IWy5OlMN9Uqdn++hNB+tnUFs01deDA6aNtWUyLkrjPLQuM7Hj
82aXLM7piagdQE7aAEOy5g+zJH6bxO2754pMOtNLnGcC0KfLeDC5ECzJ/rwV
aSKEkaCXCYn8z5c5bJ10FcjNMTZPSGTwlkLS2Ox0Zfd/IrZ37F/XLxM0ZZUg
+Ww8UxSw9teWgpFJtEJPdt4Mdi8d8QXW+xCfWiyDr258xKsXiCl0/uqEYkGF
2FZrOVcF7CBe0K7tTUrNXOpGb6mPgebTPL8kXI7DQhbE1acuguqTUxCiFue2
KoagM+UVkhkQoMPutOWSpUXFvQ8RYY2dq3J+zL6sq4rcw3yJpmJpGfaGbvrt
+DE+q+sxhtWrHwnM3AFIM2muyZYTUWjCAXhjCTm7OcEkGQ4aF2gYbPOP3zzH
PRneawwUolVcBUXWIJ7JlUhigzh5lxvWgtqZd9thIhjHMq1dRzJc4maOWBrr
8T+lAp6MuVbgR8YWAq0sFTq/eOotLXv8cPqyXfvzlu795QtFeSlT3LRmgDc/
roRvpqZnRltZpio2mgbnLY+4osCbN2ykZhV5WK7pJswLE+393pxweNbbaMha
xoJhjRi0kKG9r5k9eF7rafEjkO0Tdjhtdq0UJ/RhLb203azFWatRhPEG8v5+
Px0CXY/SXPVzsUrU6i1uYK5D6sVjErGgQ7iyn9CWCZYQ9dyWszQ3e0YpvF5p
osrrUhbAZo3KuKP2ZhPZB2tYuVTFS+ND1JnFidY3mD7UzaHHtXupBX+F/ynG
G4xQNdA4C1ulntpSRbz9Y4VXh02QsUWJ7jOl1B3b2SaB5P9dJCGIFBmcIYSU
jtsh2CkTHJJ0OFGZYVfRCOvUA8dG+VIH5B5NoIaWqbVnTLqo7jr2dcyf40f1
qlhN+Z5AiXT4x4CdWcdYIRuVMJ5z2A7ncgmnzfGTEq5ycyrX/PlfUPiSTmyY
veMo7jN4bemXTlHafX2tYUVLf4BjPGc9sAm0BrTfG75IXza/fVq7KNuOevRl
mcKxpjvqvaIbonqdFVn7eSSxwtSrfPXxsjLgXemmPQ20Bo7suxNjS6xsp/+G
Ve76I3BG0BRgYsZ9aTEieDYcT5JcHGqaDDcYfBe0Mkj+SATFESHNttn2o9bn
2FjnoNemwBeAy0WdEHWVv6AsEuqCnpw7viHNOyux27vPtiBRpjv8LI7S3tdu
FptgWKWgMg56Yt0N37x1oQJzXZD5M5NIcuZCvkaMgs90APd4Zj+1D8eqUiyY
AmIK8O+xPu8OSH6yZooC7CH64DbzM6U9Q8GLPq0d8/BL7HFc0R1TMp30uVpe
KRggvbr83A8i5bFVaSajyaKtzcp++uNDFSantEqLnGXq+ipHqt3meR4lBe79
UTeRaxi5u41lcUpEBvHngpSkOxvOAkZqxo3B4dgvPENfxgOgxVo69n9fyHxK
SGot0FSXD3yTAAxBqdThXMJfqsbsSGFFcIfSiJW82mFj5IUwgf1oLyy7mCc3
R+ugmS/GkFEqjg1WJB3izedcAuZPYYGB65lP9KP4CKZS5kq4C1THv6QnyiSS
3jsGTYh3cvNU+RSpRjaJg/qlK1UdMrWUEIzvbZOkgNFuusMi1xpLSDWq2uBj
aEmHXY/2zuXjebJHzvyMbadQGemKk1WZ4lKCdWcPKhg0rupqefataJybKmsa
Y6XKZB+mwYegdJzkLs00xDBVlhxhcN3X7wORF4Us+hOZ9/ZzCWy4EVm5sFAk
gZ5KclVmshynq+2Q/EwdiEsIcv+kfYVjjqv3YvaowFeMYrpNX8PpVWKdjFF7
qLtNPuwQbv58yxwb16TDFEigsHXdTw1xz7Q3NNfqN0HJyI1RnQBP9mjn98zw
hdJSI4Kq2OcWZWgtXa0+ORNrZv3kHTZ292kClDpN/sC5KtP/08xOn/mP0bpU
XwkvXnWGDRwGGj2BDELbaKFeCrnlJhlRgG8wNWaXzs1Hzi5AdY7FALC7ns8n
VJGolaX4vxb6xR4vlhNsFwlOkPbW/ktCOO5bQA8hhHnWZJtKXkqBEoIFqk5t
kqU3VlJYlikpjok4BJFTGSLp9IMBoDLHC/bhDZi40Qx0AjpW95VcCakXA/JQ
hP2SyvSBTVaFOm+z63KHVcounMVhAfP3EZBKxfrr3izMRZ6XvrpdH1nOHvL9
z7dnuI3n5h6M97M2wZIR2ekhPIkWeB1TVbPKAEJJRK0QNqPHJYuS/ovYsspl
BmCqDIx+2aq4NyvcgM5oUoHomyNxFiziRbNG8Ha8wgdxcuyvceeLxe3IpiQz
PxKG/juIQWvqotSiShVNBr6HGfbMqHtoUB9DKpHZrj6HeNqoYq+zhYNA0AT0
vmnpQDJOO57kDXug4vdU6DQBphXgxKDd9iMsRsFrgT3ALdImCiJR7jubIVbm
tL4AbG/5Rg9SbCMYQjPKXwbyEPqeME09VDQyyZGGlyoj2h4WNadvMSTn0yO7
pJQPZ3KJFfXe0KgCCc++rNC4Org2g3Jzb7R2IyaSo1rg/y2GfdKebNRQMcEl
tA2v3MzVIWyfKDJeW9TrXut14lLJOr/9u6JEG3+2wwD1J0+TuNlC7ldxwMut
rvEf0bI3hjbrvTd7IWQm/ny3AXaPHQbkTR+cCKkvSxcyxW61zfKIq10AsLXD
/4hJz996bVECHVqPNYb36c2rwu1MjR7mW8c0+/RQX3tCYhulJ+cPVf/SOt/H
uX9BVW+EJabEc08jpYasel28We+SZpl6RzGcbkoBtEuDnW/ogabr+1XyBkLn
K+/i76PJHAIXkKHb8zRiR1jYHGhJl7SpnWUoEefznDceL6PwPRDwYF0rdgWz
QccN7xc7sLXg0fI2HLXbnNnb57kc5q54+4Ax/eOh0FvDRVMkuwYvf6E2cldr
m1J9oRDYUfzX8l0GoANFHwgqbv2qh8Hok43USI+1qAoe7Jl1rw5TV/w6j3yt
TTBGlvOKXiLk9aVeQukudDWk9BMGafiKXRuqL4f4ACnjyDw4mSa5S5gdwA3H
G4z2WKE30gvCUi1cSFINU6n3Yb9Srd4CeHlc9enGJsiZYEM4AB5XbKlLohzx
A+8PMvelSRH0k0XtMQfKrO3/WS4Heu+L2ZpEHAcd+ziEwBBhc354eiKEpq6C
XqgzU5zmvOQNoUBxhuJxjKuwMC8kuMOX9fc3M8sGZBSRDh3/UyG4id7K/CDF
EgDGmm5zblz3pQKz7NeXFDmzaF2OLPVkGWwBpSUjDp+T+2p93c9B0klfKi2V
koJ8++UzDsJ17IcKxk1wsr9JbYHCsWCcm84HlZRoYoHHRht78sip34h8EdHK
xKe05+0BaqH2mkn78JTC0CDrCU4Zoc1gpN3nBJ+LrGpm9gpiVm5vHQGpTzj5
aE6d/6RsyGgQNX6Q7y5AEP3HlH1i1drTkzIqKlVsoaVEciSn8hQsavtycNqi
1sw5RxJq7G7XD1mV7GVLvXgYediZhKS9hu2cHvHsu9UF3sEi/EmPNhlR6KHt
wuuxYn7U497Gj5VX2NXSY0PBsWTg7/3qrmUTaPu/RJu75ShJ07wVJEKs4cer
ow3OV0X9dt5XL94h/kOx1xCE3YpPqcJ39DMLtzexjZ/60mPR8LMBtc/GeJte
0mnZZFAZb7PwPd3vNhER7bsLMaJWCtr/Y+BBpo3fkdSM02FCDNnKZkwOa3lA
MslC+3EY05HTfkO/W78hguLLP4FjOMebvv5or3rTf8e2G0ZUFM7+7qfIqN2x
kk5w2/8WkkEquBi9bGzByw52djMACMvWJp11fzYsf6a/KMUMhosqOTcoN55W
fuwSr8TtpSyHMbvK5bjlo/qAjfu7uFaIh0JH35f3VUL+NuYUneoKBhHRGnj8
Sd8gzDzenOot/54ddyIBkg6z56HgusGdnbFYv4N34VwoFFNWZJE82RThvuKc
DreZmAfEWm/91Hnc/PswRHQpgBwfqwgLc6HhshthZl2mpqcPgeiQhxcNmcJJ
/u0ZkSzF1GVQVpgJ5HZ7d3qN8foZ+1Ehfptpi4ZRvrJFJvbQjV/gXiXfB9JQ
h1EjmYU5fLCYpl/xyQrCUgXBJJyKh/dZzf+MGMRHMueewsXXD8UKjrN4Fw/S
Y+eomGcHBy81slE8sD1aD2bOMgdT32zuF1Eah1z9MD572M1W2r4Z7PTFL0Ft
SEZafPNTSX9I1WzfwXXWeox7YqMtceP1LBaRqMz7oqRFe7Zw3a9EHhSNIjFi
IkA/+VlyIKIwN82SV79YUc8eJYy0ske0Ih1kWrtcdvZcU0I/7xDNkHGaPR3Y
6mLhh70hoQECMgDm2WFSOSjAFyppZUkkeTg/7EGRwTK0H/WwVIiGutJO4OAc
7DR8dQ2xH++pX6+fOly9Zw9FTvajI4vGh/GVyHfqERyKXcraSSgnsFR2gnV5
RSV34vrJ1WF+aH4hJ1AxQn50q9CZfZnt1/ZghUFfCP+3gqeMIFTefMqnU3yp
2MGFuXKy1y2HdQ+GYAP0TRW2nEuO3f18RyJo4BvfsDHSJBytL/r6fA2xZCEz
Y46kYdccaBXwkiYMT4y5Okbysp4ToDOcahIVXpWctiaGNryNhQshjBzhGkc/
QhuL1sbfAV+LoPXbKjX3VpygWTp01I6hReugaCycnfGgHjwyLRrq0hZHk7en
IJRXMusiU223dU4rwEQ9Tcj69TaFB3qvEPaKl46nde+LZgwh9K+vhda0p7z0
QamUE9+UjoBEZbLmq9HeC8eKYh/zHWkaeISTexs+fb49wITiZPTTlcmU2TEu
0JHdJjziAAYaecUdPdHIeQroL6C6gskLEDb2cPAwL0PJ39shkOghywuoqwBE
1mtwjW9zkKNa4L0CEu2QDaznFY9xQubqbqrpM+PzOrDAhc+HYsclL/+3kZ/0
Uzqjv4VZZEFirZCrn0ztsO8NWXSg+FHcnN54dyrFSkrSoyx5JMg65km+nD2C
9FojVyZCrMaRZB0uA55G/8vLx6m8OVp7I6A3SztBX97kAXhYjSxeXK6U9+7q
0TnWKtw+NNx/YjdCziuBkjfXHPf0RlpCUkfInsYNE5VIyr+7NqBnlMiaqUKm
FwMujQShKYIBD2/VqIvEoX2HsEVrwVTFoq/TbIOvKXsVyd66WRPv/xyM0wfr
LoLGjeA5s42PXyE/b4392gXWBpi1AHVXLQpMuUjsNAUncJVPG525w9lQ8k7S
5wmugd5RRqRDKPLl4wzoOZpvQuVGpXGmLe6eI2AM+3YZ29Y2caN1hLUbDd8U
W38t0FXRsEtK0fAzXZKJplyLVJL0U1eHTSj67YYfKNhRik+71AiBAUZaQGGg
wuFaRK6a/UxS0k+54gMnxJZhV/DT2/FhCneAtyV6bS72Me93nM5zc8fh1XiM
CfsEK3Nm8xZznOFq+FziqvxUczR9MbaRLY5N562RnWm054jfZ8/OGhKcP9/W
3gWHlq19oDyIQUtnYmQDjyypUjV8V8VngbIbXTtDgQ+hz/Ol657oZ12W3A74
R140ZRsvJyFmhT42u4yA8UX+LM8ouP2SjtaiS25IsCA1D3FSHDfj/5Gb7Cxy
rN+GctiojqRPAbMJBiqK1RU+keEXG73zReT+Gc5LueMSFVqlNl937uWA8s2T
0c079z4E9McNbHCcOw5RxQCoyzeT70raretX+xqcfOdu0AkNCkplbFvcDbRW
XCgYbPviuR+Kb9kZPsAApBlklYq6eQ6my9Wd6kjLOPfTaqMBohQmdHodiwhd
jUX9dt3w031H3lfVE6CkM4fPYqTcJjJSr/rY8I1olTUz5pCH4psIiTd7iMSS
RS5RX1s/uExJe4wiy6rf39rMRTRkINJzrL5GoUxqNJVLvQEWpMFeoVj8KUxS
YqKHn2Sg1osoRiadJvkJGV0NudPiGw8aRcqfgpTho57Ye6P+KRM6q8GIS4uM
xH+mh8+tE1UGC8Yn3YCLvt6XkqvVUrYpkA6ki8ge/cLe93kVcz9l5TqfIdtB
gOXo8+knWhsmjB09d55FcHilGPVHgjatA4KBKi/3CWyaN7ofrK1O1AJJAPMM
HMkMqmrKUfPnq+RnSH0i3b7tEChiAQjz2vAJV47uiZT7YSjW1Ja9sD/LGFDn
a9LqV+L4pCnEj0JwQEK0dHJt9qaU7iSiB/AtUME38Ump+CuQ9hzUo9Z1+KZW
XEEExBG20raIgrE8S+8Jt6onYHHWbGUu1grSBs96kn6uTkZJvVywE1/dMS8/
xP3RswdwPkS/BtcPXqjcTXTUhMeatHRyprILI16uBzs8+1E9Bp+l15i33hye
EYCavotyOY4ice2qasxJTBvAaUx20ono4e/548dCkFpXxSwBUQK7pBmmiERp
ssNZvzV+hoki2HlKBZfW7dWoVC7uxqHAPi6oI6SMCgTNt1c8aVHkGmiwa9zv
C2g/wTxBoPAnN4rLQwetqw0o6V/HAunJA5M5GcgNmu0bvTn3masFtldSGm8l
uz/eSVnO6Z1vmUmG8OMFlur8gn+T1aHall2xbr/0BbSDnzjnP/QMSMsINDyF
mNFQK5sSuN6C7+hzNX+R8HJcAvPs2KlqHU0gYiMjOBgg0vxMRbOXHK/TX98T
WM+YoOfNDdBmSLR1puIny2Q/RerpRkXJZtanVbv1hOYJEAsAgdem06WZcgra
VSMVsukQws7yl+6gMwEQlfEsRK9FIhm53LNNuTvL7qMc1vUQAZi9uwiWuuqr
2M/q63LDAZuOPmaqGoubuIjfKi9wVlMttEDmTc0XjOm5eH8CudWObUr2yKvU
s69Dv8NgGA+xc9Yv/o/LebCHmJI6zmdLSkJ7PapFQUdlFVeC47CBuD0nm6NH
qSiETu6mnIUMFWPpQWKxPe7rBHokRIn+7qWh2kw9/Tw3ZZiJ/NawgGtrs7jv
0gXpdeIlNzKKFH1xa21f7kVZsHoLAoKI+bkxlqS3G3fs4YD/FRXnhYJMukOM
T2RoQ9Eax1gTqF+QzxZD2qhL8o2y9ZjzxnL0rYOugWKF32KP3W+8Ogb5Juok
cSnSNaYvU1bogGztztiqc4qYo7T6xfYZk+gcPFfWkpW/V+Fk7ZWLQE24Kxpv
vuORfQWWsjqMMlZ5A6k0o5OBk2Miz/H6EpCKCaIUj5L3v9/7XUMqLFlbJUAP
lOzERzYnlk6sdYPgO+qDEBeORjSZ0II3dy8MGM/fPI+fZftXQ4AH02A+LuOj
S+X4BlOX1AZ2sSEVVPuL9g/gegT+BtoXZLiZXszukK4iY9FGKje2zQPRvk8v
8GZ6LC4G/4Vivw9T7uoM+mvtK3YrJ3aakt18M2lNxIiHWy4CD762u5tlxVCc
1R0DwzKMChxEtlsp+pvAX5fmvoAM3OG7kHVP+2ljQ2pkPcns/fV09QNYLybP
0lnuIaDN2vZdpUE/AguCIVI0ufcbnjuexYSLsMWy3/JJaAj2uDwaI4eocQa8
VcRebBdbyuuDie9aDIePncvhf3hIEbZMzNkOrDbJytiXuJndWOwvsflPRFHB
El94bC3Z6eWbqmuPBj7RHKXN3YlJfgG4fKN1up5KY47u2IQ83LJaEROAQUEt
qDnQVJ01kKUd1eqEobH1XJ5hxWiNlf2lnDHdPfsNTiEJQppI3/sqCOoaIbuo
yqRCByYnVecZCKUMg7LzpgYLxSqt3973K4oHEAt/8YnPDrGjigMKvRruJBig
Y0HfksqqeqpjULWvBo2RivwWjE0qK+YQX32x/s91UqSbrROBoV7JGyBvqLU9
59XPRTG81c1bnIO1sX6oSANYCjlaWVenpMqB+JQjjSu5DH83OLp3Lobj3Na6
+azPbf1R2vhhY4cC8VCxcxi6IHvtSA2tnlziBOO+UwYX3R4591exGoEZuzdP
dHkzetI+BlVZndXh+9Xb8BKtEzHDF3TWoiOZTF9GLhIGtW+jqkSZ4yikBAOo
UcT9t0DAPyM5zIJTUAz1ZufBW84itmNgJO69SzEsd8iqXcOPL4Mpyoc5Ps2V
fYyM1PBjo75iTHKz0UDLFAnPspZg6OLEDv2lTfY17P7M7aUtjBdXJxDgExN1
iHvsjNzfDjK6c+cffK9oR7Qx8zS2bNJcT8hRtwHO3cO2qkRea+q8f12j/P6e
o1Fy1F4b2gQbo6yzvftQRpuq6erM67w8yrBTfjDmQaznKcTCxDcyoq9k7Rie
z3CwL70Q92ySlQN9W5ZNZm644h68HFzE+wP+sNuyP7gvKx2qsENG+HLXMLzk
whXMR6jjdh9W7vYvd/qEjW5KfGeclMtklNcFGjrG5lKjaySZwp/sq3YFDyYn
3mOjoH6ZsDwjWHTW4ZQkMHRbFJwb27Dbkac0FxubGzkurIsdmsqnr5UfO5np
GIxbk4KbvYP9crZncwF4DIdWml/XP/kyMGGt00j/vT55C3tFL3dTu0yYKYkb
MIC7m2/6/ip38XuzGWbRa9ldzv0rcR/3kP8Qba0YdDPjZyRyvZ1KuhUBT5N+
Q3sHstrhldF9e0sJvBkQTARlP0mHq15VdOELifq1LnlYN45Oublf3PVYHti9
fktmKn+MoKozrVrMlknwG59UYb/mmbtIWIghB223B5WwGrQz2rozIQST2zwR
1jbASrQ9YBLcLoSDlX9/vhVghS/na4NA+kBkrWK9l49boi4cq6E10Pt8Ec/6
prOshcG+FMOlW6JN3OzWlHcmc/fieW1ATimYAMbRbxu8K0xab0i/t/fe0Fp4
0i2iCoEutOdxVUpdH1lICLNCMwblXcrJMfhwbCZ6Blt+M/uyRv3kNB1lKXp3
SYtjIU23sjM2NtT+68sicSJ2k1j/cTfdNx7P27HRv8mS4WjtxYug6an4xExt
0JfQaBoQhu5c+OfDZpYmCzs/pRs+Gs/iqCU2fNE/WsLhEKbpmjkGKegRVFLc
/Cm3CPm4sr5xnIo8/474kUce9+ZdOCAcyqn/O/SVukAfKmBGzwxJwwyikw2M
oFM4qywsCJpPhix5NRkkkJlXMijARP1NQNLPS4Y5RmVGRCGEuhkYXycydxNx
zlHAf0TU3BT4zwR4HVjiBuSn8zq9renaGAds1DM1LmiPEABunQL25Bj3TY6R
m2dDbK46JvXZIdPVfloi9oiGD/C5lt6oqG2IpwFWFRwSkF0YDG/8Pso8ko/l
vIBYOdUl2dkopbP5+odtL1wQBrNKH5L18N0CEOKv8/9iOgW2C4QxvTEnvX1w
t9pzgQWR2JQpp73bEa/mfPSyjQ+bgM5a8dyu+dqL9yyQw61zfux75mGMlV4k
gm6RB3xg2MQUBDxUuEuD3NX67M3o9pK2M6A8EufyXUinBZcZzXVM3GmWoI3+
u1ITMpD8YbRVll8G3sK92X6JwXTG7g76EtatnNONH/y4VtwrIezhdORQTpni
iMHctVMelg6i9Uu2Bfe4X5Fu8Vk/mlkAwtCSV1RW281JjQXtq33wlqMq5zFM
J8t6kf3eqaPYbYdf6L4iNd1jDOHWDADGlV605yOguO/PVzbQ2y1fO5vWGkkI
/RZqubXGHO/iXxhD+ebdbpVqMD0/6zn3aXjbK8dHD5oNLNXe7XMe/zh8LbcZ
IALecTzJCDktv40t0vUHpyXuHlCq3hiZpHe0x3TLSCM01ZI6UuKG1VY2krrw
SN+dL6lx0SQxq+C8Kj2DuZatXCb/+aFaazalX5J10iCiSTaGrwISR1JLsAUp
pgAsfNIpKd6cBHhytTn1Yu4A3CI5ZBwrx9rZ1GikjHLOJU0w/BtCcIelpaYh
uep3Xt8DMyeH5dV3pb/rhaOHlk7RF9R7ic/pd1w8rDNtESwgdcyr8Ky5MhLH
T9IJ+w7YzV8xR+QfJDwRcoWhLCRVCYD3E7qgsIy1KLTkd1qm58gz4lfGgAlp
taRT6rto6NqlXllqzLgCBxdIljNwvd9pUIpijORDu/PEXBoy0f/r30EB5BaE
wvqMkv3TvH5+SFRdUP9DlVFw7a+U9c68cAJYRNiZZLZg5WBHH/c+F2Tmj2xM
d4fBvo7kc1yGYVl923TLn96jwFYpYS5s2mZ1cDADKnevxc1UE69dL1iYuslW
IDId+idDswGJ2H4/k5551oN+kqZT24NSrwo4FTX09cYDkxWNUANpUR0Mr0g6
kvU/mHpO6HLwtn2VtZcld9VPQD+WzLl6AtjNg07Zl6gMRltSoEB4Y6wFM7WF
miEhg7fm+oxc7NuwJCM/1CKlv4NZUl30leQKfw1ONOt+uh5IX74JMFaxo+lY
O3Zfwt2k8S6jRWJlUzmBgtS05btx3+/DcQEcfYqgCcpKGba8NThYUU94a5+j
pLIqQ1Je3ppAyrUIEQjDkxJrIzOSWv2dOXL030y0FTRcfOD1zppP4wsx9J4n
QD+Vy0xSE21RQJVZqBrBoxIRPAyuuj2wgqxC7UTeboLheY/JO4GoF1Hsa4zR
n+tqAJ2sYpvNoYmXQAdZhCwd6mCH8/xQZMEoCBTgBve4BZoxof+9iNaAJyOL
RTz7CtbePGGAd6lF5fVXf+AraVhAegC1VLQQ0J5mZ9Svt9MxW0Uz3Zm7PdVw
lCn7i+caP6xp0aCZ/BJe0CR8MsglZ9J6jw1hKVyRnPxyBT/mf+yjJm7mi1B/
5DgubE3n+cxxhUmzrkxRJ+J0hkzRfG3GsLw+9ggCtnii2kerw3mTfk1W+nQR
mwzFBnx/XE4L1msyhWb3Vxxo8sUqH7pBINZA+sukJ8hpXsD7eQ18xSjTSsZW
n+crXrpMafTHMx2ODT3Vb0MdWiUPWeJxlM4JBI4Mmo0h32/z9B28AIq/Kf5k
nnwodPA1j5bTgZEm7Hh1z4wKyrxGDogDFmxAQPs5RDC24i16vooP1sTU+NfR
FkJCq6iI5NFQpvJU7jVR3rNobv9mQtoaJQ+52WIJKNN55p55aquV+Kbl+fIU
FECQ37fV1NrIcZ9vprkaranyyw09XrcPXbcz9ILuDc5desNUgWg9JOsPqHj7
FuNE6ep6ui7lPONhqvI0FKjuvfuvX6SSj4KwQZjel4wFBEJ3qxFV0qBhH65L
AhwlCWmoFq+iN+A5ayFt51amHf+bguYh8hBJzZ7aEb22WxYjZd5/K/zj+xhG
upNi+QMMLb3bjO4Yjp1dr/8W5vMJgevEtuMSwDI/BUU/bWCSacyI2c7AbFOA
D6vKqoUJGv2pYdwpQT+6zgfDBhXf1trjFF0jxftKH1AawC1GKaAVGQifo/GJ
liXiMMRG+Lr65rOlwwkanaUavzWIyAgTJpRZ4TZlqh2QWngm/R+VjJBtXIgk
75GzTQQ4QltP5ZStsOftgHuWHlGOzFa8ByX8kb3ng/Yd7eRzs2qypzpj3nVE
11hD+SjwCHOomhFJ7LNTvNEODL4uLhrCBO0CpnlNq8nXa+EvLpVzRm1RJ3vv
84Ez7WsDpftFRzB0UHW6Ij4JclLFpibK7JwjOVTdBa7bW63sIne9HP3J9O6K
jGdDdWf3TAnkH4OwlyfHRq8rZIhNxbvBsvAwJcLo4WncF5jGhxJMBtOzOb0j
BsX1mQ+qtQbLQCPySMjs7kcVs3jVw9+dC6sEtfV9h0xEJVZ/Bdgin++9tQ6A
Tfv8aC1kUMw0T7V8nEKtL3ZwJrTSk5eqUHGHgm+vEJH9CCNs8Q7Sb3TC7jz6
UYf2c+rAUDMUDpMraKaMu7C2lNut5OUo5vY+D8WUav4qbpoVc8p5+dnaDqBN
PRxrCPpzd+lIEoSRIH2Vxh0SBHWjFDIvrviq+55T6TzDtg4mjp32W1Y3uHN0
hbnbrZH6i5b3bp5C1yeTZ0IKWbOsbOn2k3iRh/bqsrTDmSYT7Jd+b3N/oRAY
JNJ4RVEO6rQSrKbpizNVI9A0sqCtr8iut997MDXPlx5wrxPjJD6H79ryVTfb
/pSHgLZHUP6F6kjY3MMeiso1PVgY7S0Un67AHz/P8uHy8tnAEjKlOP56/dQo
fmFSK8dDQ3T1W7RDey6s7dvxFD4G46JJw/lNnhM354sHGk09Rcyo2YSskdXF
Xv+aUe/5X/BiIuUU4EjkBX8uCObl8zkopP8WZpTm/qWfFxmvfyhx0Qd/F9T+
YnL8gzwKVARDfur3tAXoZncZWwzZzEa4XOFgXZAvkhDi3f/2WF2jnNkcpLm+
Yml032MX++CQK7i/PuLUT8Fddz06nZz5p5Y+82lpExnAdC46akvqvqU4FhlA
7UrKicP8IPQG0yIK8ej8vlLJwYQqLNYZGS4K5trIBPo/Fl/aZG0WN1i8Rixv
fiUd2FPlYVW3eFcG92jcxBa+R98+xo4bQogB4kxnnreuzc62mG5IWbnhL0jm
8fiJA2xSHYM9M9kTkUJpsg0Kg3u9BLtXwadTrQ1sOb2pzl1ITEu87Tn2f9y3
Mim5w4OHUtEP68lO+7VKkq7Jz8uSLML+0uClB14ZDyVMwJOKNlTpBovtXlCB
w1a4AhhwLP191/xK+8wEW6bzz24MN7SGThblzS/O4K4N7GIWCagtTz0WLG7t
vwyvDdbvO/+75Wic+Fwg/gszf0R/rlPVz3xpTVOjOplDL6KIme/n+Q3Hmyna
V7bOzgFYnMFteXmUga5mu+tZA0zrLAJ7o0q0Sz0+YHNzPmT3r+PzoPjsq2B/
bhHi2effx/zfA6Gi/baAQm060StLZzO9Uzq2KDADpqqS+GDA8Q2pHezvRhks
9L32pS/rPgGnsWYtweD9Kk7vzj22VwtWgrGYpIbvKgp6KP/DiY1GYISM4wlO
2KRq8/UkWxMG6k0EUmFlViSTlFTHUQ3uhcSKPd/sNw47mpntRtcu4K1e989h
E34wsNgKY9c/D1sA7JWL8uARyO7REdw8F8oQiB44LdeioC+v527IEoLBCbXg
QOy5hsTLsM0uLBkCe0NMUtPb10h9gX99ihNZlpVUSzjDpYLIw3xNj2c1I596
swl0XG45mMls5DVMpLblQ46ERI8kM/7rpdKQpRxSMgpwcSxAylfVxqC/8W7z
6d1UiFsg48p0rmhh7maUm6jlbnTYbKKGH4WtALEdd9W9e+Sgwf/D2mV7ZsqR
CGM8chRiBTvX7aVJhgg8y4YJwayDw7ytLt45VRljZ7x0LzKp3qpRCt302Q1P
LrKHIoK6BmqqOo1uUw34uHlDUzbIH1Rklib0vfAtJ5FT592557/JzzIyrS0p
YUlTCtGJ6tk/y3yNzJeD7REgxVo8/FekjDxwxAs109OJqyezcG11zuc9NV/T
ITTmuwVYTEJVzSk6ivjg+/hQl2jjCaCxWc49g6gqw1GIi22Q5AKkqv79g2xD
KH8pxwu54M2ronWJgKOm2jVQK9F/Zs4LFIrFQ19pPdTqDxsapj81VXEnq8GF
1lDzpE3ADw2rrIpy4ob7s8KPTXXsaoYlu9Cbxwj56cA+mDZvFz9u/b70O4t0
ySN11LR+dVjWOO7r6f4BHXtKYOnVe4zjWWkCzsA5Wm0mNKN85ZxUVmTlqiD8
+Eak/AsOD/1ey8Tt/oqG4BAYwwebKqesR4Z8FbQ+DTL+OliB91jK2k+Ll1SJ
xgm2gv1GPF/LQGM3oadYouArvsTzETEv7XMh5o8ry6TyfxbhwOT1pMujkikU
YIsk4qipnLQPc9sdW5rX461QTezcG6Fe8SNokls4KfjMJZoqa86QwJDB3pZT
HdDOhHuCx/yCfz/sMSuTwZEsPdJVPweXDt39JiLV333Z5kJOaHW9BiYY21Iq
VJjBzosA98/1gVlwqV1lPN5oeXwZyFS0t5Ieh/0nLmj9OWeaPrgo6j1ujHEm
mxtHGQ9xrwsyuR2e7YPOyDhXB/SXZFQV3NLJTNe/ZnF6lZmvm7Xh3NXZsBVD
nuXupNQ8yf0y3Mqh2K0d49TUqsVoIi7AZiVnR3riZ33gUUeJWFgCsAWiiJ9x
cDm1TWvdgicROI1dof/Gb8aVvJAiYSwdYTMYRiiZfZ8hlkKFUNHMZoBOyRzS
o0rXrV/seFiZ+myTejURpKyziw5gpcf0zdP0W4nEuySgFrMYgd9AqP8G9WvT
KaoUVIzTWo+MOYh6SEKxq8PRH3g0ChlpvZvr7x+fMMbmwwt6rlSmNbjMOp9w
+XwOIBBfiCuuYqAmKxRTfekVPSMPCMQWQzYROsy7vNI6og/LjaIwG4Uq5fGM
orCzwHvHFZ5hPm/F47Ifg7buBoZ+qwUlZP9vOyDy0vCqzorseThaY//bgXXl
+ualk50hQcFn0fwdWMeU5uqMR0n8Gkpe7j9Dt36IpFhNddVopX98jqIDEzcS
78rFKsEJoAq6QgZEkpuk0FnQXzTepI3mttXTrmidGLAS6gz4Ta0fRUSt9Q2M
UinE6NUXehd1++yyZbSYS4ajOnufAbJD0IVcfoWTveM1PNK0BRTqqzBVXiXw
ReP6Gjr1C/x2wUdrazLt7zpcX8mIVH9VyhU9MjJJTVpyUZmHBhaVosgGrEfS
6sBqw9iSIyJi6rXJT5HdjPEUmPQOFai0gd8zoNFaFUwcH0bJPFcLthCFF0wf
x4vcS99tzqzq0T82ejZ3AbOVLeWvJL6dGZYFi0Oty8b8X1vV08ox5XmdpxZJ
LNMQEVfBR2EVlSuyB8d4LT09MccRsm9PvHEteGwLn14+YnQaxxpLZvXrpYsZ
sjyHBoEvF0Z44mJWxRkFbBBptqyXK68lZDu1a2tqCue7iElI+71GOzK3E1H0
oOy561uqrnNLNQxAg0166/Y0x5obB5kjEH9GSXw+dCqsWwnyR9ErvvS7obDQ
jaQ/2wTLRiEM7ARTMZgvIDx6Bi6zilj8w5N/a57LjC40cqaWTWl+Gdu3AsGJ
IoK2yrMPtDUx0l1IKoiPdze1ij5QY0wqFsB7v5YhCFjgSPQw8ICLbZpLYtk9
NJo3IkTQdaKcMZhcYV7Ton4ZWL/C1Qt/iXRqedDzyYGDdKZFzz0rjLOvBxFz
gKmXJtwemJe0yt7Ob/NRxfZIgEhCuysqtV4P2HrY89LXMdGcXzXIZMuDJZIM
RTrMrlfz57OLtXo6xshk+i8jsE+qo4URCEhTyVP46D7tYSn1YQardAjjjsjR
ocfYTqWYdHphSe3qszQ+UQ9dyT0HNbMwtJR/9eogs3xsuaP6jSztdQ6+vy+v
HY1q5OmouPl1MHsyxKUVvAbqviE+kxisr0IdRaS6MCmaG75AUb2mDgKyD8JR
Ulw77xPQX6YLJQV2gPgTwRjPCGqvfk8XeC7/vBmFMFNqLtqDoDjZ+mkZD3Tg
4IWi18RoM9om2y/q8zIVuvgO00+qrDZMhSWKgdOUhB31tmVwWmec1QkhHYqJ
dQaYy5r0BWOlu/BgnyBI/ZEZt1RptoTq95nIRJ+/yJgqAmaWFYb+og/28tcM
KC5A3u73tat1A8nxbVJ6w3Ts2YatlOyRW+pABjufvxC2w90YzmVEHvrs/1RP
7sEjX4KiorKNC/hBVHWy8SjGjkg+z7PmHLMQ7SqOK/cP+lUmfA3ZbQ7y2oIZ
XbcxXFYfhq7HAs11iZG5CV6A3bcyrRJ4H6o+GR26NE8y8U/2s9zHldsTJnsE
zh33cQ/bjE45CkMyWMPC8TwV2kCSg2TjwMzBM14ff+K4vJeTRhd7HLeUDc5x
C03KtSrG9Q0S47MyJzAyQpeUOYA6hW0oTXPtBYXawcNTHNGHPao6W6VsFPj8
prRfT2jMaSHipDc9C3xS4ByIlbu2nm948M2/xUj86gfkc2YwFPQXBFT+t1PM
N9Zdp81svK6JikzKIHFKUDpFl+6wp196uSLrMUUGcP5MG57ePJgH2SVZdb/7
0h8c4NpTEu9QL496iHz33xfFb19LFTn7Xns5QH3v8ZQ812+bhP0ilBEKW6xS
27Z8Ga1iRw4qRo1glDylrxUVaDD1g+otv4njFx38dT8/MgaoXwkLqj/1/v2p
wSK287Yrvvcn7ETM328UZH+s8pi2z6bNEzefC214TIaE8joPNfkBIB8dSCBg
PCBvwPolwlE7yNups4U1mLuWfxNBNrKUOD4FaDKzBQCNL+Wqy1lrU6RSXGv/
I/kBFCV9GDEHHe1alwYwD+DtUUyCZgHiEiYsySb4ySWpaequExzgdR4hLfNe
DyRQtIrFcHIp3UpDNaxf/O4rrK7kzeuV2yJm07Bzpo1fN8wJK8xJRvWsBlfD
DtFJThucbVRt1kU0XXMUSOaqdd5bqIq71eSt99uswjKhymbejp/40Jau5fkE
DmdWe3ohair82WuGS5A6oOZEAlezO7eIsmCYQ8Xta053QNZRhvvhOOv+Rwgb
cI3QDdKjOO5wbOMQOFfh0x0lT9E0Krlu1+osRI5qhxyiEI+XWM/MFstKIXUk
SVpBE97yXE71ip3ZKdw6TzMvfTLAOa0pXhWv0FSQXdiLtTD7Vt5omp4fVVex
AumEwLd9GJMGPBJtdUhZYk4s59M8eSvUpBz8aE/rKXRflvbTRb8REe6wZZ7w
rSKFYL/dO+U53ow5RHPcGqyzShXrSdfzzY9nLIoNe+ipwY2sGI2aLX1Vcv3d
3OaE/AcM6AG61Re5tyncQVMfjhsZODyZW+JxZBwjjfOSp/wIXfK5Coc517gy
efw4ZRfOqYXIBWpOTyarm6XD2lex251Dc8mwjpTmHO6dffN2i0G1lSF6q6Z3
H/MeTDiaZ2ohbtjzxT6dopI1nvChz5ncqx4IoWs9s1yaqZtl0piSP0dkelBR
4FVv8D74G06+C9VgpMEgXWih2qVK9foiPoitD7Sgd7dKU+GL22+ynxOs0Xil
l8xybjyi6lSy+XcmtoqvReGR+3WE8CIIa3GqCkaEO6r2GM/HM0XjdfgzY6Rl
6HeUUYtYE40JRjVk9CPjzvP7CAcexlXKJHS56OUoGI6TIREqZEJR8AEripJY
9ixg3mchFZjs41AfYfdXJIlhECOANV0nlbyNlFiR1057tvNPPRkiOWUYXdoB
MZdN/LFs/E0ZUiNdNkjqOQ8iqwaULFb+8kD9JE1XAr6LBdllTEQSQ58Mw8nL
OPpfCQEkn9uGQoxP5Cnq+jAwYMA5jztZ+97akSa1wtwpPQHq3Muw8DWX86eT
acQEcO83ByZZTKbIHTBda0ahihzofjeU9hp/EKZkEzB8mgojBvBi1eYrKzZR
fxPI571L8OKSIrrvFiTcQdCk2W07qiMzpS5oBR3bRe5rrze1LPf4cMEMiqPA
2N+QQlBp0KgTCJmHgVZSzbKFBK5ks4qMMpJd4cx/OcdaGu0encU4EnuiU+EX
++uo1F6QphRxrECE+naGFsx8zogxwCn6uro6H1dSEZHqSSAE4m83gLtMC87h
pzr0oS6qa2rA+U0U0yFoGp+//8cqmHw/ZLYmL9Nk+UD5ckLoE3uYOCKaf18v
e7f/JJ88IDX7Yn/z+sinwtQsGnKFZwO4Gkg7Z+QtqNKrYt8BEtEht14lU4v0
PrYi2I6YxoNX6B9EC3l5FnY4F2N/ceAfzOw2aiAN3zxVmF/2DQlvyEIrluCd
XlklKn/l3+IS+8hR9vhKYB6hlmfmL+0NiVpxq2Rxj4ie1q0f8XsduEjHOZEc
V3V1uE4aRSEDYKcCceY/mxWvQC9dkCcU/jNTaLWjJ4v7XddKmAq/NCT9BK36
zbiJPCEsQfwMsNKxAgCaAjm5kPB6HKJf9g1w3c3n1E/QbdtlUsynbLQ49wi7
MQxaOKojT7X/2hVMpbQyoBIz00vLF8OsYBXPSpFYDMOoaiavU1Utsfp+JJeW
pJs0LH0BjbYhV/BTjegqAIzC8VRUHsYnbkTw6Zvm1s2sCiIHDIGcnPfTThVW
zllxL+DnGVM48NjsoWNByznvUtteAKBm+tUzLPcujn87XM0o2THgHg2ULH+l
o1RBkHwhoPxmFi7WKT2mtXPoPXFSPA2Vk+6HBpfVPi7On6wZwQiKixRvBzEC
oNGP4x+TVyvXTQfSoUBHNnMGEPkIR5nwUaf5pjX+g8x3j/QNjbWVrMS2eyX3
AqHihOsNT2McBqoYw+bCe0Lx2M/i78x00aT2WBee1V0pp+jFaaK8NzYEflmy
NC8iFemPa0BkF+V++kn9UJ4+emVBFCn/Eg8xdgHIVIKVUWjd7u5MZWlQrdaQ
N/IjHmpWhaeboJhihw4a8AqyQizpyiOH96Yu7OBE9dxeCCHR2J6OUZfg0HQ/
FUETaxZHTXBw0QuVROmjQsTBfOssP/3byChTW8V+iekRg/MHMf5J/Fp19PWc
89ZxPhHqlFfAEE5OINig0RAeNYiO+M3zEsi0mOb0Iae/4Uu/ShUoIcFekUJC
Q4IN425UquPGB7XaPehNqxJT5wfrAEb2srNu5tW0Wdnd8f4dkrjW57LKuQn9
UwiMTCLeHDFwM3pryUUUwXuJ2gOZRYSF42/AlllOybqk+qdGO50E9OKDS0r8
12MfHTmusMvRlBaa1hwrbFYNoLTvx3IKIvL0tmrp18pjG/9avSyecNPXMege
cqL1wYOgoud54dg98Ys2JAEtPkJdKCGqBDw1xfDnTS0XWgLIXgkbMrNqOtCJ
9FdoD20li2Ki5xuCVtfwttnVi0GAGtKm8emIukjTai1ZB0CBzS8GsKnwsVib
kFZRfFbZ7LX1sgGlDqHiJQV+iUBcUhzXLcoeXgwRfjFV/jmMXaO3rW1V3apQ
vFS7fpieqXXHvO4Mcem9unwcx9V7IK2uoG2JczNIV1iEiwZ2Z9XViH+j3j0y
3XPp2BTcK6zLZkuQCPY6GQgCzEu1eIH/ocU7+GuP5+WtgE35wryUWpOKwcU1
6eCsBG5LM8BE1ndgceEgApUdPIVN7zGHSNytGFUMOGYPtnWIrnZDyQuvgCxm
q4PnHDieWTf1/ZPnXjV4klAi98nfAeESqlGd5JQAWZJvuMydPn6SbbMEoW7R
CaUchDeZc1hHTNE/HP5ThTvPkLM2gtaTdnciOa9FPeqCx3RNXe0EpNH9Y02f
ygObNIidVW8D2ueB8fo3XreV5pSbEpgI+uqJCtp9aPzS7HUGs4lVz65ZOqLE
srcXPD13QC8nTD1m6NfQ+WPvAGHMY+qVkjaSwA8NbKrACHbNvK9zFAyb3wyr
cJIXhwecOKX21/AH+l0CAJGBoiJZHJPEI9VVYHjnoz7Sp+hWZZRcWs5zqyaE
zoupTFwC2IMERocLgWQayAkWtm1NBCWR7emWfFfV+eqdztr7dU+iAtokpfLc
1cBwaMAENqtEouGO7rO8nmW23M03orRBTMUgPUPhyQ7B33CspwNqTTdGtL7Z
Fr7vaFksoMxAp10CdmeGLo7xfuUqwLRBwu2qKsuLxvtyCYwjhF9G+2lAPqJT
LJQl8hjsWs5sgQEjb/Wn0DTGIIQvKcH7UEPd5iD1gZv4vRu9SAiL4r3GZJpm
zJtZtm2iElKUe8AzxIgq0zWGAzl+QPDiSlsbjqVwd1L1JGMzAlBCEZXvdy26
Sp+T9cvsEZkXf3kZ1kwJCBbki/B29yU1krsIRXtKaA0hWuWujzNT4l3zhwY9
kufr5EPlE+7BV6Uipz8B1s4+QGXzeAIGSKWP2kuJcwiMsflZ/ez11VyDHS1Y
QdB6C6hKfK50APJ01Fk6B/+cB3EIQg+fKMlH5OHGd/ZouV+3lhKcyfqnkupe
Yt/h6ivjMAYl3W5j+ahaZxWN+q6nXxHDP0Bj2f2YkW4d791ZsU1nENsF5CAe
bVj6oE6TGw4z646JmRq+uZf2bgGZKOAwZ6WQipHuRpCJ7EfTOmAdE78u77WM
2HVcZMnVHsxjx3CwRZeqkYlrcDyUeoCR+VGfVZ5EvGVQA7kpywdqeIVPWj2x
2bjigfRmEquCIcWo6SSjtNP5LJKXiA0VaVVaQctvWVfF3uzqi0peTBP4Iaul
oS9uCFJ760JQKBLwpUxzh/AHUllZ0aAXZ2APb6IwxWYbqE5x9/m67hynbaR+
FV5QykeaJWVsNKsbpUO58S+PHiS3QowgSrGrbJ5W6KWw7JMGd3f8hOCS8NRK
XtLUffwFKlpH8EAtNmLY77SAt6LpegIjgZjfDOFji07ySr0KTIk+aDqAjufK
G/CY8DEVjXqPnb40AvSbaIYv65w905SFjE/ZTENOnf0GSpWk+Vx+HVoslke0
NpOwfTLeoxEUS9uHdF2aoDwBSNb6mt34qu6uN99jlSB/Z/BFZFuFwI37pSLt
Xm61YQYRaXpcFmBIL4MLLJ/IimFrsDjUN7Tg9B8a3DxCETS265fifUeLACLb
sNbbd6ltYuZ2gJe810C20Wpq7X4bWMPc0JD6zy4P1jfjOiDYLOEbMmMDV86v
lEuNFFSZl/urdXQTrVHEyCYpkaI0p5XBtg2PIUBajnw25alYjiyfWtExmARg
MG3UMsgBwHaI7ljB8S9clSqWdBuswI/IIlST6sL1jW/+UH+yBX0l0+mRFFmn
INfO0FmuGsYlMHulgmSmf4WT52r9wbK82zPt08x9+ML+ZGMauVp27fB4wXRU
0WQAzvFsbtE6sfbtcLWPPj2Ii+3UD+MSd5aovpqk6whXBSqsu2IpyeXm7ya0
p6Y2Q1kTLOjqgP6RRoZo5w8dxthtVFjIwHVlZY2t+DQw/8vr0zNVr+l/yj7p
sIlvrLWxMgnq+7uNA/VWioDgJ1QSGBdrswVdfAFfhk70//Kft8mN1zKEB+/H
uPt821hsybIDOzFz7WHDnQ38zR3xdcfBo4ci6khgiJEfSvGlwcYj+/0PLJFw
jgmbJeN1ebIJRo961Ca2YObHklxnM63DpH7ZC2jSFBIWKGudwzCXb0VH/D1H
TrC6i1Pxsj7ZANDNhuafSE/PC4X3z2SzfKGOCpbfRF9NdgyfZiCQfbyAumlJ
YN8TD+Wczz1p/SR46S22N2HHVitO6ymhv0CoydblzsVtvlYJYeKD4Q3hESBk
0MuT7nyZxVN+1HdFYyBoPspWE5Q1UBGKMaMjiBlRN9FDEoPzb1m7e8UGEYwo
glc/KEqyjBD56826/ed0R9jb/zpYvyhZ4UtpNb79ywvxPHQU6QUyl3BSsQE1
2cn+Gl6Ad2Al5y1i7i47F/8aIuJzJ/4TzMWkZQ18/hEkwdBan6oT9bd9Sqjl
eLwmanL8ge1Z2LB7hRU04b6/6Fg2Mozv+f7bZb97/oPzY0QPwI3s0Tp8qwZ9
VCWcQK4nsN3/6H7WZW8wSHKoO4h3TxXSBQso9ED7kN9ore3UVqgObIsT5onA
oZSNnD6dGbtfbv6uFD6qYr3/xdchVzKPUUgVhiY5w+lJCA2bGDnPw2/+xszt
Y2jHiKkIXDQVqgNysNl6A/M6Ih9NQtMsXsx/viw+yBMs0Fjy34CCiKC9EL9D
9doOj4j6vF8V3BX0UvBIPahL8nrnm3XXMiEc6QM4SIZYWCI4+zOCyX7bsKCa
SxxS5qetqyoB1xCS6faBNUz3daIxB005YhN8G9m8Y47Gs54DjLggvKDUa4d+
TvRuspeQE8PmvfO9T85fP1MQ3aWniSzbbBJSmq1f6um2aKW3HzLsE++zM6fI
rhDUlzLtErkRe3N6xv5NowTq3sL2YRWt8OrHQFTjqw1erDHN9Gnyo/jR7/kp
Mr8LvTlLvB69Mm/eIdNJ6o6oVhhMpVM6R8Y8fXgrSt2iTOU0jSSYPBGRTESR
XhTSZ1GZi4R1Wbwj0goABIAGrAHyGOo/2rg8xo6geXkQmM0VJXl3ASIe/vqD
crTwLWod+Wep3n0bMOl4wosNwuvRQjcN5jwWQgHR9J7MP70fUXyC6w7CnuWJ
dF69uQd+uIepmVZQj4fVxyVI+DCjGZ7UBRg7wWP8E1IEdAulqkpwQNVa109h
jbHdy1nGHC41SKBpjnnQaWbK8V+rl37vUZ3tGh7j6mwcCqKTee+Z4371tQ0J
amTTKP2jmxt6iIQDEY3XzQbrTXyGmMaVZ2HPRms49TZjNQlhbUnPYKlmk3wZ
wxY8MLeWvt9r2brxQ8IveoonGxSb6//99qh0S6WqTZDz4J3hK1wdnJhyQJML
2BfHAhsKxaKN/LOdi9r6eBeGFD5hiXZGJwFsNuX1Eem1f5j1Yd9N/TQG6wTB
2D+y2xi1h/iq7f5wbUD1ggwsFIklikKFY48Pvc7i171MJGKhf/9CuYqSmVOf
e3FVAHGLTV9lNJo05kB1IZiIzr4Y36+GMxpOevzQeDUeMowVyXrXKeQw1Zky
BzttQi0b1gjMJtyvQV5vSpQ1J4krVxNLon3uGMk+smN+WPXy9r5hgud8eevR
ukUIRkcbFTf+2TNnwyolWfSwcJS4GEITXyojb9M/DO2h4Y6xyMnREqltr/Ai
ZF7lvmSGuAzlt93O/Uvff8woVTU75z1mSuYHDjVMjk/bgGBkzik5QoC4NEqL
5VZlEeQKlmRcbc0mnhBryDmETfW8iNkRGRTpAomGtsHJ3YI/sNkvT/FZL3ZY
6Xw/KPh2Din2F9ZhgXFJfLcV8xTKzu47ZkWhXhzZEpYcaGd+aybKkctNCHed
8DdeeqKZFi84rCvlNhobxsKomLmwVB+IRF84Q4DYFKhV+6dGjxbE5EDCMuvq
GC+yNQ2k+74ctY0IT4tmnKOvkRPjRViBp5Pv8v6Pkc0Dt2WuPXYej6246ZN2
qnE4ZFcATdiVf/gGs7iN6lUBMj7v64eGAw57pq54GXwzqcblbpB4XeuxMPze
Na86VCGFeXoyfIdyPEf3s7FKU+htWBiK9vpco7AH9/aUCgtxztXQbmKdG2fl
i45O5PSujXZo80Y012ZM4cPTlB6H33q+y4HQzA13vZRLXVErjfgAs5KsQopH
AJXg5moocSN64P6/WTL88gI7eUKJ0HjLsEgjlpR2thiUwn77VJUTYyA4KHOn
xHE6kulfKv7rBfneY//4557y/Uzu1kugjcsJfi8Mg8+9H4Fe8gfPdidfKJ1O
1SB5vEF1KAaJdopUNfP30gJv7s5Exx3McU6mCpV65iQs3uqPUn1uWc2w5Qh7
c3Vu8ru4UqaC89aC9dpI7NMmEilE8gYcVVWn/vkRykP1RngAIN78OsZg0Acs
xcMouMkhg3PD8+o1TCB3XowQGlWPGHVCI/dZNMSnTYRcXKN3++B/R/qxZMnd
FSdYP1e8crndYeb8xOG9HTxV6OLB+9GQ0RpfupH4yH6HvUu5Ap6KnbZTqE7b
ARfjwHQakLjbMi4ZzPymLgLcxKIoS10OwvF0/fwPnXNr7eOKnqGVkX/67+V4
vSgdFSypSxjj3F0NEM4H7H5z47N8iMkYkYoq7NKCzlwJ1NwXc0Ktqgcj12KE
avMj4N/6mc8hivp7DTd5qtFtMi529JNWeNUOSAJu56jfVt3nJV3sHPJJg9L5
2B+diM1dBJVEtGZMPgoDfEw6v4eqO663hfdyTrE7nn+WuGXcAhr0ID2dwrl0
4MZmbSpKSDS82X2bU0bcxUeCb7J+hIkBI8Y66hgth9kGuOB2Hta+Kz1uVtfT
BLqU1JGirHx1qz1UCHArw32ZrhhBk/h7lEQyXoTlkP3B7DPYvrMAigl0pj0Y
LBfDdaC5Gl5K7h4W6FkSHMxi4xKRhM/fGtIIopXvsTq6KSL+lTjtkoiySsfx
NCJw95EVA2KPj59uzJx69HVTx4U710ZC2mivCFH6dQOs2tJf69r3koNLjhCA
EM8LNk4L3hEFqkk3Sya2+74CFmfBj6wW7Spo7Uvq/SlnuHGUqw7vT+07eDSv
gkcerB7RaZTMvP89FJ9HeXjxLrvpT7sSq4SKc0Zdr2JRnBVdofD8GMR7gYNs
rf3LOUAeVbLezGFUKvhWUKoE34LNntprbcZEzdh54cZOnIluwqaznN3x2z9O
DciBIL1gQBhVAQxYLvZiR8O7vv8zEv2HUUDlHW4yz3SaBShvt5QygQbeZwrc
0VY2btFZi8x9LIMvDLoQPi2MAz3SryzcFDJ7GuYYRIpZpIA05hojwHiwbujl
cSP24m+Fkoqzf0/wxWC/wKczAdiXHiLzDgS4mIkEgOVMX1AEcGv/B3l4yPju
i2Q5PiINnqRKlDlQCWJquaU2F4uAvKKaM+TLy/PQ1gKYf56bOAcS9n1wqOU+
W2i006vf/vXnb3pdHTJY6eiO5odx77283HdQqxbAGD4iWG2ji2i9KMkALXBK
+hED3kN2+/RAeAzpmSAun5DayiPevfx44R3jj1lLPUQr0x6K0Y2Fw6b41kB2
2xGnUCBrxEDfy3YASkdC3A2qnFwpTtdOZObzQDlc5Z5LfYV6ZEe3BEB4H0R7
t0uAwofcWzErcc0X1hp9yPUfZ94cSR58z7k1ctb9wLQZpO7lRh7FZIuW1A3B
ItWaTpr0FYZJokod+U5hfu9wmBkgwC+F9NkQeYkeg59pyK0GKSxVHVE5imOH
1A1WxE7CsfskWr4PpYigVysjtmb5lbRQlJqPm8sID51ovsruj/kKfd22qF1C
BE/qYoGmxneGWm1Ba5KHp7IPcPD/b5tUch21g1M4+21nd/tx+DDDanN1DZJv
WiFUJrqrf3BS1qUcW8TojusfCRR0g+wQRW+nN58rJnDBKSt5bdwwuc9eDQNB
Sj3MpA6MHw4rtcqESYoxncuMB+V7Viog5z7Pp4Bjz5/LS+bWJxPmODsnsdLm
jGrFMDf7eh9zzfx+E5iVBUoYW0JvvDooMVi3clr0vFBhMkNJyUgNuRjvtnqB
Qk8gGfJObFXKuUE/X3xhsy+4eAUTRXHi1AqdmuXUXP3O6FYPgwGk/Z8G+jlu
EtG5qckNXmesBS0zAvyRWmdjYdpSMeigSq393BZ+OY5l/GL0O2CrpQPNGp1b
AbvJ58vO8emMhfwkeEMu+7tKAWD6yAH4siv75QmBEHDAlq41ih2kVpo8w1xc
YVJeyDO5Ha7MS27BHCWL0cBCuOZkNPvGI1FxfizgpzMyH8vPv9d8yaO0ul8k
sWIijwPxTxRu6Ul881M3N7DYdNs9c+Fn2qyDQlv74n889YEqkliod0Fyrk+B
gquRw6TEtsJutGg6QjDF2xvdPKJOdRQeCIJz1/HmODl+9idvsW9F/oAEPc6K
fboptd9j8iSlLwdJ+aKQcREC1dljta0aobHWSdJjl5gPN+8XX4AonTFQ5K+z
jACxt9HdQZtMzaQWlS8UIjJjzRY7pzVGyY82ZyIUqGNpUX+ESOG1AIOxUcxT
KrVXGKDk9vOC0AMOl30toekpJw3GCR1AlraKxDIv3Bm6fceVvZPyj7VvKC3N
zdCh9fLz1y/mZKdGEaMdHk3uYYpYyi4mfg3Sd+FCT0D2Lk1483kcJmzf9Gf9
g9yXektiojBOHU1c5SOTlmBWc3ZlmAfjQ+0kIKJJLxifRuQBjAIKGanxJh6c
Jxkw6NfBx0a4npvnQOddqnuIo8NO5cNZQlILgEJMEcIwzPeLz4wWN4F1WDWJ
kBMGt3Euv1uJgTvjfoBAjHxPmQBUYRmO4txsSBvXBf8mIsngXHkcpCj+DzVz
Lty6AFv5/vZNpaEsOZuEJog138ZnCtvx40j6MJUyXV+zcCt4Up8lxaQH/EoY
DFxwM8Y3V3VJMZHbMAeXNKJlcoDkEGFsR+16MtFWh4gp0DvikCudlPzgz2Yq
k/n9+Y3T3xV+Gf4rYY6fYqyyf9vg2hBsdA0z9IaKyxQJnkEs+l45BneHIQNV
woR30LiJ1DOV33G9r0MQ5vZKPODiHFsrt19n+JrKRTs4KiCHbpQD1NiSkfBC
/M7KvVqLB8BNZj6LUFDUVoKcMWiJS7gMQUQ6dTs/ybsxfSp8vcyY9wtWxhuE
5LwHpazhre7MfW21cQBNsrSajKA/vYhtKsG2IPWUzQKr6jfrWVixyTt6zxj9
Taa5h1ZCqghtEas5AZofiZQOCgkOk2iMLI712bp9jd6Bky1g3+eo+1rztk1z
w/es2Qy6pEzr4hEmRVlCFdHF0R1EosQ4yUvMAk3aghaglfzFPXE5sB8Kptpy
urpPRSpldQ3B9Oe3MToF1KV90NUmW9iLwR4xR3Ter3xZsE6TK6Fi5HOJa4o2
r8/ygkZUUmNqeGc9T0qq17u723JYaGWINNFaxYycSvLYoWgb+EH4sPEaYYrN
BDSoaOTUK9xFJixbj3nchxh/dVGwg8pRai1tFLUnXmRNm+OAN7Ul1EqcHiyN
wUe6SiPjwb3HaE75t8ciKIH5Yx33+qnwBOgWlu+K94K5dpcILG1jt82BJBn0
nfmecFQAhXxif+9f8HRJX8mlp/tDfDG8O7n7MPMnKYQi33u6TpS8/61nTaxd
3qjd57y9i9239uqjyU+WR9kyJqQid5SzNrS609vmT20sqhVBo7tc9ZTGk1z1
TUPmtv3GNckJsoymulTMLRzc5Uh1KwoyBg+pX5jsJm1ThNh58U0rFVWjfCi4
uY/Bay11MiVuSg/FxvtiN0VO3gEAQTltLMOPx+MDkg7N0FoRXMtySoBsezJw
Q/sOdqzih+didxb7/Z2sElmvljDv3+3SZzSorrny0vipbh/NByQD7KPF6j1C
6uzdfl8VuNjkToilAAaCGsuPG6SCCI8Eb7bXrRHTJL/aThyRiOQKg57URYBD
gNIUOlp5M3wwnnj2dDGMZ7D8xdI5WK8J7go0OxlsCyFnk2SXFfHwgbRSuHno
tJ40PMPvCL5/Jun4GuzxiCUO2mODGiKFHGULENwh3h3xj09bd8CmOO8xZqv6
wRKs16Ztg5142fhAi3DZP/TE0vv5kMnNv16C9AWANlaLczD7LBmh32o5D6Xl
+SqITuTbqEd5cj4BV3yUDh928nEHBZagi4fp1/j7y1kuNH0uuJ1yDsATPh9X
SrJLIMEr1XBwrxOBqwWnV00pC4F44MnOQca12Mw9EVQIpICpp/4m0ukzfPsO
x19Pso1tZPYzrWKl7SPr3voO6EWpN8bI2/vgCXfqiE7utktoBIsnVC71aKyg
EZuh/fmY+hi6kB8NZh1ZpWgzqP6AeU1liIUyGhJWGzkQmygFv9JpeLFQ24Qa
ILlwSW9DVmwyC4va9XL3ZUjkrvHJHwI0+kD6SJ/FPbq2+S7QnRkgI/tHC+9p
KKz9OpbJ20V4I7mmUmPEAliBNpQmtrkTt40ccFZYYHct2YDeer5rahogX3SB
PsB0WuMOg4bIK+rdP2RxkdtUaHpznaPWJ7ckBqTDi4nG6yIlgYi40sdzsXd1
V7MANWJ6Pt2hgflDFf2vZjjkpNppiCgTu5qskalLm1xWslLIQf7vZMiEIBR2
u/BgNWAJv38JmScjVnb2Hw6cW0KyEOEx4Lz+rzLHWhwFDN+ZNLSloBOXKdo3
96Fk6jVVLXq2kteWmgvu1hYwtGWlqrhG3zBePdebXEEIGx/L5NoCShKbm3B7
2l3w2AF87MzerE6XcBBDSnVrzSAJCxfO1y9bwNRLjWViA4QH3Lu01e6tKbIz
egfjyetQAgTz099nwh1YhRPTVC7gznoaPsqwmZhofMxmov2MS+YPEkVvc9Zg
PcMuJJ1LIzUREnqqBIwqxI1WH62Cym2I4bClx/x6rbFv0R1X8/f91Mx+nMGK
peiRifh7R5j+eNxc7BUYCB1njhWorW5yeIW49vohY3ayJaRySgzCslKjJwjU
AgMA/AbTVauS9cP6bsv5AOIoXbOtyrfoorz/rSLXYM0yhV7QtlgMCaKDyHB5
uGhAyFEikUPsrz1435DQgPDCcx5e1k8Gh6Da/GAej6kcpim4DBRUGA6hyISH
nMPEVFGkDA7F/LNTTFYTddRERIFqDQgqs3pnBs3j9PQk1beCWnrtVQJdaooP
e8uvMWvWLqABgDtNJLUXsWIRVM9BiEEtTAu2ZcNbIKNwB+83dbuDMduwzgn4
fLdQ5Qs2zLVNYSSZQ4IGi9SFJhwyg7WjIX9d0PtRftD/neyr1kn9ufrXquBD
9quckM4MmMVGXdbP1c77C0mfjHTvhm9fip41Kk3YADgC/Iy6ogHYqV6Ciz9G
qoBJjwb4uodQjl6Ipc8Z9kTl0fxafeAJdiqkhfzxKFatzp3sew7ZhJLFW/mt
iNdSSCjDUCsSXpv5g0iOZ76jKcsaOhzvvkTJAefkw363rXJPvRpd59qksiye
yHOfwLPVkrC4ZaaSOIuWc1i8PJmP6efEl3Vjg3/vZ2BmsedLWZ2YhAYzpSSe
Gji0BSPwlrl5qtzhsJlNVeC5n8SxWeI7E6j4DdR3BGUA0Ng8lkJgyg51xWPJ
JYJvuRka9lH45Yt8ktCUblquS/pW871GRfT5c5JXXccmqnN4ZaZFQ5pDrc51
rk0a54Uf2GYkllphglHtFyCK+LXSMJr71nbFHsm4tg0vvF2RJu+9Ko00rrGD
zFYdq+HUWDbXV5CKXtva6xPxZHufduSuJbJNfFymvOT0BQhOeHC538Pi+L/2
7DiQ3iTXzxaSth/1UTjXAambVgWkqjsQLoRLb6rhk/cA7DHjcIZK9DsOpaU0
1IpJR3Vhq/jI6oZfAYWBaDfjExLZQowAVurHcsOdxNC+4Q//x724X+0xqLm7
Z6EjP66OCAFkn0EFeHPYayQR35xB5LmYKd28DBiI+FcfRDDntKqRcsR2gHZL
hHuiS0TpuL7PJCwl0A6ezEu30ZrsZ00OlnA4c+DwdisnN2Y6mNoTOzdqk8/l
k6TbNsC0clAckmryX63dNMMgM+7/Ui/9jcygnb0VeMzr7hz0J6bJ2T/qmxjy
kzGu0miWPE9qRJbWF1NHynl4UYoicDWC1piE72KmA+2upTQmQ6wGMPCDK5Q4
4zzY17AhB3H0eh8zODuwSzhowurecpMjSsEV2gDM6mt7vzDiwmF2bfDAON1i
rqtyNrPrY57SmcitvRC+BuPtAc+QdUwFLrL/58aY89A05T+JtPekEJnHl7Ad
/5g1YK07JtJWbMEL11n5JeuDB/PJTFKPIdEmaGfI68rdfi1O1p1+bRwxMmTM
BIAnK09uTSrm7oR1ypNHdkVIbXrCoYMD07pARdOwaxQErkDbCfacDz5RK7p2
IHJjo8T19mTrO1/1eEEAOb8ONqLujngA3Osf3f5PX2YHf4tj4WRLHLc/I8xQ
yqlade1/evxO+9sQQfboNu4LTpu40f69LJERQ3250Ni+lj9ILDTHWpdr6h52
u0cQLkh34G7Cy0MWjhzn8ffcsMT8FvjWrxKHbfEhCccqZULKkD0hhidB8naR
a41AjAU3yfI2q6Epzq3ca7Q+K2OWHypj72Ze9j4RsyNEYbWq8Vqb2Xz9y+qj
pyEiK4vlNigJ9uWqQ4KRdWrlcNA9j3s2KSfnVa6I1MXxWvL9nG8ltMqQ0JJ6
fZLwDut93am5OVtE0krt0mBlDOJwhQ1Yk8NHjFl01u1vAH/q7vQu/4PT6G4Q
26NpbxSz0J/9hKlmyy7+1fM6Ale8jJIpV0ZIMn9LuAUGdBS0PwmGtmimVB/1
XrRavYi8EOjx9MUjxV47llJ9Up1VjsfWjUQqNSAKKknVGe1qhYFawpljWV2r
EIhFpfRYQGC9SZkvc8x6gMS2aRmF73gDokdFeJa1uZ30YMxNP/VceSVCrFHI
1+FC1EjnGQPHpqTy/hUWkiDvWgQGo1O8V9epsiOnfbZDFHtQmgvSR0bVBbdu
ULPuEBfoeM70xPH1QGpK0jmyT2qdp90+40x0skDyWH4V3tmCKAg2A3eIHADL
IOykUUQMzJw4Ey7x/tqRLUrwGbtZcU8yWhNSBw48CnSeqFcwJjr21kwLVsqR
bLHI5CExPursY135v/C5DA/c6EGMwP26a+N86a9Hu5b7OrrgZhd2SaqOQUJF
tYEyPIG5ZnOCNn6OtJ3eqwEfi/icVUtIYZSGaZpavb0QwbCAM5syhk0y/Laf
loR9HFwFKyDfo2jiUBVEsMUXnzCJYc8UnrCACsKZVUbT4XHug/mr51Un+q84
v+/QkiatNa/N0Nbfn8LteO1Fk4UoMYwwF7NjTY1qvFkyKyvbynzdIjpYgFW+
tyYV3kXWFi14IyR9UNhPXxRb2/3/CvXxldweqbx9OI71OlkVXaM5liiBgxi6
aEg6MySYUwI8LP8jmr2ZpvnEHraMRl5WQCA1bKSUUm5unII9mP5JidTeiZm3
9yZuXATTkwKCf3AIuZmmnweu36LEg9mAdlZzoKqYW74ZOHtM6KvxkT8ifEOj
LwLkDlwm8T5WU1NcnX2Hsohq5qWj8VefgYdQTFulTfJGgpsPCszMK6C+kiOd
DJQFTiMikMHa8DRHrJ4iMAYl5zQcZDjdchwJy2MfPWeWr682CyxCW+pI3t7B
hjpQz8UK3Rvn/tGxDfoZ6k8R4EnrZ38tPK24Z9d1VPxSyc3Twzqsm5Ck50zi
TX9xLes2emcpUK7Q9gua7XmcqELJjywaD4UOKP+WdmBvpbrUBKOUnl5K2dWX
YMx+WlSomNM9d5nc1ioPNfiVVIWI0cRQvhyNt8tdZYT0wHWlCqH87e8gelPe
Aqpin3KQbyPT6XiFKYyL9jdmRWivL6zLwrk1atNoWgGTuF1G8laQjO4nRVY2
nutrzlzeEEo3JHl0dD8rXKblcBDt47VWuhsZAMHiLWjORm/z1OWxvoYHOtfa
2cTX+8sXuMotqwznm2TVBxv0Maelvt6+5vkB40hahutHpIrAETTdZTOYyMv1
qTM9pNkF3ugJ9C0ydsw1mGWNn2bhy/rdT021DhxfWdGjlt+okDRBIx2iR++4
kXonY++p+PKIoTgDHsBONgZwcl/mlU8ljzuCkCOr0v8vZQ/G/9re3kuaHHQ9
LHah8XkvryZHYPPfmJoOTZudGNTOCgoI+GHi6AJgOyTeLgKFsQcgyJawVjUs
I095cLtpLCotcRWsi3yVLci+Y9DwkpdHZPuRPR+MCkdgAC/HwtbF/777niV1
ge212klFpxntRRfwTnIUnmCpDLPxDq6NPz5IbWT0uSwFRNpdtiOBIBLfe3Pt
FB88id7t7M2BFfhzzi6ei0ly0y4lxYpITqoRdQ0sI1VtD0Xlh98CCbYd4d0/
ObDIYhRAai1FcLO2g0AJho4UEIkL6Ff0wxgOvjsqSCCzMVhNk4bWPSUJW16X
X9cdofBlaVIl+XUG5lfQ5JIplcqaxxNvgP4jQMpgQfh0e1p479SatNcMfWxS
YXZfNrl2PZLXS6p4I4+E6Yh3vngJGZw9EHV9oCnh7tMdK7cYHkULTr0SSkx8
h7WyBYnXI76HJ61SV5nnJtQQ0XAOldTAcgNVceFy8XobZTA2DMXvDc4Xuq2+
ppNHZYT+/IxlbDFI+5FRBzVuI9vp4vpf7mp/ULW97Ui8vG8AUfypBIxjiNp+
GqHhwnA6UeptcbS7hV5+QEZM3ve9Hggns81xgesmXiMvuVm0nAXDi1GH4e8k
Gux5UbQ+Yk81/LUhv3SxbC+zOB7AUK4tpMiUMlIA0buyCeyYycsbcTQ7waPn
ifbzOEDNswMPAg17OsWBVoWwPBEWEyapv0IDee/qsibwltnDi2UjzTMyvooB
K44BpfO3+6oBnOryppW4FPpZ/bN5cTJ9yKFzyyewGGk3Zuurq+0advgDXTxE
MWM1ZG/f9UzYvwBPJXW3f/AVCYr7FwP3NK3JwJRjZd+tZE4pNlGurGMWftu8
coZO/Q1YgH1Y2Mg7WxRMw+CS4Vc2cjDSWyqtoz/3oWqIW5gzvgeccatm7odh
0a80RVGPDuVjdqTTzVaIxt7nLfR72hDbhLWROCup4htlciUMpV14BI4sbTq/
QTSHGryGh94dLdYrOfV/1KG/+EuMwql3kBwDQCkY0jE1/1x0gGEV1ZI/vOC1
p+vD+gG8pR02z3R7F0lB3yo/Gtti7hSdqNYfLCs0b4ST/YZ/osN6bpiLGYch
W70/kzUtqi+rE7hom+P+Ik1e2zxCUKFot5DOAd8zi0DsbRVY8jBh6/rGKq0g
JuHVuWN5dtHc5LRdGh3b0ByiJIU912f5phyIv/2ltoYjQrgZg4B2hBCkCr6Y
QY2reZpi4ZjRP1ZLlPQtmRWDcN0EIy6fvFvl2KSi9jmjKr9vI/i8Df/Ku2Th
vYEVOyOj/wNpkXanhb+zw6PLsBz6cKK/lg3FS7TUq+3vcfu7+7JGBJ0Zm11n
EYbwnoq8xyuxkkEoKBjgEleQwMp3vh92zxqs3gID3XcEvGklqsO+9TU+gUke
WmKuKxs9/KUJ2E3IlZeG7t4JPbD6a9exrgj0xKssQi0PTo2L6XGb9qc/5j3Q
3/Z85oYj55GrNcG7Sdud5FXjpokkzCHp3fm/ALNySdt6odeUNkZl5FZZdZhx
VoS/eFDiaGHPKsHF4xuTYPLvzIWki8twuGKrr8Dz8yu8zG1VJFAX1x6CISdp
6Bh6bxCH1UHpmnJ4cfHgo8QpaPZ5TLgwdt3pBzOVLmm7aqnvMpvZh5SJ4LfK
xkJvYfYETz2stmWVfxjXzY7s0rZfP8Vy7rvHNjHJERRVEN4An2EHOD/YDUHa
8liXjcGKkDNj/JkiXBF7quV0DN3IAHNPutp1fU8bf/qVHjJtxeT2NmMnWGrb
XlzJjV1rHtbmovwJIo8aoXYjBx2G45/3FqTIZDGZSiQ0x8wQEhK88VwaRQRW
takQsOXrzsu9xMgQXMyPW8D1A+nSqY9owZw+LnLflcuiNM4zYy/cAnc3YJSh
aDApHyAqmpZfeoHhJWwg8WZQfxLgXxo+cg8ey5s7r1MO0RI8/8o/7dZK4CZg
9dwdxeHqo1ndy3WWkHhAvcEVEE5OgLMNh9NIeSHrKFl0IY4xJ/grK/DkViDE
sITL1DZOIQG9dB20F6uI551RSGcJZiLzFMQE25E4FR2+Ok4d6atNx9chK7bO
YMNNpSOArJjLP72vzMCJLDyZIAYk2bGcBwK06Ag3BesdHcluJz8DQcxDeSvU
hB72D+i14rkLR5uux2a0YvMKXT2yE4SdugE818siM/SVOYC4st97OZkGHLQu
9jslsa1siuBRibk3VsM0h8CE1JxMZZZWeMQ7ZPQpfzZRASm4AD1+gQjbxQKy
t6ow9JAfVOCJW+eSQigTq3TZbJ4BYvwXvszuK1acfT8tWIXKCRkDLn7h0m4y
6Prtseqr+FEBp6Fj5hSU3e8xr43J6LRTjHzrybRHNYRA4Ny8DHgl5OTppFR7
F++XzV14ilEgGB2jqUk2ENeWQzZsbeYDLnuOHuhTjez+9vfCyMMrrknwetvz
bcywT37VV0V8X701jfGQKRAg/91IjDQxKrptYqI4wJBeCF2avtXR47LPmB9+
kVIxsCSVe92NvEDA+VZ6xtSV5ViE8c0c/lk6mFxyze51oEl90v0lwMh6HlmO
3MUrIP4c1LX07RDGWl/mw2A9sclbLB+yoTvjHA84zY2hJ6DbmQTmpSBSt7Y3
Xevw+ss0J77YZ6owaDy9YOy09SZSvi+i/Y/HOSbInjePkqdD7MU4i6SiQvNh
2qRwjDNl+JL5fJwmC41CopY/6neOQdt6ODNBxiAe1zZnZcnDqi8ElI6543Hs
MsexkdCm0WUkvgcvz2v9j9goGE21WZzTNUf3WhMNuc39ECDjpq3XXt7XC65l
ssru4BD0eAkv07OrmupVPsR8rwvTtYjoo+IAcOMtF/nr0OEMIgZrtmp+0Pfz
cU1BHY8vr4AYiUCiALBRxyk7GcIDZtBWH0hAQR7+GVWZ3wOyAOxCBWw0OMqU
2yF7csdvp217ACT1tUppqonpU3LrGeQQdpvxNs0z+weu+K33wCtRQI9wBPEJ
KYXQYicy9nR4mDiRwAy+MGn3GG+cQmY2lMWaZnTBFXQ99QiVP02fM+VsrkGX
GRq/DeJuw171OWA+gRLtsWOv/dne7pSd9Jc3NrEXkqwUO3E/SwxhAkQE0nLs
vMj/GjfPYJqAZDMqxWow9Y6ji+V5hwjNpRHhxvj+IaOO7JbsfrbJZ56eudiu
+DqHYTClc3s4d4sd3S8LIa+1hBDNOWqYYQBSvE9rGmYgxA2bb5h2uCIRsXQY
fYGfoBOyGW6+9Tw6OZincRW0sXlt1Q8F78XEoVLr2p9uGHC5FmMoadIzPVDg
+BLlyXS6cewVZx/8zxbdL+ThA5atDidZchDxThPXID5lDKRJxh0vlS6Hw/C4
E54ldovCIlg+ylSHh2cG7Le7kK+FFonPQGV39iVINiv6+s/IGBzYFFIHQ8kj
pnRfKpmBlJpDJKSUSFSqmTGFFmN+oXQVrNc1W8Vm9TA1d25f6ns+Aoxgqfae
l2Sw/uPbr91oodrK/hIQYRgdHng8mP99El+zyHSk0Ndu4UQxZSoVzyLaF4Xi
J7piZUY2FZfqgMV4T+zuOwHBTou9gTyCMSWwKyjc395vG1cbNmxLI1aAh5Cb
fOWomSlOPn/DebDe3b2G4uyz0HTnN4rvpbzk1eTdfhWcqKQ23Lezm3TTTP/G
pXMUP9xYQ9vK765ARDL1tGT42FimlE3gjOYLVpneCkKQdqMCFD2t+7Sz+Q1a
mQj1mtvKagjLoaAxmb12ZdD7kRfNOkuPTXBj6JlU4uJkh++1vCnFHwivsnaW
loDla049Dwoax2rFOwCN4CQwktYgTI1YeDhmhMrC6O/koY/oA2iHJZaWHd4i
MAchTxtIg7t8dGkRLcrKJTu2LStBd/eAHAg6pt1zTb5m8aJjZSH+rEbK0Rc6
Dy3Jr1ACVDw2Sjgj4IV579qukGembDEqvk08VJMxs7bI0coCEHSh6N0XHXI5
2tjeA6sgOZwMJc+NKTv6SqQ+41+jN85dF8p00VG33z3xuB3ZbFarB7B1kuEc
Nt6iWajjYrq/dAgvyzK+qypOruxwKuAQaQXyezNBCrlTP+qM2sRIJv4im9Dz
KjoHftEr/b7S3qJJ+/vE3hIy8IC7inMH9k+c5jTcgBZqSm0EeU0AGywRpUew
HKHNH26IP6XlBNaEeLW+pEZM6S8j8dJh3ny4iRdySxdAc7WomRCT0Hw1y+Ow
nE7sAP46+/UgMLNK4ChVL1wd+1qq2qpunhKfn+PBxZISUFmVXxHEpwXxkAvj
1lWekp+jTMzumzLfrAqB34THdpeV3XrQQwvG6TE9lw0BnZOMWH8AVMBJQW5d
Z9AhhNBU7vrwIkfa2S+UUuT9uulyJ8vBa/y6srdiWxK8sGCIzZoJp9QJ37kB
Z1zMVcMxW68ZFx4F7O4o1pFrKBeNosxCpus1Lje7Te3w2umg6XtkTyUXAaNB
mNeJgWrWu/Wy/HRjrf50VtPGp1LROfn92DJIJVRPRhTtUoLO/Izj2r+JM8C3
yGjHb5K2l6lN68HszAFWgLGcRAJynqne/ydIt32ASmt8YY7qBk54eyWxVlRA
j7NnsjOUc0BWNTWLiD9vsXKjNCb0uSVcUIPo6nL9sNFBQGbMMNjTz3HeyBY8
PRNc3beoJSRo7Uz8I6ewkTtQ/VBab5AR08dcxHYfDT7eVOfc//o8WJW3hD7M
cl52qpcksPCrOxAd/LDp9WPGXfuS4PylJ1PNZYdeHi95qH8AUzqQQMEJjQYP
iGmZTjSbOB5pVmC26PyzL84aq55niaWP8XBJNZawx1zrwMFdE6jYOqPGPJW1
5iNE6i+ZxvCj15U1829eonEmtuLQM1xUxjeT6MqBu82Ff4DpemB1eeR+uovl
/5Q2l5KidbZikhe1sVWmX0RgW8NXJF3XRBmh6p/1LKOAnbPpMzA9/gI4f2rL
w/3Zb0mfTJ1mOfMBHFTGog380SdgWP7TxoGXwrZHpFnC85oeWaDmw8zVwo90
kKGQ2Qg8AAOUixgsEkIHJ80x3WClWJNT0VJ8FX9IHDP4wDeCEI/KvLHUkH47
nxaea2lql54TYuLJyZ/1H9zV6FCJDJzY4ovrHjsp+hOoWApNosrYJTAX4dNb
VVfwbcHpsu3/g9ICIg4fVY92+JXnHFEwwog9wUoWKNxfU+nK7Rdvv3g683PZ
lzSKfXqgab2kSs06RTM+GEP9j+lV8ZtqVgU4LS3tensNF7bkrAtl3JYHVK+7
6JM8FPENnFrHp7Tw51AahTpqyUgGlL27r1sB86QKG1bIAkFLMApIStIdqFTI
c66+njeQkSXp0HPEmiSeadG9BIZ1LoUm6ZxzP9Mhr8Z4gxR69WoRHV4Wbk/e
EiP5xsGYFmAkBa8yVKF0RtNfN5CpZwJYauq+eokkuj5xqpK2kCFG5JOXZ9Mr
IIWi1az+91xeKgLo+KwbKWel2c1G7njtrwkWWhQtUM0Ne7UQxV3ljGeljAJ+
D9NOzLkOWm9K+PeupJhesw4BAwV/BakfZk14azVsh/qSxEVFdRC5caXdZnlV
3RKDTH0EVcQ+6kWDKENrnNap11cukmcFEoeePRhzpnsjfByOg/ANY7s4YL5g
otrnyMdsx5Y5xJrV7V3Fhq9IASj9m3DbH6hH0Kbji2pRyBkOR14nqR5rtS7Y
9ZrBEVWBKuHWHqPtRmA2uQwqHqBZ6tPOSuu57+X7kFSx+zpBCvqhfhgB//RU
JzD5U2qbh1g4nMzUrx55YXk1j48tSBMau1S9DElLFFWNQb9W8MUwAxSLZIzC
R2f99iQBMwO28uu0QoD0AcPYlaWoMBeZTuaoyEqZjcgCyKfLbt8AAjYFPDGj
hnH26EBoGhqmpEZPsEkiw1NRv7mHMZ5X2Zk6bjIbh/lly58VyISzqN7d09tn
LVS9BGPM84UzAx8SPLIgR1TbL5Z9rvTheqJysw+hAlDu7ikqXOgJc98ErnlD
tmUxo2t+whuh1WgkB0pA5V6HOHi5L4Ku4N77yp2iB+UFvLXRen3miif0/8OE
3QLbCoX798Secau9iLrpZf5wZg2xdNP1oB9Uiu3y0P1ElIz1OxncgDay8UkD
it4Sv2T21CqQ0bTcP9o3MI/LR5DCoozqXHs6tXuhlYiTjjh/rWW9//IdHDTK
O+3MMmlc6+8xPV7nNYP8xfvyyWH8AwUPUcGiqrMH6kd1p2X/i5nVPCO+KIng
hkbhOQL6/EVQMseiQnELE1/PZpp3FATc8W6efZXUsR+tyUS2kLhR7YYJ8TjE
E9bUWjEH6UMkkVRKPW3r3OT+tnsC1V5q4sTBatjPowJ5KN4M5K4Z2UTyJBUb
9aDh0mNJO9eWD/uME43+vyjh8UyS8idLWC0Fs0hmOOaqKVkm4WWd8/fERKjN
ZV2SoAqASHJGbm6c72OcsLJJ/j7XoCgNIowSKbvdRqGYFoJ/k52oPY6vBd6G
y9amZG+qCuCJulzFWSss2JjCqwnTYJ46alKZmQ5qtO6I/mwjGNWWJ4nLFOmQ
XEk1dntRXZYYt2jeYrwc7CGhMuvpJyfgkXOKH+G31S9s148aUS53M5H/OiSk
4vZzr5+6qwTiuoVoI9yfNdSJRJxpvXn0uBwOPf7qekHeQzSiFINNr+G7LTfv
RhSddKUqXfvqzLxnX4LENKD0aApVQXnIY0MWVYtFJ/l/9uL3sOqJlttbQP5P
wevRzB6skhLtWHLU5Tp4PW5oDYd4IBJ5zgPEnjf9a3B2b4GT/+ytRw/e8TN8
p8k7lQksGCxMuxhliUr756/+uY6w+3fXud4F0vFjrx0yjv9ilZ9sowN2XDH4
Rw7MqPt7KugzIz7KObgurCsMHmERHe3IJNPwSEZPprMi0jGNzaeyo9BVBMcK
7Oa+YW5R0OBvybreBKQb7/m/eB+edi612eFWe+NfgdLt885JyV5TU8kyM0IJ
FZaMObUnrHYzXlFpCAtJ7FGnIETF0x/XWb+BjpWN0Y96B83qEohZuOx2bUcx
cCk+PPwILnENUDTwozYFVZqv86KsDBY92HtDEax/w62J38KL0xbh6JEeVqvL
whBelpIUc7j/x4HRMJtDpwgl26d87x9fDiUS9S6rufeE7P6sf5ZurPGFtajU
j+Quvwjs/+OveMyx+Hna+k5q/PTqXXFqYBFApmzOYf7L1okztF0yoTQlzj5l
0Se0CjBf1d0VRwO2DQ/Vt9fve0B8oyzssZrIGA/Q4qj9VZI+bmDMuWjy0iyc
6G5bWzn8IfYvTTNSnZS7k37jK9OY1OWRvoKvJ7ocWCn5JwQ2BSse2MCcsuGy
j9eIeWB3qQyBRs+x5Pv1YXMRwrfbXffEclaJmWFgayGF/oXJgDkB4s2oyIMp
rFTZvHaproyYSynCIiK553V/Mtd4+WR9YaH28Tbmt3/RGEFyIj+pRG+zn8iU
LCqqzOrNDEJoiiNealtqlRqgsqHRBsnHboO2OnwHJmf2LjTJxSzF/XPuRERU
s8j0tGCnv9FHI7Xo3pJCa9YStVR3R4p5RFoIX04tljt95mC5T3qArbqHm3NE
6/tk0ouJVcaQo25JapStgdv7lzUo3lTjOzHvU0D+UfSQQ2MDsyjfxwTTCICX
HL2cg4EksFj4d9FF/pTk+PwpU6Ow7yP1aMM9OVhW9ziRgJGNcu9eNkuqS0mG
65iaKiGkNvlAHBUiEcrsaxTwmXn53IUQRVd/ugy6xFXPu2MHuu/s68B1lu/f
C6xennvaBPfRmrvkc+BEhxxxJfo7Ngfc2W5Ifw1V83Tq854WuyCDykVvZgPf
F7sScML/FWVqH9vXLeOKMmVorG1O5r79y7vSIyIllcEiVdK1yTAIjZssrviB
lMpgsUIXlPr/cMlBCremzNZTf387YFRs3GaTUhz7m9ETxgusy+o5fDOCqoIg
y8X8J7v4B7SFRE72zAqlJkQBgsZpMX4oMtAJB+A6dMJeo3HtH6lFX+2KxmGr
7uIpX62nSOsjn7jkRwTXC8nK4LKLfEK+WcsWJssvPIstvafZMgls1rNSUunN
ODeCFgWSu4xpyPHiGGtMmGD2afMIYOAyZKYEe3iBCrEQKqcTjJlN2xMdwHRt
nwqXho6ytAwAahgn22BtHaKEvdidykEeQaGCaHR1QsV58xAlLsVUlFepR6Cy
BfXiRQwTUCWGJRrpyNmN4qrPjmAkCz7n4QdzVpFDF3aZVFo5e8JeO0DnBQ4J
FQZe8qfXpJF+XndmmqgPHPmvGcMX5svi4YB2mAB/w9V1CcqEQUQ4VHghF1sb
kn7IIsNbqLq3FuvYajPtTMTo2l5HVGn057fCqkb87Ch6K4svGNFtmCEFE/tc
ZkLwDP+pUmtueKaXDrdzWTzOWWpXe9uMfF8pYhSgGqOtcnziAgabyco+EFb9
/PcQ8D9RKtoW8QkG/eSVwcLBHEgm7Ld4sd0Am6FDBkK+sbljQQj5TQCTKuTf
HKVXerSSvAwoheeIOK38NDegQJ13FuRDWsWJt9p8OUEuFNeVZOuvMcBgRDrE
ACPN4MuYqFeu7r3DkzFLMydyYoFYeQAvLJu0Giv1cajTBz+VFEZnryRtC5vG
dKvhfNbhsWjOgwyo+Dpffj5rpnhSCxvjqy9U+vWM3NP/VTYh0V1KYhXwoJS1
9a9v3AMBk3X9GkWsVGf6su4L0gCZ48b1hzy9RUh0k2kBhgZb0h16Biy2MIBv
qVG1sLFJ/uQWKT5UuRP464OdtJwzqxNHQlCNJe0pYbFKA3Zo7kVkBrp5ZBwU
Jmleo4J12YAvljEnp6fV6hLZ2nwcywRV6axzB/VCNRGZefghA+31fhRF5RW0
tl9LXGAKoUhq1cSV34dZtPts4iq4lQQMXryZidDfncqGH2orBqwOEPbdtBrw
0GPxHhpCuitlbo5lijljGcOW3Z9nlebidBVERvoHJWLtCgabapeFf9zheyGC
7Q5It/CvRfU62bPhkDVt8yz3COsXCgOYyu14VaGyXhtraUcpkL+OrD/Gghss
hfo7A3QvXB1e23D/wibGSMFflyKvd/NJ0RjEBDIVvkJWUZwtMrV+UIb4jlYU
1V22rl6qYFOeEWeEtBBCseriidsM+n/xeC6XAWtOSCrmirWsp/gJ4+crOete
Mc0hILlaepHA/EnfvFqYKUgFs6un1tjgIl/Let8GWIwtBgDbYBBxBrtDFye5
rHtYddIdjA1mnnyaU7FCRZ/SBIfza7T/ZaIzfN4n4FRXedGH0gONNXrprbDG
m+IX0F3LEDDP3DPUlXuAng55Bcbz2hbKF8k65//nIxqvozgvnNL7pVQ4yIoV
RmIV8CiFjDgYgcOwzTOEFYj4ttvSggVgcyy1sV6fzrjkHvtASGZvEHTt15Gy
8efWfTpIHQWoAma3IyGXYX+eXltv/N/jQZI7SInJf6kEibRHy2oBeTbnOYw2
vrMrbC/qOr0qRzSrHpOwUytu7vHT6oVOr6xQe7v/4tJ72iWkoKAkXzDD8ZiA
hiIEWQT9h23LqxeCcvjBvBkDQ4aPiJTH4UhvIQk5CZT7HmJiP+PSNS3f8Fau
/TtQQ1IRhC6HuNamucLGe9lNb80oAuXPDgmJjNJIOVU9hD7CoUr0T8FdsJmq
aPZI3iWvQaNEIRwJWE+fRp2AqU/QJ/arVJqfYm6e6QZ0FGH+p7AvdHx3i34J
7AP8tqtxGweRxbKKbgzv7dAvpSwbk5WJMOILsOLfj75WIMxXAVFeIEJ0halW
5eyEaahUO+duETR3Gz6HN3lFCzR1V6EF6va/UiA0y/qwawVwrAQlrzmEj93q
uG2YnCrJtIQJ79R2GfQHRVARWCvpDL3rJsWBC5pPtKoDVkgpVifQQFvbD055
p8sqaIUp3LH2twTfpE3gQ/r/022Y2CPRt08GZ1BYnG6NPZnW7f8+gCk9VPg/
NyStqC8aIHZr1fzaeRCDWznW+zgiWFtfI3nZe4ZdUlWAZQDqCcdKn2J2CB1b
vVselxDOu/Z4Li8IZS2onwu1NHJcIheiVAjU47/Lk62qc7o89cK62C5WqST6
jo/Emn8RHly/VB89O0b6Wq38A9BsLEM2/GbXzuZ0fU/rZkAkHa3xhWXDutB8
eW98D8Sa2qiLo+Q9j9B9ZK9taM/UJsllKIVbQDCpW9QfrQV/IjhEGfr2sMPP
GNyX8+GzicYA0Tw7f65WJGbPDAYAwfIi3ZPicE4ggnXXP6Nt5bE6TLtC0Eun
VMiLCmE7nCkXJ7mjLpAidHzMyoGQ8M0rJOPdM04jFOiB8prEdCNFfoKvecLI
FB0lOQwnzFYUXKl1yJm0WEsDb9Ila2WI7GBwxmcrOQfrBs0upfuSguR6/Dyu
FSucmxFtn/oJY3reoYtlzHX8q0VigaYaZ8i284cuVzj/xCKXt4Xd/nGhsVx7
ZxivRUy8oF6YUHhc7u126coZnx8gUoLIH+p0geObZCba9RQc6og7Orn3h6xP
9zas3tA9DGFFlj3BmMsV1HyZ4d9nZ8vkFvLPdqNYsapqEt2joHMlICqn12Mv
0bniToHbeNxQL4rhOHNqNkItkn0pWdm30Pv1TIdHIzvpUE+cXHN52oOo1KEk
6mhX7q2TTsA4W9+GZsqFeGHzhXjbR0CYckPczJxwwBdc4huzUBLAXF2NTv5r
D9YOXAA4IpwJ4V7kgieQQBe7FmnjOBx9vBDjkZo5JFdK6JlHUCdiceUn47Qp
p3MH8uUQBzb2PZZ0rXplDRxenAoxNgtCNAW4jfIWXmh+xHh+v3cOqr0z480d
I1EbCTYnqRB7K1Uw0AEBAUkFbFBW3i10zuZc1orL8W2FlWzNP8pQWp9lkWzH
WYYoPriKnt3DCAoLM+W/RBs5iysUtRKxMSb6FEAO1pSFFebSjDtzU0g9haeO
oVav9uy5nfcwGkD+BFzho3KF9UHC80nsJda0lSP1RdFDhNBj04+YmBLQ0in7
88nE1XPtNVC9UsCyvRQRTg+RsUG1kHg3jyT20EQbXeDilMjQ4xFTF1yvSgXq
9peqrboGgDJ0vJVC14BDEbb+0OSnueJh/Pb5Fsc2x1JM9u/Y50gpRvn6elwg
EaEK6EbZrreDvQqesiFXlxcC5UUCu172Pavsdxo9KrJKXqJ1b4MZT2Ugp1Dx
XcHu8QKCzpxespkDPW51ZiNLuLmTyhcs5DW/6ft0MyNFjjr6SKoF+17TYrOr
dilIcmi95rFpkNA4OayU2pQkblKsgXH/NqcksAZOtHR3idakvHRuuoZR/VIW
B1BC76KpQb1/uufbjyoGUr/KiZn9+3rGQ9mtmuJrHQQfX7c0WdPkoFLyiGAp
COUivSQWrEPcayt7zN9/UQo57t3cWXRZd8yZc8oyfnmOxDAHRS5YqyVqFxtJ
V36C2BfNabpqkO1C6cDJnZe6K4QEuYmBqITRwqiIRPwqmDfvIaISooDvatvZ
DbyrFoM0WZv/CWq/asuDT4LJSKWVlSvr2U1Pu2nnkOLMcgzWuxF19rvLMTPt
45H+amtb8q9RuaNp5uxHve8T36F8WVsFoEHCRKzc3arqmsp1h/rQ4jPMpHwj
CdKL0TheA5jU52oHWeRmWypm7lgV2CA0L2C1lDSayCw29DkiPKdhE5W/o6E1
NsMwj7MerbB+HKB4dLArKcgvpZmeEKGU0snP5ensNlXR6VCubdRz0pq+B6hH
mwPqMWviT6QQnislo+z+m6TDSdxe6QvjRJv3vbeMjR+/39GFG/u6nu1+nlNx
JhWP/gOOpSctXMLT4ahZEutlfAWtxpImghI+SNOS/kMQvxK2KpdpoV6TdoR4
/tXOdqtd3mXJ/FYHy1m0AZjogoehOfItZ2WmHRebq2/Cz+sZEPiosGtQ1qfc
ZNUs6UNxgKyS0DZxbRyeVHo5Mr6f9VWQx+98YfbKWPpu6hyshbdwsA15Xk7/
QFuo1LEvkJ73qTw74fjdX9kEiuu0bKVSE+yzsDBQAR0X6YisRr1gu198jqwL
GeBPqpC7ffJBrHCvPq5ZHcuOt/05URF14q6LtAi1UK16rHNiEnkbePRfvDHM
qb552XSfVuzrqmERao4TMdl0o9pOnduJeck2Lj1TEVaTwEGd/WCySTsD49+W
UpZ7wm+g7XAmAX4XjjYQ+sYT/QuRoyz3j8K+vn08DP/vGWtQZK++UglKgcxX
t+doV1NmT8enUDhQ8Qlr9M0BpiqFkpAtogAZH7DAVjB7fveNFIufpwy4SeLw
p+BVwTa7tQAj2mogZhxeJi3B9qrFFP1RJuft7t4GgCeu2PEbd9hCxlV469Hi
gpkxcrLGcN/6+9BcL7iWHjXZ/ECJDwR3LULX/qkgl9VFFZlYsyqsaMqoXniG
kiN01Qej7cgdS1O/Ik8AVaKTGn325rj9KY/HrZzWCwn9C2zBCbAXJlUihhEe
qJlt+8rtTs4ND1KteXBHiuEwSDJvM61QnMApMXblrp99S45HNyLG7NJimmta
j951qM3U4peOK+rn5Ehn2eEBvkk7ymmlms1RHCHP044Wxm/O33+0QUpJmtmn
/v56Q0nP2Oiuk6I78c96B6BacgLjhBPnZPWNlmEzOQU9jSHKOAlel8hDBbUY
ykPe99L88Lh1Fsb7rJW8vXA5KqoTl/XuphPC0PYHWp+4sZ81nvj3kALGr0rl
PYVM4+C2sH9VxyabRG5kHVpAy0CB0upJqLoz7Y2Uu9/mENiMacRlgvGVufKR
mevz+ap/pYCL7tpuRfFT+7WzBMlfrd913CHyrLdwUpBoQ920G6DMTntXQJ89
3gRFtn6YJGYGuaPHf0l22AIzyZQfcRBwQtKm8cdUXR9dle761kcBAAsDzCjF
uhUJiW4XWmEDEcxuwaSI988J9SvEQRn/8Vzp8StKKQ6b0c+ePWy+QCDlGztx
uTQ55kmL3ixK6LqBN8kAKscnHD56McBZ1RFrDrOnv/VU7zCnM3JQf4ICl5JM
MxPkKa4S40CxSNmBz6PLAWyIW3SDOhGteEwBYWcRYpeJUH4aYnF1izsOmdKc
7yTU/OmWhRBvb4m5AWrZ3DkLtP04XlBYGNH88nWZvfL3VWWi2erTLDj79pSs
r/V0kqgucoKmf8TboeNSZBFDV3AqJUNOwHmIbLH6fgmBuDp2jkwy2MnsFCBw
j5RNb4TTg4Osk/oVIo0h6lzBIjTSY7rMopWVciIw/3llt101O1oOVWTj4D+T
RFoBX8ZghTLDtImQ9s013bhoCHXrTgQk2bXDvISMIhl9TGSSTCMpwKGZsvu7
8I0c9ORiIxoCYSBd3cYNpyfmcyqfTjbC1EXqkmGIExn0Hxs1Q1z2gVxyEQS4
P0N8a1K2TOIGr2xvowRcY77mWyIoxhYISW2kWI97zr/VzTlNpsHSMP5VeLIY
FayZbg2G2YvPxVY3WiIe1cqLsgnsAWomoXF6JgdbmbuYUBrFAw75OeFOCU6M
ltXcXNrKMQbjM8uDS8Zt9Ofb4p8Lh3MoTsRYdIkz2uU4ebNXwuEPAL24Z4et
UGQWz/a33Kim4cnyMeTPvlSbzhKiCGljucsydyy1W+Gjt8H3rhp+3FLtptSg
pIx2M9UkqXaQE79maYJjtA0C7Pzm6ikB4rcNvBG5gepTZmv0V+GvTg1rHuOL
+wM3hNfdDiLPlyTI/JXmyySTN1GslYti6osPxs66h5Fe2U4Yx/fHtnerLBKv
gTv/Z43/YBDuheeIj6kr/Xk+XkeCj/uQt1c/BlaOGOdxZ75qOW8D3iWvugCR
mPyQxPoIM3J1PUz4RaqgslxRM8vAQbbRKuEcCQqYHIYJBhVyi/pVh+w9tC2y
kC+kXu0k/5DYwVDwwLjUxjJzuEwyLG34RE85mG4+PKJ4UrzjSCDwv4WVC+DZ
BUjMmnPfBhqW/jPBgwdA+o40hPxb4mEnh6AzCrNrIl+lDxg+yzf5VKeiF90m
Vs44DswvkQCtRFEEOvQyv3tccfnHm7xJ2VvrgXqgweKKDBC7V+0Hd7yD0yhV
1SK6XSJczma0F4XjWOokeRvZj0APKg3V4/0a8bMZ36+U8qAwNOTiNANYyWEf
6TvLXfEtiPefMGET2olRQpOehNgDMEyDjT+MyjokTm1KvhtivkbUD0yEro6k
Go92ZKpH5Fzo6TkyxWXn9bk4ibisZLiJ/KrRLBqWrsk1phvOV240F/lPQ6IA
b3lqlpLrKVocrWDAxtXlniv1zK0cXI53Wk0zPjIH6XKHvtxRHfTwr8uL0j9d
L19YxA7Kq6rE3fA22kAnMNR1q3sClcAwc1r1Lzv+6gQCSyfGtqbtUOjTQY+y
B5Ppik0aPfvPwT+TERs6D07O7AqgW5I/K8ubfRA/YatuVh34g7td2TyUlABS
5D4EGQLlvuEDF1UL+kVZwfgkpJYT7QNBG7fs8ooC+8vZLMV+qrJTRpn+HE+/
rPPvMyTMn51udAR+ARGym4x0QdPMMwQayz4aKCWZcZo3122CFFlHTXuNjHps
u3qjpqSabEL2BcBR2D+VlctaE4OlEUj3wSf7UNKDul7z0qi4UiYu8g1ZA3vH
kDbD67oV8QN+Mf4/tYnsRIycrwy+RSuWuIrzUKJTrDNn+4Y+XvV4UtAk3Vwx
bqeKt2+GtN45DQg9KIeETIraYugZVIQQf0SrAMPnIAKPloBOVVOZQ7sQuoCm
5kuwVQPAhBQXFbm22uaBIP/vriMkzUfpyxxLTTCNuqBvhBKolPYCfG6S8/km
10d29uuhqOSKY53F0ZlUmZc53Pow4YmAvX3AdnqnieZWn92I0KnYKZng2oIW
rQXLElMsZPsoBX7pVw1GWJRiUBfqfKoWRrEJsBFRnTeP/Kn8vgProfcRdf/h
tySR4LGDlrTHQD3imAL7v6tZPppkE3bV8pMFsP3fzOOCV4DcojDz7r3TzTXM
h0Ii7dp3GrroZV1MX77rnPShUeZffSbK3CeSCfep3fGwn7C/PVZbyUzZMh7d
BUAP273vGLCRBaaPwbUa5Mw/td+lbm8xj1VMy+apUUxxpceQcT8kCqtOKX04
UDctdc96mS0bKXzOZ3gECJygaNY4yFVC2rS2bg2qw3C2xConzFP1Ht1I5M7Y
cZC/RMw/GWMkW6eMCJc3PkCK+Fy0gxPBdsvQzSrR46a7jS3gznGPrJ/4v84H
iZCHNV7d1GnISwFXptle+W3a3Zxwv+RJqpHuOedP1TNVQxXsa9KcERdbD4UV
yELKPxV3wGzTzHEET+kguwxiq/WoxHJP21Elxs8e2fGYIDTLIfplF32wZ7Pe
PxitK+d1G5YNMbmF7edBjO01ogSLTqU7Migg7Upltt146tEIEzjXhbDp/wPZ
m3gNz7jx04Ed5OL/nEKIZ6Uwz2KGd2CWBk3UXi93iebDRIip9D1y8RCqNYXH
843IDklkDpa05dDaBIeoKXfXho1QA7R0T2+uT/mjOj3JFRPPkLucON+EMj6o
+8NuNWszwst7HxnCtvMW2vpHPzUBd0M5OGeZE01EY0fkM02BfhzBz7h6iYvu
NnLTUJ/o7nWDlXdc8E6mSS/vdBz5zsTpxdbx0xt4fk4O8/x1zyybOKw0IDaW
TsZEL44h4YPQGL5irNoaPoK30mkzCTwEIAC+b1E9mwIRgqLEJHua+CHAhTdA
P59Qzn85mK3HFr6BJ2xmYMeT+xeU0f9A2NpAVbHEbgCXWcYCvVX3Uv5nfblt
qNE9C2IGk9UWxCR1rBdwJy++lSr9pHVdO+Fk4MbPMx0ikdYULP6Pau1EOXIh
kgBzq8nMPXttgsMiby3TsSbdaORrHZEu7zqy+hXMgtK8pfZZVy9eDZKhUPvD
nEpZD6GuX0MWusK5R1uKGrWU9m35SB3hAN5ZbWhW89Bm39hT+iIwoToUtzjJ
Z6Ry2ooF75wt6tg5qL7qqPZOS3Ln2YVrHlPt5ZdR0GkqxAGKepGo46KJLduA
EH/cNmYh6tj/ruN/XXXL9K7nwXy1+HOZIwy+s0H6HvJXhj9n4rDEjqi6NZzD
gKRPDkA/qiKNAeUxFFP77YoH9L80olGv5lXWs+1w6RIzukK4Ih2OBaHekiQf
1WjBd78EfgyvaS84fZXAaWHm+6+DHHWGDfxkOgai6vnEmlCfFe6IS+Caf7ze
ouPxkDUUNi801RAcsaA1OnxEUSYzB8M84Q7cX25Prhq7wdI92zTH06os6TpB
9Q0SpdG6SnRz8VwAWr7gzJPiniwPBbT6futMTWZllQJl1/3uTHRoiAwNtO1a
Ll0o5QPxdCz4yTmLX9hBeQ9XTgCgEBQz2UMX1QXv4HmYNEtff4eU/vGmrooD
Wpakn26AS55N1HN0Wo4TfLCblQpz1wRphRyqsYm1BaYxE+aqPEPS0QvzWl1B
yV9xYPZUDGyO0UFe0xnn3iyZaYjlXmvwC3uSJdwuqPrW3ZoKFHhYWSz2Bopf
yFGcVHomB/yp+UUwNyQ1MN2umZ2ge8XaILaNXU+/4GtJN6eL5z1WdAjWvOP/
+m3S9oiddvZ/1JWqb7Z0WhaJZzrLC2q/Z2N9VopeNehs98Q11NziGJ2LaAHZ
BkzP77zOG4uCg1xztRm/yvYMSnF640ILF1GACpZpxPt+P2GRTPaoe/rWrpyy
QR7o0zowRgl3dtol3D9VZDp3JwDttOVZG+qhzr+dmiCMKlIO089IhCUPjZYJ
n0/FRRvdqIO7wltk8cK8wGhRn/a2Py/YKcdpnbqpJPTMmIVWsl4jyRBAmdCy
edw2h5vLY3wF+MNKECwJF4MVk1I9aAeYxK5ImmOpXUKS5gFna3sR5bTArv8h
nqAV3wZ8pVu1v7YTR/h6TeI+91ICLzB+IJGEnIX8yGjP3g3K+IESuWqrrwMM
Ppxmx2v9g2V9WM3dnpfL6anw4ms9LFyGvFZyY/2wJg6syxyzo15wFTMKsMyw
1amuW/+3lBy866HgKP7ZDOUaEZMr8pKtQydGe9q/fZ/T34va21CxYAsRrgev
Bmuodj8iMywaAiquGnB8swa4/9G4rG7jdxFoWQnG7xfbVdzTI4LzbPY9SdjV
1dUuVBiv/MQDrF6hDclRTpWc4GuAzqGle9U9OTOgUxSOzInka1EmQUepJg/r
8hWklZnBkg5Un/Jt2KwFmVTW/gp52OdoGFRAect20t6CBP/2ax0i48Wsx5xw
i25g8rliSiEfk66GYxzQrr2l1o8tO9VEMbNcEl+rVzkFCAX2gEsvhoQoYJu3
5MVCysk5/wq9yQY651+O4TGZm3WZrJxW1gSgHwO+Is5MlEUCbL28WDyWBYKc
8DKlfiZXW1s8yACDy0Sa0KAfJbkemW2CtgR55KruzL3Zq6Df+8LS9qoR6e6m
Fh45t2p9IUwS2ifVwWzvJOo+9XxJgbBmHf3zRrmZBpdciia36CH1wPxSbak8
Tp8KxZ1BK0gWPM9wAIpMH8ewy2pmww31PS0OnGuYD3yETavTroPC4mKobYUW
UtKinkPzeXOlufitYuj2Dicp9/upQjgLdpXRQdI2+cNc2mVbzaCKw2s0nMc0
YEzU9XJe8U6RkVE+QwnWDwH8EL4Bi0YHug0EXnWv8H2FhYU5ExZc22ojOMLY
Wc0BzmRB5Vaa9UKN4g2/vffzQK384B7ahGxoxd3PPGiHSXeRcza578XPvLfw
gRj+pL4fNfTM6RKhZL+flC+k4JB2x4rICxiEkngKmY6bw+16JLU9zOkIhKum
oLkQAHd3FrhcsCYCGL/semz1JerWnrINcqZuTJ1hn/zM032NFC1/pb/sW41s
5VGx/crq9W1ftGua13XYJ/Y7dmtcBUCm/va9CRa0bENKWb40TCLeEL9UMLkQ
k6ZvYT4ihie+v9+7leEp/i5s+Cl2M287YZIgmi+dF050bWjsGjTeS9tX+hif
Njv+yKS/sOXI/8x9w1Nyk6e6MnB24vrVk2ssy6E8BYuv8pI+I1+v2KKMIKCB
5I65OgshYenZ6uorln8H2weFkoyt0EiAhVUGelXjXrYprJXQ6PIKHIXwaHhl
HNVPffphQt5JuSHDK07uL1POZas0ker1C0vH7y4KTQ0iMp4sBLrV/tA7oyCD
bv2dSYYsYFpQstRwkcSBKJwFYNPyPBfi78A0Kg91rKk9xbfB9RS1Eg2uYC5u
R19jTRpBwj4POe88WL0WNVBt/0fWdZf3JAipyp365G46M3V/1R9zMRiNEkNO
+ClczyQk6slw+ggHAx6qAMSV7/nNvLDHB0GK/N5xub+yzWQbZccMynePw17T
ky6M+QM3XG9EWKJeqxKymywUehEpmZGexoeFCSheHBZNqpBywsFU9ShGvne7
tEKvzXwZO3BdZoUuSEX2LTt8ZCY4I5B5+uMQKHTjgFCfIn84PDzm4oZ9ZxgL
3oAhNuKhpQxpCgABLpu4Fc1z6xQqY6963VO2M/69tg28zX+EvNO4lJqz4xpw
yDGdWog0PPAqKoqX/Obu+JLQ2MFqyy/v96wYenRkUU3Al95/25zwTfh7LPwE
nxz/kCFZVoT6NqRp/h4YTO35KkjwZT/9qQZqK/1iziSjqMiYbrhyb9iOwWUS
pF6dlehzglfjCgFm2hCXGEdUyWRpMYMKN80iFoBhT5f5xWIU4pf+NOEhTo2l
oJO18RKo9t63o3qhm11UNALAIpPC4LXZG8C4ggXdLMwrVT6XExzUPu4PtOeX
SGUr2l0sHBs3nVSCzLS6DCCUaaOQ+U3IoNYPYe4L8hdB3H7o8rl2GotQkr8X
oNu50znCJE1G0tHFxB5MECodP1NSUB+Qs2wHEWwPKp67ApIqp9zB7myRMBu4
rJEQQ7YWxaBkgiP8p87kyGa2V3fzm9k6/O+9eCtYr8pIqjkOwyUp1n+QZfAZ
g5GLKseTDIdl0VZFXOvSZjYWBKnbEbRIN1trV0VO1SC0bhgV6ZMzGS7h0XCA
uc5O1Dzmr6RA/4i5dPH9JOopwsUqSp4xZ78ePOj+z5r42OjH10VvTF3lOPoe
g8O0O8N0thKp+cHcCRGBPoSrdNqV04Ksr5IK3L6nfmbr8zYMo9VeC0tHF7AR
/ajHhBA5y/x5kuziWrjB8dtVCVoDLv5wFn2WTD8D01QF2uRPSMhXW1LowWJ7
ErIXWrJMF8H75VPbcW6nhlqczerCBqiN6gmSvmU8UDWRlpt4Evr4tvobPEEe
1OoNl2yEFjPHR4XH3vBG6wtxcC5f9mE8Nn7TATWZd8FFWhWrh/TCLzBpUSKz
apz7vEIJBSGFGWXdJ6/gLMe2y0gxATeWjCEcYYcIFNihE9eG5wgZPGHTG3CX
p264EmKwx9TSu2xW88sZBHcT6cSTCDWFtnanKw+wkJFc8iJz6TEPdyFu4/jR
zeVt/rkYoMdmiukTymwovjcsDYuCUc0qWAMO1tQvt97B3BkUZI+vs6DeXPxK
XnhHociTEWxUBQAj5v4FEtrBsKqguvwAETdC41SG/rHbuQG8t1ei7y+4OTLk
Xswo0Val1Qh1GyUyfxGGnyqFBBoD1cnQsJkXzmAmOp1+yIAr6cbkiIsOZr3U
pxKq3EO4O5ZqBBwLIXCRiFhEiQ6Q0oy49KbrG4QMf5d+hC/pLjLfj6ctZIvT
SGHzMsRoyn5ZCO25a1rqg7QTsLnDRGUf2jQhizUuiGRr73ShiAXwFyUFXt1C
8KX8NLva9Un6XnxM4dTlYg8FNIH723+s426aZTlOn2Krx2bl8IQ/yyOM8qO9
52xEchT78sT8sqAcs1fxljmlVv77TAuL/4lhwxMoczpQGfVeL14zU41VnZSF
j7scrTwwuuShj9v9nILUkiAksXyXn0y+m60LCgAVq/jPpkvP256oHEqggqOP
cfWyqhHl1cPDHgCEjkfbnmdXyIwenPtj8xqJwURH70pezKo11ua0Vl3ZU/2O
kpl7DPnrHurkdgOMQzlio3VSil2hp2fywA/ib2mv2vHOhDIbQfBtY5Wacao+
Ht9adEPsVQp1k09Hsrh8voUyKZhkodj3ot/Kn6u3CAwZa+2rj1aMtP9a9FhN
u1D9+s0sm1ZGzdNDWuH73j0LCDtWBNjxV6l2RXxY+QSJ23owcpgM4jke10xU
UVHHOsJCnh87e/BL4dAI5QQJheY2KAJ4ak/+YlHGPM2bNSWMVD7chP7BTcb6
FTBw1O3pSw8S3UIB8UEBqL9HJP8TFkwoSiVyWxvJ3RkRC3juPZ+nrFfxE18Y
+B8PvyLvyl3pNLxBhpWwzr24QChZLG7VPx4IJHAyiYFPMgIw/aibwVt345Wt
BNkLdc5hABppr6va0qh/if71NJaNxmzvJ+wwPosPOJJf5X3fudA7QNa6Cewj
LA1BmyKPv801LqOSacdlUVpaVp6EpMuhdbv4QgPMy3NXkRCwPuhKiX0UCfjN
ZvF3l0UO3QdM1ejExUTfcbj+ntoSfuX7IcuSF6WX7rmM7r5MXSt+feQbUtXI
Wk1EwiCez3Cp2xbqWDi6nfxHFkDNdwpWLo9yZj4o2Z09gO6u574IBXuThOn6
tMC7n16TCwoSA099s0vn5H/yoEZdYnF6ClZdOgP0yqMt/Q3e0WOpfc0Csvvk
s63FL1GevhbvvgmJ9XmXwydWM1z6wpSSMw4sRLRNakZlFdSvSCZnHYuIieiN
L+6WA+qBM+AO9OnX4XcpsEnYrQFJ21o7RfBdfhif6K/XwMrW0ulYMrpyD1kE
ZZbyqVJ/tIku4ets4Rj981uTs4ilKYOv553UJo/wa0i5mygBJ/a4EX3y3SMs
MWgt64AtiktkfbJljfV2+N+xbMRBr+vPd8XNOoUHs+ij0nLQo21PaR5/EwqQ
xN8ATrZIJ/qNfOd/MqdUccJhkUUkh56tYj4YNzeRJN+PCwAWxgkm8eEzMIfN
YPr7lI+owkqKF8NB4GAsMMDLtcxoERxoPG9Ic4iDpWLYiAocdBZpqgVt5ic9
swYn9Ih3yV6jxlRStu8s5GySzWwQc3QxcKiaWaD73VnQr9B+dAh5S1iodFEk
oktLOa22Kvu70NszCdfEcBAnNuMs0iuhOq95UKsBTT0q5wtuliKwrIl+5ZQv
hxhRi9cJNg+OY3HV91n3+U0BNh0pHOvcLAIAuHJcaVIWDQJlpvRPC5NAyh40
VyMZ9Um6XZHeLwkQJybARpNfzwHKF8LaUBqcd3zPGEmqq4bLMHZjoUmw/ULR
nDXo0MSxM7MgQiRyzHNdaJ5T506wryOR4suQ14MOSJLapx7H+NMl6A13dr1k
p4lvmKMwlvXZE5sqqCaX9Z6/kPFKjrcMRf1mbIenAdaAz8nGMgh2BGNjmOKX
z6S59msQCpeTBgjUJLjufpVOHKNDZ44L/vY9qSSrnBWvmD1E2pMKfLTUhgSd
4tJzSffIeeNHT/5yGmbwWkqxLa8f/FXUGO0ELAwkqC1yxVICHtq7CYj2wLai
6QwfdWlpytx0tkIVcaEUfnTuteMfILkIQE83+vFJA2wVug7Ek35EEIDEMgg3
qbq3b03ZJt2x1uIG246b7N4xBKDp636M2a81c2gkZyQ8e46y6wLpNqnzp7Ix
IlNksKTiZOUh4ybpcdgwFVwIX9uL+Nlz/nMe76MCLXVvY+Ip2Ps0DRceaiHk
b6d6N6q9SiECQZWygnOxjgUzmf6GPKqmzHTHvvY7ClX3XkP1GvIiaR1ZudRs
iOC2qTQR5w6RmlNR58RtBlC7UH1zvXbibCDRRNO6nRn3Wct4sOD3+pdoDWpz
OhLjcTUdw9kQi3FJKP1r8hibcTP34OuFgpw5e93JdkEFcY5I5ebcgNG5XHMY
PYB7ZG03Zq3iQe33/tA80Ece29I6Rpzd6YterM50QcXaPo4g6Hoim7Kovn6P
zP4HcuPteL4cq3WpYewmskynLz2U6lgLfrrpWrLL/QxxPdFeYDWc3w/Ct8il
zLErUgIlFLOo8oU+cFvLKi41bzyEzhWpDoQC4dMKEjRrKtubhGWJOXk5pUKs
Vdom164hr35DDwQRbMXQk/hrurFv47EuzlwtG32P2cdwMcm4nHbLj1kFAPcQ
PJFBPJQCjLk4KzTCoZhU0cq3IgItyZtWjByySQQyfJYwD0eQlSIjw/8murMa
JFOoWoxwurRGcjly12YMuxGpM00EzMgJJVncvfsxYsIWxyzvbW71Bw8IzT82
FJQttbAzbUilnBzo7PKMwd5tUBFuEjjPzK4ttSyQi6Im0TJa1BGR+e2kasPT
LPRID9sfoKAJ/i6FC6cuV+eQ6+Oj3fmoK+E7r7huFAhSVF/3L9DGdhJU/VYN
3nMcIAvlhkfB9o///suOVgmtjRu+WsBwt+C46mHp0Rx2nxm48XT/sRJtOfKZ
wcSqJEDmTcYCSRGAGaSDTOhvfNAcCAbk7q9+qyskjSwLT07/OUmjydBvyGUY
ihftyrD97wkGP/TYlIEgIFg9ecgsed0qF3JFSyIes3UXetS9SjzyutdrOsDW
CsVZw30tuMjXbDi1DyaFjhMihD+Th2Xvu/Vz4nrYqjtkwvrU+AAAgzJPuIIw
izVDZ3Sw68WQ4xfhUo2mNpHGx5Anu2xeb44xJn3D4VXCpTteKGlMumlBI91+
LCbzyq7rYwyMRtODxu1EY1M8PFsHaBmDwfX8+181RpXeaDrdjNIqdODu3ZeK
mMsLOB+9gPabqlVEaSYYfMtOrMxU9ZGJjpoY1svtCh9g/LMNT5YIeK+VqNlL
5O4t4k9rbuPMYfe9pd83U9JDrulmKNkdrj2pAXatieQa2C1Nl6lwYnA/nTCM
zITL2d8UKZrvm0NhNfFP5kNON5jOp1GOjk2gCRfa3+abO8D9JwTSGH78ur9b
td0GFOlOGJFAT2NoSxKpg3tWB50nzdkLJmndCJOTzTVk5NN4tex8oDK2Dgkg
yYF3IaIL2647cReqq6lavljrcXuhfSOfIaVRQqZvUhfzxdeqowoYPCTG2rcK
z9w+P8wLAa5VZcpeMOSGthsCibO6a1B4+o2PL/+KlebA/g771Ha/DDlf6TOJ
ywm/xPpmoXzYT1OIyjMUmeiBTVPs76ft4u/z4wpNYOJ2zm/ifg22DzTf+qEP
Ey8miBBKgMrXPiER7NQgsvSAjCZbLpgHBCiFFTwrywsU4F8Zqv+z2LEM8KwO
wsNeIEF7FoFRcn72zQdzoLARn63u/yPUP00JGSzIFto7nrmUI13WrWgTYWZX
PqoRQeiHOUiUGnxz3CXbVrrItNfk7VRjlb1uMe00dYszKEmsqd3a7mzgXzdL
nos7QAaZu6tyJY9Y6Yfq/oMQ9G4veoUbwTBedfZE+OMz0uaSZsgdTjk4XfSp
eDMqJvyivzawFbddNIvr/A7yaqj4BmliFXnqxYOkx+HWgNuDo1uNDAIQp63P
ys+qaA98hm3xEKSL5Wg4RoxvtDKWVA6XxJcdMFxjLvPDoeDZtKagD231mHOK
kjEibQTg1DbXVmUc3uR1li0qgsZ6fuYxI6Uu9iJRWRaK55Xhc5OIzSv8iBav
EfBRxdvQ8v61P3FXKip5uzef1IlXiZmWr+YsZD8mhl2rjJ7roFLDVTiwKvLp
Hj6Ay4M2o/me9tlEaibONIs/I2N1TpwwpEM5m5E519KiWefRGLUySUTERyRX
XLLYYdtUY2sBef8Pjf8qPzyCg9KoweGYN6SbThq5e3IfFeZgnWk/TW4s8Vph
FG+ESk3VILK3p4AvvAtC/zShyXHRxmv9l39rlzWE9StGo3XoRphwByRYAO+v
n/0rMnTQGdYy8x9REetMwAtPYdq7f/yQ0eKmbbuIiqja7WqBa5HIUHuTAyP5
QBQDeDGR3w+PJJy12l28j6swXHtL5LCnSWF0A3BytF3ZdB+a0oxZaqaeWUJv
Xhny2kusNq/yh1No56T7cYPuhPbsKK+kPKRLtSw/TYC1KcIg2Jq+4IVb2gTo
18KStYbI/mjddDeYBSsMFEsaHBniqIr+GH2W7HOi5FSDy5nRg+0k/tqngg/N
6oQeM5sUu0NavHPgqC8IxAHxd0watWJKCbi+y/L9rqfyvAilZLIy4lyi8jyV
694u0DzQQ+nY8CAeCsmpYe0kVpdnOm6FgL0BhekHTxt5d7Wep0yaZ0Shbbvo
SelKQpxpzw36Sr2zt030akOVdJfuy+PbyMBDWalEEU0JQ9G2Xx4oJNbog15w
VYYhWxLfosMr6fTb9PkYAeAFxPqTypfq1rgPS9rf+aX6AUQYhinLAdUSAlvP
x3oTUEWmxSI81+G02XrMml24Xtq50z6JAVwD9c4t9gOVQbkADqDMMlAs+6OC
EIhg6V3fjvJvEZ4zR26sbj+70bRhs289Oier3i68DZNEPtZJeFXunPaH5VNU
rjJlHPxDUSwV1mSOnnLMogGt9hClPgokF1+MsVOL4+cYjagV+eX4IocQUcBR
IDskDzPiEZOwotWJuqcju+5STS8cbANfltl/2WedS9g1THUrxz22LOCu5jn/
DbHmavKV+bSMe3E6vEmuIy7O5W2PtZbtadtd2dexYSq0CMyAgcwCxNJM+laX
IzLCu9p/WD3j7NjI68XgQCOSFolzRyDv/QSE83d9Lm8p2CiZ8HhLoP+knbD2
68HlZLjkHXvJ9UpHvsNn4BE4xeW0UOo+g8DjgC0vgEgwLc9ail2UiPydch4M
FzFXnYcgEwJFzsVQeLb32gQnd/ZLWxk5ywjGMeUP6TwZmhWb9Mz5zcd4ebnN
xA/Qlqtav12j1SKmLzgJlz7+X57cT/z9uSXto0Dn9YJQ3jFTJW9nYStB3NBl
aSBN0VHbaCw2TsSudcMwE+/NFDGXKxUEgtL92Ka9Kp1R+UMeuQP+JpMCFY12
3qYJaaNqdVOjqA1C7KsR7QN87QWB0cyEjj8pakVpOKFlC8AO8LIgkdDUojFY
HDPOWIJrS+xo7ec2G+9cqvAKTN5WdMOrEAp71S9HZYzNLbZ3VxK6VS3WGvbK
Vf6wNVemEWNde8BAWX3haypQBog++mxEzKCXj58jQVsbULP9FkP1qUJ8nGAd
csmmtBnZd4arAvDZlnp2FoHoVbgPLJSFRo+0+Dr+PKFK0v413iMYKTb4srwx
Kw8YqvZGPmeUKzZUClccI2VzvBPBorKI8KmVGYKRh8OzhS6WJ+o3wwg7aLh1
j0a7X3NvvDy3cAUNk49HC6KKYYqSn24L1QO61qFlOodhMu7esJKblsowCYYs
e4Kxn+N8u1OgtIdi67P0GZbeMjBvOAJHE+7y6RC53j2+Ucb+lmJluUMl1yuO
N80W6k6rEZaY4FT1TUWAxF3vl1EZKc0klULFQbBbFxPuY+1cXZeOpZ2fopU+
ZjCt959R8YBHTHfg8VLOrFkQ3hQlCyE0E1Ef4hWncF+GCSG4zUqezOn4/DTr
pqwtAMja/LNg6287kid077/stktmOxYpFmDiIyaKRgrjiMmxZmUXjs+O0xRt
0KbtsNRXrN4i/dMyualWRORSMlCwRApe0vHwOjCtVCEhgTj1abD+Iw5yEjkY
dFXfywynGBG5GVWvV9yE6wPwKle0vwbqR8Qbv88aYT0zUJohUcDY2gDqE/vh
eC8oqewbIz9oUhqAMiUIMfKuwHcaOCpD5xrpJfK5bhs3gwl44Szjw2dyIlch
4vgF9LD6K6vNv0tm4hvBHtHqSUfYhpxcNeQFz5E70oRlPWEr/zjKv4K4w1TY
/s52nbhQKYqbGWQh8zJTgTBL+qowaD4mdZ1Md/q6dLGa3sWSKtuyNWeAQfJq
XBRU2O+wJ7GHHlCUQcLuag6RtMstJl9A+XExSexv1AQz7vFJdM9/MP37FZSa
02o5dfRTxa/Z6IgNUcdc/O2vyWQsGlerPBfGFZ5anNupq9I8im/kDj5A+uBU
rqAU0fKFhKuRbKrXDuKsFBcXz4d0Rb4mjSkGheN7wLb9ET1CUmGHSSAIB8p3
acrYJ21SQZM5ZpmRZzxn7BlycWIUNdmpdGhkAQyk2NiBi2+hTnhiybfDVqt4
Xsk3xfhDzc0tgpv96cloH3c3c24amb7AwV2qeaW5NmuDkCz6a2+HTt+iKkzc
p80yHmOrVoA1GdAqiNp2XGQaP727kOSJi3LKdRS5gRYck/+NYkzvZJLB0eB1
f4sNtNRa4FdOM1koJXbK319Dkx2RflImp9eIM4mGDfx/JjktTRizVQ9Wj4tq
m3IH0fKx0k8+NKp3YMhKdDSLpvrMDCm9qKuNdD/2LwwI9P9+vboWz8k3GUY8
U+CAveX5xK6p9j+/hS6JtI2zCCJZ5kNe1DeRgLceIYwvPmuCSaHt/p/w80WU
VuFUj8rwUKFO0S6uEf4tEVR5P+OM2dm6VSto9Lm76jhv1TquHgHKSHc7MXiL
nBnwu8e3OA8bAVpYmD+HDWTSNy0gbgl7aztXAEQf8mcAkxEMGEVr10o24iiU
1amF77W28gvae8r5pwHLgqGu45BfQuD7Msv/lu4pCFpPJLihmkkVt7jA15KH
GN3/a1oWOv6uEUa/cZzQAi74iwwi2gu3w8WqdogZZwt88X1M1MhJ1xI0MJp+
/ZbXtJftA0IQ7TqUMXyF2k9S8SUeCa3wZSZ0+OpYzlNltP0zB1VpkxgbWpOs
6ZcojE2+RnyC/KB62camec6D0KBEq4WjX0Tt5wAF4EhbUeZW+r5B5kzuzUW0
dCCNWwUmirquLayRM6TRwRSHXY8F2ZsiAJ9KHpSPorr9LBwWPBL4fSaXYX3E
sr7j39B8HhC2MPfDWxSR1QBIO8BcCtl71BmPym9UzCbE74eRBAOQkQrUm2GB
H6hwfadGFTCdoJpYuOpXIFWMmukldM+tF9e7l/ZiDTkmdnJJonYd99xt099n
S1pwDmZ9miwGT71w3sv0JpVfbzvQsZ8yVMq34YPcf1svESZsjcV2pWs49J8d
gk2BsTpORFBCoaN8pMu6wia4its9NY+0OWlcI9gJH4O2dH/6ytr89wXeMDZU
CWFv9H+IMFFOe+kji7era1ADNMrXPYn7W7bCSd3jKZNEV4MLTN92sMIUmaju
gJxDP2bVx0GEVJTChbN5woUGK8jVM6WBYz8XsJMVxyRDz3EahyvothkQNRPN
Dv73D6kbVHLS+S3DQIX9LJ6L5MA00ddgFhCPWWuBF/eO/ng59a39x9PXQdSo
xwdXqGrjivNUSCvBhx1GX1hKTUxh9VgOgOGxVPRYUhCqosQMEinxS+IZjJQe
RBg1OAYPpXxhWykOfyJ178esu5KEB6OTMCa+NsvpZeBdSiP04kt/PjUYPd3g
/mVWZ++mrJ1rU2kNEj8TfRipe/HIBvSb76j4uCHj40lALQTyzEVwB/b/M14b
F314AnMzDu5U7ARvIGN0MnT9TzkpXQf8nFMSAl8LJpbkLKOZqu/KPYCsp1SV
UkfsQDpXrcwXoxBW0veuSvtTebPH/dD9Px6B+bPxvMXDrdwmAIQd7wyIuTRA
ms7aCYYxYigtfEjI4nAlyDGtw3dQT9oYatqMWNhRPwfWMxQkuJvM6p1NvP2t
TmLYyYY2XYnZB943Iqjd+JKKuABD6mh0SxHOyOq4sZsb75pnsavDANa/Cgwk
rUdxnNbtAq4sQ+T/QJ0lEflywgKUHgrAuwO7AvJ94DjkAyFGlvE9WYvEpAI3
4wONExE8J7qEMLZ/VJ+qWc5DDVOts8vXI+/TNNJJHQYi/V67DxTnfgmsvnv7
PlawjvsGUjJqaoSSbSFxCSPqqdga4ux/YoFEqg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1JOJ7WklsTEoQvhDuFZf7EufNwu2om2BKL1rjeD1lhPj7xqKN3LGNs28FrIubcDEVJEKwc04d4Sd3AB477Gwha1O3T7VhrQbppuHKeJFq+8JSDQW2aPoDDJQ5f6ZRzrSmTU4oexFPigYGq5FzM5JO8XHx3+pXrj0F3IH6k3c94b6rIMK24ZZ2rDBefBO7oUv64iJP7nJ02+660yFpsHh3sNLELKD1s/Egqff/Tm5h3Fv2Xl58BOJCVBgYZML0Y3EOWlPWsNF3F3hPICYEAcwhcKlBR4Lq13fV6Hm/0htmoWjUgXmgbWjU2pdjsYybH6/2dPvIN1VDlLPdzPevwUky48Cacm1/MlGb3oFbV3Xh0ZTG7JY3wVWYn5rsfVkdSUK+K4Ln4Pci7zkOC9FsmqziPkfIPrd1/edZmLwe4NH0FPWr3Rs2TFWsgOvy+/mL//VOM9D1cUi4SPxqS37NmloU2U4bZRNzDfBPoXuFc8JR3g1AnkTiobAYpGYVd8O4XLGvBo66SRHv0+4+6FBDv4EbNqcv82BUn3PgeBD0JGmVeW0CnnsK1A6j/DLHbgCSyLYk5KHeeeDqaF46wzG2QfhC74wopscmaYqyNkO228LWuhPpH951xq5JNkuN/yYfoZufUEKVKeE9tYg4Ar8ibDETevpALelem4hdrwmPG9k1e6TNW1HT2vBi6pSp8UW1B7Nu/2XBIg9BcrBjln72Uf+9R91VHU++r8GiVU+sA7r9fyjk9tnbKiPoLyrkzLpJ0ckhjTyvGrYLtCBLHIya6OvR0i"
`endif