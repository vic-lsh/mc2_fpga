// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Tdra31RWqYmq5Qp/NBzx/j6STajY8RKaqmi6JyKodicouigcViHr8vCgIWh+
XQS63gKHOYjDf4lZpXnK74DXX787qUIlnj5gnshXYwZiPKdeRKa8iz4ilNDA
ZQWinkfJkdbmD6XSp2KlC1Rop4gszHK1NFgwGrf5VWQK39mU7ML2lRGdjI8t
iF9CeG/wTxEWKvYtT5MFShigzlNkVoOFSH5OFu1XtT/zwCvR6sZsTUJz8q4p
LuG7/IYCyG2kTYNwvh+TusoGgCM09Vg8ThtRmguWfPHavcN9BUU+XrGHUJSX
ztOpAxWi5t6IJV2ysUupD0iF1B8TQ+Co5XwArEUQdQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o2ZBgwrbMIuSmhh+1E3heUYYF3PSSIQoa2YP5+Y2aE9FcqiwDvcmF3fkwtrH
xEqtSkmzRZfpkaeRDdviY5Lwa33so5WohL0iS8PizgYuecZcDOLfTNR4xuU7
YBOv8uArhHqZnbWv7/MBLoEfY2+VnQDDpBU3wBUGnvP3fheyNQoMDmcRy6/U
iNV3ngdQazrGeuWQcRZjF+ulDbA3TSQPjPuXBaychfVLOL2zbPFJQhU1jTWw
k90bvnBRBPYtQT58HcbHkHlb7Iq60G4GHfugv6d4N2G3RA7FCZDT923jxeOa
agiyRintC/9cXzVdBUZMheLtzoVfDYCbj8zWemsnvw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sm7an70PS4V/6fZnNqMYfhnSvGjDo9POsi+eDh6JKOJOY9IsUCVJpmO3oX3J
E0sF6Dovq7BKzAWKWR1ENW07n7DzGCK0kPR+qWSkofqsyQcZg4pgQnuSSHSk
hdt3gPQNITjHcYHgbosDGAgiz8rc3V5g4wfcHx1J0t0zhTaBU3aMVOAiMEXK
SMytGASxilBnkNmeUvbpsz63JFBZQ6nCiFQ2NKwSoq25nu0IWMsjlY63Al7/
5mYdxZaOW3sdiDn6eWnBuAh6u+qaDP7fbAMx6v0Aj+tt78Mr9AICKEKtFK9d
OZHEcGFQhK/YbolJFpSinEc8N4Cdp0jJp4kgYZcU9A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cIiihcKzwMGNWXY4wdmRlHgLULqYZRC1AcVLRrRnxuxrC+ZJfLh+dKcaLjV4
vsYQ7l0bSTYbC1j6AyWGQZPjyhfwJlwk3tWJFhT3YjO8LwiVmfCISQXVY5vq
qx9la0FIbLGya0oY2+4mNDYjOaMBVb6Z9cmeI9+I1kYCsMkSSaz42mbuGHfV
i+LdXa51ar7QGIyqfeKgGs7lrjo0e6e/yHiNpSF0lrcJJNvdJLXVzXaUQo9K
uFdymT44IfxAVwd3iYX9POA2T+b+Pp+QtI7r0VyD3udJKnKjIwVVlmm1IVJ7
3ghiGq+RfrDCSx42Ggizqg0mop3ZDhYOl0iCGAjyPA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eg4EU+oVVh0XN7wlBC2C0lfe8uFA0dINhlku3NJfR+jD7KcJVlCGPOXVvySw
PupVd96lWKzxyq8zo0hTYdv6ovaxm4bhxCYRM4ygpuq/o/bExEkqrrwAs116
/G1Kb/ZzHz1WULoJYg4/7VdtiFN/AnLgpPP1C7bfribxddwyRzY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
l8SL7vKKLj0TrGffeJ27gkb13UaPT6ad8vYsIpi7lqrZXz69AY5Z8TfKJTpt
IESSIT3mbN95TT3KDlUW4UnapmCuNoXzOOZFrdSxz5jQITYvx2Ix3k+udtkz
/BlzXJ+/UY1rux3c6Qa6y7xMi1oIozjI9bedZEdjYHK7ebgH/FmFmXBVJOBC
EV/PJjx4MyZt4hu7YsFaa7sVEPUiRi68azVfk+yJhNk2PfQ6bsHgr19iI0cK
jrfqLM1qTHKTyaGSjZn620pgA0Tqo6jb5lBA6DfyLClXNzCWX9UmniehZ0jx
8eyZ9fq6Iv3QcU8NXyJ4gvxCOKnNjd4a/xz6HUOGVolk7D48n/XIjsXkU9gm
qn76vpRM8yLt3wph/pJLehoiHdrZQgZO8bIceFOdXqCU0pfx1YjWfh3Ch6tv
1WjCNF79DNKLBblLpBaGMKOB26pouRkjx4+7RKe6UC/lHiH16BXE4oZAhLDt
6OciF7+mK98T9iH6FgDCVIG249laKjzr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d4K7QAdiWTCg+B+K8/pPG5vvSjNNTRSfDfG3jIvw12Z4zS5mhPhlhPEirhnw
qjIdrMdcySg7hLfDP6Q5BvBDsOcdZhVlQLyl8rjxVO7J9VT5UHfRVCbDt0sf
zfMlo+lywUIcVU1M2zsPZtA1dgfeN83a4Ce9NL+6fr2Q/7cu0M8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OA65ICoGPkbKu78cAigUZCM4WHju6wuOYvvFB6OqwNCdBtZRH7Ny4e7t7iOJ
WRPDcuY47Ve+Q9Uzf9mKilRtHvVOpM7JkBuMqdF9QOevpKIeNtKkBNhBDPS8
sjYs1EbJpFe64n8+0QuHFl5P2nNkcG9MF++7j39eKW9707AYNos=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21920)
`pragma protect data_block
11Q+buioE46Z3Ghv8jt2ijKvZswgLTr+sCbZXlKy+9KMuKwfeMHSrxNZRssd
eqAgxc840Yb2W8FtfYXuPM8gMMa6ODwCvcbZstT4QBm50mA7P1JIBNxc9MqA
CtozlA9/oSq1GDiCKC3rVxDlfLu4iIREkzDHURR1zxdc/1/EAEbKqvBdq4HB
LzoQO/RWadaWsNZthHkrelezpwBpVaHUNQbDzrm2HL4s9ElGEnTFUi0p6M9f
seNWumzw922I0bFpvTbLKGySzqfFMHzd0COhfqE1HyZTxh6BLOIcsxTgQrt4
78hTaoObVZ91MxBSgpNw1+gc7l7K2G0SKoJCtpEVgbn3F8VaLzt1jDFJ4D/E
miTUkXteRk/PWyVNSeQicvs7JJCFygEulvwWOz4mB9EhRG+Eq/nbMx20E7vC
6Ak9TWx1F9pjECVzKpLAZOT8kj7ezLSpiTguwETiac+VN31cBLCS3FmH9P9F
Ecvr12qFRsRcltJzOPYLCoAzXf9c462E5F2AhTqGL8DbLAcwEzdXw3tLvJQH
1zReYfrwUH8opNYCK2Q/9Yi35xDBqLoyN6HLcYxwC9SrQ/5LLHSwfzjKGlHv
+cFrjE8kbcsQ4fw/o6XA0+sAWSXKPypFvKk28kw44o4kBlwa+GxdZiofqA+q
boBVgWelMM/rIjtEK6K279tUFOZ0HbpLbwVF7ggdVXnobyi0PUXhVm10NLiU
33sR0OIb7vTXcVZSKJHq2a2z5aUgGU+aJwl9rDfFwcc1EndnHdQjFIXWPjSU
g96IUqTV0YawlnPi0WIMMqL6q3c3xlmFlPdnMrRwrrAVPyn1yKTwaYvqNto6
pJd/RVYP73MfSGbxbBl+ZbE0u07PRUMviOItc65gXcRwroLniZcfU7CV1xE+
biEEs2Fa7MdhZ7WvZvNLet2IpjcFpgdisiOq588C4I563MrxMgJFI/UbtOgj
8SiB6MwTt9AY09K1Q/TxGPwjeTwkTtFGI4RbtbQzaAau0VkBkfg8/dCG8llS
AxL7wWo3bezMQiSCVtRB8iyCl/9C/Oo3vW6obXVnL0s3Y0fgchmawRXxrlj8
98VeFeoYokQqOlpEIpszkyLQOUTI7iB052mSdiu5SwxCBnxH50H5baau4QuD
ERMZWZcOMiFoFCKDLVBIbFupiujyDSZmK5Q8B4+TBYf5SeCFP2BAsuQEO5x1
n4SY66Do83PDMSlGlNWLPxbGfkIMeLpVcoONWAh0DxGTS6uvwX9wrFUJ5x1/
NqkCtLubY4DjXZAoIyX1wUEU7+XCktg8A7EYPx2/MBuQLin+QsuDwxjbpI5H
ckPj38O5cHftGgkUxNqmZBRzCgrr943SlfhmmsFYQ2FF2FQWNy9DUyaULnq2
nDYAcRPK9X+qht6N4JPXahu2Vut4X+8HuDnB0oqGTW2B2BlKK/R9RMQnQ3gm
RYWdkvrbjcf0/t0MhBS78EnJaJncDrC5CK2+qOCNdtKxw/nCsp2jgp14O0YQ
W7JxtsmWWgZUs+6Lt5chp8Rj1uIpeGhITp9gej7syl0rUE5ftgLWXxCruMTt
cVe7VGYe0LiUURTQPUZbybEWG9fhFOUcIaPBTxCQ7IOMG+dVPMBdDHVioQL4
PX4oE94NaYPfh0EmSV17Svp/cr1zqVxCZyflDUw5qHYAKY52pOx3w4CtaORm
SL5W0cCfq9thZKDWDU8cBflHZ5Hh0vX6TYapFQGZ0oCozl4OCJDg3ugv3MDL
bX7r+ickPlKI8MeJgW5I1zA3OCPiY0QDKSC6/QGpz9Af/6MiTBASU1yny5rs
3H7ESurnsXEwGUiO5cr/pmO3IunQIHNzXpv+sFV2RxD3NCXv8t69qg6Eq9el
HdcZX8fUd0+f+nB9hn5mkY1XlWxxRMMKqhMsTW4LOz4JR/jP4toiXgbddpft
3LZIR263/UYtdqwdkyJvRlq947OLovC7rG4TlQLZm6g1F5HM5OCHIiD2nt55
83JbC318ore0f9sY/j5pRKVVMOjGaYhm6+rFi1myiEDKpqxooXWpSL+lX+MX
AZIQJ3hmNshvkztsng18tF7NuDckK5lG375cDCZv5fEmVn20DG/oEvle30Em
gfZsMIbGIvdMcHkwe2bVGXrlvH1YirOSIRVqipLZQy8cCDrBDwR1kIfRyxwA
GLhsFuHtBTsE3kSJPZ5ygqkwAfJYn43JOOwlG6KtRtqLfd9A1ijOxYH6seDu
5RkmXf7HHzm107mkOeSW3tPd0YEjrm+C3fUecpn3mC6s4N2XOQhcVZ0NyTcN
+jIFiNlCzKHI0hRi+bZVrCCX8+SWIEXfnM47LRB1BIEZH1KhnoJzv22UgVIT
7Zpnv/QfkdsVZVgkLitjtg2bnuS+kXpkw7EfKUSbCZdunNVrZWnfmTE7b0od
AUfcXZ21ZlJhEubphMYQl4kWv5vFnhybvqD60EyHJfvkqnrSJCoxlgIJRTqm
OPsdfnTxW2Cd6ZdGmlN1U0WPcBRWGFyy0rce4EUrXTKMZHq+0eltNbUu2lCc
2t4MnVOgRhj1/XxrW0AcsOEYd5IIMzp67HZuvum4EtsJOfBEH0X219gC761f
QmIQaq/FnAXaux5Wp1fiDbyAfmpNdpSdXH1gHJslbQAxLtWPBqAFl3eV2JyH
nJt24HxWL2xFrpe6JXuI41NJIsw0hNIYxPRebqv5ArFPwzaBsNUvIMaFN5SF
/rbL6LwIUkho47XGK+cTJ4M3W6wouqR5ncmlZ4aa6rQos4E+SPoZXtQ4MvYV
nqcj0ohx8+EUTxUipI+WIclyR6KgfZR9yx1bud+XcblNeHzIaBEGs7csZe/m
gVq1gKXIwrmRET7C+8X6+YYiX8byjwLQB996ljAWyLwLDzaDdXx8BmmZPHRI
gf/qmpUYAtiS53Eorj+CIQWD3TTj//03wBxP9etECUczOFIthOhAplWoCxEl
JfZKG6Ekynef/rgeiqsnFlLXOuWWKyEEH3VfPlvk016u30hoS4XrJg0RCHh8
4vIPgXZnzC60PDqd7YwSFK53wPBQ3Hy5/4S6o3ZelT1gAHF/xKhbtBbouW/q
UnoqXUuGQhdRc5fnnWs2BzUcP1qX9/529heqwKyGFpDhUt68TfVRycwxwzZx
SJNJFtTy51c9o6HpHY1O6pvJKlCj3Ku86Na9U+6UCwEWCAdWCuTGaroXIkPj
o8d8Ay3PbSHEhDjAk6NnnJlreG7/nQwidSgLCzPNP1OoxeYLSzmcuqjLZuY1
7od0YrtviVN2Q2guuJgPAXIam2ox8QYUhhEMy1oY2HwYNUuHyntkzknN/Xjc
hNaQlcvOc5Y4ksjf1KTw7NVb0ILXgD10R34Fn0VmjNgO7kjCnZuWEOL1CMdL
ZVJDGgZSbmavbdHxk6pZyvxnVPyAOQofYpl/Aa4s+AtdWr0AGfzzrPFjWSKt
5ezQXntHquJImWvE5aV2jVZxTfXo15wCYaKhbLZ80rjS69KUA81uORHAhJym
UVkxxBU4Mz0XJAdZwo7ZLDQemN79PhzHt6GD9lMsyMKPvzLTCzrK0h4+wLv5
C/tz04XRP1jqB3HMg3Q/PvXVoWLnmnosPHjoSn/PTFjXHOO/mBl1iUiyPy4e
q1usYx8T6IZ9ugb4RoGZT3zYbD7NRju4OFXNvcDRvZeQL00nahcS05Vqcg8K
nGPZfxdGPsTIG4ZqoR1PPjRdTzAeJ7fdxYipmVqIFUIBG2OyBNC5nTYdHhhK
6TUOz4hTwNlLIEoyK1IZ4rH/7wg1AVioVtHF8UiY5SXMOr4p5gEc5AL2GwR5
bpV9eIa1jal+aVD/o892/CEPS9kvmFDRW/OHv3y71OpBXktYWpsIVtoAx/0w
MibiPL2T/G/vV6lMUxu2i++7r2FQSniKjFoEchia+Mi1k8AwnQe9IFJEj/K1
Q6YgKjAwPGwXMp9d45xnWBVfTTnzYjzA4ZrCMhSrjCUzLk42oDhG4gujGJpl
tqaXbGr7Hxe/wWCigTUB6m7qimgF8JUoSkYABCKrefnAUw+CuJc3Ln6cteGW
YSzMO+iMJdd0+LswxZgd0KhwavNIq0gHf8m7Vv7b8BwKmVuT2to/j0B91fOR
KDdtyHw8lgO9XWErvB6p+3zPlMZa+y63zx4b5tvt09lnER9MP8gISYWElXaD
2VVzynpsoBH7VBiAo5bhOyLpE/Ku7Q7gyhM+jyjax4kHhDyNufYEPjpUbgEy
Fxw4gamqzMNM3CNiY3jkX2ygxdFW+2Jb0uxpNIdakJBZZdUw7GSmpgz0Ao1L
R1GHUXnqswVpYWmspIIdS+JRZr5lnZ4LhGD4CmeEu5O5hD2Hp87yt7KB4Yrk
LGGnpFcOSnxhBLDLWwdHWtm1IxcL1U9f1uRqlC4by5pDFFxtbI4I5hTlFEzv
8dUwPG2DtjHQNRjXw7JisbJ6bbL3osHg1YQgujugfK2zyikYHH1+ixX+2b3P
39qTjMprEmmdL84vy+h2C+7LeowF6JeinfzA7y9rmjYsrgJn96EV/oe+IgxH
zWmq+VKRb49V3awcsY5GPL/wRsJwDsGXm/OPPlzvfulVWUgzB8G6R2Ik6hkT
Z2GJQlTMNEkO/tTf0iH8bAEMYR3BDnGXflF8rA0TUvW7Ja2WleLeN753xMnL
Wk7+Ym5zlTHlA72hNfPt4GncSVZEP3fzT2fGEkiOa8E0kJbPylSvC9dqU28R
Iu4xaxohenvRLF8rfwk0NJxapISjjLeE6KXho3j7ulkK5+uMFi7NQdkOWZ4b
gBmsIXr6EJOktQY3QPODTnhshAF19orvA8MIeKurZIzsB0wSIgVQlh/WHUf0
UBNIPLrydjqmAKbSJobluf2wU3sDE8P0qa/ukxFBLlTBTKFehEaitXxrpglo
WlSzhcyqYDxdYOf5aoqrsgD0MEMnX2ntNacZ8/0Wl5OCN+tu0TwBJLQ+wFon
doycSM0qr6lXNjarfotgc3JSksQcRREa/7HJ1pmfXv/WZV49RNasmRNps7od
JbIVjfLioFGUU8/1e5TxuSZIlTkJ/Y3uy9w4wjbqtHS3l2Xh18Zx3E7uQQRA
6qZT1Jtsq6gI1s6oukoWnXaLlzHelJiSvEn9wIUDaTwuOttVitXSL8gOyVd8
s/3l5zz7/iNyCGsOaZBD3rvOqbePY+YUJS1ZV/Lqs4chT5yYYqEni9uIEV/s
X9l8aVOW3VttLq/hlpqbUg1TvzWH2tFmlvvnuUwPxHTb7FGfk+nZJFZbJWbv
S27IlWpNG1jXaZOUmmUDqKCjH6YJn5BZNAOtWmqecrsfif4g1ZiHqDWLZvg8
9hn9+zheQN0f31VUP0c2I5yro9iCnj5DcyuytwuBZ3zpyM6gSQLglDh0Ehx5
tHRtuTVXl5MAM6aeNGYj07X1snWRvf1ZD540rSeCWoxXcCODqofa5p4c5WFK
75hEQQIyeHBX57ZiUEh8AnJTYuyOoikRjUJ80U3IYJ+1t+0T3UuVSFOWJiuo
0BEK1Nt0Kb5OLNUuveMvTEX/bpyG5ovSw5wcFIHxzSA9uw5xl8SHhRZNXjbS
MAjqF/xC805lLUUuBI/iBiSRxKdhAzlYLfkB1HsxubIMJZ9nLChpCyXmOgM7
MFx//0UXiw2P6dbr9aFdg+FyoBhgK3Xk3LEsKR2EfSqDoemChSx6pewipjPW
CTgmwBWKe6wyyD9zPNVZpiGe9MmU72pEGM+iOgVjuzf934VMzJeh1RkHjE1u
Cg6bQFf56H+WV1Se/mC/qMmMkqZvNmk+jJBZbWArZYPZibYOuFXagDw1lvbG
p6WWb8RMmjGdKbq3SedeCIlvWUGEKRbTHBumIycM4BQ7FOTurfGLz2A+ln8b
C/GJQokuBYBxF1QdSjWQZ56UX6iUXghDJGYKyLUKmoeADsFBPDmIEuPlxLIu
jmwjEEHhitcbTyM0BwMryZSDEyd2rUVwQIpAyWgouH2Qq0bByMG8TAfZF7B6
59AdZR5VtcVbAyZqVGtp60qtNgNZkI8vUFJkxUFEIUIakZUas9Di8xcJ532l
9bYUmCKzd1mzgZQ4zMYsjpWRbQY79YCTwDgBXKFXqcs74hsGklWoQXq8Mz0B
te0Vxr7XzK/zL+4FQAThklILqJc+Xy8lYU2wwUsrwmGGnXpUAktZkg0TNVp9
nn9rJqACM3yzQidJVbMNkw0uGeWirqmTyiBFDUjJOvhCSgcGL6tzbSaKm4R0
4XZwVy3OoNEtqmeZ2Xim+sJNir329gKFUZ2GiWhVwBzyN5NbsvDO5kfV3OL4
ZFYDnTWjibs24re3+n7x40JE/4yhuepjGmH9eTvb4EVJ4jXLQ5DAIBMa6K/9
vRL5bW6yBxtiowE56HWRK4UbHhQ4urBc8m+o1CVaxY9oEGyq4jnLv2VnO0AM
iZcSArj5rLt8b+ir8cEd20ftEz9HbO/C8w4S+Tszg9Ls+LbXtlK0g3KGLARi
Oc1aoMt0noOEnZjClGOmZ5J3ZyCkrVIufptSk/VkRb7MuCNUifMKLWMogoSq
uTrach5kQ95sECqvupbdHi0ScitTlHhImvSt6iuy/OsepSeZm8RtZdvfWNyN
OjjtH1H8FErzB+LNAM3A+KQYRNp3MZisYvaKJTy9U82E4PcI7+o+3IbD6cmK
mVurXO90x8QpFQqmOMvcmfWMQISKetyZCw8O8hGUk460ocXH+ukyTlILDvNj
QViF85HfEfjZzdjrySPHFRJMicAl2hQ1Wc/MfSyqO9E/7QOdxd7fqcEXrK5x
0VTc+CpmD9SmGlNd0FVEmZW/RSWljaZCbdhuTYr6AUOjt3dekAhjn0cbd7M0
+y+3NB+SYBn0U13wHvyMoF+Zp5UZrX6jBUxy6iT8WdNyAUracE5MF3q6fIU8
bgD8bhFNp0f2tjl8MfYcgewoAI6b1qXhhwwObKJnQizSAFuYfZKjmZ3+dN+U
K2k6NlMweWS27FbaYr3bwnJ35m4BkbcIhLpHEUGpqRaLzZaxi5iWixxK5B8d
23LaWslZWcbGR5Kt0wO17Zgs4XAlNhch4GtDdbcqwu9QC+daIbon4uMgEpe6
P3LAH8qIzU9HGkFsp32AaVCwV1QR3bYQkf+HC87ExZZn3Pg3FZrfBtkm4e8B
HYeDAkf/VwUgNMxijT3Q/Z1f+bN1IIP6BqlBx2UWX5CspHSA3FB+mGRoqWWN
3WU6mc87eJrGhiI5Kn1tutD04TvPDCzKMpsuxvjtYqiO3NItvtOB5kFYSrC1
l5ITsuFAlbxmWIS4wJNVkdmPLgq3PUtJOlPH80HacLfsjwu6TnzjNB0Xg2IS
p6xayU1/t9qddoe5+rnoBZ0tWzRBR8hBVn1rvfBeJNaJAdkQUnp9Snt6qz1K
3IhByKASCOU1Us9lDJaRMhmJXBzp1wyif3+HRyBLWk5JETL9ygmsU6B62X02
GhRg+pXbd8g81L1iiO1i5O9YUk6pi6pvEtBUHwBKp8qWPSary3KZ8PeWL+bC
CM8rEKcUZSRz/dOfN6y6yZB4ZbqlkkTyMc2jNE8FOQFKWxQzX4chi6/QEVE2
t6Luo7lax6iQLHiZiiSKl4fe8iG0SA4X6asBuagaMy9E73B09GBrmNwFibgK
XX+6QSdjRXL1SLYsP3GPKBza+3xSIr53roHaoh0iHGho//nCTnTaeukq3TES
fk7wD9WJS+iKBLmQ+EDAyJ286t3mRqJRHWKEjmCo+Xy4SprlRu789THBUOCs
/Sze16raY6vbvKEwp22IisKDCT1htodmZOQ5Q5qx904hJIHxMMbDn5Jk8a8N
typ2hrZXZyZWW0A27lXEPDponAUcznhQ0RXaz1vXa2ypg7NWm+gpp4TZ0QZv
sNXPbwUFRlEPECRRbyj4GbZFjp1T7zT6VjZQkl6hMn5u6y16v+fziGSKOeA6
OKQWrrSuK0NBTmCMxjgP4xSG1P2tqpQE9wGZ4rNzP2lwXZLsZyaSgVgIeUW1
O24W2I01c87+SVkq5FAvZlvWnrw/u1lNRYJX8R0R/1rRQt3jxMQPhq6QrPPK
scy9ltaxF3thpWt6TVEdMcC/gjvtzxgbNTbBj9jCjSUWPnnZjZEpa+dVGO8o
q6wNrJ5l/JQ22E9UVXDGyLUB8+InbA3Jfz4E7X8bKUuQY2QnBXjMzo+oC1f4
y1XpWtA4OOG8S6mf1iyDsRcLAQAx1Z60Z2O04aq35aCTtWtCaVrJnroJqiLO
uiPn5HCfP4OphWFoaTc4rlL8TYaBTPcVRDlJD9K3WK7BH9wXwqe1nbTmEl6r
Ka+9zqT7yr7mwghxdsLEEt6Hh6gbSa6LRb+OSyd1ixTB2+ISXbAHqZICwRjj
Jfzomh580mlqaH+2ZgL7KjNwJwkeVvL+3lq359bbA/l/LYD92u+7/8y2B1wq
IdRlllqTsuKHwzjBpGCQivBWXHxnMk/gDmyMlO8CwHJMo0A4HBC73dTLzaP5
rYGCbQKZa9SHf5Pl/5qYW8sPMYpVH7y2iFgrqK31YPKf9q6TM7/IlNPmUfVX
SQBuXTHlLJ0IABJAz9FAftveanxSK1a0g5zCOFkGmQhs3syW35Ky9bSNJ7r4
uwCoiiupV6zKWk5emdFgVF1ZMxWzaC3xBDUpLFcz5kP6S/OBoV2oXlZlcVSb
Y0XTNAsOdudK2C+8gORJVaNUhDNReS25vrsdjn2qhId1sNBTfsoTKZ1/ijxz
O5ik0jZfNTog4zrC3V+zFtlt30GjxvfusheoiLuNuBa61EBwjtn7m8DSGPYs
+N7qZGkPyu2K069QcUk73OzvHbXdLz843C7YVoByFvbrURaktEl9Gjo3EA88
bJyKDMLcbsvd+TEbXyRnJagiXkNtjW/84cZ+Z9S/UcnULUhX93fVRx30X8JC
M5tc8BLsRwq+wOeEicDT9IfcEvcazZIDQ76IuCvnw7bAGEkZUDXxVPzs9ErQ
0pUZJM4xedyl9XtBgtrXBYsqXz3QB4BZhl3uZdo907xCqqHNrjsTmFaiwQls
hVvrv42+IFiglDB6ogHUJIiUwbCiDm8YlEoPWCEkgCiiE4DC4LXUKaROjXn8
ltq4I6qJGG0NzaPaqR9WUpFR6EhiUuRnO8pDJprg5IodRubIy+kKsoXO0zAt
Y0jCETK5hcQfkh8KzkvoT0TlQZjSKhF2FfYIvkPKb6JTUEBvKJ2GQj4W2ELQ
bAkQvFKhRZ2fCP4xnRPRcpRH0oXtikP/z6Wjz+Nzsrw/h9kzXEf6DTsZ6FwF
+EHGQyzszwpMlKri6zGovSIa9y42zOqZFcQOUbzFUiXMO4z4dK8GQvAdXKQ2
wACoy+15l8l86+ND2vo6uZyq7YA+pZtOyzvyXubW/oPEBR42hNE2Wykt1Z5I
CpaLyLTdLNk0tXHSL+8AhoHWSecqHOtgYtgVodq2EQv/Pasxm0O7f2YFngs9
Q4zmhmS2yW5mF00Iwujyp7Cr27cvWpzSOZ9HpTEKHlCxT3264HNDhigfvv8A
Rm8VKIwurkmvHS5KVhPR5S3fkdteUibccbY7f8nlcU7VWR1x+UIpreJSVZZd
A8BU2gRNfpGxQ8y6IECpsOskmdT1uq3MwTJv1c6ge5CPRjLKUjjIWC1m+Nf2
gyqYSlduPtNwM3hkL2iJKcr7ZUMagRVqhxZ35jehvsWxzeFAD2l/s/6RAMQf
hu9tzQTdnMAnZMADTz5WgJ2sB/wEFEFafsN7OishiixfPZ1iWvpHvZcjD9bn
O7z4v6kXPVgvmGctoX9bIKN9isJJPJq06Dv/x/Ngg8A3M47O1zba2clW/Mi+
fq4DnNGy+2f131nmBThBmzF1i/0HlLAfnOUL3cOtyZnmAVAmcDwY8K3NJ0rg
RsPuLCB/MZCgpFSBxBo3WartQ+aiOd837C4bGkLD7QJbPOBSo2kqOCxBe1R6
mJb7O92vYXLbBlV8Hep7DJeTYcexzp1jwTZUEPk+0fvuL5yzMkh6zTtgsFbK
jeXnh8krbDNyXl7UDQ9KNd5QJXUToZnay73i0NothOq9HvPA4N3+PdCXMTHL
j1UxV7QC9rMOHD473OBO1hojKWer+CwdJFOku3HN9Jc6lR71NjTclQUjZTSY
MFR8plzYsxUDqkCB7YfOgB48UsXMMTlF3RlyPGiTa+fiS0r+gn7hYpspXuyb
rGQNJHZqdDQTUzzY/GxQUAg/7fHwJsAhx7ZDesii8a451b+uuHQ9HCVu6itz
2hWwl8hPwagXn6i+pYmRlo4Cs4DncQyI0/yjY8LyVqn4XepSRwUNBYzY81Hf
qUgxduBeLUNlbLGh0r7Kb51Ou3wEOy6GXDdyYH1P6aq5V907yPB99cA8SlaU
Gf4Ij5WzdhiTsnEZDalhHyUFfLq6Kwp6RJCePn4YYjdE7Q8pR/QJBx8+6UFc
IJPT8awIS0bKYCacLJtCBrevvQ/de8SpcrUJVgY8aM3U+JbJO4iNC0xKk+8J
bG+khsnyJnr8CUsImntFaP+Y3nchJ3h9hrSjRHDYq3v0YEVBtpHrjjOZ38NP
JteAOajeI/SAanLPEg3S2hWhWmsa8/QqoKSNyTQzPrKa9NHWdknNOmcMuO1z
MXshlI76tAezuz2PQ3q15YOo3uiQ88jMZnebuVHNF4HqMwSE+GKfdWzDEmBm
J/fptHIMPwhwXPYEdIdXNKkSBn6pDf8BmDDCTVSgsWR40/NG/V90m+GLYo0j
7VH6yFT14ZmxwScbYgobFaZZicQPl1cUN7vRV1xo4oohgG9u8FbaAk+7azP7
AMUVhPAbebX7g9gv87d8mgsCF27nmg7EtUZFYk4Hr58Mg+ikH8v70Gheei+e
18FELqNY9Jv0ZgFHB4QjLd2lVZrBlliup488uff7qTfxf7HSratEkhO/YlDm
T4vQyhC8zK4KM08gk40s2PUDoBTp9/Az6h3g262m0ascBf1sa8FgcJEFUJdk
ac98o1pq0cDBeZwBf/ZWTG/rDbqDkY0PbRF5MJ5v2Pt6geKpIIpgROohkSTf
hEj4Gjk+DuXPNDIsptey8ibap/ARJzqAex2N6m6FiaGzQKDS7U5bdp77UnXP
je+0rNlydhdagbVVTtXrT5/VhnWIdaXuUpqAxwMVDT16Ly7SF2CiXAGvjig0
xJRkyY4HY5rsznbaBVTYc27Ss4xBuRgrbwKWF1NiLQk+07Xl0eXhxRwINAKX
UBNP6fnvf5wqi3zSxZc1D8j83kPGe9XPJ4kWYrXbOJhqQI2gKP55DxeEV9Nn
mIjeuW+RHi/iFzxAUuIcZFNLJ705EbzOkfwxuRcA3aR/ho2y/VcaL2XgjyjB
yixR4OXgIkLNlLDgEs+V05iKi3ow5DiF9NnBosXyaYZ0YvzLp3d03eH5bAy/
HevB4jvSSB2MARdiGCFlD7P5XXo0mu7d/Rlwqg+BF8mZ68oKpjWeZGy7ZonT
qZ8jgQJWyzXi3otffXwShA9wgET0y9d9RdWWU4g3N4oNrd2SgY7+wyIxvdxJ
ECm7JYwCteKhUyBnX/j907kybnIi3oO0jQVflMiMJumUXR9szgyCn7i4i0x9
3tUQ7J5uvhMD1KL7YpaL5gtGyAllqcLnrWXvQmyomDL+kqDQ1sk+i1cIPkHl
fn/0iVe3z+OUxN8cSBXCJCs2n0Te9KSS76hFMyE8q0PR6MibwwcNAEkhFapz
WbTfxh1pIOG1h8CG3Y9uoh/fAvDL/wdCaVibZk3xuaSF/KRBXThgKiSmh81L
qQwXK3Bv2y4CrBLhi2iDd6/6U7SfDGVl94clG1687+qAv3j0zHiXwFS1ICpn
se89/N9UuGBhUJEu80XzBJGniW0hlTS2eZxY/AzX9CguhbYciAUR5XOJbidL
RWadYRQqn5X7vXpotkmDIBlOzlrlxxA7IR8zI3VvJTRw7C/uzJpGUqvwZYL3
0fUM1qxI6vN5bLrcxyyJXM8ZT8scS1+TQxSXtPo6W6jeabA4GjvwAYaZ8l9x
eenVjuOZSJn2jtEXvYHzJcXpn21yIFEoay+5X7ZY0F7zDiwSJ/P2XifjkLXv
9KL7eago/rvkdW8xOtZotehNi8aQ8cPeZMdnGy6HSDntekUtJlgLCy1JLxVn
NDeRBVHYSviMaGmA/ef7ReOUtKVJV8LE7VvEiGGJWS/kOkqYr5jKr7AdPqHb
coRqhx0rfq/xOVZIKI4oUyaaCvcdHGtQxWwmNr3ahsQtUq59iaKZZF2RuUu7
ZApcOWwlCmxX4W8uXvSE6B4CPG4tuV49+yIKmEqOk4HXT9+ucZJFlTIL2/49
0CeYPDvqIqb54cJpdNzdKu/HeAvXKPrR6mhwQiV8IeyAQ8TVhW6rjUJ5LD6a
W27bjbWYi1rSoCnfYKEEMKQSULhiXdR9K3gCk0C9aZcnmlcK+U4GGwJ/Or3R
9lobp3qGC0pOlyFJiZBx46I3neXyDul/6Ovxvlkw3MjTS/lqIadryVkN9KhS
mK1mb/YkLsAw6gFINsbm0KhD5h2mIOZTABULoSo9M5G9jLR9Rh+v0I5ZbC74
nZ1B2HuIZPNcjbUpU9z9NDSbJoEaMoEVrrWsLWcI8n08Jfx5l8n+GnDDvIRF
jLknzeb1VSLnQUYMAdktqiBqM83lbg1EkyOH6E3McXyOfl3qEm875P7Rfd49
MldqyQfGeOcp2SVHRtmFYbPkoHH1IAJ4lzjnm0bFTPCjwM6HqQQOrma9Vf8m
WLg/QXnc2mVsOw6Ebid3YA6fFHfowUzPYZ8WB365+kClPlI4/+1YUb4XrAaw
perW7MoIXwOnh81DHYRSEnSdb2Jg4I+xhV7B8BzZDMxLVfcEnb9U6cgB76cN
8+9+1DJSe+oVLovJSc/nKxzIrecX52jbuBLvYgrkSGUowchEuhmaAgnZuZFC
8VD+Jvf4tAau3K3WkQgVKVS3qxipRYB2QaDfeThj+kg/jQ6xRWdo2ftbZH75
9JleYq0EejzLc5Ee5udd39w5lBpr0vOk13s0pTLo7aZTjHrn26YEwYYrxJne
D06x5WoADAIH6qf8nkyL6SKE+qz17XeY7rp/8dKATUUg9rSR9Kf7fY3hK6Mu
F1+CQkQHxyhxk0HAjrHd4BA9UHHqDJSx5ir2n2AYCbuEXDtEn96PFluXxG19
Vhs2TeGAHUroCN1ncPUcsLV0JyKGgTP7gn1ZmSQXjCO5iklQ25yJpU5zmASg
FGuovC3zj6v3pfREd/vQnwS+EJ/d3WZy/ux2omHazTofkkML4Ub1CN2LcvWt
rxCqVQWOLOl1sBd8ZexLk4+KtTPHsy0ZMGGvk5xwEA4N2KJSMlo5QLgDTz5E
LByaj4M49slwdFQfcKNx/LG53kqYcB0aFZIqmEQfP9tZAIiUmqPUWKkpoG0W
W2SeWjYB6QS2pxipaUzsGUSwv2EMrloKf5KI8Nb/BFs+iXBgUGY4AeyrjQx/
VjYJZuYkAt6OsY7IgW7e1+XGTqU3uOrH5BeKThmI2VLp0g59dziIVZSoTUE6
TsMDvgX8lfgVpI2W8E5D7qB8FCwj0HoL4eLtTrzNhW3FEeg7uZ6HTUdesNOK
nBb7LfwKMHOyhwFl0nyEY661u+mDKJmW2/2Zb4PjQh6LI2NW6gXccRWnWnmD
mGkPcyZ2npQlfHoc2TEz1nh3oOfShzoo+S3WwU/7AY3P98jobtFRgY4yUxLY
PfwS2k/X554bbRSPzWMNV4nRiEZ7/61cRXPamt3tp/5QnXcXJMRlVvLZUaZy
LPD4FrBRCp5a8z44CksgY2SqgM+Rl20T/Xx9k96R0VWpAAkPrFVvF/+8aC5m
3n73EucL9ZhnU/LNmDs1tobn8R6vTZ0xgaHSk+1V36C/kDtA5CbDfp7b9ImD
Gq0VvWo+tnqU5Jb//1D9uQX+XDxiu5pSZ+me8hbGCDK0J5cn968HcFVU/pxr
oQbo7ooseWu81Oifno3bWncX3j1U6D8xG7BIMpyUrqRAnDtKhV3+/9De97o7
oMyk/McGTRrjGhZ/uGJud4AY6CxeLj1jU4KouXQUQdY5SLLbQSJhgLer99Lf
mDbeN1Zf3WukuJYTf5r89Fnpjdyz0EWz1HBsTsoCpgHNSlyIQttRUclv5ge+
VkMpwCAYa6Tw6CIztNYtpC+24cKrvFAbBXdf5BLOjeBnJEpO7c79LRo0DnLR
wEsI4N6edWupR1nK2ewf1wKwI4eVA+g8dvQQQ1dS7wDG+ZfyiAmiNGy4w6AE
Ichv2wTh8w/iuFblOw3sDZvpoFRPUZzV9ywGwwbKanCABPGxXdYsVF7MlC4n
0ieWOJ08R+hcjRyrPzhid5OdPIhw3yYVg5+R51mP+3oj+i7uY54VVc6JraWx
3iZzi9Om6ldUb8njNSEjki4jhuCnVOAzHJWf9mX3z0zGUrhw1l+B6PRB2lJ7
smqMesUvB899aYd5Y6tvduMfCY5pdB2qblNJOKxb+vjxYVVeudcgUr2MQKZm
BWr/UsYMiC/Tgp3adOr3I6qQ4sHUByk0iku+EwpruhsCqf5VJWTxgLEckUZu
TErXKGOhHcnSM3hwI8vKTMiIg3ZsSUkbsh0DTB4M82qmWhd9uD5oIg2zAYa2
j0uGCPIPPPQ+uWQDMLH40EwsGty2wVCf87+Orfu252+TUr555EmfK2zrHkdQ
qQOTDLaJ5+2opsS5x6wh6alo0XgnjZKYF2mqDxK4+Qu2UzVUeNo8QDR4qq4+
46wLvBreNcAgZXIQ6nHUiIrXdv6vHkWLJkzOx4KtBhgRRxygpIKqApQMjwXq
//pNxoCcAYeZpzn0AZqFGdwKSSuAbYUuQT3WLGF9C1mDhYxxFwu24mwKyUY5
kIjS2c4ZY0m2UounYl0vWgzPVrm6AFdZo8bzdRTtpucvO2fFpjQP5aWC7+Eu
fxYBcfM/NpLCjQcj6X2ErB6im1FDheUq6ed7EjyDmN/u+iGaNEMLqMY8kBst
BOp1drUv3gU+ESaMnep4eZCnjJztT1tKl+JBAfPv6DkNqpcMwAR4POo5fcEP
nmOhZmzrGLL07oiAdfRyG4FvxMHdaYHnN2pIMaM8XvIkH6muWiAuSV56ABRp
QCqap1dQ3j0/AFV6lE0BwF0p+Tiq+4vv6HffPh7RPiLdbkxsEjvkH9YB4/ZD
ri+lZlkrsB93xjMu8NKCOuhgS1J+BIdSfA2xrqmZdfNpNbfIBBV983yAp++1
F/gd5x2dQeJ8hjfsNkjD8WR+PXcdZ9iwmBqiSDZrB+GWeNfMTl+RrTUBOVXM
NLTRlIHs//EsGpJnr37jN2b33HuKG0qLaOZlyHQuwBMTyP2BzsN1josOc4zo
2f3x11dLb1htBEriK48Zgp3l3Q/wby3SVayu5PR5W6/UE0ZBcmvG072UXeaN
pQx4rN8Hibr//cOBIJtdRjqmWjvy36kD/dgRGrvp3CiVfq8V0BX6MGtQm5fM
lJM8pVH0FLftFQ+okqddLU+M9fQ/GMsy9ToYLMrCvVXNx3HToZ7aYkM9dEog
0S7THjRVkZT86pWKRyIZcRLzm8LN9bsWAbPsgbUIdkjilatH/hhLf93uglav
/FT+s9NqxBrXoyaCJfenkMa4PeuFraZQtpcvgEm800MDtIZ56ro0VmfUnbch
Onx1BrJFoXtmCmv0nJX1jccWlO/U27g28kB71zLj7Sn0/8PUEQNOltgPrjfq
5hb8zif0+QjHancDwSI1NgvLRhhQ+XyVI4eDiHqik2D7MxPCGc66bM28w3ms
8N3C6TbandK8x6MP6paJ6ylOlHFAdEtThViBsyxtiwmf7NAqp/5+7DT5Kkzk
k5AyQn0hjrF9nzj6rilo6lUjug5n8R5dSMmxjVVF/aHz6cYDxMJi9sVhrd4p
wto3Ol6OoMf9YJ0JS5k4iCs3pBXJHGN7O67NQ4Ng3sWvzfFhO/6gWL/zNe9E
T/ebu+lXtjriystFJKRjAul9C8O2uceKNbBiUXuLlN8dAQw3c2T++ka/2Aiu
IA1mk5wfgNdTaDQV43bK6dWGnbDp26DwD3aEUXzwGoWI8Tjsul4ywN1YWZZg
Gd5Xl4jYBsavl5tbrzr65FAxLmuQM0D4xXWlqzBLw4J/BRgpjXjxNKWB0xiW
Tao+O/BZ+2gOJ01Xdp4HYGud1boUYqcKSdH//f5MYelJdDn3b/mgmC8gw4XT
c3N/1azL4EtqOh/9mU8G+bVmfVEsDBGTYc6FvBKnn4JVA1WOEPyCeEn9FsZj
F1WLK9Zx5uqgbbx870cxWkLjGDiFgOfvBylCFu5CYJt9FxWfpSGQeTMOmSMc
57G78OD/ahmkfL9aOOHnmgzsFhb+j3fRe2oYcXOhXyT7986NJsHYZZB//vjt
hhCx4UwwCxDV4fZaeKPKm2XDGrNhCgaarq+/BOJqjWYJhgzU88JWaDtVFnyp
DpS8HLE/YRe7bej4Hkw/Jo92MHo5EFTb6WgwnILcJhbNxl/qDEue2og0M2po
u1kEIhfoynEKEICRe11J1Y61p61i7riYsF78DFvwYinK8JimKoWZST8hg09s
CrIOr2Flj7L2DuPvbGuI86rY4yuMPoV45JW3C/v32moyMFvCJRNmkFX5mOu9
t7kg2Jw7gc2O7Rt6l28qzarON1cHo16hcZV7nGK2dL+EmuLyIC82UrT4XsTu
dlMjFD0YTD3/mpT5MSf/yXzPMotIaJCo+IdAfetMsNjvL4iAgjG3GArHhYED
i5WsgDbj2058ykK+xnapMOxh+Dpt97gjyOUrHzvGyMcDYsOjXs6+sUg+7Mg7
uEQp3jD9erVsXUdnK8jBZ1t9bQxXByEwZfUQHd0HFBt+b4fzsM1dVWv5zIxV
VE7uxzwnYeNOAJYIQLM8ETjix6tpAf7n88ErBz1PXK3jyuFFmrNttML9MJlf
3biUE7xNakIU/dBgBkSdmWastbYYHZT2J544MXc/P+Q7Xzz/tcxOw3jWGki8
rLD+wt/L5NZI/Dgxp4+VaYgsDKqSfajaLfz0fYycJ+yNqUk4JBjVAPVr5nHT
ky5sEvdNFrQaxYNCS/jikFJmB9mwIwS1o6R06roPV2ZXHnboInLKgGgPbQj3
W9256d+3Ygf55eFdD6YpBzwvXN5vtqv6vHVd8wOq+c20UekRm4Y/ix9foeH9
ySTApS/IFZKmc9AYlAviMMcbZGE4i1vLeg+0x6m0kNo2jpgDLfMdmD/EaDWY
ZHi8iBpS7TrfRE4Lu8poGzuCtfBA3gc0pAKF7uvaGrKniS9MJ2pwrE7wmpMu
aVHDkd4ean0enLctFz6fkkYwMkUh+s5oy2aKEpA3GhTkCNoSSlcY+xgLAjhR
wDbPhwLV5pos0cQOTMC8REkbvlAwIF9uXKpZxprJvinKF9e931c0k+0LpanN
FN2WZTkbX7dZFgt+JJ1JtIUBbwNfWcMjnik8l3SjhQ3oD5598vqAleX0m6ae
bJIhquab0W6gjOI9FRGt5Gn6X2Fh0gxam+rjzvQwLoqh9R1PHJrn1tq2d793
huORd2795BzLgd5dpHHEBMLqf1O60TuVOE3NV5i73UK+LuEC3tDgkmq66pF8
QX0oob2188EGLY403Z6hQS6dPJAUwJGRjCVgeAdrUSo8W5g8PgRUbNXz6zlh
6hPA6QfNXMWATKpglddrE8RJryEQmWQk6IrC13yGtbCpPvZvsOJmtm2P9Nob
aKXWep0GhD8171qPNbHlnajnLEbJel5qy4PDMxARfNEEdDMNQuirU66Z8RGe
1EiEw9n9A8LCTxL2LmmDISP/FcchqZTj9qF8yUjFvWmQoUeaIJbeuRxINftl
JeCYd7pE1P6K92NF88iYYE0QEQx2MdKrwRZz2dq1xNDO3hjIt0oLPpsdMJ3v
NwhSW71CqH0d5xjJVtYEhHWab4G2ahWKIzv1RJRmg2ybaEVvmsen+viJjQJj
IU+coPIJvdCDTMiaeskzU8Uo+0WK+iOG5JtJHOyc+ZacZ6iy/Eei/BDQgUUd
TURfVv+UCiva+6OVnHCfCDrn+sEVw2XUwpF168W9Mkf8QDu7jb8MTXeSWFQp
VEOBPbyZp2cGEBTB/DxXKecCbZUxmYi1qrN/Lza9VnWKoDQf267qtICKdEEP
QEGnfAFtxwYjxdidCNqI+tCazX6VNnnjjFSzRTvG/DatHJ+EKVRG091D8bff
F9WhHQRnGZ9ke+PHhyu8Fsff6ahVquZe5XouzAyybFS6teoYiqoMsF+ce6Xu
WDNLRF6AFdPv76QWQZCQaScnW/HZ736FTPGRBvln3AtHCdcN2MJnwL+szNyX
nk9/PhGgd4YXbfOrZrCtlEGL07tUFiooMDG/Bgyx2CfzJFEL3pOqWo7v7w4P
mx3dmGESpr8cvO3G0psfFrHm/t8nuFI35jNadqsCPSdxvix7uTW5r7g4e5yR
H4MoNI7xKnb9IG/OR/fjYMVWX1cLozr4C2JH7uvuo0fHmWvIlTMmPbVWesrx
GENihAcSIaIjfyGwC+sxcfvwhYJxXSK4dSEUUCUDwSonw3t4Aj1oLIKgFFWb
Og4vajL/2ySVZSqwvIztysFNxf8CbNrlnzv7Z2Yc6rWFoLzBkwBdwb7F5diy
EKwS8bSfc5C2CwP2s9ZiVEBs4sxOkgY9PWrXnQG6rYVC8f4eqM0B0lUDvOV3
/sCnDnXO2dl/p42gbHKAI+emzLI/VIJD0veL0NiMrkg/fSYkrZFglAf0YRGW
nsWPBZwNivwFB+hnnonBk3gjyimxHon3q71v3hPxnEswX+jY8E/fFz8HlppV
TTPDLBdJzMUHpJn9yCU+xep1gphQeJOaQY9QNT/V7wF77koXc+tSpjK72lGO
0l6LFNrJNDrenvHY+se7r+bGZB2hQ0Rcof0/lMj17ZMW1grj9FQ/EN5Y7bQZ
WueMQ9IMzF9ktOTU3Y/5rjqLZhCkz+MaMXjxt4CKr+0lqqCUiahe9dSH88JW
j0Ce4I1aV+ePWiRpeQ9nLIksfDQuTq5aIfIvxCHibmAd3HBqcaJ+3K0VhqsT
fA+n2fHDyqGfg+vkMGjWVWR4+06oCwi5xDxm0ek7HQD+i4giz7D+wMm+2kx2
tk+7h9cr6hBg3V4RAyGm+XmuwTExyVz7WuDTtF8GzdhUbpJylDcyMLqI8fn4
up6JsgEpMu3XUK3k15BcNK7BAIT6ES+OpbdsyWkrezpXqSQ4uVP4fyf7DV2/
R8+K5KVbLeGL9x6dhcR+hGfNWTd+LozFuR3nCzH3NwXyLrNZ6f7r4zpfFarX
VybITCA+bQeikbjA2Dp4W2By5OlIZNjys1IgipYwkvMgEOAg/B7IVb/sVOIu
EkWxP3mPNijVM+ZKHe01lHPaLLSRG1J3bYGgyZzMpK0R1138jyoSf8YSOI8X
RfE1E+CNuftz8iWmdKfS5g9iuDgSK+asoH2jCAG7J7pziXICjqwnx/fGPTBY
zy9f9zx8jHlRvxfb3bSTwtlKQaVMhCIlEpOjTo30SPw1F6Xk/AB8Kbqad4Wm
POO1C6MXrwGux6RZ6hROfgBsp0Mxbvw415XBoXZdxHfzdo8FdBjqHbcLl7JN
5qqRbAyUI93VxaENFlIlauKbBFfH/e9MWCcXKFomMHpDWhhWFNC2h1PM2VAk
maWZNX4ZwN79WPGOLqC8GoIJ3zcgCnekxaLRNTTwCUZubUA25EzUyeXNTDnP
arm2Z7/ew9WZ+vC0bGy9VymvruyhLOWPcRDktLkHyLLpjsr8UgK/I7QWmPtj
Irutodfrqv9fKbup5sNFnTiVF/B303gaCqMhdeGxUKE0DSk/HncH82IJdd2m
w05wiVMbVC6nMbHWFOTMq8XvNwpwGhhDSADnEqw2rnkZWkej5Yd23PeCeDlq
vv8gCFFytoFdfas9AZgaeE5llAvLo9AGwlH/tAEwWq7QIUYcJc8uY3F1gG/p
lXb4go111DXCbuV7dIEQSZZLiOOCkl3ry+nPLUAFHMfd54E5NfgEL7OLdgea
Plc+yksCXTnD7l+Pf3FotLqre4+WF7tApP/DHz0yoE5jqAuI57T8d1pW5TBb
rbTP/LgQBxxWe8nlSwW9EtapVGOmg+nuFrQAAF4P5O/BTTm5hqXyhq0QOSjO
Wv1Iv0myY5PC9e+onPezDykPzgZw70LzJcGAuEcKexG6+DEXRJE1ZVp9yEEx
GAiEEyD4N3hqANPkW8eCI9vn0o90O+B1zC68a6vDgSHieVj2AvKasHghOS/Z
AjY1zLIUx1uZyPvEDC55rhzuqfSQEs8xmcRWfSLVez9PgcD5ljJ6F/Q5bDil
zgIaf8xZLYvpbuEMiOn8jsYkbJxayhhNX/ylq0iyyPBAQU6AM4cm7T6/T0xV
GVekeKzHznukGvPsofL22dnluNloLHCaisU4f+JF1l3OjbBB6uzx5gxgCxDv
1bDMRIi9Dibxcqvs32Xfl42DQ/28ZATS+vy5GF8U2h4x3GaxhWcoaXf1+Kir
2S4j/u9tvQeN4If69KESXjR/1QIZ18S11W79z0yqswqup27OZ2FYBlP0G5/C
HFYFOUVi22kP9C9vNsikAoKEne6ppZoQRCHwLd8syCyusuBrsXc7DUdtaCcm
0lsHMXyaQK4J0kF1dwjfRgyk4QgP5frTX9zJzs75cGv1TAMmvzD+hdAKzBXm
Go9NT82s+WmxboyxlurPmF+PX7WqqeheYDRfXd8SyTMZIbU+vYZM82sIfL2A
k6v08TBT8Ka5KyFzWK5KrjTuJ6mkV7KJvWPwyp40n9wwQlX/giIuSjoqNryI
qGeKiQc4PDR7L+nnjnicnYwBoGw6QDraop3y+42L0vNSttFisKtG+yIIncQo
3vV4CDI+uvTDgHjW/GnEaxlPaI0PsuuVc8rB95sJJDX6QNVNiiwFbTjqy+CR
Bb33g1UR1t4tQKCMm0YI1DwVUUpxd6jUZ3DR8K9WtuhXCWD2Qe28sdlA/RSb
0G6ioTH0Bjja68pEUEfvJ3YiDsEws5+Q2KJKruYaomYP58jG5xMc7OzBgqmt
9ydgsPCjfp7RZwOljHFd/duLeRAS7yDtA2baFOs2rGD74CZOkY2aCXOTlcbs
2fNG4lQsQZA9vcqUveaGYzEUpWMTvQlTeBvx5j2EvDTpSl2Ab+Uw6sqQwUbh
X0D1ijT6sRlnDQTw8VwO5gswV8rff8MfrS+PZDbEgmU82jM5RAPu3aRcREpI
sAAXiCRJns8snCJWSJvGTfup4gpMvD5ZfhQfdsty1IzjeDig9Ry0Tz2U1JqC
RGn3ZSPV2kWEzuQTa2fNGlRX+Pxfppzi4KSrmvgeMzQqN9adbloZSclOJzoV
lNTXleDYU+iEZurL8r/mshXzXyN1XS+2iB9M2dlkLKJCg7d6/KHtaFEMh0dz
o58bPpY7YcNBY/MJERPNLsk5ElHGkQCh1X0nUuZHCL+CzRKPHBIobFgzELY+
PqkwHnh5oQIQbH1rZDP+Ug5hP+0/1v6MjTrbUdbAWl6knyh2iR64+/zvBYEc
SS/iUvD/7sC37yAmiHgx+RiDKowNwbgweDcMRC+IEuShiNADNvYtLEa9+/Wi
Rj2GZaRV1gu1r+gmEru76NxP/xEq8kIWpKokrxfLdtEqdhpX1NqhHVTXmNxo
role5pc/nMgna7F9v+THY0s4KrdRAAl8jL+rBzzpf3aQ1dnlp40QWvZfeFIN
+kFEvUTdliuPi7qb0PTD+Wj0OPVz7sScHYN0TEQBvHlqenC8CF2T6ZCwKNO+
1M2+N9iZJJUO1b3lwTxmCbVzVUTVqz36l2e2B77z6tjN23pK7Sb/mKOsZkc9
ogWeigCob2oMaUlrkmkbryAYHILEOma0zsmN/3LRjN1doOb5F08SDppYNrSC
UpKYfpP7s7UaOHUk4Hi8ra7NIi27nSIV6wSC1B15Gs5L5+7bp3fo/gWgBiPj
YJBt246yJTOSG+rgDonxQPyLKYxgl/vvnh9JtckDuzjAzSsm4yYtNqYCkm94
eb4gJH6Rw+H4FHcKoSYRVrdETnw/Sj2CXMh3LZ8Ut3fdLxGbcW/nxbWF16ks
2XLUkvpRFSbltNJA2hA7QOspaowzWR2M9auCTaWrRZfSAX3paROd+8Wn0bFn
xv+a6ijqyFM/AtxA+7QA7txm0kffoJeyKCJRAdJDXczjkNHoUyxKwM9mDC5Q
ROpxweK2OI8/ww0ratom/Q0oWuYazwqNRZMG9n8FCANWtFaVPwLlmzSRNMmC
qJU0JvXmSyXrAiclcvEK5tyG4RJ+B8xY/MBRVsWvXvNGLOwvfhuY3Pmi4Dg0
j9JYIC0kmsk6BSk60Y/Zfo+chbe5+lpA1+KiSfr8lGMOmjC3MQ6m/R5aBuYp
D8MZ7GrgLHadpGlVZO271A2yDJHPj33eh9Hiz4s5qWSNTMrFxl9M9iAgwEKr
q4cSrkyMmFTlUugpX1Qcw+ZkBux30u4Zn21sC2HoT2iTJ2vVxXEhj3KB2Pt5
mQIS246JIl/bYjDNYIxkeQgM+dgH/a6wBXI4AXR2tiN/bShHJiFWhxZKdQd0
T92b7p4tjxDqhfsFUa0BZIh/0XE9xWPoCH4O5VJyRrhtfpXJDFKuYOEZxQNo
bikQl4EuoJIsqU0rijpWOCT0M1PNp2uO0vVORzfe3iQFZhODSL8jGj/zAxtP
JNUlvle/2STrDJGAzKnA/S7T6uDpXrNpV3qDGa6qScMM+A23ZIwHuajNFXee
a2DONuav4EG2VTAeFLB7DRbeiAWSuXoG2sDYdvnZ02NRyV8K55ZaGObHodZN
9NAEFD4YVoG5zk0cEQlMLDvzni9Sg9aDgGFjdPL3G0psL8cIvqZ2ec/PSKFi
ASpAH2XNmjPoLWyeNGnvrfN3lZP+j5P50/DXBzjvp94+dZxQn80LFxN+vXzd
tpI+axq+0lxPCpWOLR1vK5cAhkWh5Lcr69GqM0GcivBgaHW6Vvl3HzIq2HQS
sfCLC5TCvMSlloPAXuvrSSiZQbXCNsjuoFFStVWJbHbc2TMsjHjjtIpa+Zue
Wul+5drfObk+da5me8lTAaIVl7CXHDupvpSw8+Mf6FLBJGcyN7JhLSoh0Rs4
Zi8rf0OWLxYCGwiM/gjqWdJaOz4Zmc0E4AfVHUKuTXTJszaqRhMoSyHtvPgF
UnRXklsJpEHImn54oqZHDpBF43istEAbzKbgoFa3+W9Wrhq6TV4/T1m2T9UX
4pPR0NEN/9zu6+AeW+xhDAznoGnyvqcEP7fHbjyX06EJh8M+fDVTKHQet13E
+1wPVhv+TZutJfrLFJLR76nFSkDDjSWmQE9Oo1hcYswAkqb/xdOxLQwu9dml
GqAXtt0XR3WcZxORtwrje2UgOZWP6xX9u7leypfjcGRAqTU7YCpdjSmaBvtF
GDG8nPJjiQL/sUL8s92yDVwJL7GBWfGCwhLJxBdsu0w18XBJmzWG390yoA41
30IhbTq+FYeWrjwrbFscnuIJ7YNSJnDkzXnuxL55fcPc3RjH9BICaQH4DnQV
PSh4a82T9+ahFdfiQ4/7tbtKBy+9RVEEbZC34IOW14+Uf+YDofVhokoVWW69
FZN2yEbiWJPFffh4Tk3vpsbC+k1dv5HTJESc5aCURnL9tDCM7Aj2DQOZollk
uUIFge/8feCxf+WqEIF9UgOKEklgi2OLTwmuQULJqcfNOpAnEyNKFyMA1ckn
3xyFdLEHlvWUL/fPAAzAqob6tLuaT4kxX1UgGyj0dAj0o3FHCgbDS/lqEPTp
gepqabcPYQwx4vZSDd+d8/xLwTWI5viaVznU2jZJBaAyCNVpylkweo/huq6f
um8DFBADWl9G0U6TuK0FzH8SPJfBfy/lzN+O/bf8IsC/uybFgae+tcKmjq0a
Kvi9SJ3kuPtAdxN0OMqpD698uA8AqaVVrIDolynQIfxOOTvdJ3LPb2URW5eU
6Pf/ZPnNQ6kkTPV7Q/lukwx5o70b4fuweWsqoDFX2CA9K+vaM88YnmXL6ckw
d0cJ28taIdCnMZW88/RuG04v9vgWVvctuzC27z4RtUr7s2nv32tolzJVqWMe
GHYsGdv+N47pJBG3XwH4JUdm420X5100KgDkTgkuumxgmrOulMMCMMx5RSeA
n32mXTQdtPeNyXWizGNfOwQLtq9nH9D7WvM0oWGRF9ZyaNPL0QULiB+ChK7N
o2dqOdEY2gmFrvFnBPGdJwEWmhW+VPEfJDZqtGbpPSgMhIVXnOD6q4AviXKv
U5GY1nLI3F1EdDTjum9MFdS4kxj5r+9Sr2mHP3BCXnops4NUGHBOw+um2X6y
ttW9XITEzsFAZh/eD/P7U9vKghS5eRn7KG+2PKylvlcXuAxI+u0cL7lFZ/5x
zISUpbGhai59P1Tx4P1LGEd0T9wJaOeXCiSz364+UpBgjNV5YDhv1VjE8psS
w52Ey6aG2KIHnU0LCTJxCwMB7C7iOYH0siP5XWBB/DGP5NdEQBw4xbDUHAQV
3zxTAfgyIhg5KH0zJLFDQDkxvm6dxT0qQC7LpuByRwrJPAu8WtlN3gJ6nnQD
EQ8aAjHkrMBUL3O3BnvVi7YYyYwRuXaECQrzYqsX493jkHt40EvscBUnQOuO
qUz3S5WWqbhz7RWnqtRRBq8D2xLdEODXozRhZJDcaRljFOgPoEPQnIHvDrat
fT01wNXr0uUKkSDBI0vec26xxdQGD3i+JODmYB+Nr0TtTbjlFFMOWdq/ouFf
lcaMMU0cJ5keJh+P+S8mbFliP68QEunXMotM3lcqnmv2vMJipmLI3A7m1B/P
Alx75C399V+AhGxJ/Z/DCuRDwCpHPnTck3b1Twf5EKt4XDNrUDHLExngc0fM
ikW6ddsPwQ1z3SFLPxlBr7yiJUj4muH7N6TmOXTWu6doicKOvc46YGUULjvR
XstXtREYdIHrY5weO6ChpqoSIhAZN0XOH/eNsxvxGRp+VuR6touqwRDHylHR
nq62OY6FXcJL4v2gtup1A7cJbiCsRFOycC2OL1tSWvrPnuFydWtjxl3EkeGH
hFMWBJ3Sq2Lr8g6Ly4AtlTlsxxPZxvS2mOAhrshbdJtrkubOWJMpO+dVdnBG
Fk50t/1imf6Hb8cK+p2PkL0OndYYH2sljPLC6BZicHg3s7GQJfXfB6oT+2Wf
Th2fbo8o/mzfYNzRt5VMM1eS3TITBOKfu+gQ7m+22RvvxSIuFeGaEiPyAMKo
ixFPlAsPJT/Kt5b5znJ579xZh6u6twhtJEkwzelcXclrYd2P2UP/fIufKF3D
flcF8/KOOFWvXaOJF9LOinIQSumkEy8IdCSTDr7FK8+uauSInRS8Y/HtGAIK
tJY1ouoIy+kA7EHEMfEWQdigV+b6+sfnrTFEQmSktdJwCtkQCrngLQUZ3BsY
Jo/P/i5HZDJpZ7t/CiffvnIZWgK7gS9c94ICnLbv3DSSbCefe3UXJo0JAPLP
dVXCBgymeRpmlON+n+fcnwZE9UjCXc6LX7iA5xVZGpUu8authzMQaq/GtOKe
uedQdQ1/AO0LFtt27ZeW/SmDX1l41pGWLfrBQ+DQ/VpPWOOPk6j5UnjVf8Pr
BqtfTUmxbl3cgCw/tk/oq1kilvoOEJRNJqjbb18dOUaeq8ud98/tzUxsKxA2
dT79p0J4zlDIk+kf5G+M60GaMgMHOJKjCKFxdSjQobQqPaf5pxsJ8vzBTUc9
31u+HeJrFgIOGDqF4skS0MZ9jQKFWnE/wuTVoiLxFTl2d7ENh/n+Zm/g3O4v
oTgktmoAR+9M7udlZXzHUIx9K/BcNN13vl8u+uBkR/V7T59NuidoJmv0Wr8X
+v0MblAVbMq6Psw3BQHPjfmLgc9zTIXm6As4kYD3emvZcXnR3z8XhkxYM6tO
XUjOgj7O6t4mL+sP3SCR/cC/6CO+hVOLUMf/vPjVgxdGEQxA+FGEGBPeAn5L
yDbLZDiWwPYqK96OWPt9STvrjdHyrPm2oYCL1ChVpl3XdBCGRIGR1hAsozVo
XIpFdJH82fUQZLdTpg3Jb5JMmrYymkqrvtW0ldJZ7hNEkcid9CbVgAqVf3mv
v2l4GX3+nzMgUOyMsfD4vFvniib1hQCSpQbVcHGDw1RKKTDvfIomPEFZ2fAt
r7La5kodwACCG4l4KlCZLtSTojLH3jh6/pbhD7mU0laW5ZjJcPYe9vkL4Opn
Xjs+Q7y9kIM9Eo8huKxWrcLgIovFe2wMY2EFa+azTtNVJ/Rh4o6Tu/XQMI/y
SiCfU10gMBpnY5yqrUS8helH/CpyGkqlKNByhKFG/h9kVOnfn+Sy922rw0o+
3Gnw4bt3IlsFXoqL7VTn9kZrhzVyAH7ireWAv/TyoJijOFOAGbXBtr5Tiqjm
cDt0+LoqRx08HJZ9ZAVX1AeIr9wjrUy+4ztr7ng+DRiyvWvhg42ACryo3sXe
C1sDxeOnpfggiV7Yp2tHJg0WWd+dnPimzIkGYx+KNL0VT9er+8oQryovnyAE
9ArGH+V6yOicFTc5ourKKXszvLypyk6NuEq8NYsmmtznvLjJpWVSCssYeWap
VqFTIppIYs5JzCOHoAIs/Opj/zy+v0stUwWQ20nrPWBp4+SFYjsReUWR9f2K
eglsYWggFvYR8LFWRbjsQY39QRhD1l3oIO/vuQJOX/13jZlw0JKU2FZKaaa6
KnjvjyhTmbbnEid2afWyG8hr9ayuPC5VuA5w/BLIzMau9JSQYFa7pazitroJ
11Dl5oQsGrB/wOgEnbbtidEFXSxeyHxZHXvKs+hphzRP1NgzU4ML0QRqaQxP
rQNexaTukmZyUOwINX1CobzypuKo+WmGVJ7dzaRU8Sfvxf13GCi7nxG+LB4V
qno0og65U7zU7Mep30BwkJlyIOFWrq2akzHNODKXFOnU0579kztxYjlTtnyq
Rbc8q5aGmLFLctbAJ9BByqA/IhKp7gR7w8DqH+wVt7EWWt+5448ESF6KTv7R
dsazAXE5yQgBl6bk+29udI8DG1jGiLEstBPrgbn3kTNQ+JbzkGR9lwRURSkf
pNR5GFvaT2JIBsQqwblqfwh/90ckeEVOFO26hEeoL3l3S4DQTpEKIWz2c8R4
xYIXSmzgHZoKYk+bnqG98OFwGaoOEOGFxKfSYI+92oKyqIZacPwT33TA6Srq
bHlb1NW7nXIYFOICZVDuoXro+Q9sL3gCa6SrU1Rhr4rOfQYNl53pZrDq2pwm
LTrcJsmz4ruNvjV/hgGQgjk/QBj0DR8d9ZWnUBZFJY+d2qfpDmlvpDhblSsL
ti1E0vSwXcMZ+cI3f4tXQGYvsAnknCuzPqgbvrmQX41Pa/UfvRO+RT+y0xEi
vwiskt8iihe37mlF+0GSa9BSp1ozEoJDTjDO39yj4N5SRS4Iqwb/5O6Ddo4O
bFEpKYvJh7XbF65a2IfT/qTanIFKi6czo4rpRX5i9M05GxtL8QE/1oOZumVc
QveLa6qQRBVUZq/wgG3C99TwPUXsjgeUWcfLj1Y2VP5z8FQ6YB/YFimugVOr
kbs/4leySSFJqHdhiNDgJ1K/vJJRDzD+hRiWrw7R/GjwXkF+aasPTrXhGAbb
dLaN2RpbNBadfwtKOemEo1y3Gg83+jrUOWC5AtR/+HVMOyv7o34Hzf+sgPzU
h5vmQdT6bsGoDHOlUv6BtONlTQjtw0r9ay4852UXzJQXkzt7FUqYRSAwCzFr
W3snSvyFOQokj0dIb7L1mo73ww4kpC4KxqcztwUHQ1/5jsDqO53bA6vBWlPZ
88P+LEjykwnrp/ycu87W2ad3Lx42t4tQPEjuNsM2b5Zq71a5v8WTWrrYevMr
5LuqPnWIlXB5t5kcjK6faNssUPm9mBQ8vD2vkLikMc1ovWsqhwxWi6DPTvAY
zrZjnX8zjP1VEQfZyMkaPDqIkgnvYQeDNET5+4jDmrD/F3zzkaShDjFbBJcK
S+22CN9QesKLWS2IFtF0clr361frgo2Zc3xVYjONZVG0jR1gJeQBSjCTHr+Z
pzlM+P7vA8JbFebHUPsJq+7VnkVK572jjrCky6uA/4EfcqD+kIfHqeNJMPK3
w1EefDvgbEx/bHrIzFq0uxrWRH6fPj5wym0KC9NfvqfQaSRyVMEoc9JOSoA2
VVbUc7/5BMdIZURGHagFI2JMOUSkoHnzHtZUGHUNRa1iBaj1fZPIGZPHN7IZ
mNpFaEggVauU49QxrwP8A337MKxXT/HSOM1CrCN20BvmF0Vo5GNM3iUSXmOm
+geScr8w0fM3nASHPgC44J2SH58n8o5igZlvSQQnvru3IBpVtlYVuhlfU47z
Wx7T46C1QXo9XWXC8jkh0v503ewWlwPsrqB8yZ/QzlLKJc0EAsb/1hI85fNz
hB9upWKYqmPO1R4rlFfFEOHyG/+6RZI3UTkROCoVOPAhWAlYgurKQjbcoEgC
WSBTDkbgiLL8t84HzJ3kVCo/8ArcHyZEDMwfsINgSL49uvbiEapclxSijyin
W8NYxrT/CVshsiI/kH18JC6qP9QmNgleXB5Lu++PjjB/wraUuFHePjVO3PG4
VxKflu7a37KEYAIl7/NyMt8tLdwHjcc9GZQO2BdqOQXs7NG4vODdWUxOUYcj
PqNznVC3M+hKuCimam+V7ehRrzMgqNFDGFGMGb/N3VzHuojkMrgfoQgPAtH3
Um17K9Dstq6EiMWR/Oz9LycGeJ4Djq0KlbMsUV0ZmMj1fcidI8mqD9x1pIFd
Rp31VvgiA/UrQ+iXsI8qAfDvkvkEuGJ2oiCeEA/IPFJppJgxnoMiScHHS2qx
ht0+azS+fEbmM/AoVJuBG4DqhO9EsNqPw89J2zqUwsZ8t+Xd8uxcigDkgyz8
24hgaXixmvk4JUFnDeJVzRWB2Sq1b8xLfGIC2jMIB6iWVrtHJ+J5LG68VnvU
Qts0Pun8ebDqoOLUGVph+W9PGxUURJiFlG+BlUVZHfDpUmo8uP2H14i1U70T
NOfYeer66uML3VJ5j9VLHoWpvhzhkA+ZNKL1H+wyWgdyDswoSmf/ErMaHs0j
fC/OA5+lAndlRSMmlN1EAe291dah+l63v5K9xDJ/FNHPZTAXO1CnIxSdnHmb
3kT5X64JjzXzS9Ewl8pmvSqshnmKKXPBMR435v9QI5yvQNYEwL/d7XC0rzIi
0Cbg/tr2RsyHr4/VX7H+2HkS1bwxQaIEXSKrNWXOUSWKLyJcM+IVgcfZPJvA
yHKsim/VRLBTVAI3xDP0p9pBhZgUdW/KWixnqmrH3wwKjz77nsG+3XHmT94B
hYyceNj32yxSt/Gi82cN0qV9u628iLvHKAMyNe8wzv18Ehsfqk7MF+jfTkO4
OHnKm+4lfiF6vol8yJQ43bC3/oSxm6E4y0U8QnXdp4WvMLRTQq8VG6OLhsbm
seM5UU9CnkkXAKuQiGbxIK311la1yAjeFhXF2uas+kYPIdB7XXOOX3PZzbQz
3EYAnw3yffHiSPsDeA6NZenxlP6T41IQkfFsMvGqcJWJSpYmvd2Wr4tb4WBP
OcZSi0k=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeiMkKoAmdRKd6a8lVYmcbZrjq8RF8tWm1uiVpYpXDUOZasn5xAE6M7Ng+dqJObhEnWSq7hz1l+tJi96t3p6pj3lYaWs4E56CkFPLo20Y/cVcqrWCjkajGSBnY4dvyKVunY4ztPGmBef6bTSSSaL5ERQ1y/l/yJJlTNLgcRBD8Cgnb/GEkE05Q9i9yUeVbH3jSw6RIHu7JOvr4USBoLonvwZQfScrJTKPBaTf+JxmlesD0+i/ipyKLlIWJMBmXU6hVhWF3s2lJDhlQUf4bpLRShc2mfa0ZvWjBeYDLGyXz9s6UilTRsw/qQFeVUaX4DPCdkOzZBQxDUyMpQdhtHDwp2ifUzBok7+OIJfIx3M92ph4EFvpCTm+jrSnuod+2oo3YFwxPBX3pK8EYhsf7m7ssNOaQsZjx0V+fuiYS9fNjKTzWdOxrHeSJ9Sq06rsCiqqUp+T4yS95/2JdgGkCzFPY3iuSO/X7WydEIUqZhc6OEPJ6lJeWCjT/zbYL1Yn3NIdWaUhLSgq9c/Y5NlBi1iNNYAYNXo1jAs+SjKWpr955A4LdfvLac69Ju9+tAqXbta31m7oA63V6i5La1ajNXsYci71sb7NLtVFEeQbZJDnfZwE+6bTiF+Hfps9EZcC1OPch6oszz8CucbWOd75Mw37+k9hMkFxEE1XvjjyhFXhxYJl+7klOwYUQ/+IlxEflRM7uLz3/0ad+xT5mGFlEIs+Mbme1EMjv53XB+hmcZYibV9FU5XarK9zdGElwh18BTDZS5GLjJL2OXGS0zWzS1GGyya"
`endif