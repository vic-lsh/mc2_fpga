// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p17POFoncOO3IfZNqAoCfz1h2r5i3IwH54ksew+NjsGutHbdy6dNAFFu1K29
f5GsMeUfhfsmUDYx9Pz94OqWGG7uBl5zeqzOokVNAA/qMdFJR+hWf+iuccJK
mPPuOnOfc9sQTSegs8tx2E4I1X4lOYWc0i2isgkDKSA5k2fkiGofz7iyO5na
0DRGq4uKjHpb4nMJC5Bs3nRTJhKMenVSw1C2N2MNVzqksbCqwBZtxyTYUatA
kerCWAbZsJsJD+UWej3GDlT8PdkTatg6AfhfhLIyDOsUUS6NaIm4FiMLoeDT
RPlg0FGoynz7d3WRUQeYHV1pasAt1qcegR63yltk7g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cYAldTwquSni1XzUYXl15ghKkCXIc0yxTJzY4+bPdN/jvstUKErP9JQ+ePFf
3tkktl0DEJtQUIoo57wLdDRhC+sg/paJ1RGaEw4Zf2Sn52yjOnjes1bPI70X
t9HNi19Xo3IJQO+qBJDWCQvcNo1CJDyrgJtDbmCAe69o7TgqlHbTO7JVwbDd
pP36dnGpG7WK+KkWtnGelmNV+wmOmSQfZj77AFPQt0M89XZ8PcDT0VHiwnvG
mO+I5BjmcXJEgNq1mIE+00QZlTPiffwJ51lg6nSoGXZ777uZYBN7rU82Nrqu
ebG5kqkt1COsY9Uen6odemTTrWdl1KlK2aSjRCJy2w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sU98zMo4rrsRhrJFz85mnpWpMh7VB+gnOxUV6m74Hhmk1Iiiu0u6XNmFGDcy
MpPJIsSPNTkXUzVj8edfod022NKaAe10Rh5NkKnVs3hhoD8ks/Vr9mKPd5Vp
gmYBEx7N2n72gSgUQfe7vzvvBjDl92pE+0BCGn8HfM7jUhQ6aumWLvauhA6a
OSvsjGvoreGOjgB/fj8YBS0yQqJI+I8JQjlb+s1TrqnTMgW2SYPkCguHUoW0
6y+Rozq4b+vd7wDBehxKY/oWXVmoIXI92rBZu8TnngVravR7mdUe89Qj6KbF
IUEc/d1B0+5o8/Lk9EfY6tfXWSMe17Ha3h3FQIAZ9g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GPVeEQMQoP+ez3MvDIMsozD2NLMXyJdJMg7wGRNKxcpdhd1pLNgxfRb9lf5Q
bXVmcrsk3GmeEP30mVnnjjJc45cCQS44Qfxm7wcCEmuhqBcdzJsZnq0DErcw
KTwbUPGeB+7CXAYqzPBAbl8aGeTwG4h1fgl4xlQKiy1BWZe78HnDhTerqDkz
lVwVRm0tpHObEsrcWRi4OIVH2K/AKwMn0mLALFg9lx8c6/vArV/qWk61dS5G
QOS5C1m4tl7Rd7v34hCDMYSpEKh0Hk/Rj1oNOWCp3dCzuMlviPilAj2vRzy9
YA8p0uXU4YiUB8Frhgn8QCH/3bX7V8BhZSnxZYhRbw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BeeGOzDgc8MA/vEUYso1xx34RZf0apPZ2CAEidDkG4FP5zREiEoD44swNQ72
6LYFMAmhx9rJ91NbqiDuO1jge3qUZQXAaN1P9dkPZUOYgn0F0rfrgVL9w/+M
/Ts2IZq7WCFjG1kjVIFeFrUwTJrkf8Pzzi1KtnLa4oIO4IRPwxI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Aoh9l9tGVxV7sXwwj4BozhEkCYkIt0C0+9Gk3BQmSVNYZKGDJkfk7kt4P2hK
Tp2KBijGzuhj7uVQwoUlvqmw3Cu6q1F0FVBYGHnKchnCp/phaGnYgTpLBj2D
3bPWfYo3hIxTNG45NVCdHlFTNobFHE2aZ2fUA5gjC+kqu9zJlX+1R5eOSkPD
O0SqECHe5R/TLAkQGhsFz3ACHiFGPH40iUm4ymu3RAhL7XBbkAyWG/zYPekS
zkMz2KkIiobUzQXAc10VEKeTm8LqKqr3ciJy8Hb8NVtl/YLJjqDexiKeuK91
luvj2dRloBStInSaRwkQklykYVL7wnxqSVL0jCwV8OjX/Hp5RXz3UWiTvF3Q
UeqS4N07+cO9NDx9hnKQXTOl060ChJNtAKv1XpjFY7XftemSm98SW+jEb6dp
8NLHxMR6OWUqKAL1XYbYke68rPfh63hNN+5LC83cBCigTKjZdItwHcMQKHfc
zGLiLU7iref8dpnaGpI+MG5FjDOnsy9r


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SD4ICizW9WhLVmH4vTSnJlY7peD1jhD/VDiMXBYJC/iwMA4Djy+L+aEfCuMt
ehV3BUfrpLLU8RDE/MywyLERrWeZa5A98Wir3bCnkqAFjMOhfal0EfluGp+I
NGkEpfIrk8yMMn3oTGFS+Krg8TUToN8jmRHyvC1gNqVyeUjOtrc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mQItqBSFlqyUyZJBmx69IPMvofFMfTIWGu527n1BpgRj79BruLNF57w/B9ze
3AXN60Q+XXYPp9j+fzMJJx8aOVhtcpXwNez9+Um2+Zny5sILcXAhbNayFs0j
hutaY47RdfO610SgeE8E8mGoVcoyeEZ1S7tVH71ezCO5wiNSknc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2784)
`pragma protect data_block
n/sPv00YMjNTZDbnJQHS7RYnsI9m8LjhOD17GbPvS8+5C8BuIDJe4rO4+fcq
jd6UvWft/gxNC8h09IFKGsjVrAxk/0RSqeotrvvNWETZRhKr85niO+26BSqi
MZW2NivUfxEZ3AxjAvZLg6d3k2SV79X8TDInuDOZpjAxbQXOJ/WtVsubKHpB
bTxAf4rjDKsv2hl182LHMR3mQI4Wwt5S+ezVjBRzilfmOUcG4ya6TXEo1rWq
tzJpJYqU393RV7Z3lpPF1uEg13SeHtwKsrjD4+hYTUFu4wMmBKdSUL/nwtP7
8zJ+qASH1nJAICmRrCEJmVx92bKA+UOT7/4Fc63hagHQWMbGyKF+p6XbPKve
mpc4qfnbTJfPtPQWlfCn6Zfo4pX/cvdmFo4tm+TkkxcAqjxztDo+HWgah2mh
+xZrq4A2D3DUhharIaUT/IdC3XKobYxIsmLEBzjoThSfEvgpXWOcUDbuu80o
waYtPlmmRzKALuEwgPhDkrKDc3TIe0+vIP+FrbtpMylRCYRhJQZtl27MkERe
e2pe7Uz9d2LO/yd7iRgEFH5uueh/ESh+0PSdkhiirzTcLgioiMFXVJt3OJwm
meJgUM01ZGPk+Uho/Xa+Y+vVSmEGoPb1muGULm5uVJ1TvGA0XecHDEI2wpCh
jiIPqUI6xks+VsoA8fFQr8c8czIHdxWI/AwTqKRAsserNLtEONDp8ElLmYAJ
G7RzDFAM2jLcIGJYMqiDHLJEvXildF78hS9bt4DZtdqwiOMagrsrHr8quS4l
Bz0kudRiytIFKH83CaQF5jY/My5c8n/gMmuQge4bTCiiCwWH7I3hkFxZMP8Y
5WyUMbEVFFOQxCMdt8z6yxp8FiHO7OshhYG+k1jzCyDXz58WInffw0Yc6sD2
7iKZDikEPN6tQvVC0vVQQeQ5af4P0fuzILugnr/zjWQNXVQXvTH4BenHgKiX
bIzrKtL07qwLkAQAToElnUN5cDKGi3J8v8wVYMA9fP/Rlx1fz+Fsi0E6P8yu
P/w6zD2adj6PNEu4Fssn8HzN0oyLsEBr5W/rbNUV1i4fQXUOylecD3JQuYMd
a9dgNR7mwLw6TzvSWnjWRk2R3vctZS2IPtTuBgEiMRY6xyo6LICOQa5Rl51o
H/qSD7d/y9LeVtIPN/KXSXeH1H2wekDphWhTs3CN1kQ3fYyOHNZtFHoLnBT2
dJr9uVd0Och7rbwfb5JOqTJnwPIDeH6tEgQohg2xpo8sZviwz6xKfvnByU+D
0wdHjmpMNujkCkKJtGXuuCB0H/k0NkYcScM7fB43+imQv8zbCQF2C2za+XdO
hVMK28AycfJo5Beofbn82iHj5FlBGcc4OrBcUGaXopzf2aNR7KFhsol6SEMg
aWVviYZp/eIcPRcSiH24wZDnTeIJKyQ+Bxr8VtWSnQzMtLFbLpzFoMVmgyY/
Cl+iApbAHxCoIXRHPPJiVua2C6P1oXLLAMA3NGYneF0qHHOOXtIK4MKkWy+l
gZ9+NqUUY49iH6hRgDzfRtn/v8TUHJ7hjeWtRGoA15Ix4/kunW7rJ7PcTY0n
wpdqTIZMkZB7Kbtm5qGAce0oBWzldmbINZ7gstS4OL4VLZcAigd6fksL00/B
EcGijMoNmHG+CCtuYfxysoh//F7IEAyxkzWcg/lQ36wmx8HbLMpXXxtKsvfT
CQFBQadGmo0EGaKJYCOIgmlvY6ivT38kzmabwYJbM1wr/Af71GmFtIyi9ry9
kMBSYOvTRjHKnmNxeIddWOUR6sqFdwyuMod2DOGWKR5+JBJ3BVYFLYr/gQj2
exlXTQRhHgOGGOJjbu7aP8FymHutkvt8SQcfk/mQymizbkwalOmEjJBX8csi
w3F7lsI08cHtwbpyaWXd/ACd6buqROb10qG5YiSLCCO9w6T1rebgViHV2Wlq
5dDBvHPfAMUpP9xqi0dk2YIkciTOkqYJxk/L7BoR0jtqZYUtygSdK6TYsUTd
qD6sdL5JPqrRy3Pd2ylBEP5bnYMtGGxBnfey1/3JYK4ov1bOUsPOLNpSaoMZ
zZl/z3WrB3oE6OITL2R9rMD93bAhcUeu2489hEVWwAFQ1953mnoRWKk9IEAH
YvSoH0X8PfAmbH5GYQeujjgx6m5Osqh6b/6vwJoZgFUcqE0ycJpbiqpaymlF
bOyei7FvKiSAzkzztQU1Gz3Ry6lMNtwwwc5Gkx2VFUU7KgXzygJdsd3rwWce
sRyn+xmCduueEEMqR93PqfG5VZ0pyZOj88rKaGeQHBRO0WaisjB4Jc4ltFRd
5eWhHsM7nLIOZrQm7og0VMQBeeXtYxuVA4f8W16cTz1u71gE2A55L1Ru4BjA
qAfo43H/qj5jaG0mZ+eV9nWCK5mSO3HbMWt4XuM+dacF4CteDk6pdxTU6bNa
6j00O4G5Hgchp/+eUbWwXxT9yuMTk3fiOXE7HMd000L3go8ZO1cH0bWLZx3h
X/ztl4jG2xRzAnaLZPB6pXsbap7mL+xZRKzk0CJrQT1upSrwnVFD0eXZgj3P
i6rR1+s73DjFOG91/pcYi6majcjRAm+jO7CCDdMhzkp6ZnzWQljUWjsZ+G+m
usdqlZXs4vtwjMGXCjqsaaYkZC5htdghM0JSyytPIeStGYFWACBOCUa+l+HX
Z6QYXRw50Fqlsl27QqBTWjAAX/vNZfok8wNgAWlYrW1EVHre3ylHyKpVFo7P
qZBLdwbKIAEBN+yW9Evu7iU2hyU2UVrgDYAvs2ZPyFiaMZNv0x2lT8SCPB7y
qC+9jJA0+Tkue5kLfvZttrxgmwWRJV1J8+UkvF3cXHkY+g0urSYtUmygq09S
os3cGAmLe9sUlrnGp4p730mus4OaO8SU9ixu1U3tXp006xDA1/mocKBhIXEv
TS38N55padjs9f7O6hd6JqRD++OzZfAStvc0pT0sshvywhYCVxu0nBTG/BvO
3rP7XlrooM1BwKqrZHDrJhPjHM9V7AcdC1+k+tL6NixHoqEFgD++Hr5s8A56
9eJfv4dODvYe2jef5EHbVy4Hy319zO7fh26Usc4FKt/HDXH47bOkpmklwba5
hJtw4HayLVoti5fsou1qTbbN8Ax9Ly/0dYQOGls6xm94p42sVcWZcLRNS2Gy
ZFJZj0ASuux11H9uoPOF72D0Mwl4wGbV7FcmwPkeTOkK5Ntv2EiJtH+4+9qv
tyxQh4t3gyWUJ3HA9Ie/vBM6dVo4ClQ9hbm72yuiNKaGQUm6vn+tbydpFMIt
exQ7nOYSymlXt/9h7xnryoUrTGu4gq4DYF26FJkarLpwN1nMAEBsLNx4ZdOq
Md0Km0hoHUX3dbH7/nVxVH32HR46ApvRmr06W9glbC/nRe6z//3ff4HZihog
2LZQefdUHP5thPwLsHU0owZLv2ZXXUvKqUO7/N38CdIVZkFvcGasgRgEgb3O
/YKIQqZy8X3HXvzNeZWtVbhFPRsOvKQIV+cekjrTVi/wJlSYrM9BsRGiQiN+
gZRYGXyJ89pFcXu9n6GjfN8YIhBQz2w8fL4rLhDBbP8EPHPO+jIuX+81hnqI
/sKDY4/w3E/BEmkpH0wgzHCILLCxgAnhIunQUaiMBQfJdhFCYoxKXf+VBiz4
Lanx6/5jkIHZH1P+fHqx0GEpgoZlZD7X49uRzVGng3mjsQ3SVU8M4V9acbnt
pBrJXXEgUk3A1uGMbJy8AgQG1KiVn7Q/hCT9i/ILAO5BiM207n6Q

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeiUaiSb3mg2cslZ4p8NhmmJiOWwtkI/TIN5HhmL2iYog/FNHPGwjznGGX3sn7HBuiF0kIPgTpKD9YE9XFRcM5HOHknRXM8bBxxKUx9sq+HOVuErjAiPmlMLanguqpqyeOR2kzTKsZcgT7JNC39wnZVXQIxQ6djnl41catMMSPPiGdooEbsDeTF5sy+fupF4Kjg5BE4r/7c0q7gyzPezFtebALFbNLxMSHdZpstQSb9S7ltKjP7/K0GY4TZKRawtZVONP2D15qgj51Mif4+lhAHVGunmBgZok+zk5l0u8ZTOkQ9dPJIVV7MYgjZnB3HeNK1TtqmTkEibTaOToBL/XYzbO1lSnsIaYA4sSrSHIctN6IeC/idFbTufUfX5SsMzOyW+7Qh4Svc+/T9Re/CI7n+NnJwMJsKOaTS4MCbXKojAfEUCuviJNPLANNvZX1djdz9j5tqp7T/RoQ8LtiMOzQqOrH6DabfnOsPHS3Uoo3eUrWkfnUd90V6x42YwbVIOSpcCEFB7C+6x/Q9jTxUBa4xfwr5G030fBpsJjmfemwBYuCxqJX+p0BGrcLoQ1GY0hkp8JYypCSME+S5gqjwSdKn6tuGNnTKmvHkwH+/5jFWze7EqdnODrBj3wOPapJDQnPvKBuljsppvkK2yYlBdjdluVSHatJarjjyX101sB88ZkHAMUCK17kKgaRO+A3vdlWG939Ihf2H7kDpsNfBT0Ii+EJNlGD0M4lpoBMQ9TIvbJwGybFCo3r5poUOIQxmV/D3YC5TY52A5n4V7w5Ah7MTS"
`endif