// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
D7jwuF5z98D3rZmzA57B3buh6kTVZNsZ+PruxAK7v8k86o3PQ9MO5SRudjPg
ctR3C0YXi2iTdVbzg45Lryzbn0pwH3YZmhPvZtUhEEdH2d1HkKAql6AvlREu
zENowrHo6x0hb9gtze5ZKm02cpcLSgPNELLYTobA9Cxel0v7sFmsoJKdtx1a
P7fQGUkGh7NYAxv4OIIK3ZWwso2ZnBX/zgHxuqpXeYYACXhtHO/4oUIQpj6R
llb4+PKp19hxYSbuDhOCOjn0zKt9QTQQapTvjy2pzJUrPt2d6Vai64Y8TTN2
fb+jX3dNkldI70wmZkjHLqGTboJD2cVI4IhYb9bO5Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qU8Xu7xqWlE6XXZ6A1xL7vp2fJSeu7aVTuWiq6+tP1TIZVnBakCJroLhOWCP
pxV4Z1NZhPZL4Fl8kZk/7m0L3lQWWEXAVTdgpVXNjUrATQXD+pNzsGqDT84/
2vrMiuozTNytjnVt6uMrSTWRJA1QAene/MX0tB+rwZ5q/MhoAFD2YWFaYPTW
suU8+a/q2Y8t5i1zV+Yso451mC3V/Tvqurul/gWcpO40TsZlXRYG0VvmTq2h
k1Ug7xwuCjceg9TtMuSyupN9wGoJqTqqpT7cPCwRMV/SHI2WNR+B73L7frcO
okB+ue6J8YC1BMTsa/696KhRXho8e85EOQBgEDxDRw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tOTbTpoa/oRSFUdJvBDRKAZzS3eg+O8FilDRyEL7c+++/ryPon0vl7h7wcT6
PNU3nPusL/VhYIwAGll1dv4mf6kJUd5bXR3JoOd9e6vB6era2WBYFh7XT0bx
3HCbhzhtZ5r3iPvE6QlOuj4u7MrnwdZmxpg/l4orZPXAu8pDdJN77B8ERSb6
S/Y2zMlR7qa6i5Zvt5elTXG1qJfn/Ye4gVDBVengZF3oycnUI+ZpxBW9aWYk
cLiWd3KEKd0dEysa2bPJJ5IcN1OwID3c90oCGxi/9zyX67D9gmsSPea26bsH
04Q0beZsT2QOj0KGcqcZXZMJZa4Ak3iaoVyfbPdidw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SpyjXRnbrG5VjH1ZbIcNqfEt51NXV+7f1r3+WTvP9Q16VxOYRyJ0f8iSITXy
bfIs5Hto44UJmZrVVZ3vpJxukOg4D3V3lJjMJ2UcXvSNhjApuN9BPIGWhz70
Rd3QvUVwMq1/nf/ZuCdniGW071Z4SIoLC/SruFb75wAxzwfOmQtrQb9FE2p7
Bk6rEtk3+ggiNxWPtwvcslbx0+lNZS1LAEjQZ1wIUwPi6NSL4sItmnG60J2t
MMsdBLdMciTxPpR0GKpMeX7ztQ5ZbXYEzuSS11offiZqMzc6GbCnqWdJlsMI
QQSi0y0E+7qr5IpVbusQPXXdrV1iYBJYaesfeAH50g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hjBnvgfVz/NrV1UVt3MzFcxFqOBxTkW5EssKuR0skEmLUITv302yNFaW2nIL
lDXPKMrmx1SoyRmAS2jFyQ74LAVjLzjr1MNCbiQYJ713c8Vjs5fChbAurGA3
yp53/DwowZ7Hc+kKSE2W1KgsiMM+vMP1LPcBNDfvGZf3RC5EhOY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
vcyNYtQ3WDDYTqWzel7Q5wVVQo/OI9zps/Z5PJwOWrLjmnmQG44FiAuNevGh
bqV/lk2e5eTOjVLjrnRjuLIYVvorySKWwWVVPUUixnDsZkCQUQ2XrSoktFsf
NOAZwRjRSLlA9RaJpoyxDLfLYg4INsVoUb+lUnd67mQh0W3kM6Bh/mgGyt19
UCPJHDh1heTmi4hvCOFFiv23T5Rxjt1DEXfE+MOK6K0XJlYtolYM0YEEqxKQ
cUZwz7ur3iAIHnUCk8ZRLI/dxaDpG9BfIDs5q7/Mms2LNG2VmYTAU5F4DE4O
KNft7ezGkOzqN/zqFQ4iqmgJJtFEUtw7xxjp4/NXzaBM/Kttkf4nRJesjVgB
Yv5eB6MqZxIbwgsDpGM/NHmG4OLrtDuPDUf918IYldgVSlfPM934g/onvXMe
gIuFVnb3XeMTzC7n5RYSiIZ8RiZS69vXEgZrGHgRp7adhY9Srgum/4odDl6j
JNJUHKDj9f5W1MfjoHd0B6AT1U3k/aVz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sMcMh05LgWluEUBy4RExcLxPTQxRHX0gr1gz1QDGqUIsxbZDmY3hus0tmYd7
4YZ2ooTwhfvrROWcY+/ItqaYtqFjzrrdyeWfEo4y5+/8FHzQUc2/dxOWzkAn
fcNlAaMK9/QG3bD/k8ajBDkGdLqph4qyc4XI4L7rJl4jX+QTP88=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dipItCN9CvByWYawHeXY4pir8nKJetg7zV+uJAt/MYFYRD0Qlmv/WuTZOTJj
blfqeVSYpIKB88/dlwmQgLxqq3ALS1gOJlgW+4lFA7OJdTLIzZJXeSLBMMgs
E6q7fNaQdUGyfTJdiBj1Lr86+eijldkzDFOgkKIN3x3VJ+uqTVE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15600)
`pragma protect data_block
Vk9/IfNFM/dM1SfAHeJ3bjs1pKHz0sBr22nmBRSOt94PrXxWVV9YTQR4WGTd
fR85WFM5zZtwK75QiQhPaVF69dN0pBKaodk3AXXiQpgUvcwS7YAA09nHznN0
Ds2HgTWQ3LWERmQRBHkjH4ePMhpJJNpQ/mg5HcnnxjCnnkS7uCwXjhRVlNpD
TJZiZ0hQxAgxRlJncUy/yBs14s9blQbfgAKc4tlixJPHZ14xahHHLcIS/MgP
zBg1jBbjYT4c/CtgLyaVgiZkw/r8+cspwkPkSKa2E2GxgRJBPSfPQGH1VeEY
gfgJGiUChjJkHXeCpVRegPnSHmf/spyQF5nkEnaYVjDFn6joltuXtI3QJZgc
VspG72iKuhfVA2sUx/Ui0nh7G9KYZexxn1vCp4oZPxygkKk9qVairGEuT4Gv
m85WiR9IwuR0vbNny+gU5dJ1mgiOq3aZovatpkw9oCpBBO/IBcBZCa5W8JFd
245z46oJFZlA4F0s4YkHBXtSIA0KFe7q5l+pdwRGSYpVZZfR/c9DdVkCsZ5u
cCmqdznRKrViZbJK8dI7GfronnrwDdQ3o5fXlJOfCP9foQak4YRllt21WdEb
FRviUWCgFzSZN+vPcSSoRECfFuyl0vegzg64KnIQnGQ80UOPw3J5WJRd/toc
0w+J+jD3T83H+3wcLH4xb7IAKbjecuq35P0DuYkEOm2Tc6imRtMEi96j+Gtn
5RWYbiIwhQgb+t645emT12uWwmbm19VNkhu8fx6i1fkaOtuJxp7UHPymXrb9
Aa1ktvcfwdWx5msKmeN5TGf2l1DGsBzZlAEu9QfqVPiq8G5pqzbsJghYRRhJ
/Q5QOrwSyvH72aWvtEK2BIjkKrTYa/quvDqKgD0EZRFkJeiOwETAim+KphVT
or7BctlCH/1i/C3a0ghObQqTEaLej9GmyC3JZqzhfdCgKR2oBJTEZaG5M23X
GBxQBW7iNxvAvngpISwDzqy3hOD0vBRVB/LHGDW5Ih5f+ygld466ncJilYcQ
XNuXO51ywTKYuR2SEaxB7xFKmOH27y7klxwPn999JJKqexv0IgTYbE2D8piN
usRfdgobwAfXLObiixzENTFQXaxcn6R6++Ty6Gm4+jvdCasolxOeV5gSwltk
FqNWv9Y0X1Aq7Cxy5lg/Xm2Ovi6Up+ezI6zS1WsbBvkPYVTE1K+FIlu6owxy
ZyZebKlMbRTGYfnQ8XoRVOg3Apr/5BCo88NdvsA8Cqr7wi9+AAJpQXb87xcd
yBi/3mnvEERmvk3EiBkdHOJeGYOw9GEWFOay/fWBevXJkuHrj6DPD4eodiuj
0QDu9bG2Nt4oyAk8o9cLKMVN4iqxzHddylCXEivheNyRRWo+GqlRolui4x71
wA8JkvFexPSJ06PB238on9KFZU1mv+hj0agB0k9dpts9v6PJSuiolpV+i9aC
PGy9qyZG16bnvgtIIjXdwM0W3JspgqW8gebDSTmRjZAo4UXdR7Uc8e0HVVw8
AeXfJgO4lFtPnDJjT4S1jS0pM4RaaH7bABV9eW/t6vbgFUiwdK6ZgKUZMdUN
b4Ash3l/Y5I3AevtSRtOGbPKXh6za90mZV9xxyRLNT+Zflu7zzvvWHDbtIyl
U/jVG2r4ra3SblLQi+3pohOYxmL/awyltiaCrzTmPOtFejaolXUOtb2x6PWd
/LAL9+yMU8YoFKE7kvWQaagX6dmjfAS0MpdO16EQJVJaTBm/XnfnsTDgzSWG
8r476qhFB+p8IpkOwvZjEKxu0e/MI6770w7F4U06FiV/Nr3oljIxpNocQ1rJ
vRFee7K/mGj1AaZPCZo2xDAy1Ow1Y3WUyrtcaHD2iCWjVRmUwXy3hqi7vUi1
+X08raY/2J4dAk+pSuHuqLawvZGf/1UQh0NJit69ZZ+pk/F8mo9W5iLD0TQL
6gBkzysGVulbt3ZO5NgLFjEqmLn+bgO/Iv4HdiAuMoncvYPz5cUPOB9oJ7Ub
phw+yV4rs+7xl8mWIAux75PKZR8cVuDVPq8hKHm6xi+7HgWe2nHHCLXANqNw
r6hLigyuo26l1BuB024f1w30rfvzltriqj4kiYipdsVjgZaw086OEheWMYus
M7K4CVoRvCxM/lycjmQG/8kLD7sZeCkLqalW0yFUO2hQPBEYUX5qt+97sHKH
VOl1DhDIn4hGh4MkdOFA8vHeUFnv1W58ErejMM1S+IjxUT5hzCfz7FuQcQ8x
XXVlYr/jHSK/Fij2XKN53TDtz6hQgOrx+kfE4FrYnIRk+fL2Bi46FKYWX2Sb
DKDpT7xEYmCG78LJQgr62vo5Gmic6HVEBzkd1zzCvsuz5QjE2+bH0txuAMNB
LLVaHnqwXe/+yQXs7lmX68CfwlXV63J8TmBRgtykz5/88vzxJwlqK9Rf19Zt
T2Mplhu5IJZZV3k4dEEAi6lcxB0rbW/+cXB+uLk1SbA+OpWxcrjCVFGXnvLs
2PBOyUEVdpuz3L+74HKFRqcVEqA/Yx4aWhesQOJNu7BZ1hgBdfgmYChzZMBB
88VqYrSMBJ5AQMO5+kxn3fiKHnOqJoCD9e891FzplBgxNbTO+DE/1hVFlXpy
WslCOu4hNmspUASJ4tCx5sV4pRHE/LsdnJRGC6rc32q5nDH8cSCdzCNMtQ/w
ojWFSjH6Vj4zMZhR8hI+gjVVGLIfybTLejxjOahwZ3Ql1wnXhxo0CJNrc1S+
sZ14piRJ74rdJ30KogGEM7MWY0ZCty1QaLEq7h517TAjy8l8i/cCVqt7IuZp
RmocZpe5JHcE4IUDLhEdCcuX+cxuODNQtRIAu33xUFnKNE41VzYPwbowO1si
F2D1OZKBCHzynVGWSmmZtRTqXUsrzbRmRUHgffeDD9YHo9aTNa2vPc8chlOi
AZtwhq6ELDKcdcct8+6ytepMb3n6L2XVQDrWxOvzX8G/mo7Meq5AAvzeX8iB
3YQVkCnQsF7NdYgSWumrysvkv10Bg8bhIFyVTknza5V+IRE59kbfcmo+TbnP
v3ILjd67XDqVRtwygLIk85vZYhNMMOHTIILim6Fv0h0r2iDvRCiCz9FFLMcP
yNlWk85rghRWecmVHqROx68MMm8H3Ft5odNjVLayEBk3pEMEB7UDBEuQBdC9
emXpa2b3MjD8FyDMNzJXTVZfId1ZeBmP8Cm5E1ppecZtuDafS91/ZTXt75uv
Ct7Cj4nwnZVwMEVXDYK5BsUudPXklGiVpDH3E9N04pbC7iAs0RgF8H/adnUD
7KSxE2J3Wyx1ZAuwFyZaal+xF57OP67kWQi9QlXztbWh5JP8tFBzgbPhCu/+
pGZ8IFkDAlxnNbYhYEdd4qxUQJeiVUzU1V5Ed8WgNjas+j6yKWtJshaXqdv9
cuQMkigaOFMFAYQjpkshcdaDmp/ScsJISRz3gnl+HszfIkJiLVCQZ48SYe6y
rNP1+6lPfbH8cNqbEBlXtkxDMvLgp5fDoF5cDml8uwRDKNr1xazJfPBHUG5K
siW/QKp40XKGeYyZw/ir88LvXPmcefu063RiS7ljqjM7oAwNV5TBKmu51czc
aFOaILEGrSE3E/bVYWd8UHYgONfo/6JSbTig2Nnf77tDtf5Hul9Aoep8GN6E
NrKkobQBwuPgVNPBQdOgBihOo8ov+p8pJiiXXVkhEXoeVIntIL4mAnhnmmbc
elstnT3/V3brDfCoYJXn0gl9Kh942OBCHc0OQ71mkn7LMG3VaU3RhOis2Non
SH0icJg1w8027wcjuD10bGgeIcLiPKFkdwC5Jl4/Q7QcKtAGYj+vhbufdT+8
VJhl3v82q6r2ZUWz3y7OV/k+gZYGwVu65KrC3Rs2q2miuKwMTwY/LSUv3QTi
R3YhrF2OheNzzOzCbjBcmPQoSKJ2BfW8/aCTPNFG3BGLPexK8LNNaUF3XsA0
nmusfjAPRfQmrN45Xqjn2yP7pvMWh4ngI+hmrhwsQa4LHdE+dnNEOvAkNoow
ii4MPkAVuMQeD/fFgzxOLPcXg5oc8sQNsRsCIHmPHYp33LGWZ1m0f/CEmdRT
7yQyAC2Cu395xH1jGktSyqpHP9PmAag1njM2G7LOPI9eB9bHZHj310RTTDgd
Ws4NA5tH9dA6G4MKPtnnnf5hpArjyCMBaP+XsxdpvqWaBDoNr+crN9wYSQj5
EfYsNmBIp/YR3l9ci7Cd02U39BFK/1y7InI+GoOvA0ayGp64fU8kZPpZefmD
Ee8mo/b8ov65Da4vxc/RFwWGnoSnE2kLqzAvTeCeYwTiqecGXlCMbqKJzqdp
HAmscM90dwDSjzsIB+4galCPKkPwkip8j9LxG00TrJuzNsah7bbNxEtU1Tci
gXi2YpVaPKhljDbtMQY5h9UO4ZJeoUBccI6U/f3HezPuMHjgtNOIV2G5gMXH
K+GINlKimLIWM3xnD2ZCViG6PoUNBaxKBrFbWjhSXkG7HlYv9stx9yw7Z/r6
WzVkaQ/frKatF3xlkFVLklEOaBkOfbfzfFs/5Bcd0BjZS6cntBQ2kWRNRVUJ
Mu7HgWJSllwkMWDlQrgGFiVdhQHzkneFieaUEX9lXfqphAqEsvvg7tcZjWU5
anB2qSsNbVXo9bxyMHEesBAGqc2jxLiq8/6OEBvfcalombsxyRt6gLAUhycn
o6wNfcaESBqtYFKQOUeuFfMvA3Mse2izgobYNIg76BRsD/S06GxW/jRR3QZh
tuO0NtCFDPgjioQDzHZxP2GHTJLj9x1Wy70sRbXcggPwT+9rxGvR8MdwsID3
/w2J/E1KKO4UB3ju8HVcnG9Qi/pIgBGPyGnPRVb4hxrTZNgGWFysw9csdUU9
Kh5YRsVUzscnA5Wx8mQMiGa+ekllvQvY6pABlJb03ESO44vKx+2Itnm1MQEi
1MdXAWMyBUa12L+A2mYEBMpT+99t6iQZgEcrJNmAKMymlVN4VGD2MGgs4fL3
rjHdoYtg6btrCsrs3R0gHgD0UV+wUoHb9U1rKuBQ0DyIO6lJ/9Wvfeu8eQ1+
X5PSfwdiM2wbO7lIvI5G5x6uaZ3FTXc1jkz8cQyTFO9NeRRbK58pNnmigm0Z
eje/zrpJsFrepj2tcO7n60qi0Q9O5CdQytOSrDMrbNKlHkVO19Ou/nyMesUU
uwMvna3zxMFApd37kPvmt/IBgmSZQSTF++myfsZmiyytMrtyC2ZvTWnZX8bM
p1XB1NNJ2qofDYfOby23302cRdwtbwD6Ev870kkA7rA/i9Ufusz0j/dS4iIk
NF1D2yfjb8Px9qcm3eVpYX6m0OcqLATC6mZ3jvEx8OIT9JlcmkrZ3L5/SXz2
4FhsuhLxZSvyHZC5cux/gFC0+lKObl7j4gfe3gxYnSmtwl3zVcYoirJ4E/T/
4swEKHq4NiWc3MyVi9G3vqkMwnAdn+f3jG1+WCdCAS+yAAgfwItOvm5Zjbzc
Jy28tZ4m1GRuZtkVWly+lrsXOkRUi5gK4ngmrRYwp8QflZR96Wy6zQwXOuyH
SouCLKXr2bfW1jiDOZi8K5D+7kL3l5f1Z40Bl4PkmlLwv2wwY1FTvk89K5vq
GLWfJW3uPtrxz2Zt0SMIeylhLg4f2pSMEqMiJFF8tgRx81cQnpej5ocB/q9A
drCdxB80BAPKXxddj194vVMH7BRMEP78a2u2Nu8cr/3yXc1nImIzeqwZaXwI
HIm2TqrYVtU6tQTbj8P1fo1GlAeQQLkMxoFPxFgcjZrXUpXLeJMnDXsOBdCr
rOfha2c5P3mmPtgIBjXkkOjWTsASz9FegHTJbObqOZj6qdSBcvNekax+vG2A
sXxfxR+hr3Qh5IRZnMWChnEB3O7E5HFBNRPtnWz2Tdp1GBDdti7bVsrc65hi
y3uB/OR7H73G+6RroqTnCjk1+L23SZBMRVRhtIiKyNzhZFr+OlQHTyIf6AhY
3LWX8rjBWihhZ4/FZHeA816YLVehF/fFnoGHQvgzePt/25nNDpI3fMyi62je
W1fhnbauzefd0omH9LsTMjlNrSpKaBBsHv/f2s09Z2ExakYxZfviskzijbUq
QcZyBXrVhQexD61RWX2OmzgsOZVmmpJTJB2JVx0/3uGYmSAK4aWC7tGTteTO
6jxlzOFEoETX/e3gNNZLwbHkPKzAFhohiQaXLGfKqyW+T5bPOJGFTe18WXPz
vkac5JgQk90JE5vcpHcF0cvsuOzJzSBkArhGU0z3r++KgUMOSVojc8je4OTH
BXeyC35VWqr6vUU0NqEQOJq7FamFTI1yFAVkHQBb/MtcXQHcOjsPn3MdZcOj
ibGPOPupdUkZuMwc6cmheNP3C2qxFxTVzOC7kKnDwWbee1SQPn1FIMPtAt7V
cPoJHRg5Nl3gAd1HI+nKLKglK1d0VLUt31qWJXvqmIVBZJDxOv/PpjfUY/iM
XVOcu09dDtSUV1tUjGRDx/ayckP60SRkTxUd6A1w2GWG+RyBcMRyPqvBhMlj
/unGEyNPbEHRb7qjcfJgLWRIbhmjqhtsPAFLQfRgM1eJA3A+kXcwqek/lFIK
1ZXr2VniGVruiD+/bBLtXCbVuHZB4tI+YOVtDU5OU0vqZDl4/1WPfJUDUeKv
3Yng3G6QVkhOi6wrVnbTcSPquNOXAq0XPMXdE8X5ewbMDhfHFflr+7DwaucR
CpVcc/BRmsHwUpOIB8q1l18wiq2XfvI5RYjvrlXnTZvsT/bO5CyZ+eqAm1VR
GrZCz3vQUn2/9lVsDq7FyfqgKGsHPvaPUx0eWf1DugqePpf4rWQaptEAcYpr
rmanIQJ3Dt7wE2z4tjvulfY/dzLlaYQsRpM55w0PAqtGB51xKkRcY75bF3uW
fM44quxMct+J6+prAss7zNYKKkChto1W8QNzWM7Rb63qFd2yORwCVpfnPrN1
unL4xe91vttY5MBHXfPmH3i8AZGxGW2EU2t89kqbY8woaqU0mwKPmj2j1HIU
I+MQBIr0/kUkdckVmUA93zTxpdTFR12cX5u0FCuTt1FdN81zYAEkgTNKZPe+
LbcfEpx/qY/cR5Rv4EZwT7CV6/ZKQY8QuUXFu2pUyVLy3jCCD4fFKptpDnxT
sw9giE6zxcfis1QTfntf6Sn/pggVQkUveu/otJfdVW/bn0Vyvbl6wbzgKC70
qMtXFYYTkjQgjyqzFm1VVqCHDPrcx+ShkjxxDENzxi2lEFuONO2tFHS2HUSX
0XBCej3qMEviR96jWp3EetzQ7Llc0BorWEPsFkA2Yc333JeeFXWGnU4vZV1x
u0oJb+rxJAFUYf03Dk/tkCQ07Jii1PfgNt+5PCzuebn0JldYimywtcHdLK02
2urxL05Uq/YlG7teuazXrdFlx3C8D8YM8GPaMln8+qq0xQombegtC+T13rkg
jEybie4tTxCa0FsRbwrIkGzyRAhQiirpeGM3HTAqaQDVMDQcE2s5vvJOmbso
tSiC9vs6nsqmgUcKZ1XJw2PG1ELYeQvWxo/X0Bjvb37EFfJlmyhhwNtj1GG5
IBoF/xpzqEXbL0titw2ZlRpgXzDhsAOgdAuMNPH4j2lfKTpt+t7UHBW5+Qjk
tvcz0EkXlW8raphxJdY0RgQD7mMWAn1Puh2G93qvaDdPo9xzoqXnixXU9iky
D3e/ROTYgcuRYtpSYZmBCYYzmoMf89QK/IprAsbXe3YbPEADW8XN6wzPkEVc
dXSQYKmWIjaAscE9K4NA7lOAJav2xM/RBcklrhJgKwKPQvcLDTenI01p2ZC7
Qel1ijS93oza72knp/SyZ0FAEBnTkp95X2ZQluKcLfWng2iRcMAJGcg0M+fs
WwP/cAHgvo0QZF3yEGnXN9FHbW9YfO+TyofrfO+NNHJU8yfP4VpsIQErUdYQ
btafPg87yfObpfYwrFdUymDkECQ4AXjJgrPQ0l7FvUx4cHVrHzlZDMzYie7o
OZ2AeZZ6XlI3Qicg09SZr5EF2z93umomtmPscqq8CobTNLwh9WYHtfNj+Idp
sZQ9VsU3rNN6zvK3DDnGhA3eoziJloTWKWCmea4EqDceuchInrBI6QFowfHI
OcinkAawh3SqlXDElLp/aZ5w5N2aH9jaiHanDOXd38z8LTH1F7LAJCTgZfTM
l7cjgFJhKmaFoar/OHLVRWNilRbbO7/hhfUL1+W3/T+/+DymqWx8TIc65LqX
/hfpDBMDmLviPAzHYjhp5WtWYGbEeNuS43D3hY4CS/5Le7rTu6Xrc7+TFNLW
9MFmSJN8+IiHR55zPPp3+38foPIHnRvP0qBVnqi9y1m83y2fvRwtTpiWJP0/
oCcEyNJcYeRssI99A/MVFVWYkK9bpnxQCDA5PJm9xZK70bIKTNY6kEtwmzSS
M1+LubmTcsBa1PDKG1KE9XjNn5yB9GNuTnSF5RwE+EWV/pZzGy2nMy0zgtEt
zInO3kRYrY3Vta8U8ylrWn2rDpEEzTXVnjFtGiZM9WKpK2cjTidQLuj54XXX
pMLUAYTc+u5ze9suN0rehHzZ3ps7tbzuygeHB4rHf1INPp3HkL3oNQHPmOMZ
0L4ctVuUlOe8s82v+N5hEJIA90g1FjcEaATi7267M59IMA1TNbxGV1mb9iFk
d1Ab2ydvj84oyprW1R9CwCFZzKNk0UIKO4epk8kHM8gv+TVhxOXeQYRD4yt7
OtXG8krpP7cOpU0/oMvULLfqioum///2N8lV+3MVOKIAMCWshlbpQ8b11mHO
LrHuPsqhY6XiSDxYOM5VGKkFL5U8mC+cDs2C509VLt1neSAscl0rVl7nCREE
kts6riBQAs7sQEKyXD0jpJ5qO1fhGzo6P8rrMDuzE5pPHdIgZv17QO1E9aWL
AEbXwSnrxXNSFPpf6/lqssgV5zYu35oOJ6554Luu/tdbFxD2EasEr5h8UbBb
rkgXiOqagKX28Nn63D4e5sl0O+rEamJGdqlON8sUV8s34XooXBc3kR7r0zSc
QfWm7tH1UMv6aF5dUlmoXE/2+++8PGpKaBCFNQy77nhFmriqoii4bKMpId3X
garEaNb2P3eVQ7aLW3zwmiEVcBPg+1Fy9aJB+O8zKCHfxao2IukU98grythR
2Zg8SlEyT3rhSubeCzxxtvJRW7o5LJOSQLw9l79STT+8UL9MCPe12Lqghv6B
/mtOJKk95aUwPamMvFTdTSd++zTQ4B3TyMOl2VKMF8wRJl4ac0hsXoBo6N3p
xm2CE66Ws7Nq2loCiZOb/yixj2hVARDnCP+WSCwYz5a+eg6VQ9o/xRuguGp0
j4pwnTcuEaCUrUK1A2BMzyYxkZjBvkw54ZQHE9HfGBweuzbF45Fmv+WSv5FD
TPasrGRFJ14ugZnznCG+CfXwDKQXFehOLTKLGSSJxAs5Ve+Q1qnuHMnKZ7zC
DQH3THSxLzQQRwHobjsIX2m5yTSgk9KOUfh1mv6dcAOKBTQhCqoVmIW8jqZB
kdz1HklX7ze8kOZ/60Zzzv9JAzoPGDEBW/PFeRa16KRzU42tv265EJp2sG55
WesvaFtmY+q7ufM3Yk1y4+oDLdZXHvulT4FKvPe0b1aQK266zq/5lIdJbnFr
9z5T7LTtqjAw96LVZX1oxo96CNwjNWti+0gT2cIpaRGgG3LDKz1U5t4TTZyJ
oE21r8C/72J7MDxdp8lq+EYF6oY43gXPAWyF00RT+/A8gc0JNvdA/SRpRsVn
lk4YY9qJ8nMNSK/IPt4FbHTlBegZdqKHkSWkOkDbvEh1Dtodry/oLxYnY4C4
yKZOVEzSO8x5CgZGyKufFtiCxaHtWmif0+QrOU21JhdL4ELeoY0CDhIOLXRr
ID+UW8Q+aCD4ADztUWijfMEF+RLxUCaaHTm6oeG+YNXBiS08bx6YtibRRPPr
rUI7gjE4qnj63TIYEC1irmEBS/Q+9F68M8XPbNdGSJfM7gpKF2kh8ucpe4fW
JRy2KuYR4kGxDbikuC+5LxeAx6SEKfOHisoD1/ZYKmStNorKGQo/X/yQ/i8B
fM0KFknw9MLTpfgEa6eWwoeIB48LDC3TIY74rgHBBxziF4DEqtvTSUFvDvBl
9Kd3D9Jhscz2r/uijb+Ye60Qh1Rb5qaN8ES3Uxnfmaffg5yTfpTamnCrf7K/
M3Bgg1ByjEjcyXZy0Uz20PmxbqM9xOhCZEj7qkW7aHsqBzB+3u8ZOb2pkZkg
gm2HGjgJ/1OIX5N3fPxMdoTfINVBflv7d32Hi5E+EPRz+fsvTL7DKqlwzHOb
fS7nY+fCMERS7DCKhBy3eVO+0/UyqHK24GVm7WhdbpM/k85MIJB/Lltc1IOV
ZeSKULh/zaA2++HE3rsjdL1uJb6WuVOhh73X4zJLWo44/nwdZ9tUAJuWJuf0
0rmORc0V6ia5rZKj+lbqRW3EU5dWX8Q8HWdudnwTbtRnIH17sWxSaqmtKZGE
b758mbwUnpG1mvkvK6l1ew6nwd5uIAiboSt6MvFI9f/jDTfbrR5nCJtjghAY
VpgjeSHTxdEDEWAchl5ZLWHlaIALOXS8BVnN1Qja6bJUszBGVSOraXw7j4ov
iJtOWFcNJvkFeRcyqOlwnAB6BoQScFxp+4KoS2oLG965BXFCIhpMnqegDMa1
g5NP0ZTQTlu0PeHi0dzfXvhLahihKTraPh8JkKkKvv2kOn4A3oCIESBHHF6r
IM1Fxf0NipcqO3KJs8XL7dsaIhHc/vwK2Nxki/Of/A/nvLw5CCes16f5ZtC1
qJ/zwkq/6KWq4tJ8m63KMjv0lBTSJC4XWpHA44nvTS/DlRzAx7FH72v+flLQ
l+Nso8D9T0+Ph3bGVcwJBhiGGZcSn+whyGgKCBeO2mJ4xjtmKrbWmDq/df09
B3+H5JtyMoWrSS3+Zj7/9IqZvv6l4TKip0VN+CeeDJcsfGQVyujzhgVjl6jf
DyKloI1ij1ukPgn0pZaRmCw1tKNs4VDulBBtDVoSMnz7zc3PBEQoYWqCWKPV
Z3z6lyqHjTeLx87+shP5mZVDYjerLaDXwv+T9oze+ZhmFHFyzw+ubVn13/uT
EhNwV3IuwNSq3NsPAxm/GhimSK5iL27jwaVrqxDJ1tZxMstJ/D0+ncgLNYbL
Zz8i2U1PbaEXNWkCoMSX/mBdI+vHDQBimvahXysz5XYfbCA8oN7hHDwCdC8l
DN5mq1glMXUJ3lMOwZE3EsklwgsYe7tQDtLY1e0g3Ed/HGpp4E3TWWMDHqks
gMz7OroRsoESiM8cqi2NtKoypHJq5h0SOxsDRrF4nIox54ScVM/meSS3nqiX
2EntkTML0YnWbgWHsfBDcgRenk9NhJUt9iNGnYlHHNCa4Y1eZJ2smHscqDK9
BLiFSrkR5G76bsBvZeVlC4ScD1Z4JmKPgPGZtKdvSZCV6UqOIatTsNgfJNOe
GJjI1Rs2GinGdn+DwuGnkbOb77Vb/fSZiDHiYkijG2bvgUTz5bpZgFXWkJP2
G/1ZytCSnpWlcmLw0upyBa1UYAYAKkOpqUunQ4DrIYtRXVZKaaMuDu/iWdlM
gMB0LKTqqNwK2ycqOBk1JdKB4qM3hvQLi2QtWBELxi/rm5Ps7BN1mvsc1Js0
aWgNuOfFD2aYqtzYE53+jUxOjATbkmW50kkb/B8w5/WJszeFjC1+E2Iz6LQ+
fipEfN7zcF91WRXKpq/4vccXrbbI40Jjyg7fhQK+FfhfyLuUZYiMG0k2KNCg
jK5SruHpcsV3hhRhP3gWPuAn7NolndNesl+WFOV+I7y1pqGQ5nBHJOYXoGbd
OZcADyXuFa4Xv1Tfx9Z4GBZkNcNgW0MWQlH6SiJxdmdq7ElXXsXYjqYaBYnV
7878/lYL7f4uMO8l9I677K0BdMFY7i68S8ePqsndDbu3O4fmJ+bpRew89QhQ
zoqrGEaSD3+ngzdBnJjrPl73D6tDDd6qFwLfdRlN0upepHDuufAeMnK2XC9G
+X52mP57BDkosFYFAFt8vEEwVp8FEo/unDoDycRxLHimOPvqhZKVsAi1n2jV
GEarSKJk/oV9sb7DwdVL9cpW+Wr8tsACuj8kjrRs4Yc3grdtXBxvCNJgR+uL
6S+cwCWNgUEQnwtfb7CO9Ph6PWz8BGcJJ8hONf0aH+cRWdPwKx+bxxQC59s9
gIVi7FPPZsg9MW2altsttyJQ0Kexn6ebhaZ0F2Te/fdqBx69jrj8sJnQHtZ/
pAv94mHj8ZPIubh5iyijexM0OSgTQDsRRTPPZQR8esL/u5xiiCFQU0ZFgUEM
trcAaI6vh8Rcz9eHCUM/SfwBQPm6rycMHnSg3HmscP1lGTUdixPjGIT3EnGn
Wv0jCe1UtIJygwru/MZhY1+EMLXLAfwXjCe0LvdQ5J7kwMex5L9TwCKjVcG7
nXivWv5qIu2u8rasa5iWco5My8gv8qVTbFO6/Q4LmO7ddGnjlwhgIvnKpctQ
iS1Ka2xYwkmchLcxZbTPwOju9pisCXZJKVZ+uGZsxvc82vvuKld/k7848455
5iSFWbZkd0pochbPGMk9vpymD96oSiy+8DQ+PsPkT4pk3XvBhNwIyak9N1TM
328u1in400mk1idxWdfYe1TOIwnaFT8wvvoEudXdjbwX/yvQvh4seSodE8gl
I6v9zTpp4x678UMvEc+otWXEoBRvKNpEuYkiUtErhQOnchMSx1Q7MG6ANIXv
NphvBpHLVdvvx8HbE3QyrCIZ275fWJV03PSqc37UoAn8FhdvVDCOFOILdxOF
eJx9xQa/XRhn9UUOpKW//1GIML5Kd0QeOLvUzvRnb+TTdPFu8WsKH0z4lE+D
ap5AupeooQJ6FXIrD8tQRfegZLD8V7WWIB+hU33+qdyBIyS2lUBILP9cYQTC
ueJlfCejLpC6mXsUnF9L/xYcpMwk3Ay7XMrr82Kj6IauKV8x5ztOdrRk/3+g
bBpLFxq+0+IXpZ0i7vbf9ziP+gsHQVZ6KHsytUbp53C8j134XsW+/eWkIIgB
QTsSBcx8VRcf15kqZf4VH2UXdbUTb3tWlhhv3HlufVb5HNi4tQXe4PkeYbtR
gAyIy+OeCrtwTQ0YqWFC7tVonnvSJwnTEt93daEK1shJeD4D89LZ7sy4Dx9P
rpmTWUTAO04v76a8q3ZKvqSD8DomhzE7WJ2S6zmFA59CqACfAzweBdJpgEC8
eCp2p0+npzBgXJ3Hg3X0GcQIggytoGB6us3wsZp5wGLZTRZ5SNedTtItmOyC
7T1b2OsPyFbprpvt1NVOoLLqI9JlEA+/HZYX5QdZTCwQ/8Gm8LQrfYTC1iVh
V9kmzcQDxH2ncVFMT9Mmuu7GHX4fTcpifKgQbs3NW5bIGtKWMQKdjzutRPBk
qK+ChZMQnRSQLYAV1Ixm7nJZTFuSj0EqSWOgHXwW1Fgg6/vHwNJlCDkg28I3
Wc1jgHLpbDh8msLzL9r5GH3IAFgI0nbw6ba9G3gb29lIxg9rU+fs/S+MBYlb
JgZYEw2loJYXd1iCmuITo4Nrvrn6gPd8qvSUli79E6UjujzdMCh2fywDrutG
Cy8WRZtQk5G4DqWP4pcLfEYu3AaL14mW3Lak3h5Idn3tWBNCn94OXwg9UNXv
3kHDevIKikRKvExvupl3jZwQmLQ6qhflIMtu1IoQsQ+bU7nLOdtShaRxMr0C
ZhHNv7dFO0HZFUabdzTo/pM8tPt7EvixyDtOKOVhpp+c9ry0r986WOgPH2kE
/E0EpNCsggnzNYFm3ltFmq73ggUfeh4GFSz/OG8v+4OM2IIkS6Yb4tv6g5Ay
3iX7OASXm94FRz4SGYcM0ezIEv/s3ZFqSFatn35vxbNaTTSmdk3l94sfKr+4
ONJa1UcahhKjIUK/i1uTE5p/d7eW57bv4E0ZRpz4WFRm77LRo8DwSxxvEA43
sGGVgN6NevbqAnZ/owBwsPAoT10r90hAJx7be7Nbi6zGWQljdsnBLjrpGxE9
mb8+fsAD0xTFUE7d8w7RDellCzXVf/ByA7oV42ggWqaBbJNEGx2bvllsh6Nd
LBg7MPAbH7lSV78jHaNymLW7JoJ5f/syj5Gw0eAiJZ82r47afSn8Grfit1Xi
btjxh+5ewVaK751nu6SZrgtfealeqCybrSn/HocZK4w9tky2xID8CYNLYq3S
fHbwrZma8AN26yPjembFv5TMnJdISii2j4SSxYNN7Aft5jlsDP+n6atySX19
vRRZSOABD//dJgT7Vx0Rhiq3t273YB5+Vpz//ZLS5IeYKE51mTaO3pnTQU66
w2tvtIwlpTT0gbqk76U0BG3r2/8neZe/wY3ScryotTUjIi9qGkR4cqV0sE51
rpMHMMtp/VVgo5NZ4osxxHOHB01aT/xOO8t6xHkWH7tcaxpwH9pRZH2n/efn
zhJXvqF2eNMOdNXUwuP34PGpVFGf2PXtpKDpiA5qa2NV7WIF7I9veRjJtK84
RZuAUMpuchalVOt61vRxtB3b0GGfk5pcRKdnckcvn3DjiyiQu1pfCpY8oI3B
YPAmpPWj99NImACA1x8INlgKQCXVSoQVafPPR1N/woufxS1kJLKzx0zD7AoK
aoXNHYiTnrG77bnmNgOaebznFGSzqTkELhEB3eqGuf5jIyxFHlyKP5nZk1bT
d7Q/Nur4+UkqMW2f4N4+E3E6nFNvYlTD4con4trM/ZxXyHVqMPWk8QMxxlsf
GqRiACR8igJDcK7+dazzlEjqviY7jtm8k3O3z7pnEljjfqLZJz2dkT4Gsnp1
+TzPGbTXAqze5QaMRQeqwmD2VXs3OuYZt9ELp+b4VBG8LUmere2q5vNXpkMG
p2W6o7YpdayG2kOGwItNBQzmHStS096zuZebiM2vJ8t1qQdz+PpQnJZPIglk
vZ+zQYXUOLA1kpsDvGQYF5Un0TzZfj5OLFR6DNSMbPUlZHr1KYTOgT0hzbys
IfcjMepCuBQmIXW26OUw0+oOeskSoTOFrBjBAPMvQCmkTwFO6NFjvMXO9e2W
ZAX4na1u3HTqeVzdfEj08orTFP+KZBsP+ZRUKZ7WIgH71RHzBytW47J8FAbb
EJWf7M7lGOYbp4bXoKFtxwrIVmW3enHXejmKADBp+zZPdqauzDxkBX+8YHGQ
5Wx37jYwLQ7JBPkPUJ/Yhx1V25LUXRr966440y3H/MR+PxYuDxtUsgeMoIUW
c3ojUnCETvYDgCQFC+C875CMRUrnkQyOe2oEy3CRkhcLq6oAY2AEp69crOKz
dqAW7Ym0ao4/WEnWDraL6DrdGrVHpTpJIwwJAvFZ/nl2IZp3hkgI66geRDlM
jOFG3/ntxLd84rN82+TC1EVUbIVlr2unxbeRVphTU9z7418BKsjjclhDpPj1
D58lzlsHa0XfGMoAJ/hTw9f0oT0sYqFg8cmlttTShPf1dhUoYIyd7lxMTUPW
SsoYXZTFWSy8yWLWO70kqTivV2freFv3h/ZplN4nT84XwOBZBd5HfAr5OlaR
2Kl+WobM8lfzGyYNlxTU32U/fWJ8IjpZIkT4mwIGF65YNMMEcbTE0MeZOFex
06DT/pwPSLGKlSLHQeWwQg+Lk7JVbOLj7zvX3LDN6mXm4E9p2ixTj51lWFGH
MJJW3FzDOiXq4b5ed2vdmnKE2xhLLNrBp77Sedxg9GzIwfy+uFZ3b4Iy+ywl
YeXUF3ONqPehhFa5zHHY8iTOII2IFSjtJk0nFgo/5BPetLLPCq/OQ871HmsT
OLLx08HNL3onSTBaoel9PDmPm2ysalIETfx9+ESffUTT89vUbHvXDymjnGfK
pDHCSxyfwy91lDVjPc+qKwVyWq77Uo/hoxjlAuxOo6HEpqW4piPaSdIIPy5+
gGsZhlG0kzEkpExX8JJRFf4B7SA4HnIlF/t/O0TMPJtKfNp0qzGtznEUF1q7
TgffmC1yd9jFr9ZClW8R8loOQxEnsIDiTyPUVmbKsejtVyXQuM3rDhrycVrx
GiPqlUsnRSn18sh5R9MeJBJCamxQEPA/Cae46+yIIUta1pHVCKLneCV/LTrN
OlsOJe6tYYKYRbCTJdPXkN6P0wwRYn6Jg2h7nO41hkYF4J3zyu8YJJkcRpst
hQ0gMMBAHrvilwrvnxOo7AQzfczb4AFrubKJp5hhq5Em5M+pW/XC1jOuJcef
Fg1I6q3oNZtalbe5wH9/vBVlrTRLy+ZIhNqV5hSmh1tDCcLhUCGXU77otnvt
kDDm1u/21nTOJ32/lhDDK6xk3ZChchtWgPl8ykt47afYASSVoSbPzW3gDB56
AuZh6dlOJkxGN+6jIh+sFO33kEsX1wWRjkNitHJcp/HM48vVK+n6T+pVCAuP
ICJ+K3oWdK287GzBcTmoq0t61z4IPflLZT20vfun3XJxYQWgYjP8DIc9Sy/n
3Mw8GgRNelxCN8tsPCXxariwVxNoDQ4GGXJgfL2hP910VawvP4RFGAkC4Tki
qRu/XyJtZQ1H5XCjkcQifxOg0LTy3zdoJ0OZaUr4CkgjpzSiPdZlpizhzzy5
dWCZlQgH8mt87rY4j8J0k0qfwzGlhnjrwvrJwVr1wPzdSpSGSe33FNiAVKGe
2Zz0n1/KGHGHg4OfwIAN8fTIlTJHH1g4Mv4tMH44PZpxV/9ubyX9xNQbl2xf
isswK/8419U5VfHmBY1rmySRyRY4S3cTfpvL6qlG3TIGWxTT8wskYXUG21iF
6M6PEpZe3lJSr9f1Jz2EG0riA3n6GVyMTOMoee64/4wB9JPxQhE6WRtxloTo
cdORdWLmpJ4cfGc3GPYkhlNRcZu2LBqJSxU+HCw096uqZ6eaq4sOnXtIQuae
kLPDIhjnbfrnu4XnXArYr/Y//nu9J8eR7z7Xg0hmATxlVGtsaDhENJ2cPwzv
hQWjIRAXL8yq6XPvzQkDDTmEFqcfgUFV68LxA0QwD4LMp6zxyKll83+gMVuF
1777EAZHQW86Vuk9ouXXglV/DJFHlnb7sSO/RIrm+6DEQdtzISSgLxZfiVn5
UwhOmu6w1hbPvrWPdv6PGq/GYv/FSqdvz0woPIgCnAL0AQoKU8tkVvUxe6DG
kf1v/h1WsnNamXjk+6NWL9ITvXk8bwGruskpOvPYMHZyI4QgD1sz7WNnjSXo
7AvAxNQ8AhUXaaJ+tcX//6V7NtggRu1PGkL7RQ5NXiayo2yGGL8uMcq2Aakw
A2RLoyri5N9i/kOFBm0KqhbODPyYbpbY2wb+wpF4/NLRomwOlCEveEWXZyKx
6WnEY7yFEL4hk0At8jqV31rn7gV0ZMK3ddG6iMmhBEnYGSTXoo9tSmugVnY6
KIGTGdyvf3ZxcTQIPx7d+1V1t0D9Cf3G4fivxGRG90S+sHwE9xz8S0+X+brr
stRgyOjaIcpGOf9IZJGT28TwR6bF+UBnIpAx6VS7a928cBjCyOy5tZ5EfQ/I
lYnJnqhC3Vb+ccJ+v2dMbSD5pHsZ+/cn64Ma+8WJEWNtw15t/zlDYAYxuO+0
Uc//isRBJKhlmRFthClOwwu17uFdppb5v0a44YJyLa8Yr+ywSO3rQnQqQ86o
N6b/nuE5zopJGSCH5jmpq7Rws0wEBTJfmI5tQMHTLoc0aH6GmuAOL82oZ2uP
esKjjXRiPme4LRQ3FqjdLyPra+xkiyeuInwDWtZWXZG/iyct/J/WxXyMrMeB
mepd5wzQ1BcMRKm5MGfi9gv5UqyydR40e8EojQL2bz97he2uabRJNUfHnYx8
5NUldZlVxG3y6vBR/dH6k41YCTqrtUPBOnPkfcUhH65xXueCyg+ZYDdI3X/c
TpgL06IPDIz0cTY20vC9ehEb27keS/vZJMEsa/6cnOYlVF+9d1Qcjlqoyro3
609aPFOXgPq4aQ0LP6WU44EFissMpepC4+AtQ6/RIhZBUYtDEIAD3ACQQ3Wv
GXwOwoK5mCjazuhX9R7HfwM+KZmTnXsYJ8z2q0SwSkPga9FmKxEUtyILedfI
jxnsbwb52QE9oMUM6C+uYSWNlFuOmcz961SCNNNFMiZt7RAtTzVeBYP4llh7
FUg7z/875NMIXS1WJfbCppDxLoc3olHwqmgEZ6eS73Jl0Fn+Mb3LAD2cH40s
qDklVg5hFzMUMNfCoN23F7Z37Z1RfG4Pp4QUEvSJJzhKpD3LNYbUksEEmupr
iW8nVWvGLHv3n0FhKlBUcThhs6NDyy03emsYV5ql2BqsdrBJb7lfwuXGWwGk
9+0CdLuCVRx/UuBb6zEb2+VOMf8GIRG0TflmiIfeyKD1/eocyjqWVAYplect
gUZ4Vqzqsfvt8HjYITBYWmh1SlCP2MTGH1ZQ4MaDjVN4SJrFnPaUrk8wkS8U
AectBrVyDPnLLylM6pY1iszT01K357lGFPAZwiGO2p2BtPkcGg2pw5XrRODx
a7V2y+N8TV+vFmVb2vWmyo8Rekq1Rh9ZKvg3DAJh4KyD2QOY0NDrWx2y6tB0
rvYxu5NdLnCKd1DDD5UxA9tL//ryl5y/1ogP2NYjedaPq+Ja9TkhL/MkKELl
+w+aicIxcFY7SlJ39E7YZ41L795Fy/foLZ8YIY4rgr8zaUPPX69Z2FVpXe7v
u/4PcQZ/N2L0m/JBZMKnXUKrmfCc7lOpO77ZrCsfAXX9N/VmPffPL8PCaPs1
uJV5+M1mSM530EZMwP8YNc6w7MRlNVMfiQwnPH/aPfP/wMYiAM5k44Z+kE9Z
Wgyj0ZtaaKDojQY0YFJivymgFvjygPRTUZJ46T/QjtB6vZBLt9Ju0zDGeDWr
k488/Vb5/iaSPZNO3pX0OkbYA/JfalPnjKJj6heViKPwEOPx7Fh8HZnaS4FV
xjGviD2hl9DE6HaVi3CYvVhQqu/5FJG7+Of7xhuVtW9RG9TV2L8Aq2B0IzTX
IT5oqwhmALpFI5g+3dDfKtjT1iPFz5Z1uhohk0EbDNw9UUA//VUBkSPhwmhA
pj3HdDDOuh2XrKoZ6EeK1TDzcjEmUnYP9/ook9YW0+l0NJkcR6o/82YxoEeQ
RrVNCtOj2k6gOT6EglSvsIn8wbzypmYFAet/4lvl32grEnH5Weksph77UCWT
hhrDyRwMeYRp9QLtT3Rp2/uS/x1eFxgMp7o7IwtZIP9YhJMrqvPc9oQtaoTZ
Sv8IPGzXaGDAEiEA7P4vhDX7i52gTvrxjUOBWe8xUh8qCZqzY9oHsFY5UIIh
a7yUv3LVrS4l2skMgiEMWoIF0UQC9udKkMJ6G3PFGdFvZyZdMj7c96u/FFiH
gt8MATIfRjNX0zWouFdBHfeRFndEQe1Oe9qiHH8RkKAgxgqqoMxMmX/Gdwzh
K7ph5DmXRu8Pci7M/gBNss2YsI/TyigGf3t3Q1txo+OFUex8IYrGDooljS+m
QuyqpLe8pBA3vNkwkPbRjf+79xVKFIgpCIzRBKkkLXcU+HzPuwAmKL9YI1Hr
nk6eDAh3sdmOU/p23DeR15R6s4S3A0P4ZNvt4R0FGrNTY8zHkK4E9+sZgkua
KmBwLaGwcVW/+QQx4pusi/ERwZx628VPtv5HenKYl40E4icV0l3ncyD6FCxZ
iFrTXLeM3/Jt+V4epUFJ36//2AnnSQ9Cv4KLanGoJTNd4iG/OtKWbEYmM5rb
oBcSAh8bQzbTspCImLYB/jFB4pn1FJs9SUFwltS84pVUamjybn+8W4+u6joM
OFi/xwx8dn6WmfSgsl6hK2DiCYCLb3fbFDWK78cM777O8OrLP+82XL7lfer9
8ju4lujmJ2NjZysIvgEN7dcyL1sBdWPWuMVKOHPhQWHuzxpiTMQsrSLaMJ8D
1Sn6ymr1jeYACeaYF6WIP4KtGzzYpeNQGXNUggskbRgZz57xe6K8yL6XdpvV
gFHsNdf7sNJKk0JufnTlMAu3vN9zizebUtNRishC9b335/sMsfIFBQYacGsk
Uw2eIlU+pLicIBMnXVfNhjYe3Q+N7fZRtDO4bIzfgiXGjKLBTKTq8lToyZRX
UiUIyFSIHlxHnonq/iRL2EeEQrewEdRXHOgzAHIrFEh2a7Ajzf5Z1t7wohuB
NSoyvi9ziq3o5Q0pUvPnxeXRRCo0v0ZhQjoDhouRy4nX2ik9d9Xs6LI7Je7u
CI9CbP0hcjEGR6IuP6AhnKPV8ROi51zh6+K0EVUdlK0cjOsIcviUVgXk75UA
pRaYAOWBAxIzN8HLTCMmgotqr3gZwvQ8VfA6th2LZ851jtHQnsUetLH/clLE
xLvnTC0/jdDJyt8F2TeIlT2PGToWbyPFwDnLrS2NXJSkZWr46aIRXKS7iHHl
0kb7ecO+0VaFHUSXTLntMOgMSOUNTHHj42bLWZQvJGddmTBMp1WZy28fe5jA
MkumyA2YkuqA34qrBr7RH5RgfRXvWW+FoIMgLRi4dloinonyZ4RydTWRcAtj
JOJ2+27brOS5yVmKaPPFBnv+XS6MUUy5fZd8hhuuQbLRyCgoWOdO0kYLlqDL
YeE2HYXDyHJS3mjqUKEoY0BL3yLT03uM/qTGu+dfBtogcHHwZTeVeKvIEV1j
G1IMlWfrlMbhnTHm2woYkuf1DUkKTsMY4hIG3a046z8k/Sc+Ttx36TYP5oq0
V+H3r4fYArConj81S02/pNdGGQrU5VIrqsGXbFrHx4iMtDrEmHBYGsi4lH/7
e4jQGFH4LdQAzxA3M5Vjj6WnbGRMcED8qhhQoYx/1lqA2LW/OiuV8tgMdMHi
VGbd1UWEsbm3y4eNYE4qUiEOY5V/yrrdA8ssdWjCRlrpZygbohHZWbkUjZh7
/bk8MJ0KmZDkuwsy7EUgDfEbAHI/DZ8Tu38X47lSIxFvbxEGxzJOZ6SHICpi
jtNMncSLTZwY5hwSrL+OYfqkXDDFLrRF/fVwVHJBiHCD0yHYUYyumYH/vnce
Mn+m8ER96LJSOux1hwVTafKpa19bL/oXZbHTFkcY5t2JXhoylHLs5qeJi61b
xE/pm+ct/twcrcQD0SDlCIIyFfvHEFu4W6C+X/oIB4Tueal71d8umY02Futc
8Ah9UYEc9AWMoWXexU5uJ3DbOFV7cnqjxhUi/Wzp

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpehYYU0xWwWP6iWH7WRNZEEORBkO4JNS6OAO70SdYvL9K8wu4HTkQg37U74LLxpZvmXtA29tY1CGyjcrjK2f3IPNQZnamVd4HCW9iuYjahhZaniluhXJLI7ckzxg6qJvo19F81wW4FBebuIA3H41oc4txdNTxNljZReuEJaOmRsW848O4XfYslGhL1f0827JVbmVc+QyxcvmJI08tYZ+fAcIYu00x17INcSI0OxvnlJR1UUNwBVMVbjgx2TWl5yMZgDIxcm6CdY1QZBxMkmNsc9Bs02gttjA6v3SAHN+GAGqf9gv5nq2riPxI5wKPAG5zP9+vVDu7rR0zLO2eck0JPMOIgTwKMEapNe/VCQKVDhWr7kqYq/J+WS5jQJKFjoGzL+9LA4/OV5VwejAcTk3ePoM7/fnASKC9D2NSTD6KHHTjFvbsCrGYIBy9dmwVAfg9QWPRA3TUnOeZvT+XiJ7O7+y2v6cTa9c+4Tt3JX68km80jv445EOrAncrvg4ROuXlC5kpxVagE3pxRyJ28FTK3yxxFwdUNRuCRpj/hkyzXN5iOayKl/BibEPh3rFxyfkGtGvfkXvnVWMM4456p7qe22NC/iqvBdiTw+iQhw70UcIqkfCYXZ8vZZArgI4iY//h7BiC5REaRmZkdbs6Q+qEF/ycClGiui0Z0M4ocJqzozefZqjENiXXGhK8IW+LS3icV92cSrrsMs0a4kYAVYEIFjn5EH6hl6khEmt9Sycj5MKeVnXGF7fpx1uISe8s/J/OHr5IdN3Wg6n5XPHlIL09NFF"
`endif