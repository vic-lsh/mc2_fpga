// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SNAVD1OmJMwwsCdl149T+vuyn/GRhFI+9eLqdOtYZeIwgNcHy/SdCxiT02A5
eQ614PzSxto3zRpMC3d7AZH0keJT1eKWJZO6BGUL1djY0oSeJxuTZKCqQuuN
rNtYFcPCxc4xEwDkYphyjQGBxsEmeRHHfqRM+WQyxDOINIhhq8GanQCfgkAq
4ngFsD+HyaMnpgQ6K7b9cQcIG9QaMmaCTaFHMCtnEyqOgLO7tH6J/yftNPgy
TtGjPtuVwFIpV8NG1oKNvh10Hp65b3u3c/JpPrn2V0uKB2YxJVyNDwioFQjk
pIYme57HmK7upWkZGu3J2PwJm+V5TCPjjR4f0MMPOg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZTt+X4AoEbAj8ZablUwxdHdW5kordYT8ntOI3U5lOBHjkd/ti82wJMV/vNxv
5QoakGLSECGtVHZXGYjenXYYHXAv0LReQmk4sc8XTNKvJTaHwherctcIoR5p
U1cFxULjP6avktqwFV5o5uMW4xtqufqnBzAYoqKWiXTzrfLph/mkZNNvDV98
O7Z+uIBqG8aHqAkoBF2x2RHTmqhfr0xBiwFfzN93iJTLYs3d1sjNuQpbLdPV
mw4Wl+FlW8Oacg8G2s7hDVVIgzTWCphjQ8aCaYJ2ueVngCYN4Ok1K15sgIBu
8PefEOLJKgyZgJtO3y0xdofB3LoMqRMqWxVmap35mw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AgB7DBxp1PTkni3QApyNvCpd3VOR03C2MynFNhikzPX/g8y1XpW5WCVkDFo0
KcTDHgwu4nFQLcIdeyXygP2CmMWXY3uqM0gQozj3VOgtYt/JXxYU+uGgLVA0
iarOBmsU+2aoLealZf7ggGB44oQC12y+TRySwlCn3t5KCv2uIFffwJMQQEMv
yvvbmNh80F8dun/2EqGEPmeKPbYi2y0LrtJQ/coSWcXqBKt8HdnbWr0cPLJC
DVwss2/T/hnWmN2TMnaAdLcNEJ8LjEKZ1dCAYlnHmvitCdvCXtS+uVzlH31a
09CeWYrMjCHGYijIFd/fSjwxtqJ3AmtoQna/BWYqyg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E4GYE8YLVbUOrcdfZE1Ay+hTCuj2DDV3JQDOs4La5VswBQoVkKJa2RQA90vN
ikFStDV9ukQQizSpQwWhaiiJ68qOgE6KyeQM/4Dd/PMpy9Uu3EcRIpr2Yr+j
B7ii/cBc+KnWrFGydzRT7t3FCKOwSC/ew02Vys66TP259yfmGzqYJ/zqUndA
X3PklfoVeEojX+CDdkO69/x7LG58gseaIva+LUdmHpaQ55Z0lO3q7e/Seo00
pq7j/uc4KTrK6h5n55bOsan/R4WhBQp/FawRESqS8yL9SArlGIbauY7LRZkv
UV+207y7Si9i6JWxXDabg0SPRQB/G7lbKa2W8YsKqQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qXix9nCl4NcIC8FkdyZYTKEmnTBXYiyRjFKvE4OQlabnsxu7gPaudfPEOX3D
2uNDgh1lx5yiVV3mR87hmABbrXJEz9hzWAeKHJT8zUkD728o6CII/pWxg9Ps
b87tKO0lBmSOXAWJZdJJbmutvZEwkpCxcgWK1x5SeCJQz3bTTe4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
gM2QWAlgFhU3LRUt0CMqZIaTCaVNlUeX54zw0DCIDWZxjbCdW6Hx6rTvaK9g
c9X/fLu65L6a96CBg0tdolsAIQA3w5vI+ZhVaLKD5goEbR8zH+UEkwPCS18Q
8C3AK7HigsV45sYjAunCNZdbgnApJHItyJLhAOni36nSmGC2abqaZ4QTtUyr
EIoiia3kKPzi4I31Oq/VFiE5uar/KSQRYoGPPeUEmeo3VC6THcofYPW/tmuh
6KT6sZSthCYTBuzdJZ0E8dCK2DGZDBQ18M/1+bh2RvbvHtIeQdTOBw2WwixB
nMs90KP/Os1TV4jjw5DBOFS+JAVBGyHDs040XpU1jNp5pT8xtLcPr1SDS8LA
p7aPImQx73nsADQx0wCb5uBHBU6bGisHYe2aExjLNW6PjDcD2nf33JToDWx/
ezQepIgultnwGrqHCssjejtLyuaVVJbyLfsuGDB5GngfiFf49I38H4OUyvIc
68qGioyXoRlUmLJ0ii2qEGkiqCfWoR/Q


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JNIxYiI9MBKxYKbKEMc2NwLIEkph99GBFg3iX9eykRGlysiMR0cne7q3LauZ
dlbEI8G+ElyXW5MGQ9n5EEvRtIOtvtWS9cQpije0cqa9LxIT8JxssAqGofA/
nnWXr9f/2udqK6e7NsIAR6MuTdulXM1ngefoEWOFlW+Evj/MDZM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SHpqgYvwokpdZXpnPpYQUc3aveBvoR/1nG2R+khdTeP/FTvnCRTRlVMrRxPu
pRkdXKCCVt2JZ3s8BQBIPCkjKpUe3Gi0PA/s1s9Q6v3heql75jq1c99ATQAA
qCDa1XskLXGIYE7tj0WuaHetz5KgLdUOotKWn7bVaIJnnZbe7YQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13040)
`pragma protect data_block
zeueOkpRys/fCCqWpOlvah5WJf6HeqTtDFmtYqrWc7gt5sATxBnpqbVkZbYb
GWYlZGI4iaPh4Vfi608aNu7MFvPEIjmHMYFB0GFB6aZtUW+pDSYB6ObwwHfi
9bhhjorVOckJ5LSYPcXMQaNrvU5svGtcqgCWifUnhmrmXcVW0Nht/P0Zhbid
GzLFiyqot3yjNImXnQ7nB4hBL550eg9kmAYGw32sm2lq1A/zlmFQnzXVgvVA
1Pnt5Ve3ijT5ZJB3b/OjL5/jVR1mcbruGM4BmwmVtQ4woh7uMXoML+7qCNIO
QyA+uR3IrO/nEYjmjnEzM2IXkVSVLHOTVT1wT3aSma7epGWoPO/U/KPFQuhP
i1NVMHBoCFNnl3CMMHGJNPVmPBL2dP+x0m0NRj8XJtMoZJSNFudSnorxF6II
FtdWV48PWuMzH4U/OmODpZFOAasNkiO+l/VsE8aHDIVWK+eSoqakRJK6J9td
qtv7G4L9pIPvTG0t9aTpQoSswdDuuYOG1GEMjG0h+unMOnkQxJzvprn2XQ4z
cSLRSvyVXDWl9OfF/sI4J34+dk6pSEyx+agJe6HzXgUpZjohPFebvEJrMogT
W98mlBusC2t3OXiZWgbj2b3iy3mPlTr2K5DMddv60dYhrAQuDwC1LlHkRAxO
kznrANWIn3BkJ0wGhyUM4kahgeb+dRHcAFP7ijw5v89Z+k4g0sHSQuN+Cd3h
HvcNEh7pDcVNfpiMBO0v0Qiid69G33Luq3UwoIb0gr2hFqm34cGBYMiPangJ
MZnhXoFB3vFQsmh1Re2GQ27vcGs7G38sWVF4RGwGJhakLV3Od9154EhgdPnF
0PxSnoYN0D6zJp0A6SFDYn8//WAbi9a02Glt+Qmm2aftLJcvqjOCxanM2Vjc
95JHgI+789zwjpawyH/9Pw7En/WLOENl3RyOutAsmBWViALCHy4TEglBYTvT
YqpTNv3SvbvLL8yeNP0E77BRWNqleuKpg4FjsOom7YbZxzOxzDxdp+LBzXy4
yzELug14EiOLLltWZOYv2bE4kWviIUmaM6yD0kYpUMqu72t0n5P3qmz/EuAO
K+3lOUETPySIQ5obh0uREpoRP6Yv+JGtbqeXt5Jz7ZIBuXqPRKNTbub8aOMc
TAUlEnzZ6o/XHfCM15INqF3uvxR/hvE/y9DX6cx48tEumVK0gG8bQIggJyQV
9jJ/PDvpicpXEMxojTvdC6XAMXO50SmiWMp0eZS6KWYB2fcL4veW7Tp4/i+m
zf/dn0GqrUUiIH2FLOgS3GfqAuMEUYFjN3AKW8pYO6/3ADBy2rlC1EpLHzQo
/zcxg8zqQ09kDaUQhJA66x/dp93vbzGY/OCGurJl39wqFHBF2u9vW+kR8tGX
DTkDd8xJuTd17NIuPnqlqNHA32codF97grni0fmAgKlWJpQQUczedwXqK527
VmjZVUa5Cp9trNsWQdeVhJsCFbcBKd3VldncSkZda4HaClyrgNmAbhLxrfki
CphhxwxBL2bhWAK63XpD8KsEa+rYN4BdDT/hMO9CnQ1o4MbCgznCLgfqlD6S
8WDqjMW0hEXBEY9GGrk3nqMy1CA0799rGFmkYPO/ZqIxThS+C5F+rAf68Y1K
v7JKDzgRFsgwvwlXtpCZGNvvcRN15fnHbSCi1k3yIMzBaXznR0AwLT1qrnxR
OZrJkhJQbxtbvoPezD9fMoFmofErN+bPOzl/lv21AIm9TkepQiTGoxcLrYmU
QhEzwB/nYGcP6oQxYopGY9fAjNbGcKuad7d2tQGUdYEyZMae+DCctIT0LlLi
y2roCsa27PjN4WcOeR3PAJQNYPqai3APdAXORXEDlQ544UiD6Rxv2KuSFCua
sMVQSiO763w3ro8gY7ExH/4goj5rrT7isNXnTtHSyxRdJhn2Z04XsrjjONHZ
1yjnAaRme1/2vnX1MufH4Rn/kKOqbpRDwxo+PWy8gP4ND6hwOowxc5Dhtpxn
gKytRmsHl4485LGRE+eOg/W6+JLinMBMfdN+duwmAfNuybJq12+MxxxgKbKv
EaZiDa89KDHkfNmg09S6PdTIl2avWGd8n789eha2VdGfBY2kJDxMvlNTLNOX
htmPK3MWhznXQod25ouOxYaIKbzRBxnMb9a6aglZADubRsvuJ+N7iWY6eV+O
bqQoe36iWPvtIOph/YWDFld9Aceru0YhPkr1dt35EoDR0wC1sjn4b/UZQ+0t
xwVAP2EUO/FoaxM6G8Xe9a2DQV1pzcPDTaudQdRckrbJstmpUvDTADIoEQMg
GSX5FHgHQ4aZTrnG7eOyJiHKSfIDzzm1j27mxJjSxFt+7nuI8thNEiXZZqpa
dGYXkUTDPpYMkny8pNPJErEGIePuPa9jo+RA19zKh4+p2TmB+TME1iK8HSSS
hWEwPGs4tFSS5x0zSXCFjjP5Yn3SXQnlLmT5t3HQheLcP6Dy8bOlG/Ahi/b+
40y11T2MXYNn+WqQW+8gnyzChtrZcZhqo7ds3C/lgwskav5NNBEczlLHsotV
idlkw5kIMRaHUUsgypiTy4e0yY8QfY3RftLQ6yFtpqg64si5fzX9lkV2QTDM
WEinz41q8KeHvj9HVUSYiE4maqSuji3ybRiFMJ/7pLesukU2b2CO1E/l7GtK
+3m+0ZuVPD85ZHFheo5WhRK0L/AKQ5tUWIM0OQeedX4QxVj37Cs+NMevjsAI
+sPKS116e2mueD+QfCuF3SNvzxA+W7+Ii5kYYLt38yPcZJJySewfzO1XXwvm
hwRwZQaSVIgavlNCRhnwDuBJnQRuWvvje0swYyoU3jihX3Rr080iDqtqdQP4
9H598j0cneMCck52yg5873odV1LOyELkyWEJhi6IRCenwkamvtzU23lLfquW
jjB5vLQQCVgo+kr803GW70iETl5dn5UKbMW8IRbk6jsv0+pZvJznruZwlemJ
OLfORWiEZ2MhnY1YtH+NDLKbgxu+jnepnJMlu6hMcUES7WZRHH63Afo2nu9x
H9hJ9eXUnUzcSePAIkpSkPrtmyQY3Bt8p5um+PAIJ53IFgEL93y797Qmg5fC
ooEv53HGzkzMpdac9taHVFEf0BktO6dY3/vsdQ1vAdL5lCX73aCajjpjJMgL
CskiaEf6x/DBKiBbSw+f6ji0eo6pawOZwYMjGYvCw9ecaJiSPi19atC0CCaK
03C3WH4NfEL2uOHpDk2nsc8UKCWHgLU/Wxsux+B6yP3xuVzmHVJZCdNXL8+a
j4+metGO0pS6Di49JdBMWbHBeB8+IRRyVQZhhuroSOgTZxcZ8bP2K5ubQHT5
CtT5j98+/Iwett1t3Wq9ZJWNMgB2DKQpYsWPmWepGDjVJoCigu9h54JExfxd
Pwz4D4Jnf4B4W3mbnG94Tofsil1JYnTFM3MurE38Vj7E/MqhHu67Exr0r5l4
xFRo/AK/E0IaZt2jILgWN1Zfbw0vvs62LMZgrPhh3wsAIguwG+5ScDx80pWE
f+Zu5OYuqrT0ZBn/RiP3smMUwdMsepqhok5r441sx6dYSwrDpCh9GGDgVuEi
psYb+Ibsr4/mMUwJcglLk8WM2c/i84pZYoMw5ePdjKLAmBxoqEd5CPdmL33h
PdT6s0SeR+oRJ90W8EKpoxqjhsvtDJFdKe9dOELLeStKGMm0z1eSBagorSfQ
b+NUurG9mBEZaXR+FwtifmxJ4ivplJYsmBmQatmhCWuCm9dnP8f/EvrgrGIM
05epekKkVEpkByTAHWqNhvO+TIgJg16YwOU9yDYbGyX9j8Z5TbLnkv6/R6Og
earZPCZVLJYJ9qkAJkTVHb+dTNVGXyhtdboADgaHo6oGw6aXSfFHLGEqEJiA
WOaegNLS4Bp8ZruJ8j9LGWdtpYNGAdE3tEKx9Sf3s4NC1Yeart8/HVqUXgJg
MR0KuErqZ22wEf10tNEcfjdkKcaWigQNF6WHIJG3lrwWieBjW6hs1HFZcQt7
bA+keJFknzK7xp3G+VkLBqWZXQLZc6pBZ/QBCGJ0mWEffT6qSHnc/+VPIus3
fOn3ipEkFzamWTeZ+vrikCslVYych7BeHxtGg/1yK/tjr+SqeCgBU16x4XZC
mOxJxGVpiqGIuQaLR9B+wmxsvTkwQLVdCas1JEN85dFIb39KWPC/RIq2Oufk
j2roDvb89gOaNviQTu3vkfOWKEo24O1uD3+BAESLvezqz5V25RzV3vTYG46x
B1RcB3eItERIt06dJDkDPxI28iXL+IZYOTYpeyjpYJ6hI86C20WALPnTgr1+
PdyuWCiHWRuIOAwFJ+GZAUZu/HH2fjkIDEmaZ19J+1xp2wseo6nCWJ4qg7qu
xbvWVFatuYP0wwk+QocS7iiHcrsbMWAA0+B/NxuUqnTG9CSc5S0ZQf3kR27I
NspvRzSt8FeeD2ChomjsoCXBxCfuvTxIzAen5m9rD75Hit08s3Op1R0XE9nk
4EIeM6AA92UQvhgz6V0qaZ4Kw3PE7yJC6hJh2W/+J6KS7PM8VjpzsPCMg9GW
zPzvznKVGTwGILLIbHVexCF9J5pkJAWCWddRnv3pORsR5Iv8eltyYD011dKV
U75rYa3nuOVHtCowxedZAY3LkskHuh4kh1BuC86nPLak3DeWD2YhedadEFxf
2KS1OeqOC4NOChFukW0HTcFoGLfw+EPSg9CgmrGU4Zd24YqB2uq2rbNtfPnc
/Si6oDtSiuhsS5Cz0wsxrpQ1BIhx1VhD/U3/FfoqsOhYBWw55OeQijL0K9h4
rXbbhAKHLny/2/Hd/AwLQ1j+8Y3WRZajAdd1zDCklO5ntBdbQ3D2ebJrzZ0R
xrypLfJM4hGJkUt/TV53sfkrpgY7YS9sEkXuyotK2z6bP/4EBug6P/nCiFsB
sm8LhpFu2PJSKG8bgunxSthseTnEzq4SfNq2KWLuMdwDnK8FnSnURZ8OmgE4
BNV+yLScim+2Ov8OhA7kHygXlppt9E4FozmSY9f0iEfWdcqssOymhP6rCiAG
DnwG06ztKZtOBvKq4n4hJRHaVWYTml9KPcM84+EMwBTYS0V8OIwebaBtvS1k
f00Lx6yIKyYj/dmzlxzncFJlijQJt5Vh+6TbjGoMtYBijl2QC5vMUfdteokS
nIrwPKdWxH9qKhZN6FXchqDVUf4cLmIyGvx6SQT2fvSTqF+Bbjp3uWUwLYjC
WatL1P0DKttdC6LQIQ4NtoIRxxJPqwHKn4YcGWYOUSkWCHM42t4iZAzR7mwd
jMJ0D1r+eymHfNOgmTe/xxcEei7Wmzwy3YRPp7MDKENTvTUSvT/pAZyks0bO
faSzXM+9h1V5EvRvH5DM6lxTaS8AYbXSImE7u/neWv3+9aQLOUEbXyMRAVTd
9nw59Gc+EQUE47wfNt7lv4rQejMAsG3dR1qRtAu4HlZOiFHNl1krQymvHDsL
9OQvftTauDHwAK6HCyyqi6taf2kynOrgekpyLxxHu+VoG/IPYt4xD9hKPPhV
wct1cu1vLZe9LUUbAV98Cn+CFuSXR6e3NF3cXJ+nkJ8FbGVceoPzOC7XDYEE
mEltPDb3aPOv8+L0GHNBSOEltD0FOqshDTuKjEzveN19CxtQtI0+TvQAUjVh
vD/4/Ycbd3lzu6bYVvpzD8dxshkgnqHsMc9KWZ2wCzBC6LO+3bfwHKdletUF
c+qaHsXrBkAu1Gi0OGDezYOyEnIE3+mJ3VQZtKsU+mx7Xq94Wf47O85OD5YM
+YQ0jxXcyH1sTcrZDZR1YYQv9/f+w3raMpFECwEEzXRM1fij7e8AFKVsGDqQ
n40wpymfkxZfgOsk0j2RzrGYHDbMTGnkUFPXgKRVde1nqGjwadeLvVAVTQS7
g+0DN4euXBt8XCw7l6di8tfFf+Y2e5gpODMsVz2YQtQHfzAEog83Vxp+SQMN
Mrep+oMJVrjyORAO9bxKpYiRZfCKqBbNuP15pv5tT3PFxkh3GTGnR8BBVtwa
KgYgZcyJuToNO4AmZmzLW1Dvo4wV3uQ3SZBytQv73cqREK699QGR87X+D1OE
P5egrrjII+6WHQB03yXhdtifwG8GAaoa2B0onc/YnRggM9spiBWuAdMLCuIN
AGw4FmnhtjckhqneS0GYfZvonlaFHHkRAXr3Hrn06cDrguFpq3flYY/PYtJ2
PmI0A0x05PvDvHogKsppLMYlYU3B/D14QFEtFVIZklpibpB2/oDpcP1NsG43
S29klmEIWlaNGNyyqGjL7tbOoPWWiHGxDrpQ4o0c0rUfvIthCtFEfclFJ6qL
geHkAhgG+9avVwyuU4xwyHO+hKTJXYHfckHa0h5lGOI2Q+J6g6rgXvTt5C6q
+ZPDhfxxbdK02s0Cczl84tL1Wu0Odq37hYqAriavFyopMbrWVGM+i3Gve4Pa
OP9MalkXQxOOgqMWHkELSXVtbMuhXQCMNL3N3LPoA25hLAoGVBPd3FAwTmpF
sIheYf7X8Et92Kp1QqOx5LzkfmSK9mjS3ccl1t56kqh0dU2FwmCP2XL8ikVc
eFy88KJ/umYBlOsajHpMl2tRAmdWNaYnKsJZaOIMLRfC1LEmRWG67BWSJ/l0
aVfLuN99by5lny7pIeoSm23yVfKwknVgPZMfRk49F3whaCjXXuPcE1cOqqxI
l2V0moq3EZ87PBOiLUkcg8gFb1BwmomtMaTxqIpMZu7NfgXx7MAZMDKCusSP
FBH/RWZ5ZkTbvzi2Skm8LHfHXLTTXHx2aHXcWi7NDJcMseYw079Dk/bHhnnt
U7mOASHMb3EWlc4iweDBsEWzEiqTgyJnaLlDdnfpVm0/eFwX6UbXYr0OpsE0
E/BjiDFSXrnyUt/KltABtiIhqtPB1WPBVqHTNS+QjsRfZ2JJFKs6BS05M3c7
JE9p0N5e3AQlIqbZjzyBFZQWCAQw9abj6AKt8rc4+n0NdyLpY49MyaoKUFQh
r0pu4Ij5V8Ca7MeXWhBuxhz9NTdOaf1ysX4w+a91ADj0foXEosCkKZCMoaMM
Ai7ed/COO7RfuY5KJJygDktpkMX54Y9kZpKSX6QUOBuTFWE2wNG8u9MJsWAi
pIZ3J2DbKwgTWQCS7p2T8IrfnLgD/9p5vPgYM8lRg7BlwoVhqLljAB64BQ7D
ol9p41hpjDFhACMA3mgh7g9I39ytIEsMg4ekFpqjHAFE2SbwKI/qQBxAod09
B6Psp+qYozUtxA2vsdej5itw8J02ILho9tvbaOuNB3AjO4cWJ5wv4b0Sb6n+
CRjNnp+7dB2jYiCY5GWOVFK7R4wL1K5u2ijLL/zGdr7+spw5uEGwgTsRYwtu
aAthe9MgOIdcCsrZiGti2+54zpMmLYa3hbppIf9OkGjpCPfYkirH7pqvGbJd
bEUXGsfaArYcrJUkfas1ZfIVceWc1E5DhXH1P7bMId9mj0c9tT231KW69f8Z
9O7nU8N7ETWIhyNaTzyr/6JcJXM+6CGhharewli+b/Ob6kpsLiAEhVr9rpIe
ieahfYpFEPk3rZSk6UKMhlVFiFPdYIJvPgystp+ar2OdpbtPPyOi1zMDJSMz
LG8qGY/CkcwYGXxpKyyrE2n83LKiRCM5ifmxFCikpIN3ycDQcG6nhY+exXu1
wchtU1dRLSmF8QahcnLexWYpByQXN2rRgTEqKWGyIszRxKYcrwvZb6/6KMc2
Q6ETqR4ZAporS2f5iamd1oNPcGdhcqakDtevP09jD76IS/WDjSC9ME0q7bDP
SRAm9yRx6Bma1qitqx0XmY2dG7Ip64Sqg9+6uPcoM7YVOjd5zuFxlUw2M1ZW
OHDjLAdzyGlSl2aPHciA/bOijgsMrAXrswe1BAEhhR8iYbGfQZft1Z6nzvkq
C1CyXL2L/xUENUYFVv78YGA1PqyTjVBsmEDAV9PtQogfdOk9JP4IokseewvY
bOnyRjgbV347ccsagGszDpZLLQKLSy3Y+cz2Ivknw+HgSLZt75aTdEMKpzpP
OL2PWOQFvw+bOM2g+AiDeR2VmDYce2j/U1PZWnOITEjFqepMRlQTy4KJY7iI
8xpbWlI3TAGDV7sN1f2YObLjfOL1c2zavm+ll3hbyWBXnpo4l0BSO6fPdRc3
OiHbVje1z6srKuMQ5vI1Yi0n/ccFx9AcsQl2ITmcNtS4/66wdl+IM5khitri
WTVISeMP64pFd5396AUu3LT/4mOZp8ckGp5XUBTA4Ku3lHI6TMhyj4TBGZMQ
bbpt1LgpvOD6GQKQNgFsIF5zoeuRrQBrXRq7NjgPJm8PLq2QhpNqcQGEq4ko
4hI9u3DufGqw+2GPdHaEVzVYFLwaRSyPQMB7eQwcqr6dgKCSuLYyyEIjFTWb
dIlzbCYLFydjA9c+tOqSbFFs+g6Yek/3jnUT2svdv6fhxAco7fTTaouupHnq
00aHz2MCL107brRmT6NU5FlWrOK1rh9Mszu/EaPVly8DlHXgjy05Ar+Rv/MP
yrDrTTaTJRxkGxUpj/QLn2g60g2CT7UeTeKZj4kkbNhekSuRS1wyUSM6aPgY
rAu77ZymYbEDEW+aUbKEYYinkCLg0a5WRhQVa1ORXpINPx9YrOtG8tjZpqxw
rvT1GL9bOW6Nl6q49Rnd1cb+9bSdbzfdRcwd/dZoYoUUrZwumn3oZwgkTJaG
7AUw4MxW/i4lF9z4Si1fDaogtwMZ3k5QPHjg6gCBe7qq9O6Q99fMBU5FI6nB
czaNV4MPvdn41hiSzgUBxxeLPPnDaHUhAt0hTkteYpyGUGpIBkj9/I+iR5CW
kFPAmPqmbRJPme8DZcGrW/UzRp9pA+VCRwoqubqkQbUNTGBkj5Uk0dS2I8jH
50DTdpf79+pJB0ITMcivMwU99WLx3qfy/u2S85sTSHvhT9j0ZrYIO5/JCVD3
v+YXOpMnocELgb924umTn50/AyXCnmcdj8roiIaklN0SUa16i3Em+GQp3Iqw
yWaQD9usN8KSdBD9097hJxcw3Z6b8bWdzemTmSDx4AlC8HU9/djq7B4z4aro
eM+OrtfiteMVPYY3UL5pKxrZssVetIyMDWCOMDHai6ndx9M4fvRAXYHmA6xL
iLlECaC9Bq0w7IFm0TuAC7XWLETfTmiMaTO2NN1q2AFCtOQCsDFM+rxTJHgA
ADXqSzzyHDmbyIVA6u12A9u4g+ZJpikWqk5y6YOLFE4NCmyAYOvevnHvkN5T
8jpNP+QJ0Tc+EbcyGjcMAl/+9kyNj2x1xSbVWc7W5cqUrRY7G6D1G+KSRqut
1qCXSqoVBk0W/X082TY3tQsJBo72ZsWVWq0oAea6hPx01kVqpH1nIFohfoS/
CywL3+r+no89ImrJSKEnIC13vDW6wZYvuhslAEDvwbmn8eKrWSre3Mz5ENxQ
Oc6ENuSdFmmr37wzIO0yVw2fIAUYTN38QpqE4IqkW1altIL5gdmqDH9l50rR
TH8r5HwdHjOpq/Cm/8Z+Szsa0ZEcgp3hv5y+dh8dbNNuGotnL7OoXUat1wvf
WoHVLSLkb0G5KogoBl06xs2Se+/zUXGwvTJm7ViYwfSsqN9WbqebmiO+VEte
FJeI1iFE+X6IhIk8BdlZVYt7BSQceAUlvWSyaSkZoQy1yINzMeJe8k9guE/D
1bcPZO3fEruVNTgmw0dt4jR/WolBcgqQ4dO/uvbwXuMXdHmrGSnxi1Ldx0lY
GHwcNXiqd9IqUnQZqQzHj0FmEpyumAT9TMMzJGCGyhnO28PjMv/kS9u1FCxP
Jq0+Qv7X/HtXdAjRQ3gEMBEcs6bZTOMQvf6okkz+XiqmyQZ0onBQa0eF74eE
r/Hq+QMY0XX/xTgsuHsPdLohXBclKBSngOMRi8GkSvkVyV6jTmN4NIqzNgJd
jJjN8uMOcyiYcevLmbeeQ5yY+NbGykDVoGepTIfFzMOE/Oay64JO9Kr4wuaf
RR/vrlXpdk8HiWoQ3jCIr8sdO81l6UW11knNSnEtqM56aMVdFXdHkv4AeiaO
GL6187Ec8rtjXaGBTcDxDUksHFiPA1/FQfpstilR9tAzi2mT4Cnx/0GewceW
E5lfFgQ3sVryZMUpehkW1Xbo6WDAGI5YDCcIfpHzvqD/lo0sHL2S7yItQjYY
WeWjGDt6J0LeiDKLKYuWhPzicDHxKeCzKYIS8o7LLu6izhBvXRqoyazU6gUE
9/AVU/FysRDsJc+HWonzC/tZq33RMSRqrRIu3CdjRmewWdMTOJWELKXYQ0+n
YRMwlDDWVdRbA62SqOeyHMzoV+SQ9VsctU4cC8Zu0rA4kU4nZAz7s/p8lmeq
KEWMOZXl0yQh/wxb89aVU1t80wk7TlcGR9LF3NIR9GOX7lS3YUd8d6U5W3WD
bpgCzHEDRkkFlJT76JjqqKj21EPStUkXm1l9fl3ioWMIa5AB4UVm9fSa8csv
P4Ybsljdza5e5WLf1DNk538S0MDLzmOVcxRgOsh7GIIF5nAO4cAQxlq63+1C
SEVVUF+vhaJWhznPG8Zj1d3bztBBUFkWRB+I6BJ9EBYBSZNF/Njv4fxgq8rC
ggZBnKFe8WVc2Myiby25qQKGaSCOUFuUFOghVv6JKRvdHtMrdD9NEdHfCKlA
aw1a5+lkN0q2aw2ORn1SR8c94YKuqPJZlTxJQHZE3RrsWN1Rfgl+WFZiZdnC
QNGuFgfMmFaB44DKtLmXrSDjBnD4SA+AKO9R9k2SEcd/9cbICTKOQJqTrB+z
cW8R/XKDz3hqWGC8jKsAl4zs1aRXm2IUEku4Y/bSTlTiei5yQnHdyDaAqlZ7
KIfdZu6VETgAxW95t7z95L4+MZi0xohRkaQUKM9ECDX7wmAS1gtUIGIg2tA9
/s9DEOj5REKCaMn8hrlnU5jaCODraBSvovrBfkPIRrX+rm8/GeqAzUpGHWnj
lc3S3UcLndFYRKMm/xt9iYIj3WSFekFWKuK6ou7uXsODs/Nrzls4FvN11a2M
uUwXhp+GcKDFurgRQZE9mx5wc6RVdSdJMmn3kd+BW08caXSxxUmwEFboE4az
329ixqVIoh9n74mtvOlapgWiMShBBFkZEqRyC8Bh6AQRglBnGSSYJQ+T4H3S
Ok4Vf9BaMtVXUDO6/XsCQZE5BPBlzXuYvA0CFemP/671A8nJdarVwM2KMsR8
f7nwxzjGUH5FXMVQnpD5Xli0Bp4LonmLUhYzB9/pZc74LKvuL/+xzcJtZzDs
sd8TD2OUxhkLSk3o19AoUypdr1ZF5vbkROwH8XwI7qQoC8jQqf/svBcUBvqG
fWxH9NzbzXwedre/qZl/PQsvr4PVoF3PCRDirbDOzn6xRT9hNpK0H0aKWx6I
FyauzcKlKtfD7ha/zsNOk6ZxcLGYGBQTnuDARpjZ7awPbLvPftNQKc0GMAoV
JYjXnbPamkt3Hc8IFihhrH761B8+zNzLjqplpmti1fCm/Zlqr4VvRRFubA5R
G90IAeEnFFecqHBR9H3xoReztFRD0JpL51j34Z+qJF1Szes9dbX+67Jm9S14
M411idcZ0nMV/9CLzRlvV6+lTNwUDoML6bPdVspkHHens5zC4iSvi7Z/n0hy
EgJfbn3Bnop1N7JiZhKdtxW7roOLGnv30yCuzeKhH62de+gdyxC41oe6OVQo
Xl2jCZwxLIjqjb6NRlJsOjJvc+7Ky40tOexFgo52ob3LZlEjQ/0TFYx0oWpu
BQSC4afFS1es6tI70KkqbBajjQMnupLeMNoiNikFaJV4j6nubVk8my+0mAwL
GSnkm/sELgcBAVO8GOJ/MzATVK/oNaQJZYJh1/7iFZv/ECuZDi0L+YgGReaw
7085TTXZtzAA7XJXBL7pLa3ci43TwLo/kizJexclf728DCTQxYzMUt48rbw1
k2OSZC9f2b2eTUFP6kepzPUJfOCgl9MaqEIbZ534MTv3uIgm83hNLPZR9Eqy
YKIYnDY794sq9ugEGV9V4CdRLFO6lVi1NXff0U3FHWxL8F0Mic4uQzbG0fQv
2B2OkUZSdOQHA4qLVSyEkSH33torGZ0aUb+3xh14F5rHjEqHUQaBl1+Ot5Tx
FqghUqfiw1zrlKtSxKZBnX2vq8e2Xe8PMJ+N8n2mSyECkhLG08oX01V4Es3k
kL2jUvOFkSbvUBMnZ2Z6XPkqaI3vW4aXLEpg3MuJUMT/y7lPteUIUSwTckD9
EKw/i3/t5/f1C3Cm+j0qRxrxLq0Mw3p0NEtGIagtzR8drJpsaSSv19pCBhXG
4jdOvOGT3tjXmve3nGzqXiE572ZDObAyBETcWmMZ03yx6HaE4K2zEY6KRtF4
CKjd92ffwfS7UinfrT9rY/pmBriFpHVwriC7aft36+x0AQEtS+agmSsBd6JV
8AWv5gTOf7rXivB3Z2LZHlpnoadZIfhUKCbN2YyarFodNX3GjCUulyF+3u+5
U0TfxNj0qa9NI/3FrBFBKfowkOO7WEEmnnrKpKwk0PMZhORZ8X8zStwapAjH
ZsPzB9zdki2rN09zitJ6yytFAPacXiR8Gi6Eg/WDKPHexXu65ybtxcaW8YVG
NIxsIcrTsRxkjLlzRQFh0NDS5bRtiyOUFppey80cxXtithBIFiHtmVRNuUo8
y24ZdlkHEszDK8RQq6djBIYsg/qZelJv5r2xJW+vase2U2NLgDg2Iwll6xFd
ZA6cmrdHAgRNDT543dMsPAYcr6rcwhZGX1eZw+AUHwEnhMyckb4aipXuvHOD
wYgNjfYxD5zAzqi+GR0quzCb9rQPQtfZTPF/1f2NhELTJey3xX/2ZBIaXtun
6I73DpKmG3kqzkc1HFXDWEowqdT0e4XVuFcbVVeqY+05SeGnYbVlCmpYeUfC
mZFgJ7FehfmIgX6+YrdwC/ot/Ud1aEakhi0yzdKjZraJ3L5LzYUmFU14KqOD
9EU9eSMBjztVuJ+bA7FCQNK1OtthI2VQDhjpYMlVRqU4VN4dbF/Bw4bUrMfl
INlSy6ogPxesjTUJGEhjP3eFE/a7eVo6cIQmBo11mxZYYnhu5y5yZchBZLN4
5i37J9h4JfeJQHxy1PzRutkEdvzcee65Z82hRNqTHEdvUEw5FxLgfxqIlxYa
KHRXMXBWJtjzy98Og0fI6q1HobPk15HZQa8P1wyUz7qfesjE59Ar48hhwv0K
V2iHvOX9qdhhVLkhMTB4ngKuLre4IUPsRYtmgw4itofKbu9uhTF7TfdPZMRc
ntoaZXe6HoyO26FA0DBk954j3t+HJjhijhx0NgngcBy7hZby7JraeZ8+HDkd
DFc8RXvdQOdEIEy7sWF8DGU1w+WksGJ7ECsP9deWkECeW/FZvBqlZ9GHev9y
Y0uVvxmTjnVS9G14cgu3Qepjbg5zZrtT4cBUwcD3WTLuX2HVCmqA3PmWnCJF
eYhS/vIn92vAutPt1fzWfNZkrrtqgUrBdVNMcO/M7ehKeWG2qkMmiTxnddHy
RINiVtFoaY8pH3aUWrGmb7QXdpT/6e+PZHdm6sk+KBHvUIBOOMiwewgtHBtS
j1Lp+MSRUZ5ulHUrp4IECLc+mE3ddUXTR429DfVJv3BpWrs+XLphJ8DhHRzr
QjeZLKcjrPQr4FYeyWXXxp1a+i4xCcFuwihblijvtI5SX/2as6claP8jK3rz
MQGsW+ls39QXwXxGUwx1gviYqbq4leUDFtcWBEbTm/i6+a7CyuBeC9KSk24l
BkxHKhl9TF9gTZr/pqmf7oBVGCuqE+tclk60+CX1IbmdxZN0wZ0gIIn9kOEH
nOrBEZDVn+HynJSbpYcWhcYcP9H2nUeLOxCqPZKSOyYunTkhXY/OIoMnYrmC
Qa/zaEtu773KKif2iwVT8TdreuwneiS5gNIzCs4WOoVSdzOTpCmEZP4Zt3hb
eMCh4nCZeLeX7H7qfqZqopBILiVBy9jJoJMWqxwKjDOPkXuZbBx03RtgcA4a
T5qyc/yz8RiNF8/lI+EHtozYAaYfYsJ8nuUCI3Sl6KI9f3bFbedJdin+OJCV
bF+XxK2ChCsUQG7mRKA4WAe4vng6fqFM3nhdA0+Avqpj8uChiPRgN+0h8PeE
wYoE/vjgDlXiqcOZ1tHxEd8ppnAQyOgb06yru6NWf1tt1wxLuRlvelQ3qcqY
rxk7YdzIjF6G7DEF2pKPb3m+CMpXapoMMnBp2et2/G59I8acE6jffi3RMOOk
8HFtCQ9J+sYFMTLxmLHbKdId409jBrVXAMv+Ss+jdCnNT2Zqf3p+XB969n2z
gVWNmf0yGHMeefkK26aC6UEFcCWiebTv2NCeh0YKvTkZ5dW5+k9RAdOvr7p9
tb++08hLocu2KhSIbQKS8cChrS87XFhdEHuzq6HP5/ZCwtRSaP0rSKdmz/oe
+A5O9VYSdbjP46sXkSrb4Ef9XMJC93+GYRVIvswdv8MPqnL/wFmBkfTmq/nD
K/AQU+rVQZxolz4jS2k1wBJMRzVdB9NMG1xlstnhF84e7yQgnYOr64FiavBi
GcV7kzbNUqfeJrPLLgL6D/nIlxdjH1bvARWJI6lX6RhuOwxm+a09mQ5aAdDY
yuS36E4vxL/CgqxWWOr0s+Rr3pxS7QQxE/CRcj1r41CAyf0zw0dmW7TL3nTR
u7j4X5+sp1EaeZoghHQS93aLn73iFMeQIRx92H6C/AGim6p7NZ8VS9q+Kp97
Q4uYQAxeRrBKuq0UH/vsr8SzJsKNGZ13cHbyOnf89M+/84MOx3iaV5yAkUME
Cwwfi59gVIGBNYCeUF7DyiiRgmrZfHngsdTukJS2PPOp/B1JX1QV5RXRNMjG
qW9G7e9xKAsAN5L61BJZvlhm+ywyll9LI4Ir/bzGIfTdWIbPC1unPrtqQVqc
TXC1ERYeYk+Mtn+zR9JFS+TI2MJ4ihcksdT4UoPu2IjsOKmKbljvi4KsaCOz
fkexhz9g3txpNo7qSiStOCkckQPegGNDGUl2oIj8Gwnblc+50Q2PYE9Sq+07
xoM/FDO8mVhMb01yVbvxMHCdgf6uvuNiPdshfpw/U2XA2UCA4+2l3XL28gfb
yGovqXU3rH4bB4TNJN1rQUfOwjoN5zdlihS/5k3GKgDOOvBoSUwH0QnGhcpm
PDb6oGmf1gWjP26U5nDhBgwVfIz1WmLgt0AhzdbozIB4zWUknQq2nzs8h6Ri
+fNOOXfBARdaVfO/2vdGkWRxVR+eJFLyaxzgENv+Bl+XVZEuc5mYoYZ7Wq/H
anfkERWtIUJjYcJffiCWFVTheXdLJSMM9C5H6arcLC54qycJB9Hs+qgFkuD0
p7J8SzczXCLVs5svH9yzLBmVokgI6uTijsPwzNdnVfSBv32xJ3phxYaeQjXH
0RRT1DIGNDnR5b1G0AgGl5qfG+NRr58iVA3jm1tJLkBP75TwGlipAWtIRrZ9
jfhY/GApEsdLPWhSeivUCcXRXjhjQrO6wCc3KgYAVXuQ2LT4Dx8L5EsLXh6R
O/WNPA+u14Wue23RN1wmwGL6oMOZkMEhkuLaZWCfFDBETZ2l0MwkS/Sr2uOB
NMm6TGjOenwZOVfmptFK57zoxrYnhaqEilfw1yfCjiRnWcuGpUZOgPGNBRmA
W5STxMEYaKRTqDNOQ9Elgw/XiSF1Lc6kC5965ULlE8v3f4a4CgERodleuh8G
RTGh8U8yC5puveHTe+UuCA6fLYc2FQygQNu/fKcrC/FsNM4XK3s0hHAyy8IV
lWCgFagoadP15dQ0NQqGZzMNGMwMHUvFVUoZeyb/4hyPV1nVvi5dG1/Ef47B
WRljXAP3sX5zhzIf8rWPggYntj8hEkW0+cDYuaY+AeQF1o2WsUoX3qeaBXsE
S4DzWzv4Hw04naEU1RytsjosVodNDDeLcOj7QfNyuj6uWpWtwxtuua5Pvl4Z
XW50iHyv3Dg3gU4ZkB1rgSMTCFupwHq2UnxfeTihy5Y0OZYF+I96eKQp50kh
zwweYvBaFpNd2320HnLLkwqgeZEYVr52+e4zec/rEVcBMkEqfbhyQOFzvpOJ
VvvL4MMR3byIXUT3PuTx7/XTbL8sHy7sKRaeU3wWBV44m3moslMq5SGlQO8q
cHpq1KJStM1CvnONF9H+sDBuTK3ijoXerJL9HfAegJaVHB64ATmu1HaWgl0X
ZacRcBMi6IdPH/R0FCJ9wUxrsvMBC+zKzMcgUvyeFV3xYvzcRqM8XR92+26V
KbkQMy1+Gi7xRpq8hs+XCCIm7MNrgIjknMgg+evkot7lQDB3Ca9AsctHCCiZ
R65sQQpkXzHBgCZQFlepyOtgDfxV2vwUwJAftE4swgy0SbLgdDfzIFxqj2P1
+AUT81Chl4MPfJE4UBf9Toy5EQcpg+KYnyDd+qwWLUFL0B05giAcFsRU3yZP
gRrolFEOhushz8QUcg+6oJXBpcu8qGDCzFEwt3YGItOhIMfm0kmm2mmOoUXn
SToXZOjyvK+F/bMhFAikU0UIELnXIBvvU4Bx+eI6pdN+E4A00oHcHNQsiX83
D8g5np5SmED2FQnWsPRM4x20m9uNXLBJ8DF8qMGKHHTdYo9jtlyg/JK4Qv/N
vJ8ti+lNUU7HuLrdsm7I3snb6iKvUAu3BG2GYBzMXb3GHcdIzvZBxyTgAswO
i8c9xvj1JTPGkY4CNT4s0m8MHvGbv/Q784w4PExZjcA12KTL1B9aiiDTUn5r
QJtr9XPJmq8jSVSPPMz149N/jeD2z0Dm7/00J27H8cXIXVxd/KHzeKMnuOzf
eOUjimrrFykPSGcKwBqe/Nd/6JgyLSG5P+yILNwfHVFFCQ9k1NERtHwH93v6
IWohpsVGgcXskkmdhV6AtrzTsVQw9kPTbvncawiwt2eEFS+vxZ8PIakbS4KY
4JLYwM3JUjwIjkimYkzOY/cmIxeQWDRvL0MBckET0A8VIkAu4+fLurdgBPFl
0FhB0JSxsqNm36RgxdJKsv3V2UMErfzFlMG/7VcucrybbOoLPRNXFznRuKBD
sCwk6znQrTk47UpwyNuq4PogAIWaJWR7xcgsqIq1hzr7xLPiP3CpR8ogoblX
zvxwNw9JKd7U3qDuvgaQ18KJYq7nXJ0p1KfHvxe3lzSKz/3aJazoHUhpZBx8
RrRVADFI3PmMftQYunmyqs2kezHbTtK4NNI5oj5RAqePVRnWPrDrcZnif5Ix
dTLvh1L+C7FwYJvO9yg3LEg4Qw8jU9lB8Juk8Pp0BZ4CY4i7VtVHkjyH+reX
vRVgOB+SnyR0aN+KurR18sLKIJIQO3dUQ4oihZaeVej5MWQrEHxFQUlBhS6l
q5EExLaH4AsMDClsrT7NjueCs3ZZ3xh4oy2A1yodUBy4RUPhkCxSe8QmDp1N
gfUNtIPtfF+hkRQsJbKrzzNNVL490hWw+6hgm6feMryHNWOB2EAjDXt4dR7Z
lDGA82APEXI9Cyj3vBvgvzjHzjSkLOJa8bRVECEaKhUR8BTOY/rPko0oE6HQ
UkJePaUQBcOZQ7ODQpaiOxx8TYHLeBDoTHjrnArgJ8bw/N/L9VmdmKFgIgeI
qjskDV+NbbQoHZW/r6E5a3YKIiLgC0YeSOeuhVtsp5Zlz5k=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpegUSe+4Yapibyri7SNlpR2Wx0NjY9/wofmdRx/UkuqBJJakoJjoQLp/OSnR0wmxySc3CeOxGvC+8N9yqZMVrV50G9uzXYaAI8ENv3E1yvev0JjNGmwDisbI5utI4HcDQopESv+3aZrpmbJGo+7yf6qjBAjUdAigC6X51mdv5Hp0E2bmzLrIHAAPTDzejDLbMh1+FX5+0DYLOaLNJVVkH6VKH8AQVzaLKsGBKxgT1G7nUBdFCNFd7XeTCCQ68Aa8GBVi891xPmbZMAm3oDV/jROrjv30EZmKswr3pZf5nGf9VP3xi4B6dl5T6Cz09oSONcTiBMLUSpwDsFan3NDJlaRYwVEY1/R7XYgtOnjlVm62uLfiRr5exb0goAkUb2+55BMdbx3KuaFN91R3fpyqbGBZcHkUxyWd61A6X7AXzzN0RZ0RLolwtj6AdeAzq9bZa5Jc2PXnO922jE1kDW/yfgsKHIDMTI3Zm/4vrc1+9jFKjzuP19F0qnpCBYjUd00HTDhbylnt3y8D3fO+Ow6YnWyH+K0CTUeTiqLNFL+QbuUk3p5w75D8C8Efl/UuZWaYwQUzWO44sD2ivYccF8A9vn/tav8y2fBC0p44POexDpOiiAC973HYdzoemxN6Ee5zZzMjl52eKCro7bJO2CGtto7Ja2lCWs3Yzdh+b5qhJQiRaakxeGpL5L6urmSpeorURuGrDHWpENYcGFFz7urGPeMs6LqIoj9DmZdDfeIGWftzL5s/qY6Wzq4mC6wWi7YWdAIJb1/LRWJtoGkN2lzYQJ0g"
`endif