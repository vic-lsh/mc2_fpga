// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nfbq1umb944EpAogsCurC0FuKMkWHjJ25zF07j6huFG1Zt79xv1enI6ZsWaN
MBKuUXnytOe7Pj+/vTgoxN1J4MBV1LghmBtDUclfXgP2zxRU0Z2YCCH6srTL
7YZW5Y1E36a7pweJu+QTUo3lOVInhuI7Uv9m4s3M2KfGUlfJreG5+/ch0VGn
UtmX7+fqJFWhsVAjAyUY3N5ktdEhubYqgZo67W4RZFCuzem07GDGwEtZ5Y+g
I0pJdvQ1ZuaZ2mLfGGpkS78Hv8Y42ekQJaelwrfA6+cZE1fnyGH1Hh/Ogs4l
coOreTX7VKAJxY4VU/ybuvxqAnF3s80C6tqfPrUu/Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Szn5v+QE981Nm0eecHDvdmrwO+LYYmdcE2iMV9l1Koj0byrci56J/BnTnqTR
OqGKGkDfKCWk++AXtaPY13Y48CeGTAMINHAjH3uylKS/68JAVsOBslpDHeAy
mpjmIoUq335Pz6u6z0cu/XYnWqPWCR+WotIHsVWIpddIOMElHzbucLOzxiJz
6xBv+P9E5lCCUUCpcBAj018oi66cpxQIV4zMA6ShIHw37a6+ii11JG148T9M
Sbny/7nlnI9+G6pWpoqXiZaVi4+4O/JLEqA4n8TcnOapCLw2R2+4X9BL3kcP
rQRa+Tx7t3jXF5E5UE22thmccRw0l3HsyClYXkNJzw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HeasqjEwVhWipbyqAxnDXCWyBjeOBA9dsB5V+QMQqtirp3JlNhQlQ01/7b0r
B8s6iQF0Kj3e10v3x8WQtXPHHoQrJBBHKxYszH1Q9Q71vcr1C+Aj/yuImQxB
djiZJ8RZyTaZuhA1tbfyP9cliUaMlIDKye+4usqm78I6iRTu6HFu8F0e6J3j
016VtgcUm3cYhWVS4bm8z3jFEFJE5bHlUAj79z8TZHhrYEqMvadRW2ZtibDp
V2RFSWVIcvjqWz1r+qqSCCIhSUWlblJ420KMRA0WHRBVX/nzuEWM3K8rtCHb
AVky5pb9BvYRO9q+ogxsxVhpTmmDtzS1P/8vReEIcQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gdcbDte7eR8jWSTD0v+mPQaX+trk9ex+JXRah60aMFznKePk/OklZxCyLila
X+jNy89M8DZoiCJroXlgszQAkbyZUXySfWblfaR4LUdG1UzoT5ZJmJneLXwW
9cQp+o4LBcC5Fnjbjjo953HemWxTSRHouo+YOUzRCKp5hw4KQ7jmWLj4tR6d
eyBEEbXHnspk+I4VEo8Y1eYcfcqPxpU/DB6O7b9VLprQy04DrVWTm4pxWw80
aMsvYJw/4+tZTM/oSwD1JlnLizDAs+9b8IHbI4ZIWXDPW4B9mRCIBWBIyAum
4gNeqhfMrzoYedYNEFlJZkO93G2lYCWNEzIsU+CI8g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lqR1EwG1croEEJH+TO2sj+VyCDKpsXlYRXsmpwDHEWO7kt9SDfEvMSYXgFuX
mBZKLqDebuq8UKWfH/5uUqqmefoAAIGkvzIlGTn9oNfBsapZFDGDEkFkvglb
tjniUD8LmTfeoNySuK3XP4+I97WvQKGIBLqoXMOH/4Zdd8QOVVw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Qd+fz+8Ad/CYS6Y6gW0D/PuZ3A+/M77no9GdDRgJV0UXDnHeUydcp/Kf8wZd
rfujQQUk+Dm+NMSkdsbJel5Bh9nsIu7Ox6Eeqo6nkxHrctaeIh4oG4o/dL8s
YB4p9ual3qJDqrltG6OhgMFcje6c/V9zQZuWclTgiJCZ5iGyD6zQyydnz1Qp
YgSCVWYRR4fwcM7l4cK9bR0MrCWITOp5BYYs/rDb34ClS5WEnWyNq5LPALtc
cLRYstRcs/9tDyYDo3xOc5CVy93MxauvdaLsMOBFoa+tiolRcu7tRVvG2ayQ
VQ1ZxmpVCq6RjNfs1UI7pFpkdh1IhEcRJ5MOqZTFuccFMVmiHHHq17Ny7V7i
1QogqqGHarKF35nWDrYNJVcyQhXVpBtfuWBQjxdVOLhhtP5mYUkVFaqdcX9M
HkfnF+JuMoT117Dh3IVNjwybhFSdRZJhVcFzYDPDB/Tv6d6UEdVb7H2fOiDL
3Tq2xmhnwMUt4QOW+wbAnzri8KoT3ulv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lODvzCpps21jUXe56Xm0GwOcOpobI6f4aHQEzW1TpEwUrqJ1fhTzYKF6ATPl
LLPPT5PzjcMSPglrSXSTetMFqWiN++Aki/01GdRLdNkoR4QzwR4L7TVBOwAU
uXofsqhR2oUthp/UyqL8Mioo3SDRb4ns+ST5J5j5tp3OKzo4OzQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XYpVIOczmagz+X8sNcU7QIHbwY64zbpEiUOzEnEgqix03kUHCdbPlHqNfJHc
9OPAmxLTXMiOnPKYY8AL+P+DeXMuWLeg3qkO0Xd2K5WEG87AhihieN+RYYEw
C7wRTxU1ucdT6hxNoZulEWaRk2tcnlHO0mKPt1tPa871MhfSa5E=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1216)
`pragma protect data_block
IjGRmuBhTNHlVsV1PyMF9UrOP6GSOvtUGoPmgK/iqDyKVaETbCI3LEnZcznn
QY5uVtXqNKTppzaOhj2osSiVV6MJVCR7bq5ktYuIzNjok0TeiwgZCTf+4yN/
51SCoS8hfFAVDS9znTcxBsLsIAhzKA1oGwoTGS/FbJ3lkRImBKX6SexeVqcJ
4NhUCeNJ/i+YGo2RyG1JH67Zn+e1bE67hcALi1IuzWcM1/Kd0INslvtLsDiF
5yyInreLJtqJLuk9adJMPnujNaslR/GbPyy87yvM7AF2yNJHilvbB6s/6Wah
+5doWcUgrOauTT8F8MV+3cNETdf7bng3sdGtC+fz3z01TJ3fCMuLH1RPIbLI
t4sqU8L7BkcxAXZiEObXlYdqSkpxjt3ZUPldzDrQDTiAH1IrHkmeNEjxkggs
GHH3w9kZ+MJ/QSDFo7cUei2RlNZGbsUVqgj+Ra5mL+MrubOpHYrwieXVEyTD
UE+hHsQfWkCiO/bpALn1lJ3EdnYXHKCTkLQILx1dP3vpRFqak7pUwaotwsM3
DY+8Mz7Ff7TpXBj/jryFTKK3ZfeCdNv4KLisF5ysNDwRrGYc82G2HvA+cNd7
L4rxZXDNRFLe36pdlHUVUy9tJ5j9F4uusykaXw4wMS/nbw/Mht7HRVIg/HR7
6u4ojndwAGPQblFnBhtqtRcE0knLwf+Zq4MKQ76mAosewh1aHIm6Q0TIIq8r
0NgiVFF8lK04siUJWX4V2nkj+F87fItDo57SeXeDWFj7I3X7iZS6b2zKrmTw
HZTbYO49uQz+qxDIWqxO1kQzipxHpck+dn4mYMqbx05oSUDNFNzx/sQoQuD2
DS/NkdP7KhNu2vMmdDhAPR1DzO5dDk+18vyOgTRCELsG3+Qn+DXSaxEZDttN
XOTYn4oViK8joSK2ibPo88jvQGGU4QtByrgt9i8UlHzXVGnZs89IL2dkwkv9
XVYxg0FK4HpMozsZ4kNnVIC1rSZMB0uGNpSgZ1ylRooboORNp70hpjVdRPy6
y5+nFJwS9HGPwT1Qy7oPHdbdsq7QMs08rvkNlZ7EmAYMD0nOYLlOYwigcGoj
pJ9XfOE9i8qXjN1KukfWfIPjHvMQSp81+P4ZnHyMbbO3OVB1syWO/ac+G7+F
TTDpzERBYReDULywTQA4YJrf0HFchRHhw1uPTFkcloCJ7xcM6Js+BK53+Vey
kPACZChWMP0XhQYyvVM4X6ARkcDW1ynNww1QOH8BR6QeCBPQqZj14Y9c8E1D
+7EYB0F5849L8aEBO/q0kfRHpBEPoKhpk6C2rCdA1oXhzn/fB6JDFs6QIuof
/QQDG8/SQK/XKqrUHsaQSwCrIPM4aMG9IrqwrqEdHYlzIarFbYtVhHHP3uHt
okiJVyVDMZqciBqmudVejWIuhNbXzaNOU8m9wlzAZNU1+9WtFAVpUGusE+0y
UBcL5aDVTUAk2Ssr3JSYsUG/i5yAj5x+VXu66Ju//BlNl4ASBIM1LrwCinuR
nfSI0/wQBCwm7VOiGn+2mhQ/Zi4yURdDvXoTOlhy5lHn0hNQfmUeAvOqr2aL
2EwqKfKF2VNZPMpbvtym+Po+5TFTQu6Ork675bi0sTK5fcsheD9ke8n9mb/S
Cg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqfEBdMKgIR8p8s5UTKus2EmbNkza35fjqNV6yjm7H2R6811ce9BtjHxAOnEiBJmHS4dtIY01Zg2mRBVHwlUxaCRD5xMmQPQQ8dKYLnd8EVDcWh7gvyXmnMaFFOmF5IcUNpDNZiNTJHo79OM0uNNJ86/3FIOkiXxStDApAHC4NgxsovIay3xOpMAwzPSaSRIsSv+X7hmxy1+OBY9cYVb3GerWRlU0wyi7IfrZ747thRVpLI88O/RrGKeLeicNitfPq+C9hR8Mu5e3cxakhniXGjHvfnTMf6ruGoSYunFXQiSgxPP/cNSvRkdEIDeOYCn9TS1gPWm9RKWmyaZFXgRODxV13tUZRDwQihFGu1ezeBZ7anTHXxy/t64Mxq5eRt0NOpST0M0V63x/pSyjBHzcE92pnvkS1o5fgmjrx+M0n+Dh8eTS96nHEqAL7KDzlXeKcCw+rpWMgqUYX1yLZbdC5FXs0Jym4MBFObsi+TIq9hGpPA79nub6Fk1C4rVLXJ8tDslQTJ+snwJTFRyvtoyrBKNX4LJ8bVI+ZW9VLUemD8Xp1nBG5yICXDxKP4wZFEgT+fNAKrIfY8w/SBkehzG21NgGKee/62snhfuVNQpqObZIzT/Vv6USPWJW3cXBk5XpL+2VopIL95nCrdBbmnw7nXvoGYuFO9Qhm6ZjT77fpc6dRyfUEAt5LF68NyWTi86C9tTvMMETPnjhDdiunDLPOtzi4UCeQD3NahaLFuNLWkwZxWCMI1uPXOXXWJAXPBTsrtzXQ8cnSr4rcWWYGydYARZ"
`endif