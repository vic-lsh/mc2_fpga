// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nJi8+4WV6/tPaPw472FaTPwTBLUcjoW47zELgk6ahgay8XP9y5skUnbO7pR5
I+qfmAPS2K3zIHpn1+hxxO0GLwk7AhDdvgv+M2vyi/8mJh7NM88hvgIzILKX
7vowus4uwj4JsHikVUxzzB//+cstTEtDflQ/eXcSbd6Hb9N4Bo+tIVJ9j6pN
JSQ7wxh6J/+S1ydEsVATecBxqQQvD2C0lbhO2pMqajthIv4n7zbVs4PQ2D/O
miDec77ryLNbC7nYUBu/jTQyQpsxZHCYN73B/8m1q/f/O9AbUQE09F1frf8o
QL/lMDk4DMhPG7IBTZiLdAxfvnaB9c7C9W0qfKvCOA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Idy78mR9DOtub1xFEMqsChQTBleD5/+4dAhsW578Jf5dTSh5yWGbAfFYmMtV
RFS77UG/Vse7sdqJ37fdqNOwrDh6vNoYCRa7SLlXk1nNPrfZWclXWQc+EAXn
0OeAf2xg/VnhJrYdh09TQNpv9H18pfwI7WXqXKqhMPVfs/rnGmvBqKV3mg7B
/Zd03nbDAkDcx4uqQiXQl351A2avAS5bCLrberab/pCMTZpGViqd9oOr0Txn
jJN8i9Mx0MUVXSn3HqUUtFZmQL/k57J6gnROsUvN1kmTTsRzuJmwMFjOYyrZ
SpGDM5T56WcDoMj23QxK4gGgUjYijDDjObEfxfo2LA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
U1DGHsK96K8sAKwBsa5F1gfOpMuEAcnq1M54LEqExxMZt89ZKqS09DySOclq
GhAzbT7aXbTNKACD6oB26RyuABnG99BQbJpBsrIEe0z4FnlPmJQSz6umHZUM
XrwYut2LuaRY2IyEjqpGynyfEWBJrf06khk9st0slZP7+uXRjK2ga/4WRxR0
CrF1lnvZjZ45yecMl1CnU2QBJdU7uBjrcEbLkOGqRUACrmBXFPaloW+8IPvq
Yh+BG97qSIhP26tXi8iQw8tPm4+F/KpicH42nM2yS/8Fdshe9+hy/hdXw+8z
9onVnyJWvlpDbPG7klPT3/PNTyLhhBJmtb2Qu/XOBQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Mr+CnuNmKCU29qNDDJfZ0eqG0RZbfJPPlhvok3mKIpsxsBom7j7CjBcmWm18
spGGtKdng7MmoqYDdhquCi8OoKtCxj4rOV5GcgZQ7Fe7LxLiGj3ybKlQW8dL
YklL8U5FSJ5p6wR78d91nOGxWeWKABa+RvMeJpQE50bOzQ0Wo3cZGEZehhE8
yNYJIJzZA31AusQPQWIwMbFUkS+mMvG3hd6jbYfpmBI6YJ6frR7mq5wEojKP
ec4L3I3/Fj/afL0zTq7lTPekcuJp6OGYxFhQDwOzmmE6ujkh1QjBd4DvuUry
mR3Wjtc6dloj6jc0JI5gB6CWdYyXjE9BImgyV3mU/g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ipEiSIRjLEe6u243pAXIJIAR67mEIldyzFHJPGwMXAhuJCXKStHzMmcAFtXR
dDHxb2kW2fvarJNE/GYmZ6bJR/e62tTfZEVjYmgjN9Gcyx07Cjjb0z6dT4/Y
WRGW7bMFhB1YTGLo7mYMDHAIk6RvTF9IkpyKsLMpHU8AgN5wxIM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hmbbEVXShp6Rzcq+nLktwA5SVxMYvi5iVqNXBAU5mtCh0iqPIKUEbSV+2lc9
+3Owk1S2n6HD/YJMb9qoZeY0UF5UkCqsMLHbjhg7ql+TV4OmDN3jE7sJjlxA
REeEp1RfuFWCYTlhvfRDj178CW11WVul6yhbZP2gPqd+Xu30pGQ+OS9m7p4H
LVHLtALFm2p2dyB/0YlUwAeOfFLOofQ/yWecxkaFycwvGwNlLNmqox9nwHE5
+pYMY5L1jx24XIQYzwJ5BE6HNcsM960bXAjluNj3tBOJt3adJBW7JxFM8gnw
LVSq+1yJcfmVJJrCJ5b4b2RwA/ayHOTxjL723NhOiFdHWj0Ca4l3X8PgnvMd
UnIVGheTN2G2lZlPnTYcZ9BH3reu/3f1zWqJ9mtrB06U+6yz7Sguum+EQREG
NfEDq78FzXUBThkt+k6L9+y6QrYbD1jRtk8/OcffpmpbUJrRu0XcrJ4hD4mb
jmUFxrTX94wjFpmXd5UpBcEUWBRciI6Y


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FLAco0nofFBqpUTt2/oZp++PYwfrySRrL5inIY42sMLcpVcGhUrGwuSij9eD
z91UgrKCidBhoKucamUmMEQRzmqXZ6dGVFhngS2Bxsq3QMXx7JuU08/xMv9s
l6S808s2v8np0F0u7ktVEfVbQdoayCOY3gIAfodHMl1Jo5/VW+8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
D5kguhnzv4jLaPblFb/2w0rHp43auJv/ooA3Qd/2XoXd5Btz6qK6Yf3j6Ozg
23tzJHn6NUZDCWbpKz4ccAEItZZdvyjZrV7t2x4gJhq0Q1ecXupPtR9cBcMp
jmtFalM8kk+LRfc6gg7/jiwhm4foTbheUBTRf7/oNh53thmYrQ8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 93472)
`pragma protect data_block
ZgwSDr10AwzeTHu48mhxyuI3RueLn/uZbpGJ96t6dbsvmKO5TAIy8ICd7vDw
wrFhNRRjArJCaMlSvxxxv+olQh+igPTL317/bHwgNOZJqll74yo4dWxi6k8Y
4BO6rkT6q8iGf1D6cZbqLiBx0Ywn+CGTAO2i+VSiDClELGsm2kcnfx0+hf8v
GhxBum7BA1Big8umJEW+bYQbqdgs8vRgDbvlDzDd/K2Xus80V4WDvMCjZ2+4
djJeJtop7BdG3xdCL/Jq5cszepelmU5I5JI/J0lWvbN0H3aKzVZy7TIBnL4u
OkDcM1JesGCdOYhO47w4Ae4uS1cWYn5ismpSBQrXs43veHRrmcSGTUmqCeWH
poeTZ3DofeU0AnbzQfCvK541gip/lQ2RGNKbAkInM/zMNN9rKa8XNDIEnIvB
949Ux4AAle+g+m53YWuzCm4WRq1K4msSmfGaEQaWuVkw7PvUpP2NnVpXQ0EB
E4QSPK5AkEiVozEOrID32PrGLmy5eAYMnOQbWMWwq/qhoTngJJhQvw7X0H2t
0XEc0Blf/x2erPf9NvwtyFNNjROsRHtHv/rNE0R26tKh4BGWOtW+QuRWF49B
6ABq5+eUPn780FUykgFCdKhwd2VWX935BeixHQrQoFar9xeUk56+oQAPxhHj
v7OG3EfjosL1pmkolrA66K0NhBuhz74pRjoVIsyf0jRCNHuqWGpSvLyyr6Tk
JSCJuvHeUlhrTOm+N1oQ2ryXs0ajAoNZZVK0qVPgPfGR9pb3eCuP3WO3N9Zu
al+sw4wvo2fCDYxwAMlYYeDGJlOYEbemWjCgSBJSNvs5rKB2CwLvUJKHqKtw
4nesVD9dfj5kfAfU/o6LmSK4MD3hcHWgxEsCBH9TnnSb0VMmXUmCw/sO/FeD
0N4StSgQCtPGM/bWi4sIINmS7G2Fop5Wpi7//w1Sl0l4+WhI9Wt0T3sLWYS4
jfgFGWaHssUQ1NJZl2ijoGy5IpWZcOTtIm8ykwPQl+Hch3nUP6v/MwqcqGou
WEkAghNu7jHTp3F57/guqd3LVUvaC4/8RaG8gX6E3Zpde7IdL5BDGJF/xb/M
uQ3MqGL0l52Y2+5fiYMf2QXrPnxq1PHrJm1XDlgLkFNcwI93ri3QVcoSA9eY
qklvR7CELdSSv+fiPJsgRivGR/mWJzGALV1OuRM4YMnpsi625ubLF7VEquVu
7La/cEtcoMqXoQSAa/2rtjpxrWVqgRX1u+k2UKRmMNUz4wVK/Rt6N+FcIIea
FxgRczB3AVfFkHBM8zw367ufSS1NtMkMIKOTwdkANcGGrx9BlQb8tG0ACkBX
CWMypmISa3n792gCnz6B3Mo9oUQU+AJxLxs7SpAxkGsgTWrMnlUq8p/JTLW+
tlwhmS4R/rnRQMwWHCMsKATDApcGJONifZTp4nrQevqHWlbxKJigJsoZGZX+
Gs7K7Og9rgTanRxofKSlx5M0yXqq4qnI0lwpCQkWttBcivGBccXYp+r59xFI
N5rHFHGSaUwZKxidazhaWOnSwOvdHZxN8OtxH2rtixJaXDvf9HKTFJldfBbk
LyM3zMBzSSAXyxcT36yS97N+I5AYHSxozN4jnG9dRSubl/0zEFL0F/pi8VoJ
VoI/mQO5CxDWYXtcU/iv4AWLthY3AaC2lM2qEMMUMFexraf0mQXkdAbuGwKU
Xkwj0BZC9oZ1O9BtBSJSKhNY7qH9e+gWxnSilnN+WTKIJHVuUUpNUpxp9o1Z
YR6UP8+7CuKmpzIscGgYY/QPvT//KKY7vl4PFypsIzyLUlkN5rR+7e5ZzUSR
frde2KYjaLEbnTqSPN2GqC/U34h3LOPiXvdlLme43V72hGF0KHS+qU4++dN8
bWZt6/eoykdfaO5s8UA5ssecMxWKi0rz2iwEAvEU0s7klRU0Vd5BAdri5M1c
dg4hpk5HTW7gFqyIECeNmP4fdiXRVCGmccoOlUdfOsbWZA1IlSEFzSMdwVEa
afmO6vcHPm+raMwZGq+1Ui5fM4bwwDcc2PPU3fPGff0Za/9+vAYmFhY4AKA3
nxa+M3XWEsUXS14dlNthZ+T0UODJ1IIOI5RcjdDK6PhVqPfbDWUpN9kduR0M
0tm/ZgC29zkjPJbvInrCt629MRHZuTsO0qAKKIhfXH5YRu8L2CDDj/Yl9JN2
VpOcYXstCdHyvrkD5JTom1HQ3w4+NLzsy8w0dN+FXywPB80MjFCFMCPoc6kJ
PGgbYPafvf0R3wYR+FqNZbBqYizF3Q4LaG1bAODD+wLPEKf4UOtl6101P5Om
Y3kLAQytv+GI93NKZWcvph6Fk6WmfLHj/i5CWJTL9pudmkR5j2KhoTg2Lhh9
Dnjv0kmJRDL+ntqfT+VhcPlSlfaN2gstsAwGKfzdsbOJFrcr2nQTV+VsxSXv
7Jn9O5RwDpcdH+RC0CxjOKng/41aNMEpkKUYzhxSAUYk1xSakjJ7RT/eEcTx
Pk9jiTV1N75ib6+OOh6+eCn3SsC+yWOQZnoqbUTJM1+dMohj3+wrvUXLQII/
2p7+dq/ILqrq75zm35DUg5EXGWjUARzA6slXUHexk8pVgwDxK0D/wkp7jz3h
8mrnp7XkLj4BOSUeaupUAlf4wKlYtKMenKWHAPWkOgQpVNaD1Uxk05KyfdGY
bfid/zKSgwZz60ggraP13Fd+h2DLGGE0AU4kgyLlJnNXaNdBnpLITY012CI1
IWrXcWqXWEpzwNCNd/uVgCef6efpdTppB4DAAtBi/k/NSRFJ91DnsXpWxA/M
Y0ThnlbM+Dcaq4QGtBBSr1qhBbQ5r47kBNWfrQx1UuIyuk9XQ1LPMc03Ox3i
+Klz3BDhSZy7dMDc/Urf1JnGct0yR9faQy2jKrhS4yApLE1DEuEhDch6V43B
+Q9CflJiA4BEIxhPb8gnGumo9PnfOPzqipYPrjmdj0staamNmghTDZEI8Jmd
K/QTYwsaEeYP+/bJWH4h04DtLEIg4soXYpKYymP4syF36XA/UIZ2JmPlNWy7
Wenn5S59bvdg4+96LHPUch+QyqzRnLuOiGfyVlWUQMofh3IhHWwgaYsl6KIV
3FyNTbVL7n65NjiiM5L19NpKppyQUTv5VX83nhCC/KPTUGWFhMpOoNF4qhXY
G4PQ736RSlprKGhetCry2gngIxU3bYTc1tTg6xCAYwkKgQm7VvCW2JXM+82x
x5rAJaEErYSdzsBFP/Ar2Puu4hL+pudmlAl/HzqrcrAx9BjcnjTiXe3+fzwJ
VAhPgB3jo5ek/hhD3KCeZEus6HwYXxQJGbjhgT4md0kFC2UKVglmajPrZmKE
KHV97eWyWrnQp/97P9yMC6vc1gJEReE5TyLDsn3HuM44hYlOqBOP1IqWDJrD
rweUPGgQIPLMuWkYk5a1yxGCr+2YqoeLMD7Z0FNFRxejU4GZYy9kaw1DgTZV
xE3QOCIeG6YxaSDQhElMSllch3F76TaDhIotarFOXXiToa1iw2hqhDVR+rM6
uH4THgoPmtbX/j7rnOd+ohwHvSkWAEk4YQC6PkSMJIuQMO1jEKPyM6cwAMd/
00nXCp9GSbCTKINfgI6BeLCNmemOzqIHzgykEbE9HSDpfZI206I7/IWrdZLb
6XCWh8p/yyxddKeBij4iTxzIS6SuhCMMhaNun9LKdSVO2pZxPlhNES1qdjJF
RzJ9zcr4hhTru/TG50mENJxbnLVPeCEQ0bUTEl68lSFSoE7V3svsckGlaMRH
3eAvZjedMe++pKiOQSFyzTkJK7cOyMycJJz4beQVE2snElyFB6CbX26+XheN
/rCCPbsJX8MFciid/WpDVMtr4LVOE8kLqe3bRQflualjaB9LZJ22g92JOCvG
EeGOqhiDT8V55A/084wPFulXcQp/M72lcAsK1h1Yc/mR/O3yrvbDvjnihFn2
GWyqWddjeKe6obX8GCO62u0Akm3AtXyQsPTTPZ6J0AywWxGeL0TaEejdJSH7
GcP9hpjhU6FiDxMIOYbnAt5IR+QY8t50CcCLmS0sekWX3vyUI+4Jo7TH0Jqt
We+Q8Brc5N5OMBvp4nNNp0NVwQRrH5k2OFQPCkFZbjD2cXSKXGQ+U+DhBAYw
XLpK18LnDyznRmUK35dLDv7u0i/LDrRbrJTpbRUCHemI3HKuGC0ge1T9nFi+
/PkPmgSlDYjYUs98LT1qtnSSlS36xxBYsoHZ6UwzTOCrB/Sd+4KDwXMdeH1W
Vc8cXQoesmlSBU7mdAON6ULK3vVhYCZR6BJZ//olf85ltuItMUblqo34++vH
Rz6mHFZIUGRoGjm/76t4Tk82S0G11j4isI9FMYg3FvyJZVm84aoEfXm1+xat
ee5rTEjVUyZQ2O9LVvnKkuUze51IHYMCjeT4EfbJ7HrQBhMLZ+/YnYYeJkMi
i4TTaoBZuDAupNFZGcOHhzEOpSMxLOWpdLQq1E4n22zjjAI2MH7IY8XFy791
AxX8XYYFrXB8eBZPPnD6hreP3K0Ap1CSfUJ1/iXuDbXx6/AI3MRooo+a7ojZ
V0QNoz1YuPhnv8RJZhXRkLK/qVirK+5OXwSAMXtvHm8RZoRW9qaKjr/QPmfi
XA50fMCB9EcoEUIrSf9590J4u5sttT2opD2AFbuveIKuG8KU3f815ZgXH9TR
m5smkYXsuSvzIVcXQJPxTwglbHC0MWupJpWHtiE/GeCVcuP8nleqlzabuE60
ZAZd1VzjiLlhCRJuUlJiAQsa5vHdwCcHAdANfXYf3aRWvUmYG6jeDMdlwUbW
WmYqkPm9XzdqYmWabvbiErLmIXMXXinA82/76m6f93Khafb5GDV1h4Is2AQz
bnJSWNiHiJPmgXz0ManC/SXTVpiuKNcj0o+lJTWNTsI9ykJP/ogGcOYdKCYy
YOX5bX9fYkp35z45XO8iidpoZoRKHMBmrCZ+WXKy97euemXlRbohmYLNXE8L
d7Nfw6DwicD164UPGtelTzBue5ZmFTxdKbxrW9NDKtMySqFwfFcn8bXBYrJp
Z92Yalx2sea6AA3OiCdosDnJ7Ey3a2dpBnZU5jostIMTiN2mUNnrrmp6eXbi
gG3NW2hnt+WVCnYUiabLu8V3Dt9qg8GX+MFv7MJ3z6dAyMn/IIg+uI2l51q/
tmY2liklo34JpPQ/hrYRP4eklcKeTf40okK6G8pN3pSwNrPLd0rZNEhZmHk4
JNTZH823JGuTXhEhuom+BQ5OHAG1CzXIPRgkG6ADf8EOg6cTZSDFEZoUKZX9
y0UAFoqdRik6zqnnHNEy0mc3o1nYY3VLb+mO+X2cLo2fkqzhzBE8fOtTGkPa
UDTxY2IIKmE3cs+7nPhAXanfGF9weTaHLzzJnf31p6BB8M8RkNJL4VtpUaD9
mjT4qKiJ0StWfW4DSQPSyotFyseY4PMtv1oNog0zLdZCEjZLoq22adCbwfNA
hz6Ai/Q/wVdXJJLhvWCFuvKnJJTh1I5uaq3d07fE7RjuclgKDC87QRBrvPCe
xz2WW6jS5svHsUzj5uQW6hYp627/y71J6Vd7AvTScHLLNVKAKR7sAOQLdxgO
Gth5CkeKo60ojLDBzwmOhM73hKu3ZhTwH/82EawQ8Rf4oD9j2KwWXElEFdqV
h0gIFB2I4e81hTisqHzXbARSIF7GK8opWKHJLMlQrQlXOMK/oAZxW+z3v1h9
KCO3m8RAa2OxuKSfuNC4aa+W704d5AtzFWSIrr481Q5LtLz70KcVZrIpkz9q
97jpsgeyoibZws/VI9P88LTzclGepwCH+fPl24gxtWfOOm4Bh2/8J/ervrad
rMnlSIb3jf2lSrvmvgi9kWT//cs74yJQ3mUl0EZ/xaEj22/XtSE+qg7HmQyd
pkKFD2CqmT5NYcxDD6TTFkRoBgaZq2ZprXxtTh+GryenppVY441Ctlnw4Njs
lngQVnJ+kMUn9xQJKqUZcJKf18E49WCPQWMkFUXMRqIuRGF02tLjFjPT94kS
CScF+YN3lqFzKrZqrIGW8ygCwZzV4g6UC+f1Euaw53rUBeyj2Y1jp5jKeChZ
8uX/rUeZcnCsdQjKL+2pgaWLUaP8C5oBMg7R40h07a7s9ol4d0bx4KOD0PBc
+g/wS/oxEENsasPnStIdNEIDlXD6NlnL6lnm0Q5ZEr32xP2H32uKceYZOlLW
4q749uuI9BHh+7EV3njelx/jdultF5mkpMz8d9eS15BVATpvUro6nshSvxOa
k2uUYf95rraeqcXLoNBHTGYhpbWZU4zVyRw14RrbU6PZFRul6v5eCKZhL1zc
X8ll4hEa1CsEkuC2niEBtJsGGaSHC8lvVxmOdu/2YoY+EoUR70DCffKlDxxn
gIDTSccXg5EK3xljTsCR8O1ei0d4S/PlMOgAW8UQIPREJGFtxWMH6IzT+aPw
bYvJYGl6SRzz2QCZC1BRgb9fxKBTEyu8RIKXEWaOsB/HCFrgutZ44JtItLR5
9ElnK9viyhUX0Q25Og6gpM8FCvKKEylDsep5utM00cYi0WQw1lmj1US3QYY7
q3oAg2jyBQAi1WQGPpAYz7ePHGF0qq/e71jYu89ot7eWBwZ/SLSuhVLYuBpZ
ViAEKcj4NBFbUpkZqZOrEhtl2qoDU6Gdh8FsLmIQXAQnlAU9Gw7xGqrwpHXl
09ZjwvY7gVnkW6MF2JUAgLtf1V1eDxfPNE9TjLGbr0NiISS1QNSfNTRPxMh8
kk1xXfLynU1rGWEB5i2zwlmrEp7mTNijZBQSUnBS/RWDLfcYiBbXDfaS8D7X
HTpj8KlC5+MqnOu+CKrUGjeJ3qqEvxdOoivROGafT7GlJmAIre9GTmxz2s6k
IyIK49OdqI+REXrlWmBuWm5XLIJ5Bh/9tQin4ZIU3hFz0YtzqIohBUBWsVSi
fFG6S54GFvpK0MhNU2aQUyrrd65bUAjyPBFatGqLtfqEje8JgBRZXy2vsLgF
lO2TA6L51QFEhV7P0dWXLl/EZb1ucYku0RisF9JTkxoQ26y3G6JTuqxLWlqT
rocqeyQdqWYa55OUR19ttM7U4SVBF04TCw1Tl5u2ThytGfkGNTYM/1TR28Yk
9/IAUrdMWBBnqg8N+5XMWclWJn6pDxV+prsO6hs831IGd/gUGOoQUlNmzaIU
ps8eMmpKB43VFqpX4GX2leRmXH0+IDT0yVbmBYhl51aL8iKUAI72pvImjePy
9Y55k1wS00ETtDDVFe3/028YRZFqNQxDLHdBlZqFvhZGTCyIX7A7e+SFB2ya
3OXRl32CDFwzZoU4JZQqrgYonLRhIv1WcTq4NpC/qY0MN17p7fS51yz0HO9P
CdR5pKX+T9m4HKAZAN9ZWnmAvkR7hKM8J+EPOiSflVy21W5PDXiSZftMQeVI
g1GwEOOzFq5HvM41HEvo8HyjOA+Tah+rEUoxUnoUWBkvE7Hr724lh+yqFCOe
qQiSj3WiErG8ET++UXF1jYswhleOIathRT04WcqAlWepxsXImaYKMBKlTtgJ
Pdy5moPBGA62Pv96O4ddHWh3hjwTqv8iMiyeRGZTgEEh5wy/TCmoh6hmEbAo
4eBh6NIv23uIp5hR3WaGqiyngSc94k6XipNUcHVZr6YsEdRiPRUrpeX4pB7J
db04RDcN/D/3s24LKUjy+BIAXRdUKkMVJLv5UbXmmFfnB64ttHvwfucKJcPG
gyX0UTiBuuWAtG+0T+EZxVT7J18YbJbReZ1tRcSB05il+VP308dYNWLhMg9y
BNC3ttK+En4MpTO6SAkaZ9C/vnoxvVFbzIsFB0BQmv9OwIVuZRgLf0in2uuc
7MOOSiRm5mWA5P8D8Qbgux+go8UmMciW+I45cWOWlJbPmFFLA/lj9jZkjle2
HWlL1LPbK8VnEdHHsAvegyiZk574rsQIPuiCeqTzt7vdjjMOPPUcYLMAbfx9
so7KmwmJSqxjqRxDDfsqdWW0nIntD18jtz8hpKfUP8f/COlXiX3ZPwfvHbaO
WJSrZAloW/gQNtCRptXm2FBDVyG1zn76DfPSHMEpR6NGOfallto9FFJBmZbz
tFuLT0XaqspzyMMS7QcSkWDcvq6XEje8yBCM8hETVvrndTLTnsuDiCrpLrPg
LSKT4VtP9SwJpthtt/ImgVZptRiU0SvoudlrhgUJ3XmDuv0NrM2ePst/V5Uu
/9fEVfaS+IWlAUh8hPdeIHWXfPirZ8vP8pYe76UOc78nnj4+rj+O3rYs5ys0
1ag5cUzGnhokqCvePPeHBCzQC8kLHmn9dhuqNcVoRkez5BzIJ7lFNu0wSJpI
OVLosZ5bNgx2RLKtoqUK7XBeZpeJXut6fGrliZiM6hZaWYRqivphXB3GUp8Q
5Ge/ud3R7vVMTeNNyTz9Pk6lhXvcAsGKu+2BPvv7uzQXDkronBJaJFM6i0uf
l26GbXD1MHv55OKITGxXOYOIbXZSX3yt0lJoticT2/VSa9Rcfg1s6nVV2LoU
wmp+oLbyoaOhuNsVHxdZ7QwlBiX8xC2/cy6cnsfLfREDInKGSXxp10/Egr2u
fgbmw0QRlyvDT9mshryuFJTrdLmsruZzP9p3iC5+xMeiRXihdpvg/lSf17E0
E04LAtAgVVVXMK3YmPXM1mBHiGWqZoS/xwp3J3KB2FU3Pff5YBBPCJ7aJNDq
MNkO9l6/D/tHcfl2x3Wuq0tdUEzZJt8hFC81VrrGPoTLHGRHGD56KqRbO5zC
R8BdIQp0qT3o+qYdGCNl+qlYidxPse8tPW4dkEUn2VQYgRoLDrlO+9djEysO
ROgPMNjN2GJrLsN6Qg87trhQtcLcygWFd4I+1rimqVglnVlaxZpMwdiHS0ur
jN8V87HWie5yY3fySkRQ5h6TjaXGsp6UIsXP7j3f2F0QKt6LlZPzaNDzNzbQ
adCPC4RwyoPRybcdqvTv3i7y9VChyrgHPZIAEBVirgeKmME0hB86Tj71lK+1
35eKNMLOk4nxRRxKm9SNdF8BSvEJsCG1cH0MXk8dK5NdqbAS05aGzAcc8liF
KrYW7jerHxkE6miSnAFy40S58I8qdJvflKYJh41Zq0evpD3Bj/JUim+hj7EP
sIR5NZ4cO4pHR11ur1pgqLitNvA18pZTBWZoZvByC00A4TXjL6YOHIwu9RNp
lOIKTiCtTOiLpymCFc3PSvjj+M5gqTj8gytWLwJ+eHfRAvQ+RcKFim0OIaFA
cSShI2IQ+aese0QgG0QSTeAvQ4BbpwgwuB9JqWgRKhJg20c4QWCFUiRc/NDz
ld8x/5MQDO+cfUAYIRBYmDk04HkvnktnqCNtVby6cea9ojJb8rjRSa5pi7IP
BsFnDaX38jyX61JXSJB+BgsXK2UasWFyBv8a1Ldljd/pjL5XbeGJZPxX4FW8
m7TDxGOvOF6YH7yPt8Svm0w72oB+2Sbdhyuik4VPdlBqEWgITiHJY4elyHk8
vjg5F1zI4FVAzvLb84jKJv70ZxVhAe4w+lJXnGdv4zpygPHJX6wF57no1NR2
UPb3ZP6sOlHtREfF85Olal5e43IOMZpJcOd9H/9kQG9Y4AAOsFtuwg5aJQsy
DYrLjL6yzt8J/Sa0g2Lz8aj9zvYASFFwRWPll3uKcq6orjIT2nT0PAHH1fFB
PsU7sSu+5G+pEss4y8vz+XckVb+lgjJhN2NgiYjNy7fcA6vSvSJO8IZ7XzTU
LeGFRicNIjUia2LzvdCNvfwY3QPXuw1PhARnYEdoKaDl6R1Gu0BwtK48Wwc7
+pFHpj0xXNa2pI6di3zYTVKnfYtxwmvTIK7b9lB9i7Ck4tmzAhrE+Slq/ypv
+T8e0q/0haDUdHusgZ8N8FSIRjItLeNQ3wSfqfJ9zKAywLdQFEjCLeHUINu+
3TK1A8R5fZhT7HWGJP7cAzeeatwsJX3UpXPrJqMpidI7I6zXL7sM3l7DnULK
KBIGO7MaUEJJV4IPJMhFy6zkzaP/AFIAbtSCIFKRuMJ+AZ2q118u62gAb4rj
vTknnA/7p/8mJjMgqxN4LxlSVL6HF3MlgSOYrNLBNHjsbqqLpC58XLBKp8bs
wVwHS1fXVc9O9dzpqsdR/vG6nS2OkaQ1SyfQztP2ehuIeIU3iVEqRcfxO1fF
tlOS1kGHoTIJIACcbEUSiYR6qqPmv4rnN08uxJnVjaKRbTkF+BocJ8ZklamM
XsaHdYSDXjhdxF5BfPy1VCE9vWyf2zoDnsx49ubYQ7NvK6r6ttPdHfFvrKyh
tjDa/7fh+qa6MCwBypyRzfpC78UL1XqHFh2lDyxghXO5jt2FOgLTRCZdSh8g
2z3rQFz5ZO8TWQAEj0Gd6Jn4WBlUqX1thxSdHxa4cyLB42EpWCXGuWo4vHXi
Mq7xsT1bvIu5oFZAmkba0KvsF96eTshUKQMg5/Drv0MbPfg2RRa+VFdu5i9r
rha5QYthTjTYEyrgzMeErgJaH2oK5csm/z1v3Ub0Idf0gs86y/lWdVPVdO/F
JfxNDLZe79xrU9cjyhJOG9OiAgLQosgSjYSisVuAj60MChgAnIZ3Wb18h3Fy
wrhjNaQp+x1w2pZ9TycxLs9mdVDVoGi/4AL4o46JGMWaBQTpJ/aq2O88S1/l
atrZC7yFtqmieE7Zsdt1z9h6j+WQQs3weEqD77Tttyd/aRXeTQznzg6b/qU3
eUPVFDfsZOHN7jTGoBdwWxE5LfWAxxgmJ5w1KgICLQCNo3JZ3b2IDlkLGbeT
jmbgZtzRfSYHX8wJN4RoYr4nXDK7Ix/AuSImMHVLhVGC3mhUybaN9DL4/j4C
e/DiyPETtO6VFboSUY6IdKF0KE0gBEjzvth9UphAIWlQBL1AMn/TZckAowO7
qjuqsHFABBV/cvd3H1S4Ee2oc5cQ3RyH/BTgpSJTmf66gnyh5ed4Z+yLoWML
wxrcPzc3CPTeY1ZdRgKTmUpzi8/WwbuK0VkAnZXBoPeL3U4i9G5VcAhaSnrY
Vr5eZ4znWJ9H7YwwnkRQhOeM3fPK5sBftAIrIhkYzxFjLlSK+Rs4KniaKWmz
a1XdKbk2erqOUUxAiHkPLKNZm31w65aMUK0z1DCwEnH9N1ALTocqrhF0lDk8
oZNn0hOSTA1vKHNhYzGbg2BI+/Awy+L9KpaDKw1orIxLw8lDm7BiXev8b9yX
co7m/jvuhOSu89T6/LvYG8Kk1atlldd3fKTiyvHupO7DGlBH0RRnb/X74RtI
hY3Nn/Io4qBsh5PQSYMAKlYQY1RPBhBODXWFLigSxd+4KXAVtI9nfSeTBxwF
y9YyFRgDqStAlSmm313O7V+Uq+QB0Fq97vK0UkneDUhiuPz4rB+5eig9cbp9
VIOhOgv0xvjk9jQqUgTtJ/RHXIw45qMJghwQJbfRtIex/hbHHyvk41eg+21M
RKp+BqDFvV4Tarki6h/BXW28XZT+ZeKxLDhoQOqe/H1KHmvXDVSXGL5JjSUr
joRcvUlJIkCRvCcdqhghTbYqHSYcXzywhkrhOvjnXNuwtgpuT93gcFp/mT0W
r4cXTAIqO8rPxlNeUqPUFXdfYU0q2yob4/85XjTmnCho0OfoV2yJFv/Axb9S
fuzt99bTzsq5IWR8j0q0PzbH9GI6QGir7Gulc7EDMQqoufCbKdl7F4rA7xI/
4IyODLcL7zutMS331G34QJXjXqVul11RAK9JInDLkedbos8GqL/a9YgSashz
PBWp8+aj/LAQQHm022bXYCGmyKss2pOGf31vEU0s00rWIxm3bsftBIbaeCIE
JkgXayxMB4hBDZWt+AGJG/GmxM29kZzqxryTQ/+ot6a559Rh99/hrFVKVXP0
kFQ0aEOvg9i7IbHnMgmfvetHvSnRyypef97QhRbsMGJtzYbCaT/siz2PGfCT
uBNzP2p3yZmM9yJEotqdIlGxF06JNDl69LZETQierr6iInmTyBA+oX9JLLsO
+FS9jhHQtj/ZMqTdRC9yhEIGijUleb+Al3ezsBDq/nJp+dFXKLKxMx7h5BXe
FXTaKWfsyopC84NFKWRcfGgeK43FZ8IrjLnNAVoMilYvxMzXY2YGytQt4jd9
ZVbg7AGo5CSZv5nOUaMhIKs1ITK2pDFei4MCx1NqTpRE+byhbjnCFv+rIE3u
vejeqmkkF/u72dm6YbJRrvfKyQWwwXhqzR17EMJ/3Sv83JpR1xN3ZiSKUA9G
sq/ZSjVnSW1zsQsdur0ObbQtX38Z1GZKLk2MDUmNzxwqRYDmC3d0nE0HNuZF
LXANNguO2ePnXvdU09L7nOOIuzYcvzK6xmLRF7sJkvcl3PXqRQzLQfjwFZUw
iXH8nfWD2qYeBQGI+2HFucuZvyKFvHeOGC3+wu9sE+hBBty02USjbo8yh5Le
05ezLVoidRTgp4HaouAZpjasWY12iWGR1CbFDhK60oZS8RdljMgdDF7O7sMj
2M80uSCrn75NEtnqQFwJIw7Dv1qEuY2y+SnbHU5CQhzZkomRUNfwWB9yVye4
NjvkeYXfBzs7/Hot4hOrad2YLhBMXQWTnN7zig78Q86hK0rHDHXFaXOUnhV8
Voeg1jRi/5qPbXQORiFMqb8dxubaCVXWHtteQDhal3k8Ep7qQ5HH1IMql3G3
a3yfji/IWFTPr9jvyMhjAbBEWj+RakTANa4BKp99Yej9sBpWb9IoBy4DIUlh
nNqwzWgk85E9FrH7Yjlz6BpD2j9FG/vBzt22NbSRblmA6QEUerZFOccCrUpl
d6FiD9im75Li002dvSIFXAJ59LG/pxp51HQakVbAmSVjic1uGLytmXKVIs83
K+Ldjzvx1frOfoY2v6LWXBR9ZBgVELHrbiTZ63RVXBViuTuRsBpQp/cu7uS8
MXR8fD3qx/3wUtXTvh2Erk390m4z7x5be6GNE3uHvInf1/KqF9Xvx+gw3Ips
o52uGeu6Nd5h90sPeknvSl5vVhlnFF0+QEOzyGoMpSTO7Hb+FTPcxeuXjXKn
9PcdelclTQNyMPxV8gYuwwN3hijFLePDrbbY+reDf7Pi6/ohKb/2MGhDjRz+
fw8oe9iQj3C1L5BpM38rl++A59/Da9M90QWraTnPoz5wnV+xVC+kBJBGJZJL
r1M4dr2czDt0pqn+Kdr4G3LnvVYFjgrDLkBMYcRQUM/GNxo/M7YKhRV6RjyW
3fH3bIEWjab12pomMcAT2KbJXBd+o284EXtRRPHxjv3zo5YfMxc83O0KZEpB
uX5fuFA/B5OrNYzjpPoynfEVO3+B3QAT0p7vIc3H0vuw2/2e41uAwDVf8HAc
7DTZzpasCHYz38FigYfbxbRUh+/+GDkxsPkyI8LjOM9iGmCtoR22huD0P/DD
Jh5i6DOWNRRrxmNqAdGePbFIO72hVlcb43MjgXaS/J4tlc9FmaM1qt+/dg4p
woQ0y+IEgs+XM+qBxdC+vqESmvD+aQf1vSdl1fCGEASndi+KlNFxKqcpfe+l
1oK4WTzmVHEqUadS1S8u0l25wdcHMSEL5D998cHmW3Cq4TYiTp5HcXMKbL0V
ckvcLbB3wCS33Q8S+l0j7lzshsE2lkrC/Do3MzSu+gjZLU9SRRi5JG7CTyYv
er4DpQZz5diffrbYw9ZHLj8Wv4TcdgVirufSqyBc+XQ45GXMR0UrBLi4Efhr
GTrEJiuahO+raWZqFOHCGsepxqbHgO9cYNrG7ePa2fMmBhyDOFegMhKJLGq3
J232FKZA9E80J6HwKZeeHAbwTy9rssXTlvbXpKAUNUz1X6x78cj816zvBkAI
gWohaYU/JXJg4Lg0QjZXSNfKbBhwrmMjaWIh1K+hW8AhoLR9MH5UIX8GMGtw
h1f60Lh+lIAGFrsfQ0d+UKtbKc9irXR2ke9OivnDqMKI6wmXYKKgok5I0alk
+T1Ebw7n5n2Dnxf65OWiWAlkopcfHGbcVjSjtOj4JjQJoIgv0NQjOWDJzPIl
Qpq6KLv2l17rJBbsddY5vJK4qdMoQqtZ3pdmlMAbrOLKRuWxTa3rER8zZ/1k
SyMvXFu+MsJMMlbJJis/GT8oM7EB+fmlSe7LGU/uLYC8Syh/nBTnlKScsxEB
4s/fmClRvPEBgATDEpkKwTt4UPLyDLls0i5NF5VaVYji1IF++YIxgVEIxOUi
Fhhs878bzh6967oZ5xW22AT1jja6h37CEZp7pYIIXhcsybvbF9Px71qVxwaW
e103Tt/JpZXX83VUVNnt2bNSyNYiyy4Rr+vKRCJRIx/pw50OOMQN9s2kJy9W
Wk0EAHM1DhoFyERraSEGxUtPGMIt8L7dkM7p4sH1ByJxnQB6VDaYAy/6+z9i
yTo57ue2o/zR/f4m3te4PwEMFVJkpsCWxDsEZZ/tyWyWmS1ZecxRWyk7kI/V
5toSNizpLpj8GI/rLXkZNyhBxPlHJijbUsrVq9ensrm5oedlgODLG15YTNWy
mvXAWRLPIQQgP/d4c7rJXyG4c6mpoYQxV5diZ8INBdPK3aADEmv2DWRPHyQD
1tX95ATUi7ElOta2yVFAsV/Ltwm+ZsRpJyGb6o5/9VGuw19dFtP58mw0YV8Y
3u8WIgSbNomP5anUTlqYMo0PCS3CXA/bu+NEEtuWMLzf0xI8AKkJb/FiKdBc
8zSX6RYmrfGhpxuNTp6ZrPk7Brdgl2HNMsdhlizvVemASr51l6j5cTGZ0ZJF
jNHAYFMBuOD9Txir9ZsWJchFF7bIFTtUoUD645FtFE71HlXSR8mFLcYh8yCC
Nrb/6IUoRZf7j5rg4Tzl9TaX8C8+1DHBaCFd2KmInoRA0tGtQ189nY3eJYm2
mh9ejykZ4R/SZN9tg34VU6ETwpM/4z6AZ9WuSbwx7MSv2fxKF8EEQPiYgEDW
QdouC+IGtol3c0aXH28EFJ/z5vB5nBf5sKYj2hnmigkOjXbO1PZdkP3v8f8E
X/yUKsoOz7P1rUtyUWSvLW8o6tE7a5cXllnAmfAZ3/TSRHAidPT+Iw0KrSGb
0o6K5nQo2leriiP0OVzu/HJAkjzB6rMSTBw/fBjjXcvvVqladpTV+TwZ//zI
H7YJdKwAXcS+HH1vPMAOAyHQRdADbHhEs57oEKQR7dpD2kflpnjOB3brRon7
RC7ZI/Qf740yg4sGTX0GjfBTXjXq74Kmlg1oA2DPK59IlFa3O05MJHHOLtpt
L3ooTDwWTSHynnr0lbJhWZcKWVdlicvQqZYzGDtgmU4oIN6f5XyDNabEO4Y5
9qmFZYhAwj+cG8LK6uw9IUQGFPm2egWNdxpiTEh/VufpPk+cNcUGWCdvToZI
dVjc+ocvc1NQrbtHEldTcaPtYbJmKPmdhWd36U2cq4fEf/VHhXrWogt+UAYD
3v+fWEvhPhTcb7Rse8RuIOvnhaM3FgiHR0oioUnwHPBguLyW+ctv20RnDc1l
IyMoMzLjScC25v5vKVwhXKUKYCctmwGvoEb+5xMSHd/hNC1aKmhf7CLbChQx
MhU9eVzF4K8SzlfXxCMHI4S7m8+XoQFPSlKs9C7ClQMJ/LIBxOo+qsWRvfbQ
z7MsdG3vU5YvKwaZdL+CIQ+PwDRRdIkFEKFaWTPwfIOD3exfLYXU1MQP2by/
u6hq5MCOveWMOf14zkgNoKsJwzREUWivZcBc04xKpAxo8Mmt3IBXOF4r6iko
v4ADqGIZTaRqDt3iFnTWh5SdpMcGbHewP7kqblIX72hxmMJwWtkQDQ7QlrzG
TJfl10NqDYREfcfACUDxH8GQjEcUaY2MK420rD8/PhVgq/o3poFS/VQZm3K5
vnV+STgT7gqCwoESMSeeYBBSIUgUxPuhLDe9Kao4hCa3rK5vL1paDGy0WXKp
4raHaZDysFwdV2cJKCiZ6w6SL5ANbNJcDsigbMeINMTRhVgDJx7WIXNu9qp3
BReE3TowxwTRwSaMnavlRClrUpzsXtTYnF9KVoXm8OBDkVAKly47wYR9eb6M
Gqj9c9E2atdgfL8DoU7ufjOQppmsXWSAQXOe9itceB7fMtiQloXyOUdr+WeQ
hD4N5zckaT5bIDAEqW3zT7eHH9mvufJTDz2o8oKaeUQ5Y0U0QCdlv9AJhxND
lIZGfAoWDJhnmH/VCD43KOOAG1T2NY8tVNyTen/K007lMOqtXw91iONoso1G
0IT4LdfiE/xNXRB4OeOByoz4HqEeNtXvoG2qrNHv1y2wArXNXlgjtDevYX8I
NTNpdV7d8dBr0EX8WguOk3X+k8BKLAlrD6Xe6wi04OlMTpTUrJFpLmiJ/IP0
audeJZEfjyQpqvECrH0pTmlgzp4n6uOFFIWdF41AIAYM1dKDgNR7l7NHwWcg
hBFrR/t9x52NR5XsUHUJ9L25kEGTSA+z7qg1PHde978HBYKADuVQ24tlX2OD
HmMgiHzZUgISW4NpbGq/yvCIo6MIaFJOmuH1zIVC3v+9MvZeF1hKNW7tlIlR
PUfvfwbAFQzRzSXc/oSXehhsVGQ26eqdh/+sKjepGl3+gJH10wX3bFJrOk6G
a4m0oZxd0yRlZajrSp+x/jcEYu7kwXAfJIGLkJfRA8dPi0c6aemwh8WBUAgS
djZFryELhO6zNi+X5q3WqFHVJCeAIwwhipoBuX/DKWjcA1iKImu0KqesglL6
os2ieH6zMXCRVlx3hn3iCgw1/1J6lH5hgGFTjmEuCyZUkpVm13i/jUgh7bZ+
WjwP1eyjhKvECsA3zTxPEa3RsBdOotHP0TlL7FIFuSehaVSmQ5SeNeEydTPm
y/QS+grTtBILVVvjz15fHIpGx+ebyGWD842eNw5ArUipmU6YWGJTw5kxFIm6
/iOC7kEffAp3w4Vnv4DpFHoUgXStS+XMv5feLfHvSQcwmjV1aVHUHOP3Lxae
ycK/6UYmtuExp18t6U+5jZIv4bt4D1aRlvRVbb/yz7JgFhahb9zdrjqdXEhG
99D0VT27JUgG0fXi5rp1mQ8iLjAU3DOnSkCi9EPtKAtGmAn9llWwjMsNn2yC
JPt8PF5PXWIJrc87Q9XMkyR6ngws7tWWXXI3/DYWJgKrVRyT/xu9m4BpAD7o
38pmNaA4hMtx11vo61cr5qJ485kY9071bTgMSyuOBGtte3rq0Rx9S1+SMqb5
meqLCuMJp8gaf32x+cVRyk/fntyFzg63dMly3W6qLmVDMig09VXy2Iz4ipef
hqVfGXElL9DMKVGNb1dNFnd+zvEYpYzi8ileivsRBbkJDasMe9GoGHgRnKZ6
YlzRBsOWIzKgdxjX8T3P1YF8CHWUSnzrG72ZacwrH2xEOWjW64fTBABF7Axa
VnVgarndaN0vxtOguxzNAiZReQlNzVgv5yuwigepPoIeqg/GeNxB9ee8sFhO
chrQwY3dPTLwbEPEcEErztqZg++8BKBdqc8MyU9pCG0bG7ls2qvyUkkL3sl/
8S4/8UVV9aEsbzyRRHtX3hOVxUdS5iDP7TaWDG7+JYazLYSlGAFKU6hUTBhC
Z1cAeo8VBLFb2TBIOa9suTWBhJ3BEKRAjUFHtumcVBj8SjpbyeossFnM6bKK
RjDiPTHmdcCXmUifz5gPmEjjSfnoigS4/lAAI5XCAfIXfiB9eOzGeM0e73if
vjCyX40tdwtCTfYtXsSHvCKQyezCgJg8WUj7/U51eA/kxKyU50FM2dfPN1ZM
Qkv7N4KpUtJhPCarGy2KhGtDQRk2oV23/i1tkdgw8bhXMr6rjQUH8P1uQYgG
GY22BJ4kPzYjxCps7QqwbFkcT0IpmfD6F8MKfG5lMOw4tHlZrDfkfzahoYJB
9KlMZrA/gkznsUfSNJjhTQLGfqq3XPj87HbEOzZS0pCd5R1594R8OMPV71zy
Caz6aScacWNF8M+SSxwx5ERzYn4vAltP4Dvu+Fxu7UtfdD84RtEElRb/i0Wh
W5rFizR6OxGJAsLdEncmd0vKlPMy3wLGbJDuEZUVVRK09fRNxXu7QHDjerAR
ITO8hEjbKbuddqSYtso2cmDLEl/JU6lqQGlRKb81JLemdqe4+BtlfTEp40oL
bFbED55fTzgkJYRnOl+6QkR3v0aOA6pDmZgPOsp1lAqkbA/sOzgr7YDk76VB
idR+X7BKSXv1g6paJvsRF0ML74LVj6b4MlvK6Tv/986Jhkp7XlctaQw7f+Xk
Qk/XujCmIFz0umtrvnG8G+OYjGAWkUAdiVgM7VZBgV6+Y1kczRSh6vJuYW6R
1wrANDCDPV5aajjZ/86WGvVT4ckV06q4tz04MxXpdvdRmCAI3GesaJTtY5Z6
ClvzegIKlTAuze5S0XQPZhPhrELeBaaqLWMaQ07FxMnbEorxdosJjialdQ0u
lV2zeqs4dBasWHjdDC/E4iqTiF+CQboVnMozfO6Txkmr46GRPLXbwBgVyAep
fELcIZ6CKREkp34v4fJAB0W2opj1l69iix7Fdl2Pt5fa16xn8ylGXcZoYKB+
dBmYoM5XhWbOCEt9sA7fh6ql9EnKrOxrigp/672QCbnOA9FCIaquvjftA2xD
rht4HKT1WbtXlvQ8m/VetQ7Eed16PnnbMykhzyUjjzDjP169WGcSBYJSDKBf
eG259EYnenoqxLJz/X3PfAOscw2aI1QwnRp9Fw11HLaKkFzymGjd1b6Qf1Cl
UQUdyooXFk/emC6/DHTqfbrQseWJl4vibfBRZOZZCaAHal0VclMM+c12Wl5a
iBjpnP/Ylx5FTbIdn9gWQdg7Wsbg5UXom6/2dmTeHsjj0FAkrCelOKK6ntMo
oM8s0MuFfxUStqsJD0ZEm92s4iBdXjsmBbE35rQDelYJOYYW3CTjenN8VUih
FbhKhitHWo67txhOwou1/1zO9qxLuIK7yryPQ0cxVbkXzFl4Qbu+A6g57/BW
qXEcF8oPgvCtYe5qcO3GhAHftcsAt2/uw3A1RJmTFIKyw/O9wmEnGXtNHx7q
SIkQMGoGVxaAwcmwYVk1Wy/W7vHY747Tyaw88T8iEXHvF6mcnOiGjvcHuO1q
C+7KEam9OOVyKqkBMrHryWOqD5BjdL8JLIO56ZB1NyqEnQFC1npgOOZZdi9i
Fki4+ows3e7m6kTqi6AlTpy2kiD8SjX6xeeDUxuDVpjLYxj5kernIunWcNIV
pi+rfP+vv1q+H1i2UOeEuw3hjBCYH5k3sVjD/QBmf5oH4Is60dTG0oH4sqPh
4dNBKTY0a/zCy2Qi31ELHcKDX/+mu0rxQ0E5/d/O81AQ5QcJCSxxodh3ELfA
erf8Ca/903L4AUmqE+Vvk0mU57vntUObUqkXj+C7wI52mjmFVrkA6IjuFiKX
1Sd/lRs+/c2LG0SaINI6Am2Ky8kaIXO5ToMRByIeaOhXBglc+Qdfigh0GCFz
0jGbTKPN+fS1pnESjOudbWbZS18vZ7xEY1nqx+d+RSSI9qVp+3cxB0TE9X2D
ZZZ7zL2xu0/Ey7K9RGB1pAatV0ePDXsQSZWCCySecNPY5TflKeG/ehEvc5Ad
m0MaDqvO/GeWTIJXAqDguOENhWLqvwiJK7Nv6tmM/TeeYNyb7r0USLkRroRh
SwFt39eeLHP8LPIAeybATNpnTwotQGmaLoelTuYcWwR7IH94pZdt7t/UQr9k
0KcFyOB3tWTzuwBcVoNjkwal5jnUYDoe0Q96zz4+1WVxsqz0ZIjPXfMCjoQ5
PN230ZN7MWbuUW1MkQKFsPlxx3oNlWXvFf0V6p5l4I3Y5wGMjSpoZ2elHocu
Dp9OBad06vlaVP26WP+FHlOI6i5w/wJPdCJS9dQYUXtttnw+4/lNyJnG8jXO
qXE/80Ayb+nxUdG1EaUQQuOH9pCPyAt6tNhglySgiidVGjR6XLSP1uzYZB7l
Sv0g2XjDreKpWtXaMmR+BEa5St4S4ZRXxGxzZACqGbbOaZS+MbvTMTTNjZXj
Rzi4KB49nXAwB92rmwNW867cMjlKvpkuXQeotpYWbWuTbSvyG+ELZnKAjdjq
915SG0VgUa8L2xuczZx1C/Ci0ctNs8RXM8zvaEAxiDAuEeH/HaFN/+0xsOW5
VULGyyUyR5qMavF2s0SamwhAcZ7NAvwrbp1+9x3OCOmU7PlWPmeTaBY/2Vgu
fYxaZa5FJcX7DM6Hzm3dO9cU8hod8uL3pMflVqeU6UCXQZiJnfsbWh4qemu8
FCy9gJnyIzNI9xFJ+3n73HyqDEPISAsKj0gcIPm6TgVjmX98GdyppRrmB54h
7bEewHEzhOu65E2qd4h8/Jt55Emq+xNlg2YYSMdTqdGZG1IzZ5bKoxVb8Qa+
W3payI4UTUObHn66e5DiJJwc0gjTRg1rE15SD4HNn+4S6a27rE7JreIcie0A
gOou8B7xmtkmCABumQrdtBtr7RLQmJL0srM6sbTgmwoZ+LuCoiD/dul+VrGq
+jCDRW6wufX1SwmF3MnT6RZRpCeY94Szyoioq9ljq3KTDIX8GfgSSKF/a0UU
umLs4uFrni930X+mcEdbV2i4JkRNdrBc0DudTTDZz7OP/piHs3sqc4XksYrg
T3JXu7w7xVcM6iReaZ2bDpY4h9c+ZILjfqxFknCHqJi8EU08C6NmOAsBC1oK
h3waaI27iqOfGXi8vxJB+lAqMMu6N2+lmFovd5s+DCEsUDJ6tdSfnhk9X8AV
Z5GBqGNJu6AAfu1+h7kzHy+l047q5nSAUUoR1M3ycu4Aoopl6rHmnJjTcsbo
kC6OREIK080w/dcwFGu8xNhlBk3v9zyqPrceLVqpmsY33DsRMjf1448LHjfi
hxiZDXjzi9FqkNzrh07km7ONdPw09IqJKcVppz5fFBHFlhvxl/UNxu4x1Vdr
reM3UsmRy7xG7BJaOue3uvgWO+Fdt/669dtORNRQNpqW7w88S72YfLaK4m6a
1YLDxgiy1RoOhqkCs1vp/dY0s5AvD4y1qOMAsr7Uneurm3vYVWMP4S+91/OU
/5LKyvu9d+KpLCRfG+QJhLkTyrzalVqTD2E/qK3EkWBqL5LI4yZ5a0fl0vYB
nyUhbXQuOF+GorsZFOl6/8thHV+ziboKXRvfh7Moi/t0H8If+3yCsHiC8YHG
xr9owMCsqxau75bryM9cWF6tXeqfFys3GYKCUHwRHd+wvnsC9liiM9wFZjBH
D7OuGHWjsdHISsQdPWp0IKTDph2ewiLNbS/HU0FBxam1G15bnQM3VzoJgVda
7UOoBqdYuvMObnqj7cxy4F+hJQapEkgI8srA6gvaV+jBFAbLLQAfsn/kVFwd
+KUypyhklokmgCHVqNup6UaN3v5Wzf+qSQ1/POZPxr9K7/Hh+rs6Pc/R8+ts
a9/vd5tMxgBPcmwK2crYnHcjr6yvZ8XSdFAn0svfrw4CBXeixPq+37LZVtfk
6KmV7GteKXneQLZLzS66ut5Gw1J7Fwu3jF+n+73vrfjjKgh2L91bWdHDYSnO
GIc/8/cKlgapCz9lpRymYR/ncm8uFQ/eZJ3M8brK0WoeNoSsBFHs684JRky4
6uZIC5j0WY6XNrmS4XWFkSGt6aDtkPcHRG5oBd9ykwKAj4a5QtW0w70vu/Sp
YKsO/J6Q6DwtyOd1P5CzfRghzfCM65oyGQb8Tngx+EusvSqudsQk82+aUpyj
4Aq6t27uGs0tTHqt3VaUlrfOg8xZI/WsCx0H7uLXDEg+o2xk4VOLqPXiPSx0
eNpSvywM9CyKuXECCGbQTnAmWdWTcZSGE+J/mJKUlatTPooZMKN/kvxCCAu6
QK7fyoUAKs3p2YkVhsqHkRpObq9IxO4yANa0WOe99qfc+adY/AawXAeN8+zD
X8NFRbHZqDqWcbmP9fK8ZfRz5d60OFD6b7zmN73G9icNfN9TeqFQAHZ3PlKq
/O5mYaM1Gus0CXiEU2DKnIdialM6E9qAl9g1k4wii/BlR0bfYg1qmFdnlfL1
hGX7P52sXzy+DAKuo9MmAiNttO6Md4bGMBDH9B15R38vQUi4K8XBlbOQ56FB
yhxYwWFwmmNXFQHmpLaupR3fbGgHzV0NdFXP88PfzXEq6KyeRUim/GHwR1dm
+PQ6Bo/2emImn6UnvVxggDRmbCFWMacocUFGDDVk6Nlb80webTuhMeB7gVNN
eowynNomSczHIHhEBgbjIPhFzhSa85RriEL8RLsUYGCo9sGsF78iPRF8gYQO
6HUWIhScsT4fdvqyXyem4wwM6kv0a9A7ZnwzNb7OV4mEKEuDOoPVyIZNOlYD
KeJ6VNt7lZmOvj76IbLjhxwuiHMEAIoqjxLxM/rppWfP1apx5Nxo8xLVAFuL
RMOvUXnGTwHbeOq65BJGcFmLgZhzxlhahc6vYpSpNFYLTwV2e0bcKDZvezSP
Cj3+RcJjQHcrqXDM3tDTfqMZpB9q70Z/KsRQgjEiKoo8fCYNIZTjIiACirra
sPFfCJ4iGN9eC/iR4nriESeWAorq7GpmHUCccsegsDP9Vxc+ulWP0b8TEAU4
yzCB55Odnv2ekDUgCxklklLsHj0UGSmGvKTRc/6kRW33wrAFwX5FDkoWF/Vl
FkNEp4FZWUo79e6BzSTqdX0xuV1ZnIkKHRfp2KZqwQaM9e3JpDwBU3b0fxqb
MHAA2zCzCOdajOW0nhOnv6vLJu0SWXaMGbQdrHUoX2BOCiGBowojw9U9LtTm
3rOzilEq7+8Ic0cKUGNcCTbJlg7gYKJfZzYmfQv3h/sduGwLutrTSdQ/jRdR
4RVpA1uqKOL+adA+DturquUlLX7fQ8eoYEKwZxZUlB5MqbiBj1sOBPU9LTFB
uB3peuvmzonMVAvuX3KwgnWkPC4utUypAAdO7w4+PKcXM9y4Dj2UrnOWqtzu
NKegOZsH6I+xaCYYSM1FRgVbyHlj+QHW3tj/2S5g5TZflqXVY5lElRX85cvj
kzTA6pTBC7CQZcOdYsUtX1DRQc6PPRQB2k65wjaWRCAmRx6Cv8JMtslQImXq
i1fcyqDVxRmr5nPH8sWDHxvosbFtiSJZJfreI22GUVQ/v8NKbTsBED0gbcMb
y9qoxgaFhkB8N38QxGRsch8Fz/YC21/Ip3m04cR1Vsp2nFL9skwrvr98t1A1
Ddm78ytst4HFlHlyI8r9xkMHdCCVSLLgj2jtHYB8eyeHqJF3iUA0Cf+cJLkb
gjdr9EHdrTJgdemOeA2mEHk4XO55I34K70nEHzbka2jJ+f3pzhGIOouIUK5X
CEvYNj589xdgwN6hcOUVKRhHME4pT1uKwyMJQDQ1qykqHIXwPri3RvmuvSoS
K2cpasYKVMz6wkzhLdSA5xjWSauQMUpSdW9S/qGtWB9vvxsNZQ057/wAyJAR
sEGMCfbYdShUisS/GicyYp14V+QsU/qGyuniQVUmKnjM6UEpZV1Zv2j1ituL
O3NDbuCvbw9aJfcnGeCtnOWpFpLb361pFWUA/FfxumsalLegjruvWtVUqUV9
ZShLtCnIb+yZfCN+8TpfIiI38YeCRsucXgmdR3YY6OOIXJdwEcmeWM/9qHKY
M1gO+stZy0N1KvWBU6ptkVSnRWHEjQGqTBrm+nEE3ohAd1qBzLzN3qqwqcHo
sneHlyQr1B26BRa3MYhvNaKKM/ONlTih2UrbBGzHI+92b8MtbWLYcZOiC42g
MC1ZT7x5wWuEl9iOSz6PLkrkrjeCslDKeuowkuU/E/Bo16pbr5MOq0wOCfU+
YBOuUbPu1lwcZ4M7MF6JhlZk6uhVxPSPL+3Ki9dggA1d0O6laSMzwstqfFqj
UsaMvy45s3qM7CjOQFFNXz3fjovx+hifWaas7UNoMb08GKlRZGkGg8qUq2EG
HaU0uLiq5sxm9fJcmja4Q2R7tyvBCE3ZSMXLzvQX5OGgY8Mtpxapee01jM9f
r2a07vVHQD8uNHnyD/8ZclD8A2BH2QdGdiDqKGxcWlvbKqKfdqZiOlCp2nbc
Djdm41Y0WT0nydJgtT9QIoTq/wLwzE4+T3LnZHwH6lKAo3CtfHWUu6B7lHMv
HnbhCdxiWKUGeyux9/O5FzkPJ8sVl+PA9JSKA7DEqggoow8dZmJkoyTSkFRV
AQYaB9FPM/EsrtRv93efIVDKz8Xn1CPcLdA9RpBurhQSZuuCzSAUNZj6QGqh
e5/io4qmUN5hiQFG5Ydx4sOrO9MnhrCePelxp4uNw8e6yYGJVQ+eyBrQzLY9
CTyJTJt1xiVpQ8NZfMtKAxwIhCcEc26NLZQNZ/t1RUs8U+tiHzNHiZ/QdoNW
1Ehgb2CsmugfHtWs3mZi57DZPiGa9QpFbekGt4SUkAyLaCiB/iMTqzXHcYiv
/FqvMQYrrJAjHDAS73z94FSxPn6F+JoE/aiS75+KJsGmT8JWtDReZgaJar6D
OytzAkaZ/dCacKwhrFTrWVnV9EjWg+SlZxi+FMF8tzzXIAXVL7xthR5GsRNL
RVKxwP0yZU2IvnpBPn4xUxlSODl/fNVCEEJCNwGtIA+WEhvNmq35MkEC216y
xu7Cbr/qamI96g8GZe3B+TIZsoSoJCPKf1xjw62RSh0OSuocVccV8+51uRBP
JIK2bssJdVua2pW/2njhKqJ/Wrr9LV3A+AkLxc7dBumG0fnNIQvBZL/iZLae
+KrBKMIFDZOQHNE+zlpKjgezcnybUHlgFaeCryHFNfF9uwUDtPsx5s+hct9N
vkpwmKaNIiWHKczZjIEZyV/VaEoAIodFxm3yFCiTI4HUD9PJB52948SSwr3c
e/ZBl2i5BjuxDhoYAF9sYPSDb4ccJRc+C0EBxm3YbNhxjpmVnXlmL43U/GXi
8Hv+iw2BB3rI5Ju+npwm4zZAOCjigrxRMx6ceDNvQyLbHoPNkqz7zxLJ2/Wl
zc1+2Tb7MowrAS8Y5zQtvajAGm8N8n7SzA+7Fv7zvxLxOYCXy6C6EuIngGbt
CToqsZpwEtcK7dLRXlmVi9NPoWG0xLP6HY11NObLNuR0mXkgJtv6gFCWP7jL
xzBInUannetVzSme00n4pBmz1TwcAJQONjpJfRBHww+jxcfjwVGq9AUYNMdi
SlmfwRYzOc6LUAV3+op242bZ9GPJ0tLV0nzPTQpp7Jp5UrSLXM8xu/aYPb56
2NVVEBsz4irbj1KRQ3CORmDqJLiZLOqc5hFrT06phdKYX9ZuM6DIxEBdFnKG
7hRX0ulAE/d89YpVItvCpbXHcCUYrwb/7nyDVVcTElcmAXV3q+iDRRsHwXyP
YKi85JaXri3ESbMKPGttbvfeCTQjJ+Vw1mtrhCCEDM5uqPFCAFBE/Lh4kdZK
43g3X3LHd7KUN7ptJClQWa8iuogO2d07KSeimBHgNJiMsu2Qf3HaZ4OJ9i3Y
Vx/pTmuwXbzl2mYRs75Aw32c4QX7ROebI6+J2UZNSd4pFq+aMb9/FhJVrkOt
7pua+wkk8/ui9h9i7pEbRx/+2LIXe7it1bEYTktHtgSN412mT0YjdWH9OJ6S
DcK5WMf0k4bcmnLRULS1G463wGangjUBUb+iUsOV5mICDVmRAaIvLSB7F+gx
HBIcgpbJ0LgOZIupOE8yxjiDMGmxb4M61OrTVaxGcfjaL/pWdtycqhWuiMsf
vINFgevvH4aZ+X/0K1BMEsH8B4Wz6KSjgQ9z6fnJ+twCWmQaO+pCZsr1kkdo
xqWIP3hdfiAJ82a9haDHLiMQneSTIysk/AbNSo9p+7PmkxrBy4VsV7I7oQEB
OWI/xArKuClGTjJ3Amja54PWkUDt75QGVoJm+4zAdT97Te8Uj6Leag1Ha5dL
6P18DmQHvpvlVPeCunaN1+vzVcIzHjkbZ60JGShvQo70m+XUEH/IvcgL2Y48
bquzZymni2yG7Uee0s4hrdsmX9eDYWAWBFqBfNNSb0w1ma3h2xV7dE0j0aU9
HJ0dNKj/PyzOhdb5ZDIcIcfXv3jrscN/7IETvmzzmvMcT/8fmGWoCstfd61l
B5D2LDBeKzH2Iv8IEpJODkP/7ysXdn+SWzl42V1x04D25lr/D3njzsWm0qkS
xUZsLtgxLwTS02afYZb8Ek4nKxn2amT2yZcoJ+Dr7ZKPxkVX8yY4RVWj9aDk
iC8Uqy8HA26TbCZSbo9zkiBIwotiJ7uQCXcgDYNhN8yJRPtGhMatBBWkxP9r
EOZOjePwRT9vRJN0VZtd5/ajA6KtAEK8xkEXvqtUyslrJrIwU7XTGBBOvjDy
AwlqCUv67GgMYQ6mEnM+vaICdRsXoh0DXkljoF2rKysBtK6WEhGDRE0wYp7R
3H5o7ny5qTpYG4J19WRDqXkn8ToLvmqCx26SOAAtb2TKyii0Wy4NTFvxWzwR
+VYkUloRT1CCPz88SyvkgNqFeQd3iowxZuulDBAMxdKnnqEs2M8JrpzYVBJ1
aV/wAAex4M9aU6iQkxZspiNWf2LDxs/7YZBA/WUXNzOH9Nahz/JqupgaoIeJ
H1nGJMpfokix0bxYk1MzAGCQnTeVttEpB8Zw7okfNrgHLAhoOjEMtPUVOdtL
p8sJh3LtCo3wJZY5vxEBOK9Bz0kimk9Vp2I9lWZ9V9HF8ykBymkfK14FKcUh
44YIIf7VQpzSwIDeJAQ8yj8AoceKDAp/KJmJJy2Wf3tgGOVj1bJB1zHJo37+
REi23rmY57iXVkCCffeN8kOLB1uLbTnGIoXlP4w1NuWiuFJXTN/3vFZbugQ2
ByUYWVbi9+CisW258Urbw4s/lGVmVGQ87pyUyEc2kLHao4UqhY+SqMXmdLvf
heGZXOj2j4OuLCAt8QVvbFJPZ6hzAJAny16K86Xg75NSYKKTY0z19FpYxTWp
tcUyWpFJos/Iu/eIqSx75qVyiCb5aK1SePD6dyqUACKekgX7EykEgRWtD6NS
I7EPgloFtHAUTmWApxF2s6q1zU4jKV4YowMKK3wX0hSAqo10gM5lFSgKvWUk
qAkTnvk2QvZhDG5C3Rz3f/vRX6ONedFOqWJIT4tw0xG/sBsnKO6lbTBcq6bM
awKengxpypn5XjI3wij2s9tjXWz8HbtEow0/lxl4KG/XaM9NcuSEfEGpK6ZI
XRJUbFv+LbibiQr1z3Pd9XUmRvW4EvGs4iTydQgbI5Dz148on44pp7cSoCv0
eZdWA3gXPASSTov8kjdKYf+Cpk3W6PplxQ4ThrxQ+yrkPV3YV6cgKefFyChZ
KWcRfuo1CHev0KqY2H4vFsa1nmSsf1YRAgVuHmUi5Ip7Oycz6nj+eiT/ISAJ
rsqyPn1d+Vl1G8ZbbpgOx8F9d6hjH+GEqPATea01h/7OrlvF2THy6jHsl9Ww
3r/KY7jbXEefpwx7uXatr4tyaelxW0lKeRiN01AnYQK5nU4Qu76C/mmniQvI
4BxSYOaK8/OmXew3xmrHV9Zw65AjAt0DMkr+i9xled5UiSj9WxmvdPATgLEN
t79FjCZZKnH/K9Xy1yQYUJ+tSI/4x+833v7LkCMxPzBvuw2FjGz34ySr/Oyo
uCwti/1lN4/okx/Wd9oeylVwLFYCm8EvQXy0+YqMkRdwyprp6YPl/mLEwIL0
kCnwqbOwSUrm1aJUHlTdDuqWoqSrr/+HBdtES2AVltK2ZBhKLy4CsGZVZmI7
+hUjKYmJAB53Klm46rb8SWYnajq/4mKcp9TDTQtTzXKfYv4S+42HCjjXVQ/M
xqQi5TAg493PTykHXHWTY06fbqJ151inLgF7R8MAmcILF5eDxn11Xc0Xu7J+
8H0/ItC16kYB0BNywj5FT+/i6QfsFff4lhk8Fs2KugoCgnyz4FG4AuO8z3Or
cOpA2Kv2GuFw1SPOVcIidp6VDw9OtSBfcAViEt5eh6sGAdl8PAeZEwxzVwwW
cgEA2/CIJ21Y+vfcZ4FXiBmJT5lzrATzTp2Q/xxJiNkjWg4uxDg/hhU7rfSW
uuCgE+Ea/GpPRkCkAZuii5W7OpH30oiishkXjhIbfFqKExJExsdJk7OHTkDa
jasGpkdhidCy30L2cmtYIynyGlAggNmMPYxn0VmrduIYUypIdEruDxmA60MG
yHD4gznK5BEviILz/YHi/acNu9HLVb1JpQk2JRjBLH8nD7pyQL2KQ2wCGlUs
d87UCYusRvzErJgnE3FuqjVNfUPilovoc8U1vbaJVb35RFFKTT9EzVutX/+T
PV2HYC23z4RYHn6aGBZaV0s5m5TXd7OcfIceEFPmT8xLceSLJ2qJKhoOjY9R
BF6jfO39QumpkeA0qDBdq2foT09gA5H4zhvou9YEgr9gLdwFvrO8h7Rx9TfD
AfZV8YvFIBoXSHXJqHPp5A31GQkAiXcSiVC8+mLWQzu+nekzJGQFZIAe3ABP
SEKHKeqNWfX6c+GDswYPzIngt20aogPplKp6TQrqKAbrB5DXj2BWq3CQZ9EJ
cMuFrPUZj7ROyXeeRPPIqWlp0elaSpD9cG/gnUVJmFHXy2mHKqTN/iquq5+5
F/Fdc1dZDq326HTjyFxOS47QlNvhNqc/1b4aExHdD/gOGr5Lhl12/URkfaWW
hPwbzCcotQ8MXCcjXeWLdcQ1JC9hha+ANcy6G1biNpTP5ok5WhAwgS/Ago2A
S2FY+FivG6iDSvP6rANxun6TSPK8ghtAH+L4wORaOnKO/R0StwvW1I1I3RzL
y6PZ4I5Sls6uN+NzRivLTIHKWrJJ66kRHsW6/+pMWLq4dzslkQzj2gLj4Upu
N0L3K/Y1m6xqDSDIn7NqzdJCPxCRdBjls1fMYCtdHUSiG9122IHrZDDVZpjW
N1PkfdrgWZ5E5NxmbgK35aMN4korayZUNGOOnGQU0rR4L+2YxJ4Mit5JmlcQ
cR4hEz3h3oiZCHNiK/kNvJvfg2JVmfdknhy/icguaIyFeWbDDEyBwUuExgU3
RXmaYS6C2kwLG2MyH57Zpq5aiSaDz3JWOTPLhOApmhEzsiLqqBUbut+flx8U
wnmisl7Ycp2vr2uWDQdLBkfXsS+8ynRSUV733yPyZL3nFGJtCT/cratq1OEW
ZUsdZ8NDWOLrR2zpLcyb27PBK0yCMzjHsn7+zOIY1iXXvNVlbYCPdGO+FlJm
JfPIDFoTpbXvIBvO/yNYfOdV8Ttt8LNBcg6ZZ2/sXXH9XgeTWwrTjes+m1eY
JDyp+HmdnvX5ZSW308Avn7wSKk/fCcQQWrpHp+psri6xtHqFI7jzRFlgOOra
GzwQgALmAHAVWksrECSgU6IGi9SCUYvIMEUTSQIYH/wZ9XZo8io/0MF/1nRV
xuK88r2fluGlPaCWCwgQuHTylCdtIcU2ewA4jf6OP8N1U5CKQf8FfimGRM8L
JmTrTO0vfPV2INoiVgD24O1U8vxh2aTvRzhp/F4it76KfnVsWwERPfTsrY9Z
CvKskiCuncGFev6tNkNFuGR7ecnvrF8suDo5IiYfphal3i2i30Rz/oBJ9x6f
vhVu1ZXXYhSeUAgVpkKIs1C6+JHsglPkC2hxzmvoZaaRZ1mUr9Mrqfk110To
prw8VN6bJuhSqZTxE7+WdSqE5csorhVdnFod7picQjU4UR0cf3LJA2laAAEX
6bHNjRgML0rYwdvu8terYoWQzATWhIHLK+7U0TxSMH83G22qhI12FtSIQBax
9kuAlmM0bAXUf4CUJxlfVcF+y8yIcR6n/bZn2mfyIzd6veIGEQjDtQtdMFV2
TTVRQQGIocPiStOHaUIBSc4/fFXUp/yQcmRjgsyBH+m1at6zeTNm1yAsaUbe
geWny+mb8zmg+vmW9VHgJZlU0dTrl7FQE1b4lqa69icqTcj5nxJLVxvN3Tv1
C2Ke+vLM8dzU8Dcy5IfWzwBOjqtPtW4mbEcV29RnDsD+PDFx59s9H85qAfr4
GlTBj+edRO7sr/7HgfLRirGAVHtg2wP2fd80Rst3/31w6Sk47gZeEZRZY2KZ
u8ElbkuTLpK+vV0GbcWS2FpyVNYhuDq0w0hwzAaoaONS+jM/mATbicdAFUSQ
2USHJtcRgc9Ut6JRLdZBpvfhJqvu36IuyW+sg3B66aJnYbqiGv5R3B70oVsX
tEkugvcFSBFtcCuhhnPTvPVXFAcdu/O+t06CBsQ3eIj099m7gXWGIfeLWKdT
Dj4bhsGv8D/tDmUH2Zgsdnngq97efWRHFMscEcTC+NMQ4T55bFFv234YkR7A
qSUUKVbutD7wcjGwcc449UZFA5tNIYhad861QxzdF6D6k48IF4OYx0VDT1j1
lczIS3O4UfKmZgF2BHi44d1FTkRkKQa0PAlD8QPP1AJUV4vMJbMtz0h+KIO6
HqtrfUDLJyOZxlZhydoovs0huW/DTTiS3MWoCHTozOlTVFxm9fux99qeeNpd
eDJBkZDDtOtaQjEVRWMmFDzr/azQhNwuKwsJ4CvQ+nLpin5cqEdnAWax4+cT
m/6beTAv2sU9nw3bbB2vfGys+22fcL3VquD8RCih9nO+KWk69MRtdr75FHx7
YgSsWLzZURJd7CjorKFE5GZFvSiS+0Kz6qQlBP3qnyTO8Go0VoSFurWdRYq4
ZMIj1tCgJdvtEScqrApNwYYpOuLzChGEH0et7x/2WmNbi5jGgk1P9MtRhjqO
L5kDqWaDuEs6mRTCqW6BzXFs4yZ7J+PR2lA04M3pk7Rcf97IjxyolU67yiSp
Fz5Uy1Xq+Wp5myqjCg9YoAkHQjELrWlnHcIsJEEs9lpgXg0+fKvIZMqbAjMk
jAplEhNgRDTdolvC67auqhAzMZEc36U0DH5yLYwquWyGn6TdxBB95uCO4NrO
+Bjv2Zy7HQvv2RfXY1n2VMDAg554X0iPd1g9bSv66jZe8OBZGWlS0k3qvsh/
3zuh88r3jKvcJsz0HgD4H3c09dUQRAoUYUg/MfbfiQ0XOLwfH+qZi4RDNOyO
EkXUzttF7KLiVWHJ5tQkgEt73yrpuGeTHiAbNS9BRrbj/3gezcdlHUWOQ7/y
FNJ9R/NbX/cpdDWZEDjJqhU0eb/sCPStKjyl7yAIUc8QA/xnZiuDBxKIkCIJ
8V88oOT/dIC8EkamgWJnWVvnb6inhnODsp5BkZ8+sFksSa+A5d6hEucmEmOh
dc0Zy75SzlkZzEwA6U1NlVm9RnHaFDyjqbWCH2pEO0EYU9BBnWTPTGDJOMrP
TAn3Jh/M7epwwrssVs77TNZVQT105GwAf4F7hKhM9Hp/yd3Y1o/HX6Mo8M7c
lNtfWBO0oGcTelyYjEqSQrOPDp/pj/feTEmYuh7jcpdZP9syjqfx5i23UX/L
G2gXyhi+7PJpD3T2y/fxdiSNI+FmtM4umtgiAJBDm91sh6J/ZPd4pQA6oBkf
WATF9B/e161z3aOJQnNPO229K/pLy8+ls0bEcE19c9rzL06w0j3wDYAFpIha
gmyLgukbv22pTMklDxthCSzcTk2AOJ+LxD2Ii/YZ/gsahUaM+bPb8FRhV+aR
VP6kugYLYB5zj6dGRQKOYCRk09H8+lGCjzrBKKVIr2uD4XYdZFrnIs+XBvxf
YYZknCRCjOUc86wiQu/y177ZQ5jP4ZVPWgvTQvyDANajv83Sj7AQYvNSdTjQ
oL7sMwRmGUC7pHVLjb4MrXRyV6qAP8XFH0BkkU1HzwzWVk9KPnRlm2D6Anzj
mR98zulGjoX68FZQg25fuyIuSJt1s790zJrCQavprDrlo3PwGcDNonxV4LuE
NOE/oTZeRsx8Ak+xEpxrQZnCylIQqFFX00QTYUwM4suS+3+5HQBqev9rgAHq
jMXFFwj1LEq8aIoX9w45Bsg2pMEyswld7Kk4IkLcB9ikFtnKUNXvgMH5nhLc
2Sxw031S8u++zjzU62wwN0aM6KO8i1rPQdTaHL5utnGPGAX4ASDkWqIy6kIx
CaMUfyzSguarxJwK8hCekU7ZA2mUz7AUaOWjypePxuwm1HoUNQFgMcYh8D2J
O3xl841GL8+afIMkB6vjZUbPIGZWHN3XO4nvLcsi6ULvJXL2OYVfdrOjk+pR
9Un/35qWay1CbtX8bwogUlRJcjWfKq58h9s5hZhBWC5wLYTNQjexoWATOTkm
7cVlxWZXezriYOw4C8Qy/btgmVrhJ1O0XXDXWivCnODkVKYuV5Vpdnd/dPI4
uroVIrHZLjjuxQBALYIp/HNs3+Dv00NXpGKh2I0OBhU2IhBCtuQ8Gk7GIdHk
yOK2/uqfGej9sWdbNK32eNOZ/gyoXr9stgiiz8ciYvyNi1tWyjHniCkJLTpH
4CwqlL5G8RW8y/aFimFYIr/9w3cERjmHNOPVYysAc/Q7Mow2FCRLHWPwHlo3
MYRmx0LwLBn9yhbZYyC8fWf47lCd/Zh1RUJVFqzQ0hdiiZt9IFKKsA/ff+hA
GZ2vmS9DMmK9z6xOlM8SviDq8GA6TnPBXbY7WlKG6yAb+QpwvjpvPEfbeppP
hOwRB9N5St99ocBWuOZg2672ocqsgWGKjs58R1y9CTISW59Zm6l8pZFKXytN
mmquBnNwmCdV4dC8NN8kSP50JcJ92Wx3O843ldDVnf8ZaL+4qi5k78eqgaHa
qcQ05D7LUey8t6CnDNU8eizJDvcP8EohVfN1DhRhJMfgUM8eTKdSuokC/K+U
B/EwdiUWCSGyjzT1HWFRG++Ye4MrdgLI7Sze7+ANp1+NVqQtXxIko/Mdcm2h
P5WRUJWpWkLWCWXiS1Dpoa9LvY99eaHC56FYp7XvUq/UW377rOaJ48eT8zvP
DzwJxm6GBtSaKFg0mcaLouVGF5ygLUXirbfgCs6WWSMW3YOICl1bHxTptESQ
NiuvzfAq6Fh1w7C8qlOQxVL/fLPRTOECjizNRTXT8abBtJRo47vG+31GkAv/
fjz1+TPbd6vx9eY+PkUVCMP7hXre9Olmj1oVbwElQhg8sFe6M3o71Nh6rk+r
P4wUyBFt3jXWDSbs2F9aVu2rtYk4tgyRe6owIVhClE3plq9DCoQ23plCvOsF
omT/p2swoXC0ZJiS0IHo1gnuCoMcI/u4v5RHw+AwAUR6THKYv6y0M55Brhjv
alvJRmHHDCXQ+iiylm8oZ5J0Tq7FZgTnjpdRIXU6P0snmcAI/W6S4fC50k1X
9t2485edjpk4Vp37LcGatWBXGTZ34CaAPQxd7cTOTmNfMs+0pi1g+/BgmVKN
uhQNtn2yHde62rmG850aOzRV/NtFLMYaLqN3XalZ/5ZfHNFX8Zq7+Hgg65Pa
rItgnzF98QiTzNJ1iVNfXAjgEEcy44QDRxXBbvaZXPFpF1xLJgApZn154peY
oK9Q30X8o6TOU3ohaGsrPVFH1iljOrS+2fADMxqs7tzvEfNfDmpiYzrUhJfS
HJcxStxR+bKCiJaqKi+kRY07MU6EB93T/HbzDlWaoRsPvKU559JyOLbOel84
XW/iZNOA/kSb7TbbMMpPx20JeSAeEUznA56E3HCyBZ57jwzUeuLqyGFnt2mm
j+Q9uYqtR1/a1lfBtjJJjJIepfXTLIW8p322z29egTI1Ixzi/3vHkgp8RRAP
WxSWcL1CuzQJs9Xhu/k8jRnujLO+wejpS6VOmRO8ibNv3NfygQUi0dwU3hPp
Osja5ssQZfvaall/SI8xdHocJRJ1BusO+MoHo0T6KE6dSphDC8nVFXRrOzo1
+U5sBT7o7PPaJkz4erE5ff3u7u2HMHxqtXbPusrdLrO6Dajw0vXWoGTBxEvp
W3CDfaXJQpp43+/v8y1pjqvS8uysd5VhLNfL1RQj5FW4G5h0qV27jzY7ZmPz
oX93UfF15N+MZZ2XCDBK9/6UtQDTvkJVvsTD+f37bd4vCJicUMmqNEyerCG1
qkK4PFms2+0hy9eoZaTyg+mZT6fxTI1c3IB1l+511TdTmRVkSsV6F7dbqr46
Z4S5x/sXnUiYjDwULMjeDZY/+NGWdPW/fH7OrCHtHVut1Jf7SlUxMP5f65C3
dOddOGSv/L2mGF0nk4FYso6qQDzbuqMYk1m9uno/vo1DDisH3ayzJgf2TvVI
nsq/QGepxMpHV4bZCF1uU4mYqBi3p5fkySgFjCp+/OI8oaxFwL2ECJ2Rhb84
Yc867FtX3iD6msmm1z8AKWIy/6vDhKSwde9H2jCYDgdGhgjMhQYmcFpou2mq
MzEJrk87YS2vWn8NrhZN+UFi3Gf35cBCrncCrmqpP8jFWB93Y57HHbcTL61X
sLL3rzSA3XWiLgthgTpK63K0giHFla61VmBw0+lBuPB5pIL184gvjEJHge38
W3SmRVALhovOW/HdfrCMdc4rA0GrDUL/HdoTE2Ic9TDmsMI/tpK4LH6F7qFc
SiHJVqR3bk9R8cdUoBjwC1cYuKH0kCmijQgbnyq1V0sebMqWzefDB/qxNhT5
fMsAel3RUtkMn25Qd2RFNSSVSbCSYavjfHLOTi62RhtXI4XzIHTka+cJMR4D
9NafLFfP5UPAxd/I2MfWexDbus5ZvYteYWoCugRlB+5NgEUN/LqIPyS9hirQ
jTwT7Huf+pxQbrzHgYV4tSUAvA8NAOkssSkVBg9+Eergt36V5McD+WF65sjd
RRJQbof33ag/dugusFcCqfRBHUOY9/XyMjf0gtmjtwTfDxUku0nRk3AnyNJ1
P795G6GPcTX6l0ygHDc0UkaacAjs9s7MG+ores3yf8OJ6R+wVT/p1U9lhADW
kpWs81aZJ8+pf3Q/SWqKi9h+bJJrtQzC+2CYHt2/s14Dj0Zn7tpwyioVtnGF
nVwlvQvtm6lqaYcQyc1LAP+IGe2B/LzmFsL7e5TWpxemiDMa1ajksBpfSkMv
fmNzyMNccOrWLanhSoTUGPjPvH7sR30455sgaybn9+2KXEn8pyjS4asLKLCP
ABooE0MmCs8YlyDU4aKxQeYTv4WcsnmMuxPtqvthZaagb9FiHFsc/vjOXEbc
hzbFSrpPsmSUQa4Rl8qy3r/ocLJfjmmnxmH6zpWPTzx4U9scaNRkokYa2EjC
veJ9xAIzpYdtyVo98HzQJuIQmTIk7m+CD+twHPytZaWrEpHbBNeYSIjhV2dT
R1jNSCWvDWBctsLOvb3sOSeOHd0WJ7tIIjYdIqDRREEog24GWY92C8cofJmA
uCSKofxuP7bMFkClLuilcEWQufJnHl+7es2bmPHliNi5uxEzLKPy0uNTZBCD
+C2Vs0CPu2JhtB6K5CPdaTG9BKdEirsU63xpRndg4/me1rKSYXqhPKSvRQjN
cDB0kj+ueaOmLR9zDL+wKlPQFCBul/GqcYXuHo2MuljqAgj/AAcOxULB6Nxu
1s3se1EHW5XYIJQRDGMqU9MX4CuDkW51gzwq2a2GawOmjBweBmEMLYj24o54
OXRBJ9O8Tt3u84dsoeolMvjxv2U8BCTRLCsxk+mMZ2BsfyuZwkFaHrVhXEvr
ZKUGC3wvSGe+phiNl2tjBG2n6boKY3LncTGrExkHUK0MpC4EfVTD6mFmnnu8
becG7MlQORnlxiyDaEQ5GE3aNMa+YVyy4qLPh5GXOA7BnGTnQWN+0mwraoGa
D+XbKrekzZPnCxrUUpFcJMMx5gAXrUZu/SeHIIwxJRQTWGzHQrA8dfPvxOYS
V/60M1uyjL5wl79MsTwt18qzKtVHMJPeHA1Q7/sJtk3IAun2h7v/LPzpITUd
xVeFAov/FfMQDMGUEwv3J2yW9B0TAUqq79NcWE2OQzWMce6ttbOZB2C234U4
N9NTprm4H2iUQUJOLmoQXTzcydxOVy3qKbD3PykaMORCKkkbSpRM4orCao40
x0LVjl6Oki2uFojbqjLCOq86xor0yMR7xccEqMDaMGvBCxu33UqJwn5RWPyY
IF3FHBbrs9YNsA/3XP2Jbwr9XasMFTKyPccGbCoswAHyDTk7ZswhbfkHTb5C
joW7Q+rxJDrOfBC6ObXViydfDSEJ/es9JJBwKRF6yyGZd8y1yUt9eQBEJ6sX
e7hXlRxPCEfcQkdfubLt264lkTeWO3r+P1flZqgJLVOII7ghD+pldyxn7OVF
w5zBZlVvFk4iQaq1sfg2cO6IdqEzJVddpMdQW7CyTYURsDeqLbRP1wZsR3dc
Q3i7JZeBk7Jbvtd1djc2/huo4R7zsotRdauUcZoTiMebysu4vEpbrBaEM6rh
Ji314aOoWnmCWe1gkD6K56iqvgoLnngm1CxhxQC9vjtHJckkuRs8RbQ5kMbn
4PqiP4BIIe6Kr7RWs5Q4R7zURAOBJyuHObEUmInN6prVAKBJSna6Ge4TSJsb
EaaVqv4efoaHYH2MsfDkXOzHXt8LEpBI5gm1bMAZDlgUvRcBI+yUpn+GNKfR
i5sxYgp91H/s2SlCtffeSkNSOwp5PfOjVEIcMLigQFfXfwbI6ntM7ISkZ9vq
rvycYGmhX3mnLPLZkvznReg/b0ysH6zjrtgwaplvc18tuAVxOXUGqupjL+Uo
OfUmzhBVmhKCio4UWUgh82gENklCUbyhPMGmBzzDC0aTU/12HoMENZnSSgU3
rGkV1GCkc80ZNjljnSQvYfLltHs1XkqMNwPSTcCC/yGnCWkFHrPerka3o+Up
kXFI7nXFwPRUTKucxyBOTNNXaIKfFgnoK7uk8GplF5RmODogVkRRkYnGGqgA
14azek+YTs0j1zajuxGmGf71I9WwJ17k/7gEHEZ/CMY5cHFfUskdkSSB/n7c
+2+4c1rDLs1AbQveOFpaNh1WtoPgA02Wl5ranNm79e7hzd3T4/Wk+k1spP0h
Vy5X/rq3IjMLMkNwfEJ0pKHyOtq7lJ2unyA9PImyeywyfQKCLNg47F0A7iuh
zfjUrSWe/IlJXx7Z5HI4ypQZyvWH0tFWhc6I1EhCkII0lEm5IvzmwHgVp2px
41E55tvmJRvzAdyVpPZ+4JA9SpIitxvjLeuVLcf9ylYpcmu71VDdUMCqWoKR
5H5fLMi9ecYnsQFTkkhPLkx19bbqzk4/myWuBjIrnK6WMgjP29vfX9YUse47
PB8pCSLaJesxZier6hUyaZw76jVAwURRrHMADMEfhTo1SIwS5phMfbSq/uhp
uv4GR4yESiVhnoz3rDUmR1SgFyZp0Xk7EyiRDXTHLqjZf+I6vBXiihWuallj
J13TTIi2KC1l25dKIicEqdgHqpuYU39sxUrKvvGPIWQDalp3CREF/9O8Fewi
zvZGmLxQ+Ria06ZLCQymhdJ1GNLwfO/LfYhdFggQtSwX5e6WdPygcZhL17SD
wl9zONPaesRp7tPIttbKvhnoVBU0ZWEi6FkK7i25MC19HfhFQ5eW9yG2wlKq
0tFEjQcNCfkjucEY78d5rkMUjbkYuvM4RKg2K7onCRvc1FTNF+c+6tu8dynV
iYze1uo9/oRGd85N08h7HOSR7Jau70Mn9Yf8UsH01/ygG5QQyqamxbV8hi78
B5rol56T65Qwxwg/pV/UGGgfehhvSlGVe/LOMKFkKy0GR7vyV/Vvry7JCNZY
FQhUWLCWHxeQYDva4a17IjnaWK5+EkiXsyTSRUUHWayObJFCiekPOYk0ncjk
90rQwO8RxTYXEhlo9qqtfYTYuUNJl9B5jGgD2l91DKzWVQc2/eYO6N73Wufd
eQ+KitAptGpa2tQU6TdW6ssdaX70wtzNECWVaUWIn+3JYGGztcDb4SOMV5xI
lMRcsEsgEr/G2u3xnHQgwoPYckS7OP/Xy4p5044bUh1ryQfhoj5UEiRgJmR+
rfwlDU9Sd/XVDBSt4KjvgbnWWTATGyBP+8dFSyNzMf+7Yqs/jnEmaHoQ6mgH
LvfG5CMk94Fp9X1nkS2g4qqBire8b9dn5V7odF/VHFFxguD6ELSKaN+5ZwNy
ATyEBGb6MinWDz9OpxAKvNPsLcokekKoABrDM++Ur0VPZo07NdA6AXeIOymg
VuAzIXeWlOWFyWTz7QRyQOC2hhBjgdKgSxupfT1xkb61Ai1gP1W7k0+zp9h+
3rFS/bXP7pV4CbEov7nGA4ECclOT4susDHMEvcEd4LYd0Ih09XdyJMI2sY6L
G3fINHEu4+zR6J2wUHpz1qPO0NVp7tVl+4zPu4nZGg7OyUGYG7fYsFFYEPGJ
PkhzrRhQz5MH0ImLcz//NnJ0Fn76tj5qMo95fZmPJ7d8Pl9TmOKvc3clCeBg
nbA//G+sFX+V/PsGUdBxrNZTCZJh7OqVRVxHLRuV5wr+tvN5QSD7U2Mx6uR8
pLn7XD8Le5v9fKRpxOz4ygbN5w8zqviwizSJ4kOm0MLg2UCISkQyoqI18YEB
4Oxn62I47XOQBOQPmri0YArNcCVmlU33UJo4a3zPVCboN0bBZtSQAf4mNnbi
Penkhca4avjr6Z5tGcI4gRC/KM+JEQ82ZNK9DgPnBj1769zXQkq3xY15JCsj
yRn8OXdAkSLWgJkp63/jfQCUYOcCETRAc97sPSfJcC9+hkWxgMAM3JxSgRtZ
n+2WL+Jouhos3bwJHMW1szlDa8ckTCfekZjH2+nZ9+gePCIrLALjyWao1wbf
lRfMS4g8KXlvzLBzSi7GV32KMsQO2Ev20DnACYz9ylHJ3kMx5HX9MVirWiLF
9gJBP6C1uP/uToMrDxJsUBbxhwebWKo2m3q0b+iUrMqQWlthvqUTAXM5F+Lc
g67X8/vOeLhI2xxMRNn13QfgzQpAU3fQKhKou3dRTfWvoYyW2FMTFviZ2J9u
L8W3/Uj0kht7+zlthbem9BtczAeaezs/KUmbSIbPk9zBN6RuGNKECV22R98x
2NVXTGa+ijIT6Ijurk7vgTZ+2ncq2rt3SKfQzNco2V5uw+Ir/BRKCCiN2+d5
htL4J6EuxzvYeteDhXrytX6eOqIyvtcCO2hA0yptDow5pqqoL5v6kFqbjlSh
RoncMYaG5Ad7dFzZDDfcqMyNxsgBGfAtZSKkzHZE49uQyevXNC4xzRQwO7UO
e0EbNiXKn0JwSXe4DCRsGk3nTyo6at7P74H8xFo8scdYGTz1Ma1jZXJooZq1
tYYh3nrBKVFgy+bteRWsO26nKXkKPdAPhrPt4INCW/R72vN3IVImwLS8PUsA
q6DZoe3AHWE9XLtcna8vYnJqSQNcnYfKLVkJPcs3Bpj6EAl7UYqk8dtxfi6a
z1+6tvYdeu9w4zKjd4Yxa+JdbVT8lfsS9TnsBCCuub41sSq+w2V6N9x1CqCo
QBSV4+3lxSKXGh/VhN/rqB1rCfwwx578C+H/2jHf7eEXK2Oq3QcQfF8oqT7F
JTfeD63oT2mHDMD/qMtcPyuMS/tJx1lIMtvXkRPc+IYEAXzeM2Cvs+9BmBNj
ThKQKTYiW+kMB3mt6hqzMSgzMSN/i1mcJtBdHPCbpAPqw4jq9cxxQSHAPaBi
8GODdQQaIiSF5coOhXpZ+zLRTR1bLFBvK8dbr/gkRBSy0EaTurzOO+e4wtUC
gpS6AtJ5/ZE3K0UjpZm/MfmZi4zmeLxgggXyd+nYLkLFfc1PsbsctRuwKXhs
FL+WQtIlXQyOqBTMhvSFBODlf8kfJfKEs1CsaV8mkHtPT/p1znwMZ/AkJpac
gwSudSy561M3VOLvp0+uWIXlJ+0I08lpKlpPIdCmQ/ZcEKYepg0NXiBdlBe9
69lPLBHZtmx1tJ8RqGqkkTjCJtlwa2ZTHB/SBQMudTpgfuMbqPPPX1Jdx+Ti
F2+noO5z6JG39SBTMDnJpyKAhz9TetvUTWJjiFFUOe8ZhF+uxuNzzeDL+1nz
+2VuhAeQsqn0U4RoDxeM2bEIfMfENgir5bZ1Y5XQcBatIS/DbZX6/e0SBYdJ
lh1l0+wYTr/9P3u/dD3BvH4T/LtVR+6DyyUR36u7JVKeqcnlHqS0B+n6NpoT
Cm2V2xP+1cWcmhPrRDXXb7Ip12oNKn9Wnp6qTvgaGKL5tuOPu0S9+jUai0K7
TI9J85xzwb9zwhUijym4KPU1xCCNlwDK8nNJkzmK1TExyDXpmfI/c0F7sDel
Q3UzwJCCdtpVWqeTnlCj9kMPA7bN4vMdJOqqz+5fLZ6zsZonIm4DFGMvR4v9
xD5fO3u2b/MehLL44E+ZyZCUk4m1qLpmnRDls8P5A8bCXrkUQuOSQ424waEs
1+I3locFgG0yePY9qQfkwsVHBydyt5zgBxMZmCuZB6/9HLfeWFzWRoa7AvK6
hOEvmIoA4DUu/zbxBl7nvJ3BSFJvPx4hXbH0KfZBH5m6QBnzO02WUMQl46T6
9JLCSPCvv4ZMDenk3IsiBvRPXbPXMvrfKj1hUnx6jNowm5IzAF57KXP4QHuZ
Bdoj0wIcAOoGL2Lw/4bAPZVRJFeeZk/WI3c8y0+KSMM3gxSnTkJn6NiFR3hK
qlcm2I6PGc9OeBmFTk0qSqQdjKo2m6auYDNMBgS5cCfJHaTBf49svIUDHYrF
e1YbJM4y4M0SfuK5iUqAOyF6NBkG09UfxMIWMTWCRvPhnkHYy3EIHmNsq1Zx
zesKcmI8IOp2f4+sLjQH6KI559fNMATL2N8dqd2lTkZaNBjfyBkVCmb4Z0NI
2ACG/iItsnfIo2GWdX9hQ3LgHi/fkIa47mLcuVVWOxkUIzPhPDEXX3gCGMdq
7W8GESVVEkMuPplqta1lROxHOl81j+ESxOlfw1wMFC3sZwVcxXYtmsHAT9+I
6E0Sy81Ljj9mIAT8QECajOFw//nxtIZpR6P2lnXCW7ILdANR/hQNS1zTgd40
yQTqVKLpdtgeCo+bO3Qtp7w0VcMjcLD8OVZ+MW3sRbk/sgK5cygeFt74XV4j
IpIKcnWyq7+wud4ENsYPYATngMHJWa62nVF+3FosxsWDazscYkMvi9/EnM26
dkLI55LTS/TaX73Nt4qpSm5fo/L6nGazsL1nBcl1xOO++y0ku8mXBE/tuxGg
jPHSLwyFyPYtKeNDwLMwWWzIBfKFjblCwgVVUgcky4U5DzuCH7A0tKqH4+M3
0/9h/BM06cLmgVou35W/V6PS8YEt4GoVaeGeG2VYVD57Vwv56XUnSseSxQ8k
2l0s/k99PEkzpaOc816gobaQ/ZLMWs8vaQAW4TAaJqUwETDo2jnPoc06EmWf
NXVBidK7yyqUgNfmCSIyUVgQtO+UqBdEQXoVvCFwWPm6ze8JHBjA0gR2/9H3
zODpmCTJLSx+cosfk9EOhVlXzVtdMoEn/NV8Cp6YqeC2/V6ibh0PjOxykoU/
QSMgZ83KTEUhFJmtlsotzT88rtkdXvB3Ej5F7WmHEsjWMqpYDaVTUIl1KL+B
ePZ+GmZgzQofhjd5hal10H2Moc4m/5B4nTKfntldh3g8HtWz0m38XO5zhdDw
rFN403S8E4guCGNOevBMjVX70AvLdfm+juD4O6ONmsUVqZhvrlN4QCynLc3t
nqQrX+d1KihHlWIkKxIvqanwM3CuL0Ll4K9ujmd9o/u961J+tdkVuvzmEAd7
rnt9UPVk87UfiVSc+VNQzB2VFoTjX8P5V9tFxbczgEdzPxwWzz810UTSSPfr
zjAwP5Ol3LbkN9mITl6INk0mI6ak4Y4k2oY7hTdLjGfJKdAmnIhXP7WYz7Vl
fXFmMB2B6r80l2VLZCtcTbq8vIEKeRNNg9ssKb95tMjI7bfiU9iu2yjYdPfO
z+LgrLflFVgqxPoN5Do2IkXHdbtd1xN8WIknEB7vW5tj6SJ51r4cFPbR8xIy
tgK+Sz56Ip8qe9KvUE1y6vzR1jLARy0kIR0hgzKbokVKYfi9JyFu0yuM3qor
UYlTUNO3OIornWQVlfvR74mlrV0YybmxBU7bd4sIv/uPStNyLOvasM2wTZkv
dxxVFmahDN9O1n8xqPt9YWbuZcO8WGSkcK/rQyRVBzlLPL8JT/arsKlDExBl
nefLyBGga7SetEPiHPiaKtazJKtlKdQEoVuDL1HH1VTdEYG8vD1etSHIhM9y
4GgZOWU+7TpyBiZsG8sWmnQko4VLcHE2L3pHc41h4kIQzMLeCfrR+1c30tNx
OGP/NUSHHNhCXZaZhVKuzvJ0gF0L+0nBpReoAStS8mxG997/lEfXuvyUn8fy
w7bncVT7t6AmN0uiIJZ94Pf00u56yT/sXFlwyPUgU1l0jnu7/dFBWpkjgXxB
L7JVrOjOD9YEIohOXz3m9/72ZQkp3TY1ZmD2CPyszJ6g47TVfBVxsDuXONVd
f0K/63PYaaJo6LixlO28HN0W/L7NDxnIMpKabEzqacbQ/jkZxLuzffM91Twr
ht0OsNSZEm8AZ/4/SI81Is+oLaj1Wntp34yJflfsKeYw872OwgrcnzbOiWSQ
q+pivimwEJIHCx1wIAHn55HvfSDxA196sE8Nxpnn0WVFECYOSuYWvK541xLa
lMsYeaBDifn+vUaPXl8Q1Q1uyBwkibEL5GFYb/XIyOsKRJp1IaXM66rWfD7q
nDTrWDGmUbS5cWgi7t/NO8Eyz6HxOBVspfUm62WCB5LiLONjUkvurtDCjrrS
mvXDdk2rRlmKiZA4Z4+7+35XEbamA3eFLneO1re38JWpqBrPv1V14HGkcbdc
GX4PLVeAH/4TdOm9w+8QkiwkLALS0FCeZDF9Ysn90HOA2bNm/J3VgeCH+N+O
onwZsLI59H0B3xz3/ictNOQQny5PiiNzGqGme96rfcqNJmlGQFs8CpLwh3fa
dN5/gxJWWQMdhn4vLmu6FetP3LcxEvVIiribb9ZgtWc2D0ENGyp00A1Lolu+
iOMCLffkv36gU93TQb/zYdOEYCQ4OHtMU7A9qUWxIE8CVhYVSM+eyW1F3TJC
R3/85WG2riG/czaBhVNZyRM9tBkw5b0/4mRe0Qa/xPeCIR3xucA7epMZxBoS
M/vJhB495gFybbE/HoTNq+WNkMhPioUABepAXUF42g18ZYePp44XpjRD9TJV
N05r8pnELMqJTBLd/ZDLOI4CD5BSLsrnmVZxJYF1CLMdIhVW39h9ZdOxhp8D
tIDWT0lZG9/dOQjCqKC7YZmE27yYUihfT9khHSvGgrfZckJ7F5UI7nl8ZT1Y
nWalefdolfYdClAcQK83cDXG4Tp5m2YQzrNHhncVdppGTkr9XlXCmX5jWHkd
Di0pS02oLmUKyVJYSifrwWDlLJx/grW5O3oAmFnVI3ZgZzpuJpLW4IW2mpvO
4WmPdjU25NbYk4aGKUL86ozFkdaQv3tcB5mdWRHGA9/QNlZnEu7qMJEXGVqt
itXSjvtXTB7VZ/1rAlzt/8XuhPzX3+Slh1qTYgkta3YQIEqu/Rh01lPN105J
lU1LYtUNKR1Fdl91/ukJhapjpwC5QN3Kv+bzC7TS7c53NLqRO5Okbd4EsLUm
saOe3Apme/wFvZLj//tXIXMXpT1mTx9dwmxwO/212t+lnSJ0OzP14LSYjyRl
CCqFP+Zf3ZSu1lePo4o3fTlw0qGq4UaFcNveknzXiOSfXa89X5kFToR+xTf+
8nCCWe/ghG1FhjAI7Co+I3w3d9owM5XT7Y62iB9zfyYKpzKw2T2+YkPTKD2B
bTqh2UhE/J21Z/2xjoAmS8l8I8s5RhddYlHr3W6ExMphuuXL+1jfiB5rXw1n
vSR7KL0N36dnDlWs6oYl4T0LACd+C+TlrFBpyJ6Fl3jpnXFR3A9ELWlQmwxR
NYorKcT5oEOqkVE+gUkMl5iUCL1vgFpPGT7rGoFk4JQBYcZS7rbUj6wSY6mQ
Jif1d4KyRHXMVIRz6xOz7cYhbYA9vwnSrGNrAiQKCvB6etQJexfYW62d1dE2
+K4txL4FZ4kP9iMQ7C2Nfd+CaxESLfD3AEJz4bveRkOWllIVPA+0hcbfa0k9
+pNNHh7qZE9K5muVGy0BLapHf8n9SBCoOmB4yds2VnjsDxRdJbOR5BNAlR5T
n05qPblm2nJcqZpS2zVXOWtU6NDtJWTk48iI7tprblY/2QciiNcBYvyXpqzM
f1zzTiTslapfvUvz5hyTTUdUZZ5KhQoN4s0ept3jdORZF34cSfzKLkXAKMZr
0Vc3W1VlcUF2YQ+TZ3Xn/rPc9OAUcutYvcRWIUR2amVQbtLEpHKO4ze1j9on
x9BQntmwXq+uU8sAKQRX2ZkeiSnRZCR+8ORHQWv9ZTb6NIGPVHPPcJ9z62DF
ZjMzMkY04VTuE84qhl5rvPMGwVyLWQueCZqCPGBZvrCKHabmCuZuvTBeoJC1
QH7u9JVOnK+u19p3vecfmh23ZGxQP9H3OLBAWjmGREaRx3NCOhTx2T2UJi4c
ShGc1QK9HTt8J2mLUABogsSFfzBUIF6wl6rywtlMMHThzMElTJDPJFwm4hcl
iXzaysF4rfevqCpXrYyIq1AjDtoI/L1xhaRtzsC78iCDl5cGV9vN07CyBre2
McVYb0heu7nhtA+3kuT1iVzO0WjJmX4f+W1bZIosSguLKBHLgDiJtdlmfITh
Fo4iX5d2tuJnqpYJFGDfvB5oE1li2ulWb6TcSpsxPjGb4ugAOGwxlNMqeG1y
10v2YvlJ5ycPnuUjOP0xdBccoR/0jo9nXDInKLKFwoL2pje+D7EIrjypo1v3
GpiKdr71C2G8nsc2WEGuwSFV9x8CNh8gM/jh6IfYUJfF7/2fzdf8G4CKYNbX
voC6RAfU6fiCvkB9pd4vtArqripMYHjQFdr0hF6dnhW4MFgnvU0tdv4m8QIY
U4IJ9WbMtZ9oVQptlN0/xrBWPzUSr8FxcukkXbULPVslWL4EavnPIzp9nOpv
SFlVJdBEAaqe9NGuuSaW8yo2NYcWhS5HRL/GopOMNoPOL1YQDAILsTuWK+Kg
C1OSig/qV52tyolynm0opAeDspRCU+QzlyBQTERfz1tTqkVqCE/L5eimzt2i
JWbh2JBIYngq9b7MFP+NSoPJJrcjIDTuWwZ7yv1OdaITe6ouF9sO9wV8HtDw
p+wjkhrlegK/XL1yIRDBaLhAEzjhu5kiLZQqiF8F7bB7HurXEuit4lJPBv5o
NqF6qu/4Vt7/dqGuLOqLBuDdKq2LApegJo8E03CxT8jkeSb62MSANzK+eka7
6vGUKcmfDa8ddYPeS/mirszXhkvu0+zU0PfCJ95rK2FTthtm22ME+qA8YDir
6wraTApsRfjnE1flIpYDXvUrANiRBdVjV2B06GlIZgG4qvJm9nex4yQPeyoW
tpFf2PktQIV8R1rD6vAwEnKFulOlZ4+qzuC1j36tdxYAkHiFY+8Em1Ur+Zmf
f1o1uYHj7MLR+cu8qlUDtldnOwO+qzzorURcU7bkcFaetw4GFo5U5Sldhd9Z
isccpynP06V0mu1Wu4JrIS7zZYXTfgnrrlxmHqj9+YcYt6XwqsVaed4xbbLA
aLDEMBdU84WUIXvQKIaAYDM9JJqRp8fQaaYUwfTZ3seNIWlgmOmVF1v/KRei
3hgwK1U4g6qRlt/mr32YOYoTRTWJN/qxoNKPtYO8Pqk9jk5OgEpHcYQQ+bsi
65jvMW0iCv1QdiYzPQ0l6s5XtgvGcJMTo0DT3wsTCfJDaL/78U0MIJAt40Fo
b7IB9n8CiNl/dTWc9dRKLfXi1l3ZvJSQSL9jhq4DtMgtBkLrcYtc3XI+3mOl
W2aJLkGAYV1PoCTNFhXfEBg0WJf91UCDoksnQHTI0BktT2xSk4cn8G9uGIly
JXSCZvLRPUiyWPcSkyR9DIWHYnMGBB6iwgvycHJaU8wT5H/wXvwwrcwsPoYi
V8N4DO434W2azjECBqNNeRGWYhNZNkqlWQ4yujV3hTZ+16lUxmjg8VXTpQOb
EqegWEJBCSPsLjAXT1fKg26M/9Ae0jWnbanBdWafFFJeajxzYrrLmchHWr3r
h0buTVy65Nci6rgcY/mf+9aIpGHjiWSBsMP1uKRHz6aGQmQgopnfoG3eOo5n
yG7sBENLRX6abbD/uuJKmte6ln/qzFqcQoOeZOhvv9G0VOVEAumpBZPNpz/s
TAK4q2DGLwbyD5/yxisAbTpvghWD3Q/5tW7Un7+RK2cs/MjNhLV/nkiz7WK7
jmv/tG1+mk3dY/6NroxFgom4Rdu8b2bwFKzyhmC8rKLb766yC6q1vIthLKKX
7NvftTZ4rejysijOUU0+T/UvKZUEr3PZCfcRDQCf7X1I6QLzNYIDGuXaCdIq
JOZdwfXIqixBxYw1neWv1VsyPWht8lKKi/glcPpAovfPzY4dHUVm/mK46iB9
02yUTGsZzgcn8mVWeImNvHqxBB/hoToGBvdS6pCsCblu+Q3vlh1jMFn+0Llr
SClsOG8efJfBhlvmLL8wb4WSUO10yISp20xBknRn2vZhf2N8eygZcLb9erQe
TaPUUayoBHgK/zapwTkfZMh8OePT1dJWNikvOp2P8h165IonAmnAJ5dUojb8
hK9nVX9xC+95wwPZHb19CBqrrjpjzHmV3oCXKccvOkbhIQRma58Ga3Lg6qOs
Pqcv/1EZRhNbyE5HlDKoVkPCORouT/mcIi/IrkUz7rZ2BC9HKXfg6xMMywwz
YqY6O+FJcuXyw8xvtStISILokMQcMIvk88AoLmH0ttggnOWRYm+4he4dzaxS
cmCdiVtm/JGgbcpRm9AEVhjjJwv+3frLOE6Ux7XytutprEd4B9vr1RDJ3AlO
kbxRN6Pvzv6NjdKncabXlsp2qMIor7SIg20IJPkDboJ6MOY3PEbgkelOaLgJ
1o54caxkn8sReLD6GEIBeaUFks6nwCjyQ+9FXFc9EFckILl0APUisUwUq6HZ
CY8HoifKYtYy+PEPXDljGZ0LlLawpcNHVy+CWFekxup/36cMsOqVgeTB4KL2
szodfYexU5AC+ZWolAE6P5yJMicS7BCEX3UWAlV2yD3PnXoylEIRO9WRKncX
KkigZNP0PMcho4+av3Dt6hX1zAGi5iHqKzTyxHE2hErpa+DuGtTWzfnekD3x
gujnAm4hkvk2ZryfoBDLUU/jEeNLey/5U2qbF8U6RJohPQSUf6tUnz5VRkYn
7Yw9qi0ln0qD2JLTKoibH0EjWlK0CdjQjb7VStfOFLOF0mNbjYtommJmdvm3
j274NdP6UyxvftmsjzHA9OZSxXVUQeh81tUznMZgnFhgJA/weQwuVS6iJzIU
1RtRAJv1E9pwvDk6FHQL2LFZNPIW/GvoKzEFRJhtdlT9q3epEBMGGjefIgif
u8Uje7+KV+ISiI/nbndpk36st6FbHOsYRhDJHS+JITjEcCEXxjfUnvHb77ES
oRIMEp7NaQD1vrFkFfLjLc6ZGm1UO3IFQGfZ+sDiEw93lUxlqBgzsNSYtPMA
KOK3MmF4FvvZfz4D4+/kPTA0ESNzTw9QHyHWK6GUSm6Plz2KsC0I+XKqwrMi
uHOScpHpVDEIPp93NbAMlHK10IxiLahL5nTw+tMG5QqV65V+2gQZc2mrSjzq
pVtg9nxIsChAjOO1j8Rl21N8ThPMgNHIsnr2UfSqBLL0B6n3cnxv5ODmrT0Z
DflTRzeTSTIPlQ22Q9y6pGyZchewYtKet5YYJuH373Ous7QY9lbq/Hi2D1k3
hUVwwgoVuR21u5ly9C+kclxVIRXuyOXeFrjCgqNI0PbjRvYQnskGEbw+kc3e
+U6DRBDSktcBBiGrI82O5MS1yCqIXmXBK5PmhzJ2p4Gf6039UdHbEM70n1N+
jxi6FyDjoUMts2ESF6tbWdO63dk7Vy/i9Z3pKvrMm2psczT+5LxSSPiGpyUv
QKNgg1wQ2QqprUzZ05mf0K+mp0GiA10XeCax/BUm86rnjUI356p3gRT6XJDe
f3Pg50HnPBAROIdhfUWjc9WppUXD3n95gvR2+0jPGNE3nc0qSVV3F4wH56fW
AMHn8SN1h0NVqAk9FbZB3z3B/kAROKFFAwtNT8Xlyv3/C+XZfReOR3zr/Pw7
hvzbiO588CUz4PIHGkHSAUe0rxHADXvE+2IUJCswCMzuLv3M7qYJDqyzPGp9
784HFUhkFPAsRAhH+Wk+GFsWTsWtuJk8GVjk52Y4pdstfLLVaK/qM1J4p1ts
/fZ+XPhiGhPmnRWmSMgmu1z9MUEFgUeGRiwrYfuSXNKD60NMU+XSxyLUZJ3E
AGDKDh+TTdCgdy1FHXOAo4hLfPZLs8qZk1RyXnxdj8MbM0qsuQRd5hjfepmN
46gm/yhfKgNK1Zu0XDv/drGv5IBwtQIfm/CA3GAkwjVws/dKnTBZmhKkxZ9n
rgUM8OVmwTSvDTQO7Rt86F63O/UbxEI0fKoC57al/NLEuCoVZru4czipQE1G
nVlBst2eTQGZcMRdvtZLPaOq/WRLKAHfkIaB1J47HV2JU2F/mj8Cl0JZsJ4w
RBS7FwbUP7NAxDAwujCezP2m/aKQGPfwiYitAgm/rDIj/CWsntvfg3De8YVi
Trzl3/P8IrlDNiFDKSui4NBvfSUiHrC5nGv9VYscBAmmr3hkZ675YQ0Qqqxw
Qt0h/w4XnDEwz4mzgqhPW6oVPyFcOgucYZNg83izPmUthyxqiev8TXlSc3Tt
QnteqXjh/P/WShD+1Q4RA4QhMQW0EKJsZtYGlIY7d/MUgQhCMWyMRlITGea/
vS4RzxWJ/TK7ZE6udG0fPoFZ3tb9b8+ZQa3+quvBXHGdpcMu3Tweu7EuUbAA
p9lGkmTcQ+CV67BEg0oOLVxh1a4W2/Y3kc/uTxHVDZE0I6aN1eIpZLPIuHKr
B58bJEO0s5LK3i26PMUQG20ih7Dxpubj6xgE6XU5/msteZIsyZhYzJe+GnCX
s8+MnEKuSeuuBSbZvPvC/3efS5vNzKdISKWVIXvrb/F3uyuGc7kPHvrvxygG
AUfvWmr3wBMK+VLCWzBafkLfGOmXVKpuTlfWmFTxsQTdihHTLkKWx2H4+85+
JR1XPqiLp+6XALwc5fEek0gaJ7ym116JCuRIuGizVCLqy4uka3T9LwsR0iXc
fmb1ZnNPZaitajf5Z/sX3eVsSY7zHb/p7gd3mGzttpd3mVLZRmkyczfdTKdD
ZEgkK08i3TyhgHutirVi0KCW4TgyOs7awNnJ+JPNzA8VGfQgkP2sxl4dJpfQ
YJWy/OMhbjWSKLaBsVSiizdD8Zez/KYpq7v6QtMfWaq8dECBphwV23gkABa8
27yl11PTQUhFygmpFFwq/FqDvVVpsROptzlCDuFDdVIjZJRR1ZRVZOclCfxn
RD39auPKFVs+2NEyCzZnkPUzC0dZViaQL52ZQi81Buf8NkVpNxNM2l7yULjI
q7bgwTGwa+RAMd0c7JHS3Tne4HxT+gybi6/g/giwHhV5dblQEb//Z55aa6Iv
bvNrCojE4gQiW7F5SywwdUEMAUWwEHnNrxv2TTvsPP6lp/540V8GTEFd1c0c
JAdmyS47e4Xc8MEOro1bROPed1Kr9GUeNhD9w5nxxbv69Q/5QR6y/zGbq998
Hj/cxKyYORb3m+28OsKmvmyF2F56XRX2boB+OlMUBaNj9N84D3Yry+p+v/js
m0ROJXhQKXgQBfKJwYko5U975b/GEMRTlTl0bBK/9RzsEsOe1YKpJ8IDbjky
nIHE1WmTIAECJ8FtySPQTaOMgl9Z5WE6D8K0xImLpxhwtNqVboElKFE6eLgP
2Fxx/HtIQkKGIHwyysYhMH/wyjacwLeir0AhkG7YFn2vdvstV2J7u8AF5Ubi
iizhkPHdO12MN61H6tz6Rkr9W7pBacX1U2PYggmC51w6pjGKI5ZYg8DBJmVW
43Cdxw9MWQaVk4pgBZJxo55cc8zAcFgdYrd5AkX0+4sPpcErW+CcysMXRafz
d6W8NJJCIolsRL9IwuMQmThRcUgm2KDhFZWDhCMTRb+uYsmaWBmGu85clEpo
Kiw1q7G91jcSvPLXt2PGpNmB0fd4x/zUTOa6+CIeWUOD+CsnjAk2ee99DD/E
Hbeaqe2CfPyuO2Jk5h7gcnC8DlV64cIsALjcq/PfZ0DisjD/gTFFaNVAKtWG
+uOD2DecXQC5WcCey2fGJoCGnU4qKOSB14xWIggEd331Tb27njPC4fC8cR9F
M9ehGZyNj8plrRuJQlcoc6OYUA3YnJ+vlipaTmRx/mRC74kDbMJqm8OxxRD3
mMqAVjwtEu/S49YZBvce8zl89t9kGUKPbGipy+d0gNXkL+0TOFsVpk0MHpjU
92JqCrGiumEKsov6BP9z9etzEtkZyJU7MWAv8PrD6PVoYaheFQMJfTS1Bp00
dLYbzG6JCbgHXIkrKVfdpxVhWieW+BganMNi05p3QYV7WZJmI9d1Ksd0evL+
0bHNw3YE8XGBgNAWMlMpa/N4uBlvONgVA9qP+xIjJdR2E3gexGlU2erF8Y/Y
EOmhUs1id3ivm8o4LENd7c0MZJyz2c1algTIoPe9go5JwCNgJflpdyFL3CEF
TVOiBaOcWDpT44sHlTo+ULh7XSRX//0FwSh5JH+ClpPlJz8+wbY7ORkQQWgp
84XP7WQSu0HqvtwdhNoj/cX/T5pzJokf9nG3sI8wgqjkHDZp4Srk/E0XpkE/
dyCLCMZbm7dO6rBNusIDwvAJzzrb2BQ1AFn947ZX/FEOX6j2XvPhz6jp7TDF
EG0Am8nsr6PMAk4podhg3Y7J/VL5fE/LhmXXDyKBsAe8yyLBJKnfBryc530s
+ABzRa+VcagDP2Pqcy5RvuAyZv8aF11Jj4IGVEFilDLMJAJUtpD5hFDMfhq5
7IlcpIKQWcOu/ZgRjJBxieJhHmSUoJYkHv1wixpw6ZQCO3a5JmuZkJrjO42h
zfiP3gZZsPr3E8KHIenjHfFnnsWF87ny6qkAxtC1fiDyPGqnZknKMS46EFnM
hOUPnA0BtHPdPCe8GEiAv5hLUM/Ey77nPQMzou9kxJOcXcJqSEpnwB42gW20
+JowodD2+VCAHdzxjuMmIOaad1l7w2u5OsK9apJ3V5Y/4Efbgw6RCLrUeafP
KbvQeWbpFWqWy3ao0ek0VmjWbrdWZmkMkRkLuISaUENBoIiGDpHsVqLC5G3Y
nap6/EB8AysVz4rZUzIrsQK0lmnT+D0/T4YK8TkfcwiV6jgW0HVaLEXrFYw7
rHuDnJLZ7GktGPgTrXrqee6xFv3AZUFTygtTDC+QdsKblLk8y4+ChkqRyuYp
sONIWYv6UuZ29Gi2gjhUT2NW/cAGcWlR6HoceQtFFjMp0cQdxpIt8AdaecGY
D826gAsibGxZ64yXAcpY8Z1OrjMBKvkDMeGE057tHLtjpPAK0aEn6GYCO1Rw
b8GPo1AYsA/MPMwM5XgaD/98G5/nCl1O0X3zHaakett5sWnV3a+ufvWAX/ag
nNJuEh4t9wxpTNmCBUvZmaSUaGw5BMhdpnnt8YRddzq2HTtBf5gULswcazm9
vNYyrT46yGV0VIGhBKB0aoJ0gl4B7hnCKwf230kqx/Op49ckh2WhvCpcljSU
Rlaj9OlFivKddPgK7fyFXRU/hqaXqkMg8jcoyYTgHmZskyYqNrPNFAZ5fFB0
mXmsy9V53SWp/WZuOe6fvhfwlEzGiiLgF4z1xU+lvuz2bC4Yv4xfLRY2Qtk+
OMocly+wDZX2lpf4wckUZa9IRA4vA/aVCA2clbbSWTMMnLQy+63QUST6Eu0F
7uV1oFdbvMFjIhl3PFSu4yzBL1C9VvE7rsUc83VXsYfAtef+yJag6TtIhodY
o4bMSHoNBYcbh3yUFG7iLj+x61YttTVm2LyxOaQBrfwFX7YOwbzlJ3TYJeDp
EQozuvPPbQWLI/vvcx0Cv9BBrARIk6IMuZXiANT6Y0IoliqmAWSvtDoFB1Vb
f9D12CTR41QJejq5OKN8/e+SFOvf7JQQIUyQHHZYJkCscoN5K/DfsTDRiAp2
GxTN4UtalU2pBS+JgaK6nGSzFA3Wgq6rbaRHj9T17lqhv038TPOkoQLpEBDr
32Z3QBOZgI2+cjFMkuYiQe5O6DVBrpmTKTPgWsb/ai6L8K/daWZRiOZabUzI
lwiBDMrtZvcaBEwFDU11mLQ5uGzorRX8NYxY+BlUBuJZouL8K2fAj0ST56pd
MgPCWGKRciRqlq+gOhcBDpOBqZOZvNiYyLaRtIMKMGnyUq2nY9W7KYlivMD4
CtB1xKxJISN9lAM5lV/aygTSaCeTpo/3FphUiUFwWFjpnkfeXQOlG4KX7mOc
VfqLIqIBWuVEiTrwK8ChY4WTOQTZZiqXRtv+6dYmq4/1gYz58OREA4qjN0fR
1eHKI9UcDXQWXLoQCAocvnKjTcVIdOJ+tj5hb+W7uwOd0eVDPtxe6SPi5XIY
K/3aQWFd9TygLyUJEhM3AF5Kf7MONgVW3MytQCe9GobUQndQ+mAAj5aJN/j1
eqqxG93T8mI63dVgd+c0VZkyF/Ea8Qh6E/THcpJZGzGlDcFMZGi0gQeAGMqy
hiYE2WpiNK1vztbardWolzV+xHZ1tKfyv3hFeMEpRV9inOmJVelDFLjjCYVt
dC8EakbvdzMSNBUU4i2dnVIN1HV2QsX4PvpCxC/xfPerMqZEyGhK6X9G4+Gj
chffhtJmjhLW+tU15XEH6aAwrdxH9Gx/GM0jUaJyRmOfmtNsRVowfjUjvTYu
IBmH/2HJDWgn+WJBV26vVWnZmFQoRjTNle7gx6ywSZUYYCc1GGRmowQGGvfP
R2k/0Gpp24OGBI+AQf12I71XgqPBMulWzkOzofB2g8EP+SIUtuwFiSuXis7C
a5cyAgrNtvfBedzfQLCpNkOsMy7pWI/cPobMNRPdBe333kMVB1OHXSynWwdf
6Y51as3K3qYaE9WNgNuJLvAqXLZw7qOFzu0B7WKyV7O2p4JlaKv6Jm3PhnO5
FEtICG+GfFpgvFiokWLBAmcaXK+A94Y4lWmUUHVDbxk7rEMgzVkjtwaStGKF
/Hh8vflNdGsjWRSCug/3BGTeDYfcFRFjzDJsKtC8uFEgS+7qPWUTJClHuEZY
J4k49gXqB7fmoXHG9KY6hkSBJ+AWV8+c8QXriNFEP5Pr0NTezQGRj7wm9UIh
5N+QDoF5TQe9m11MlvxcZDFuHZsBJEWsb8Z2MfUabC1kZLD/hlVkCww1HP+t
a7fHHwMFJgX2UuN/VMh1NrBoMCR8WgDr6VEzGSDmi+JuzeCZHtHEgyLit5ET
oWRCYcVN2mvO2HCxQhfDqSbmKtEuhu1tlwAcTmu0X50KGuq7djqr41ECCfVm
ujQyAFmkGq4Hpor5V8JR8fvqDRPrFkUvas0m+3Pgj8CRuZZwh6fu7wxYRski
s7MQ1QAtYTExXNyzDB5166dOtmlZ3ByNDVHIym1mUcpkXMQyLRYxmlQ8HPMt
sa2z096FGBuQ3tzQy8hf8v0K9En9KrALctsrQA11NO38c2NWzf369rkd4O4K
JKzdP1SKp6pQxnU5M2VlWLpv8rDQrQQcxM2n0awxx8onp6LDW3Uk8PGyPf2B
a07JSOURPHkGNt2zOBa3DT++K91d+fSdQ8rlQdrXi82k1g0yxSU8eXfgqxzt
DFVa8sTGc9oWInNeYhDbG/PIE2t30i5N6zjdXp66UXy49Bj9YI2NzXk9OMVm
s5BIiU8two3Cy5s2w21u7erQx/unk5kKEDbecOUnRC/k8GBAEM9+EHD8einM
zLeA70YeyZ0X/4zmwmVmpf19+0Ya3aU/zC4nFIX5NGBVfDc+xHLPwty95/4e
K1lHA1jt8BMBChTSZdBEtrPyGm6b1M7Si2WosAKvIGQqKmh0t6GBbw0d3rDT
bC4XC5cHH5XWABSNE4Jy+Yuln0dQwMBJzY0oW961kLzZU+oBzn96NNyEI7gc
UC39iRDj/at6jqS4F19jY/KqCaT6YZlb3UmSY3aEv7ERdAS0c0+/2fdLy2m8
GVSFnZL+mRNPCS+aTemo/MxNw0VQ8sU/wG1aXHRlYkzexD/lDb9LlI0CpHYR
EGJnkwLbDpkcN38f7v8lNIvfHOUh7DMtUUBCK6UPjtSURcSlPSpivc0yxzjt
XuAIOyW15BWjpDlOPgzUsY2xXnn4M9nrYuXdCOYqJp2CTZ5rXWUIx7MlE/lc
H9Q2kzRvN+59GOum6aOSdE6dGEfFGiHd4ggMZOCQpbKHkuvmDQ8BfWR5JURS
dXjrEIUZaOXKgksO7t/36DpMieqMqek/LkRGg5ShT2EfeH2QU5xdtEq6Yt8i
/68/8x5cF/Pjz6El/2rrYVEnRH2dXMPTSpjXnZjS0ufvYsfgzLQzaSA4d+0L
3dj9aiUDndqqUDfUEkpHlyAT3Xg85Y6g2sTu9aiY8NNLMwEId7O8Zy/KBO+B
dNDHoo+GnuTAfOAZB3wfzaGwo2HCyFtDqH8qmp7UJMCKZsxO4tQSAdp7Jf2Z
IDtZB7QBJWjlJ1PB2IQ24n56/Je946iShlrxhUdz2u0a84meIgHv5dhYrH1a
gq2W8GkL9LP7acKGwpPfxXxzXnEQ9pMGiPTa0k5+GyRRdN6AhT5sZ3b6Pfa+
qMdaYTvrSH+xzaZN0aYkaftJnU6V8y8hUdx+bK53QyXVrVTYaqXwJR5Cljas
NrZawjxdAEL0Qxg3tojUMmca2WyfYKyED5e5uuN1zK1GgCVkpAQLiHBBoydy
pmOYgR/s6TCL3w6knHCXbu0qd0ZW55anXURdrBGOrbIBE8OWW6nh40lDpI2Q
BDG+yoLS+UGa+4u1tk0yNnDFTCj84l//8PkScQHgNIWujjcG3wGnV0OEAHqG
ptH5W6Gio5L6vYC8l1YaE/sWasnfKXlpeeYKrNAkhkMAW+uVwwFKe/Y0DG9E
oodmtlq2H+9tsrfL+ZOfOz/N2F7V2u7QOeTNtZ+aDO+d7C3080sJg1mktOnj
cbt+IDiIeWTzh6306YI/iOxf06VkSJOjOuj6SKMwoRp//cslbqxosg/7Mhj1
V58p8C7rbkNIcemNV12lyq1eUrHSffFiVMMZxGVIhu/V7RzJneiojuwObqNj
Xl2u2YznzdfPcLJ7qSC4cev6Z95xx7FcYJ/hiVN/zgbvYAPZY12VVi/6b/H/
qndCcCWTxh6jdmGgITIfHDguN6ISs0vmoiVgSTh1ZqjQhtLf+N4ZQDCs4BwT
uyXQvSfQNT63cv+HoAgZh7bsd6y3knW60TgHbGhB7mOxmbvS6cBO1GQB96a1
uTomJEu5yLcCAXue/UuTuSQ3HU27dwV4GHJBg/hpLtU9clr4pyfvN/CL/JJK
kNE1sOexkmM7GUS69o6p7M1ZadM8LuSPZh+1SAwYpevunUiREQysxAFFZVqt
VhfvHTiWiecE7TXIigCbSaXQxcVrdFj5HYFM4z1/2usLolyvE9of2DcvNpf8
JwHwNPGeLtMI9ZLKAIl2zfjtkTBV9ouDjJ2+Hm4/wgYzV+vUiRGuEgHrF6zN
10bcha80OS/IQQjJmLAtR5RgXgLzyDOtH6yQbmZzCcuCei9zGkRb38/yZLQK
pl65Iyl9oPNDDhovTI5UsQzXb+OFoqEIPBNultlRHqig7GP7U8tEeZw2wpnW
ia5bqR2rU1SoDQe1UIx2EOag/B+wE/2Rh6BCDm3GJL+UHYKk5LtoDnD3vHwx
AfxlifhxUjH3X0lJ4ruQSy+4ux/0AA2W9E1LCf17jtoCz8K7rKQGkK+YsB12
WR+6AkJGtwm4dWQ+akIyO5AvwNsaCQxVR8XuTtPNAtSEUHm+64aGGS/Tnwdn
oYc2ca7NWpvVTdmVnZiEkhmmA0Zw5/6OXyC1eIuqGOgCk7cdXkVYC5pZf9t7
UPsf74u2cKFowKPc6hTfE6fmR0rjgN4RaqfipgH8h/649bbEkKBjUoClCixc
UZr9AY+uj/KokxRpe1MJUrtTFYsR8UTSF/NzUsSE4IKDkDE3tCvyChDKbgaG
uE+uWqZaAtHxkNRG7HqT8TSURPN6pQpjZxfPtdWP98c+dDklIb2iDQJnpoz/
XWjfLBZUsWZPHauA8MK9Tum1xgTubbTsJpyFSAXq1rsD4oueIjuQ/GTkJrlI
rCrhkr9ZKz6KOwH9j/r1WYUrxuSUNkh6P9719kIT82ECxAax9enYOtEhAWZp
dUSUZetSfditQgD0AhnnMfXFo6ADmM07YvsrT2B4fksM/gkkzYetSsYsrGFf
3Cq9cs1fqtG6jujyaeOzl1GJfhZSu/tBmHnxnyAR7Xp0o4gR3dzP3Si0mRa5
tEMDelxHMJcOBo3icfPphy4XW94FPI/P72rkM6NI37MLj8ptFQVcNbqiRWW6
z4seZJbnP2AI6/++3EJIwE+tx97R8ln2VQDNcr/6Vk0Zm2VuG7mQboHierM2
ALgef3cMLsB1tyYvOiryAuYIjoo4d6T765qCxFt1TYTxiQk3HiLBlHCiS3sk
/cK7ySt75eSJ+gPab64V2WHW1yOf20+Ka3Ii023rfxPUN3urZ/ZwvkMgbBrJ
VFpQ3spifs34zztrWlmCREkvsVSxGOnkVUpvl0LKLjq2bwOX7g0G1YgxhWRp
KWoZ+Cc2eD8Ha9LjMUbTX8iCwaDPwEmO6K1mNgQIHqsQK1NZZgGRejCaSPiy
Msr/dUeLE7AvkZ8mqDMWNGSxPsBNLBUeVe2Tt6lpIiNQhH4xyz4wG4hK5HTo
5I4fqXVxkya7GV1eRQXXq4fq78MgvtUkIy7USIYRDvErSEozf7RmIz4CWxoC
bjBWmFeP2RhvPuFR5o49WWAJ0e6/DXfJwZ19q8gZpeK2qckMFCRDeOIuqNkH
t5KAroTLRW0gPB/9bHeJqTY/SIskVGQs6Bd5iVTYNJKtF8MQkO2TCm9ER1PT
ZxN0v5f4zhWqOIK3CE05Wq64a5xbVrg1ZqETjxQ5/GyFjLPFyLmcyBcwNYe7
UjRuqZl9TEpoTINhHreB8vAnqGXbo3IxjwYT1ShLFYqhR3L6pO5t2Tf3IhZJ
slxf6KEClgKs4BP5MC7kzK5M7EPvliRHwdktMCbSd2WaqfuvFBDEgk0aHwO2
ZMSVZ+WBtfQtVuGDGhl2QTfrbXS5lu1hOgIVKyLMRRIjizqx+246fZr6dtX1
/mXGndoH8v7gJljxal1Bnr1d3BTgz/L2wr11CZBb6i7K04srGGP+v8Ltig8/
nInW0amQPLvLYSXAkkgN5DMge/kvaiPfe22iB7cGn4nqpyu/rz2M6wtU3M9x
8XJH8X3wEas5SA7Dhb9hwiGYfPlerX+x35sCfTKB8AAbj6USDp86qe2jm/sa
Bs9uM+UDPjIDfv9asTt3fi6aO/eRFBsbcTRfTt0qyjlPiuQAI9HL2CpTxb4w
mLczbNyELS3jNf6jSf2CeRtRjrO+jFDSNe/AVM4n/nsVmh/xfs6T/ayhf8Fr
xD1Z0x25cdZDUFz6DqHfQdEoDa2v0k2IClwhBNg1MFXT8gF9blzl1eSNzegl
f85fnIOeasuQtZ852LPhCAT6NdAZn2rR2Z28NRo09pXOwPaJL1gPro9ClV5D
2PdG0HMiM4HfRlBXTQSszw+IeLc2LcsDSkezhdC8i5HscT9Ae9qMeQQJoR+i
USFmxiWC7XY+GCLiupeugzPB3U0Vci9JoPqb63ucHy51fwuORGTqQWvIC6h1
Mzvm93obS7XRFAjiSHdIGWqmliqz1+cASX8JBaO1mtNAW5N5ggFZwCY9MAmm
AnrdIS1A4O3Qcts/sYAWeJdQnUIvPSWy3Hc0CAsMJeGoqjl2GRFxOQOVc39L
Sl7gNISnbbaKBg4iK1z6GoD8nnOFh8FFgdQzth2R+SIjgAk7WawRuAuk+uTO
LAYJJ7Fpt1gcG30xGgafezdYZXAsywk6N7u6R29NvDmSGoVyhJbMwN5jH9hH
uo/c2H9QIQ71TmZQLiDao7bjDpApXS7PsBJoE9688lkkY/1LnOx6AbtVUK5L
xQ/bJGSbIHb76cDOc9WnAIlwZtzzvRAYqT/EO44ceR54nTdWnffmnADyfEfc
xq4HsqaHI5CWDzXvTTJrvx/PRkFMblLvOloMD41PvC4BUH5CkQJHaQrYAoWh
buFdDatYdirv4rtCiar4cKRYeqMyF80DUDjgY8JeSDMeUEv2ESjMpEuPmr7v
hPkCkY125N9HU2Cfbwb9a46KIFgUVuAnIorkXec+mGyi1yzJArkXUyVcCksg
0LGwbf8lPtAIhWdxNAk0Pe+cwSBxB/ZjwO8iJoApDBbKQyYw9PXIlkTOrKW0
Kg/teEKkdjGleVWPqMRWVKPlehH05cu9l3pXDddolrb/Gl9xcyHZVrOEXuwy
p0J8iFkMowLDQXmGHAEDDi+T6uAVx0pKRHprKtDn0iKSw+IDlMbOeiuUJ4kk
E0JaNFmSOky0Hrd1H21C6ONbJGzpXcHh5F546pQV1EjdVfD1vtR0yDaV1Xqx
fgUwRM1iPy45YqZY7LzGapwufnZgd68Zc+yaZ5FhvplvwdmUKIoYc/m8tfFP
lmK6RNlVsuF216cyEV1XA3xuZqtlFUG+8BevqxuTmHnjHZgN+6aRVtExzckY
VbrBH6XDztycj1MjDzha+AWjpY8+5zNE7EhXVXZx1Fktbqz8v1SUMWpi6CT7
4M0sSyhIDt0C/TvAU2/TkZGeLqQ32tfSjuOLsbO3+j6jWHiAM/DKanaqQrPt
Dg8oroPB8zIXoBxzpsfu11UmArQcYWAMLXy7dXYCcBqoCXnIYI+paLrBiyUs
0MJqVmlZP+5p6Mrku/ZkbwQPmSUOAarvDPWj3dqClXfBwNqSqlP9+boXc2Rt
GEStCn0SUtT+ZtSb9af20zrPh+zyhI7loqz0HmS8oD62XAyEB/upOPJ1Qtgs
oplquiOMX54o2RmFjMB2ULPF2utuAU6O6gUnrL69J6b34LdoAOygrGl/cjR8
4YWdTGOssjs3/+EgW7bHwk1w5GhS5hIBv6rmDZp1p1bQXdKIDt+zIox1Vct6
qoDwK6d/1pZ0Y9q/rVFyCf2hjZ+X3FT21B1sMJPvNB610PpmdzF3IUvTkqhY
sDwFkfFv4K4e/uo0QfXhZG2h3It8nwNc2dVo6Ykde34zzsN5gULIR2XJc+Lc
32hocqx5/A2rKNq6gJE9gfhcMnV+5bFzdPVQ6Gj3t/uICSwOTB4Z7GOsyVRa
65RLcb1geEtT8qk2haGYMxhKgHmFuGhYLhSx1o5KvbovbQAZySp2VOUaV+hZ
mQPRzSqaGvSbWNpCmbgoKf2UGh/mB6InurP4Yu4V6qFmp3fuojeM+KIyTbaV
StM5QD19oZBzjVAYKybhGtmQcZrJpRRPvo9Q6CqAsnZikHxa1ScMRo+PhWNF
SDlfsYYHisP0N6WXP7/RAONwwjXA1G3AKFpS+ELrtHnmHy6m6t8qAXh6YZgy
Cq+vlgJTI4zTWOcCayAZG0sTocVwGp3VX+/UIFgw1JrJOc6jsBIYD+/nYP+c
xdMBc0XT1vhqRXxF3L2eGNfR35Hobwhcn7g8ChjOqDUbDBmevosLNl8++Zae
1uDQbBosHQ1uwso4wPM85Ev+rWPFaCOr9/mMuCfSLqgGaH/7YNgo1eL9GehG
/u2W3haOqN2jK2ZFcWdO3Wd+O9asTCkSFZrmpwUbMtMMe3ekQrnSYf+J0b7+
AyEVpW0JKiOQfGifHDpxWooFeIetYUrdunFo1/4xr9WNoYXsQvjMgXtVRzsL
B1dIiHE4Vdse67ZOC8fTVSzwGzK5C8qDiduqbmn+yB5JqTEZB37yq1mYqhS6
QW9whytI8dmVvTjK6GCnhjHCi0DW9Ao+Ij0UBrY6trq+Q+A3QA6gj+u889FN
HevwfLs1a1IwcQX3XLfjKY36MurmcOR6BnYhs8jsIgpUCz5Smgt5Kw04pTLh
/MDBmIE7L9guBIxu3TKHew4Op5hClMUaFcVxCiVVo7LCnTnLosQFu7gs6xdN
GlDnjhLH9Rww1mf0wRo0Vm/jAKhW+w9HCaqZyv2wZQ5YBPPTMgt4pfbZsPc7
erdZivdi9Yz8lw4/YYOsCYKhMhfsvAgxvmHfn9CeT0/otPJgRsh3yuFGh4E9
GoENzYJqzGoHUwvJs2zITqnAE2tuytDad+O6eKptiMLzpF2MMnuLI2tB04qf
IRmftM9VKGv4Yy2F6NPbgCDxzodEcqmb39bm39BFpxvuWTadGIlPrxXipAVO
OVUyrSk/pvEAERfdE8+49DrkRDhuqK/Pqtt/xzZ/b7YbOc5gJG+ANHUZpjYz
qKJmi/JXRYRdAyhvm657207kCY+20ngPf6gFl13lopWWHkNn68K2s/bH8Kc0
HF+jh1wHf5T0wG9LQaDNfxooelS/Nb0tRvUD6tJDjOwgfpmBeNu4daDDeTaP
Db4Ab4l6fpWegMF7wtqUykPpEvc/s60p5qb7ofIMzwHD+7axvPPwJDHTqrSg
krc75vdIIBYtmNII9karWM3aoITkGspg0OjCY8E8HONhNzEyZF2EY9WhioD2
AudvzXYZwoh3lWTo1yAdrO+1tqW2aOHosJ5TJxxUfH043kNDu7UXtzJmBWNz
gO5+OAlQDfIFS6DSMwPd/D9SfDT0abUwEtHDfc4rddUNpnZcBECtyGIrqc25
fcLCY2FxXqakFxzqag7h41kHXQEv503QUS6MjaE2DFB/JfGCtsePdmAlmUCD
YQagEtO7a+N8TLf35RddN7BrselxlJ/W5LltWHw0+TPUO1QC9/Awh7eHRFFn
CLwYksrnYEwQCM1W4/HetF2HicvkJWq7IAAkuxpDXgyGe5/SDeVTEmgm+fFC
KOCPercmN1iSrceSQyUUnrCusL9SPtr3KNOgsk6SaA1C5VGDpEuW/bI7bV/7
x0shzhNkh+P9MaWKHXbA1casXxXSAIuRHU8bB3pYU8NBodEYXGtFW3gVFNVH
fVelZAKOVQbohYS6fgNxY4Vul1e+Paizy8hFTCFjiM2ojT1z2YPyT6ULXTsf
wdpohz9EmAqJOVG6qq7ZEh9Os5tdk5sldeTXmrMmrdM688vP70YK/8f/1a9H
eBPlizaMsE4CMGosFNA6iC0h9YXzhlEPNqRJyo7P4+QJZgYm2GJx571Y1xZG
AYtw3kDJ7PK52bSNSinKKReIh+A6ntKZDgUTHD7YZupaCh3UYA5jd8G5jX/p
8ISM4klxImZl2FScyIW/RFUN4msEQVEqJ0Psj1338iE+cmssrYuo8i2VyMDx
oCtUfh2JCCP2xbc2zuJaPOHsUZ6ixN7XVLi9lwAiC2USBHdF0YhRhZY7YsD0
xpmOesrkLoorffuzApFaR+LrfCCLUlb39S/0wl1qa5xS83UtWhD6YgaKEQG/
nSB5SEEYaLC65fPnQYgmzViN7uD4fwiiHQaqVbcGr6pvme+Kh8sIvQSyyZtW
q/9slDdzhvm5QU7gVmQO+CAusV2g7XoXBx8YPc+44gObEwHqtVgjEcbmDM3N
oIgJnKVZ34MBwkM8TWDJP/PK+NnBEG/h4LkUL0wtFQANm7fSd2XtvTHrErMx
VLNhywDHLSU9qnZCOsS3a0wDFO7qry7eH8/mS6ZbtJ2jxcQxgbLCW6z/XhvL
8sN89YYe8BxiTlUaqQq4fN4i+fzlcAQ3nqKyGNcus9G+pAdC/+aiwLp9T7cz
UIl7EUjGab6Zu3nH082rM9L1fyZ3oYmQAX69zjjFGk51B6kKM49Y8Ae1pMHC
R7o2dNwIOHA/TgWDp6FEc6tjGFJRr/aNNpNHCicpHnn0LiQouWofGW+J5W2g
XtoS+eKscbZezDLB/TaXfl2ALdjrSfilSoenn/q+s+2BNxzBzjHjmYg2sSXZ
6DiPjIPCeGfKMmjV3GZzCyF3KA0oq20dUr2evUEYslXXSTw6wo5a9qXehax+
gwQcRDx1ttpAl+EPiTSrFQgLypSWc9y3ihxMJhVdj2XW1gAoRkWvqbhmkaMw
AuvDZo+GUq37a1pxbjcmRqsXYZxT38E4l5ALy743YfNALHq7hrbTh9DdoZPw
BsgdeKtXeouv/VzDt962Nw1SM5H0X6IV1AWokgRM4RmzXxtq7QLmTmTe6LT1
8gkq49D5BCuhYAYgFsaqSfyWE7vZ9pH9I+jElDDuqCl5h4DafRaIba4bpRAI
bKk52QCH0lf8FgrAmbLoeIHsFBcb6C1DSYnNf2fhE4u/5qyRKkEHaQ7ShN0Q
KZdzKO1ewnW7HhZsIkIPiW+qmo12KGv4ZcRsY54rEyXzpdkiH37w3AVnLyeZ
l9YBcg84SQAyJhr05PTZt167YJLJB1iTyoPmOx3O8RMdLf04RFIUquuRFqqs
i0rllbXF7Tn5xDspvxmtq3PjpPu6CE5UZk5ETHAx0RYB3fo+4sSxgZ0p7Nsk
HRwHbVgrUdx44YdqFYYLBz/nt+G09VQif0w2FUNUTt9JFTFVWKDJHQDeVfAv
DzTw1nymqoafvs/2d+236xVubWFmWNKIiM2ROssg0RUr9QqEKEPS9sn9IdvW
1nxswNLjpdMzrAObkNLpxTIDMXYU7RIU2+RNKZpajzlDQOHvJaO1GgnDXxFc
WOURLBsQIqxARUZgauZR9h3ZIZ3AsVW06p4uGWWT8xiC6JF6tLc5qOLuRf6K
nWM+7YZv8Zf8H/tXn3lR1J4neh8kj1yhj3h/ruz4Mdj/1yGQUad7VyqBW3kl
dsH0KQWju+I5q0QSeAmw4bC87+XfosUMopikCSytHdt57REMu+yWwxSfqUc2
SkcGXay2sXQXXEuY6RQe3alEm9U234KGU8tv+9cLnsRduXfEscL2mix0oBsu
rzTtIxOgbrocPoEm0NrfyxTa4DlCQEFAcvMqkqsYlEANaJKJ6bUbrBzwQHcF
jF+CJzgleTI7mZwwAwYTvcYZJAjiup0o2a6kjFIS76HJdGkDmd5jtSi3JqCv
Qr+aZNzES84YjMyS3dsrY60STv397RSRT8ecxGi2VekfowOuj+ARxYKhbLFe
rpgl+yBAXEn2/njlx4+PtKqodhlDtKlCb+ackZS2xYz2eBNbpXQzNlz/glu2
U9mQLbB9RdehAhwxVPcbum0iVw1TKeVGL+CBJQX0/0V6TbkcYQrvBwI8hOzM
DsFjYteOOaHHZK63f2kAmzoNhRvM8YbD7k2ReOrmQ/Eqc9mgHt9zW/CQvaQs
Qt208vohT2G+FcXF2NT67V/fiIolKwMV+PdV6Ed1GfEfxQi5nNr5ioqhbV0S
UGN5QB4YYZHxsqBxWAzIq4xS27sJgmdMdTobnf8qmg5l3/IGNIt1mpWepMHU
+2wZ1gsXc57nNgdFVohl1W4ezAMMFDcPjYcq8/6sKfKRKpDZor6ZhgCRJtyY
7OBbzSo+3pAPWJVmESvgQwvCptQI5B5YXsae8F0QGkmxEf4NnRSgO6NLkgaM
ZujV9w138ILKXmEf8ZekR5d3xmmHCVDfpU8Bg0bKzqUuwygLaBJ5pIz9Kod6
umfUbo3afwrAHAY4JDQoV4SVqzqg+KdTL23tZLXeb5AIewfE2NAzDT0rcU+J
8bAAnuLjWEjSMlQtDGJlZyLoGQHy+IFbqoZlb4eokklPQQ/L5Hq77Cs1YIU6
WZIM/73e+04cI0BFIpJOPE4UDXddrzDnvYP0b1yaI6s8XTuV566l3HeYXD3y
TJUFLFI+vXFXjqYquLIrZs4ihSDwyfptMZ5HqT1PTuU2IFitJ1dXze2Tj71B
fZBdp+AN2ymMK2pCAjiLNCxQ5SmJP3HwzGol3K+iCdDUgK+qdQ0OhbDrGH8k
nnrRCZSOENUt8FFbfwl0iKkHKR43ysBOISZzcAWwfnn0UnyMGFb/Z0b3x9Ra
UJ8yY3vfFa3Qt9OOMO2dN0CpwqZw6/tBmR19fkYV67vnDCYg8ednVypNaMgF
GRxXJDO6ROtO1tSFsgK9Gvl9h1yDR70EBxGDPkCTyBnxpUY2ef48gGhf1nZo
gn5dK4UcSoP6tS7p51O2gBJbfiI7BtHpSE3//DeEqDGxnuxSZAQ0U2qIrl52
Mgmkbegd9aEOQ5bT7WDjHZG5Fq+kzRsnJPAe5BoPP8Z/F1LiJBxA8of1Sn5c
n6GRnVb4UmsuOOGdhcqruMkoD1KIoesAFODa47KmcecyTqIwY+FY8kz6Vndr
up8Mu8MC9lJFA1Rc4hzlbXcmCgeXbYE6iBUXWFa3nbmbEAqFCLkLF0CjJhVR
CF3Ohi4TSMgEKSPLXjCgN/LdHuDx7i8AI6eASyoqCUvlpsfVwTQ6zHuSa+Z8
/RJm9+fbwJLIY+8fJOdix+PS/uPLbVNO2+AqSOBuzOwJ1Hef53Ma+/GwEYc8
SyimRlr2VERrTpWQTfyxrEx1ww1Jv2boYVv0eJWBRr8iQQFv8FYIkAsS5SWR
KagkUrmudQPEaOCRqXbV5P3R0iASqH6VB0PgkJqaDqOJDe7Yd4FZq8AaE3NK
p6xbdGxu3zPxOHRw3Fek7hVZmayJJ1Y58sQzdudNsnJfbzrqZ5vOdvEBpdtW
CB99VQtuNYo18v4+lmKDcYS181Sr+Vz0GwLrK+A5Piw0YPnx3keSMUqdlhYh
hf4jQ6pFq/IKsQssVQ71MN0CI1GGX9KUMD4pLyPYnw4vOUx/1etvzECSXaSu
aRA8mraWfzpnrJpwC05SFLCTvEIqwPJh1C/HI5zZH9MXDv1SyQ6glNMFq7qW
hyKnp0xIxTJoWpFI3FY+d1qrXoGLxBzXNez8L7iHIKe34kUw5JWqlCNtSVDL
aPmBwyLI0dCmYeK64fjTgFab4xNRqoDSZfLX3ROJtA69qVCaf+zci7bqCIeb
BRJnCIcVxadTgA7YClrNoMT+zOxPfPy0ZHZ+xRyiWyAhcCb+Yw41w9nG/Li0
OXzqGiZ+74i1ZVcdjL3QJB45TXQMtvEG0CyfCBiu42LHdmNMrj9WumzEOtOo
mhbkpCgch96gZBXCLiWNVBm+4PUV2+BKkcdVLlbJsiq+5ytSheW8hRqJ4VLJ
/qZnQvHhutvZMlVYTgTnfpn52uQgd13aYoCCoPuKZTaOhT695JNumwf89NjM
I8E22l3q6D+DhstQgGPCnCch3i+fCmQGZUAYHhjkQ46fNB0kF8soLuOBVc4t
MuzoL59vXFuhYmpxwP/qJ9bGknDeThuvCRC+ltZ9giw5bA7i4mLyD83nGUxv
6YDTXNBMr3q9Xlb7Pf+sgkymQM5h9MihbuTf/mh0ecWYBGtWvP8hbgB9J0hz
zjMlws5uE9zuqQjOfxNu2lKIgnwNZ+oGzwRo8IwWLrfn4ZJCLfZZsd5owHZi
TPbDsi5S7C15LNshfu+8u3rO4YmIDdKxOP0TMrkjdFijzAgg9Ihuioaqc1Se
Bx4ccUxRN6vqLR7Tsp88OA5bMABG6kQcFy0Kp/zQrHdn4Xj0MDV3XjOADkai
wUTjxo02Pq615CmaNQpkQpyUVULFu51BiHJfRjbOGF9CfAh4O4CXSpwH7oTY
TzdhLw83RVi1wDxKAWdA9kaB3HzJaQLMqFVkCGbO5C/1Y0acVkhSAb/fIQnC
liqQyBCJ3dnbAKrj5i9toS7uk8uzX5ulGqb5aeYUTk/2DZHClweilZNwjgh6
ua/WHS/jbb+Fr5/dKh4m/fSRUoezBa6U/HgrqLOXkUxiYQhnAiQQbybE4CUB
PU+FcEk5bwP8LH9JTjjKKfCO6pGi1PS5TZjB/LXTSxfcnoq5HJJhAbDKSeCA
AR4oVJCeTRYWqtK+/eNjRUcao7SvdM7644x5GYW9d+FvAg+alNy+y2NGvge9
v1k+MYiXZZW4izZV7ah/zHgSC2pX+nJ3jVj0+i+s2S0GOZXf67JyLyqQwn36
Q8KlzVtk2dO021RCCFLoLqMIBq7CDp3JLUtTAwcR8ZtHrgWhCDo8w6xrLDgm
0EehkwikJDQNI2Vcy3WCyieOTuaFWtUuFBJN93VUmjb90yvypojb3r2owTn6
B+o3UlUBhKK7X9PPUbEAv211Xwi7Xtp7IB703tLJsMowesPIGlFvnNspBI0U
2qEsWdqHYz/Tg2HfvOIylUeYw3zhOsANG+QZAbLl0+NcLNndOHhc0u762shk
TuDVMZwQ0TLKRc30C0W6VK7cqqzV4DZKDrJNdRgL/a+HmayKkYfCEEt9G55q
a29fq0d2twu80jT0jacGbkkZ40zT0PyFfdmlEmp0U44tTNmGZsWBfVkwK+zz
dP8foT6XOT4fCLw1kt+2R7j9jfPGCOar4pT6LM3QPi1H0CvivMlcZFhz0Jvt
62h2Egib0xcgM7DjDrTyNbIUdvIecwCzmnXcoC+cH70q0Wxmr7B7hV3CRhxA
TNfwkCEMoXmgVIjEDNHXGGyeYWdlMKg+BV0Dd6X4o2vZJRQsXDzgmhzKMipY
n7Cn5nl71Ds9dqvloIoi6xjuBx1gihlEPHen8pdJnLp9D/mjy8MnhJhaSlb1
IFi1UCoPP2OKH5oqdqyLNOXgUtJfWQxkNphN60+9sbfBHZ+RzN6n20dz0Mqd
GWhvA4nKfxJPa8VPmXpef2OB7lBGBOISn2Nux/DxhQkV6SLqXZ2nRcUX/muM
Hg+ikWqOY7IpR+1dCPNhxUzdbpkIa7dsLR/HHWSSwgKARnGWctwe26rvYqGN
MaIlwJw7H7UVJDKtQ052HEbWduOL+LfTSFJWZMNXlV0zYHGH3kQ6HwFSab+s
lptnXAtgAh+HBe5QWZq/3pNvH0ilgcFu9c3R/jSJad2OaPX/iiP4S0wFaRMO
fKF/4dPTvUORnshPPM4I+kj3xAWQIyolz/COEDzzXrqqrVZCUFise9Hk5Bgo
B12NSu7Dflfkoc+gjuzX4QKrAzqNaQDNXc3otl/HbFzUUEl3NvMjnDnZn0r+
gpziBSwag0GKza6dTZDxYzHAGI3Ew0f4fc07iujC9Ljn5t9h6To02V+C8sIk
VWS+T3CRwo3EtTHvb81oUJFOjnW3a69heogx4otusk566LfeN+YY9mrDltma
VuZ7x7Pzg1Q4Z4+WINNa6X9QfxxbFyhrZuqy11lOO940EmJvx1dfEJZNxQsk
cdMa7L79atGVrp8E/1OfuNsIp2I5ckVMzeRlReGLpnPi32BBFzksN8Rk970z
uJKU64j5FYAtd1I5yJNw9SkpkWnv6m/woLvebYHy0Z6TNx5Lg73Iayvvx+M5
AnSxAfQIuMvETTQxfy19FujCIzC+bU8AJGQqiLMUTtkP6JPHAFo6eQjiCzRK
k289r6GJW2JPff0057kIarZvFlhHaTCjmOzrjK3Q8XFNELoWhFBKaGkjryN0
OjRSrRgzVchLVw6txSWawVFbor58rJJDFeCHGj3kVzt+/LBKBjXYr5R6ESt4
pqrX2AIEUfFK9+tSLHB581i6nxpn4kDwjPUWgpMgPQKZIYRcjmRBzF6N5W7n
623O/l3dNoos+JGU/RVf1JmCcnp12igRTqJwDxyPLHXZtolkW1BHIbBflkch
hjgP/EGl/CfB8g1xJdTd2/k/uqtiZSsxOcPFQPaLfZi8hwhvUOxMktOsTsdF
qenLa07/DP612/zwrjLV/jI60d93L/cMOr8HQ7YqHCJVDibCRvBpSxMARNCP
8PvdDS5UX8Ek9hfxlOFy6weXvha+LI2feioPDhMObBlJ+IDEK8dOxMBI2E03
OtxZTqbPw5571/LwCWoPzknmkli85FNTEScPeMaOzQWyYFmuTHpS53m79sJ8
8z9K9kcYjI+yN7YC+af1IO0Wus5TKCh0K0a5G9beA0Prd8EitIUu/zDnPGcW
oKmwWtTz9hdQktnHjlE6ghlwKadl/Kk5DOg7pb/gTlbQWuWZDX6yKEQ/do21
pNqEeSFA2XzJuo9qxauyerolA8mibPHjXjVmu7d5FjgVTB+B9t5p5lkFip6x
9M3rSZsCOB8fHnQb90pniz7Q5XGD1tvE38gJZoiKIj3HuqEp7eRK22azRW5R
xbLpkMDGBQcpeSn+Tydzqf1YBGNcl3GcHxrqeJbuOYkOHV2w48EVysUi9ehR
JanuHqVMDmmcLuf/F0I+sPyhOBy0sflzfAVanUe5m5AZ6282XxZN3Zl+owPp
HKlgbpFmu3uShwgyux63KJNMaRg5hEOIbjGVplbHDJ5l9w8AcS3XXeYL8F5U
0gMtBijOlEdnImXUfkro3/Zd614bra17QYjUhR38+/9KAEVUw0imB5J5b9f6
aVXevcN/O5XuweOjARSOPahqVJiVNcopThUoBuOmxpGPOBVN0m1LSbBtmvxf
7cYp4JyMMeyY8+X1lCgC+l5ZlAg+T2kh3n4IFNnm3DW/FpI2KFhvzkSTXG1i
PhNJuiuGklZFatofG3Qb64OnOJST4WOy7pnr6kt4JrBc22p4RgnC33KLRgsF
1/QYyTX+uMJvVrXR3TO3l7CtClyVfbHPV8W5XwCacTZuyVR0jKiytnDKYEtO
IGNSLiyHdKM5nXjqV7Kp+uEuVNE3JvGqgIQWZxlGwFh++GH+ZI28NBoCFd2h
P4bYVGqafAESFpl1+SW7xHlKi/aIppJFgYi00Uau+FofJHBa/9gnLRpaU+gT
WverJ01+6nThuHyDJ3/BxB6cAEGtlKzNcm8Ler8OOtS51BFfuh0CSbRrxNE4
Fm+plPZHBaOsXqkcKVB1S8pjoF5Mz4LJbSTwPv68Si08qgsdfc5rt3Uv/fo2
ujkboBuftCVXLmFWHEoirDaGAiw2Pkenj8AF0BEtrXshCwx3ukq8VMijTv13
jPdGVS4s6UdnJPMgN0UwwoPbKW/rvTNjW220SxrhpEvPlqmeeQ8wqD/wO/Z2
mCZiqKPtlAFJyuH6aNxmf/8GHEoBW5WLDlb1ptAuw70tNQFA1bsRx4mFvwyC
PDEatwKc9/JNZpcblqRGfwOL23dtsnZfw6HkV4Dt7mAJBkD72ZQaL6IIhla4
Y0gZ6j+QQskS7OAEZyO0v2hk/bpY7tOiiI98YIWgMQh4gG9YB/hfC/b56Rqx
hMiXjXMYhnbLgv42mG3Vvj7nicZngblHgvyaG7C0sgzNqhJSu6dBHqE1ggBa
Y+Y2GRsf3+UEvmV9a9kX88ReD1+JI5w2YVfFJWmAZKFQ0OtM7M8/daTlIjaw
wsGWyYs2+vWnXhGr8aOCZFHijgCPbeiWqKQ4NEm/WDQbuK09wlMa4vSmEsKQ
EJ9hsiU7yeQWYEiC6DB4Vq46I8T4DsLavYC03xi6g6mIuorCdgqHfUcC8IcC
If30vPf79BxVzoGT5gFDiKB9Z2LSnYq/UnL6T82kWIGEfBcf3A9Ul7kdtFiU
AMG5+11FqFUjqP4H1Ncs0iyVtwKfokOyKtNE6wCD7+q4R40SY6M8znlY2UUA
3Q3hLmK3kfQOvUlFeKj6t91PygmafSDKKXBkSoRYw2XlM6AH6tS4nLUveG0m
43MzAzenJW54jZ9VrosAEs+iP2OyRonbs7zY8WqDfBT7hJZjSrCmMPfbO2nD
EhcMIk5OOR6o8wAZoNEoUGRlfd/xo9cGWKZZFn7y2EaIsJI3YXuirBBDhzif
Kx6AbugCux2oJg/02yCOEkWIPzcSyGhl4fsG0Zfpr2RnCE3SNGwBqWxOEw5/
2DTeVHhc+DrkghLqBRKeXlsrAZbaRT8b5nnh1kS9Bfa5UUnATqOLKNIuWKcz
ue08wiohRpDFqwvB/31s3fzxA1qI6z4hjyPvIiTxlbWa+J+lpV3n8ymYvCXk
wnoz2mIilFtS2ZJ2TfrEl46onw1WYAWRgCTCbRwBi1L+2psHsDAHMGqQ7nHD
XHZR3XocCG1LZNDyojW/wBhd/HTg6LefvojdC4N2OSXrWJW2Si/xPXkH4AXo
QIvZI3/3/2jJsHC6gV1ZUqP3rQLuSv/V6OP8fh3PlObUpfyVnq6A2rGk0ewE
VV5Q5x1/o7xY0eWedamNGxff1M2q5LCq6HkSp+RzQAg2Z8KYeg3tEHTct1zk
hWegWwlVes0LKn+QuAfaJAFL8V4vb7YN1gHllHxRr2gjzYnPzdNkfRDDNSwQ
d6Fv0Fgjtil4e/El2AUbzf5gDyPE6CPHRFHthzro0BAUVDsyCxOLiomrSLSP
+mia863MVfCo7hZAN7juO/7mzBs/PqqEMxa9vzZNTs8W2E8ezIhUmX442ZQV
WmtQzEPfNgO7gd/ATbJFmZcPlf5L5u1+VamKzVJMs4SZFodTorW3ut7dkEtf
Bmyy9TxNB8cLbJ7IvP6po6YCuiDiaz8NWmLRvsYCFx9iXaRznfa7ztG7Rc09
Uy05D22o+Yuvi58IVHsLXEmifvw9P+CrIjU+LvxaPSSAYjQR3cWZWnlFlBqZ
VKnISE1oNQE8C/gy/lpnVVbLd6eUMbVrST+9jWf1zPgrjt8WluKx0hvH8O9h
GXY1JuuBdnuWEJP1DnIEZIyl0mQ9P8L7GgsqOY7t5puqU1bwEfRST4zkCD4r
wBJv37HsJm46bdLzyRkFf8hcmDYwtoYHApsYIeHM7KAqBuAAQra7bUc13vvS
TIhlOalS0slycmBCPUGuEyQqQi/cEzcD/sFO3ARr1/QxWNhF4jHYQh498BLq
qVoJgAGZ3uhEc2AphYWLkqiv3MTV4vSEXDnRckmWTBJgn+UpCOVCZNsBmB8y
psTOgGh+P22KaaHHwSV/XJTwYYdpHMfRz7wUTQ5/Y7VwzR5+bu8Xf1M+Rpjl
r4MRI19HoNZYiOUtfcCtHdYmeOEjKGOsReUSQOkwOhbRjChDWGAsM6An+Wkk
7hbNyqkvaHFd6H2gEyQnhbiOxdBFh/Pyhd57Uw9WkJdEgOko90qRT45nPgr1
S/3Bo7mNfU3FeXkd1XvwHh39UTzI33BEb1xpJhID30nMmuCRDLgXrRJ+aHtt
W7/MjAosIFUkVJxoeKGlEBX98ElLA1VQIymBXcgS7eD2o5wjyTFkk4XgGHVo
C3mBV6xJTKIukjQHv9roblLNB0xXxOqxmAk9HU42ed7xRcOt/cz0Ln3tkLiw
+udvFaMk1JKmXyQzLbBB3XX3y4+oKVOQ13N/xbtclRnya4ydD0MBHWmSVkCq
PETaUkFiOiG6pqrIA69hYNmHvCSlQ3GLzZQRIYt/PZYVcXlMSjiOioapuHH3
/GaMCQ9Q/dnTB4gpUsHiTcVwzQrnfkjIH4fEk1CVD5dg5OscDU7RJMQLeOsw
Y8mNj0SDY9yVDnl498mD+6AEPjKJySL8yt2AopPq151EdBs0JfDtBE7HftVo
GWN+f1xADemwABxtJwD6y6zNUZPBlgYg2T3vVPDdAcLGjnw01BsAe5b6I7/p
qn6mn+MBazApJQpc+tJONWPdDdfSiIh/PZfK9Vfm2ogK3hqoPFvSokdC9aZF
HK7/Z0V2sShOri/CPBke8bSTIuc7EtiGWTj3TAMSd15wux/cisx5S09yI9QD
jSAQLifeyPhdG01VE+Z8BIg661OZhUWitqpodTYIvG/r4c3qyObdjgEwTFOX
+Hhhrw4w1V1BPCfvD87tw1UpbGc7aQuHfEUjMTAjV1jVvKwdSO6TD6/VrtAu
2sM6ESHNt4hCYfd2lGhu6VcPl7Pw9e4UuGaUSEbsf2/UEZIZYGmLloKHcmAE
wVq7RvPKwUOTAlSWZBUtejaHY60RAlN3rd9PXDBfsrzProGQEqkj2FLE299j
7FCjiTMiYF+LgZ+GoEhaafFjgRqJ+16JRkOWDya74++raK+B2638in6fzwEE
LqlJynXJygerwzOLzVoMt0bALHXIlSiJZ1ap7DLYBYgpwoMmFKynnnGoUcOr
sqe/vUREU27g7s2OIzmVUY3pr95fnSMw3ISxoSnNWPhTdmomYiGkENkESzoo
5rKYdw329gNo2hCaCdpezhPgY+Q5sxc71W3O++VhEP5Au30E5t396cm1RueU
HKzWvRm6DazkWNoT4b/9IKIMqABx3k6GFS8TDDLotx4zGoX6RHIEefWNzgu6
HWP0ccw8usu7UQula8f0ZBLangvEDgrbQpR1BbEakGUSVPer9cwpLMQnOjIQ
WN/MkRbHBqhOmt+kgJcab213TI3arcMbhGAcybbshH/RyBxlN9G01oYuRP7B
FuH0UextSgT5nPompnAHy/0SMw4V+wnCachBcJTbfTHP+fjzKxD8DIG3Xg71
1B41X9826eyc5xfzO4aVAIsLZfVYvIooVeoiG9WKlj9HbtHYSZhaTd9h3Xji
QCmeAZObK1SVxjosO2llTU85K5/j4v/lWoH+lSGsGOTA5mbW6+xzTYMy0N6c
ByGZosXoTrPeUfOHfNQq+z/RJCaHhsu/O3Vk/+DDoy1tCErqnyiJaPphPbh5
5Lu2i1+Ssi0yWr2JiR5xvSMRqhXUIfGWGE7sjWA1swHIDiDi6DkAWOZQojDU
kg/+oTBL3jADO1eJdlhPhaioXLahSebeJgP5JAEk7TrozFVPLeWCMVQ27LzE
HcFNhURfghbQbm9Zl/4dGx+tAI8pQ6MGGrc7qDRhZ4rC4vXaJFtCGyMUyslH
0guVg2NHqD+l9bdmkrTdxVvcKtQjcbBdst9NOU/XNGr+SHyNGFoYAx3BPYYd
4+zYHLn/3fxAo46met2ugF2+NCPM+QzZQzBsq0Ycx21ogFQsoEcHGVVG8dz5
D5ynhj988zAaa6oKi+QR2Ws362+emB6zHv7AnZRUBhtXrmiBVxSy0qgcUmvA
ZxP5MzS0g0KkkYci/EfUXn+vQdPTym83q0hX+jZrQF8aTCxiyYHXu08Cp2Fo
lOG1RlsSSQa4jyP/v0+/PBWN3WhoGTLKO0qDz0f4Y1vs7RwJnglsepTTSvba
jBs5VM2AHDFBrFwWhlmzvUzce5KsqgF+lnk3p+7kzNdc+XBPpS0Q2IPkH3vB
2RGrdXp+rebO9OCtIvAF/GoFWr1v1krTfz0GGvPEulhK9o0f88WAS+ecCkFD
/0P97SIxBeawAnWsyy7r92EeWvslqMzCVQd9l+ZvowHZ0V41/pBcDnfBT3+P
uXsgxqsWcrL7r9gl4oATBbXA/MWwQdqm6A8LYon6RhHu9q4q16WKr1HxoatV
3IlrjWwS5uJ8jJk1cqDrXx3lDG/a9/dlJAlN6doWjh0i1haSwxrrYXvmdwpB
bgeBXYX2AGnk26IELfhlSyXG2Kn/LQxALJDtOqta97LdKFadlAbcR2RWsgBB
xQdhZxk601FM9m0gAKw379fDO8X/AfoHyKYyJHMiNqHDI0/S3gTrIggGV9MU
94NL/DDx27gdmXEn9sJZq3mt16vRsoFM5VtpVe2nI2L6etj2cz03Wts/xD0F
l/cz+ynGCVekbB3w5ZKameg/3L5KYS68boFJo3oCL/o/eAaxoiQcd/BPw4h/
qDbOGN64GVtwEJBTHn4qtyPsLNh9sdfS4WQ/I4Ms7CPZa6oxC+ws/B72hdQb
k8Ax5FV/4vtPwYyvFJz2NrQ+JXutvmSLScArtmI6uhKq2xAL70dRCkwZ6Y6r
X0OEWgjRQx1Up5DIFY6fmLFKm054cqeIyJk0Yc6f/qO+frDxGRJ59EnzN55c
o850J8CD9TFyvntqAq+ZV8sg8DHIH2X/Hoq2cOv+KRTlNvaq5NnK8NLQM7G8
sx/1ySvHxthXFcBYlX5pISvCDYP/cYv21FMhebFvrpWqzK/0+5n50zcLPPyC
lJhndzAzbswVo8eGUN0BHpLaaYzmoQZvG1uBXKek1gQFpi0sskPY/TlguYXi
mpar2Ww4Pn08snE7dLg3R6ETyE3YIWGa1kQ5tAVn6RmyPsQaT1XQt6ScrYxn
43B3Fb4KyHhBfI4Xjh5tSe2D3gkxBoPC6f1cMgwGa7uPrwHMkaOSxCN/Ipts
6ES2YX2zs238/wThFHcdv6bZMEeKQEq01gzPD3BDa/8uD8D0hNUEfe/bWmYB
29+lmOL4E/dXJ6wLolbPH5q+j7FTw9NOssZr/PVThnDisvJh736XRdxK0DoK
E07x/wGKC6vz9QSQOPo5edFu8dhX/0hFDRvA2KFmfjfkwDbPwnAI3GDH0poS
wgiLe4TPL9t3d/7sb18wJx/BDkToULtZCYRHbMuhdvxcxjSGPTLMwerajtpT
gosjFkGxiAZDx2lODRFQ1u2eBB+kJeRpWtJ0yzcYwlz20VVgzwNgpkjmO8ff
r0oizp6MkHAYfepgzbbwypFdFh1CZCB6XSarvBd1iTCtFTQH/jR+ZQ8SxrPA
MfZ1CCmw7yPYetvQUrBRXujRDosVmjar/pOfLvN37hy4S0EzUbgrHSflDqdP
z7BBhIWXZLY3nZ9QQypq+ViZwbIThjrsbH1pnbhBg/sJM618YxK3hLz5YQC8
IgBbCABHQRcPBxFseNrPLd4IYlmsoJmjgDywf1ucNmAZtpDGw7vmmsyksulI
/3wok1ZdzVd0ODs2eGgq6cVXoNL688gbzMofLOJwLfs8hRHV6JrZDRVfWUZL
hnMIzrkW+oOARhtVx9Vi2ZJDQi65vcCJWfWb4+H6fZmDgVyo/JSk8dcAhD91
kz+mbLCnPa0Ts9Z/2tUZIZlQlSAI36k2ArigYyEkgXe2dJZq9lFvYMga8yDw
h7KNw3KLJufdZD95waGWzApPc0sYQgND3Nzm0wu7Rp3bQZ944VflcIxeoGS0
R7s3DNnstF56UJMeuZ9yH8W5ovboqLjVDpN/48OXv4c6NIJjnHwQx6ITR+VE
+knwQtclhYFIGF88c9t++RrCgXKst9Tuzjm4kj+1EIS2hXhAfo6SW2zGLgKc
Je+LNxvMDG52qY6gII5KVo9ZtOmWZ6XqUF8O2y4dktT7UruKdUOJDPrXHiAj
yWn/vsjRhI63RkzNOLWJrfiqIPFhyHjqUWlVT1DIOb5enD3dn9JLPawEfZrc
cvTE1AK277WQQDuZask/odLgS1GIfwB26hYjD2Src4EEwLCJgyBoQEx2gGvt
wOuHNZohMEmtpTY3UMBu/pr9mFEkQNxHyixmlRcQpwCBXEN1FQqHN18h6JMT
AbMvxGzOIqoiFcczS3VnYebUMU9zAhMwf6x4WR5o/C8CTl99FIppitblM9km
90rF5GhNP67t33mAJ51i+HFMFNnN5TBm649RY5IfOyvMgzay8AG5d3IATnh9
j1qmOFmDWaViBsG3uQPUmGXZ0j9VnqWSZsnpPSQcrWjqcovSdsHnkZgcLh1o
szeOj49/Q0BRy59GVEH8epB5OA8wNBZgdAoSXSu0h1SX/vmZnGxVF9YWLY1M
CLxzRvjJ/eqSVHuA/96ALWiXU9cm6wOL9Y6YHbviv8R90HmHPrIzPAIJIK8e
4EbxoxWkg3eCiwBaEufiNFWtyyC2GdV7/YpbB5qvkQHv9qaObTOq/P90MYWJ
bRQhB1GbmP1RPl3chlZ2Gj0iWQ5DftnLO1GoQ1HOApCAegxm0oDgSseVDQ6D
aOqKrQjrAW3VYlX6b5ii5INMRv2j/nLgh/KRt7wHamnT+r5k7HN1MBmxB9+v
BThGxVo5qEqdpMAgt7fc4w0/qsC/G128rBq0eLBWKLF0pqnxjfGI9nrgjmif
ZAvUsl76X4Mq3+uuEo9uw8U9emaKCRcxV3r/f0I4QGTlsmoeUscxpvEVOyn2
EGPMbKH1SXQ1yNGsp2ykX468jPR/J+uARrFQ7kg1TSlSzYVLSmINBq9Dcaw/
9RCuyuBCYyZ8y6sDnm8WOOtk6h10KYN6b6AeE81YrdmkRZ1mFW70utH6FZ2x
7Fc+utu+YNMc1kd4yVo08P26RTu7oDE5jtjX/yKClEkNPnkOFScZAGIcLdf0
JG76MGQk0KqqKEaVv0PXHOFcxvYQGjTj0yInFCOQPJBuhTw27fGmNVtj2wS/
s0iYOqGvWgWhG58ulo89GDKFPiFPnHbfG5H1JR1DtH69CEPS3d8iMbHm10++
HTi9kjzojavjaoyxmqefCws75zdvry/Ile64co6MaHjOmMGI+MI0RXI6Mrlf
RvNlMtAqBraV36Mbynu89W9YvW3XovM4XW2mc6NkFXAHTJ2SkvDHU5DoUKff
XXyoVlYUWXDQbiHqMGPmoRd7lB/CQG+NKUAMytHiPcifkTn90Fpx5ntQszuJ
oAdJAH7JiU825LVgu6yMOCK3K95f1X9864c3H/LjpdI2VZ7Q684o4ju5tbBs
r1r+V2YIgikmyEU9r+UaxigOUCMWZx2ufityJtqnB8Toxv5nCGxoY9ozaqcm
9T7IyZRUYCn86PCx/ZaOnhtNQtUPoDCuMPbwmunbPw03EKZx4p0/XJS2jAdZ
wG5FKv2Yr53MQuJUPw1ZG4DoUTtGk3rQ1BMisUkNYMM/Jrei+P6puWbJA4QA
jlqZYF8kXoWxxHJ/sQi68RGGvL47oNHher/GNqhQ4Z+Iirwpt/RH3V5lUqhn
jfYgH/vEUNIuvWDJrs6awrpBDAQ8j0WEC/5vuMMtOZaZyA+ALCLTkneWKsxh
BQb/sVcLD7T9WZeCLAeXRZeX93dH2++NPwPEQzVu4ZMbUNRuiichjHBSKpU8
mxypbor2LYLXKKgti/ExKMK7ab6qFiTkl90/C95ltRUhsbVq5ZpQRr6/Hose
F5sJdMsRykWEmK3hrsaBJ7NJlMsAjWea0L2AhHm/qgUcTIRyQdtL7xoBfy9Q
nXZoXaG5QW2L5iZnipHmsqQmXD69+KoSmvhICzp3IMCbei44SAf4vdTzgPTi
QlVdqzhBjrPrimAt1tbZVrn8IjUXmMtn+RHLhYlQroMRaRTXt3rCvPRm5VRQ
da4ztw50a7OkEAQip/Xptva/2FT+TZDrN2MnnPQb63ft+PZzvnSH6trnuZGB
QlpG6QB8AATrwHWETDP8DOm4hty1koDEcwBirM0Tf10Xxpa0uNtLxMn4OnTH
/Ndt0mllsJs4U3YflAJLSBT1yAEO7ZfxfKHF8pCkU7teQh10y1YNWOU/RWVl
SZ1wULuOfHdRR2vDGrfda3D3Z6bFfJvNPvGzQ3O36UHYVPJv4cUoxwFYQpPa
95sRUL1WRGuvqieCaLYzT8Dgz6q5JQRfjBVmVvwsDOuTi4AEA3YzORGcMUDx
6N0klhcw8b0a68ENkbkLryWsoyRQya1ke+1p1LtmFR3hkrfPFQLwbY4f/K7c
NCE4Qw7nIWoSEKNiDFRrLD+FmcwLRfBZj0zWqi+30SHLrJuGg3j/PbcEdUuy
AQbN1kXb6NTavCvaXIJ/N6voSK4/vjw2/CYoLuIN1UdGT33zPKTjiYZllmZm
lTHjoMdeI+TA0ftahl6HaQUpcpruOCzlmm0b+iM/2i1yo8htS0GWEQpEbH4D
Ff7brwEpIU2IKuRdWqvj75yB9iFX+wz4+bgakcgLzcRbFi9RA9uBpY7C0IG0
RvZXoiL5xFjTvMzuZxOhBNCaR/uowGeQnUVqBYB+UviI+mxon6shUcTmL5gS
ZLGf0MX/AUPCyHVpwGvGidX8O+okihs2TCrRjirO7DuzCVcA1FDWfFkGFFUy
4QqDW3yXAM49OQNB7K6nMFn2qcpj7NRb0/WE5cLRpQmVMRz2UyqJivKsXYrn
addcXWDPCs+1Ys3RLI/HjlmZ2Fv5DqPur3ei4nFpM098f+JoJt3kLzHR4SIJ
XExeR3eRTevZpUvzfDjZu1+Y4C4l0rzK/uCTBSymFKLahdCj1QH0w8hwZ/Dt
5dNA5PjOLZ+6b8TLxtiWmVIfrQL325PVqFAQpLdgf8MRKNYIw7tPjinOAl/c
0+wS7f25rOsE3pik5C1aoChYTGjX4MyFD9r2rGtWQK9eqcUVxRjNfyt9zB5W
DV6hMlDYPIrLAtc91XwVyu76KB2RSk5/EeoM6kPLlTIEA1oh7b1cRAfCCKRt
9RYpVrLujhFoT69OZG5t2iUhSaEMOBa8qQpRwEheGz63zyF+YjECwSwbVKXp
yQlXBod49mAsM9hCjWASoRJZIVvcFetJo1NMc0FpPOkWW18tSIl7oufXuqz6
0NBS9lCUkWaxI3nWEFeaK+rQqy2XBjX1cWTdB59R2pRmlDHfkJomk/2kRsvB
PZ6sC/bCZBzpVqqF8nHsAZBcsGLng4iun7owYJhG94oQ5BTJXhXoZexFzqgP
m96fwE1mzbhw6ogUe8QscOjwk+P9BTGBwWSJxr8wJrgu6PbIQFXsjVBAiptt
EtqHFJe7KbeA1G2gGR3G8P7QAPGjZ+xz1BafoR0WB5wVC7OaNSvwf5M+N2w5
rBGkyu6cNvoMTzo8DWf4KG0fgBYa18lMIGfpIjKkiPGlPa19QArlhIdgVdAM
in/Hp7LzvThloBWk3jGmP4eh+ViphgwF8gReSZi+9V58dIrEr40mAdJgzBGZ
n1BISmx42x99F6wP2VBy7ReNvJfTuL7Sd3Gpxzphv+MdqQR1KLnxewP/DXFy
eLKntQO1jMxjGreJCsUw8VAmixY9q4Jf9Lktb3r2KriwJXNvW7VPDnAutFVf
MF9uLKUOAuWqpMP3LxNP5hUZfshoUeQ+c43I2D/mZUD+r2T32C410SfbmI1P
pCU/Q0gkwEXTBxRZXg/klrpw95i/B2qkppfG7P9jfIuN3xg3podYAZRPqO5a
/ELPiPCz575qwv6LHMLKDSniB95eQSCoWBQXVJhhGWBWK9Up3YVYbEby8hFj
RcP0tZ0vrprZUVX1Pv1t5yXhPpXMZ0v3lk7x7ibUtXmzBmiwUaK7Uo+d8yzt
dsOCHQP3B8uff0qaHQvUDIP3udtOe4OMo1Wv7fpklq9nv52+WNuwtHRX7I9S
V8JZ+8a5s/GFIqyrAH2J3HHHmv6QNNtVzYBki86To7bT9GW2yErC+vL8W+U0
zFm6wuUpSNjsZlKtjrGrL6n7zsn4YyZrTtoB42upOkSl4EUxapqeYM6K1ZGc
gvc52v0p7MN3inHaOF2eXAQ25rPDoT2kQoOGDEp9KYHf2m1Px0e4hwdbQfeU
FAt6LPequzgtV5+aG+d5guuYkPmP8GD+Hv603GXQLhM9yJdPYTD/r+/jJvef
1xxbzvR3jp3y84GgWD49DRMSTwEW1dZabeJmy1jd+N1qtLdBXcxNMWBby1yQ
2YdTdu1qMvP1ANxDAPgeh15wAYfL7i4EnJFCezGEVFbmdaqer2qAcHFcypBx
7IjClotRmvNpypHebOdQ5w5rPcp/YNpf7SBvGJ0RiQfSxxormV9Bu57RRfjL
+q30Z6N1GtGlw1963q78vEBJ1zbmQc3zT0HtnU0cfctxBcxpfD6dxK2lcyCq
6GjxpImTKevr5w4F5GST4b1/U1UaFUEkyVaK3RcHHK6ejfP/mXHLjfUGD3o6
aLtcWzY0vNO5XGm0ZaG+zguyAjr2gam/sHlNpq2fNxRiHcsZn6Z7qPe/KhUH
qyubGXCCKZOamK1YyryOkbIJ3bQCIWyqFxpEELkUz6GFBtdhyOSypcny6XU9
9/eLx59Rn89Q6rxD6q5leDwbfQFLJZITfdnoWIUb2KjVlmVs+EhSFjTidKlw
UlB5RrazkoO58EZ1U7mdmGdQj2ifWL7YrVxFRj7HM1hyuKGDbuBxHJbLe3zv
ZLDFaVpkXgSiVdIXX7GyjZF2ciPaD3sgFcZKxIrGHEwONVTBcoTQ3g1K+Rn8
EttTcMrkPvQqSFPtCPcd86RD4u+7F5sqFTNoNGcAko2gB1J8oWk72kFCa6/k
v7ljCOx0T0lH6WRyW76fYmxUPUjXPU3zGs2xAXCgmLG+OKC8PDfeixrpHU45
bA3a/AAka8RMMuJUdVp7Ovetjx0n/AhYxjPgX8DAgNxbyqJx5lWGUkLZbD/u
i1bOrFk2AX40YSS5dQLD3QUiwiAej4H9jF7eJadvymZ87rWq5Aaz3/eRQRkd
zEEgjJoTTFJ5vonORwoU22RA9egaWQ1WA2tOhY6vcT47xKStRl5wdZosT5uF
TFjWzYzPhwH7RNoF5nXNPEt/xL6849dkzD1xtb3Cl+hI/L2YWOe0Wpj+S6W+
o6eSqcgZKD0ljhlXD2qxP9bzWxTXIUgz7wpw0QSyjtAh60/d8d8g4AV84uoI
Rh+qPUZ4M7A8/YN8HV+0mRkdCoR9fCbMPWI4IOn0m/EWGeppdAABBGqzOXnQ
UKVoESCQ/djo4xZOAtRxPciOWPwDZkWcG8JJh86ipQyjJBLgCGHJyFNmJHCJ
kwg6xtTwDoZgTN26YXTn8JUlzjlxsbs6+frgXt4XH/A//g7OkRHB1CE0odFE
VWkfZBm2g/KQf1Gdls5nuOwwECCgmT9S76WOQppCbdYEBo8WFK7RSrqYIwz6
/H6ONo0c22ICvgeBe5pNFOlchKkPPppoVqb3QTKLewO1vUqK0kRFTRqaBDUL
+l3yIrzaTmjfNLdc5k5jyy8xhtjjifI4wWh0O+p1PfLkdsKn5hNfaobVGpIB
eZ1PqNcBPKu6uXPgk8G3f6ns+Xwoxznv/DpSZa+8A3lqJZi1qKy3o4KDzHxN
7srend7AQ/9oBAQ4pK+E1o0XJj0+GMDAqaOjNiyTH0Tr6wTbqhkDo9S0WLmP
ftZw1jtyQqeR4L8Kw/I3bpcXtcBjpQ8Mz4CtRXpacHhJQBXEuTKFu1SpIrNz
J5bJHVxYAHjRBlH43Vrny6bOuQO97Ov5nFb7xphUlBTptG3ZeRxHs3rZ8WR/
y3rjj0S4vf/Isg/VM0TajWBPHlfpP7dzrUSrwGlw4zypVvJWNGB7M/cikJEt
ImnQEhonzWT/tXOjvncwuZhrNS99KuyHQmSrcKnmL05tALGi4/GqKJePwSwB
H8dAYodzFBbtDa4INmGSMDarmhgienc6qfY5lwAgYqAB8auWhaQhZ0+2xOfT
aQ8xvOzfljZv7Pn/GoPhXcajVqjlgFyV2gligDPp49uPdJfPevo1IZjyLYGE
OYm3+UGfsXTAAd103KW3Sz9kSjOWSUhTo5xF+6NuLvGO9PQvi1zYmGCtQty+
IY75HklEvsOD9SlXN1NrfB82lepLVyRzkd6QPOsM1VBcw6e+FPErCU4/ksMy
ay+SywxEpAVzhBzRX8vH8jTmkk2kDX+20ls+zi+88nwd64efUWT6hMbqDqHr
BwrQw2culF6jqkGKusugB4LO4IhhXPArwKmDAILAHSiHrbWLxXpVyZ5mrVZU
u1h2Z/QG6jvX/b0v/yQanp2emB/34joHLaLQmkaFc0FLF6heePQUU0Jv+T7E
lWzHlpYRuw27RMDXmJaQ99yTqCHRpP8G/QfHJL4kY8caYHMy2TaQnjeNiUoC
R4yE/MrL1uv9YVX/tJBxKf6CR7YAuvRwOTeJXaIk8eQLt28Iopc3pcN1tSuJ
gkzqgI4a4IV3tFKHfjd9C/Bt8i67vOL6Wp1clIKWwzhfweB+PAaRQz1kGvrt
L4CZKK5/rfQYAEYvf7x8xxCASNQ9EV7MPh1Q+GDo8NOATkRpSPIT348aNhsC
NeJPU4kzyrb02UhzxhLSYJHyh0RbAI1CMPZQRtSeQp/HmUAvfQA5iHRpyXcZ
xPn68It+HK/yTZpHvcbWG+5LOsB+/4vRlRKD5HBwNKKHYkVKeCDOg9b4UzD1
OyUD075oDPaTHX+GYdBXHXUBAicfVAm8hhkuuHU6Pw0D5+eHuVem/Is/Tvjv
GjI8u1vOdxPnL5xsCjuCrLOL/eniqVR/BCA0lM++OS4LLxAu0P9VdBGR1GNc
4LmC1BRoEQR5wScmoooLytqjX49pAGSiIWQlmYEcnJbGkBCwsy+Um22bIgj4
3mgMCRHSv9ycC2xdHQX1vksb8xpeGByxwVc5gV2yyBGWdvwWufvaSTBFZLQU
yggGOULCx6f4XHHVtraRVQCdOLswQxZVFs3ORitXEVIVWyEnZiH/P9zZFZr6
7zoPlqwwmwdgT4+v4Z3hzpptRS4jgx6rHq/xim17a1NHPWLsVCDvvWvg84/0
6jANdh9BHrOC1qKhotZgCopIToJbuxuxLxOGeQQnl1gFGDLShTzbaru32oH/
dRL/RiZNYf8k+TJsltMlwA7/XX21V50GvsPciMIBWQt+S6RY+/IK2h2x9ccg
/0oUeiSTMAR4d2boV+sunvaS8UfzSf3w/spMM7oExEbU/yzzaXdKqMyRamJJ
DQ1WVAchAMt61YM5ozplOnZCaMNG4Rzqfwd0TgzPB8se/drsULkpZhr7PX/N
WD7wv0hvUFq92O7f0qXoYAjdqe1xiaVXPiftSlNTSfdAqPv4Trn/CRWZDYtO
DlNACFzVwVvipVMy6+Wr7w/Bd58LAxTj3FY2jDqcsxYBfBCUY/ichZTVS0Y3
4y1sX3FKLwQZbDumBbs20n/BNq5K9LgqyteU5bS6knToRMpW3iYMLSboWH3a
5DsY4MQqN+k5M3aN4DA+TI1xGsqhegfyRQHwTnPAze7jZrndq0bFZ4zVpUBC
Qo5fAq4v/OsXOv5984SNvK42W3CKire+YSjtECNu3m9qeuVJ8AtFibL7xxI7
ZROcMyYzf7PtpaRSXSKCQ6IHiiNJ916C4R1QjA7DDy4BPxtCBBkpuQh1xKQ+
JKAQMMURFHDiPKxou/5VwCu6JfVV8Yu7/PLsdD/UvThW5Yp4d1ZGXVyDVuUN
GwwEnpFJtwopiF5gDyZxUnL97MdOHuyRKh4AEwxCAOkmSYtLprq1r+5hjyWa
F32Vbb4+PLRKSn9ESfPlks6QtM/tfrPtJV+7C8UqIQsp+Apqwh0QksKoGnCR
vgcrVOCZDeEy8AlF4BJ0pu8XhAeCOopvE+FsSc5960Sbr9TXEAEFbqoZmA2D
NQ/naNysuCvNYz0X4AL21MZU3wd8Wn8Kh1vHQHn96y5rxrzpofPQSWCV+YuQ
FTgE/V2qUJ6cHshDzjqN/7sguUzeblXNriwyBZZJYryp6GWO5S4yIub09cSw
2b5R+o9L+0c40eV/61bpt1Q+iXuuYGiP/fNgqbjtpVkAxy7ykuMYrB4wxwqY
q6wV8PFlMhauAbNeyZeI3itPnogdXLFwCtnuGKSjrqT1qCm40hxxvZu+fFRs
7XmXoyU1iwHL104dDfRcVABu6OP+l/7ABJZjReEJJkt6lwKQLDAUMaeLAz1A
YWsCiXJyFB97V/dFomaTpegKvedushtE8sk3zn24PTe8YxsfxssrgLO30SaN
etJ2Z9Fa0r4+Q3gmmK3jmxDXqBtOdy4r1Ciw/u8vcadNInuncKl9S6ddxy1z
cRMG0dF2LtLgz/KA2pqeN8vFMyzBph6X01NXsks1N5ijROQF1OHbrBQVDVmZ
BO9iMJvKC03ZQi3UeYC3IXDFaapPQDVLC6Cbs24FhvR546YLB8gk7t7D+DVR
eMToD6BUaCsuMWSoKLGja8xT4rXgbdmJvgTpDRZaAWzAsW/RKoo50OAOwALm
K+28XyYku9Oh5yMBE9sFCTMjP3aFK7XT4eA56Zidt2dzasaaeQiiR+/7RflY
bZbRogRG2kGjjPfFzTC8dGoJIXcU1E/WeNS0SFTFPR/nWYO8zYm/mXVd0axr
1gsZh0Mh2NKtitmeSaRdGkCWGaMF7LF70UA1MB9jFnVkNV5xppTPPTYsoQFM
6ryB8WnUC+AoPM7hDpzFisJ4lMIqOIJWKBeR6s4Ov5cB03MeR3RJS/gmL3dC
2lpdqTvrWjnB2QdrRJvo5qo5Mzp7dAmysGnTd79qJ/6b0+NepIj8w1SVda2e
QHIUkOg8TTEGKjZbzxoTWdS18f+PXUuSmLqwi+YEB4YKQwXc6FvDTbrau4+6
uxdq8ye3yt4QIQ/t/i9aTTw/KYD8yQrgYAqSHF/696pCcNRUcCRCQyKMIalI
oN5rv1UE2/jQ/glUzbpbRV4GC44Acwr67PjmoN8BdcK0nqSwH4Cmw1EcHBFL
KVg/fWoGnFgXXiiM63YcByzP1HHJM+QF627ho/Z9qJOjFngyTVer3i+JtJ3l
rLoiuU+P2LAqNsTqHhNwIxqKKYQM1InY9BZOLe7y8CraWOfo9OHf88zp1ISm
XkxnX3gLGjD0s76/BtRDtK8U4MrJ46fN5L47WS9fsLfgD9qBvdYYLlzLmeOK
jjP/WLPHNOYFPzw2Fx77D19Hu4X1VBbmR4y6abDWOyNkztTfYE1vk5bHt1oW
qgDLZdFBIovOQe0OWCcFDvHeFzFOIvL4KTcjGlAbek3K2ZWQgUAHyCVsaXub
7qj7dYWhypQ5oNN5I7wRZlllTTmNE5KcTqGx6jjcIj8EBXgYHjIKxam41wVw
vtsgNNiM3Cn1qBNVcG3kW8h2NOTH2TBnAj3VMszUpc22jBKZ8uQ7b2cVEpb7
KAm5vN33Tj7hpJD9rd1P21s29jf6WW1ddH3+J4vxYfcgtVe5HEDZ+svBfLkp
G7TjEPyVbsUq5xnx6cOZI11a/nkJnZKcvrJ6aSGYTNr9Em6lPYhZxcaj/JrM
QBEcSj54TdCJt+Vcw1neptVhGylsmxQ/Ib3l0sz4OaRalm8/7C1P8LDe802o
qEHMBP2Qu7Kr7G8v4Petg4r5P0Fg4fCTAYuHS9r+NOCbP0S1yUE3EvJImLe5
fFhx0GCDCe+UN/ZvQYSCY5xnn424Z3Nne3mbsUK4Xxi0i5kIp3+6W4bFjQ6P
DkRvURfNB5BurEi48+U4v6HmGUQ1NKanyAWvtdROIwZzFL8OvXmenL+Mt+zD
HEsTEOiaE6dFZ0r2XKAmFHH/IThDon0Xxg3NNHpOIeNCSH+0yIO3V3uobH8j
WwZVfbm/mVdaLRHNjp4YjSMLjCq2V5G/468MR+pDP4C2yETF7SkrsGDwA7QG
HGgp9gfkzBpU7W/Tjng4BjnQ+Ou/jjrYXPlYJEe9M3DGd29E05I7QmvvkGjs
SKSYf1vTTyLOpYU/1X4ZZH+sJQMkP293yXhaxjegwJ+lk10eeuM2cKKDW4eR
1YH0GSUYzFS9xAqALiR0q/cnpt/t7huug0kTrhKabdbAIS+sBHofe3TyTAtP
JwYXwC09a82t7Ng7Z+h72mC2MPIxZ7+cx5vTt/KmlS69JRZMOaF5oEinRtDG
/T6rENbcWW4KX0jpH8BsrFH5pcyOoCVu3faxtT3k+yLinnAAWkbGPaavh96P
CSIZ8OPFQGW3cg+wu6Mbpjguil09AKe2hsfxlaDNfd/htpbzLZyR4/9Rz2Fm
1CWpKqaiQ6jOAcTLnVyKZUScTrHtw/4M9l+UadhODO7PSzPeck+Sg+zfq1lc
tBxDoPE382Q3Sq+zKK9JMcGTqBK10tc9ioBEUDLaOJPtoCXvTwBbGBhbSiiW
xGGWsotn0YtKMZpq932u7F5XQkI9Ja6uekro6DYq9GN7YxTxojPP4ENF8ueY
CWSam70CszNfr5mQi7rWTG3SA1d5boqC/UNGGi4LWmgIeMLxP6El7rAxs1yU
CWKbDwynqy/nhVYSheNwBI84Yf1MJZDjf04L/EF2BZmPQx/v4UN3CMHbMrKT
Ll7A7124sgnkBpE64efmASmROoCX9gt1p9XDu0917L2zWrmsgLetGAyc8O7W
D3kWvbZedmXNIu4LTlbyr/UubfoEJpQ+Klk69AVvlBcuR7yWmmP/HD5a+9K/
DA6g7mjAfj5ZtRqTPAJRp/3G6u/jMWTKuG7Bufme7Q1WcAyRvMHJRxnHmPIS
JsuyzewIneXgb+BEsXLs/R5sMPYIXjdoYddtdMW52VruH6tOLpbRGAlJbepR
HjpuuzjMaJz0POEW8b0OLvoKVRIJA2AZoy+mG0wpdWEBXlvJEMsrxS5BvaE/
QDomVmvuwYPeMkWTepiE2h3Lbme4N2m2k86zocxFDHApD6VbwDy5yKetyCGP
w7+RmgFQaUQXoVP85jaTOF+kNQ/ybo3wasrZZ2l4UKom2H3ttDMTl9hYsJGr
qyGBdVHZKoZRzUHhYDDiwMbTYpt0U2OsBc8//5dD64dnDztQH0huZyeHSxuN
4xxwBaIxIfACAAjEK3Wa5BOg4TRnZWUKjKxibnHScpHMbskIlz04AIJTApvX
x90nZGrKbSZO5LNvQBoSiZyi5+4If744XiA66xqswv0Zkq7CaUgCgWjmZ6ha
xs+4mbl+WN69C926O3o6c8PMg+MErrcXPKTTHZZZ+6DN5fhoVSdDXtOWQmfP
WUqhYLJoP0HVeVnxNLeP1MPxspc5J7d/VIrrS+5//sOOhmZTDFZpzFaAgGTJ
ON3BU8zh9Bp4B87cDbxP00P7tW/bj1LRfbslMfWi7aXeG2MEtf6u2SST82ev
et0kKku/UN7QTII5ULHN2Pq5Ciy3Y08TKCDalxFR6/5S0pq1RrYHZEz9LhiM
61iYPPVH5nW6yX3flCXCMIIcrZVe/n9cHk8+B0/Bb71WX2vb6fwhYECqxHKT
xTu1KXM8KjxBa2tXt1rzdnVShcKd+4t7FecAmIdLBVnKM8f2MX11kLSDPRhf
X+qQY02Ymv9GvQGWADCpZof6xdTZ2ANb+Y/3oo0JnotZKy8hfPsSi6jRJyRJ
3SkPMu0dt7eFMvD+YaIm+RVrfGBGvQPy/NQgI+fwbduyrc1mIxpOEcwVN///
ApWFhYxs0lKetXmVOBGxeiW3hC3spnbTfRd0jHwOnjwD8Lch6znrfID033KQ
nFbPJxsLFNN8xaqEzdLuhDP1HhP0yzTizmUA8CAHsYxqhUsquj2BVcJTneJJ
eit27bmpONBPtEjkqr6Uvkj0L0Ww69+aF6DSJ3l6m1uHg0lGonAfCCjLGdAY
Y9g6eZxJfnT5zaIg3K7CR1OTyYiI/2nLcdnGlfnohHliJvM05Ds9s4tFSOXj
VCqnOdt2JycmKICycLjal09QAbspdmKODfq5jOBJNraGIFj/9Pl5qlu0Tt9Y
8dJ/uJdD5ytb47XkQEfqxf4BWTk6KT4CHhjYlEFkT6qPiyjvRrX3VQRDPd1z
CcGxcWymNOk2muN/3QMWi95ROEO91A22IIb/Lpq42K2hskdCkDiBkLKfNLWV
iRkX315PjuBREuY63OAHOAE/EbUlid5T2zuzQ0/f/ON0LGKRQSQKq8XHrUcx
ZYKq/nXp0GHXJy0zpPcLRrw0TAPlm6QmM6q/EW1BFw0qSlrmFdjAPG2cvyg0
yksHJ1I+nABzWjvtD7FoNulSXwj3watmnFuGWHCtT0RxxpMvsxqDz3n3H8Eb
V/4clNGg6t+mNpI30KophkEnQpfk/maXLsLTgXSwxcBmbSDuVdlh5uw1lAXl
72xVDksERsMfEZQn4h5xMD487KxG3NuCdEpAb8tPL/RfWmrbyRY/wVWKGzYh
IIBX0Q0FhTVzpjHvhvqXF0dcJs1C4rNqf2YClp1Yzga9yda/WW/Izm18ErIW
+aCqYeAdjooaLRSRT+zx1lpSQ7TSlLjz+UNu4l8vYTf4mhhw1IYkj1YiQmhH
e0tCEqn0dLtb/APsxMpvb1oexqPS0399YB4J+D7hkGb3d4ClN9N49/zNHgF4
pnyH3ub0nVroapctTIAkIviJjKoXHAzsuuoEqFPw21tv0g84VH/cYE4kRGS0
LfzV0jxRFmRcwRrev3iyfONPCys3pEPAQa3VQ21d39DDb2KhLMfaChHMV/jg
sZRDeO6NR0RhPyj00xER4GZij2LgviXq+1MdYku+hKJ1BjJfYkvSevXv5JNW
n3b547WXRE7+DEi5Kvs2zUu9XJUbvpV/eDTncSVFaBK0YfZDd8Ya7VFWDpLY
fy9uPon8GPjCmN++ecYCfWlHvehlqcoJoNksVZPQ1ak/wZ3SalPSgR13/Tvk
kZXUjftXxlNiWrksRZUbdtcia4d28ELCFDX3zNFYt+iL8Rg8CkLi15Hcofu8
l1w9zfxyIQ8FLnne1KcC1EbbmiqzY7v7rT81ji/zNYnIcsJZC2btur9bR8Bs
T59NFGUjZjemGG8smnJ7yNKbZBUQ3zp0NyoVOaO+OsWBiDJ6PRKv4TL7CY1G
b+gFYk7LVy8gWtT8LPX8e2UaQsuH1uKxW9Nj/wDxdaE8kr2pBGpjAWhd4FV+
MDnwRj3JaDmswlgsUFoB4lPCnEHDT0k2Ny7eB5lFRbL8VMX6k0T0UMJBwB+z
2Ixxk9PgxdM4QwNAB7+uVr2jDV4chMY9swjCoZobvyo0Z0lcK4jC2CGimDCu
2lQgMOKPLl7V1tOF9uTFIOK9edB2A31uZFnYtZf0l5yFkUSroqnTKdc5nnsb
8GBaHioythpwZ8eLz1Ii4rDCV6btj3iQgomrz2Ht9E1ryehxCeXTzxGvvfgo
dAGXCnQHgaVwMzm1jybILZai6seuBOQ8y4FO2g2gNaIWl0uwzj6S2TeIGO/4
1WZTdROmUITU6clcBSfrkgKYGlz58KXDqVmv3Nwncv9o2RoB8cXiyzhqx5sS
rQRYyl9gq/YkDbJA+IiLy0kkDMX8iY02dHSXhEF7VpmEEcUUJ8XSv4+H/xF/
sW5N/T4qt3/QaivF47XOHNUbyFCopNDyNWrPQwC414GL5KYd1HhC8YjM6x6B
mgZS1G7j4pwDfQxoiFuvrkzvbwnAzZxyuTZg8UbK9yxMKUx936hflenJaJd7
J8YRQelgmCiN0EF4UZrRpLkQsx1Qwp+yyqyPmcWA9gtgsGEdy8eFoh1U1Hua
r+bu3G3YN3NBAc8/OWpCLZYIA5H4343nupJlz8dPAWENlQ03GgWDL9mHFK2U
teb6q64TIE28+1rKGBRUeLYwkSO3XkRCRz4uTqLrE9X8pCiGbFHT/71mubs8
9K19+nlGffLoh/eS8USglTd+gIjDtFKcS6/K0U8B9zwEmbXjCuB7Gy70ERsn
lsh/liIYZnYimo/JeqZ8wpIEGTLG6Xow14ga22O1CtCsjcqPNlQdLy1096JZ
Izl0nqhJbqN/Y8wdmglgTvlNTwTR7wCua1kFn4Q54hblEIk4P5DCbQYBzgPq
4ZUKTqcQTYTPOvXczsTgS8gRBguWamN76ixPqBoJprPspj4JJrtNJFL6LS02
7AN/xo+v6JbuqH8R6910QiAX+NPyne9gSgeUlGfg+UDP57pWxK6yaacrkRN3
FjhF2KPysc32fxT4cMERgQytTKXplrogzYKeWxPGxxJl+B/I5axXKqfq4ejq
lSe2D/oAl7KNQ3yjjHyZidGmgVNv2KArrmBlIE/za1zpnYz6lkhr06hdcp1y
AwwOuk3irvevuZ3tPPCFy1KrWsLnuJg04rGY2tvcoXNTrOwULoLnPWRE9m+k
ofRolO/1E74Q6pkIffCQNLvzyw2vdrOUYeosJfCTveFtCOWLmpJh49E9vBS6
uh4FMuj+A+sZo/9bzheqXIj0SjA+2/u/GGZJG80NLuuUfrWbDsC7Xid6R06h
zywmty0oy8PRPgi3gfPuTTSWgfOGVGf5KRRaijrjvGnjBJIZSagquCM0RmHF
/ADtd+M5ABNirKihfRCY9lK/DO/6Nc8qkk3tzhhsjJEI/L6GN7YkbAguoL0S
yjGVNWvE+sb6QXY8mwDjyg5pwkaJeXPlglxO41fNZi+SE/W7XMZBTxOA46OO
T9acAl4iyBwEG2fsZh92g3NTsdrQ6B89qSCcg4zd6TIUVipoTiiipP9ki93M
w8QyMm+rv9gycHF6apX9akzu4vwJl8SdA97Pm6I+0iNyumAYGugkbQTjbaYr
KLZkEqrGPxsBj3ox6xjuT+3LBCxwx92TbmhjjJ7bW4iQ4dkAisCE6dTpZKMg
LoK4eZDIl00H6qgtfME5X3PUBqwlYmbLxUKoWvfpAQxSufkQVr3nPKsHkVxM
5ZlLptbXfINpfdBvMm+MC7HZXcV2JLLpiFfXsnrAJoQPi8Bi8hB/6ihsyW8P
QiX6YBU0R0Do30plrShClISgbH03Q/MzX0AcoFerAsjn70Yt7L1b1n8febCR
j7hQObOf5k0wKQJeKTKgHaEDhvF8A2tI1OviSARMODOghMR0Q+SkIOiNLTtn
OBPymurip5hT5O2knEFfHBKX9D/NXAOQy5MC9uFILFdmWPyIeG5pRFsQzdZK
CjmuiqKs1VHa2R2UJa7gyxD4OeJLz2vhydQW82cl5JYaPXW9SwD5uWBIbJPl
hTJMSNhj7TSrduBOfJtC8xXApVYzFnfQb3LV3ThvKhOHMHCvLYrhgaRZJllB
O2rTwordYcQM2Sa58Y4LiV/xSelo1jqllhhnzxVqKIsv3BsEWyI/og537Dg2
1DbdZjKLMhXkBM5xTVKm2D29XFBBvSt97J/2PxDbYmhPCMD0MiCkdsxFXAjC
Nv4s6vnXppsVGsa6kOvcpVWubTleZ1fkFV6+p2tH59pxSUBYx1AccPrspCBP
5pP9kPL//XbJ6pAiDBiDT8O3JJXAcWWlGHQaTjhYbs+OPCxX/J/qqAm1Jpzp
98dAhBksyPUp7Tv+9xVsBtogIKNN3z68e+8ZPIIoq+3iGL5HFiF6IUGPfEZW
JMK7i1JCdSiIVQToVi6Jzau6wQ4P6MvVjvHiA+WMt5s2qfV4AxktTil4GrdG
9+oHa6nUYrbphUGar9G8oCC2QT+2ejugMvmSwSAJyLGrrHvdJTnk43aYQFkH
Hw8Lnt5ftJQx+77u2C+fC98u1luuH6EM3tO3gps+aR0fpP6DGmQAfJStGDDZ
Kmdn1S4TJ7bqz1fU6MLta7xXWzwCABQpx+9VzMZfHX6JUAXRiknl+yXXqvoi
GruAedtOEodJYNzpb5J6MJH/wGZxVI/JN/rinegttlK/a948GR+Crpj6a22i
sjP2zrxlLSyBWYTtmIUlMBYAkHakE2PNO7S0YE/5Oe01fXbZPFstejdZknXT
hQtvN3s8oLu+haG9KujutYPlH5asDJHrBpSpsnCquzNQCkLYVpLlnnVt5wpg
n8e/avQN8D/STjYgF0Xk1dmaE3aGINxDpPaLmPjUsTADdNe0Igv7AojUvtvb
bwa2RgQiK+fRZ1u6GzCnqB3XmSnIAAezKaZQ/IYYD8l6H9u50cOA/5Ee+OwU
VeId9OI3x5Foltgw0ZUvVTg7wBwwR+Ap9swk/qhrKldWhf69xvm/unAHdYUM
3ZmyC6ntAaVi2XeXaEsP4BUkdhWSMlm9tldEFyGFNHO2+FEtnU+qspT2MauQ
I+THm5NseXg2Ykzc96utXf/EAbLKv5tcGMHtGAgRNxeLVmGMTVBf9WMn5IsV
+MGnRtVeFaUbXku91IzUrOs3vP9pNb+Id/4CevK/46qC5BK2YS8RF8/RRW7d
OQPH5wXmAHudJZgDsq5gDl8O4Vmrk1ESyLeLb3L8p1GR6RRWHZamCKllpYD2
0BbmfZaWi2/9ovYrk1M37x1ir7aatkCpgIRWAETFco9n7T+4sK7bkumQXyxR
lh190thleYr/4Kc/uCMlQVxWF9JcegzR+S73lNpi42lhKhvRKFCp7rh3BwBV
Gep8Rs411qw/ifo3IF+drKWTfMcXi+3FqVQTsp4FF+5/sSsYth94LBc4j5hb
+zZgYyKIXMuXnITzkUiGJgSij9JuEt/QKMV8M6hofNMu8GOQ5mVvoL21r8Oh
075Qorc98SWfabsgdgXwFjlhn3ClNEvvO1wwdBEuJ3UcLNobXIBmws0uL+Fg
icm0om84AWbKBDbYmbZcpxVzxhOvM9GyTsdEg0/8fQQ0h05JZkv/dqWIwwSJ
z0Z2e+xHMWsan0FJW+I9OR8P8ZSmio3I1LWL3AET0sERqxQG2vVRjxm8JLaz
ne7/pfvm9xv966fQnkTOMaqXLDS2WAT5z9/jCtkJpDvO2DG00yR3e6S6tKo7
5+Cjm0jweqGd0zn8r71XCP9z8N1lOfcrsJOH7ili17swSw6ivB4f8gX5V5lC
y1FnU/ZYAZFGQMzH2bHa/hTPW+5ozVqTivTn0BIEALbUAlC8ugN9khneGpnk
0y1l5QZtPoVLwWcJOBQ2RN6eRpbLea15WqzkjIPHyruTJluYc4XV6g5dfK0k
pn4cDGsXGeE9FbOcMsjchqN1XMHLU9KguHjLc6ZBgAdo23Q9rY17RpP1Bz0E
mmod2goflKv5yvV5nXSY9G9OVrgkDdZnNgf5eaPReIdOhl8tiSxuXXIGy2He
QOw3hvSOosziFQkWB2ToH7BTOySvZGSTMdSVA2TYbTtXRl+APLkk8B8aEb+z
0i2aiL5+pc0rTC9Qio2wgi6WtqUhm1NfNtoshzf6QZPwyBPKBLJuafU3S1ep
eDAHRfcoV1diUiSFRA/DKuThjhADyi5aq7T/xV8srILx0Exp4c47EM+2vdMh
oyNSaymFUE43As5F5dFF+whJoeUeRzJZveL7z5KoTJWN0yqJzx4qgtUifZWB
C+/yyUyetrB93mZKOtljB32pHVX2rhQzcAXz8+tH3aLZh4SfwS+Femcyral8
MBxSWz38X84eg7xpKfP5LpEINgL6qLZr3nbo+nWSMLD3cAyj8N3UKIRMyq9/
jBJSslHrLXiShBTEJ5k3qnpeJJdQg/mWzkLwNY43TfW7sDTU72diY8rhh6ol
pECziLpu2cR2jBKdwLPSlaBG9YsOAGp75azS0wscLBkCAoZMFJlTed+WaQe1
pcx+5VebwgZjsNuLRxfS/M14/tg1o7dbR1HYcv4OhwmTJ4k9NMf4S297wexa
sIuKAXPa1m17z2cbfxarPesBq4xnkUyrZmnz8Cvl64WLuTHLm9kJmxK08PMO
/fB6wC7ar2uAltyzcMNZV0D785G8UEaKq5YmFbmooOz+XkyC/hU9kiUK/FcT
cq10UnU9rabToHP9LfIMximCBw2meLJJr+522/zUvtgBCP+T9LpmF40ree+n
fZ+sYdOUn6SOu6onNO+jLqOwj+kkDC2Xa7MORTyQVvnWNjBTZtYL5pMDd7zg
AV4K7gscFadXuxdZ2K3GB0ZgKkuTG4ec83fqv8pMdwMtAydnA6LC8sPjxCBR
Ns5hECPeb2UWd3RZDtKWjOfXyJTYMe7Ikd7fg68PHQwc43Q/9EYd7IMMloiR
fccMxuY2Itur3GojILxvHUx5yKVks/5mSpqx+eChRdaPIxbZ76YdOLWfmoyP
jBjbSiUJwforjn5j91qZYfdU//I7Lx6qdQxUFDUFCzh1KLSP01ieBt52tR5j
Tq0aasFFEmBwLtRIfjWpCU2TjR3M3A3gGPKStFYEDbyhK4LxkIJn6ukULOwI
Scha+UCbDIOox4MPzMnl4mrxSwgzlPIjUNCt45w17Oo18lSjblZbV9o2DUOK
h4/aDqb8LxinFv7o7GLXomjKSAdMIEM7wFBmBZDhEwNewo5yoltizr6IXsAi
mCzEuSRrx6yAraoyT21ryJmo8kXQENghX79LE7afGBWkcq/kW1n/seRnwRLX
YsPeDEzpemiNGDebTy+2y/Kc+tsjrQmzzgGDlEIMwiUDY97JIs71yEl5iskA
0jTthn9yN/6RboonRUHXB7eytL8cU3mxMLZ8u8SpLNm8erMvbr5ldW/1ZjkH
5293LudVrgSpKnJndzW+bp2KrozHz0Zab+WYYG0dcBlrTlDrJOV1IW/3g8fb
zR3lNZQV4I6UgIwU8WUsZNeNIHLch3TjAsV8QgO9hW/wdxl8M2aTrCNf2WwM
fF25vgqllQF+fJxckkC+5sBOD+I4bjbKb4ZDdFSZqPcbO/O0EJyNgoemCXhp
n2CpXJkM/peRZCfXaSerp9XhK2KWs2TUOZSPvaHWWYUtxEWW4Yr8lGnZjnnC
uiNnihM86MqEf/M/crXhKx4GKYYnXDViftznzSuyTxVTdaOwOEcQ8mjPik4s
6/+ABoONgY5ZIcZaAcWn52/qUW86TgoWZH2Cf8m/9DORLZqvSKB3qf5d2/7L
PltBffgRHmmmSIj6TjnYzIGqyLXeAFH5Xp9sGJS96z+YyRjOCwsGQLn9kBEn
kcZZ7sGbzMqgqa9ZgGxs+VNsx0CZtXT9CEsiOGRc0QgpxKQYjWzgLpNjuGDj
kRlFSF9MsKMW2RKHnKt75peD6N96rR/ck28LPcTbTj0lq5AjccP6P6DCwiyV
JLhu6FJHFwplsJvVfd0qRp2S2QZ4XoZifK01Gxj6s6o+4SrSyZ8TdaLMRIME
uVoCnacMcMho7XFlCD0nsq96rfGLJXVwkYQP2IIhWWGvLIUjVn5+qJ/CH/X0
Gj/k3GwMvWvW60HkF8L9/0WfF4pWUs7u47/+2XszUzkatHt0KmtbnxyGofF0
nEUzrrxFo31ot3WgBu0PwJrnDz0XSZCAeFeidIBWwk+eIXHeVbdl/IPcoXyP
8ucc4j05u54pJZUTPyEl/xEvE/+HhEQeeT/l/hvuk8N4y2qnRK55iytfV0y3
SRkA2xERAZsgWz31c+rTqXzndiXLZUr7HGLYtYmjpq8OTy06C2iATVwwt0zh
NHOH3/ZOY5TBYyKWRgyXCNxWio2xPytQF6GdBsOOfOERsuSIHl32x+wjJI/w
TQjQp6zFXl9PZ2wKGuwdB7+XOgER5unSFTJi8Brs7Vx1i9HHRSu3KAmGEd7u
indQewC63uVMLNMTY0Vo7RO8TSdTZJC8yppnwpGLF+kw2kcssoipaQ8u9XiB
G0gl/h9Lc9Zb230Y9h/B8nroFdBqd1P6PxaTEMj+lHxBmt1o9ZAMwjnPxTtk
JHTGUfvzILNyMrugAyWLrpKl/shn1WqCor/CfeVRVEvMY4/vwk18GfLfqHc/
jAFj/xiV4z6Z4IzM4OunhIvXJ2EsCkyr1SByMpw4XZYr5OpdDdaPpAs7ZvwB
hUfdKP4WNcl/FkDVHUYYlFsxdV8RNF6K3VPOQMcFZIvQ1kp4oRjcucHnwcb8
5Svxkt5EGHs13ZNPIcNjWcvpdVBxb5k9E15YJCw3RQ/72MEaD2G9g3yI9zpH
fNyrDhCCozAZgiTOLowtgEtWVPjuDzDa0tmOlAkUTyjHYCEDP5mXWJ3zINXn
AZ+SZWS0xkQAW7aP8aZFlQuXkRdiDZdmE9QK/iVEnUvOpMwDf3PogEPVPAAN
Kk5isY6oqBfnev3hFh1r9bu5WhfDo+n+S/vsh5M4k+mSFnik21LdVeOtRLwv
t507HMmof6OyV7SG977hjVgnoVvl2rc916AR6GS0JdYauH6nPSqQCu6FUi5E
u/8IkOxVW5XSacjcxaXokVKL5Ix/SDEXap/MDhLGe8pAOD2qj7t3knEh4ClZ
Sc6KofjlTfriUMlqzyH3Bz1NWm02t6eOM0XjvaKpQeI9zY/HLinNOSv0nnga
WStUeO7jzyjRS5lfb1nkbSHxq2TqpgsceOH3IFPWsBQfIvczPKQqBZUIqagY
nHZ2DBtzU+vvXzsL1C+2bxrOPbifKjdmGhv/KrPevU2raM2Ymjrx/s/YGLd9
A3JISYBrXP2O/mr7bkVSqpqNW+QsYNnrkS1qDANvqVCv9iVczMfjPXfJ5DBg
0JERjt0SdxOlxrq8zPkxpjRYo9W6DvP8xzJisGqbofsOfWntjJsip9/ieezg
HlPw1XJ5tPFmTgi5KAqwHFS0pARufdudMFfu7oDDhEBeiPTA05sxZTKEuFwP
7JXeEdG0xV3Hd6O2Kdb68Q9PBRGI7aMZNnxxHENU824uOVZrCYhkF/6265bk
T19yR0UAOTbTjY0A3yUR8tHqePSa/Mv8s9woV9oEes/EpqRifCRth56Md6GY
hFYruKQNajdcbhkOJDwIqqXj841SKMQXgMMr3dDvvaE+GgG398gOw57LlCKk
29SWy2bwHfcB68IM0MJRJEY4d40EuSqtych1SARnET7Xvgj2q2q3uAzR0ZrG
DrlM63r6TKJrB4WUke5UpmpAPOuBEb/OgWMmUhuifO4fMMTlyVBkZ1kDa3SV
FTMhmjW5aB/jDUnya8DV3iXSuNgtjLJ4lyw4zDQaBm0S4HTFDDq31BgXF4Wa
8peF7RkUU1odVGZqxr6fqNR9ZwxaQMGTeEv9Bopfb2kGp2qsR17+31nK39nR
YQ+bRtYwsAKqBub1OUNwtbKxpIOfUZc3QwaPbgak8DZRg2gBbkvu26LeJ7WL
Krxv1QVm2v4Q1aHqEtl3eLXCOAej3LahmZ9SAhcfVuzbRj8TCHdVAWBL18hz
b401WmfZUEUnduQGWtLmYbvj+OkXMUAPPPQnc+oIPy3Plyv7pB+9kjG/W1o+
jyMcnvw85OB3WgcUEzc/eu6AWxBjJa4lyCWjeYdhQplmLS2QBGlB1v7pyKjZ
wIO+5TjOjKKO65nWoIRDlLM5aOZCBRlJXoeU4uWvipeKLZfcQqdzQNKhwt/M
LdmFRfou9GoXxom046E5yZ8A+cLmhvOK/tXvbFdQihNN5X6F5UoBUHvYJU5c
JMQiB3DBpG/WtbH7djTjYWSvvSkvWmP50LkLrD0JrJSMfJRe3EZ2exMFPRHk
xkIirB7aTKWkb1zMZSB4GV97gNw8gycwk+3AaacVJ0Rv8+oxVWKMuK50sg9V
xkTrZMUtpGraEo8LTvigX+ydyseghxngj8iptR2L+Jzy4MBHz/ZHafNUniL7
+NX9zNSte6fNhrkErgZIYKBVdAxZ+RyMOcIQgngXm7cTYYgMPFrQ+99+Wcu8
cDz0K/34ylbwTYRiszAMZN+KCTvA+sE/Yrx+QhRKAzavSqfhrpdn42Rpykc7
YR21uUSotV8qttLQcTMR7q98a0KUtYIBEKAMgBf4ccqSFI6vW40enr+fbkR6
MRjcmhS865P8EbUjFrVA682vutgR6KPwWHZPCxzPZaIfaEj7TlTfVXTn4K4E
P6f8H/A9wKRWE7WsCA7CdEZnneAAqHQ+irHlmpQ9z8zTc4gM+LtMEROuXO/n
D0myylpRynjX2gmbwYlrxg9uS2sTaaxyLEJg+O3mQEAROBEHVY9IDygV+mZ5
4faCVo4TP9FK7v+vPRARj5/aUssmUvN1CSrle+YVTDE+NuxlUo3Ydde8ZFOe
tep4NiU8B3tS6Yi6dBsB93KYLj2KoJCnTpaX4OGnydOgfqGVzlCBDCvtBN7C
56DoYrBBpjX5fNiEp0ddzZ5LZA/k4WAByd1+RndJQSnujhie4cXHRNWthDji
RE5Rerz8lbs6b0FIarJ7D9SgEwcITV+dUOgreDbCuiS/qE/b3JgsE3OQrv6z
UyYDBqFAYCcyA0ALJphCypshKqEXr4VkR3akd8v6/3aDykLkG2ijhB0LwQ2c
tMC1fJjcfGDOEfdFQpfHFpTAuEgNGZB9YLfkm8MjyeO+5vHdiV5touBtcbGN
8bYZlitjUTaM5WMJ4WlA7ex0tDiprWF5YgUIvCDxGo+PYiH4A3f7Hoonndtq
VFwvHyJoNsYZFUsUkbYoW4tZZWdYwqu1e8mMxLqzs6bN3wVpQwmMqugoUO/W
Unj0EA2gYMlHpez4G9Y6ufrmXU4Fk+9WKdNo7pZHRkUE12rCwF1IXbMHfDMr
orIwBSYI6kNd3Kei8atTpJTtlrAuUXIXU4+YRcDj1RgURjya78brTrKsUoC4
5Pz5NfQOspnm5dx8CpbpxSmQy2dnN8q5GQbVOGhFQjEWC+FFqtAKmWYjuplW
n1pGXVRd2+aUXqzpLZVPSMsqtxRAsW8LYj/usaKnzEhkS8l92hCbV76pq3Q5
RQ0m58pZvOSlHRCNY00Li32Dq9HCdbVrIOCRynQFdULv699PBVF1tqJS9HTV
Ju0oMA1N6T6YAfZu+wNUw2D7Pon8vWMeXAL258V3RsU5ivC4H/eh/VTl94zw
kfuCb6hwrR/QaNDau86oU9PSAm9C21/CjHicFz5m8Gc9fV5coPfjL+VsePGo
+t5PwY7D3VV4OxkJ5KDUuth2XyFncBiVoHl95uQopXXRVhFWWeNOTp3Nwqq1
l9dmlT93voChoCFly81T2yPX/el6F2RtKQj7KbVMiCweU7VIFFX3IHxzJ4Ao
4tOTcezaAwszxeK5q0VYNSq/r0EC3CtE9hI0qRlfqeQ/AlDXBsN2T+YGjkF9
wc+Buik7m0DEK67pKN3fzWKsA26OEp2NRQK6LQO8uLwJBqt10cfnPKqrhDie
IxDcipMpX6uBA/LbdjKpTU6sv6c86TwPsTyKdjeTQ1FQX3MyzvoOs2p9WAPW
d78yMkiYTElDpcJYcVROMq78A/DzVcHMez5xadLLs+0ZoW6d1nzugFDIoo/D
gc5v8TRpe4wjy6HhJLbAwZCa5H21l15+wheskpWP+OgC1a3OL6J5/X/C3rl5
ZtbVIaUD+x1UAcCxGwxnsW0gsPXDMvXv0YxlCW6hlNRr42PE10cfFwyXVMtM
5/6dsG6hSVkBSv1U/Wpz9BFx9L0YVZhz4qbcUbkbz82rPIKEbsH8X+51GmAL
GXKBsdQSNJkx55EEP0wYRSdQUeNNnCfveK4vlOpf3VfXunS79LQUIQx+ygGT
4Gdazstq9BxZpC9poGFoXsT0JqTSP2q9Uk/pR6oc4H2YSbAX3qe0X8JGUfxQ
JB7sSbc01bKyVmCqotxfIoY7VIqh7kqCGrv+V+zJyHlNvv0uoF7VoCyF8uvi
da1jHnY62qYq08XNKiH4nihZbSnZc9iEPb+PACT3tzZ+JB0gZX5uipn0b97q
ENhRhBjlY36IU0j2HxGwZ40ZzO11XxcX4o6/j8AFUUGiT2Hu7m/JfeyNyoxQ
vC1sROwZ1WQ28xzoOATLKBixhKmci5PxWhuoGw9us3IuVQaHPMTXEEAApNnH
N9Cp8iM+wxsRb9YAeg1l6BWCOSBcZwd2WUU/EObBfnRNgXpxteQ1I0rGk4rb
GhwvfxVTsAwRun0gvOIafbYQGFV16rH9sjM4uk2YaCUZOYhgdxWkym8sdvr5
P/jLcBHnPWI0LcxQu/jOfrkfReFPETpHYnYdniKiApib+Gy4jk+81BH2Cbzt
QxRKcY18elfVtVBK0hkQmyjxhnQaMxyK463RBdKVK318Nnxk6dZEVI2ux3QV
kvzn2gearkxPKJarhEJ744VhjRdLH1YsHp3ZBTnGHSEHOdB/2d5cPWPa346i
vmkrcGEP4tMoaoTKP/IJ4gJp2zcS/EsCPkK4QMzkQrivPbd8HHA26+K8+Qpk
jLPRG/sXNEUZ1PZnz1V0C1a9JjTDJFeCcODTCAFyJVycyI8ol2bTxwzRM7SE
jUxU87dGJV9kFWMNpncgPvHZDl9Gkb+M8wvlTalxlwelyB4/XDm2vz+lTnvq
AyRGZ0HZCHja5girG+JPcaVWDqPFZLS0CNy+QHqIyAuRB8pcbLljypERXvEu
T6mgBA6QdB2k8vXCDS8H0dvOV7MFpivK8EOWEP60MxoV3hAneQ+5nvFQ/YGK
B0k/8ik64SV2TeTz6o/B8RQfODi5A013epB4npIOAjQNb2xeuqrKY9vZEfin
SYJKH7ntSzaNAE5EVHO/Kpqq1qwfmOGs6MXDDdihlpxIlDImXxa7QzXhrY3a
XN94EDw6gykPU31rqzgWCotd/P04fBtvtpbO/AjesrtGy9J0+lDDc8zGrFeY
DU6G3yQ4hXpHf+keDLKUb2VBdeXqy8gJ4RlPUMF8aYdMwyzfRx0NTOL8KPPa
YOKETbbxrq/xvSuKse0vppw3Wq2GQTlr7dYIfrLaauNtNIrf/a3KxG48XMDW
u4SURn5cpk/q/EFkCSBRj13be9hyZeCvnx6gLp2lMyQ+XNq9/fWzcX5Sp/qa
RqSvqXwV/umA8KZPaNvtcHHNvWU0XB6iYHaKYKs1CDNHmF/7jEzzQHCM6jTH
lYz4RC9jZagNRnT7jjGrgvrNHNAAVDjdX5U4X5amOl98TyAy0Qp9K8nMMByH
cWUgmUZVqcsX0NVUkhestbwcc/u1KKw2OCbG/LkMNB3HO2BGqRAfkTbQbbBe
NQsTC3/rR+ULdoACGj75D1mTta6ONwqZovCaqxbPdT8yGSxlGLsLG7VDzjqa
XMKZjWOuX7MpjMSzmKfN1qCIauQKZaYI4hROG9QQneTsy2oeHYpbtyc3CNAc
DvwcUJaSSR3AKTpkaTFb6kghVm7HItyKr90dDsOvnEdK+7cX5DWW1NoLPW7T
gcazA4YuNCZILo+NTWcNbliY7BWkmSwinCtaYuP7UCHGllISP41KGU6jn8KZ
IoJCbEoA67SqbRMevI5xnm5aIwz9s2eEQ+ROdMpXZpX31V12uxiA0BNwdNyp
lFvaclPietM+y1JtP0oc+cHo+Jcnb0dxlDNaKHuRqeF+yMojhdgI40f1m47D
As0uNvsK4xzC2RCwZHrlq5ZJTocoOKK8TVO4kpcKUakZj2yECX241VHLiHMt
IPYzKcwQRbvMNhIY67uS9MerqFXakBLwoO+9Mr0r3imxJ5W0YIYFj5Py84FE
a1Vhh5CISShHxS2GaU/spFLXcMq6Q7gERUSwtmcUaiTYizZ7bJxuZpQsr2tz
K5dHqchuSfpZewUO7tJYYJWUVFoPJ4ynm/FlHGXYiQnfFwsRDzvfGUUsXj/d
YF3SKvfn2sBABqldVPwO2XDJO3ew+SnnoOTyGSMo7LQcWQFIAolHj8nSnYMH
V2ZGPE8yEKBpMV8O6Zew4R/A9vzFQF8DBAP5YcaNc1RYo7PhvMpYSmiNQyS7
xA+YmShimzHuXGonBRXlytW93M/2zIMph8GAF5sKFBD/IJX0ag8hxVErhQbE
rARYQrsIjmXHt75hgdhKZEw8cHh7r38LKn4YPlWcr1vilUu6nNYVXBuiD5Lk
yo0BdFLgq0Mzxoz8wzMdY09dXwiJBJorcxNa5w64SNGYFRMTEonqtuqtt+Gp
eQ+zfLiVHiUUBWQ1MnKDtJyUByJaCKsgEn5YE935VTAc6zS02u0xuD9DXUmb
zIxuQj7VY0RhNZLuqjfv3J3BfubZ5hDrZ1cGBwgt0IeSwDi2o6DGCddub+Zl
rE6ZZbmoMlYG+EW1EdwEVNXXq75St3K1M4UbYH6OpJKGGn+Nv0eZOV8x6h6g
poxk0ipGABW5OH5EPvwtzMiejJLRaRiDPegd1vJiOZ8oS0vvL5cljW8WzYi2
RVDa9uyK2eYBvTf6RhK0NS/0M8bl4+0/aqM0V9lUEAm1J0Twb7dQn6ce2erW
KnDstQwfvmM7rjiE96g0R539VuNo2L73jMZ0+dKVE2p9NQ/FMgR48F1Rs0Yz
ZvyD+uqgZ3EvE+XLWFHphSuUqR1110tX2QSFJ/KVZBKl0xkVdhxSwuu3xLHa
MciSmj+a0t2iGwKPcAKZNZbMwkI/nK78JyZGSy6WvrsPoW4A72YcQA3oy4dc
8egltjexnzld6jVxfyqRxNMnwbpiir8DSY9Bx2oy7I6xsgzr0IJuWzjDDYkm
b0+bLFrU2QlnZugSirYjcv14S6mPSjC3dwHuagDdPYepKWHxOZLkBmxN5jTZ
xgb8LqCrMpLD90Kx9wUoSF44DRGwgs6hx49AvFo9lu6pzUvv57rleVwB6UnD
0N3PaYcc9LYve/UhL6jB8sQNktNRHT0KfFe36ALyvGj1BA3aCNplr/OS8+IQ
k9pGTT/J8RdIZGAoNUs1zOUU0HJqgQoxqjwd1Zmkdqo7Xc42xhu1hIUOfUBJ
6wj0yknfjdHWst9NSv2qCLtEinN9fSUVkdI6DjFnhwU+Vm6xn2zRUCimHqNV
QtuUPOeEvtYJN2S34JO9TRSTsikpC5+gctNThPGJw5n/BsMkSL1iv3EJjsBa
Je3yYVToNRMycbQsWC1NW82ueo/dlGVJDXYkZiqYgSilPjTcTSiKz3KLO43Q
hn2uSCsjRzmooycKe5uqbq8h+lF54ZimOCCjzfQ4VKDCFGgRalSHhJ0HuQ7K
mWXGDFn14jS2s9s3CSJiT95QOQGrEQhmr+ALPwULeGF4Qq5XprPNIjcrn9cH
p4SbsAGXsF3NOqll4sJ2v80Q+hV8CJ/j2asy0m2jd9eYgY2dLBi8G84/pyZR
8wXLiLVHFrUjRvMqrdPN8ohdLxe4NKSgAoMhvpJoOQFmZ9lEKnwex8vN6pM1
eFTUwIfe+FKlo2IKh6YJVo6VR4AEHGgfs/J8vSLE+5qH6t2ZZE203yrr9ZwV
q6qmcv0+9KfJ5IJ0OBbCKbEsR6r4s38ILDipzuSqIpokWQRkit510B4n9G/z
9Lpd3fKj1QiXy2rMsqYwfBKPHqkQKfSQwWiNzRurznZsBZD7lYf/lSx4TOJg
Xgt63ktu+E4mMPq0e1Ty6jj+HbskguwHyhtfVpp8fnjDVOoQNt10uJPNil5r
WU6NzPzBEI+q46nSNZsLtFHrhpOGsMwT6lCiztyZ46PlCsLUvx5Tn0saFJdb
n3i3KlYMr1gO3cVvCpTZ29JuDRerGlgZW7pnt1cPEauAxEQhFWwqsup9jnnc
RC2pePsdg4lM0RNsBdPZur2ZjO38wY71sNA8czCbmOZ+gMfNWalt1ztaLOtz
ob9LhNyyCpm+0w/PWcPMybjj8S809KZ+9/l9Y3ACbRbdaZEgrEcJGsO6rEGy
yD4vE/wS5psLyIFI5OhFIwBGKDQk/xJ+dQn5I9tc3nMU7lWJYBHCJcWTklCI
QGiLPFxQrPyAaisvHSowk31KgaCiRrMY+0crT2LqtA8jxkyDwjDNRIc5fXeE
pv83KMO8PsOvi1ubPft7b9/9BTf/hr5J4r0qvQhyOUGSheh/wabkrfiwzqNo
94wAfePvZPckTWQdAqtC0cXW3DnPFUXV3XKMIDr2ezoRf+z+uFarZ3a/RXCg
uuLbB5JKStYoTU6ouigb5qYD/UIodOjRIc1C9PiviOyXh1kONhqthTI3zeoY
SLM2kAaE8/HKefhEqaYDkxN3mq371hQ1CA8f42nB8NdCMauYlqeyXUb2BDVO
mGhzBdypoBVDl+9kRaJhfnfnqMKTMpODwXSMq1xFyGbM8u/0sdIoZIICXlt9
RbkZ9CXC0kxP/vzzxaJgC2BIlaK0wWAt0K7KA0J+JgCYt4MyYrnzpoOn9g6g
uUmTAMQ59z9F4URWrAC2k6vE4TSn4avyBvWpAavu4wxZupnhf+lUu75HYDf4
U4xrVJg/RiUu+weZCbAY21fL7ib8Tyb+z5XJNhWdIkYn1JsSXinTWW1Ehhom
CKzajQoKqpZW3bMzOzVMPnBlyf9HrHjiyKe3OGQedgfNlWNwk/yfjVLaA7UQ
xEXRlctIP4pHDzBgsGLSGFc6XjHdU7zJwtxEI1HXUdg3+SGGv+YUQnX2Od+s
9gUHcIbGSMc6CJN/g9SilyYcR7mFo7dm82/0N52la8XJozlq51t2j3Gtbqnj
0Yn/lElnHW5nhqP+sFCh6ZsNmPmL0v8VNiE0Q1IB6g7JhEM/CZD3kpAiiuG/
DMRGBt0SVzh0pMHg7eWi7D1y1XjISPGEaKZUAdRM2XVIlt7SX3qGYyJiob2y
E4psnARk2hugytcoIqLEazXp3bO2G8y2ykMwsXlp0iZlxDLDanl6OE45XvC2
GWg3K/3HU4nba5WHqQy3KYgwKytaUMPcuerbJUJ9fjR6O7MUAWxXW2nZUEs1
sNoEpKOUYVLdEtBvvbSzsngYl/dOOyQbyTPjk8YR0VmmXO8piqeXNCS3H5+e
RbQv3i0uUGtp/QQBcgioodm25cwwUpo/kkFU0/APvdgnt6JUol6iukE7KthS
eRG2WYEO1KntY84xk6S5Q+0B+OYi8h/Y4vApm+KsCXR2wleo/FE3VIJKu1Ie
Hb4uL3PsjrY9EIAKQPj16LI+B78pQ8e+Bjujly+L8XUwKYAzUYcYKXpHnjjh
8jk/zRA9qfEaLhoE6PF6qyTzxH65Q9NOhEg900DZc6WwLyfRPygoLFSCQ/iP
533gFwcMZqY3VPO4seJJtR9R8+3BIsGK+6Vm0MF7nNejcdiHGqYb7axGXq6Q
sCXQ8ZBfomMzxmdz3CfSHcg4i6KWev2w6UxJWHRiIpQyYvE6Dph+/3J4twom
vsT9OxcyLHzLArL0o061A+a4FG+/de20w2P3teYR6GcP/s1w3L1f+UwzcOUX
Xr/zvyK0y+Z30EdpuADrGRFqYE2Nyb5oOytxbptFVTu27joE/auAN5DiDKE2
kBRh2dw4joVgmEjxy915Au570a+kl8Y56bVXYLU4AOXddsUXiXb+qCE/vlOW
jsM7CSsVB6EcV+8uzYxbu3751qnyI1ruEIoUL7RJfhAuqTx4N2+L8O42nYI6
4XTNIJw606MNor5AwGSl8uXT5sh868HnDkmGFl3yUqVTZ/Uab5UBgfn+cqxx
IE/hgANihoIhY2QbE2ZYlHJjz+7GKk5oEEfNbJPL5JI7G8y0Y5iLuPCM1BNb
Z84DFFB3Vk+7nXZsXzR91LuxCvX+DX+JnpeGWdF7KpEz4LM6Leu0J0x3ms63
nliRqjrAcYpdVp+wDQsQI8aSdlI+jMiIrGy7Hrh5RqCVwaYwLct9aujpqCUG
I1JLKGUCxf1vOTxPylXCbJxcWtn25+P2iN8Vib7OymoIUv/WUnnqqAyPITNz
fT6rrqoWSu85CQgslxrYszyhG8qMXUQ86IUSlLJ1pq/5DsfYnPejl/t3IQcM
Qr4SjzZl3MO80cxl55USbJLC/rpu+1oQpVOjyvNRnhZvpQJdhHdorscQdzeU
OGLX4ZdM63Dm1hhMClwhFDUkXnQfzuNnH0TLh5x4Zvh5s5fL/nsQ1hD0lJCp
zmeHoKrAwTKBVBeAG9hv5O/JlxhI4qlR3tUKah8uh06p7jeAPu5V0xGI/Ocr
QxyOosUDFBM/jD6hXjnqO2mH57T5DWJ3VSzyHX9Efm6/4cTKQEOOpjSHqqTi
iQyDm19WXg5RacvrTCym+yV3kLW09PAWqljBbnjPiBrdQC1pyrPACeyRxKGn
zpcdRFXZz2nwyNkabnWu2y2PqpRiZkoDr4QaViSW11jXKq0LcxdWefEnvvq+
XWlXkuGGK/J+LD0MNxR1OUi9sO5/4gk4FegwSjH1mtf9yrb7hpLNThpG6Sx4
Q2FZzrDw1DXZ3Yu6Z5jB+WXSaiPGU9PAkZoCs+iU8u4aLe4LtUlbYo3WH5zr
dGheNF1GDFmJbxSq2Sgfiw2tBaQkC63PBkfnRd0ZO9z8ccNJBdFboXOcYlBy
bKVJ2QoRolopxSpiKX5hlbIa306KhozZwXtLwFVaQZtpmDUr7HpmoQ7+7SvJ
TVKqTWEeENsJ3dJhZfj+PPXIN8RNv+cosKrUuM0SaBPwyDp/AYN2OXYoyGEA
DHuibHG94J11US+DmiPpyejXaf8I4FxWfwsmuxExZmdXS0q3aqDxKGI+SHoi
1ofUcrqDRZj2bOhNHfWNHcJiUGCvla+pCtL8Yu1QehwSDBCOeDJvnwbyrBxj
daSVq7fB0mNMd/Vv82hu7ESVrUrrAH/dhsH1wPEnQXycY8+/OO5yQArr7HKw
JXJqw5j3BxA9yCVywCF4Xh3K30S52vWk0VhYEGa0ak7pD9RfYxCcFORUlLU4
tPpo9ddNmQvAnkJsg22sblOl61OXGN4M90mQzUYa8Z1CHiloJTRCV75rdo9K
p92YWt3GtbBr4y7H4725Mwpg7N0+z+vFyIxIyIw0oFSl6gvnJYFVJ+eJ9HvH
kWuCF/W5+Pvv2+/D8ks3YXGBSk7BOCrc+oo3QsSnGG3vBYT5AJV05cmO4FS5
svPOsmuOWGUiEAUU6k04avFs31WWANa4QO2JRiH7vdwiA9m89/usDfflFvCV
cBfVufC6rcpyILkdf0RzfT/sus8lqbE2h2oNARsKPc4JlJ0tJuXn/OnwvF6g
fsLYTBdEWQVATYbdhiAGSnZTiJOqOnez2HeSXVwNh3bcrBoO5TJFUyuvkDox
5F5t1Mn5eI9qvwFsqK7gzF2fuZyJRU0/ksiwFFUlpzvAtH5l+1XYTgpxYX2c
+rZOVb9O2aYKRSvrzdc/Z6JorWu5HYmFGI/HPz3ooXbA7gadX/TrpcaULY76
jI7A1ZuWo3sChH8yGgqtKbINsS0KlhcSDvu+HlOgVM7ZTus2SOgs3/+UOrs8
jwmSydtKvQ2xPw4VEFB5q88/z3grQw9HbF4ZdOOnC9BnZLJBUTdbIIXAJqpk
oIWvJX/gPUrzQVIfrnvfSOQWGnLQvRnuAfUOOhAS3RVwobEaTZKJjBwUc/uZ
Vo2fxrEgrVLmMNgaQoP+Ld4himIL7a4Z+SgClT2q0MsyyMZeWpSjEOs+xFQJ
kkiKDS7cZl4cRjv5IkjKO1O3bQLZpFO1qVKvg3DVvAilxStjXHU1wQkAK3J2
Owf1lwlqSlRa9jSjv/oj1YQWbigR0BImu5l7fNBXgaYU7JpOqw5kX+D3inCH
rOU8mlY4bToTVEg2cnJuXUa48fWbhAho8SiIzLF1hDOyPLQC63peSFaKvCFj
bR1/IFGycdEo8dtG7ZbabcZ8eXaRnyNqZKorjNGZshvGbytcuitR6of732jn
Nu1uXG9jPkNq7xIz8ji8rL+NOIE39I2ZDn2yzHZ8xjdrgCmhGeq2gLI4je2C
FyilLD1jXAvbo9U95TcyFSQbWyYsMz4BtKcpIicvAyMzbixLCZ/r8zRBDAs5
zOdqOqENRRXYi23wTiM+cRrbMhWYfpPo0p0YgX8LwWM5EV+dQN79EY1EblpX
HctBCowgjVy1NqkwfVkCb3pSVuhOQ0DON3IZVJuYtDX8uwGFZbtw3d0Enrwc
42UOHXScZN+v7hezxG42UXnbW4rBSIvaJYSYsZhDtzWH+DghQdr6thQsG+nO
lb63MXH7/gI1x9/5tajznXei4rEc+u6BPX4UHntq7J1YEf1tP3UF2csj7sVf
SzkxNAm6oTW8SjB9BSGeuimD16OXJgp8wwMrzlz2Sup4KxPW1M/jACc3rd55
5YSXjLA88QyLF0lDSdLxPBwWng2cftAx21AqrobO9vMScZjIKDaw2n+mRKZH
yIpZQ95r9RRv3ZbupChF9Kfqk5tk4uFM3RNvGhN2xRIL99Uy4oYohELGOMUw
Ha8bTcoju2moZkLeopcuCPJz3qp1ksl6Wef+h8pKmsZ0ZnZOnckgXbzH3irm
+MY3mCR7b6RjvCwctzyCUIgMuLdVb7m7f6uc7M6vnabdPUMaz71BtX69uj8m
UHyeew6rsqLIDGaI57cCSFsqMzqd17qI9+iYaLECoe6HxOUx4PQG+jtzvY63
e/gLHa9pYja+rw1ULCkyt6cdPDTYMda7EdfNsmGoY3ImsQODrgLSCMMc1ywn
Sn33RTupRtc4XnfER+nUxPDhl05YfF4g2Oktvsw3V+GTMt10+zjQ8A5KlV2c
2dfc5cuH4ARfq14IhfFyIQD5hUhGBLlF+jzIP4GQRi2k3u/A0xzAq2dhmaYU
mF9Y4QfWVA9eNwLHH7FGkNpms/PXibgWHQDL4AU5/PmC9t0mNafWVmNId2Wo
b16ejvArGjFJVRcOezRXvNBsci6dRGR9f8UkiR3WEqNrOq93zDYS3kFQa/md
KtL6vbhMB6fTqLFJwJ+SNoq3gs0BXIaTv8vSlNXSiw23VWMAadIFFPMgGtaO
JUbFeMb8Lgt1bbVo95ucXdf8CONWAzo0cibeLzs46oZKYq2UtNWvukYsb/88
xVtnTpBmvsRFffIbyQn3hwlG0QMLF2+bTRGs/g9+KqydHWN72q7mZbty31Is
HE6PPXfY4iI0TynzrFGn/VuTIYmGm2SdDYZyGqrmepJZ05KURUi+7/F4YXiR
ZOMeqOQvydfXhWziGiEYeaK8TFk9P7WMj7xTWaymeDE7bd9AoHTFSY+LeK/9
KgP3oVDewtz1LJevVjP1ZBc0xnrRei4KW8CXNIXyOtcnMDAUlsXCGO1yYpEM
w2hCFcJqpZkL11oTLA6DkNCcE0uBSZSnrwfgUviEeXmIst+zKBTbRAaHQGJl
YDNLi9SYmA1h8iPruKzvnt7b+D19IGYBaA9OepT4qK7kBHhg023qDQ5hvy5z
jUxiBohmyjoGp/ejqdGFa9uPNGCLgbEQjftA8pL3K1A3rmMeAnc0873G5KcY
MGxhhjDvrTm4hQcRG9sQevbbuOcFUHhRMJKqRXgbSx0UL+D88AU4q0n7oHe7
2ZrVCOPmso/IQTyewelV73AGCv7xh4Z3IYfSLgaPz73TlVYq3fE3JuV3HVUK
B5LwIusWXRcYpfPf75S/Q8QLg6AfrTDd8TW50B0Rh515X+Fj3+1W9isuP00U
7jE9xbNiDSVfqNtEMfc0tc4DE7libWxkv1d++FfXBa2aK5uYiWVK7v2F+hRj
cZEPmwOng86J21J8oUGKwq/pw6/WY2RrCPX4UufuWALAI0MxnNVnkNbzpGkW
73yXR5JfT3TgfFE5cW4DNLtZGlq/+nSV08jOaVBYvQM28V+f0Bm4Wlb9wSi8
mSKxqQ15TWvoZd/YScxJmHDVNp1FeyPT571//G2qTkVpgoTrdSyvzJ/W0nI9
T+HQIi/hqnKZNKXBTO1tRSHjf3FXQopRXgCY2K7KPRX842StQfOJuUbkpOwP
8YBeqxAA8ESnqL0TIceHHdeJBWujjanzKJJf3FJJnK3GvG6WFbgjl8yliuyB
CpLC3Sw2Ik9Vf9Ge4om6ueduPsqQ+gAcs6ntbDf2HslzLtG95MgQn5xaIwzN
NGftGm+/0go5PcLK6uZl0WJoBwvl9nL0T9duO+8yWgMOLzA6YGsEsWH4OmX3
LD1bB5zeag/aIQbg9q/q8YiOeNsYxEcz1QF4x4F99ASrPUDsIQAKsKNrUhNq
ygHNXVwv4sETlmxCavu8SMJdTGvw8LJ/vyUm6svM8ZfKrHyN0vb1Uz88E7+M
PkWR6LPO4Dp4hX3wKG8+fcEik/xiwWJrp1qrY/uFQ+9frmMf4t1/DpQ6Wfn4
7sehZfAnbhStpFsk97/3TPTrMRY06KM0zpmlOp7+B2njr1Al3tWvsMUg9bbx
qUb0NsWNu08R3qgrUu48x84chCR1/hRk0rFoeZ6ymN3mSu2ft/q2iTmwZr1Z
SNpTQJ7uRaybQXoFx9oKWbrAPx9HocVZd7IQnnP8QRrhHd6+B6VkbdluDrW/
wTak2SOeUcLKvtqkbx7RJH1u9D8A2ZaoAuVUZx8FTDZsmG8s8K52Wl4s1B0B
X436ibrhQEr2vCEUTo+hPwxjdcHWCYnMqbGm4zdrnQ3ED0YEGTm/d/wyu/u3
EaYNrKEKTZ+0ubI+zLM5+4aozSpxM8R856PBmz/fxEsfn1PlDTrHEeYPvHlI
/lnRQzoAwe4tDwVTu3+Q4a/zR6VRYnJ59wQANoUFQX69eiqvFMNwWsexsDX4
Bh2VlY9H22esrZAcb2QnCoCcuUs5qfg+trfy46LygRUxjR4nCvHQzb5391G1
1t/XA7FTBEA4zgqfX9J3pqMos6BMh/7buIwRb3VCWwWYd+/0TrqKmbZjD37e
XiyC3BWvIR3rIbl7TnYeRfWIHOZoEi3dd003hRATzDDSIq/Nj2mAcRUFCwN0
L76VLwocGNyhWjzZWsE/CP9kodIHiR6og02+e0K2Ck4bFBlwA9T0iBvqAdJW
b+ppxRWfi2MVBPn2o4nG5aAKMWYgLj3CEcc8pDrW4E+Y16KTthGs+X3IIYR/
7ypQG4w3Bb/nXathi5bi3sHN9i3OGuS9RHUcosxhYWVojaG25Fo6rNA1TYJ4
UIwnQj6rVp98glffHrx0l3DZSSwPhhOm1ZQ178bDw29Fg1BqAg9fyiwyds6R
c79asEm/IMS2PmxoPL3HValWELyqVE56f3utpWWKJPTSGIsjs5+XKj+23tsP
dpubIJPOe14yPjX03qUoJuWPaK0H4za3HrK+SLFaqiLZSWf/7epvv9l+B72V
YB5QzArfuWH6Lr0SRNCHBqWwGgdEDYiNgmzrmzk3O0szvV15zLWfRXcadBHV
mAQRtoo5H6VLDSnhVKjAQ4t0ejlZo2P38burP3P/LoRQBiqvw7xbebEEUr9Z
9uD7uQNghz7dHvqiEiJ5+2dyVyhDLyiGcybQW553JF6vq9HjHRIgEr77NexN
21N+q5BMFuIs0oim6+y8gSzxs2bpw9b95GqJ0tfhRW5qw32ZFqHcb7iQDiin
nK+IoRkOccDaKv3gnv/OVeLf/ueUIl5SZvuEgu5rnaX/F/XBBAqX9hf77YCd
Cp00rfuKpy8NV+bnTzIV4aOBhOo0OJDK47Azs39qOUCvvtwTZ5/SWk5nF03w
T7zhtlh5PoxocKU264blWOX16SlZrh6N+ByKNeK3gjCCqn1hyMolBxlKCS+l
UBKJtLHntFwry/zWk1Xz/rQ0HvlbyGFAVvFdBJEPb9isE/Bui9AtFNzAi6pQ
A098IDwe5VwrccqznMJV+gYxhuqJL2rlyNA+ScG3JnPfVRgZeXF4B8DJax+X
Gxxg2G+hxJMzbbjONlHXveu3qGfBtAEYh9CbGISD8FKoiNVzG+6IlCZo/1q3
TYhDhQKHAffdwo28obnLb+CiUxRBAe5/USo34a5CxsUsgRHo4UkKteseY4KF
RF0cIFkzFqL2wn/lwIuKjWrat4TpUZUT6k0uKrqF+b8WF+2hGvnz7o21QDhX
R07sWF4i8lOE+LJAqpRoKTwCyhKszjRWaf6JnMG9Qqa2gzH8PF4mSGPSOdhx
SREVo2Xrx9KTV0Qyv5reVLjhjQIe+JFgY9I08LsRdfopSRvG0XI23MOlOthD
ODAZfQtDLd5rd9/cUeSJKH5qQDoIxpWPDDluAjKUPmPURFqYiPYYrS6lgbep
27oKHqS7O/+vwblH1zZjuBXrsQRa6Tkt2j2OPkQJkDjQOOmcGb125YMdWEo3
TQOTlhKr6taW571njjtyF5JxCOc/VwsZeMHbefFqwN5+lHFF/mBJq8miMW6y
aqkqeSDQT6beCnpz/I7uAuCNzCk1n1fKQ9bafuDXo2dxKn+an39UdwCK7PYq
StfdoluU955SxRstD8DNfNSIlSClkLhQ2WqzfMS6GaKDYHA7bPkTsk3kYLc6
VUBnVIMih+Y9+y0I7k4ZIeT2omb7GRz8YzGe3igm7/lpRH96JaBx1RM7TWvs
a/Ck114xMdf81WBepZWChSWe5EWSmtZFivgupLkbVBBvkzEzKNi6Hd4jH5iz
HTmwrkPM6LZbA2uFXjRQxXr6aeY/+NYkiF7r6WWInY1zRWOYwblIW+1FBwKm
GbQ3SAVGKiyywFEvX47R5DN2hBlVkMwd/HeQnszOZI28DbyOxQ5eO+5AHLyg
p6AmBfKknhdVRISNd65qKIHdBP4U46mD1zO16kTTowrQKIPrzSZokjrxpzev
VCU5ICrmJMiDupHSYeLJk70G8FlLeFUHPKuv2NOeB2SongWSKG8WTVy854g4
k91JHu0WCKlBIZdW5MAy3L7AcIu33+wrWU1KfZeripKxIxdEv5AZPknfrXVA
FRqMkeHuWdCn/ScdoYtqQ0Gqozoidmq8/il7Eq2OSkWC01O3MMef7Kj8hZ1B
VCFpZPDagDTJYPCo1GVW+4KHI4sqcyLqjjzkaKeXjvUQcwEqexxNfWT2qjTV
uksHgT8ubYAOieIuXdoK2DbQqPvemppl8imsWIjiKVSn0M3qrjJXNVqBQDRd
nmNtb/bPuqVWYTQO20he2VSM6MR+U1vhyC3OkmFl+64s3B2No2ubwj4/0Syj
sHfOmpefn1vapLw5r0mX8uptjZxSCV3g5oJF74O/yrit2E2LTr6PmTuocAJq
qND2EKP2PkPtE4ShVnnuffYlK7RRQyJJCtpJFE+zp8Pf54qx+LmfkNDKkf9N
Wo9V380ZneT8f/g0+m9XcvlVWdxdmktwsz0QeKfWWpoEr7JMHo2Paj4Suslj
fnNUcSdzGMOFNPsUG9jM1aeIkY9LqY/F5Y1iw4rL051uyt6190pyxyG4drbX
hZACnVLZxjpn0qSqiN1u0w36oycwac7k6qCd2dC9sZW+J4OceB5pz9dmJO/y
DM7imltBT8a2+NYY8GDu91pPNlI9gIQzXbKDIQg7KCvehJVd0S82BzoeDbG6
wVtTs76LRazdQCgOmQ0jdSo3+iQalbl8QaHej67c1TwvDEiJUXuEmjHxP3Tl
1HHl65fCu+B/43L4qBcz5ux7phIEMY8D/4w77fDiGSykKLUHXAXpfOYi2HLN
zxZ/y6kfIkKPc2yrzuMaz0HQkGQ1uwAqleB/yY6Gnj4eyaR0pm1yto3qrud5
BVV3PFFcnNOh+H1Nr0KF08Kxt+kmo1zbA0z3eYG2D1llxMyPXambtxqa66DJ
gJGc59dr17TCOCl1UQRCSq56MbgI4DwxoEPzebiR5BZ9F8YA9UMhxbjQ7pN5
bAqFQSIos1CNO+k9mEdYERpYmDK/Lz9QXhGsdGVPRSpARIOgyC99ePa+GCqw
DK/L5YamnlMqhi2obs5mQLEAk0D4N0jAurrkH1sY/O4leO8oxzGMLHBnltsP
rro1GridFJ6bxRqGCeqo2vBI4l+xtfuUggY544KFAb4/ajM94q7Hw3reZ88G
Mvdzbc6VNZgwIPn45DzPGFU/qX7e0nQJHqyY1Ay1+dHD3cJ30970W5wFwgt2
YiyTJx+WlaSMzVs3+trwHIgSTal/ptkCLDdjuBozU0IYkweW8JxESGmnaTi3
yK9AIVR18xitwHFqu9OyMZbmmpdczdcKiZFmIXSTKpDv6WDL0aLGo+YnXe7B
uANv80OytwilMa+WB0XbwBBol8qncP5peOsef2owX0uHYSxeXrQlsKlh4pzB
yLSDt+U+qlHBCAlWJaiuKV5PE6K1VPgK7HGyfijQSAIUN/ZjJ+zfXtT16VpG
YtHawwhmHB3Ugw7OBcQwqGuKXq+tyMO0hB92mXL/7lnb9HGo4fT32mpXB/DV
kfGejCYkjY3DrMKTuNIyEIc/1F2fx7+PAH/1+KeyPO8wVvtg+DyAz54wy3RC
7Kfl99JLOTWmg4uVqFUrTYZMyjt03HoXPmL4pO/84KelenX3BVLHoGsLlCcE
itXpvGk+n9bH/ydAeHUjxqWVqUqvI8TqI/x137jBA6c9amURyy6/+lcx2v8X
MuMYBO5EKKrLKHzSWIaU/999OmAyE/h23fA3m1aKynxDEnPLyogGIeyjEWwN
uii6fVllqg5TvU/oeZJoks94u53GiAqA6YAEOTLthoKp7UjI9zLXhagU4KX0
cvIgoBNgy+H+5Zjci1y7jrNjZwZKvxgfKvUjxXCCdMDie/57r04JbZnhMOTX
7geBkTJYkZjylxqwzkaNgbXjjruRg3cJ++6Sk+JJmiYSZNYXzrJHL7LIhLab
qABk1PjS5efqP788VZvVJtNGDV0XrTaYDoiE16pxxdpGMZKrecfn0iAGr8HN
O+Zbr1XyNia4q4lQe6iQngevm3TwxpGzyQKWdentL+jbzPuf3kxa/ddJIxoA
PVWQXh8Mq02FFHVaLcyk24RKSCtw51xyP+1VwwCQhtqproqFRdt0gBhyim0y
SQ1r2MPdb2VikQ624lxBsVQ+ENrWsRCHOISHb3ArrsnXUL1E0pu9I2ZxLINx
+2vQt8SaIu3Jh+Y7Jvtpv5l7tFl58RKYoaOp4MtvdP/P4hAEMEihZguezayB
Q+xcR8Xn3gcNLxyGOEjvMAI4oi/4jPAPx9f3fGpe7YghZkPHB88RJM6zmRKu
qjk5cM9xNUnpMUsODpp1Id1Y4p8zVuk5pEh3q+6tJMYaNmk7LAZwWHPtVuZQ
pDRyk4nyjEfvMkE/MJ5UpyM9ucmWDqgcoifwVUBGR2LENB5nzDcOuzwrEaFA
S7NIowcizWqqaWTOYKy4MmN3tVnWIXYM5Ta5/frS7uxiXrEGP+SiDQnwel30
a1r5RqOu4OCNHZy+j5hgUiRG+oM0IYwPLWZhQRrWKI0Ic6v8XfgXsZIBe0zi
DprUL53HFzi+Q7zj0HW6c8DB/+FQaFCFtotDCMVBSrk/ghGlZXGu5PLPBGM/
+7Rbtykuj4V7y0SAhlEVcn41ZlOyvavlx8/PuMzBAqcJQm7hd+LiWLgHtAlM
eHHP6qaNboFILFgIz4ltEWFrVGUQoHa43nfQY1fjJEjC+8WUdQhvI4uSSio4
gbvW7cuoNq0saldC23VR2QJzhqzbBDMF1zx6lO8GzmoctHl4Miz98C6c3m/i
qbKO1I6dyOjicHteVfaVN/Y99blSztnAPGkSxLPIux+UKI+kd0jFLvc7c3Uf
r6FFgy4HuyRrdWlwB33X3ykRzDhws+jlfsTtZKgN3nUKAWwa9pWUnsGS/K3m
FSD5qU3ohCA6KuxbHlDOMlYdxnh692jW50v84W2lSGm2q4RULxwbAArZ6Yl/
tMPxh2SEXKOtSK6PKQ3ovMaaeyr7FH6Ynng5hZeXZbknyMg0AURjDgA2HIiu
GfiJz5ve+odDIeutGgeZMB6zCtuhAtyXl1rfy8MsChuGpJ8NsZ6j1Bt12HXI
n+otS7o9AH1KsJMSQlpzqbgJRrQVeh+1YH5L/ipV9AQVRacOjcRSLrSLHcwO
wVx+khODf64efcYuW5JZGfH/UbTXOMTtzt5jtRmhDKHM28fiKqgIW+Ns8WHI
Us0B+++BBRAu5QjdTUk19356ef3BQMwLKXy7BKTa9MoFdwu/99cXD2IdFfsq
swQ9XH7GDp1ldnWo9jQTmoxxMtUUDpj6Lts/Dla2O9ALCEVct1/k9WrUzLRQ
G+f26omz08sBS+oenwNBZaYj4RmE/fGauXbWeYkx2ELl8idXed8pGqQ0yzXJ
fB3mljCKJRbfyDOlKZ82rnBvODVpFS+Z0pRepxYQKHyefDAqk4dfd8/z+4S+
+FMKSBUEhEOs9yya1mbYk70QfIowwCOa675rtcr2TCBFzjQUXQU7u5X2b5/5
5+4tWkw0byCQxyLss9X6gFR4XAYccJJIkMDSTVKFW1+iIyqvtWo+CWyfRp+v
PElJR2t1v7i1L/zhaANoOIU0dliAOTrzY+Zli+KZXGYR0xBxNAdTwhgCRyTx
Z5obeLyZBBxBBVhaeRCxuIT1s29bwXtxdZP/yR9LgDE3202STlqi4LQuL7Tv
ziathgy/hj5vqNCdbldvBoLA2qXNohcb6UFDRLyCERBeuJ1nHHNUBZpuO5RC
AXW6HUUYCHAJ/FMGcHVWyPkdLU4WSYtkE3PUCAXLBHHdFthXIp7TYMCSkBLn
b5QDa5AGIpzVdPh+3qlGrXQ8eP51BCOUEIvcN03duZVVwng/Iefl62Ry+Rpf
FS3jwvkUCSA1rlHHuAm9ivL9a69Ys0RMB7bgaAJceJA486/aPFwxnEHkfVK4
e3eTeyYA3XOMTq5yXdMxSE+IOflRXhT4rk78K4ueUA5ALQvZBbuaYIyBTnGl
bI4/4wiw3+v3WiQhvgIS6mCV2DlqTlwYxQCmRT7gJI4o+ZUC355fLcps8N80
PhoqTUuAwXDJvXGQlKiO1PFPKUtMIiCt/yN+p81ZI33R39Jqje8aByx42m0D
WUhrDpEQNzfWlUl6LWVD5F1xepEGOpvHYKJLBTwe4wvnsK6d/TG2HQURq7UJ
LtZELlAcMFlSUsKi6yJ59ZfXssutGQiZRKJ3kIQZoZZU5buHD7uY1wivOr6i
8R5EY5dHshJRcx1160Zy9HmwMRAc1EWFdA9nu0kWaeI7ZzSrYmWUEs6yN+Eu
z+BzQTOFH3eM7eBuLjYsWAPneAnaLpbHVRX2Aa9oi8NImPnoxdzmNivuWQoF
a9JR0USOyIv+gGeZ5rWap8lQmLljubePwNlt7Rdr/dF+AtQ97EDQjinL7jty
1cwvv4ssj664xSbc4o2ZPQtwcWOn9KedSCTVvO3DnkfAoT1jOd7ldG3uikxp
yfICwlmjRirtiz4l2vhqYkfK+Hk/dPgtXZ0oAnIlqfTt/W6CqGbSl76aQiO0
4ndLamJY7eXz08D0eNujDNLXSdac1IA9wyTGcHc0GQdDg9jN6+ogMgO7+ZgD
aJujdZi6uFzMi3GJOiCccQniV061v6kBJYuEuVQ8xinsB6PFXZb7Ze6Wwl5s
3O2FuHNULNLVr3Cm1DmA0Vk0TguCh0BA1KyOJaqtU1rNd+9AEqgHd0KVLJmB
DbsNAPqEsGvUU2cExOGlEhzdQ4lNvBvWS0xHWxxNKrPSUl2CCmPTSdgJBtzs
oTHwDGZrCd74vnj67ywb3D5FEu2ZSqr9I7blq1Nd1HL+nlAqAnw4vlCSCMgz
EtodNCbAB+4hDAHv1FDAaUe064RHUwiTYtGLJOI3jLAHvO6wl47wEpniiOLP
0o2QrR3GyLgWCYokEhbdXL6U7y1f5Xf0WvpYIvAKj/NvjwYy3ISlmnsc0QKe
KRxVhPdJK2PEwbCLDEsHa+1p6z4WHPD6Akp7XsdrBIBhAt5R1G0U+L2Zdut3
1VIIPLJG61ey4hUJkqpnJcylCg0aFbMZ14RSKvkzJs/QmlkIJB2IRTdujYPs
P87t5RYbfRxBjvwK0Q+el5sdYlB23792oOORbmj08qbcUjy0gixNzyozztR8
NM7X5alO4Kk7mtf8zv4Cza8+J/eI0A3zkQ2M/wzINsbfnN5+9klak/3VSj+n
epHCsWC8VjEskRchrdFEfNHuOJVyyqlpBibyWyRsu+yviRnfNIIizLzv8AiT
dJ2g+hEM/uv0mbDccs5r6qnTTDh0+WemQDuB35nqKg+lh5tftQS21EYcf6eQ
mQKe9kMF3XxThNALbyR+1HL2raRMd8BmbfY67m585+k9PRLDnjSRQ9ar7JPN
dxvSVVOysjuNwSrzkBgL+pHtq38F9ZPaLgLkwlEDscNhw61txydYTfdtwZhR
c5Dz4wdbqx1/cW9pPWWBjBi/eXnVgKZnXCz1LLV81K5O6mG/4ayN3gb878H5
gNRRw6d+wOHysjgv6qWyePmqUDARZlnG8AgNYmlD6G9VD20kkUw8NLnq9pvc
5aUEAXBovvbhiUJfxDav9t4OUEB6FMm8xZRi50bHzDUAL17jUBEY9/CnQc1m
L2Uja4XOsR4uD3+w3CK298piIKjjO0aEBoKSrcubcXDIdiF182orDbuZeosZ
wKQOMr50OWxxGYSPFUX9ezk/TA4Lrr5+AYfcRB2LFlJyVgtc2rdJjZuOn1Q2
0dLZekJ/BJiB/mGVgz88wYdAovzt2xtVSrdoMm/AmOO6f5aauM01LLjD65iK
7oxo4GdHpvLi5cSFprOxczdTT3AbdM9Lb8bo7S8LuFUJZNnSWO/RXZgg0Ajl
hQqmfK1oAK5sHcAymRk/9Qy4CUBgksMC+sYqNpN3d72ZwV/1NPlcI1ed1gCd
ESCd/kweArdwGbH47ByInxwl0zkPH0ljGlLldNPRlzShgVOXuzYf/8eqQSJX
Tdej6TVjiNUbzreDMog99FKKwWZ8IIBD0KZ5gNxlWgCvlgJi/lcKobWkzX+L
3JQv5h1p82zmayMjXR2hNakNbatgljV8aBbx5n0mCWMpUCIO4m09HZaJmcSv
bkX3IOx23RpdUlo+JX/vQceQJR76tKXx/tl6ST1LbcJ3/kXXyGqy6BGT/b1t
jjx/5/BE7zEtefaDyF8ep+Ba2e3XxwT9yi8K00xRJSE8kK9UlmBvuHTow0p2
sVuDROgOGNfzci1bTQBBfzggjnE0H3m7s3vYZe/tXtOHdbtTX90OlbEkbmfR
wrTDN8TuBqdZ5dkTZEhqi1/la8PDQKp8q3r5KWYi7wWwZDmc1hFw37xEEtRk
z1iw29/ddqYcI7PsxU/+ylYesmBa5QshdaJWBFsADINCklnBWwB0ORnZENA2
Jaagfd5bJBe2M+zb3pw9IJG8M84iPNmGeuCDhD9JLRqys2QdOl4lBSl75Xzh
oWcB5GdIcxdm5lNkpvquJC330BbsHzn9XpKvxokdN0aboxRZ/wIfWe6swO+t
50W6yhVGMsIKJD/rHWJnfxpLo8c6eYezdzv0ebVHaisYIa4gxdeOHOApzzpl
mLT01abvKrHm24nMjq4q2+EDV6autydYdCmGn5xN1zaP2YX/DYvcLAJx/Lpo
4I+FYgi7ECde+Oy+WIpUW43H6mbsXIFXftbzZ6j1n2Y4UeC7s/nvDWEKYhU0
JO//Zj0E/2cBLYYCGWxN+srE2F1kB4sGssyT+aCDAl3cNQp+FT3eDggZe7zr
7sdNynr5UDtG4vzvuTtR4juIX9IcVg8EK5+ZL4S9sVe4qjmuKdXv69YzdgsB
9Rc4gJgKi3vlCyvgIT4fHmNiSMZUEClqWdUppt4eHifmr3JogGGWKkVf0cqr
FlHSD5JIBxwPnBcEpMVikIVCzIQjfBPdxW6mM/TwdYq4L5nBfVLb15jYG5Cj
90oD2fBIbsY9U+2WBBZ08Ojv1YvqkVLzhMGGJTu4WEYiZp4JiRYg4xMW9F+e
hEydeKXh25w7Ybv2OscYpI9BK6blJNouNWTZsnr9Q03UiwC6wKh/Ojr+QeLp
+CgGJSCFgSVVrx3ekQK8JDYti7nTnKHkloTwhSI6Yrr43JunR1aGux/ZdjwJ
fbRNSdtbvjIch3+Z8756Yn4uyBdnCpvjW2LbJ2vbABIAFTQYhp/k66aEGvAA
E9rmsocstHpiP/K01iGddbZOQDUBI52bRM3fZddNRkmmdqOLSlD2eFz1ZwAd
7uwxlvHraJy9QvQO03+yVmhyTxJ4YqjNYuJT8UBx6oTVxZNJI4l09U6F40VF
6LClnCYLIVR29QHv0bprt/zVo9oEhUPIlFb8xA2Id2HELKraLmRbRfkhukp/
j7PqewYYcgZZ0Odt1cbsmhGFjU8QAlNoYAHJa+/iWtOR8rqLoQu/nBxwA2N/
7Cs81qhjFSub7v3pcugWZOst3jwxDti/d5rvTy2agTElvAGuSSEQ9t/66xPR
SZUfPMyF8fn4+t11BUf9OQpy1E0zad8Z9YmLRSNBi3mEZfqZ69whAKos4r3A
/0wBE+dx9mRaYyhjjPg1ub78t98yPXzeZv88E4oSEmFdTYiWlgQFQdHi69RU
EBQw/1jExvfitTfVLlo3g0HopLakn8pMQrXUsh9kTcGFSnjM6w1DWuNQ8sLU
j6wpPN70OuxaA3jvhoiveeM6eNK4LuNL/sE+Req+fp6LGYPl23qptaA/4N9T
OgXZnJb4rWV8Usa2dKn29bdwnWHuxmebBb0f2rbGHS1nzJi1Kxl2LX+gzJRc
vwct6o4MdkwhH/5ItOh4KaW9qVdUqkXbJgGsqLL6FmQuqbwhuZ/0x8/UmUqV
AIz2LzseLbq9HwRmKEumKWzHxBvlqp5NY862nmVoEaW/POWbUNCwstZJXctP
25VaNnFyfOkRG1y81wt05M+2EhVRRsQiq/wUK5UXNRpJoGoJIAdpUv/5G87U
f/E69DQQXmeDyRDuC+vcW39T33By9EXpuMacD9QCmYYW54CaUKIgWhyDEJLd
fHiuMMZVu70eVUJbpL1KGD4J/ZDc8KRMOWY76S0QUume2fghFbohEub5UIsw
bC8wEXfN3ALi9ms3dn+yRzfFlhKJ+cvvmmQn38zRzWIdv/FSY+qF4FuwVap6
DUkxGnbDegjusBpK9JpwjCzdxmcpMiobtYRC/T5pyRBZXCO+SZGVOTXNluB1
Z8NH2YA55sw/og1e/nYX1SrsjFli1zfxoQAKbQXJF/uXRAWCUCcqJZLLr9gm
BZ1u9vlcU+VEUNK2HwH+d4nsBz9qINNSiaOtk1yg4VrRb9kI9kvQiKth0MJq
1o3z81PC7EQLdiLiShDVX2OXwjuSyTKOd26SCzNoMOrhl+ekT3L7yIRk0dBy
EdnSWGzetEI2pc7vr3NksDQptRd2RMkT7wjXgdAi1c/sP8VMb+oabHf9cgGu
EJ4xIqa2nj1aM59tYRCavjM+/3Fth9tnf/HOjouzpbNKd3vc6U/T1ha72AC6
SW2RalVO6fWzUb+h8xQRSmdwQi7Mi9ol3Of67MMrp0YqC62F9MDktb3KWUo4
/rDFgSI1uNn0WluY3Ox/XX/QdiSh3ugxeuzP1289fJbxxEOw8n8iyR2YBdjI
BVOt2IiTIYMAq4JExffzNGLYd4qhjX0eGqstOY7z5l8QVE3zI6DXV3YaKcvi
1bDqjkGeMsMILi/1p+asnpt+WsjsjgewbJF/hRi1yrTrmuAnV53q2XgaMKep
43Ri88kE2vehH28RTW2353z3zPpqDfngdCmmOK6ob2Vg0+HRqifHlhuxuqyK
2OAmbdoEIxXA1pySPkAUlhtmZJwrrVvm9P+4pw6z39HxgWuYc2EAjD0MJXEf
td1dzLIIDTi0A3fYRNfh6TIkeJu1kdvxMyY+/51Y+fbbr3fhtmIyE1tugNBA
KOFxMnSaykY4x1Eslf5hn5l2aKWGgAbrE8hb+206DtrYaLMUb5UHD7B6smqp
p/M8Iwdezer7wuE5ofoE6jn5lsObc4jmOB84DXnUxd/APGFCDTiaye822Fth
gujm0lLcId01iSaaBRrqNNOj047CtQeeh676d/KUOMp+z5asAy2DSi7dlfcQ
cjNQmHJlpYKzf+8JKno57VRl6Q30WAgjRfZzrEUBsT+6oIYwcBYtitAkho2w
WB5xzAgEaqO6PrznE9tJYM4awzuTsrPkt2lH6FEchR4As96B20ulCwBFV4Xs
6xMEuBJfYUbbxjRLvSTUAk92nlkYPveM3Mc9mCU7S3Eins7ajRZIUSUUndkg
SsXoyuYVJRUrcB4tJ5IfbmN4kRR2G+stoOb4CbDJBokH8lfpMBEBkNnGp5u6
RIocoHOoFEMKKTa6qzpuoSQ2wK6cBdq+1aTZXIYR4pQtVImezf8epPgkqCBQ
kfInM3dXPbNtHmvvNV7bBO4WRFdAaaVelTkhCGjPGT3/IY5YSq2AStRXj4R7
cMtsWD6LhFghzsuiig5QRFPizTmg0ksoZ0j1I9gOcyXl43ntbENF+ncW0TGr
oAF6/uCHjdI2D3EgvIFBDiDwvxaF4gPtTDiwYb2h8FyqAYfrQR4vwZ97dpCq
OgDJw5fqeVKxkK4P9mK9r1nA7p1Gf1TTrSCMP61HN08dTi2NZ1gQa4XdiTM4
Sij/j9joujaeWeja+M45czdAIvechCHXsWO1ttwuSDupz56gACvQZ8dU0IXF
8/7JlWR32oxYtywJORdn1XlE1oMuaZnIbrdEUxYlxx9D+TAqM0yKXkFK7UcB
IJYfqxs+hrITTFruljICTK6Tytp3jkxLBDITLmCaa2NCdTW0DsMErCyIG8M3
ruXVxyCIj4aUrx9L2BLiti1aa2vztuss9AtX0wj69RHKg2cdLY/lXRZBMtZK
L2Nu7gXAcz+wAiTxwidV8i5O6ShKdpBYUj0yR+TJFM3gtX0hGxl66wfhZ73I
IOFmBLtkD6xBeEhPnn3+dxy4Ar6jR1LutDaK6KEC7PFHdqEE0pMO2HJ/PrYa
w67n3nkXpPlC6BSMPI0PptHf1vcw3rX5uQZN8yD/ybAQmP8U1WkF0tzTMWeS
o64+x/dIY1I3TKeRTL+k0wsiaypWrZA4UDk+8ytqumA3KoBWAm400qbIz4wx
3VU0dM261WlUQ1vQba+8OwN/hzgdRlIFR+5kQV1JW10cAT1PBtGZiiATQEx2
YRo+cglnHocRnJC0Z3GRxYnT3IcrEKfEeA4hJMQbZqvEiJEK3plTlM/XnPwk
Z6cQYwdPSHlDFFxiYIBEFTVsPwS4m8u+WNJde/C/l3aUulYpkpTBhkoGl905
tjcCvNn0QX46K04s6FkgmzcIRLdQnGPmXQURjWnHy60Wnt/UnxdXRlNVIrAH
ZSPFDFhdwL3M9NrdXln6C9ZCq6ZxZmmkNDaPf+6wK2if+aPSWaqdmON3MhyC
opRgr7xyg1yCWk0S6NxIIp6kpMtrJoHGyrhPtfzc2ofGkPshPfLEb9d45AkV
PZRKm1+hvWySI8aNv5cX9rCAJfcu0KmqN6wGUewQnwhws/9hnDDJ+MNHkM/M
a+ZapxZkh3VoWb8mZFnte/jgJh691fCpirbw+QDFZKlpyYlEV20bfp+YsBg+
AADXNSuSnNd+3Yzox5ZB1qe2om2SuT21KuqMwdIeFV0HtUztn9YCY9Yf0TfN
6y2pgfE3bi6iKESOj7j6voIvu3U/KYOmd0LgVbvUgAILqpvVvCDsurVBqcUi
Ikup8ugJBxq0ohGDKiySgLHFKp3BlrcBpc/GT0eD9qgpNATv053UgEiPlRxJ
Wb9t2gu7NdE+98IszYmGqjusGp0uifrmITNpcggNKQpvA1CHScDsvcYHGhZ1
oGia/CuDWIYNSdTwe8dgH0eVC8pBvNjKWNoWZdXdpR7ufqJSIZJl7lPNaIOD
WBOkftOChi19Kh8EYeYrwZDxdy73vKnGG6bv19iHIYpFedPBS9XE/W9Yh8Z7
j+UGrRRvY+k7EnrjvRaD8XHOflX+shuZXrRLlljtnCRuhbicgt7b4eOUrZw8
7QCZX80CPtM+mBeM/vP1t0QKXbXUp+Sm3TxrBXj6Rt006Kvy+dER8T3752fU
EzqanBKOvu1BLr2q/g5+iaJpsBZ30k9lujW5ma/oeo97noQoHnZx85k0XRUl
8JMiZJwaA9jXIdmyJxMhVEXV59NFWqnfxZcvB6aAaQrMSsp+yPr94LlRU32m
Bca3Nq2noGu6XkHwte8c1Au12Rky6bAW8A2eMD0dLxoUI5ZFNPtpzzBf2eeg
LNx+3OFzeJAKoMAM+gSx4RCmdYhTalmnb2JOnom5Tq5ibh5QQ/kX/4EmSv8q
kaBEG/0D5dNNFmpEjWxRbZ8y2pXTE+hKRN+RwJMqcQxz2Y58uu/VtbQAm7gv
CIB9VT97/r4Q6TxX2yNhEpSYuX4kgzlaxJbz1G/0mLyLZDGTUNVQV9r6/G37
G8FV3TBL8aWHwoLJKFLY3Qy+J778AcZiDtUVXLPg3paKEiKElWAuw4Ukd4Ve
Wtnr+zvcbedZWuC1F/sdey7gfs0ROkSopO5gHKL4Dgksj66Ubb5Dixf1UgiP
8YADCJxdm5jz6TbLJFTpbpb7/R/JRskV4eX46kgSf4ww4SYag1+zX1Kftoo+
RJ7YpmKtG0VHaN2VAdQB/LQpqdkU6eNKk4by6JRInsHCIR1bwYrO/uZLML4Z
305Bf+jeyIdcZT2L9oH3qVF5r9GVqzPi0IlvzXSqu8gdDVgSPN2V5jAttDL7
I6BuuMbdBqPG86+ChNqY6+I0wvGkIh8t+Ow2pwzBS+/x4tkBNR3XMLS+020t
ly4+YbQUhR73NniIQ2kf2yKjabx4Jflho6LeLExuKXt8+m0suWceeeQcudBW
EHH7sz98Hi5zEUw7wByNlPCdDLvRH8lSiuI7HX/R6++MMrVi2SVhi7QgophS
8kBezLYwbIUpLJbOZ722exzPwd9NhdZv0SnUNWCPkbRcW4d3RJezu9P9MZjA
MeISF1+8B8cRTi74J06Y/uOIUD4EY7dGlIeOtvt3+M0fFieRdDhtIPmheXdk
08g2KzYa41upHSf1OQuHOwbwO5mWIzf+VUxPxOKKbMYCSG877yZyqqT5fpGD
WehAWtAYgxmeDZSLQek4fxBILL18KwBh78yc4CWRqzTPZqNej0LVc+Xo1pH+
EiceJFhE3z1yovHQ0rEDZfSbFpWzib4StZjhnaU2eL0LqAGJFpLIyMv+bB3T
z3hKw51cSdpu8lHvm+lBsMIbd13dBx+n7u+/HkSAJZSbEn+k1riDj9JkkFw4
MJeFtqek0Tvw/FAZJpCunVhq4pr7muf7RBBovCszKag0OZIRsB/Hfj6Yole3
CE7urBxTJGcDqGV3U6LznGXcLBFqZNA/FdnTytJwapsKI60RTS8mC7hKIclK
p+Xu2/slKgCbfB0b5y7ZXTCrEgel86OWwSk5ZcvkvwbsVpShB9wwNfOS810l
EGrfRREMHOZtY35QFrvLHBjoqrv80GjAWG7v7YF6FZ1IqrvMfgR7wgZjq5YM
UwrPd9LEEOI6zYzBCttISkpyavW0W4colcFYUaRcVzlCqWLCmdfvmIlILqGC
YdC8/PhoN8NHLCv3IB2HWBvPpsWUa6JPMBUL4dB2287Lf4rkHbleRz/prW7u
b8W4pmudmZMdq+GuQ76SJQGCZVxaKjSWCexB/9btqJc4gbm5yumpoAOqC+1i
yXpHKN7H4lYCGrlI7zFbhGGo20nCOIciG/G6mPNrV0py7tVBGmGzK4Mraqdo
eJ/iPLYdhUXQXx3wzIrAWPgLXAIyEAZwHONDyfakJRP6izdSA1nfXl65Rd/u
MVNkTsOVRDVqvYdU6uopxbEwlSSeFkoFEHHsZsz7MKuv+KF51avTWOyCkfZ3
a+wqCJKsG5Jz0bMqW75nUVYeydMhGvpbHzlIZEFHpRfz/7bI41gxG349rSY1
vN2ZCIU+aPQ2C2fO5eLRwaYY7zGYgxjy+byW0ej7Nel8RWi6SwGT4pZEu60D
ed6PVgHwCYr8zIF7p+EwLSTPDbwLRKWs8Mk7vHDW+4INybejVvVe+zHps1ZN
gBZfVehK9ia/59cH+dklVCOg5gepeC0QdV/gTCpKDVRYFoDgsec9zxDQkDcl
mjwpM2aOdm1XlDP437mVCxnyyFZqC0jiGEua4bCofAPBNtlqSm/7EdJZaM3T
782Viajh4VXNADpDk3c9K5iAX42Du7TEiW3UxjauvNxYtDbXvgjaCbkdqr5L
+2x/wnWe3sYu0r8q5o0UAxxM1T5FJzFISW6yjlnfSy+nhzqpQ/D1VDMFDE/v
VWe3SDR80VGk3VSlaIkMpNMfuHirsbNxXqSacw2JnXvAsZ1hlC0Dx/FTjwCc
9tzjXqc6TziObNFyuTV6hWiXOknvr2wZW3mgDbnt4Pkmdc2HW9fCT1KaXnip
GqqYqlsJTakfxpEQoMfTwqMZ2+tEvxLPwRYn+efVIa1kdZSZWnVR5pMdgrTq
EapNVdKmnNsxaMDZXrxxXNJRGZ3Zr6JhJuaubKHXZkZcgg1V5TI9oCFiV7Mq
5E8m8efdu9DMOgfUx2jeFQCVwU9kdPbx42+WnKDaeaIJlFEVCINltx4rNsqF
0JNxWuczyrLSi6Xz9w5YSx8RvAQ9YQxX+NUvw/rDUPC9fsLoLuqiTQf7mgSy
R58t2grCJ+BdZmV9zt4GHk75sTw7NsRAKkt7Tg00V0rcvuYH8WHUioF8S4gY
ZlZHWs8Y4g3N2vIpXmJWyrINI8FSo4/aP6iADP+MyGLRHd1xF0Su7CpTjgAU
DPeNEj1LWHryhQ44BKY9dk9ulfZ58LmbTYtcjD3y9ylPHQDfzNl0lkH/bojq
MxhA3rerwQmGvcL3u3SxmXXIyBMK6tpwqiVyf7DdPhDN0h/1r5UxKfD0+h5t
6H0je+uQKDoz17CC5mK8OIetOBzbj6QxqzH6nXtZ4ZSwVRCmmpNxDQBr8Ob6
qSUcIGHbXjUOgJBHuAYfqoJcVMs6ue5ayOfR+4NcY3cznTSVCj2bdobYfMfX
pKPBKucx1RK4Q8XALed2INUmf18G+IjygopJKPKhmM3YzorRamiwoMBZK5dV
or6xq3ff9BrM6fXIxEOZHbDiQ+AR7QrbI2/CbeCUCwR2ms4/F+7tHVPv5EKM
cR7LsQpGAyb9Zh8t5qIv+FYhAuqn9QDl53rY3HDZpS0rYI/JIdRVUk/ExGYa
1O0ZIGDZ9cA2J9qfFMUJCoitMwiUPwtJNuhKJNTzHYcsgqJ6lCUKrg09utHd
E9Elu72J1+BuMvcRxs0g6AQN7Z3TYntb0XXTCBTWLmHtsc3Ex+9r0YuoX+Cy
wfqrk5FOky11NkLV39INcsvyFPiAZVMKt+g1XA+Y66WxiNQGrnzTiO6cFa5u
GDo+GNRQXR+x6eyqL/FcER4LsELctuLL47B9TYto+uREhPQXykNk+xwuS52B
B4uJGg2Jt3xp0cZZIifgrny0uud7/UJbgEWSdPH/aUxkukUb2c7Kgp7Qaal9
9x/Zfz2t5G/h0aqKiPJMIQYxoKUj9/m+q9l5TjAQUMn6yBwTDXfXAE2RWBjO
pNqcz9EvKnNO0emuCrRw9tK884F+Q04dNX+j3kL9bmjmRqnAlhZEok99xMlR
xTO2dUrUNjA9MYbOiKh1IU5gvsCJNRugLotdfros0F9WXjk59zggJ6wSbuZO
8S7A4maY8SibA224aIBCihtNFOhj/svbJnN5xuiEQke2sIT3+60jCZQZ1UCF
fuJNH5X8d9aAEvAyAuxJrtUorqVBvKqF3lmbnvsd/U31n88k+hwECs9S60Zx
3exYzesQurrYzrXNwbH6I79XKUYTvUw0URpfI3qpT80aXea4r9ruv5UKFaPh
b8GkocDhXg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpejp5aCliFydguEk96+z/phtZGEbjPnsZDS6vx+hpm1LMLjm80wRyxiU694Nj2Ax0iFHPql3b0tes9hJC2gVLgDN1NpXdq+fZ8WG4PQ6lRt138AGxxVPeqAkRsUnViMzb1NFmAhqEiqfjDxfros+P1yrWPmdf21Vyao3dy+zwTUr+t8IJmXyTUy22LstrRQV2nxRzNjlR+M6SZ6EZzFwBE/nHpS41jv4wYjvMgsSMdvQ6zh3vZkaBJbt7gb9MD5l4CKXVaD/Osy2AKq4RUtIKsw7uSXK3pqcwlFU8Vb5VZ003/eQ4LfchCr/WHqUygSMqMKT2E3x67NunxSRYLXcRcGo5Hy3mRGcZB2kbznaGvvELM6PQzoppREq4HNp8plmIW7UfysH3uwWDcsowBCLiq14mZPgJZC2ALol7tp7vLUNXLcKPfpeAC39hc/asGK+2IF2cmFbyJ5d9fN9nSoXCpTm4KiPSQtWngTxpTI4eh+TmFBSiLsmLXgS0aRl2/80FQYGZwVflJBT2tG235QvblJ/wfjIPh3b6pNxeqVqpCK+VEY/nAESw0ypcaUig0V42ZW3w/7LKfeOpQNy/8yCbJ9kdyC2dSh8iYfBioqjuXHWzsQ8suZagLo+kQ5gcOGq5mKY2JieRI0zFJij6vv85dVsGVtiTooEw6zq9Xa61ok2lMvWLRgPealbFiRuPyUeaxiSBVUhECrM93Q4DuAJKYQyLGTCjIOHTtk4B7F1dWMYMYwdWU/vWJHx0qvwT1BmTUPTK+MqNSna1eTn6d/XgYSl"
`endif