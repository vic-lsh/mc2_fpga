// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FWc/WtYb0MBNCQ5sJWHegSAiEKHY2PdIvO1M3k8ZL27i46H4dtK+ee03Th1i
RpX3vwV48mcCcEjPqC4U1Z9iQKJd2pSCbYr64/NR/iHVIiVze6HFajxirLEP
7uEsFxi7s+y13TgOnYM7RDIH8ucy6eI+LDPTbMC1tMKZeI7uzBU/dNc5g95n
DVQL8A4LPXMF4upq4ig/YdEmSV2BrkKzicc2srQjmV/fF3aLkkb4fm2OhlW9
FEicf3m8Dk6ZAY1GvDWnpT3W8Qh2R/jCcI8Dw1ZdwBVUtBSZStixTfncwkOp
5jwDFqr2I9dS+X/JKIb7oAxRgVGXTvDYWyaecoGkAQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pisy0Y9cnzTO7f3RlhQ9aKK3p7BDQj5I7iDFM0rTaoiK5TUcmGyhoOSfD2Fu
C6U36RXMaWSveXZNExClS+ukg+7ARAsesBLv9BQcgFz4MV+7h1qaT7mT2Kvr
+nSeSJI2RiVir0sx4/vIfbex+eBTQXMW5qsumDE/nSTKlm1M1YFf6t0MC+g9
Ssq/JuLzaY1An6abHnyEjyoZzCXBbl430CwJ9TxH9RRATx2po3vMhvsK8T0X
jzqv6Sd17Cuzbcw+yed9zUwwMI8mtxxFZBPYgcvkkbddPLdpQEpdjXGNR8kg
DbvNtlZmPv4M7gjgWhm0nr84n8zUnkQWspxlx2szCg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ifgkrOHopMm1tbjWLeRrLVjosN4tjn3Lk8MJW/0pn9H3xICHz0vyLZPl4PMy
pdvi/ebdp4cYFSTUhZVZ2oX5DJO/RcduneV3+qOcs9rGX4oIrt8UOswaZMbv
NpwI0IupjwC9poil44ThBKUJD+nu+CPz83PjbDsYDkBKT8uvqFm72TdDbIKi
egp8o/wegYfyktzjzwK9ct67muePVOd+Gkzn2LaKyfZnQ+n/MRzakFKvgiGh
rdHki7utkrExhRB0mpq8qcvy8PCzfDYWBUiJKh2NxFIPS7ZjQN5Lg0TXQM4n
3RLx+p+b3vk7EmE+8jJ7zQ7ggICg6O5h1ktEgrPCYw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RPaZYm+bqHqOqKcI/pYQ3QJNaOeVD+JQhSSplbLLIFfw0BUJpCNfpNAOOHrk
TsNPyE+KvOsbr6TUDXi05qbgy3vGyC213vcTzlP3Px3db9V0+/KFJCKchG58
SU7uPTPN7pNjpTkne6LRttOyZY+cuAsKqwiMiwNBFdnA1X1BjKJ2o1NdL6Qm
R4F8iz9+kLvmr/mvpuVe5XAzR+DSW/9SxpwSExG+7/yJ3nuqZ83kpXAjGBH2
dG/SmH0GdSoa2uwLbN7rUo667HwjUOvU7tlvKr9cYUmRgPmZvWVqFkY7QBTv
7kPQr+6l8DzvYUNW2Zl84yB7KGfgLcDJ7eNXdNbTzg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ik9fRgjbQLTIkz/KsRoVTHBVCUrnfYz0bOpK30fBezNtQAFlp3KUJqqbZGDk
3b1VT8McMLcUvbaBO7plL5D/gOdmjcJhNQBr9wiO9Xpmv750q8JxCmCMqW79
jbgugwU1h7gxwJrIXQBjmaLH3u8n0kSf/R7AQt/XfdwdbDaHbOE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MbSP1AAtektVTQSX2eS+EzXBV0Zvssgg97lH2h33z8QzOqwvw0T0mR3d69vl
2EihajioWcCK3aPO8e3EGU4QIcrOaaf0hX3P9h7FgqNmhvdpyEq6oP7c5nsS
yAy4NbufxGDlmciVpmZDo7Iu74JyUbmuYvJX/OdPBTVfJzsQA6UmSMZtkNT1
q/K4ztlunWKLpm8+h9RKc7LdB7trtoSrK2nOAiEmoSIpHsxDGyzcBAntg2Tk
72MALiBiuv2eImdlA0Xc6ayr2lqRA4N1VngNca/KFnptew6jWvI/8Bz1/vDI
WBmINKnv+28ykVCUwNwl4LAfCgde8LtiRr5sxedYxoFhsPlL3/Fn5u8GbolZ
Rnpu0iPSaQgqsRA9A9BkiyyJCrhopdU33pNDAiJOviAsjP35DRPef9BQlULz
NZLv3M8nJTntKn3yCyLSQ35paLvx7EqxeAsYJy91tLODr5BChSDEIO2xB/qF
qBMl/uc0IIiObj0upMFJHUrpSEEoumIa


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ETsqFvQoxycoDpX5md7rPAAHsdJp+AjO7f41ku/VrPKqYrWjYWY8Zbc1v7CX
SYv4lNRrcbdQXgd2pusqPzQ05vLehU4Lf1OLh2Sj//GXH45EAEDnTQge4l3K
aE6e0ZavDFGWpPwzJBn9c5syKVSOvgso980mnUA6zXvGUBtSLVI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
flN5te5cU8ZtqSNUMANPhvGo044KUJiFaywTZCVbvCrXx95skn8+B7pBnhTF
MpK7LtG8MrxRh9fcSyfkfSPCXsWtXjA79oCn1ZIRf4+a6gBxpe2U/sjIySE9
ZmIKyj+cMMxmJS7b+Ty6hQUWxZonVxPrzQncIhmg5NBzJiuaUJ4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10448)
`pragma protect data_block
Zbx3VjC9TmiTGFgH0QE9XKXGNYW1l5+QJFzz/ddQKEDG0AoQSB1ZtI+2j04n
28suVp2u1cZOuY3nMQqt8yBDwYD0guTdZfzwtMctrvBpTZQlrOXjWuBkGQtO
rASvbUwgZi6inOByWhFfiaL9yUdxLT8wfoXXPAWPrUG01EKV0FvOkuKzsB7t
ZGgVRsDjt82dPDOfoyTC3F3qQ4t3AvRu5X8a/5prpPe9DCE7CDoRIkC+T9Vp
MqrZqs+fTpVguO1LRwIuJbGslr1QeyfrSXyWuAPadlvEB1biuAxkUyhzFHUp
Gu8oMa82FAYbUwrg4uBvLrjw7KKH3Nv999YFWlrYDN+NZtmLLAaVduadiZDf
K5QsZ6JqMfUgrtFPn9rLv6Nyz/UAuKIx+Y/kNLQHzfMp0cHPp98GrFzEZTnC
C5oxUg7G4CIfy4El6ykzT+/tUNh352g+oapoS+BnNf5t8xMpmOmLfML0Ej9L
noE/GbS6z1b/lACNWCP3y6GgGD1LSZQr2wZwcWgGaqO/j/m8cUP04D1C3qPU
bf31N/J3tos3iOetwruorldaXAElKgg1sNkfxsalOqwZwzgrygeoAIgSCxt9
J4zQiGHVgz1mOzhfV2jXEKiEWZmwspQlavB+x+eb72uiD5zSjycQwHhOatsZ
5f3zBrsJQn+u3mHC1xfnZDM1ZSEFbRec3jyxPKo7n8yYXeefT2iJ5kdF2EAp
D7rF7nJ8OEq29d/COK0cw8SqLpD73vBgnr9NfF+M+Tfa8/KQCaIruCCD3tfA
mWSAXVh0qtJFh4BSQ/cEAxlL7ituY1AKJYHdzF5jjEhuPz1YwpfkT1huSYXU
jCkCOTCwX9QvY8959cyp5GJrwErl95uojojaACxg5UEFoEHiE1UwC6+VuMP3
TlcnAm3Cz78N9EvZH+Ey0nwdW06i0zTU9nsiMwQJzbgKvQowAQI54Yr4UehI
N6kWJt4uzBeyTTGZhctvJw0GdVg25wDlWfapppX4DfXx8ZEqOyzRFurQsRUP
JvpDrEdJXDAS6xbSMhIwP1vaAHktKjKaBuy39B/Vg6m3fHEfu/b9cQnlDJ5I
r1Ao56t4/DZAnfCOQ6Jux8l4CoYVJ2IiNQm7lagurLhB7W/Eo4MHnZD55z6b
aLU5Oy7JLz3cvT7wYzY5BONJhBCnjJ5lzZEUILRxdOYS9S4AfmzQCLPhTOo3
Hhoq/1onNd6cdDs/NhFCB9k+jSxIR8gjSOaQnu+UQQPOkoJbDJq/3Ec1vZ1q
2FR/5F6TF3kAw4DDYor6PQCSAZ3OQD0xZOX/C0nwosw6Mitrog19NWdADqiB
pXShmlWidwN2rgMLsAscdEdUK+TwGNG55VewGylL+LiTf+wgtnwUu2CVHCEy
kkrmgvegCZ0w/Mc50y8JJN/mwSh5NmpBsCEpanH1WLUqXh3/XOdP4u5hhPoM
jcWZAmOFTNEyzqryrz4rCi4TJQF5O3rfN7JQyPvcAFW7MdJRsGKm7Qp61Kxc
WMpnPdvAoPsDtbsNOzEeUtIBvz5wyeMUV0Wn7yZvc1ASUvebm0VhFDaJJv+c
qFrQic5EzmDeaZQefWWMReQfWuhoU6K2yzsy8tPx2UxDA8HMsgx2/M5HGvuM
4GZuVV0XoBUveVO1dD3JYsjZbRmxYwbeFxL+dq3KNSyc2SlZ016kCTBzUV39
OXuQAe5EOW3AN/oSqw/tztxfUZr3d0F77ETsBajsEsdckPqAoFYXxJVN3USs
yThvYjD24HxQhgjJKrX7qc/neLzODbWRlQFjoibq+M4gZw34B1HhKIXBhhnK
F6dOJhqJUmDhOY0iMt7wqmgfyg5dSx7gQYc3vqvw4UGBu76dsiFZikET7E+K
Vj5RHFc53mDLz/wu6jt4Mj1YSCj6Xwz06hxsnr87mPnkzi7IMI+1hB66vrk/
RgElAZhfWxCrup196zyPMfGJ+NNIQ6AI42+oPn+rHsfo6PglNifVvJh0arS9
KIadOVtW2RzlxR4ktFyspP1BhwTImjuy88enBXPGRS2C+7K2MG1DItenm5bI
FrYln+q3gusugeQAghy06DxR1YnQpXCAJgjJUZDmkNEdtZmqv9a7tTYF4bX2
UE2g/tZaw0S4NLrOI4vzd3SJ+FF0Jo5khGMbTFMMRyEhFSwk7Q/y/RnVcQe0
11Vv4jsfCsqGgpKEvUISvPJOlV0eHisOy2HZLQVWTB9AqiO4dE5uyOYwfj/X
b1jRWYo/u4JyU+wZUfyzhQwlS/Alaw4y+7a+GPlzU2hnj80B0Jmq/jaaYCwm
ikIh+dy2SNbR6ivU5fjgUP3hvjp7bjw7SZIQ1ob5I9nZv3+8JNhzbG/CV9QZ
16eWu3A+ApNBRNhsVa99xZXBXtWbxsiNwprkEc09Xjz91jeDAthzWCRVlMxw
AClF+R09bKIAeKi7C5nxzdOn3+PPoXRgQ3wCCCK1POAaAAu3sz/BjdzIDQS3
9f8ypUtuZAS0r9sBr7Nlotj5BJDWY2UQal8sWuB8nGcSsYw7EW2FqY6Uvhkp
97ULmHL+iX7PCikwXrrjU9AjPjUFo16SM5DqQ/MJupT8/boi3n62Ps9QEX7+
eMyiYPXscD3Ntc9lJwjfepEzEQ3HGY8wAvBqvLCbWavKkDXSGdmco53oAYTf
YlQ4dyoC/iOH4yaeMmNrWLFmvn59CsJgM42zrefmsurw9vzE3iqykI9PciYu
eN/eLL6o7Fp6rSYGD2n+fu+kYXgQb/XFSgUE6B8EwENMjlxnpvNms3YGVJ42
zSkSuOyC1FqYNgcYo815SKVrktTHonZCRfML26BtHLpG1D3sbksu+L7Uwbn5
SP0u7PSdDzkah3kVbjtQCXNANf3vIpMzvy9FnyRjfXa3iQVdUPpc4xYvnT6I
BzcIi4yIdmRef/DmP9wZ10hFRbNAraA4PjxaKTVM3sDZKk83V4seT/qWyiNO
QM8Xr3eBe1QRTnhCWUNEYYQMpChLtC/4ELdfhkK9PAv9PqftqeZJxB8oHdeq
Y61s5/+vh3Ai+uoB3bjiOtKjqyBiSfBkRyUyUzIR+2K8bPsoFEnJN5yF8Suf
x8t8VAIISupVzSzTFm9pDQ3WRBWO2Cow/MnTN9b9EaB++6GIxhX1wx84mbg1
t/dbrnMKf1cKPBCmcJ2/0lHxtTISYTrbfyPUOEEvHWwGVDWheMe7paRI/LIt
q+hCe3O5LIAu8k7nEOGcnJkBkpiV6Q8WpcCJkqmYWRf5POiMvhx+g0FrPeA8
VOUOSbbB2bjmqGpVM6cVI/rEx4f6iNwBb7cAxVnmRd32pvzuTaT+sl6vJ13V
UiDlrGwXrl4j4/AJnaZ4AOMLDjeSu4cZzEMEo6/opvJVh4MWSlRrLnip7vD4
haPzly9TexkC5d1+sPad5LED8oQptftN8Dg3FK5OGgVV5ubpADwb0oYAukQt
xfPI2LwIKSt1QS1dQZ0KEFu5UQUZixjQAPeMD7DoK0s+ZBZU17LfS4CsvvLe
RWzLHTwHde4qi6utD7h1zYIzfNN/3S/bgAa4h4u8xJaXipGjeH2DltXf2Yzw
++2tBc+0JC2pG+3OzivnluPDSeXvEu06DLkhsjJva9mVUtPMinBMgUmCoCcV
6NkTBx7Bh3nfmVlUD14MBEP1fxxRAtBvddD7d3gcv/20GwUVsX++6J7h0BPu
qxslmIjF/V4hrWDg/IPK9i5vr2NU2WALHPgwz6rNw94YlyqtRbtD6iOS6v0i
75zszzCtvmHQ3higw9+mhIjVkj444DvJpVL+1f4ToQ6TWLGG+KAFNp7Ojlya
xmWxwGFWyzrSkGcbVTxhA/qDoNMsZN2GQWaQIyie76LsIO8gD3C40/qLubzv
yphLAhmigRcUZiAcjAbnHfeywurng+P6mwPDOzVLXYZxZGXX8Ox3CBUuMaxo
iMeV6A8bKwhV+5Jg3VqluG+YKqOT3CmJSAHQxABufw4wYdYI+Ix7YGJ+dGHn
SnY5GF7sXeQIwjacHAPbYNF81M//MMAhJjTMy9Et/H2zfJnjMXcVPvpnBTls
WyxoUcL0O5yv8dheilOuZAMrbkSvtcNq9AnWJDf86/zuWbf7bfKtasEvQwkQ
tmbGtA0vRi6VxVRuPqpYhLJnUYdc6/dAe+NydoBG5pvRIV87vGIPluckNZBc
WT7DF2Jh3x5z8kOsKZMyraZw0j7jKjGnpdfTrpRwMX7iHgcP03S35aE2KP7j
BlvjbGH4cm32Th0n1soNFAJTVPzt3cHD99JOmH2GSv6Y45RNndt7uzsBRyMa
r3cgcY5cIKLtVOk3EwtC7GyH4QTgZft+sSzaKb90NfkWkwh0FWCn6l8IaA5H
nIUG9Rm0EsKv8w80NRIqosfILGZiqwsuh91+vTnEGfth0wLgodcm8/fhQ9jl
hTEhJwdQEUdM1Lh2WzNPvFJu/qEdSIBmTi3G+Ery78jkIYYEAhlkTW6aQuy5
IKsHfQcrdqFIlG/IH/07hussi5zy9NnQjsY2PAGx8tCJH+OH0emknf4AqB6P
FV8iPBmXSTX8PmdZB9ynTB9eXSyGgK3y+JwX6HdZxnKZXflDHea0DAIEAsmM
JbLkJmb766Mlr+JPcFzKHZ2pv9ZDBdKtIiWmrSsqZUPPkS0WwQQ+GNgtz+Hs
2FuLI/3/W+DWU5eAY2XnzwzGzy+IMM3ElkVUvXFNwxhl/JvTQ9zuS+2n7FLY
ufppfDAOiEMHuZbryl3rS6Rde1FFHs/ZARn5ZsyPS7u6Q2j1PyaC2TVlFP9w
UzJsM1vTsSJqt+/rD9dcnVwH2ByEsvptsBa9XvFSk9cvCiKm3QSX9HjZZt5a
xTthqchn3tkkZNnlgSx0MZEjJi+TSYpVHwTeQ77PcQe05cp3IUXCocIbHw4L
offs006Rly10ljjudoOtXc+ZoYLG7YfmT7muvZbDtqxhjT1kQzbbWBaNut9V
TfX4O9Nonsr39i5vUix4NpWmkfCATMdggldzy/NOar9asPLUpr6XuddCOgg3
TR/ekW3H4a8KMVrnlKQ5hQn0LEIMyRMQebZxzODuVfG94fOQV7tpPwxUJVSA
0z5yNbUFPqOQZGqrZyCIESyEmKa/T9VUhYOuqPXeqYUWRTHufgiGISzah02O
0gjaaPBE+u/FU2CYSEomNv1mfcN5isHGD12W1UJu9Lv4B1bYZGdQAO8NDSwC
L6aMwvKbDkIL4Kx9fiWqntHXBc8FXGZR/gt1GG7D+fw+lecUf7OhsevWRR2H
8q6Dgs60wOi2iHaDArstPWKUXoPbrD2nieo4EpS8lvAI7b1RyBq7DOK4tNry
qHsIg/ejnLcv8P17+TyevK6Ywel1lsUqXT4s1lBX1VrIQBbRz8fdmQFq+x/j
qwUdNfVPUWVQqMni6RHgxHEiS8GWTfIfTSnoqRA+ErlGh6C4lvEq9WykAOGh
m9GrecxqVcp/NVuV7WpLPqIrTJZnvqBmtMcWTFbArDBc743dAQJFLJlj/aJp
6Lij/O05CVifmMNbwFqboYmrJJ7yuoioMQ4Rk3NkeKIzQomFtobOIs++LNRB
j/hTwvopFh7LnLMmDiZF6oQKhdOFZq0QY4681srYi3G6xkWG625SgTXHZ7qJ
wxI1SFwZ+QNvmgpsPn7jVq7mL1+TCv7+st7CMtgCxmZ9Mkj0ldTEdw/zJkIl
ZwBjIDllg3PCgbH0jI+Qx7c+/uOzjjnsi/DGhomBSBy7GPKvfA9/D31j7uaa
O3vn5ER9VLn+APooxUAyVI6OcSp55n4m/mm8NYCNV+E9HUL/tyj5nSViJxQE
d76B6Gb3w5i7STsHL49dKceWw4mPv7ekDkT+BOVHRRNzqyvYmAJtypgAZABT
H3bnT7rpD9ePLDsZavLAVsrJeGJYqMoX5osxBBUgIzdVgHaqf9a4FCHTjoPk
0f95oR1Q0yFtm4i7Uxs4xf3E93FL8ArvHS1DHRzNFG9B3AgfjIoxf83XVtaL
ahuC+j2Os+NB/Ygu9GnSbDYT51XftWnHSIsPbOPa1IytzTLpmg9hUAfPiZRV
Lb9rfoTfXJ+mcht8DcgMRA9DqagIjYnNUKdGmEHzOShB8AXBI0cC+i/INh0Q
lTBuPzfmQA4R1Dni4kGABkDI/htyfrxVPBBQVcmM1lCQNjdrZ4qV6WcuRMbA
Os4ZtRm+HR7MaYuQKVvcLZOMOznBjbPGxstKO4S91W/KVolGinlfNxBrJiCO
0rp6SF0AqIgLNj27Ccr/v15OowpmA1p+ZWSZis2L7qAMzxf1WiKc4aLudchG
5dNs+O7TQFBFTaivdXiBaaekCtONwUUSDLA4Or0bkBcqnJQcHBOV8nAnaxuD
tdjhrVbMS2iBf7Y4HwWGIaB7cM7DaR2240b1CsKmGx1xoSbUMyis4b1ErynS
5NGoN28kRIS9W0T9cAijXWzSqrnrEMgd0XlcYQcrvhhyV9pUdJignu8Bd/Is
6QmZiATDlNbIA0f/5X1dboftynl9LlCjNL4PVMguZmpKH9KMENWHQG+8BDQu
PlAYtANpJwW9lbfs2Oy5CSB4YXttwq8T19qY/RE3QbKAC8B7PNrYPpuljFbf
wcVYUznB9Zbz8A6GTDnkkAztO8V2nf/aTWPHxHJ/Qam2PXjtFyLLa6XeMj1X
SG1lFHHV9HVPAI7jFA98P0bzdf44if1tgee2NstmdGsRXzY2ktPVK7bqO4z6
IC/pyQk8RoG1hAn1Fr2t5tboQb62DgjnAq6KTQFWf71w0wHMR7qlfC7IyMLK
mLrTg1RN0kVKANfhyJ/QEMlyr3AvzzwAuf8ocndqMQ0Sslvi/U5A6APnOYK0
L1lhdPkgnPU2OvIItsuVytUa+hvpeJpVNAQgF1EAMBX9LlYAXmY9W90hy2YT
48LSR7CrLClMsjp4wCYeuIKS8qfnjyj00Bu6C+S7xK7p2NzMco7Gq7/6sjmM
8sunqOQiWODhFzK6XKHrk8KYILT8WEUiWYv8O1Gn6E4YSyCtNvIHPOBO1UnV
rEX3gCta6TjafMYkiodGZx7X+w6QRVd7VmQJDl044Oq3TMO2SPb/Qgnyto49
K0MrRwOWYJYflF0Pd7yzNklsIg1QXQAsVkJ0aExyTFlW1Xa8gljadAruASTN
yj3sYWuEj7jaMv8QeJe2Dr2wjO+s7vTkL/+mQU1LeGwlSc6qphQyiX9BCsD+
d/jFC8176D+62GnvqRmv0Sg25FYmX23LVbSjHxKvHauLEIpkhQoYNd4WqrsX
Qs8BjVBqrT9LmLINWj2WdV4Awcmi2AptaFntguzOHQZfKanWg1isTeQnS07/
LSidMsoNKfFMfiBrJsBW+k6dUV7N7rYNvR3vnbUQkV9kX1sYZOhmH7EeCm09
ET2pxs0x7rdI2toplfjGG+VVcfV5tgS+8GqU+AQeNBBUGYW+CvJvaCIE2LQ5
roZWsl5JZgx3cPupJ2C4UExOGRyM1AmFp0LdGx6xIlqq4jOgjLg+jMwlmbOK
QhtOtL3iuBHu151oY5N8dIo1mMysyGCHqoJtp1nmc1NsMibXCnc9VXetVfBp
ljFVREJrPE2PjjN08CqS/b5BmCHSMICj/4vFzenRWxD2ztriHaUBePD1+cCn
d/e0484FNjvag9vCwXyvdtpPEDa0Xpl8/iNYYewIqY5wNIBpMehtx2AKQgbR
SOdWBIaU9YlIOww2DDJf3E63CHxVCH9XALMUc7Svs4Qlt8ErqtmlpDPyfskO
n19eYxI+dz9bqsEZEPZobe4q9zEIv5xiKQlMF4kLk8qGSLK2iquMeI6LIaAK
UYideMiptyQRqgL0AXxj4N/4kB7n8Ir5b1VGqeXgM2S4zrgZkePODuZpZ12N
424+1PCKrBuQAVz4nGMUv4ts9XMSBKKah77Ds05hj39qFKKjcYiQDk11HBuP
avg7qpP93ZdO4Lua55BYvuJ7VHYMeWXI6YQZGvSIreVwO9ga09WFOsU6ks58
gA5R/YHanrExiv4h/qr1C8xF/ib9uh4JUn1LV7R7y4YR6e3WuxvzVpM9EpLR
ebrJ5SB6w7K/1jNF5sSxF+G+Rm0UlqY+ki/OzspMi/83bgq2eMQRoRIkQyln
x3J4nqtGebtC3DdYSXdxd6I0pSbHvY/k5AnV+tBRx7ihYpa0k1EK/91XYOZ+
NTtEHyY3clmp2gRPreXRCzzVSMMjxpWFKaPS1ZSSwDiyE9hayIkzp0E8ja69
GkxLLR3jVe/IP3/SKQkMigXwrJnh0LZk94wUpfIThffjSAne9VHHfXEK12BR
IobVjBcw/ONIl2oFyYqdEe6Bi9KMFszDkuO0Hi8a+0AsXbPIf20AP2Fr9QTx
SPrAuWLg8RWTRbl9zN51uuOll1M12KN5hrh7RcnxxMKYubl4eYo2XR9nU+Fe
08D9gPSAl1A4yt6V8fzgznjZnx4u+DJYaAlN1jxiAHQRRv1fhQs+DRgMj8G1
YBNsa6I6oPzqmFJH0N+iVFS075ySLWuvJmcDVAGWT3BwtZY/f1BZmmBRLgt8
70KsgkAVOzoem+clXMa4egCTQbDK/LAscRnM3DHk+7wmgftI1KcgHnanc4TW
f29y+B8JC+KnDP6o1jvRQmoTIyjM3tQ72KCUn37F5NDh7ZLv7izsTBTSGT29
HJgKXHciVV/s0i5IAB2tM/56wbRi0pshDJzH2bcvmUkXSi1bCdb1NSNvWL5O
uodT200dx7UVDhQOyYmCT12qehBuISynw/qnecz9eKw43G9F1hD/ZrAkLEbM
zBcTK8ebSVSdjcURjoq2j5fCIBQOyicr3QWQfMqkRDHl0WBb7Taff/V4nSkX
d5+mV2vU1tCYanUu6UDA+fFHTpiVBk3EGeqZVcQTpwB0+QCvSpqkHL5Gsk3f
mxQAJeenmILd3AQ1HObtiG3CvtCz+QC9BI3e7pbUsRI27tpQeAqWLxS1HgbK
u3b6lwyvFyKC/z037yO+UT5wcNvmuf9F+os5WjzbB3CnYzpNpaSUcV2vlrHa
xgZ2YzKw1T5/t7NpYrTNCbUDGCkUIwhwycVQLmTy2De5N770+3MLRek3yaW2
fojZecNOcKSM9OOhBJpZv9ZtoddLTK6CjXmR8bK1YCa1CWCanj2lgy3CBEiS
U9FNUFJ949L1CfGt3mUN67r7ke4VIxsOceZlBSC7OS6OxKhmdJbtUP6l/Gwl
O8ZN6Ty3Jq/APqKBZp9yoHGWwz5Y5kNEpPu0fzGAgiUeeXiG7Ve0Vha/rqrq
ZdYDrX8r4j4356b9S4hBukVeKynLN7vM8eDtAwBIzOTg4FGASWKDoGrenp26
bJlwaPTnca6fZoGwj4LOq/KrWfDMRyfGg/76VTmh9m/XWcgSiDNbkux4B7X8
p7wvzN1iM1QZ2v4uQrWGj9z0UDi8rNJet/rnWyCFtdNVlN89B34NoAB41fK0
cY6RdjpnwpGmg5xlqjkSQTiGyl9HQtsf1dNTWas29U1fYi5n4z92vT6RFYS/
Hggp8GfjRxV1nDEdupUKX/uaypqVTCNKnXqjRDa2kAC4Rl5UU3bnR90wd9m8
ThiymqJ5Umxth1be7gynHcbcrSwIpl3QdpUcCRzEKCRbdVggx68Frwab9YO0
JRp3EGvNxu/dUS6drZ3owdF2KkrhtjoVNYqBwIltXK8N2GULxs8jpd6cSFPh
hJwd2VP36zznNPkHHJXRROOZ+GilIHNJ1S2lMPam783M31XNFrpNqG+UnMoc
effC/eRaiSlmGX4Lu2ejnO1hXyEe/MT3bxaD5w8h9GspPrbvnuiGFtbbQeF9
t8ZtOVjpB/bkd0Cpus6jDMXY6vKoHbQ7JOKjWDYg3G1cjHcN1oTWFzKORWz6
zdXFCfQ+WKNSdL3oD+MFsaFELQwxuu6r9IAA+FeDaIj+rYmqFEO3cpANR3Y4
lDBqNhB8ysc4emSTtb8E68fEac/vyLb+fcCIfNaw9QYerHtF2qrcubVeRQof
peVF1cYX06fzB7DwF0+jJTW3LHDC8wPj4Gck6kwqpSmow4dX5aMi9SMSoppJ
YBAVfYh2uJl6za4CLwzICjTOKwZiBjehHMGBxIsdrQzbs9YO4P4P60ISYaWW
ACqv5X944+OrSiGJkRMMI2uAB8bTwExfpn+h2GSoL9iFywAduSzLXZW/q+yM
BnsSXN0CXp9u4+xJKj1ulDHPTG/0d0GJOV6aJ1m9+gJzT/hco2FL40NFKMO3
hjvNIrWkDWUpapPPD3O5G2Z0+IeAgJfngO99AjEZsjSoWAnDN3fRve62Rsnj
4zi4hJnaNvdUOc5Sc8HhhupmRhRElFfGxY8YJ7vJIVU7n/N5ewbk4CmoVL/Q
zUY3xqkxiyL5FiaxEqvi+z+oUDYB91FpIo/EDAs7vTtNs/zzVfRrdaZCKhGf
RD1WkVCLnCZtSHoYiLD5iBL+jwQRsMk1v0d5EIhsZG4/fG6fCj/iTauGa22V
RN9SFcSISTXjM2OPbPpY6AMB+4P47IzHCk9iDsf9D5pA22Z5PoSLcuioJkbM
EcLCgMfHr+HwjMeKTSziBd5z4RcpTvQ8+m+Hs9PCCvCQRzozz4ObG3jqI62w
yLkldUWsEKkN7A7hAswCXlp8ux/sGYFplKdJ5fYnKYmKERoBMw2kEMs0C15b
YmXisHgKDTlvASADAodumoa3ROnhi4cE2pPYXRBlG7roSmS0X8oMKwBdDS0w
37jQuJW0T2E35HvsQJBpwlxQHQOVtkh+flkZB69C9Kzo0NS4ZmNK10rgbQj1
RSYLRXa91OU5W9qQ3u+R+YGt3cE5G2/XO6bUYSX93BYeXeJKpu+82DNSxPYu
Va6Z3cClFrv/VbqVNW1CiZvXzYGhSGfvKAB4zNZZmMP0z7tIxdh/5FQPcwVt
xq1vpfPdo7P6chd3y3DLX3xE8ip0WhIE7K3HG/QQTJksDb2CiSz+A2Bz81DB
NNN7hdPyNHX8wPqifNKS8NhlsJis1dluyNkpf8TBSCO5BsycYD2reh4z2R96
AukgvnxBcP/D9nl4aOr0rPDXQkn6JZOucT3eVM+ilu35k4RcgsRb0q104Y/T
efjGbWSLgVpN4EYdvQgrEiiv2fZkGuFzpugmdD3QrEcMgwW5qih/lm4234VA
kY/LiQSx6d/msftPFrc4vnHs2ItCqsM1g/qOTe7im+UCgo6xVe6/ptfNasoW
m1zL3mnojGzZAlHLfqWDCgPJu8PwEneMMe2ShxOkfpyWfTSiYYRuoEsffega
ZnGkWAWISMEVRGH15ZKAYbLDvgX5qrKvw3ORL8iekFPnGuJ0IVPouKqdxW6o
dBKPx3aqdTziZ98RW3yJ/zZD232XgYD4Rmqw0OmRi0iVULj/NHX1GK0S2Ba9
d+PLScpT/9vx79MWwf4oTiieQqXcI9boTH9txOC1WjN8BmrhtWD3WI1ucZ7f
PrHeNzbuU3h7K8dSDqZq91+OszXOe7Qc3MJCDTXAUlEpC2mOZbOrdN+2Z5/O
h1SWbLlmYZu0Cdph5i8kzyXYYnWT8wpu0SJdHCyLpnz8VHtyTewNSA1712oj
MGW+8PW/ZS0YQXwCqS0RuFEmrgJWexEkYvmUWSdgJG/rms2xfhNwh7Ye4xcK
frKLicnnapqyTzZhytHO/OiK8+foln7ZlwKI0n81mwdBqR+BrrdIbF3ZKRUF
4IxP2KivLrWHjGZsiJUKIHrpPG4szZ18N/lrZtAnpNfx853H7kdYH/KAqPc4
j4VBi/5Ln77wzVfSwsgIvfPW9NO25IoGZ6TOv5DdZX9HtMbWSk7nf0dHdiEy
XTKqWKAJu5tvyCJNXN+DNSqzZktemyW+4r50oZiEKrmB/I+rd4DpDYIAL24m
Fc/9esT2yjBvUN6byD5DwyDn6jXmOdgfndDbCSSBRXD3XKVYuxK33R5nYodu
Ugse4BgJC9yTi9GFs5KTqRS14N6W7OlqxVDYGzhvzSxPTClL8JHCq2C8fl55
WVqo/Wygx2NVDB1g5OtVakp6zOAfG4/Aq6tVK6WeajYDXvzhoN9oACfHEKAa
VgfGz2fWqtsmpLV5VXNyq6E/Z7V9Wps0g8odZ+0CNPZbdEraMFNzNyTS7Pwi
VttdobquZUEfTr0GwlUV+C/RKIh6LwraXu+pY4afztT0TgdnyTE2oTzly4z/
rIxyK+21eY3ih1CI/+VqwiN9aHBckABNGM5T9YTZWplpgow+3jT0QSRk7ZWQ
+9dPWLZ82P3P+Lo2NId3LQMYuH6MFnhSqGgEn5ADlE+V+k7HYJvW6pO3XUwl
RtOKzOHWRlYkI9LlWHO+aWVGGsaLgkiRgTnUdFqf5kV3eimzrLQR2g+OTH4B
xccr7LQdFaSAIyA8gTnyMqWw3N7HvT6p/6fz86XmiwfUpisfLDZn7EEjXE8C
VIyLKV8cwey6RnsvytGSuT3vcWetrzXmgLHkz6tRjM91fGVrq1WwbiLzV3pG
qi7O8lA+M1SycfmYiFLl0pFiOLXxKJXgKGT2ERyRYnC8/JpbbDLtDJaD4F1Z
Lx7n4wK/dJauMFtQZ5ArCCwO13aYv6PqTsT3f5DwyzoKsJMfNBpx26DzAOX8
w7r9RcgO4x1oO8zhr8dD1WtwM6s3LOPFYS+VybD6qK8sH25t2yF9NZE2pk0H
sHAJRuwxDtHAkPuKDEd1orDVK0AxrKZrXaQilx4gcS2Z0AdGhachqg20LcgU
4vCe4ji9mq2oPdxl1Lqeanzztz98APNTrfLX3SrpjL64AQFBbcGRfzUji1c4
tuTaQ5nEtquWyf99Bi9sm5j5gHuq+Axsccymg9HwrG+zONgCjB6/AOGZFDQe
imhjIh1fT+Bhr2QMnK1dVg6mvd7Zp1ZLmpOypWxhZtapzoJ2OjrY5OrQ2HCB
8hMALZXeRRu16GBiXmWYBFlmmlrG6fsFZDc/ZuonsSggwH36MNWRyDaN3JCZ
9Wm68wMQQ5K9/m4Y/qeypQcbtt+7CruWlu1ECFiJJ0Ma4ZyCbN9PCw6YTtIZ
bX20nqfdoM5CdsBRec2O3bHFhl6PDrIvORUWAfEm/0AP3nAn6FtgUBO/sbLz
YVBONgQ0nK7hLin5aw2PzV6c7ST69A+vngUf7I37k/cnPXtIJFT19fOKWxcA
RRoTZpxif7ZQ4C+nciw7mCKKzLUO1dtkEgz3TWAoCXFMCkezxZGX28XQI85U
6p6CrTMQdJa3/lPZR83AGewyPNzG5z73Em99WHp8T+noZnoy/xuB5/WD0QNW
ZOdSra/cb9hRivNgOhZJw4uvPBcMDen6k7PjKaRrUeWJTAQjlTeLyVRtKlmj
d14vOVfQqS1f8XfVFKFcAvnovrQjJDybaLMFn4EN7fAr1mtSTPWgqyXahafB
R4FEs/UxvRIr+m14UZJ4M4q5jOQjbgMkitz0Mq57UszjI3Ji7Angnsh2oxj4
WocrC7Ha8NRui2OSO0mE3qihn8eU5qtjL+E4H6faWjylsuH2eHsAR3NuJpe3
dxwh3dF3BR+oZr5QLtatrkZsBhMsvKrWyE54IjUa2TqWMUUSas+BLs/bYh48
qNjv2TzdMbaVR81g27Lf1VpwtHli4ifizd2tZHgfF+iXCwxbpkLdjzFVSkiI
unDkKP04cASbiV4JiPs0jnGmMuIlejtpEb1+VxcPDrS8wCVIOL1H+hfvfh5d
otQjVpiBIYHiqptGndUpreR+RXh7enPN9BJse91cB9ldMTNCUiFMPdpOZyvm
HtSwgiLf617Oh1NEAXSgFmYP07eQxnGA4S+rYds48euCygfekCXbZeigsZjK
mAA99b/G2sokg2jU3SIUFjxnZfOBep+4NhxroIz74Ec6SIsgaIeGUaQejFUX
nrBDC/chkmDyYSlN1w7YuVizrLyCxae6uvI4CoSb2ptpjuwdCJe7uCtHvyHY
gz7X9ZezHFSgZhQOphmXRGqnRANCC2XP9dgloeX+B+WC4a/tpaCWY9ygcBwr
fqrmDKoRriacM1gqeaVU2dVJBg02/2w654SCMuwZwtzFuACwz4UUUYBYhzta
W6w6fyKCojs=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1Ix9YjjJEunnLJ1P8w1LTIUO71d7dWqV3IV3j4pWRJD6YgaEEdrcLkm1XHlhTIwo+H5wKmJoMuAkjjC7EypIW/AeSoJ+4PZ5vJ0J7MGRAseRuw5Dlfmn1AOLovNao6yThF7bCkg4TuDB7klWpehvzJwqLvZG1KitHKUILeXV5Sa/mK55xqVxBIJOBoogB/9dINbNySq3C/EBzFLsAL7nKj/HX7dK8n6CCrV8BMeU4ACEPr+4TzfQzuymt2CH9iO53GMGBYvHTXClHEEs616+XJx5IOr6JNnJh07/SinpCGDl5x/kbZ1KLpQJMzdwKiR2FmE6yMEbkG5MLpnuMC1EostZAPo9PhPyIGfZ4BN1HDBDN+cAQsmxiTNgGSW6SlKwCFzl39OwMGgPbH0iXU5JzHNt1GY7OAcG+ZSdAUJXAtCTor9H3Pi3T8N/LLrBEDDmBG+8c+8SM5azSiJpy56dsNl1/JM3x80nUjhS+EkeXjGlf/IWEqwxu3/kaCCNvCLddJKPA4gjYgLgUJVHW+svSGOImamLTN3PbHwM5OoWb1iSsMcRum2Uxt1DaBj2lJ8G6Gaegk7k+NxhP9hu5yVppiivZeDsx4yb5EFlLeUTF0gIbNb0QAA1SsH0CtIYyzsOI0eA4uixj6NpN9p+WGTuew4529o9MNv2VY1HIcD9llmwKqtOW81qliB7FHHv4B2wjE8OYLCzhXWiNNaARICihPxkAQwGHLbs11ujqdQgJoUwN56CpSfOSDVHal9Z2pHpP3ot0QrvcZTPvKnn5plG0+c"
`endif