// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uGOLSQZ0NBkLmjXenYFu23dsAaaj31qWh3AyJFPm6PDFkFfTb/Puz7FBN5r4
EYaux5UGEqxRtmeI/SAG1WXvlF2QyiCXJFvAYIR+Bo/dm+G1olGynonsu13h
+MQrvJlGhN7ihJVtSMJEnYrkUeQf9zNfU3e6009qfjnfNmpxCns6AwGzVMrp
bnk70eWprFWeIA50pM0Sp4hpZmdCcUaioStILwQoKQbRSKStDqOgim59DuKZ
2Q2Ovi3jmo7xiea3Y0OpWeTfal/6nVxhr97ACrbRaZtcgXMfrZjHfcRsJZH/
U5bTiL0pxZD2XULDRCWNIz/sSZ56D9eQnSfHiCE6/A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qzQ+5ts0I0HHhbIVDQAKnnP8gulOLItXOlwrAjQGN7CXj+d+DA/2OqngK7Yb
riqtCT537HE+LlhZVPUNmi6yZRQVt1xMYXTIkB/FJgFZlVqOXo5fT4y4RhFC
3AwEoG8musYjtenyoyW2VmmSqVYLCit6EVv22XSq+GA8NGxycGN+jRZRx9bs
reU0mxWwb3j5BvLuVOnZ7MaT3JCcw/8qvuaZ/KmSmmv1nUv3HiDxq68CSUer
KDMeB+pdn90YnQgahjgyNveNGt/FV7F3hgtIIpNC95QADR/VShHcnuexznSs
JKcKnjQWbk94OPzXnbHzI61bc7yZOWalkg3jRJVAdw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
unuaZ51acqg7ecLiTJhsIQrk1otSn59tco9oTmXAMatuduGhanSrBI+qqtUk
JnAmsB0XKfl6eqMZso/FRSGzdecSPhPWy8G7fpPzsjD5PAHt2hGYOz/KT1v3
X+jE7dQ2++dTkBnvCCkpk0HnvDkCPT8ARYc5omThuu1b/yifmhmuYcGKEWt+
LN/a7O0ceMLQsBG3jTzx7esXKqhaF7cjejzuxze+LtCZxCwe+gtJ30cWLVv9
XZED3nCIC1S0cYqQIqiABl7HaWJ3Ni7UyN5YMO4tuirt6QigE+gbWO0czRE1
y58ubfCHC6HklpP4K+mm1AcSv4tIJQIKIY78+lU01Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qUJzKEQQAmBTlkl3JTMCLzeSkC+XyGRXy46eE4GWk261tJO4MHYJjk6WHgun
giri1I+TcshJzoCyF9+FqOEQ5P9UvxUSkA9mHJsDy/jqWBce5QsCgjiEqEje
LNwU+Wt7Jd4Ikexyvky8yhNoXbIMY9KjWIu1o+goVXz5K7BSxM1uUMFfeVqX
wrOySfXYxD93kErx3x0vdq81lF6aMpCKcCzWSlO5UOZyB011SfNvnjldiWoM
M9HZIzQcA4J3Eu9OTiMy5PBxyuO519ymG7QKV2m4GpRhpAjuAqIR65Z+aG3B
3/S/4fHQTrGLrtaNTm73rWzUb89wm/PaMcu/KnoKkw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iA+wH5HlmmGU+EfeGSM3VlLSh5/AgR9aAkdtKXHd14dqB0FsR/GMmcM7NYC3
jqD8Aqkg8BqNGI6XXikccpfeEMno0teROUPF+3TC5iQTMt8S3tXHmMnqoFkK
saGY2eza36mSeesUUUF036LVxs05jo7aR93cxQ1esX757zV9f0c=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DN5OukqUl+Sq/qtkrmyvGUPM2xQj/mO7BzFNt2bSV4n7EtG+w3UeE3pmE89V
Kzvlq3ULboE3CgpYlk6Y0/NT6tDzLu/qGwZzUt5guLzR0dpmv8SpdCpgpZus
S8uA97YyJ0CwogvO0e1hbfDsv0a8ttUjtpdPwbkZh3M8Hec7GaxcByA71OzJ
MfjZieKuqGP1gLuujbB3LYQHFrDx2y6KorGQQS7GlPLqZp8tAFrwehtsQLMn
y45j1k6aCNhaoyF2thWEaAC7f7ujOjTPI0wCpVIUVVu5JcQmSI8YcZ5heR1s
/9WOBIQ2KP8gtY5gAzI18V4MBDHEF+CB/jJpt4Ai02uP1PnXFVnVPwnGzAFx
ojiJBbNuRqzDe38g7KlBzPDdkb06MPcKj5HDQNhEgFyFZnaLfwPNEjmbRAPt
cYF5uyAiCpW8rVKRJ9AueJNpVybeUMiXFOAXlkEn6d0pjXH6HK1n0Uu5ydQH
dpKMbs8nJb4BYtJKql0Lq5hi2IIcodc5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
odukEHf6K3uwl47EBRrjkYV573HZKrBFgrOKOMrFruhq4iLmktbMmlJ4dqbN
2xd1XByc5c3xQGtDLzXukjRvxX/zRyVThosJPEfyf86+zeluBaJEJ0n1SM2s
LCKtBtaRhmr52+EfbGcd1qa2OFWV9LxLjXHW3G1lBCPoFmcmFp8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rvVb17T42e2hdaDjtB6gEbBrbqUPpvY++199jZ4g4yvGub35pI2oOwIbw/DR
uQSTciZQopwnyjawDMauKgXEV1tWr/9lNxV4zsUk8fyq1Fqc3NNjxAfilzqa
Yb/kHDhK/TJw1myCYbSp/eWIv7fSZzxRFS2V8RN+CxTspMI3BRY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 66784)
`pragma protect data_block
Z+Bwlx2u49WdzwyGG9SEnxm0NuJbTxmN2eALJm2Nsswzkuwd1AyNfkravJ3s
7BRbevfXsqQQvHkdu65a7PuLeqgznO52fly+oMK9G4BKN+FZgAM5px2FRzzC
vCIS1x0VSajHPseuPUOQbm6Wl2Za0YXlQIsSrwmnGWAOIlIxuk5xHSAu2z/s
rhYfz+cG0iXeKZUGIf2AyvsrVcoyzoNMBHZwfQ2mscgKHKNqCG8h0lg0FtKo
Z8pRieHS+XaydRjlsnm1do5MEuDnHYyNZ3JFBd4AuS/P5kVc5sy0imJrv19x
X8q5iuNGKibwRM1B1EDblR8+SbOdIT0OWeM15dJGZCeqNcV0LDDXu4GD6Wy6
By/3KqaS5bmVngjUHWEE3c0jKZ52JOEEay3NzHRDNUACwTGee8fEk8BQv6In
DjpZxyljA2jJ3woG0UjtPpw6xKMaSMrSBOI51qMz3ANNo0GgOUmSr0ue7TZy
9v5S+NC3V6+UnpWsLBYRnr56vumnHP/cdcNFybwxo1ll03isxZ/M/GS1mdh+
G/SJ8JIbLyr4nAXGZKM37rlhhvORaXVR2FLMmB6yUdx2Wz7OmqaYDRQ/kV1/
SVuQnlPu8e8reNB4pFaN86quYUY986Y0w9uQCCMSW2R5f0TFOjb8SI2br1Wf
HeNdgl2BAh/hGDgKU/QwwIqd0YlNSQCGTucw/guylD4aLjJuz8Z1Bh3cjgOc
On/NIJONZ8dMJ3HspQmDLJVegmXxC1ETuX3LwShttr2gf0faNcGdFgxAA4Su
bfOoP3gfLTAKqvrF9SyWigS9Z+i1sAiG1gP3TqjKSsVqAXgLIMrC9beW1GUL
sAOB3gTccLoYOBzP/7eDqRCL/g771bbV/BirpzInViGo8d0D6J7OLXcK91/z
eakCHcQttWQdAG5Pi1xXsM7GmYAw0F5AUHDG1RnVEhGkB0Sprf6AqzlfaH9G
lfcZ6kqit7Wd0IATAoZn07C4bKCtp8zXC3YghKMZFbtiz8gDyXFrYSZ9fo/x
5jbnaObiJidkNw8/Vs9AgdlkNbyvw9WRU9wSWlezaxo8qh0g/xoFmWWXqe6a
yk1ju05EuEPD66u2eL6DNdgJTj8PIiCtRI4XNNexZbqlPHuJfYwF4crUqKww
Cdsmhe5+wIEHtSxFWKP0Rqmafb311UInfHZ2OkFwNvom5kLLx8aFBroC7SsS
BnqKJ0KDIN0G1wxk5vjTl+HUY5JUUX74MXTPv2obJFYRnzBKSMmNJpoEMKW7
/5e2C1T3Qclo0gQac617WelEoPd8KyCOjXhJ8fkMxtCBGo33/ObVxa8TZxmF
BBaGBAbh04N+auOuSuln6wjm6j5CtkZt6vxU8FoTTpm6NopsxhnnJGvOSDko
uRAMhkMrtR8VXDK/eAs2apsfrOQa9Q/WZeV1g5k9Tp4gJdEFisHmjBghvPM2
pALAMjXllQ5PIcZD7JcJBdZyqLw6GGDXcbnwXyxl0m0suLqnrzSXpskYhnuT
yxO97MTaG1u5xihWDVxekmaZz0IwLXjWsPHne0cj6WFANSPJRThOeTD+jqJL
YWXX5firF9uDeKX+KF0q96aciLAMj2isOsCXHnPwL1v+GjFx3uhiZ/QGIfq7
y9Fm2pjVuFGrA7VLx4EaIO3A9OE3pHT2FNgaw27r9tgIXTXGwz++Ig/0gDeD
frJv/2eWCZD+w1SLJZicCJtTZSt6av+uGxN/Tdgt1YZorqXiCsmpwkK91jsL
6nxH99X/f2gkH91xIm0fuOo+spYqu9dY5C/LvJ3iJPN7NFrKjZXc2SLBrk53
76lNwc4qdGRMqzkf3g9eVK6/sAWl6Qkg7tU73q2/uyWpg3zPfM4IFLUUPSCk
I/GZIVQSRurx184P7u+XUNJ2Zv7jqVd284Hq4rQfeO+NJ8pIPcwpJatnybTk
6iAZCnqiZWPmbHl4z5cU7qz06D8LCG7okv5SvA0c+bMz70CsSDZVG+lQiAP8
9vojzEenFmv1p8msfWyTUNTMBMDDvAGjYeOuiJxxFDnj92qtLWOmS8rllyHx
poXy1yrO33ieA4LbX1NB28ufup/Wpwtl8ViP13sSRPI7atOOE/bIEpMzaiGn
Qb1AqYqvn80TmgOQaEoG7/+4lHeOYAv33vUaKulWnrcdaySzPBezoW5JHFoB
rf1uEsMVOxNUFHbp3S8bPBGyLjzX2BCE937kP4Imwv9+2ELDIKl4YTx6FSrG
sJLPFbWSSJcjJxCWDFjbatF+Bpeh3UrChOhdOPC1fzXOuVqzQR9FfzlEMRJf
hOiGQ2AOo+DMglhwdEOREwWhLHlFv6t4oCZokRRi7Uu285pDxGIlUzD30WkC
SLQ/FEMgo1luEli8xoFlcNOMVYMBcZdM3PO7UK0yuBWTTI+KIIENEL23KZGj
8NzXM4VrT/oj4UEGpUJ7EiMwXoCaJYQcBbcns2vy4b5ubnKL1wz0fE/8jp1E
fwEZOzpedmnStg7WrzoAq17Njq77aQrGHKNX12pBZlORmCA4Q2nSxZHb+Ot2
EyA50DVD44kqbfQ+E12aYuyaePvQHsVDrJRUoK5tK3WN5wx5mOESNnuMc2iN
mmrNXi1IndNym9RiJu8mMz+Zc8wnFTp7w09Z4cs+jVgMGP8RF8Xi+aIzhEsP
nNa8XEw6eS2NWWj42jn7KMv0vKmMjGKf301U9XchYv/xZoy3t5t1KDuXC/ei
rlGsuDiSjUp7jle53AY0XsfVxPXi4AlSafI4bgAwcx1sbC0TVryeWgU0as7j
E86xYbFC6rsODi8whfebv/I3sHouwxDsAWKW4suEmzLJ5DhjBB/IyIuF7uML
t2BN4b0yEibKuE+4Of3LweWsrUZCmyGerrXU54RagR0nGfdtwtZzZssXqwbS
31+MXz4ZvHIX+baFYrmK8aRBUEqUbekEcByBsum/5nVMuDnwdmlLwvyHkZpW
ZHhl/gee9J6vlhbJO0LJ8/3dCvskAlFYaNQTZrK/vPdyR6Cpbmaw+JjOMUgz
IFmhE8Hjq2hcbVHADabFGfHbktEgTLMVD2IVrHI7Stq45Hflws+NaKiNtgdX
GODR7+Wd0NYH3v1LKSmD7YbwgxeSKMo0eYmHSDNYKP2Zwp2hoVO4sk8Jq5yE
8N02KXc7afPpDhL4fYjwytboIPKLwrd2N2UgVYEhX2qEsvzfjvBu6dmqorZb
dzvX9TSmFJiKR+csr8jKCusaJlE0yxA7Frn+5wr1ThLpBmpv7jOkAhtvSCg0
DFTYk+L/iH+BTaBSEzRwDrvjJapNmklNuIipZbKjizJhgLLCoAqGyk8M6ll9
Gh8DzSJZy+USE/D1zxylyjKnDnlhm2simn/81Lo4x84CW9KzqQfwz55WmaNJ
P1QnYFODTtiHDTCYUrbTeAlTkBTxMS/zmh9tpldIWQroSk2GcewohWJ+2ZY8
eCv1/GytM6iktPDuX1987SZv9QxEAq8IpzKLgoEZL3FkKs3/gmGQ9FV/nUnJ
+7lA+mMYyNfux4S7LERpG6sjHgOz3eCTwRUajrdRtHJ/lWO7v3cJAOEfLc4u
5M8W1saWvtkfNVO0TLYBTCpECxUbQPtwQ/lXwDNAM1kmcJG3ffjUHeiJv80w
uQb8h90ziqU3kLJSgXdisPbclC1YkdIe2I9Gu9pOv1mQBOx13Yv5USSiUDpS
XPI+0bD9PVJwDDVchx0HrdRtCBOPGwo3F8z+8x8JqF34kyCffpsBj+Jsf2qn
KXTefENplEj1AvSrBo21DutDcaVjGDFHIysWnXYSpmAL3xQ9ZGu1DIJi0P59
lmFXjaj7MHY7Igy2vNQ3aDlMPLoj4DKuTTT+6zIGfRc4agvpM4d4Y3UzWkzV
ToPO1vIO+7rrmCD0OIKD/orLL3KEnn1oeojKsrW3+dN0abouPAgeRimNs5dK
nZKh0y0tpcIQPHpAvVIbWNC0Ghv/5JYHjBX60bTgAvOkZ+oFrd29GBUbr8nX
LTjiqo+q2kwbT18turyT/mJykZJPOlOymtgeTR9hpPeRcbD0sQoskFmCuH++
rQfsOGwwsF1A4qbcoWvH8v/IVecJynQmNPypIqhlpvCX6+++K4Lb97EXdSYl
xP9T7FqqwpBChoyIyZMiY3jEwWdR7QgfjNUhpOXri/yjL9tBLQM6YsS8xuOp
3f2tp148sTc/iuMNQNujapBQNF4tt5GPU2BMPKM2bmyA1hZQZp36BcTZSBgR
eZyKoycFzIPO5hZ/GCt+NffliLRs5Xa87tnaWjxn4GxpBh/A5NYEa65dHIWf
r0ASaWcfIlVzYwhJcA9ZtKMHCrvCUiitMkKRAbCSyJvTBJ9lNFJQ7iG5e7Fr
nhpKvT+DJKZ7y5GEyqkvn9QYAz/TUd0K7K1Kjr7Tf+hS/a/AxJvw9IOa6P78
TZOBSDYPK3SLJD+E7Iy6b2fQ+n/zADkoMLs5HdDlUKFAs+wIpqaAdCLcQT4L
HRcJw6IADU5fB6dvadBQV3S9OSgWAblN6ItILzch4yjnewySXZxmwJvd7dTc
H6P1PPZhE+tERLdtgIjbsTKOu9MRhoZC7cAkmmTCnygQQNAuGKgmQZaOcCot
wL9ImveX+R9hlWdZaQ7xd6S9r4StWCLdidbqnkRUWzQFuCT8/v9m16ko+JAc
8q1LKMcgWlWvDc51NT3knHWc6SdWBM1apIX5E/X5/ETWvErS0rJKAbB78Hxu
nTFcANKF8lxdrNY4afNfZ12fil20sc48jTCMPhNrgIBqujKxKBk9hY3rnrYE
YNBH+H3DX2xreZTkOh4GtM5xZiyApNpd6WtUZytS7YVMj4PO4OmA04o8QPxl
LiLzdrkWvRK5feoMgN8s3Q/PrONgrdVxNdblT9XByvkZ+/GqdtdBfRTQSQvz
0NKRZr4jpuYaywmayzUtM/c8xYWW1nG2oUMfL3utFsU/57jCSR9Pt9pT1T+W
DO9LK108ioBLvl8zD26Djxj5D0/AVolOkzD3N/765ZQf5iomtoNrB+md6OQS
BWyRdmeRj05i9+ESnjQK4936d19wdMqX7d/oDMKHoOo4rlnPjlReP3ixlaT0
axhfKbe+eyyzX9l6/L7Gnq+XPHv84j4KKMLEkq/ASFtt/2ErqY6cf0fsYOdW
B/5w3B6eMJfnvOHNiAUrdo3HoH+PrdWs2fH94tpmEQOmrBYjjDtbCbyZfGeJ
vZVuZAFL7RAw70spDVjo9/TxRgcv+myOJOQLx2WxcyxK0CNoJtDKik9HVOph
49wzw1aqKUEaBbmEFSquDG9yp85sgVnzeXAxkuEIyc7/RI+avcCsGA0yfIQn
Ds0FhLcGVAQQ6iw74XFc3bRSOpOwEeyhapVWy0e82JjZGsCq0bOoySvXOMOV
qT/3KwbTwCVpqSUM1T9EnCjPXvPD8B91HOSeSbSN13Nvk7Vgacrps6AVUKaZ
PBwzKWWyHTP11GJyK/1AA91UOifFqOZbqGSNxDLWN9iZbKnTvQhCj1z/8fpC
aJs69Jqelfq00UPpzsHJwNEBHydqRNiuE5BSf8bB0nY/Mqf7XSedQnhU78Ul
5O/vZl9TTh6P1k7N/Aix7ck2vJzXHKk/CPpf93F36prb5z6i89B17oXZFz1P
7P3m1xIbDE+GO3dIzb3wy9o5A4fJ/pd7kSd8KdLASmdZKmsI/oVDDUUYzDga
wIeM8GR0SeviekRyttvMU/UnHBYWV7BZYSnBOypxr4WqAo6JRxb+eERzWhza
pg+nUf7WQYEkVgJ/Cb7ZMIsVqm5NeMEpxic4wVJfcY0KQ6jxYgc/xqHfGSOL
LFGrekqzTu+4gQeD1KPDO33seW3BRm+583b4FhUSbOqmCVFT/01ZJdQFyAqf
rgZTxegn8DXQ/1kARkHIL38jSWjoXGaoVpbAnD6Lka9/FGn8BfFQPUHrsGWp
aLKT4x2AbimRmGytOcGz0vjjoAc3EXMpq0i6PkigS1UzEwuB6XwDq7b0Yvxv
p8YlfG4cpTqF16U/5B9fnsLcqwHYNrwVGv4ybO/QA2gWQOPor4TYW7Pmtd6u
wN+5wFCPouxfJWjXokYN12XjmBT/zoa2v+FJ/sGAeArZe16kpzGS8r/On4mh
WJOITBcig3kDeeDejw+QSNxBrumD/QLUvcySKJ5xGJzzlBnYEb7FXaEfeQ3g
vEEb0xUYcYchDOFrDt8fxLs/lKQPWibbYufJ/soo6DoT9YAVjO4PJZAab4lT
G8R1cHtLhRK1TvOSwxBoaaRe66RVcPXVFhgLD547lF+Y5KFt31OOC/VkRP0e
OCmYQLIdnvIFdpqJuq20kLi4v13qpqokE8/auF3KBBKbbnjYS7NvJoA/fHmx
TExuURI0RYcHT55tIRifqZWsYQp7b61tkz8WwN6iL7v705GzwWM9OaRHnxuG
5twHldpvA1CdjBtfbwYrwQxTpoguhTowfiTi8xonRbyeE8anaaWzpxguDn5u
gC6/CUqc1FQRaQjge3+LxOyDfmv3Qf2iiBRoFdDnyr3wHsGal+xCteBhVmJF
++qhhgYfAHIm30y5shCvthBSabsVrUHiXoL3DDfTyw2eqVm7XF8SLCBmm33o
RihSTJQjdEdydlLKREguzTJOnrU+iGCnY5o/+L4x/9j27gVHYzgZ4ax4uP2c
m6ne+lcEGKdNoQ9sP1AC1sQ1r74ZK9ZofAwlT9g9tM9iCeh26PoW2FCIWOJR
qHLwi8t+nFN3f9QZijiDnS8b6kkXmP7+VseA0tiJV4n91gZPdemwhTdEQvB6
Is6WnvYPqC7Lkf6Ej31CkHCbnqwj7zC7Z8h5XXmAW2YPAT9Qp2vXQf5GYnq9
o+TtdrLsYdBe2IrB6wrPpnwFFGD+nGgdlsYi+sSdRN+fMicE6wLLHthpJxRw
+WCKt4n1Qsoi/4BJA2QLQwuzhC8QxlPd8Ip92JD1orDOTM7uXaju7xm7IztU
HiLz3ZS+qZgG/tEWuhsppWLLzqNFdvqJ1s0ETEcSoldBRIwsD747bEwNxPB/
/VccpxOvX5DW/YwLMQSeZ7olRaTy/9NmIz3ITX4q+5vrWbCByIKCq3zXnSnN
O+hchy1tvZxDlvP+9TpVNKqO3RhjsKTql7sQloeEU7f8fPhuo6iFYW/GnZ2k
GkCrAY1m6SzBNIp0nl6DgPAYTM5pfO1cY8QSkgZ6wUXxadHpt4ZpHku/Up2C
TbeFvtvqjNSJF2b+XKXG4f3EvTRU02MyijG9eLc0SQ8YYD+5ZZuCZKhI1gR4
vouuoZMI6UJxwr8G+qfsRiOSksoFAAQr70bXXwDfCnTcuEiw0140l4Lly72r
m70N3rCT7Eu6Nv+Qzy2RkriqsXFkG7iI3RzT5y6lpuNCD83R/YXtq2Vi6Mta
c9lQy1RziRsBsobqgZrO26Y/8y5tZMdI+KCvlGVWYg4mxir0dY5vSNJSDog1
EM8Y/VNlxao6w3GGijCtXT3b08KpmhvXRfcKT7bWYSpQwTmVd9crq9lUsN6S
Tr/wD8+H2kzunD716Sf03JzCxHMdu9SyTsOTRWunGuuVcHxpWm/SdsJJV9Tx
ZyoqRmV9V+tRc2pd8oB8lVR6QImqzdViMt8tSvo1xhpRV39NhlC5eRCsudmN
ybgaFCv3ixP04nnSDnj6jxqYQgf0/PO0OA8ezWZ/QIuzfx77aC3wevLaaUJF
tTanrs+SVLLSey4cgWcpVPZnSlfj1pIozerexw5pGNDO6TlcST1jpzokUfBm
3KiffJkPTht0ggnozlPIYZu7eeFdo9Nn7ThQxd9rwESWceekWXKCx6rQKmpf
LeVfK+91rtzxjIbdwiNPA/KY16FkrnJs/WroYXNM5yRo4qa2MSGn05jTeZsV
M3UWS7tj5YMETTDwew5zEQKMbnNVTb4uLT0ixohctCPEAh5ve0uhJkyVuNnP
lo5c8KhzHWWB/RsUCpctzNf4pMXPexAOWwYP5tfV+zriNhaqvNRGuvyd5SBF
te2l6OAUK5eAN6hY6bctRNeMCdtrwNZkc+nXd7dfg6cZPw79/GwVV1EzZVh+
NK56cESjKRYXSk5CQPODqSUeitqzBLcjvJVCosV4f3zzjzYI3fn19zej4tKp
YEopolzOV7qi79InjQe6qA+SMHS2VLiWi8ykaRD23sZ6sGeZpdzZCTnsg8Yp
0Seju5d8xKfUa1oH5un+IYAUFXTM5Sn4tu6dU3la+GmZz/ouS8KfCcJ+7sFJ
3ukQBEs45xC9IKyyKKnzFDE09nXbZ7Rau9Btfq85S3Li9jofoBq0tDmUrUid
joAiz3PV7tXH1AgQSaAZEVqbNaWk8OtuxOmhYgAz8PmpwknaueiGpqdj94Vl
5/rwZ5WGKrvpIUNc4x73bnV7Sg1H+L4JOHTjOk0rxSZ+PgUVRoa/nqZ2dVhD
vjucKp2pjDOwpktExiq/YxhZEtVnUUzyqVeza9dNzOjmyRX6YjWd8vKkFlEO
CsNrdZId1ziTZl+S2WAtP8U5TmQ364Z/3zlblZqXhKyOaV4wrCtEptKc2NXs
fNjKmGXx+0NWmPQyYG1Q6cKBS+HaX4ZuO/Emc0oa4tKy9iUFPpkXJK9GXCLM
Kk66IPwAQRmhyvVIzw6zohhN8UnGeEAcSM1bL5AVI3+RNd2wty70a3jtqAAi
xrfHCfPA2ftXsBjalg2+gPtm1xip1aGQhTl7DMWmv2+qvvv6C3AJWjtc3RkW
r6dpFa8SHp7SMtRnKb8if26xeNMP7XQD0UlCj+xKi5EyU5KdKLKAkRWc5JH7
78CqoTRmSzhX3WGTQDKVi0mgo8jcQqtgR5xDjLr/nmMJUxbE1j3T1ZPs1Lho
z2J+8F36IB6OcOeZMz/ffAxKL86F0kWLG4fLtkuRMrU2XWqhq3QadlVFJUeY
mUqsW3fv4J4QdIrLkTkJaVz7YZwo+gkD4cra/l973AZhgb79m7PuMJs6l/ZB
ebnXUss72V6Xd3T8R/a5bO6vjiU+gpMtQj/vXEOITvzB+YqRv68vZ6CfCT3j
4l19+fPlPgnaODBajtlnZmy5NwUsSkOWUSD1b7jxahTL5u57GDA7o6rXyAzx
MAT2W+YOhxxLnxUAJ28OtJKrkh5Aua7+5ony8QosnRwY5ZjG86Y7mVxvJAG8
cxLyShpsyOj43mjxJzWTiTcSpD1w9JSVpPeubrnD3kLNTofJMIQuuyiYX1L1
/EnZGu7P+JNexEI73dF/TmNZoydqui2bE9iq2eC+mSdIpCzKW1RK+YnxZsHA
PWEYUwyl8Kxo0Zn9kL3m+hmKRjN4P6I/gavK4HEIP7fd8esmPrCwdBz21+Cr
B7zyETSjbXVq2BUmMmv0LqlTB+tD1PtC4cheZ3t36kGkJeNJhdLGyUa+hRX9
gyD4fcR7Hernu1EztAaXgNr9ZWvO8F41oIzcQ2eNb08SR7LF12Y9l6aw0IgY
LRs5bCGNv6fZcZv0tpY3W6c6fBz3G00tDDW/tCG5BAQUNnHpZCsfEcRdpkuh
JC3xdCMcHsARleb7bo/fJMqYxNYwPZ5nQe6xjGMKmKaTsNWiT+Exzj9wyFJk
L+rn/qzbykXllV0WNOGIhiuBjWmL3fDLIFkn6oQ3dRgz0TC9sgBYUZYBZuoh
5P/RglHsSth9nNFm3/+IFldMD5LoIsL7yNG2uGG2l6psIkXIK3M6Ugn0jIPX
0NmTNNAFjCzbvXvs63Owv93KWc+XsiKmI+mohsmO/BE1/Uy+ho7zkxikUsDr
n5eBBN92jfnwHFDfPAvUCgXmRdoRZTJT+3zl7xpKgba1kMRsJqCKSQLQSTr+
HgawGW++fV01a0PRCquT0vdmJmcGZBEDUMV6BKKh6NJEl0KVvTrILEMxy92z
hoHlo0DkE8LL/mrhHokuwL9EL8ObUwMmeSGXzEIV4ipS7rzjTuaVK6d1nNff
/cphBJgXJc0F4yIJrQbrocAwKAiMiJVzUqsrK8ppMeDQCcJRYvLTaYaLwDyq
ZBgdrHX/xWQKWuAajdSJE+DUpF4cCOC5NondWIMOD+hJKPcvouHLWArtAmlf
kBIQr6cd5EUzBHkTq9z0SP92xmV3uBrDTvNxIzkHgsBU5ZHRS8+rYf7TDAGr
JzLn9jExAjSA4LmonDrQdkXCLq4wz6CCKTxrGiZtSZdozO8sfsVvJC9t64aD
1j5yeVRja47vsme4oFyM1Zk/KR8Va81X8kFQnu9jx9lFyreAAFaR+25r9LtM
GrlDxALywLsUN6hBZUlvbIi2f91FS2N4Acm9sPD1eq5FAm7xP2RYTr9pE9Hi
bMJdb4edz2j2iPRYHT0RbMcVgBs9iauBei3eWox5fWf9qFNB2lfUgbLBrGZM
IUVix/zCBPbS5f0yryrLR6DqEE9KAJs3avJ3uqB70A4Q6DCZ2s381vC1DJNd
orbPBsbudtCBu55A3NqB2s2HU+yvmCBHKsg6JwNrBnLiU91erA1ZfjlgmZTi
fIxhCpymPWEnnorPWJ0CKcHE9+PfSvz0RqgDPAMHLhIixibxhpoKTKnCSu3u
+35Og2TVpIIYw4xoASxULBjhCl4GLpDbwJzACWGmLYfOE8dlyJVIGveiqB2k
B/rAhu/7dBb/OwDesgkE+Q+WB1PJAFSBPNkY4zbgYPFeghpt1sYq7aLk9cfc
6lp4zp5pQKlFfDsHB3aQVbbjwvJQxv8MfyKBnjBaf+QQ8vztUzriI+NrJPpa
39QDr94XUhOqKCsxujtNtSeXIqq9oTEcVWWzn4K1cCtoocsEtJaNIlFVDILg
PFq8DNxcCjcNpbdhNG9Hgifiefj2n+yxFqNlrbc9x2YbM/s990WkxLM39Hu5
M85U47MnWDQy0ml1Jab205ZW6v9VlneMGxO99WnzszOxPmfGrmhUc3jUWkSa
UL5+9Vw07C0tNZOQCwnMgv9/cKsoCbE/Nf/72w90eKqZkAjSymPVNWRcYf9B
4jc+pRsgGHI/n1qiqN0TiZziqtM6lmzEZDw89Xf70SWr+hNMw1p1G0mdTwKo
mUnCzb3NumWXkqz1f7f3YJeO1f/hAgJfsmqkrFannqT5+B411NWa5uj0X7Dk
pG53IUe/U94a6dp6LjKJNCB2SqTUXXpQ6uQSzPx9OsyuTAudiq+9meOaY6G4
9cuH6BRqGxTB7MafrtEq09EEqXnChIV06meliTaJAlKUhNjrmzxE+goyrtK/
NCYuSZB49f0uYG/AH4QZQntFzQf2zijO1qYVrNOvr783izKA16uiW3XUqnyc
Pyr/P89gYRwaK5LJ+3LRvcG+YjxihovvTneBRZOgYjIVx6pzasVFr04/CDAo
fzL6fg9rFon+Ml4vntgiUqBjD1N4qsT0Mg0Len93CLdSt/BTdWtTPWjtvLCY
HNTFQQDViDR8vQs/Tt1alyazQLPY+ZLD0sGsABz/tVjtZYcLWWtpIkyOpSBq
jN3Ye3E0As2+vdQVU9gk1CCJfSpi/llr9S3Yo2fWY7R7a9Y4oxMYw6/XS3wp
ic7+OUed+R4kyqAkMTLTV8nkzL6GNAXzdtaIv4fOYd/+TaCWfWqHcwDOI2gH
HWNVmjQc6puT7sV28vKUSn8yrdWUBgJ7+SO/vK4f4rHnNNTZvBm1OHzMeugq
Ufdya/3shfZMckmfV+ZYptsKCYj6UQx+2+dgweXTutGKBF19VOBA0LIZzPuI
9h7d1uEt0impIlMh02oPU7hQzjaIjKZh8dmY2aasci8vDUWfY80VGT1n1OTz
Mbra059Y05gSOnuzULPiqDr2bfa24WCeQ/WdQMd0OsPb8s3sxjMnQKlRzGjr
StzRdXZLiP5QGiOCGStN1sSOWINHBm18ftvpUhLL2aIPASRybJRe+7INxlDo
ZKzko+nrfiUtUwN/UicgDQRGBbxxbi8RDHLKmjG+bdR5+VhARVEvqnUB3NzK
kw/qZzxFuvyGhNBAk+1eC5JrVLsSSzSwbRP/2MfPd8Y53Om3IvbzOaCeNg1U
PFErqe7B3f3Ki2hiuPfSget01RJhY/XfQjczgdCHp1RqQrc7PWvCI6tLE7bL
tMzQ1lGDk+DwnOjTvYOu0jsE1uiBfWlZjK7ou+NPvopG6eJnoL19jnUqzagq
AvyNvjAy2Qk4nISRk/rWdmF1fz2Zdg3SQhWqvT0IQ1gQBLxA6+g+Wb1rTcC9
mEug2FaYtLD8LmkD737i6MeHoWPS7RAAjtTQ0EWTw6qZA0ea8SrziclJVyCW
7rcIl84gmcf4o3di2C/C8aN5bYZa7/4ya1dw8tOP47p6PMP+BjiGPJ2cpPR8
gAPzZEXvq0/3fgeZczDFAh4/HjujiZV+sC6O35DbHQYtls0A4Y+4qA0PJvKc
bqeZdBtJN6VOpnMkcPFWktMBvxyWMCwAwdKMSGuFnHyy1T0YHyq1PR0x+Ji1
8YHlMFYVl1N5wyYuqgJltLkXuZro+hpydfTJlprG6j/nMtdbUg8kRokPG+fy
Eh+r4HXyS6/X/xmHSGA14JwU6nEPWhVYdhL9leDy35wgBX2ysNj5jOfdYv7t
KXXkf9kWBIKvIR03iguhDv2mxDsBWj4jppXGKZTxlQxAarTUaxr6K6XDWvEa
6fnm1/AlbyP4pwQJxaqkWsrYwMWr8H9H/OTPbkUhiUhB7JlkS1lViFPTLcxq
ViROh68AaPkYD2XzwaO3umw4fOnjIVIqM1SmkYENsgrnbx/xcFajok2J2kjv
hqmaxEWYTlA0v6OVGA3lpoTzDx2+dSyRKLhdIhFUCNc85zZEOvzKxOASG/xt
SR8nBzkjFXqaLZOLPQbREbrtLlmMXb7EHzChDlsF9S7Vx0Qqvx4xgGCKZLCF
YoL1NZEEJUyyexjdE6f/V7qqJDWvtdxbh68Tv1KjkSe/QgDyVOd8JJPIKpXi
ysYmQqnKVyW2kVVkZB2QHKG7BEnHAdNKeXXIsYSmALkMGBb9YWm1Bmrk2wtj
ZXIFisxtNAlTVB2p59elWpLsvKXM4jdlyiDai3p1JtPg9UlD8Vtb0rVigWb7
BfOLF3XlYnHvNIU4AQgUsbta/AONBspCah3Iv81mQt/oegOxdU2Yq6emcC8y
Dm5oJyXs0RSh7xBuSExb8VSb/EvYxArsDVJ6HbuyUeWWHTZRf5ITr52+Rd/4
UIlG+OtEFLgJoLItiDcFlkHfrK0Ze1dckD5vmcNfZPAnndrvY76BTlVkT8vE
BNYy81OefYVAPxnQz19Fl4o6rOoYX2s7uJFTClS8RZbr1X1sDDgSgB1+RkVZ
zj56Er6wT1MhFt5KJj2tj3MOd2gKxS0QSdKBV26drKZlzy4t3k2fLrdz3G/D
3ZYrKUmFore3d2Dojxf9IEVTf1FqBeV52mrbwkcRXI6aw8JgaJs6ezfEb/54
GLcL51Wu9//d8vArWRk8cq5zVT3A0m4jrRCxtW+F4vsUZmuBd9rGhEC2/5p2
VyXsr71f/sQNsZ4lXBGNxA5+rSe6sgpN3/5BriTWmMDyUGv5P0la3lQh6CJL
B8zIV0UOoIoPcDFo9Bre8ZzNxQgsorVo1rQKIDDSYBUhe35YxrGET/677LDV
LcNN2C/UVv92FEh31ZcfewUzk9OJq4f7z0cuHpa9yqs744dx4nNoGLjkPSeS
Ti/6vq6HBVdVXecxLW/vrcn38w82DYSaxGmEhJwIXZNBduqirprWl0s+UN/T
ElGGuNaPQIF3mRh5KBEaqVYusbLWK82N0W7KLoldVdiDLVSUXku+XyL61MR8
YXolSijwQPo1b5fPNsDMcuRcwOXzTYYkUlWv5Fpe6zsQUoy8xyMT4D6eOhjx
DiHDUtBDj+ZTFRXXXS4W6yh9Ji6+FvmFp283X/Ed+5zhNMPItWNje+GB2kMb
qcypRH9/svJS8QFwF6milgfHhK8cw/v5Vaic16RADM0t9Cs7OWft/kAvsN6s
J1YOG2DcAINrjixRLC1PmkhSOQDlqD40sy7WgYU9aI3GRKNgXhwjXh4AlJLb
a7v9er+/glqPuOVSuE/66de68DN8NV5goLFBkm6kCKfjDEFJ808T3nFLzZLO
YeJwPABADxHz+l2ht7zA3RQdBfsYgpBLqdcYr0smdLlPt/3pQCS8lMg2FTex
Aarn2cSq05ntZn9PJM3gJqvHu5HBtkg3+Q1npphlfDUB5747+GQbwokSp0lY
37+sjwz6Fn1AjtlV3FTohGC6db7NEFUHB9QSwMSYA/hp7vmbQeCsf5W/20gw
jD9qDghsmiE4uKAz+CFndwsanfU3mVy9uhdZ0uXBJimTL5+41yX7Ep23fijp
PA/XJf6C+Kfg60pwxTe5YUTcLGARfyZmGsdYqwlveJwRW/1ueoi1Osz869JE
YDtijz+6VhGhA7quBRMxbqsCZoGVmj8CBcvL3zKUc9+8fnnLEOAT1PRcwhwA
IX4C3UlHpT4Q6TAFu4nVy/frH8fymlwnA363fpYle5jaG9MPpi5luJGdaXEg
iFSAk+S6p/x2XxTusUsRxfjmktVTjgftkVQhmfjfZdk0SI6RJ53tX2cc2ASy
/P8qcwMQpja24+dMra2Zh8PPai3z8FmF1h+OyipgxQm2wrXiw/QssUSobqjf
8kvqHUZtUhH2HR6Cn5g0bM7oaOAoihPl2SX3St5Fv7d061eS6wuelfIgPXo+
5lOdDTRB+DIf/WoH5/u7VorIlXHvsvEo4HGnT+yzkW4e9P9QD4ulNoRrvqzH
72AJe5MiSrh9tsYqLItIehMpn4zeRa9f24aRLB9Cg2cI5S7EFdB/RZfr2Pcq
btJ87baYDJd2vy4QvsjnORoLAeJlpI7bqVWfEZsDIowvux5MKb3UYZUGXVy0
VLkXPnCCLYRekDchpEtQCeQro40nWYiP06WgKGnLh8ovFs0N2QXXcoXn3DFo
t4YxRr4HQzzlBEBU9xa4YCZuB1Ff6X5uQcIU/KTX5JBmx68Bri3I4I40pZFc
rc7yNJnxPOLWt4hTgZaJsvZO4efYp8KbVqsOqWnRe8CXTP6eDzj4mKODCU32
Tw6kN0eoMhQfwwJGpK63vyC5p5jzHOe9rZAx8eRT6mHJpaIzKybLqlb+F6SG
RLNFGjO+XdFzlT4jWtO+SEatHyRa9gdyw2G1sDRvno8FlabJJ48sRg5i65Ad
QduC2JRU5+gBnH6XAFVVk4UofhOAs5tOHmOF/sftBMUKe4Ja0TYPI6qg5mKv
Twl7bgW2U1ENsQFgQk6fQ7MYD4zjrVIsf5N272RGrZ9BmZgp+B0hkWJ7pM78
OcM3qfbp/aw+QjPAQ+rvAQToI/q2WjhF4Qp5cSOjNVvYsVBJ6zk9tUG25gWX
Is4qBzojlCriyUKoGdpuLc/hqhDLA6DLDJDVaEUuYWwkCqS5G6iQJfKkJ29C
eIU4+SLd+HvDJ7ZHV860WRtGJJ6ZiQTQHFKIVN/7LN5rf9HIUTUDK7jTCj7I
DmjelGCOqzpdB1tWdAwojtUPiFKjtVJ9jjaG1Hudbt1jaPVW1NPDsX1iWwGE
352yyKFeuIqHYcFe8P42krhWgJhcHOMQkfxg78hWMq+jGic11y1vXiQo+niW
5RwMXTRkEEuOVSwUHQ2LJdgDbUQim0BQP3EwfFng/7OnfYao6tIE4dUCqTSE
jpoIf3JO20wlmFM1xTxd640/569X8SbiWjCril6iqDlaF/001OO2eT1J5F7G
5RSdLR5SVKtx1XivPd48aM5zFx2JngSJBH5FmY20RiQRmwI70qbUMOYAdv2i
e1Hj1KN4MRP3fO4LQD7QA23vRYZI/XtlqPqpHrpjX149hSNTGtHeL5H4bhx6
jinCpsYbCAkmJZdXUPH/lVqqc4+z1xKViT3PUhdELPGIAj1Xt12oS0cV3KEq
NpZjBIIEQ62sNCGyAPPuKQMraTCbnFUmvsWvatyCYOl8Mfq0H7J6vW45EhDd
SpL0Qc0HmoygOO87LaUfFDH5mWK3kKl4FStKe3/qmdPHhJhl4+/U9EBBCaNN
Oo01x+4QTGAQeUGuVLQ/mVJNwnvegA8EGM7qe1KavGYrFXZpGGtIvNM2UprB
2hxF6uBp1zd+BGkojjyLiiWL5NG59PzITGRP8kNtyfmgTjGluIeaNHqDmP+C
ufjk4Mu3COYHPsiv9Uw/SAWl5/9gNG1ShGYbSA0JNVC+Fr9uu3FYl9EsJhBH
WnH8GSIQobwImxdlyGSoGq2HGNmmKbCp1zm47OTvFAJKEyh3H6oGSe2HmA18
xSpoKvmkv7k6JrfZav3f0C6JThwTbJH4MSdbKnaoa1Tpmk9CC+p353LtqX/H
G0qq45ERgbk7z6yGtoLr2Y1Gi7LmT4I4jKdIe5huvfuWPYauyy5MO9s0HAzM
roPTrGDx/+PBAMn3OXLS3v0KWgblcCQCW4fQfMLu6AklB8A2UEWNJroBU2p3
dPt0AF3HJcZlGchObP5+0D2OpyLlP0C+kdIy3Ehw0gPDJf8YE1iIgFIMFrN7
vcYA0irGVT63kbPnQ/63HOUknGohkLAG5BeasGGlBGlkwi8nPaEMzvsmTtli
tZ7mNfqb0ci5AXMWvbkhHsx1fFo4KUxkaafFVS9ZJ+dgWtYeTXAC4fGnw51r
kT4xJpU0uOhvf7Tog2cIJwLFVNhirvX+UKNz2vpMcJxBCEpxKlCko5hTIP47
ExhSOEgSydXEYbaHVQ5xE/reQvcXwSxGxw3fmzmZJa/nO6UDrVF9yF9DZu+q
Kj75tvxsFhE0ogeH4/OV1monVaJlSSa8mz1dYsGta+N+G9/8B8Z3UBp7dgv8
wHKK395ljj2eNZzqJOM7mjgiRXR0bs2FT4a8SOlRCw7OXn5VQs3yhz69Ews5
VVI1w9ErH6Qet8CEcqa4oCu795bSN5vLL5xv3oXzCHDZP3QPTbY7y/J1gMU/
Ld4Dor/Pfl0NZvoqLaRxwG4F1TPxjUY7ivk1fQSanW/DzdmXD963K+MjRdFY
EYEDfLOWfHKkHOF4J3CxVhHzJoB32fRS9+fvtR01u/JlvcOddXqW18d9z35h
hEmQfoh5mqz8o+HlL5ugVORG8RrxmaFf0QKiOxAlRRW5Kvd+VHZxgASi1+/C
oV2kGqq92t+GyitSoFYmcArm7PzCc4WEtBswDUk9zdKjbrWdhRz2A+eat5ll
3L7voKbnj64gjQPerUD94nm3/RkklZnG0hUT8EopXhKel8VbH69tnbjKGrrG
jHX2zp4h448DYbocT938Njlwpsxqn+WTbqwkxY+VcogxQM5XShxWtPIRhl9r
tDT75dtMdXAqLN5f4o2HYn9DhHYOunCSK0sG4CBHRkOTZNm/yfPbtQntVkTK
VDCMEbmpnPDfo1XSWlr6gtOc/P0hfgNJ616sttCJ6CA4/3P8Gto+UJAcqQIS
eQtkfkKTTkQkCx/wDRK1QSQ/ChMoOYXekidytoXxPBBoKm6LWS1UiI62PKim
5YEyp30p52B51U0RobljDyG6nlZGkxIa01wGm/wEWhunb4IwliWAHE0gMxBo
pWhH4XBdAO4UWVsttCiKq0hqIR08OY877z/+j8nmrfwZ1mbsRqYfr9r7+HMD
6rI9id1tCA2Q9jc4Kg2iWMKE/8mns+/CsJuejax5edGSV+nKu7+OeklJApPW
h5F7l/KU/78vR1neIFYAn8hEyzCNx1dUvU2MYeMFoAilYhwsQHve2GIcpsT9
cF0oniaKXlAUAGrwqLAz9JeVJlpVCFOmKFMZkmf8sd9uB7hb8UDghvspb1jU
NH2oJDBPX+/if+x4s2UgZhJJP+IrdfK8ddt9JjF718F/ZoMJ2We52hZdda/i
wFAafKSMkn7yzeKYHAvaeZ8W0bzYm+ELkIPlMLXxTQONFOxyWBZ3xdCr25rW
BnRUEEPpRXX6C4wKpWKo/Z+gCpnf3D4bE2bwe9pIiTevqzmMzrEwoIBA91dE
Z1KgkpLV11EONBo2lpHAzJ6ZqJBKu+mXDaj7C1BTS7mOg44yHnjhgagiFouP
pPqz/IfcqKWwOifUW569W4/nbKSzMAgMZPgQpvzJl5vjNU6GXzCZY9FivZ9E
WDGEFSwOMAy5zwHizHPcYvuCySVlp7ekOcSvSBbaUPOJVBhPCXl4TPVxfKr5
wpaHWFdzLjb3OwS7soQUoOXBy3KbsdbEXuu3lMfSQ+t+sv24bXz2b0RWD6jf
K0RjgTb3hPzJAsL6eoopVVqpi7S110u9siur56j7UHja3+OznncWKmSF87Kb
N+JtiFnP6t752vKn0QsJwZlqyzFCIj0A5O9flRLFLGnHSSmAqIyXyVfa2sdH
4VITvgXTW4KwqFuTFyc97lQZ79EEdBTHQ5/KDqJsRf57JEkWefEY6GrAHrJ9
+C3Ac1/dtOTv70Dx31PxYZF9rwmGFD4qtKi/APn9NdOAdyxU+4QNftHSodAy
xKub8fR3Qt+GtEFMRWsw3+KF8eYbhQy+/GXFLDWVCAQDl3+3NKAMc6xnhQUp
fEWiXTHLzrD/hzUv91fAfNHPVMsKa2RQDjk/8H4aynp4xyQpkbrrqrNNyGOK
Hd3njTkfcnf6tgXDH4y8J4Xo4XN4H28Ak3JyjewxOSeF3MEfEoMkoJb7Bvi5
q9UiOKPjEvit5EAIolgdunrURssGLfiUbs/+Fy3shVy8OIWj3D5kXPQN4Le2
9lORV87Jx4VGw53wr2UTTQYyUBCzBPTDCeVGhp3ZrKZDjZDcjGgXEh9JBHeP
GIUNHCstXqF4uNNI1xlkTWTdKcB4zfYQ/5H9SCBjvEFPGHRx9WZS+zz/H38N
vUYXsMn5qxzi0OtCnfsGeLwD+tlBL3hvYFTEuvHpI40+qDT+0XpJFG+WyQMK
d/AFdU69dSgjgNu2ESqgzzimkSSO2Oe2ISamOAL832/CPksGVLwgSlDns8wc
EkAwMmckav1/pu4uLEjdtYrs96pD0NoZcjnkdRH2FPaCx3ZI5T1DTBXWAndZ
7no9AcZp/q2DkX1ZZ5DcwDGJM/X/bspXbkKixPZ2wqFXNn/3Q0aberfID67d
3MlfGfuAAy3O0uxda61l1aBuWRjhbmMimZ0iPNECjMgVCVfKPVH6VAzYi4Jg
rxm9zyvR+8BA98JmyOMr8HoXOOpBSAM9npyih6zZ6xTXasvuxvWLZ4/6q8Iq
LfAXP0E3sTcOcwG7y59AvPvrCplrdMrZqtihAzKwjphXJ17NigT/pdWIpCv3
QD5ZNglOK/UrUCY9CSx2iN7sh08ZGVW6IwPrL7TITu0eqteYBK67qhTTeJxd
62JKZcs51EshwQI3qdxzikpnVr68cTXyi3jRZhSAsmwwAar2cV2toRyUjEOW
ITN38bZ2JP4G6FN52CUx2uA+r0bt8vJYJsPCdOTQrKtDIbfn39LIVYswNMEo
BUXwX3h44ZHcdy6Cf7wSeLQzZ28yPPiXD0FBOKf1oGQdMWw5+yPdlha/JWpH
ohhvq1E8SEoyco+Tgw21rcfcVgp2pRfGdjJTXd6wQW/efTJng6k9ejJJtTZ8
jpZVY2qcLw4PXuExc0QjeG4uQTpvsY2KdP8TYTGRMFnUrTI4+eM7/DFwdS+K
S2jBqZoWa9l6wTzFtdH3PM7NsW9p1kx1iSUqw4CGUSW1T3uBSDqnam7PeBZw
5Lnb9XCTf6LrA80Y0UxrNByaeicvuPVcm2MJk9oxPOQlCjCgT5n+n6uHjD6B
KcHifHcnIbHE5Vd4yX6AVGlY7p0WlabfBipyd/H3NYKB2ucTiXkTfQsQfGtB
ib3UonBDkX0uVZgp8I7lpWN+RNFurBCwFRdZO6ARRdAKXkYfOApOqMgo5Srx
CpCxNPTN5aj4sX9ALq242FKcIueJhjBs/EQQ4CJU5ELrYYBHys9TcR0hM+Xo
c0hwLJQ8QDuEUgdYmqGlBTMiMBFIb+1+LELwD4WoUxVgEow25sB+IlZsAumU
k5PvytamK8sxN6QkVOziibOAdN0n4uGV7DPU2558IFIMR8WAgY4QbHudJvCC
ZQ5n7OfwkFro1Q7Cv0g5hN9A6xGtqBg5vxmDV2cxkY3EXfj3KmiKOxZv/N1r
KSENzi/egmx0cCBxMmo23N6yhOFLpdoFF5XANxUrJAJKWKjo9un5YylpoNZB
esFbmuVWDp9hWyINi71x8MjQNiJE5o7seUvB9W2h/4J8QU5LeN507h8DCwgM
FNE48r1u+hGaRlErILsMrpZNxJEH3hGsEs6Tr/iB5Mp/DUWILWaKFjeRJqBz
ZMHpFqxtvnfvNyohm2phBWCpsl4rySfOSHRkAEE6Tl3hpVexSmcSfAHyyeuB
1O9+8tVzdwG2sp6jwSq/ViS/kVlRIuo/ua++VBxX9Zy6fmdC+uDLeLNlwXPr
nahKEXJWN3set5n55DdaoZL05FdnpY+PO1S62Koa9o8R680ubGIIqrLQisli
hUV+fPMinjB/cEoDroipVb9jfx+itpgoYHVQ+bN8j2MFEiX+1rx4K8ksEiYQ
0W+RXZvSK4XquSBmUEQE8kR6kJ+dewrzIpHgg9kxiYko3Ks2hxqh9LZ44xQc
nvOWdv+K40z0bSnqylNLXYyijycwnK5GuuD9FaJ0BuDQXUZYXNk6LP8qCpcl
wKR38OUadsNMqN9MUkbK2iJWvhHwx2fruh5cuXWBYBQ0+K5LfTXh54KS2j+D
RSbLM85jE6V2lokFECsU/V5+6JrwqS7eGjVte50UJhxc4rq6PgTno7ITWliX
xN93w2Ape1pKNownHPCw4iqh9F/LP0R2FiP67h8cttv7OICIBRkBuLn4K6/1
bClxjSKnjE6YzXoxDY6MPDUj9cKJtBwhjHKY6El3Ujr+Dcv4Sp8I6CMTmpiy
7ubpBS1R/y/eztqEuMV5mBU8ZKHZ4v8xH3MGSRAqnCaipDLNpVUazml+zYzD
AYltECLPbqzwzAK0f1rkHEZPywcCyOGk20ooJ2HTp7Fn45OUeOHzA+7MC/pO
z/PZepMqJv2myS64m7t2DveTpl7/md+bNHd2jXE6FperZ/FA8Y3k17X2fopU
5pqXQRlZLl2G91AlP4pz6JE3uAdORGW2clJKZRaUM+Ighy8MP0maNyg9iI32
8d49jS9cXkg/BLOC3908Zi55T13SGRNvj9wO5lhP/zt0OfITII3N7/t4iPrG
lYW5d/F2d/wK1+wWk7UXju427cjmVSj36ls95w3AyhFshcRE66mSWrWBcPzL
xI0Fmne8/O5V3yrjRBZIHNAMU0qsJiALuhbBroKqL/+5eWhu6cY5BLWS/Wkt
jDq/LeV7jNLxFuK0/IT5IkckVrhLZe3BDrtuYNAZSjF/4QDh3KJwnz4s8urz
7MM6rgQamTMaKXGdfRvFR6EFGEtmVZ1BTj4GUQmuicPFj/XHovQetECLyTSz
G9i9C5l48cRvKSTTz9iLGJF6SfcXKmcTHT36tw2dsuTXx0P1ngnxqSsAgloA
w3XTiQG5MbCpniWV4z/QfZGJr9xChqi3NLGY1n8OZ7J2sOl6VbLe7+pV3/b4
7DmFQ+rsaYwtsTnWhlS/74zlGArfHP8LbA97IDW0KvDz4hKe9+njKbRW33uU
+lBYIAwTOICdJz42pL2E+aTth6DEwaqAw6Xo50k14Pd1zSwxyNJ5wB20d8I7
a30x8Iw2zXMxAqbqcdDFcoZN76orHzVFHsWAVjZQNMR+oaqAuFITSrhi7keP
r7X+//MPpR5izgBwNENTQikS9a8LmeDN33nQx0l/gKYK3RDDyfZZ1/8nvOBE
I8qWslSh036CuXmX4TNDPLoREwz3UqXCKkfM6x1wKSG1qaddZcC+WYAr1lWC
8jeXfziVPSE/aSFr3OesAIk799EU6fiUoYmb9AlH3iP+/kNrd+S8mOmf7AHs
wEDqwkRq0yjUNxLgxohfF+7UI2nSRuAfULQ27A6/pohmUIIWk3xPEFRaYuK6
DD3mWuZV4/1uN3hSt2gMrE5xf7j8U8wBTrXNhgCywOt2ePti0ilpGB3ZXDB4
4b+GSbwWdsmGEFnuXz3ZXs7PlfJl5S4RxMRTyUUfraSl38oevL/mNi8oK0H7
e2nzcLsuwrtnIM3c8/JL388jrJGeQ/6Oz+JhBEmogcjmggysNnqmhMg+8QCP
ziD2A2jp6KZQ1c5g4IvBA1pP804jDrUBjPadcggfdhOByIETrRPU1BC5WU5e
wTM6RAGg1WchJZ1i42LAs3kzgzVac1OghOR3XhwVdNKw1WyRf8AnLACkxRLk
+WpbyZYjZsRpZkvQDQuBWLaF5+wsf9nqhQ0F1OYtHA7DCHo2ZawOUAvo02yl
cAwGvs3UPxjCKYoBQQ8VL/weIYmQY96grNO89ijq3JGBZZzXyZSONkZUuAPz
S3AHswGKYq8SCBLVGBy27wAnBIJLB4DPmt08YcUBDGKDsM3NrER3+4SLqniE
cAzB1S9zYXR0YgMXQmmdfT84uwOJuYedeem59nk90p0lLFZtOfogzqAgKdzE
dkLsEDV2daQfBlPkBvoeLGHa/q5tVAZgnZKb2meZQupMJ94+fUnkhrfSPVQB
wRDUOsd/uVJYkzRePdcjRQHiZlYwo4qhz93Ll8baTAXY9yW2iwYdjN+Q78H2
6oSiRIgGjdNkcVA+bH3QH5uNVVJMw5UGaBv5P/3/saAG/Me4+WGtNNDIBJoa
vjP5u+/lJVNF96dqjPZwM7Yv7oW+QMVJz43opWt/xxfn1zS+qslJnSCeJh5s
ZOOX8e2xwn+W9rT7ag4OeA+TDMtdG+pC6vHnplXGZSFd5g69zTBCK8HMgndP
eVaP7MplgByni/VM5DQ4IjInNJWa5/uxZ47yc+krbLx5zlDMRFvQoxz326A5
q/7+cQae6+22fxEIbSM0YFk0p6u7irB0wmheJ+oWdvewpz8BU8cc4icRmZBc
vJyJ7mR5I4F7mQ3TrdmhJOIpQ1O5MSNaFNJzESW0TIkUHDh5F3Ij2rmWzDVU
M4JxQXtnnxarHlcYu92D4HvabY3n6qS31GIrSULoPmo/CKWTzf+p1DyWDkEX
NouNnaUiO7TSnlrNk0nAdlCbRP5iD7Vhkcpo3ySxRLHnMGnDpnbzm6ukVtya
ELMPLrwa8WEaWnBUY4TsD2BQxCWTpthyoE1DhXJOJPIwYlZmv3WWRqwSTun8
i4gPaNbxfBvEx7dadtsQG2G7otqVAUd7a/bJYIHJP5m4CVVsXVNuKS5P5cSj
f00D2Ojsrm4VKBk0rIKYBPxaNXQnWPQvOSw8I1p7MNDNCyvmSdZsP6oEu7Bt
/NvB98ke2CnYNhoRzyFGrDQN051yptJPW68XA0F1klmIiOXubC7efeF6EYXB
w1CQ5XIM9ZFDY0rQTghoMfcqKX2V69XsCyAFUKG715MnBz7Dm3WRiDXbg0fB
EBKfypjrU5ILb27krllm+Tn0CzuaTPr4djN5pViR7DPuGCd0bXBwQD9tsKTE
cO1ATIWAVcSk2m0iNQ/yRp6ZKgrPUcPwpGdEzzSXAoMzHoBEvFhl5lXDOGCA
5n58RfVdh1uJH91LJuG1X93R3eeKRMiHdiXX1wLzBR2aEInyaQT8M+5mD4xr
wZb6KxI06VA9v/qkWXvYRrk8bG168yN5fXvxz54aqjp0VEcrsHCmmrpgHvEq
PAdKJaxpoJB0F6dt4HhYtD/C96uBJDYr/5aNNMKc5Xw2Ocu4WY/N5+AhFQrl
rdYXMaA7ao0BgtC92q+LG/RckUlNj7QYmXAFVP5BeeSbEdLJ7sAgScpiN7eb
/3S/4OJwfmR+dKkvqoOZb6Xg7A+vgGiRiTlbc1veYuw/mAqxjJdCip9mE3RY
J8bUa35Uyq6ZfWMYZSRvaxyoevglm3sxexhODCI+46CYnIDC7R6dLYRySCaB
sEmWYiMV1lXcr747cvK6qlXUALlLyi5E83piZrliPIaTm3bE+ZyuTB9/OW/u
CFMpv2CrLqr0v2ITiGDR5hs1y5GLI+jPfmlQ+e0BH2OUI6keeNBz7K9NKJ/v
o/5gYThxz5xin1QC/TUqr5Ao20LruuNbgN9FKc/IhOeeET0KqhS2eXKFELWn
ryCQulMiNaWUcj3plyK5aXQukbEILJBE/WogeQ7XqLDG1dgwAJy/m3S6Rjrm
bPRQ5O0yxwifDOiRrxfJAbDribYXmlbBknFKleY/6bYOFsrvlvF799KhTZ9z
+4DJsTUEbpl9umDpg7n0e83KEr3wtHrqCQqaUTlulM0CBNUxGruLKGrJz/NR
cArygR1cDvnF+muJw0l6SErmZHx52p52Gb4HU1ejDytXSolxNOhsDM7DJ/hl
Qmki55mzRR9Icqni/TO2pH7dCo3htvyjt0kFkgOJ2vgpXZpNrZbxUJgsBF3g
2mTdW9KzncqUv5XMWKFaZyTOE5vyQ4buFoWJWVRMZoMIar+kMqc20XowC/SO
ct6zBPwWUKEUAD5+OX7KVdfmCsXcUj8ZHiD4BRGnECCM5bBQGkPAIvffYUmv
dwEkZW8Ss9igXk25tSI3OICAw702FjPMIgYCRU2fU0l4DSUs7ic5AkaNytCD
Hcy9z+GkvQ1cNjcu/lOvki7+N5bWbEVD+PJWgybea4xikZ55fIXrn6PjfynG
nxGlQOL0LrfuWg7TssgcJd8BnJ9wPH1xd433sGBjU7Sg3/RrqjGqAUk+xD4J
E8DcFW6TvHttbqbvWY0uISAM7j/AP1k6F6f54N6MrOHp+FX8NsAxJMLsfgn7
7ltPw9i7mbSYtTgMbDNsvYsINIjyKMXZsTgS5dZQ3ZrcFrTpnfDoq9UWCjo+
kwo/gIqWEEyrMKwNfSG2e17cKb3crRTpzzkuguKoT7bS3lt9cuQD333Y5k3X
vfraPa8bO4vCwYvmOlelowG2LSEag8V5nBEydl6DysW0euC/qadElyvhLQw3
uHRAY5XjIxdFliAMJ2l36MMByzUHD62aanuQqz3M1jwIXwvkDzCBpkF63+ao
icqfydDROjK40EAvn7JbJ2I3nWpoZUhSE0YZwg5BAuR/7oTlOUYDyKGakcg4
TZ65pVD+MVvg3/GjYzM3vEq30+KvV4T8GniB9XaYcVuz/mCwokhyW7EzXROW
q/6RAWiSvgXhbiucvruxm6zzEE1LiKyGXJIhH2xkfoVTWXydem97o+1BkUSo
8kR40Tmg1JZwHtJeHbtQweh9ifp2pzOHAM9FewJXocHJyMzpvvB0P0qutSSG
QPqvouHTNQn7sKGiHuGkfrrdV9U1L6s9F84xKf5RYXdaDpRgLe4ABCcutYXm
IT9BA0z81Dtw9uztpc3dyxmjZOA/6ppSI0j/3Gz6RNCz2CTAeT4Le6bZUnId
UQywKc1fhJ+7S9W2SyzMLh2/buEK6rXW2EaLfcgybMHvPY04Hsa+t2SUnB0F
pByyQNKE3jgYYj97NVqpdm7mtMPbwgMVSEt4PYYzMwUKfrB4UiWq1cZlQuuJ
MDSWQW7dIbsk746Z/HdcqFtLT6mhQaIdk0567QMQXO+lU1rsBfxym5G4OcJ1
BjwTuWkQTf6jIltIfxFYAMVnjqk45+DvXiRGVh5ywfu6dfoXfVgw7QzxJXKw
W0UcP8eAbeB4uCEqvQVnQ1BGSSLKkOJjM9cXP/gAPVUfMAhEhU9ERv+bNqHy
kppEdPcfJI+PcLR7q5uojU2Xeut5vQrfoL895HQ4wAVxkVyGY3SfthDS+Lur
hiAh3VWr6wUMXWQVeH45/Ff5h0A6l5y20sZZXalM79kcoDcFGBDe0R6Lxfnp
QHQF7hv2LXc4FWaMGbFUs43cigq30ZC52KxgvQjfRpKixP3f6HTycE2jtJOr
omzOVbgrW/lp/UOaKupX+IWvdcDABBWqQCrTFjeaReZas4cHcNt//NDkDBBy
kxOwRjdkoQmzD+NmuPOJPxBYtg0hasboduZK6kXACID5pmUtUso/d9asQfxx
bEzuyax7v0Sd1IbJEczjH4wUpTbvAcXB5Wass5UXFLXkBALXgmnysq7NCFP/
pw5eGS51pSomdq567qmpn92nI1OcBzZY1CR/re95dRN1/8XKQ726cnQ5FzDU
zK9F2HsWn9dMBN01M9r/E0Lqjogi+9fONmlQvUWT/vBxFuC4oQH6l0t9zCJz
UxCDk5hMib6lR02MSoY7UxlSxRXlSt0Uev86OBX73AK5tYQab9e0mVYhjIs3
4dvxrN24+6+QfOjsTrrR7R//mwU1OkL+0TQ4LLqmxwZuy2wsxwc281l12Dt6
P9EAJNVug0eljo1WLfQBLIGUALqpnk3mficWvgudrhGVuQ3tuosRNAbi7aBA
fvN+PuxH6hsHkBLYp3cv5J/G4tn56vaR72Gty/BzRPaRgWZ0VhMxUg9mS7yY
ra4PYVrdu+FNvvqMjiS1Ximp3si9QmU2YSAK67IT5Y/KqO9JPI6qNw+o73bH
XG2c6fyeh/19TUjzRLdSv3vGV4UJ4Vp3eI+2zwvJMtk5BMT/PHTuX6akD3r+
TwRBbWcB91vxlYGqMOIYcCKloyl/szOmzXSr7uFDK0rAadhE1F+9F0ZRAaWw
bdi3Q9PB9bLcOE9YhXluKU//xYBjkfKPqKVmWS6Tfh/UbRA3Txn+IXNY/KS/
wS9LowzaB0ImOqWpF7JEdtv+SjifqULNAzymyE7N9rVEv4jZkmzvA1386xpg
rQFGc7JyRXt8tTyg6M1E8ReESLKyVVNBY9MnIMZ2QYhNDIqH8jB5dSFqPAr3
gHG+RIbPavBZyGuNUik6AWCNDj9a26hG9t5SyRh23H/9gdQ6wLQajEuV92Sp
5ap2qbNe7geeL1TXV5leq1qpzlQHhWBO4qdmISsKH5H5UMUJYPY0o1nlSeky
TITOmDEw6/98OUnBpjQCaSUkQMYgLK98PIGM7/CV8VqxYmYA+k9WPphrwh4o
QKZ9hAm3MXgoU2EB8lga2O6rkuayNAC4sE2PbPDuhC9qVS6V4HAw5DWPfkEf
33VOaVVshIbf/mQMdB9scyKaP5CUbMXvpaIPUQ8Ldbh3p/wcRVyNBc9tSzh7
WkkuPgaE7stvL5z6TFRa2iSTY212XmoatjQgWO7f8h0Z3VUzspTDfZhAaXfG
bOAuQZigsTTH7CjqlR4sTfBWy0biJrYB0Xs0uSHSa5CGAxFwamSgjiIiena0
6Se6bH9nVb5x66cAgpXLspOcntJDPwLu8svzeFTO8gZnerWShDYa2NaOTd9z
XzwBNuf+LjeLh+XgbHD9Vm0pj9gfwK8EslKKcyPWWvLe8DN+oLRlpZ+DC1CE
8nFdL30QY5b/gPfUrwf2/F7giLAHFvwfGTKTjj9OHlz0bHO+Qh3ZjT2ZqRFv
/pfK2PYGeKv3HGxeE31jGYU9HvntkX10bydeMUneiCywWaRqfwj+nNTZ5R+n
pyQhorJbtZk4dcRAnxZR+0vrgWXq8Lo8UA2octVTort+ri8Ip7NpDLXV0Jq/
kpfZ6ziOeFFAv7ZyvvP0cigZazY8+gksUeP7+UM+kQ4Z9bob3cDjYpmYJBFC
rmc8dOlZjisM745TZS4ZGurcp3KbuWfiilYqQqmBC8yImjDFRFBHVf9uhiIg
QovxcOIlWHbm4fna3/nCmKCZG8yEoVemcXh89rEQFHRwbPAuwConJTklbjFK
yxqnZ5cxzz1WO2EmWIW5iFxMsZ0M+r/C3S4wPDvEwf3bVD9qbaOT45XfmQx7
PpPFCTInRYX6707uxbnWVnxjFzAsASQykWC4cptWbcxfA45G7lzK1vCmzbty
o/thMJxg30HLHGYGLJQoOwGR16Ib5JLywBSWGFcQLM+q96f3T2UZRZ/mSEYV
kN3IPPW9ETj3UvZ/lMMiZPhnn3hxhGkOVhMLb85mnQ/O88OSGfkS5q8kJFbU
iRl/rTYRquwLnjUqO9cG+falvEbBXRN7iRQGhVomLrGX2kF3e0mGcLMTsI1m
PK7J2QgG3gK9UJthUV4qfjBi4OrZpnr/4czGmx5PLwF5V5QjUihIkeMeP641
eySSO87VjKNTy4R3zltxNRKMU4hgwwzFrsDs/ler3ro0vy+3p5b98OB6ZU7x
NyWZ7TYoTeUCpPf+0flR8tYyvxWCutJPnAFoTiJC26j4KGVY+HYF+dI7Po91
AAAdPFf4yDVYfaitzK2SpUgFpr5uZwzYUhmgDqSvWJD4eMrbJ947wvXS0DKF
VK4o989uAJXsDl23SFGHZPaLITO5eXMQZMFfDvchix36tjzFThxvSGq9csbC
3AFhNHilaZvYLD2AFBjX0+C8rqyVL39AjIOSJ+a93bNqIxqzf7/4tHv++R+e
OisM8h8DwH7//6b/8cEnZcTaMdh8/KvjeTSPKSpY4kYeCcEgAht4p6q9ObXa
R16NK3NB+BVkH26ljsaFf4xeN/SKM57nZ4qQbp3YBDpORYnzpi9iXsb1voHj
Uqz+hMns06vlx37s//2ONcG6cpctFpm1VCg6tJ9LTzTelZM0W9H+FmsqZadr
hLnajWt57M3Bdnkd4OS6Cs82mhJ8VEzWTgzf0ePovaYlUyfLmihF/M6ZnM+r
6lIK8lksbvKen7/gDgAmislXhJFA7DxkhV2FYqnevGCMBXOJtWpWru0GkR4s
vWA+ryplWsdqYkdSeVKQmedn2JhMDHCg/HpI/PUEs+r2y8FiCZcwL3XetxlI
TBw/J44h5HxAMr6IUd6XHTDyRb0Hj2wbuOgOA6MymbyuRCf4IS4fSlPtz+Oc
U7r26ILMC09NOj3VH+iFuU/H+yBf7IS1paC5Phm76L8Q6snkYAcHhk4BlrI3
0f4QowzSVnjkR2c/Vo2RGDT+2Un0Ue2+xCo/pQCnsQPUSQW2perQaLNBBNjH
mXJNW8EBxqYAiRsYdIRGnLa0QM1F6LSyBM9BJc1hve5aZ7cDcV/CurF1TD85
H2lvTxhoYXvyKOW6u2SMjJFfmupcMigytYxHJkMgCD6eUwddgJ/+ljZeWsHU
9nZ8dI1U/7xE5oUin28rW6Kr9r0fOF3jTvDnKpBA9zUxB1cJBE8+UqVMPKeQ
fPvruJYmh05qO0+OUn8uGKKIz113uMh1j5t3TMXYbpicv50R380o/e/wTr/v
iefK07ArCZ8xYhWQLJJ9E9Ke9oZqjTHT9BIifP1ZOdKC7wew7W15/5NXii9F
jH2oduXA9Ry2xrVxXNefdHgi70/TqvHCUH2prg6hswLvobUQIUFYdVde4+ha
TpOLzSUe0b4avs8PLlxBAcygw5fvOjp7T5doBI6DqqOJlg3a6N9CKS5a3ZfJ
goZmPpg0soiMK6SbWWhdCburUXwYYpww5yZeZ7iuxPNl/z7sq6QM39nK5CCS
sKccfu7RU9TiYj9ZKUZ9hmV0kx49L+kmv09YrsY58Z1MhZKKqpWa4P/Shcqp
eW/264I0IpNowe7c3U8nCqZsyxqaURDBD0Y9eHG8eBxzG+fzbmO65yJh4vY0
aXT756dyczutjHJPIghbVGvj8g1w3E1JaL6lBR3jNwSG2NcfVwb0RlnbodxM
ZpJN8lELPzHL7tSxQMlRCCBcv+cQBlwNNzVbg7FU+IlI31Wc2Xplk6ja2PEr
QR/QTCa57OBOlAj8w8kpMkCdwgAkiAhXe64noVuuf5aCulZ8HwbjwLCiIopW
1UdBSQGhVU9dD3M/oY2cR/Gv8PHhkDq2L9FBOlSrw7Ve770MjvLT319xt9WT
j16jdyaiLr5p+FO+5ZVt9ZktivCPBYE57Sx7uBmNiF1Pg7XNL4MhHGKqx74m
xmow6mMKEA5H2k+JShn2143836OTObnBnBNivMgWMYLm34dbVIoAoccl5nmw
zPmALT6BQ3AJ34pl4I2P9KLjzNY3HcsYkIKRIR1j/azUIlbPYAUjIWUn2uO7
zgCgvYH+nezNc36hHZx9xp0fsfLO8sb5ELKLyA9Djl/QLKZERN8Y86v2nQHM
v+5J1HyAD9XIsUOTCECvtwFdTfTzlVq4S2+0s3ue9Qai+9bDdAXsExbLacoI
ah7M2ObN9V0nK1kTFJJ09XA3yetZUCKgy8KsMcyTNhSJkUn2Q0DdT0EzEi3d
1DbMD4bYuNRYgsBScL7w2i/jK3RCPkSatNNz8SpWpcnOykyt1kE/TVgFOe3L
EkMyCRQuOJI0vUKomxSTvi5rGaDa1AaeH1lQtg1+v992XuJSOENeR9vhSue7
3vaesJAESDV6xrPcqIqf8yKxfszbm1k4e48hWu+B/Ylcaf2sHLngSurjV3i1
JhiFqeKTRh4twgoV0/Og7qSfDaQuSvfC+KZRH9//0edzn+32IeCHYwp/YXAQ
6gh+0L+UgFsEsXA5uGFlJbT+6qesFWMqpJfVgVBI4YHNcSSb8GmCmt78f7uw
Xe+fHa6pqNlNFfMpkKYIvLnqbKnSHk+OS4tMn1HkCZoBW8Ke9HvndailuFW4
l561zUg90F0QnoSGsRAnVpxdC40IptSQ8e37OJGLoibG1oV8kN8X2e3FryKP
GVa5YooyN3bDkg4J1bkIcFJWfAV/tLL4P6gBKhUJBAjySCxpDRYZigfxcsHF
/1W9mk50Px/SihJNfCWJ1ImfmaZH72wU1lscrQXp4CxiXQ1k3MJdGtMisyna
ODQ5+q7RuzKmWqJoVxEUqE57hNy3JmxWEEXhiwdJdTRx2hZo/fZMtov6HrGs
pK+DfgwD34S4bPRgb6DCbiPkGwFQ3xBxkz4ozMMG5ylpY2UhxWrdAG1eFNnu
QEg+9cFSVzl7aMVz4umf2DH+OpyyVJYrVHTm3y+UUr3vrf6HXe0RksF/U3CD
lOgaKHOldTQXiwK6A8zXozMQq3H0E/tVYpmxuQil+dhFQP5XDHqQ6bGFRZWA
tadrLxsYqhoMxZK03jRUDrGyFq1j+YLMemss9CYom6KIhPj5rvpsQt4y6E8y
/hTWhQy7FhhydGcJ9nyt2RAyRdbq4OSb109LBz4U2LVIJeN51Nl4cpsWnwaF
j4Ya2ZFkTFq8UmWsBV4vit9pg47TZ/VAeMa79MCJivJwqGM0IpkmJKQZLVC8
2Rf0ysYbyR88ah6/rMue/DFXxZHuio1TFNF5L7xdOuun/2OS8hgHkpLZaqOA
J8aOpLiGkVkywaX85V7da/1ciO0QOgalLuVaBrvDWolsDshh4IDcFyNjB8yj
0gpOUVtmkkcR9tYqlWp78OxEzlgpK0lhU52vc53UyqrFgilqN1Rwqg37dEzj
SvHJOCHpNrb0ZYCDHcT9oOgV3qgpfQaTCab2m3v1BiY1uHSU3kcyo9Nnf33f
dtdH66E5jbCuTfufwPlE4i41WBPyWAuoL88C8g5DdV//rjqZduMh/3u+0vbC
odHYFP0b0KqhrA73xVFKpOPikgG3eaenoA7v0ee5Kvcn8148IxeeZw6+IGkp
BOp3dNmbJWUF7d3/CkhDlTHgtVyuW13D640Wkt0Mxumq0k4P8T9ulYUs5Uoa
8bS7KtfO6L/GDlMIrq2mGAycVk63az0ZENF8W1FsTEIQm8462yKnt1QUtAEe
xWSd809/aQ0NUQxyRqYtfJ7FMk8nfaglbk8yzXMfcy1rftgVcN0uKNq4uAnZ
IqiQIBaPTrAJ0czRXuPvDj/QfTqnAlAQYFeySvqFhj0+m6SOB/ez4bZq52Kz
kAyFuXKhOTzONXM1bzt5csZBrB25J3cS92hL0bvKPG0bGQRyGCFkaM04TJzj
83RB1CWrW4VWHOQS+scysvv0fHkeJmHyPIhW1PKBweQTguryLeyKSXOkM2eC
7hNfY/g0IT+zTxSmK6pDXPKilB5tV9QseOBA5LLaadBao5735/1a89oUluXo
ZlatbbYbBXOpwMxFdBVtiWDTxIO4t954uxK11tHuWJCL223eTfengjz9lsUs
zngK2zz1rlIxpEuXLDmuJZzvXbH7oKSeSYRFUGdPQq3Ibr3+1TltIvoffV3X
4cNa7UEcZNE/r+6yCqnJoounUQ1qxqBqCm1oUxRiNF+8hyPKctK8e5PS7fBn
urOCk7R6BSQXwl2i/2rfSR1//8tAPwr6yPWdV711YGy3Rc2WFWj2sntW/gV5
CBE7ZfSU8ltrGhmPm/NM1qvSQdnzVcVFVNTJneg0nbkOiiA1QbUTx+S7qklj
39nCoiJfOE9hep79KhkGe4Z/afsknp0CAFwy2nmzdcxkG5ajnI3aJH1xHKiR
N1EwiaVhncbauGEtoHa+kQxKlIA4aTd97DvzED3vzXD0qvvpkBxGGrcdcm9k
8cBHzkfCrAmG8Hv34vFCqD1L8ZC/EORndvSINKPl5l6sTIJQey99hN3xe2vp
osvnPD+7IJs2flsgRWGYipzZf5Eq6GFdhGX76kXf3+lUICP3Q2MjS9wxtqgf
71WUH4KUVP4GbKc7IUcZvx9xk6BE1EpV7gtb5dzPX9QGujdi0iOz/YCZERAD
NrJPCgIDmEepMXQL442lSOlNeUABuCmUOREQ62BUqhjNxQ1pSJezf+MxKfNG
G2rwGH+NZzjyjF4r5Ow80jwJKQwV6Fcz/Z1EbJazgM6YrwfFyDqbX7kzA9D2
W6NoGX9UfgP4zNEGZmzlD8GX64KcKmV+A5rSym6/PRYG9LQc4JJsQmT8WqSF
RwZkrWjkay9fit3pDw1dPvd+OVFT6HZsVyCeMDrj9aXlz5xoPGZBv+hvYSUj
U1bxwmgXQgNtRflDPEVguIDtkj7+Fe2I/fNp4eiyskKc1Zi6xCjN2+IR1YAK
rYN6KnhWM7zlE1vjmoiS6PRhYYEZOAWQs3zv1uuXsbuoJeAN5s8vZbto2SIN
McEOPNhOagzRpetNIfxjG2OvORVnAy0duoHobOTQvaHxUUBKLYlzHCqqNrHJ
PH1GaxB6QeRWXQeqVi/QC35kQblH03jb4r4MntAfLdLKnh4VciMHlQw8hIOL
wdjDKiqKlmWXgBGpLFHXqIDb/q8shf5yLVqULd1FJpiK77A4p8jFGSHp/8CD
6Oeph1Cx7KFRkj5vpFkPdAxyYaWugyVmhF7w+9D5Y5gJR5ZU3gElBGeJ8lQJ
Rm1EGC1iI5DNwyCp3tT/3pcKZ5f0NsWzN7NLgkzYk9guu+N3Mwk5B+Oo8E1+
D3e73rnHDiy/Zb4LQRsHU/PRTCGbCQZDwnTdxcmNUj50O9VHdIPkvC6oQsVU
H7dQvhpEoYob5OkF997jfgyu0My90FHW1FB75mK146pDDoZMxu/40rzes8NO
lGcjkoAo/Hds5XsAEC0i4l0iUHkAQLvlP3MTtSaTSrFIijw9VgRluFqoBUTn
5zmkidMSExP+3G2KQt4VAOrCw4yB2tPABjb1t51RZLiL0K1ujtpVRp+XdJws
SvkQvr1b6m55TTDf4Ygf9xXjrb1+GDjwmb5lGjEOUlWCD5JWk/Hf91SdRTyi
NWPMdE/ugne2oYz6cePsaKAH3G2/Szl0rFK7qEHVH+cI4fAymhs/DNI+bxS2
JubDHz58p9Z4J2MsLLXt4SVNjod9xZlCLeIjJ+OmWeGJi1JizcRrU40/i74K
FnBI/F852iZT5JQxd8Wu0S4AODRWF/vZSnSiKJ4Q0UR8WSzi821lNzdQvkg6
dJn5xG6TzGPw9P2s+/xLcaDcKxrUzeKsbmURm1ZfJzxSEz4jSty+LaWryrYW
MG34dOd09bFb2/81NgGarm9t0cEaxr/wUxM1XMt2N9p8Ud+J8biE/qwUMQnm
LvhHC8piq4Av8sGZsgR3+op2W32DW5K7NWGtisw6GQhJ8mHdcKGrEJkDnFDM
dYXGX2hJcVkX6iMrDohbI1CJH+P8Tu0h5r05pIQ8lPD0EvgRhNe6Jk8Xt3Q+
DBs+oKnG61GMFYiiu1/R2FN0+hYxSLo7sSiYmhfhJBEfOEbfh2Z1t3CAGrJF
93GwhXMzanEgIwGuwj0TZ8ludZ16ISdGWv9+efdGxAhEeFyrGaCjB3iswp+w
ciQNuuvEVMo+wcl3zKYozjnBn3oftI9RFWwrJzCYSgDzFtAwdoeaHc7sLJ03
MRYzGp1uC1V3j6qwKLLoJCH0yM0WrJLKuYuf3U9HiixbaJoaVTAFAlDUiTUs
9njfG+KYHVC4Qbo3bGGFEBWTU5KQAa4HRq118t8Z/Rj/quwp1tZMTv39yqgH
NAI8XkKuso4MQGLyE3CDu3N2Ogm+BG76sSEGQvabDOZ9cBp3Ybyf0Ze902kM
Cl2L782vTDGv5NzWb9A1RYilkDat2tNpFgsecE9Etepkjs9926RA6JkMb7ns
9fIrg2sD9AFicnxIzuBPnF37tDOt9EHjq8GGc4opbHGeGKcvFpCfYFw0ITj7
Cu3ZJESKeLyKCirAp931Abeoq2Wc9uBZEApYFu2t4uoBXOgVPuQ7c5XZQ0L7
p1YpHPOE2MIfajhb3cBsypNWn9lLcs+twtylCFMo3jq75DVbljeQ3K2lazC8
KczaTPFYz8eXfs4w2Xc0VRkApJwjcT2uEKtvGl5jIYFVNBfX8zhuPTYWMhHI
Uhgwy957YPkUGU2/N+bFb+jmpXCCy5SyvjCu3WiMVuaCwWeS7N9RFZK+fueE
MID/WHtto5Sir4OchYAq9e0p02nVvqoKpYs/Z3MGUo/0KOJkyBb+z31Xz8mO
SpThAuE+axi078j5cPW90duehrhp0Zxjc4SIKVfbhvhZsDbBiBWxCuSurjtd
GfisqomncDGC3XtWTbFl5vR8eGkGYR15svH6iBvnedfNpDuNJ5pFF7oFQNu4
PSsJrK+2BMEQG66qRUXOCIAVEPnSgbBpWyYcKgDj7XF1EzrA2FycyidwxGjH
wOysFPPYBD6hORw1mZgzDePh8zHzjMuK3kdGmA9//LrTn0+FfTikQeCS+TEm
ak2NVAXy5hAn53pnqyRlbhggHxnJNUPWi08Rwqg7IWkpEgUasdtYFVgxLANd
DTiEbvKL8seqpLDGhPrF5zYIYILtdueA31n7GLh13Xn28TLBTbQHpPbGvOTC
XwkDr9pJHInW0xa5CMSUTjpQwP5NHX4ERJ6RPTlWPwMW90G65Ky7ZW637eo9
M768SHQnUAP1aSQgKC0WbQKgIiRmidksI8lITNuo7kdvBf/mXKNzcvTPG25/
CpYDiPfqqatyYwN7ZABw2MCLPAXgA55SsdEpnn5QEtSk3FyrQwmUUGEtSuXO
eQ7YWtrPnUyzJ7jzBa+qZYfGl+vsT2mr9ehrKrG9LvhH1LffNcXRcXF+dHb/
SAWsU6tijh1T1XdlHCV5HAjIDRw0Jpext3iAcpnV4j5Q+7f2N80ls3wXZvgb
xX6dvNciwyEf9HTgpUpjAHeotNOk4M+8pOk9dLhfjs+LmuRagUExbX5/nTdl
w0HmTLux/wjP4OJbVAaytS18qjx5d0RBckmJY3rQra6rFg55PrzlM8VlIi5Z
Ui+uxk5IZMlm8gO4+sJ+vZWslXq0iDnTe6cyq5f+9mUrRnZsLYJf95Dzf/rq
7Rr5mt6mCobzI52m9E2gTqarN2QIPQONB888rByHQAODnEeYUNGJc73pA+2j
9ay0H2X0/AdzfRzyKjBAIsixmC3M60H4AozZYxI5NyTDcl8pCiud3GueIXzO
KhdaJPv3qhTy4e3B87hQ0l1C80PF+Se5LCNl8buUeogtdYyitPGUU2DWPuyq
/pV3Di0u1YCIvQSJUW7CsR8AZXPK50CLtN0vjgznPn9DeVlpt6Rf+uO+zL4W
GpFsAodnTn+rhUilv53+2S4QZ7vurmSHX3mYfJRUiVFAPh3w48j0pZlZvNga
8stCfvu9wJ4gQXmfnJ7RE0yCPkLYqdSKTro5vZevnJ3yJD6OkClsIdNAyJQt
OW6PQbBGgQOc3/N16tvitvRH38yQK2HTH+wc+mN3m9j2/9CTdx9aKITvRZDh
m9YmIckxdyee0omELoniHDaVKN99xdn8rtleXHF+VW73HUDCs7RMrbgKBG6+
nh3y6Gw5QNOI6znL4mCyXvwD4JK4wB6LJHUywyLJPgMKIYGn+PpHb5zc0pLD
fkRqQZtZgvyY7vF9YA9yrqFJhvxgjywtqY2ro1gjz+pLmF7CEbirT9BkD2S+
fP1MNka94fwSAGxNABj86cqLQg83Tp+FT9T93GEp2vmU797wdfNqQy9/ana8
KxspxGw9AybNPcAl4lsqpCn5TWtzlxFrCOuEzOxan7s7H21Vgq1ciH4DDMqh
gcEZ8ZuQ9MRxs8a9XgEKZ6BxPxiFGea0JetkKucQlh1Pf8ILz7L6fEEnaV78
X4z6dEw7nixF8jpmREyo9bzFx833F68xg2CtDm3RluiENiYQtBQBrO78KZ/h
0ExZVc6/iPxFZi9hP89lIRPOs/5TjW/0xdsjRVne7ZTd2BtoOrwO/akALJ98
Qq7oZ4wfvXnSm/qsjiHUc2OoudxNC4s7EW5Q8R+YDyYY9mGZZOZwSUhrGZIu
55B+/rkIHUtYOJsntr5iq9wmcNgPLkdFPBi38bozBPipr+JYOOc4lEagcZiB
VLMvWH5pLmTWe9wk43hN5oe4eyw8/vLLRrIg9n2wvja/Q0AM4B7SdAeAYpIq
v7zjuGGQah5E6ZQZtQAzl1gUGZnyzTvGP+26+mLtxxrHEzqhIPmAXsfLpezG
f/3tWWbuCIN/bnLw/haJKf8zCn723ch2W9MeAhsGkqobSzOxooSqUsJ/gOze
D+kIsONiixMddA2LgfvWaQZPO1YlLPlFgIdkvFNThF3aXdh287eFNC9UCRBP
y/MAcqa/yxikVBokqtMbkeoTPVCP4nDQz7OuF5WCbgJaWpU62d8l/WixuurE
jvDDd0LgNjoXtMK7PgJG88Vau4NnwcZInRMDPmDbV2z4o/yTCcYy+eGdpW2x
fIY1SVcUhxY22SV1xEy/15xfgcy7h+wxh5HkKhUIFKZOTSKrWKxy9Q0lQzsz
wiQ+f4MQQH38EbuofeIw7dPDy9//CPsJYwdsB8iVWLkelcmhVNw3Qyjydmay
1y5MTWxck2oa4cMuS/NPxgguqdR3R7H5tUjkXuZbvN3K0IuvTPcwgXFrCGf4
CorXKtnQKJkL7KFOsViHuUSUiKNAQpW8MEdAhFISA/Fjpoo9YoV+ODQwNlNY
a0nRjTgxzOKWcIdQgZaifkRtqH+M4vaUjZ4uV46AFyWO1ako2aEAKLlTnsK/
y4g4tmZczYI/HT74SU0LhNhNUJzRcqenNJOakDRcWfYfCxuMym7gYJ59gVB9
4fN3iygM6CZtZBZuxbTFR2NvPs0qnQyA44WZ7LrGrB7ZPcHB6psNjSXFCOUv
j0mx/ZnBci9lAIQhab704L6O29bXt/JE7vr+NS7N9iegLmDbExGIgUPewIHO
S34vd4EpWy2++tnlFnTj7bl8eINNMazTj2BmjuU7GwqtgYuJTJ0xHx+lMqrn
iguJKGuTUvyvlGF62DqWWqd55xWdt5++evnu1Y8v1kGcLWbNoqrxZoPXkh87
3zjXTt/RaBE3KAFtVwCuEpJGXJpZgdsF89gWUO2KD1cRJfWbfJ1FZvhOgafT
Zx1Jb5K/gcvKXpHdR9lDEwTyC8kcCljsTJVokqYQ3EVg4Ue/e1978qsoovh1
ap8JQEfJK6OAJz0cDSH9HfycOU55cnGXZ0GvuwQHGRfsips5IrBuCssma3+v
HfewY4wHGEm2TEo3c8d6dF5PBnXkZdsvp00uM2jFW/Go+xv+qC9VzElym7QJ
nLISqTVaUyEUtZHtmmvCtOFE4eLDQY7mVMfo0QykSTbu1GmzebuCtXA/4Ba+
nLVCovh+BpMN23j5+c0aih2MsKYfGhY3tu8Bd7mPjZW7ioLBQCwQXWw7Ik5+
jNhjYG/ZZxlSF4BqVbBZyddYvGqMrMqozcdoqOqiATU4WfcMFV1ZRnQTF3a5
xGJKe6mBVgaJkz+kMrejlY532+sT/BrNYl4cHDhDUUv8qzoeNK91IYitAKXt
XmMIkMD9uKSCiM1oUPjzcyZEBUknqjzzDXJ2AGsw2uIHwIJdQ55g3kh10WTN
aaDxY7OQn8SozO7gOBb0VVfFBk1hkHGeIeMtqiIbM+1Pm2ehmOWiRS6CpJin
NX/BRjKiPcJrt5f4/SWHPpsCbMu0maui7R/HekzAFfY5Y+EtGrpWBatvyIHT
cRVBcd7AmVCKZkR0gSkNhjtw9MAwF6TAFdplrqi15htRicKCcuuUgekQUcGE
urJ5YxYy3tS2JrcMHMOA81Y+0xfdL1iPjIx4fgi7VUs9qHrguUEnJ0OJ1Fls
pwXx9DYF71ibwFFR7lES6U3GjjwVzWpf9rFe88m0iIJvCoQXBn0c8N7u5Tja
gt2F1C6wTmHknqClNXCUtDpyhtmda6FB3ezotxhbCZSqAr0oFc5zn1Wtz6gY
9HYMgVIyx0XsNhSfCeDLcVt5fkTWFoaxh1yQeL4GSseX6k2UCUFPYbhHwlZI
PMDC633uUomafkru/gx9jQhDJm01BHbnNJZSTSP62gdZ2WGb45K200wRCIYQ
UlkCvyv7Nnht6FRfgutkHqyWGTSArqJNfgEeRXBasXvLo6TrgYLW7wyaTRn3
RUprL+aRH5xkH1ds8RNex9Tvlj9RhOKqpAwqhmStyS0UcECU1hUWpoc9Jo7L
NnBTO2S7qZpAD/rCLJgv/EgHxhstMCDxDPl6SCCEcB6GRYgyasElOGc4R6a5
XIn+Em6AE1fmm4LsF8k1UGrudyCzu9DFjG5SmSNxNLVh86zdzUuogn7kxTKE
arl2m1u+BzZdU5bqETj58BAh4fsqk+94VcVnQCrnigRZCLfTcJpqfZcUuw43
L8xtJSkGP9GU3mA8h6ZlQRO8QgJV9JntQtOs3FoRt/mvvTxj7JhrUjgbwTjN
ljz+HYUmq7zr147QFZgzLLAELEBY7aWVEeVvQXSXuA/R1klHzoKr75FrAF7E
rbi/yTS5iU59xsBHL3F0U3Rh7jKrWV4g9R9fTjdkYJqZKyW+vC/R0gXjpzA0
sSpvIeqjhx5KW0B0lv6wwkNmKPYopH54+W5ZEwJCWddmQPewXPHPPbC/7UOk
3K3G2s0R9aPHHF4TnCSgJbJU8DlXhCGYcPd2fEL8mooXaSPx8lp5VREwSVAn
p/yZYU2jCuvD+85NsYmyQ6eihyyX0EA++Ry2Tp52t3PfwMDiirdZmGTSvhJL
91rCOFmTxo2aXK2wokRkuC4YDR94LvvqJHkr0PAQnOB1mNxv+RaPwzmFWJ2v
acJj4BIidwLb9BmulFHt1HcYz6qm2oGFkPFHBIhpnR8GMxYd0ZhQXmMtkWWi
KK/cpVHg/uGdej25iaLFbTG69Ut2YHF6wJPFvHSE439MO9lyJvetgtaEXLfa
3WMGjvMSZopqs8VsY4HGEGKTG0d8p4v+OVC97HcORp349EUF09S4gGEW7obV
B21t5SOCMuUU7Q7LFBKQpocMVG2H7Po2mtQ5Gn+9Bq41CGOckQZ2ksVQEfx6
MSZkMq5m1rDZc4Ny+TdHGkg4bgroHMXmSDmDzBp16JnYB3sBdcCJ4nA74I/k
5m7sZOlKvIEsGT9NREydA4d0qg8mFKiOtKUyFk8zNpYKc0zv9u3lNga9mqbb
2r9bwFEp5vaqWmInVkAUPdTCi4StaFQJlfwm9DLeQfjoctu0mL2nbvEKfnUE
w0buWBpPxUtTGlW8KxCfbt6BFKKZzr4sjkPeEOgcZwDyKovrBv5pNzn0m6qv
poOHYBGwq2PeS2sz941sKS/61QeVvZJpvrkOhMACEje37n5tjjHRWx8OMK6d
Y9J+DDEIGYw7lJfgFMoORU/si1UxCN6ZMJvmQuKACOT1XJiakaEPLabudIg2
2AKYR4UAizq0ehamr0aKWqePUTBdz0qkw3AsIvRgv+WcC/bGwm3BKY8M7u3/
wWRo+h6JqHxx6liCgjVj0l/8wHZhbTiuX0iuhhsRwQE52x/uZoYb3zDO9AOu
sz7woxsHcv5ti3RXvyTKHxI2347qhqVMtolL30RgTb+smzvsc2XwK67IZbEz
QqaRewnN8l5opjaiPHZWnatlrlNmRsDcpeohR3CDgYqHZm/rPeFiQn/So3i0
1xTGgE8ShLJbSPSALoDCw5L0KgMy4wHrGKtpTLAiw1d4SM/SVxX7VOiGDXyy
BAREXImxNVD0kv5Yd3oKYqlXjD0DCU8shq2UMdA9+P+UkKShXKoXZsq5KCUB
r2HE14gozVY2MSOYMzcrYMmj4bzlcuBD2xHy5zNC2DorBlD9SnDiq7xz36I9
rRMCgwYm2F9JAAtrG7SiPn4kGjNn0Qk2+yIJuyLJjApuDsV74vrufYV+9May
Dd0b4tEx530AwOZnmhJ4h4hu+EdBPPhEqVykHCTVev3eK9FT+lcVt9vofjdU
yoRrGkK6BiDbjBBPKPE+8PWz3Mz/YnyYIfPo4OJOcxxGcMSslcJIEK1RBTtV
/NTP5jzriIYZki1U6wGHdm6yCWRSVWjmdg/mf5CT51jQONkzjIgHXHd69KN8
oQADAltKE6X8mRgm++iVrdEEPjUyAfR1zY+UkYwCQ4qiyxdHrizUpH5rO+Ed
lU4iaRi6KSjnXQ4ZpiyXnh8SjrdwgEIwPQewYKWJHThuDlazl5Eo7/sNv6kJ
Z1vb3fNbxKssK8pFCMcOyZxwu0vPnQNAYAxE6Iw6wV0yGindiO837FZ9Uyz7
eziKlHLFCIayJfFGb960SoRx+Qwyf1TcB+DatvjNWHR082O9m3+8nBlw6UNm
BwhYoD6VD7gv+KxtRauCiyU5RfTYEtanPb3KZvpWDZiwR4sAhxslOO+DW1q9
S9+KPUihfB0SQZM3mLwFxQ0tt3cZhp+UQ+WiY1IkZOoamoPzOGbMhEVEyFdi
gsc4G1Qo3MPPQMWS12y30+GpiYvuV7Fj6EUtBBkK6Vu4YuzDB/UG7sfFDg2L
YDiatxYs+0YBOII3qIoDpFvjV8Nyri6+OZsVArPN6VfuYGcynmxswWbXyLp4
lAF7yihR/xRiezdtGrmksvRKrT0gVDVV1a/sH5nBZumXtvaO+Ce4QV4k9NSC
RCTYGpIizBn3aS/VaUn5w/LNxbotN/HhsP8SMlcXZ9O3zrcFvmgQ0U37uwTU
t0TQgpbBKqv/5OIdjfnYy3TOHW3ggfNoyGCC7XTufihFsdb3yJ+SRrfldxsU
Cvy9fqmbadl1LGyy6D/0aBPi4RAmllmGdh1PMrmVAyAJyExnR2YoT7UlW3i+
oxbzARxu6Z3b5EpfNu7vyGFSkConBintHJTa+Qont0CzLtgWJ+rQCvSqvU5u
7d/7tKeXzLftBRnknP8QuYMBsuHa0u2HrxliAVb1pUF6/ZwJ07IaQ0WmWUEk
+P1smsxjpKKCB84lyvmCgRyBLUjKCn4KBiypokmHq6fg1p68fQ5OFIL2SgAR
YQTO+6n1HJ6o4F+n6pauBjUVXATEbkNgjc3Wwv7aLSefjNaWgXNarq+v9+T+
vFo3CgX3hYumyLN55bF4Sm581iYr4yuaCRI9zuNvagWkjQE/BPcoMXouz6ob
69QD1EuAhB20TcbExAE2BORXD08sT0FCEcGonP51VWccflDKFLr7Ym4u72YH
TKzvMfsrFWjPMC0HlqYfMT7KHycRSiScbhdFt3zytns+oBXXXNawvkcBpE2G
N4AWneCdvpsXWLjgKQ2WfJJrietBngoi27LhmCyU22+mYdsirkAN0qtNXBR6
7Ag+n+KwWAIc3xjGIDp01OHp3pGoQlWO8nfQEb9/j8fSPKOAs/n1jmGhgIVw
B4oWob8GanvQcqdJRrjt98NRzQeHXbB5Q+Yuf0iCnzSdQfooMy5v6k5XMU+K
jGMwU00wKzx5V7FiUk+txmkMqAPIY+mjy1nPccqbPPNwUGQHcROIy+AlgqVo
VvBtWzaKb3oY8ExAAn9qh6wfr3+YH2mxZA8tbJ+HJWNeBwNnQsTr3UtnPqPb
OULdcw3KLfedqukSEqkKHmZEBOauNmzUJ0zeOMxMOWpBWaK0ceUdMSbLs6Vt
AnY9UUcTROOMcUu2ahIWUdD6PbqtCRCLz6lV4jsPU0bffNdV2u5LBc+vgc1y
UUK1R8j47F2cKVRAhtDGJ/gG4aW9FL4pQwhJwg6m1WvEu9eWfCjZunHHKnSZ
X+z9C2TmNww8tL7m3zkkMAwmID0YM5Gww2piWKv4bjP8TGG+2Ly/U2a789Rd
7g+dOJsyfLTLSMN7I/ucJnf6764PSUYh19cE6VGwjIFDtCUOOwJJ1loEPO96
0HefTydmkmZwWVGpMXEzXK36qGgV611Oqyd0ets5eieWPn+JO7N9dvKw/Ayg
5ieeIpORCLfqh9iP9uepb4O4pKvbyKuT8GXjKvy68eQD0Y3mycMYojfkf75f
UkOCcKKNhi0CJyd+KHRi90+sOF4EfJeAomcHwaPoJUIDZYhnl8Xz5pkp7axM
8bzzNJqZQ7EWN16Gsx11aANvTRm4WDuKTaOZZNIRBFDbmGs/819ItN98FEOu
6IrKatBMjaKet5EWzkeldTgPCXPKHceuF/zKeg0HCubkNMWVIkZ0jG9joJB6
tOzE382DiYbqQMwJ4y+Phac9ngfFEZHYttto710uz9lESXKRNN6lkuwPn2vk
PUbM6yXppHmFPRw1vu7ghS8laBeQ28VEEFtIVAyA64nUF/MItbMZNFpgvwFl
gCZfhJlOebS2qMDG+WMGNkzDt88x9LhB84jzeVgruqVUwovI6Zp9VPWM1y00
je0S6SghgEpfdeIukgfFoSBeuyIJHceiyLTYWM457MgPZR9bxeiN5WLnZi15
rKTtbctHpjES8py13NMF0wMJEtvfiwEtVqCm0WZ77WLhtx7dEPm16AFU9ddU
X6hAGlEI24k4QgGrxkMad01wnSD3m+7CPD9n+khFyXgoYJWyobTp/7Yk4iE8
s8cABkbeDpXjcdTF7YAxhidkmJ0UMHY1HcwMXrmhvmHCosoiG8VNeK8mslqZ
JSnvoPuPw/mQfvRI7wckqJpekGTupjZGZdHdTufQ+BX94U3un0NRxsYU1lM1
vpv7gMCarI4dQm6VIi7RrriFF7vl6Zq5XB9tyK/9ZUQs8WmwkqG82hRA5oN+
4UA15XrZgsNIow/6oBMWIi5RNyn6QVDZvwhKOB5uTgJ3j7GsId75oUe3qFd2
TEiFGaYVNAL8hd/oLEqrbmqg3i4GRyOmVjahiecycZ4yUoupriuDnHu1nIn6
witOfkjkv2+CbkoO+moaCHOHSJxShfLCG1YDZlUdBIy+P9yyGIKwIZgIsndT
8zjozD5ebtoKRg6NzzFCBYyOtaGClS7Ot2mNCkbtgeA1RSHPHuF1mljU6U70
uhqEMDszYOn/ZQ/bDpmAuDqEam36Ja5hWcTpyFCHgtWucOH7i2h+VLMxINSw
+cSnNYb7M1oKZigwJuT8q2p3aZFTNF2LtLici53R+oFL1cYu2JsK0OT+ykyW
c4BMxkfkt1sPJ4CR/y6H7S+D9CiOT1Am1Iq5yMJF7fefqZPHX75QHlsCv7jf
1MmoayS36P0rSqTeVD4F1/OhE0WY7YgFUpdSW2/T49d68WJUq/0fYaCch5Mb
O1i/j8I695Oa6DLjZU7XUKCp6/x2J8vEi/yoJgiqStcDF9JHDtDq9rpf8VFB
S8qprusmowoOI3faIHedsBtE2mAGm480boob2zyJo5HHSdQsVqIFjzd/nX9U
cRn7l2B3484kKVF5A4xryrU5AuKnem/sjQJeP0KmLma17adxyItR23KCqoLp
Uazlt2eK5uMowL+AnoeWAGr/9kZEQ3+bhGyWNmlHu43CwaESKBUcd/EnDIox
JWPbg8efVRil2o7JqjKZQ0oq1dUHIbsi+5nATqA4v1FbiqKCpnAlOI14k2ec
jJW7o3OpF4z+ZudXMJrvm/PAfe2TRA039QexDP4xmwCKaEuInGa2k7eHb4eX
G6WpaUo0MVe7s7aDsTpiNesgE0zuTFeL3zCllUnAAwBJmXf33Xg4BfqVCQvm
CjSfMJHtwuTOGxAtZHzpxWLJbOQNF8w000bpnh/pd3u7UdwSsTBCtbrFXTGI
KqIT/ko7AOvRGwWLEnS27DUsNSAnbLHdaB0rAFqGlhrP50kzZf1Ddt6Yjhrs
kW3m2+hbBbdnFOY5UU/uAGdTAYk/pH6l1BUzSYuRWADVwlwZ0K1BAGLHl+rD
bZop7lNd5BBsfK4T5n/FS6VmT9EGZWBItnaToP54RmnphE+A+4FabVeHkfbp
USQERy2aP8oibr56MjDGyvz/tYDN4Hslq6iwMK1KEdtB4Sgc0Ngh/hGh7A5c
wvnhk6v3mQzTE+AurJ9wuWtnDsgfnlPlneW9umaUvKJ1XtYzT1fVIUz1kF2E
9ItiAsVM77ble3y9PfDnyYSCb62Isrxv9y2dGsJzuv0K7C9sno2q6wl9MoRU
9h/IyAVHt31WMGFidxksffTu260ERYTmv2tPTj5TpZ6C2Gzji1ZydRLmZFdK
j4SHbzzgS0Hv4kN6N2WQV2QWDncK3Vlywz9ygdE/G+DiMabRqVzNk94x8GyS
aa/EPtKm8b2mE9vb8cAb+JaaJNVR7T+uRTKKoyqZv1q8quLil/oV9ns5rhj8
D9h5i2X30mbMkkL2xdjYiZeFu2gjfD/kyy+PmQMuKugwfteEX9ctlKKMNL5h
AbEsl//5zL+Sd0hutzocPosHmPPuYf6RdEl0FeMbZZuZx+XO505QWWT9T3Sn
DL+nOs5bc9E4DLt0ACE3c3PYJs9bNIP/9qOQ+Tv/c2EOk0307ONTV6RUMMFG
C3dA+1FgiQ1UJW5U35dNFMaQrmIjaWPTmO1/uAcrrXkcdDJqVnNBZbrwxO01
J8nlbzoHPxaQ1Kbh1Nhtig/HJrQgeP4f7guNIiU8KNqcQETPrMU0olcppjZu
LJm/oq1iFfkPxZd1pq1QU3xLMShgU6iF4qYPSZ3dmxHb9LMAkoWp/WChR3qt
SPedNM1b0sl+pFt63aKGStPspHjkjXRx3giDxouSLPGKPL8dg+Yxg1c59T1/
1ZbNBBvjFvK/nnnAZPRHYb092+5SGiOvG4GAyS8rFR87PAqMtE7WB4NaBSxK
VSBXamQcD4TjdX6oCVgLA8OlX/1qGy9/NfF/CjlzVnCEpMgtgKb5dhXsyYSq
/EjEmlXKo2/kQm5PSqwOmzxNpkkt8iG1wKf4LT8qNmS9ZdnVbz0lxBjSd4LT
TmPdCH9dD4UbAM0KbDgPRx+y+aDeiMwkzhbxid33SV8pEFoEMrBu8lHq2e/q
r91nx+zmth1M9HVEPpynh2ZjakTd5/SJW92SXrzUM7+OPq/lqoYvx3OXqo39
6z7mgy9WtJhlIlg3kUGDd9fNDNzQOYUcl4viAs4lf/jH/hjdJdta52ubCrvc
W6hDLew1nJFH3S2vP255L5VSZfwhBYBIRJRjZJyfzPkcdO9YkrpWkHS+7NBr
pxG7rRKfqqWjPzmhCBcwDaikQ78+zrooipvYfvwGevIgWIcb2UJHud9b3csU
gA6NxP1Ojo0KZdP+JKUBVDrL1g1AY+E30jxJSd7+15eh0h589SppNCXMAN2y
RADHackCfNb/y6li0FFJedslK9H3osY6R5oOE3OhR13Xgk8I7nc2jTkKk/pT
LG4DNRKEw8t/d215lHBUDT4wm72up2k2pPcN9x/FYRkxTguZYROfN7sUlYGe
P2MFdR7k07Xip1f5eu8/YQXqFOuBsPYE77QddwnhxY6uwwfw7x/PTvRmEaQf
TtNifleQUuJj/a3UMcxQkZrYsLzgx8TINenEBiPFTPlYpcv40OfiiP3pJ1Rv
bIivhL48qdE1NsoBFrk6GDtrwx8+qbZ3R3Gjl1hGxaICfhNUscqOsiGFc2Iu
jVQhMeFLpiT2mphXzaPWi/o2wppKwaXHl79AnBnzMxNY3Wr5fQ2QQ56wViR0
vd8orBWPPi7nxlR9a5CfA5PX8pRz5ANNKGIaed9HgSq/ffY+q/+BqfzGYCc/
B8E/4cFoXqrzBky/TrZvIu3v4v6lijdeYd43rvz9V+QBlwPqbBtX76t8w+FC
GyU2tJ+0IAV37rd9qJLZN5ymNGnEzB99LikpvnFR4dEyDBfMKRsKpTojt1N9
EG93Nci6H5gjoRR8QNyLYRzcyNF+UDJTaIjinegENk23Z1vQQm54iycSZBGE
KII+OyEbcBKplTSktxRm5nN+tnfAJfvtRBPOsujX3aKhUds1qV768PcOuu/K
bP+wPHW9RZxytkN3xrurIW0cas0qk6+cHSN3uUiBf3/2tuy37Y986VojmHCD
Cv80lNQxHVsdvrwKiXAeMUlHHf40DAhXbBahZcKyWT48pTzaUkyygFoj89e1
GWXdEyVgHWolvGiahFf5CjkdVY23AiycaUrsJdyTdI87XHzxGtkJuzbPRQUl
eujThZfbFUXoLgYPBDgYYFXXkcKfJD6IMiEacJ75zJglvvg67eScVek17XJ4
KbI1WoWls7yfUQahb4DGggnScIvrz2yFab1yqVBjhdRFIvbL8QWzVyv60PJa
S9LTd19Y7wonLr1emufXBMLd3+2IICYRm+09Bx18Yrx8xm8LUy93O3hYWHch
JXCTVkL4XCi0RfdOIAGiXJHc1Mjf+iq1pfokSfEaxJZlTyykjbn0Ym3+OxT/
6KCfZ0Sq/Yq/akkYGaPRizuS4sPsX2kZxls9Es3pAgoDlEsidCHipfXkdrz5
oi0igIgzWbFfD6KYI2Sf8RBMlQJYl6PQw3PFF05a9RzhnDB9Jv4Y4APCMFIC
tV+wW9jAUw/YKT1h6hyUnOjb3wCiJCu0EJ3X62PQKDpVDTFZt4kKfjnxbls1
Pk7KeuQFhfSuriTJTxQPcXG64gxW6fp1ZFSX4aOmU9ZmgJJ8/V+UB74Z3qLx
5PX+VkmQUAEwB3qBluByDjRDoeat4Bnz7lzTH4bfLenzWueX95lkR9NNjMqF
Wb2Va36QJNsufATDhHbiw8Dzg22ktZkL0v+QXAQPNV6Vq+Am0hc8g56KAmKH
4n25g1/5aZROsORx6u7FEOG16vNNwZqhFU9GQaG8LStfNRvBk5pLp42Uszji
HZv3wqF5f7L1Jfj/E6W+RNNxtYvHUdUiLQklngEo70Z7nmtwYoZgDdEhvpml
r+WKtb7MAoe8NNa47Ko8cghPieG1TfS2bUi990y6XPzioEdsxqTmrG+l+pek
N4tpsV8dHzU3q0xYBcNiBoB7yUo5Yo4U6EsZPLbj+N6OGm5Uxmp6Q3OOFG0c
RreVKOWr7qQ09lf9I2KTQVgZnlf1DWByYydrt8cIziiqMYvKNDUjiuUWFTaE
fD3I6Nz5K/tz2wwtY5wKwyOIaRHRGbRTeL9alvlVe2m3kuOY/x3WXkorIlzA
IfGuBA8UnAr0wUt0KjkFVxqbOXgXoTJYqEI3WjZFl0tULN2crH50VekcbDiV
9UyzM/KT6CFv9UXIlhSvJa+j/VFJXT9Gg33X12JcO8ttcl8OX3MVWtgeTzSR
x80xVaPiozcRrzUM0YtbfoTKKTfWBCvptXj8PD5t6euJ3FTTzEGKPv6kezhj
adqZsNm91e4bio9DZebQNaF7vcyondLMvKAR03CSv52f/y+46avFRROWnx1k
fPZseq37BZhIIYRgHOz758sKHNIdLEMGDnZ8Fa+g1GpFnm6xLpdno7zn0t1r
biDT47vqhVTUWusxD6b40wSw9bv69py8BBOhO7w7Y7wi2/TnZmtYfGb+ZzrY
UDasNneCxZsN+hF+m28NJadjEBAZ/KGhGL36n51Np8FrLgimT4ieubL62UXA
Bq2x+i/scDuEmejvqL4rdZQIjvNCxlYWaXMRhMGjnzMIbjJDjLR40BTiqpQd
5gxwcd15TZS54bXdfYTZGQrRfayPRll2E7+o3VB9Rma+6mlzzaF6rzl0ez7z
WXlcqQFL77GAkV1hlrmFXYTZadmBTH15ZtsDjgOgjyrsj9hy89BcVOkhBOV4
1fpskIIP7J+Rr6Ehe5tYAiBNVpQq+j6ucGhN8n819A3L0PBez7YNrfGF1now
WGFGqgz+NPX7gV8XtDAfpzpKDCdvUQiPoFqqN6UQGFRlCfqv8RxTt6mkX8fn
vUBnBQUm1elyT+GDybH6fc+eXRYBWoicfMeTTNoAMo4D6/fQA+nMTY573hDG
dnUMa6p8xZ8WqLV3mosE32OT4xNRdu1zbBMBZees+AfDVAmXdAH1FKsbEryj
Kuw3Ld7uoL/gPEKquYZV7JntQUhnT86oqIzrpXGxNY8IHx2Zq4W9fH5nEwac
JadktTt78L6yOkaqlJy+Isa1KqdQ0qZZSEj9HVAvILS7pD2r0QpWvLzVInnd
2HoOW3Wnnj/yir2NfhsjP6WyI/oi/r8PelfFWAk6MxZWMNfe4SXDU5qaLRIz
9WseEcaP94QCNshi5fg8+dKZ2so1dUiUvLDEnoiWHEYq7BD8vTo8aCkH+uIU
myPGD+l+qbp2OFb+Nbq9mZG8Bi69FFRYmCgxOC6RSPKePQ3pfhsrH4GG4ryp
cWWe8DA7AZHSm7gAeUzn6MUtVDUBoKLNWB2VSfqStlKlMZsXLIuHIMSQYiHB
eeN1bR4YmdeAuimwUBbj9BS9h3HSIbBFzQQP+ZFVAP6+Op7/n1q98+dcmWAf
E48xJQDUQw1lRcAfT7WExM2/O3CpSOJKM5kYQ4Nrj4E/U5N9deazxfNf6nDZ
RzQzCZFvbwySxz+4LcwNuH9X0miCtMGsFdDhLn5gQmS2Ke5/twc1z/5L6LdT
g5Yu1DOjA835hSRZBXJc1FJV9VKNzbrHTJsh0qj8zSp62qh5rTTmeZj9SRb/
EfMAR2qUA3McEz0Qdfm5FhMidgZ0UnDMKdl2cZmHuDf08dEn6Yj5Iw5SEb6s
q8BCbY0brDACclQTSw9Sx1vPcK/t/6VjkcC/r2ho98n3gM5jrdkLR5yh48kh
DjDYy9gAMvmjLkFqFPRG0GQA+4fak6lL9FmV0/z7EY4K4RgwtQqcEfpu4tjV
PU8KEoV6aY7Rmp7f6QOhR23ffz34Vi06Np9A8sW8i8p8xVhKsgFgHh96GtsS
yHe618l5Gjlti7Asc/9hUsouYsqtBV/MMdw9dLN5oy4VCMpQueTnAuZos3bp
Ktr0ImJOzMnzAzuzAdMHb8OSvumXAx5kHQkTUZXJfveUOXbDDmvcxfrdJ5Wc
VqzAMOvAnNGgnPbLomvhdB+XBP9yYFz0p8Myzqo5M9dd/kUp85D03WBz8Odi
N9utznmony81GMJ7LDHCTbDt5rECSMe7x9xhq5F3T5dW5QgPOSaJg/GaUYHk
kt7eRobXHhDNH1kzeePdthiB6ctHKCsPWbXXbopEmGuwyAOVttAuJ7SYwAT+
S2Yr2F8UcS3uf73wgg3eQZrEVFUsgYqgwLxNlhB6535ckpOK5HZm21l/eORS
mwA26R25Wfx/Y6txePkKN7qaD2ZLgvE1lKW88s1vny/7VwTe9vJLAvkRoQ6Z
lzsYsp9jRVHgifnfsX10sHS4meurN9V7M0FJTqX4rfUrG1c3aGgNd5XSPBo7
syd0mqBScxs2pBifdm9GnXrDOgVMjdHUIMOwQKB5bEsulHd/svsh8m9ikNM8
CYcFoQ5ALBnqsKKSogNrqxL8HdZVdhD8rp0vwJQL7wLzBu+gtynbQc7dmjB9
HwXL0y+2A5XiBOVWUjLRrqFFBkCLTUWLDXQPHAOnIZ1ob7IrTgW+oief6GuL
PKOlUHuqkrpcRu3ewg0Fl2uK16Pm2qeJGNnRZxS9/z67WI0GY/u+a2/lEGFs
QhoBcQSJyvlrNdHWo6LHcZPiAkEtsetc1S/9sM3nSei8bHosx0SkQb0HN/aI
hC4oPjXzjNZKTL7LAucmfAW0SvXLEXj3e9VkqRIJKaueVjgJQKRzJp+Uv6C+
DV2HXkKNcWB3RfhvJeIvkhQrm3oMMCcWvUSTxYQosjP8dYvalvJWFf/cc8EI
f+4g+mVFC2A0T3sbXIzGaDKxX7st1xPOh/vSaszoPGYwI92jOjUNvXYKleV3
ix5JCh29z8GHaHOR/EfxoyIhPlJZbz15Amo+uL/UKlxCXzetlDG/3bRU7kyQ
t/YDl/ozJOESvvwceeOFoQoKrbot84CTSVTMxhqnc7K5R+mmynH1OF49yu5N
PYjKgNv7E7/cgjPvbW3QXJH8pWYV+JA8iIciU1PoGrCIq7cAjnED6ejwDuuR
ty43v9K0jwKAZJ196niL0bY57Cz/Mk7pRhxwSjz0f8JAl73w6jSwA7sy7dec
4GMhVFBOo1uKVQDa8T3Vr6JlhxUUNJQzDxGiUyPr6GNDUnI2DslmlU1vUDKS
+3XM9XzfoUsqhutXPI4MKVu89teZ4zFOAhqffPpd8UyUWMJVZkCaoyVzzaau
FZmHcK11dx6sA+j+mP2Ui7BsJCy5WwIOfE+GFweVxlqipMT4ILgOG5aTJda0
fWDRW+Sx10VAq0jPy20Z55zE/lCiJTNSHs6jTf0531xXYAPgdwMeR1wv+Rtz
9rNJGLuXbbVGPaWFaE2aZde2MWG20DkcF852zeqO9jLELZofTYTG5ZnwlahC
fEZ8rjO16xXvOvTD310tbA1c64EkEHGZ5doJKKHugBVarbu+ONMLnU6evMPK
sKmcZ0Fws2u+c+ntAveVSEfr1yNo9ZxdVD1kZyi3YMBVMJfd0bpg0mc+yBWz
0ZG7YsSvoHY9BfQU8dpysXu09AgBx9uq6Fbr+pOXpVf6yGcI5l118Uq3jLty
lEBbQT3kla86OCWh1db9345RO7SAeoVjfF7navblN1Yko5XxZUs7kPo7EMBC
zjbGXahJrcXwXonw9C+2PqeTIH9xFHBwXCz5bdJBSBXMuzJ6jmDS2ooON3yr
Y4VpeBiMsNYPi9aFn6tJVI8oRP/AtfczR9hOHl4yqkgfFCObvYHYwBMRmIEO
DliPe24jLiGIAsRxLDHGePfL7T+nPuPMB7B1ccQTD13O91r89E5XPRo6xJKH
y0GBKChfVkwrk5/J4SpqROa+JpSujypn9DADxYPYlYJvUNaMA0sQW9p62gyy
93uRuHrUBapLqP0S0SSygiqqfTsoRBc36Jj8ObaFiEGSq/9XLl0jR2t/KY7P
bQRqOdNqyFqjECCGZ7ULbUxBJuVgiHdkw8hjdvKdy/F+a2u5vQ9pdced8TPY
oYoraL3U+FXfjcxQpYwMnIpNcrfyPTSNG51OtjEd26snZC7WxMct0aL3eji9
6IM4O3WDZoyGUrY35hz4VIFLyqnmh2Qut3Dahet4UaNvtEeIlXNz9Q6gwjKq
OSZb1eLHgtwxOQjjfQiqGdvDec2IPtH1S+M4dMZ0U+gdWL2ijzjdqPCSXecm
bFkj8aaqXR+akQY2f8/ZhWTskROjyIB14jB70aQuNUaYTduCIQX33BHCEQFU
PfAIocMJSv7iKbqqPmKcHOA0I2JciI0/zjUDraC7X6atnt9V2Xt079eCiTQw
ekBPSzqkE77m2zPbmrWjN53NEkvI8Vb17S3sHjZTyPfuooy59aVwzcCNecyR
uaxSummVcNPY1+ctzvkTP+m/zSRrF6Jb+VemS+yx7/9RvUikK1JH/nTu98v0
wpakW6afe41sK6gtiypIhkGu521xqzYWFUASIGDAJBQUMKLWfCHpU1yVLg1u
om/k0gtU4edH9fzYpBbfdzgQ0YDWMuBlVeBJihtm03FI0NxW23CsQqWexBBk
+VpiEXMU1bJL1kRfcBBxrM1JGo5sWGremQ90BLaCINXkv8VUz9EkXe9oOPY8
isqX2FOPhdRmbPyKXrphXbhk0JKRxnIpUg2422F6dZtBzJGFx+my3l/xDNQR
Y5dZiTeZ9DDLpYdKIXsuNlZPrtZRPwWbuPIMZaF86MIlrKkD9d+c0xFvsgXV
EwyIikVM/VAxU7yAzwPoEcafx9L74jByE8KUbtBbRRz+NMjeqq5Fv6xhy7J1
6S0TBtjrkpjLCNDQBCMbHAYnOZrXZKRt6iFtWVCjq0l9OLgXA0M4kiuyzzd8
n10UjzEv1yDhaIpgbt5eKfL201M1UjCZZSpH+2i8IQTZtQd2JwjlM8xdKbZ/
v9qK4YucWiVNQW1IKjUuBk7SdUMO4Yxbgc2Ztqh1GO1NXw2mym3QSnAswjFA
HWGqYgH1+6voreoIc+zsXXYWrj9anwcSpw+p4iV0nkQkQsVn2qC6r66Sy0UA
CKqwnlSHf9MpPRkiGFnrBEVFzFaesH/hB+rVGFDgyMkCzf0NR/OZFR3bh/0+
uprblEtiTWsKBRpEgSZLo8MNqLXkCSZhH/1XdE7sI3Rq1WoFp5Fzsl9B4++b
TEdkkZQbDr5SUGxL0CbXmzRHobq/7siYMbgYiuARwAosFt0J6XzfbZHPWSu9
o208R8pLupBDfyLIAlCzJz5BUUpY+77HhHmnxpoM4iCBPyA+ySnbM7BnTosI
6uiODQshA1lB12FuC0sMu6+IfNNwejL9BXlc0owM68BJalgo3+Dx8R1Nyw9f
KITkDBy/9pzn3E8dde0Qvdqf/rvObyDAKlaY1PXS1X1tV0g7RlgqDWC/xEta
8um5norPEsINfBgxR3pAN2EQ0Cc1t8GCjHa8c0xfNYzpcn3JJUI8BVUSWAGt
CH/h3Thx7GgiGZv6LciwsA65jab/SIj5P5BJZKTo1e+T1L6TlZdjEpPed8wW
w2GpwAZmKsBYP+lTlY0NLgH0eopXEGlieekuQc6L29q/2DSNTa/eIt2B+Bhz
bNAoBKEG/zocylvCT79TIjpc5GDNMTY0WaZY52RfQkASyTOVi0ID9GyxBpmy
VQUM43uOJYaTZ/fiuXUH4IrBSlIErPtsuo9+VJLUbEvGWge6hGKbtOu/nTO4
IG92SOa0ZhEfWyljO6cSR+sqOxZO9A51PrGKHfoupxt8m/g7lAzFUFYQE/ES
dutIlY7Tq4tkMNXJfTUWB3lzPWIT0emrphyI7P7wBHcvkfBvJRl+s2xP8i+E
EVezszTEe0eFLGXay5c+Vp+J+wK3GP7mgI869FO2gQCGlO+k7B+8aCeW5D5L
v0UXhlXhunachqX0c9/x9XPOvtVLVodo08CERj4Yq0LtIalJpcoR4FlhG+dt
AV2BbumxLPJhdC3yME+TlWBfcQPpoQfixs1/D8UvDyfn8TN6fdKS8ZRE84hl
QCxj/v6vYVWKwl/FsSuj2PUtaKXkA14/vnJAYLkF3I174acNf2vJW2mGGxJZ
tDLF8y0HccpS2bkOjkdRMhb95T/P1xCJyLb53o2juFQXAa8gGoLMNEvrOM4c
m04QXxdwmnduFlr2M2+m/q+s1r+sIIVqHLmAbwVMZkpi+n9zjkAYwQGSQeaJ
2g7pChzUg1tM6g3OPS3TaIjneNvWbifXsKZNrOy/XlfVqviwqxunuJ8Uy0Ri
LFMITUFRqz4ea5eP2xuFehQhXdlZflfiPNvyS//7D5927lM4tyyun6RgzSAe
fVg5CaCsWiazC7FaJTasgnpY7vs6n9sURSVc9fdGteXvz1wSMB85+hGg0X9K
xfqVRqKBqI7GYtJRZSFNwyHBLrDg87KFXXQC5Brp9OgRyBooZA6ww7Scg8oK
qiVO9pQMrWpM2699EQn1kkm3ncZo90v52ZRw6oMr030IeDZNhvTgG7RSUY5P
YxOu3zw0cXt5Mr5exjczM7gVBNEaU5q9ql1Tx28r+Nj+B6XEt/lcOS/JkuBC
3lilQQcWfqWSO6nFOPzukRo5F3mskm7xl8qMQA8IjPFg+MtnUFjeeVEtLZb+
Xv/JyvdmRLfEwDfaF5ymBYNWG0kfR0Cz6Gs5SxEW+RWHNodj1g9/C1bROmTl
NvyQU5UeVdv4DwclhB0djV49HBleO0X3GUP86UnuzC3XkZDTb/n5yfqyIuux
Cz5E1fzmJsfqZWXEx3SQ7u3tL1mIDo0M+2HHa+r3Ysk7O8Qltopj7OWvMKgp
vc/KfTovaosMHkcZCkXmng31R/1MwxFWFjdgzlYF/DNkVy3Lxwt6zz4f07EI
Sry6lWHSrXHoGVFkoJAxQH+m6fhkLaaCdh0knlSefgasb64/KWgJUp4FXbW3
M1o3sTuqGJkzqXE1YDfdtup54ZNMddDwiOMVw4das8ZaHA5+S6mXPgMt/FCG
USmAx5hSQ9WWm2EMvr39NMwExU6jibOvHpyLbkUOCtLQmnj7xXt7CuhI7u0u
Yyd8inE21QcZ63B0C4R8Dk/PmdOc+AaDcjDIvXrSs3je7muT/MxABzuiFhYy
DM2RlIjw8EbA7m8IcjAMZ2wgGXswo3NhS8dvDmr2GFBeW5lOyaqCRkwWIpkC
tMi5ac1NlTFzwTbrBbN8FH3cdVsw9MtrvD7YRndBgTU/FHrTH2DAmdgH4d03
62+wn8AP1BfJYiBSndEV19G6ZTEKf83C+TNNV1dS0cAMl2APjCvonwF3Q120
fIC6UKWS2HC99x6gIhFf8OpSlVMcPm2IuZ+RKxXOiM/q4fuVYYvMJSC9a4b8
h1yhL14sfN635yRpVF5+mBwIqg1n4sB0nYJH9OpiPOi/bk90/WZ//7rPv00f
0UdR09xMOp/0Gzr8AVGjtMzcMcIpBipzO9kFhLbWVYCq5auHHJ2uaclECx0Z
/OXjEQACr5PvU9BnpOp4i8eH2u8LKUOYOboyLit5arW/MWReWpc2vK38vNUI
nagZYFFOdhcWvzQcl+V5vM5X4TIiBtY9HPOC4g9qWwEbT3RrSPOGUXhKWuJH
sv7y6pKo9HknGZvpYawhWcfUDA3isQU8P2q+VdiEQow2N7aMR8Yw5J8SOvTW
xsORYoVUsjwTNZjwOsTHcmrYbFmjuv8VNxXZ9cWLcA5qHjMdalUPJ7XO8z4y
5psQB7KM6dX4ymVzDf2O6QYPwPIA94hDpVparMhZVu8VPzxBAitOENLfl9Oe
W/dtH6/hf8ikRwxYkja4GLmFDvJ5NChK/EEBbI1m6O/BhFCtNTA7kItF3167
3Sowbzsg7oXd46n7aWQ3eDczRSGvazkhWIm/Yl4jkXuNP6Ey3M9phO6hmrij
Fh9gv2RRJ1Xknzgjjkf+r3P17cGKJkbWwXjl5S0LhgRMqqDJQEYXRtdkvgPs
oFhbb7LuAsnJtsyUH3+gFUklRvEastoYkKE1GPlOVWTBMVghbGQMY/c8XYFe
TXQVFc/ccnf40cxI2Dsoyh3/Ph4wB+0eg3Bji0hbaLYMjqh68M4R+Y9SFuDe
HI9P+RLyN+igFVSD0nr+vZ321ALKlHjL/8Kcqv2h3xuuR6IAjXYotegJKnu9
HceULH91ld9JZGONw8cuOvcm6vhcTAjFGct/0vfeJQ+tkvj08dyYLXvMAA70
D2OZhiSI5V+NbRQhx+/ArsbK80cZOYaQsVuecxwCglORoWG0VL/JnClsseB5
bpgnxzdSLijQkQ1j7xVuBHuL1t0izSYMZTnLQhliv84ZmBA8MSLb8qFQ8H5X
tuKiyPAFxr9D9ME7tCT0y53rhWHlTCeHQkqd8zLr+Fxt8Unykz14x2a/LIfC
Mb7OIEtPL0ZOBucm7eDVeH2nn2QabRUNoaWu3nfQk0BeVmeyVzXxRYyfJe4b
/rE4jhWzCPQ5RzgmNBVVVjj1iQl0kc2WCuYkYUcGsvT+Vaglc+2LexrkNgzd
+I9cRfmgSYQWwcoHA5fFkuFqEekCih9R6fNbyMOn5AX68Igpl3HOhKY5WStK
r0ezuqIOZW9jjuht3grDqiwejjyK2uFTVVjI0/ywMLXfK4RHZm8fQQRkA7K5
Nxpfum1JBZ1am0dYRydMNePeXieCjNjYOw6SjrFeEUmiGuZiG9xUadq6Eory
VziFPTCAvWG/hqhpHe7yuP6UPWrxyRfWDCKcsBif46Tbk2lKaFB4fDe2N3mN
Xayu3aQba7MHAgf/j55gKts9F4GZbfO1QnryXjBkhqlZ7WqcmXCf+RhiM+lC
fCRNgX/ZLuuOxxvglUqOK4VEq0+LRL9GwcO15umsh+LbhvcIPk+ZU6mHRHkQ
58Ox8EmvDGfFSBJVE73WhdYZBQGv84xn1Goi613/PHoPwKi/xtxXhM3et8D2
FhECmSg1XP7uESue//QvdCivrPZ0HkEAwfinxV07Irj3zgEniGU6BJ+qS23K
DE1tpLUZxXMhVp/TVAk/gyb2kM+UOywLPJb1Hbo0Q9tJkJt40pJbkWuitJsG
wsDh8jR8Baf/9ozMyvpbOOhLs9Nq/I4I0jYRoZeR1FWDcPve16o/EWQ+d6m5
sQ85HWVatqM+peEbn8xgPx2S3q0YvLX3KjbKYoU9iePqDMuKSGmxea4+99C2
xEZb1twJsZmmhiZWjjmfX1C1HKqZsZLdUqMHqbO0jF+549fmHLY6/8O4MZDq
7SVzTcTk9XrPULcUr8C2R3vq0ZUcJ7V9CtxP/FpL6OQIeVNjIdku9jSOZHMh
Cu2hTrSIURf4vleCmEJmL63UicGsHuM7kO/CkPqgFFFAwoFNtyTIQ+FennA4
TPxViI8FJdCf2bFmTsKw38PnXWA4N1+XdX1Wbs0nqlPM3Zliv2MbOCuAAINH
3pmGcohmAxsag3qMQlIvT685kvNOcQku+08io5wq3xuqDkXNwDcnSrNcpWSA
Ma8lN/rqBj2P6GGYRCbw9uGwE2HzmG6p2dgY/oQAokh3rZhb3epdGUOWS2z8
FxIwt3qqtp8QqUY/ykVvS5GFq/3Vz9A6bdjLDRLAzmo4CvtLw6wPGYgWeZCy
sHo5b1od5eUsnHK+trxsC/SLYHzR3PYMP+9V5ddffwpwyeI2B6O6CNrKo+CJ
wZKjqvXZoTJtYfcA6bx3hj5w6wfC6xgT6IimWpPelWHRb7laSX5ty4tgPNc/
N0wUtR0ZNINQHJG8oYLkErSFxUvGyp5zcBu1F87Hv3pbDBhzPY9NZEv3TfDL
PCqAXA/FEO0mVBV9VbBe568SmdFb0LixRgGCIFa3/fJxLSAXGs2xll7VPnDF
ZOXN3EecrsJpRWnMb9dPG1HMNNZPdboIDM4CtTcSFlvbJ2WO9AA1De9voizU
W7uDW96K0vV943rNhyBZV8kRqVDPeHIF5hEf34U8cvzXqiqPuTojxVLVwWAC
VDKR8Ook93FMutksJoaakhXVJdI45Dsucq1sw2tVQzRCq5NZC1YWfU/d3cuw
+l7rbreYbtL5LbUQcPZSFzt8BV21niNWYOXZzXkJUKgp6z+7z6a4RzO9kM9K
yDis4qJNQH83felVYFeFC2gEeT/pIev12U+QCLTwlDpGSVrrDI7cD29V3YlB
gsEkYWJ7MAJfEHe2dRSJ8PbgIPRtBG8g8QjTslAAC7YHSxJ9PEqKdKweod6K
jWa1C+7h/I8J8bY/bWkxJR0gfCkf15vUOO4cKAqbeVaGczLeRDiAkrp/R4eF
0MfkjExX3sjsCvtlEV3z/HUxN+Uan3sMht/Ayk5lQlCzQ//YWH1DZrGWGY2g
/+YXVgbHMNW+jVxz/AvvX89eW76UFhFXQaz9MX8jXIIdiRGlXNkraEhTruY2
tdgn6K2vA18UKjiHY/CYPjObNvVbIVCMv8GfzRFkUjiYsBElj4dqTRoDgyPK
+1ZMviiihS/3s+wES22slGwuwCvzPUjWPaSEBZiECf3quDnfMHV86DNmiMw9
Im2Yy02kiVxAK1zTz1muqoEVkteC8+I8vfsPDBW2rMzcV5XFvl02RL2AsP60
Hah167ilfZDx8X8Avaaw/iKMd8GVG1GUH2xUruwppWgwtevNXk8H00WxAboT
HX1a2LAQ/iy6p5Xs3IGIQJuy7U8na+JVa/7Tuyd4HcdbIiI2OQXB5tevY9Lz
kQyYL470qeBAIhYn1YngLoHishIUXuHkxaT5vbv6ltiRMVL6NkPFIZSGeWPi
t/gKoaYQfaUJ0LME63JUrPKjb8DKmbSh6lJxfaSOXrkqQVETiPFWFy5JNrUE
T/6VmB8EJaIEh3M25cYSwPmQnQ9wJOj/8qC/JMhHrNcbtMhsEQcRtJVJtTSm
a21z3lF7Vs/+wlFlgB2mR5lR1iYyHT0ysCN28wSxctLFbyedHWwDIowL6E0M
30RhdkYOaKjwl715c3Qk0X2iNXvC3/PHhqKJgY1kv41GA+d588X0CwG9XxK1
U40/5oaCS/NC33/J6BMJizEJepPXUoA+6MOdrlCK4+SJ0hxRNJvCEEcruYAP
+E6YmNd6LYgoJbWsQqeFJElpf1hpYugoz0PPcOUezwDNlcCQnfzF7BEvFq/+
0I5Y1u49B4w3efQwFGXzhTJNKmAM6y6kbMKRZ3OpMHKYTgTCIr7z6DiPujnV
GoIa5q7JR1kLcTVw/sKdJfo39QiCXJxsqYQ7jaIwHQIee5D85Y55TyVjz5/i
1M+oO5QIM+OQKFPM9jhx8vAA/8HLr79pTLG9c2YQU9fIugsitfGeSZUZuHYH
Wiy/FLEU3UUgYB32tCQNzj0YVNZ0qAjqKAJNF3Zu5gfgDFE9ZGopWuiErBgl
16TiXUzJ/4YeLX2GnII8FFnahVg3vLSWJC2cfnW0qwYZI+X+6TssFUJxvsqe
aSFX5yqnNllSeyX8jrnZbO8w+lZwESsjn+uJNaiH+v4wnCsZn6llfXJTFM38
m3cTFLzylsOIQOoC2PGzadPIk/ZyzU9tchDe4egFYk3hM3/aDF/iMw0mx+j7
u3nk9cDs6CbfF+AAtakpi7arRiQZIxfbsbooDtd9p/ZHtanWixd/lMmOFYhY
yG1mu/C5IWJ+fuGlbNeXuDJyTfZ2HLBmFlGgebRzb/+PhjIrDioh9+R0y0HU
kDatBwq3FDbY9uGOPEfs44kKh1HdDr1TN7neqWuDzyICJRXSDxZux1jJ+eC3
bdgxbvQjiCht8R24WrruXPpxc/rYoboBspDzSsGrrPTMwFsJGrCYvLA2fnoW
73uBC8uhN+A4gWlNVGs+qT46booIrTK3UqkRxEEj9UCr4cpccj6wwgmTg8gP
QbrBxYOiSX95SuIGf9ojAw+Q2tvhOZQ1q2TMzE3FxiFH9f/BarKB7W0hJhJy
uqPsPrVRAqFPtGuCsquRYSwSAn74UIJDydVfifmyETFOvH8kVHrZKVJrlQJU
BrblNGGbQn92vyiGiqLH3bAmMSWCeSAHkWd5HXqV777TnyK518f5rjt9cdPD
I76KCawOe+7AYYyqzQZEmKW+yPe0Scx/jSn7/jpzv30eCK90+n8h4Tqn+9Py
woerpUpLs/lDRtcZGpAt8Ptu8N1sG7oCDpeJKLaZBal5IvbqD/83PMql8IY/
cx9jW/Oq09M7hAyQ8yisDoVhX4KxJdGeXdVleorZbzgogffUs38/A7gnHgDc
9GN+gqVXuxevhksapfTEzmW5AJmSbhE4nogMo9hpEbqVPbmQOp3wROInyUIo
Q6vXSsLsZmtByaMOdQBA9TSHHfioVLdHyoWjmMByBG8rvLO9EpPaKfOOiQu6
tjeI2GLmjhQurOHlbvjBaq61tpwAklWCil2HtpduXfBH1G52UaWEpqEseOnj
+vca6Ax8FeT40JT3HuB4XS17kRoknRAWslXsqxM4kyfNxUxma78iIhhTR12U
s+QqV7tds0SpEiEg196gb+ke0HkjmeFjCQex2vIP0aj1zXiP/x7ALtlWygaN
issBsIaKR4JtharjVU3JiKN+RQ9VDIlnvK0XiyMpGp4mOfoVh51fSUR9Od3u
oD2VWNdhR454jxN8Qrg0WFzVhQSVjbS98+7WY6WQ8d6rYX/K9mXxIm7vlWXj
eCGliI6dA8K/GO4/AZ1Z/EQ6+0Zt6FVWeZfqIzXRAhsJokvrUVfyVvaXdRfg
5Airi7A9uTzeDlf64XZ0xMdgDaXpFNPpBMaahl9N/rrJRQbFTlKfTL81Ay//
eryOZ5mJB48EADkyXX25KHGu8jLTmWna3tQemow147qAsbKD3+dG3fziCc+v
k9SDNnxOtXBOGB0aMEvh+uE4ENdVonvmbg/9S3PNy9qn3adL+LXpCZYYIk/Y
P3UA3TUC6YB9zORIuQQrB97NdDGKNcVgAozI7xrdrgs/JEJooTljJbGUMPfx
8P1OQRPmA8K3bTLdqGIZ1HcQ0fFBnsv1a2kQV8n4ySGHJD5jFXwQAsZyg+Fc
ECLCja+cldlDxkT0UdcHM2ytsKeLyeu4xA+anT8r+1hmoqa5yYog2eFS5WBm
FevJSuN4JBgIBdq5Nww5RGkwjJOofpnuX9osw+mVSYFLQ8Vld13Hx4jMvem2
O6zxyh1GTIgz1e5bUt1kB8YodcHwyukoEH54oFynl2mqL63yGk/YT+P/sguQ
GoS1e0p7lek+lm7p9OCcThiXn7m5CDn2PnhOuyAxX8E89jgFUn/eQ1Ntzbja
UOwqWmTnVAIXctHypObhHwdNRlCyoyuqMlngyhUNrgYJkbcf1Wwjd6A3Kh6j
YQm3G9oJw2sv4lwnVAqg/reEWW2+MjB1/gChZCLdRrRHRFl+6MLM1zQgaPRn
nU81ebfxXwudOIrioKM0DRy/mTzgiAKLxs9dxrF67RKznbUyM7Xz9Wtr2zRt
7f4oTgs+gI3UGCk/n7VKv9wGkY1Vs1zoK5eUbreG6mFtFfzuG6c70qCpS2dj
XrIc8Jj8SKG7yeO9wdduq5oG7pvYeCwtK8dofRmwP8qXJnv94kzaknJq7oni
leh4Ei0mRjSPCcvFoBIdRxvZhUYyhm6jh5f60KVcws/E1qPGHrEoVdbJaQJS
uI27WBNxHcmFVPR6gmT5IzAsNGAQU3/fUG6RG47RVAIj4n69HN2qh2BPegM0
t7BSfdI/iOaNRCNc1I70S+KRqLOTSsACEteuzmBft4LoO+YpHvrf5oHa4HgD
fXHusAoOoRZbtMy+zVB+jmMFaTm1DmOtjApiz8sFp9wPbePCZ1CmfOu4Rd/B
qphQKZIVA0huGA/vC7NrKc232B7iNZh0DtDyeKABhHHm84b1pmAXk6MmqB6+
kx1hr/csB4AcDvGl8rQoj3M1YEgqxqxPp60bhUFm+ex8CSF24Gg257sLEOAu
30ilxwleLx3vQY21lir5eQVAtxMkQO1MCILtHL0ztymT1jmujcq7wxLPG2LK
H9ZsqkTCxQkUGbZkL/CckNnwwB31ORtNg1ZBR1LBYILTxp1eUGmgw2sk4OtY
qNmPvr3xeqLn8/0jWqdKl/pW1nvz4bssApYwRX2qtYPlX8uQFUXinS+VJ52j
iljRgG2Gtzrnd19598h3xUcZ1/EuLJHzQPMSwCOxMiM7aTiW9br4SjdW8JlT
KjZx35c2dR3iDBIbggOxE43Ua1976CMDbO0axFZa8Y/LdZopOrQXMGsB6/63
75s8n9jZ80HzbMvsawNTXWIGPZXD9HL/ADoh4alYah04J/CvCHrCEsH16jNP
kW3UrNTQoFUTU+B7fjwTqXkjfrA/Cd71vOIFTPQYFlEJkg4cxxU9Al2vfuGK
cXEFkZ/RLdhlGmBGUkBg+wt02OjwRg9NKpQSSogziHktCd8Qq/nXp6QvSnYN
jV0M8kR8jzwmnIc2sV2smiyZY2NT7SYwfxjOFD0ISjc5QZTWbrfuvgVu4iwA
F2q59RdEwasX3ee8QvThvadMVfZbDuFoMULWl13KTRlDSFzjuPUTO2AtpXgu
MJ6kadaFydH3rSfLHI5RLLz3JXY4Au0Un7X9lfqUWXw3s8zgw8gB5R9e07Tx
s0ueIdqTc1A6eedTHHFLA7WFiZb9OW9L/+poM0bJcEA+orpMwlAp3MFlnagW
4xkUCSTUAeIxs1s4UNnvwfYvTOwoOlbl7yWvDkoSTJGLScOAHA+x4KMocuBX
iUGBZ826xv/gtRbAHgNr4BAKlTj223Qd7iXCz4QyK6rMoKhns1WcAQVxrZhT
9YwI9C4++PTlKfOAbovcnYSpVFifJQDc2EBlt0A62q3nVgBuvu84VOPEtbgJ
bhuVnTG7k3pHMmC9qcdhaRddkV8LoT0rri0gHOBijXlOYYC2Hr47c2Y5NBbp
4wmeZ9Lmpvtg5G6HSomJaiaOQaInJe3SBYMyfr3sRn+Fs2WKXdFxuInFZi8v
0kOhKXqTsvsO3dSexvBh9Ide9BahWGtbene6oyQhQXa41ZEkt9neLteIXu4i
iM6grqbiwecbDlNfeJziF6S7EqfGNKKQj/1C7NohY9IAJp2y0JRHs+VqVhgi
Ak0Sjb2Aapd7ul+xX7dLDe23wdv/4bP1WTMrvbvmPo/bc+raII5hTG1CMDZn
Qvdowl0Gl/bCkMMK65Om74v+JWFkKCt3R4knhuMTBZyjEWH/uNYFrE8pxwup
c1DOibATVJETgFDwMz7NWKDy1Oj5ZgqdEszCZaMlSpCnecAJCvhYAJ/rGfe4
o91oI1hZTUNpp+N8GEURIYk9scK0HPQJ38vCrm03ve+lGdFCU4PUxb+beE5w
t/8frcvQvrgBC65zJkcTf5u6hkT54fUr96fP8u0PBqP4bCdhGCJ6ElNTOm91
SW9arq9+zP0uOsGkMewP8rZ5bxcieg6Z1uIQOjlGRT2ej2JPzCmJf4w19EEi
lniI/yLagl8rT06RKrNkDKWtfvMFxWaxhN3qI2R2SHKP1BSETzyWBHdJbbxN
RJlzhaQFrGM5u/RarGlvtFOj+b9BypjUUFWZEFBW+l8FKne6w6eZ2Ho1xS83
y989cHSQr2n/eRXw493ggQDApJGWwRrELNSzyyL1kO8ZkIRWTKsg3+95TsP/
wE8G3GnxXVzYV6Emn1dBgx+JQ3R6sRJOFsqrS4ljWB18p6dsXsys0vPPTfc0
+32vxdL8SyoE5N+0acWabtH3BUO5xOj4DWjeKng96KODEpCeyh877S/gUthH
yCSpFWG5NdezfEW59S/QXBAUmwnNqHpf/NyBzufr5bJdMm+egmNjKUNGW3Qp
6VzH++gknJG4OuYOOl+2L8a/gW52l3pFKiKbOBQOFDthk03P6FyDd9Lvmc7X
EWkvbjVEw+h6Qd4sBPIJ1a9UF6K6gnDA4tjhz3Ub4Vql8LInH5BHZeXDzFdL
4FFQubS2IHwms12FH11znJ7b59SFFhO/joDV5BjoC2oxCIKMAdIIQmAJP/OB
zvOq+aT7Aj0MUGIa/mgkGHy73fZvuXINGZLqFo1pC96OWRHF1wu7HXNGYHn0
O9i9cEk38oc0iXzntg+4MlnVqWie5U2MU5Hc3DIiZDiq/UUfCl/xtbfPCW61
Pw/iyH4obq5ndoYlSsM8pqhjRfHYxb5fcRHMtNvJrI6nZhNy2OxoxdCiunN6
mnVTD2JAN9gkYwWsqn3DrdWWyNhtGJHsYnWe3TKKs9KJd+wuVHQGboBvOZz0
QfWE1NSGCwlv41cJ3hxoN77d6+4XBOVvHtDFddr/16ZII4a+k04S5CBPWVmK
pUFQASyWw4qg/uqfvd1sXLvUXGqJajjRaNtppgprZqqMSDZ4y7N3R3lVBPfL
xTZeIS0XQwlPGm2M/PRSFjBGAhIZhor5XljqpWKnFD6NmfoIXIs1dxAvDswf
G/NtSgs2XH5uMnDcDiK1wDNmPc2TfYa4DEyBJeolJmDnHPJQn9ELZCnK23u5
hJCGUOZgAFVSnJcUBsk3dTrfeAJ1RO8Q0PWtF7upyP9zDX+EdqOmEamPDghW
OT8p+M/mti7vTUNVoSGXFaRI9BCW7LpCFGEkZwUaeTHoQfgyt/LrsxQ9Vh0S
0uzc1pkrGv27hh6Y8M25+GC2lQbqWEMQwgH9UoAYV/4huHGBRgp4L4qsfK2b
PGrgDc9KV23hQNUWkUoYpkYjmpOhrLoYiFTeT1rjgNCtftVV1HfZhQj7GIFD
Kv6NTuvcigizr9k/lk8HzVQG+/7cL20OXvMqyB+NxwCEQzM3fVTPm6viLyeI
XXUhLga8LSO6eZg96sTm/BZ1CtYR46lX84wJvNWEQxd3rxMXNiYwRNYl44EM
Npgyy64KH4n1FZlzVs4yCv8wOfBkljwnXpjjKF790cufKMRa5mIalckD/9dn
w16BCHMjESnKUUo4a08C9wAhEQUvp1mZoCOh2H0zMq0FgA5a4T+TuCQRjwp2
FwhdZghxye4KR+SAX8ZPHOseAuZXZduXiUT+64qq7PvgAeNeGDFFiCz84O50
CMii6IBiN9DTwk+gAaoXD/jP4UfJSr9Yw8XWsbPSsiu6tlATUwXKVvKLnvN5
WJ52Nb6lwpP1MKvwgyR7JIK3byr0SDzJwTL/ZWQfVJo2/CDi2a4CuA6xLgqk
mdBTGRYJuMyPcYxDACWdQ4cmTXNiLz+o3sbt2Atw0K3+eWH/5rc/EAn0FOf4
3nVvLmJ5pMW41LL4srssaEYo+uPHKYbvSu9PprbSz5Wil+JaOcvof+tT51iz
MWrUQGIDiEjETF+7FreUKAy1f8ofcb7PRuCUnpShLpCa3cbrbj8WGedfv99S
7euyCup4h/GLs/+XwmG17EclNaVn9wGp/Xdfzzgzts6fcDvpj0hTYrx4rW/q
i86xHHPahV5bBz23CTeYPDCMk4NhSvtQa611A03/DRCw1yE44Hqo0QJ2odId
OjS/A2o0QNFslzHNdd7epFflXyklHgmI6CSXSNg0m/PmnSnX9TLflVIxzrWA
v9Z2Kq1eyZrktdVapq+j1szDOhUlFFiFx4Ysa0RsqKU5W5OfseT4UvkwcSdy
anfEIqwQ5ldimZTZmxsLYopadSSv1p4KCFP/KjumyXhOeWYBQfsDHAowRHGd
ey3ppQduXDYJo4z8lKjnYVDK3BU6S0gMUR6ZvGq/yxen/9sXzh7ZCaCoEb8A
Iv5XOcd/U7N0QN3r25XqElZV2fFVqEVzGM/lbjkoTIPJb8tWrpvPGLYjz/SX
XdGzOkp/+T6sVO2qv40iNiGyElL8IDDjV8MXxatxegZwZovKNgXH+LXPahOx
pQ1QU5lADmXOHn4KH5P8wdrHW9OwCMtZOr49cjW/my0aHfM1vAcTuwc9PhZW
brFqcMhteQFok7f1knI5dIl3CgaKylY65TwW9IGUCqXgs6xiYesSt3dfVkyW
n1R/cq1T6Wyu5KtfKVe3kA/luMby84nmjrtWKwNUyRceE5UU/LLuLv+s5jmj
2jO9vABK9gozKxMMWav5KIa32fwE3HLOd2FBiW3HHaASpQZ0BREdDnTqBtJp
eMXU3lB87mZxMAZ0tmhrZg5bBBHqNTwYtXnY6D+O0TFpUQoT8k1uJ5ra7LV8
LLIkbefbG7RL9AosOGFMknBmGdTDwR3EZBorqWR9rBDik4mYsYNr+aNJ7x+U
2VQb37TsCrQhpJ23mMnV4hcH3pAxD3jw6aupHVG5XwSLA83fEH3O3awOSWAj
TUDRNUTYQmZcgDcOJ5DmjBNXue/lzGNSmOkm/fUXPvbpVfqDhRi4PYImeIg8
f2VyLmBxv8Z4CQM4QAFf1f489dQSMnNr1Zo96yUKar60vJSrYUfB6hjNVwhf
rovPydNH+Zdz0VSw15oAsROmE2wEYaO7oy4UGUdVrpMOKsYhHyJRSZthEz7j
CNh0udlc4hacwWIlkjro5bZ/+vUzisbII1UK/66NVmVYZAoO5HXuskAcx0eL
Q3sd6H6tm3yzox3BhTnU+oUQmnE6hYw5wHmQuYWlOLDzdl1G2/2bDeFwTvv0
HHoz4UBLoYbXRZAsETH4+bWZB+TKgO402TxdRsrryFdMesDJ6r0C+Pdl5Txd
BmC6aFBXGrYSu7DDITBeYXMCgRzjMjQVz/svXGErE/0Ij6SWHzmYywbjjPxU
NTffKqeQ9eT4mVCPCWq/q1b5FxXHsHkWRVKTAVWoAuUhuPHExSJ/x4gquOU3
1Vs3V8WZ+mEJ6RhwHZMehUkZ31kJOXNhiI/mJhtzgVS+94GynwTkZHMTggSU
v3vb8Zj8U48MjDvhNiOz0hPKBPhE52weNyot9es0zPXU8+rAwdgcxYwTtaa5
mHtSto+qDvicfXyyaNVfxCvzQcNJQXPk9cXCsBxTaL1CEkBcYrCGSXorA/TD
BxQjEImUxnBrzgCyjyMU3whiWQrKDw1jhR6O/49xbLW9J47lzk4hpuQuxz+9
EN5qjc7u47tQTFHQ7vtFDe9srNQS5+KvkNpioPzyCOcfQJXui0U8X8S5FQqL
9cXlfma163mkjicFeQOnUIyMu9znsIrgE27pONmY2/GWfUrjkCkdpOD2Ffmu
oHweA4DjhhaWTyjhIb51ijvb3EvspiweyyRFh4WOv9zWeNAm5GYWWIt2m51k
u48qCpwQVKuoU8fvwgHCMGth3pMdDeQ2GFEYYm1oC23oSBMWRSF3jfJz/6ID
q7Bv76ECOqGsbV7NvkTkI9w/1FCLHkzfdxcyXq/m2Gi1/Eoj+TR9INXOm6MM
I0s+gjq8nJZTk6GIL7BafxCatyRU2yA2/njRaIosxN+NV2rUc35Ur1mDWGzo
p8JoC96GrrXAW5vRqdWwLP04bwLGjABHr9pA9MH1BfHilwqH20+N163BWGZD
PJQj5bfFd8DC2Md71b0uILiZqI9pAX6NizubyAXihyJ4kmHZQafMFnO9a2nc
ftIKkwpdDOXsDzGadn20TPoAF6cUQI9wh63Y+UoVcczIIsu6z8Ib+FYyUUAI
ZNMXlfv4B3Vttzi65XGaYlDk+2hcxLVVyRdq+YoYdPXKyPt27vhkm1UD7ckr
wQh86YgXqER0poEsCJaghnUAEFVloa8VwF+x502/MZiBQ1nwMsPHdllovIvo
lzpIBPmzMpJgqFyIbSrNiV30PYQlONA6ar7+Hq3MmismJzYcpv9gUOXoX9li
C/vM/z3QP7h3KIGuc8STL0+dqe5XXFTkpiqZQl1eD5+b/XYpoKthgqAkR6v/
zTD2a1aKHRTJx6h05H1inKK04fgEMX4T0pEo6L9vJePV5C07iGK7X6PF6e7M
mTT6PkziJelSNWA5DfrUPEYX2P1+NLIFRVH7oyOUeL+DqiINEeJvkdMlsZ4O
P9wySRar2kPJPBs/TyXoteejadB/8I9F3/HPoR8cht5/pS4vClJnUr7eY6rx
sKk75JrkGgyTST9d4tRdUlSJRctHm0rgDfjwBjTewtsAD1H1mZUc6oHg+U8k
eGUZTgKYgMzvgQP6O7aCvFionK3cCFhckrDJu6bOZdmsDFUzZp1eocT/nHzS
zrme8PcLzw7+eOXtHh9sm6YiHu1ygxAwZ0o+vmWkJX3jJ/8XBzM9zCSQAZ3R
+wRnnN5nN8dJiqg28ihcJKWmFtyF/p+PIOp9vj0/G4qmXjarjekDLCdk7wDd
vvMYl1b8zBs6J3rR26eig0a9oTAVQT2SZ0u2dO13cyZzi4H1x/1R/PbCwTre
FoFYEWA4IyO8/Nq7PAn3SHdW97u9aEcod3cFlhWMGHUWCc8KeGK2TPQqUjaw
L2N9OYlDw06i/X6u4Mq/HndosXdIHmoaqj1ns9wvlpdTMXjHwdch+PpGZLLA
uh7VMc/XVDSYRcxFPxZPH3h9Jesvwf7xOsYSGY8M4vTHQ5mFB/tV0EjKpNY7
xShDeUusVpOpuqXsH9aUDIhUoiPA0k9RRlGhdeKgfTnWEfM/p+7G3uihYTbc
Qm6ycyR+SYX3ao779uQ8Eqky7lHW8allodCFp122teliOp13VJibIMnvtT34
XmtA8Ad/LnD/7S7HmnHSRvcS1VIC+qJiYpMlZMUhl0fIg6xU7XIo1XPCr/RH
givUCyhCO4LwVCWtO+6z3rlg7hTb60SBcDjUiwAkiyhwO3GFV9JWtVjkCagQ
YX36rIScWgLiNkIDpcbKcT6XYh5qcjPv84RN555aiNGX9xTon7h9zTHRcwLT
+8iojrKe+yEMbqXxW3qaojp9DsjnHCULOyWofYFGWhqDapcdl5tv9AH+SExO
2LbY66A+wHyFnwy/EsYzid10UnB7Vs/6po/bk4ebOoYPHvfLARQ+aGgA2gH0
gx3EGtVk2myZYRF27W40pKbd2gGdsUoXCuoqLuWkZ8L+0rXINMvFq1S9Hc7F
b7Bem4K8/cVG2KqR6+ZO8HcrdNZbDvt/qWxyUho00vdZbDA8u0fAflI4kCrm
sQp9smq6nNxlcS5UlecKz3CIdyxC0QFRgHIEya4L8lH5PUbHGRPBM92gXFHt
C4YfD+OGwRyrmqE7Iw0YbS6gjfEag+Om1ZB+OzsPqdQFCHx4WMUKflqnbkoR
f6wZW1STWXgh8v2hYRgal8L0U2xNhqi/is1LMSXA7FwbM7QzpdoYA0G/aR1q
pmB6245k/qmjYQ05NZzUerqK5H9WgaeUPtKHNS8vQTpGn1GHvCFB/Q/xu2ju
fEn/XuxERL9pRLDzenV6CCuXVXFew1FgSHv2Ejs6yqPV5JbhNBFQritDq6Y8
eauIAtrDNPgV4f2ZJnKuWdZBEzmDOqlPAxDSUTcMbg2FI9B+INNnQ3xzj0R9
AFkxb+28t8UQO9nIlbZ/8bb3ORXCwGvbAExUCEKMmkNHp9PJH8HQlP4Nly/W
GSEQ61+pz+vcmHnCmWsbQVOOFzmBQ6mDHM+cASCNtVFz9IaJzc8QDalmv+f1
3gnglM6UHj8RSNB6eAIMixHoT0oS7bQKzzL/xSFiUVVCIHK85CtOmqqhhH+g
+prUeHMGePE8TPEFXyl9035zT66Txf7/4k0tjTcsUqwNXo1YOnZj/+5N1ysk
AhMamHWpzDAfTqI6b5uYbDwIArCXdukVWfFyDUmwpFxDqiBz9zXpehAeLXev
vLRM8ej3f8KCFkL8ScDmsUAPcdUoLgzrawJC0i+gQMy1ysbKqoTVZLahl1Vy
2kasMLHnMXfYmf0v3Z2AmGLtFZwE0BOI/kRJ4x2DHqTgJqAEYlrRrIIpp5zR
5JBYt6oPG2gFyJGQkK0NSs3832kyOFfxEVDujq0L5JBJtEJf3K7+XE9TUrVj
JtbOlWIzgiQUOe7JCz/vDkWoc2D0Uoi3yJoDeEpn1yEwCBSrqf7JCh+ccFar
54P8Y+CpnKRVbwSzCdXm8wyZRIVvvo6sNS1sG7RdUJ0rq642OrFST5JPqWvb
2msy2K+J0FSh/cP+zvKrhH1rAZlJqTVcB5jpWtVmM4em43m7Nc0lRo7mhF/S
y7DMrr5CmK5CzW1dP69275RI+q9XrqKz71kHgYiHgrS9N8hsQeGOFA/CIhwZ
tVm1vb97GbO55CkFQkcuPMfPJIrFTccccptC1zC2GZuiCfW8rE4l0RR9Rs1l
wooSmmapJATJDwXQTByDq4hKDn3C1JtblKc1ET0nFsbnrow+wRovcH7qDOkr
XA6xhowHGr8/MXs2+3uF0Nv8OfvIuaFfpWDT9amTFPdltjzdFB9dyTrIcLx4
cslUsUcjQA1si1le1bmfAd+RzZYvsUAeb/KyDCIASZwPdxAQY55dkDKRVlZm
/MRNYmCGwGKLx+EjKsAAY6RjcAfLKIckdix+pRgmTrijmBjqWS2VaDQVlodm
1/OJcxF4DCYqY5n+kOj2qMsZfz/DqkJ2GLkdRKKAUYxW30o1svGarNuTW5ir
3s/diRbEP6P5Xpwzv43LFIqlYp5MIEFxve18nKkyac7jFOOHFGSeVwoxn+1D
iM8D572hrIlTzXhGUrn0uML/F3rqjBF+BDLySrRj2qftkeKGCPMjRYKvdDbM
DckpkPdnGzpEY7bFtk2efdGoLdvMJaLV9gpJgOgXsAKOWUV87OJbpXF+hW9d
qFH3aeZxZzy7F+p1p2WmGUcj5MJrL9RmEGEOU4vwSKkjhngqOgJOvdhCHkPW
RYQlNnmISuAuvHUfOofJwJ3TxQUyQ7RoYQe/Rgj0180ELoFetNobcUzk9Eeu
OtDZnsr4gStjY++29XBJzKTINq33pRIP4m6hVhwfDHGK6lhPU/C8+we2sH8z
7AHpl9vjAeidgnArJq/4ySgE3YPwt573Os4wNX5IzwlIzeiwWgnZMtMMvIFn
NXfOY5voCPbb9YXkqcsEH0bn9otVmoFi9abI5FxZL6U0Pg5kT2TE79Uu8a4Z
xRWtrtCStoAWR12moF9p+ISnFndJvPJx2mYUw2mqGradjhSAnh6vE7LxM1Pp
h9RBFKvtfFJnG8Ns4Vjv5OgBjw9xUZ2VI1f6id0D8tELPnxpgkdmT4Jg6+LF
QESpz9HUQLp7p5kdcl+k9RSuomzwZwz/ZfGfwuGiJLYl1wyWXktXp9dFISwZ
JnDOKFW+sjfsRaIwwo/tUf9fM1YZqMpUCAxi4oM31XvJbspHfEWtTQVF9QDv
UlDFSS9i33u4S8mpcpMYNPdozDI9qiiDCxckO9iWYG4TpUkpmlsx8KQZ8jMi
etvyiBPlEy20jn2XXIbVX6UqJuMTRC2R8ZrQ3124nfELhobdjcjF5Zvgo4U9
cdffJnGPmrd3Zp+IFyKXFqcGjp8mmU0FoA0MX2L86lXOQsdeEZhuuElrcCUP
x88JKn/mFFMt/tBfNcr1MyvRHhOZR2RgYY5UkHJk6umUIxzGYH4V93au7uYQ
/4Ll0TYJrhEvV4hNm8GyDBLkLd5h5DLnH3z+LmCUd/vNXkfbhHYL4MfyWwJD
wn072l+/pSYU0Ps2AeiQVOIG2SMqXZUYwmGufUrSYHEum4By0I0p2Z6GMx3f
2oAEqc80pvVTALrsiaIXXzbzOLKnnHxwer4vBfOO2H0YuZnbNX3n8RYWXWBg
FcaDKLKtlriZNhUxZGTVUut3FB78lnrnBY4XcxjuE6sNQuGXF8cST6It0WyT
62PH2VrFSd3XUm3mX5E/+vQxpj9rZI/aR2tuT6LcSgVaE4vttMpCpbL/cZmB
8tUiREZ+sAJc4LmfNkvODZPtk+Wp7XGIPzbUauvjx9vEL16SETO676B1P8Mo
VkFJT2VPE8i/dsntHVoT3hg+XnXRpacF/iOR6ojXxLK/xnvbiSJ+XAAwps6M
fRWzc2UD60BH9C7XTXnKbysrE8RrhEdrNABGcrcd5Cd25JZs+5ne+/UWv9rh
Qgs7JfVMyZ33CQfgistHHRoBh9xFlTmhkR9Ka9vReUavBouJ05VZeHRWxXz6
uL06MX9WAh7MhyxofBLKnfPxoqQeSbtaCz2fVkYrrZ4E1NFENa0IdTd/1Wth
7VtFf9eshr6nRXbrstYtyCzOxqK7DpuBJdPDGHU9hTUVYxwlessFbDt+14l5
xLI0Ti61JUnf9TB0ioiWf7qmH8rEDms+9Kqkl0LPKjw7A3FNWoO1e6ynAiP1
fASIfHd3SVotfviZAxwDEvwSJDW6u6i+lTyPHtzf6l9XeMcTjnY7iUL3YVjW
ODgPOCPiGRqGh+F19+eTla2+PBVlDKw04C1hZSJcd8vxtKWCd5GkVCDwiGPB
XoKzLJ7ii0ji2V2n9DQ0+8JQ48tj9lIRPEs5dqDEBqaFhShwFkCaWuAYKbvw
iajIOJr6V6SKdle5xKQMHDVVcz4OUSDKqzyKX2gTLKgncMjd1Ecwrp6/uOhK
2iNFMGa1MoJJngfKLiSHJ9dtRQGAYORDbTsDOGGRy1FMoEQ7qZ2Igov42bsq
G3SGHm+Uk4AUq/NrYLY7KTOhnsJTtZMsd/iXcuX7zNvCRje0XER96OrNpa54
cUDaa0v2fhr8mh+kl62BcMwwdmAwYwjP+E1A8s2JpaVM39bdcGEwf4w7GK3b
KuyIRXmGepJNGfpW6OcF/Jdcg6zR8JZmlH9KQkM/9BnBtWay/biwSivDQ779
IlOsFNlluvpS2oWxAN/aIrUrYtiR0bnUbgaR0lUDPjhFGq/6eXUdyYzhYI8/
eoVgiERFgFJTiEeUOkoG2VtpLK0lIcZJzvEe1inoho80I1cJS8pXwT4WtLqU
sY+9n4+OS7uNbOoOVc5r+ZQWAfWVg8dsY+vRnKYgociJvc5wrTZgtJVIZ0Hh
vIBskIwJoOruQUdCUoPcsQ542Rtt5R19D1XqOfrwwnEO/pvTG9Mpm+0rTj8u
Xqj42icAvKAjpiUmaqC1VvGJXEp8m5dbl7QvnH6w4AAeIcFhJc7ZGeN218KL
C9H4cTiX/1S2p3+mZY0wQVj+c8aRCf0dAsspAeaIdfkgaoUAlU5YPgnBZrr3
REIhY9z36dvr1d1sF1sNQ9xmREdjjFxzu9U9UeCNYTiueEGZiemvx0vuYXUF
GLMysnFvGSSEcLZQpvkyVKa0+AjJ2weWDpvMi/igmXirzknoMjBDSVMWo/KI
i6TqhvAftWu+U0eLlvbnL8PJpuyrd8A0XoI8XEQOj0WiL6ONofL1e1i86k6V
kUb2HVB1Oce004c85Tn0Xn6uQA5rZVpZD5P3OgfqEFGNT3bAsBgwjD3fpDo9
MScweJHsEEldPaH9F3FyoVPYCrBECCGEvp5dBm7m3kJ7qVycltA8aSRgKHHf
UT2E4vCPw5a8gXTPloTXtHW2e5fleJ2VdE0kq8TusHV50hxb1R7knXzCK9OK
rICRPQQx1tMhyYQV/0YwAhyskaUSBODyuZ0680b0vDdRLvb91TlJFl+GTsVf
4fdYigXHc4lP/K1HsZDERP6TDbZuHQfHWiZHT6zY3XMOfzT0hKNpnVOzoQYd
/uatZAKuZkke0meJq50iq6h/CWCFWnGQdomC1cV1lmAhoOAihJ4nNFaFrPgy
NzLDugjvcXtTA8ZnyLqTJ6xwj1zN1aCod2cA81XvmXmSuWDOOVi5fP0BYJIx
o3zOB6U9BKsrffrFWVD/xJrFvg3euf+o2CLgjXVHYxCo3Uw8D3lN9KJSXjdZ
K8sUMVkPc2qo5P0icYKGhugr9PY0BtV4ZAFt4QGTQj6ZFN9PLbemdmKhmrpe
74zyNxa9ejztlAJ0tWVT+9cZ+310GcI4ZpOrFYBzeC+yMEyvMzf3jE1O28mR
O3qdWj4GEJFsAGDcNWNLd6UPgTfHZ3Yo66o628zlr61CNHLZLQkVyRf+Bx3M
MhEFmbl6n3hBOm4s5mFThrMareLkk8zmIIueTwgUO9NwCDxOfxHBOpBUSNdR
+UJIEjXJhUmDTKEvEltOFRCxEHHZsuoCsVu+sbKUeTsB2IEM9IJB1JQweEWT
5yiR3Cp0lFMCHsssRSw8/tQ6c0e2Wsxq/RZFfiUoap0UWcErD142iJxmDpr6
ywZpVXpVfK+eHPSclxI/8loYN/927KLAbUkp1O2c4U7Zc2z38vJzuSi+77OH
0bPq2WDBy18ZigkNBBYMmj0q7oZQ4sDz04DTbvyPE85CFu+miVEVdd9Qne1S
IyJ0VJm0ONTAVGAxFpIRa3MIaNt6MtWCVo8HD1U5Hp4+QmSJEQha1fJSmAxE
/2XZTsFX6VKGzu/XX8XjozcR/RWWOvjYOPPD0S+z53UK5TklvzNn1Ght0FcW
qEPVAw8tsW0OnbLhFTj4YnwVKCa1396aQP0hakBNSghV48+gNdla+3oX1ChJ
W8YnV80RcQBBq/OcxHwnc8scmddzwvsQCW9Ta3HGKq84VHjNSWov0cSxWokK
i1eWn6NIANNIdginvF+0KmUFT/zlNP4K1pyk5l5blHft5rrulfI13T5b2deW
A+gJUinrYJ+yfrGozgdX/AjUMMeYvn7AYk8/ywA4n+H626c5VgFXBESABQcI
s7tPaAOSCQFKnpX9IrXOWnqg+eEWTV0rnkhwzOPXYLVq8QWlCGPogd/IsUJU
FHou5pZxdZRjMsKzHil5hK5408ToD4Q6nNQNCVqq481b3yMv5sCUu6FPYMkz
5br0y5yt99VVhxY164jbIHwxhrnplp/wezaspEekClBZXn+ID/7H+bm6b+fp
hTp5SOeRorR65AmDIz2sWKVtapBRSXyZmGTbuLEIThBypK1twkIbRi5w1XDk
N0FSHexid03sJ9YqWTysL8Si9Nz5RHtKwxpfRYVAO2BUN5aSQ8ghgkyjHqqB
IdGnpKAxrgcEIh3LWQWm7Ja2gJYJR0KMdSUQC3sELDBY6LfhBVzLaAATNSWT
LkLnbd7WsVhYYV50OX8WogOAlEFovF/CYLNgIJQ0UJghrth5ri35wEAYC7rx
w41mD2/DHi6zEM6VBZBl2rZ+Qj75HheZnLZIcJLspRihN8/SE4GGTdkH0Jxt
6R/DTtRl5TdCVHQRiew02xCh0YA0pxrUCiCEPiVISTyeyZ8D5M0ttHYpa1Xh
td4HwDIF8Un2/5ZshldTg2PDRDrr4fvtzx3IqgBfBIs77leBvs9b8CNLSLR8
pvpknL9h3BbOViwbtFq1J2rjuNIszcow1kiMq3lZ5GQglRweYDWHHPVO2kuj
GoQmK7BZJ/YYeOZsNlk9qWk26qQedXynuAGqKCGJL+jM4PA1fq2D85AWHr/U
TNFyWf3g3K0VGVb1ukFhyHIPmYsUrs9zAeh8hZk1QBa0JksRENqr/xa04L2L
4yxvgXY8wpfl8SainDmhLCFgXLhvdPq4Vo6MwPmCfLw77Gs8zKSLc1/JDyHB
pdjpJkdk8047tT212e6IMK1WkoApTr4ZoieOnvfgL4zOPorOH+PNytmVhqfr
9TBw6t6xJ+r4c8rxlkoZFajSgdH31v9TrP7tb9KrKGaCFQRCJtPKVVhSy8JB
67pY3Q7JYUQOsahC5saXEde2uOlRAs3Jz9ep9cRsvksJmk9pmOnpaO/xGKPr
ywC6MOvx76oAfosrAJDpy68od03lQdihrO4vRaUWy0skFZ/FLW0FDu6ViEoa
lIUcWfU5tcHloZvxG11aqSY7aEOag/GSw0rMXfMUvHO28UAjPdcu4fp+PyH4
1wbSapJGMWQZJ+KUcwJmwpJt5GLxxooey6PLMso13SEIJTtmqTiVxURQQJ7w
vnzxbgs6UBueCsTFtEa0lynP3p8ixH+tBNnEwtEz2yWV+v+3cYh0dFZjVEqC
/VHd9R3pSaId2clzYOrkA/HUPCX2KbtB2EUvNRGQJ91NxlrBl8TdCnTS6inv
KcCy+cObvR33KX14NZixdKymJo3Z5TpPeW33tcQpHNU8BHUKM/3oqeEDwtb5
B4sOmIsHEfMkGWjiv61tjLMx0xrcoMeG4tpeotszj7Kz4BjImrigQPhLHIcJ
+4PNOVe/r02ZcBHFUautFsHpYPW/tW10XIvcARWbAIEVDavH2ZxuJXJrlEdi
d4EQ5oe2e/EB/B7u6JIKfMbFXoB4ELRAPzmDBUsNxV58bg+WKhukKzzMrZkz
JQl/IeW3wvx2K3zpcIznCo6QPaE2gDsik2ctATwUgetlatJmlkLLmPV1+HS0
TJRX7aHRUrw+HaPW0eUN7lr31oCVR14Le7mLf9nNjUFoXtTweYUp8+VW3qRa
McyxzFpfDTmgN0NN5ho2+22FWxbyLJtmfXRYEj8duvkaf32T3R9GdFST6jpr
UTJnZmQuAunKTdRlbKTIhM9B/UawnSfVP0Qe0rC+7QxQlCz+fSfLNi1Da61E
CMBYohx3TU2Y/cMXNCRDH391HwQZNbX+BKscnbh42M36dm0lMHJFqY2DaIPY
LoxW+9rBFYEZTJ+iKsdYRI/7dBM4P1CKl71AS5fwjlWrgW5suwEBR+N9k1ca
ZY8mhrM1+hCqeMJQ7iocdsu+00wDikrnG01ZC00pQ7RiFiKNV0LntvbJ1PXI
On/dGkGExqw62sHOXGnR8oqxk0LTa9Ith52uihe4GjbBoBMBgk6WQDJXjaNM
ctpdoYuvZ9qkDq9kRzmQQZOOS7xnRHD62WVbu/5zZGX/5Hw1QNoViAdmfQya
C+4A2v4wQr7yvdqNQjdVXvF5pT4T/EQTV7LWI7zkfrxdcnqmu1I7r7CmS2BP
tmsd1DCJbl4EKaNxdFBE8ebPXrYhfUlTrwDwBPtIGkOIG3MVmwNqxoNlWX4C
xSSE7JZ7FGgb7uLxjMs3f99XT3GWjMebeI73KAg26iwlMjSlXlfq9C9QHbYq
cConmBkhDNYUdv1plLj+Aul1cWPD5w3P2W79Yuoq2X5bWJq9gsfgp4BZDwhc
2iA2r3oI2KCJ3mlhEpNFH2YUQ8WkG+OCiZoybaHZqsNmPEiFYwcvXckp2nF5
HWerkLigAQzlfx+iNqIIbPyFlYwxEsr964zHhUluFdRQj5GggHqCokn18+ag
pEtCNl+jn/+0+mUgis3pzMDlNMEQq2++43Eh7BB254KyAYdcD1TQFw8/HbI/
RCIsKtAIM0YmRspN2hHn/yXlyHR7qq156O+NTrekCzNoQN3dgqJFrNskK/eD
k5WYVJHPCDT8irsKV6tuyvYp+Rq/oPpR3Zuhg8ufLqPaB0xeQ6dOCPtXtVny
Z4kfXUgwIiIMB/LXwFzDkKLegl7zBXLThY1bkSWCwf6gJvSc2yvPpH6AKbaQ
7IKXehUOxHYHhdQlPIiQriqAaQl1oGoPnP828DlHs1v+XOni9G/zb3XDnpID
BBap67MtIzGfANjwGbXoWCU1S2NCSyrN02Ao7wqzstKCHFqTfLDCI7Ddn8er
bid7Rzfh3/B2L/Qk1vSRQd12ZJrarg1Y9dnTYkdrWHwc/USc8u2YvhasjhIS
NUfWVYgoapY6NzvKNokHhlT7pIwJD5zYzsMIzM1dapLYpeptGBW4TACFt53Q
h1AaYXlM1l8ewpGGg+koLYUVwO+4ZtyNjaAu035sdVDiNzQhgeYNK74+dIN5
o907i2nv6F1NyLoT7q9GEEG8VbQM/zrsKW+qWn6Cbcd9VHjyKCL7dIXF5BIX
Ld4MqdbNMp9NvPKOVx6CEeduqb1ARjGDK+uw6FE5fL8NCHA7ZcXsIwDud/Ce
S2Uh8zyM8aM1DMY6Yj1QWqIYg4sNyxZaHE/m8cMrny4orpwlnBk2xOIvSmMe
yc4MSPDG3VFGJnwdfCibYSGdDFR4pLbifj/6Nal6152Z52ISQGqbVDwF3uCV
XeiaBF7IsxFRddz04Ys2nCEA3BujfX7wPpMJs5hVDz7T0mgVPQ5hUieNX7Cd
5YyncxEX6fRyEo9S6sKtSEvVl5RvdSaqrI0iTr766m1Qzv80ooTPKLD0CD08
S3GRQkMvkUqTHAHo0xBvmj2iQRD2f4awgBkOmK9GaEB/aYBtHMZhE9j/AIiU
ms618i+Mc3vsItJ56MtU7GifOv3fLmpzXLscItzyN+kM28jJG9E0ZcpOeUyv
Xhj7cL+whEmr+u0MurP5ry/rWK8CpDcPcNcZMnvbPV6U2CbsyvpqVsMXZO3b
wjfxv7leWN4dt2psiEyqcGhGrbHFrDDv6Z/tFeusHBmrxzMHdN+GOzbgnKMC
Ipl3vikfkUmU/z0etaNWF5Yb7XABNkgncTiK5Hu6UBX5Uy9dhiUxpMMOIqrG
1QQx8OmJaQwfykX4BILjXKlz3ZvUmqtO1L2GVEzE/5FgEkqXslNg3OzGtcWe
Slf8rcs5oFxpCk5BR5LNviz4n4wtMR5cwnf3NgM0HiGPdj23vSMxEmBzbV3f
m9kEdmjv6o7gjqBkaPugLB+Zii8zWqdn1xgH2WN8erZCWY5FRM9vQEsKG5dN
6RSzOwG7RfX+hxpT/0YxxP5ai/BjnWkvcauJg4S1fXS6zXFsS6nvxl/mMxgK
RDLlvbV9V2CyPK4wKBl9FSQcduQLkOWdhQDTqd7KV+M3CSTLrZkvtBgl2jsR
rMgVqQ51kqr9kFz1LLzmlplliVRNPk4xJ3zpdArinnes1JImlQEPsx0TTafl
SE3X2vGEt6BTKgtVzTbTvEqEj2Aesb7iEjeApl3Dh+aog5+qn8w72XAielXE
Qj0f5FWwACOCbGsU3JIRiKpyzDptavi8arotvfX+Zo06lraZKKnT08zoyBTZ
Lwn+18wGoaGbQmVQt88eC6Nb8oMLl/345n3+uzr1H9p7lheKe9l4WyU3BPJe
lZ6pLhtAWwi/QncPgMew+f1mQx5Rtfs8a0eVdjfQXWYpPZKHeoKMMKoZFkvh
b0KoOk5XphOtSReUr/ePUwsvQdglszGUd2m9oAptTL43LoGby6HJ+KKsWbWA
0LPsOVE9iQWvG/5ej1Y77qGVXiRfbYKmQ+s8gUO46wCDLO/u9kOa/GhqwxPD
1jI+urScaSaci7HM5Gw5gBz/stX66EVFrgyE3lgSsAIohNORGdxBCktPIvcE
0JcpMYb466WIpnJD6k0A/X56+nCWWyefc0lQ01dJBM9gkm2yyQareg3pCVPN
obvKCi1Grx5Og4UNyI/rw4GxSaZsbCRjvhFa0w8aIQM8lMlvqGRRX8MBx93P
jCtdCVf0fMvTwPcVxFEcfkFCU0UA+E6r6YsaTrYR0BAZ5pmejBZcHuUrqgIA
8eIJn0xhRrDZuZB9cOgHoanuDBsMskX0rLPcugMozb6RWZtoYL2SS/x0KIk9
bO2RHwSN4TtI5bz5omuq8SPBzrChz1Pd8D3OUq2wLqvoMO8ohO7Fd3fAw3CH
2lP0oTKxDmcyhuoJ7lP0O6auPHNl+o5wlb8Fj+d0PEzw/bDhgahGlvPHCJ06
W2qXBuCf8mC1ASRDmAGsZSR8BU6XaC5XIMXohJXxZgWsHf2CRvy1Bd7xRQqP
U8LAAsa2kOdfZ3MUMJ+PpPA/LN4c+SAyV4OFbgLOzRyxe32x7LrL6mRcQsuw
E1kRO0VBFHuR40I//1cOmdaf4BG+g9n/18l3sPE4d5Qlf+AA6WIGPnXlIos5
+G+a3kvSIdqzxypXrA5OxHW7VqiJQa3ZikxGlzpabPOKAcsvQoyPPA8RE1c1
q1H6zTQ/1OmibCz9/+nsEjlqhZdJ1RXK7cYeXEat5w+eXTxNnAfR5tNtZtPx
QcbZOZRKpSa9ciw6kr2DQZEZzOuFNt2Rhkv/l3uzp0qlko97YMlCZfGrmQYC
AEz8nu0XXmOSzaiD6HyrgaW+m4SzXg1vaDbTV+o/vBREMvaZ6kjF+CQDKLDQ
PnWhsiNCfY6T/hdIZepPABkqaj02PYtygwGFj650lzFF8YWjF4ek7ngrXSAj
QHj1z5nX8TXovIZeKTtPhh8SytLZRqm2W43nsyT25/4+vR5UzRgozwKsVdyk
BpFoZIwuH6hwo0Ffl5e5jlbuEIAuwlezxiAHSKPmQ9b/U1iyb6HqRFa//9rp
oh89j1ZFjv8zJA9pBpSD1/aPFH0uAfZJrszYvfr27H5mb7CTE/SUz1paCHMf
J/Do38wgnr8PkhNRvk5ROv4TALyqVEsgFLAbkS9/4evVrhgB668wZm6rkqg6
jOrSWCAxqpNQGrLcQ8qVgQIlnD/17lvIAOqMKAeJXcNqGu4y5IOvkyrzyCsq
H0zugWJZ4QKLENJ4bb8Bi7sEan3NzyCqvOqlQPD/68SDWx29+mi1OEwdOqGf
dS4tcizUsQj+CnxeNdYumNgCKQ7MldxrbHo6EGivAEF7p+1PDoT5tajpsEkR
BEiYIikwFr1t2VvQ3o2UYm5MBIMhguTlcauCJ4HglB8nx7DwhIaUvVCpwRzD
9zFHGWNOSsdYa4LGhRx9sJ39OIoVRwEQp+YOWlVz+np+SvEl9y7f0HUgSIzv
Lg7fnQSetzkVypc6FtglnTH1AUZrvKhbryGI04A5YBbxbg/EPCxVPoIUBnad
HMuJrPdPUVC1kxzABqHn/cDFa8ko+keUMSMJ68GsNVbX7kTh74EJpfOPDtdZ
GHh3Oc7ie5XouXkonMcR+YUQiZyWoogzP0/bU9qZwfo07PNjg1w5Ty9eyqxv
oqu8WRtGWI/rjX3qGFUvYMBt0d0F1kiyXEvwQr90a3lRz+MZZqYoeP/8XRB8
XpEAY0cL7Jfo36PsyAuknWch1OAgCl+oe2dWcapDCFSLHHUG52iRePCEJCL7
kKRle7arJztEG/rxT4ksm5k//aCS4BQgsBLamEMMgNLfCiuS7Qo1qtQiL+z1
Xxg3Z3pAR8MFOpWyw1Sntq42AvfYWyVVKXxWfP0N16o+VzJ8khrFYiDz5xBs
IIfQ67D41uFX9Y4pdQcKSUFZcdHxlGYPsU3E3RDFDKj4mcQeJIS2PQorh9fR
Eu+B98qV8PAPSXfYOfwiySNhgs5CSt6OBmYwzKVTXQBpTY0nf42Q8zggIcCx
SLom3pdQvQCLY0js3qRKoMJL9ldqUDD7Q9qjV+C1yEAsAj6243vuiUz1lFQ9
3vKwEsy9C9XTZXc/isG5KElNaaTqFF8X0KCoTITPgo7ojg7FS/avgQLc3Bco
A3bWG/bfGWsFJj6p4i5/BINGTZPLbT2vKG6oiL6Hv9Dsv6rQtuYDV2RezADh
EIqPUxrQ53aYKEY/jBSZ14Pw5pl75VEg4cg7DURQBH8eqBHKg7hR3nlUt7IU
dBRh9E8VvdNsuZiqW9HCd5cSpWK1ESZpKnLmxx25qy0Yxro0M+0pMdTTBMzp
c+RUiJ8iumOceTUAgwGtA8l7sZszJ81UV2aPFxhhWkSlgIVHD2hE7lx/bvrs
9e3cpGOU7YAExNqR9lGnvPiHyn10LQFkEOPFo1a5SGNCOx/euM2fFDZxRggq
jEBKHdbpOsPjPGIuJbmyqDpsxBj9d09nraiSzvWQ06X31GqDrtH2Ip0aex5v
vqHb9L/49l57+5RXV6i/6Jm3180Qzr83UMNo19wd5r4KrTjlvUwiezt3oSv3
YKgwlG3xQI5Bl/aq+2PQYHSLmRDHeQF0dhzJEqhRJVwikS1jfiTGKhXeECzx
POqiTKweUA7p8wsed3hCVzt5xASuyrS7lr4dxljlY5gqW/FUfZ2T9GI3Zlei
WWEfppfaRuuHeYXHgbCIHioYYwWG5GaXVL+aK3iOpcdPIbXb2hq0YxJ6KXj5
FqSMpXPz5yeTP9Ku9uyTlgvWHrSpQT1itWvYiEqxfXcFYOghq9gJ8EJ+yotA
JKh+bZaXD4NDwIqs4rH0H1cQ+NLpfsS415Lrkd761y03UuLwo6tMvk1utm3Q
B/fvaQvkFsoyn5s/RJcoqzEv2c5gehZnip+1S9XHFuEr7ylhwvv/5iicto1h
OAu6zmBbKmPmbyBVYfckwjgxKmyp/LJPR3pZoFjy8T0ZPntwA+xSrcINJifH
gYdF+5KT6eg8vLkNfXAMi+e8xQvEYSihFzzFblRfelkQz//GB9kdT9li7uli
7IRS2cOMTOedlEF5pLw5W9oNJBiP2NcDi6LXRaBime6TIc3KVhzisdiL6RHV
1phb7bgr6xRFqfmjiNVZtKv1xO3OsEqR41CGwq/i+JYQ03BxumEIcghdB1wf
eauoyScXXTwedzEZZu89E6KeheY4plamha/B05yUscjR8nCdm0ZJT/Y52V8g
ssNkFPaDhECtVpoCBFaKqE6NEWsnUa8S1wOGTz8L/H9v6zfM0K08ArbTci9b
o8/5hUwuholMQe9gm/goUkU4tlUI45fUaaz+tSH4pnJ2YwZtlP0ygOWvMPp+
FhUNTeDgeedCA/g4KMNNFlPH9SJwG4L2wqVCrHw3USfGEB0qP4BnWLER+WvG
7h3tMsptyP5Ndn0pFiHs096Wut8SjgAbMc6a6yJ9bfu6NjDWscqV+Tg0HPVc
svYrxooqfe8cWyn5hoH81Lk9aKd8xQ+lEUzcNoSvy7fKpUq8ZmqW7OKfpfW7
HFG/48fAQdPMJvvJW3x7udaE3XdqwouQww6ZA0+jmaxwsc2U3TvUDeZRMaOz
Cj9d0faGvF/yEd9BqJ3at9VeoW7Q7lW94/UjGI2AP+z7lYOkf3yksW4bHV2t
oc8XOoOtNIwGKmZvL2GJnoxzwRAK3d0fVMRiiOUWtDNYOcUBOVjhYac/dTmA
Zc55ia27nR1QJezDnRE3q6EcRFFzsn7/i5NReO8f/907J4+fImVZvaRO43L0
ic0Cbl87J5y3b2zoXc5HoZYw+eXQcnmKdwPZaOsEiJU6ZgcsjyCRaAnbj9fy
Bfnimwn3PpGkmZU6+E1AJsXgGSSA0vhC0oFsiF38xwhXmEn/nQ9OngOZeVb6
ARp3GRofQ+jW2Oyx+WzmdYS7X04BpLE9QcLs+LuvmKAOmg67ajuYiZOLZjXn
40Z58GgoaJCNaMh9sVV7YzSChRTpiiq6eKUR47Q1fhKHVIAVxjHAmTYBkbUj
vVdCPao6EXeqlUtAa+CyvmDaYGUUYtiOoTjGZfSVLRIWf050KRFEK61T8d8r
st0TlTuxmeF+Xg8nJ9FN8RwWcrHc6sWQFxgC3lFLxPMaILtGwtJ30kcom82l
TY49izgiYa7g5rzYrCiYcZ6BOnjVlJN5CidQwnTYXmVI0/V5YmckuA0v21Ei
JOq4BqK5pNhsFyBWMnF1XlAFK1PhBntf/bpNy0x4YtOD+A8clZucV5AOhhs8
8s6oTa6xl8MGQIxs26fkU57fHOSjLFzlKTy8HZDEOsa0puLFglpdUQnAM2yg
IVbT55ZeWsKrDPezq+sx7MKEW42wBmtCWVHv/d3wNNY18h4inxscEDInSMb/
JBJh+/jsGQoSwddl1ADGpjM0bl5fb5EDqhxqBccdviTZQzg4UADLLw4/D0Yj
9L5ToI4FiGkJaGd0k9aBnh6T7X4U8Kw8uPIwAVVaMe1WuZRO+I7TSy9rkudB
leCXm0WN59IR1UMbr5dYeHDNLr4cZ74bcKUK8YOQOF5CHewGbDkLv5onvMy6
la0dK1XrfS1tT+jHiiFTAcmZOPAeM0pnCKi7n63EOV2sT43YMN4Gz/tUHO0N
nG4cZX/mtCMsaMvEvJ6s3wYAxs4dGlwV4bKGbD9kRmu/DeZka7ZiYKZKaYh2
IApcTK/3s34ANst00K94Xkmt58310pT/VowiC3aWtwDOfo3z1LRYCo1ZCAsv
k4TjSgNMdEd2bHJ2COXj7x58VuNE4sbLEfYgn8kbnfcycf/Id4+tVpBpIAyw
76Y/3L3DqAH3aV4S7G8HfSGhhQQgApuvtyHjtlG1rnxd9BK6oOH8L/bVCI65
e4J73ZQ+R4PuKwRx3U//7aYc168ZpJ4N+Pwe4NiXKzSxUntsJdhu/pywkWQT
TbNZ0et+kzx7pYvOfWvOsy/DQxpZnYp3i/P0z7Em1Ub9DU7bHvtHZB2NmjQA
w36X+x+b+hGd7wt9jaTo8KrQTcMlOi6/LzCjHrd/U3g9KzPe/vfdsGA0SKPY
A/27xKzxW75sfJNP19a5SphRByb4j+30yAMNIvGT2VYhnrjcYtuRoMpNnwB1
ZuokyawG1VKYF0m9c1zxMnqy5ZtuEojEzjFH+7zurmd9v5BR26puDsVXysd2
RaR9+G+gxi0WmmPwmBL2UpWUfPIsPFa8X60EgkvMbRz6ApntlfGS6EkKCf4M
0TrzdRAqG7LvtS+0t6PuVc4vqjHeNmvvRKDH6sg6WXCcTc2ik4oxmDOcLird
wzcX3H2RKhK02pldgkYG9CUfEtRDQjQdML043CE3ZgPS1G89wE04bza9TmgI
OFGChnlQ31+jSzgz0I74W4fL6sqaeDPjcUV1P/6lTvZoIJro9gE+q8BOd8mT
+4TMYtfY26f1f1oe7M14lzXzXpG62045tWgBukEWdFb/bOEquqanq3uIVAHh
JIKkPPxi0TdFcjcJiOGOhDLrbQpHW7f9z5V7Ci1j7X7zjWgfBHG3R83rKH+w
GanzIskQTcq6Ex4Dnvoq3AvtIKAdPJPDIozMLINUhsY4TZuFxCD9mX9zVi8c
fbtcGXTgbH+4tFjCDIDnZy7GpceGkqf3rZD6NsNuz53SxZPRBR0Bk0FKFMBb
/WTq7g18LpzaSYcJpkIoixnbPA7zw0RbEHlBexxM3EDhq3T5cNyv1pYvCQdK
PLEVJN7UAW4M48Dc167MPMV2ullLm0cd73xSNiAWJcJ0NmjiF1aUBlZkCja4
VzYlaK0KUAHzaDcQiiV5HgOjz+aY9kbor+GqUn15bdbQPqEK8flSZKeIVCU4
rXPjfgplvZmoY5lg5XU38BDriDc+I4+GH+mEoYykOJLub1VQn0TElS27VWGU
xjezUVNptJp0rbhPTMFG6Kfl01I38jg2N3jD+Zfn3HLrb7oNUYhybMBm693i
wSsmNaQLwH1ScfPUo7iSxm2VQgHH7i7DFfOf9jP0rshxWj5Fm4b4V499nZym
0JdUlWdBYDTmpiYc7DgjDMjoDju6AqlxEoP4Bh2ACDGeUL5iIVYqDFo/DQ0H
uhYYT4u2RLx+dbnTZ5N5j8C6pWLlotAbX+SMxRr8kPjtHH7AOBg2Pk4saEfi
rw3GMBkGi4mveZcyIauCYXx9F/5YkGMRTOwm7gj9wKnjZX4Nh/QlvQqhrz6C
ioILpBGaiSb20il0J+vw4j3WPmm16sn/SClOx2Key2uqp/L5x3aM6MEvXoDY
XuChR0uFrHugRcKHvvZiD8zgvNuDsfbsWuJUpcQBXTIX6lpvrA88b4saJfPS
MyVRnIf0ZYfzB1ki057aIKagSokVUujAOcrCQn2TCd7IvL4OVaLkkWqNY/Dk
H1veL4CaMDZg5RY9344/Rj4QiERVEf1tEzOSIYgsEOfL+uG3vm+Gg5VPU7D0
a45ypchXWsDjcrJPJp9VJruhzmUzR23Nv88MqYzZZrnXTg+NgbxqR93ilFGa
SsDIUjUhZTQt8MB85Gaej0UCvNOBerllaPY+D9bAcafYMYERr+eEp9gJk5My
mf3fzEayJlzL5c0+cVpGc1q6nxN9YWHumI4h6zpRPu20g/0jTDldUxq+uy28
zpsGscjzwRxguM7R/11VPQ5Gl6li303MOAnGRdfhEBKF2aYfa0iYVgsnWu1w
0NkIEXyWllupPERQQ3qLemx5eCRB/exKBEmLNGc43d1OZQ5eq9VFlJFePa9Y
SRVGm6GbbydCTvatDIllr5LAXp21z91WpA1M7uwqc9sko9M/c8Ik5KZT2MWr
HnpB0M39Pg2fFGXg0AP1SPvWqtzxfH5heE+F4nkFyWwscNPZSKgY38HOWPXe
7SHbosdkSoFWt8ROwUr9xrNYYYJrfhZdCOav78w5r0KoPrKwO6tGjJcWjboI
AN5i+o4LI7JgSVhhog+dkifLw0oe7BDJazKF+3Ra/KHVX3DGVqKv5K+lNZps
jf5XSuf04lTQrlxAUcIm3DZTarZy2i/1JN6v4vAWITvypupJL5ddWRHnX2Qo
JMwzdotqTbaxSFjCps8zQREJ1hv6T50feoh1Gz+ZMonuOyEMMkG4l46FfL0o
JIZM1cVpI4ouYZeHfW0gcMMubpOe4aymBK0PpddFzrN+MmYtykBw3yPUIk5t
tWwpX/xEGUEumB2s0hqY8j3Qq+Ryivf5m+61CNCnO1ayhMc/FP0xwcYqCT06
7yVDBm7ezCrZ4bnYCt9SHw7JefGtxAQ6BJprY1/VDbJmnJeuwHjX0nwPJrdo
AVmJ24e1+qWEfUWiTX7/ui9kfV/ZZzeBFWVxd36V6Eu7oM7IzxyUzsK8Ho1U
pVZyWj98CsMG/ifNQvVB2jjlmxSR9LIAvOw+JWHqBAJQLvVcFFmCT+NiYNEb
7sBBfdjvpRx4Y49tlMAXbG0+RLaHaFK4cZ403fbOEpokbdPSSbw8za44vCz+
ZfhcH6OgNNaiPMsWIOhm2oWIoF/l/dGZHfKzbfgu2UUHPvUmV1ksHD8/R/as
HujOPNTQVaz4CUR3XrdGmYK8aqw3we1krapNguVZbvas7hIbE++TbwEzmyNe
B/PODH7V/0tn9L/H23VW0e6362fSCXGTChgPJpjRdbnZhMrqb8Y3Wqgz1Jsm
VW+8NuumbxW9a95wKcxkCpnlDnMiLAVd/QMFDuDEBvbhh+rXlSCouJs8ghZN
HG1idt5vMNnrJLodeT2q2kgO8Ov3gkWTV3WJWADIYft4N3dpM4nQh/71Azed
r/ruMjNu6A9BMmioL1o/QODbLhUBx911lAGQuLuxOrsG2lALyIaL6Iq3JevZ
j6Lu7XahT9wdHo9jfAqVACt1n1MSZDnLUkOHrf6EBEIaO41i4XG2rshwF02/
Sq20BwQY1+OgmoHWPwC7TjWQ49xLYSdRhlHwpdmbuZyH3RraUcbNvJoF7cpS
4eXchvcu4WKxBKVd0UIHOVgXKM5XIgB6nBZ9O+230IcaQfqteI4oZrjv8aWs
ndDaK+9BbNakxV0eVZlWedMM8CLp4ebOl9n9F/e4P5981vtos2i99ygUajOq
wkpmYXOp/mq01igLesct+q+ZOYCTTmOXFwKOASk1KlSewGdkwIy2YlRo5vXs
dISahQg9TGpN36FlcpXB21dQ2pkt8C261yaSqVyOutHYNHpORKH1pSlELmDb
ePU+2K9ArzGWxqRplVCg+RQCDXWj0tIV5/OSMSgvuuSSviNCtfa+7kGKHlsX
BBA5JPgpMUucQiqaxKSdrqTycTvccx5QmfbGsUf9COXH3sWd4qsqGdORZdM8
XO4TuYhNWYj8VBbim6d1k++4xYd6Sn0IKx6RZJNnewW1KuJTqqNMAD0NkPrh
15a0ltr/f7F0StVhEhhER0DiZoLzkgIUlHMJm7wLPpUHZaCnVG1HLIBiRbjX
aFZ6atFrdtQuy6KfCzugLIAsoF/q7MYYwyTtroYugPYzj3JyCNu3ZMf703s6
/L7hKgNQyZBbOC/g1f6uWbyYwQyNfnzKK0lMmcD98QSw5wmTThkxLSytTVsc
x8Oiq7/907wbduwcKMce3oIZ1XxNFeRl+6ZQ7DLhAwqtyKFiFBqcmXWV2hsP
xlcr+uT3DF1Epbn7uBxioL3/1IsfYRRFm7Knx0aZwMnZBVhfD49AeBNhwtV5
UkDJhX7v1zGqkkGYFlvanXonwmCq8t/+kCOkJk2xvIX/v3mgyFWS20evgjrD
9yMHCNwSLqH/3odNimjsJOQE+GI/qFpvgcicgPsnc4DUqKpJCvBMfj65+ABp
WhD5gV7hitPxUdS0AoH9UAIa/NYma8+wjrn67t1OmQQFxXLjE6RtiGS92w4f
MhuvBvPfZ0/YYPz48EGc4qBhBL6fXrVgcXFsefor9zkiCjnky1lEN+FmtmZX
mJoHEKSgHeUB3Bct8l3PGH2OHrX9Sr3/N6t2OHe8cRyhPOUs6p9TDr4Rt7Dn
QnBfN4e7NyshWB/OjsjdkN6rSFpEqQvmxTqJYQWC0CzYAZ0aH1Bj4TBkcrKM
Ib9Aj/jTZRg+PmVlDUd/i7OF6mePbg2dnSrQWJOJRkecLXYVd4CWj04fsfRR
Hl3g6LJGlksMHi7z7UnXHKq7rjQDpWexOBhRKXcddGHXIPzqB2k+s8vzhMxw
HzX4wqofT73wJ6MsBYLPFCyLlrcxcPHTbQcTvIm5sKuczI6Vs9RlynSyz12X
sNTLmvoyF1Iy9iyXruqu2TG34c8+/8006uw/PmFCILDBMWQ0ce6wZqhNonTp
KIP0RzzeU0aIb9rUcVBVin1oVu6NuZ96GVy+eNJU6Npmv4gHyiFiHFmS+vRa
l6zysYMhCL4dWJLK3xNkVoee+6cWLKoK52xoCvzfFyeV7YmNIy43RtHDxtf8
fLIBk8swrkwhP2p9shNpSm/OsBprQkfXBJcFKQy7slIFd4ydJEVT7G8fWZAh
wLAGn3AqxJlrKyNH+6lh0IPH4HOJY9nSJIHCzqwpkdbUrnU7QfspHoI49nSe
LH609rwz2itX91vsR8PwBJQ8cPziCj+AX1mRTrnDydVkBfHEX+ISffdnTAqm
BvXsSwQfC0bqutc+JL6lMRDWPQjSaPgCK4ZoLMjWFdYeKBNw70s2gkGvJU4U
6cvwy6dAFvbyFY6wDNF2MvAgY1O9Y0yL5gQ5qXxhTpwhLUUyXrUEVNzt98lX
Vh+NVHFcYkLaLIPI2eXtTur9FWN8Imztz88KeQSEzLRL6O7M9enhEGn1oScm
4x99lulMAO72Keg76mOhvep9cA+y0cC6LkXCQxoe2C1fvdunR7VMtaOUGzMQ
1qpu3TRID8zaoukfU2uFgkNG9YVRbrLp3yN4BX8DvQ7ZG+qH9ejFhOzhTNzr
oAJKb3tnAnKRTVZUz/wG00V+6ODWytmODTVW0f20rIzTs+ypgAXOGpZZPrFg
gp/cm4mZduV+OhknzcPz6+aCqXZlZlHywKMIvPEimYDm6HBOqsf+c5P5Ns8k
vzFdcamDXgr+OlcUoQOEViFBEBjs6ipxQC4R2QlRWyt2pu9CpdHwcT7jj6zK
GnoUPL9CkX7oMx2AbMOUf54n3Mq4usNAtUYlBqPxwlXVpdCspthLYz0km/0r
lPlksxhMR9hzjtRlqRuXo4TN9FroYfl0GrwXCuShA2DlihvKPZxzvcNYdreF
OtSZ2MIkOet7+76Df/jkH9Cc+vmCoVxzlGkTVrsJZHlFnu4pcFoBkULQtK04
sb3fhOPTA7ewmRg79USIYv4Ch/GhNiEffjWotSjABFFygOgOc3X0QO9/RLLc
c0F7bGzk9uKkGf/RHbLqhwo0IE7YjfkkUdVA0PYWkrZg8RWmvGt4liuyt9Ar
8T4J7iW8MQW3SPdkEKAORWjKhuaxkcoP/IsGX8TxIBkx8HTV8zAfo5nlP3jQ
G+TR7/2it+ZK532Ayy2Kpci6LAXkiz9q8hXQ0xTeVg8a+TBETU1tFatO3wWN
6utFXATxavByjJdIM4Zgq0EEHGmA/3Z0zV0KC96glRvKYR6vQmrnUHcZujSn
4a9EKVIklFV4jcDqD8y9ZCJssiA1gSGf1zZwUtlZRoDYsTLqLMhB9pZtGz3G
69G3922LltiZrVfU+qtbaIrCVKe58fWxrsiBj4+chwhZEeFl5OEciB9nJ/2+
4cxkpx6SEj9Xn4uVOSyE6MLbq0+Ah58UalJc9lQOSM1gW3MEH8BnpeOFH5hn
lA0Lt0hgB1zcphcXWsQATrC1lZkx8LsqUli7GVUCF1nXrSzWVYgree5BUPD+
Cv+To0d0I/jmFJ2gfji36jV42MlkiHlV5gt/7DtFv+6EyJKRrucccefbwa9i
G2PzchAVnjsxt6NahBwm9mb2xrknxQKGWHunjKhJDx6A+YzHvJOa5RXJcrcr
pES6YHtjHrWwuiDE9eMm9STc67Ks9puKi1FWfENlgGA0IxKNsfuZdaQ4ES/z
hrlTanf1AqQIQGASWLRjuI6yCJQ/bTCfojbeY7DKHpVj4sgt5jp0tGjnkiO+
ZJMULcbhc1aU0Dsif2I5FNwIvStblNioE7getGLxjsA77nj20HkA9890sqEh
ULCSM1CxDkyHT1o/gP8xTzncl+/IEwgeIbvdDwyn+K9nHik01Ohw7qafWdcs
OXxGnXjZPnSb0crc3Q14cCREQFbMvy7n5lS+XO8W9dm4Nn5qFkJKMgsypIXz
tglWJWHkR8nshsrk6gZyXnpY31ZzNoBabyuKmBzOjUJJBNUVyNXPnyi/S9ov
et6Rn2bcC165MMx6R+VjGpp/Ksm2V3F1N5zW9wR/LGmGgPzeS113aBKZHvjW
gUg1tiEusSD//TRgUqThM7wKtNn3CQWeDzIs1gspbxIBAmeWpW5wqUGEsn4U
taZEnR69qEefvgLK1/PlZPqbxdws9JEOFi5ykXH48JqQyubIV0r84IfivYJk
8X41kOM9JYkZennF9Xkg2W/KYc4naU8gzYvjH5eyRgXKQVoX/uxeTlgaDcC5
ssqdUNj2KyQtSQikxKSik2eBltGST7qQU6YcVxbNNDQO6I2eEckBxLT4vHqX
KpE3ZwZQrIRbI9c7DfzN5vSChHZ0DzbHx8UzOgamwMzjFuKT2hPFgP3Kmxxm
KMYOG+0uX6rxpBzAPG0LiV6kBSGreNgVKqZH+32+wjcnRbKppIvvILX0iApB
m0DBAxZaw9eR+f9EaSkL868JqTTd/22UeQikWm+hgBPoi0gSyIL7UzKeHbGY
mFeqdZyRlJnqDWGA8oXz+Jm7Qz+kBx3CMSQa5YUX9wlj+dscebXQxE51+H1A
lXoLkh4yd0XHNF9D9j7hXdjbUl0o7W8sT1Wr0oYRrEhHq4dpTCyRNSHIKCDV
wWjc+Q==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpejT56zjD3A6hVKff1bPy26HM/5KeAQCBOlCWZZCmZ4wO9ieormW/PwwBsDYarZpFhBsqfvDl0sv0Gnf/26M2Hlawhdxr7liAPXXxgH8qNS+U4AZmtPfnhEAMuHNwtAMhOmjKIEI8JqFzJOmPQMApKJLO/+GdnvUvxu5j52RBR92b7FJU4qfkR3Otu9DZaaZDVs0vSCctzSLTOGLKeXx/gITIJjJM8Omj9yDjcOowiLP7MTi+3sHEex7JLpX4MyJqU+dPDYsgNgy9P1MXIwaEWMot8kVuA8WQtL7LxACc3okelKMheA6RsiIqf6gs2uYBIm0a8ybeHehBz0kqLZibyNK50KUDRl49I1VX9Zy1lxHP3wFZZuqRcsMLuz7M7vcQCUz3WZNi+BHp5JwdojtwwZ0COHdCjVQ59eRko/0ULA79NcnxEJ+Yfc+KPf5dVwCN0GAFTgEI7//L/Ra1G4zDRyEaaQN4EnyfgmO9xhsj7q0rpXNEk0v2M5LX7ETS1PQjsnXZC0e870nBtL2fwOH7l1yo5TiS7e66ullaOXWX+AwMU1IKF8Lnt8HZ+dS7JihmLkGMVermJ5HjSEzjO7bkNZyo95X69q0Tk0gKN1iMJLwSr2pz0EPXrluETb70NC2PkNYOXiUqTgTsoZM+E2MTfmvDX4oN5NSCzYZm1I3PdXvVLvXNT0dKd0wd1+jHVme+t0rmeJy6N4b+BYnkkDnlgM91WwFcW6NzJkh5IcTG26NO1ABXVFD+4SW4OEwJl8JBylF/Ibk0B663ZIO+8xgtQY3"
`endif