// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QGsogdmTJtwzRgkd0mliKTo7KkF3KpGYEOYZJ+ByOZd1LXCzsQ/ihjC/RbIp
n3F0Ez9P1WefAVbFt8l2iDTNNYx3sqCCWXrZlPm0wG0cO3Xud7doNE7Gz5VJ
eVGfI3GPMDhxBIHfad/EZRMHC8ceaqOtVwwSDbsRKPlwsBsJXg9KLXN4OrqK
JVBtjyMu+cjeYUHsF/clqMSBQgC1ch8xSbw8Tay0gcRuS3NULwte+zF2KMw8
9VbIalkXnkTaLJEh5uza1KxmHl2LIx5V5ILV4pqL4ELa8R9nP2tNl7/Uavjh
kwzbDo4rL95jdCt583oINPkOvWoyCwZYzqN+7BTADQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
omH4nkEWvmJQY0phtj5Z3Opz/RC2y1yHeRCaLdScPmP5AW8NzwVJwc2YftZo
TQ8rUxVTbsBLAWCEvPHvODLCNbEG2TGOWvlm5pUnUf47wV3aKAh0Nhwmuw7t
I9GE+oYnPJz/Wej2QmhhZ6qq9898Humig1f23RmIqnjY9cKdvb86rDyX1HkI
uLhqOnVfNECZsP4Dx8cz+BjcABtpbUiyK0EnSwEph9YgAkj0IoPeoV4X2Fa0
fvSBkOf+twvw+h86G5GoizJJf4+lqwvmFfynlS3FQoq153onHzIc0PCVQScC
ZZOLzH7NdAJC0Eyy7Hh7vdNTqriw2OLK2SiQI6eatw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UuhoxiJW+0e62RVzhhQNnFMqoOMJYzXd8WMTWAHgc/EJmYwFe1dagzo8dcHZ
Va1F0zqxKjsQcnWN5P/GAFD9iOqPKBf6dc3ti2Gcw20gisiLtg8f15t6t/ld
t4FmC7mvgTEfP+wDkxVV5WThHvI9hIziQfwyudta2wIELaO9iCVxSnAvTddN
DTRo0cbXz4V3GU79tvMbJkJvZPzlL9qgQpvnrlFTsZV7tMlr5bDknsRarSRZ
wniOytlYhxbh0G9fEYbAJ9WaPq2GskBhyHc4iRb1kP6NflrMJxqpr4DY9UBT
0g6gi6UqPuYpKZHWNa9+kh3Ao9R+LapJI9PzLf0a9w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ldZKGxrB22p6Qxh7IYzNkwCG55Q1Tz+520dxXnHGw44PAA0/JLfMSmgTzisT
3eGNeoMElB8v5TzZObxO1CkFx+UZ2L6i/4a5vSRvR2wEyGpsbhjFp8caR8WZ
e60VJpgEWPK0TCde5/U5HQxCGo7VFtlDffrA40dI/RWGFKR0ViiwE3K1laeq
g1qRCvHphskYSW29nvqc7wEi1kUX2F+xlH/BfCgniuPl50NLCDBXXy25zfLp
qVVyXUzlZG8dj/Yq5NjrKSkNw9Ot2M5zLwaBh2UgsvTTGa2+SN9b7oEU5pv/
bJae5Ki0TG4jIYMfKem4a2YqW/NizBHWUMoSQUAvyw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
enHgoj7TWk/ak2yGrKEQdfrtvJyplkYVdae86wB6xnj2xj87pg+jL4IZt67N
8I6O6N2aeDb5dsPKKbFE4vhOKUyjRJDRqFksECsP0SCGRLstMsU7nc92vvlF
MzUByhk7htMxiYeKTYAfyNVYgyd8qcpc2m/q/m/k4yLGYQvz4iw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oiOmu0a6Z9qjXSyq8zhux1POYa0ccz0jCI5cMNdTOVvCxG3dWDsJ4sT9wSx+
1JOqndr6vZcqXM+wH2kPd5/RKdKBnaFczAjeC/nt/WlrG5Qz1piFL0O+zzWO
wgVXOwJpX96UpgrSQWUAf+8nwsUop2JE91hr1qxK1+btBc3uos6pTrSWut5i
PDBQIhqZoj3U7nNdlteyUcNFGfN4nrQ7Es/g+2SUKd+ZfwASt16kCNCerI6J
gLerl3D300zRsyT/z7imMumw/MlVoglSjBzEAdH3HLLhpSZW63dklwwfYUoj
jl1OtAyAvKBHrMXkvVmVTpiObmktORdYoAh2GbpM+GJrvpiTP1z/AYOKXunv
/Md+vpbwxQcf1L35OHFCSFXIr+hYiGE0zupVOPXZ1wCfHBeXcfQvt+l3yRHq
duM64GvHrBFpN7lvmssPuyZTnqwcGAnabs0QD3IAUYYJaDihdS40hLHIsvdT
4fFD89F6hcLaovDfmmUY4jhjHSbLlT9T


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
k4scJpuYQcVo35Y/Tz+kUwiAny40qOfibpXlmNKjQgsIGvl/g5mJ5jNCqqOW
lME5DnYu2kc5K7nzdgWUs6BQVBLrMBw6i4bmeJwfxTr+wQ7eqAX4g64tQB/E
3+Cy281EOGxEnOxl/ug9kp74die7fecoz34nUTH0RmBYDkIfveg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
c2G+eq1NQYxGFQ/tgYQDiAKzkKA898bCbuqpI7p04Wj7RwikXtAGi5P9E1gS
BS/5H7NL0XlxKr1mwCXtYM4qJbnhh9XyJ0Hi2uWQAJAdOSCy1ITHhekvKTPv
+t06xr+tcHe955XhznulN+9lREIvaFPofpslrPwDy5zRyYeGT+A=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2160)
`pragma protect data_block
Ne6FP0PJ/YBO/bnr8lO7y2oa2M/UvEfTTYAZV5OjFMmuy0Y8hBZQWv/ThGSL
N6kwUqPdKbnTnp7MvPRQrOQ9aTgQuPnKGIk4qeBV7p0GYTj2JquLW6zH3jx4
lcNPYOZfnCmqYctPPfNo9o0Bog9RD26Hcmm34Nd4wNigoED6bKy6XWM9fiVW
qWQqBR95MiA7aVc1yyi+kWWhSfB6lDisQrnEoMgQXqSKXQywLr9OjdM2P1bL
gHibg2NiVPro2omCl11NC5tA69Gj6nkYO3Ersaix3l5/zv73isyMStHjkJyQ
YKLdo7krveQt7dNpk6oRRVALe96hr/W7aT1OAiFcBmuJIb1wmUQHw8nmmSN7
t7WAyAqT0NDY1id5U2Y4XL6tJgDer3SBq3aBOs7/1HSJ9Hl5HW7KePY4PJBN
c1tADxCLp+iqpixPR1efuEJ9Vcuxg6Ryl4jd6ihvdkaLoxTX8dkZZM1++j8M
RAshutnzxFxAg7iRtTRNOppg/9UKE11XgIBd6i+oRcbABYqFobtICBTa3y2H
DB9I94eLUWhvPU2XP3kewFUwskILZipRRNrvIYYFPO8aXdd7LccibQGW6XY5
qDGRYX3FeGusnqGSQPfuEMzhVmrTHAMT6QA9CsZV64GR161rsZcTMG8jumTY
aiq23nla0hYKPC0E5gNOH34DnV4JtXdZRFgCU9vrOr8pEVZpFLlVaUx00cWX
CiAaYweSaJYvS6KS75zLU5+5Mqb1orbUirkIkUJWhUpT/xu9eMWO+gSmg7pG
T/pMUCsS9Iz4nnnaMekzBY7HWbEJX+k21gIE9yW0b89qNWknCXkMZMCTUzWc
kpgOflNEXozdey+2gbwbeBH2Erh1qL/eEEn4fK/QNWENMSQi6ky4SLY68RBG
xr4T1q51mC7yf0w6lWtFERi06wT1HCtRU0rSN159PGuh8DdYOcXf9NSQPb7O
nA2fq6pyZ6xQFOAzNb1w7sCtziX0A+N7rM1mDbvxa/hn2uc4n3eA2lVu1emw
Y403WCt+pHwyrXCfGmT61g+0/iW90VIVOlhRED6O8Xxz7afwFV1m1NSPrdFC
75rPrYFpBoEFVIOZeTSc9N7Bp3BL7zKduabJrjWdek/52YXfXP5oOyLzdaER
kV8gJQc9XCB1Vvmq3hC8GaLrVbCQYAdZXEpytwwg9jnd6bf+hL+3nHJKY2c0
/QtXG3I2zntxbVIwm3f8Cz6CKiv6SS714uRW+A3ezFOB7wt15YK+C2xCHEne
ZJH6xtWsb919rkVU4mUPMZg3MOq7wNH7ph2DmAAwa+AnjQCPCTyy+seZa+Vz
bYlnV9MgF7IdtrIwIVWIMgdqoiXLd7LsVplILYDYSLJPY0yANjccSHFMzsCe
8w8xA1Q8dQbmtyDQz3XjzBhiOJgGEbMSWCuU+iWYGEOFipM/vMC3KsiASi73
WuN1ocCGHNtAb1XxKkmocsipssGTSxhWsEob6Ab8xrDtD6Ga+24D2GLLtSCN
MscbusgBnLa8uXMuabOKdSj67B2Z3LZlhyA4j96mie+8EydgXlOKVFiuqZsD
qWhilnyAcFoPYwYGzJzMih+ShsW0YIvRwNgK3CJz2yl5Ag3fPMTHbFccT/LH
8EJVWUlZyatjBJ4RCG8g1bvR4FWugjfs34EKnFhdSCRg+9Rc2Cw3KcG4nrxZ
5lO8sxAypfz1zVfq4o79QpL7ZEwGsO1YkEh53xt1Wi7lL+kFl3I2QWW5agYp
Re7lmnzpcNO9jP/SYBC7oB7nTxNHkB5lX6J6FxNVYOQ4ZZpr+UsAzv1Q0buv
XL6yxAqeJIB1lNUhK4hoGJjKeO3evcIYIRzz56sLom3+/btlgK4WN+Vqyw4Q
9lmFGj/me9xtGNDe4Pvn+SeC6DGTrQIculGulEau36w4lft5xefVdMI8Vm6c
Hon8FnEx6b1kWUoIS16v+pWwy1yb6OnzHber3jtR8cYF2zKlEMFUbbr8KQcP
vujiPabnP/dq57hCHINBpd/2O6qdlqOev3cc1oRUwa4DeqM5uO0n7dQbQCEt
TG1BGkPXJbj/F8r0fNj7TR8Rkv6rLcwa9ipa6isIqNn0Sgj7SMqMxi5Z49b3
41Dgsct2Vanu28qf04HIrw2E429EaObLdw3q7gCM9sx+pI7JpDjQ3MXN+/iC
Joqhqtl8DD5l5f8iVkLZ4rd07JN/Vy+SxACMX0Z3dCX+h/ptjLTnfYO9EJq1
TrXESR4ChSKOADBoieDYw9/cvq9kxuTX8qwXyTN/Sza1WyYIG/sluKzLYVeY
PbeOguaE0nu8NQryB5ZoALixhFKOmMkCr4VtsqlJ8yc9BRxJ+d9VXcWooXK4
DQDNYdZZXGbnRtpQM9xuv2B/M07PMn5iCTD0zMYKAWDojAp8iPXG61ENqR+V
5hEQbfg7zVou88sDkuQFvfgQP0GR+/pM36bDzb6BmH38Fa404bm4TVF39S4l
1mrrZeu3oPMrSXpO+XzGbA4wSBfGY3d6QGWUhxd+0/1dhgwccgikDTdFEaOk
fwgYLuM2KEUXKLjcnKJYMBLhpvSkNMdC7H4Pb6jhMHpWDw/8LMg2zpeJmZ02
5Oug/q3+VSEl4jfs4+Uchsec3DbTBVKTw0qPBAhTHKYy+TgycPQ3oowcqIB9
ZIkSRK9l3LU6/UvWfkMpW77rh9+voa7QRaKEgNc7h+qfmm7qSA9srjbRKCiX
z17HNr74lZIWONlw3v5oFMA2TERgsq35hb9PyOazBMUScZO3axWZ0I09zp9r
0X1K9qQOILhoXj3dD7zlPQCKKYQwCJe7a+o2P/2p4U1316BRm9nKTPKyqhTo
12UGzr61UaZ7InNMMK+KGX3oaH2NhrTMoPUs1Gu5aA8B6qaZIX4Ofg2JIQc3

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzfWBu8kX7YX3pdMmY9YumhpnGIwH3JRWXgCvayJq4y7w07IAsCSW6bCsDNdpoYJb1yx0FPd+55vNNG03J06kQ23LMc9ydVWYfGgdhEg2nE1FZ7uS8puqWL5tzbAIx52SEJZxVt4ymtgHeS1byQE0NuM98itjVmXR5tDeRgOFHnHzSmvQqKOTfvXGKHeyVWhGMiiOx1oeGe/a0LAth2C5MpyItF/w9v+NtkZD3EPWoyuvH+oBl+1CmRpHiYoaVNznEmSnQ+zJ/Y3+x6X0DiCl/ZnCjZhq8BRjXR7ZMof1QM5QyG6zEdxh2pRhkEhJjrkBe2j6QkAfeIrs1pH//8EAJLcvuIe0xpdbIx5Ffm9/Ez9ONO7sCOZT2rc1VTrJkVQkI3BvOz57PTKe8q6uJsmLREbKCc4lQaJaERt3VAbRzIqN7OHV5s4cAr1Ez2w0R7m7GvX+KUp9ouGWCAEtTK+fL4lAjOBIO4CFT4jAsNCrX/yjtQCkEhpgMCH2Qy8T23vMeU9zwLq/MJTsWu+fcO3J3C1tWOf//u1dQvWPAKAVMaC7NCsEUpv14n1IIfoi0JzmD4dLp1b8RrKbqvHcWHATC/EOIv+ilCLUItqZcPBjONc+dhid/4hf6zg3IXwTzesXadKSZpEyUbz44fRsTYT3cVCjme3eHYRGzqEBy4vXLqfgvWLiN2AujpYkj+i8aa2tiatxC3bNFm0KaDVuV2CSy3JM2UQoZp8Fn9fVgf8sMV3kYzyjQ+A9oHGKMMAYFB8uxZzVYmRJL6rT4t253H6Bb0N"
`endif