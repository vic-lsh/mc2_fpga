// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
02ehyIccMCYvenEpEASo+6A1zbvBmFjxishBllRkWzaxdyi4APTgeRlzyeBP
ZRjDsRifU4HI6VpadHwNMpbYAIAjzurpOuNUfTMe5rDOfDOLp05nM0u8Shzs
nWQ0UCMbmGkX+MmUwI6GmFS3RRU9KS9RBKm0bu+em4HGy4ruSG9W4JLrL59O
q5OGXr6kP/rh/JnJuiRX/S/ltoegI/tLGimCXBVcpB4N9GlaHrS2yiFrl4/R
QnNwj6+vhE6vViDAAXbuAT4LUhlzZe5M1TEO9/3lqGXt2VpNEvdGCtEVJn/9
178DG8EOY3+HpoEb64tK7D+y6zeCSn6aYXXWHlhN7g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NG9i3w0HoLNqqIKKVYCbzkF96AJQGDiQbv3A48z0TXz5T/6YXgUqER+Jno29
LYAK3jh7HoXDtY6cizSXf2lV5Plytdt5n1ZoecJK2gA0ZIuFHFgP0PYqt5FG
RBIE7y5TNuRzgTK/NNj+2LVgx4DnlfGhwbaUnpQQuoiKMwwBx29Tg/WvD/0R
BraoOUlk/9fO6xV1Dlg7N43Qy8FZp0JlfC/PpMRDJm9HVH4YLUzIuJ4GElXa
s6y3tUfY+xNHt89Dh5/PPEy+hNU7UxNvRFqhjDyzxLEW8bNqfLRqxOkUeadZ
sVxYCcWCcDEV6L36HvJcPkbgNHquuZxyIqyjDoyOlg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EO6WqqrSdZN9OuT9J1HHANkRw9Y6l1CYl8P+8suTuqxs2pTPnM+v27Xi8CYZ
7IR8qkOz95R2ih+SlhsqqPFwM4XOeihUwyJc0G7OJyNSyMCNsfbCuUPCTeq1
JaSmXSXm51wk6SwIomZ79bxOoGaPYudwpO6q2ZIriHu4bKo1HpGYK/CHWu3L
ynyzgJLsfW2SQkA6Uww3PvJqO7xO8KqBLBkqjiz4DidOTADbNJ9c8YbZ1Oe/
c7zWLdyl6SMDOywS7107XcPppt7EahYY2mpkRJFOEydhtRsHu5xo7HEaVter
/Qtm6EKYen3Snf0JBEO15+nIcm2+1uZbzNM7aK1zjw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V+yYTTmU/2svjd2EtI1fFx/rN6JjaELNi38nC4KaMhqhTtZ5Pj/8b2p0YS/g
Imm7YEuqM+hixgb4H7hVvlZhWXUz6mh8UVj+rmot16RKyEClPi0T97dIdweW
+qNiRHp3fTnpTLXjJM1+HXC5zxAqrR9pE1usOwzpYTXNf1qr01D2gfoIu4q4
7nyzDsEea7CwtmBdrMkTMWbTd71N1SM71i1NtxCIK6UpKuiqA7cyYyI+UETS
2qSnk0wC17xRUswI8wK4++wZeUEVvXLEqbyk5OealgcWPCsZKmzae2XgJfOy
r9kD/zn6itEPzNZ+8UM/Uh5xc4gjkecH8YDmhtqT2w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tTk+zy663YW/zpJYCCcAw/cd3pBeE9gVCTJOFEmGAdx4gC907F5jWzMzaGKY
elW+vG360EbnH5Bhbii9uSWzg+uLNMGh+JwEzCcWFm14Xfg7on3l5NQ6ly+K
pH+A8/2KW4/2cjowBeZHY1oYLUK1OQrgOdye0Vn+4XoBi3Uu+S4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JW2f2KZjTOHlIy+DHEMEC2vXgmS7VcudztWe8fD7XldDesptGdilysnrjErU
mnBjWGU/Ksowc3UidIyuYC1EmBPgyuui4808HU9vsyTrN5L6v4cwWNxdQdWf
nMF1+hFnfRDIKLUm+e2mJZjGMPe7OFMvJtfiTrKqhBUYNOq6us88AH9/oGbA
ozvI7qE7TUWQiYp9N62mBty0WC9cGn+/lr7vgpfWu+TAx7W4hHLtETt0ixvt
/VzQSsIRXl0yKoRpn17EcCqtguTLMS3s6Abn7F1dwt7F01cNrb7Rr7Mip437
c/Hv5pS+18NFe8l51/BSHsNdkCiSX6b2Pn0YkIgYliXfUi8TDAvQEK8vjKn6
5mfhvALSKg6L2WGgiGKv5s62oXMcEyg01Xg4nW2tDbVKOcG6Vz2/N7sV3kfc
YBK/aYcB3WkgAF22nvSjS3Ye+hqCNXiQNzniH925hiGfx4B+0RzrfCbhrCuQ
zBK9/K5H2VZAPMCInIosd4UtzLmJ/5Is


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J0k2rWqBWHmqBr+RKGBXOERfi0WOI4U0jkvxrODVvMkZU1FRRND+EOEpI3iA
kfbkPPsb7A9yPpN0sh7aKTmHD2RVj1muqchfnpfD+K0Kg+PyMWafjbffSPim
pcinQPysN2yNXBNSf4eYTJ6r2iBv/esEelgXUmmU8wr3NPz1BIg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LFWKPDoZ4J4U0bNo77fXX//WEtyaD4Z6D8GfaBN5fKlWHXE3H0GdjG7nrotd
TT3j/h9YAVIpx6UkhcvSJk0K3tiNtoNpEyeaj8Natg5Hj/mazq54uhiKlY+/
XRxjYJibDyMPybHNG8joAabCh47vGMZyoxdcZwK4J3LbtByIHk4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1328)
`pragma protect data_block
+iUh/eTEA40oh32PADGuzo51p7ZwSV9+53cJg9GNgA23hDrECqQ+H+zKR7XY
wPG+V0n7i9hEhHVTwUVuuOZYFWjwCMoYdkoY+YpuvEgmQZ3shyqkcOCQ14Gg
hdreOJkYIgq8RC/RR4zMWjGLMBoV4qdc/3PaEU/G9CM9NWfS9IYM/Qrk2ZbF
MYtjJN/IW4D3RDdJiizY1f4cCsNMDR0P2InuTyDVf1BArMPsPqOs+ASOnHH+
e84SbQXAXvjdsMZ78PBRAozHQXI18cu6WvBOMTFQavtDslg/759V0S/TT417
NqjvlujDqF9zU7/DFl4qlay7OlrxBW1GBpiVJ2zeGUKhRTzbgHJJjgmYCKZM
uxAlpsxKPQkooub3ogxEMCA0ybFIBldBlZGMzXVpOeRznX01Pb6OBnIgTCHi
E8RdIbYPL40rJIyR1njQd+RjOR2qVzgiuQBWfp58stXYf11J10OLyIrtZeQe
lppX5jPHlmbkdot5iIirEIn8drZEDfXHOdCmP0zeMvMFValHWbKNINaZ6T50
NuevYZuGFJqvZIcAyDnBV324K678WHX3I8kuVtVwc8jK+v9ASK/rkJhPwXwZ
SFGxBbzKYBQMBP+0dSP0pb9jm0ulZy/1UIdpf1ecozVurXIbhODfEaPXPd/J
OCk/idvC4EbCimTEwwfGHeGIAN8DHu1Lz0QMOFg04wq1iXhhucY5vLAJaHyc
1aBxIdsWx+8JsJEdviHBX1MLzMgpCgfgJvhXkScGEQUvYaGZH54JWDb5NIO4
0MLq5Bper142Z20+js8qKoLAl1BT/fyWS75IQa25c80nAVZYxkE1myL08FdU
tgmWZwOFvV0TBn2RvT4r6g2c7r+yp1A1/KryB0FTP4bnzvx+TPiv9Y2VRuoL
hBhDj8qHBuzzk/NOCZmlHjqx3uHLiWjF/yonQxnWnwdlA99xQFMHBVGAEwUi
2dGHgr3Xuu47ip5ZZbE77TBlP2bsFhGHvyVNjn/gY3UlneMneTJMoqJ6DxIU
VOUUTT/eDAxSpETeFPr2VDnpUr/BaMUBIgrlCCNAZ4wOpewLKl/Wt5PZCcvr
jmNm8Rnxa5rhO2L+y9qMF3sTGv8z4cl6Y6sAwuLvvQeDxab3SF7CM6amuTxd
A1jSboNYyNPDSlHqyOOUDRLBL0RDaY6hKM87nwPdVz45Ntz/uKxBayz0RG/L
B6RhBBy6N5tDtEcGmeLMVlzdytG8C7OXpwl0AxrOjRkQg+KoN+1bgBvyw2AB
C4iz8AHUh9PNRDDtcZzgm6UYr6XZyGk6IrduompaMrLsOYtzR36/+wz15hLs
DVMDDNN48LqACn4G6xDZGKi+lvBw6u7XHvFVnyE/YfFCyH1OQUNqewrABoRA
O9NmIslpY5/iUWib2EUUJ66FxWOaClxsD7GcOQ8aCARtxeSZwvd5fYFPxF2U
zLXPPCiRAcwcHQ/PozQ4vXblGoBposTioAfIogu3zfDNjKwbGB4k0+zsc/GJ
pMCS7aVeqWNOTE7W1HbeQTO1s9hm2tgy5Tnc6TXtrSfmX7p6FbVSTSXDXwWN
7z6XOPI4xG3xKXcVvfM4CndRQBg5W1z5YBVLjMrDFMMWzYRbPNiDkO9rgX0L
r2uhnWpw0X5JJdawuaqNnVWfGaUwaEvUsyGkSxvPjbwMjfKJRHFcSrgb1vrI
WpbDR1Qak5dl9l0gC63szL5UhGdDTgNHDEEUzE6BoHR/agXis4QmO/zNfa4p
B98/Pf2/FAYeN9TMqECCYZCTPqUEHUA=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qTmERRtPYzm8P+9u/hp/5ioBHpnkPQ4aFVALBIM75EfgG10ZVX5blMS3bk0vMYtL4xUyWxWwSHS3JYff0RTPU630fJH6v/lPiSCW1Fn6KMJYnc+hht8wAb1tKkuKP2ZTeAckTTM5ZUtEzSYCRJJUgvuiijC7E+SKyhc+1eS8UNhchqX26GVZrqqEGy9ZXhIcSO2z6YjKM3p7KuwVrITpK7QvQzd//Fehi+oH6JYGmT5Qdn8dT95RWtoNz3zZamKDRhrhhXpg+1rkArOx8l+LwEPRCxX7ADCO2EUP2Dq3pxEkjUtSKcFZh8bbR9k2Pcjqp/qERLv1XjbH3snmicH0EoxIsLgbsmLB8nA45nAGIapYKGeqndmMoIMSe2FZosiIjbrW3NAQLWyAb2fWwY1n+wRH+qEFqlYss6Y37Qb+iZ5J03e0FlHtepPAVit51/+wz9xoPyQJ7zd4qbCKupvmRDUt9w3AwvXFXpmRbePBVgNP28KrJw1gU+QlGwueL//QbIz+MZ1ogqgFNEl0DX1+xiXR2nESvXX/wKY2L06e5qSTu0Y4Yj6Z5WNGm7TLSNhJMVzAJA5AgzGEq5lRNO4KP61oRrIWLAnaYBm9iJjJpQMIHLyKuLxncp9/mar8VswaWf79rWBGj6VVEoX+6Xqtht1FxP4E4VQJ9p++n5Vk6DCNanV6gYZJOk5uTA84HV73XZsbLUAxrCBZr377yqV6rSPb1xdlL4XDrX1lDNEIkz+N714Gtt9heC8H44MSEDjyuIoWt6q6BcgqaLaKGlP5y1l"
`endif