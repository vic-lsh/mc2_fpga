// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UJMkfw9Fzi1X+csuHL5oOMRqdWvAhjz/mvFvk4gR6WV1G3GYOdSYVO6tkShJ
BQhBvOnOCUI3mqCDid8KyPiKDKWj1vASkJhOP6ufTsJ6E6QgXhhKJnsv+Sge
1po4x/fXI3HZl8qpIlXgGJbnzka3JyQj8Rle0lYnvgwsmsK1xy5Yhj5du8vG
jWZns4XYZRtPdVnL9uJcWcHzCs1xrz+1ciipngzKo+/0pcY8y36VFWqX9k8Z
Kd7wlfvJ1vajIv5kWOcf/QEc7ia4ELaB59ys5xC6dvb8jJVRrLvXnXevJxQ9
HqdMNRI6w8sgKsUgvixpl5vQNtnmJJ3cut4W7XaBhg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gmFO5aY6rMRp5NvovrIH2offFhCsr8v9Uvo0yAzozePUhEJU7wawQKOZ5ojU
d4rTDQyKSRjHBb3FKLeRqKVZIMgeE3WeWdm8mFcJ5FXpx6Vz+OQ83AulROyw
N6hTDRmLVX43SUC13yW7X5E5wWUgbPk+oPm2WfilVMZ/8aLve8VO533MN7FK
S1VWr0+ojPz8HWZjkfSJb3CJ58gImPqctoOLwQ8pz920D/goBtfTCqaKLMKN
dkEEuiHZitHY4L9oE8xQLaH+S0EwGS874mL3ZTeBMvNPwdcBvsvdsDw851CB
NvlNpiAp4LNEmPnDEZUvtNTR4bS0qjY+xfWU0RI/nA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J7nFz0wdNHPXI2MgJ9iuj6SbgVM90/Uht2+Yl4Rgtabb1REfdX36usTzvd1p
vT3mHTaNsh1Hq4j8hlxUvgv171CcVHFtIB6FfwuxoHGsvIf4uuGzX8XECFfe
Dz/ZBsWau6R4dLNfa/aeJay5NC7+K4FB0kb/iDOTuuQAtx7ewl2eGNRcsAkJ
8TZFPaC6NjExLVRcf8zHVSaLm2+ghrqeTxRVWNYK8DyyBwiT8TeNMY8CWgSf
1bwa7oXJtrjQ8xA2S2Ip3qHSDJh4yPeMitQ301qXS79S5YAfEreZCA8rYVga
4+c413KY2OJHIrmYSNkfRlE0/PuBjacUzWOoRmco3Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J1/thSLACom0zJrfEuza6vy/HSitAGakEwNuc2G+4Xin/WdUv6Y8r+tJdJz7
3R4ikokJI021VcoC5Xc5ue0A73uKro1bMMHe5BT+hAqTQKKplAbJKyeuGz7B
4kOsBTYOuTOrJl3g05Ej4YAaXwTycuDf2W5AfRHCoEd144WYP9dgLQ/UzDPW
fsTbkt3x7tYW9AHbHImxsNJ1qMqNTIsVEMlCFmQ8iOmxYhBqEH/fAWwPQYKw
J9mYQH4SdPrMcg+RK0Au6u2vaeeGCWaQx7vDHxWntnYG3ClFQIG0chgA/kal
3ogd+4ifzAndD7K9YrEzxribOx1jBrpJT1mFLqo7FA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bEZVLkUrw/8nSd/n7C4Ze9VG3oPr+5g9ZulI7Mm2KI1prRNafD76RehHn66O
R9XePJ3/QCqzA+c8ne68Zslr6XPeq54+gOUqGBlEDHQQcneM4UpRd6qcGC3u
BF9K6mgYvA70FOg90QbxQ37iQTl4EWYpQbEPykveHSHVuryOi18=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xHDl5ke7rLlMtqSdzFXy6JYhrQqVKBPJE5CJKautJseiltCNoahKh/yrJRET
759lxSCwciGV6vZTu4RkgJbkTwkT/NV9xn0DJQJuKYk7Ddu1hDXUuEHhCqpE
WdcBjBk08kUucS9hRFodkcZ+H6u7wUEGjmsqt2SvMPnwQTpe2KX+vSoviGLd
W7G0NnBhPAx6FcWUrw3xbrZIHeakt6gdXod2rMMH+3bwoRh0/m1EXVT7As+k
JvDsTCM+CnxDaJ3OABCYS1Ccl670VAda49Y7gr3QJHX2ITIcKpbtLzahy8Jt
Kf8+N6VRqe4O8We0s17T0KDA51mqem53bnnjKNYmrA8CVKRwbmELMkTEIoNf
4ndk8DL6T1XDjg/5bPj7l3Hm5K3V5SOLfgTknDBMSWk6EvyI01RI3/BENT8Q
POE+ozuu5ryXdaULP2Pwbsykh3/EzVY2Ido1iFXmGcH6f0krzzYUvq0j9x8H
Dp5C8Wa2STu3DCY0xQDKK/J/HXaKO942


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
O9xQ5ndkG/lHQu5jA7SzOnvojgdv8eBnZXGe9dtvMq/p6/Fl0RZ4+fgeDz1U
Qqy83ztiHQcTv9F0S3LT3+4zPpKcf7ZE7syaXfsFPeROVmkDBcIRNOvQ2mG1
p9uaS/ppHzD6NraTftVaFjSZbIuJXNSlvsvWzDoOexHY3j+KDSQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HZ0j8SxgMoOYl3hn1KIEB9c1Xhy1fDxYAQzTndH9ZFqr21j8moxkEfJxgn1V
YrlwzKxijp8zr/X64yTyPeRTi/15AB/Z8vN9O51VCf4K9KkqlNvjOzxyNJMg
tAzl5Hd7AacFQmuXHt+CPEVTkuPTK+3spUOZjV3OZKthRgMcIUU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2432)
`pragma protect data_block
fdAf43R9qBhfdMk/H0QImuTfxm6FKhKSRR7Sm5sCrnUkZjdQhVBN27SbQe3v
vdtiosRbpsnJTlhV4mhPRq9/7nOXMr9uAMtXqO0C9l35RflosmPtmjGIXRb+
Jz11hltZ9MLqZEVT1e8HUhn2Prw0DEgZKbXW237VrJ7kI8rAWMbW9J6tM0Zd
wcFLy3pkTnsk/nft+p0B3ZWbyS3qgulLayrsvPQ23vNDf+BtaOiWLppd2JFy
f3jT60nGqIUfC73dYhd+sFIH6vBsaSxqCf1h66IrEW627FPmFEpqoyHCnE/N
w4JoknRnhLK5rTP13jnZvMNgpDzze6AxSHxZ6BiIjYF7sGnrC15HvSuOjQu/
G1lyIzUjzKpniIko/NWrkfaoDRMJZ6d3kpgYoEQm9vNYGxdjPeSnnFbl7evA
10BAPo4JK2K6HFCsMTg/VH0/M5O9bggTlV2qs/XrREBgb1bjbhsYagztY87A
pIbzS9qUdesR/BrkhfsqIqm4cD0ldhEep9zY7mi51QTScSBoxG8N9vVYlfMU
qspZ5pLGhvXQZH9VIVSRO6v0LhA8WcRJYuQlafQibDvOpLJzA4YCZYT8l6lO
j+url31GewGweN2cyNY7t+VonZyKgaiRfglxTtK4kfyjhL06SxSfdgjpcn7B
sE1+QfR0LCQ3kgwpEKPgky8iWXP3pPz9IDL5dA5XNqObcF6Iay3IKMKubZTr
E9FJERMm7ODlBKAdDZHRSHPQGEN4iaItWjOkVUcs1lxavZXBNLEsGSfWdBQH
m7AjJMKxeDpMuZurEysBvsQ+ZcJHN474hfrJsuQVj63jm1tIkCqRIqahTxWG
Vrm160wiHKeZG/jT8VguOAWrdfnpnfKwIOW30GO3wrMjT64yaRtOL7gnHxYC
6l4QFKrL0BUrYIu+1fH+3OGAA/2au1PH9m6AvZRl4BFhLJr1djkP7+wglecO
Bq+3hSFj7GdR2UxSfJTuT7TrkiO3oguhnRxc3nK/MPD+26GvI+F/dnGfano+
LGCvDLRK9sc05lc3VJodv2KC15unW45ZzO9F0YKeAGZIgG4q6bD16LaSOZPb
asSMkgz8yIZJPTmg/UIXOy5Dtzt132LQEWF41XysMNRlhfFbXpJlsyvzKed9
mlXbkk5H7rnl9x0Uvi6RafoyS7JQMlkbqC2/3a9yqsh5X+uwG4VXpvc/Xgf6
XnMdarKHLGhkeJ3CGyDBbclulDhdmhSreXgtSyrTXp3YIBfaIAcGA7+Zx5ZG
zQb+rukdv71ItqR17eCjAn+GK/mmxlGm1TTD75aBu7YLdrW2C4/V9jULK2BE
5i+5K4Wo8Ha/7jhqaC7AOz5T87eOtougYODa9b02g8Vn8X4lSv5Rhx1/mhE0
if7FkIkkgy/31W30v6U1814XTA74EHq8AjBk4iOMn3elSPDre7jndXPv3AjY
weDBhVUkZSVjqpBgQWUW+ewjchqkv/nDlRjOZ+E72fTTJQlDLRtaulqQrngx
SODccPydxGBUsHUjZLtGohF90lbClbkjPSuwOb/CLwEpaa11Gzc53lV12Eni
jrK+aXsdh2OvdaPGhu/F9TihcPikM1TuFqv4bCdWtlbWKETAFZMTm945NHlX
POjoWiXP+dWaLuDP2qd7kbncZxE/FeWL2LKGi7G1amSYhIpq5vh2x9DbdKyc
6EfGfAyyepOmLoZ29XqONGzBsgq0l4Wowtsaw1R/C97rSCOoRILQLJL+qus4
CG+LvvI0GyS/NNEwxcim2BBPMs3Ia5Rf1bVJ1XTE6O4R4a7VQ67hMva4void
LVDMk5YcEUE2CAPUdvTj1F8kAbDOSmNy+zJyITd0WCwFxD+eRvlVCmXpDk5e
tNUocb2w1fOvUO5dAE7HVz0GQMKPhLwMcLEE/7x8RbHpEL3tw64GvujXfgLt
+MSv4HlcINQezHgZ1pnJsbBRhyO86gO34ShxsJ8ieQLuG2/G5sLBvGWGuzHf
73zH2Jk3p07wuOgK1ON5/s1p04P6sKoRRZHD46CSlAloEmi6Gam+kZuDFP49
3LvG+G90UqU6hVSWNmPwYlNy+in8I6p8e6/oH2cRRk6K+6aDNdM8hdWy02/f
e9k+mw54fMiMYpgaaobyS3JTj1sCWCWJe42SsnfpiAKTKJ84qKn3N2S17lUI
4gipePZ372I6t7vKdmGE6+3/dUIGVq+98ngeRpPzFmvnw432mzSA+tlUEsMX
isQBnTBwGQk33E3yEa/LBJ/E1m9wFMgOBC0t4Sb2OotTT1uHzaWmAgOdRFlz
vHrryqalzFGnoqvqPaFghq9OeMPmGJiSExXWnAhm9rFIX2de1X3nFJoSy8e6
ZAIuQrkBiuo82IjbE90w+8w583aCV1FvJU55Eo7/h+HeW5uiZWrsxuQp+xdt
k2XGgeWyHeekFE9utziMrMO/8Dy2tM2iSGBBROm8rcoohuPItA5P66skUby3
GRdiNUu/WsPyKZK6H+6sBr8RPsOjDSJOJ5EdZVEfNUwS0BcoBX+jDBwIVuba
Rpnty8QNIs2uwKuVTONahy2nsIEqRNrZ8CKXDor6xF30goZL2HiWNyhQgfu7
JkfnjbB4CVZ+EEvfFibebTGmcwGtvLUHF1kgcPmA8dFxtsXcQlcOWS97piD8
4rTn52pe4gUCueziAqIunYzWGB3qnMbeeG0FVOahKEdbd3zui0E78A29ZsaC
mowZ00FyQa3NmBZsCsHDwsiVita6b6Eb5X7MQvq7nmCB/qCUvZd1Tj5eWBa6
wOSjXz1+uf+LzaV0DUdxCmcrZuhsvRk8qKl6TfiHgR08K8R7oRMltcGPRAy5
4YxMBv+L24u4oFknxA6JmE/U38L6Kf6GlZrmgwKLC0AROjNkAVlclKX56rAU
HXaQgcfb3Xag8K7FyA4huxNUKXl7CDl1JCXGZR+bsPG0CLZnlAq4hbpN6rtR
qsQ8bNxm9G5iXZ1dwVh1QFQ7VUN2AEac8cwL1ujkyTC0nuLyp1CcguyJOcw2
UOOcTzQNhGKQvq2tB/8g6ci9z1Gnt/YZrrai4IdstUlm66GdqCvKdG/hxedA
tOPOV02/gv0fK8M7JwEdocetcU32gTP4lIL3lLgoZpvtPpkw90L2CV+Weoih
2ayjBx5qZP+ES5yrdz8zr7Ibf1LSfdfy/Hildph7r5wWSv94y/9lKNRtmm4p
OpqqeDHkQ/JvM+ixFp9H296t68GO8PdUA09q1CkHYo/kFsZsft5828bpUdXg
7Cc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyJLjKZQrt3wGAn4YaYK/CjZWHcRi+QiTAlUPjz8YV3wrjW5mqEZyrmVOJ/kioHA/tEdMfzGCxpZRuN7/lcB5ZsLX417NrJMmqNqQ+/V8O1qL0skNB+D96duiEIuLBLgXh9DgXVtpbBW6H/g5qTZJTyUeN4HJiSOHjCRq4ZsAf0fH2ZE9+Onye5nBMAuSkabJRpxUU0++BSHBPKsfnoEhbGOYntJdm4V9NtB85JG8XBPZKxOow3yAOk7WcQNjsPuSKa/k8FPo/qVA7xGhh4ocWTcUCPIq8Pne+Iq9tLAG+8lieehzlZGdVV9sAx4MnXLxGoMlP0G8J1y7BzrkHHppT/u5/DfEY5j1Yc/+W6px8GJEjZ6biMAs8Jpo9B+ViMjD9KrHPcV4mrJWw5xdUj1IEWbpqISK08iaufIXBusJ/AdchAts47CEONJCO1TDrWZ4DvGawfRuYN7NX26wsEuU46uT056HdXxEG3a+czhQlRYWdM+jNHCdPLlK31if7+xSS6S9GMp8d0NbDUCKnUbfJxjqn+rbLrLbLyp7pxEHZSPWD4POHP/PYTJkQh64Go/6OyqoVAUGRpwEmqImvkeyUG8UGDizKlsTmlVQ15QP2ZNXS6aE8dKRMHOexohzY3ny6giwz29NJXdtzr9Foz8MhkUozouQj52TqhPVMm0PLI1wxg2cnJHr5IJ51l9/Xj0FVPGIoq9lawIwks48Vmdfk/i6YoloRK3ULfj1xC70G139aFnRReZTvRLUmCs++6dfM+PwUewqW7dk0bGJIaJ5MDB"
`endif