// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ABFyF7TSosarRcAtXI6FkJjWREPpMh/z0RpbeLJF13f3/wiYj9UohhXLmUJP
UbDz8ORpoKUr3ugMxMslHPA9K6mw856qTTrg4iOKedCzkGYYXwLMow84nFq2
zaP8WYD0OIvt9b37gGmF5lLOs1Tz1fjE5yB94K+XvDOH8bNpYuBNI7TZwoO+
pOwSVFfObR1S/cPccd9DePSjYzUINdzVM/FdCf3sLnLjYaSzcA9zWvGsKuGv
gIvU6fXjbTl8vaRXCwcLEuXLDywqClumPPfhkxJ5rfcZRYYE8f6x7x+Lh5f8
dHIh5xzVSIRoZmqPXkJHRoY/0mrWCQ2+dbc0KgLnOA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BSC0pA1I2sHmcdnE4QapIO1QS/ihI/glY3AeSoqaVpKlbLu9aQtazspA4aBQ
OwJHD/wYpQugzfR69lSQJ/sVe0BpkhHmLWmE5bLIUfZ7wNQPxMscHhu+ZsDd
eCDbNCsJenRt88sWgrzTDYaxKIVAL+j/Dm1A/6777LWUbkM6bcA4LgW2LCBj
VSE7YGXB9h0e/WbGJBxOoJ0lFco3DKQu9WEtHOotiP2U7LuV2h9dcU0BgfLx
OzckPxMEkhEfC7ek45p9bp30gjwffBHKmrIXM3DfLWbUegZfoPdfMoaIFLNy
ftjU3XXte1Wvp/nVi0SamBOn387uDV8InXjBsa8cug==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Od7F/gpn+K/KoAGRV2kf3W+VZ9vMgN3uhN02oSb9mnefRXAqeVBZu5MOEH1r
tw6ojqmJVFI7sgyC1+oS7EUGn4mQ3sqtP+pBH13lYXFeH8KAdk7j73kKLfgy
TebszWL7+xD9gwHT2/+wC3VgvArSM+sFGyLrcoXfuizU4/cri4526WdCGIjk
DzmDTFxGwHtb9zfBPhHckGNwqaUX8TcVCLuCwSsLTOpep86PTFZHVs6qo4cE
4H5Gu0yIPOC/hxqzLBtoaywdq7qnKTGTBmhpUJ604Jfon1LTdoJOwIXjaf1/
QKwpEjCs4MAucjMvjhZXdesg61e7ZxLIyQcFVepbYA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qrG78176PSmNTTIuaumU8FZlY9Hdkwmsg8cPVX1sJwgX91thL5F+sHg1g2ZG
cnh5xQicuJfYPDV3hyn7LGuO0BTr/qZI7eSWm5SUEano0puxgHCy1OFAnDsl
EXK2Z3rJLjkIXyt2Kcn0BLS+CGgf/ZoK/dKXXwqeU70//VoIwjeNrEiXA7Et
Vt8dUnMdFSPB0g9I373h3lFfvIptYV01MwfkZQsK8Qi8ekgC2kVvfT2O3GFX
zsHY8QC+XFN7u8Y55IWhlE/up77B1vXFQjxYyQpOeqiDFHyjaCf6gq9+0IlC
PYFQwgjFvZ2JTlZ0Tbv5WPO7LMDTVFIg5QSWYGntbA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Y1LuKVwijolW8KMtzHzwtnZBVShru/xBhAZfnmL4bh30RzZcYvD/YxmAnJLw
7hJ0y0r6jmyQtlad5MJYkJLHPlvRLqIqPYU8B/01QAkznIrEi/bHKjwKesnq
ph6Lqz1VEBOTv2JEthTU2q5tRbdUlyCykCLKn0dGv9U5hUNSwHA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
p0ta4QyGIjgKognQszhXCaZ+GY/qlm5L1hzOE9uMzq22zvTXFw/UV3JWEDH7
twp6n5B8cqih/HXHIfe4AfBnTJ/aKXkDG9UetgESiVY6ur9vKm6JkiV7WMD8
KVWH4C72WAIfbHsDMn06hkK/soJ9Z2nlApksENG0w5u4MYVecgjiXNzp7ap3
IjR3nNe5pnwVh4XpMaDHO+DKOQBy3pi05nYphV7Bw0r/8KqyYQShsjHoKc+i
BvQyYeQcgYuQo7LXuQ732OguWF2DDybMOepq0rxxx5zTqklEJPtzGIA5XiKd
j9Kv/V9opsJdlgcr9ueeKbaRX7L8M30XHR4osHcCPbbKhaOAg8nD28iL2qub
CZedbZlaCK3Dkhm36EltEHe/j/Uxp+JxkPYiNCQjhuN2TOWK8cuS2oPUsBr3
SnFwc3ZkZyb/V1WgjMbO+u+u4B95+DKmQS4RlbjXYTa4tJmzX8iNWLVA0YLD
D5ausnJQEUoQmYE49LqvyQngYo+uzkZj


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gwNl28aN/ld9JfsxLFm34Lq1Vow+MXLSb19WEl1hia/ykhAtycDvlw/VCXK7
cbUn3xIgFR1wgg/g3FiYVPnAR4rMao76OzczGoseG1Wam1EzH9j4pbsu7WJg
uBo0nkZRGfwpyw1CGybFc68ZgMBKvhnnJpWOKYp8qU+O4iDYdus=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HJNQYiuhIZjap/udv5ss0tbwdxZYjyo2cwcUOpgGLgLplUtblNEaNNbUV4To
sQtOx22EdtMXT7OyYa+khSELljfP0aDo1+RhSBbuMaRA+4unxR6c7aeBd6Ic
KUeOMf9buYGizQd/ULhMpDxDY6BygsrOfQdv6wdftuPfo4U4DXw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1744)
`pragma protect data_block
kqvXfh14zMtd+OyfeFGSqZppN1ikBl5UyIk0gyeDp8b7CRJ10AaE2gZ3eeOL
w3O74+SanNl+5gnxcgFMk+tl3O+MGAHhoayjnmcHvytzmyEUE/MMRESEZETG
u8UR+hrHx3oZUf9KbZTFTQ3JfrQ05Vso80Qyl+39833OStlmhW6YxEmgjkRn
OlGMrtI51bQuvRIurVd+dvLzKthWnU2QsdN0b2VN+PI3hlcfaPY+Hj3qU/tM
uokgqxaF9TTnrC2J0k7HNJHr+HuHKeGp3iyBrWzTjLJxFSEOfm68UXKRzhEX
TccJ0QHfxtETu8SIYYykH8yPy1pQgJdyfxLaLrfgte+qqO83yctniwc8acMi
yM0JM/FB8f9Twjgo3hFQgYiLrmzlWcINRGAGIoYjFRue+3E0dE1cbf8v1Y7f
rIlJKUYxSNn3W71ToVkv5BW2P/eZJgqIV85pa/qe5sgr0hnYFVO5ogk9GM1q
QQdBU1auTALqGPfkQxxv/ENXiJiI21Q4O5UMAf0P3PUZIlKCQmZIBO3gLvNX
hrmOXPbD8GHeoFGyg9tsxX5/ryl/HJd7QxMbgRUU8m+xk0aBerCG7gX1cKlV
/oLISb7tkacZzVbte81gATfVQHobd6M4lc1tNILBJOcBDVnapMXExwd2nFnL
2LW3RnpJ4YlolXVsBKQWJt0rQR5HFVVudM8WrKBApoSueqJRFTn4Tr/QRatD
E5+xM2O6+CVyJMBkBKuHcqI47n4i/WvwmTDJR6Z2mf3dpMnSBI1J9EryHFrn
gLpEtzfrb0sscKzTOtCNc7zy7YYP/r/AUqmqMWM04Lze86Lmakv3wMaODkPI
855vNRa4xnl3yfqUoWsuUfUCRPdn2B5sNlmxYEIqLfvdAYI2WWn09EO4390t
OIu80MRoqSASIj9h0YUNZ5dDY4YxEKBSBaTwFSZGk4EAeD+eca3r9Yatpj56
H4WI972HRdLgGOONiwXA/Oy7bCwSVpI/ctYsiRkgSpkp+hen472+Sv599iDn
hG9ZYuxfAmBIxTmC5TExsQeutypwFTLCgeM734gjTBJT3/mbsujaE17zoAQl
THV4fY+9x6tyrZFbyjf7v7JKwCeXI1XZmoBmFVcllh+z2Cjjl06yoRw13frp
wCyL7ZTDr66U5H4a0vj81Fj4Vnt6Cs5dNb/zYfc6BGvXFyuUG3dOQgXrxATy
sAezcfYsgy/SEDnz99+apqZVTbiBguilIqEsTa4v+Ypw01wZ8JJJ6rz2YEG2
4qGTitkl+hemgE+Q4o76oF53r9JHNV39hpWfPd3PZocMBmeZhjm7qwyNQSj7
4V43H6Ff5Qww5jGnTq3r+VIUQA93GaPROKYsW5bf82soqDb2Bn9rkYBpf2dx
NZzPhU6uLW3yU4rT5T30J4yqtTFIgpM8xxQtmww/uHy/mSmapy+RDJTv0df5
u2tMB11/Yzqo8fLuxIoj3R0wLQ9RU6lsrjdBR2b5xdv5VH+XURjSX9F2SQAE
+OfiZS2LXqo+qGflbn3Ul4xBBipu9GEZ0GtyFvmquSXZxMN+axej71cGpSf2
L1hB1D88xnSl7Sk3EwlVlIbJAPb44Zen5H1XcN2HNrldthXHuP2x5S7ifix3
KSHY/KiKT86OCGfEu2lTXGVeGcQI9j9hL7yhdCGK7NheyVK7MHbHIYcMAQa3
E8ocXzvl8sXEAGfwFqHoYcUiu0q2kJwre481TUD4PdtGWjaOwoBK7983NQtt
248rFTo9gBBqFs0pBvcN/Y2qdeBzso9USdXYDhv1oPdwQHGeCO4ziJZkyJUE
cYaPDDComE3DyH8CN81SpAOpl54m8RBRpCreUQ1J2VYAaM+1vtXx5c52mLS7
5Z+PbbyGJCWQpigNdClYULfubipThZU9CnrHEgoKnkOxJrRMwiK/gTxqiar2
OSy7plU1nMI0MLfsma/GOfEVICf/6SY4qHlJQQZyd9CTcpsxb2A7DbD/LjGb
yOX9Aru97OUJJUW3MgPSLdEb+kjLnW2lLaJnjGsz4w6Vs+5FEAtCsF8C3pZ4
wwhGJrPntXcrLzJMXG2YX0EcxyjpaiL6cqRgTqaWGJ31C2tG5miwwS7iZPrH
Sv6c/uurIhlwbTTuDgMhnGdjRiOUQ8R9dqdx81Qnu/tRn5793YQ4Y36ZNjba
bXa7uYL2G7DpgjR6ttUWEgA/01UG3AvFS0wH8AOmgiwLzZccn6TItQ16yy8S
xXlQ9I7uvBU6Sx56jrqvYCZDWN/7DCFlHwprdfwdMQ4ixWECZ4eHkxxuOS3q
xjbeyvg0rHLqretrwmbrGC/9UHUmQh2lc4D0eA/i4t0NvQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "9RW93T28GeolckbYRvHffOsKFRFmORm+azyCUYhudrVC3P73ufaBfyRVMCXUVPfCA/gVx4qupGWo2/MTXHrbiqujt9kp6+gvryDIvlW8esKlSeDbKqIxzhLY+DL5yFAjg+mCmTKnMSoiZ9J0N0zgOO806IAkac+OYN9FbEIEFuaO+G41krhhxrcYAZ7qVX+m993ig0jH+TdTkf+bgk6VV++svRquWf4VNDUj099hz6BzqUVu95eqfdZpOrTGUMeCmjP+NYR+hpR8sw1RcGr99V65qo2jOfwifVsGamPenrWOELatNZRPDSV3wKE9Jz1/EDsZ5o3eOa+0YivaGKuthVGmBuyujTDc/litu+KY6YVM3a0YNnktnkUGMR89v7pF5fvJcBPtqpYRMTz7hdTxH77N8+QyIW4QYqyskk0S+aF3SQamXp8Lp1D9zwvGm8/b4jk5PzKF6GgnXhySLshBdxKtDGxc2OD6ElolqmYy2UEoiyTdsZZoTR7on7ZobviS1BmvXQV7bl5t9HR1VtJDG6u4kQiJmadBfHHUZU0H1Z6/git6rSqWcKsBW94SStfSrPNzaJXvioDpBvnq7Sx75SnyngWIY+Dfgi+/IIz63+Rh8z7GyhPfleHfYrw1vJQuIv2BdeRgeashxr7fy4tr5fZusjUPaf+TmIr3rlopjF4stiHlSWKKik7CkiESQk8dbloas9zlUjgsYjDbZflWJ1aa4Psj+JMcoM35x3G3DJZdgcSVV4OT3ZB0M5ktK7NwkqKu2rojNrtOBcZ0gDI4ed8bO+XTz0bojoI/jZyD+lwpwpT6Gbd+01+L7nQtM+m/9za39XK59nTQC475+SMbCAlCKE3n4ce4xGH7wN60Ozl+Zr8RXawkDjy5QDWd/0lHlpNXoChjRzn3prfE+AVUNG48uK0qOmPG5CoqJY3RopZ3bQa09ATTQG14C42b14xJef7WEuLiH5mnquS8wIXDYKjzyF2Jv8rAHx8tq9TH+CZd377pqu79dQdwDS2CYKJm"
`endif