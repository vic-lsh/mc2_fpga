// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WIBOjrSc5bsHEltUEI5CRKkPvxXcOf6m8AqkrGQKXzNYdIvEugticRGqwQrl
QrKPkHAy1owOhpd1lstYp16Wlh4Y/LqG9k7fqw4THSUirMagOUiaYIZxSNsR
FclMLxlzEoPGHwIpLX7+JSk39dh9MoOdUZcosupmLgUIsLEbQmYIulK1oZWH
ax57bRZWvETcADahrcqmzSO10eTxqi0y0RWVGYJwYX+JVK/k9wW89tpDHA56
RPdEL3/+3T59yezBkUxXQ2YBjmCPkoNA/Igh/pkkDAqAt2IZoasxpGP4e71H
GKEB8TA+kzLuq5gcm0v5eqMKiDCpa4HEMwyZ0XVXdg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Kh7+gORxpaaSDbCFRSHS9SCFikDkC87uVUI1g/FHubkUHRUt91f/eK3eQLJk
Ra0XeBkz+RZQ8vDwb2/fuK1+ursRBkXq1kPB91MXAEwyMK99bRT/CFEfx/E7
8UrsiWt58QqCEd2cyjq64MUd+Z3AWxLNZwa6RnzT2TeYYO1/6ui/ZohhhDlg
jW+4GNXtKoXnqVSN7J1FJLM4lmeVcWXZehYs3dIn58wV8UC2aAilgEeoUMGp
IBDUChmG028vNo9ap0Aj7w8uxQ0tVoqJCUUfa7bPJ0LdaA9Piun0us6Iq22S
EHRThi5Nx80xHcjBQWvCIgskhdFtXI9HBe/U5pwi/g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CGIEBd13nM6PMtn14BrAfztxQjplW0/VZMpeje1jbfiY24lvTF9qVcwA5Jm/
YgG2fBgoWkf+UcuCRRzCJMC/iaRt5sjWoEtba2PrKCkkTC2zV/5joQhGIawY
wWgmIPXRc09Tel+pY7RcnUWzyzlRjImzXgHsGBPRKNst0LNikevMUaVzkxA6
gpg72Sw80R/VS8EfwL7J3tD97D2K3oSUGNP2Dkr41NWwpxgtZHnLOOPoL/fj
Vw+Xqe5JbR/1Q3Q0A+2BzurH95k5QjcJyU3ah6IjvxTaNJpdeqjlqC+E3Hqg
z4PRppHnnqy72kdGfUAJn2dvBzq0fb/mhspj5YvhyQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qb+HbPob3jhGqRsExwzezw0zxi+RL8FL/4c8J1/VbPdY7yMpjEolsoF+7cU4
DFHkGVmj5MOE+Ko3gjSeSAYquzZ3Fi5NMHBRsOdhV13Hiv+qlX2JhrD85fYI
+WUYHTDxA8Plp4RQASHKaHD2f8GwlGKQgg8hnvqzBStYUjTTi938jFhShCHH
lPUHfVucQWsTW+IBuwiwycSRYS3YbwkGsQHiLjTzFVzf7YV5TpR/xJKNGgID
thrPf57JD4tz5KvNJptnGX1mrrD8Cd6WzGqODchiPsxCvBKhn8D5SYc1z/Ia
N3Q0Thdy1fq3AEf0Mk+ZDAm4KwglKsprnbtODZiUkw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KaHY8xWrRbjxsMncfHzr85+yfYNaFn/cBr43kneAkmQ/leX6XFpVcoZHAVEg
3bSpodkoQCRtE4DVzqoG2rZe8nu2mPxiLp8GIVbJK+hQgG3EU4mcfPBh05HN
wdh7D7HGhY31ZIG0ejU3K+ExiSpizInQYYWEN9Nj1nqSSvOgjhk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Z0ovbisZQ/1R55sABKyM19mNUSK5ikDfEG1SCcZlMgGu9TUwCD6jk2M01cB2
vgknrFBnVJACvew47HjMgJBZFEHjWFoIBAbyekzjBbFo8Bk7B+K+rI1FDoNq
q21VRkkFauHnH0DBXOyLMYTnq8/qprbJGmTGpU2EJMB2KmMzvEnY490R1Kx2
BhsBBby+Hw/MQz6XJvp6gc2dy2nbEfsbXZ+BGEioJf0ndu/nZdmwgH2rTJUr
vjyRusXmiZWm9vbQ7Tb2qc2rUTJdnQXF+46Cu6Rdmzl0AI3kACJw8u+6QFhO
sr9EIyFOV5Nb/Pw5bQqaptgupu9UbzKDnQtk3qVgoYUxCr8B2so0kUBY+902
hiPZkiVq+0foP+gqU3nnzYJECTdk+N6iN4dpis87k91xb2jOlpU+V/wDPcPK
AHRc10F1wpn1V+zwuk19TY/5VEruBcVG9gb02G+fpHgoPLJlyBxsYLBlsf90
BygR8xzOi1yBy1zmfeLJTflnb1vPqk2w


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bXHkT/hDoOpNOkQALgr/nI1yQi8t60jvLnD0JtbcjrovqSV1hyoyrjM/TJuG
+qlHP+fbgo/095tqrhFbHerBnGHKy/t9xwCiJ778v7/OMkBgpInLXcBfY1/w
tHYYawz/jLx6hu0dGbo4o7Ri7JMQEfWkywWdbJtAXjXiB5z/sQQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BN2/4YLJRyqMyAFZuSi57DN5vbPXk7dJCz/ce4L5CMVGzPke+BBsTdH0ry5S
YUEArIFionpxZNbFdbvFzHou1ERFM+W4HDzJVPPVa+/7Of5FvIss8krcD/Nv
iqIN9kS7fqBGyif7V06/3qMUEvF46YGU5E9Qet1a9nxpFbcY/dE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10576)
`pragma protect data_block
bAQoqntp5ta3QsYKJoqMEjFytIfmW/zsiw9H+CLpNrTWHeIvw+zGO1YpFRDe
soBT1FQnAccvxbP4r/rUUIPiTZs5l2aqShlMlHiA/ThQdszAVKlQm4Dx7ICl
DsUmIS+xxusVBbQtAhYkAlBLEM5VwLw1co7Ug4upLdYJJGqKvA3Dk7y41QH3
yd59RzDs0TMxJEjlk6ym+XKeBE1tuseOpWE4J4flhyx+E/4RQ7WEfejggEbU
HYJkVPQQ12ZjsCLBkOghnwI+ZNWnLyppbeFBsURNAqKr1sQLZaJ/9+9RfCmG
29TnezI5e6mlZDY94d6k2uZm6AY4Ca53MGgpydtqJfPpzRdiJmfslq5b1H3t
9l6Qla0W5p9We7oj6bFoOZf+R9OyvsgT6/BgAtGGxuiP5+fwy/RWpgLcpR2/
Zf3QWCwtbYm+dfNaz8LLzvPPCekkK+qSX+tOnzPfP/EvJAcNr/s2sdkrOili
6Xrrgyqp/24OncQLQeQjTudKs7sk/c3Vs3zNERa1sfNoMhWkB6EFNpj/+fTt
rCXkpB/g0/O9ehi3omvXiPjzHwvjlcWicAvFbcuCH2Ty6ZRz208t3EB5P3I8
WKJOveQwZhJ7fuI1Q6kUpfvfum+PsAy7Hekw+MuSazNvj3pYqZuG247nkTIR
zwj6SDPMM8LdN7S/A+ct1HjD8W7ggrlboj645J8lfjUZbr7J2HCui2qFrJQ8
K0GODxVqeP+G246YmG0R+epmyI2Nz63afoGOIDjAGg9SQ54xo2/udTbQj2fY
UdaPmdV/g1wtQaiuo9DxjJk1jbpJ0LesbHVXVNPTSygcY7Pm3tTtyK1bEM8t
FfSlh2+GPsWo20+XJmG4uxsn9T92X2QQAC9SQyPUfJx7lKpi6b56/C9yvbcF
n8/u7DM00jvU3NOFM/jTFKEN/C7eLyIVP1XF3OmSagSGUl3mN8zsaMtzRqZ1
hNgqQV22QOc5DZTKsgLbWh51PmepV/DoXmmODTtj37qNhC+d0sd4+J5QUpcj
X4AVBrE54BmeZQYSrf7X7Q1+zSqAUzfoHjxSMrX7crFkurCNvztUbP/hOqHv
ijcJKkTSuGC7FSWfdpDpp0EdywNQ9M6yTzV/FPJIvhNpyGh77lG8ml8l13lI
ENqZYIjp2HXrDKJERnq5mKd7KxIiMP4zykGSCnnt6wT8jqLKGzlaKbOFJrrU
VTQC99DkSunKznmygxmNl8JpjPLQH80zorJdG0tf11fLfUT86vm/A1gPvJqr
yquhJzpVQslg6kf7iBz3InjqOktE1XsHACfb5hG64cT+uB6TxZiiOXAGep//
pTjs8wlJH445H54cnut8tBK0KMzCo69oFQ4vGQZBP3CRYg2zZssiGwsf+M23
gx/H3F0Kd6xX5KolMZppWm2Z6ZIf9C4Mo6j/0CCf90MQfCFyWCF0V2+iOtpl
GgDiloZF4QZAxG4NEaxs2qHAfg/0fX/GJ1qrIL1bFQSWlU5pEIyueo2mkBpZ
mQWzzKeuY+2Cx6XiYvAS3KHyLYIBwE2B33VBkjkR/ECt9giR7evWQ/xFZ0t6
gI6DUlj3nXt7tWKlZv4gNFTmCwqafS8j7TWtSN/I4E0TFNtTVuk3IMtL8Slm
QiMN6XaExdo7Itt0RFJWEDnOE68jaG0dwuD7/qPh3j63URJ0tJMu8P86bFEx
rs2sGW9j5JXjiZU8J1mDBLMd6kOKnuZdXeu+7sXP4VPiu4P9xMQdchADMm+l
4fXCHtmbXq/DhvpPUxiz+yYQ5bESicr1BWRbEkBOqBdPxKYrF0u8LEtw4Zcj
rzsApLXJEj73wj6uypnkjid+DlfcCl0df07qnZDog0bCoSn2brcTctwsjze5
gctE3yZw6+WCU9Li+KXl5p65mllPRRi+sKdi+3SdYhT+i2guvix+qhMCFi7G
yhNR/tMdEd+YFug5WQ/TNMOPs3rzmvowztqFfAG46Qy11ch7h5ORv7YtkdcU
nW0bkPty+q4FZEdo9sfRAWWw5qX3S3I6+xT6GrX6a6V9K/Fsezm8JOx5yYmF
EVzoAvnjXd5JFwSE69XmZRJUlwG9XP9vITTkSQVUZE+QRsVTYAbmnXlNo8dw
SVgf8TZpGyTt4yXfARoQDlOzBd0oiGwCPsFZ33cbBwj8UT+uALSLpFm1XEsM
ax6eXXmR366hQ7HRET48ybRYEzAg0oc+wP+kNQvlEWq6HEG/n6JJc4vVWaVU
A14hu927vb0mUpSR5GCyv2g/aon5kzHrhH4mnz0AFyGnboa1zAERYULl7Z5S
kkirRcAubRwAXAb9SY2ykteSEZgYK8TUHy6hUYAwmSbSownF380tOCaDVQ+2
hGoIf4hlqjRa7LpAkoNqdYUSxOYi4cX7/hBf/7fw1lfNTZQr9iLkte+Auvse
hNuxiL+NIy1bLeVRYOg7ZDY5RggRN9b8IzX+8vvlrfbNR88qO3vBdmkxDiQ4
f4Vp7YFkuKfGLRi00bgsnH1KqJEJHboLDnM45t35KnXH+LKkQazJUc3bLlmr
h8aEZ1wOoQzE8ZdM42qrZxUQJH/gMkKolKd6LKY8zmqer5voPNnP/o8MH9af
JtDWrQCa/0kluMQ8DIJcRLLH6e0jICSlND0zLEmJdApbXO9rRXiD9T8yM/G4
pJeYdOUqHY0RTewKuY57ow+zI3beNR7UeO8AOHLdZlnl/6I/1qu6uAQ0dARp
T6bVWf6i+MJJKxfJBk0HYF/LBKX8XLApyLcfmds++ue9zlUL8hIQamSbeR3T
Kqc3IG4e0YPmldl0n24k1TuztqzVaHLvfH0Bppbi912ywBUx3DhOItnFpEke
kRbJZ4wizWr/ltj7Oi4yuFu5AfPQzPtjAzrpY+dH2zOINZq9P0cMc6+K1uNT
Vl8o/Hag8pqxg4yarFwcC9U6v+uRiQgOfdQq9coX9HaaT/YFxlPKwXpA62XL
2tb2N90eGDN+yC4pCE1inqYbcVvxb/z5154V4Auv7XTC1McTu/JGofYdEKli
MZTwJmq2th6J3/NUr6BMOp0X/EkP+ETz5WEsb883BDGtMMh/0ztWM//NnKdZ
FGv8DTIvit8jrUFYvujTmQaBar5w7kMk/IMNCo8N7hF7qflKCrc+MGRq3U1k
8+ceo4OhEfeVyRxM+UMRN9ZLG04MZcMd9QAQ5nFb+IsSmeI97l+3kRXOPf12
/o5jhMH71XFhv4PqqK9R2ZfxDsI98PDMg5O26kTFpWPnZHwNDRuZUOcJDdmw
2/6IfjeEMc6Ui7FoZ3hFoAQtaWxE5ASUC/oU4ikhNfkKH12jlqYK0MbBqoGM
UVVMCZ/a1BLo4Pjfr3RSXxM4lwlwzXCgdJHSU7Dunh5FrvG2Rl2EMhxarbjp
xJF9pCiCBrgnEngW7swd+HRImbNoTvbW/AiZKx9rHBl1zcVWpB3kuXLCGPJJ
esaaPRzqYHuxElj+iLhhIoat1UkV4CJCFh31shUZXDjfkXrv/ZtE/v8CeZN/
rkUCeR8JJeNWQSEnvC9Ob/HZ1Sy7DxbGWtEKaoJ0RIsyNN1jR6MF69LTA0NZ
psxgU702JgTOPXUEku2ErW9+RvDzszgMbpzeyEGRBMvEO+KjqYcVQaTF5pEv
DPuzNau5W2oRVlZlh9V8yP7Uac4PsqG+l9HdXNi8/dM5tBqjHDeDU49Aackb
CWUxqusaw5lIu1bjfhMwmvRAGdduIDUKbYtsvPFUu1o4kPgF3JB2ztmHKlPl
qREy95+YsjnvuTQQTBf7lxMsczuA2tqFBsDDNMOwFlyKHmC3N/GwKKooUv8H
9sZ3m60SlsRg4VgAJ7b2glrF2iBFSpqXxTZD3gpR76BLdBsGRbKix5GwAvXD
ApfKeCODNVtLY1KKFMWy/hUcqjJnDfao+qF6DKmaknmnIZX9wsnWDzg5lCXF
yyl2hq7cGhMLyiv+ARNGKn6FbPEsxxwjVJRnAZAObZtOliN7wbzcvrttgXDK
Vx4XJn/MJbp+HfeHZRwDK4m0GdQ+6jhfEUOlnBrxGNFu/ChxlVLm8fixHQz6
1kSTpSzwyacyW5e76C+OVh5spQZgg9m1P/zDs2asHZE4eeMwumqgXee6D1oo
Qn35Oel8UmDuPCmcLUmxNKc+6m4Xhaxs8IdMgUIu7DzMu4PGzwz7j7tRU+RA
JYce00OY0XW7NzB8tef+flmjCZzL/kTv1sgO9pv4mNSW335cFYayL5SaYnMI
2wzyD//LeZQmoeIjHVEq0brPgq2XWAoqknecNKGm7m1JRbd9SaSMAimHEAqZ
df5XZw0ZDm2jlRSke52LDOVwFBu2GolPGlnedKWERRP7ImsfPK2ASFTv3jCt
v/+V4Twm323kaRT92D33KbrhpsllEV9fZYbaiZ+NVgiVM5WySX+2CB7YXSTN
hj1MCQDxSjMF+5h49zgbCL8wyq29hFf3Nun5qFb3y0h/sduzpGPihLEk5Op1
iJpyiO23YibGXd0e6oD/V8ZzT+MPAUNuqqhVOIdLHHpndSzSIEoOg8iNjjPE
QqM9TN91b9Xti4RZpGZ7fvwCkxsfQ/xG5IYSSyCaJ8VQfSk7tqWKQln+ujnZ
nDkkM3Wwe2uaAhgdNigJp23UmtGLN22DK9OCJwTSlyDndwqLYBToZrCm276C
KIZDzjqJBXda0rzqHPs9MWKqjrqZpMvTM80/uWU3TuRE4gR0HhM5llxJvaWl
x4l1SaJskqQRF7K5ODsYbWv6/3+7evgXCVm9wa9o0zxp51lrFcMho1AUvjWS
oxQtGE1YFUyjTui4nDR+pJOKtXISjgmuZOOiDFy6p/C4UZI2DkxF2HXcu8LI
3EF9jAclfQvBo9R229+qJrPZoArsKClKhQM2P82JIyVmzHnByC3y7kIAoDnt
rO7ZjlRGCEH8SQxkSWbW6cZdC6Wvl6JBPk1hSmx/l5EUV/ky/Vcu2zkTr6HS
X7bNWYiZjGinXyVStZ4DAKWn8r6L45lkiiCSdbOy1SV70alHRMjUs8eQBqMX
McWZOaTzxM17kWN7GT5hkTP1QXUI8WixyXy+eYt93u9AWqGhg69nf1MWhs03
qqgjdmLoHRgUzoaqKJ5VVl0ZE+CzYR2xA6+Ti0ymTGnbVnVlktCJqSz/OLo4
4duwU1rhCT4XrJiXCOx9vFbf5t5Ktult/yidcH5fiAG60ldPFpG2Be+BBbKb
8TAQueVDk0Urbiz9GOVnZJUTRTao8WyZJe5/GaDZNbCcE5AUkKlMiiT6HcJE
DxoHGk/k/alS+zp7KxC4KwwbBux119qnaFKsrBS9CuSy/6bAHydb8ET9vk/X
ZypIOPV7/HpDzesX6gbLfeSYBSETd3WXvtYHNWFfD4ONi5QL10MGFIXZt6vF
Iv53IulsCU+q96DOkDXwrdoBcrgP21kBjwEvwV0I0fqVhhobNFuvjEsIPjAz
9ydAJ5sZvfiNLk7crYZV2vPAEr0rgUDyCykXmPtYFVZTJP1iFENB+rx5vuTV
JA5DE3i6814qduQxPVyb/hxVD1xUoELcskiq37lWpenP2k3415Pwb9rtLFyL
pU9KhSExuWcBBQ7MbWA0gcDyY+lf8DHhTCr7EoWRQmtzSd2hxVeE2tgutB5u
GnUEIAcH8SSi85GFRDQ5znCCRkYlKyTo6zuiPZF07ov8MUQC+DI4Ym72TEM4
3sbI+nS5FcRnDuBU/H+/cnx66HYc5ifYa6f/UA59+LbYvhNbtRkNuHPTwqr8
aOQvyQJ5c5/8UBXJ9idtpJ9asidfduJvSAE9SxQUvLbb1dHNBM9xIs59YUNc
U/OVB4NFOVbmS4dODtNpZ+O15ObOujzoAS8COkmXrnbmssbgAr2OiwCJ8UYf
I1w+MM2elTL1Q34t/UUh6J/IgzBEDaBH5H/ZvP36fYwRbcA9KixjKpxBQAgz
ZPvIj9NmY15aZXdsoxNw/sRKEDcEkOBh9Vu8/ZGg02DDNd0ZE0w/+n57OMOo
hiE7Qtcvcp3U14wzNyMeGiA3/DCzhRPC01JpnCfwmv/RcVlqvGhF1/HlHkhP
wwMnFfUKmw5HKlozvi8MxjkBPTWeeYdtckIXrQPbU6BOZIss5TMsp+pmXMmE
AQkN8i0hWtJM+KSUBjuNpN7sVEvLp1Hp4Ws51f9MKAQZzDtrQ8DDWrqCF067
sKr9Dz9uXxds2+jHTUXOFk5bIaaOm0VyiJYHmC0yAFkL9lOlEp8tPAwHVaCG
9iyscaF1eJx9VWew/vnpFR0qw/sKGs//3g/eI4ZfUhvarg3VoWA/auy18Zd2
xtqCaCh1NNtcaKZF9JkJ3/Q4VK2V/i5mt5+W6n0CZRH90NMBsaTk42cllatW
9y5dNIkSA/Ta9NgKY6yS2OfQgLODKXuwQnGmxnh+UrRVaSYJeR5zM0QYHtmB
25pn/xzv++B1cWBxGP9xEOpz8CcYrc71qCeffCo2Fw+GBE6K98LEty+RPPQe
BefSrOOSEluu8db2gVHcO9R9EkFCnNnxgyqmhyF4PNTh7LVWzcC6NU66lHsr
IjuEEqASQ3BvjlBrQg5Z5wT8/XxdihX4Agj+PyroyWVyJxikq6VOeLifSXO4
9yRzbfqH7+1kmRR/H/e5BUeHLLwlxX3ovfhtyZJ6PfnRwxdEiLR4DnDavZCp
VGanUC+gRF2GydC/mgMsnuobBoj60GP8c1Xj0Jo+Qw4vEXb7OCETNLLeFige
vD5GLvIbBP6FwTbkBXf9b5mm1yGX6P6BnBXWWEN75HeeRSoromjdaV+ghY69
jmzY9zPpjUiNsF5i7Pig6cLIHNMoA3ekSWcAjT6XWPvQSe3dLbP5wTHMAQV5
LZ/Dxsfi34ZjUwb+EISHDutfuOGJiRPFh0e6MhKzD4SXFFdiY8PumkTzin68
wQmbmcWyV8ZyzwUB+vL5VjL7oqW2N0I6qet4c6ssFa4bUS4LyoihwI3IW9QR
TeQr5ev7Sb6QqGHzJiJ1r/+GoiC6BuoFVQk5RWZ2i6cF/gcyzm6JPR197fcD
rLhSsImTOsbrxZauVEkhZkvaalIBr2KqktpcZu8xfsGP59NECU9Mtv5OZThm
7uPTOoFaLHHDzrBgr8VWc1V71uGDde6U82pO0t9B52OC6pv4JE5wvBpJWRQT
2yXlBII0KTW3jBeTDVunGuVWMkuViocwM/SPs5+JiGBuReMwc9yFG1pyZGlF
lU72yYrYg+JDvOV1cY7iXzswPxTu9y7rJNivtJ/mxryRKT/D2oZ1l3w9E9Qf
eC7Na7tljKUevd5gxZNMv9NG778bjzFxwqsp6X6Cwqffii/ghGdtIXcMZgcT
owbamql8F0+CxlOc5/yfBn+1L/YBDv9dXw9N2iQ8DB/Z5yz7zOvdgc5M5PYR
TWbcLKGrqQErpojDrkA9w8a5G20x6mqRo8ytRtB7gcdjtX8iKrTFcNKvcxrs
PTeaDpriY4qYiG8+Wrj8wvRxdfJDPjZEmDgzfF6mxpsnGLYU/PV6iS45qgkq
eHDEO1ZACaJH4g7Irh1DlNst80qjCtOKt40M4EmK61I+cON0TwXnnfqF2f52
n1bnTp3PIA2jURwnWodLIXhlzcvFAHDUQqeg7tZeZzSzSLevX1LRN2nx9y3j
2etwUrwWl6B+0g7SVu9dOpGtDStEcTu4LO4kIk6stxBcpTwmqW37uWEQ8/wU
i+wrWBEjHTZJE/ELgYm9tuBerOgXTnx80IypEmO64ADlDsorS94gcm+qMQnp
TGg4U1CUVfoiCnm8faQbMKCWT0b0+ihTSNACsCQqsdoa4L9dfzQtKtsK2YBX
0NDRTEZRYRVA8GmawBGjBPKNuI8s5S/wwVlvZWoOBUuOlJBG4gR2y8wOzc20
KxSOWnrcZFwD7RyzaqPFFO1TFaNUCR8DMfDrkQLUMgAFEs9fCJib+bV2eAzd
thIKLgwC1ZPW38UrR+GaRGfPn1L4/4fBcbpLJ1jXFWB/dEI9KqP+3e5V+rB0
yeN99+zEkWxhqdUA4zMWXs+0KEJC0MiWAT4g+o0w2iKftCIAGilyX1YN9PGb
3PFc+3yBmRKMjWEuR1+f+M2JA229YWf5+1q2cxGUwmFf4wetm+GBrUyZTZsp
z0NTvmEo7K6yU6ryY3J6Evbjm0enwxFhjjl1k87GupE93qlkLFVS/I7a7BAT
PiF6o1cwsarIzBQG5YEO9270gGgMNt5sANoUiEtizC1T135P8ku2SpDruFP+
qiJ1t2BzAquJF6JV/cR5uZIK5Fx1GDYKmhypAOfkUgv+x3LOWj0T7KjLN5Tm
sZr3KEQOJB6IJyd65BBUk6gD2zo7S5SvVoFCeXdHV30KpvbqtUec+64bwMKf
yOO2kjFXC2d06Dvt8vrt2CdROEkmKkgPQ20AUtOSv4080ShigNdleigjt3Kv
055sM1QGIiJ7OyLbaIQfuYey7TX3lB+DVmlH46sLGbs4pXGnqI8LgOTSsUN4
D1HRibIq94IfBEmvTZMzLbltZQUay05Hk+6AdPrwzgtcTw7iarSE/W/wnRxR
X4yIK4Ta83zpjmT24kxb0hLD3nPqyMNhvz+tubpR8jjAQdcTXhHcpuOcLPCH
SMeMz7kEQqTuA1h4KS8yT0dodvWERjJ0qyHM2kORKraMmNPFoU3kNBvbZtlr
yChOO1m/82EBSsnUVqm8UHsC9AhPnxbYV1WSoXDlcgwAn3Di5xuIoi8JPXjm
SzRR9kA1F6Qq0YTejEo8P8f6hAeR4ohuzlbw/Ve8JMdTgdhdBx5WVUWQuh/J
oOnN/vNrFO6f75UoKprG9/05cP9zlKrQHkhH/MytXBI2zZraEWeAlZqEj0He
XvrEGLyEUGaW/berpOUc/tmw48YVHbCSFdfKnIExdcSdGx8Ruf+1djqgvP01
ZtQ0MhsUB9lmlSo2pwg/tHd0j05UqMcFcdRtvUvbn4Mtq1c1KJXPZdhNKhR5
YuUl0PwIuP0e09f4pQA2PPKKvSQYgKIKcgEO4pbLvLl/jMs25VQsdpjW6lIu
J/XXcmjHstYxBOuBNi+idf+XzlYO8c8qUSDwixnjiGOmsj0MleG6gWs01Biz
yW8Cjb9EiqRYVkTm4QSwKZT5ji2O7Xi9OJJIpkn6iPWjee6Q063yPN0YTklH
fWIFYeX7D2rIYjdo0/z/uEp4SQbM1yiHkmwf5bB4v8u+6LGuIOY27sJ/cwFi
hewJfecqPHK9kTVQebcwqY6zvMK+8JaVE4OWJCDqrEK2eZj0g+YTZgP76dXp
C99r6tIdmZeQJ8Bje2IXlEefh/GmZTz+5LlXpL5YTu2u8n8GL572OHN42qkn
0EQ3Z4yNmMvToc5I84bJl4atbRNiSg4t5doTfuXxURQdZJ7ypsnrz7XZVCQj
ciRlxAZn6JrPsRd4YdhJY4YIWp7xdTtrjV89g1elZo5ZVkTTriJIGztv7YNY
3hJuhI4rdUuQLIq6PWLHvRm1BSngdbvhuZQSh1Q/CRs4qIPiiqPjihFL8svn
x6WP73WvZw9WVKarBBFSXeqMcgq2mf7CZ90H+zRXt8ShCwlefLFFe1QLoAXp
ds2Bdk7iS6LVWwthPUn7njV6Y0zKnlerx8cXq/mfnvMtZ/cyuvIsDPxYY5ZP
3f6rqiypeY9+cj9tk4Hqqf5jq1BOS4XCIt72OrEJH4m5KnVOv35iyMjvMBfI
SMaqDvw2k/JTdIoMoZ0wAMbOUZ8HxlsEy3omNS54mxzLK6JBTXnO0QQvI6aY
Todh2nslbr3RTF7JT/6Dnkb96AYeSsUH9OiBgh1i+u5kmbpPjnV9CmV5fJ98
0zAHxDXlZPrvspxmag6txZj4PQMdRZWtqBsWrZhU4ePwQ/Uiu3c1FiJH+byY
NekAhsazy39F7BMiJEoEVlTRZI94mU40MMnfCuLQR++hWLDenmuQWqcOjl2B
DNBGNcYO43O4s9n98PkpHZo/wfWTTqGKsbiMWZhmm9BIxA65cZHHiYw8wJfC
dLUaVmYDu3uZmRk/HPwWbwBog54QBVdJWcBgCK/OKHGA0loGjSFdKEUa9/96
Hld59+zs0RtPqsqMl3xDqat/X1NktHuoAjnQyUX5MgQaMS/OOwOYUv0Z3dMM
ElpNAhufSwECT78Mtmd9GSnb1L26vwkITfvD8iWDGGY6K/Ee7M0IxZzealvl
psFJfmt9T0cJkXa9PH4P+hQIbMwUJn8q6uT4wb7W19WY/mDLQfoETEhnxcCJ
4YOZdnpwTafynoflKH+DyeqIAOQESnDvKStP0NKvxdbjjViKjS/buFEkkSIb
+CWIRp5s6qlVul+Dr+hmKJoaAzKxf1n/vttcWGMkXRtbVRzVfO4or0NyAe2f
v2yO9Eqk6Q2lfcJ6FOIb1LWaREBaWynuZ5pM0pG4zpQ5c5jWZvx9n+VKPr8q
eBlmqwJij/z+87SjDpH07daIPAEcuYFhQY2aF5J7Jtd/pSdTTsjKOZBZio0G
4GAjp3UCQyJdvroBoh99oYGRnQZxxRZkIzNrGcnZsJCMI3eVHiZQ8vandQ5/
T2HOhIoU4dAzEn0AW5/gDiNzFoOh+JhFmTcLPpwS/Yn4s1188RJ7W+B09cqu
15G9XV9ADfz+Q6Vgbf3TpMGyWrwe462FZyZppTUlLJKISnCIgADOTiKc5zgg
fGcyCusRX/RetAPPFQjVJ01iAh4HjEjORzIP3ky6mKzBT1L0YGrwsgbMEE7Q
HpCD5UagYFNQx7QTYFZsuYIBxObX1Z2H0jODUwYkZpVk9QzCHG7vmSlwXk3A
gRu3pmXfZgvu+yWnNlAsPWO3N+YY0Rx7Csogz69GO3VmmqqW5OAE3/iP3I55
/Fl2b0NoIFIjq0kR6iFEVJFTlUnaOA+zYj6UiW0aSPWTSSqyZIh0/smaiFZQ
KAj/V+zkxt1eHi+c3/d+2sIJ0BCl4bFbOhkt84WsWTWobWUJG2kR+w4z5Rsi
OHOB0v4gaNy+lKtmgApluxaMh9NU0ylXDzye5ylgnHsxLi96orR/ey5P05bK
bsxnmy+aDiGxZktiRxDkIjDpAekibZa7IE/phYlYYxyjL9n+9Vnu2sD3trlZ
fFiFupkkI71fblio0I5v4gH2SWhHJp/d5uHni+MOICLxb9u6e3pPb4vqgaLt
mTf3KQP2xiaO3HokJn/G3VK6N+pLe72QByK333CIA3rEJrH965agH/Mz2PHQ
LHz3MAYuEk4EZWTYqKex/+N2DdohAhdyNjQbdZaKBBQwAOjrvq/kZOBLS/Rl
hf91zG9IGzEDRgHd62r2oPjhzBxgnQTW1RL0mHgBjo5QNBP9Znq8ftm3ujBm
Sl/2a3+0cGdm50Vk1A6kOmm0qOGV7MpcCaJEZIlew/R1DtphrM0zWS9eNdE0
epEhoLVG237NamkgHYt5vyA/96CWYJyN2kFj2SY4M3t0UizLNLFctj4PrBjT
hrnM6v/Igyhc2aN7sx9SF6j3ZuS9h2I4VMS6554hR4+YDUSHVC5biPrhWkSO
SGC0VsyVF4rO0dw2lZfHNO7+ydzRDoCYDMLIhXeaW5+l1kID3J9gtXnIKpKN
C9JXPmifenOWmhnfDk+URsmeydeSH5Z8C14zvT2iy3ASJqUvBjm6/sIeJ9Ab
yuRA4YyTukhRB1jc+BVADpU8Sr4N9bZUyxBWhOhRHYYk3phBRupBhX5BEyJj
SDSrB6T5gMIAw8xEx6yv8tWl+pxTMLL/5GTKOvxg4Oye/kNmV9dLzgedDDlZ
EkXiHgv+NaX0bHOR4K0ONbOk3aEo9+VyEpUDOuKRH9Cj4s2hRTgfAnSin37K
WbJ64FNpPu8GY6WISTNAuj05ZL5s/QL6Ib2IcPewyGA3+iodE20KGaHuUQdF
qOgDK+d1tlbxvslSUEPxSAuxNXL69n6PC1FQsNEY6lbrvfCNMM2+wg7d/T+R
sXF0FduaqkbDScknlDVsxbf8IsqLQxtBTbCxym8Umy7mnKnpb32TVT5qEE9N
iBhujJ5hKVjtbYyhjYSgUSP65YX8gQ8kHfGnj7hoI2HBVJaby6VsK2OiGWIC
w5yUs6GgkzeqMqmNfXJq4a6iW35kVFrLZzA1GsR+HTGJxPvzASZ3S77z0tRq
WSz0d+fq5s19JUYq3AQ1zdgl5dXKPIg6ssbj3Ad5XlQ4hsg8UzOXT/RmtoQ1
T+kqx7rcatfpOGUxgzqrFUheWeUBY/EaP9/MbReiCUHf7zOVfysugqsfxFiL
I5tN8OpCqYcDa7aQPD8QDikAcFxjF9MHtjjbVj/vI0TEEWyfPJj1KSnsyfm3
CXL8qBgDStF1qa3gR7B3Owh1kK8lMqX7Opg9Jo+G8XMxWNT8xVr5u3FwTeEQ
0+J+o6etN3pfeby2HrlRPuRpPUlMPZigg/7eRtG71vbURa3kOFhGAwh/nHm7
22RkKyAi4AoHXxhmHdpHtZjnjYDFJoh3abuE4acDozGIDEJc4WS26TjVQPJV
oo8ggO2VSgvthe7mAwcoH127lBg8dDOAHULV7YwmHZ8a0DuzeOZL36APTCBq
d7pXPTQulUblMaRAmgISqUjT2UF4WeGQgsUobp0oEn9BmoedpYEFSIXr7hVm
91lwh9Yj0DVhbVA69rggc07oMNSDDenlY/c9WWwemfdwjjCyprA/PeoZJhoe
/HZMUitztwmsjnys1ukvzpUsyzfIRrQDXERucEon3MydbLWXuSmHimaweDoF
T6jTa+tiBhOvKK16CYhtP8p+u8C9KMqFJR/ofItff/ErTKzGZ/4IJaaCOj1w
bFAk4TxaqQFozBzQ8X92KaLWyvcjLI+iZHtT18uYPPJE+ixBr5OIU8kgHSL+
8Yk7+mI7jX+Kucay4hBeXU8YPkeYdy3mfZfgtkcBNSv5SjWQQVB29BkPmgQk
bHyQTR72FMIHht8W9qVV+8Rvlb7w+QpMQYSOoKexP1WfEai0pxqZcnLFzmu6
DzYvo3zojGgxIHjdJZAKswK0v/Msoqo7X5G21imAQL5Iun9yulemIz5Z4S1y
UbrxdOkUMqb+h817CpIOLkSKGGWTVoExvFn81Y9HBmh6axGbqo4uWbW+y0Mf
WG7TtbMwRz3tmbodZmqLnWzwvieBcC5GLMJwqVoTGX5J27UJFUxNjhBjlAPW
0CU/LqF6g3B+CWv2f/nnT/yCHNglrupV4YZ2xkhSl9WJp3A1ieHVQlDKG+ll
JtyNpcnXJe0H6B58q+d0j94x6SbGluqgrkkxpxhPP9dOQqum685HZPihhGD+
iweOMoLg7a8laABI6BVZQvS5Q3mZn6HXfXduwFcKcQv0D1RZo5uLATypoUBR
uaFVazsUF1CCsvliLejxNFzsodGKpfBljqaE5gU5IqCIwkdWDYLJr38QonVU
vht8uQ8ygLiEJWEVhNSt7xlXiMb89//RxeUzqcNicZ87jvlJn7buNtZ3kk+9
bZl3Z8G7seGPYO6fDuCybuhT8MAAlCgkeyv0LlOPx2N9n+BE6DHVJASCXOVS
ktOqxrSsEEEp7zkEDo/BaWejRetFWEDxn8ifizinKRE9I3WTFjLzddS68uT1
o4UrC4l0JYdJSNthQGnFULY8N8SFQt7tN2QWGQP+XDyiZHW36GDo+WOdJAwC
zj1cOGd3n7y0CNRquxP/AkJi7tET4shp12EQwnc4jRP1aLfOAuxhLNx+3DU2
3iUobGg8GKnWsw6jpUKeiDsmwHfDuMKKr+s54Bjr77Si8mUgxMoWopuqrwZ2
LUl8KCYf9QNg6SI0P8RnR5vajfn6CYz31xBKHudAERRWnE10l8jfjcO2WvkI
vpDWQC46IaVvU5yHp5wFoqzKbwJ8ue4LMwLQw3n0S9PQUrmlJB4vvnzZ3q7o
7kP1CMhTZSEENkDxptgaZsx/VJHM/3f3ZWVAaHZcdWaiDxwz4h+9awUstrAk
RpP9FElbUDm/esLrGfNT9X7VosX+BQ5SQw+lNJvQWSDKne1RNQS4i7EDZw2u
dHU3tkUVhqkYy1oD16rPY9JaMdKsRSSuZ0T2n5gYOoTzzCxNIr5w58awyj1l
7e/7rQsMgpnEtKyxuxv434P7Ortg4s8J5tn1H8b6wt9/G1qN/SriBV08NgvX
kLzbJPUr/bgDAWT098UPGVNZmWbAle+1CnsRCSHA+Ya+piD7TYGYR/2DcKvd
TL7+O+NOWNKmtHl7ehj+ALhXXcAvwjy/y4Dz7I/crtj1tBjSgUIIztiEaxAI
kQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyL0RwoYu3ZHgc3in4UxOmmL9gzWyIsEGT5Ma2r/DnVHgVTAq4VOqvg44/YCrs9j4CcbLpxuB2YiGYFrVr78KTv82oraZye2npkH64/GfWzpatNrGP4Ag6J7TaUDjPMha2Aj3miRceRWiqvjeC54wsdR7XzIaffLKVPr5KGzgiv2W/vXW+SHDmpR1Uksz4zdz/P+Rbi9V5ukmgwi4qaKunOlut5Cppj34c0v5MkqNO6ZNiR7UYl09FNlZujPsASBF5GLaalCePuaWXWb7H4M7E/1CYSwfcYFWSRGtpB3STRA5x8WTvbKzi1/8toF60N2MdoR0QS8P8RfPSGEmUzEPcCj5dj2MI9u5O2EOor2KVy41/iRcB0m93+O1E/M7mLEtwj2EN8nEOgOgc8XzqBzBoMszCH8r1XKAbSGT9hntHxHuj8auDcOnPEU/tyeVOQEZS7/Opu2L/nIiU3YVl5QCffIZrdfNc7yML3URWfK9nwD18M/pEg3woEJ4CnKJ+NubmHoT355drXf1iV2MWeBwA4cQXqf144WX4rUuUPkmUzIbxt4Yv9r8ArEq/iLwYNBpP907iWsgMhAES6hHQ4xLx9p/QQwBzZpxtp3oTszztFzgbFEIuxXAiwWGI/OS7l8l9TKWzViAqSrBA2Mfmr4T/1j/l1hFewWpwWLVgfgP8UvIxRz/sYythx8ZZjMOO+2uuF8Sf8aCqHQucrsz+81MgMYivBA/9nHasfSutVIfdInK8jHsIgh8vTZs0nH3BgmlSYdfzain1kWosALr3uMt8Gz"
`endif