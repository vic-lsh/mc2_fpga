// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aP3Jg5fW63ZPtjwgY6TSzFYzzOavLDZHGsQJi7LxOcKooHD5fSjhs75IhZY3
YzG3TQIMzij4HjWZ1XItlNDVf2HFPXlUul9rXEL9CY7xIs7vSzy+v2REBNJY
0E69uP7AeSAXajlX0McBovFyjIpaCbt5oQYm1GpJ5nYFMe5fBonmN8PbygGv
sf2O7FGi+m7kaDgXIT5yDW95yK1E3MwgPaI8GUF2WIU6TSD1gy7RDXcisTH2
FWlTUIp2K042HgKCgkk9J6vBwD/jDjRALK7+gw1fZZ9ltP/iahc3w6c94SBs
JasEiMjAwfEk3zN0q3spJhd92FKIx96D7Vwarbm7fw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HhU/OjgetK/VKLfC9rs6g3X6cKftp2cl9p7uiK0hWRS2tGCucdBmeofZS1wc
WFLrGEJQkWr3NRgMNuLo/TiXmHAc7jfF244rXHSq2nncSXWMQmPt/k7+zx8v
rAMWWQl8VexdNM0Q58fiULRG8NNZuE0/JkEi0K1QAtJ55qWljHZvCNKBlwHw
p9989910D4kajuYbG2jo8z03pVcQP5tPbaOnKaNjPwKNzXar2iUZrPC0Unqu
idmRskd1VV+KpfpEfSQFLv5uDv8UeTXns1oGMWPwzTTfyiYduyZPRGYORMmO
bcCF9gVbVkmzgzGSEtdntPDA6/KrRaiMeoNPO1UNOg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Cps1HUqCVWWHg7aik5asajPiT0tgX0ZXRmHg/RYf9SC22L3x1SicaWUOXp7P
owfIXvwKwAhACvwzGoRzbXtKfL1u3m108EDt2aknmsH9BRscFMaU6QCwvF+x
LuyJNEfMtX5m5TaMBQY3TOauwkcjNAJRys6NfYTTlL/VU3UWXHgcRQvq+Rx4
ts4ChQro5xfHj5WxWFEZ+O5zRl/q702SO55j+2KwAO6Cd/jI8bGx6rJgs+H9
MXDc70mqDa/YWIbbVxAHHPlmk7NmX0n3ltZF66bqOGuvuvt+EvtReQ7JePMn
WIQ3T2RuWNO1owmCZhZK+/5eiNaNtIIJvaAssrvw+A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ElGP8n3/cl+5m5hqlYW6GlDljwLj8PqB5GGi+PEN9DmnU4r8Ib2gsBshLVO0
IY1VPX6PHLButxTVFgHLZdY/DzRvXQKfPbpAOte1O1CebpehbP7nv0lmVujB
z6qnAuAHnZLbYXOh76aeBmf1vlECVqntB46F+RkZUMIdfW4jXYyBBiMUy73N
HLRStPEVHPFLwVhXFIjUrfZHXE+FiWoKCwSY1iwS33ocambvL5xaQysRG7W5
cJCE/bfU6Fx+yQLYigQ3EOrChHYIFhle60TOWkzxevACRpy8TVIXMlX1fiBc
gjyo+/TADRwkhdBJXHNtBHCU2rD8SQSKFKgvZuZZeQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fMMp656yWaGe0FTV8Bk84ALucP2olcAe9Jvon7YycocZFnau73W20iulP0ep
2p64c0VwThRjpN6Cx1WuV9Vpie27xwC7p+rgzp+g4gB5nFVGCb5nLZs1Js/8
4U+63HQQ6fp8CNy4SP5nwqUI5eY8bsPeGQci+255WvqPeiZkgkQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
dajKIP3eqA+ceGc+5LzkpQVMtzXIjXYTwCzL42vVn8n/ymXPV9RiKtGLPC+4
qgXBd+I+UjxGly0p9526in8R0NAOWCiZ/McaIMpjbiKSe/hoZc6WhDXtWvQK
zhVBOHhHJdal1LDx8fBIlktHLkRifpvI/oyC5KJwNfn8VnxWw62O32Hb/5Kf
LhyZYPGW7HO2ZrrReWXrx9TePRGraPL6h3pt3RBtN2OU0YZcwdHZMIv36fzl
HVgtuA220fCVENoCuAr856lR9gB5Og7K+tDo/k7dt/AmHcXTfxlKiA/0Xkm7
LcqKrfi69UN3qxXVHPmcIFk8pKVqgatmsiGLzDqRsUyNj9KxT7g1WJ0KPi+0
oqLmAXYy9LEkWr3boWbuULlJnJZKa//wePycmOJ3R3At65mPDjanZG64asT3
QhVEBZvYOQ1dv6uI9d86uHuKrP8ISlVwjHVUfzMTmMDfLVSrrJZBtBe7PEsg
tBT5IetwArbulb2yUD71J9bL/lc4KE6o


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fUVtR2kXSHiQxVmvwPq7B2MCGWNe8l76P/ZU0aYh4Pu8Oz6O9qy9cR96O0Hm
b7WOKsYunRLwgw4By0zvCMNKCghcd4hNqWapQe35ql1Z5PfLw5ZEOr4pqfHn
vYCnhVUuk9zbIibEHrt7kCtZdyi86sOoeY2YclMAPbMxisA29gY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
a4SHLhd4dw9OHm7XYDwMu4tPv6ol2cbJxR0CaWFucSE0ofOl7Zn7pRKFHy1k
b5SN+sJDbwFIFxlkcWOwHoP0ovRDXeixMs7rd0/fPXxDDqDpHXmRdFnqLzza
WkTJS7smjNZSUqWN9qokSo4DfCvBb0AAS2MYvYpm3NnC/3nYd0c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
iMmhpdMjbZM+fdJ8jDpad4E/JnMRoTgNzwu3cKQJwvotoQgWhzxNcjopneOG
8iQu+RnL2L5rT0RQheI53O1WFqoAwkqVti/+tOa8kunwy5KU+FEY0QhTu2i9
uozcti3dsEi0dNb6/qbf8vD/2hpDxb0hwhlX+3xEU1ePZ/qbmDILuOPaYj/x
zLz7+XPzbVIfYG6NmJDdRdVNjv8aIRO+XDb7saB2I6us4lchtkfF10aASFCr
fQtUf/8qGO/neFPxS2iRGTgcX/LvtWoYYesyQtEbLQHTFwBbNJWsxC8yEHo7
w5proqT6EsHyP4F8UXgs0UTqxuio3cJwZE+dSeK1dRhYnumbpPMfN8PAuvet
t3fcuHLekfjgwWZvuQrHqWff6YdlYR9/f0/EyFJnKHM1Mvz1uL9rU+gI4sKC
iyf+8KDy1Mm7rV/4dw2xzKTzIRuir+vK431N9bTIC0nKsqF+fpRtRsSSxxAZ
VGNwtHIGQZOM+7UnXW5P/FivU7VJIV3l4pByIof0dfQVEREpZaKI4BHK01hI
i3jI3FltgjRI9oAngga9DWR+qTqGpPleB1Oo5TL9BDxefUUtIItYEYtFMNXg
zPtS5nn45WqlDAZ2TNAR0LBdcSsEkrU6y34dd/WvStycqosjQuWyo9JzUs5w
DDbCtkNPIFm3netJnGbh41ktx4fmWMa4Wf1TpvjlUi/RdyN5gAfTaGGqrEQP
Ykb3UCvmZWxOlgLVSkEx0uowI5Phnz8Vq0ZzkSRA1jSTnyVpefqGVokiZlny
BkPxQ83o2gQUi1gkqp/KudAbrmw6KNrnnFJInC8218QNnTpEqFqpkhWLdGa+
uxHJQM4/pJLhe1Q6xB5KAp0nGxCjbl/zm9m6S7ft3Dy4XKKOIK1Xc6Eq2NqV
F90W9aAYXQrVKfqRjVnnDVRrBqatN3t2ke60COzny+68vNtKpDnTV0+kCkmI
ANJJrFoaXJlUuCKypDaK86cBqIqrQkxg1HuP7xCt9UZhdF93/7CY8pOiledA
NeCKZM2rAaEFHFfxk+vbfu2p0qbEvQFS+N7oYomPXIHFcMEeoL/xJZv9KPVc
NKCsTaIMCD1O1JPtBKvM7n35hg49gneSh+I9y31f75KwXnOPREFOskI+fLGz
HHlbS1nOUxNQ4U8ZV2frESsLU5FvQ9K6RU9wG10otTF5W+Dj6u+c9hB6XUyM
MKHnc+41NhF5qvkifL1gIP29JH7TUO/IDfMHQzIla4ON+RrmEMnbzawe2NKK
U2fnNZbsvxv+FD6UHVt/KNGGrilebzGgdidS26YDutXyT71nUstySQYXAxub
E8UoeFRbsSjEoN7FqrGGterod4nstm4z9XfnDQsee3VTzK83rDXaoCviSniM
7dSF661XfcVA2Q4K/0AmsmzhCFpbtg3R1SHrH9CngZhB5vElbY/IQ4Pq/YGc
0rswOEmkFQOEcXXM3nPCdA5x37YavSjxPvS1IyHHGVPXlem0LQTNpaRkanTT
1X/e1KbTJxBKfZvm1HAR/Pvg+pAfxTFExSlyrSSyeMfdGBB2jkLEx2ZmGDKF
FMitvx2cm44tYlVvvOafh2dvKBKCTejgxQp4uE6SgDhYbSPmUV2P0PkmboXB
sFIeviUQTsPOp9cE9L8SE2NK7CMfM4p8iYdmHQMH+YCQtXvpQKi7WECRtyKX
s9in51QIYQQhFjC7ZJ+vxjXspGY90X6+Jm0vqMVDK33blgazDrClTXMBpM5H
+4UMlW69Mw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoyN/OX96gu34/6BcAcZCBR29W54LoPUnbY6ao1T7EJcy36Fm8jreuLMrGUTYcOB8X1xKTQVEAY8G+dkOwZ1lKbPUUqZMnxC0NsWaBytLAKM/oiU7xfTKByZFfPO8OKxT2kfZmtbeGJ2XNriZbq8Qqflj1YGQWSR0ZRILp/8OsEEw3GodgW1OVUBjJMlP7t7uNZyDQdmVy4VFhFZpRNtCCtVkf9lLwDpyx4BimSmAkL8ufI/lYT9rK//ip0ppJZDbSSP0+vYmLmQiDGZYPaMZOJS2h+C2YcDgfngQ+BWpi1WL1zPP6QjbZM1UVwsPwnutA54rKlurOcUC+cWkNRz8Fph2uqHj82xuuopL4lDX33CVhD3KATN42i9B0rAK8BuPFH7ZZoJTEYpZJ2DgQIdN+6uV8+QyaBTFP7TS7oGa//RagETdYm8RADd5H9p+0+uMztKv7K8ZwiKuI07MUCNaI1KEtfreTLbEo5QE4BwPqeh4kFgZmflWNkXrGaHrn2puWvYvLpA8vdwbE8pFe3y8A+F+7ejyuZvOzLiY5OfqN5Y/kb4IkyYeIUJAE6+qGeG1wX2JIWzHa3THD3JjcBqGsk8W4AXDLcJUZze0KyOBAOKMBqxOxpDgq7cFgQnmszhWClrNTuISk5rG9BWiIxwVWSSAlxwbH6nmnOWTUnqiiF5uWDaLLzfzvqjlbGLYIHEK+P/yFh/K+HEEC+S+YgzOdhFqglzHk3xhumkaLqo/yeX8VXyPt/hnsiqh7DZ716xOH9J2YNFylXc7HFs0eqbwWBS"
`endif