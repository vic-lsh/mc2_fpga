// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bRjdFKDEbpAcx2q4yUh//+t4F3hh/ZisAccRfWZBmOyG49ZDrmDwMiLwXJ2o
tLSV6lFX4PQb3gSOJA9Pank64C6Q1qdumxnx1fic8sWPD8Es70xG665ToH0z
NQv/wuXwncy6nLgmKD2cZW32zw5Tjb8yfGgUc2FWplxTAiXvQz9VsMGVdt26
kGzYmj4DUMnEjp3P04+srcpcEdDq842SmTsFfQmL3Ho7ul/CTolT1qCnRP3s
m8/se2O2iGqoZB4HvwlggJrnEsAJOIMeLKUWgdfpXHHfDbZGsVIq7iBo9Sul
awi0F7oVliRhMLdxP4m5W50abDMrzT1naEeB80KcJg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DqDYYDNVtw/0LrLT5nPb4zC2g+motbluvneIGMPMqH9KI5qlvjWEevpiW+l7
SLaq2j9R+R1aqW/fv67GZ/bfpZZaifgANl90KZC26enJtxN6oXUz5Oe20Tu3
iNsSznPysyg/pEiYNSIo5q4Bbl08magc1pgFTYPF549YbT7vabzyHJie5OHK
R31wcO8YetODXHQxeNvlK0pgzNzl9/435rNe+Xz61SVegX5EM40j/ywLzrSg
Ln+ctEXWZV28r5LLF/CnmaVV+mebghFIX2tPEzQz9oTqUaO7umj6qDUGTMQM
0wbEFT0Hw11DnTX+am02Ro1/U+vD6M2LqGDd9tWf+Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nX40m0p/izUyZStDAiMHccE3oXytgP1YxQ5mPfz5zzTQNU0czF/wegZzf7Nx
OftKBdpf1GfKWmu70UotfQ/oYk2om3w/W5BxXfNO6iSe7KHfhod1LR9Y4oWo
f6OVD81p1fh5hVw9wPawgeT34ya92clyWJh248cA7uaZPtx2yKrCryiDDjvj
e/wJTT3v8tk+gRvhTTbPTHrp5pSvapoiyJLcGJyTGzNKpVe4jj7HbKETx3xO
hcRbmf4fu/FyTk06YtkNri0yao0rpFNqSUQiwev+osUddTD/x6l5FspspfaM
jl0Y6a0xqhqMa/CsuMvm8MtFm9CuZHORcDPggVrjXg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aDMiJxzhEVbtYlsTby9ryqVmZpoqlz/tA0sqxT5R8zxCSWHC8aXvEm1XoBRA
1I2Xml86BNer6N5V3WVHiqEevJPQP0VHX3fF2YQB73Ly9vzxZDoem1PymaaV
HUOLp09n3rWcxWy7NUDvxu0XKAYvVLmW1eO6Q2yEbMewr0j446CbNWFFi6Oy
gjHw/+msUaEU87tU2lnxH6q/3cUjDen7enDu2FQXNHcOUz/RtYuQfiRNcYV3
fMY+l5E8TbL9682ruo8RP9EdCIT97yDPmv3RY4yoCELIbE2OmRxxjj4QfoXr
eSCS/88cQJukraHbtH7SmJahQgud53cGILiavpzA4A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K8okRyaHXvDKGv9hMGHnCi2jJ7nhyAhWBupUYyEqMV/eI4US2V9pvyxyuHei
ngPZIQrCq21lLLB9lX1XJ09VVoXE41KotTD5Rlie6KP3gApWX4jRXGXluroL
l0zorSzsksp499zsa3HzUt4U3tYVb5nAgUC0Ro1NN7w7o73vomo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
m/sWagf/VX4FFEJmEmVK8Y4nNc8o5oijDWhIdsoqAhHXLotzHtXDAK+YWM07
06DoTd+ETP8Ooq73OYSJ+WMFLihibu1EQgF7Zka+H3olk0KjUawIFCpoMZm0
Z1ex5HAB42juMBH18qXma4fSY+eCfIH5o/LvoPqWC8cpwoUUh20Z3ieSFEBE
C8oHt29JQetZym4VXYI4mbz/sp7LRhIpNeiFPteAoZT0fEaP8HIGTfpulPo3
CzkNxJc2CM+uWqxPGbGagsoiaCgHFaUV9gzuIRhzEzuNlG/Qb4nGDSxNmOcq
s1PzNf6uyuZnAcxvIT9y2YC000MiUNGyd0sB4a4ddvB6NElmWSBcuJbSNVRC
N+dpL7LOBADEyxKyZGQXV5ILADraGowuTVQ6h1MFcVdjnLRHcnE9iKgR3kGE
jUUSZ77ijzOaIV3yOmBSfX1GRayr2slsmjkTDA2+u/TntIDAPlJkLedr4Pra
17bKT+fNZLb9tdH3NCKDlHkJvDlQ4W7q


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jOmlkZ2oo4OLsjSTZJLuEN5BPgMamKShTr9Oy/HYq3l/u/9MR/18jrgBC306
/taDA4FaXaqFV5XO/X+GlR/X4mCis71UVaiECUCYtGP9d4mzABoB1vrWlOGr
Uwh+CEB+fSorwmTvIYuehKUCv5lyrXYYg9puIVxdiwahYy/a6Pk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GjTj91oZUbwlFpdp4mEvNAOViQiyQZWzhU3pZj8i8I4xHs+1i2CMNUn0Jz/I
ZDeOOhI6cgxFIgDlgo6g5PETWeq+JxGt95tVOv/zFiXexyDQRCnVXD1ZpkbY
oSWKc6to4z/U4s4tDmW7YqjCpZxfr07YfjwbgrCp/llCKpiBecE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46880)
`pragma protect data_block
BijpAO96VWjxky8OqBpos5i0iN/XaZt9SCYFN+poQGy1z1i//cGrHvLN3jWq
TL3wR2eoLnjYPCCs2mP8XDKYBO8/K9r6HasDnLRBpnB8NUkGiwe6oqSH/RvY
Kk874bCNmy6lQESAe6KOZFC4R89bQjg31kCQMkNACO6aqkSid7W++/JG1Swe
jyKvuYT5H5TAeFfxThkAawwxO4bl7L1+Bft/041FPXAjuLU7oYwNmb/OxY6j
/2D9nDsePJ2Y6eDqL/SMFqC99Ckb8/viX8rpugly4KoMq2botlg20JUweK8D
6BS0EQ9MKVpsntWexWCJuPzDOxDKkroAZcuriuU/fYaTJQsAYjDB7Q1TTDIL
Q5YTNlGL9v5eeYhCx+AwPtKli+ACpDzbM7L2uN6LA9rc54qIqqM8+wnBCxQ4
1oTKY9z67vR4r0W7BsZxkC6yz1MADpiuRS2mKHcVNbDPPCPUy6Ig2eqKMFwd
fWLGv75SK1IzHHxM9fbTOruMMF/Oari6KgZ0KzO+6PDHt1B3YR9cDDCP8pkF
lc3pEkAaC5GAm43YVfo7g6LilceEMHeQBQIYJbkkV2qvjRZwIGbZ59Hec8b0
IjusKqd+pZG97+aOR8mjz3nW+sp+nrIxXP07ODA7sWtajZKjBHROGQy73dMj
NxOfHGm+E8ugzlYaiUNvfULW4muHvw+Rhbq+pAyHbb4vieKFmemx4EhHN+yt
V/xvWRMirhjTnUqChszlI9YbRY9BBzXL+gps18jRoh1BaZHaFjMGP1BD/Bme
AdrYrMHqY3buGwO4m1LedBUaoJGwQhgIzEhtOcp5SE5o4pCX693i2gVXKwji
i5RegDGz2Ozc92uzp9+pDGM0n0g8xkp4rhczXFj948XY0XMKjiiLU5xwAn/e
HnWhCxksPIDH2JnRcvsoo5V8L/IYQGe0i/dezxdKhG1PgOQcQTV1deb7b6/1
XESvyw8pfbtU6GmTaW3UhCOgFf5xdzjIlCou5m65ahrYNTfcXCTUCzMwfhzF
4PcbCVSTlwm6mzyMAEx86TvpCplXriMkNpFueRrIDDvicPAjNrEaTXXlMNvG
6hIHfjtHeDj6tWv6jXn2cOsqEeC3INokw4vbo7zoPcc1fP3f170LQpfdpL3h
/xo50cVddh0XNBkwJPsSZ1hMow0lsKdlisIvZ4E4xbN6b1x/Utwc1DtaOP4M
itGM2EAPwEN1NE5WwCmFr8fVY0nVlGDx3HSGtYDTBZuxCIV5eeRbxmwBkYmD
2MVrw9Soipp7qOBhlvjjFxApeB2Kc3YDkwMxiug56cjlt1cBRiOXq9hzmm8m
XaOizB/6ZvChkJZ2XZer+UVWQwlifantWC6D9blpDhSgg+wfatmAHwtpg9Sq
k4NAXXDm7KoOoN2g8Um0uHQxZIS68YRRPrSUk9S+QiPe2u7isMAIiTeIIuFp
EuFnGqcADslw4XceZYfZgOVMG4BPjA/ziy7AseFLZV+2xsn0xelowGMZnKd4
8Xtk6aJwgTbvVvxUHb7hYAgr3OuLr7IEIObgWses4kYC1eVvVaLkQgULX3Ze
9cKpEDghk/eJu3H+TbGkadKtFalgif/Bw/mDgMlmXFW1vZ9HiuEncw3f60ES
cOqnsKiFD6nlNollW8DbqgWQVZO2BTaMvMyw3guwCp/NXmNvRGoY5ivQdUHx
n4jpYR016Mdw+0bkafWCEEYPuxv4aTLgazh9Xb2pV+RGoJNJnrJM9pijG8j6
gST43K5F6bnofQ2USsiRQy1/rfR8JExr+NtalOPCr8rmfBArDhelUE1hPdwM
/XOrNrv42Qi3iGRX5Vpgs0OGc7kurw3NKN+weXuBZ1AEnN9v6F8axrkVr7uX
kJy/ZkBjlrwWwR94rDLBej+ROEWTYdreyK8dCw9wMZFfZq0pUrn8iTm1Tp+j
wEoyrMhs2CLbtqA8bAfp/QiSGL2wnxOR+SuKrym4WJ4ttYtoIbg39uCHT77z
S5ixN/RS1Wcw9LchWS8FQU3fFb3o/iRcq5OjMiCYWYrVYyh9NthNJKHqaKQG
2pvzjmFohzjXd3egGmHc4igw9ide1Bb6n7cVVXJXDnLOfKLA2eA6hvqV628w
Mk6UVRRhXcoCp23l/mqReTsIWxHZjbjqt5OpdE94hQJOm8FOzDCvnAsiMpbj
R9baKTUz+eNZHdRgrpPEXGuyGmU+ZtWFcG3h4rBeh2TkBuUB7OHzGtL3StU3
vuih8uJYnW9WFYyNl0NP+olKA4CP8JLorDKjClGxIjWZ/QbsKM4oX4TI5yxa
NRpG7SVi5Cp3pKkYEqwWabzILLLYGGqLRB56gHfdEIbhygRdTympOP8+iYKd
rVXVEWfvgJEAEc2zF44si3hxWJAOql6MdyrncNdbFP1qHgrx11fbHiMjd4Sr
WinwCc1DD/zUEOtWiJh/p1HZw9Dxz8lKWEBOmmtkMkGYEphU3zHHEdhx3ock
MQtmEJU9hbASrPTd8VwwL8KuonShu6enSR+LtXF6ij//v0xVe24ECxWGs1F0
yR/d5aF768ewbQNG9gX0Rx2NnGvFTZYOxU/8yudS4fzJht14vu+lpejNvx/f
5VGQsD8y5LBh/tw2Mnwasu6IFauY6jIdTAW6gC2HaglmVEkddgCvA7bjocsc
mLMeLCsPGPBEoFpDAjA3vEituyGVQj5vflOj4PCQiwqj89s0gPH4gbNthw+T
mGuc+UhNYwHlQXJkPY/3qNPKgvvGhWsqGFqcPKTf0F3m7+gW2Zev5DgFgYdQ
Fo1WAuEqtENpsytsD1k1NAn0oJJwoJWB7CbofKZiGTccwJN/nUSIkp5xjktv
1rYN/KKVXPfvnK2/udYF+eq3HjhUr/DLextX5zjMpyacXp7NXyTz+a7xNinI
vW0qbIwgEk/icHtHP+Po7IcJNLaHY35WfYMn+X0ijdSsWmOdAHgCBE3p7Fpa
IgXLvhAztl08stn8JF5Pb3hRjZZfO/kVbVLnaWJKztTUKde5iDP/kGJz7Csg
MWvoSvn0IUkMEdXmfe1GaDz2al3omFYhBC6u3kSmJJGjH1kOzTPyoKUcPeYd
ya+YM+LpIBwhRuV54lHV5T/DNDeKYfxiNxkCPy9pPw/MmH3P0U7fdAXm+FG1
t8oEiLLTQga2cq8bAUBNPypEm+r2NGCA8KnJCJLVvUgq6LLWEQ4TsjWrSLK0
TILSZIGZigZW58TEqzbBAKvcLKf7xRgKQln9PaX9niaQUwewjeraE5dSD+Fk
ipq6Ia7rzdP4f/Cz6PMwPVlo2+SgZ7QvZpz2eKNniyBWidKy4IuikgKE65iV
I8RqBT5WWOsYw74MOXc6sfi765PsjhER/G3jrPEbJpodeSQR37ImHxf/XaJl
WHQMnuj7SRG6CcdDjemh3o4gGl4vPsV1Fj5wFusFMQ9D5kN9tDas9XQH3Nzh
xY9P2t2KTpn0MbDjfibAs9IgthEEv2scKL4TBPb0AqTOpuuMnGp+EsUox9U7
wCa4iKzeInUEkd0OFCNxYD5I0rQ43QUTmKOs5ruQkEM+Sxi5gb9btsyojVoZ
RSdp6bekMGMCppMAEX3adi4ztNaXDTdSBeDYPjDOytg/vhLI6N6Do41CtEq9
zprXloLG5wwDh0Vyckz1sn47gvuIZG8Catkw0gfDsr6dP3PQ0p16oi5a+xk2
tEXdEAtka4Sm8VkNTQ2mB61t6+SzY9kAa/kcyueX+Gkgi92H5fAUiSNlJar5
oHch3whJtJHK2mabzAdOZ6JLXnWYodgM+QO5huVj60pEkBG0loAfhyaIb63v
+oC5milf0Ql8EsW1BG1Gp5t2y3yZI/ldKZ3l6AkFJKTRqDdq2FKe1XdRlVjC
d4zrPo3/1u3oB+gsC1CbNIX3aL7eJg11lFLdr8YDQJYcMhDFtW5YNsGJQ0SA
3rCQyeib0OO/rRfwquT0j+WjjzIDEdciF1hbRa09vBmXPlhxMUvNnWEotnEk
XJY8QF1g0pZYKS0dK4Jq+B1BwsBgKsFsh9gSr5moJj6MxSVQhjouMQ6/L8qz
ECrBPsU4j1D7Q+0EGiYJporQqKopeK9X1V4W2Ui48fDx1HXF0mxiEY2+uVuB
I7WJwqjdjhE4PhT73T3dXn/Rcpcl6XXlzPSjr7B/tkOelbnMeD+1BD0rgXNd
PnhAUxJ5vp4h0gagIPJ/azQJ9LlIS2sGpmoaj4fmF3HO3uUaUw7jG9GNGXNu
URYKk3yAqZAmFZFAzqKKQRH64bw0HuHIkV9JHfqBwvfCEpT/8hTYz70PmbsZ
ATy2pr1SIg9yZ68bwF0F1jlzLaqgXibw4Pj4HBzGI+jUyxQKoaB5MM7XSWx7
ajFUe8eeTF/QIZP6L7CvRCSV2Hz0KayTCPqdwlNNcFL4Op90lyTPlz6mK1oa
fsv99W6YbpLKfKtCvlkhm/Vmis8g7F1FCmFtnuFQbgOCrqg6SA9jtBG1Y85r
u3vM64joUIJZswc8uOoxfUPKNVaSP9DUKyv7ouYlZN7tZgKMUIBUiqbQluEV
kELNqBNW2flBiDyFbC6p7dQ5D2cAfgU1545/PMzP34FMwzqOKSQqiN+SBhxT
4YVIiVTQnr8T8ljC5kEKkwEflOKS3+6q+LrdY+S+gbRpAtcGwirEUPgYO5G8
/yGOowTgHy4XHJnwk0qT5Tmxp6DaWmx9EK8pWA86c9vKJf7BFr+aS8W4BHsf
orcjdzaVJaMQwyXzZD9gaQMwGTqZ6iLH1O3HqPj/OSyihaHoHRv5PfqrAS2J
nB5NKpCjttXbFrJE50+18ISYbGrQJeA5jD6RP5SksIY6qnufyYWBtpGHhhiq
KC3uFBFB0RHaEw9AYim0PvuOSvutsgajqMO6HYhSM7iBuvrl8hnwEWKrgS5k
yZqbZc/5i7v7XkoRXJxhOPG40MMZDOY4VZwlaIX7O8acfqstcn6RG5Ekueht
SqUzFOUaK36qVVKn24EXe6RtdSoO7TRO3EU4jUtzrNA7ZUDryuBYZdxYOnYe
t2mUUBOCfkJhSaTFuIeQdkFms9Kk0ZO/7/ovlR8ik/bW3z+67gXQiqPmsH6f
AdnstiTlE5+nbuOwBXqlaSnxWrRwJa/Yd5EOPgYO5B/glypOwTiGqIjxrEJM
JrA4sqsDw4VwgqpRH+tOG8wCQ2Wjjl6fs7Uzo/trg584gOcgaPSSmvayHlRx
h02qN4E+tp5tT/yx6OJTbIoQcbw9GR45wTcI+sbdnYh1IzJtq9tmVRvi4YBx
vRhA74+ce04Loc9XgovadJbkehHQLvyfv8muTTkFjzE34tZaGN9UkA2b1TeC
zZzUas3pwDNID6xZCfrMjBriEB1YBg6pje0x7Fj8FDgWJGdL47BEwBlCq4wU
C5SiS+uKellRpKKv6rRpv+5W6R5MC3iLJdzMzUAss1gbxjnW4iNL3YCWPVma
asIXs41SOPmn2DdXizgaYBjrcIUHpYWEt8f7xUnoTux2y688zdd/GBLEvUcE
Og3mQiWVntkJ6y6CYHCP+5pLYixs/3IVZW5ZVdfIiGNoAtwQdwLU2Lm0xKUP
mTyKVlziScqzBZKS3lyC8QenMeq57rJ9FXAYV2945nufb9KndRwBboeh4zuB
Euy4JmHVlBlTPCcrycDJYtrRyRiIV3NCP+xDYwZL5jhegoXr5ZZrA14INJKf
6DeEDUAbRdXjQ+eDyEcVvH6zel7myg6HgOiGEa7zcRnm2LF6RfKSrvuRa/iM
w2QSuK8acVHDzVbLtMDX6wtunpW/p5r8QCxMM5VIrIUYZ0dEgGQDBl83R1I4
tLjeOld+SuZN/oMYqRcJTVpdmXja1lIvzGWmv4A6OH9PvBchI+e3b4qvsIKN
oC3xiaXef2EovNG3Ktz6ibPPwoLj1oOephjOFBJibpbz/o5fG3AGbDBFbOOQ
brZVfxVcnzaii1W/uK6msVIdtxzZFcViuDW7C3RkXRLT1fqjvkKlhzIQurUb
OEyPQkj9ioNqN6oq1+sM029K6b0QsLw/ZBsnFiMb4kQz0AofH9XmHo80sVRS
tw9Jhk73loRSOV8akybwv/uvNadAEF+stAECR00GBUGUoqwQdQVVWyNVKshV
hZMaVOtAnuqEu/j9hHoTycUznLs6xaarKiu0/bIZbBLPcbEklEn12JuEnEjN
CEmCFtROXy/zxTLXmymwG/GfvxivmZniytnJuDO3k2yyVrnQe7txM8ZA9qPe
YemCh4yyZFNfe1cyDKj3jnSt8OL+6bH/YfnkiTGhYaIJsV3JdGBWTjqU4xii
/VVTywPdjJ1zmzsz/I9z81s3YTRf+TrP9hJ5d5Wu/dfw/A3GoLBZZKXbd+ou
IYCBrBG27S0tYPO44+WQTYbURkfiLxI7ONqGUwuSNkrxiutzs8DCZIvBnzKm
EDXqKRolFHvh3qnXhWbaElrZOKbrAhwAA0dYTx5CvNGvala9wnbulTQp463z
bFj4mp7EVyInVnFVqAn3buZPE/FwmT6ML+rNAeDC8O3t+4fmaRfP5KRDUF5b
TRDl2WS3b0W25GLOqRED/o2pg3kd10ZGia166mIo1EfQi/YB9Q73RLe4g7yN
M2GlYeY4jXN9FIJ06Qgfxt5z1+G/maP6eP5KFnamD1F/NvzDZhpVv9QbgGqo
7P4+eFt1Zrn251PlC9LjpwuehN4AmIFYigZgHFzUMlfFzNB1oLi/jXe7pEej
BOt2x8S+2nEjevCgUMDzLyttG2VpsCWiSar4IDtUrxWteRQIfpqv68qyAnI+
+a5SU5+D3gKY+fvrvZK9AQ8fgZJaPqY7Gb+kRN5oVCw1NESGIbuT8PqNhF9s
9vvRHF0p2CcCt74SKfIxoryeI4pv27k17Eq96sJNOfiIjBlFg53JhoP4l0pW
ZXlyj84TpZUHkT25pAfpYs19Q8ts1zUM5w2uoibXnyWxLPoyP+Qi7Rc2zn7f
6Cg2PXGpLPUaWfbepISfZ2+kqfDMlS/tpIHEfqunbXBOpNSSTGR7N61ERMLs
eeCarffYRXwQlCP/kxqChTTL6vJjawUN+tI6djpTnT80yxREI8ON3n/sTiSQ
2QOA7n/KeXvFjZNB4fwhVFyAHvWvL08CfmDv0VeTDqlIGoQTAGxkbxTTgSCx
Kv5mQuO0KpNx/O18wurT5EXLZrJKBlKsVtd/iN2RKHcJxPkPo8goVodPmrRM
Xkk9oZLxXi6GByCuSzJ1u4dbYBkERC4eEJJeBLN28UqP8KSqy+BzEMVrFpiL
A/J3hMKkt+vOEMr78oKPXbI1j9cNnc9iVfk2USsbrn2fnimTpAp0EUyJLcIH
dN77tVRi8o8THQiMMWvUuB6nf9Ns3lN5ZvEORdDbxRDn5Ue5iAulUOfEyj84
BUY6G7juEuLnfQg5ju7enurcc1rPTQ3Q9pRWxuHEBOx2YzgwjfDZfu9L0aYs
106eInC47BiUYBvsK2t2ZahVqbFgXvzY/kxYH5yctxtP7IE2Br9M09BF306D
Vjt7ncSc04CJjrKcVkZEip8vyfYFjTZ+5a9mgbOKeYES0yj2RFvXev9uwhMD
k6G8gzgYanP6v7GvSrXmUVEeezL0HOq6bjw49yERm+13B1bvc9VHECrsSS33
GyHXFljB2BonZ2xnKNaeHPYDaLXq37UB9xtv4e0JBQNZjc+uVtGy0/VqHkOV
3n77tAO1RK048fBACAhmVw4xZEbfFRYY9upz+BeLRu3u1KTX7kKTO/LmNs9P
/8J3A70VQxhS3EFI567O3qIy90yZybqGz1DRsHSRHfIzl8x5rjIljuAmczlN
2yhny3ugHgQGy5HWS+GuZspZGk1YhQbIwWC5ZzQz2IRSb/LXx+4NLs18UPbS
DzAw25GCzVdxLzETErxtOYLdPIeF+TwNmFgcnDlPuTgHLSJ6IpfmLR3HJLeW
C9rG/967zPQGAfeTiuYbHcz9ENnVdazIRlA+60E0srmH1ctnElR6JZAlCFAo
xIHdjp5bCRC8EAEZysgyQ2q7/GoGKNGqSM3X3UdMcyUEyYT6ZG8+2/Oi5ICk
bw0xBPxlpA4T8BvMeKZlrH/G+5GN1I4DCzTGjqiE6Qx2hHuzPk37e3PsRK2A
3IWdFMYpbFLUylRfJy7OLN9bFJ4cIhcm8QwLIHXUMWPd6cv3cq3m8gjzdDjh
iEWRL8/fj9thcylxx/99ExzPQ7nASEz1kQTVSJfAkLZUjVYLgw4iNyILmJUf
FLW8P43vvTKguAJQPTmZx7EzSq/63MiYPIuCC91xEi1Y7EjfOoYaDID4NZ7I
zJobzSz+AXVwaPW4H4VTtw6GrQkAAfwRnxXwcupN6T/CZKJOW6yWMGci7rQG
2BX3oeFL9OGvNQefVBu2gz2Ie/7uIyhBf3OFC0Qq+S9zSXXQT/+kmEdWgC6p
jVAuGKEd4HbWIn9YKeVThkPY0sIatVpA6KJZFXIk/arGETKZKhBbiU2Q+BOx
cv1V1gLy9TfYWU3En/raT9LQwRF9dpEiq1oOcA8jSh3zP3xaMl7Pdbd8Z2T4
BO2ne5UMIg7dVhQj0hHKA0koZVjSzNm/pGPkq8LSiK0this+tILoh0QmRoA0
7KrOrNRjNlr8rtIAnmatEiIrt44qLKBEHmOhDjxVOf7TRXI6OR+1qnR4GJZq
Q7qYZF2jWQ31zv/ea5VPTrDZcL216O0gfe3+iGNpAaGoSogOg6XPuo83aEY7
r1kYPhE8OSB0CcyPXZQPDWosM5F3397UKl48Cgj3zOL3dehQ5ADXhJY8ijzo
JLk/D7Qcq7RMAtvvfnax3Ak0T4IYAFt8Mb9l37tmC2hti+cJ5N6bf/keoPbw
HPFP7cOeWXVH3/UM9mMWA5QluK0BISu+Ko8a8soMd0DYQ0IJa/wOsl1XgfY9
poL3lgZOfXj53alGew5N1/p0GAK+7cFYTkgKzSqxaM+wQ6e5abAh/WVJ3EHU
Zx1wyaCum/9EMRgFua1eT/NjEPG85XNZgMhTEq3Q4UuMZ4Y6zLPE1QvWk71U
UQtDmRd25xZ8Umt55ARrdNiPxvC0t41v8HmV1zE5Vb78WLMwXRrPuM/Xrnc3
mDCy9gHAQ1ROhYC0TiBnFW4APScv5rX0CHFrYCkrLcI/S/QNzNf8WYuSIe+Y
79kuLr2xj4V4nTNsHdDsUg8IddQzOTqE3LkrbprIbdePzIHgz8gIWt6sP7f+
uNYjV6jFRgSmzy+RqSsGEnjT+6/eTnJ598C1pHKIkqt++doKMhHgwI1ARcjF
FGijdKyVnZr+l4d8EmT6K6pbJ4BD4wO2okYNfRdIVG3KsFa2BIozy4f6BwDX
FVni2ka2ip7/uT7TNB7qCTlZHonnNbOB3Nj5SEZOP8mQUyhEsKMpJIV1OShC
Njem/oYIu4XATHhQWQlbZ6yK1T+T09jfNsqaujVK8r/xHwdvzsdv+1ql7KYv
AqupPiFckMyLAA+2nSQ/IrX5Ee9Oy0HdXy9GWpWxD1itefkL3jaWkfThdC73
GTX1v/YsgaIfcs8qgqUCkROtAIwCvIygtKSEXKA1SsG4Zio0uxS2kaDEO41Q
gSocBLB33c08/vdKawDZxJMiPl89AHuRUXwcKo56CX2AyVU7uag6EDrGcuef
1LwHZ0PVb8+95fOqKAqE4874M6dU0UoSlYBOpSrzO9erg0h1htaBPSpMqw3t
OH1DmBNvJpslfzJR//F2ek0vmZ+JTW40Jn9o/2Hd0PvXGYK04HIUtrPC+z05
4lLX97DGjsy8k2ZnL5h7kbrfj6P1jRC2vm01X1ngpxfNYw2yTXUmA6T8QBsf
OnPgYs0f5WVL03Oj1fwSkNU+2fRGaUDsJflp7egtS/zq4OaIYkHHkBVNYfGL
fAEIkndg1RRn9cNrkMQpDrb+JteRu+zFGYB9hr6dhxTS6OArHKyOeGbGJrjr
Cl9agwOpfN1J/LRy072qsHuG4hZVsezcfGOB0o5/+rwsQLbw7Hox7t6FbLXc
k4ZdQ3D3zz3kLOS02HrWL3JBo0xoWPY5i/bveHsTJQRXkVz6hmCirm8eKAH9
arzoD6Mm3XC9XiLOxEHwmqgu1Vaxl5Hf8noje24nDd0bvKb88epQ3un4gUTH
iGeJ5H5l+DogMSOetwSzRaMZcwHw38f3qUVEENiupWNW3lcfgpu0jt2tCs+F
UUTZd6bD2SwbSd4kgy1zujq3NNUic5t3qYxrdwkJGhsP1g62VHtr3d22udoI
lrMX3ePRTY4EUgt0WuKbbkoNnV7I4IEZoDCHyV+6YCMNPwxkf/jqe8mz7OIZ
h6rAi9CLyvyhYmlb5q23/TDP3DTDJGHokY+BPRr5naI8ZKddlvgJc+DG0QMY
9cbQlSMhqySIvja+UTwUNlcjJmEoEEhZ018PFyTxjDSEBwPt/W9ho7S//cco
hNuUIJhtrewbq+jHMIjaKZWPPn5npFBvH4ItLx+aV2zZ1KWYjFj3h7Cq01bP
WeJNjMhTIckeB4ajh0hCBYO9M7eb+l0SQGnD1btb4GUAhS05Tu/Yi7vpHGx3
a0jKLkPstRvAfsGosJ1xFmKYjdS3Jd9oFVbJfpM/sw6ccUb58c21jgZ5v3UC
LYH5q4pH+vox2J926SCyTLoPCNhgs8vVJ6BEw3vvpXaQe/rmGWsghwCkjy/z
/MfnGRvCFDDNsj7x70MDtrrc1jHGBWZ+vL97plpwkUwT5oQy7HTJIE2YTj1K
i+zzOr7S40VzCDEJYs8oWPxEjhaoq8D0Fa9arJvFjIZTrZPX2d8VhEMC0fx+
p6YQWv4Q7Bk3RMuaVBvhw+Km2tNJpMFnX6AQSL8in1Q8+4cOGcjGuqE6dsLI
6b4lN7qFLw+e7zOV1DetQteMugRAn164eoYYZnFo6DOqujSEr6Vvf+Ot6bXc
9nK0RzP6dE/HG0XUiER5r2s9fpOUITfkwpQ5Ct1UsUkFOCofgXKxdPaLib96
enHIXAVdOQGCkqnz5MGsm2UCogLK8qHGKETTnOOWJ07YumjWV4IXWyLO4uXI
ml+r9hI2DvlenIhtr0IHp2UJ2v0PH5hsmr3Tm9uX0kEsBmpK7s0hE4RO13Uc
ob+7lMj1U8WvjgTEF/6UT5r0UzKEVwXsmyIuTRxpvqb0TzAsYMBvYzSgTnHR
bSnpy5zIjGdc5etYxpso2hWZ0PVjhMwJCmHoZjJqg86i9+xyoSH0SWugJz3e
mlku1jEi5Z3ZWIdeaOm6Wx/hSJ2bBye8BuqzvKdJ1/shY6ptXjXdSXChZ4FT
A4e4eHVQiKosIeMCtmdXKsDtZw3iY2s6GDUgg1yUccAqR+th5CK1OoclcraS
ecKe+fFl+4Lnp5PJCrwGVUYznQMb+baHZ+2i42TnCVNyU0K6SBsJevwF/Cmr
n1C/8l5tbus+cLCu/CmmYrj5qtWPlLtzqh0eeT11TSEbabcwEo0UQRY5lkDD
g3P/Fc3IjXpy54FyuElcc+OsgEy1mDoakMQkzAxbgMfacJCz7LDjXEsEpyvV
Mq2ehwnRczViVe8zeiiJVuJ33HaF1mgf1m65uNu3QSg39hWGud6CIy1nvIrB
dkJ4GwgZRYjjFE+ndIa2onZ0kvdNz4pmcCw5YGU8Vo9odEWvxv1TOr/9CaOl
HvDpEMuBk+FO0raVUNWuO1ZgxMJbmUcyvUH1KKeqNT/2f5ZjQHEtaLi+xYXQ
wemGNPKhHg6/NeLMeG06HEzQrfQd8xbyA8Sx2T51C3e7TqLxSvuSgp/KbSiK
noueGVOtW81LYBdwUJa5TgwtcX5YdsLrD5iCpNhbvtqTd1+yn0b/VVrIqT2M
yIm3fEGygrgvp2hvMS8FC4FWog9uhSI4fOjjyMD/69+t3/jaDpdWR793y5mG
J9ZRdT4mwbRwlFUQFZXpgAyGYJz6yaAHn9lGz45C/BOOX+MCj1PuvqZZQWVi
fm8WlCN0cBsGuOe4cC+qQTQvUHKmOFPAGF0RBpCqtNQchMmIqoTy2CtZEEuD
oEx0qlIBCkTk2JPkqwMjaw6bmFujGNIvQC3cclDSxYuP3UzXBaEEZJnVJra7
hWR6vRzFXHHHUbImlUiF87KvYMXX9a9OMApuy1H93nKlyMFO+QP/pReXMNaG
TPJKQNlhqFq8t7aBPOoDWncm8FTwIVafCt+pJYLUsnkr60q8l7hhvuGFTmkY
4pKLfDIOyN3p8Jqvkx/pkD7UT3WErpCTpofY2DPLYypHnPPfK0dKPrlVSk/R
q4pCUhE/6ihQzn4Rw5/YmArlVhkWtA0oJQ6HCT4WocusaBTiRbMhmOPs1jp8
+hYrTF3i9plhfQ4O43Ga4F3VfgN+d37ByA79guIXX5aAPTQeTQny0z7RlMe4
t1Ij5SI8PtvWqiI37b3QOOyufNPYxefGDHM0KA6YMrs2YwVMwQNG4J23spem
ZJIZBeQ/lEzxGHO3tjTfcZ+VSE0uokjLDNjVInXv36mGpX5lzVyWZt1SqTwW
DGXYwAN/1zNYLxn5GdIxJYII6i9/nbgeHjW5YWzqQPsdfMcAeefJPyzK56Rh
xJluFgZ0UiACO0oM0TxKs8Nz6zr0VWIhIiK2UEDJbEU6b6TXoQ4vY0pTz3gg
y3aTiCnKL83p/1umT0vmIPOxXsZugL6dVI+8wCyJn2MtuDj58kXn2hineA5g
WQF1OigT5ZmSBUZdY4Gb3CI0mqhooaHL3ug45fVZMHaMS720YvaP3ukFWs3X
bw941kpKcRt9I67OIKeKJka9VakgMeMvAgoinYl8/uJvbTqAqM0w3JF+KXyJ
3BRatnH72xlQn83Pgi02rerxW+z7/XlRBt6HvAV3TiYjPi6WPV6tWCY2vPJf
kq1+sjvEwJ0GMVpA9CiW91l9yTBvVVXKDiGYdOqamn7qRMEktKtf9lqXaGpj
Kc/z+js9qMqS3e1RaE/lZ6mVttK15lirx4f23Jorj51P9iIt2gi3EhAB3AkG
cXYaQmBwxzL3PEkm+0z5F8upzgOLR5WaVSGE1kf0HTfnNwin8uIFi3yGr6DC
NBYKzKDCsj0dYj4s6xwmzPrWoZS3+JPtCGs3+7WIpWNKIXLkBwV+oj7V+2Sk
zeDyrvZ5u/MUyb+M8cWmrTESBPv67xlKP9CmYYv8H41mmAUWD4FPOaFAgGD1
tbMkyJoMPV0kwZ0IBE6Q9h15mQBJb291cz4JW0ElsCojDrRUyXn1Nbu1xWl9
1USqKXZUweOJr4prYQRyzZgr3QQao+8Ztsb7+c3ejaeAG8fFYJCbrGCB73kb
13RLQ8dGnrKwGImkAoTI/Pqzvu9StWdh9KY0c7bagNlADVPqYZCakzRjqYT3
BRLcqKu0J9ra2oK681m9LI2LHi7GvQjrFYk+OnYS9A94rRxDFYSGd8qn8EV4
ebLRHF7TEE1LGJYZ8UDoOWZn7IBt+sTG0NgxWoRgVcJVbIeLKu02NxBDtzwM
EU3gOCStDAvweOyi7VS8zLRIr8aYaXFQtE2exKHdVy8LwoLkf0Gle9uVnauA
WykcUbPmOzON6xZGn0WtIBVMQGi57w3Q9LjE/PGh6RZtfTElbKaHQ0LWcxin
DlK12DeRt47uJct5feMbS/bVCJIG424xjWTosJuhkxSSfDob5V84pV1nt9gl
lRsp7UaDZWeKvGtOVr3lqTP+JgVdrTNV5KafMSvJ30d5W+7vOSUsPge8Hpd3
zwAjKqvcQSZCuwiTkH0Mz/nHrhW6p0sPwkeK7CvynuWZ+I5a3zur4CfXRDmh
wnHhpZE+7UjTRVpoGSBcTGgJDcnQh4lQ8UKXRYSQ+wveiAUt9ofFiQhopzEu
YSxo0uvvkeYwjZl9rCgfyxtYx0Oj2BaiqeEH7w4hmc9MKMuAZh3/q+1GA1zS
4ZVTz4nV8pO4frT6p1dZoMDa/fmEJG3TKHqAxsGHYJ2c7ZqqrfQJCItjLSfF
mPcNLKYwrYGRGfdg4usnbDtXOJlakHXdUAdpWj7+W79+D8FXISOVltixNrWi
D3YepFhlk06LA2LKKj3eNhkpT4X8B1YjTOOzudbMcJnfZVWh37ZRz82R2FjT
fe59409aiPqg27Xv9a8LVwnysg2WN+H4rMDNJXjrx0qbnb7S8HCkBYSGG2iH
BDxbJe/b8E6aL/Lk0KYFiRQlVWcqZfqyF2bIaSoGuSfi3nQ+94eZUoT+9SGm
NXImQgHGuk4sKKb6x+HIpjMrHexKMn+Fo5sx5kx1RRLqDMZB/7SGDt8WsbCR
9cTsFaQjJcSi4Qs0sFSXxk+IG6Hh5Xi4e/CjMO7Ad4XquUhg51KZHVieNJyE
XGJQ90aMxs4lndTgke8LCKF7Dnk4reowy9heztAnekt0P4XKSU2eocZdzo0H
zsMRnp0XS0Ucd9X2uveEAjwqeCVFDKjUXMRtyjx6Ke1OgA1RFHk9JHCP7Z6o
K0z9q0LIXAWdLmdvQ5MhpSWvCbYwtWibc1f0h7KUVydmFCQCEmB1UihZ1iqP
wQO68FIeMKJHIaRidAbXlmIB5rOSU4O+zjsX+mrvwEiGHpsXeaS4YlZUtzmU
2cPn2d6lDXKMPk+UMq8xZnAyG13qqDbXx3pQM7SfbDk4EitkEqsrkoTmLSwh
7TslrMizcRJj1ynlgAvFw9wCPaWGpxJPx7KobWQONJFTNgCiSfu9vi1+lVv5
fW+cS/0lNgWdvX+g4ww1nueWx3I87O5RBks1SQSIpC2JZNTRNBUpQcW715XN
ggtChPL+g8yEnqKonS/M5a8njy3YZpyT03YI1xOv0J/wxkArAhWGV4SdtK5Y
QAaXk5MaADScv91mP7wtRcAtgSrPe5EvghjRQE3t1ZaUbiZEXPi6HNcJCCEk
dwg2qfmxN3apEhmRBX/EIivtuUTg4kEkU/cQ5aQ5XC6A8m5SWDbfYLKcHL0c
9XnwfxvIaFulnVV+NtKsJSXEpjdRrit+jMyy+6Kzntlx90ugYMgElzxFvk4b
RoCV0TZeHikvrOK7yLnND1MU7dt1JC+Fd+4WGvvVwR4ruOF/pOPD0rFhCACG
mRerJuxP5UA5/beQKsatujNWMkCl6Dq+qEBsKWhz1+u1OZ4+X8qWA2c62FmM
5LvRd4fx6CUglnwDnsZ895ezpntoup6452OXTLa3GbNj7vjrArbsI0FUXtsk
WXrZjcFXGLzPpx30wmoUzGssqT0q0qiumOs4AY5DgfShRpvqxQOtAG7Bjj9C
dZ9LUNtLR8PrrjevfW/a62+ZXBZ11MB4B6gBDg6jALhfg8SD+BOqEbofhY+d
5Ank0Xt5ylaVBKbwBjv/boLHkg274WrQTu9rrTGYF9Tvn0HdPHfnEpSCDfI9
JibzQsKTDcx1VZjVBZMCreBiyNwwIxDTh6ztLSXzrSaUuxHda33JQzo64DVS
K+qH2q7p608uwPwRnDHOCrliitLlJnlsPFQDv51qYjrX5ctGJHnz1GFP213m
bj7YknuRwVwlUAtEMVrer7YdGXQwBvtw+Mah3zGe+/dGlte7YGl2nNHmGnEq
/ojMzPHEjX7MVdMDgX8Az4YyqaJyY3Fd1nzNvAdeVPs1t2ECQsZyI6zP6OQw
shksU57vifN5Sm/7NYwqbaxvbp4Gld1Cb0MIhkAoRC2u/poCvP804QNkKpjo
GKMBrDf4POULOjlVFOw117o/5dlLHx/N/plvOl5Bws+wBb/ZRQBAcuAzVFz8
jk7XAg8irV7xKawVk3BKH40rPfuHQO9SIyvq/LxXnEbvh9B1UiouEn33p//U
XCcW7Mh1z+yKsN3J4fjMbcuukZpT8zVgLsnwJwR7n+Zve7h3K/nd00ECYEBW
+KwRvmjd8EFy7A2byFa0nu+TUhkZY2NoiofTnhJY50n+CFMMJZZwpg9h2hPB
x3rbs8X+SPypyXQ2ED1H/n3UpInxOo31FZzFFeFneUvDBZWCzhr9s9duCzCd
gcFWGahPKIuoLQG/J3uvYhQXnOxyFXv/X+cN5d91hOpd0RxsXOtrhZ5HnRyx
fpyEjVgFy/8hekcatY00GNkvJLKXnbGcMrAMI93A+Buu1TsXzA6pQyMd5oDc
Hun3B6IKOMlujV9VGvuNPX4vp60XTIYsub0Nc8E89lAR9X3R0isqsf1FdqfO
t8FeF8pH+3c3DRAn76FxH8nO3zj7wXzYzL4VWZhvZtv/8cW06GyQerUkC9Ox
vmwCAOPcQ/of9YWy+NBELFxz8rHb4ghDTSwStcn2ZVPrMt7H6sDlSRQ+d8Ha
jYcB8qBlI5DJoNzzb1i1gTWTBDyXASWi9ZI0UyYFrJI3JpVxxOjFzvgg9/ue
wIBSEyXi6v+8KvWGnYugtO7QkKouZviKPjVeR5GlkPgL/HXDRlS6HI+JTqsW
7o2u/uYzkR2ipkh6IfTt+CGY0cCVmyUS84jzXRH8LoaYwadlEQlvvhj5vh3q
GBThB8ubEdCJ9sxd2awvC3MS4HwxMX8N7EIiAvclzxjrhbeDUqGQ+QlpZBTA
lSCqjj5+lv8CTcOuu3fgNEQwurxDsQ2zOzTFodcfEeQWFmcbnAUyf4tBDILg
td74+5diImQF1gGOc5XVz2eGf97sbIK9JqVKKQH94g+HwXdwPHYJHDo6wOqb
8Uh63+XHzCGcAZj9OgLjNqA5yRxVdI3fzneZyaimrcV2RsGy5LdyKPKEOJlj
otV5kP+VwVL0CinGtdve+1G+bPRWLugUccyrrSiIwLemuDFcIEeomn4xax8f
Phab5c5itUJMxyY+UQ7KJR39nL3pqtqKt1qiQcpn4bhY+NRRzPHUiofPE0gC
eVFu/LylKkyf+C5vRuncr1jLyFlZHr9RZ44YBYpRwzkwuFJPDyVs1uoFEOJj
VJb04HuZqlPLU5dEWYEM/+vjUr+VbAigS2Qa1oecBKa8YazD9qUsGTTEYe7F
Jbq1zCYVqAvb1MJBPreZdEoenWaPNgNJY4q0bo7b/ZhAm2q6Txv325cuQ52x
Z0ASUEBlp09UisUuRPYgoCeL24iLgd4exzV0ma2uY5cS6dstU+1afpwyaOGn
22B8P3MCYtEvLOoUGj4fWLf7cg5Qb75CZB7mZD/0Xr4enZxQukHdmqSbWutn
9SoR53LJFrJb3g5KglGGCKmS/JBc8BeD1Gt6JNzj/IbmXJxmslwn1xKaF4om
gWEapKIy+VIMV7CImQ8lOh9C+2hviAcltvcc969PKFvcb48H7KVZgkEk8D39
QmVv86cGl0fiVnV5pEpl7qHCs1nCDx51uGFLjTixh92CqBHqZhNjDPz8nOOE
RnyRGFy1QgwbZMvUy9Oe0YaioPQ3UshPIOuljGsgXaQ6BQjaJ7el+D4edd7u
LBBVGJWgOq9Jb0n8g1KLrjTzW0P9rZ2hJvYkutO6sUJIaR0eScgEHCo+2woM
5/ZYSbLg25T1JbN9rNrZvBpYjuUz3sHqP7nyvkUaBEFxfDR+V3vHCH0llSQW
PYUod4y46pgtIW8u17vcvB4Z2DeMJoUXgFIAi6S2f9EPFHS6kMO14yn0X09f
4qSDqxw3Zd7JivNL9fxCSTpK6NwpyD6KV0qehHJGrFrI0EJ5mPxKo6Bv0Wvk
5a3t4H+M4E+LM+0JTJAdmcPSslPR5Ghujs+3FA9OEMmsAmDOSBE/eqf+CLze
+Kd3GK655M/SqSAwhkRJZwtJQ8MZ0EI09uZ49i47JRDN5VWIHMxOWr9h/O0r
ksd9bYWAcdCnSE0eC10h9tt13bj7Tbr0sa0lMmE66zn6BGAoxR1fHANt4wJa
BArRc0G8uuH/eFcFh0Sg2G1dpvrS41aD0u7YrCarxt5JPNd70Wlspiojh4lR
EPYj6v/l1QvxQ3kmRcyHoBJSMoqooUnBCQazavm7eFWpyy5aVSgGSkwmfwgm
nBMlF0p9APnn/zuiAuvqk33Mm2xDdSgDfFY5vt2lnaRwIgE/79ABipjbHvFD
4NgPHuAOmvkGcHelNE34nKsMmuRy8LjPgWcI/r+zvs/0fbnkvKzKwdugK6qB
ogH8NsomeIcPEZRSYvTVJmZZ4rPjmdFBV9yWoY4/0yDSIwKmzkML2ztflBE2
/+YmP2sSgglYm7MN4+l8cF9bnrxvnV2OpOzEhub/vXsopUnzDEHoKJwBtxTb
uVfmV/o01nLtidAbWzxGj6h9lNvtBb32AGWvPZo26wuFHloVhEv369R4l0K9
pC5YhkwR6oGE3pS/in5tc039VBlqptakOWUm1Qulh4h/SJ8lfqV++SVboIuB
e3JdwkKNF7cviCLQWjOUgje7F+Ptpc+xnCTYvOOYHIxS1mm4lZU6IlbwNGEt
BsHwl3tC8+6TuTKx00u35wwu6HAmfAVEIpuJN8A1MtQh09Bzri0qAsJKP6z0
YpOrviJwYtXqp2xO6OmQi2dPwP5f6f9elyS9RcTQdwrwIFp64S6CyJrx8DyP
z4VqOCtWhtDLdTGlZe37M6VVxsKOWNCmWnaeJG/OqKXiZ7dCAM8QjxOmnDQF
5u8wrplMP849kHybLN1YIA6x+PYY2sG4gqm/qIpWASrdLzebUtX/9LESW32z
QTbQT1Yc/NOohvpLfPuVtDC47l7j+9zKTcQZabPb7qAPO3jm/e3zD8zG6OvJ
eAJUIKvoyklscJGJKuYNE6YWhOTUFKFn/eljd14kCJP4ugqE4rnna4+R58vT
tYHCK3uGtxb+pYqwhu0RHfkg/IfY1X77ccHm8YYY1ujzczpkW5leFa7qsXNj
DiYZjSTcfdhX6R8cZdvdVKgkLU40gJUBU6/Rn3Y5dBqTt3WSOfsLUgf9NLjp
1AtPvT7HOvJtWwSd8cpdYBw32CqzjfForrTvdA23Vg5rsQcIBgn9oDQxQeuf
kwUfddI9mtVs54vZqWTvUWK0Z3FGcqzTwxbt+wEQDswa5tdnLqXZbgcnf9CQ
wdf4JHogMyC0nGpvRzhYPz8yt11tDwqTMHcSZ8zWnoq0TMg+ICCWR8Q3e2Gv
uIhy0+SPOH+QSTtb4w5oD92SHU8xAb2CPVLqcOFX8R0lfP3MEDUaSM/lwk73
g9LLVAVutxIyTqY4oEBJD8yFEz+BOKWU02MVIju8wIB7U+N7d1fgbiyYo4dr
lRU3sRfffkJshcN4M2D51rHzg9uc0jU1UAuvk5uBRp6vgzjYigxYh3QdwKBF
sFB5XUgEybPY245YIDjEBcn1yG4Wgdk9kcO2y+p8YWDBeIMU3J7WhKrFPRIn
1x01sLYVtZBXFA+OmYudbOGZQvauiq4bnHd5ewpJsvuspBbxzmspJLz7OheO
0f+dRcpGrHJvPBwe8X6DRmufWVQ1JSXyzcMajyw95kZx+hHRNFEdUpG+SgGX
7j8pPP4snX3Gp4pV2rRcQSr1OPJrJM/JCnkaTHmBfr0P4PItHZbYWauXvKlS
Ry5vLAGI4arvKYDMWNtRler8BCNP7D6+B5TjnOQ9yEQzwl9+e0Hp3tmRoRB8
ys/+YIT1xNGCyfePtGxFBiQ93fV5EW2G9fJseEqKHTCTttnBb7R7Jrj2YtLO
HE1iYe381agxJWn19jGoCQGwojwTaqAF7/bZMfuznj7eBxqAF6WsMU4iHYPV
agmINuhG2Y+BzqrtKtAlLweXKnmI7MuPsWmJxwIlFdp3CHWiZ9NZBcwMGfjx
o/9EajxZQEZLcBx0xJDVKIBp/MFk59JjKP/l+L5oynvdqpOCeVgygu357EnV
9mubj7PoQZgaPiaymQcIE7vNJUM4HNQ7E/NZd5mG1f7pKOCG5ZudoAF4IYV8
8mo8O0lFnG/CHuNAfk3ZMzuZX33tusagi3JOV7vb/fyiVZ5nmedCSMKmD8Is
UYaDt1b/SRQJmfmo9Baw1ZNV8g8wmx6ls121odkCztbdOh3Ezmx96aORvuoq
Mo/tGnnhdiY2wYZel/4QimduV40gRnWUOJcGF316mcaBjfTISkD5UQM2Pqmb
7x78+6bv3Spr2zaevz3mYP9XMG/hNsgEfF53gtKrOW5YI/Uok+SUiP+V4k2a
d1ARGimGM1uALAtIjy0ycjj0svdAEgRQ+su9zqd7zNubDU5ze8OG9FpjmGF/
DKl2ITfjv0at4fxa8UqRtxnA2qvnt8lTars7nSSzvc5FstNB5QlH1EccjrS7
Ug5cBWP4TyaC2cRL8M74mlbPc1EE1gDBdGpJ2myh2sh1W8PN1MQ3ummWgumS
eUZYrVS3HLg9UOLHFTi76b69zUoD+kY4RANUlUI9T3O5V+2VMowyFRm821UZ
VlhKQhqMwKb3JTVGcI/JphhnWpRH6DtwzQnkUWbkj1rwFEp4Os5JeVmhcJEM
aUvnTjziBA+HWvCyE8scIgXeqoDXT/vRp5F+lb5h5R7SW4YWNpJOCxCoBV9k
yO21AmeUkG4vrIoCVRuuNLEyaYA4d3fTnSDdET/nfItKchofn8b8ASZ9XRT2
WH/XWT9ettmSmpM4kXgddcaBIsAdoh7R2vSLgLOtlu9XiuT5qtymFcVenx51
Ta3cErPnOj2Ddcwr9jY2Kbd4uvG05tkPDtmS9NbUPFr8ZIvR8Vl3Xj5YfyeQ
8ATChpE+b/xr1aiDIUvzZQ3/ZkfhokqdsmPAFyQaBl0LPhnwMhxoG7A3/gLn
tyPdRGIhf7/xxEduLPKUnpzKktGlEfahDbRUi2pBj3VUFVn8BRk6rxUVVmSj
ctkhCMPxrQon+S2fXOeC5CJND+YpOzX5lHVBrju8tS0x6dO8kRJPoRJvIOtI
qlWkEVYrowc3A/wnuZlgvENyWNe5xoS2qi8JiWagtTQJ9GujF6WBOwI3ajCM
OJreJGVhQedwbIYRuR+3+U3xWI8MOR+gpznUuSCg2sCWvrCGInowLlDqoAw5
CR6n7u+UZ987L7SmRGcDpTEFp2KBr6tQdTFpsrv1a5s+n61b1/6pYujODp+L
KpgLI2cO5MVeKt3uyWVTYp1MpG6JhNyepBkIMx2R9+AiLnxNIEw00qsdSY3S
JCYc7wXksF2sm8yRJQR4FrSyzfCxtgNnZgkQvIZvxd70vQrBqMq6ncvZ19Js
CRQ8UYQhEwqweu9TyD0q6eSKLxGSSjdsajMufDT2aMUE82bYb8UHnZm6j5hz
WHHqTTPhC1cV+PA7KWbGMagCicYsB3mbpqQBT5SCNoLPUgqhxwCTaNpLqHSb
bAzrF2z4FtY/ZJVaEWcH9gJtwAgg0H4MVRbsfSaPV4t2CNce3aDSQKUNIEYY
XNKdspOEAcnSSt9FyO/i2Mp/Yk3AQXzshaX6wjsBMhmyiA2TNVE9HcGjL2g2
4LU3nKKLMb6XSBCB3wcbg1OGRCs0zhT8dGDwXHlQZ1e/p+kh6wkyx4SSe1wU
hmnwUWFkZ98e9rcffkKLsEgwvT+/wMQjGB35JrVx56HUr/Zma5hDi/5phDEf
IDjk/j7k0eGJmWByCjMPfRS4AZqRp8oWVnI49PQqm0E34uaVH8fcvxapZAK3
GJAGdIE0gIOopLQ1eLeFL1/MRnjxDqOPxefHCOgPqSOx5w7YuF1/0oEjn0g3
041ErBMjtQJ5ZRbL0uI3RVdQ9RwKJgGFyTS/QPVSV0h4Xe07BvpJSgs4AqwW
/AywVGHDHeCj49iHJD95Yy574XwRBfpUM0hT3oRTz+WFQWDeZ7OnTZ7nP9OM
GhUDlaWQfEf0hMXhTmrrTmzaoWA5DdHPnmxaiMPisTwGHW5aDzPbN3Jui4Gb
bBmiXd/sKVjnHFiHtHp5UHR1W/5TPSoNT5R+emuSRwwLNLaKxI3VhaVQiP7i
Tf/8gYP5CxlNQbCyJJpRODkOZMAdC3vjfLkw9wjiPiUNi8fMeBIR/+bpQPdD
90IAp9yusCLLNegj/X5i5U23qq+m+MUAsZ29cM0HsUv5uL6oMYqg+OhMSywc
bVtNawfO5cnEWzOZB0vX16jXbshRALbOzpePJTRc9d9Wl0nIJNE6nuqR0/V9
c8R4VkCqH8LQpmtq2NdWSmAIJ3JXBSSfViOy3WPkiWIEch4CJebEUZtQBi/D
XHpdXI5VGM0T8xsuXjg8c5uor03dFBFQbyXcUiz3mapYZfyIH4TEn+/Zw4zC
wGrZJ2nE0oks0lOizSCPVdtWkVeVHcclMh+ceJTH3hG+7CXVV6DlAr47DgyH
mS3NM6WC6Fxr9Fdkwh2l0afw/2s0L3H+ZemnJ+U0eiPfEzyWsvnFQ07GO7+1
tckHeeg2B37ip0L3vQWZGuYQeIkbjxNjSXf8vNbochNQ+3vJadT3l59Z2ux/
/eQXprHOvzEqoMip7mF4GGjwKuwkOv9s30rX3cjWJufFnDr7S6aJOPYrqfaw
50QtNK1GrLa7ZOFufnlrQjes91pqUBdwXmqpyFTGmYtxmfKnVXzAVx0C61V1
WnR3lM5GTyUY9zgzMA5Gq/zbXwyjXBuGIWFFqfcfaK6CWYN2YiDKuA7fmDv1
env5jEb2DhZp87PLoI4mBAlwOVBcEsuIwaymA54/DViBkqlzgJGPhATN1aon
ENEjKBsd5DM4jNHeLB1k2Oc7DGpnJosDuK6Gy4Yw8ZFzmiOKg+72DfypwVq/
hUvd7UezkB/KC4sT1WTYeuHe4rAsO7PXRrcrLKYFrV4cYiYeTwRQi5A0hhHf
4S4p/VDOE7/IrB0ChkZdLZ7azUWyU35hKOTjR+Ajk06jIHIQIEzrsgvV+JLM
oNq6tqu9aVXkPqCfJKCOUw5PqFLGHcEvwYNn33oumJKbBsZw6Pn2/KN52oZR
2+D7MvLQZsAP413FbWVeLg5bqrYDXPYGz025jQsQ9kdNCCgFVhS8HiBoT4QL
/BDpYtMeEEqYah4Ri+tOtoCpPbRb3gGnpt5W2Z3DbN1xiqK7bTXlawqSbbTm
k5QhjMZ0a1iBbhKvqawMx6zqFPL+6bx9perjF/+5mayaee0Ct/8/8O6aLwOR
X0x3crU5mvSbkmckBIDoi2/VuqbSH1XbR+m6S+smnO85g8yB6QIfYTG6ijQV
LoXJqf1F/c7NzFh9IZuSWVYtVQmKK4Ma/IpKO/wz6Ep6FLZEpOW9Nzsg+Qbq
0AqmFlFngfTcGiAxKKXp00Y2IbHhZbLTPQ7aT4nvzx7dUDFkwkaJ7epbh2y6
CT1f2RhaDVMi1ZV9VUtgDOG5HOBoOrsIOFzyR0Wqt8jiisPF8y4aCrOdn9GN
vWrP4kFWI/xmCnWP7YZexHlrRPcbobt2wRzXgDux/D+I7+RjvvvBSFTmVr3/
D6XiJDs0X7QT90nPOVUb0w/UHqEmGQ8AcLKjHFngMnQsxMq/hd2QLDXKU44P
me1kUPr2q8hfGEjTv6AS5Bgj6PwgEkNSDcwR+s93F8bIMX5/rkD5wnivaqZZ
CoAy2DM3ypiMx4ZIdT8LhLnMvxSlUpq3LOUCUTDezjcNkDF1t9/B5QLMUJ5o
38KynFyrdlRECAvuOOjB6G+ZO9eFf+oNuzu4FY+kMkN6A1R7vb9l1uc1L59V
ugmi6E+JPP2eu2ZuCy/SQfJj3DS1mY0kGFul21A3gIIMd72ZTrtuAASqm1ru
pkH+AtuzgU2CQXFsW0ZHtuNV6BcPKVlTwrAHwzYzNYbJqEknvK3dyC/kNL8E
Cb5KSFjc/meNNq8RV/G9IzZ22O7sPMJUa75vPjyaqo7Pmfb8qleDSEVscbjB
CP2qxbHy+0I5wYXbReJ4RaXZ7hZY1SeMXXdNeqpJB6REgYr78wEDrkb9tvew
59AqmKoTpbqCl56oqLW4VhgM1ZgKrcq3fcX1uE7gP15Y75jKG1J4heEBoKyV
uuDTjAWsydq0vEQf22Rhz2LcNvsKBL1LUrTcU8QqGzNxhgvsSUuQGjJwjGsy
EvrdjqeDdIn9/lWDf/aNGXUVJzcLhBEI3KhV0IEMhmkH7BfMDQi5YsUrJIDd
nPHCoWULSfkLcjWfZ16SZaVr4LjzPhgI4FS8RqwLVMULmpHlpXIxnPgmFJhf
TAiH2fmQ+uDoTXGB1KxiPPP0a39EtQ/IlXhKfhxjPO3nmVgPkpciwbu6T502
l4fPeanelZzxcmCFwjhbc4khuYJ0ELszUyBa6scn5Ug1wtmjuHXSpmXBiB0o
HugbTySRjdhEZ+Hhsu4rmU1/cDundsfspcDULTsqM4yBleO7aNUV1zrtPz1f
MbP2MheqR8o48YpjFEka3iJ1y764eXfcfgHW0lXJQmmUMxoghlDbCYggQ+tc
1lIsIjvH35r20DTCL/9dbzf7OKiG7hNXaZPyUNcYwmstLzcp9nSGc8t+Uo0f
nTrymo1CQb8MwsIoZ2OvYdDfVqlJ5I137vSiXnsSAiXHwk64gdB8balgCIGH
A/In7fcE7lyPsVd1ch3TXOa9xi2U9QFIazEGJT08bhSZD3XU98mgp5Y2x8l8
QCdEhC4e+ZGJTRUxqlNkbBsW1Qm/qFpm9dzozDHjkB2F/exU48eW0DBg58OW
GEQbBkOHvjiIcm50jkhv7FV+3XnUaAZ+utDjLxFQE0qeVCBRQ2zPxxaG1xQt
l4Wupinilasy0ddj1bol+vavwG6nXGCDwLiigda/MHCdZk364qoHBj33CFAx
HC71FI9FtKYr8yWu6QwUnAmwPuVnhafsiG1Sc9B0Ea9RFfN04/mAPhuPhPvw
oA5vSkX5VMjIHnrnw0RAewsWEC9LhgznkjAOlW+LrRjEjInJ0kKrqHUz13FJ
BQxLVuozqlZX22mkPVDVKvTXaUzwP2lVPyh5FTdxeyDj4zJ2cipHNRltQkve
WXk2nBsZovkzqOADPkWiTZrQYEb/0y5HG7CA+JfWPJjrF815wvnJ7QvhagSi
T7FIH9ntcLmiCtUqq1y211XN5JeFSAVoVaywe7714SBu7wreQxZN/iqq/ihu
7G02T4g0O0KUdeKVeMqCsYUh5AoHLas3JJ8nveqxUgiF/WbE93v+I45gO9y2
u7KwGjhj8KYPagYOWlFMoXgHMqVLekcoP42O51HFuARH4Obx1lHdl1OEMCjc
qmUHIyyiXEt6XlhCyaVClMNOlSWz3cZ17zFgK56P6PI/8EfHqjlfkfcvCQcD
BVF13kQ/diEn2uR082OVdW/FdtypyBOsB95LSD0biNV267mTYDRNuRaT3VK1
CxENLjvAdQmQ9HzhX2VIh29ptypgFeLhZc0K5NA+wX30bGywV74ZLarlH4fM
OtSUFsZlosrDMfrPIum0ERHv+WqUm60EaG9eT57jiCGxdH6q1xIJy9C35wax
awox6WO1U0jmcBIpOf1Ht0NgykZ/eDgE86qelDsM29LJa5+UD9Aue7Dwpi46
ex+9NncW/lDr5qgWEmzRKNSMq+r8A/gINEkdsikffjtHXLjrazYA/10n76pH
t+WncOlLrinKEcamxfVxU0dGjTPdjeqaZVydiK9Mz2sOht9H7mBwnpxKM4FT
yIIsjiDvUsCpKN/C/Km+2mjL92mAs1aeF6BvExX66R5nxz3FXlLd/LejZjIT
AL+tfFIMrNkzfrXxzykjxJB9y2UJfu8tFeYT9s/j+KUv00QZgTBaVfCsR3nH
RmKuUnHookQ417bP/WL2noze7LbMxFcb3zOPzSbk1/LEoARNHFIxkm+RZV9e
fStjOp9DMQEY3aRTBh9UPJGrXMTbeF7lKtqmfb+luvWwV5rFgtJQdCDO6gvC
UVRD49lYhNwXnfyd2Kz40NfcX3JA3Q/4glUnaeP5Q097kuY6niIOEOUBU2Lt
zPz/UDWXBkHyk8U0Iix5gjNOBCgpjJjAnr4ArEO95GMMvU8KE1JhjPxZZV9z
Ib75NNdfd0ACEsQH+bNVNuHvXCNgZM140ADwAdLTDpkYVg6wce2WPxcJ+/5U
HvdTBWvzd7oz+CMO+Z3Si7iy918WDDr01KqV5Jv0wFw3bm+zKzCfd+Xc/uyT
QrJJ5QxmbkaV9PoqEAn652tYCIVJ7MCxw4Jtje0K7qqHdxHa3aMuEByD8OLG
r9ZL2UI3yXYXCM7vp/+ppcieJQljkd6+aLl8pIwV3gC/4Jv4yY10a0o4qYKU
fg7DuuynV9v7WB7ttU6vqTWbC4PdE7dIq4yQmVeD0WaTPMH3rqmGur5bZwlG
6GIyUDZdbRpEHQfYYsPidVvkDacdw0kEUHOu4AVs4gNso9QKd6O71HMRTjz7
Vj0Bd8XU+zotba4h72ypfpwodswdmam4YgqQlq5yYC/wShAuxt0h7QNKVSXz
sGDkkJmX5xfQ8Y0Son6T4xJ0F/MDpr9aMF//1a43P5TQznuv27ROU4G36zAj
YFxUZbGhfIaS8Rc5XzvlbBr0aYq3vNVqXcXyaGzLNjjcE2UA9Gc6GN4NhzJs
bkdmuaLRJqZpivNJvTkPzDAj8OAoRFzsJ+nNIx8HEVS2jiEKb7pNiFLle7BX
FVfG2vpnlqL91DJwgloJkkFbzwy7X5Fkjc/z0FErLNKlwkR2Phx6qfkyzNDW
vQCbnm8h8GaqW2MAwdL2wx8reQkhAXfD0K18HCrNGqrJrrYCrZbdnAnVhVIG
sJuu2YXpYkT/ogYxj1g/d5BjhVZKVtD0mKJP2xv4AWglLTcrOULC1f1X9bHY
jGws2mI7iFP1NA7+/T2kN9TKhi98w8JCh4QM+9bQ4Sh2FBah1EFy3skw74Mj
gqxkVKdzq4bcG4ele1jlWMhA/sfi0BNUTu2wQEHHw7oqaqf+/I7JbqQRb8IP
KRY3nz03ccwKjxKXTDtiRm5fjgziv1G5hcN1Pw0tATdj6vgBuYxljKSZtPFz
MiOteQVtHBV9ZV9rrswzQobs2JsgRo/3jG/PgUNrnISIfjnnEFSuLnI6H666
VL7zzY6PFsCfXXvlVJ+uJD/ZIz4kLOHg2YPJnmGAh+QIs9nfHYxKXaxTj76F
sklM3shQpLkgEcsOw8qcpvEaUeAcMWoN4k2PXur3XpX60RG6DHwqNdXEPTT2
6fDdLL/zCLsF/vOpTfftuXgEx/ndtW4vgowzr7ACba8lXI8rrSXVJ7N5w182
w81YVJp/e4I/1qxjVOkcWVxqiX4zPH9mCEuzboVB5IkMuDGYOIKFIbrgQnxQ
fna29KGhnqu9f+MGMq78iyucUSRhDRf31JhEjTgpKyqV7VPW+YcsMNzzNMhl
u/2wqL22kwWo+ykWGgsNQaJ5JohYdq4uWxKoVa3mm21Z1Cy8wuVBEasHPvcI
SOWAvUQF2GzbVII0Y3VIkVHh1HSI0Glbnug+Aepz/jLhwi5VLgUaGBu0GFjj
q1mjlFohCYyzo2Hy+waidxFa/TZjCrQ2+j57OYJpOO57dKWdaIQbC8Pe7wfP
/DpX1IxdSYeS1SmClyE8f9T+FtXyDOHvnaki67Ix8j9B6eBBcEyV35xCVk+Y
UL1RBL7E7vBCBHZsMMdn3ZJTyhfm7As2LHbJCYv7bSuOVuRJYTobAiX1iWwg
O/GpSHtjFuv8vr83u6Ap6QKWSP5tv+d+5vwI7qEESL5jSH8mVZlpCeLUa0fw
XqL0KRHHtdW56ix94/SOgHhBSbmhlWX/s9uq+PH5DvIhpQ6+0PQn03alKo6y
b4qPZ7i9g0qsaGqqiIFbrux7IeQpghsTGSLGda4iJ/QMkXDXxWtXn0DU3bVI
ht7XNDVjBCKxO2OG3qtBNvQaAd3LEBxzjEBZ++DBBwtZDhPOsc5qkumrrFjA
goaH/VcKZMf/L1SSHXEHu9GvHx+3VnYjqnvkoFXnbgLo/o71kLOHSJ7Su13U
21cNUqtieDk+DRvrBoH7xr7Mq08Fm8GaTZFldc/NgMOeAEJDlSdwNRcyEMiG
XzS/4XzFraY3eatFZ7e7L9446WdiX7+rNCBJiUV2od4612yCObGAlb7dGBeF
SNtduAa8BcXTIDogzhkqsjTQ2e7olAHC+AnhzODZzzFvPJ2XwL7nwfSWNaKv
ymVEWZZNxUcoPC6pNvLe3tJJI/DhlhFo84CGJ8GBncIoQcAc1SOxEfNFC5bv
kiv6CEduCvrFbU5bSMUY2L9Ig7bN8WT/4qsZFs9aW7mFCYIKKkUS9CbKp/KP
Fci0+N4yaAMUubvyuljFTWZZqyVyXC1vSImJ1baGkx7C+qmoNTrqnT0MXnOq
Us1Csyy3xzRx9yGc8h07fIx19LOfNkzLvhfsIBSqsBcoY8Eq73abN1A9nQ2F
byOBCF2yy0bVLCQZLmshRn3/q5o+r+Zz6EMEJA5W5z743+MgVcO25a4iuCC8
skqqF3O+EiBtY6DMnGl+4DOing55Z6SP7CCtqGPkNxHXUF5sS2JK6FzHer7g
QH7kxN3RSuHzQYHs0p6smPOqTG6hmKGc6fuDSi6UlU872zNChZMwbQKq9B9B
cUTFwGeWdmDw0TMM+lU788ULPfGkMHA267hq2NDWJYF9oBxP3zrl+PZsvBHp
R4pVdD4fegikLZxN74h4LBknpUDkbcmYePoxlwy1JT+KLRFa2w50Ls7ttXVM
E632n/ylM6JQcuE/g4Hl24OEC/P+ZXVomataBFOEqu8/84GGDgGS0pFA0F9m
+i98GNqosvhEb6vn202EbWMbYYZh3vLXy9r/z9n8HjAAgjvgOABbG1LO0ox5
DHXgx0zKmsp7I4kQkJXuWp78cN+URqfoUCirZIjGXsrB7wwSSIl1IOMIo8s6
0wuHVbDv/4u8DXh1sRPP+uYd+ji//BHQWT3/MPVmpfeWTjfXHxlHG5Y8Q8Zq
+8hXnQwCHpI+FtX/iYVDb9T9l+kRYnGAE1Crp2kh0uCtTORnIbFNNemIWbZ3
HTy2Gw4GZSGdwVd4DGptS6g4saqnk7mBrjgaPfzz3AHN8rEGNmncJcTDdCl1
DUThTu4JrfpRDD9Wusoklh9WodeE8ZzUPJICPsh79BfGtj8K8yGFKy8Y+608
9aXp6tMB2LN2C8xnmGMNajaH22F47SueJL0OLrgf5UL0TbCOZxm3Kaa0c5TV
g7miApWd258J7hiZwhuphWixNIqpLWt+CkyUv2tXH4tWYpntYSIhCpysSc/M
tKhYwMUAMzmsr3eO31T1Ck/vnhnkRITCGdpYpx4cpFF+Wx7bSxiHU+jSB+jZ
FvZARH8+wiHGtJD9QqeEFYQQj7GuyxzbWvrgOhhdaiL9V22fv+HUF9L9MlnI
iR2WTj2ISh8l0m4E4CpjI2PZABJvfAe9RWjqtCaLWZrs2CyQjMwsuuGCWiJL
PGd7HICsffz3v+BB/3ETyKmT+8tOOGvtvN754tF5+iB9/RKRGqBNY+PITJMw
8UJ1KNx0Eatm84O4zFw6hwrs5JH1K0EYOCxjxXYYohk7dxdO+ToleBWI3xQm
lp5RvBsX9FyhTndnAbT3I7cywBchSDo5k0+R9yG7elPuNxqE4u6xeYTuKIXQ
il1mqUxU99gWq+vXZeB0uPPOS8wX3rvv/E1cq5KDSv7eiVsPM5t8n2wqD4Q+
Db9NoGJtRoZXoWjjIiJ+79pIExVnDSk7lthkEIy9gcWfsdaLPWDabV87jP8O
awI1VGxWPXvP0lxzawPw/7stOdN94PVfEUb4Iliu61vLivZoWtG6eYvnxSCH
mCHnPBsVpMzIBsEWYQhD7FN4+a9qAKF6h35csBuMqrKfTBbalhDTZP30hxxb
HzcqU4qIxTB0AWyTu932c3z1fA6wkPXYqwaRk1MnXJRsSD5KQo06w9LaxmBf
O/5HoTnicCWgBJneNlmxMsnvp5P3zFexZTKd0kdGSpXfEDVqRJqXjnr9dSF9
/B30KEJHE+zxuRZbJoWhuzLAMCsCrl2q7caxE+IOz3EJWWyuXViyLcZ5tfQ0
HtQY8fnGjbaJwYdVY2/yQLjyh9RyP19oUKRp8b1G7sii0Qu0LrZebZk3bRI7
rYEgihmsprvMDTfWGMbKXFWqv85a3PiWO5Z8NQ3dCF2lPCSbKfgovWZFO32W
7+En+XvAKp3a305P22tVVYFzce+Wvh13prHNGnL5KxTDnYFYH1zlAiu/8iX6
w/fssali0Npeb2ShNVo1/Qdm35UCF44jIGJ2HfhGjRCHeLS7GzBkhmUq2hbI
tjSME9nb9KsXzoRGG0FGUrCCJ52T3NRZltTKiIGxlQjFPDoL9UGbQHyjsdIe
BkIDJVC5TZSeZgJr/GY77duacAHsv50U3xlowsCKfcp7buIg3yt24COeJVEF
d0FjcW0OBPaWY0K6DTeJnP4CEr4kJUoVUo2bKeD2lRsYL07VoBgE2BwlnlwC
qqS9dTGyusQTXyhNyMugSwuRf2mCPFlpRGebpQkQqgSfMDa07PQ7NsrXGDfM
ffzWXt5i3roN98D56PGZe6ELQ26YY09uY+pQ9oh7t20QY1pC3KFM8nOkjPPi
y+L7ZX7/GhfQOhyDnhzhLGgzaFbLdsb+ol8GqkOshRn84KXQgrzW+2+H2hnD
x9/iYctyD446nXBx8VTm2MXCsRvScpmxeS3osvvZfv7psfeGBVMO6LPYOxqV
O2VhJZVSavxsr0oFvkhPj8DVvPwyc4DvlJNfGG7S6M9aFbxUgwkNAf7ZwR4p
Rq9pEl4suVLrmmqb2UOWUzudRS9T1tkP7qEpFFlQ3OVJuDVkt/p4+46zaW6r
4SkfGPNmi0TucZwV61y9YWQkT7TkDGeofrE99OP+OqFzYerO/cPylzirp5Sy
uTASh4vGl2zCnAx1zow40dIiIpIHh+sfpg0gpQp9N59nXv53z7DyBUuANzlm
2mWtjcGDioPWIEnCNi3iCyaIo8/xqERnOmojMqbKfRh2xrOs19MAnQDev7iV
p/9orFL9qFzlOAyuRKvzIo52mmo+mmh7IXf1W/GkGyjXd/3yCI10WUnAvrUT
HbqHb/nkiXDm1aOt8ByFB4XrEjGSR/PsJg8zT8srjIpsElTiEgml46+R8N1L
wFsea0jczAlMwnPXbpTc+afTzQYohkTdnFL9QO36a8rbzNc5qLnLVDV7ozmd
X/Il9cSY12PGDxIJHMc1zCeGw1ag84GLb0d7sQPuIqkWqPBMTciPw34Wca+S
gjb9we2KqaKaNaQJPc9jyJROySC+nmISOK2lBy8TXVGj4hCv5lj5w50A4H2s
drjCiYEpGFvQrm34ys6jnmvkj8aqgvjomH1H3N6I+fSqzmsO1vb7tJ1fzObT
HNJSoxme5K9OZbYTTSckuXMDo8psELCVBAr0ttEE4PO1Ez6rYg6cdGxu8qYu
SNRLnTi3CuKBJcFs2LZgPl3mcRqTeOXSKCP0KM/i6F7Ld/YxJ4AIGLvsTZME
E6VxXosaP8vF9f/AsOkpXXJ/vt1wennAspJWRrazHUkwizmDSMlRyMS82IUL
ds5a9bAQMYm8HjAQ0WOF8oz+b6aa/mYwRcEnjtXXvAafh9o2dI+mlEcT0+Sa
7grdzYWK5ATq1/fB5yKCqwq6vIosvRE/QB69sEESr0VX7Kr/sDqhFN4jIIgw
MnVsmr7QwEBR85sZkWxjqUWm2v5r2svQnZbz9mtLobUbZ1wtNpPq0xzoolZi
DiMWf+5h0HEpXScYLTw/VH6ElbiWSz690KZt17mBJcbOQy1ndehp0/JMk3pl
zgoMfmsPh/mjoZ60WvO1BnbbS04XG1upr/eLTWZXPkV6qxsQdK38Jb+dxjs3
R1a/JLiNpT9WbCMhRVy2OtKSGW5ZlmnxsCpi//dTtJNWVjaNBjyDgw/RocCd
+u0/hccV9jn4Be8Mp6KhqsS/uhNVqiDyu8HWQ0IBr3BfMMpS2OKyYvGKZ/dZ
A4LctfYjFBY0vSAyttFLOz5NympjEwv8GR8lC9SWDqx/G0el5ZaFXlLUut31
6Ftojwh59F/vsfvEs9xHDe2XUnV8i0OSoSyNPlneLzizsOJUFiVIChPa1W1J
NdKGwG+7NjrspBO12j3Kc1MQ6sBv2d0IR3E9xgrPWtiHRPtRNspLahVA4ytI
47wLqzRDW4YL2TSeB60WZmb2GHa+xYvrmQmBb7k44pAa4eiyxzUD81TMZtHt
pADiDKq75saFJEthanUJoE3ayujY5U+/zoGPtaZx1uYyNmDvr35UyFcP423G
+qWY5n/knXvW/8Dwh1vA89gAXW8PYn25XjjcWFi7fdW75lKsEjXShTWwNXL9
1OO/sLeYuJSx44jEXfph/mdVKTIQoRzIpGdHQlAN/2aTUmEc/1lt5PDoKsJ5
6PhnFEOIs9Jzky6SaNAnqs4ZVAUGxVLptft0tH7NEEKmzkASAaKvmFUZZD6m
IMoWNfmhWGADs4/s0jtA95lwDfuzJSuryGsYdArUdUc4sKEGBcjCXwQ03Grp
0erXYWeQvqtQbL+gJZO9mIbpXrxEBgtwfRiGDqi/h+f/Tp1Y0obFv+VG+UC5
siww8SJ4K+JNhnOS+yHdfGs6nEFhEgCBcm9YohuN2HYC4s8V5fw7Lofu+c6V
ojdo0CFpZhcmo54ZPmkWipEmifRBwtfy/4jyCwD891llz74oeQ1APHK6ahcW
mNbCTddfgfAYHftFuuojEvYc2UyWKBZK3Ud0wyVKlI4+vaZbZwjJDpn4VVLn
ojHfWeZG01TYuzy+YO4SJHAsZFHl1DTkPJNiy7VZMz3Po+O2jdTKFhOub75t
wNAXx0nJYp0tj7/bT0pKyT7GDD6ynHHyis4kLhhMwCO7J5YbQZSOq2bhjQLJ
tNmBW11rSrRKta3wWnZkrU2IKHWp3gQuT6n8yUhML1/DfVg/Pk5JLhwKKSss
CVUSlnEbQ8mxJOW0dmg30BNztXE5XQA7m/LnGML1GsIKkqZX1i6MBP1awHK0
jLpzxeuQBWMDzaMntcMUCzsf0xa61LVcqlXJmbL+lVGVe2taYvhubCfyzX3w
GseZP0W/0+OCuckRJcAHaOKj/1ZG/ILY/0/7H7gkhTLHz5wyXuaQNJf763m0
xP7UAd9fg3M3GARYYQEcgQ/q90RNKCHS3SEbLzel0zd6HJMnpUWDOW2Z0qMX
4azA+/HN9Xh+nu0YwWE/SIXlrjhf8Q1nrooN+MH96p+mkhQZDJdAeQf/DS+p
47Y70PWaX5TyBolbGKn+IBfoJyrdKag88aMMeB5pyxtjyS/7o66TZBox6Yik
4QuYSjpPEG4Ininem/xYizI3p8cbWAxi2K78CviNu8DjoZ61Ohe0VgV3DKRD
D1Tu4LVunnez1hbs2cJ78sM8pYITRCBhybB2HZYxnQWGH6LuFypFm5l/bMMK
Otc3A7gTq/YHNn0gYYfxrL45mhgJX6Dwfj1cDZvi5kj73Ggvw/M0h+u0IsvC
tIGmGQEXaboGgIhestbfIGW69IqAESKD61/sk0Idx3aV8X+NvcxKzsRe77Tg
Q9gEtHzsYua11R6+zWGhoEql3nrQIlKrjewxebfSdTjFGFn53Rtz1Dzx6U8J
5cA8I9Ctt5bR93PtQpR8baj28T7Fhrdki8u/V4LM1jePFzqjT2xHvTcTZnZY
4D6+/PFwqGuiB66nYXNl/YsElZiTEAHfxXG/MasodLQ1brvjtlvXAtTA3cp6
GFGXKmLDd8XHhv7cHI0cTGrYwluD3Oj62TvyVFRVKO8FlXiTDbcru0B33f4m
K4nQ3ze6206P6YIsMHgyCnbWyil6R5tEOy5llMuQXejF0Z20lfeKMXL1x3fD
E1AHtCjtdaq6q5rDc6JtKZmSx0EAJRBTGryEIT0/wTCcT6kMz4enfTcyF4sN
dxTSLpVNz+wukGolX6JCUOr7+KskuNXYQSdNGdnFCH+ZzmoOS9LiYAkwbUFO
2OuVuPblrOKXV7+hngS+RdVfETX4P2RWfT6Y095l/CBHuMxO54ES0RaxpsDX
AiGHzLcQt4U8TJaz/GhIrNwvX40evsuE7kll/mGLY314kiPAXE3PjiI25Ap5
bPxQyAVyeK3mOh/SVYJTQ38+kx97grAw+diF/kUzrQI+IVMbFowVjCqVLPlS
93yBvf2JS7lhMqcNnWXyt9zlCIh+J1YQRixU8HHXwvbzIrrU37H20rYVEcrM
WpK86JLP/HCFboA9hRcFwJY8IIsYysIIfs1eefzgNB3tzrTw+bJFr3bmCXCg
KFGbIr2OXopVRleHA0Ofn9/wYu49cj1MJ+Eo0BhPJdGVTOnLTRHm+O+aV+42
DBH6UTB+YyNhp02nqD7FUEelayQK7YwAXQ4y67f7Dp0Nih1bjcUx8TRmPAOl
vuN+UxwCsq4AbnOfEKNVo5sDm+X69Ds5w+4RsaLVNlzSR5DkHcl31n0SAAmw
duAYK4AWWCuieEGukKBT/fBIr+Sggu293jtXPNkfos/UONKaAwjuZq2XCqNB
qoxUcSPQ8np3QfQ2OnfxR5UBhUeP/jGbCRK94ih1UdTor8G3R7AkWdcnMEK2
GPZDDoweDACrCiE/R1mGCAENpj2XfzizLypAwTMLyiODmtkLzok0bAgm1Ko8
QaP2HXNs2W4reFm7BO+jNEoPAAryMEFr4c/t/r/dUNHZWwP5dXpmNQXbQ4Gd
ZsI5/CU+zH5FkHHSMOlDPuwxd9Ssvb3Wy9lQeC1SmKrP8FFA6LfKX9ues++w
pwLeVXQPxMrI9U5vchd/nI0j4TO1JdMzo+EgnZOqYwKyO/oceZCjwRcQoPL5
rI3N/3T4ImaynnCYuVtK/U42eln7G/ZCeMf/wKhylWV83weq60IrwUdPIDuW
7WUFbM3QO7JWdnB0dB3STVZOAuYWg21Hl4TsjkdlrXl9na9NQcf4KOZoxCdA
0resawHNxxt7NTvR0yca2s+2xCLHPNMYpJyItwXvRbyAedMYSGHANvyFl647
Rp6ywmUMT4wKOp4yWOuDRDYh6kpNQhnRNHpvyQvsajIxubeW3pjYeslY03tg
Dv3CDAF2v/gKwTOowLDSuumjAtRWA09NONxEC4rLw+Z5LVCBHRZtjznD2QCT
hzIK+5FGTqw82Y+iURxw4IYMPshpuY/gBo3aWzeuMYSqffZWZMCNMUQgsuz3
RJaBB2+fLhxesj+Dczovq3+nuo6dyV+RwKVG9ZtlcbOEjbLvocDoBMzq2T8J
W9BP7YYmQdOmbTX2M2xTMwK3Fdmdpc9MeHDjFZqGFGJd6w4iPyJps7g74dmL
4zt9B4wetj1iR9HVYzwYdYom+eunqUksfqt1A/1oazJmCA+aLWoa00Owdr4M
JuUzfffXU0SrYvEMSxJ2JJTUBHcD73ZhIEl8SF9Cva9EAWPcjmUCNR6yWLx5
Ndg9kK/6ip3MV0P7LccYID3T4JoUdz2l0ejVpoxt030E/VbZHthndbDMMYk2
qYS+40m3laxhCBusTzUr0gHYXaILJ7FvZ9lVbly9uyjxiSnDRiXYJVJEZAIB
fEu8HMSaCrMDYMIUxE207aB4h4ia3U5jg0azKHXqMV83z0t9g4LYK4dGW6WO
cUkBoOsyhVc7+L7eSEdQZojifShpBPcUzq+03o7saExrfTzB4ixt76mlVLoM
VFvqCNRjhWmN/LqYWAm0FJibYe7KNF0qzwZ6UsmrwtlE/ijXqGltQKTNriDB
QjBQ+uAWAg5GEjSVm3ONFdYgXjP8y/5T9NLmGXE2diypbTCwtvfT+Bwx9rDZ
cUdB0DhCE1kHgGuUbTBhi1+31vjEuSHQ19K8bouv1RG+ztKSc0c4HEugcPX+
N4ejuKZVFzXwKIxfyHPAxy3P8dnPx0Zrzu+pCTkEfoEp7Hwce9Rv2NKoBcL7
DE9GzobN3eQmcMnexYqeYMchlYEHUy9ulrXHv6KSHdgGXiASnG5m6oBzdJIa
I8JGWmwWCSwzIXTvbeKIBwey0QW8iJPHUWuYo9UB2MefS9OI3yrHS9f7pX92
N3ffR0rhkuMzOFV8ciIxGebfOU3PJk8r5rtokXcIm2FFTlsek64DJS2OzhtJ
sfZtwbGc2Ko/FOuMysFcEjdHVCJ5KJgzdNm+B15JPdrxA4fSm3dZDqJg0abC
QTL0cTmCRjY9YBpfu6x96j2iWTGcQF+sZHs/0idvyDDXjsMNVZDIfWf1GfCw
Hs8zs1I3N4nsuNBmPqAsFVIiNu89o6mDDET6cep36CcVbWzSFcow1Semqrp+
LXd1CR2wRdm0uMi0zUaIS0kUFStjMfocy0rbl7pvlE4wkfNKBdgbgda/ik5X
Usz5tTZOoKxKI95G7mrKVQNo8ZrVA1si9h81BFC+QU3+UA8qmUkE+oStE4+C
XjxGFWlreMRiy362z6miD3GBN5VMgdBeKNxE/mKLGJ9/OCGqUGQbsMlNLfGc
axUJGD0AaSDtCmTPMfKdA/QoRz2SGAVVwPhioLPk3fSr5GEJBdyvtOa2UYdB
XLg+lcWrzSCiIjgte0AyQ8UoZv+xmjmsVQCYd+cyX4LYohkUU3FNkuCCzQye
/IV4GJkepgVCsYe/eQmAVmRJgWaYOZrDl0WTTA7n2mBUn0n9922egH85X7Nm
DbzHEFsjhDcavTQ9yHK4HNl+eWxKvf471gVm/CSjGFKXdC86Hn0ZrmxHgROL
Z+eOKvi9mvHYuUuMxAqRjoU+elbP4WuC1HUhABb5Ea6tNCMsOuY6d75xlfCX
Swf+vXMw6fVxpJtoLlbONR4yRoqpeURPeJw7sOGqGOPaE2t/5otRz6Rm2Nc5
7VwuM8C/oa1lmmSN3tH3A1BTPFlwtdBPN0X+uMnfHAKSHAxN/G6ONDm1mjZQ
myOQ6oMDerY/mhW3I/6PQNCDV0B7Co/44TJ5z0DrCRYZpQ9+4Dd85mhTA+ps
3apOdRIntB8XeFn96Oq+IckTjpz6+e7RxmmWIFdL9A1rKZjcqgDKJ82YY45W
LV6X88BU+voUZRV3q6+cJgtOQ8PajlVcrt7iAShA7anjeq7ECDl6NfP9R6e/
V9ddXmCi5ebVaEEDR+2qho2I/aRrgm9agQ8uFBXOI9HJOT8Uo/k+yZ0pN9wb
usnYdoG8h1nctCRoufnQwwlHEOgF6yTRjOVVnOludLXL/SEuA1djf1WkA4nv
tiS8+dLPu5TeurgZ1TLZWSFswQtX5dCDt6juJMQQoWdMtmdWSYjrIZjXhX49
SGmXfQBbtEZOQkWSaoVlJpay8/6NSbjrSGvi5+jqb/lkt57bziXn71m42dhc
jWVAVCKjiNz648FmBt9WGS2cI8Kpp1Lwfs77myGGWQqEoJbJ/IQBl9qFSpAq
Wbg8ugeNhrDwyQQbDE3eJRtiVSiTPJUZZUMsP4NYhkhx8EtLmpqvCsrKMdR0
JjKbvlhelNW8Sl9DU+fQekvCHfAgHEgYLz2pCiWQbelmF+NkL/9m8L91hcIJ
AghpWzoLFUriQvL64nBwDWsqX4kgNeokEjdOjcHGMX9V/Ty6jssu6l6mTWqL
pgtYfBp17njjGD40dGyDQvjXUpmIcheiQdRFR9PlMXBjNBnTACl6mtI63M6x
oZ3ayJ4bTRppHVs4A4EVoJkjajdj8gIczgxRKd2QJyXYwiODPBh2daVRr1mM
dc63H6nnNMEf9znYnUqMa7ExK2XPUVkipnAQaycdSElSliZwDcIMdbuqQzAv
ZoOvQ7J4vrhXbMIz8yhskYEkuVIE6FsYxk86rn9l5qVL/dKXQxAYGcQ2CalA
fyodXwNIjPJmxGNIWW7bvKTj0JhOzu9TVUzl4HlVPYF6B8sFF41w9dKeKOgR
AjmX8hx+ni46gahpQuFNk78kxVHGFjzuzIHMhwRjaLHjRSEC4Pin/8BhF1kS
ex5bssYmxe6f0JPO3lShhpmr8tCmaJ3pXX2KhXrYbv4VVEUa/G2qmfgOViB1
/utAwis9cyBwpzCdU6PZ5m3hg6DUerXA8Ma4SNbRthofY7A+i+8uVaGIsT3V
i0019Aar2R+RvFTaZLuHjbhoJy0knfsULiY+yfXTpD1KDYjTY1BvPz2sbgLT
LzNzMywRW4kCwjzc06iJJiS4v+j50l9wd7ON81yugtswC09zCubteSb4t7Nx
IrLW0KdeDvcBEbJSlm8LQqQxuKilqoVGChxSA95HafHwbM+t4+NUAppeD/JO
ekmrlccY6dsmGO+oAqBHG1QGkGseJ6A23EFiHo/yaqCIrep0Mi9zENwwHgwC
AWpJSnRAB7pMTiTx6bk1lRAKeb2abiNhMjj8xFpkx+F0vGi4C0idXpe9epBz
gnfpaRRwgnreWU5JYYCRw8iq2557Bix/VbOEY1a2VxiRrCzHmWkpjxKpvKgZ
BaUvEo8I09kb7B8yLP0Sv8e4wyinWrdh2ZrnWWLhL/cpSQdoS/TsGAjfpJnW
GUzxXeOq1WgU/lZNmWdxcS6XcEui9MiXNa9c6i2TVjxWq3WpbA+0/C6e6E0j
ZYSaFT8d+fb4olrg7q5jE2vSeqoIyh8DHXCCM1tfycowwwUQSnV9nfjoQsgu
1CSzcFyFhVPNZ83jzZVjZH/3VbY1ZubZntfC2wUdd83EKj9t11kswx4JQ4NA
0QO+Y3v93BM23kn9icDOnxdVq+9dtt1FlxtsJ55B24Q6VohsUSDjZIV9mNsA
CDxD1kbKXPN5vkhEuIbh1R7Zplo+SSUQtaCIQMY9PYzFs3HHnkrFlgs0OWQU
G23CqhknzXOxyHE2vdt9WBDMcWKY9MRdCmoKaErSC6NtfP732tjzVun7Pc1t
x9Bg9RFcLlYIcaVxulJgahsY5B0AzeNiEDatAf1CYYcGRUg5NnepLv0dz0UG
IpDHGLRABN189hgIKQQYZX5vEryDwWEy0kavUKZ9pe9Q1kqHoOceOnT06abB
YOQ+kvccp6Sj54CPIUv2uEexuGw+WMV6ee+2lIHbpHZZ6GlUaAxy15iKD4Lz
p3TpVp9CHlwYBK/9T7/wZWMk4nMoB8nLv2MOMo2v6Kvu4cjqZ9W8WGAtP0Sa
dTCZswpLz786Wl7Bl0vCREzleDntA2VCgU87ytyTPpnaNgDJhqfLaJHGyJXs
eI7qrjBlW4ok4BzZlnxc1Kmb6nyK+pXxNJYOJhkzpSawzdlC0sBBzHR4M2XJ
qnS8U6LilpzUgeCiv+1rOn1zxJAuptHDwbwD/Mn+WRGLWwE8YfsOnpMhaJ3C
kG1fDuuOHLtlqGM23tpQd9t9xfRiI9WvwoHFHmFHq8L3AXLWtbZIqGI1iy6A
m7fgAMoTbKMNdvIzxFXJNbB1I7/wCb2k9fp2jjPoDA2s/AbBhemLuheKVKvj
FtPXucXooxcBpeeCoAsPrvm0/povRiFVoc3kyrdF5ChuDCi3hkHw3IfhHqA+
itOaDuJ6OHPvvRbh0nDmlVJAhY51wT34HbJ30imp5se7wvYQebjrNVYaAWWJ
+wI5jJrPyZy8LvBF+oiJd1XEydKhYVmgzDDt4y+NYY8qFC2odICiPFIZbCfQ
PAqobraLL7fUq9bPxMFuPhSqGWx9B/aOrfAIckjCAeVLpcBtChS2q7cBsf/5
wY1BGKsT105o08gLQASwGAWtxzVvKAzXv/fwnwQU86m8mmLGhYUfnWIOU2KA
b20Yp77IoIpJeqyzsyCF/Ab/ljaWTYPSw31HZ7459wAyKCG+HKXU6rNb8rf7
Vb7N0NDkniybx8LwbxJJHq4aKUgcKZNT6OkihpeW4aNcdH0c4YylYhwJpAEr
6ovIA9YDfDXtazg9VbBed2xrKdMIAdq9xjKDw9DtkrQOSVdCOW1AG/SEd3/h
UgIdBPEL4GTVpZaMRWI8sL8wq7r1v1oJ8PrlgZ86i/MWbQjHtGSGnGJNK3dG
17YN4c6THTR0i8sVfiMfLCXY+L+2ERlOKxuZ76S7g1u+Ez7tGKTi0yItg56+
xIc3eyuSjp4F5eixYprnZl2mNeJrEDHlkFgcpRKnjUwUbe/0qhkH0N2iX7Oz
4arnc6+mzJbbmin0ynosOWX63PjH7X3G0iAxp5DYXCCqXCRRvZaHYOUxhorZ
sL9bdksLkRwHclKxk456zL5W3uA93/ik2uJt7QlitK0H8D2lj/G1Zz8Y+B8p
CaoyRr9sThmtSzPn476Px8PrL7N3eZA/Fjr8grkS+GyvgvvgG6Kp6OXvrV+b
cWkG1h/4vZ91cB4A0dUUalszog7hAS2BI41mfX0BfJEVUEQHIEMOWLfmxJ2l
1osA+lk92ihX0PpnnPlWe4SxaJxHsZh47P27yFlZ3y/a+JoF7jkUGaZO1HEf
heEUxgIX6vB78T8hXi38J2jHwHZIfLVoxTcCwp+g7mjjrKszPFgxHJumLFcn
mILHYvly69ZLw72DEgylSbIcM7Jqw9E9pqZubElKMIUDLU9/r6n6+Ge9ujqB
KxygM088ilh7ecT49ijZX9OAArVXEfq5FKEE+p5CW+pKg6sedHEnUZvNYnFT
i+klD5fR+2uWQSY5ZR9mowj0HsAgEE9WSMgYO1FPNAiB/SPA+8Qgl8vKMbOk
LhqoLGHkFK99SjJT+KxpKN1qss1zcsnWwUgijoSlVtY+HWUNE5oCtJtIxXsk
ruDo/rEWqQ9vd6HvI9qz68p6BPbX71q6b3qYRTfBDV5y4vZZZV68V4LmrgC1
xZ4As2D4fVGltaE26ay5nDRh7T7imQn7Hryb1H//+4aNknf4Rowr/t7owd6a
vOQHlgU7FUyphXIJbe7Ek5f4oI/wkLqNvdw+u/tqKZBg+r+IuohVbNEVU2hm
h8Cnv1p8nTleyO5AHSugBd8NrW5h5vqUXxq9UICwE/fb3ajUF+7BsS1qd8gY
yvzCzRqaJMhDSNvQDxg0X2ZC3zd4gCjwii2h9AOvujqS3gr5FV9pM0YnEuOn
hD+qe0is3PovyCS1ZnmWtSYrHiBg7Clpbnih8yG4aWihMfBE6G1QHlf6IoFq
X8B9HtVOARF6bxDDSj6y4I4zXzd4jn6x2MWFkmK5HT1r5DvE5pr4SF3SHKYS
9KZD3tcvFidfmZvu5xTIxVlfb92D2OqwYb++DZ9lOM1lShKOxRTY+GJdByIL
y9G9ApnEDFy+5qvONaBoCo4N2Y5MgN3Fq7pO5iWSyx5OPJAehvuDE5DIUTQ0
0UJVawQH0hpmcB1CyDOOoLr1tQsxoZ7/Yi2nPRaazJbHoOvLLLsOfExCqc0Q
NARSk07bA3WdmiZtL9bKOJxbJqXBV78NAUyaoWGurr4enpcEaWOWs55twMRz
8yl/vbydOlfy276C6owoxFDj6jOQdD5SSRK+8CtiAZ/oQMkMrxaMx3m/188G
PRC3daev32qCoDYrphe25o37B2IvwUwnmfXyy1xRaM5Mp7UyEtb6XiPphNUE
HmpjXIix29MNllPgl6Rp/PDkcy4ms4lze+nH/Nw6Ztaw2OdOIZ1T/hIT9jkW
sGKobYrDi2D0QZe+M92kvkhsSqXJD5LjeZuc4nMyhZfpJz+Sz55XURVoDiob
SFvC5+0OHBtF9TgF9P3jBZf6tcK7I4Y+25JAzhA+Nc08gN/MlbxxGFmmLz4p
dlajLUlv0bdueinRDAUKan2LpXXfOU7DwuKcRLfZ84tiaOCGdArJ0GUAVHxG
+kWli4HZOzbyIkCrWRAky2Vjpd+vBo2zYchBDdw+zKOAt8/OEQQgFt2LN0Po
ul/uWqg/SkFMdEhyFHGixqKyKXs0lio7z+aXaGukK6RpwK3kMvvLVOGezEGT
ouU5uRYz2DT5aw8evP26CuXi/a/S338dK7zD+pLru32tg5gNsrkH6ESpdxoa
bntxLuUP1bAplvS9W1UEh940HxslrT4ULZX7wHH8aK3sCXLEpQYMu/ili5hz
e2ggSEUHA8nrBodiqwxpFLbpUX9b+IV/7XiJDQdMGNIAb8a58AqhWvha9NAi
+Ft+vInbRWWwn2Ki6ovO1jFpgqunUClkatEFyL4G2pu89jWN3Hbn+8ikjfYQ
TdXh1vwWogK1K8WRmLxH9J1B+3lX2dTVtWxS6AVbYlsdoVvVeIUmA/JUminV
/EpSw1ym92Z+iQv7qnoAKHlYXk7LmAzobon+S9et7CO5U8DuLIPr/vWY3Z5W
ohjqGIR/M3UyEiiz3wLBf7FvuQ23xsKXooBxoGtox7EEDqnu1g8Cc8pU/qse
94HEJuIdsFxL91rMlO4oE+FYukOlt7SBbqE6aSFScAY43TWDSQKhxnin0wfX
2HJSXWZQzDmWv+vUOlYorFdexdfdr302Ju8k73nTnFNuSSYwiRXAVISEtJM4
GX4jgZ+nTC/+bbbnRMEQaDQK5PNjEKzQUBzhEeQt1N71mkV5ZoQswCvCAT/V
/hR5n2Ls62P2H0yLhsyHBzxzdJuHq7ONAlNa/WU2AGd3ACFVIWVQ0vYPOXhZ
LdQk0qCT+Q1BzjQWtbPv9C/SQoIJ8d4Vf7jZpvBk1oaTw5xza8OikpOEv5yi
Ztwh/GlvDk1KjCZjlMORfJ6s+OaXQwsa2MxuAwVYxTZ8s8FwGhm5+BuLDXD5
LAAt5bnV51ZauqhXP2r7z/aUjumy/t4mCG9oNckCvLHlimtIn79Wz/4ZifYJ
Dw/zMiyWB96wEq2XVb3v1A+50DAcEqvZ7wNA9CkFcIul+Y93Aa/Ttq0z0cHR
Mo/sr6e7g4/of1BTslmFwvjHm5myq8zfu+8YzS+c96vl2wahxLaXBGu/rnRh
kYbp433DctAi/Z2zFYVVf4moovqWihvs7hImRZamaGWWozfEDJ9ebi4B0zz+
DP9b73ZIr98JJcj7Rfj+qBD8LFqrmHuaok11+SQR4P1p/OZUZpqXP4oSDN/g
NeBIaJWpOQy2mG2XpUvrsz2etB87R6gj77Z8nRbH3zA2/zlv76UNWXgD+knK
cb9LnNZcrNgTa3f8n4ceYEYX+CXT8KnweJdFDqZMjObzrbgfTTrkGYnk4tqi
/zm0DJ3FE5oS2yT2HnAoN+RvyyIrmjtPZUwK9mjRzgbdXKQJt3PjRXK+5Rgh
FP2J3lUDaf5/lvi4+0izG4wDaBa9rpmxLEPNc6Q4cgn0L6CLGLOhAXCJCKyC
cmQ/TNDCntSWsLQGMW0oRBgCC26Jw5aEQrVEDzrIrtaiMVIvIPRinPYkqeAS
/45l7Sf9Mjf1nju9FG74RwyYpzABoD5YGoEa921x92Di3cNDJpNSMI7AYJG8
y4LB4OkkdDlFvUsJPNs0NYDpblwQ7KLGu3lJKf03RKFgNb6ArnXuaTdSyHzV
D8rOjpktpoYp4//C6mjHOLzfeySUoABfqZjR6YfMvPFJUY0WE7F02ct81mr6
BxKf8Kskjl9muEzyviAemKgAGK/bJiXH4Aox+zD6QmM5TRz8ssVbsrQG3pnO
X/lOA2B2V38u4JYh5suFhw8lJ6dHvWyKqiqVUmBaZSqxKFjNXUvpc6J0+KKk
64KEn9SHnRtJa2NXywYiSCfFWiyfLDwWCATCeeWoVJJwxJ4Szl9qVrboFRKf
0bPymqJuQ/9e1IYSUex/8KDqqlWO0qiCVeolZbK0IKpPGIht2r65InWgfAHN
W3xzUyozCyzbN2txXYbewlBvuAxsYQ40qZPvif1sET7eKxsuRY2n4tJOPTir
ph4h8SQRrPVNgPWS5Aq9Vvt1KKeJ56dlRrIhvsuaAVE2WdKW/y3tZp8Pinfl
8mREP5N50AHdC8KwFiJ6A9A2njpV1rF2N4rqXGg7cA3YEile7dRdeHBOcPEc
wv/NwngsbPbrCWGXy2moSlQn3jacL22fzCfjRxsVb9uyM9W3elzF6l5SUz7h
uiu2AdcNFpxumxRvUJ9esIMTAAcFLYRYbRymMbttJNkTnFhcx6Sun0eoAoKF
JssM0MzPcjYxA1SVAuvr3ljSUDuN907svxFx0J/e1hk0PWGIJ13FfHn1zMWG
10XsX6spOr68jaLOONyJiXFy5Ecj64ZiDAlDl26aikk6GdFcUZBTTA/c/lre
N+DPgzFS+EByu6mEUKFgSYqRfZwPhJmu8/W+caMV/bYyiUtTphdr2hYzY3Vo
qcAS/EvaOu/FQtyC87MypnOtZqpZliMNuUXk9mvfbyv39YX+T7t+vVjLe7OP
U9RnLknWYGB43Uxm6FyAHEinLB5B9qIHWztn77Df1c+fb4dStvouDA4n9sgN
MkkhCBxGI7R70f4z3McckRbINJtzFxvq8QQ/3XrfJ3SvS9QZ8UDcTh4/N70S
AF6EnYcCLruk2yD1SMHALbfxwWxbXgvy46fXWBynRtM29qf8v9O8ZfLU+uZV
4hlQ+LwqAMTeb7c9LlTqphl5dmAaoVV2ct2bx/JxeNtHgrQ4bLaTTWXuQcpg
GCTyBy/gVScWzqZZGdZ8yUXb6rdvEq/YkfZI24iReGE5CQ4zATyb0/DKXXzV
q7hqS24djn9rQRUpX//rYjMaUOEFpA34pTy74AVbWI+MAcVY1mZA4p5Y+aIU
uS4MTHcnwg+yS+aqFcpUvEwIn0rJ80iODljoU/+RATzxje3SyFhaGHOWjUln
RcgJpJIsupmJIY3DD8xp9q7TfVJXxypJ636QGoWHzzFLvx0ihGHJ1qRCZEg8
Z9yrXkZHQRgFsPVAWTCRr/bg1S8UexADCOS+GMLjx6hUuzM3GISVuxYvAWgv
sIGyKXjCXOOMQoA+XNy/lEJGwVxcfV+hM1VnhAvL62Yo8/+bvNC5YskGLR9l
ATFiT9HxOzOtYLaEre2MHZuTGFsQH0pWgm7LU/gA3vx4U6Ru+V047zQxv2J1
6E0UTA2UBhe/MI7ab9OPNCRair/+4sjDj/LgHZ/OBfGCXnMQZ4GwINpRoVno
oYQMa8s5ewBzxDP6Y3pLSNrg6RNWSBHvL0WGAzy1c5SJCJyRj/KqcboPPa84
vIOPjgovk1gUhL2yYoD3PNApXQjJcLnmjKB8VMhY8asaGUDXrzcoTsPqi8RR
ozhn/wGLeSDqcT3+ImmQCI+KEdTLD214n6yNAa4uPnssz1sjac2GHR8W1Kao
TU85vVvEPCe9fPaNI8gpOUb1Y9xvx56hqj3H1yvWGMchL8b3P/A4dcUWKprc
8KcnvMd8DHvu4rUgrHv8KfdP07zD64bZn2GE8YaSLKyQw7Zq6XM123m95kGl
BSmSVLdFCtNrHl7cEAxk1+EdvorCI77Hwpsi6HFeuug4mHX3d37jYSvTsDP5
T57u0kDOaq2cwbFbyP/y+jaEMnkaFr4PW1N0D4LDybJv/BROiSfZijss5q/r
WO3BM2LHx1i9Oa6W2Aokg3EeWSqiG4A4JxNVT9s79UBbFjGVxzlh3LOzWcBn
/rPsdXLtGDC9fZF4OBtYM/bh/dOILERTv49KjWE1GFqZJttEvrFb369Eg6e6
7OM9WrOSZVWX++h8zAuAqsuIKPpU0/+8ueq9S1J3UYJls7VGtdpgXJXZuU6x
Wupciu7HOBQVieBYtSy4mivXyV6h2jC2x8EXTG+Zmqq/TGxFyFZ6ezQyo1aV
tL6Iqoq82oNuYdCwSsfKylA6EkFGZ33LkmhqTIm/o/KGX8cvDcBXKUKzmR/c
T27aOGUkuro1jXzlw+SLLK1IgzkY0wxYF5+d0Rm6lj9MOAvr+Bgs04lGsNAB
cf1MASZjoQ4KmIlu3DQCb1lk2IiWW7anCFLUpVgCoeR9hL+DgNz/N+ZOebgz
kxLWTUhKeydEmgMVCYynaIHk7EcepJ61SpI8cBAcJKQeNejnj8dwraQaJI3N
LofIl6oNCW1pCRCKdiMffHzw8eM+t0fqHgEghCk3sh3VEySCCg0U1h9bv/rL
WuXxbUugBkrY2g7anGzY35viWDfhAPtt4vuMT5E460F/YuxCUEsiWBURZOpr
qp3URg+HG3vNXuWHaZdSXoeaRj6ITkhz7NuEJa4Q+N+A7BcbDe7tZM9vOKIV
gp66ttm64gqZ5O18CFT9QW5GiCNML5eaJY5xAdk6cu3pukh9LV338PfFL9Ke
QMW97JwceBwMPDpvA/hSRUmbY/6Y8Z6m9bedbznn8MBAgE0Qx6pE16QPwUUj
eax9ETaPy3Z7xGMs/Foe962fQbY7prNP3ozUbW9ovzHm2WbapdlPevkAORzP
ZxV4pGbyWyjQctCMMfC2EgduryKTu2pou5M9Z0DW7QMaxNd4oXmkfdQ8qDzQ
m5MERd5s2Jcd3kDVwPE8+8SQWhBFwBumBTp4JgLyDZa6huxlhNPR35IvPJlH
0Ynx/Vm+5A1o0+UxVmyqpVtsJcgzAMdeujjmzp8w0nTbTMRTwlisbWkavni4
ccbBqRSZaym4IpMruc3aBKC5bj3n9idDcdSt4DZgY1BhH/IKxto58FYh38D3
sD758glg1VyfH2IpfwxWHS7ocmrjg8u9MymoyEBdnUH2wc/hUwTfeS4stgoU
6eNoBn7L737pBwbINPY5rEpZMp5iQkc6bC1kc3m4yKvj34IZS/WrViJG389q
LZenLms/jSpQCVMKY9taM5NsZXCQpAOEe2nJhYal0A5DbsvnBEh9Hr8LohmZ
DphJUSCV5L317NQfY+e67BYUiDWgqegMMup47QP4dx6LshmJArW6K9D2vTUR
XAgcwtltJn57cm9oO7QDk/6PYxsSb04lTjSgobCOYEET+54DofI4793r7rnh
wGfUEzsFXtLaXrS0hi5g14GmUOhiswbs+zd/4cpp6RgIlbb129LOpVuZg60m
9zF+Z0fEIML4GvbJ53Zy8MLQcgIlxBnJ8+V1bOJ03LtWGeW+TSTkpmdB1sCA
b4MjirsoUl17e88RMDsmJNqaMFW+q08qdX+NOTRTKUzJrKsOZyVvicPBSUIB
6bqbmpi4NuGMjcD2vdMZZtWC1/4ecdohDty/OgqJPYWt5MBTThDBZ/B3o3YG
VwOvQtukbw0+/fMVB3l2QmR9ygKG761VogK8JFQhIenhxhvYIw/hNcFBBNgi
ANo1YXU+Jw6zHVs4xb6mBHPZBf9uzzUNaabqCxynKyN+B+Ryf91Ob5qa5IX3
b5+saB238vazst9zzA+RhesGH3fG/LJLvSKfcgzelKxBZYstDeKo0r1YWHbJ
do/lm5RiPSMMbKOjvbJlyanj7/cnyirrjRwNfcWetJgUF/Q6hfpSgZdrCOKE
x95O9A47Va+zYldDPdvO34OupkmOjvfjv39FZioLh2t75lY7D3138f173H9s
P+it7KZjvsE9QoJGi/0zelEqjqOgHwzEHvxZp+cjzgPgBZUQ5ilskLj+FAD4
PSxkzpZZFQUvTSXCsAw4dFVxGvuxz3IB4tQsoqn2sPipo0s+qTIdCDmK1KHa
2S6hoeYtrdrGlP8dVwhRt1zxlWXMVEj+NlGh2wGbpsg4ID04kGD2NScFOfLz
0iSnH6rZI32MdlW+Pl9LVpFl5kpmRPEU3XyI0qxnJFfVh5A4lUlVYO2pZ7+y
XlLIRnD6m5eZI12VyieThBP6oEl8reumOT4Rc8FAlUpHt16nl5FDKdoLhIDt
pv4hB9VqiOVXNCh8EXTJyoOgiYxLfE+LXsQ6hGlP/qj8aOt3saLbEYRcgUGL
Donpup5d2stKM6LD10Wt1pNC44KMmiRr8xPfso/8kblM/xOFIUlMbkUKCKmX
6WSftpEqQVtQHMCw9XsFSswUJUN4NDKv6P3S8gwPlWl4kneL/EutBphiQTAf
/uCaD7wRdSMkXnrx8h9YA//2Aw5CJ6XFBpWGyne1iSOCRg7DOpX/a+EQ/GHF
tJXr7KFrl0sbIusDLYrqJxaoOHl4gZbO6GQROKTziiBUaCCyKjPdgMz4wwsJ
qW0DQ/UT3pdK49jq7SSVdQmuY2WWgiQ+NGkG9vre7ReureBpdzw3OsFyQekF
9IVfanSZvwTPDezwbLphKSCERAP5tBavIsJDSH/1MbRRMZ/6QdcCzSOsWGFN
wpHAhhSa5JKOQGvZH+ZJZVxq+DVDttAHC7eTWWbyKcQ7eZ2fNYpW+OGexgjk
JqseaGRLmXmS+fcNI77Y/ci3XD+dFIIT8PNzq8gg0oHS3d0mD3N6FzDNvoq6
PF7PJej+b360gmEiMt8nR6NSPmYF6KALVt2bbjc5ah5H/78co7y95mHruDXE
qQFBJ1/Xkc3cgqW9baCkGIyM5y5+9WJNDf2naqZ/Jym5aZxn51yWYyAGfu1d
vscvdB932IgykTl/yhHK57mmtK1S3OR0LxiEvr9X4naScH0d0+XE/xOpy+WI
JI2AS05hpWROh7QynupwD7Owt2yzfepbFMxcHYZrwUm4tje1I9MHX0e2Hlox
jqYDjs1jnmFw/0HC3FHt2MhdJcKBqGmcV9TIPdCrkkxcmDuGA0EVyMRDDDLo
nU6fRRQLElwj5bnpSFnduH8KaYf8O/eZj4zZSP3fgKpLEwzbwMMQfwQAKx0J
5ZKx97mYochX+a+gRu3aITD5hF2BdSZptNaCtt9Z2GR0bYTptyh6k9mNWkdl
bnFycL2H4hJV+BgSa3+tmPCqhEQJLKqV0ajO8TjVOutlXxhAe4LtWvL9+aNc
ydXCMYo2xvuhJyxZQ362Rc9KOi2I0ItDNoBzy3PBEOJN1jXWFyn+BxPMDZvx
I7bXcOj6qTv/FwWKdrHJwx7j527q3Y1FV/v4UV8RuNvrbDgKXdlHuIDWD7nA
m5pRnN9Fw6AzLro1CeQ5p5QPLni/22oWQ9cp0rLf0BzbUWas8LEMwAZ3Urhs
87RlPxhEY/e3Dzgh06jKwHo5I9kF5m4bq+aFRYr+2Yjdee5J6EuQ6X+2dDpr
fvqRqDKvacK9DF3C60QEv3POQrsmAM8JanYnoANUdWVz/UmbpZMaisg1OA6C
EqTAeN+Ghpa8c3LTMtZbpTjWNuBfg+CcAu3D4P4sk2+0xana4TYxn4iQFdAf
0GnKKgoGtgbSIEPqfmjdVoeRxrpX0haxtcwdz0vZvZZy90AyZIF8aIltdeul
ibey/BQiesxlhm4A0w0CnfK5Pncr/quDUtsXRV+MmtjC8CGcTjLP+ZgSQ6fY
Wlzm8zwPidPCGtdcs4U8R35wCFvKij4iCPhzhXnvVZyucgqQC6JdqYzvW1+l
2SIs06BehqXhYOhrvmxkacat8EhY1LHinlBRCNzrV4aRWRNPUzGJeLwRl4/C
R3meguU0ptJ4VRoEJUWhTEbRovvEk0dVLMIKKVraWcbeTQ5qenlx3nDUPXvt
JIYP3L09S36A6gx0a7MCcWyWo2hnIpzmBPbv9AwWp0P1C071theW6XFF2IJa
dlQlPfcnkL0NNwj0sGBsW+o6zaaNy3T3P1TIy7/1YE1jFP3HsGzmeBc6XamH
AdK2OmsI18l6jT7Rt2l8TD1wfMYqL7GywhcZmH/oIIW+uH8r1jHGbz1PmAbd
tJHWHO3RNy+ORJBJ+VpQw8u7NpcTfOvbhV1wbAO2Clr7qI9E/ilEWewqPLlB
zEhK/Fr5wJAwcuWhTXtDmDh432ipxSzazaD+hvRT8XYdvX3FWa3XQvHyLco5
gJWqo9w49JufXu44auLn0z4BuS8nLxUh6gGcxCzSRNRM0qa8Bgqgw21KjqzV
NFtp7VOoxRIS+OD8XbZQjfiaFwOXPqs0i5pb1AL2H6jENjm1GLTzmDEklv9R
bw0arUEGKmxFUMPQG4N55cWpr4SGBPyQHfsEJjYnnkajP9aY65Fmr9ea6zpp
qHMH+btrPkaQEEBlBUgL/mtV2PgUvsQtAGplX4sbPnizsrLBGV0LDW6tTx33
Wu57QZcqLDBo/RLiXM09EsQBbaJAB2fXbUGPNWAsUddicbImwb30syZbpVKp
NacO9Zov01DBxM+Mp3BTp6N440l8TWZnyrTpO6gSzBxQhrTO1827R55Y7kWB
nx18gBuNlMc/lg8RUQqdFhxJJ3Md2vT+HZOcrMrRBlLxVz4tmGuyJCxtB3d3
tb21XM/uIQIt1pCq/JS8y0f9dLxfzKqA7oWclYmok5vSEVk49ojOuehyCGUi
r1KCcDXtvKn2nLoQkzCT0pqo90F1rUEK2NT0KWPBaeq69E04gCz01IoYc05e
q8bKhH1UPh1VHDroTXigyxvI+m6X4/IKNCOhs/DaN+R3H1+CNqJYeYnbU7rV
uFfoLAceGaU1rC+NpgFH5ET+ZX27gcL/cIIAJA4AI0aB8G8HPFAAbFFXzmCX
RZmvjBiE7Zz8AGYXDlyyjDc1yimG9UVWVDlQYcxfJsrejCndigk4HIBnCoZO
LE6WD9pTL9YD0f2jyO7I+BokaW7WcktFWIIABcpPF5wJDzCOVqr4zCh1hd50
ONe5CorMnFINHuP7YGkAKTI9sNiPMQ5Hy3EFkT63WIAjotV4q2Sr94I94Sbo
8f3V8h5NoscT44NTYoTMzUqXzOXoKclwV83iGLwkScs74T0msYESzEb8Cx9y
grsykB4YUO2GQgwdi+wCVQZ1pBj+EryoF+8UBzV+F1hCK+O8K4qRT79eGFGk
HEI1Zf0yVnh6frXDlQbwNvY5+K388aosYpOU9tug7Q6zs/kgdHGkbWh4RRpH
WOzYG9cLJcA0y9AV9lbWTr07RDNRb6An0GuJ93qLJKifK4usWU8P3iXIc0zl
kj4Gs1LaJD40R4kqayVc/WSeiMAzvarT3Y1ViOfzR4tH+PYBSN/btFgQqC7t
teqfEIVKpnJYkcs1oeBI6uVJ4AiQbMRp7lYQOHJNQF/Ozh0Wf4qTUbXaqOcX
0zO3izFgQAz3p+KfbdvRus58coenkpzRyaxtTRr7QLKdSTEVmIaEGVV077qV
Htm0EqT3SgSk1H642wGdMVLBa6eQTCx3AB52et9My2TC8HYokRrusdQquCa+
9/PjePJ7mzMJmjT95xIf8YhUDfVVR3pOBaFjsjtS2Mk8ogNi2zR/dZ6hvoEI
uy9DTFU3FJxKVzp1qPvrAC5KhzFfs4+ftB5/x4jBNjUTL7VS2iU9jCnEnIDV
3B8fJCXm5dQGZBI5A7gvnSz7cug2CkwcWMixjQ3BTPQL9XKlSvhD/qRZSXmV
5wojETFy5cucHoQMnidEAh+w1tkl65q+LAChA/5LQLfEZzj2mfCuXZcnvS25
1kIQunP++LhMKIfzDbqSp3XsxQytzE3P4vwPHVibnp395P0Hv4zy672XiHXm
e7MvhwtjEMelP5T24G4BkuOVDHsFStxl+GHau8Ncxzl0YxywjPrv4t/rqphi
vq8VGvW9hY/zXOi8NDN1QaymDNve+cugWpmjLH2sRdGdTFoLW3QIzX/MWrPc
xOzBHFDcvuFy/dqxFM8GqLr64a93wyDylEMXK5KOp3gyNc02kAdxyUaA+itE
Q3TKn1H0/drONbSWBpcIkWInoKdfwoOpZtw9jrUdd15c4wzgCoNzUTCDfN68
H1BYCNmdRzHlB8gXXLOQkur/JTeveKMiYTo6KRAwOJh66GC0p2NI3B/jw8XD
pMeYwms3TWR1bx13TgaFYbdsYqJRnZlXb4Yv40s/Jd7G9YpUZR/2HRBkzGex
s2KHjMm/8bnYFJ9aE/XX5hmqCK4p/DDW08KHUE+Xe677won+wU/dSyG75fCu
SUbZz4CPdZP30iUNCU6gWiEs+2gXclXGhijXZeKzMhHf8AkcvQ8gKJfWFBBa
z4Z4paYPJLut7XPJFUB9rp8DfyDbBuPwLZWLiFsRB+6TbBJDkJ2H8h3IHxBF
Tyzl9CFUHTfjDo/30hIHRXOIskh75+9vApTUTOSi0ON7eG9eohksxfJNFqJQ
W4cNqQv78wKW/yMP3aQ/5mck3c3JAngjWikU5JdSysT5Y910gNwB5fI+su4M
pmLOgmUg3APAswqtR68uJjcJ9ZGxMjDsx6ahz17NATCe/YI4z5Cumg/6ZvYd
N2x4qXvMpkLA1/Hgkn7N67GqeqjsZdXNc8vR1Uk7/JeXKNSCyCwquFRrl8GR
MS7DT0/3IRbiJgnd0y6ffi1vgXIvCrosq6idfTVh7rjPmpxsMhNfjxMAoyfM
XBOMG2g+NQcZ7dI4HnBYonpATIWZwnMOyjCJeze4uRgIR+DgNS4IjChDANqO
dDV7DFeTGTQiUSB5AjW1v4uDnuxFJsZvF6bcOoqe3GLr7bVoIGp94PaGdDL0
TLxSQicKLx4zSZ98dEQ9JIl1rwOG7Zd1CEpBP9qae+TqlbnFFDJJQvF0KNp9
Q2B5XcH0hQeyafN/BvwRFgYtjniE4FaVe8KTd+oyCEm+UYxkCebwwzUPfiIP
xOKUYJVyLln6/GhyXUlJx4mCyWDS2pbxaKU+jGTCN6KK47fQxO8DTXqDkx2U
M4Pm4s7TUI7xlKaccvVSEhqxkWbtPuNYjOKRr3YPYoOjzZe+nyJGsJkEBAXJ
ZOKd1sRgvvehMm87caPwgYaXbN/+fnCJVQaFPV3Ppw5tx8lqyxYdLv0N9jxG
JLEya+Dx+1wQ+USL6ziSzFLbUolOnHXBdcUAu989BVFnIIY2Ljjl1gFeTMtw
MjTOb0RdgrNZP3uT0qUKhKWNpjt4N40wFEbXH+PlnK+C03+F3yrxccfAl+n0
fhOy1je8hrz0IAH7jpK2D1ei6YSfzWChUJSof3JiFd5mhGJIqgFFU1yjdVe3
PYgcf4+iSoeuxBTJu11dGPFRNeInd/ISxAFfDNIZccVXqnssK72LhPfx0r7M
70w14koV8C8X/0lwkhHoZxEbz8wAeFRZPh6Z7+EFp50aIK0J36JENvR8taSj
GI1vy/A8fCOA/vxnU3xWpgryrm1bmYYaXPFrsFlqMHbJhVf6CWiiXGWXRcxC
JO+5MZQmGKuxq6Sm0xAvFqOioBTn+UW3daFPyloPfNTsx7H78dhBQchYJMrO
kiehZvBddS/3WqYWxaUEdGmzRFyiR+j4mHJHc6dSCGuc/KxvP0QNUDU3XZIw
ecaouQxOzpjfkCjsrtmRwfMrQYpvLenUiD0bStT8uF4lgPz/2qyX3xjBffZg
4eQYp8n3GuGJVKOzzwgO6C43qGNFt5QLvT33YeNczmV8iFJp550gEyroQ8+J
BIkzkNZmJ304Hl/5nA6jdvl3/NdQlLeDi0pUwk9RzaunoVu7+tfFUpZIAy7N
mMoWjxpuwH0mJyQ8WyLCAL4reW2+bsjCIYnx7m8kRNhRAhXPIp1Zw1WNJByJ
EpiaIe5bFWd99qDzAuuKT+JbBmrgHGO/InCH1OgUXmbjbt+P2H5T2TVhFxqE
7xWaB1XXE3yxTT/aYPoGedr5psZmMKGtA6VtDDoMV89pn95ZNzb1VHtnntP6
sjmmBkTYo69QJA9VSaHf4ef9oa6uevy0ztjYSygiMv+H2u6QxpM2lK3/gP7M
rGFuITv48pC2JafeQJJT8MDAookKGctoExp58r+cjwmXy6dxXpGQEGLlQIys
F7lFJX9DGJ76Ln6rGxcGyK/hhiJSCIYnNS3c5RoXa1SlMBvVswFNooTNsZGG
R2TC64tcrxqQ+PqTM/WgWxKJ6yZl95+OS4N3ALdLqWnX20zB5Jtv/ALcVIcf
KlYs+f43VtCAq0M1QfGxBsV08VC1OufovC3+vycL9SK6kLGQz95uaSXmOCEz
Q0Ec3j2XwDDuXk9JzdpHiys5wQ3goyIlXLP9c1bG7rjmq64OSYJACOmTtxBp
x1JQkyvdne+4pPyZPy3meAmDIIg7nR2HqP1LsFmVyLdi+TI3K8E5UGtedudC
IMeg1wlOnlNDILii1+aE5+bR/H7ocDS+/ZqReyqi+vT0ubP+Afs5x+xfhzFl
wzfOFFg90OSi+y0W0eLjpsQeYtZuPqOXmXRZ29ftLCCRYPZysxattcTRud6u
ba7zahEvDJAZS1pKduR11RStqMqlDTL3gu4WUxk20+8cuAyajL29OoMcYzNz
juVUE2zrcB+ZIuXxY0b9kII2cTe3pQReKl7J7HTGHAtFCBTae4ba0g6wOm8g
4BlJYybBULa24DoSIeLtcDJGVGXt/LyJDkz0gmhm0wz96mtpWXmIOFAw4SBg
IFidZL9Bq50ysMr5kZZZaVZZMi9G1+mVPGboSag1T7tTlM+OPqXItgSmBWuP
shW/bSuIUyeo8SzlJK00FK9EaW3kI6IEqy7WS1FtTT1zRCRY09U5qewguwEz
/kUjRBKgcoljIPmhgRxLR28dO21UJ2ZMmgQJaPjErEs2LVntDUBz4F6TtsOU
vgyYZdRWV3C8eDCq/9X4qrm9s5ga6lsk2QWNtVDl+4Dzg+qzTjyqYAyntJng
71Ufo7czQRAXZDaQYQJxLELnjCWHv11pMhQ4Tr+icaZLedfsBu0tBMni5aep
O38Ea8+HkEBdMUbByAfzsbpfV3LBJAScZoIs93GJMSGMF/ztpCNJ5+exdtwD
/jEZB5MTXycqatXdyb1q3qtql0Fg9RUPWVYYDLzkf1Y6PlS6sAngZnJsOeuM
mZcDEPGOefMQ9NEEjfvNoWgIbS+l3zV0395PEsUVfREiEAR6Pt92ppw0TABO
PkEZp6/LRVwS2yXf9/3SPwn23H6GRgdWoKPWX6QqvCO0uSkEzSsesP5XZxK8
Hpjl4VNIpNrS+Hmd8KQwmbCON/XM0Z3P8cMp0tDYZoGXv0eGQ+SeuLGAERbd
L0xZuhK8xXGR9V9m0ixU++vU4ogJYs4/t42+WVcvEaqbLf7tWgUHYc2Ce70I
c2IRM+VOF+tyKNmR+yHmYCinXFFBTPRJxulejVMN86740ecH+HlirVl/JMEy
e1DtDTOo5dCII058cC4wNHNIzN/cWUfQHjUB73jQPr4KhlYFy3Ok+nBdYI9K
g6h9aSbHhpKGy0ijZOvrx2c3lq3jJjhCKzLtigcr/5jG6yUQOp71VQWOiV2W
WaEWvtBIfwBgnwrWK9s4b2p9uGsRYixWB+0F/YsEvw8QrxSGLsEaXppivSdg
CHv9f4kSy7pR4vd/XvVlx1UUQdTYf8S3lJUl2iUCa5Yye6sKk382p5taCSlg
L2zu46ZRr95kA/bo1fpQLFwGEbs/cjhgIrYmsaze4nouIN76twyQVcOdyBBw
fhVqpDX2v6Dl69b5m25BOo7cBP88mR3zswd6DIaVbukeytIye3wGxlzLaePn
ldubXssW774BeQ8n7/WUAHBpIOsFupOocpACT+g70RSfTypnVdjSWYiV7xby
X0QPL46oYwBE9fP8JqFVbCZqeLRVK6bcWoqCOt8nxbJwlUCRkZNSfD2NQ+NI
/wiqd0cu04bmHZJOSwBDxB5e6SM019AOJ983cL2LevI9uv8PuBO6kCn6t92s
K28RjMY6NfiQadREYizdHwcmoikHLdkhcuRuDO01Jb1XCWe7q2yPtO5YtZBt
SnIG8ubJ0MyHKuFCI/oYX+UDiHC10F2PHX+AkvxNA9lUy/K1YbWmbytu3F4L
d62wMyar9G6O/swAvS7xJDnrdYirh1aI3nMPfkUctZWfnLIZWKzzi5QS4ShD
i5ZRQfubCkReeARYd/yKoBZfO5NGMk6ybu7GKkkzmvvfo2BNOLNthfJppUf6
pl+IpXqi1/QFH4wTuUzb3odijlJKQet8Ihjr2IuddnvF9o4tnrGVstcM6Pea
UszAvBVtmn3VTeUq6NGDMuwdEhQzbemsWoSODE8zt0/q/IfhP9/8Lj7FMFdp
zuZB86fJQEb29/57FmErXzg1KorC5mGwfWrQLER5FH4KH+P/q3quOkg4meMJ
qyAm78PYHLMsnXr9P9MRRvTeIJq2OJlWEzV+eo+uMveg/x/tdVHiW6xPW7/+
E7RZq7H1PJgKbzWvmVRYfLh4mICUEZtmahUavjzeG4IbYVyosvqZ01iaO3X2
Vu1RLrKJVBxyw8jJ1MNmqMbBgBYNsgLtdS2YAGukDTJ+91kQ0yUVmxq0Hk5n
PIXWXS6ggJMkBjGE6HcsqVeNYDIahQpry4BlNF1gTolHYe8daKDBMQhmCJfl
YhyCDB0Jd2ZXLzBSZblkeGI/lEMWeuXaABOLKlb3VuZ9nZ//Sj13FfJZ0lkh
cKWS1KQ1uPWWPSl4YbaLUZo/3GWoyy6E5EKvwzSt4xgcmCFCIaZw44uQUAqW
nu4FaiubYbDo71Qml4HxQADIINcLXAyo9JOzyl3yPuibWeA+W49yvrmfqKMo
2l9H/2B/Ey9X3lR1kOWkmCRalAm8g0KB00S8rUaISsJjXmqjNHVmc3FZwewM
tGLVCf9rcw9rH8NYisM+QxTN1Er1kwI0rsb87QCoQWlElV3B+RshJ5pwt+VC
u5jSIDZguevfYlCgFoB/qxSXka2ywpcFzMtiV/9Ngv2IEyEuALJzKxNh926k
QIYiJGcoh3O1BxMgy9D/5Nq9faHSfxmVN8VcSzQwWQhMNaHl2vq2QQa/xBgN
ruB4srAk8nv2PFAtF5QTabDWmQGyXUOr/OWartx0nDx8p8iL8MeknafXBPaO
2F6nji9J+V2a/ly3zD/47Mv197lHUeanKVaDLI81zY8VkXsKLCn9iHIrynrL
s2AydgJL5LaTtGB/4M540+8a3leOYePayaY105zzntaBdMzglhQlNBt1hA1j
qMd6SNHweCz9PU5KPKijyfLpfqROPZ436i7yeQCgwxjim3RlYieyIE3GLXqP
9tFFm4yyq66XxOD2wjBe/FAfoiM8M/5erEev5rhdNlwv25nWu4ljEDchk1sx
OG6FhkfykTdAwVUL8uUnsZNsicpdrkSn3fIsJqfVmLDYWMGKhoAee2aRaadt
0Y8/N4/e6p2j3+Ilb9ZeRwwtWIc1KXhV52JRjFn2H57laKFwjcef3wpz+Kf+
JrdHnFy1Z9gFG9MgXuzwj1Fuq1HotxBo1Pog6K1D143LUrToNOFcCjdMJlmi
9MtxBhFqXPdmrNnarWCTxml/99Z2mtig7qTh+OSkYBDw31EIGuxiKPv3nF/z
fKaX/jDLykvq88p357rlEN27bt5nnnF3dzH/11yivtPqjExBMPgcUBjtNpVY
J/WuIV+dSS0Bjd6QLtzWAkq4wWiuFbdaUliTEXx67dIIZMYiRiiu+XHrBjjz
SZ3gF5x8LrHo/ADNYWDh3F5HxskR+J9Fm/bs9W34Kz5HRjnFIKahlbeEcoyc
ARIWfPip0n3SDXZs88syZcihw1siEx8P3IKgNLD3u3KbrcN8QDmVOIDyz8FQ
Rc6fklBiEJXOuiRppO9qmuMeYen7SwJRSZwKkqwojwWd4xDvuK7j8EUYK5Go
OZpUII2ApoYnq9Ai0TKHATnnBBqRtKGS6CVBhC5IMXONu7208G+gLVYn7yma
M9NhJMMOPxp+fnGEFVk7S1Uh6E6b9jvoWMCpg7jrZbQCC1fO4P1hal9iXVeh
jr0xw3IZW2Ft4QsUJti1FhgTNcZD+irftcp0TjjCCsUvQobVBvnDr7Y+yaOv
7zaRC717R9Q+zB84Lw1Wy4uDMqSTU/idRqDALwCcBE48bMrnqXUrghNcfvFK
Fq6btSrI60vJgnrsK4vIjv7bO9Td7v8lUNwOgigLpBSFC/1gibnNUGPTvaKL
OtrA/HPPyFpWbGMo+4lLh8QbwCpEcIEDZrZZk1VSbzo/9/x6UjThRIwbKymh
p/jLkeNAc7lMsYAOiViwZGKtyVM72puVtswE7+tpnrQEimvnzbJ8EzYcMQ6w
7p6FYgjwrFI5ngELhAe5v6e7pKJO2ognGs2DGmnZ3O8zFnR4VDrHF+gb3U1q
Uc1sU6KyI/D0f5JArPviaG9ImxWYWN2WeT98aUNMOnUKEzBM/Bz7RQqcgUh4
mQrNZZCyR+ejrcU7oZUOXmCt+ieFfuWmRFs+IxdCvT4CT73Lk+xozIMZDFV5
WPrcaaNSi1+X+mkdqD27l3SXDwHYDZLsTuK094UpZnW4cm+khrco7e6Ex3dj
RV4i0/UaKf+wh6vqTBsCEWeibMN0kIl71mCA4fICVeMOiqAVso2pw6ZsZwkW
rDfI/htwgnNe8neXWoLZhUMJUZAzNAn9lRJg/DC/9NsDjAK5Q9GxMqmvnx7D
h1N0gsWEApCzrmkUXrdbub+DO2q4OTqkGorgF+Is/APLdojlDetC2IAPUH6S
txTcOEgiNjug9QiWfwur6ZnZydH/11IkPnBejYG8/a9xMCCNs24fxk8Egro1
IZyiz90wzIBH1EHuPCUokoGsLvIjlxqiaoAetjchWX6MWHz8bOENXcxyP3qX
o/a7aRX4fFDHEA9Q88Rne7juJrdL18E+Mddf5Ntebor/vZBzSIPCr2KW4ARO
CSlqWrduXR0wlCb0AZ8KwFVL7gRfr787/CeCKwkeXPRTIRO/c2DrWx55pgNu
uK7xD+n0cGgoVBvnyEHU2YVxRz6ncigNO/wo7s1mSklwKHywo2FmXaQO4qdG
4VdIQc9Rr1E6LuB555RsgKgrC3L+kSQzri/dv+tcfmGaHL6s+m5DT5Yg4V1l
Bbt/1odF5BQ7o27S2oufsW0Xl6hwtkcQf0pHOQe+jLGq2mWpZvkCZU5GykR9
CNP2F4ryvm3lbdg+BQtHdTFPG836pc6tmk5AdA79a7OK0/tn3FUwCWg+n0kV
3r0LNKrGxf+Cxsebz/HOMLM9sswquefmdNelTnrq9BwTi+6+ZWzPC7WNnI8c
xz6KyzlNgYiZtSxympoCOmorquTRbNJ+W4nrPeboXAP9Z+zoYK6rIQxzmv7l
o3cIzMkGPchQ6Fjc8DNYDo2O5QUQiOrgTsymihOBQt5WoPAvKYXZZDY9zIJc
qD5Og8h4wa+pHdRqA/cJK+QtNXedGGju4ru9Qi2GHrnEE2vOEYi8uHag45fs
j65xMJ9RHblnyQLHExsAnw8O9ONevDqDRMIgdhFREgL4nRt5NngprAItJzTW
swwt5gJ6ex2sWOXmH5EILkztCbmy4EXnz7yHPVqU2q4K+BgBb/zZ3u9HZDmQ
GYF999xEYz8htAPB/jU1mo/Uv0zaHoBhZICO4F9y6vUjkpOdI0rDmJV4QKNq
2lii49kKQ/Fb0Ts7dgLElCXYTzkDZtyDyTZXAclBlQsps1Iv96V6BVniYThH
+c8FDDmnnvN6meFELLD60ADNcVnSwAIp6tB1h3IYiwuGQzKaRrfd0cDlRIdg
JZSgVVIxeEj5x9MnxyYzT6ytMjVBQqQCn9SS5GwRK/fBKgyEJBRTXCyvvld3
NgO5W14hBoiuhqWXnrTMQQL5lbhQiQdu8ql4byqe+ud36x414dWmFaC939ON
VJhPWsiHmgCr4EwND+0MXW4fi8jX1a/3rdVKHdHezS0e/WBnXtQU9AY3es1y
8r8SAvoYH14+YK1JiAZkVJ3d5p8EHFC+acRMaSdbe1lLb7ndUYBTDG26Vh3q
MqfNOVIY4CCStT8K/Jxk2VnDtYJsgeiJ2XdWQN+I96P0kwX/7Y0UdnVLnLVq
/AtJy9b7Ifou9BRxZpipmuoqSBzf8obePK9l8rWVcuTHG9nCpA7Bk1Vy3U5d
PqNSH0ZlYVix1Efsv+wDvXfCMZUTBhvMkuC+yyfe/DMRT33TllsoVkGqAASA
w761FE1tOt1I3ppfXwXdDONI9pUaspJfNH58X9mN9fbVIlG7vdTpbAQrOrZv
40/XZOwUehnqUhDdpzBdtHb9aFQaIS1dpjq+nXYGQOh9XXaNbYytiajwbgce
5oNgF0KeXYufQiZyfvJP7N+ECp+qz3sGgXr8jzZT3HRv4H3sZnzfHDPi2i4V
7PIUdClkmb7f5bTdd3ihSWeZeh0wAdOhSYmErUh4aTUm1w6EXXzFbvmOpg1k
7SohwGB0fhhUuAqaEGE3oevKfMsmx4R64hqbWYppYe62hyAuZnf72/6s86Eu
A79u5xXGzRnWMBP7THuaz6c10x6Pqq8tnKqijuRVJmbbwpxhwae30r2hEqe/
fsWgn3iKJSVusfvljfaZr5sv8/eprHlMz6KODWOBISgqArtc65bIoVcuWttL
ka/x/9l+D7mQ2E/kzyY6+yEDnq1r8FV3xiL8tbHmYYzJnY9boNL9mrT1No0Y
QcYbDpc6opc/Q/j+jN0TZaj+I5FAJ6pEATai8ie3emAB95zIYclCLGnEWZKo
4Uym2aISVyPjm/o6TjkDqDf2lBXbTzI2vrLW/bbon0oQZ0SrHDP07TSkcI8U
eAOmH+ErnnlGB9yqT8wE5HqyNCt/5PCxdIqF9jslXTMf+u4nAn45xQVa/LXE
7Xm1Pk+Wo2LMEycXRt0O5eCSqd9MYgRHixhgab+HUyC2c5/hg+c5UoalPwCb
8I3+OwBm73/qBR6439GbjipCHv6SZ4+x3ULG1b+IhZbLqcKV6jZbAbphpLum
5Gn8zqq049vW8R4f2tvQqQ4Hxu1Zl6wdVVbHFOtnTPgmLObaNjcUAUSbDvve
VMRIMYCW9BKn6wRQSr79mc/2YbaTU+PFlo9CQG0E0r12J9wvduPRMg2CcJTH
5Hm67F9SkI6UB8GD6gyRYxrqjmixufGoB1KY1fOl6VuKFUVVk3rbg54xF0YZ
9cdZJWd2BWz3QjjC0j3tXkdQtTwTZA02Hkk7g6YcT1FSaJfBePDyexS/+wBe
Xh5eLiFw4KI/4I9m9oanCtmQ20Q0qp9H4ZYoz4z9a2Z4w6dg3t8XQSHYqoH0
a9iapmZ+O7ZgmQ0z3VM3x2USdiLaDx9VXssubwzANRWHmSauhE5tGEK9SXwn
5wZkpECi+vkAdjRfTi16uKPvlfsQ7yxZaM6+5S/RfkRtY40ms5lz3JULwKLQ
a5aTTKYRN6V+b3pT/84roM4s+eTo4EEbBPCeSjj4Oxp4CA6RkDI/nUIHow2p
XunRA0CUIr8A4d5f6BzOS9Jg0dFxK/1BlEOScgbMJl0+DiOpp3gnAQgWn/Xd
9RiYSK2H4cVoJ/M6GxgX8VNFFfg6gtA5oJXQHC8bkDnKp6+RstqAI4kzqyvi
h5a/t/N0frai3T1c2BQV/6GgZiDJ+nIqY8d7if9gUG59H8JbhpHvMeibKbAR
P+grZkWxL1X+kYKFcYqdKCEnEsfnaNIk5dZLjmwRHCxadT+irYIJowwudwCi
nPPU3VboKgC6ieKXuKLKg4Xz7Tu/V7H2gRPJKFoRY/qi9YdFqgoVCcucZeAl
TrAGPVlEWYZirAvbpnLNXphXt/zID4cvTp3lHtezLCYUcMduXpz4/qwuYhOh
ZnHXLQZ8yhtU1++1DrZ1va0DkBQYqCC550Tt/k+9Q1PVSTZEwQb0yieqclWk
u0XHDOvpw6baQ9tb7EuzYSOBVcqtn8OI+2GnIubdqvfWO00bVflvvtYAPkRu
Ut7xCpgxn9k3RM5/tMxDxxmIVYFDCijv7Zkj8igFkVPNa/ia0OqZMMmhggZk
Xp4QCoDyEdWEfaU+gE2hTnUn7BMlKAeC7pAz6flzDJQ1hwovNMXD0OxPRvBV
fXfsFmJ+2Rwk7UmSF3JN3pw48AZjAo71LXti6DJ5uNBzBAOewxeBN+APgLyJ
H47QvcuF70lLos8ReoZFnRQ/8FGukoQy0qUqcRk7wpCD9LRvTG0M9Uwqeudw
9Tm8VShVHa62MV2qFbgY/akua4p8ESzq/uHCIv1/yF8Hhsh2TyadD2nxQ1Nx
SByw1LQ4OduHXvUTuXWhgoLphST7J0jU/9B9oRX66r60Q8UXoESY0UKMRkyB
+pDWHmgZzrYx+tkej/NjpIQkdm8ryvDvyutQmoaZ+uGxlNNgfFxfFX+IVOoZ
iXQviYhe+CdQw0n+mS5umX3N8J/xWS2RCDNaPgZNZO3pkjVtOdTZdPjCnSbG
VYaSuxPC3QwKoeaEqU4OByfAW9ROCN3YXh5Wilx3pQVj777zvoFJ9eRMH+rU
nPEBYMcv4ETdF5hA4UPiJLOMHWbuMjC/r7Uzu83w2OG0opDnSL87FATUWU3I
VgYCDeKBQuVKUZxzV0zZmtDX8OWJzuqEbSAfyeiTd2dsOd++hoqwKwFlna9L
fQFn90Ds3tnom+Y2naFPp3cEei5AgIm1MOilbzWTp5+XMv/3IQzTAs+aUFlY
VVmXxxzcps5LnA6oDnpBaM0UZRcEZViI/GiaT1MnNupI6FUzid5Ulk13yJ2U
i0N6NVh8LlKXlMOeUOd5ZP6ck0gUcIP0QQt/KjUrdMQaVKx6AxnufzJQafFd
dKVEW2rp4NX0n5/gW70l3E/tTgNqWqOXYzyDJIyijHgC5qSGMrXwFQg0xtoj
qplAa9ekWfbJAKKddQhhqTmqfumWfWnAQl3h4APcNFjJvvEq/hxOK3qyTF8I
Er4aOZjOUDIOKykKUMPq5biEXb85JCGxYqO57Xq/jiWhA5DZUesZrhjjoVS4
ukDap1/wROFQIFhUxB3RYvL0I55nnHgdzXtVrxvf7p/23Jfzx1eDgHZjW2Xl
UUjHpGY95dYvxUdWT1y1a+1kCqx5uQDjOb7cjfdk4uV9Q0BQc55jV7cvySZv
4EraDPNSzU7wGpWvvINPkr1tWFePg9LgjgOBnrxGu10y2pjL2C/mcuZS276n
wim5qbq1SE4uwEMpeEq/zG4x9ATj4aybSvTrNg2Y6cXkiDtQX+/eB5IiNXso
Q+zwoeOXSnLkTs0bFegMINHZss60CxI0buaDRtKJwsSiIfyGo7u3wgz/mYE/
AdNWOkjPVKZbKxW13Q6NfShBj7e4TNa3fOsH9tc70uPMRe1QLBKMBoK4tTge
4e0GPhzMz9w/wn0xFvumnuspc7jTX1+ucQyW6eOp0b6KBMo7aTRPkYD11n1p
QbsVIxLSEkgmVEF6m+4cXXycqdsBI0sAJb5046f3IAHM2Pow27KyxorzlWCK
G8cTg2bLTYOxXKnrnJJIS69p/OlImcSQLv5sEPdIlPnZHgS3dVKcrGj+GNsg
4tpZR0nDcQGMHf5b6yf5yiOCmMNhAahfWIH6MtXlZs/Q3vOSKWupOHUgBmLs
a/nOCmQfHFEPi1aoKEy6+Zf7FPAtyWvbCXHCv2NoQs2kaKFZN1YYUDSjuoJO
plB6KYLp6Un5RV71od2WYBOr1EfQS0VqkDHQfHjjtjR8nsjDgCLfGpXfmr9g
UYTnj099NEB/Y897kmyFq06GTyeJQ1qg6+WAHgJInfytlqOMXedRL6etBSa1
u19GwrCNWAwPUk/hSktxTtz9HUexE77Yuq4PURtKYDixp23yJUB0RHydY4AJ
PBxJiS09x7P63er4M7Mz25B9iK32n+s3RH7cicNT8JNGP0ME16Mtneidg3uH
JeKhxJr4mm5kUYeVke0WBi3mPbRtAXhna69b5BW0F5ixoBMR5HUn626Tg8u6
f5wM++K1TcuzvC14UpNjRUsi05/uOJXsEJq5tIimcEDMmogHU1S3jCpab7tD
juUPchQsBQ5NMdRmdlZWgYgknGaXeCuImzeXG5AIM4WyfPg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqei1C2pJKFOC2juxKORFZxqrTicUG508IhVLSSqg80m0jddDIdkVQZu8RHyclcmSpDOgQlRw+dGY8pqc2OFNphJgQi/ZCflwMkc+xUEHdhScprKJmGk0lHsKtR1NQdiM6QG+iXeNoBSi+5vXgCSUfiZYTDEJJCs8kHDpnk46XAjXgzaxOOEcTnmQFamGrHTSIxqbHG52q8CSb2shBgdEjxZgEpWaQPEPIbIouYDtsMjddWVHIoXk1ntRmkMr9uPez4VbjHHamZep5odDgeQFdtIIkH8eIqsnXD7ttACspGyR6s75A+mihOkVDcFBLldB3yINRE76+bZ0MVPqXimrQJYJPnVCQRjAcsGjF5suAhAZNyyDnjBfCzapFSXaZCrekp0QmdmYzfGDSPtAQg6PAj6hXaG2Y0rSw6AirjtJmo2FARvxDKh705FejozpZyOshU92cPGDp3kwhnEcvFWXxOZc0iVF2nBuwYtSiAeu49rWohp1HZS8V3oOlc6/aSNhvDRJHDupFC0f1YymLLQZ0L3veL9BA+cqfQ3UVNqcpyeDMtxcwPw1kfDBQY6b6ckyjQL9g1krg6KQ08pbGrZR23MOO7GZt0E7BvM7eMkuUlrnLLMREcjaDYuywdWWellly1dr11PE9GJnEfyzjPG4aoH1Lnaly/MEPqH1lWmp8ZHwa8qo+rnYWBhGkzN2fctEjBGlgkXiQLUi8tdZNLyf/1zJpTr+P53ENqYywXrT/2rMiYobDQEHc5tsvppiWBfTUHFvpBgcE6cy7BYJ4m/eENf"
`endif