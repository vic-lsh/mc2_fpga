// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OR39BPsl9gL/YH0ygqqbwt2z3TuBklfdp7S2RS4cnkww6S/OQV7KCWYpVjeT
EHlc9z5luhYSehYnmM/8ggas8cts2Vgnmklc0bJQ2gVFu8pBIoMRn05IXC30
vrRLP8b/6WQ4I2TLQ4cVfeQX8vZ5gL+I9xfpzsh9UK6CtybayMcNcw2egsun
II1krxE/cKYmlurbxN6Iv/mFJ00iwmk9tqGOuuiDnNDbbk2HSaquCe1mdPNQ
S1UUsuM1lo8ki2J5Y3yKlbuV0hIL4TOplPJh2RKtQOuh6+hwMdYBg0OLaEXR
m1WSX1rBwRd256yJaRJrfDQXAATr7IKzmDjMx2L3FA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H0zMZGG8FyNt53tm/C3vVCmJo/OQy5/l+Yc5KjGllOymc3D5TJjItJL/4T+a
nsXhu1/WYgGbH/qCVtcVUOMdwSjl4JhbudiRAeZ+EV8kRS/fFJ06sGlhYeJq
sScDPGr2039iM1FhkFzmMSD/MEFQcz9I+r5Z7eTp9wofRt6UEtTmExmdy+/9
F9y5BTjdEFjvlVoF2kW7g4w/gcZP9XuBJWsB333GZSDvxXZsvxDWgrz4C0Z3
6PMUuTTzu40Na3quYLk2nWLYch1BgHBn/b3vbMmbuqxKP37SbbrdncoWJJ72
hwsx8nDVlTw/6rMpLJ0zm/adOqmf67Tvei77dW4erg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A0YDK520F84IKfnrkdM1mWf4+sETBgmptdYUp+L60FPQNEt3lC5MGFq2O99b
8EMxoMxXTkl6Wim76sF6PRp4l/9gZZppMeS7ZmHE3ppiwzRKAX8MtMJPaaur
aESfxeZHxMJtUA1iZELCujddfTaasZOpyaf4Ei1O0Cxjfn8fZ/UsneN2IpVY
uZHVkMETrt/JItIQJRQ5Sdp0wTYToG8x2NRqpqJbq9N0jMblNKTtZa8KO2Og
d/DuFk8jv2cWqVBS6N0UpemBnxZmEodGhuXFSVoDMShjsviGrw+fn1pgDCpf
D7acR3fp7ZBwjBFMsqyc9q1+1bTZkq1Xx2XL3K9QcQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TvWFLwaAnIrayCGkaqs0gKbd+egktMKBy+X+YTSbVYU6aio05YZ+mMMncxwJ
wrjWaSxVXz2IT7J4RCZO6CmxSOUPv+VKz8OizC0oUh6OWjBwiPPxs1gQUp4M
AaRA4hcVHhutxa4CUt5ObdsmE3zR3117dolm+AnfkA6XH40MlPdiypOJ6QNy
vHB0ysr0NZPV/+NmKF4Mvr9LlLChl8MvbxVZJA8kv7fUrdCKKOh7CVfsrznq
0MuoRGMLGG6tCqecfWKXeyCmfN0Jg0g8bygLijlk8l4atUgITwm/4wTEq7ES
JOkPDxORqe+t9DmTpgunQ0YVpLw1llS4O3T5uTfSgg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KsHa58izFfSL5SbCcGnEh1JqjAzZPvAjxNMbeJfyrqu05DXznvTaD8GgtD5I
yV2iXGEBF70S8zNkAqUvtbtkbWmVLVraaCDmDiQ3kcpom1xHA3gYhADO41dY
5gjPvjCUYxY2dgkdqoa4kWY3hMTVF94rh1ecC/dUNUolgDnd2+8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
RQ5bi5vTqHmPxexaONlDZKVeSYSDiBmmfJmLjEFK8UgtPNy+hQq10BrRObb6
FexuHl+2JEaOHbTo6MsXyJ/ZXNsPhrq31DP71VFjErvSHngergiGR9+dPko+
nQmZxIUvHXDVY+koXDnii9oRw5LWp2xT/iDByucDnOquSqDvHwmZdq4CjhCV
yfJ377uIrUlU/fnjy1P/ojUgWQLZYbOTdzXAi7+9vUGVE5XoLbEfxr0VoQ9c
aRjFpp2zsDWO5zHDm4nOu23e0fM/p8QYS02IaB+Ym8J+RC8YsXCdn73eQIcI
vBc6Gv07WWTL27TapWfrcCjJ1FNBLCXsi7yzf1VU6J5yB13lm5TDGijW1BNX
CrhZFwrDKkGrkLf4wAHNFGM+gB3GSfdWfZ5HMQHW1RyXjEgt67yHRkOE2gZs
uUeVCfY59yMagwZVQYBKOP6do5nBZh5lSdLbfUiZ9wBt/FKJ02Wi5WHbnP0/
zADTo+HoT+B4YTp4kIK1rKaKLIoSk7q+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
quoA+O8mShJObXbew7rrd+Sb7myqmFOSt3rZiD6+MS2/0eribG7DZCdQKQQt
YvX8TBfMZqk7sM5iHtX31cRP223DSEwXqsdsaAtiLfMO7tmyokSUpGX4hqWL
vlmfN9EmOwc4oeQm+RsFDOWuPaXcLFHuKKMDyL91MM9EYd+eLL8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ADwItVhlemvHzPcQimiwx7MBaKk6DJp0dxz5XswtsePGqoiCnROaB+3vG4Lx
yQiMVvK9GAPNpB4odOOiE/rOkOBHb/Y29hhLX39kz8VewwBxWxGKb/tUnpbF
krGa2+DA892pHQiD8oWiAsgA3z8bwA3jvgt6nPXp/MjY23KRZJw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7904)
`pragma protect data_block
Ta0lfsZkWqQHb6Ey/Lyj14MuwEXzACDmiP26/BG+iJS0NTBLAFavOubI/Xc9
O4/fMdU/qE083b1TBg+Z04fgJnUiDtfgQ1EV4kbw0KDMTSCL1A3wXjZ81w/T
Tjlz3ZzRIt3sxD3j3ZZPVj4C3A6QfUlZwWnYfklBvZ7pA3Z/lEMEu95M5SNm
c6Vjwvy9JkfCAs+dtRPtC1NQ5KqAfe0wdxm+AE+u5tiJ0UjAc310oUvxH5NY
ySmJYBc2sPpYriALSZesejqOgwZtW/L0Dlfn8tALg4Sfi/4a17NVtR7Q+iJ1
PerO+cLy2E1ktbgExwyait8ODKjz/tVURq7gtEe+qHSu5wNysBYho3LExFe1
zNz0HDFhoMI0SvY9qUaHzkXFVq4xlD14W+NcQWs4o/dW+X0JRtCFYJHanyxY
1+/5zGXVAr9A6azQSi6lNTXmijjV4tIRl9T5X+Iv40aNjpdFZKD6IejMY6/n
xAloFnzkDsYCkfpMkNqiqKTsnggYCoWzuDHV8Y55lf79faXQayI73ghyXxaN
WX8cRPCsWfil2w3ltwFHTyxmGKXqy2Y7cPfopAeljIA089akFhES+lx7FERF
WIcMx89ojYKyHEM7BS+7rKRr7BL12GaO6z47Mdda5J+aBwFkri50JuB5Le+2
tSLr4ntZZxzbjk5tU1MN9DVFG2Wt78ypzCek4GLC9ZMHY58NgK0Co6FX+/Dz
qrS0zrKhlfLePjE4683ds6ws0qYLgENFSCMzQctsgUuUvfvGoTVP+skloD6B
w1iFN6FgQIWICB0mOUXNCxHLvWhqmvhXuARMRLyuAaCFwxCN56HlfrupLyFX
GOqEffgssmcixnnAhIT97PEbCuFDkFU1gkVFxzeFGZp64AQkxfCmXCXiS3Ie
e/Wh8sXgX8DrrydrxfXKUSS+ubf7Fa7jEW+fqZPo8MY+PZvMX54YtCWfC6kC
C4dw2rQhBFQV8C4CRrnZ5PbLoUlHs9JonzyJi6MaAzroVhfVxs4loHiHkbWt
q7ESXEkd5XPKKnUZg0FQQRh43+HrjDT7Aj5MB6NQe6VnrYachJBh980UdzGv
qXy1wexej1wGSTJvS+gmlWI5LggWTIOnu4WnKUlxnYkN+Sghx7MzD6aOEJWb
u8O1nMgYa4SBJi6sDYMr1usMBjo2S4Xw60NdEFf/MVoqtEuxO9kj3A9JxGvK
uEJ99XgBtziM99JjnAsdXUUMX7wCEkPT3AvTw5Ka0hKWUEHfwHY32OaMCPRy
WtKt3Mg0PqnA50xKvKpuunDBTp1abPAGW+QMWl4fyWgjhoe+zMzeErAy+9GP
wMIQBDD+sQ03j1FYvLd4B9iLdPRvmBSLMgcJiZ2gAbRLyKiE5Fh1KTBTswoe
PlnwSR0QX2LsJxB2nLJhPYU9OQbM0MSt0ryoPUjkYr+1eYqXgronE2f7C96D
AqD9BtyEiiPep43R0yq458feVQEA+aIKELw9TS/oAjBipk1ks3YPnkRqmmMO
5bfQOOWl/Qq7oDGfx+Ures2sYdsoeCqkhIn4ilQ6iaptmoJ0pOm4i8mEz56a
b5n0aCST+u9Np7bKicVit4GZvkweyKPAowFRYV3YDq5fXvr5rpa94vITnRmW
ZFJqCZiz7LZO2KccYcoQy1ithBqpLXgPe3110ItRYf70oEwJO0F5jh008MIP
oezFNg3818QY7zcshfRdLuXIH9xNo0zThSEMuPELZIpEjfpzgygf3uwFVijr
b2ny8fQEeiyEAipv/PGEnX1L5WOtG0UNPF28Ye7nv2kBHyATanpQmlEc2IqN
59vUbGzvkVvys29qRbgwK1mTU2jecyi5jHrZVHy+xGSVyGi6du+ZPgsPolA1
Y+P9gZ/PkrFvxw06stXmFXYa1AG6YJ9i0V/3j48Eql06nvk3s93lt/n5eoTX
1YdWiKmgxYQTzeazAcEXF3nUIdPqDA8EQl8Fx0ONlz8GDkogVE66a5gp5AgX
z0IUmyhcSHikKfl0y68/DIkgQyWC1W1+Kd3+4588hfxyAssTiawrUEa0UQGn
ke5duWL9lNaElzXWOFEJdhidT3Vp4Met62df0HA4wkm4RRxHMH5sYoLom/km
V0KU43SzJ3gHykyAehINzopRo8ajr7Jg6cXN9jEyIFo8EMc2ZPormFzg9b0/
Fr9sx48KMfqDfL541aR8WBUtf8IOeJdZJKIhljNRsorYx1AR2TrM9C8X0Pp1
D5+tUNzOOvD3bQagn5IehZ0UGnRwG7H/Vwh+fsRHzEcuE2q00z2Z0v1E9B3V
GqDLFc7a9BPXXXxHRVkA7K8sKfOSHuz5WJb1ut+v6fRFSD+AP0RUocSimN7n
6jqnQufg1/Cu02B7tsGvwWLzW/RjtCtuDKlwK5FE9sxLzO8tABniWNnViw1m
NM6bSMsDhdjh/sX+mzhS1UBV48sYRnDM+ipTZv182HkOpj0GpTkuJ2EdeUPz
5setYd0AZ68qh7IrXrcpsgNppAu+c9O59a3TBlHtHZ2N5Gwqry1kSPxp/oZx
zDBlphVZxa/qDLckUrOgQSew0+GzneRKJKIiGUOAcyGJyPeBfoyK/KY7wwyD
/zdtglwr8ystAR1dusHQV6rw0WZQILWUj6FUbMKzBeOMnd/R7565HN1trc2s
fBba6cWQGAl/u8GgPsMalW4KZ1M7yMiTSyIVW2Xm6EX2daMvD78mSpiypNoU
+CTiP+IgdvIp5QONU7Xp6vzLRgAkQw9BAAIDneOZP9JJoCpDQP/avmEkCgJt
U+Hts/h33AnaVSOeA4WlrEKE3JP7eptoMPFj9QCkTS+b3snU9auG+q79LI5H
xCGu2orb5co6T0ABVRMs6M//fblBP9voYLZGY5v+tEOTEMZ6pQ+DGvFMxFw2
SFXikk45kSybKC0+lErBz1vczUiW4q2BMSpHow7GuNc9W6favYJJD/JRiJQw
f6Hn1pNqEt2vlSMp5sIntgenIXr8+AYJT1jDz+xcBvSBShKtVZkNR4ON+iAr
+P1X1YRc8zVz4nyP0HQhN3d6oJcjiXG9Rxh9uUurgZrf0Ze3eIAPcaVPb/cA
2YfZVsyTLdcpanxal8nyFXk7SYuqlljOpzvQTV5bOruhaySYNeK7HOYjSimn
jnfe74p3xCql59+mFSety3b8yDqCab8HFuJ3D2JuesLL1TuuYg1CAS4I6kT/
JdJuX1TMckbtmBrCw2Ziwe9cr5Bp7ytG5/GD8ydB6nsdPyoFWB6M+H1hACKP
BNNW1+2+grYJa7yfqpOIZKLEqBVf7p4no2W4GQjbgptnDdnJgN8GUZzsjVOG
588TCOOipsmw0Y96/urpuzLXWq17CwsEKKp7n9E/qHCLRmd6FzeIsA4sX7ru
FX8TgPX9CVzP3+cwthbcgUwzd6RRv2s4+Y/SzugFTqyFB0jAFcMfYNjDxn7a
cSANLWCRXf3FceTS4TD2hg2pM2Y69RvgGy9NWvL9LUe0eBHEwwejoYGnkm2E
8fXP8DUXeDLIPFW3/1hhZ6niqn09beo0nIjWgCD2B+VEZRr91b2aoleoufMi
JgtIwfsDD6AeOP94j7/pOL3t22FSB8xQugMgp1WdkTdJjNYuzsTGzl1EMvSa
Am9sOZC/o2GqNlz58kvOS9qT6/nlXxjJsXG4AR5CijywJKW9GpNAla2eAjXz
o6yQeSDjWze6iaAibyWX0uuGPUaWClJlIiCMlEVLxUAclndF4/jnR63AzfoR
RTX6ZmtML6sVoeXz6dKB8Px6c29/I2iDRdSyINs6iIF1oGEamjocKXNQUzp+
zTw+ASXbQcPL9FFwruTFd22N498HiDpWXXj4J2kS/9hWNtxOnAbTD3yL5YVc
T3dfo2bA0Hx9y2h86kCEbe2/23PHIoOYp5h0Vnu3mkNQsrRjwswycssH/Ekc
aZ+FpMCiuiB+Hl8Y2Hannmc33dN4015oVoWW0oG5xpJJi5comxmxZEFroqZ6
X9WYSmosbzCI5i5USf+9sCQWv8UI7fa2CkgnzqyfUtQxlF81ZxYhA89g13lE
WyGuTml2nnbpBEzqgaZa4P1t4eBpeZm13t+yeU1I/k50pSyQWwNJ7tF99scN
3SIQ8zCo+bCHNX5G/yYBhC3rALRVC+XdMnYV0y2+bp20MpAQQpF6jMuO5cqA
Oa+Qw6JsF6rH2u3Te4MJOoEKq3FHkWFnXHzRPzvpL/JJxGyhIHNT40YkPh/b
mIachPCPlv5rTN3mDznYHU0uJfpoepvxJoDq7A3/H0vp209tfd8YsybfojmJ
QwO4tEeV7OD494p/FA7YPrO2GlaVty0fINGcaIZlqDE1c72myXpitC4nzud3
cC5sJOVdkqbREXlb2qThg3A5jQOFvllDfcmDc7p43eM23v5X32Ubxz5EmGbu
m0SBeNB711fEgiTfclP56Eq0yJP2yP+apCsI/iVXjxQbnydb7QehvkAQXhVw
xXnMLCdLrSbMOai9nhlpP704yHHIZ7sPU5R2YVqXCdZeuN37ht0iH9r/JLx/
J9qhUvbZ2Ct7+7XF9d2EWAc2rShS2lqNA02ADCLyJuCGi5vvVDrjl+g7jIil
0A8nUF6SJaLJJHfl9Q0cs+sEAtKKL/PbRam7qfbPf6yjzFk8Itpxtu7cVfw/
KvqIOXvXUp8TJ68RXevOvZrVV8D+kUBqLPtVvZE/a3YzT5Q5UuN+dbwz50KA
nCzmSQgCF6oJKKAkvD+6s8KxeAvfY8tW29xs4TXSeeQ+V/J+T91Nvh39UgNh
lNcZHVtGK1cDJkZzJVBGfNbTwfzax+lDo0OKyq/uMZJv5fkLR5TNFqM7jgvU
pwd+W+/8uxxBV6enulLj++1pQZjgXSXxQ9QOWlmFJ1kZuVv8cbnPd2EeW0TT
a5gf8FPw9o8HaNwmSbGax6+ZcaPVbNHg8CcLESqoehvcizVfFXs9LiG9pvMJ
oJvwts4dsNtMKnxPH1kwAlHIXVTT8GYo213gfAyxoTlnZp1e13pPpvHk33dX
7d75CisehyOAdJlrwbLelGY5qwQx9FjIdFIXilpY7Asi2h9XJlN0ExGGqHAM
r/MiiE4CEzr/mK0L5h3nQfTPqkz1qw0Tl7yHxHNV7Ggg8y062cOdZlBoxZMI
jxrwYSUL4lRWwXMA+Lycqs2295Re5gta8JLDkdfPeus/lvD0BJ8G10eat5vl
XyoG8CPFJtgvSpGJ9T24cg1m/iErLIgHvChi27CcWS1wKpeZ8rTwmPHe8P9m
jDgnRdubBtonamhpkh1IdcxU7YaLVzij4aNmeOizn2medb6Ax8sS+Z8Qz9kv
MppcrzqV7+/+jo5oropE2cHrtZVuEMEMH2lqICCJZIN3VtR8dlxfV2FVUZGC
kD+QpxipfR4SesZvVQG08/cs/IuRzsXpRmKb0o50afuhXyZ54GN116Wa80lx
viU+gqVSP+U79mc4F+auDI6sM1hFbZyrx5+Lkv+pfMGIu3zKqrnYPwcdEMaz
sUL8exoemls9wC64QdCrrC3YIBXyKk92rlqwj8oRLI7uypGxEIF0FYKsndqr
+/gl19ZcgfiGuG5nznkpr5Yew+ogdjmpAYyF+bMDPAib6LohBjPFkrrP+1k9
AFBZ/khJZ9yZO+keH2++AWKHvVp0gWdRQ4ON4thMYqR9YjJPiSR/wMoQKzI6
/70smMQWEzxxwxtIieTyryu1bzIGH9kyvhKu9+t53Ut6RVB2PLS4HirOXDRI
mWRsk/zovMPVZw4sP9vk+3ogPmIijMUS8mSZdf7IUvKEgdqkalPHlpslrZuG
iqCaa+sY+6q/5wrohqSWOKwwIDMH9lxDOYRXuq62JfGhY7z1g0c+Vdz+GNlu
ht5ZsjnGJT7L7cxGpeqnTv2icHo+Qut0O72I9sBJnmJc/zlgkcz8N8IF2rCV
pk6Lq/JCLcoAFPk5lSPjb+n0qMjz8fjSCZKFCplQ5+wRpcPPg9YT5Oll7O6U
ujWcdqp7EgE1utVnB8Cudma0RnPV7rDHvATFy4nJaNpPuQTDL9k3zxVF7YBa
JIpsp7PgBxfQr97V8SyZxmHXsS3iUTNZ3S5LWyQ9EMlg0OLE+JbpfXr+rLHo
eJIA9lG2DNzL5WDGNUkpWcj9PstN4ILcsm3GwQq3lOpuw3bdGCEsoNgWBQ3p
pVnSCyg//C3mCmekAw4acRYXefj/Ao+Lir/18dA48S5bvKQ5X+D0gegaZIFp
vGIbOm+/EloG30v0w+UoZDGe/gPqg6FzWfSUFhXKLq7iiw5sHzf7l5ksRE2T
hWHP7/4DFT/PfCMDZ0fjHY7VczY0lQhVBxUe6du7J74O831vu9YpjX8saH40
nBhq0g2iCNsLeVBjHWQcBQBezF+1+l7vm18W+bgLCT34ukQCWCKEXGdwvKgh
qxSPWYvwASIszINombydxZoCJ+NoV7QBE4r4SeHXeg5cadpSwlcjjeZqGy9Q
mxZWl0B5YF06EdwxGGtVPbdqDhIVFwNGJ72/w5M7B7LdVWSVfpSHCmz7KoVs
eCgV8TVdL0CJSU7ZFcbg9vLmnnFQSj8CINE2KqOqGUOnXg1JXaUF7Smbz2jj
z0SkJz5TMOQLNs3gtEg7jkIKTn4+EAzw+xGsAk60xmDBihhk5zmybB4BgxL6
ebPXTXwf12g2UwsAWx+4nhKch9EH7olgUy9gV1g8jOrePX/hfeyi0WBKKpL6
lX9CFHj+ucAIm+A3XFnakUl1GFHg/ptX0rsvk93FdB7ONUUD+zwF7+t5Uh/Q
UyKVbeJFn8Zu/xVH5URRk8/6DHExj/grmrqmKiwGZ8AYJkZE78ARP6MXkikk
nhCPFm0WO7euU9tI+P/DadNoSCh79rESxr79zelyJhpnp875YgWetJR/JJ9y
gNSXTytSMDHE0IO9YIbCJd/XuOgBDZlIahsqC7rd8ooQMOuRVUrOwpbCkInM
l4Sq+68NOFfWoN9eMkTJNENA69WFz6YeB/jf782ZM5qRZeirKrhss5VyEb8j
y3viH31zYIxLMkLYlX3sFUrjn7KNS65A6ToBx+wdnz0wheR+s3Hczp5BJCCj
C0LWsZNWlh0xsiy1tbNxUPUd7fMKa1gdg4rBNDRHS8Ob8bsFu5jhGGjSxy06
VyTgOJVviDnOfQIpQOktHYyoErja7r4/ikZQZYudiTaR8o4Vy8rrXXYDSh61
bmnPc5iI87UfjPFDAJJn7+ptN7WA0JMIfBKebblpBczA70S8tm4fp9D7jQE2
yRD9e96oNju5J5jx9TVOTa0nyVtdaRUl66FlJVaA1hY28jSN9VPN7D0FWjIs
uqRa/qqXd+wuk9t6lo2Bew2WIl+6oqC0Jl0HA8Etv5QCNH9sV+gr4vDkrUlX
Ih2w1a+U5nwHcSQ5+lIucdQvAJ6ebOm+whhF2dCCR/iWZpMz2TQaK23JgS0B
8kc4apzcoNdCeCtmjuxPuaKPYIa4RXhOVrKMFqyxUFRHEp06vdPd4Sp5J8QJ
iZXyLXYnrPtq1Joqby48Vf4D5a4YAD/ukKaEFzvPMeUwqlveZlY5ruaaSmSv
IQtfGNMHYcxUBSFhl0/bDsdmvj9+DlVdElIX9PMZVtzGohTh1jovYxhwlSXx
j3eRZkx5Dh0MAIF6UDb+TrGrggct2AjyHixwXG8gepb7PNprvQMYu9vhWI7P
cchNUskx5TsrVVTKsgWibQBGLe4VN4MHxXfi9ezmq/CHJO2BRj4CPOGEEdAv
9vslLIMWSWlHztaNqlRnlN3SatC0JB2F4/btKMQPi6Y9f6aynEuLsp0cP2LA
gF0F5uaI6G40tp6HChDmggRh6eq8ZLkvWO9Tx3S6/jo54FLVcyEVLMvwqW+m
/LLDb+M2Fk5jfBLJ4ZaWzZH2kRc5M/ACCXjSWGkUka89myZZMffe9J/abjkc
oKqFhx+xYNIR9xLnN02SQaDDsF62VVmoe6dae6Aa1G6ocwmkElcx4cONhJLE
PMLiem01oT1eId14Pcdbc80ewqKkkg/8J68ASZbQyw9GHISrbxal5Pf97lDX
eJPdR6lwXbzH4S++3DPnkLlUu704LmVSMf0z44rDSCBxYz4By1EfdAC6Etz8
78hfc70JxDTaRI/CWF5D+YEWp91E/5caPBaPHfUrs5I4+X3ADFwfCNg49ZZV
2z5LWnyBtj0ly8obRWcWzAKGvp3gC0krSC352TNivP8UIu0p6vUCjZMuIHFD
jjVb5rCtZBlwQ9qeooewo26rbKpVMvD0EmVfL3D3OM/jKp2euYsIzyCPUceF
g8ABqXqhP68NRdWEZu27Ld6184fCP2b/oVLo6MjxEpQotCUeCAIIarIuDBKO
OAmjopmEJMqJooAug50PE4M5RIPV1DCDeYcIwHxGqpCw+bMg4+LIDbB7MttF
S+llduZoTPn84yQcsPPxek4y0mEzKELhOOtlu8DamJmegokYIWnJbMQzD1jg
PoENStxck+3ATPleN6k8dnw5SRSesLtYC/VstpZdGH8HPcvJH7fOc+RJSyDF
j3U387+WPjuj8XaU0qtjOnPHR1mg13JScXVrpsDTmgA1A3AZBvTniq60mDXK
9AKsmIvYPSsJpnFfsnlrADqJYKzEVnbOMbnsPfHUMM4ygc4iecQacd7qtT5V
jBAkl2NvHVi2dPD8VpjrPnwrpMchgmqyxOKX8svemRk0fWyj5R1hW2Tl+YGZ
Ya+VNma/3NyI3eOPO64YFcCEGIKPm2QBVblK0J5eQWWMOfRsMIriCO6Od5Is
u282WF+MZxI6HcmNnKQS8QzWnTZ91CBpMo82N7Q1PwBC+24Po827BCD7sr9m
fqVoXoNzA+Z2fuDudYuU3jNXsveML35RtAvh/7ytErRadOw+aCk0+fBteGD+
wZAmOF3T0yYK4EpNShUQWgTX9iCm0oaAHlLOCRwsUT1lwGgCUVgcWscQw211
RCqpvkbkMKujZ2kUZqo1Wy/MiLMAN//TxggDRQvOJCY2CVr/RYq/WFPjaOzZ
HHGiJVpaE5F83zyx4YkhaoBBlZ/8hDroSfYHpkO0EKXT0ERGXM+q94ockc5u
07u0ZazjjSimUR4886LOaun/VC+kCOh6k76O6H5O47ibCZOJiiYmDcWaAhxs
MlD2WVRIu7plHvGoZROsqJiV3PWIbaHRUh9USgtiLBFGUnA4M2CxhP4r6hqE
2VShmRCz46mg7bacbJIto777dLmD7fJ/HQAGke1faAh1cwnky7TKtbKJv5t0
71ufT7knE8TubMQzk3AYandNoS/YuG+eA5AZFJn9iVPgpbBpMLcToWNGy33l
mVjz2WJgp8tGQYDVamN3F6b6+bDTTTfpmOUGqPFQTyXlMKeu7O31WheRcKnJ
ZGwKmk7CR0HJg7Zbc9jdw/xIB9jaL3iKaQu0DhhIlMeV3Rh1sxkqbZGz8D8z
9OfevELTIrqcvtiIZFT8RyGQYfFZiq9iNfJlElUTnlxvfW6P/RO5JdTFwBS5
0xpzZKu/pA0cIrcL8UCY2ZfVHF+o4cSyR5fZ3PuZr1rc35PEcJlSpbocPahN
eqvFd8HdyNDZpS3Yk9HRRvwuPwsNDni1JfwTh7yekdkv58TQw418GL/BGyeG
Ifrhu9xxzUDoHP+H1DusXSeDQzLODWVpjIlF8Ey9A7IMEi4EsNcQ8UhQbvB6
jWM0oo9lXl9Q/mpuL+3aj+xR6piopirLSnxFMY6muyMqh/AZT10y+A4BAYpr
lzH+jsevRuR6dZUwqTP7OPqoflB5YUfhhCcfv6wGXlsSxiqKi6bBT/J87i9T
EQi3zPuUersGlehAyG6fTir5qfNXk/QYK8rNW3Jo7z7xZcDkEnVJf6YxTnpG
ChVVnb+S8Kgf5OpRVbk6jemrUMTLFhXmq0IFYH2EMrTNAWpL7VCKRulWpTdk
lxHIhGXRdley9K1zxIgy4o0CWJB0VzVoYfZvYYLpJE+0H19+/hJCXTA40Zc+
/CGs3KfcZQQqYiIO3XI30Kp2PDWYapJG3dFAq2N2JRe1PpLDfuq8kEcQYRmO
D0MwTwnFSBxMSe5fElZ48NROgUaZMbMgDus+7FQBSotX1IJ+iPQqtZR3PhzJ
tKvDCBOr6AbY07vb86YJFHM+zgIKw9eVRKdEPfmudLC1uT4MVnAVlcHUajrW
mfTeiLu0Sf928r0kaefP9rmtbNv7ORKsqW58zq3u+6AbRCDSup1G/rKWKMXp
oj05lGiplvN4p1XaHfvxz6l6brB95gFpxVlfT3cWi+fGBKx57wWz+qMImyHp
GGbnX6Vm0ZpikEBAmqipRgVrDHyLNm+jsxCCCUNpga8urxjJPoafZYGlO+wX
gYdsiqyIGhvv1Or54oZTQEl8fqBkad+bk6trEc85ae66wdE7eJG0iRcnvxBr
+vMzTcwQlZUOOCcc5ErYo/uY/agQ6KhXyLcXw9H8YZUwqCJG6DCxvXmR/fIn
DZs9Kqxk1abamZgnk9SrjMUWBhp7BVaZt28r1YGVAJvLxPt2d5Wdcwt9h+0Y
rNKk2vc1uI5J9uGjIk2deFY3uCYTj52BnuTVup7G4u+QowVLBzVCROt9wF8z
hkvTytJMtQI8I6sG1R75uyZJ/SRumZev5jdxy8E=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EqNWBN1P9ige126WdGK2j1sGV4sho/wcbDFAWZuHUEPdvBmAINVUKDCjSnz9sBKZhUf1Tdi2K9ZD75GbsBdY0uA9NX9KjE0hkOyOrDyz0nuwTug+1kBHwit0r3OITOpgWn8idfpnHM3FaiiAvHeJvIXiLnMSFdEIf2+zGDwdH2gFj6I3qTv3P0kN+v9EbSew2X7i5HrRx5hrD+utDzsvskdUZDklS73Fhp+WMJVSscL5NEQiBgquPQ5irddqEcnAlUM/BsOh8XJUgooR5jq0m8VTuoXqPetU7yG/OlWfDFrtRMgpuywRRvtCGaby23bHuZ9FRn5ngUP5rVwCkh/T8CQJPRmAcQ8N+00WQzafg+UCX59dLIs9VXJmpmQSc0zpZsglzCVgbccRO3qRhgIcPlhEdhwmJe4+GSCH9sQkvcye9XEF6LwfHFQefct4uJGIDxXYd5uzMbL7J70Qqu6HcapjVZP+Az5eO7V54QZNxymavnAZk14GrFQJZODH18vo7UmTXJ2PYpbe3k9020tGEYXBYc+eLQOH1wiERsNL3vzxLO64q7JUgbsOqMslU4oxFsIPcR+lsf7UmoG5j501GHpJqh0/z4mUzqOvHbEnhea4skkJdsOWk6cLpOeRsTvqQShHxQwF4vVuFLkHCL9YGpkSBbgFs/UJ/HDPQFhuVu7f8YWo5gUzJlvp4OG3wuUAmM+6X6AR2yfJcLGhaZGPYZlxB2Hi61DwlufUdJl3I0jS/mDvsWxxeY5mALVDONn2dMfjjDp2LG+9BLTAu92SSf6"
`endif