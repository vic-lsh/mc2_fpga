// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HSKCKf1yPNY2zGCJjieTGTWm2by+8Ib56KyIO+2D7cfdoKNikdtPiIcW+5Me
FkA5CKa9SXeNBTZwA/O0CwyhMBceGqWoYaTO2MLDHaKblki2Uzhs4t4q3Edd
QuC1c2gUplDYIxM+GH1ToveNONmgyms4CdAvVNteS7pJv2+1MpCcTNg5/WZt
C2gqY52tdF/u7ijgzV9YW+sQUHWjL0t1fLMHAf0bQKbvcRLMTWoE+AR4vrtW
XQervxMi7EG7jFFwFvnCrn3JfrWJlZJcWkEkWXxjnHyrvpuGwx0VrF3E8sAH
Z0v1Ghlgn1D+5/vm7W9iIME9+eEiqnkvgfJAeKj/2Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Zl0XO5lodNFwcXWS1J+IFjPE7aHDfKm+TbESifcgI9FJfznkN4czFD8upX4m
d25DHIGln6eYVnNNQNMpqD+iXds8vbMhWV1ekZUKyM+ZQK0XYEqnSDwZH73z
Mp38K9mYDXuMIjj51C6Yu4MTcCQJV7Vm8nF6EzEKjHvUt6phxWzZ4B8sIM/e
UGmYQyBS+82Qq4rT01X5PZGskmiNrivvcvF+BGUjKXk8fdve3bkZxOzFKVBN
a8beDSkZ2jvjgDVCtOpYnsEK1ig9yeZmjZHdb2uLzjlV+qNWYukw5NvBwGbc
xwiUfWkbdiVoY1qaxqQHGqng7uyGpDYvdp1snlh8HQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tfYh2U9Wz0HNppLkkmsC0tUbJ8c7SRNEDlxczhemx/RZ/xEOaMJerVYHeL3h
iVkRKoDifwZqP4LJgM/VFfQhB6RMEZ1TrxHmaRF+ICdK/TcbyDk1Gr7i93N5
6rEGDtJFbR7DXgbcp7Pk8CjTxiqf4Jt36bx7ToPpnLiLD3MOIo8WvWSEou+H
NKbWTookamad2vziS2Vkx1xbqV+1Ue70Bfftl/WJkmLNrL5h71CAbtB1F+i/
v9qZlq978G79Fbna17G6NT4U8YwGQ2fGUUGDerKa0vjntAHwiRYcC35mNhBL
pWHh4oeqfprTrhLVoVnk+5qjWofbGrOs9aH7Rx436g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pDpiSBJ+LUCN/7ziEQTpGEYPBHZ9lVU3r+uhFGcWIAeHzKhHYJdNIpXJLo3O
yHjlPq2mEExl366XXYlmk055d1jVKhQkIqMR5448SjSA+2cEOZPilRgk5a0Y
wXuq6pyJQ6BcWNr4aBxwN9Yk/R1awvV56UWYvgif4Bl70g1BEnFRoxQle6Wz
raySPdTAone0YvgoJXap5eUVQFaYwC3DINciUfqDKjBFlg4Jp28hG9cC7xNM
ezQWzTbNcyqN6/O8Zjtgp32C8hzK2QFZrky31EHn0gAIEbkBjPYCk1Ohr7DA
obnwwCtxHXwJxX4qwts4qB5PfzrFcZ+agd+r39xzjQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OhghFEu27Ciqn5tAOeZHUDIEJ0iSJnWxJCogsSJoTQJISjgZKrWLrYtIjkFz
b0KqjbS+fuF2tKV7ddSWc0/Mki6ZQ5ZeUTekwlE0OuRrn4N9TuUWl7+G+xYT
XFAQzxI9T0RzUrWsGpjH9OrGRW1wGmrskAVhabp30ZsP7yMYwao=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
M4WjCSuZgfl6PDykndV4XtBoZoYN5kxs1/rWonC6g6AgAPJr6OnlRmXFEpOp
yvx11ez+PsHOEXWqGzYAB1U2MVS9bLsfX0VIIt3C8r2Dg8NBHulKx4p+JvlC
WxHDeFDLBQY/CD7KzOxdLCBl7cdMRMJAFy2p7h50/L8AeUGf0yHO6htuc6Fy
iHzDuusNAVwp48v1Uo8OiMJDrcNfSDNh08WlOPKMH8DD0grWXEQHmj5Ylxxf
nJoM1C0oKaSGSrKeshbH2L10wBjxdos+AjQc+vz4gynJ1hagxpHOK/vS2qR9
mIQYHdLXQEw5BeItq2eFvzBwOG8AV/rTE3Z7+dCKyUrh+FsyRAetf8qTD9qV
8r6FKeIsAjdWDez1M+Eleyvi5LBjx2+uQq28DszC1NvUhGfsLuUHjaYmH9Lz
wvNlwZW4tahte/b8MGkRYHwmXheArYXuQAIhC5CVbJLViTZzYZHdnhVQYwmO
zlXZcg+2kzwJ2i+tkXrtcXwYKTIb2BK3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
c/R2hWd96ySbzeWh0+1p7UzU0phM9ntXG/LjTyI+EmBkVUEp0goIPeaGShKv
itNS2wue4UxcjrTpXxSoASSFkf31MaMrUJVUxaQW+qTQBuIOQo5nyJQWpGuG
R5gaExR1tbT27dez1X3+fW0Vm3CQGI5UhSK2cx0G2ZSK8z1z8iE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KvK8DGzM2tlZY7+1Dlbc3mgDOv6ZbHg40jRa8dzJgeFvBhVaR9PKZVxPTcPk
Srzj5W0276XkibTmQ2el5PJjsLL8kHFhceEMUZiBKKOQ062f0/B5+E13t+cB
7kO1NpGmrMDX0qqrNO+aI/GFVo+dQocK/MGFK1ERDOgLI2FWDtI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1360)
`pragma protect data_block
NCKj9cTauDxYyJdNln8Ea3NUqIszhOsq3/AVN5qTt2U4amZSIrC/GxUf2Dny
u1jLSvAwPSUdG4zBVuwPcT+DnJkMIW8ZNAYSjjpJuww6QsBEoIWWH0usECmu
/osAKbSg+9WElwMC8g0ZU/Bx4b3s2XXH5TLPs1DV8DIfrqa0CR1kNDwZw0/X
DLn8cEzVD90YLfBi+E6l0PrT5/keim4hUlJNz4zY5z4V70FmDzQ9NocM0bWl
IqPj9l+H6Tldt045VBC2te8Cu2nag4ZrpO3V6bahohE3dIhDX1ZT7KQpLycS
0rFVyWIhpqLAGMxk/hiAi+tL5tovjC+2uZ+kZdEgqMs6/op1EuzyxF/tJJGb
ZNUmynwbppDw/5iPC2cknGnuZgnAYzGS/EEPvCZTpP8AX0ghrdp10gJ+UXDr
64NCVEWAkMLasilXBIoBphFSgL7rBqIQachZEiGFfw4Ly6OmG9YvuFbt6WH2
kgFSvjsCA3n+QnE0a2X7RNHk+hiW2RbZvyfWNX2KDI0Kr6PrLshV4rwAkFMG
yWhplBR2g5AQ4F9WhK6MB506/1nFgE2ENcrKtrZEKNt9WRejV6sc6AmqQf9l
sD0d4foS0NjWaR4fc6OttMDk1MFJt2pgB8c8KEg4KbF3o9R1SIymvv5MDUtW
jXUdfDPuobpCgkFZZYnSEyw5Z5OXTtcEji+AoD/Xqg8/lXjh6KFE5FJXF9DO
MkbgTdg78oponWIPvlHQMVKVTK0ADfRzATFTg+o2C7MF/qYy9NRdW815/bsS
t/BKL3n98Jtoudxpuk8ju0+xpQMe8wKAlru2eQ+/KxqgSPd67MSxAIPPUSXy
ZQ4EsH7IRtJTF9rKQRlBYRkYmuW48ToIz8NlyotP2Xxdy31LmMnxuwSLyeGi
hMECWKErXobMv/S0GYGjs2jWmxAyzUkk1+0k/WEhyvOpDS+oL5NC53OwDth7
YMrArXJSPFWob6QRuRlT5O9hy8NkXoYjqfZrQ253Ve6NS6LpeGeqG+J21HfW
T5qYaWnqYU8rGhHnQ900cETMbW08bDcALCJb/V3+F0SiZE4p2Nbqhow5ZimZ
3pqoh/7FXllp+L9loDMb5io9SeJS0fCAIpZknfp6z0gYPjzSpI4jDKoQTmle
aBwrgwW4xuJjSL275oIUf5Zj3QqXd/d4Y/lQSmirHS6Ujn6nljtIoka7WWC4
4WjYLZRvB2VNhLSchmlh1Ld9JdenuZmJNkVFdc5n1kFSspDVSdUKgZ33o1Ld
dWTM3WqSqI1D8f5xWW22VhJJv9hSfmY/pH1PViExhJRkBRLQ2rTtPFE7offj
CPVTzro+pSSDdI6DiWP86FCoEKO7p2WZjCnslXZ86suAJjM6Gp3+77YLIzig
5+QBVD0U53WjtTuaQayfWvIZHwua+p9PLq0DfbGk3Xt4HgHcVln233ok2fZa
QZOIQ+nkwCOyVhfk56edoSZbGUvufisu6HKbDkyDDMNFjAj4RNXTdeU/E4aW
kwwBWoBviuIAZo5aJW0co6Ry2/l85MTTdAjzQHOmplSPJuVKxuXuZRtaJsUe
MPLuwULqCW7lmaXJOldpkFo4al8Tcp1mjah8HJa+79+v4mOxL5y4YipPQtQW
7JWWmFqI38q1KAHeD9zBsVyRElofEFXUPA/n+cCw66ZSsVbhShArL95G3wWk
AmNUVqppTB6TC1YI9I5OoqPwJgfjAU05VGHtTsmHcDCnjRHjVFGfLMHDd/RU
sSlc6WXf8sVN6650OOWaBTFVao6Gd4/KJKZcnbrrFyOoer9NXwJt0hryu+1b
blRIugoydyWydQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoyGW0RRq+FWqEMuXoBCTPyXfz8CFut4+aOvD/PnXzn2YAE94nBrJD6HpNModEUii57xoO+i+serV/Ccar7slm409qg4B6kgmBZBs07Rj9g9cH9SCFPS4QOMopAoE69NVcX9p8XmEGfB2WesAqqES2golnUcUG7VYdHC6noREuJwZRq/+38F8uwPBN4Mcd9Yur3YkBXF8hC0rgqPdvykEmrQ2plqbr4GEpO295hmJq1pld+XlrNtJ/gbQUAfkeKjBInbdjXOUb26qMbqTl2FbiwOMy9AgVxJolD1BsabpeTv4uXG28qKk9rmAdr+CFdl5KPjyFMh61kLbAz2WvXMX6keb3+eigq95SN1s7K9yNPxjSsCeBWNmYiiUFniHJFe3lKQTcHtfYfsX6LNef8CC5+NcP2w600Pt7EdjkMvK2ra6p/49tM0Dyj3qrDUFdDlD6kcphOgx/7qZ+iknZAzq6bEN6By6+1ceVpChp62lQWGZHYpgwazLsPNjVZRSYjF1JYZMS6rV7Y9/Wbm98T/FPifILmQCXXYtp1tM3rRx9RSF53ymTr3I3EW3FS1wXW1FsP3TW5OCArl2i4HaTt35KO6VQMoZ014lqY2BMjoRyUi4EKzHnU75mvrGsdRUr35Yt8JFdDQpCHmdkid18h9kSBJdfcgmqqszOiY/cdvoSlSUnIzxK+Y+GpzMq6JsokGU4N67s2xhRXnDEtI3/kX2ge+cVvCtdifwGJTj5JKJ3zR1dtHZnzq31J6v0YmXD4wjnIlIHgzOffgk42deAemOVkl"
`endif