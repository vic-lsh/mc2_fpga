// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
q0rXrWBlOXsvRPgrNWnvmycFIP83bGP1x+5YWojFfmqRIgrivUd0oeZN/STw
H8pyXeNtOET+YP2x8nFumXl9TJ24rBodN7QB3fkyNlFsqoh6g/IxpW+/4zBh
oc9kazlXxNnPWzaowieny1KJTU0Llb+zMCo0Ad4Bzh0VIoFSmeBmTmL56aeJ
zNzQtLSomZLgcbwrPHKCxa7wM4q+neZ1GDblKetuFsvjHjHHhpjM1VFX9ZK9
rNmSwL+7jSybSE7D96r21k9gDv6YAR3mCnO+Ag7dRwtbiAoQdQrXo+u3JuTm
ICh0UnXJHCRJ0goXTpJT2FMrP6bUk/bdibOxgqXiUQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WSkUcT69vQWGYjztR7L6BzWHudx9LMJcOEKkGLl9VGqM5oY72+b8AzmOWzxQ
ZE7S2vRUeBXJcVNcsFI2v6g/wdXdFR8U+qFJ/UcUSr1zzcBnjKA60TgKiuFq
dYTcgAXmyOEkC6TpJeUstHNQWmwPUzDg7wCObgzK/2DsVwBTglo9nDs8wNfc
14cGve3wZjm+lld3EUIYNLBNsVnR768J5irBdCrmXP8Jzzjxf+1E8yqRwc5p
933BeT9s9Wt7BxY+MdkDY7flKCHkfgQRSUy7OhJYDMWCxnHV8/2//wpC+j3k
E1qAn7Ut0yAT3357PKv/JJrkm+Hst3Is/EP8ZB2ByQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jGYpoFvaRP83Zl9zxxb6YorfWTcuEedhKZmeP5Bfi478i/Bj2iehG0E4V7ih
f0A0Ob+IwqG4h9bsO1xQaRW0BGUEa+kumhfUgkVfI0EOFj6Y0A+5wCvOwrYR
iHfJNKinoKomaG9H4AC+vLB2jFPN6zOYS6CaMNnFRWEKmdLWHAsu3nfdrwxp
vExY4SqdenlYSwRrPz/7szaiQmwbjQP1UXYOmf68oHvjiNxLABLOSMMsW7y1
+7/XPq4+FpH0EBNagwfu/afmYzvLfvV2CCqeP2lUODLsKOPXF/pEtTIn/rAg
6aKIUqUlh5dJyYIZl1AiLmYEzH+vHiP8pJFF/yQ8vg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LOHHxDuOwree3dBMXYhx86iu7E+s3MdtiqX/HOzEwNbGf/UDtxc1xPhPI1vr
ooLPQ9bpPxY5BSbWYfqScaRjOZU7BayEfoxUJpQLhjDIL0uhZHW+gRu0xXf7
+Nt6DmhM9WLB2yRatyTsezq3zP70CVUOc5P/wh/HOUTuDr3udBGV+0cNPYeu
CrAxVR9oMswcxO8+k8G2hMXZ8mRHW05pEiVzd8ng/YhMrcxvFpi3kwfWE0ik
u5jlOydBeuvjra9a8KMoDp1zhCzdkytkMCPdr7LTKJNxj/M7tAcc/Y4hmcnQ
CtbBxdSKlxrwkj0wXpMnDa8oxqYnL1/UUKfXdfP1AA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jxGd869INwYCxwlvG2abvWKe578xQs01x836bRapRqoTupBryAz0ss+18JHy
mVPNa8F8PKaj4UWI8BpIUGDlkUj0+O0gp95VQjwzkTxMipKWUigtejtBAxW7
H7I9iTaz6BUG6rTbKFCm4y11gM9YlGwmYb5yKy7cDa3Kw6FSM0Q=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
IjDN/4OtM/vC3fiSoyEVNk3YiTQ6POrE+Aswv032s+r7F1BVCjVT3okS+y4A
up+LZsNrFfPXoI4AFATCB3pt3rYVIzTbrYgV8rtJC1B0s0eIDfGSpcmtLL2+
1TFoROugqegdI/tvS5tJRGDBM1QYkyU1DUJrTpIfyL2KFSpEpgrnpX0WpU9i
aO4z7h4T1AlgcGAxSNcZ0+rbky/1Dh4CZ1KshzL8VV5O4J2Bax+KWvAvmlhJ
hzdh87fXFagrd0S8gVE1u0TzUAbNAnKKfVg3EwzfEUVV8LHFChva1tInD1Z9
JdcBXfXG6l8E9kV2v6qjIWwiZtYOwA3Y+Znoo5FV3zrF5RKzM07LH1TBDEtO
1ig0nfCguWucABCve7l354IQtBaRtcRzO3BKAt/fdGQPNo2ZcCvbcK0f6k/p
qS/9HvPMsCKnF/8Li34CsXBwxC7uB1wsM3rKUtebi+h17ToYQybsZqcWH4Ox
sYQefs51h9Ovbnu1xAKMrvIBXoJDsvno


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jxePdKu879sI/bs5ne784lgpiNxKDCHcO2lI8TWzSkt8czh0U9kK6wpBjUty
ahee+5zusUEEh0kAZ1PBxpqA3H66YaleOHCfeg48dVrNi0nW4VWTp99Bk5av
E0Y7B1n5EeKRINlKbbmVpugw8RDF0iWsV6Ra1epwKZKn706Z6pM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VPDkg31rKWHd69Q21DlwrD59ypEgnWQGbCi9v0wvcBn+z5RnxWnCTcC3nLw8
JV+Kksn8XPd/bZjurf5dltdzt4fW/9dOar2VTXcWO/T/BxO3jItqa3eydJbM
ehjZnIqQMbsLKYxcenkD9Y7nW2sUzyiMoZC0eFhLPQr8BnJ7wFE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1280)
`pragma protect data_block
pXhCeQ1vl0l++pJwIhpDAdW59ILDd+WGNgRUN3WPRYk3WQriMxhO5UNJlrty
CNVYGy0is2vIu9QHtm2JqwF1avwTrlnfU+jI9kxevcl4jko0ZE87JpZZmEVn
lnDPI7dbry4572QNnEdXKy1x9Jld3a6cFPFLlRsGLCjKNeUXzJFgDwDreNuG
DR3c3utDuGMpM4kt2vruzZkobF/iJGzNmlc4ziwXOe3TqNEtvJnLD4yHGpPA
iZ78iTCA5khUeVzbpLI8L73O6xW/CcsRwBpU8Hea/RR2LYTDrqmWjmkQ/XCR
RLQY8pOdZ1xISyF444U2jEZHVNDe0+9AEgBgnp7Sa0h/uEgtABITSiZjLGqm
/NHshkNR/Z4h3otzwDyBE/yFtFyqOZq8o2dEUNx0AD778jTbjI5hCa6mPeLn
FUxn3uW9YlD7swecmxopG5Ag0SEHnq7VDbjr0LvzSwV2YHM+vfseQMR/zIzL
BWfmnrsK5LWTUxDqHpLY+C5TCR59R6hXGFaxgCwJq+q/iuCMakMHmTCDOW6q
g6i68oP6zBy039+vG/qQbfSK41RE7A5kVTcs8CdflGQDJRTc0BwH9xc/8Wix
8WpIATb2BpaSjnjmrMHr55SiahZetTi4EzFTjaCMZxje8UUAl42/uozB0ta/
Vo7THyy0ReASmsL2buzMb7i4DQCeqCL6UrxNID+22l3bnRm7V+AGSJzABe/X
LnsE3fhXarvkSAf7QkuFsVaLjDbbnzRu/YyQrw97kQwV8UyJ3cEMn8051/OC
VTZVAuLaCJGKUKU9jqIvhsMNb5MXeQXITUAlX+DFfeNL6mCYE1QGk40qAjb8
d0zzFv/3tFXML97aWJH79Nu+3WhRwtoUrfcwgvHjnPa2t0rVUfhPuU0aekKY
lLEe++XjQNc2Xy9heUfkETA+LNuHHM5uclaSfWiAJCYYXbp0i+PRfAW4/83/
yWzDqZGder3dcUy2F/DpKxMLs1SPtahtYjgYqqIrnuE4fUcWjumsvMWxlAIM
jcaom+4sdY2J2lai4MxyxljZjRTyf4su2YNs2hHgYrPWRJW20hdkWwr/B57F
SEzIkdAK+FsgqIGg16u09OAl24X3NxCwCBajtmxhZ+MbngKKVEdKEKF5pCPp
sgvqjdhBUMNa6KxteivpyKXd785zgBILHbKZEgSYTlTBD2yuj7CoQKVJg7+M
Jb2ijJ8VKrw8lRbwX75UC/FB6qc4yBQDG3R2vIF0ZtN0Wz3YlhMhkSTeSEJv
2poTizjLAK4JXGmziTOIUe4EnyTRw11u/s5ad1GBsgJoAfeJtCaj8Og6oTeq
85D+eemz8Ov+SxVc0DmAgZSp5HFeXs0LYks+zQtmuUkRKS2mdzh/lqZfsVh8
wc23lcW+cnyYFpLgkYPFSsFDSDJ4RQDRd1r4Xl5M8idxhhJjIAzUGgOfISSz
nEHC8WHYHkrOEhsPEiI9EJ8Q8S6TJu57pFRarNyh7z1jryAeyvyXLlDpRb4K
louQCK9pHHC6QZHebRGAIPxl0Dk6TIGXCJTaFfmS5Zt4jh3hct39BIaiUWQe
cFicrawpKOagv8RrLdYvjOvdEmj36LZsAzdyVKDg/vOmYFhFh0csQdLtyh7z
GGrwvqsgBB4gIz1Kul1D86zQs9us0go2ijMdbTEz32ehg9kuqjYA711yrLEg
XvVyeX2GpqK/ZRZ4hYJAfG539QE=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqc2MAMAR6exhNo6Z74OkvXcYjr/qKAcbMKIhPYL7HdoJIy2m44Qc4U729Zss465I63HAW1JlOBGt8/0qBj86V3MJ/dfTiernyrZuLfUyp71E79G/g2eD9aW6Kz1rfPdyw973kGztAAHZlMmls+76HxtkSa5pZlgL2R1C+54V+MkV4tU2CWEkJmPSFhqZjtWO8PAxS8jojNEqa7D9kG4DY441SdKl3P/M3xJgtuMXGaPO2Y3v4jPQ+6v5jSOjkNryEVzrkdl+p62J8IOlMRjGG2ZCwFIus2y//kiDhuthclZcKDxByuFSh0XBc9jFLRq/4k5fddUTokMfFi76Io0biLtb6Ese04NjKwIjVkJ+Cp/Buym3kk6Dbis5hUdeg9LAj6T8lPJp6XR6VoJg3Qrpe7vN/zn1cjxKloM6l3CxPk2GRETn5LLzxFmZqh24KoVYmTtfZ0eMCb4QaJamU0+3lHq/PzjgfKKh1bQAuIFY6AY6vK4/VMpvWLgkTx/4VrmgfqU0naQXnQ+I1EdKZdOqhHJrJ7hYec29Ldf7e4hZfZKfULED2QpjtTW3EEUt6zwXUOQ2hCKp89pofrp3WJiFee8rl8TSJKcL1iyJfbUTQBEm6yF7oUtFe6ZVVjqGmgjTO1CS+84QMvzZ2lJbAhjx1gwYC9cn2++0h+IpjGUjyJ4g7BERWcEsUAfMDqCmTg8f6yhUdzbtu1ubGS5JJIiFyzSC2zCd9qTAKCa/+Hu71H1CgDvYYtWYjYZW7HPwRvmRLd0wtFTBvNBqRuvrLm53oL7"
`endif