// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XnmcXXgYqSkFIeKya+w1wReu56OBafn72Um/b6N/+ETs2clGVnOGIjDdi6dB
7cDzHo5Eq0rr36qEOQQAPvPfJrvcYQLiqOvT10cTXf87+oXVC56g3lrWATJb
gPvlpRBRqHREgGW/lY5HoyaMsiXymX93vxmLL5m3p809rkP8t3YSRzF3IK14
QVDbnRWmtylHKAOhwtuff/zWcgiwV0a98Gox/a0/8+w3o98N7y9btgWJh2bP
aRcBvjQt+G3lgwCQVM0nbbTSz/9aQr3dlxO2GhdvGtBBtzKnxv1UbPVPpXf2
AMqoS0/b+AU3J3mF+SL+rNNLdGgm0QsoEdvZoLcK9A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LTre4v7zus5IffjkBYpYJV8+UBKTDjHQ71BhICbxVcuYu00XSucRC7rfVeB/
tAshomdbnRlwiMsaiEJhlJGhhuwhehHMB8uyzBX6qvyQb5FLkxNlbnhiunWt
SqIUSwPvApNWZsgFN5upmrpRN0SIdK0Z5TiK+y7iB2XvYn71gGtwy638FNFW
2aDHWZwggJpWpROwfHaYpN8lOCZpc+RYMaW0XBIaHCsYjufkejeULNi+hoIs
ZHun2H1wxE5T9jRdjjzfYe/9Q3126GxWV/6WgncEzp0uNPCA9ua0Tni7kGRl
KREKZRQkPDHjMgZNN7JCKmQvMSd6ew1VlJQuii1KYw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MkPUslIJtgpLG4H515VhVMcqWAFmRPX2kL11aFcKSW8r1Uw3U52Mtrh5wvld
oxZ9RtIcTlWT6R6RuVBwu7VNs/g+ha6NGxRPGsAAyGDqXk5sKjdiB6+9tDhN
+pWBKHs4SIhMsH4ZjjC/gaaaWryUY8ThQGQHd8Wj4TQfeJRFn+aNxSV5XI5d
EPH6kKMoBafRyArDBDVqNIIMYiN3A1PU9nKGzjlvGcTYtqRCpbGnJ0WxqRmQ
spCqVNiqWsPUKGQtaKpZ+OasFac+mHpkTA3uywSN6sgp2y3C7pornEy02Sgh
S3FbGiCo13iLk3j5CvbqsrBMlshJmPQcybOxQk1xuw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SXZBJVU3CUA0OTd9FCfgF0s1ySnfnEbvlkr5nMMCl2NAuqC8f8tSysIcSsFt
WNEIEEVHmagYu4fYCuATBsSNxfUZl0G9E/YLxl40V7QiaFSNDsstrykC3+lu
x52tJ2z6SNcRxyqkJ9APAUd7tUAO+uVAiTjUzRZchN/fUEvBP7R87gkOtVDb
gpT7l5U9EKb3CoUO/m7h1M5Lgoe0373FlqGUa7lsAljsxDRrkFIl5MF02mPD
HhtXLGQYYthNGYQf0uF46pn39zYpK7oVVQxxcRlhUd/O8v7uM5QqQofP8gir
cDK/uRXi5GjAs0zW3C2GtLrpeSfsQzeyJS8wpKhJSw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
moj2UQrIXbO6T9hJFjlbnIS4OJVLwcrqUOwRO5kTxsHDgTGNK+0nPH9oI/AK
iP2NgfmBtg6ewXz4/a1kWhDxu643LQA6iK/sDHwHRKljUYfMU0TaBKbjU246
n8cjyVTcPrZsJbvm32xaq4yCZCDBT5H9mO0qQfgLaO3g3lC1KRk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
l1RNoMFRoendWzJxFISrbwg+Mo4g4RiMkWh2ZtV94yuBGWF4QCzK3GLO6dRw
hxRIec/vm/zRbTfNUcV9/lnQbbvvelgG9vKGFAS1n+COylY+c4C4fXturpI7
0dhGKq9YxIjEEXbpKqdYqChgFCLf/AtENIrlmzmTbnDyELQWFwfFRTWSKgPX
B62hQnHi/ozVIeUCyRGNd6Y6b7WDUWhKsiEpYo2wl+N9oeuQ03Y8PPEKhiiD
+2Wl2VtdojWyfnILD7yTzr99boxYN5JYtV/ePNq2CeVqaMjgdyfA5btMjfZ9
GOnLSIRmihqwohp8ghRT8evYVauYtOs2/ZaoYdThp3WET2rDRJARy8bt+w3/
dEuuhvGcSM7KgoE8qIdjHgxjP3aGOxDpjlAQnGD+0nKcvUuGckbgs8YZ7vY0
MX/o89VoowYEFQKNthwS3asiwpw/xyikPlxQb5C5hsiE0A9q41BLnYpdesSB
bsqYsUbJtNElU8d0+s1ILvpiRk/mGyNO


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TuN9I5V2m7Rrj1jd7CHqRSZI8O65rq6rwVb/Hyvqj3UAUEneno9ngEH9H+ES
VRcRgawZsoWZZsUSoIbeM9+47KazNGTaxQe/DS3Wd5fB1WKj1kTNJcL/1lyN
5/sgP7LUERxK6fxeOeCVo9rAjXKGUj/S/mhwezg6PNmuwsSFsJI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nL7sgTmIw1CDbfZTdZlsgjCp56IM8ABQ6bAurfEDv5O4//tEPBO8zQK1VYbS
7t+7tkyjD96bgHq1Hlk2XC5andcWoZtz6u4N31Q9on4CqR5rh/Q4vFknfrnS
cHyra1LXAh0MDpGJMQazQQodvHz/Ng+ar+aGa+1nu4zEfjeSeAY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15344)
`pragma protect data_block
c7bky576QeY9ms/eN7Ar9C0Rp32zR3UzNEgPCeFQvVuFgS1m1eTFjWLoTWdz
ycmBAUqJuKQaysHu+tpHnaTds6oQPMydwkHv2Da31hE/WGpsIfXvQYUZlrN0
J8gmdXPgJ8oyZMnVqb+8anwt73wP1/bf7+FbZeSWCZhdV3yQT04RsEm8iy2z
7DfEbWXPTabrM5ygVYDYbIQMvRcS1C4CheX8pWhf1mql87+TE6g7TqVHaECs
DK4YyTEUho5sOmZD9dwgMdqr35G3Lx0IInSaAHU1fyn0Wjtuh0dJLUWYPcLk
G1I+UkTKIuEVqfeAOLKQEwErk+lgatVCsUtuf2nd6wuOdyGm7p1fYGBzWODD
qPVXroubGbNrudIA5MA4flPr0Aednzj5Z/KisMTJytfGPWWKilATsILN+zaj
bVONYTPczv/B83Nd1AsUv1X4GYzDBsn1XJVdNZVcdSh3Vi6/NJMvXmJPnByB
5fcNbT0xWt3TFIQOBPBtT6xYggN94sdiLhS23QwjXaLik1IYXLLDcZIDWlrx
dSznZhkEJvOuaeirmNtVXCp5XPe49SlJZpFxdwX6kll4/17waatiGHDM7Rzk
pjlgLlnS5V1J/Z5OjRfS2eieNiLBQB4Q2XtPpmcFLTiEKsELybSWVdNtolct
y2uKHZ4CZs2TDzz3/BcBCv41hEkpGYa2qDekDmn5ziPVyzkHL3cQB86Nchb+
72uPYBLJ4sQaEYmoRBwyrPOXkbsbAuaWNQ1BYjA0GgXgxkOc0u9ZBBgynBVD
J+5w2aOAaBBn9pktON0t4OH9/v+HQSBqQ3gmZp6f1Uj+GPhksqQemWWZlSxf
Ilvn4JFdeCUECKJ+AgnQZMAuZt5SEfvQRMF4zaUuyX6usQlQLaFmPi86FjJG
n7TMg3DBXiu07UPy6BGcaR9H1uhMPa8MX0Mu+AtmqptgxaiUU0+QH+wRSaYY
HxUS7HytjK6/gR4KJpBSIGBqxLBDarCkjQQhHg2kzJXPdn5rtRvZ2o8Q1NeN
RXB4jKbB+dSiO2Io8l/xKTjKXoc3UCdFOeO3mIgtmuJ4+tf53dYA834XYf3z
AI6Dc+/kHBqXyT/RNJ6gZt6R7G0HRrbllECYMoQN2/0C9KZoyVnGiDY9+wKi
JjIIppAyroKz4CVvfDi9FSCdRibWucGdYqDdXG/n4qK8qgc9neVhQ78XcmZa
peCcHoEyjfxFq6TdYj7BJtSx+M8wo5PkVfFlM5aCaPoScboMsaLw6kt3GLkS
b6BGP3MtRYwDaI4qgouh8mDSYzJIMdE6i9T53PJPYXVSxoyRH4HjGm+MIj/u
oCzS/b/zVeGOgfxbOIa64khb5HVLq9g9oVocRDgdlQH1JriGx2n+0SyjnuLy
ioOay2gsLjFCAmqwx6eSjhstb/VPsv301HT4gTTbeSxII/rzqt4ioIYRF3BM
VJDJu7W0/2+k3SHJXmoGe6dLHYnlzKyz1QKhZyXt+t8uamO7IPqfdZOHhMWX
3POOau8AQIFVS7nYuv+49iOmZZ6aWbA8HuujgPA9h0f4Rt7fxI2Rcq8zn9wu
JUY0zEcLy//IMTFciyEmOGi17FIbEc15QNbgT3IdtvS9e0c+Gk/ZJK0C57Iy
1zHE2Giblot7w9QnE7D0Vw7XzQqH5iUCPZwya5rk/Ma3qHmp5iejF0Cql1g5
t315INYSWakkEEkmlCMk3Ss103rEDhJkV/jWpBpHm8IUfgqtCZYX3x32RgXA
3KjfTVSd58daNshnQR7mUjokhqeHTsCkUyP/iUAx7Z0/WvW/inyl/sqx29Qz
20FC1ciWoIF6VyyE/LDdXtXz/PE7BltBNffJZQYHUtM9i/wDGyh53bFKGkSN
bwtFtbrtVxUZ8CSC4rAGVPbNxYY4lqYeK7jHbfwGYmlaQ1t6RtJaj/p2FNAa
w+GDaU9MV6VSkopW1cxXRbw1Si6tnghGHIZQxYTHGa/TWhXv/n/D+cDo3del
GdO03ObHNi88wqm24ZX+kp+BkJMkk6zWhuTDk0EYMl0LFGj2oCgOgg9YziVg
DZrjlPWV114EB2p+kHbWFCoBCZsPl7ODb91j21jlViN6TAmkDf8LJmzJG2OY
Zyq7e9ItUXUdYnbRwBGt+BQS9sHFnN7N+lzGk89GF275LjlCbY9q9Zpm0y6m
TO+3aiaThKmsgwMqappkGlcLv15lU5SDAGOqoM0bAqUm0PAH2Iax/Lej5/gH
RYc5q/PXEAX4snUjg7xiE2iG0OhkPdn2no/o2BFGYZC8v+e/dnEYH4b/eOBV
HQIb8Tef0H8yZ3VqhxWfauend/bDuNLNziLJfcZp6FZkPBg96W3vTXiTMMti
oBxA1dWp9+dg4MdgqYEquoq37P7NkTgy61NvctT1nvD7YmXlAMV51pzPB2j+
E/+x+SB+5Kg6sqCJ4BTB3HnsDlmb8LVEQZvTy/hmVcyG5WdXanvAjohE/ZIx
SkP49YAr3BClv8mEQ/QEs/ASs4ylt3nziCfFaVwZhunn+MB1AJTzLcDn7gd4
HAN8yax+i/IGvGl4AVsCLhi/2CZQ+gtnJZhxobYEB0IR/eXup9WWMdVtGFwi
jAa/im87/QAIq2HTMJPMUEKuD5CC2BhKJkxSU2Sc8xSvZ+GSqPqW73/sWiMw
IcY8APRQQYOgK/SlSI2VLayxOaY0QwL/H0j8TH/ItGnsPnMddD86TnWQ9i8J
gUAsEvhrQ4LWA5j67ox7EYA6IdFhrqG3+TOeWcsErRCFYiflcnWYRiscBxjY
p+JzZE4SGpLW38TBYTfmmyQFSPuoktEj2bk2l/iXP2QQeEbxSyXAWoo/RBg4
CHR5JrZl2PGtXkFbGz5w3hYVUIJwuYLP0t/pyupJfl4Sm0EOOxSHn5T34UT9
Wjh8DdaRuUiJeDHnFapNv4X5wlOuHBffc8txeXj4T82HVprpwUl8H3e/kife
mLCjhqeQ24w1rIktiPyjbKKTxDxkI/RpDIy09jk43DJcEgapIfNzQFD6s54T
EK8LOAbEzPa938ONcfeHO28dCUZNOXCFoqP32Wxcjh6IwVeTTLSiipE+maW2
1ushGU7enWfUviWP92/wnB/3oCB2lO6rZFSmb6v+MYFCNaHrsmlZKIGA4yUT
AWD6+K4VoPwBoa6XQYulRUIPY/blt3vdCOWj/TJboMqfYL08PBmO7iHOIHIu
VL9eUmM7892kfzeTJ9Ffab94NRt1NTITBafiehCSTspat6y6Y0oazDQDequH
CzE84XDXFhrqzIm5Wo1eoq2z8RxZr/NiNr1ahXwfPjr31pUuBCb0tDbtxZyM
WEUS+NsBPvqmGHAY4GrznEjEmENdwaxKo560ZIgvPuwHdg1qORqz5tYNbZRn
YZnMStPcQtfz5pRVYCCftvkynxOJH58hyJ4z49g9G6Fk5/XurFKGroC8rKdQ
Wn4nSxUwWTQLlPXbExxvvQ3NTXWJNqs0yZ15MyeWzYEl8ESSKUxHIfSfl5fj
fcpzTIPnf5kpr2Z9XtJTj2GO6BfPNGMmTOm2JUXoxZu1PJPKvsbtx4329JA+
E88fIM55Un7lwqDQbZ/yjcmbjud0Jdt3ffBW/ZV/8cbrQeAzorlY6u0DGj87
Bp9tV7BxdhbtGb6LuopCwUl4u44Gj5R+2AJU6ins/OPeX+ZTYur5Q7ssQrSH
2AVGM7XXQEShMB+dW65tSTLzqLiUTOYBrwsoVlAP8dLLCXVeTCUJ53U5Qpr/
qvO3BYiVq0IynHOauaNSYT7CymY8S3j+YtyWwvi8RBmYV2HAvR4905EKbb4H
TZXyj15PLI7xrFLlJ7o9HB2EdN6btjPN8lMPTQy+yM+sSPDUJhSE7olfMi1g
QO2lX6qb1/9fWECmcori70GPxX6FU34UV4/M9+3QiioIdDiaubLzy37Bfu2I
QyTqlxJAwMhCNo1efgFO+A19eG7b2jEahkJSI6abMxdXY4Nokc6547wFLk2D
rRlrLY1KJCT/x4FrOblEAUlPSqAkdqD0Fjfah5B1gnuPN3WVhrUEw3kt0dha
7l0BW6BcIpxfBY/IJNqAxvYEFRI/qCCB/6mjC1TFYIkBs4FnkeinXVhVbs+Y
0mH/zAAD1ZpnWXTRCfgzgiFd1+vgi3wZIM7KWFhP9AYssDSjG772Exd14Qgf
DhiwjdV/P6OodjDZ0rClV3ftdV5Wx7ZGXeSl+cC+G8KAnJc2qN7bZALTDjPE
OPBYc0mCUFGEh+IePwKDZ68iA4ANJOQOzJtZFHQDQkH4t07oMLspXacsyP/2
CFh2OsZPWVFr4jvhsI3NllTo6LpgI4MPhuuY9N04qzM0aGOAdZAIpDQHVjaG
YNlLjfykN+Vz8xjtiyY9J10vwOS2TGQt+3lpP0XqDHQo25KN1w8BCCm841QZ
yYj29xVR7zKC13eVLxUOC0/0m6Js36Zj8lrFw7NC6ZPpvNDO0Mmurf7TZRLm
tEj4HzaJOcNwrzn/tDGRFvk652XyEvu1kqJ/EtaggWZZlSLLjEdT9PVQenZc
PzQUePzNouS+H7pkalndrQ7A/7gM3HsorWv+UxG8tMb5Ur6u4n2kHY0OueYJ
OBehbnlBMw+44gT/Dc+hVOsJnwcna31EwvyiNx256IJBSM11T8ebnTov0f1d
Zj8DQE49LwE3Q99wdFdE0H73mfhWqEvGZTsqRyvRdFeFQDa4tFzSagFyk8Ba
w9D6cU1Q4zjRfV0n9p6lagCKGUC75zi72lIyv+FMc/e6JJ9vsujTPSlL3/T7
1yAjapvkWnSTVz9Ko2lvmcG8XjWkhh5o9LxrEC89skpCRvM0InX+b9UiMWlg
dSuqsJa6WlrTZgJd+U46LDXZlW5mCSfhNdcPoMhYhGfJo2AS4xrhI/ytBMP0
xkyIzSe/UObv1FOCmEkYE2lBUjphZenF3u3TCwwP+zPlR4fRRwimtqvUi4dI
Zp698h5szB+2kYwfvGs85gFfh2YS9Wlq1QWeZjD1Jk17abOFJENWK7Gi0fw/
6Qm81z3rkt0eXxE/lcJjeTZLhz6AarHjgKepFNE9jCu7Qcrc/Y3CuwAHZSs3
jApcMh9KsVt+GtwVOikuaQHLVckuU+97QSYzRLCHqprSgKCP2vJ6UnGfoq2V
LeugVkzgly4t2YPxzkwlKVvYzYyfONNbiYBf1StKEd6SRn3dq9kQ4F4t7ovV
XqEl103Q4i6KUwSofN3F1qg5AaQF2sJ128YSCA7XI28n0UVB5paIBvD4+DnU
c3yc+/2lTD4y+URvENf5M6WNQHglLZaIrdAjQ6xsuqQVSTUAsLih7AYXjB7a
zXrCu/4uWYtW5uonKE7N4mZW0NiOimgqZR6HBsihK8SlShH29+ZLWX6R0kKV
6qf5dWgLTPYG4FnqoE0OT03tO64HS3i8ATUhSEMdnQICydvCzy9/KNMCrBxH
PPpRRuks3Ja3Ti7M2SBZfcqNYRLvhMI5v4BuVUV2R9Fpdfm5NGfbOfTqACM6
qCh/GIizX6FrAvx36hwDp0gG84l1+hEFSOfm9HVsBZ7UJN2PJu5evA1CfUUL
pOc1BO2liiSAnfycdqzOdR0lOoqKnMgzn/kE7it+ODb+VRccCzNYPsOZNXG8
R1LiM9pgYpjfhwmSHSdg4RhvfMGfrnqV3in0WuZ5euzOtuAGbGi/PqaBWJdf
R7X//Hr8MA5fUktpAzf0ESQBTW/eflzMmPqKLNr5FAo1DMcdlYrE+nOVig0y
jEEVRo8F0Y2uhJ0mpqgq1zdETFrP6G8Vp3rxnDp7w0QX7k3CK2AgSwvqydNT
2PfXnd6xJUD3hnehLio4zSTXapQZ9CfbblIv0cLiY88Ss+1C7t6FqVQxLxEd
+0cbgfM0VubwOqfckoNGOyuzRyADTQa/RKyZwecvFMHdoaInMPtvOr/ezrJb
ToZv76mS6P9DJZ9DiS52sHCLB6ldUgbr+cIcxKKpP/RAJQNkvUd9PJLEP9ps
1llzsCjH54VLKTuR4aFp5YSTOqT0lBvtBMQgGy6tRjeGqbfQ+vzuYixZVmqK
zv3LsBLtlixB9/U53ebIbwsIxm3mhqb+Q0QyZFDG3gCyDAl8hyG3V7aGn+Zi
iamurWw5vHiDOnRGmCHP83wFlCLiQb56ybxru1CVdq7wQ5PEOpPAu3aCYlIp
vlvgHN1z4hDBa15fJ7Y1BpAwvVI4w+efkqMqhMjyAI808W3iQy5q3PtbLSFN
LEmTU/8Pac0RG2Z3tFsAgph8EK48GUrZTkDF2Y7Yt+gfM98cpRW2BbqEaZkx
05wVbxl2t2E0zkNc8j62LOZoBTMqdyvBDisiOtG8tm6bZ1xb7eHjbjC6JejP
xfhcVur+Zc2SD8sjZ4aJ6dW0X/9B9MHUjO16Lhb1JgaYLQO9NGNe7syDn0Jo
f/C3Vv9AAVW1+TUQ2TwnqKmk2NcyVZ8lwBEAfCq9WfPH3pLXswnub65zYdgy
2P0ZMynLTSXox/BZTYZEXAoDxQmrYGxjQsIOgb7oUfr69jDn/T9PPCIogYJ0
8EkS+xihK890EB7W33XhgbGed2dkOU65ZBPlukAn/BXthqmhDtekA3ws48Wn
Fs/kHnpDGmJnLI09aG0vH+lBmvcbXsMr0eHqOSy1QLlLA3DGm31MfY6buvRk
NBxHPG3sXJDsQUEtN+BqNqgP5Elru/vhgYMlNEY0ljdHuXVwBh8yMdku79OI
gkbKEsah621cmnq/E+SLPYjJMf4MdFgDJ1OQSVsxqxPxyqVx3imqsHsGLchC
EBeFeofNomJzf0uCp17Qxxqni8Y/ZI8NjzqVT979YouJGAK/+uJRHngGiIF+
XiUjtjkSKNoMO3DnFIolPMeWOQnQ9SvHMYaH6U0vucKiwhqdAKnQfL5CJEPo
62C29RSFkRNVHi2xgtq1HAWwwgHaQPe8/Z5RS9hPXsOISZDgDW2IED+91vo7
DSR40ith5lE5GTVcGamthrXnEp4WzLxTxDmRTn3Rt7ruIRwiH7laOuq0mGgt
QS+jDsnsEY6okLCNfTeVlsXb0n5wlBKqpKAfOsq+SG3I4XY2dVsUuk6YB/am
K81wSVadsawJWB3vJxbrAyWneI1azMVMDcScCimg98kcCISkNXb7r+w1GgHc
YM6rZ225bYFzsqGWYt/KL1HqmXT1a9mB3B7/ZoJ8UlNngorApVbsmQ/to+jx
CXObPKaHL3aZcr3hIWbG7weFox4DKlFoTlobYRZ9HuVuL/Tqd+sszQgOml6Y
z0Ha/wMhwsvXTG2slVTvFWJcJdvIHPrAnM89CiIekJYpa336k8D9TeAI7E7S
B+cKbI9d9WrHRwTx8jr/I0renityrqxLjz7QgrxwPxJJYL7d7QZaRUmAXj3l
0AQvNEETtgoQFTQ6udQwdRNcwiBCy9hYzR7rq/cJymLuWlf5OYVuRqNh+Kwf
Po7n76yAitd+4HEFHD65CJrnW0c/AfmiHd3vDc+M7spHHanSLtvxnZ6hEgZV
aJeb02rpqan6QVNbpBnQrPAroTt4FiU9UuZR5pFSf9cs5t/tX39ba9Gc8r6b
YSrJocUCP43a4JkvJI+SzzSHutwYy/CZ55YB79SXwmbz+XJ3j6+b0cQPWESF
jIVnmEZ7/L4JrrI6yCSwWlzEldQ3oiUXnernef6MhU4/lNBWOkhvL8bPm0Yb
4N1IW0oXu/h+jdpy6yuYHLMiiJauqM7WvJt6o26Ny6XY2hv49YvxWc5qnD0d
jetaQtkVybxf0DIOaTuypsOslfWdT5cRKCh+vWl0/tMQSh3XeJkWspFlTw/a
uLVwboXoKqQrJlfx4oanQGgGnrdrIIeXIAqW0gLVXWR8YQAk6vTQ6l+5OmA+
SLnStW9h4/WZtZoMvwemrugpl1AqK5wrG8/vBac7E8hrmziPzwQxy95fxhcf
OrWRzDOrQmDtdDq1rrUtcxbWnudUJcSvmZzdZPWJxJmwoRocqEHuOThlTvi0
rtGX+cjw20kDEggd18JYGrrPRSQeWZfoaKS8ADd/5I/KQ0tQlTa7/z/GgsHO
m6GAYWGCUrufGdZZN/pA3ar+ZqVl7n70obfROL3LR8jDQInS4/Y4854T+utQ
SfSndgyaM3MZHwZG9YOFATvcixemzokionqQDSk5Vk/6g9ehoXWXHmUU00MQ
w2DqTN6gHSM44L7B+SxJtVgnICUnw6tFgCYdCp4VoZzFNBmpWinjSc7gZtd5
9cZSdOzLJMdlqpR6PNhb0REzlfOPtReuApInaEY1odu6lC7t4JWXguh9n04Z
b784hsGsj4yoa1pNsd+AeSnetwEo3M6o3vtzDGNDvaZVhKRijD6/Oqe8iNHa
jvck+eNkbL48IhZvFwXJr0ODM31SpftqmouSQZ1ry/znOPRfFo11nTW04V6N
7YwdxCHQhWQRMnK8ZKsYDST7jm0hSp8sBZl5siixhptxsf93fTA966YzjdS4
26RcZNPqSfzp/h4fHSIz+OvYClVXXqyjIzkpJ9rYkugXeYRWzrxZ4qc8xniN
GNe3ljj1DbXZfTTWvMqEqd/3+T7OS+8Yv4LbTXpOg7d2xOsKs+LRvgtEDO7/
EopD+KXOmQJln3XZnZAAgEMoFYa4GGiJV3kkBzp4SpQ9qgxLrWObdFYOexsz
aGCgowRI70SU4O1E1/xnSEKQ5SmR/+PP0xJHI5xmcJvvUaAgY+yBTQfG99yk
TYKk6IbfLz1u/rufudXP48IUkDk/snDSqyzhrSQtAV1CuPCIoO+0TXmHTSrX
9hdcpn3sC+JACpDx5yywClRLf7+Uaq9PCf2yqUAxLiCh+RZ3EvFAjLo6Apu7
ebAO6VI+xFrqBorhfcbtetcYtBnYRd2kgitsZ/7OWNqP7Ba8/Em2Cc3tZvX+
xJDAdIHvkdti0PKUQJPHOqNH408zp6wYt4NvFs6Xizy0gLZ2NC/yXNa13ND5
QvZ2Swq9RkgQa6YM40We088M8l4RJTu7PGTwatFoyh5HFI0Xc3/1oBJO6OyW
x6UcQ9N9C8pealyGY5b5qDnA+iJUAkxSx4MvpgD3VBW3NVmAa14Wtpa0pWMG
iTPmc9E08mF6A9khaVlVtAwQZCTD7Gie2svaalJO2GtRWmgL629vSznrLMRm
VxOuE2xzQR+9WF9GW8kanLRsMF33nFjEBwafp+cMZFBc2icjnJXs9xWCfjZv
YEG/bbWOrlEsDuLx/nzjV8BY/FEfiSvL34Jte9pEInGa1jZ+DcSg2bHTQnxn
KHGjjLAPCriNZukNNKqpZNUj4kU3UV5O/VF1W3JKsfut/DMVRnNnObvQU0NT
ApwMbHAK88oU1o8GgOOjUFhZF5Ns/cnUA3RzvLZhnG/K8tN6UlODAnIeZ7y4
sSvJ9YElFyQ6+Xvuy4i31iWTInqIug6dMohWlVoNGmJ+opYa3SkMG9ggtUcv
DZvT3rY+hw8OvrVuLATjhNFIWPR8f//5g1t5D2rPtkZY7yqih6YOwcT6lF3L
NmD0iYV1cKTghpPmpWwAUjj8WuO3IzXlW0q2I5YmGV8eC9d2JCVBRkceP1qr
IiwmTVmvjpGZeZHvFrhYxH9W7ModlHX0Q4XAKwsQmxGFe6YM86rtr6TL37aQ
8ReREdFSFvipzJJEfOK3Jgn5BPijtl2bQKXGGDk9b32wrpwdER1cJmv1YGNE
vC4oHpEdqtRf0z6h8KcRAC8EiSiTmsDTJCfmn27ogMEzX5ybdBUb7k0jfHmJ
G+2FRFQyTJNA/ptAZalP3RHrBE3wg731ChKZ3yBrV5+K0ff0nBXsnSzaes3A
AaH9SjEeaJ+m8VYf1QHA6EeAM2gwGJO9kpJFURsncjed6Y9dDiQTDHx+5bSH
qoHWflvIqt7VvNuO3RSIZcGX1qese0wLdJiONmvjCnLE5ecD/QTgnJ53tU9g
kkZ3b0zFFb1zXCocLaCiOHek4SqnpOdoM/hlhjweAcNt9avH0tZwn61kuicz
RWh+0czcT8YxlTgt7DgkStcwZEfaNjXuRSYT5l9RhCLYJ8kOlEXuEuTq7i6n
TECP/Bo1rIpgAYxo6uB73HH9/DSccaPO77aSwUiLGwgYWRFy1Gs7v40dgZAr
7mRNPl34rk8uzJ8BJrz4WKfD+mDUCWXMsQDSozNuyv4fsTmWBgXq6B7ftwn+
JojHp5RqZMqZiWwkivNu1FdJb9Sa1e2m/WluWjekX/iz0pdsqryk7/Rriak8
xK4/LXjLiwiuGtUsTueSQn50xDfo0QYknDYAK244Umqokt7HkheE+PLo1Rwh
miMtQfSOODc06peA1Qo5rVNnsD5z0mdYdesOh4mtoNKku+/Ab9rW2XragHkz
wsVZaUVOELtb3z74t4BRim4wQTreQ6Bm7uUaGLQm5T3sdavZSPJRw1AW7TX9
WKZknij5GzqQdoWt2jK9P4HBtFCaLXf720v4PKAx0ml3+9967xDdHN0W86Xd
8TnPgc4jMFRkzpff93s7lzY/7EYkmWVA7dVj/9t8nL8bWhPRKg36lIZg6RAq
wUuCZYO2AteHJmBqVFM6QZwnkQkSG+LhtcVXkGhEQ8gNU6uSDKF3kS375/C2
a/HDqviHYGovtnwnbN9g8/I4c5LWvRZiVww2cIvuT/zc6jd8MaHQnKiyXRcb
eAJSL1QvUuMXvYlFJmtRzlWY4YqEy7OeFTNZZKbEPv49Zz2zjE2IG7gelTjc
1RzpqGjuVwVBHYbF194EAKVIb4jk/z/XEvmAZMOLWZ1Sf6dnGJae779oQUWq
B4wojvl5y5KKXj2nLbfY3sNDCAxOvlwM7cn3evILxaxNuVusnzYx+ypeo2R8
yKPYnFDy16L2FhDc2UkE1xW+CyOtC3NFvxlH1jk236y0TvCuVNFeC/sqY1bB
6fQ/oeLdSMaENu09IQmrzC4KW1ySPSGWjSIImXNK7NfknGaaftesGKtUlH2k
mEZ8zZh9QZdvQjgZUV64+REROcZZLPgjJK1+zMEzbq6FZArlyjrLvWbCRPn4
B4WdayP08MFb9Do1IABIJmDY1J2uvpC6Z6sMfydX61jcETC55y4OyVk+t1Yh
0FMgg9bHrHPhlNNkQUmyoE7N8QoUQuS/LMfnjUp5f9E3in4QPsbaShsv32F8
u7hlO6e/JZ6zkd5H2Ye37KnxN7JdHYFD4snPR9YZQW9ns11Mf8JDCZC5DE1k
c11TU6lPEcLjXMMRvgRsshWXDBEcZvRBLj0BISVUk8RghhYZ7GpODQht2yL8
nIEr6tOTk6bSgXECWMlse219eoMsFuCyiiEPwibbFrHhfsDQ4GMLimyS8dGC
gn2GRqKsz4//DVUxG9QwgMAMh3KMJrGFF7MeOu8APW7NJIoI5EDbj/OiwABJ
MUg9pZcp8kW5OmzQ2m3wv9NSfYXOJ0FrOVB5ZOEDfKKCWnDYrO7cw7VBRqs/
CDu6BoQ/8wW2eno1ACAqkCMM2VNUgS7Pb85OISPmAm0Nikh3tczmm5MoWl3L
Prmv6tpD0e2h29v1B7732qaQifQ/9luWFTBaZI+ofj3bu/XqJCYqWP6p2G2E
koFprtxWpIu44p0kcSOWQs8KmJktF9ihcZXefZEwSRWVoebV4Fm2j4Q84cuD
AhGh4p3iN9GaEykDjs6+YB6hAhnbV/nPZPY3V3sJB71RBqLyCMgc+z7OWeqq
13aoz6FUabCf5jPp+5PhXdMF9iKF/1F7FY10LrSux9esRoqbpGlxHIVdZGWT
4yZ7cdU0wiNxiIwMZenaclEwgsQjOT1Ias3GmNkH5/eNHcLDxcufBwJQq8B4
VAuR7KcS5nqHhPj9nPNdsEdwj0fT8mx2VuvmI+NxPTv/cNgmg9eUrOnYJwTx
dmAscIoD+0I1XcENl9MlrKzn2N8Ii1KqZIgTGtQlVPQDc9lb7wHH9B02CAMw
7BfhmKRBHJ5jkZXbfrUDoK7KLINm9fClIFCIH2l0QmOzrO95VM4iZl/XNlaP
lxhfLXwsB70w/sOtAVBsqe7S8KAmy8E21dnTNcgcOcoxE0eYtW6usPtDQHGU
QrjoehWLlt250np/02gXzX0FzfthKNsueaiRxkTLCHm07CSG5AzeoBqvkxPY
bux1pSXxxFXQv3js46EfeDc6Y/kmz7li326QJvnFuoTYM2zRFkTvV8CPrQds
yy4L0q3YZTeQjNuDOxEewCwqLfurOGrWDQG6cmFLk2yfrqcBOCni0lfvF3EM
0La1Xd98cXJstUSCiK3b4GfUv5dIjTRmoV59HYeLpFUpEzJmEvRLB5tOhNap
ss6x8af/O6mmwJx4rbYx8crdDitjOkYQXWBuBcP3QU49Pr4d9NBpYaHklNsQ
bIY2Ux/+qIHe1qV7w8pRz8CylrJ/TYB95zWAi0J4wBtjxmUCn1UAmOz0khYD
nnAmuMZgSi41+SVeacz4WPnLGh0psYNMQTOoBGXvPLeiFCQZ5Ke18wMCN20M
GQt9gpU4ShSh73ikgGBTc05ZoeN/YWUfrvJ3qPXy+L9RTl0xwL9Z97UbOvKt
JtF94Bny3ug2wwKU30wvhAQHYKx9yRpRe/0Vdu+SdUFq16vOjAQMza99OoKI
YEpiaU3khNkWH7E8njdlsu68AvmfKWxYcWY3xX83WQ0UYYueybqumLi1ttbr
h2sbg6evt8SALu4VvNbVm1N6Qo+eoDcmcV/R7pmULXupa5RjCZhe/Nv7ALxN
jb3uQBukGIfdBIIvTb+AafkeWbPRlErDDhIcv/ck73gGMPcqn+53ahAzjWsL
o4aNCCmu9DMhEpvUZw5RF6oCDHQn62oQ0pW3jSvxCq2aBw2fVvU5Y1EXM6Tx
aR33Se9ppKd+CfyR7gZgyg5SN3E7CSQXtsNVH69iB6aUkjuuMx8TEHrPke3W
IEy1xBMTuDugYbdg80lxHmIAbtZygwrSkNa8Ep0LnO66OGuHACXIBzRkn3Ev
sDnaZ8VAaQQmcIe/KVSJ2PPR3pu3EkACox6SogxfHS16fVQSa1gU83ctVrQV
yjJl1XlTaQzmDAiLYUsU4RMolmepRfBfFRyUr/UyrmhWCuiowCClbKtsRn56
uYkEYJxgpl3DrB/sERz9EOf5/7ZOhUPXcwx76vBKMYcAYgiiEgg+eOUexof8
HvtCC9jhINjGKo/wCh60fQXeWugt2vhSbVVRWOPTbw807axB2rjzVt1SzrYg
EScrUp+ouOg+kxPZSRi/rRJpwvvtWX2gV3o9NPDfeAMQFsTDD+lOIa1Y7uDa
VCPfXFC84/u82SYq2gt3+2XoPPKCvN6eg41l6RJrYJXk/1mPXNQeiTbCHuol
r1/dWNuj97TVGnk2iyTbgnVD1/9TU9/pBOs/klBlHZB9d6z6xFfPJ/29IpgL
6r0EwJlDaSBGfPd+eqZn9MXCKOWNGPWdBdqKb/w2hdCEvvxB5P+JJGrS6PII
T5xzcar0c+pz3WF/aW4kGmWbnZEy78uR3x7DzsY0hckX9n2AnKWRknlptznk
WXSQv/J78VwueDkOsIC5GXzckcnfgEO8ba9xzfbALETRz45Se36INxjZK8NN
O3/oP1LXz8OZZ3u5iJw8ZDVYBRUUqK5qMhBU/u8ucHyGV28YCQ2y5ORU7hSW
DNZWCQu9260v8ECxMkxpCgnjLNCtEdMSDyXscnigDhMrbqIPa4rVR3v8WJmT
kwot8cs9mqS8fi7ZlMLl9M8sVbzXTrHhT8tz80Si97759eg9Kq6Cm2RZ5u3E
WrcXTFcCeA9t5YXlC+mw9hR4Hfa3NiiTkSdAVKu8LrgRfhnGnXfrqLk5REjT
9InbClNXliA2nO1rnAyf5kEzp90YzVRcLQEiUOUh8RY0UofJStraHnrPPrv5
JI5LaEb3LlCxNwbBD8G0LagTs8aWb6lY0K+Fd33DG56jG2PeMJNdd9W1u8X7
BqL8Btoa6FCHQ8gf47R6/GFb1Vdw0FNi4nWkt4DUViHdA5Em3HSz4w2lNEq1
tuphwfeIv8gUPTmvV1MEdHwHLqhQK3ygV0+GUB8GhYaAexqvJgzoDq90pdoF
vVr+X6Y0SJ2lumPph7F2wD6e2idiyhEiOmdUEEe/ji8UyM3emoveaPz9pacw
ySyEE5gpl7/8MTxz/biSz0fN/Rbi41BY/0saKBWylHhpp5BH/jeI78+rwDxK
eWMCV8o7AeZTXWR2zdUgc+lFt5Z1XhROhizgkLhT9bvKqOr1rBllMUwXZNvE
LUrxOZ6RQXhSed2e6wAYIM8qCMHXylV2BF90fEFlosscSz4fRoMj2grjWKS5
onirlcH34ha4J3OpvbV0Q0v7yg+o0O4T+ET2rUnG3mOGIUrEiwHTZ4jHiG0+
26xATWbEepIyQGKGqkgpoI7h113zVjp8IT0xrK+5gSdZnfsSjm2bvqPEMm7x
HoLWPQROfsCREVNnmRIfxBYVbc+fFQLFb9xasoWPTYMuSAN7BWfRvF/iIPQo
yKX9pVXX36NomlvI7HCNB+oA2reZ+2XZzPaAE3NGvXjZc4e+kpOwN/k7MeuD
RjVZ9YQnFfsC5OZUjUZznP9d0EXWXC02c8SP+8+wxxoQGGCcySNRTO6PvUwQ
G+VV01IZP+DU+D3R7yF4nXiwC5ljEb/Q9z3FtPIWvnzubwxE6xCZEtKDLRn2
htojxEbHax4qGrctjT7qSuDJXWeUZd0wNAKtKpDh/Z25hr+k/o8uUnVqvTB/
OwlbhHa+S2ONd5ZCWUFYzQEDXx0ntWLJ9P3ZrAXgai4RWOw1E+5vsSPZmvpR
Z++tAkQ+++dzpCrfG/Ofh346agtyI0EG20WtIuI0n5bHR5XB1kdKWmkC2Fo+
K5VYbxa9EvXu9Ci1R83qVcwm/Rk4353w2z9K/p8vYmovO/MzQY0DpcwVmvFI
inaewPjcAU5mLNYVuUlLS2ICsoRxtvqL8SMq3eH/eX6SLCQbtKGpuciiuNhc
zCZDMZMjLCtmNXMMuNFMCPXCW5rftO1Ko8rJ8EQyXEQYvb9fhVWA1noC3QJF
6kBo+fLNiZ8TngmaQouLt7AyMKX9QgB50UbUuDGZz97WIEGNStS3XF626J4+
zvQRQvkgkTyB4ClwxuhpIEXrD+DlEG44bE6QY6E5o6Jh+orRVgPVveCAUs5g
dlMUGrhG2iTfs+pKDBfoytZjzpRsBb/muv+AcWghhUKZpdPf1cXS8paqHeyn
ID9RodfuBBwB4hbZWz/M3j0iNP4R4MVBk0QTO0wxUBQoX+s1bWSQUirWIwd0
BjPlqWRr9J0Rb8ve3m6uCp1l7Rsf7s8mAx31WZ3XAlqhHE+NYsAgVIZSKqEy
hEeiJeF8HsU5h1DyxA5dj+lrqdGnRDr8lf7uhCgkKq5J+2ViHZjETQcdWx68
rbgjhNg5mNiUbbCTf9axTeEfHuKmC4rm+vRj3CyxLkuQMpn74/XNaTZHykBC
z/DaB2s5diqnSrCpOGjpiUrEKm8+l6vbuBUwSL8SIO5/wZZLBlYfbbQEXJhG
lKoX5cl2CiR8lx6VrX6PSb4Z1oBucnlRoilMK7vco5BGaQpc5uYdvFfZ6mCF
wdcthfpj81MnO3arHirNu5R3bz7sTQrxOa/PA0LTDKu1yjqBWIGFgnU0mqck
gcALHv6CsqKivqtyyvfVv1J+vJqB8hCmCposzDhyw6HKfr4QxpFV8/zbkFW5
uZT54fswfTNoWOOmAIPZ2Iz2tZc/NzdQffviiydrEVUpFYAoojTnLUmBIOPv
nzkso3+7WZlqmKQWiowpIdMsbp6ziRG1kVSt99s1piA0U4rcPkhreWv9pgpf
BDnebAmhlQtXLPKB9bp4Qx+XnEs0Q6F6DOMmBo41d8BYf5i72uaJXUy5x8+d
KstH5sz7sWzvj+egjh6Bpw2l+Bn3HsXXK6GSxm/uim74N7I7rYguovO7+xmu
ahmbAom2F1TibEQYq/QUysr6ROfG6pf480sMIertfmn+LofghLGwp7eYoyLG
fqyCi+YJNR5moM3YijBQlG9A8rGLRMK1GR0cSh4kzCYn1LHoMzDQrRDoRanR
Bq9g4hCiMHKoXuYrUG4AmHJnt/Za6J+e/Ih1o/e3oy9yJSPfBB8tJ4Zjwmi8
mOGYPwpLGD/2Hlx97foEDVwUcc7n9ttO0j9T5OZQTAK2OJ1MxScjF31Vvu4+
CqIVcVNgfkj8qEr28ioTki08DvOg71lpE54ztKrQzTYqg/j4uiq62IVxznPJ
2MF8WaI8q6esTaev5LG689U3AiTfeQvVvJCoRlg0wckqNDGD4yT1X+1mqJGF
3rqYaYCOZxX460K2Y3En2QCF3Z3mu71LQZDALkTJvJrtPeaZk0XzjrrbgISp
91mLJAR+Fb3WZ3YFrGhuuRdGSMCkaF+w6+wOTxWiqa2fifzQsEyXn6VUEVwN
uoB4cj0crWC6yk3o7AyGJdoSR1WcCkgKBw/aKgg2sTvHnO8IGQdoa43bVvzl
PD0H+3BBpcPjVqpuDkI1tw1JlO5VEZeiKNyYfE69bCdaxggkB9/DYoVYESBa
TwNvMicJG9U4jbhqbjTpfrDcAaOHfbPOIf4WSZPbgFiFisCZ9YTBY/96+vZx
J/qBg+UDx7iqs5RqdiQx6A1b6F9x7PfTtSwObk+FJpmwPDy+SN1t1Vkk2vfu
DGYOQrG4+uu/FFHKKeLuDDjJegJ2sgyWKNroF4CsoKrvixdJfqGDbMxiS/uN
rlvsiV/WrVXY6mvvyVh1ur9ft16LqAfV+vXTfeNZbxUMeUE31fzOzwk15odv
98vOs3aNfkBDES43I30qQfbvPctj0h47wJfBVPeuX2ynErTJHC+VvUynP85X
E57Vkl1uKnDlxjWE2TttsAs8fQWGCiVD/Soik8eOIT472f1R69edn2u6MELp
2iuinm9PW7TMDrQcuoP3eSKrLE5nUU3aL6+Dq3bnmKFyxUg4J9vzMSAxzN3Z
66dTHe/8m96ba9p9b99qVWQ7QCMeUXeSx0EfCQIqY6nzkA7Gtbh2On2tG8pW
Z3FnRuw4kCVouHrc2Bi5PKQo2dcMDCYhdLExbYp5ifEgLCZGgUXBN4ZEnWgK
J+X51eowXZc7ZUcCTBAMV+czSJSKBK9Sd/jS085pzCApsieRNkGPYYTzR+Ip
PftCZu2MvjFnXoy0ImTZoCtMmnN7JWd4OTMW4peEJENvuQbzfoGxwTdo3sQ+
pM/tUoigKeRdkQzFovvULBQXSbaYY8JuEsP7nOlMKsqZXRT1tEdOKxwz/F26
L6lLG+pv6TkBFeor6C0XuU7B9CjUdHTxdVIQit+ebALPrzSWrOuH9GzAlxyx
8ljoWDB/RPlKwwyFmI2CbY8AAEwO5S374cehXdXiS2gwwR/OxcP9wO9377UA
EHfWw5r8Uw3hDQhwZYo4kOeJIZ+EJ58toBnZI8hDKVO+Aw1ExJ4JyRhAJcEV
aO4GPj1R4K0lWTc+o8SpLczNZUFXmwBODQdbgyuPeGdy7j78sCKYrJyZ13dO
mAtpOcaeRRXuD49hU3v5Z03ZxLeoxRGR8rhF9d+i+xveh8cs9g/PpbqrFGKs
Ax1lrBR0ETVMC29SaqVVPkVXJ5frmxcSFwWzmht845dhkUex4zMUl/c+D4Bp
RvG8ZnvaUpUW6EWlALo8+u7ftEnbHl5Ar6XF3IDJNvTnjJ7E59DI6zYITEtv
5aI+j1+LFJACCwdEk8J3cl7fZrbJ4gHh+dNJbbgIsiF8om1rMswDoIW154mw
EDxGdVs+B8BCic6LwE7xtForaZ6qOoypmfoodzPRKZCZdnzs1Xn9lNBLPfYR
iEcfC6uulYDAf6BpU9ENnttfIs4dLuYfkKWqqP5/UnLVNkrZwGoJ+NorGMyq
OlgdOpguAwjWK+8ztGsN2+6PNuIYQkLQ1HJYMfW3YxrXtkXMHjsgqfyv+Z2y
8vAcRDK1sfnD40MbFCzo1xaremU8mO3KKWxmzVA0tevFSdDPmSVwKlKSiRLH
vBaDjGCjdTHbjFswf5PLe0onl+hcHAcveRqXhiu8fscMmxM3seFNNcRHGt+v
KeiiLVu1S2r5l95LLXH817IWQJBWdklEF3LU4stEaZBbdF5raerLHa5vf3qx
/8FJcpPZR9W+5ENhy9+U0UKB1vAsfsxCEE2YOrNQmeQ73LnwsryHhKao/ja5
dRqM0etaxKg8HDG6oFLZ9FelC6gnSvACshW6ZNvzltZMyr1+OejEokRjSFWF
hHGe5DhVbcrwdD6GTVKx0XbKKEGnWjGTqQt3j6dNxPGLD0HlfwafXPrbF9ZQ
r9AujsM8sEMa1io0nFCJPGoWgDnYirVHYGStWXBF+RcH0o2+eqAtzZT4Bm1f
0vQkYuUN1EuFG/C2Jt6ZvaO6opOLGf6rbg40l8ygSAswAkPa49ZnwoKk/3+r
aZ6j8xTScr8sxK4bbt+0ya1JgmRqF6VmQ1j2PVVj4X9nYdZI1bJXlNDkYFAG
BACCasT4lhw/C6l5pOGytbC2JnByjrXghBPrFpzVMKS/U/Gs8zpBG4m/SGo9
aMMDHE7s71yNLuFRR0GL182qiBXEHTZyPovjjuUqC8ZqrxFGkzn6Fse6yUFY
kR9l9qsvUpohLynnHu8thi7MgnFXX5Kzs3oyW09VM631ljcdspFHSnIwCA3g
flz2Wx0aCcDFrZ5SGaYRXLl68d2k6LPEVf87PnmxCm36edwEE0Gkd/OlerHb
LUJK0rwRMiVGjO+MBs/mn+tGr0YykAle3mIc/6IXBwH01yMsQ8knWWASXCWU
zbaHOg6+KlYLuH7N5S7n9D9uhDP1ghQbOy13w0DaNA9tswqJQ0F1NuYE/sIk
bUrIxrsfxpnXHUXcr5okyiukhzA+K6p42lg1xEhLYtx9sg73pfZFn6mZvZov
pwSDu0/wrO//KXFwno2fSoN+QYhtGasx7N8PqVp1pvIQpEcpxpyv+9g49eiS
+R5aqJqdpoCQCf7mu+TBnULM1kK0YqP69tDBdVIrPol90GggWO0VvpGvNWqJ
mF9xc9zDIUVkXcb7yxoBblJ2c5jBgCjYR1sopm15DsWwWBVE976rzz35tura
MHNW3tzyySnN20Nn8GFN0+AM4x8z0yt521npPVQOtHjzG9ZnQxkiuT6h9qPz
oD9bf4o3NOLT0NBId8IHXLoK6CNM6dL2DbHejTbejbDdk7ykwMj6J1nfHcgk
fOKf5/01GCpW2/txfH6cRHvFfYDA0xWzCbWXlgbrRHcy4p8sWlSSFJ13jGlQ
TEUpNuMpHEiAdkQX2u7bz1B4cgz9HjE4A38uBvdNU1pjBmVcpKZouVKIGAhy
/q2s9+p0TCbeZe1C+S5Ituk1np1AZkxGf1s/XUj4tI9jHKqoUSZKRwD85ukw
x+VHBmu4VNOHoFDyTITG+S0qwrG8WPU4NhMZhOTtp9RoiXOSQLZSP0JEhOJ6
GJKkZk8PRmIwPizTdllOuXLsmavvjt9s/YiNdQhHyva1V0DUE0O3RhEBQJXC
b9b7lIJ/iLkl00UlFh8Vqe2XUDZsfZPon9vj3LRUrofyLWax0oqyIL9DfJf0
lOIqQmdXjhQg77mAFzpco8BZxJOgzfDBZkb6PLmNID+FWKx6feTxxJddDQgm
2x4DlT8WfwVbzCIqwn6OmZlZEOwG5HwBE6qOdvK6oxybSzoRWiloQseAy0IS
16lHyVOwVPlq82PwEhU1L71x8/DUZv6YK3RDVjV0idk7QxrdqKPqyWQghxEh
2XCzdR2deEFSq+SqjriYT5xdI0dQg1u+3loJdoShQbWm1jUHvfpwvskma8Zf
h4TuIO91mdsO8yOK9l8vAIT1VVP/21DKcdoOC+nrq4BkuypjAXkK4kEoNo4H
JsUvpGLQ3UtpmYNafyiSFd8pNycP0JmGe9TyGkTpE0Di5vWa1+PvAsh5iF1b
5vuFPadkI4Q+RxYVsErvyeNgUoYLhCAKJSCAPeZMjjYi/fKm0/X36ITmFbca
qkSRw9XfDKMVRjZR4hpKLg3hdCphf3d7QPHxMVQxrmktN8ul/a3yVod5YNTf
cRAj2pfvhsrzPatK3ygFpmUolxB/JJdsSaLBhQEBbd9K3Cst04N7ezmnaCC8
Ql89BoekZtbc1u2LwB1LV+a/E4pjli3ffeU0eNm0vy4x+a1ot4zwUUQs5eGp
iWAYF8qzBfNn8xrx3IoLsh6svYGwz3Q22imCTYOKqREU2aoCgktOazpUdWVy
g+VJv/MVLO8X7jfPZVj9dU94SqUGymCq2wHmeMvROrTZuq2fC91q1zAw8Grq
JlJzLrDrSUD7NQile5Za9B3Ey9jBF9TmoUKz9cMmKwBk1EPffSAduaclrQtW
DniIEv30LmKSOzkCKxB/ZqpoqgRpvxKTxPTzaNwas3bj42LqZOk9OQsK5fXa
QcJ9SEaFq/PjXZZUz7M+R9bbc7Lpeti1mfxX1laUMxGgsDb84TE0S2Pb6w8Y
YexyPeW4i7jfv2ayggo1T5rCCW7leJ3B1HmkQA522wf8Sna+Lfya72KNjaC8
DvENhCKoNK5pZ+0WVOT7HzXAQH2YxqWITT/2jYkn/f0/QNvAqfziUk3HR2CH
y6+Fue1LgW7fsLHtNvuvsrgj+ay4d4gi0UqA7RuXz0rW5xk98jRZemvS824=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1IrSky6JYXQeW/D4HRlYQ7Rg7mFMeStiWR4rGfyvYgL3cnxf4FJkAw+dvxbu4UuBBY0FtthxCV6x90NjdBNotLzBfxGOmu3M3WwDaH97vFKv858lmtWAW298iGJkajgxHX/zCCjebf3i2btutrOBlaYiYV1P4bJF2zDtUb975v9FyrgS5YLyrU7wvcvenOUyui44TD8Q7SFs2MDQVcGIeQl7Ud5WbRsusSc9djAFECxp8Yn1yR2Swx90D9xY2VUgUBzHfA7CQUT0VzddKhGFNpKSp1w7ep/v0VwLS2hRMUDN8skiB+Vta5HzLusCdXjdubS30rATi8BsJv1xvHWsVwSl+abgqygNEGdHoLRyd+pLxxkoWo2ZwjFqo57SuodK6ea4J3Ha3xdCDmymSVyvax69S26fkNer/hGoMZQmR3gLjIcBuyMCjccwpHoT8qh6KFdeYJH3YhnhQqK8G1v4kQ8EGhg+7CWTSh1oi8r/TYBud2xJ6BBfqbOQKz6/oNAXWD9bgouWR33MTN2HsvPnjofwyFJuO0lX/4sBB8JijGtCR0Gzkeov4JLRx7DQ0RdqDIO8ExegXQKQpAhIWET96h3Si4+rtGJnbY0SnHoRQVaL4bDXINOw8Ab2P4i1fNctMIfTGryk1HPuVvq7L02/OP6A+gq4T3rHOCU1ndfYlvVKHrqpwqRqAzl6Aw0XuB9xCKUPjP87E853Dl+VhbGmn5v6NC/wSI1fQqhL2qf/1DzhvD+QJFTANtrQZB0uQXW4ATelS8Q5XrYvWiAP8YHWkXG"
`endif