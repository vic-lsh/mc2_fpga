// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WId2a33ancvWn1TvIpbD1+SJzVd+GtGlQBko7GDrxaQpiy9+L53842NVmgoF
F3SwXEKvSMSJR2s/NbT8u7B/vh4m/cclwG4QoxAjop7W+VwcaLweQR5U5JLr
vn7qAchqyVRpxSUgxhzrsOL9NxLu6LRS1TAnF+KpYTiO5Iv57og/lv1yDErX
62q2sREqjAEp5I4xL8zf59viiOYElY1rE0RdEIk8HfHrqkmpMhoe2lttpM3u
w7ET4VyN8Zd3KWSS1PXAvXzYRLodA0Eapni8352d/q88w5Nsr6SIFgZtvnAb
hOn2VR2Q2fKgwU6RKrI4om/YxZTL/Md3O0Rz9UoFvw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SzL0qAyVw27mJnoEsWsn6U/RweKGMhsOhGLuCAGJSKBxSLHYQjC5tpGPnKAI
MFwRDWY1DzVVGnxtZHZkn43nQZVByPzgBiILHyQb9/aQ0+21PFF42f371d2v
ZZ02gWw40t86olZtuH8NJH1x+1UEnslz12LRVDpDjSJboui14Zz+KcTHJN3m
Ms/g+BgFhFSFighhgD4R6vv0DpM6eJy9wSuqVLcR5ZeGumomr4fp582GiRNt
D71biSGNuXwi1/fCbw3aQ++D7KYMUakP7nd7BsLdjKaBhlC3s7Ue8NE73WU7
bFMqx5m5ge4G/AclpIHxbqMPkErxyplvhfN4JBwTzA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oL5GF+Bcj4N9cwcmd6ndoy5/1L7OYmFLlmLpfhgaMSv4o+mCqxfsC4fIKrrq
A15aA/H1NXL2Y12c6GPZ79gfqwb663TGLIXDK8dpKnRvlsKl7aE/scMUfK//
pgLtPTGMvHYbzayYjG6EVCEj7eIIJ2H77kjNEypjSnO/iZhpTZ54py3D/vfF
/Xt+ypdVRxUrrXCMlXI3DeuxJlD1NwytO7u//HIxQlqzm1F78/lWHIM138Uk
FViiFyF2R/Yg12rQJbBlHuQjx5YnSl31DfIpXR582DiK/ZRMSCUyE+tucIeo
ADJfrHhTBAkCKm4bjdLoDDcbm9Xui5JLYlXTYZlPUw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qrLxHkP9sN9cN03fH9/6Ex7VOB+ZLhS6/lOvR+1i7DG4kGtihAYyywQFU+Rk
a/yNPmDdI89f5G0tA1Q1NSGV29ibO3LFtV9XAcyo8LXfjSaf2ICjlMGrtgss
6ucQJ7lORJ1/ykr9XoyYE76VKtkhOBENiE0KsuXuK04IFAxh7Ersk+KD6r6b
Q6UbGaZdFFOQmkpnBDirqpk/1vbqsvtCne1HyQsH4HBrxyjAyfreIUnNwGkH
l9osSY2Pfjk9HsV5k6WyK5RrHJ2kZfzzIxy5vxR/HFcciV0O3lRmDNDcCNbh
IYeDInGNV5CVig7zO3Z+ZNRWIKc/NBLZVvf/iYBC3Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FHnAkYG/XJ0qCyQPhx/k+ZE/7ofEBAoYJ1cSbQhG2hwaBpQFlaqNzWxfmQ8v
y7yxBAOKCt10HC/W9dK1G/KMgOiMbEFaRky9uOlFP0R3qSD13DW3lv303CIs
HAVomo/lR1hOPIAUJtGVj+A0oG+WRJV0x4ozJ57M4EB7unojiNg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bfIgeF5LB81iytTFd8c52ujnB7yrxv+HxIjCRv7NzBZix5+3gAYDQ716lLE9
5mxnsv6QZwGzIJW56owL8VOqWA66VaeWocTWIG1I3CBhHk2I/uTIPQzm6SXO
29LINBJH9HO2LrUoejsysHE2BHCAajEu8ojwbyUxROfRCX0l3s2UZU38CY0d
Owbwag4I6M9olJ7lAuOi/32GsBe8xkgto0TZ1OqKFzng1hkRMjFZNG4ZyY7t
OLdtEnHvf9fJzMue0fzsPuVTTuL8q9BgTQGkMy6u4VHmC9bq63Rqy7J9CnXl
t2pu5mg00KW4i/OgYYM9SWJCI3JPc9DWI6z0+66D7FSQO00zUCNtWfLPOBP7
hltgJMVK/tG+jRJIAwA9v03wuk+8/J4TiZG7IZRdankvBTmyEiTRkiwXVMY2
jCQae68QxIKtaWEqz+HbCdJ/fzNDlsfZIF9tZ9acJNFXXvXBpvj80y8VdjtX
GJC6WB9+MepfrxLSaA43SpYwH++UdvKL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RY/K+PwT8N/R67NricI0tW3Mam8oCD7A2YxmQx2Scet0korzkyydu57bOJsc
Dx1Yl9ck2n/TR5KmoSFw6nE0r9iqJ4PcE7yjs4lVDO6B17QYS07a9i5Q4G0P
zOnTnx5IFlGMsP1SUFD6Z9PGV6x2JxUPNz7JaMAbkYkxfcL6cOk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qwsieqLcCyKCly81I7ugKT47W888dhBjgkUa3fnJebOsOle0oLSrrNTjq6DT
t7h4B4otIQAACeyNoqkYyKT9ldU6MiQIIfDEjKCcSdbPqHCLYO8IiO2zkX+d
nMf5YyTamW6oQ4Dom64T2NkVb2v9HkW1d2LC2k45mPjDybT4beo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1120)
`pragma protect data_block
6JE+jjQEfAa23qxyYnoDCDluu21zaCCZ+m1SrzVfQm2zHNGuv08e635h0pNx
q0R585GtSN2GhWJFSadmSv0bQoyiu04Mw9hR9fJUCF5uXdLPGY3p3OsH9m30
DC1c19thrWiRlpeA0NT3HrwnG9unjBpPkM4EdeecE4GLx0CL3523RpbsSruz
8CPfVFNhae9eg4X2DFYDDVrvBAslLdTiTa10F5gy39FsWTXVSHxvoscGJyKd
bE8GFryr0gESCVbq3qE6XNHm59hdWE0hzz7jk3v+utSalcOOmjdmrQpIf4OD
1h8c1WdImDvfvOQNRuGJm8vn/Llgoo8EDJg27Xw8woshwU7HOsJx+1VcIDUZ
Iu1YTNxFVdyTDPYISJT+a3k7d0nVBlLk2vkEVss+zuU3zk1CCz8FsQ1GhWOl
wfD/K3kdk/2cUyGgk2PYpSsECikPP51cSLzMPpktC/ln/9fDTs6g5V0S4KSw
XbyA8j65tuK8jJmhs92aityM8E/yqUkDk++DUSS5/2iV/H6ZQ/ZH09XGkjT3
e5KWl67TL7GK6s9oYdsEE1J+YXty/bJ7jdZmPpbyiAKMbx7wqqjWONoIl2tD
6Ep80maGrxQovJ32Ibxry74e09PqBhJYrMSXRsDPy0wyEi2AIEXUh/u/Q+Jr
mHnwX4SpSsBiEDYAmMMIRPkGrJU+7XKtlHjyVjoixc2a3oiRGexd4IPtxklf
HV0fkjmHbAyKLlQJVNgFZK5rWI4cP6rHHlJ4EMUmelZe7NwWGgAJDfobASWt
b1x0toxZzGGDnaW4hxg37qyIkFaXJkbd7LeNgtmZGCCGDneXgQWE75L15D/M
btIxwKgmxLbCM656Mneub97YN3/eR5LNwgqJ4QAmU6Q1eWN1E3tAclpyVlDe
uzz0+DvvTXpeKp3ZR/lC2qOqBJ/MyaoGVqp4Hxec2R9e+H7lQhqbZwVp3ixj
F/YXpvdjwi0VTDooK9KAOHp98Pr9i4XfcX8mWKLzngus+nT4RIx9Z6hQP+yA
DTHX2K57BONY6J5RyBKf3OXL2PVvnDWKt2OY9jm96fhKGfh4c8oZjeHXIFpS
By0Xtfdn7BWVUEsGKGcV6H++Y6MpJh2f5+DvOKuTAur0jSdOB4nCyg6ji1Z6
Ii/sz0BhBM+ihjCv8mkcboxpFA0u4GnC7W4WrvR68rY/LGWAF3J/E6RDsgbE
Fh8AhB8gtIDdVBfkm0ZyFaaAXRM+RdAD3+iPTJU2Ph7fPL0W87gUIAOwmeBf
3YgwkZonnBy74rQQ9RPii6L8LwWjw8jxSEcGIKN6MJnhYqEETmmd3EiwGdzB
tVeyS1u4UmnNMzOpW962Fwt/8QdqIXo+16VFPe+KNiouICjxdtOXDnSslHct
cUvtQou/Yb/29/a8BEXxRR1v4gUwl9k0YI9TMUyLXT2232B3s5degkQImMul
70K9E85HrdybRBjQA9Ei1icv2yhxOpzFQt4DR0jRMV+1iB/c8xByfw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqeSqktt88i1BcHbeXtnagvlqSXTWidT5Ht5qX8W9udIxU+1YTGYqT1piMtrvC8UxYjSh1D+dlixE2dQltQGOZJlvEOgcyH78Ovr8t9qGRVo1AnUtvR/Eu1kfO8UC/5R5NqIuY4LN8xKI2KANVX/Zy7zbKAZKmSQ/hII+LqyEbriKMvFq/c5YMRbous8WZ3M5StNt/vA8iMqwncAytb6fAu2Ep7IF6GJD/OjdPX2UTC4VbCoVE+6aAYqdQmtp/tlPzd5bxPlVXaQ5Cj8la7502N1EzoGfOeGqbnJxtqd8cn4w8/C9WcZjaJ1R1z/TtK3HvH2W/W0Ob+qxt0MVndErZPM7gFgvdsaQbtQhOiad7uqhZuzLPZNeYp16bw8slLZcBnhHLqmSt/qviEvRVZ09x3fmwEuCWy8bgCrkmwBEUVSWuRtEVeqjMGhbNEV1a9mZalbm+guoPLGtxzxcK1voAL8R7vCnY88lDoKo3u4eJszULWvwfkZC+HzKPREVjGimexXoc7upElw4pYa6KqEvwgXAA9HzO4Nj/i+FB8My2yk29LyVG00xNBgFf6QTxPFjXzIxASeuhO97Ty8qB1UsBiu/Jkk88cPhHp3tLOwwWRs3AaJwBrq6l8yYY5YUvNjfznVFVbZT/O5r8YKfmIkmwABZuEeNXmufeB4rTiFC0hWBIpim+IKjsLJ92AY0lVsy+l/57kBR7h2mnDun1Uunccmrup16O309mZapwLipoK6gqKkwNtNrlBWVNxHwGXugSoT0sQCrLBYV6mlBUnYy4wn"
`endif