// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JcZ18qt3tpL9n/LGMqklk/QDUE3kVZeeWokPzDnsNZ/R4f/jsGyKi1DUgOo1
iPy2lRypVnbe2gvdz3GnAvdDpfysJFQcI6Rpa7qJT7lBtVx2mkXVWjbET2bP
v6tVZnSJI2YkxZpyqe7r6jOMUjH4idpiWtnDkCC3tfDwhEjBGGACMjSeFqAg
d2+m0ex38710l8j0FVITH/3yPkEAGe1jILtt2uC+CvMm0hcs6U4u1DUf34O0
7fpOhBVtZyRnXofw0I3DdT8ktNuUzk2jmb7QDEzuSURh/nFRDElTAbCnLxrm
ioUce5ENtHB0XgRAWgGsrd7T3GyemWf0WbCFK0mfKw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d1b60c6SpzjCGTyL1l3y5ncMOmWAFxgdfFHjyAXf8vBXfq+y7Az11lbLM5WQ
NOPxC4zBBW3FhYOFjy+QXImlT+0kW8JUzAUbdfVvsrFZ4jEbfWtmUc/mDD5Q
CBVIFoonjPrmyQz6yT4KBV+tqrLSzlIU97qdrAWzmI8GyJzT48QRNKsIj+Fq
swFdzX56O6s2XQwm7MkLLhpMosvbeY4+lxfYM1hfMYNh2mE9W2rc0YxMKAco
RnCnvyTqf6MiLyrT/goScXpUpdgtJfEz5TONlRfmdvxKOsJy1DN+PGFUckDq
fFDkVNhtQdFspRBg1VSCCGmgd7PFJocAVG5Ik533CQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qf5X+ng7DNbluHGdpWXhP3s9wrvJnyQgX6dycaKrft+6wZfNweL/sxnA19Vd
xsqpOk6E4A+VpKAFIbhGA22cfJUmWBTQgiVDd5l4tU6Qn9z8MQInY4dDUH/N
2XppsPkAGNsNAF1QUBzta0VjQ7bN6N5TjYOmQRt8m5Oeo3Fq6nSqZf7MPj+0
trNs4BhMU+OLJOEWN/f6HLPuONtrmUPwcSFlt3AfRLvoKEmK0R56Myb566Ue
+OBf2REdLougAKwDIC4y5HTf6WiOeMc+rmRoxWdrd39BDvxKDKaJjX83wx7y
K/v/zOUieZzSCSTbwGV7RTvPDyqfETWqvMe/YO8IoA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KoVkrt/D6KABiOlmxAtmeC7V2s3rcuzlJ0TAenNUR6vKELB7X+evuCQdDL/D
FPPpZDiZrC63g6m81tbwb4YaivEvtCYxhton4ZBbYT5pIG/w+4kTL6caglnP
FcWBoXcjHzZs77YFo2kdeZT3Yw4CsGV1KpKo1otrk4/2XNHUd7En9e2RHEtF
RyPhsBMAf+ZXxWnnQwc7hzbOjdxx2SClkSIKEWEtpoLmTD+BollrffmuxQmg
3Psnhsn7Y9+Q64lsmRq7B9xIaPKALkbiQJ7bTyE5oZEB810kkWSJvuACAubV
tavRPTEEWPaxeKlRT16RFo30F9BAT6dy/mmdJ/oC2w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CJiha1eorpzQtG3YyMdK4rny6rnP0jyGR5LuqxAeJ/TfQSD9wlh8ZlQ9Oryt
5xcYCH9A2Sf+Pl6QnS66VDxjyJVemQsz9JCFe5mK7O1kzVCDNuLt+P2AkPx/
4+3isOJwv/qkdxKepMPb+BY+YtVvOOP2KEih8FZrSDP+q1AOnY4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ijVmhCNXLdhAPqfv0UgTHH4ZeSc5E0HzbZHwHmSLAioGPBZ5Zy4XxMQZQb+Y
M8m9YSAqsLFQC4NRiRBdPnsnGCD6Ubrytp6DeN+C7Pva9HM5utfGVn8lDeTo
l1Dh16+XRWgi9nBTDpMORHVM5yBz2ReHE4IGwB2ULlbmwBQnb87S0uVRQl3I
5D0CBpf26lclupngNiGsXXioTiLsRuVJGJQ2KKUZwa3jK7t+dfSu1A9dhsuD
XcBVCUexMNBc0YU5KnfAiXliddi2O1ltFCsGuSnN1gSByvRL8zPZC+uW6ax8
x+YAvHK+hOZnAMs9q22SM8erZn81755wbNvSgX6dz1unkIAD2xy7qWNHWLGK
c8sRSzP9Yp7UbXhyId4WESmVB4y3m4Q0xzhbLuqKPYshsaH9CDBgWVJAkbf9
KWlskRrvBq6G2s3I/dQVgebwtGZqCxjzaw5WWFSr+SNIZXXVuHDzQVynA/s2
TqKukFWKG+NJ0FngU2/XgEePRKc7vH8D


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
i2e3710QklSJoJFpI4y6kea11i7PowlPR/Yi82vQKae3sxtibOfrdgP1bxOP
wmfxKAvyDwVxhxZl1Ey9JlkjkOfX5wk+8+692riKklMGwCYCM19tyx1u6U46
vkfnKS4ZKOOPAJCFTMrU7TcgXK7JQ05lzYWWIQoXmLERbGJOUDs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qSVkJslRH8QMcqz8AiHb7fGAS0niQtjWjmIk0VjSJA2DEOU2XYxMQfEqJmmT
PyZvKpyPvwj16//9Sjh0yxB4QOJmWWk8nvYQ8lOCKjiqB1vrMERMMeYKcdVr
FJCTfe5foHDDGIPFViCZduXpsE4+7v0WulwsJLQx7Aw0FDuQcoQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8272)
`pragma protect data_block
LMGI8XLKSe+y38CFN3p33G7z2I3A2WTWP2jr80v80v9mXr1GBNReX7kJnroy
9v0/JDTO1LqIH8OzRXwVCOw3UTb0L02MNYKs471KxZS0nGf+dblfImMjEBFE
Nq8Q+75vd7411xCnlJu59/qWEbljQfS+Dw6hSZjl8ciyO5duia5GkouwRV7+
PpkMOFG3T/abTsl1nBdcv+Z7p2/dV9S1mhGQ/SBOKVUlZsiJnhSq7+2gI3+o
ouFYQX8TFTf1/QhzFqszvm1WhjLHHGCGG3ElCG4GeuFsjAr6LUrjaLPMSD/y
t2lfP1y6rN5w9rujoy1mbn3p71T7XmDE6IXMXsze5sA0yBnUIPieHYIt0HEV
CHJgRxRE7RWoCkmWHbfiLACeZcyWwzCnt8AD9kQmABH6Z5L5OMBzMcLkBlcy
BFECNxAjaoIMvb2I5tTnlVe/8TqtN1WC7eCrUSQuo22brPtrrURgEz+r8IU0
FXsbS/y1n6m6Bu8z1VRSvDPUlfs7J0rT6qDmYvYWS2WRVBS98mqTHivLDY3Q
b3IvjTQIbBxB0enUBz3hEF9icQzbzEIjvky7pWnemPBOCdiMVirEgEjmxiyC
rCnnN+LDZHk3UXiibYq+o2BEPV0q3dL60pFSGvHCrhKcy4OgAV8f88dNGzKw
8gsPefNdEneYJCrbkw3nC/7b05BO0XjDFFTTuG1J7FC3jLQZLJcQE92wQzLK
rLNkMw0y7iGRyEl/ZtHH7ApPVfnN8AFysuIVc5bJBvRP3L/78InK+1yofSLO
A4D2AB/gJr/iLsm7F/Nvc1CtDVir9DgjI9IWd2LvJ++ooMWp0dgKMHtiMemK
0nQMorpuVB6RTCk2QEnFfzgYzt6urfZAMTjj0y3hwdBnF0jQWs36xMExjwcn
287lS19GzSPNgK6EThXCyHgBspSK8BRiKiBYhZIfQ0q4rQAeP3xuA6OqH4ZV
PkS8QJdXNT6C4mzTaz5sbabCSMqwt09d6ODG71IW48GJywVwWAkqqpiFXc0U
IJnlxJnnUJFv1TNLwysv8YR8A1/bqo8M/aWphRZybTS3oAJqQ4w28VQZXfjB
yW6S960Deex1ybdqcVSsw0tBkfOzu4pZ6n2G69FPhwEcEixsOX4efTYLZTdP
/J0hEJZ338vTEsAE2T8e8s9dh/2eQm/a5zK7Xe7zgX2O5ZAQ5GX/Rg9Obnr3
jcZE+Sb/HuTIbGeJv9veGVfxPSZf5D+/NUgU0DIHIAqIrmQIirBebq7ixOG7
XEuu3ZByP3DJg/LxDOVwvsP05+mS/JAnG/NO9lAtOoHafJMzy/WSPdJiO7Oo
onYaLBN1LRv2ef5I2TZPBajH0UUu3dgLHDTV3AdqU2ZSojgOdNBFvlq89NOl
aAoSpk8z+veLJHi4GO9t/AcTgOvLEKjbCrrnbumyqK1/70bSn0VU/8fgWGdk
V09PChzZB95SphtFg4r8z3SNGxNNQrTdeTNZagzrD60xB/DGzCb1i8P6E/eZ
uazTd4GdS556dVHnWOpuxQyNA3DwtqA75SJt0L7byDABwtq/aDksAWFoOFxw
lS4+ekp7V7uzOqyHKDl7VXK0Q1rx8in7ZIX+Yf+tGhVifoeFL5Dg/BCsyls1
UNOaPFFuQKUov1GjbQLIhsIy/KL27zWr1+BHXEw1M1IMUWtBuoQM0SaNZ5cj
SPgyASveOTTNf3Lv46Imm11mmiDeSC6NS+lfC8E2cX3uLFOggZmfKNdSbhaM
4cGZOXp363Y3WA2O2uEPQH5ZHYe3puotsyGRbc1IsfSTJRiHa8E+pElPnqgY
Y86yGuYSeN/RwWdvocNRHoltCxPSJqFTJNKXOxkRbHmh6TnLJ6ZJ5G3qlew5
wSYRgL6d2Hcs6fEiTe+sNsQlDQZwWdOd2wfrr7m+ZH6NTAjXRLAdOMyfo2p4
rux7v5AplN44AvV37+FTDbLn30Eois1D1vpbi3uAF2hyvGs1C7Y9MRgdlm47
cT495/bFCDn5T2IiiUUhEIMtnU+SXoeAq9P1aEtPNeCujGBvsOQ9psHGSw7i
nnAWfMMcGNLXr3+Z1kir34jvJ/gB9U+aWL2JsKIh+7rbCwKAMcqUwXupSP+w
jxJMDnKx1kvbtXYTGLuBKRYBSJubDA75sNqO0ZN6MQj2w6gBMmwmuyiV0Rhz
aqSc/2sAIXOzx91UoaXyc/hvrWvbb2S591KqxorENf9Hm+J1AfQ+ofr5K36K
jzD5nehVNmO4Tu0ZFQo0DxZFn1cp4IhYNc4wuOzRLCyyXuRpOXR17mwoXV7z
At2OOp5Rd103s5lnE/82cxCafGEfp/oBdknjMsp7adfgW7qi6NYI7/nUurpe
71OSX9m2TByq1tgdi53qH1HXraMW5C5ipCvZgbMPEsOFGzMVTeBp+4RSMDK2
WxGvffKdaLHEajnlvTUcK9ucQZNXzudwdme/CaZDXZaHXDVvfnBOrzkoFQlH
Uqefgtzlb72Pt8lVGOdtLvp8ySjdFwtgYCDqF+6S7r9H4QqvgHQ7KZC8qYxd
scqa2KcYuSddZ6qUfYOUMAGoSYObwOVWQsfFNefm6WP7S24oYbmSbLYtHXE8
cp8mDhUV/JiTLJV4x4NJb9CS8iFVUuxbiowLKm3sHx100LWn7x3dgLax0BJq
Nbj1a4iLztugSlTZXMB3cSmO7TPXgEOVr6p+HC96tPuNWQCn6jU0HF37ytVu
/AZtCCEV1WMt0xes7/0RuSILxX203BJsgCqQVYSFjpPC87SAlzj0swdtXbFQ
RxcrY5ZvM8wLYYV0TNf6yTRtTfw0FUsALM7sApcbr0KwlOSds7PXjQAzSN19
xen/l1vaViwmDmYPZ+6i7CRCxGc90+jVsUwA9RgvACqXZuhqjgalBHY3nao+
IC8pYzFiVE6PHnUrJk8msQRVKaZLz1xWuY5FDRIkhGPkKuuCeWQDtnNoaYfF
lNNR7TT95LXw5irtZFzbDIXI9CRl5lsJEQzPOVNDGmJxW1bX5u48gZzN4HJm
ikvdweI4iyIw1sykf6QkPzwiEygkR31Z6Dnoijw+Qpuk5xSPdzQG+UwNKyEo
+9jqmBJOGEZNNhJl5L+7dXiZkEx56yV1o6NZhphb/y5MtLJwfMoDXSndUvDZ
aEMK29R4WdKuuF9UGJtqSDPwQGxUeVbHaSe7yQa+SD8oaQDnpC1RNYWrqhTB
GKzeaRSyPRTo61HppqjevIFi2o+AR5ebJisOgG8NXnvDd7v7n9VGI6PQ7nj6
MbHh9i6AltKA4r28aEYtbXDhqnGl4hv4VAafwo8dyK0gtf1gVJxVjgmStgJp
sTcgGyeRnF72xQFUiM9v6UWhF8Fjh55a9Ll2krUYSoutuBSYWScYj2i+Maxp
/oATAG3Whbkt5grdmrB4Yx+y1VJ9wAB5rV+FcdP9UCi9XFBx0GrtGqhqLWGR
xUbQiJ6t29PDpmHGPVt+iBfQaBRsEW3ceLpco8AvxQ71B6JgIJba6G6NEdDd
SSBqrQfyVePlzJpPqCVAjbYWcYNupSaEZsEUiqkqf8B+5AA9i7d6Ok/yYS+A
GJIlgrGg/NqcaBqd00TbLaPsT5Ybv8oOZUTIzu23iPlVaEHQrE0AQ7gBu6CE
EWIotYkMHvq+QwO6TMffTMdEmp1+36JD80ad4+gu7Bj/QYPZt8fXCrIQjcJh
OSp9HWAOVD2mL06VzFYWt5vxrzotVEWX7Kz1/n7aM8tkrVK0SSwe9qyzhpZf
Tifkk40qZ7bWbPbcePytaK1F7YS5HZAUiVosm5D7OxE/XNCzoC6s7Vkn74Vk
jP+mnDcMCYcGDn8NeJYeqJdhikF9NiA4LBJs9/ZqV9eEewLiKLXk0mXAkz8k
9z7gxL3DXMaAxLKvIuW8KsOikxGHpZfdr6zUC+Xdy3HfgR1458uxqqqZHY2N
wgA3gSKuqPMSyuLdVWQz6hqaoIwLfGY62vUgdtwRcKIa30RvDTLj6roew17H
6N5ISZqp995UagM9wt8A0HydQ/caCW1IySVCsyA14/RQp1yhXdIk7GUO+IxQ
gSpJEQDUjLhv9/ZG57whTUKiSWqyZ2Afk8e5+eGkUNhU+IfF1LtXbuLAccVd
McepoUcZqqc6N1kNClHELBM2KAzwR+DpPgjM2UeXltUiGzr3+nqNxqOr9oLK
y38bim27BfSlazCgGhWKf13+86FzKubNewLJn/dm6tRGJkg/priM/hYDBRKC
cow/R6QinYG8d/3FmjYOZsAtuS8emElK+Ait2IXtal0FX7VxNdGJVXz2rE0W
wc7fY6xfQjb266X9IXS+kLFikZQaRkbsz0mxLLK7TGqhtwaFM8ExVJQ9rwW3
blRMqpm8h2SiWJpkDJeEcKDu68tOgiZx2gYAfEa6+5erZj4owD2MLHVR2HzW
WKYwCKMOe4MpYRcqi1VWsRY63W+lFnpWOEIZTRlNjgzDhmt/XQaozbEuXgbo
NIPSW9RsBH6HgXlCcWxjMxdePDqJByjHSAVWzx6kaL8O5ZXxrolsT0/tTnRg
f+y2EmHWhH3qV0hmDTu/crqlvMMEsP8M+UkXpAc2pKCLk1AENowYN6Ax/DF1
emivDE2Yt9+ulUea5iNS/a0Llrtjl8geLKzFDMylm/NaHRKazhm7DQj/qfN2
BOc/KK8K8jXWfUwAWtzxmRMcZxxTle5TgHuyn4SmOR4LTjP5hxcr76Xd82Wt
AtR4XIVsSl9njjuQSCgJZAY6YpYNMfCiE5MVldmOrvU8Nwj43/G7VO1MsHEf
Q4J81ITOmXIry7qwG3k7/90wPG39D5m33vSbV+rDqqrtIcJte4ixOL7KL/m9
xV+J233mQ7w1NCGyutpQ/8qpdn2bs7jRGe5Y4UqGvL/Tpd8fkHqt6LQDaA1x
qzJ1YQRm78mAs8SWHKE+CSz3nejdRk0GFRwEmARUj7+yn6/5QHv/3oFZDMWz
ghh+UGizyVcs3O0Ang4n1eJsY3g9upFfN89bOQNoX/GBGUzTqM2WUARak4bi
2373iKqVbKWbmv7+jICQBJ+v7CVwWwab6817+YWz3NNLoOUyMd+kVrYvykLb
kuYmUWb1BDbZiVeuIRD0sMl9kqCiiIuBJOmvgD0QXlxepir6uQV3RnaEKZ+H
seaB4p3HEDrP6ec3x///Wk9SxZjmgKh7OQyiGSTM8U2igw2sbLiYJuMF1MsU
wTQcKIilFztEmQ1x4wBg1QnJ3GFF0ER3aAn49/8JDXNk5BuLk7ZZ1k86SQBI
xRUG6TkS62gM+QIc8yqtmwlixAr/UtW4i6upN3jofEiF2+mHfbEoAti4FYof
34jIKD6hPI6GMJBaJZKhq08Rbvk3JaNrfN9Sye4B3wytepl/qGRYcfyBm2L3
6h0FGIf5Aqc4ZcFlcylJ6Rgqg3DDE8Az1AklCTS5ENDBJHVE59YlJDAP/NHd
weVijTmBSc1EE5C3bpzlPIBoBmfWYMiuUtDmF+fa+N3VNDxtUsnBNVUn9QD8
8XiXucePeknBchB1cIx4GRz61koYFwgeuLPCiSKR+7WMUgEfJ4mHW9b/gkki
YO4h3E8YnO3dFTxngEp1sUVpa1tAbbcXahk4c505OgfL98Ddpuj8svSvS4u7
IrW0jVTBLz8TFpeGVqc+eXOCTQQl0EIDXRoQ/APlIHfTso668JX6T0t9RTus
LK81+ZtGVDDGjFLiU3PJh7g3VfjszSQ1rVC/czkRheuTeHa6BDLe9vWp3FnC
UnPgveAAKtIih3zs1h7zzRuR4uSEy3+AfFe43qaEhaeunQ6n8pnx109/qfA6
Pqub3VNrPiRndfu5V4Qnn5u+VgsfsvR8lddnN9ojKH+PhnAJxCnw698M8dtV
HQ+OpsIkxtdfurO1p1BdfO2fixAmGJ8Z98ma9gs8SQqROJBFN5yYAVTiQWVy
Z/6oTrxLJHnGjtn/rBvLzm1jk1HpT5zbtxA7mFowzxr3UXt8bvhHiNwOLvVH
RWySmUdnzApoB/GleFt2FY5s413BrOtGZLr/W9ZCkBSLLVHO1cFYYzwjtglW
1Md4eg4ScnXPI4XWEO29m1J13w70PbzZnYlEwWsjxiaysycATHjSJllV4CX+
4IXu9IkGxn5XaxBQXo/qHI0I62tU2iv/TPfu5wVvd4otwFsdvJvYxdaOoXSF
PiJvHMSZ9qYdbBBPO3ZwTcINVv3uuZN6nF0fEieLmvQ5FEMMGynSofZWumcu
/ieVnNuEv64EJ/fh6HVMwmh1IbGVNc3DEPTEZ1LHglTzGggtQemskwrDaXCk
8m+8ZsBAUH7iVoSk/L2VqHFiBxkaCeYLyMM5KNbjAT2utC02W5ykPcxJ28MI
f8BycTXJClCM5tSqwE0j+oddws81ucgqjQsre1iesuonAExItS+WBKksQWRr
h01fs4KbonOyCPlUpg41opdsq+XiFJaKWB5g3PTafKHeAXUoYINqQwms1Mem
u3VX8WtPbvHah4dKueHipuOHkX8cK3QBioUnNFG0UolLa8i7ulc7dH0xDELf
cG3xYJBhFDH/Qs0llsB4O9eAH5jZTVqG1dWmlh48r8yFIQYMwB1YcnBMHDOF
qe89BJZ+00pquI0l6Lunyy9cyEgC9pU9jO9v32kWi7iwn/JgBrvRvSdsP9cH
9aWisACQOJaqW2lj5N0310gpI8QxF0oAKnv+rloAPKm7hfPqvd49RHWHEfEm
dM0QL6ua4h6sNS+JIcTqvNg2MCyP7rNMVBbwojeqQ04nAhLOEhX1JA+c7u0X
V4rcYBNyHNeLIHNG2uahz3c+f4BqRrUp7KuUzb8bDDE6OF27vYpCZSXCQu3k
BX5E6+9EKppNClrpv+bq7A7s3DuQyhbA9V7oy6CuPG6sNE2F06daOPO4A31z
PTQjQswPrUyFaP2DxNXspXe0sHWOL/dZAZp8oPffp33EunNd1OxAA6ufObNe
0tvLtx+wYi6lxIihEYCWV3dPRAscukZ2/qU+wjgeo2m815lmgkfQBRvrusZd
s1pQiFnVQoy43thzG9JHcehsgWjCWwxKYIuxpW7e27OEs9TZ5KAZQXyOPSRJ
eaGQLVqgmADQBhvGhL1FN8vT2b1L4DzZquSivnWKhx5CgR7us0zl0LyjwoES
ZMoiwy3q2Anprt4rlkrEZgs8QIa/+jGOWv4ixJ00iqLEKQxWnBwtcinETb73
342o8fhep76I2BgJswNjeWv3vkQkz28o8mlK5hKGo1ICd1Dn9DhrXnRnSNt+
bwQTDY/uXNWsBczYmSp1Bf+wszWa5eFmv8EvcN+IvBndIweVr/Ti4ngoiLJK
Z5uWoOoTFZkGBdEtVzSiPecgch8BSO0uHxX0s7wGznCkc+BGmh562T9t6qSP
CJ0l++V6eEX8Nhqahfa59pck22rnQLZpQJvMjE/rFZYpribC86kB/Zhy+4GJ
Ca1tvcfR7cSTVBK/77klNx8Vc+GDDMJsXcDzDfc0SGOSEg4xDH8G+DYMCcCc
rT77MquWHL2T4TKBSUpkoKEujOS32QXG6yaylk3tMr03ofgJjiy2v2tnXLYr
gl735rmATq7F6oTAcJZ/o/ENsglM9tLIRCCxu5ndKJOuMtpSQuL89NvKa4L6
Hnat9Iq1rEAwIieJz7qJsV28nE4q3ONzfGVNRj+exZ4PITrk97p3RGg9vo2i
VzVpdmH+EtBdl3D7ZTg48ar5xCz+ebPoF4cm3fLmQWmAkmlVZJtd7/CmXFpi
oBshLnCKu0yRhjT1lH8JXv4W4fb//PhdgoUZyvWO6uHzMiF31HR2R+9/aNow
ijml0FSq0N1YQBergavRuhxEZ+tZu/8aqVUvl0zOV/ftOTPdac5z6HXZt0f4
haCV4JYhjoLLYhywcUVWuflZhpw9eSuIwf95EigfqdApzQUDwxBKyKqP8/HZ
fOB2Fqxa66aNmb2WXoZckHvrKtR51KxBEupvONUaa4w2EbiNrdXg0djP1VKF
pn96lWE0eje/+ISUgLT1+t5zhxlBCMh52HZDKEqc2QvYL6+FOWZGPKorUA0t
66wgd9wfxgztdzHa3AsyguUgyNWiIQ1Lm2iK8L+DL1CfhYGnDDQ5pyWrC7Ui
L4d8yVI7Pdk6LxvTjUcv7lZIRy4bjr5Uk6GvgH49lgXYnLq3HgOQWh8QQCrZ
van9YTNJcCTeqV/npScEFc/7ilg2P/cXo3EHTxspDuceEFWYCc4ohSY5ehWN
5sC1H/OlW67QF0MIzKvRQuGZ7UehVuISyXZtOTtTe5IQDVcRLE7qAkdDHfge
CNGTq+xeqOjbEmFEebL/qL94XFfFPpUYHTwjsTBflv/22Hf+0/wSFlG9GNzX
8mdqn0O3WltdmuNRPZSbwx/F4I4urs/skNziCQnmAu7Y+5i45VIrEowG0eRb
Up4cVs+x4hQb+PEQKPgIiJEH9LsFf0aGQVKCsWcQVQ/cEWucsPgxUVxdYD81
6sxSD5ECPJoqNAj0BMxQb4JXrew0ewMbqwa9rhUwiV+cF1wBeh/M0OuVzEwY
DLhNlFVR6E8OzFCCnx8cxGqEEVzYJ2a8aBT7+9DekCe5qeibvobTpuOW/m3A
0ZLb/oCv4nUkNDSvT5TFw8ASe2aiOJELEiui+6J+wd2lOMR0j7dpTTB7zLoQ
nNLDbG2d2epwgjR8Ce2C0TdaVzJTSDPiSQ0W1SS4J3GNy8G53/ljqNsCR8Z+
stPk/DAUOKx4/Lf/w2isfDCOSMr+Twu96heis4W1lK7W1dN6fhjQJCTJTvoA
cZFySk5OEFkV29cPdxFV2GZPGbfjjG/hL6+eb/psmLOReBFnW0h4bfqvW+g1
4Recrcfyu79mLFbUPJ1i4SeALlQAyn2GDxLRGGTpWWoMnJG6skTGs+sq4wbB
d/3wzuf7QaFcX0ePRgTvMLkSkGW1Mr/X9YxaNK76hvWbVssf6MNvHSqk8UWQ
/mwGQVe8obUwqMyPMClMx1ifwH2O9URfzRgbrVFyIEsmH5w0qYwYDq/mDJRH
JKQP8k/LL+q0nWDsqIv+fvYCi8QPFmXvTsrkMuYW+tIVwHa8MaLf/tXkFBJ0
wi4AWUaDyiSJtFlMAi+rch+iMjlahKJLmj06YK3HOSWdg80IE2vth5NNrrIh
yC7cvETjbX2wmDjgPs/AF120v3YIzI7IwgDbAi6j1NsTH1ATpvGzWjmOjN5B
nJmlkGhDfadZRKpUMS8lFz3dQq7yDc58k3F5tfn8lhDqDn1oPGXCXKT4fjY1
5DZJvXsf28CDreGI+V9y2OkMfKPWppyEcJn99xNJu+VlynneXgeGVbvv+mok
IS/57y7haGva2mQLRG2OqerwqwKLLPj8nFOmEnH1zzP37yvs8C8U8xbp0RvW
71gpzIy2G3ZiF2oqCUhr7nY6QTFWqp2bdQ15H7KK0zqqzec2ezz00v9j4b6S
F1XFnoEBwNyMU5vy7QXRDK0SB0zdkfyR798m8gHHOMydIcnu31/NoLUQGaPh
lkwXc+z57aRhmkkzbqpdtCI9Tm+s+t6B1+v22dgy2OZBUjWcwMIlcn++EwqA
n5UN1iMWXOiPB36ock9XmFt2xkhcTr9H7d/gSocHRw5ZYg/HQruFmRVxEOCx
tUCD4bSbq8bTSgksTJO4oCVXfxvYJspzXRqgo206bWdbP0LFgTt2+HaV4VaA
BpITXv46FfFpEVSQ95p4N97xIxLG5Awhp5IZXqrZBORVKmLAFHNZVC3n62he
0vgD2nuHZ/lBpErcC+RlJI8hoap9MZ3egHRusqp3p5Lyq/P2iAggu45Zoaq4
eiD31zfGxylgo/tBfamZTZc78qPQKsxGzKTRWSv0ZdUCP5IU3wXS8qc3foVw
s6ITVYjjOGQKUVmG0jf0NNpA5f3p3fpDgHeyJh/asIgrPdmRYe+RwfcxPEiL
HzOvQpkJZ+bXwzCHSRP4unF36opvvTJkZx4a0gDr6K1CYUJWcTJci0jNwcIR
kWyeYo9Kob4vPehf7VlcNFgOs1Nwe77P6nZQ2ciS7p5g3EHYAs7NcC7MZCGM
rAfCI6O0YXKhd2q6AHLdKvevNkw2IlbOGp6u5p5HjfEwLxjPa4NNixlMatnQ
4PcZvOeT8RXHydlN8iNYFnM/xkJpk1y9tokCCGeHYKWT44tSeQeIYtY/b3dD
dAg7qSkfbE+4EAbUUiuKKZdMrq/oqPHfV/WD6bZu8g5CoTvbhDV7TEQct11X
h98jafFkjK+SKxHjwQBQyrbyIkLOkrPup4p3J+MeLV14K7WolJMjHy9fU+3d
rOniarrx+/VfixsnQ+0JbQNu3g8Kw6zH4MuIUtxE78D91GqBstzpE4U7sumB
znFBk5PeTqVD7s4IhSTxQCPQMYE9zR0oe0Au/7qytcKnyDA7IVK05Os64efF
eW41sEQ6yqQUpuwg75ZltH15O9IpvnMWp5te7NSddILyxSUfc2N/w5j156tP
GbINddKVy9Tzxe64NphnNPpeea/0mleGk8YafZHHKz+HSl2ncaxYHsGG51+e
JMe1TW88iuUvn1SZ1NpZONZ07sO8QXaxZ2in7IfdE1v9A2Ln6xbByAkEV7y1
RH9avbaUKMzz9CGkchgnEagLDVyEI9uSR2OAx39c82QlYErTLj2E5umEij9+
Icz9tqeyu8JiB0yoCMx2QKm70ZN8ysq6EW4aGb61ijSVVAXqxf/fJirLTSNX
A0SMiKFzgnkAXl8Bd6C2pg/ssE5qBrmT4fmNhGQlq712u+OLXTLCyMASXouD
7WslNzmFhwBNvO71TigyT/kw9Cq4EdVpm7h85lQ3fh67154+hBV0JKQUFWq4
AEAbtHG+w8Nolk18OIaHb29YakBnlzFbyDLcRAhDTvWAyklLHNdGpSpAG86n
YlcJVwJdpyGhE0O+M0HgK8tRUxhAfircykRFQZlMnjfqZeL64QDK0Kk8Sy7L
Eh9/nBN3V30BN2HcJH75PJ7LFcS82EMBTb9VBr/Y4p2XzvPLItFOH76CNcA6
zGvsBGlkSLrigMwoIIG7Cf91uAc1wAxL/w07K1BSfNMqNa9ec/LW9jovVztx
URYUxDaHyjWER7BxJWUcnPwybX7yZSpvXDdCD5i2/ToSiBxxBg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1Iqn4+RM3fGjIY+q0iEqGsuYK1obfXr0pqtA8qH0n/WXC83N/kHT1gxOAFDo8VKNTZSx8KT04JbtWPNKLQaK/pnER/qmje5Vv0vHqV5o9JU0RnJJdkcB6yKKfQW2BxUNxvBunMl5MNUv74v0Ct1gfPcI1xJIibCrwmvm8uH7aO8cErW3QcULom5oWSkT+waW+tRuZPqMwi0w3lCmWUWFXrSgdyeC/ugxZicWRBdnEyDo3XkAsS09JAm4w6YMzKjseZSwXaxMw0Y9bVTSPISIge61muYcS0YzvfirxrLtrTPOfaaUh9JwW2D7TNMtnWFlWS4Vh+75UcW1pR0jQbFWrrDo2EX7Eon4ljxMlBfwqBRFxxN1E/gO2hEpg/LGQnhnCIk84ykL6rhdsuHIUwflMhekkornXFCrdQ7CS4zWE099Xf2HbjpxWEq1UFSdO0wEkgPAM8DxrDyp5CO+9tIPt0to38X5ENxmywtEbT4C+xko8k7NPrlBx5udg2CBKEJEmh5uAAzng58quyDQ7xhnytKvVwtv9A+3xl9B+2YO3Tw0lhlwKtFPVVjt+c1sI2Pe4JtjFy1P377n6t/Kta7Qrpr9LL3NnoDGPaog7kwifDbjbuoafnmt9PIcAuD51rqiDdvTfWihaZ1r1KfCCSv6f2EOi1V3pUjR8WVYAyT73bcpvjO76kv5VcuNsOxXyNct+WlEdOJw0E9par84bZDrV//Uloovnp14uUrTSsMfvG1MchP6D9ILf23Wc0wJFQu0I9s3HNIKc8+G/cAuzkm3g52"
`endif