// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Gd8zoR5sOtva1Iqvq1r7ajqXKONeu5MC+O3L8FpbTKNDeDsdlAa1PXoXDfc8
kO1PXzErV+Us8LRV/LSuxspnKKHkWUJsigMFYUkyYDKiVM+ow6+lJo+Y5YIC
2UU5yBLhKSY69mo7bvKxtfEa3NkZXgZOhKPzJWXqE01VCsxf2jMwnxIULzUH
b+4qQqtew/JYF/01rH4cSOIGrgKkP9GFXLVg4vA0ZZctmUXxjVUWWD3YYKA5
AhsaoQ7Crl4bROEHw7hvA3CbYzLXrAUpaAvfOUca+rWzO6CwFsD9pVpPotae
ClfD7E30nsa8eUYDmo+jwZoc29QGeHTjZFR6pVy7fQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
F0gDN6uYRSCAUszxgXyDoRzWgv6gvLhzEblVb1C+aQyK4l+RAP5KEsXmSjUB
Z+YrvS70eWoucPHJcO0igZ40XMuoa/JELRi6Bb18ihUm2SE/ltVPnlkSYXqe
QvFqhBczRHvz50VYK4QMt4TtGcv9rECSsyxqO1DsnshSniy8AuOX+hnAJVf2
wzGY/jTZsRiozsPMvIvl7VpflucGyaevR1KGRccoN8As7aDXhhavbHMNsqs3
2HKTi4eI/fYwEyLnFLppdCXpXb22aOGsb+1FeDmAO7ZR9abuwtCAJEJ1zTAp
u4JiLoTPKz+JaM4eqvPbdEv+4eUkXmqjbr8y79SAHw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ALyDVvkq51dJJT/yP5EsjYdKjKd9+r3yLOSXPUk6ew7Zm9F3I+aaQHkkLqBb
eQWEYDHdtIwsAq566W0TFOzqj9CcfC1On6GPtMZNMD3yqkCg89zJN+LA7mkH
L7uC0oTwq0v5hd2cdNaQMwaBBXNYcZJ/ni75lKleeTvSPqInhijDCuEt9/0Q
yDu5NQ4SFfKtXbcJI+XjpBqpXG1GVrRKkO8LeO4lLGO79k9msoMYboSVwW2X
syWn+FLp2ocrtGBBTr92Vtbm9USF+FTiDuGzsvqnu6oi2Li/XkQ05IjaFRrJ
NvhDcnMAeaBXxqUBXFHSu1fAT0hcXVyQS5NGEXFnhg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AiG+xpTtO02Wuj0jFFYwxLx91cNlxPkqX020qQk+VFTB+iFbGFaEfrjrKDke
AbolywfJl8LKImscTGUQJwim15Hn5yA2TBBb/L5C0UbCu7NwC1/Y9MZpkY2o
CHmd8NX/5c0wHpgaO/Qsl7Ve+JfmeX/zCycKNZQZgzl+y5gUSUaHIdhVaCJd
xrm8/VUFYK6jGYQTSkNIhBXczcEg2EfhUIkjlSYQz1IHtZGAnm6GFoIeOBdQ
G3yQcXSLNFK+2pSWCsamZQRj/DAJ+yl30y3Rde+bacuLrGx/AyPZLjHLL+tF
Rc6Eh3iDA90/cisxJTz2h5L3hEN9KJgVJuD6DOWuLA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
f231+VBMyqp8rZbpZws4ZMcqY4E8obaGXa2e0nUMY8RImp97JWSHjaJ2pd+t
bRzMNWwqVw/jgIOkpx3xUoqeF5+EUrVVbXkO4+ZBlYPErjs+Bf/nRix3KyBT
vHqfSwkHlXN+TgcBRqPz8weK+KrEHNa+w/aFBQCb/+nKWDrzOUg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JPx9nYt1/iOWiY9G8NUQqqmhn0j1i/cYCNmZnRnwegIOWJelR7oum0d6lI8p
th1MT0fsni3oT+p0FPiTQCZOfY/ecd4XLVvH221CprQhHhsdUaiFOhKVqwJd
nh4ob1LqPZT1jRbwGmIYTYjQXHsaWstdYttbZoS0dD6GmGN2YIQJkHj9f3NI
8zvwhjtj/ZhukZifSNYAC3EKqEKyFwI0QnHjdCih33ACRFSXIr8Nh3xuAiTX
Ifuelx8gPtQ48mb4wOmCa5LD7rxLp8yDyz9+YrjXtk022SU3Zm3WAAiu7nUu
X8dNifyqZsVt7IHFHELoO0vPbh4HDBsJ4mzfoOH+sE8B7jtcUrNrsDNjNicy
mNHE7jrd3i/XJxs50BJponah5fCPb9okfegtGt7JDF+svOM+gs9GFOh75Q5E
ALv4BjVxnbRP9Vc1hLEbpCqNzs/JQ5EVy4gahTf0KsbCKeeRPlLprn6ujI/b
ZkXFUuM0YuVy+3oLN8xUewTz0eqYplr5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
T0S346x13keo9nyPAyTXt2vzVl958v0DB/lJCoIfAzhYibHptYYWb76e8Ocz
huGlcKwEEZltopbzjqV9X3B32jaYS9T0khbS6NsOEoTkoF1excNV+isfjxUe
kR2o8xgk3ZiR2vdeI5oJdo4+wWQTlHMBvzS1b93TB0qs6DZN3to=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FVdagijbfG8JCeLbxJu/0Is+t+M6ZD8TMClMItQA2gYxVr81/VLmJfxFFAWT
Okg9m0Eq6/swxkkSfDgPPgDwIiF4tXFREjJq+yajZ9uI0s2Nz2X7VQyyJCw8
KK25NfVakQE+MYz4IefsoFUy77Bf3zTa7xEMcII3wFHZJ01u8w4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14752)
`pragma protect data_block
oDqK34Kx4w4gMcwrQL1oE49WQiUYyhM7mTvyoWuJqRPVx42NX1Aszqzo8hbO
/2jw0SxzEL/e2lKzXMvn5WOCIf32lYaBsWUpU6lWO3C8pmfFo9LBXGCJFpEP
ux2Q5jAKWEWAEI6svPcy0uwLErmIZQUxpXszPhZMicnNUs7VvzAjOXPKTsAe
lmdLFXhtOy/p53fxxELcqK6LVgTa68kTPAVYsUniqGtpkyDPLRotTXJYE75U
nNcNq2ZahhSyN2kMAqR8jy9QmoJOngjSt3TqGNxvzKMF9bhHYPsj98OJG2bK
U/iB9Y0WWGWj1AbCUlOiyYbYN9oZYBI5W+owF+1B+8ZyPX0/c1IbWBEGO6b3
TyuVg4i0/NND0u8Bi7dRkpNmoI02qbkFO4JpiEFLvyoc6moF6xsoNtfY7K5k
sT30Layjds23JbjC9KaPopQUWxwJJW6W8c79d0fu1dU+Ns5Xe1FmaV4hQbh1
UO5YxUmkGgia1B/9X0cNKdKyRv+DQI15Y3X/Fne+B9HHoPKwFky/foasj13F
Ec0RxIoHK9z2KSJuN8XOvzuEm2t1wxsbxW6hi/7AIG3ZtpcnI76DSukg/7cE
FhSUmXFYwSqM/RZ85DLUX5v3MBAxM4SNMFF3d+3gjMekrI0DeKhi6IqMOPdI
K5+sDZamtzSpwDXMpo35yTHRZCygQmJCidB5QNqO39gXTPOwyRvf1tUTmCUX
giI3L9UPVCPFZFOmlCF8+0w1ygtuS9fVJ5L5RdiaR4+nKm8OkYknTLGaX68r
AJL7KSaZkYmgXkgA4tE/Aiz07xx1x9fHAkJbwYz8vWKaY7nFzyAv6vN9cnho
FbDwOlLX7XirFGujewi5waoW1pl3INV7nGyHB7R8t6uAeH+B+WFhxd/0OM22
BG9pHcVY+5/Hxt6yBJSq1ngmhppfF5AiFzmbe2QAyOHm40TbUyOxRRjUImDc
zvVgZZn0GQtS+YXggndAf9lvH/FVs/iUnonbo1pxLuEQuIEorZKASRNrXBD5
CD5tS0p8ZhO9OZXvWez+SvrpdozccszgXyh6ro3/yb+bY40dI5TQKnbJxhRe
vzzFJO8TivdJyNySAnhbiivB0kOSGB6kWNvzIDytVX9V4nHuYXNyXTactO1z
cPti0YPxa92Adere4HLREzQgxMWGZC9RpazclNXVmM8H5QG18GV0qitzmzQt
BQIZFGNO1D8QK7/OmqZAoA0T1/Ld80QxAlYMTYiN/RNqW8Nm9r/a+Yx29qR1
TT2gIEnNyqnA1zdCcAYaFsp5QKjuqhgXXy1EISTfevKOaMA+Wa/IzB1q7Lo4
CD2suWLGRaeq9K0uKqnL3JlpVXpS8GUE3nlNEHZVhkTjlHYevEk8yiZHLZYw
OM2QZ71ALKw4fgLGBWO9Bsubhv5WVY1Wkf9vQSvASU1+oAsOmoI6X+aJm555
JRTilgBui0H0zUTWxhKQKML1ZbaIXailNsHQ5neKBXzRAPs6vu77gBllasyL
Y+eYnTT/sM/vTzBXupsY4wGsoXp5HMZvCePbPOCxmAnv0kaJgkQKNLwSEt30
yD4B/QsWw8hVsB3p7EN2C2RnsVqw1CgsMt2okjQXAkY0pkKk/MXteFrY3DoV
lnGgTXffanXpnwPiameD/x3GTeLG1cb/NjL8pi+XrlGyTH8swfQzqbUj4pxB
E6oXrlKPB022EAL97BLGWZuCG36CK2g2TuitsBNcuEf2Qp/NiWODL6Unz5yg
WZAuvanSpyJS1EQnQT+TNX5/ZNEk6MVSZF3yFpgno4TrgLKsJjRl08DwHRbO
Xe0iSaGjPSqtKQXvMRL5ARXClyyDg5vNzthVluwFcMNVvRvcqUN/988krivY
RWntmHbi/RMv88kvGBJOvAxQJgIRj2BVZ4bnwhVMOwvnR3FlTXPwS9Jngm9x
hPRhemajWv4ka/6Xo04tHr1WY1jjskDlVJ27frgQ8+RluOsdfqibcztel81H
J6Qf2cd1PcBrKipMIywqTmsTgTUw8FQgnjvbRyhbjmqbgL18g4DbCpP8WEIP
DYNhZ85ejwBBIZ0JzbcQtgXW5pdHTIISOQZxkXJv6nJ1oq0sEXa2LlwEyb1r
wZXDIo0vRFujDX4k4LuhlYBBMZypHciGJ2UXtyT6A/aPNE7phJglvCXLWXWA
hfcQbjv5JaRIKIS+CFmf95BTYwNEH+wvozYjg5/7Rika7PmMb5BtIrRhL5dC
f7GW5V+0bY9o+B9dYhv6Mt18oRRLfAFTKSgFPRmo/pzgK1rKfkzyKmfu8hFi
4HZf5UZ09d2rFHKrSOEzRTBPkW62d8OpJ9JJ7YUWqI7yaHdy3rchKNltd9xL
FfKxlfPHUqmye5/m6Vc7UI5r92y4UUABXJU4+fL/OxFcbmUX8v5uu3CuCO8f
AVbxzBWmhW3NSTdFreYqv5PuiXxiRaHW2YmnS7IOdtg1umaj8zc31YWD2xxc
s/KKiw9iW3JoA47PuMQaKd1kKopq5JjziJDiQN18cL7h1n7mtZLVP4wtG2xc
Hjdjg91uZ10X8hvWHPqCUz+cdktZ8XowpAzYmnV13UuFY76v9sKSxAIsM6ey
UrTgSv36qN5jafUYJ14X5E4xsyOhg3sUEh9pDGtP6CwEdWMaPdV9PqlGTvMT
M2j9TxImI1rxwZGBTQQCoaRPIHaPsT61utkfkS/ZNjCWLhLLDBuYrzPZjYi+
GExP1UtOBmGjwI/Zsk5UOdttAjKtlFDC417+DNFj43Kd9kELkxgL8sdpAn5S
GyAKsp/A3hb8qqecRQe3f/LWwtHzO1j+LGd3p3aIMoLTdQuszKYQRgtqF1dD
lo8nhojsyJ2Gxm1XnXRHnPdkai5IqN8I+lFDgzjM/Am/dp3tlEXJBHX4mSuP
cgx+Pm/eKzy966WzvsMY26b+l+F7Cxpm0sR8f/O9gjCycjN5vy+ix1oI2EvL
M+uXaUgeeVJKhtM0ovR6oPNW/s8V+5rw8oPnheHIDpN91qYei/ghYHXDZJGz
kjrm7iC6pN+/3xOqNMBw+RE74SD7HkO5Tgm9mNF/wONbJhVTk3de/4gQhjvW
I+SHaY3FQgTEKimp4KRtr79ANdsEYs2VbFFfs4HjXt5TUbQ3ipmEMQKtXhUd
eBxhy8FWzuMFnQX8r3oamaiOgLZpf0VWRfksdu3Jjog5X7rmzRh8UB/sHps1
xwo4fKRi0YFyFviR5TwiPMaHzIsrEj2U36yLJpiQTarv3pQX65+PbNfLeps0
3rhrzehYotPayaUd1gGR75IKlMORDeli/HKE3ZcbS0bvXAKD3ceZQ4Df5m2V
b2UngmN2hxG8SR/G0UFj9XgDwA6A6G3DJFVlBRDTEykK7rNwfiOgJM3/J7iO
RfNg5Zzio/A/7BRKn9eJ8+R9I62eWc651/OxYQeNRzpo6TX2DGyWqD7NFZeB
WXzxDrGIP7MTljb+WvUCC0ovPzq7Ine9F9p5g1xz5Zatf1/Y5WQ45cFhEfUm
nHksRBFcXzJg8LgQJsGulKOWi2Gia/00C5rnXl3kcCmhpDiNk3Z66LhoJTnQ
lW7YzJeRbLjYlynT1pMTzASFtEQYgUO0KXiWe6noN1/vddS1YTuGgmZIb8l2
IPPwdAgp1ToXDBIFwRPnWX+VwlyJg84H8dloDfuw4KcacEsJs8qdAJpt/WvD
SzevGTLYYLHKvGo7CPk+bNR7tNPQpTEgizfQCGcSCMP+c6jdIWcAsKfNFTYm
Qnu8YOPg1JACujmiEbJEO+yxJUeYMlnoYtawlc19qkDbvll8Py0YbvoK2vjv
ep7yOOuZkwpPY5DbRRruYaNzlUlHgdlboSZoTubkuPM4Mg6xC6pk30cZZp+i
5tPADz0tURMdXTJRF6vOBQ3dklHm0g7uzAqymO8Cu6JFPSso1Mo3Wwm93+CF
Uo30xk1y0mXOpym2/y04Pja4DvwIsSrsZvhU9vCkX8lc022XSeajfcxAQLz0
YY4Dp2qBLEicNqf2sE2XLZC+L51LAR3U41TIO1aZQgRgj1JqiJi0PY/Gxuxx
KXCKaggAvxoyqawyKz3BoQkVWUo2yMQq10Td015DovGb5LjR+cfb6L2+FjP+
c2eOOxbxCDKfv7u1ygXBSsXkFPgbxcFy2T90xwWA6IhOGxe7iRC+awW8BtE9
f7yqSH/tZ235p4q79sXKKrjjWX1SEOD1+/sWMl3HIyrLEI4bso1P1vpfUS+b
n9qUBaMebD2iwRbI+GJHhm0PVcFcUGz+eKbYLRSYUcWsSXo5dtfVwBMAKzr7
M8bLTWCR6o54bXLMQ1BK5pU+E3y6VWYusc4lW3XNOCnN2egYpt9Eb9HShx3C
6P9XmJE0EeVHGrklWzubS3O3kdRHDPmszByEw5FbG9ZBrDK76Tr4h0KlZBon
nwThVuTpJfnTAyah13lZ56GR3bBKIGtfaZnSaLhnEixWpnVfGpRbto+EJKDj
sevieRZy/gXigc96gxWrGVlW3Fr2136MJBMjHSfpc6SNt3FaHuf/pHhnyrZ0
LnuXIhCiNfS7WlDGL2Md6Tjmbpef8+f2bRZCEQ2gv+RlPGK19Y5krZznHO21
kWhKJId9mVfRVuYkOo6XFx5UwlKnBXcc4OFRKoM17W951qu5Z0sAERmh4+HN
hhd5JXjkrl4dLqMn99Y1XlsFQj2BtPG4gNTOJUu8499vHIN7L0b3tlPHLXfk
+Hx3A7BH+8LoxMedrcR/HfUz1q30RIQFRjTyKNgtAFYTlFlUMj8pkkh7eBkP
d/byiKdOKFyJsRxKYuXIjhc3D8/wvm6Bl/oOG8W43CXBU6LlZsdq/L7IFokT
ujooU1Nw5Xf/GVNSTYdw5YH2gbu3+XVYuYqFxtq+7lceNWIFtrTWdhIqE8jR
LXnstPG+vdtWdb+v2DJlkAYNbRBVSM2LYQTiEEqsdoGhS7CWPZmDKb+gOBPw
7VC6zQW+YG8jAkxiDj6mlnSpHlAiYPgWvQpQ5b9WtLkB9oMcdBkL19/3geLA
QDV5GrrCLESI9bfg67veoN/UP+5zf/Qt+1Tvyuo6HxzBCY3qhd8KBosxuVa/
lHx/u+ZvdZxMbP/PO6r4VmQiOM6zfsBrzUU9d7x5ChncecWz8CN2HMQqR/tA
LCvC9KdE/8wquy3isqv/24DKm2siM39IUI2KnyAhGGHPD8S1kEeFOcTU9jix
qbZNHUAc3qOc0diO7TuuRuyVG0BmjKmrefrI0bbzgaPYMNmjjpAqW9AZuVai
YuY+77ormthHqh5vDqhyaqjt89IBfqPXCvUddWdQ02jigAKsQVduNsAg39gH
Q4YHE6xdTCM3LbjuudrSeWg5wpfUEKkryd8rDXQ7PK490hPinw5u8lUW9lIC
OwJRS9fOc2ffd9yhTZWO46H5AnoOxWGsiO4yzcvZdDxTfmp308MLo1X//K2a
Xj2vdglW4cIm3yKGW5/zdiOOKb/iOCF8PW3HEUjHUEXo73oeszgwnzjIx2lu
rm7Axcvrh6Z2UCcq8QMSzbX1ZA1PFFxOoIvJAId+akeBVaXAmISVBub++7H2
fSdSNJslWSAg8p1ZK6nqPmK3bgZ/ecP2AFem9wI4vzfiJsx8TILwLtUOPnP2
Lz1djt8V2Z3PsfLso7L6PVdhTOrBXNAU/UlYbsX3FYt2Z+CJFpDSKYsLlnNn
27n8W3f+OhfsD2KZDRyjXvLUDca1J3ozaAnwNnZbCJrmby45PXuoAdBVIu/9
omq+FmcenoKk5tNKmAAooIKlN+rTDi6JpgOQzYka4rxjEoHZfk16UgjFBLEl
dreHgvt5BwhKmFMOGVFcWH/DcuVeHqBaRb8eeBgzx+CUt5A6rWegWiXpGsBQ
tb20MYPIhViPPB/NVH2fe3nAQTt7ijaFg4iF8oQ3sGZ4KH9v7jZKInajt6HL
BCzzIuXCmr9dBE1fPnLWNmsqEsKRVgpNrog3du1KXfeUWyWXyrNmh1jJai15
9S/qly22DlmZ9Lumr/08UGKJnWnO8smOjZoCZu9J+4x8qNEZE33ROZ5GO3Zx
0yBrkKfGeD/7atkBYtZhBW9+JxwMiEnX1NmBQ7gF1qUez8TWL8e/xjo/D+Fg
iZM14GuVXqEC/kSr/1w37e7jH7mkTsVfTUELa63cpYaxW/A2WX0ESch+mWDS
ggiTXPp7d7YbvNNw5Ek/E1SeHP+3VJigM6IvdNCFKr1VF/25R3fUy5lHaZBn
nuGIJVQAF2KCjPx5NmEdo9AgDYXzmaXZUMCyaQ5XP5L7dgy9GcBqJHVig7iK
BjAR2bNL0UffayWn8BlovUvTAtt7XQaXdrkC/atWtzTkH1ZwF8UPoLmNePFx
fQxLikR9yjspEqhhwlkNU1bbmpSynV+gtTN7rrmTbYMvqFrI7Jg5knGoF1xS
040kmrXJzxGoMnIZwAjBhJwO1X6dqw2Lx32b/n1fm7kqC6G6iX4g4xAWBzm3
9DwsYzGt8hv6h6XjA3WYlXCTfxZoVDf4ieZRfgPwK/KqqZ14TFn0dmAg2jth
zicCzNnS/qIahyVIC6TeHFjj5JpzzIBVrT+0IhIoj1nQD3eSV9a3cBv+xuZL
N74ozjYMz2bS3enMD7fXITmHdly1qi3VCd11E0vCG9pMzRlfyHAYuNg6l36B
71/3OEZs/1TBlZV15gRE6E4zi+IezmLlfVDyqiLn7UbjtQr1n51rZry7KrW6
pEuv9Mn6MxvLpFIhpsr85vgm1SWxl0c8vy3qPp8zz1KfUHmOOi/pfdmYljLG
UJEkwpcoe79msL9LC34Nz4mNe2OprAAutzZ41jRBP4sawjFqgZra1Eh/dp9w
4w6p5d33Yg3j4X26jMXXChRE40cq9E0JtE2PSzmSGcRSWFt025VrcVutJ6mG
cV6gJvl22UpZAxngIfqsytcGA0wfTwS8zseODZHoNjEB9CddeHJODKb5DGjZ
KiitBmNnNYnt9GcIlTnX0P7BHfKi7YzB4h1tWprcbY3/r5DsmPxcGmUkh2ni
k9t+1Dh3xf+AKRGly2+Y1XsUBmu/EKeWRtPjFPRuKLiX/PcugxowpFzc4rra
z+JZoKgQ4DjqTq3lm1b89bJb5DHyCitUI9Le6vQCwmx6jbtWvEnFoJEW6Imz
TuzTic/H7jWT6aaX5/qt7QfSqoGXfKqw8ExzEQw+lVqtdYcd5zNfakF46GtI
9VUCnaersbjPzwHW1m2vFB3c5v2GlTrNwSpH2Z+Yxv6K6Lj+ROWidPqBfExW
r0QcB0C7A6zWAlO8NqRgEl9+f8EVX58xrDBz3g/8ZYHR2UIyJmgnAJCx7SXE
xv7FCz5gvI5EHLjgJ0R9lAqY6GsNf+htrrQYVi/x8HGK4I6dAQJKKs1Dikyn
3k2b/+H0EfHvtPt++vtBCS9pgRVJtZgzsvax9NJmASd8QV6v0h/kVo1JqFLS
OBMSpzxgLNQGT8DKgqBOfPxrDsRifVXEus6fvXyW9+NEfoRWR0UUky6Q9moH
Z553jn1U6e4lRoe7Arh1LWq+A7VNk4qyIsFdX6AokfzgJu+BmKVqz6Yf7s75
Y7TEfmBuv8GUeHZMbBpIVix7/5Uw2bziKpgAMOelETlfr7b2oTMm9D/Giskl
DDGV7ShLld0bWoOG7+eIVR6jaQQurUTbyH+dAij7Rg2L3bUjBGDlw2EnIy+z
gs8kn+j8DG354KVm1wB7oMDMqqFfX1BqbqcnFPUMsec6AmZ9SpKJpDSnqnhZ
1zlu6JlwMfJz3j4MbV/jyYXBG2QeU3IWTQLxRD+jRZQ8T5QjTYE1HQzGijyI
O9KqWNmYyrSqd3oWb7f5S4WT9RF9UqoJW4Yg5x/uUrJ6c+UWhiiElg2HVbzP
GrFWP+bQJZKfqS442VGg/dXVXNAenQU/icmqeTnXISMe+09IY442vWw8+m3k
nDnrGxT2oWAJhqDCfxWtxkL3P0clP/+jWO2LIZ2g4fMRftJtaEbByxCVunmW
FrkoVS+bGTRewVS9S0dG/bFn+fWDUmFkQqAHNywrwKm7eZqW2+CcqyYz46PH
cYZ7BZ5K2BADqm05aBu3wAY4nkvobcIEzu9MvrPKi7bJKW0at7H/yLUuae8W
0LZMVUokpahLWTfpkZohkIH7uVOgIXAEeb3LUDrBYAwrH6CKTpiVw/XyfiDP
Iq50eVwSpK0r/fHoUU1pzWiS2DgC8EHiD6bo97C1I2pfJstE2Ys/1KnzzLR2
8fBF7aKKaYl8Hol3bWVlot6VQu7LCT9Esqq5faZ0NvwxL7bEXTeTo39v4ywi
TBI0lTagS/oT67xiAQnKbmAfJaIxD8wpr9HdsxlmQYyS9TimdL2M99oLSe3E
CCnD2kijBg99LSK1OGtdPAiIi9p11QOujQW9I5lRtxfMFPbDaVvgUUbb/02s
wNOXoEsYMth+9IllYVQGSrJJYD5BNnvl3M3i7dYplrPRdUjeqwq0pkwmzmNQ
fzszj/QuFNBv+MLIhyT/iGJNmEu//kmCaw4k47SNyS9QSN6LzOGySCGXYa1m
MzPEM6D5PdozvAATCxig/fnjNaOXg71UPotBBgQpzYf5FY99opRJ0lyRWkOV
sqTWz7qv1GjiIk6AEHxfes54mKtoScDusGvPe1zspCueikcAapFRy4CuyhUh
h12qcpIvIGB/660MKJkNgabzZ5vCQ31lIgnl5FzxVeJCa7EyemshAct25y2i
hn+U8oo8UofZj04M9rLBDbQxugQtrTNrzJZlpz2upsE0d3bevT5CYsjR6u2m
+TBb0qOSzAzQmNSFE9U55Tom8W0mobRcfASBsD/mARmCzGK3HBmQHt2/MBqV
GVVuesSjqJXizXfuO2zY+bQUI7EHmAGGrndV6bCMUcuQUpqRpPVzCr9GJlNW
O1XlsgYvXl2C1bMm8eUcikaPU4A7dDlSw7MOy9WImSptKVt34R5Cg6dPYb2k
/VENHGIqdzdx/1Z9QtPHDl1lZF+zkKX+9ZHxbEI/0ubddwBaW7m+X1P6C57s
J0cWv34Qma8DUU4LKeBqSkH4/g7EWqjBTLz73miHmpaL8sB1iH4/jnX/IDV/
b1LlrQExLSut5xHMOaMiGeB5B5QkGv8bdYtXwmE4+0q7KeiAsGoQTId6qIiN
43/uvtKoinJloMG2fAoHQdPOPRcZthFnEm+r2U4BU18vxTtMSIJ3QtL6wgGZ
j9uMbXLtUbhqZZLEyBYHR07YvaopBi/NKp0EfM2rp0paOMUy9TZ8MrzWDFKa
WpkDzsGdxV6qTrfTc4G5vpipygg8FGZlBTez3Ak06tiri6GUNBK+uPhP7U7j
RntuzMrHRL/O/peSEev7JrovheOILwLnYbK/fIYkhH8QBbqkUr+sd/WpGX6n
RkYh6c9U8qFwCuX6hlZi68PcKYobBW0YzHKQDEZ2d1jX1YfV6Hr235OoQFwL
HRGJLYsG4GKPKPLcz3piSn5r73qZ7pUDiC2kCv2CAapjfLNup/so4v4ALcrf
SPYl2EZxPomVsbuBsRpt2WHS5e8WxqXwatSpcDciwxXTc6z8ouuv8Vyg18Qy
Mz7eVZpahfwXrzsBPwaiAV1zPTWytjudVJaZyZ1Z0Px4RpqvBqAIE/zZz/Y7
QrT8doONFgwTh8jEZVuiFeb+y6XB24HerUcgCG0Ufl1kXsIsAQpud8pGKIty
WInaaHYYYB139MapVVYc7RZSaXmfEm1yBZ7noqISNVy6o4f5/55jYaZhblA8
0+Jm/cBxAVNinedPnRV54y37mMHK82TsQedl1AivQAk/Xd79vECrW/D0AupL
wFYw1nqPC6CbrmsnEGulb3v06dTt6jkMVPxm2FfvagdFakWLd2XXppwde0T1
5NKQybng/1W2493uKcI60DL3k0RzXzEuEvjZXEM+1jbQcNcdWAFaTRDcBFsM
25R5T49IdJQu6sEi7zwGqjC22qGJAFuoTKcwgl+qcMmF5HOIZVlc64jzYM7n
garim69sVFY/CGFi6UXZg2cJGtEA0dfY4Ei7nI5pyXK2cEsSWSayNTZH6ta+
gPwI4VV+Qcs2yz3Q4FwVFn3phTyIWL5f29j4tWJYd82R7VVoUPfsXQlA4ZYl
DrWWgWS6AKEyMNuePgzgMEDiJyql406viW/3A5HFZNynPusPKPpSIFeibYH8
hEBD6sG/jKWn6/Ktidwn4OsXVqYM+3p2NoUc4PfotlyinjhpHulbV+FTHXnN
Ll6qwfCcFz4Cuvv9stMO1EwbblltiWtaSyizJtpQ1qj1c2fElaUAzJ0GaZdl
1Xi5eKrTQ+XUaxOcuaH7mUq1jL9GDiGGjEwN2Z51mbesEp11LA4fp2O7GTol
woVp1e4UxLYqN4BT9KYk3ZaCqAu9ulmXG1ZCtQDleYOnELhNF1rKjVg+lTLc
dyY5f+Cl4wKn655omH+lqpd/xQ9ck2Lq4ar3+lWxoH4snBxeVOUTiGL6UriP
hbzMrnXpa6vyt1A0tucXJle8+jlLPBpVBLK0igpYr+J614GIZdN45jD1Bkit
Y4W/rNtb3abx+RoKj4nKTu2x5EOa8l+qWZCHgA/RHhWxiI1+3vzq3znRI5Ga
54lYM2YBUs1l7sniVWdyLcOasqk30MhdQKgXB4U+beqL5mUpUJu/7pbXhQAe
5LnPyCTe2dE1baJWB0N+Hb78q/jvpm5RtUSl7pGbxPdWgMwWrAWXcev4s4nV
rntbXVXGmiGQ3tFgIdTYEj+7u95YP6kx2mRtqMqB2pk/3U7HDGXVrbnGZVS5
yTvZ92Cz4voQIjxLFFSK3N7DmiSoMbyXoldltpbrJC2f7gxoZWSsdCU+NudG
Calaq7uIPVdxJXI++yms+XQNIFctm0JLoz6+Sk6RTNYw4rHeSk7M2kZ32MIK
+cOAFbcQthVkk7+r4hHOgIo7xovgSkMqxLDvb28UCixCjGNFp3yCxAqlPsB9
SNiYEBRBIZ7rK70jkx8dK3stayI6WNjs5s8vPRfhfbav/K1nbm/bb3Zeitvi
+LESa0xiiVVi4hetfVlBHPpLu9eyXRRi6GlAXVCXyVC6+F/wiXVs/FTdnEMa
ybz/51p95WSEbslaH13DNMlfsPcWJCp5TpbUTXA01Exd1iJ7LCjRzWj/w+SG
PxroryiaVGb6aGO+B2Qjd7Pw5IEFK10dWhzDeN0Q8AcZBzlUedxgt9nc5Ky3
WjJNx5SM298vVdjvw0fPGrdur1kEloKaGYuiOOwGHbrm+a5vk88YULOfY3Hb
a9gO7Zh+E0IXb+Ws7uqunLdG/MRAMkDwakXyro7D0bTGLsXIThMAZKcTjT+y
bl/sLe0HDoIzGkfbEg/EZ5QA+faUSz1NzaebmA7/697G3taXG/xTXPNpgC0Q
vpKsDFPEXRjjl6LQSD9HH/6lSbzWRVwLwoHfCKSWzIiI5RXa1kbjwsXEklaT
jrIHhm/9oOtOmIqkOYRcbI9UpTPRTrz2GGtjcD7biz/M/D3GAGw2lmW/wHCQ
toPpKLfflaZkNEXUjccy4d8mUsf4KgA0hQ+cJdYitEAUY5VmSmz0irMKNDa8
PmwbBbXrNHDscCFtQxrRC17bWj43etyoILNO8VK27DVtU5DFuB6bP0A3igjL
HvaqVjJyh+VzaCHqNONrHBeDeZKJDUXe6n0Vyx8Y7h3eUI+5opEw5ngDj4UN
mRbQHAaTxk6FrBoMpDkcpzqSlGWciyr7sNM2zXpn2tkZKs6OwVsck0CIYzvy
qCPDNYHRZnBwppHekFXkd9nSMGFeBGvt696r9Bb+qfEHcylUMFYHOhNeeyqX
K8RxclPLpG74hPP+wrvFszQvXpIS1h+jHhBOnOkIRoRkx8qrchFcE7nVDbqC
4HroDWHJOxWPrlL++LTLjH3aoQjUnoZB/P5EDkMUFdFfJJYo5VfZ99xPc7+y
uq6O1OWlqx+T5psPZlr/A9Y3xOrduUtx8YhUooFUV2Hiaddm/l92I4YIzE+k
C7Zi8MXn/huhyvKBiYrAz7k1GqDrnm2BsaE9GCoXbNqgz4MgKdW+LCdB7WhP
0B9HTzAGGGSbhH5iib9Kzv0VI01bJWdtYildCMf3OAKLM/hvbw00enY8iXeY
5wrzVEldbR46x6Zf/obaytsgnzFwuWOuixZADNlIkkIj+giSxkZdnDYXMiUu
5dBXzYNum58/NzuSTlAynuhKPQAYbPw2hKabYp+fRYGpTs5oHCiK613yHBW0
L3TxBv+dHs8eyzx0rTkeyDuLP7jrZ9LRH8Jqj7zBaYpEqKhhgi5GVJPUiath
9ekU0bW8rj6aVq1WN89pAA7lBP7nBomssWpHzNJHNPAchg5wQcD2H8T3l79j
1O/9dC3KYuUlDkbeBh5XiVjuSa8vukLaI66jeA3ckCuWb4RafBgae0gfhOOn
4cmLWky2nAH9mikNW2f0jhVUr1kvkUKDHq7VBiuYukB47Hjmq0wKW4lEIhUi
hvNW2h+py0EZp4bG3DRH9s3f3q4FgWEZBu+JzKxmMfEVoZA8FhrkRTnUizU+
o95XwfnjJjdAv2fCRS2LvznNUDVUZsnPPLhH3DJMZeDTL+m+OpPJQnot0D6i
7vJmXER+duXzSB6Jwit0cFgMhb9On8ay+hrdZbakEX+7Jp1yk/8OFCMPE3Rk
yHEHxm1B1ChV+dP/zYo1fFmvQiwcuS106CdNvnieV+fQQpiHynl0lH0Fo0J1
Xx1QGZ/T2rzbdm+NxVgJRAx0mRlIYuTC1vaHfmI7JXZqy52fm+n8w2F2lyyr
QCs5Zgpai4D1U09gEQ9jgHcvFweKw2E80aWlql00cy8zrQEPJxpOkOTkOTM2
CNhONGpx4cBsDqy1QHdw6cuocfgO56H6VClS24lIfTm+ybgXUWQWG7x64T+m
R4+JlOJbYINHORobKBC4rFOycHjgshbYGT5GYVarob2rz41wddWgcj2v4o4a
VUC4Mxl9gr+VnOxWpGExe/P4fXeWStgUYPQYvj1mR3ssZQli+YvR869h95M7
syKgYoPoPfR7l2+m16cs0P94SRcosk+KCefT4+WQvwBVNfNWKqTae+K3RL2o
uKkfAe61P3asG0Pag+U9IJU+NumrF/Sgg6txCpdFuzolUoBqKChDYpiegFGz
s1VwFBUmEJdt9y9FXHvhk2YvEm5TLETrFsHgbfaxxKjLkv31m+vC7/hkPCyp
A/Ywlz3PSMNOKULRLZXShql7rAMtfhyfoe8SKyhkHwCaF7fPIr0n9s1Q0TQK
g4A62owGiEQdFeHbZQINxk5w3asF5mqxDE8BKJSBXr6/MIaIhLyTyQD1QAvN
Iwi11Wuzc7bDLMz2UkU7zy1n+lwpAJTonuSWaCfiWyTAboS/21J0SWAh14UT
i6tyg1xxK2/6CdKZiLM/FfONRSqY8m7+Pzvttdf0+WFFSiZMVPuS3cYF5WmT
6yhMN4/NeKhwWVd1i1qJ4fWX5d8/oDPd2TUEzyKjYiwOjQmM1cXTHqsT+J+g
SoUjaSc9GvTt2m5h3HCHiRvHvYsPiDTwVDhXNADJ3kQNVALPe8gcwYwP13KI
iEGNybDhTRxHHyr/Wi81Ywz8dI+6QVaIILUomwSf+HZ/1fMguOHOCplj0PkC
kzuXqMcqSSaKs0q1ya5oM9UxFl0V1ZjUktShp9uSFl2AB1cwDi4iHysDs9YS
t8zDknm3z0bO1lEGIW8dEyM3zr7Ld1roM2CbYlORMyyGmxyMmt62gt14yBsT
g4S+pCs4jjwbhNTfajmH6jQodM4zuPzxiw11vHMhjP54xuYbX7SQLSmDjj37
oqInJZJiqI9f3S2o/se0J3Rom3pDNmnX5LIku07Jn+MNHZ2byEY3GpOi2jYj
Q26L2IZOMeA2j0OogDFXLPYJI2q7bzihTM4n5O6mOiZjNci2Mq4Ts383l8N4
ACFZ1nNd3+RjYljfKhxzI/EDDPXJOncNlfsrS1aZVN+LYFYSXWHmWx3fnz6e
dMCEr236ZoIdUY68WwiZBsfKerTmQUPLVzQu8m7NE5XB4JWqaHUzAQa1AeBM
cjhQsGMWKtzd7Ufejz+SLNjxLLRthaJeCu1D4UQQDF8vduYd/rwpLmp6GQAO
9DEV2ci9fFqf25O+qC90cAbjwXg0fNmvlq+HkGEuU0nflFpBfPM0MDwHDzce
uugE3RdYWkpPxCr/z0u8nL1zttLAWJBn5RNX2B28H3oyNcLs5qVBiB8DTvWN
q9l1O4MJt5z9mQgakhOf8KH0ZskZkEdnRX+9foW+v4EQ2IlGdjRxu0Pz4ZXD
L//AnKQDrKbIAZ70+6Ex+uZ0+Vh79EsPQEns/xQTW8u6/9JSTDaZoVwrqQ25
/lafZtFcCAOROU/pzh4R5P03UB57jcTxxvDc6/wC0ZFMlvsJbO+vnYuSe1O8
7RnlMzSsCLqJLR3zCA7wG4+EkMKCXofjJvidt6wmuVHK83xYmq5mxZ1K9awx
GvzS1E5s+JUQalExubAJuCGWymL6MBJA7606m0TciN67T4QyrRVTvk/DtV4l
eWeFVl8Kuq48vb6I8P+diHHsNOYP5RkgF2n9Bi3cUNU+AF6rwlsZ324SIk71
dVhWH5BpSq5wzYJr6LG3HwP2QiwY4zQqpch5LYiVSI1AQnAt3FuNSlMmVcbT
yTDJJbjV8vO4WMh7y7RTygjzJPDMUQqWVpCzB/aSvKl5s+UCChzo7EQyGQFs
OBBWTQb7VI//9oRpkSios+/nweTP5cG4iefZluoTnDM+J8jomIY10fsqnd+1
Tq95GGYcJS5MkbcbJvPjRH9LV1mjA1j6zYBbYkkcErzkaBv/tnCKUI/inJhW
A53eGVmZued2Bc1uqH410uKAF7u2FjTxA0qCUWRmZTLKlk/3hSq+qTBKvUpa
H8mQPEq7ff48dYQWVu+l49Uhi2X2zVWo6DgePw4824H7eSggY5aTp+p7CuDB
FaQ402FzsU3vP1ky5LBDntMzHI2Uao0XG8aeREbCP8oyC39UYjy8iY3lyuYm
yPNcvpJdYrkzjlnVjMQAbJYTjtUsMU/H9YIYV6z4Bh+U5h9neMu+TQjIbHf9
nm3La8QK6R3q7yTUKOfxeFR/lvdorDqDAS34zpO31H67cJf+iS0DHhSQjZMT
mi1HY2X27NCeRrXP3WP+1BnFdWv4StlvXuyabl6X7yrb1YvWf/Zm5adSBEsx
K1zQQeSlCcZn8NT3PoKx8KN3jqYBIcNyhLonNYxwHi96kDTNzWPGqx5i/xWG
Q69Pn/fGQ3KUCd1YHLoheJnFVc4nXx+T3yMdtcM5UWPTQ5zdm6VX+2rAHX3w
MC3cwyRvchOhxiEt9m9TWGFvzVWrWv19/u0ibxteEOT0o/uYoQkQbhOjzhpU
WjDPqHlzBAOERN0mL7mZJwxkNsdQD+Ie/+FqDnSYnufnZAB/95wWsdhAfWuR
NJqDvksn80saXCEqxAYypAma0IIFk1a3gGWEIa6nUxuO4HL+AWL/76C2KnVy
l6Iay1yUEz+i/5RYRIEz+Wl+LhnYrXVsitep9xSk6Qt+EcA2WCfSiUjbAPz4
cuJqu4pyH75Ef7xD3//bjEBI0hoQjmAh84Du/hTkqzibACYIDvidU2PgmXah
YsP4wZs/yX3m0lxRtatTWcK4WsyBcbrvRrqwEL0eN4CGlAmtcs9qfNH6qYbj
b7w9B0LQGvlJQB4U8TtIogBS2JVXC8yXz53oanNtSYnQHemo/Md0rA2cIjYe
bUCSXhHse78/NUWmZAJr+Va7jW7zfCjpzJs76liWvqucjcdL3Fe9/SI6VPXZ
suxGlBgPIBLmOYIy2T1U3vVu8eDODuteDuiD8mT4xWawbk86yDbHZKXre1T1
5pl9nyKC3L90k7Pvf5SX3eiL0TuVwKkdOvPg9l3dQuyeopcDtTKsTMbNlCgr
cmTVs5WFFGy93iMbg6eW/oAP76o5a7bb/i9WVdIxwhkNFZMWEWqaGmqk0Ib1
tCYcZzgmv2MNgjj7/fqvccCSh5TGAHsAZjh6CStsxj2tJgZ/+kqGz/e5rOlO
wf7zTsKrCOeWwGf59MCUrf6tPpshSEs+qmlPWCbZZyfsO1EGxWhrdD5sRYmr
vjQ7dBYCb9szbJejP5+Tg5OxBsGnmmDXtQ4NmKIFF9KGK49bMO+gB1XHf8wD
6SsHO6XQkeqY/2YHQCbaZ4dMRTs9Y0KEgXnJQmd7Kfu2o2sAd2nehYFGzjtB
oYnROFqRxV1aQtm9UmHbKSY6QN9XIm3DNjgFnrAWv+W0mdF22UqyY46zn3xd
Ge7NQHPZFgHjydVJBkrY7gmy+N4MQqDCwoz1RAT6J6Y1OvbgJBPgzE3M5q8W
xeAuoS5Y2SLRiBAzmUEeKXdstwdCEXFIKl3QKMFucJRtvC6vHCKytXEdyEvl
jK3ab+BZaLfcKRob7X0nZmlGi8Mm0DCFRutPzwMDTpwvAML7NxwmeKeFQfZw
1JrLF8EZuzJmthrVyFIe8G1VbZsUgp9vZpV8O/ysVZXbDpGJU98/kGjMS4JV
s1rjKvZI9IMHau5rOwvArNImstMw1y+AJmAzHoRoAMpc93cod5WLkzjfojTO
Ac3WR+AjGp69cbrslu4O8mDmA+mEUfiNteeGBITI5aM87LbQ2LDk2EvjHDBY
DTa5QH5Ic+DZb7c+/M0SWH8r0r2t6yaykQH2HmCMjL0Y2I0d22FCJKgVyVP8
gSLlbXytTXF9uj67bjGXIRhPYZLh5O9yeykSBdcJ6rP7n/Zl5IJUotW6yI38
Goy7K/7dLjEHaxC2i9W36v7Fsoq0gMcOHP4YeVNb1qiqxFkJLQ+t/VgMYVOT
6vyPLUrA0J0aS+p3NDDWkd6QqzRl3UIx0WnkyVVewdfwqwl2ouRWLBO6qZdX
fvh8cHWPdfx9+48zKh665wmAtJy9qq6uCEjoHHrPCocEKpn4If+mZmtl7uWC
Oa+IlbgPRd/b8KgvCHI8+aLq/CEBcUKtMr3eZehbm1TZjZBfgZL3JNvY4dgT
BSsyBosZyPF1w74E8LIXkJY+XmMuVVXfJYfec9MbvxzCPwjD+CPaMypg2HEL
gde90Gu0S/dVr00UqqSzNU4+eFpmClIoIWZYbIQ/NYxJJem0SrZkYlnZAhD8
eO8W/2iJ1/MJD/1mL1UwsCWRegIe5qX7ZZ+pjCA/+WEapT0s8gKRlO8KHlqf
G5nKXZvci9yx8v9thxHBHz5qNLDiOYkpW+JNPXI4/gVtKo53tROREyS6ldQu
KsQ64DgQN/66mxmz+FeQ1K3ZmCRXG2Gok9E4YWk5UAN63/8eOFo5JeasIRFg
LDI+CVDR7eLhOdIUwGV/C0oZnQdiH9TOA91bN6dyIvtstml4+LonDhnIcoyd
NKtR2DQa6oJ49JYExapBCWSkjb2PlMrlDxbu3WBiIJGkT+dZqLLthHBef7SW
Hn/5EgZa4kJSszP9hAfOMlgqLzZi70vW+xffTD2oaJSfIK8ey1xZ35OU3i5g
n8l/OXPX1ecyJ5sZn+ICX4XgekBbsyZ2CPNWSJ1jtqcFXaseg07UTBgimmkc
49in2rjJpB7BxY+vDy1yJYR5t2cK4E6MCXXPl4msZAay4VUaTqmiT6rzBJQR
CT/vVw2DDoiLKrPpykVlMxWIhCSZFQCIvJGr9/x1pRCDZlc+TEc3bzTgkUQe
4Wi/rKczErvA6DwDWmfwftmdZCp2GIAhBq9EitpaR5Iqgradch52Xh96jxui
jGAW+WK06/WdyvQVNsPCPvIjV8wEQx5UIE0pIVOqNpGyhyZHSUwwSYbIfFz1
xuMdHkLXNHO7exjRsXwbirHyPoFI8CBxpS8yuYfofJ23ZO1RJDKfNvAri7XT
4qQeror5+E2GuzTE/+gxUrSZ8JCN0Uld4pb0Esc/HU92HNgWpIAJhmNqWhpR
AS3UAETgYJDxQvFfCVAhqbnCEUbgUCIBJpqEUVvkwLcv6XeLHkJVhQP7K++p
lta9kstYbHZeJF1SphJ9XKYnAa9StByYPF+JkqT1uAHX/ObiPK5MYTgZf1Qx
YFKTpHl9zkFvHOHmXeoMOiYv1PcqeIklYMnr6jeTtsoOHoXyXIaaaQD57x8q
2fiFW2mryfUQI94No2OZWnaaLJwR/0OGGd+puQouRuIy+DzKYY4x8w+MaBDg
HL2EZGo3GfJtvwlmAz2nefoM+lX7BMyeIr9WuGA0zY3OT5w1U94g4x9ecSxZ
2fPl7WjHZmhZc3ckjoe+q/cX69qwbQFSGSzvmHqTdcx4QkGes4b0oBh2VPsv
nOxuVZJvyTa4PrxuznT+bk8Qv7K9CMmH8kNWcEpkh7S+xD60xRX2Tv/K4Ft7
8riGYYHpjvhSO3DuaZh+vauQDS4pfM5bc97K5Tv53erBLjXo27Tq4ECKAIZS
ShVgznyIYS4gZOb+D9il1MsKa/vYFrIFI0gTzHM8fMb/HLqnS4QYc8j6EZZy
7L2ROq4sSefzrCval4Ys0aFFIfZ24oVRlzohfQNhpwZ+igY2xxYJ9vfPpEye
FFvhUtZPdJJR8df7z1jFjGfGPXgKYs9Fa8fO8Dv5Tl9DEKH2uCxvikC/+fUQ
BLeZ84xrqaeTb/FBVqYbZT8buF5NgfkuISVXXTk+HmekR9CdjddxvS4ICqXY
6Z49Y8VBrfqXL3RlzavAYOlgC7tvAl3yit13M9+aTNkwfgZn5YLr31wPFDo9
m93MfDBV8CILAuMELuda+O34Yv0uXXuySd+gbQY128zEIFD1T5FyYRdw3Sbs
0EWNfznRgOfm3s1/TzDI7xhnOShSMwPGEL3jNBV5dnK8hsVp28RDz4MHhnNd
54vRKUY/OEdT5QXYk9kTK5x5CGx8h673djnCDu/O+c9s62DwL5xPVM2ooUD2
wJ/Hg+0Cpy5G2/cckHE9WEWpekK7e9a2/MB4aGpmjgob29IUq+p+oFUnXSjY
GdrZnARGfz/+VZ0CSPJK8mT4TOkIzpnKOSf4Q5awYAbD7b1YsRzh80e+fPKs
ha4IWoYE7SilJ651ZTsW6V4Ir7c+jfz7qCgFpNKP5vDnks8Zs8li3oNu60LI
Lb1LNRowDiF2RUtdlxmzTsTbhW4rSqvASFD+HFRnErjN3sHtd6FuxobhZepS
pN/d5yEMGNPZmdpoHduNFQpPQt7p34KHAQYs18bvZWFa0GrhVeoQT+07O9x7
gdVXt7uvtHFB/Ns5dpxIMvtTj59qmG5zpGeosPnDJY3TAhBPcFKCTE3DbGeR
FeXJlRctGGWo1HYpHkuuQDnRUpEZbUS5Kqd/X21Nevm9eZGFMDgbLYj+9FFo
9Yhhb9qxgtwrt2IfNmkR9baz4N5Lm3yiG+0/oUZW3AWnAI2zIrJuRwUztBm5
QpjwHVc0HTpF4c4zWlaS+14EG4YniHaqY19ycP+67EdhmjcHFXtMstvDlafy
Rq4aYI8nkCZbyyVWNCpuEfRpvBsiVr1eXagWGlBU6AlWxIWdQ+gj/xxwwXof
hQtW0/4JyAyRN2rMx85NY4qnFSey+P38uKyDu3EG2FlTzKAksYTLAhEUAZN7
FkpbpRBXTX+i22IYFx3nPAaMd7bA9eFGO82KryFcAWpefxZSuFuafeJepqyG
R6C4BEqC2xav2GtQQz4P291uni4eB2FGNUe+bUr1m6399XFXwuLp30xljhG6
uH43Egp6nd5elpkJdwn+QPOQlxpuLG033lZLPg2CLXj9e08MzZrgF3zNvxDv
u2kQa0N6iT0C2FJD0NXoiqZtIB+ps2t7y8OeXHFuryT1Gr1UaiZR2iPeHWRn
GZ2nrgngxlIDwq3Zt2bIn/3a/KDfkaRY+rdmgUtPhC+ANsxphA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGOiOuTZFfw00rpzHpnPGWKFEDd90JSGD3Zdtv818pn0jl3GCB7MirBAnHyR6B06tOkPY7dw2l9w/hbIyDYEv+fVJeg8k+OELnFT+UDG25eaOU/N4Uq3YPPFFmU1Vh6cgy8IXW/LZh43+wk2F7m22GvsKjp0JgFiZ2b6Yv5FTcbacdBtniD6yW+ruSfJLb/ubLC28ompIdEHqFGPKIEHIX8ekA9skkZtnPkcx4mW8kZhxSeukb7c2k2JImrst58LJkeBIxFEID2YFO1+hYb5pzCyKexHduHtKVN5cjkRZWYSTJ67VoaJLf8VHb2ntHRsi3IYhpNELA32B4a24ygSWpBB0RhQECff3OYVONkMQX8mnafVY5n27Zo72ErZBCMrPpB2Mu/QetirUVzp+n6OKO0iYmQZY/ZXkDTesFyhOceuL6QYYO1qxv8U/eflwgnKm/2P1I7cy3qPjr0eE9cbmSMtvP+71IZwWITKdf2Ra7vR1wBo5TbceQVYyhXaIBUIWTOJKqfZiCM7gCZ5eAY0+AMwrpVFRl+7XgeuVtsHDiLsaVbcpiRMySJ5GImBIKyzebUlD4u3gfBeCK72TMxrG9CrPEuhGH/1Jj4hCNUtEToYco0EsixQuvifWIX0S/aPll9ljReapRZd4+GJ3Y//qAu19KLipvu9VxCZq6uCU+z2cmKyI9nth6aFV8k/B7mRpbUpJDy1Qli8qQoUerTybEgGkmYrudsTndvV3XvoS9iuy3rbiW8+QcDYpOOO0FYJ8zO/EB+aduzv9ehDwhqJbYTX"
`endif