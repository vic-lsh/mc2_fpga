// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wAETUUVyjI+Rck/8H33poHD/DObWPawSH93n6tBLE365dg8HSPSuoEspoQmi
ZNfy63xrC8x1H5j4AgrZFYrvlChoPCg+O3dg9wEnO4B1j067BJWi45LoGzD1
3LtPlqNSiBtJk7nb4KP5AKN1V5/00HdMGSKcrijQ8hU5UYJaBIw7GE+NFgeF
N7Z3Ohd5NvlBIDpYnY5rzgDDgmc+G0mqU17VbB0DPVyuaC5RVPrxUrOMUgQ1
xkyl87uEvQQCwRl8Vf+UQDMWRLM0aWqBrDCsnW8b3oXUBE2krmxcYk9JZvAj
2/l9FlTPUkTrIws8o/yjVAjrpmXeysdR1+eqCJFAVg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ggntoyJ2zYD4X/m+8dD90d42gAMoJfOnIbIWdAjjocj1JEh1qtobV12iIo9f
Y3c2J3CTWUS1mnJ5A+1CN+gNQe+OrK8pdHXnyKIqtuo2pSMOaWfJSTGRMP8U
ShPCDIvLpHTO3ySJmPwMOIv25wqcYKjpSHu1WR83lRboxripwAkEeOF61W4j
+t8FVyNspKUHWxB39lG88dJkV9PtqGEq9a9pHwRs7s8r7bOAiz6y5O9NCgi0
kxgdCvDUwfE4BwpfjMwTVuvk4oM9Ed/8ee8Zn/0XRCLQRKrbc4Rz4NrGE/xN
/sMhL92AwYMeeJQT56ctH8zINMVvG1pCtIiG7W6MgQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TJr1cuHqk+7F+P3taEn4QahiMjLVHnXEi19jttcLG10T//eQ0N/0k0uUEeid
+YqUWDB28Pb8EPc1d/59r1qfDXplawUbFmO7DVErW44nqq8Gula5QPZ81Xhj
nBxsGXXEErLmUHfv1Gp4BdD0niN6FI1PGgkYTVAUJcjaskj45nRs4aX3mH1J
sf3JLq3nYLeVrY5Oj37iryS79kKj7j5TZ4R4sNEkORLuGx8J3qRy63vQcTwv
JKhBDsEASMsUos4Apk9wSxw89NJ74EXPRHPsivZnCUrumPaUoeYEZ/KMwcSe
QFTx66d4PAhofOC6duO0lJTlUWvV5VcOvPljIJKrag==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ASQYgvv7Jh8zkgo9fmkGXbPjH0Ue8iTlXurBv3F3Rrh9j9qr5iTifC+Dc9Gq
ZGcDtr/pkDmI3ErqC3KdErhC0/VW/vkMk9zfuXIee1M8K/A2pK3Eq222HHe3
ElRLTTegoMEx6P+ZNl+wPu8pGk1A6g5M0pREATQoQigkqb1Q9qqZpob6tLLy
+jTzPXXYRphsD+S88Kq+yWHaKhvaEp0Yi/5ObsnL3qbmVPcY4qjS8CFQh7lU
OOWpLE6EUOATVoEzh0hzPuir00c+p04bTsn6viMgrcnLIeXO3ARfZMh7buhF
gYnP/yf82uF2uLZw5lnEH9bLiPG7bvzFyTsIgiZMoQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aZOik42Jgr7Z9ic+Z8Xcr+kAO734gsu/yn8PxtNFLIALgt+ollZcs7CaTMXm
mIx/BWP/o4+QdlDaTgb2HWBB1r5WqdatDQomT1mcSo2lahyfAdi1MXw12tjM
8AsHdoQnxUQDfjcwtglm9pDcSMyRto1yHiDcg9/zoV6MgVhanHo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WC/dWrP92NeSEeGyG/490frLSqStB19oJzKMmXXI0Qmkxy2kO/s4F7gLPoCv
GG9MSsycUechXyxLPNN7JpAN4jUdDLhyZjt0sC9zowMDuCZDtAoFLt3xpP9W
Dg6+RykVnIF1jMczTDkO+ZcsKta3JTpvikhZRTBn8GNHfCtNnAm6X3U72eyY
KDUi5hkH/O2MVS52gwnlmsJXW3rhgJBirsWYyRQlygQ97WtCz7aHtPNUVcxI
MGWZhxo1QJyB+dbNC9c0ktgqY5wkYrnfrI4NkxYEuwE8tLl6Sv9jmLkJgYzX
vah/GvhAtk16gVONYd+7j2+QZmKyFSLs/uaWVmLOzdQlSYtS3xxkAMagtqIY
EEX51J4GlCqiV25mNMKOUA2D48qB8twdU/SAbz04eXhkKSi2fr3qmeZly4i7
dXQdX9Q2DG+MufEURx8we8ss+ec+uMbGo8FbVDAqewKJePEuQ5cTt3DG3Wk0
HaYyWgG7oICyI8fZe2DFIRCniMhC94ja


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iQkk/6CTm7e8qJR9L3gQT61f36EFxFieWDGIupN/dOv2NuaECP+UG/AUinfJ
o3Rr3uxvlbqxyqtxok0cCoCthAuMvjKIxHfP/3fiU7N9I3u3hU47zi2UnVi/
jGL0xO8BVQ2NbSSbGEkTd8LfmU1s9x+sucZA4qGqZ42q/wrDE6U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QvFNcGe2mMNZMAwH+eRgF5P/DlHA1rYD4CV//GV1v+crjfllegIqv/jFaiLP
CYYbk1eKvtq57AQXuS5CX7Gb4U7sebuCz8mzXOgfy8VB67zvMtZcxnAlcEbc
HBd3KjqDC3qv5Z7kAY6RH3qtTV1YaeBPVn/ZY82ta4tX0TpwYCs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8784)
`pragma protect data_block
LMjaBcfd3OGf37E6ZSYLwR0RnGMbSJHNj2ABRSnhjHqphXCv9bUC2PGlhfX8
PW8YED0dmmDpe3d5zVUiX+d8yzn+MosTURyORRSG7SgvppXQt5Ced2v21Rn/
6IYGtjcqkMAZJIiKLQLLAr/gZlM9LtKy2qRF0uL8i4hw1uVzlRXL23J3xjoj
RRMD1DyuEPy4s7gDFblLnf4QQNIlVfiFrz6nJ/qcaiXB7t6pX1DZEi+plMCz
1B9rDw6HtssPHa7z1I6OsnzK+Y5Az+Jreyiv9AQGUgCbMwxCXAZr3j5/aNPL
PcPFTwtTjLB2r003M5mgfaOgVIM4rYjmPJuIzoY2KoMol1+k04Xal0RxXsbi
TwtkHzfIQBlMrt24UL8vsp64Q3dc8lGcfGeuI9cmYCc9VSdHxviLjsFbVaDA
OOL3FiSRVJ9GIbeH7oLQ2y7R5vyph4glfzdSqrX/HFu4i9WofdGGzN8oh8tw
lgZxtnZRM83FDmoaslFZZIFhahPHXPttj96yZP5aAxzrJc75cTPmkxSf/t9D
RPp3XoOz3jPxLQ+J7sJKDzcUEJSSJVdetWbAjq0mh8s1UQf4iQ20kUlQ5b3Q
70OcgEKyUAkrCL9nFTWz+xPXdOOXpJZkfdvJxxK6fg8q0I+VXvjqzbvG+XvF
NBOue60O9ZR2ODyJkCk0hLrRnRSHt4UowwKVI46zs66qoErWFJSvpgFZ+aBf
Y8BZSbhN7tVCJi6rUgemag3kEO0UXSdqCPnE1wIJO5FoB77TyM2WgG3T6dWL
6eaX2KRxTTjKY9izCl2pMhrCLK+GQXZH5MOQBIKNJZ2R+LlatL9uTL/cdFKL
7TD0KchflCE8IBASQXx+Iy40UOAK1K5W3tHt40daa7hGBsf5wogqTraa9HHi
mGMPZzkpyERba9bNdgtn5ms8zu5Y0DkGJkqhFrD+x4lAllD9tguuQ0SZLN6G
gFkdBtuErH8vft8MC6jmdcLODoAByxbhh7p6i4PUWRxMCLTuPQItOU7GIitc
c73zT5c96z75Wy5E7npTPLsfwyG0V/xCz62yy5WjM51UEczHIWbCSCRbp31h
Tt8wYam9tUkgDdy/Iq0Sxj1slHzN0Q1jhIDiqOFMbWD6paggpGkZMFlIYTPt
4/vHZQwJ+YRkf78HbHJhBfzYjHMMZnL7PinFDZlscbkAw0SbEOV0sOjNbw6W
gT47hqXyugVFKisGDicrEMIpsXPZghoUPNnt0GOWHuO4LQLCABmBhBTRpBTl
DuApvQSYIQTEvqe5UySFyRrvEIKogbHcticCZTqbYZrsWFx6CZJB3YFUxh8z
KNdc+UK9vVtmT1mMQ/S3j9684TLmkCAIrNj89cqH+QJDLEPTeMgns9PCSgEX
UcuSlAHuqnMIE/cH1I7MeVocGWccSM6/61YxLvYWVnpSaDZsUpL1VHVBgJ/s
xfxPte3Ifl0rYYOJ8vKgVOfKcPvQQGc8rHHtAi9MtmSoQRzlhVE4HOO+cb3/
WfF4JgU0k5qpzn76euhNQtcWLv8lfhYY/Qwzys0DdW1K8p5rCy0vl+LaQwVs
ZzH86R86t6i8KLR8Fcz8KKv2sU43YIwc++nXv4Pg5AsRGCU9+3YVcTgtUVbQ
NzhdOc+m7vzMzrPuCrAkO2VAQSmwRHKeFmmRl7LTy1sTRFD1EDAHz09MS/fm
OqdePda20r4SbOkJ0yas5k9ZGSy7vsSnjYZCpkkhQDAofS8Tw8Jy4Q6h8Iuk
NshLU0FlDyq9dfH99JLakzYsc+kqNhLGpsANxlMXQbc3zNJYvwdZ2rClWicP
RGLILMTIBWpn7+cr9D7GYI9ijK2DGqnwCmZMLazyRtBud9trrpbvK2pYNN3O
pApFvSFxregh/OgSwSn+n8H2ztvM2qxdVk41xTyD+oalZv8T6JhXHo3vBgzn
ecojGqd7FXcjVOTScWPEj7KxupS4BLNqpqQzpuX/Jkmf9oD2VHBfpSp7Buh4
io8kFwU032u+J0Y9Vp4YTF2KQmnRHKX76fTbZ/cwv2G7ctCYRv6hib4Zgkgn
FlEcGdd5jahd7h1WV4dKTQGU9YN6nNTQOXh1jbdOQ+G7u9p/ErXk4Ka3tYW5
7qyQc3cb1nMOPZJYE+UUpuwsglIJ+Q6EREXc21ouJ+HYOvbs555DsYQr0R8W
iBhdwE+QPLCXdMsZ1B2ehZUKSWl0KWm6HIVZhaOs0r90V87kUXm7lc7rB/DV
u3xIhVbkvv6IA25yzxpNxnoP/z2IEpbyN/rMvTMtAMzIRH141vnr8KQJHWbf
47IWBAGU2TksSnSYWk+Qj9dzWncygOA2w6dQ58BSa/ZreAkvWtMsbiIWRDWQ
nyUTX4UOgurBl4bLUp4k3yMGDMh9ib3eIFPZXOXpMJStJqbXWLRh++CSRxh5
BdH6amrfNrYbvzuZbzI3z9ypZrRXXf3tmxM1KakiJDI5MDYxAm3e82bB4uvL
hWsAozciZ+2GifUzOaSQL4HfJ3gE/becqTmI2hrQhhECk9cxuupjvItFarzO
EffNxO2w3wRItlTud8fugL3+gEy9Tei5oi2HuW6Tigngq43QGcn5qX+koC6D
Lq7XE+t87obGji2em9BoU3qyLp3G2FGwJzh95TTBUHvDNKl7J4IcHMhrZixZ
jGr7DDclETHPnzMMoLm0D7Jt7ISOD1vPNFXwSFf39L9BqC/i/HcoWAPhQc6M
r5016p68QQ1R3e5PqSuDkoU8Ugjo/f7IsOBC2IM4aCsyZuLMYC4fwLDewvZY
COQXiq9HIkMD1Lo5t1Ch9Je6x78BLXqo44UBUglbEMQZUOFGWKF9TUTZQ/jr
ywm+Nk3EAcnPGqbTzapvF7DmRKwf3y8dNRAb99006Mrn/rvXHCFdrCX8nTYC
RG77dj0BOUjXYCYTtfH82QhMu0Pst4DHtSDsK/9Xs3ONrdEj3RA8S+21Qzu/
qf6a96UA2o+/xUM7W/uRHdIuBS2eiIqIIWJmAL1PiiJ2T7leAj/es69HQwhB
q0Q+fkXoKkbWn/KB102/y75MH4u7CEpomf0DUpCfdz8fPgx1d17Wuu//rt9m
ue7L8e4KFPqD2MA1yZM1Y9VIToMs4I6/RaRPgWcIBiwGqpzZTW2a/4NcTDC2
G8erJDzup3kMuQm6H/92ywRkH+xYFGC/kNOpVmNFGdRYqmQLyx0n+iJcw+LW
haUJjf+DGILzSIzPYOcSKsf6Au0FAfVc7o9Zim8zbjx0xw+1z/2Ii1rar345
eF4EMxdFLhF0zNaxUuMRJKNQo1zjpWAASR28z7ka1jaD1GFWUdCk894JQSHQ
b3zUmxgetYInYKXM7zKr/kXjFVSTniYF7bdShBOc0NJ26JrZjdvJfAMqUoYS
6ZeU0v7CM3cFDq0YhrBMvxC2Jxl28S3k1O31A2Wt+mX18i5OXOs9kfZLa3sf
1N1Quaw77TjjmxESnYHWbgzZAKw4UbK2NvH6/L9mKgZ4xLIO4tw0VV7pFlK7
ZEVNA7sGH7Ef2auyJrcFio5yc5aL9GDW5BwQjLfcY7L90FFddkpyDCBKIhq7
Dsy7D5DKx/xL8eFrVBXvu0UZ546f36jG6/JHpkw2OpYxgBgYkUM/KIO3nDPF
YDQAHCgWBlOMiBWu19sdBSv7VDJbNzzUNmT2A/AROQ5t0Eahx+MZR07Q3Bxr
le5EvZoddP2EPf9kejDQoqlKdR+UjN9fJvoz2l+Idk0X/KdUOESmej20AK38
p+g6YkdTFF54rp/eDomwpQbKmgbIZwytxVIdtLN3V1VEQtxs8R1wuvHE/zRG
cDuO+cHPsDQdbKHYr8pIdj798nknyZhIQy2+kANOQ6Ic/bETrQ68WZbCZw0I
2RtbrG9sCCzlgCF/g1wpdQorW1ufIyDLdv2BoxUubatx7eRmtRYYZiUjTQUd
WjtsXuE5Hyou7rJa0NbZMC634UUHZsvq4iAnm4+htFvu8XmoPvkSiHYVectd
7WaeXYEo9uZzRnaXKcQUu0hcHsuz1A3/KriDoBroHQwDJgA3MvYuBVuvWms1
kzCacFGTpDbkxh9Hpv/olWQcpdtG7mSpqCR9p6EyQ34TpjBCQ/QaBKWFiuvE
1060uci1ARdogyLyB7NFY9XgVcCDEersAkmIDxxr8oUzrJv0Rp6RbWeY7WY6
w24gacSq5FNHx8cmq3Em+1fLDTZqkNl7m83AVWtkUjLe1CsKMRceJy91haVE
Nk9uiY3VR7/3X9qs5qGrTijiI6SURw0CXCgrs9VtyKPjh9se05pNTIzsGf/L
r2/u3+s1NFnus0pg/3SKVvS1re3kc800iJiU5srC5RMxNnz4vQDJBXzcDNEM
TTAKkheCZiXHoZxJJ9DiMK7n25kTBlHDf+B1EobWl4FlhC8npn6/OSd3sa/w
mynrWo8+7u0X4TDTpS8b8lzCDGsmOroRwspoLVNr4XKytCEvgbtQaO+i5LkG
WMlcO5VnUUmIWXpamkRxYJAcgaJubn0ttQ9pAt+bE3lcLEMfJ+zJsMHretXB
sar4/QVkYldNo/ceHnVR5HXmzpgrl9X2efc8xlSclCqvJa4wDEWN0rKTsigs
kw3nn+vj5xNrbGOHnCwrc9exZqocUj/mTxPq8Td+u1HwDP4fcjtpzPX/Yfts
s/1mS7hR+EVKSAQ7DPfBSJzXjsSyaGWON7LTb4iUhAFEx54aO6r9bmwmNZhi
5SQlu/enpdPmd9xow1x/Uer0sOTM9wntL26gE1pKxM/0G+EAakUVdPC0ssec
/Z0xKv4oV78QJmDSnB5lV4op1iZKqSM3oPH4VHlLmA0MIUv/Z579LdxcHrLX
zmEkbVko75j/hC3BVrfNpuhVsflcw4OZJllRt9i2c4FdNjlYPGxL9Jrkd8xW
aiCFZbgjNAKFI0q7GzQ+VQrjW1HRUBMbBrUKySpmRKVqvXj7Gsc/6XBzfaRL
FGgZ5cQgCxrkQHZoBS2dDZ/Ln6hNmUsot2DJehMbZlxGfg0xnMPXSMDuLy3P
AG982JBhsrStx6O3yLGx1mKcuHJ5i3++LOTkAOB1I+zMkZcN0WdCbpSi6JQi
fWvtQPs7OovXSxxzZdVa/SALybsGfZzGLA7SFYu5Nc7mup50O2XDQM3dXKNM
g3xWwrBu6vK1kV4yR9o6VR7ZnwUMgffp8JW2nPgiYplDsSyujtW7J0Stfiun
wTIlQeikNHkShRCtIhJ0jIdClU9vXTmT22FrTCKKXXCatKBsqHRrAkne5ECR
QSmk/OAFLFSKLl/Sdi+LCHryMyZljbqv4gRWenwLPRMrE4G4W+gYQ0lfPIs3
MmFmmTNXoDFh6rqDjUlVRPEMHeuKS1cWcNbna29CwDYhCR+CX0zbHgP2ilVb
d/pwqTFyEEgkrvGzqRWBD6GAINl0fb5KAjAg5er4JjfsKIdJkLZ2ujgIlg8g
ne99WHrF4+Sx9Bztml9dmTEFMuAk3t4O1R3OKJGJC/Vtw5/2dcmx2w6Y1WsT
z4seQg6U6059JzJLai8CSfMnGpTzMSANODR18n/XbP6QrnFO2lCVVWuiGiPd
+ZaaIALaxgY8QPaNw/YyKTjQo5o2taMBuf2yVsMgoAUiTJF0NOViL71BSA/I
MEUYa1arSMcTtmYDGhEHN184/MwJiIKC3ZasdQh1bFUIUlktFhpF7aqxHHpG
lRRK5umn749CLRyr6hp+9EQbVvaUMjojj4u3hyknLNw6Hkk2vNzuvADR0kj7
bHPaqI2rg8R7OfodsOEj4iH+Pwq2VU+3Zdo3SUfCPyZDZUkQg9x5GItzyDJ8
XI5AIAP9+LVF6Z1tUWFGnitCU6SuTNYMpSpf+YjOkRwBJRESrbSsQ1/aJvZO
A7p3mlDGjFvOPwIVMUY+cVsx1cDUjv39FM3oWytcHWyJUyRseQAZJ67in1z1
2mAnja0V+t15rddmi6DwcjF1AZHeRSxPQw7Sg07gDZfp4nsiy5QkiHHTAW8g
/khEgo4oAn7kiWEWXzpAaFmRJ10RBO8vqqT5/F16zj8p7MY/VbdLvpJvfnof
yeqisNc1ubnVj6vumHEzUoYsOIbOg20MLNl+O1mJoHBf3lUX33r1HTup8i5O
j2PmlRyakFi3JW0idSqsNTIsKsDkG0shziaiGTtS6MSv42M5AefcA36bOyub
Z4tgK6ABgCq05brDvfMPFlfncLHiiBHdANmx6XHR67gtEBDMGSvwZv3ywmjY
KyPE+Cx1oBPkhWf0pn/bUITm6Z0jDPZu27iYlQx+jqIqjYe6ET/MYC8iF1kp
5Enz5fEJf0jUzPx9o8uhrDW5XRW2YkYPJFj8sUURPXNkisrETFFaEWfI5egF
HjOdC4EqSoy0IXUBm2wgkEX6CtibOlM3vAhdGIyoB2xPt/MjYwF8AtzNNW4L
IWRPwskXK/btFYfxvMYEcUQ3EpfCfhdrIKbSX6hyIL+3EdyxRfrL5yoZEAHp
BW2+6M/b/6V7/JV/fNqllD3ptymWiM+28GRKLwld7dSNU6bv3rif+73ALICa
PK4+TrwerQ4JZGwPavljAClZw6a2dXK3OgHWyD+5lumMug1H0ND2kSw9WMll
LOMiqys3kAF47vEdhrcUpXIX7FK39GoqkJ3sVDeBfdkt4qER2YJv7pc+E6ui
U9Fpfen0eyJLGYZrgFhOEvS9KYfsSz643EY+/V2+iAKf2DOkfl2QGcvSbmcc
Uqh2NsaXusYOxI2xrRoJKrmeT228ga7BmTJHiRtR3aZd5Sm7mudSi8gr0uiV
m2VKL6nZ7c4/NY1zPhfrSOzZyfjzRE5EfQnoA0vCmev5jliN71RTIvySZoj+
3G4qbSm+M8n0P8vvf1WlRiNeAU/szf8z5o9G2EWFFkexkSvOpsraATb2tZbV
d6hv471VHxLZiAB+MkJFuFuKI6EtxHaqoKBRodMfWPLxPIhDL7U2QSh4LmAz
SWHHH7//nSHQ4b79By/isbMVS1We+rd6KARhetvdvz/Z9wCtMu7D0Fs4ZQ/U
JJleJCfc6aJ53tOEhAnfrIZ03IbLjz4NbY16SuNhmq1ukJUlcifXMZadQoaa
vKuyGq6eLx7VcGjorR/vIv6sDET9Mpc6Yy1rg5xi2cBAB0eQZC9RWI3t14Vd
KWDBYv1vhRlTUhefjM30tR1oq/538IxzjSrsgOlX6HDqzqBtoV8XyX/XLsop
RGCnw/7YOwZcUbzkmSNLXgFRMzUCJWxZz8YFEuJyTm4jXxIovrjJ+ooIWCjR
G1aSkHYzwxpI6/8Us06NWCZPOa8VSJ7eGGZwwiq9i5s1JZSIjPOpku/Eusbl
PRZm4HzIEbFpuTstqND02i0KWVRtDY/NRhUaYD2rtHmnwPbyj3/LlD74AzFl
xcIIvg/U0bH9nJ8z2MjgpRS7JP2KNZwAhBiQwltZRRd7+z/4w1FchfoPJdom
XDaXERWY6TyGmvm9rQKehqzlGWNOIPQUvlrH14fCAKzeHRRWDJGR8Tw3ljen
VJWzV2gx7TmL8JUOvH1GiepvuOwmvyBFWQoX40Q3ht8SkiZWt04k37QJxyVr
pjAV7kMSSf4IkUwnzg7ndsuk0dLlJhv4e9lE/JTj9+GVVjRq/nFMxslictJm
JXNxJvAxdsYvDkQsuMqP85qmaQP8bCz3lSP748vMUlcHgqSpKBqVeMYXCx0r
VFydZG6I3faIxbYBoYqVD+1TArPQIyBFdf3FRnuN33AAyUUSoYD+M8gEBc4x
1cuNccSqkbVWGyhEeC3bxx6BqJAaPR5Y/svHWPyUb0PEQmTq/jzfOD6nW8bd
iD8AwcJ7orQZijEbN3nlB6OX0KbMRzg4u5oUX2rt817LpOQvR16pwGVodvME
pVXcYviiH4IMIMLcncGJOvndz8kZEtGWO9eUQOX0x8yfVp9v4Jhp6CBs/aaJ
wi1Yyth8F377cfG4bG2XN3/+pBQ+lDYOq67fz+M83Gf2W1gGEcswGhB1yJSA
8ImwbaodHw82e65MbOf0C+UutjEqa6PzLzSUxzDtcaMw0O1aNqYwEE2RCEQs
mQeZHb1r67yHYSlye8Oe75j8k0xwBTjRwmW9MVIsmfN417WELpESBx8NqskZ
18lgnOZr3wA9lKtFNL6Dk7gzGZ4mxEbyxvwLF2ejU6y5wVtBHmjRfofwwz37
zpjRsm9+KHmCLJuAD+GK/u0Wpou1ZriqHPsazXfMlyNEAfLiQrEjkAE7bi31
45EfonEVGd5Vf0fXeQfegzYn4LghMS+nl3pu8k/83WZr6JFV2MFzUlLLrv2M
mgi5sH99peRRC70E5UyW5t+XPO7uFidt+8DA+AHNGfJwS/c6ZFTK0uuDBk4i
pIcdWAPeRwgPzt26B10Lnt6fdtyH83Uq0xdyiLQ0yw8xF3XUVILnRV68M8HL
3Vf9d9mp0yYRJ8wol+Hhpib7HoUPw/irD3hUrrjKVDo2eg2h6vB2ZpJd5Ee4
d9qKxuQJyScUIFggdCpydWVMDmKvmLe3hA1izVhsZQjsYxtaWaOXRCRlUdVK
35e0IeYQPVhgm3DpjYc7mYX00+5dOQLRqAYH7ooP3C8FQWQ3crobD8Ui+y9Q
uZz0W15mNUBiUNf2aCy0JDrVo20dqt8h5GxvLHpxzLkgfKjRTLZ5/9VTYM6l
u2XjjAlNU+pO8KfrOzLeKiCrid0WoTGyq2yCtXVtz6dez4TkG/CH0UFkdpMy
wxrOUTWnpUawF/u8LNtrcvhWiuJqenXCW983XPiYYHYgehx0HfzftHet/fej
/Maeh4qd37Vf25p6ttJFsW3STPVUTOog+yZLpR0RFa9e2QO5lUvdBGERmk6o
0qqNva/0oc0gZKV8FGgLM4XUF+9mL1iry2urjxqWaxA2JX/rtO8JjRWQ4Psc
owixpIoaaLLGTFnNOzlG6HYaveItXXyGkQkBOu1tnjp4BuFMDOf9GqXtRRrf
Mx8Oa37Lh85KCjOrZpp51HaWU8lzwkWc5cCYEIe2csLn38aEfiEJhRHWAjZv
05RbLN7NUvGOIDML0/skhY6XuerJMrzj4fn4uKEjr0cGOHsLVj5SQKHmVgWq
ulbBsT1r7bU7gFNFStg2oKwe8ccdAQg2n8aEoZ3GGKi2Wsofs12LaHw25QbW
OTGuy0KamDcu2u4c8DEHrJS2PW4+PsJG5EuGe/88Q8cSkv4115tUQUQ1GQJp
FLD2TCz17FOGu3724ePIxsSYVlwtdum3PMyqqZvw84f3Z7hFWOTi76st4hy8
sHoNEQqoukKiCxJkW/CYXiartrJcWKO9dGPz7VFt9pfKfBRsn28cDvXzDz0+
OXMYzHDSlrLwpqTo1+XoTRHS/yRlj1dZ3uBYpRRw6OCqugaBYxmNbKQRuGnP
RWEKLsWasYE6rB0HvRI5pqQI2KLBiHKvjEzX34RhQnmZGeD9NLV9TXEkgvtX
cRoCchlgXqy3o9cevGjiiDaVaoMgLXbL7j4b/hcIJHvkqaCVEweTA6zAocfr
iQNpWzUC8LmXqTI7onyAf3l4Cl0zwhCo6lEO2o3W8qn/BGzz9Z/WhJl4CTYZ
aS5yKgLqScU1YqwBClNO6Hv1n+Y6AOY1YuRk0sWr24M71nUHli/d9VKbdTCP
qQKuNTnm0uIpu1bzC8N01raehrx9+m14obTtorwJK5qhJ2TxzouNsHwfcK6B
Ic+5fwiBnLc7iKiGel+Cf/1feyATKlMNlKb8qe/nXv+kfzi0ALDBjiwCnikY
w+A9O48ekm3XbY98paSYKRs1KvegmKTwRW8hH5PH7TPfxKYSfF2pboVfRa1g
YIs84YbCbymD+58LXXHDifNYt2NBLWIfX9vJQ8VRr7rVBcURh4AQJ30+UHTB
DLN6fcrZt5PTuWu/v5co0us98tz6WpB/SKYO8owtd0m6pUTeoEMg+mrK8Y6u
REV6Jzx6klBdhFb4uFx0otdTE6CybGqeN5k5ONz6WaYwn6z9X57Wyyyz4aVs
keMBZMwQ1fSN51CzqisaLmagkNI6d3opgLVGV058RON+4JFzOEYW918tXNSS
+jpOZpvUO6444FuBzO1nnwGMoVGcLa75+q++7ICeToWTBRTi+YTJTZ+TEHs+
Hs+9im/r7Prtokhn4RIkwKVY2NlQFPX2PakMCol0A0kgzyn9qPHMMi9ixZmM
gA4Do+XX4w8yba/UyTacDaxRB+3YYh0fZTtyeK6U+U8edo7Jmc23DvAiTCHd
tmlnwD3Xj+eReqiZ5xbqI1HXymfAuKlcD3iccxlTlEAWZSeb7QMBCP8TVEBb
TvwkRfQsFlyvdJx0rxJB8d3WM1ENOZtrT3/elsPRnOHMlbhECqw/3JDyCna/
6pMbEWx0oNpe6q9tW8xkPkhlNTUWiBsvVfrXtmCBMtuzx9JirBO9FVB9Tvel
dAb6qzI9xkFO1Ztr2xPIHWeRYD5vqkQQiWe3EADsxGm6MxWSuwnLJzUktNVV
PcJZYXsgX+DSEPuEKVWu2SjwxizFWt5+ik4HkWd96RWDIX/QYW2K1FjpL+7H
q+eH5dDfRVWpt7wvoWU7SD9tHIs/zZJOCiHyevRgMBkp1A8SfwtsSJ3BFVJ3
s9tGqRsh0yn21qgPAzbCaL/VXBIbADYHn5C8kCr6hCMI26yJOCYrCrNc+keU
g1Zp0pKKboVUNIy3KRzUQDBsKliNwr/wmAhmoPY0/W8MFQYcDMc6cq9GKmYg
inYug3mSNJWR68jW9LPAMtWfOAIDstdEe9p097nhZenALuvC51I5OEd1kTY1
4w1UJxiaUiEzQDMtDPhTnON8CkFYAB1lbE53DWQUEaOi1b6NDUZSc5qa0KOM
V4MqWde3W4RQgSAIdL5XI+YB6VzMAHgLLaLkdAGNrBKj2hZYEXTDaq14PKdE
+M5Yr8WpBmW1BFOZtMiNwM5dxJDv2S1DQ4nebx3CMr7kPcadWty/A3bDrqUe
gcBg62OtjODEtj0jPHRTxGqIjXYpHZTJs8t5I/hBjbv86IhL9R4scpxFGBEs
/yUM1TQEcMgHw8xEJpptiwZTW7LwH43TjCjXD39KEWaMmoBzb/s0+l8MmlQ5
ahHms4w+765HyPcCgDF+YQ+FnQ5onBVA27guKy4CPLRevJ0oXMx6k4J147M0
XE84hFw3N6LuehTfKp2qtMwgcxUUDWmQyI9xeGmtC8O8ChkfX90z9hEXXlsD
eibX+Px+9gm6HeLM54ghziki5G+IXlWBAhOOGNrrzp73y/V9yeQcySDOV3e4
lYS30qax9z90BBn6TCqFBxpllsQ56p4baZOGgQeSY8X9rzLwF6tJmlZrR4FM
nt+yKkgJQrkMT2ld6d4HKKXXPW7NYdBNVpr3nzQToWW4s/4NZCi+oEkFTxSM
XFdIK08u72gCqavrnoRl6/JiXrzc9+F0fyHK0fNSvP8i2qeZEFlkdm8aYsT3
ZCJeAQl340ncOoM76BbUItk63IDKnEyzqf4n2BHQoV4qZZTnLzHiHtSRdoV6
CqsvcrjWY1RuZ8orfU+ZfMlH0nfhL/VxCBV8VmUJmQEKmpJajtSLxxq+ot1i
prmlKuixg9WQd/u6a7htZkqLbtxWEaRAX+NWi73yb4bJKGjYAuKTnauP3Zef
4QXwl80w/UW3dglqTlV1moK2Ip08CmBWacCut/gBTomhYznC8/y4rOQ3dfv8
HhUJLDTwUeQJW4wbsJvp7IzhdJ0k+pEvzw+ve2MLJZJ5ayya5Qkk3BTxI5aj
9sOki7ijbDGY2xYSAyPv470clkSvg/l02VnWRKvFLpjTKVF//LR2DuOFvZL3
SHO56v8HrVVg

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EptFedWyycaFZ+NcNvurMTCFIcbW/wqM0JkNNfMQZYD/epCQSWl6VmXAhjDZ/5Kwgsbq+DG1sQI1uMSl6bbcejXmTDO0ft8/GhXQQFD8TszePKbu746bT4uyZ2m5PWIm2Zcv9eDvIsouz3gaHxaq+8ISdWD8apaJp9i+sPAeiD5BqdMkPkvctkortIYgx9pp9Gq9vV+csETfNzacplu7+cxPcLhMsj5qZZSNvxtjRKOqm9dw86SyY/b7yYd4VlLcsTuJbFsEg0uj4jrw7BsqOXYgvxYXZeP5YO67U73+PAA6KIjj6eAQu4LJEAZavvG4UGjc4/vsqnnbFbf/4dunYKlwoATuOtXHpabeusAiXqF0Qt1VnWtZQ/L8MNY2sUJdKxkHU5jP2z30DESYsjzrA51L6T1bkvqb11ghRLwMWtiLzbmSW+ReuMTEk5wbJXd9N/H4G4BmUT9volQ2xqGjvXGfmEh/AiY1cvsJxXb3ogoT1oGDVaSSqdSxMqZHifvZyemt/gy1rdUdYhbATVuBi80m2TSo/Pfk2UlI9wB34MPd4Nk6wBjOLf8ctFwXmoT3IKxJdmwlu8V42xztfbGtWMhgS7UDDTL9EsOp83hlhWrdvi9CF899t/i7DHHHJBdg8Zg7V9p4h+FUAUccwEfpZGHr3bNRYJx3yyM8G0duYNozb693wupz2TtpK2SZskI799BNL/c8gcPswZPeeMzkb207ivK3+IrvGSo0xzYFXey8as2itcQ3RZWahWM2GF01qRxb83U1U/IhYrigWhwE41d"
`endif