// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
yeUOJ2ErSfNIGSQd3Zbxx/p2yrBVie2VD30vUsiuyj88naa+UqDr0Gm8SC9v
ZeeMWDRShIq4p7RAFfl7SHvvXwy2sT2SKWEBOcujTmpwd/J2+CXd5iTq5731
9LvsCnATQ/zlkgTELSjbi1P8i+3Mwtu9sdiRvI7vHecrpI+HXu5q2EJaxAQW
Ni3unHMapwCdgEx/ctThv1wPZwD8R5MFB+5ULR8GvNa1omaL9MRdecG8WRCP
rIMhfFXGOAlKLXIhTnq2XVkWRBpWGOsSy4nNYBXhHJC5tlTz+ZwFfQmCZKOP
n+fyA+t/Ev69pHa+OWcXrBLhd6zxPxaqjeQfmcWksQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OWhwxVSjU5mnwjHpm1OkNZ8f9riGPFu3mRln43Eus+gHIqr1VeIjATGVm6UK
k4byz2ugCxqVZOsqE7nege4aDDNIU2PLZ/0Qphd9JVMr4t457LbQozZn93YB
QU2PykY+cHyeYzYhULohw15xKgvx25KQ1M7+bRfNjZpaCnmNuepsDyQoTD8n
nC7XUz1rZ5O6oYfmkwZiogTd3/IvQg4I6vonFpG/MrwvTKthMlVef0PCvo5n
2zzban07Of61+8BCeDgpHSgXI6k1LSqDVWePqe3kopW0qwKgcoiFxK5OuN0J
myfyneuwr4E8jnQXT3JlN3fRPDER+l3v0D8T45daZQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dECP+dD7QDAEsOOzG8oyrQrr68rFqUz3Wlokx3VLcD3Ytgn+EHuSJZ2bCfbM
IVnvitN/Gb8ntxPzayMJNJ5zJJdiA/bJPAbvVY8eWmfnJmGGUQEj1XNgpvE9
Rx5sJhsNHHu3Ub2J8jXYjNwwNbLUhE+OHw2zCuT3GSf6TtNeFJED1HB/KtGQ
+LpNuQLQrbsA9XU9ZEP3CG2eGCfqYosNCll41qZL+ccw0D5FsQ2j+ORkpVlG
tBSm675aidhZRFkX5nRhZHoJvPrsaMKgyz367mW/OOkKp0wJQ5ox0cJ6WzOx
9oIsdKkfEV2HXnZJm3MdxxywkSAcuwMFAmXGtwlL5w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
odqn1d36mqua78AGfRiOtSfOJb/mGQ4nzaDROEq0sRKt+TOdxYEEFUNZqn+B
nc/xNVHzfNkeKwlKCSJs+nqUpJOs++yFNDHkrmAjXimCZYAdYw4e5ZFFr/Pv
Ym5aecjvjX0+YCYHKOyZSze/PNqI1CORlFI0PJ0cwIWPDTdaJ+avjQI0p2Yp
2soQROYBT0ew6dVfrp+WEhfm5S/03fJogMJqjr7bZODzJBEwf8z4oenj65C/
ScycGWDotN5i9Rm9gb1fnUfoXhfLQ8RrvFmCJGdVWdLKf+tu+Qg8eGsaIqHn
FstDA0zXWhJYb/1BxW6F2e2XzTasAqQ9Z3Zh0lKa4Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CASq45CKr8enTy4DV8SXigqbjC997of+ytvdY+98I6J+yK8b52sDcdDyFh6z
AhOI0VWN9qWUulqD26OXNtbUA32HIZ0971w6++8BAl3GSSyQse+mjVgp9zaC
hLS6DD/mzB6JN10sGJIG9VSTyRFl/TWLoOphakxiBO60mIhuQzU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uSYZmuEKMk69lnfEfrJY7gEZUxLXMJWnONCP0IkA+u6l+MtA1eUYSHRMG504
a9iPlIcfxC9y1EKUFf8QyMQKXTdBk6/A3BekiUtplMumaZBiqCkMfrYNAc6E
UlBNajuQdn4OCLHEIHLAnYVeEoAwIRXT9cYo8ULplp/LFMT+cyI/ukpjnC/u
rHhEyGivlO17ChujE0BFrma3By+tB68VPW+inAygZkqrICpV1E7U6QBtQN34
iNvuNFUsWgf//NqugaL3TiRMGYC1PAPyHn40W0ycYe61Vgy3EsEpQRH9mvBG
zwtrEIgZi3pFPn3kTBa/Hp/t+JU6JXn4x0dNE61RViwuJaaihFYWlWS5S4VF
UH4Yif3QUlBZ9SMN9+YywEhJuV+nvLktyWYGejyWljn6GfSLcf/plUWE9D9N
ngpwmUVB0IvQDuZQthlehY1rtKMJboO4gopmhCB0JkjijP7BKccGvBmr8IrU
ig6d5aCuJvVJraSZtHve3cR+s4M3GVzV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kq+/635ddWUT/Cb9Ppn+3B4IZ3zcs3CHQX/eNlFPrMOjLq81bUlN/A7jJaVu
7SR4HXa/AE6C+vmD570/s8jd07y74fkzf8pt8G51FBTxEgt5UzOIzUVnQ5FB
jwJkq4/qHgGy77ToHNe6VH3tF5k9+PaN6xaxD6Y5XrUQNn7BqAc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e/59LxAiDjR2zvCsMVTXF/0DSNvMICwrg0DVE8XpKvv2GUFOBr0QmcEFNQh9
gHIA6TvUoODy2zpdVwXkrS9ylkS5AimQscWZ+xLFBNDYjNjpdct7aMf5jTHG
AAAEuG1XJd+mrvHOZElkpPE+53MAtLgcuVdq7gqS9i4zeen2czI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4736)
`pragma protect data_block
ApaeFdUfJhBzvZMCJghXe4ozuwVyiu4hEmcZ0t4zikMVEMzbL3MEqCJ+P/oZ
ar2dDmSWn30hAuh2Peg5aessIDsOOu6RNWnq8EsQmo0rpxuGSVhheG2TaI7G
IkVh94cudS3AQRYr0yR72evdE8e8Gf7ljgnxpVysFTGoCAclJQ4qCIA2rCB0
uEe7LKI+t8UXi5oRmrMetJI8Rmf3goGwl/DuxPfXGIAVgHRTIIwCYw1jjXcn
P3MqFz5Eo4FK5f2x6DOgPwjQVuuBKVSpnUcIBp34wF9qvOH+YkmzP1XaLCP4
bVBJXub5tHaIQO2srjOdd9FMwGSRCp4aNtTviSFwP+dplCFyEvWFkd7xEBI1
GCWMVA8+ITMdbGm8itI2hiItqxq4zcucMhbmb0FKsktJDl3+q9QeyIO6jwa+
rkEXfji41ngPdZbcSMIHrPteNI/jPDHOo2hu07rhnsexjxBW28gezOlfR3Zo
94UzvhjgZFIKJlIWTBV09mk1uwH+19MxqSRMoDGlGrt82Vt7X/xeew/epUvq
VWt42rYDeKLzxOHStHyEHIJ9POCBeLGJ5FlO0X181O72kLNlw8RGzAWRYk1G
+I3JuEaoRPjwtMRSFrm+XGiVkaREH+sWQDIKS7mEjkw9JTprtno+dNhFtw9Y
9j4Rqggu0nZRVieJzRbr5Zfx3t51rtNnfVJgLcVOmQ8y574wz7piyTXUtY6I
0bLM2IRhofzf8+ZmZ/zlwXoSWYKIO3yXl/5Xr+/7uSSF/ibmoJFrijuVEGDu
P0tILhaz6KkQnZedb3I0yHIYuxG8j8/4VnQObJPXrzuLsHRcBzM7vlkGUhJe
kowFMwN9kC2Xgk/0vO/GlDvfi9RsYwt3K3ztO8NnTJyf/zOhhB/QSTrVK1xX
YWNHR8eYb+FLEDqFe1jd1rBdev7bHszg91eoAIvS9YIM90aekB09GfECd22k
zWJHlrKbKsSmHq5TQUi4vCtoA/fJMNqdS276qI8h9J5PS3v9AsXAaH6ecQZh
mhxa9hfuMJj0Z1bkDcQuwL4DL8WK83nYdR5fZVdTXXGfdN9XOIzlY/nz2i1A
WB17YbXkMiLxYRdWuONWDmRfzcdQ2mUbRm/lysYzwQMy7gr5NxzF8l7eIurl
/Lt6L91BCXmfy57twFPl9pmgKwXuYuaRzu48DTkUztFZnYeQeELmrzuUlFEm
+xZu3JRlY3z8ewpvn0pC4Rsq6OUquwdCWxpecKyCMqt56UiBcj6i7VCB6tMr
bPadJa5FZH599V1lg9QeKr308+8qIz2vUX5/NbOTUadY1NyGY58bRIWrc87A
DD2upEA7tDC4L6xBuyMBGGBVnnWdl0Hy1i1yW0QOlVNB29SXaUewAGtmv78I
y39+WxqY5u/aa8YFF7JtJsu3ganfZEv60ErZiHl5mQlUmFsXgvn+tS4hPSIg
lAQ0OFK25z1QSzR6ReVR9SSqN481isaebCd9Npsa2bwE2jgbhiQn4/mQxA/x
LH/eY7CF1YaoJesT0yrMlrGEOye8EATyHbdd5Grfix7jK+iYF8e+wKfIfAYe
TOugtrMT6I06mc+6uoE/F8uhHJ4NNNasY5BcKK85lxxF99ahG2kLdXUXSbJM
+rWtexVKEeX5b7ACCOGtgf7A2gTyT6MCkq1tHaWYXZ9vDfT3z1cMuyKHK6UE
GFwT6O3xdiV+VgTHTiSoWtnV50zzuD7reY0/x2xdzk99bTGuN1E5UBJJMnk/
F5b7+shalDX+1qyiY54GFh3r6W/C4OwlnhWQJmmgiEo3HVNVF176pE/U9sO4
vRalSM+9+qVf6d3Fgo0iL/nQwtYC21RLDptNyiBu4PFp449PImdnGqAcc1KP
m6SQL0vRHBiC0KwD5Sh0ui5D9NcpFAVH8IuleObdSjI3jWDw4kK5FxG2Fddo
pzinSQPTWFFmmbkN9cMOcxSZIoxgRX2md5l7W1Jr7mge7Wh6cApVzP6S8Qxj
z+qmUUjCMbeO03P3xX1nsdxBFrBCVB6tdYE0f15oUQLStOl8H5cuhYZdaq+S
tEqT0XTwJ+Tr8v5GQ1cDd3P/P41s+oRN6sLIigz0uR8GiDnSWLXr1tAXIg6v
/mwRY3vmYh4mB4QihWMUrMCh2Jk4uRDVxmq/udw2dRlQrAdxKlliCXkHiBJp
svDUdxqxrjhPfN96jpd0xlF/9U2tT3ESZVxgKMNqRhD9S00IgKnNkjZRyZsL
4PishHgiX4ixOVpDA2jK5yTodexqqw+qlsl0dOVFbcJL7S4HuCDhKnpVOQvf
H5mVUDa3m5v0PyTSaF2rFLThsNcOq7KIWxgwKQiqcktXGWgkvUG/YGpvVLta
PtdUeQNSJPZn1Wux5ld1Rh5697+vw9ZiEiX1HtSaSGRcz0bnfJplh31rFjGf
ubk3SPYB8KE22xy8HwREvc4/mxyshF0JFW7zrOiezVGlW6PHw8yrJXw4UgJa
VVeURVJcqkzXBacy4uS0e9abeQOiZ94pfjpIJdspoqp0WCh+l9T5wNR5kOeC
RH+LC7kHUK7AmnQACptzlLNYvpIK1tiS3390gPl9BRFwpT6pooM26h3GJGdz
UlsUj8oZooFDn6n5RPnRozLzYDyIsfuHuPlS4YsDRJDXJX/p2729RSj8fG7P
uEI/3k8WKgHrZZE/ZadQdVb3o8H8YF0aid+o7SeDb82yY0YXkqth/6/ETGsu
641aTeutsZwAPPmVaXcyTEo5/dZusjRn8vR3j9g3lMfUA4PXvDxtFTWSm9tQ
Of2iunQbQVFF6/Bhq1Btn55raD23wyUaC+GVZyFcucI4BLfk3cxGNveJhmTC
UH+ItHncKXfFVQMfMk00l5Cl1Zl8CIwOTqVXrvuRk9wss9AjS/+KmcCc1zTq
/G+ZpUwqfht/Ukw4ouEnq473wnYDWa1Mi/fekzFVNbMFYVAOIkgTobl5RHwC
H+QwFXv/T3stg3rXeuri3XsBNZru1GfgH0Fz8srhH0Wlez62SV3rF62RnJc9
nWzPXNrIIZz/uSwl34dCfhCtcpIgrKTgAIImLpBD+tUZT4UeIQWPBtCJL+2g
NepByy9EtEORqVI5F3iAI0RGtMOMZvROAytUsiAiCfy3obXRW0hViRuVUCMI
SmusMWbCbBSkoMaZYnDFBKM6ce7GcMb9Dqmg7ibOpdvBhGjy3BO2DodtDlD1
et8pkquoG/W9EAjHvSk5i2IqDDtCtCtmCTY0z8p0oDVdx5vabnGU+4nkmisx
Fp2z7vIp7C8kpRSKuUuhzT8cgCQheEQxbJWGrpCsDW8QLhd/GI+Zam9Y60/f
1+ePuscPCyAwHHGWBVbkVlBX+wnQiAevPeye8BSwivrlUpQTOMhfEqFqpMvq
wtT40dAsXXZ6Is5AwpH1yrfUuq9ifDA3s7uIcg/ZIKGche+hKq5d4rKnUZF+
cQT03Sw20qPjrtsgCgZSJLSDYqha+Q6c6eOPOvCDGVurDUb99hwqbT6tFyDa
qnGmx1rIlgQcu9vnLTJ892rJDu60OUfE5zvRGAOUQqZycTu+vxcLv4X8itHe
msPPmHKRdQDPnJJZBCfhdmENMqSyxGrTEq1yEp56uNis/KJ7TfTY9nnV+rss
MybgXwjMDxG7jWtbWc7cQ8SWE+LRNnCsp5c+2x7HyUtVFaRtcZlNj2bRGk1V
Nui5D5JxGVUaZ8TzH98RE07Q1c2LE3pJrcGKVgtaWZeV+Fg7lcNLAc23fKKa
+Oo04q406vIXMRi1FIUOiaChLkBQ+fYp/V0Gb3B/efSWNWdcJuZ12ZMAQXi4
MEnCoSWZcl/QB9LMNxjkBFFcIfmSTV8SZbIH7rOZfB0Q4sr6fxvRV+3h1Jj9
m5io86CqN6+AYIvPJ75leVMGRjCBrDEGK1lG1uLaoVoo+6Fun1Bung/dgEDM
7KC3UMFnej32GF63B9yLM6VOzDjXfC+pTw9OrHItAEHVSDdInEhpjMY2BYtW
425GZ5S70ZRPBMI/ljpUxGh4drniantaj6AGxZCSJ5qpAPeP+1Bm7zVPx+0j
FoBmt20qZ9C6tkiWPuFPiEKVhrUrwFESmlfmtuOBSY5LaRFJXTsY3o2S8fjb
mRSNqnZcviVIJqgYXET+AGvOB2wirZXjfZUsI/qMB7eHImKc5TydhgvuIh2o
00mK2BG67WamkO7gQ+FX7xQhAwVAn4nGw/iG56Pigqg1BaI+bU+eGsV8IJJ6
wurlcUqmD6S8GyVhO7KIdBGiYXTMA5Ioq+H5cw6dilfDawuiuF7Vtqerriou
/tSafIPQFinNyoVoRPjP2hp5wRPTPaYp9mci1OXSEKVj8zvfHRT2zuIKP6J6
e9SGmDZIbgNRDKi9yRpFzQQHhN1LvyHcIyBdNbaBYnddMQd9+jfInky1OOyo
A76SWiU9YLMA6mmNcGqJyOKszTvd1gLTACijcIDeVOAR3Xu7KuvNfZrUED3G
ucFkWB92ql24tK4U4wdDkP3SbjjBkcZBn9gmvKdjMFf4p3S9DtnmvqHWr41P
DPiO7J2fdA6ga3i498Hoa4Lypta4rtpUOggbyQVKUZyz6dFUopKi28sQRfto
nJXf5lCWoOa4UeahOKpho+Zzznj90XTrgeu7lt2R7F45HA9yiBorzDmQlCAz
VBmGCiZHWDFR+7i3JOfDpYALzDTFo5x+ANsKj6M99GSp3VA66TdWgB49LDNb
AHAIkyedYXlBiNi+w8uYCpNDdwYRrnVq1zljnvW73mO+NyM6qq2dcTijTsBj
lX2FUV8RSGZ45XsjEOUHJfBf6AulF9MZV+fbZdluWqjJgez4TCuk+XrWYxDR
7bA5jVWrRZMT27gwz1e74+BRcrd2RZJQBv81XfwuaiYTdofOZphtdcEmNpPt
CAv6EgLSfO2xKDJcnLo6ovrSX3OzKpPLnCwVO+9dlXPudO+N00F8P2gAyz6n
Lbek9aCwrT4NMCB7VcRQEfqF2Mp5St/nLHYXiQkSlNOR0zBd/HTJnwGxxAlg
+HV8FcpZ5m0DjccjgeJHVxhF8aysRyOb3IH1TKGaQq+tr2VzPX8yLYcE+Jea
WCNFeMUZurhIikHpsgmaWZVJmkvkHgv+rUp91RD459mXkKTdyOf5VwPFeg7j
0Qj9NOeupBr5Jivo+ov3NW+l+mRqPg6td1BqhINQ1vU16dft/MupNY0GcEZ5
AXENcge4eQAam9XCD6oG+i6A7AAwMJYOFCoPM/dbZJa1yv6112ImoajC17b9
JVI1i9UmCkDHjcvplSQ5Ir4RWxcEMZ//5bq7F1h/x5WgtSylLSBkYQvzTy3L
a/w1i372frw9TF4ZYDsDetgXdY5BNtVte9vVlnm5kmpLj5RrNW7yMeo25N6b
3WOoz1NqUYN6Jwlcf60Jgw56+0OK+m7sRMkLiZB+/shXwnxeGMIqv5RzFzi9
hoZoTYoPANsT8bqa3sg3AAAq+Ht39JxIm/BDqNl2D4F3XhXfI2syQwhxx6kW
QSvDXuBUtviM1iWGsxCsARDji96/JHoxUTBmfCL66GuRy1c6eGjxK+UwpBhy
H5RhxCX5Hfkah4tZH2plWpBm8pO3BVLbhkQz8zfrpNpGeT/ml7jNVhEj1Hmt
CZaC3bJ8aXKNiOEaPIX/N7c4ztd+TywocY/59iUrc3bw0YbnsiGuttSJeJQO
XLkTXf84EQ2x7BuzRUrVRbpBH+D6VKQKL4JizjQaY7ORDz7cJ2yBCd8ukCfd
oyjsseZJ5F+z9CSzYVqINDQtWo+imf/Ru6SS8nnGWDhueMGCo1x+NUb3RGeU
N+LDRrEew3DKRshZX0wDTEJDiyHJH7fpQXRF2vnLn8ImXfP46x1AgmlkCb1O
/2/tpBALDIFmFeIO40dXsl/xZYfKvKfU/c120PVFmzF1JEdMIDo7cjPiV/qM
Qj6PnAdwe5zPeBajwVfew50FM5pKiedVMP6XmW3UgOJgkv1E8FZspXRX2jq0
6nAPiu0wqFWWwZXgigJIaszIiO8oF3VKJxUs+xMRAHCzwQ+eRKlSEqjHTKU9
WjTbEMT53qcKfHRSIcrs9/Sy21jtYr5tzkzH3ZCAppQJ2gZ1QyCc2PKA7MVk
DbD7WHt+o1agD+3RffQM15i0oRCF4/ncqczd/ToWQxDYvN3lAGO2hmQqLz3v
QbTZQuceyi/CfKCabrhPkoIC6+5nL6etLiUEmnBOS+ms7i088SSy9ilKWGLk
Y5V6z1Dj8iia7ckXJHq7uiiEsxF1jDl97v3K1K3UtB4UjnC6pGuy82rPrhOG
vlBz0Hc7+NCE/1GUEBPkZxEx4csOpp1ADT9CPC8DanuksGWy2009PtGsZL2e
PkY4DQOCXCu2+uY=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wiJC+7c0uRxQfeX3b2YzhIuiyIbo/hUNKn64qCJNGP+dBoAJ0fohhuRPP5liIS/dz8kpSUAUvEJ5IocVHg9KzEOpq0eYt5SRgT/Tr9FLqhVdt6aUFyDviYP8tK4Rl7aKMQRzbJpK00spCGGGNN4crSqUd8U9S42n1Vw7frbVJF0joHQiVL7FFKBQ7qJYobJq3q2j1+dKDdaqiLbinSyOPdGbfmHWoY6UAYKbzRLyVdcwjK4P1tzq2dR+HVYgZBn7INF83ZjEb6F0Ts04GWvXrDp6Xi8o7RRuV+4dv2jfkzMWnec9MP1qJgu6mOfn9nybeYtWw7Pagq0yJj90zqCzLLGGUes1vAIa/b/ojAx1GpYitw/iVrdeRPnizNzmJ0TV2IrHG8VGLk9JqQtjxXIDFZyh0cuiRWqKQ2jIJi73bRW9GZsDxUesH6VpYrR49d0TTKgyp4Ko/91Ah9wjheCL+ebV5DVN5k1AZ19o13WmUAjfARWh8oxVjjkIcan79OyVLc37azFOynNxyMQXbadO02VCRMQ2XD45i/q3TsTxIKgcFTuQxEws678++6wAnbp4qsd3+EvXxPqR+Yu8vBzQnS213QcotgZc2dS6XGQkW85PQJ2qOOZQOBbXB4aci5mEMI+5YBMSJXfBKdCaT7TDJBQYSS6PXWPrjv/+DbjpgenT661ychVxQyt9msk8Y1jo9sm/+hJn2C5u/CmOn8f20+i+C1++KhTLE0/vvZ7gKGGR9y6Jja8IqCqc65vbFQOXtJBOzLyk9ZHHe7s5DHNheSX"
`endif