// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S8g4G4IBtKr58kpwrAGYaieddmW3taSnSN37yydmKJJhDwy7W9++KSx4EwWb
i1jvJrxtXbetXZYQB8FecB2Q0KRDlBznN9wB2gAoKdhO/Z8zz/eNm+ohXKbm
AN9hQBta+8k9gVDQATR6Ej2Gf9dWfqKkQDef3OcyTOKiyGKJ9JDgUAobUHQZ
IJXx6thydqJCjfD3xl7NnCeosWxWUV2kXqYGThahVtyNS+IZIkMxLLXd7lYG
aVPBD489mXVvNUCZfLXPPjyx2quwJZi0ABH81rNO5lnzckEQG4mP1FxSUeV5
E+XLqQMR6+zGUqZSlV5uYaTVE2SYrh/3Vp7fytbFlQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RA7282pOOavdZjj+gVt0EyHzYnUKnH/6pHlh15XewvL3yPZ7TaGpKqi8Rlsk
tyi5dG84CzAL4lPwnwmQTZ+vilL0/ayiYPnhs63AwgKQ74US6S9eQk0xooku
qBWgBDcwmztHEN/E3g+GEe+cE6WWP4xI9SOPyEb9jNBq0X9pMU1KTnYS+jq3
5a1VVoJWjyFd2kQjDcJum+cbsc+Lym5NIn0z1rNJJtkwauRSiiQVgxerYKP2
cBxLsBNCqod3laSom2bclYGUTLDPG3aRLsKaPyFCQM2DiiXawgV4/0SsgoJx
ao6AuZfaOCgiHduykefujV23NJlCB6r5z0YUH3YFBQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jDifUjq3r6deKEQxIc7e7HTFZCg4UaN12YIquKATjfLvg6OmaBczFJ6BwtyU
KkJvEVzUi8Cvb+FhcOSopdgU+i3reigCMc9742HQAK3wshD2r6DQKZ0vIsMm
mVsDRVQMuygB5HLYv47Zd65ddEEyhi/1PbqGk2k8LSjIsIXDlgvMI9ZS0I4F
mVrs5Ns/tIVO/ERIidNAFdJwZeo8etBLIrMC4AVf90GAuVkhCasWkmOoZHoc
/3A/4XNlAmYmQFq+YSg5qgi+n7pXAHsV13kOT9T5i1BKjYStKrdbzrM6Dnpq
VCXFotxX5en8pTW07wiRcdMo2ESSPW0x4P+b0piBrg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MdtMgSgDLsWtJ2WXo6/aQ1aXzQFWCeSwlSeG1xELEY0Rf5Q8/7tvakmOqh4d
lqO6SL7rNq2zBMbvlwCQD3AeBHdsaTsACFs4H5qPrT1GkH9juNYnay2UySIG
JblQnzVkoOIbSZXAhk8pn5A+FK6V06whQOkH1ChPaibCgG6EgvBtdvlXQhS5
gzbMwySfhmRSUwR0BKoxytJ6Zh21XT5LzyIe0TkwJ2PXgBkGG6wM6/32Ita8
1Nw0LnBO+OJK2EtCg/7G38PctTHVaL8FtZHH4sM9o1ytlA/e1vF9EttqgVXd
nZKYB9xcao1WTJbRbfTRmR0KKRCE1G8XNr1IKbo73g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OVy4S4O4F04THKR82mz+Th8vH1RZ6/eYSRvfwFNYtP0jR2A/OKWtTGzj3Zq6
npOVXdX/WqiMtUG9fmlLrAEm4QB8sForxxcVSgRcuYO8Cg1fxakJoTU/9zJI
osb/+zuOsMA6fEK8p+BFJvOYFvnrFupDr81ZCRDH3e3OqqK9aPk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
kaIUAWmT3x9fDf4bX9H0+dH/LSWi80WIRrIrwkW2/HX/J2A/Ydz9Keoy8RQ2
tRuF5gMtV/mAFvF1zj3iF+3riMzB4TdloFjtFTgVvvOUak9MOKaToy1PQ0j0
HVr6IjoxJjUoP05SiJzAcOKodEmGks1okXls/0ZAwdoX9n5EGcn3f1XMQw5Y
sjb51n6+nx1zoqeHzTNxaZ0zfdI08ayMYAUqzr7nLF2S3qoB73bgNIyr9j+T
NkwMhXOH3m7zdDz/megWr2ye3zgJL49Hf52Eho/AZTjiXSdhrkE7gCRQjcVt
5Grmg6KeA41BcCip0JjTc3YAb8F1mTkG2fPz1FpOKUCzi7Z5gD59LC9u6CJk
wdR1wu2s0ShNilanTUbS51l6WUw0CKotQai89NnfUgEwt1NHEiSPItncfj8V
0kxDvlW4iGwzJW7trTMjCQfwYBrmDGw2DPw0vEhBQNWi6LLklheJaM0VgqAp
8jW11iDlCuzpridat3afUTqWGvkTpB8d


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Rrfg/aCCHyTaKro6k5qFXkm6MDZy/izyV/dyIU/gzaI1cvBDV2NHAshKMkCb
5dEK54Nz0sF0aLTscztj3N+ieZfI6Q1zVgMJPEigpRKRl02pJvjVL3jv2Ngr
aDHHkXaRu7iEiDHQAJD2aZ7bGTEE7nhOvSphXypDyHQLBfCXtdo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EeEg/gnYsbkiF3g0CVpqVXa0kAOCrpCiSsMQ+fcAgY7c8pSHD//mk3lPJB1c
FPIKmPmv1FIhbdQeZidj27BbavxbZrU1Q52gOOcp9gi91fi9+jyZ0YPrC51B
PZP2HzAw9lqntJ4xbN4vtoFikTKJ81afuxFB1dHr0pARsrfQsvI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 50640)
`pragma protect data_block
zdDEJXK1lwrHPrJnbwm03SsCkQfNjPReF6YqwKbeQMMau81/ZAhdgxhaBplP
bQJFanx2qaHgpJkRQQgJSReiBoq/py717dqKD1WVMCVVyTAL4GCLAEdDO9aB
R6VlBfwW9J9uUJoQ8jj1MY4f1f6ZikUTGW6hHrXzwP84szQY9JqVFNsThh/V
+1nzF9COUYw9jwARpeosUCjiAdRxmbHBDZqNehdDefzRug5FyTk3/4AcfKah
0jr8l5Is25QA74dOJPUoLU0g9As9hM5nGsF4JPIzzN5BiVbN+VVWY/FnLh88
xCLZbNN/38Ia5nPrfuX3S7LezlhBxzBPv6aDWZWhtdRvu41RaIiZBaAUY/uR
NSKp5AzBd57iunfDeOsHbgBKBGhz8AsJUk9YoJRbCKAyy5P60tFZJUm00Qb0
SBpZm/k36oZ+tMzg3JNg7ciMA1yrBHZuN6xtbcc3tk0lPuVJkQusUVdKkx4+
dmVl40AZORvHXtZ4+9bAyhQvj7p4AB91fvk9Jehtem4tdQOjtSDRQZiQ85VT
rQqJ3suDdO8NpA0Uq3CEVKTTADDRTgmcaEZhRiKcs2S9DaSAGqLCjNAqT+Ot
IXiJU7y6mKEwDl5s06AVfhPRLs7mKCd0WIdjWz8CgXFLRFthYynbCFOQ6vkF
SUkQvl4FLn4UbWudXOxTbjHDkUxwxZDAAcCM86msh+FHaryYYeWi8xaM4Vvi
J4Jz6K4tqSkJ8FoDEwuzhDW219xv+F6jgE5P4I5gmueoHm5hQz1RkpHnnNb2
VQIDAfTyqkjfLrEW+U5fEaKBuI5157xGSAam19JgLEbMWaPvK/XPePvUts5A
pkznVqtqQhix8/Z1tI6FthtVQRV6yQ9hXqr7DMrrMI0ASlXArt7o90Njs1p2
OTh7Xw4nJ+PsU4pPydaytpEQva0LGrOIFa7MBKWPB9XgQZh/GOXDBqhsUWbk
GZ4cxDXrYj2lFfiWyesQ/tjAhpM5A3kTu2dvI1cLXe9V20iaSuC6ogCkDe2G
NiAK2WtozPXzz91uS9pqRc1A0Ly0ejkcHAolzNk5Q1uZxDoaVmxReU8ub3TW
q7l8wgZ6QVQgE3p19KXPHuDHwymqg0lLl/+v0/067YfMzvu7PZO8O4dnB9QK
OBFdFdcBPVzGVqv7fYyfpIJekXBSDQoUEUblv9VNu6Fpgtzvbwt+eWtGzS5G
E9Auzt6MGFWApmvelogVVTJT1k/hqoNaAr+CqPZO3Ya29zypdp5XA/6RahdY
S8xCM5yiI9HPnE+DJ+o2HjB+mDcHmMjaE5sejqtrs0lBDPZQPTda/QzgB29S
IzV4QWp+1D47odtaXaoHdyrceefOctSjEPLP+sUQmbsL6Y3/7tn/DoHbFGxV
s11cZxCVnVfznPn5jKDJths4yTmk1W78x/FiTisgRUdaCFh/XrOUacwG9Mf4
Z9jBtkqnFR/1+HibSuVugbiUbVY9ijEZRs2l3eqr2FpmUOKJ5qNBFKfozO9G
yJQ4PRpSDbSH4oaI950JA5lWaUQnnyvZJVDGVMtyKkUWNZwLEJ+lRRUOJ8c7
XFPtL/SsRe7g4+WCQd+i+nbNS/3vFjmMahlTCn/7A/GZPCxr2d0YBNiElTZa
QH5izVXwb8YUhxz/w2N8d1EPnH4LevXjKyGUIc7Aqe93shUvVlNdCLc+Gf0y
9eMS3qbXJfBXq4gYd/ERy0JWIVAbaaRVpytgsDw4XcySiEiWjl/T9TzBU4vy
IjFBKRqxOpps+HHGeFBhtJfyerlBTMT/EnvY7lf8F1sxl/IgGTwlZLKwHcsV
danByCbJ9q1JrsDzst8uq3x4hX8jeaASjpV5heIyPA3hkXXSFmy7yfmKO2L+
mPnpsqZCNKdO5zrBsTonkFflx3B4IMJw5y6NCCjhPKY85b99X8yEruHkn37O
mZLOq+6u2qj8T4rOvmDFLwHzR2V3gSPxBLWZjYjE6f4qqNBcSnhI6nbQzMZZ
1G9V8uwHnweVLkV+qZ4rtH7aaBazetUpgoBX+IeylVSaX5Buh89LrfAniT+J
uBfrro+Af7jci+o/0/rN+xb5MU8esIDv8dQ9GyLsa3Zln9a/yDfO8HKBn5tC
Ku72mgOG6HiY8HC2nGSGmxW3I+Nn6kXDxdC5WSEvk1PyE5JC7Pj5PJkmkMHE
7BfqOqhxtQUxHGYGCGbflCkZYJqhDiWGy4wVLD/y3PFh8VQEGdT+CqKQhvtf
SDNufOEAvBZRjs68HV61V8/0Wvm8iLY1eaMBukc+SKyf8UkpdHwLf4nGYsdg
9yMK4Di4L0HG+rxoSz7FxtUhelh/vRSoL5gbKxqkUwGjdmukLjQ2tRbOXZZH
FKaIzTm6flAZJwCa7HdbR60JmwiVglb9wb6f4m2ZmO35KLVnz9RldxmIHp7l
yYvW4FEP1qCmAiahk0vV7/FRjF9HBmn4oRQD8qJpO+bEZEJ+SyIeg43A3nRE
eeHJoSZNoevjQmpmmaCiPr/DBnpfXTOaev1bQILpTk34YnYiKzZVXI6ZVTUc
Tvwn4dROnpHNZOQgSfobCobJEKoDbVyrcFLXfVWY0rhTZ8zvSXPXFylVxHYI
t/fHQbpKxXTBi1tzRwzpnR9BhZnnc7Fqd8YaD8ubOPmwe/jA0PNcvleym9nH
CnWUmq9hyXoVqsCwi3J/saxkpXklWHEVcXFzNVmACc1yEGpzwCzq7ElRT1Ii
f//QMNyr/bthsY6A/sOaqNVFPNhgxVXiYL6yUVDfQ1RILR3DFv5xf/kVPN6G
Oea7tiTKJi41axE0vo7hvZnHvfDZ1AX24lpanK0T8WWQQpJXPD6f7INbKGIc
5uiME9if1OEn4OMU3D2RQHCAzEQqXu725aoOVD2/PpiS/LF91jEay89CpKDe
JSMc9II5Nj67r0LjxCx9XRt5Yr7qgFu7/Xz7rH5Z5rFHWzfQP2Ka2xx3734w
b2q9GsK6h5+GVkfqrysu+1hwrnaMHbaZgLGdSIBRZtxqp8JBa7kg5T14pENf
jsWJ2FKmc9ON+VxlCAE/fTx5A3hTbyLzms6ZWTEyQ3Rv/HLn5XWhKdfRZCUo
tJG3jIpKqnhoS9V7zCeglZwEjL5odQUysH+QJl6x2S7UrMlvSt9XZMyJL7BR
yDllVBEYCLak++XBGumDKRLBTCXNTrOzzDh1AsBvXKED2g6XGlRuEZrvAdcs
6oIpP7BKsQx9RfvuGbFDI6tYBRg8I4MX4PziHO+53gEj1NtN5LhGq3fBXvaT
TGMhKznZTuf5zq1gEFme07YkWRXm6HAi8e3sJz5dB+Jt4HE6dh5leVHbGgm+
kXuVIr+cYS+8O/FXVFJHDDhzAXlBhLK+812Sqb7bV3TvKZotIa9xZe3r4dsB
vwS9BKQ5B69dBIUWidOG/cMrNPJkoon+qNixkCYOCRd6Dar2bBtdqyzBehuo
pYjkUU0HRUODWFKCyB2O4gSlO5AqNl5hx5zXJZWb0q/bo5ZL+S+bUZfnr7m4
sEDv1+RVcPxLmkj7D/SUMits4IMoPwBqD47oQIla1toRNM6xMNteKQF4GOJR
+BUMaRZonbMw+K2F0GAotQdS+zTCovra2RZN13DX8Ltvg2IJzYym7Rjm6I7i
R3IJQTyKGknWIZzcKJ5jZROEUgF95zUtgSBH+bYR/W99BiGgErRTyDuzEltG
dJSm41D44kRCp9tbkprfSbgnfr0tb8oivsJCDYO364V4t3cHzo7BGsWv4h+P
zcEJ7RgjUSxzHZTI9bs/KBiLhGgtPkJxoevkSGBhGQ8jGctHrd3JQa7lJN9+
+sE95+6s/pyfIEBlJqxVSqbHCj8Tx623ZloR9rVsHQRqO1vFpA9+l/GOovhX
bVPn0HATKD5CbXewCcAA+69SoEAy3xB1eXeBkCYg+AssM+9HAj8a5SjTuwql
KY+itVOBaoRZnhvaGPlrvfqs4+96DbxCHwjdOyBDOZf56msnT+tgTfShpSHz
tYHO2D6OjUrd9aUB9Bkl/KV83Ohxp6/NaDwdCHeaEE8MppdpqZjGKHoT/hIZ
iak7WuB2j6FcbGvJD5dYxOE4qWqsLN1TDPmM72IT5255bmxB+h0/yg1M2mKj
Npd9Joks7G02weedtY9+p/rYyAJZxXz+3GAmJHgjIsU6EsdAolfwNqxd9NeC
FeL1NLxthlw2thSQW6TncSFgnP0MqZa4GnigI5NuXxLnho/2mrjYeNKDceyK
7Mr5ClN798PJ0sBvxS47ff/FIQwtutxHfnt8v82stIjp0GawywyqynKnO2XH
IZR1JvWWbeQ6YWrh4DQrkjAu1pn29nTLotJMvvMzkg+ezm2ndsc+Ds6W6/BG
yLXo9dEMOCA5oPJAp7VyqsB5/x1FYU/pdW6M+ifW3piFMOLpXctd65QHfSy8
8e+qmL2Pm1BaS5CRYbpFYyfszgqh8i5r5DO16bjbAIxE1hwVCcD5kvJP5bx8
TJ3ioYUv1u4E/94C7WKrJ6b9sQoxJ/bE4PkZUsyapX+IvmYFR36vu4htmHO/
9eZ8Rft6+XtO3hcM62Goz0Yv95igHm58NmTc4P+D3llwU9mGBpwlI3yYre7X
uWF/vV6oosM2hvejRiMdZifgUgFpEGnUnpP5myTURDNRapCmhEYH/cObaCmy
evKUp+9oeZEsoFNlUaLpYkBqTVReuWgk8qadff46fM9LEQhzaq+UKmqB5aqG
syf3dji52vhmo3U6KqoXEuPBJkBBpC0TI10MiXdjRtmwBrK0zL1GGQE/DBHU
8ir615c8q3PTZ88JdZ024eEIu5OphSIAHLLMwsEO4lr5ADHCVgnuOQfgvw89
4N6Leh5sjGoiwbqv4AFyzpGm8OtNAPM0TPf1w/ChcxnvXTpnS5QuSu4GTO5M
gAd0psN2m+GfEVkSg9SfSoF353mZgaJGCzn4fRX+bgbrZianRANP0ieqRyCN
w4SaI6XmKhauIUvYzde5lRngDJ0yM/BmOCgpeGaNzXoGWH5TPeCzZaBKHs1Z
sTSpbmntCoG4GEZsoOeJ5xxZ9CQv7RWw750EihRXJ8XklRUPoJNNJbTV1fb0
JMu9CNhGcWw1NPXReHHQnGPT4K+fWHy9lB0KbyisjLqfuHZ+1iHs6F2n2xSp
1+1rgMskyYbTm6NwGiGkTQofyUu8PU7wTlhulI9Z1Fj4Rtqn4WkbfFxNCywa
gLgDpR+0xsuNA3lL7NGvApzDQUmdylACgsO/0kdVc0Im7aO43Df//hyp3XNf
M1ewhRFuwPDqujUlneHaGYeJZ9VuE9cdOD2q+bY7GxsSb8bRQK40B564Dr5C
Ln+cB74fFUvQ0WhSYgSDcdW7XhSrQKI7wb0QqsdR3vgXBq4kxIEHhHvbXLYk
KX837vhd3rkk0QMIYS3tvU1bPcJAc7AAIlZ7g3mZdhVZc5r8dfT+dd48EP6P
fRI//jq3gSdZ83k1k0906TV4P+aeIkAZuVjvD2U61whc8OnIZkF6IsX7/nd1
OMxHRk1BDxzybDfHmdEA9SCnLXtlRl2ikLZwasWy29/2VPTHwuLf3kznhZPO
c0FBJmzVq0+o6CLjAPSSDKEMgFyufFlFsp5j2PR5PTkh4az4SKXGzqRwHkto
Ju3dB7SRLe/oearwUwHZqtuzcAH6JKuQH9dgLK5P41uo1WUa2PAZ/ccfJxoQ
lmu/gM4vPDeTc0avimKw4RPmZwLCJXFAVo30E/KZqibIL617Tbazgosg3rBj
+0EsDM96YYQYo3q/rO01qHJ3r5TpoS0qWbPeCGZxrsO9yO28UIkAnXNhkSms
LN0HNNQpNMEU6x27Z7iQlheBqizIj4vnNc8u2DoRWfEkRUqnKC9fKFcwan2a
iKMxWkNISX9s6moT+NRe9vDUQ0VOdOrglnG3lH5dJYK3gqc/1OGIeeopf6oK
Wvrc2CeiiH90av72rjkln7eXoyoWcgqETm0p3g0ljgldqrUGatrWuS5fJn+4
ajSzLSjMvLbhIDRBIJ+Pn1aOo3tIy/3N5jBXoOVuFm9ZsTICOGzOruyqlurU
zmhidRVZL3ONovbL55Yj29o7hPgjEa8M1P1e/yWfQ0jH3bkBtpES3oU0sghX
GW2D1VE+winHSwWO4KIXPFT468DulaCC20Of4qX8zMmzU2dTp4uHpsed/2Vs
Cu7itOXHKVDTR9Wi84knufRSJWs+pnJ9Ruaqt+CtYVf+Wa++sslCigO0qFh+
dhbm24V8Tre5MynYookJixNAUwi1HMSphlM4XqFEaFvg+2LK/IS+9XDZDA4J
0qyAEsifJqRsRQ4iRco4a7d+jSaRKDhWZEouVDNLo5RD6b/XIIQKt9q8EIW9
Ow5TtjD7d1FQ36Gculxh2FgfiibYwwNbkyOfx6hmlz2RHhTRx5Qu4/PFus36
z6Ket3oKWieXxPz5IapOBeaHP2PwixcYB18jtFfdFZVK3ip7J7L3dCC0+eNV
BxPzdcAMaoywXVuzRy/FvaBkdYDZ+X6uu0n22/hzgMt12OjFLI9IG+FB2eQS
fJoJFPERfxyEwGwvf+hzP6WL+ARHX1/lQowtv28dxD5bkYJ5deiv/VhEYqB4
xjsYwdWCz9SDSiDle7enzP46tWniX+XhCsiIW1ba9KW8OSea3RNu9vkMIA59
EEIGlGmbhymD/OwC93kAfRopoxDEA69a9f1Ck9olBbbDOt8GxHjWqLVqW0iG
q0Na0XbpG25fQoQY4a70I4RiYInqqAW6M0ZNXhR4UImlhnJ/3kKzQ2viyDNK
bEQhq2vjSNkXaVl5fVxbbkfP3CdgkkHbZ0UAhoUt3bqTf48m+zqs8DG2taAK
QHaPIHtz6NQT3DqcbDvVPRpv5wfI0JZIESY56UeGSFimkp+54y6iOavsXPyF
5EAwNUd6/Q8mmSVEWHrJxu6GZ99mBjo3Tdde98rlPXRQ1QWtQlIXC6KRrLmg
komxZbwDMsFzHWy5oatfJWomPxac4MV4MSTZBd9htAVTJKElMH/7z3QJqsFb
1U2W7wd/aEW86svsnnXJNwJBLE2PgjaPH1rVEJGm3SIHaAgUJlpvLDQcdcNX
aKKY95ws+taDd1icaXDGq3vDXzOj6ResC75rwGjaC3Bu17ovf0PHVr7OiL/G
3F+EbfkeYUIlS4m/isXJkGXM0IZXJV+Nyf4F1Ma1Gxs5OwwTPliKeYVvmrQC
10FkNPRkjManxOq3hels30umxLjSopZHDHBWHiEDsu7lZTwWoIH8Rr3Gr5VB
PDt7s7VZ+8ik5tRSQa2eHoFENYHNrYAyDGafcDMucVs3wAyylZNzqOfj/lU4
fBHpOcG1lyXxPgDZ9dfOZ8s8sHASRtzBzUkfEyobmiMaJIVFNtJ+X0pTVXGb
M4ibOc7WFswt3wqtX3qGMsMaWXfRrHZuaGIGlEk9ek/Q2/NloLSstBNo3Qol
Q/J0IkH5AAWYE7Jb4rbtu0CLjQemoUciQOY697FWVUFvHW9b9nFZvxio4qii
q3TaaLdCqbHe6IigekjlDKhNmfetnJ80F83WolyEBljAx0CxizXLTvkd0lxr
+37oaSeGLkzQKtNg2BDVudm7qyHmu7LGkSpTrvy8/OU+WmnLdUV5hT8d6CqB
vae80B74QD/Gjn+79PTFXzdG9XRgTFmQn7RaO7GFFbj9fwI5Jl1wW/QYbb+u
1Q+Nd6g9awb5FSpKT1Lyf7EWO7VhAZxvYihHlaIDJGzg8HCV4TDDMuViVYPP
0Rt1cYpOcZevBOQDP+pI5tbznDdCDXgn33dIbuKbnrREJBxDGOWwJXa/tBee
x9vuOKRGaEqAbsEaBd7QETZrKs7PZ/LB3uKjTsP4Sr0ryz/w7sL57lZ6l7G/
C3RXxpUQNN7pTwUq2xF4QCr3ggqItiIDskbFsQbRyUrT0GzyFfvozgnFxgw/
lHe9C3dE3JDETFH5Ev3JyegtuFnzpGqShdTYohEmTzHluDhw7B3j5XDAQTOp
eRhD3Q4gmQzeajjsXBYXFSUSwaQoVBJOyDungo4AGm9VAmTZ+GUvuwKldZun
4h+9b9szxVdhMR3Z14/WcKom+/yWT9LBw6qmCIGHdRrv/y0Rf2lGCQ+VLnV0
XwS7PqlVBLYMTFZlf2pVJ+De9qfHzaVATXxCqmnVfV2UgYJX2R863hHNCw0m
0CYriVgr4r1pWEgYFtgMsJzFYDsbt6KGyf6Pj0Qc4gMqlofaAenC/J71ynJO
PHMMgGIPTFaHNDp+nAKsC4PvL5ZYFS7lyTi9G4uKl+Diy+SZ9zk50Rz1E5ZR
ya5Ws/SR7cTc7iNp+UeJOSqkD/LrUKaiQ6j6HBHZ1FI2oOUztWZolZFo5/jb
/whrTa/3INMktyffOrFegB8wLRRiVpAlsx4eg7PnRitgPg3hLLPXpMjvbr7V
+SrbMltFUUbLZH7fgr73AP9jszHW3/aoHFhfA3KWR83joPshECUB2As5v/qe
WBkU6pS+Im/5D9ydtHXjHZ/vEpCLgeSS6OxYttmqN5fhyN0Z7tojmTkdXtY5
BCfG7xDdD22a3OOnQAHJggjr+BfHR12n9ckWiRJemNYyD0Fa78KwthRN7kUv
kQuuUw05yVNRstwfcQnZiqftDV1s+OPSdGVzhEMP9HIsFe10WMynFECY7Eek
UY9NoJiQlfdBVGo6NXtANPEkg9hRFH7/A9Ispsf1rrnxSuX3mQeMyoOcVk5l
7uo3lads95fKhmlv90YbpINMhMiR0dGR9gVZJZQhib8vrmqVSt0/uzWxZ6K5
BDKEtmMcPNnc8/qC8oqFRRAROekgUqx3FpPHGYJlxa1YauikwSfuJWObudBc
X3abjX0wLx/mTD8EtVXn9Z/u8pOkTxAIBzntodAPGd9kxeYB4Cfq/8M/Vk3U
BCucUAllvXynwuYvnZXOUi8xGZedBvNaS1UR+/tBffcP+fQmhrnQ0Vs0kwpA
kX5RYqPEbS9yUkQH3o94827a1HCDvXJtEnn3y3yM6h9I0BEuL24PfZDS1VpT
cXPZzn7LDiDgBq6QqS2EoDqfqdJoeYUgnGR2+Ho46YkcXJKI1AbDZuAn3pbp
jV1ci/kLz64Xb7TW9j5s3GjLjr4Ci6OYDQalguKqxYPFM3W++DuUaH8jV3kS
MPvY6GnIFMh/4Wq1epBq2yQyGvyYuyLLZdw5kFN34UGpeRWoPgqRJfzknAVz
CIxagPKsj4BZpSi3kRW0bddCikF6r81sZkVYeo7qLdhjMos5wJ5YBEFeJp8e
hPAVAksVvmh2KXQww1kULNSo04zd4tn7WCaRbXHc0JddSzhJnvfMg8L/ZXMq
UH+z9doHWpye1p/U4Yf4Vb5t/RuriYkXPwDVlxRBUcXggMLrSf7On97kRXiW
q0NwFQWOCwF91aNF5K4XP3tlGh4oUt6113v/UPZ5K6QOC3ko/8l8vvnDp2p3
13ZlXT7WuMJyGayINluHqJejZn03DQQj3QOd5ivcpQQIQP/BZxAeAvPmANEZ
blpu3TfBcQYx1FuXL8FK/x4LinG6dPlnnT43Suz7aDPdjYGEytv90EiL8tju
on8Zkkgiz+SgHA+7UKxvMACbJCzqr4RtPU/eqHFFZ0JUA0pADelNZ7HgBmv6
+fM1quD4JtssW55axRv6oa1QMwCRlY/aGcALUY/sETuRIrZndyMGYl7TdcFb
DOmFHwtO7WOfTW/OwaK6+1epvTKy+pnx9/Pq9E2+c2ZXRnY4RrutzhoBfjUV
famhMDTxAfBPIstPHGj/2a2IbzBMEON7iS0e9gfP9CrMau2IVVM88RSsqIdl
1+F+M6WG//kwuCTFC6H2eMTa3y+7zt35YcohH0qM6+iX8jr5tzx2WY2Ud+uh
8MxtXIo0/dVQ5Ur2x0UPElWaYg/3+kyL4EGfgZnSawqRroqbZRSHGKr/BRQf
JJCeLZ1c07Z16gU33r9j1NcjfwvdT9Ox0vVznGQKa8jSkLzkUh9hPxt6DwCm
IGRlzGZkEz11/KzDKOOlZYFy+dEnzzmQGAndzNMKVnhceJ0lhKObhE7/ERMd
WfWsJcmcBh27Jwb3IWja2Dc5D7rsPbbGINGE0zv3ouWYHR0Yky0Jqh8mUuWN
xDZOx/FIqrYdBsfMsqpoOH8wWq+Jku2kk2TXSbWkrLaJS728EHaC59/G2gji
kEfCnXOsa0KMCjV5b62BLol+vqEHQqe6DD3dQJ/bBAoTTjEFs7qWdSFqVuBw
H1nd74TQ1j+p9t4wu9llC5CMXbd8iWF0O7Pe1qIZZgVviTduI2kVjQbBVsrd
SAUxpk9m/wP+lOLk/ZkkXRlwi2m7iwVLUT4h+UphX19hsd3K/WD/LTskdgh6
pOErTmnQY7HwX780tVxAt1PZNlxKGsJpx3k+JFrIbw71fmJqbjZE2tmG991B
oXlCfYm60AgXMRDUSyEAQjjcj0sKAvZ4kI+jyQLY9ByAIOVvEYe5vb/gv+01
7y8vfJakAUwUtY2p3JlbIgnMamld15JQRP1H3MAcxMRhdnX2xTR+8eunfBIm
XLUiKf0/TVs+rw+9N7/RkVT9J2/offLDJV5oDLP40lkaSjIiuq//mfcfL4h0
0gPI6ErycxlbQQZHUD+3Vbaa6qLiDkLe4vKPuTSEGRTAPX5SBpDdNMTZG5VU
2ig29AWUWcFQVffiQf8LaYbryIkNfKsf8VofkP5UhvDErJf6FS0rym8Kc32N
1kjcH9iq7Ym9e/TKiuNjII/mMzBr7KIW1cJF9RCcsMDAxPCLXmYB9rAZg0UV
eoz3xiIe2b4COxA1PVrBHKyLakjWq25eN6oo4SrbLAKF598RgzaiyF0IZ21h
cufTLuac0YLuZS17ezKF06ozSMU9PL+OVqoZoMwRtBFUMbwK7fqbT4mMtlIb
iNz1HTqeciLEWROHenx/hsfOWxhnd0GZtzvtUfb6cXyxoP+ZD5E0SkVgctLQ
Tqlu9rjcemBO1KWdsP7vQxwiKkmhHLsM03z1+1LuUsFEWDikon28nftgKBsN
gHwGXza8+A2Kdzki4UuRjq2yJX+vcI4IyNd2nGl6XGtPEPGvurK0WO7q2Zvl
/Q48GQ72wm1Iss0fAFQULANp0pDZWLUXszWYodtLx6inWM75pPQYHXf8Afm3
SP/SX8G0NIvfRKj7LzL//WycI+m4NTuUeSDIEWbLWFqR9DHjUJQwMqLbYQr4
pLlsSCkYo7BOW5KPOaq2GJ33C0YWE/tQMmh0gh2SDMW7xjQDDQZEyyuqmMC/
ckd9UNO5LbfuNzzzQJdW1SA7cSGbsA2u5kXtHJb2HuPqogVHjwvfnqEZK1kV
97KBIMQsK5E9RpLdAPaDBRX1jwDWZYJF3JqofWeeZX12Ymny8Q+kDN+1duOp
F3HUFKN7hiJuh2hCJC+QXL/E5NQg9xJ43Iny3fvdDbHQ/aOT3hAJQpuZkDoK
voo04pvOS0q3+VSrIkceQ35eakabEp+CkUZ9rACJGHkzTK9YDMvImQTUlz+Z
7g0+cIaeN0Y9CSMGWUMfK+MRQnaTBBwhmXpZ7d4l0N+xFQFGGGIbOqvvZfna
OaqSyDWiLsw8IYI/EEa3yLg0xFWiXBbsb/VJjWHI0fVDLslypppszZHiKkZ8
s/zC1PkV2atiis6SIYeZDndoTrISmAS61/XGkO8nYlxUHQ4GcEP+ywRVSYNX
fRy5LVL07kaLEa+ljC0OyurcwKHKnn0ESlNSGigyDLHVOEf3k7paREIQiHHY
bPKP10ri5/Smin3zbbAnOOVACkT2paPS+tO1RRtvB8aYCzgyyv7e06NmZwzD
ph1+F+1lFmlwOHznlzmwWdIegAFXVluAqkTMJG9y0BH/yCVVaHaBOJ12SXcj
T/HqPx99TU+wd9nG4KOEVr21Lo6JODlCISg1xNkom9OVdIIsIq06jqmbQamw
NzQXs0pM3Uer6aEfafTG6c+0+nUsAQE0PeXS3xH8N/XlPSjoTaX6OiEVG6wB
dsIb4T72QLDNeeP5hzeIVOuauqiuSU9RWtCz5v8TnlSpWRFzka59b7NtS5wa
Wo2YMXJQNDwNMYTq6O/w7FHUmfWFXgAoCZ1m5YVazdNG9gszFBc52D1K1iDt
q6aoZhY86LDPvXsuacSlSl+D2zSOf6PWx/gNfEZUDt06lU//ndiYdYFvb5rB
rhnSBJcFIrcO39pWanR5bqNv5uvETMAkjrnzNyU3yppBowvQbnYT+iTSH97A
yzMiMbehBNGClVehAT/JevQTD1BbfL+zwzjmdz82Gbwx+NLmgDO6rMAe+azv
iTGjAtUTWgmDsY8sKVvaOuip9rAQD2njyL6i1nPHzsJ9POoLtsYVNvzZ3C6Z
5dsTVY6kUJDiFWznAPm1yD+XfqMW09lxxnug41OF6O7EM5ifu2z7MMl5Qs9s
f1fgfgRqmQtjXONTS/XG4mQD0YewVh34jDM+YM1DBuos5EPIgzlL6x+R/Bgs
AS7yl4Hzye1myNmwBK8yUbVeorsYXjCNNsH77lD7XpzqBWf7fOqOx9DIESnN
7hcLMmYzSpUa1Z8XZtVl8/9CoF6rDeKzrfLHw3KvLUpk4u5eiZISnwjK6cym
FVvqxxAIc/u+sl0kuMKvs61Ujv4kk+Mq7KsI6nTmpvbZuxbctte+nxnK18Tx
BryFFlfpGl7ilPnGEnNyngBlghrW83hQi13fIDTSdaoYU+OP0mIZW0aQeG4r
ilJSwnZdNKCDVoGCAtC/mABkJipgjawBQ7BCUVg9Lo8xmK38MgUlHt+jrtxg
zU3hzfgsW7/+cNHMC5XC4sHRupLJ8RxKwhvQF2R+IOaRDXnBQEo+QdmfBYDK
TgFhklmwzln3Htlzc2HVlvuFYLjE8gwqfj2J1v1L4ujgRdiikhrkcHYRiG5B
n7dJNOX5XMXLEINOvdBYncky2wEVZSQGqoUkFsIJ1pKPS2mNWxq5ff/1p4If
0+akT1mFx7UFiCqAeKz+7PEswWXtOJDl1E6U5kIFaq2XmWo6NSfA2kUwFWj6
pDb6NpcXf8jnVAB5sfM0L04Nd/Ym0C+4z0DYzcF/7Qzs6ggtuawN1q7yXbl8
rbgvu7z31y9g6x/CXrjawxQe6Uw6W/nz3S6bA10d0K5z2ghUWruEiZwjuG36
rps9oENIlDAGsItdxUHAKp5lrA3AS0rsSAC9GsnkCiSScZjp5gpQhuUtXbnD
ozqbcSP7D5ugKfeCtuXKJEt3stXAg1IOTOOBUBBvktF2e1c6RTFDwYeSh3n0
6tw9ZXpPUr+9LvcUtK+u5mZuG8wWq7Xh4rCRBWWnol8jEBpsPhSe3oPeC+ki
x+VKgdX1F+4sr7IzyeDkUjASRlCA3+wT8btHcA5w/vBV0u5B09/d/3RFb3rf
f86sZ7CmQ5tdkx4rx0+m39lfPhXxg1Ei/EQ8gey8C78URRqV3niExdA5cocS
fTzkGsYq1wKb9kmZZqvwWGOBORIOfB/PA/ITtjoSSqJldZPrJb2xrKDxm5/g
d/pcn3xevEFrxo4aPeEvGpBLLV2cqrbTR3DygeYXXge62jwj7HGNoGvzi/DI
jCeUXK5saAchM5ty5zV7TxtsAYO3/fHEKk85fuowllAnPz1Gvc5fb7dOujDi
y77j5B0ahFdjDIa/Aikgwo1ETQhzyKlyWfb/LZsCY5/WZjPHTNun1SojUD6v
QxkuJkGiHhLZD0Efk5JVmUdslE3raRlWszSITBBOd9YBswSiesREQGRMnvqh
WnTyEADV6Um1vylsPgmsYJcoAkUCFWnHrnpVCXg4F5rbQv6aNglKjTGbUqWn
0OB4NMUv/M8bHkv0EhYw+q7sGeue45lueaHPfCAuvdeJOPzEnMPSUxH5AWeb
M7FeupmQaKCMR+hYy+rTrKEdRmJUDL6G/vmpjE5fcC7dTEYSsCdUwmBz/OTD
EqatFHbPIXoA5afr1npfa2dhMfVS26H0OVYROev+7HguND+MQHZ2SUJv3zu2
VEVoP6SZCM103RiUUCaWD6dhsOgz9qku8PWTmT+tDtn+evDAMgCgLLD/wyCk
yN81GbCm8y2PG7Kj5YQeCclz3o3h1Dhm3P2MLNNnGcSCnfb5iMoAQXHwYtZo
cBFS879llS7dNfBPFpLvusVxSxPV8wX1m9ICRnk8KjAXn0Ew4MiNKSEIby4M
jCKVWzpNcgW8OJucrQBtymOwd//482NcYMYeUZUbAz07seLprBxjzbeXqCfw
t2SKLY6b8FVNAw8EQu+YX0OshUWiGvRnIhyeTaZFpiCzXt5jQeTSaxJ/bKix
b4gcGkh1oiyseCFKTMsWPC46WG/5DhRy6VVM7Yp0oZr6PCVfDBNaQ4fHak9l
0GBYyATyqK9+3FyomQiqsYISLiL6KHrYoaTRpG91KL99Cz/YTNIYNIX4OrPe
kVwf08yMhObukmecnEbIE2SM/WnkRX+b4iXfv5OXnLVeB4Dq7eo39DvkNk1/
aUW+rm5XwwWrlht6JZbVJX3/xqyicTxzLJrkkL0XDQdfF6TBQa6hpfTWrfBY
gazLrEvW7fAUfusIUAU48W2IDg6rdw9xMzvMYGu87qSSzPhEbe9lX2puriLF
emZFcNRM+9kxbp2ehc1loGQw/mSRz+nJvu0Rt4duQUedPk2MT8ED6Q4BYJA/
OYa90p1qpt1hbktLCreeLmlZU5j9ASy9aExQLGbGMT05U3EOdqq3ld6FW1Ce
bReZI/mrEKT/1NhM11ds1REqdCCAYFCdOiLE8i6GWmiXpjzYKkJJBUeTVpCO
irZaiV+Go7sn/5+pqKL8DicVlV9mrOk3a6JWlzmMhJO6WFX5lNPcD6CHwM7u
YH8ZYsWJ/CLP7H2yal7NLNbTJ75w7l5DHT4C4iHMmxObj12nO6AProCSottB
mGd9biPhnI07jovv4wK4cGyvr+n/Za8+CuIjKTfhhmwyDcTnDKqn8Bnv7GiY
31lzUnkFI3l+35oNxM58VHIqKxYl+B4yYIdekvipffuHLbs3Pkk8PsYy1Oq9
VapVDVGu1tFTL1ZohVlj3I34oXnNko5jzQsefyjScTiCLwXVru38lh+2Eymw
TnZV7nvvcFbWhOObbowjWJ935g3c7DeveDO8mbxYcK3v7jYpT6We3wc7SrFY
uEPiJRPwx4M8kI4aim9TT1dFEOtPE8PWasc8BKN+9FzYa26oVlNqzmgREvjP
qxGs6M6xC7wQMqYfnGhTj3qrQYpRCPf3/6w7VNWssjtFYHt7M2/qRTVuHWdg
s7VfJcnnyRBkzVP2SeuAM2dN4bJSS2wss4LT/rMMG476zauxqP3GW9igSPU+
Niym3SNOSWlolyIXM+MPhCRL9qU2LYTCK+FInZsafq1gj+U9N4Z9ZqY6tSED
sRTl2T68/2GC5VrOfC8+WQVqHoDSvYwt+egxANe2DEqE4UEa0VDv1cEABnHg
v3JRoYQj56KmZ/j/FrW1LWbKll5T/PV2YEOPxaEdW0ujSCD82K09hL585fXj
5SFFJzVdfHTFEMZPvYJUMn6J1dKfIcoV7WtHx2V/d9wx61Q5ASmrNkLEUryc
XK0IfJAuTb3qOZlqAMzSoVtPOEF0NRNHUefMvVMtHcGS+6Y+DrHCrHE9nlnW
AopKXg1edcUTKHQ8G/dTNy2SoautQoEqhebFDAFHZa3spVcgou4dKqEkIfUH
DLQw9Z0Zz+zg7shnDIXZyzoF2+fg1npNk8OUeIfdlRkSvvzo5a4dtXkDuBkn
AwC2gGClpFqmrccM4zu5MTCJy7jQBIoAMSceKSDt+Q9ELTgN0+UInq2p28Mt
I2yLAgogJm6nYuckuWxj2LNIDRjk9zYlXomIoY/FgrHQtbUEKc2OT2n3IJTq
xjM/suzLzRpK9XuvRRq9S78v90qgWE7ei7J9Mz87o92QIog1eI6TnMtqVLY2
+5ubPITNP9FvghY6GjjHYA2LtdOddcutndRNcFp5FHFLnPB4ORtg93Nn+J0h
47ZJDcTgZsZn4cEkHt/rn35LtUANBx3Ouus4BwR3VURuQ3MHSNiE8kUiBlLC
OkWXg7lBMbWloUgAp9T0JGIwUv68ZMHFTHL9Q9JLWna4FP7b67WLaS8ujeCX
Z9lg/S0EpxStX9b8WpKv1ppXfxH8DF2/0+HDRb8hY290Ln/HsRdQBcMNYtND
QIPay4GMfqvUyEMrN2jIt02qE1trqVVWQT76+jUFGGPkG+3gnuppWYSiHhEF
/JgkAzkxDsfuTT+eV2RRvwyrAM6c0wEVyIEfxFA/R9Pw4+GhwVZeTBwWf/Td
V1j50Oc782JIEoQKiHnZI7+pdiuRuN0dn40Y1yGwlZtIz2/62ONULiWm0uMG
H2amHV3rzD1R74M1y96ysNOlUsbz4NeyZb2LaRljmqe4hbWk3/ID6/pvtemf
/cXAAjl73qWakP6hcWuzrlLGVUs/4gEPWJPgxG7yAVe8B/b9DEk1F4dNPu56
gmeVoulxiAsUxEyiA1ep58NmggHJa+RCKMljPVLcTHFZ/B+ERcYZtzWTV+fe
Zr5hADqVKcbopxj0nRVwiLviIqpTeHorm5vV7NkqLTTLNh60fwROzYpWRWot
RxoTbCzbMrCOL5nz3hOJ/hGcJT12C8bLrhyY2mSaWr5ueBZiAbeu+8I6Xi2x
e5+Qakz+jme2z6dekwGOikthD2nd9VL0HkfeCPcU8oa+EQnt87/Gd4mIyGCP
8oIRznwFyHyBYXMy2uonORV1pVej1qoHQBwr/3AMve5+QkE0j5LwhS/U294Q
TEBAKHfR3isr4cS598yMzT9Hybk/ml7dNMY3Gp0XYm2cBL3xr8h/Notl6ecl
03qX3E83+Sw3wMP7w1JntWMeEbkTRtvEqzxFmYkfVecHDmZnvfywpL1G8qc3
69Iu/4YrEdEhXk+AgbPiH+CbShRglzSGFeuMimbWi/+W7NiWWCfjOvKDKVN3
EB1xX8F0l7K3mfE8NkTI09nTloVbmnUtgM6DcjzV0gLxkZeCCaiDsSsNDPMt
Y6kfwPhMMWJ8ft1elGyAGvbQCbU1dn8ePkM+YterNpuobu7jrD8bOuEKXuvF
JWCAmkz9afddK6uld1VlJqHxVt5DflKnGZ6jONoK1VMYOj2A7YeZx/PbKjEk
MYz4473X8Ct/fsTDjO2nNtNAiGA13b82KOfbrSZ7k8Zi6tCBsh91f4NB7/7C
9f4qj7n40XuLpm1w8zKspRZY0y0UwkFTSgzA0/UuzUR1QSuHAIf9Hdq+0Q1v
D6dKLSfwSwjNAnVed/ems7qjjUO+VRFNDV4kX4t9Y67yz+KaoQ58ly56vXvT
x4eHoG7h0TT5JhSFUB4NG7yP9WNeFxCpHP9nanZr/rOTa1TvRhHgH3ZKMj0R
sGwkMfkA9j3Oh2bv7QGpzGUgi+DIlL+PXFX9FQyqRoo8RRy7ZyikUl5rPjaK
Myp0M6kt14nVJ02KBTHA8a1hQl4JMdI+hCMVidtGqjr3RivxUCxpx013C5C+
m9x67XLa+St2vX8mrvY3VIOCJpTIqQKDTYBs+tm3nIWOJDXBKoQZcsUDz7mz
P39xg3/+CWZFdVoXAOwCSXtBP1j+8kyroDhW5H4AP/2YRWgF0THIF6qR3gUY
tMoR0iKbv1IjycLCuALW9DfAKElpWHSVzgPWIzJZajzBknPaYSA5k0uv7P66
FhtNBIpcdbVtIa648HqORE2jw3FSWnKoFxEIkLHIj8fVGbBQ+tv+VBF9bkdC
XQ/tBD+V0gSjv1nZOsAZz9rDeHUKRqbWuVZBWEt60pDZknd0ynlaztt0VttV
gH1G8i0GytWF+gZflGsFmXhISciNlU26v15MapSbOsc526dVraHJ3iWE0t9X
guBt0Ao1cw87d68oCL4oJ34QBChUyz8j404VelG7C/DBuesO/KuSO0j/zYh0
pObPXJS07k4Di/w5sjFoYsUhXCwCR7RNUTTbRDY7lEwL40AUD4y09KZ5k/tf
HalFbVCOlaRRqqOhnX5/EtVeUyFffuzJxn85MThL5cwnZiytvy+Uu9NYbB2n
DkxbQgKLP35s6oh2SbtzNczZR6h106LmIX6DnprEtj2iO5fAk17Axzhm4ewh
W4+6u9L4qRenCmgQtrtAoBm/cXnWw251AuOk/bpjgEqEfYmBtmRSXn/9WGuM
WiFODujgan+G63TTAsfip7VruzMVxjqSEdRy73bHnkwKsd3EMwg/U7rwnHBX
pBsi0Kcoi0GbVzFOYnk5MHUQA0Wqeutca/4/1s3KI6kvriKdTL6KbDLeY61S
WyWoYrxCvZ8Vr8zwuhhOdXgkiSYsqZiQHBN5Nke6NiuZDROzQEW0ZtJqMDwj
Lryoc83qWYPgkH4sZyhVYIlU7KQKD7DAOJrNTO/LViYbi4dSE7G/i5FfexbS
jaSvv0IlJESoXprmWWNJ3XVQCglM/jUrLewn6gj59gIx2fjshtJMpgnkoocX
sAbUeuVIxSDdzskwdR0FrpWwmWWVPPmHfyMqxGOmYcT8HRqkFtfKhzjnfrsJ
TuIoQc68Utn4htyTOKwfgrzuO7NeCxg59CAo/k+BsEQDXcsL6jkDzs/N5fYZ
1uywmjy0AExE0TzhC30KP96DjIM5J8IBpE602SWXRAHf9H9pJM8z18ZSzd7B
x4l/lvi7hVs0XSgGcOuIetO8YkgrXSJXjYFub3nTCFRtlWpge+NHIZDtvVXO
hSs3+4xTw9dH9+OW+o/0EvNS4igYv24CqM1RJNKTSpoP86lJw7edv5j9kv5D
FY6pHAc7KDfXGvyoZHgPYNAxNp67q+ZF2Alo5IHgWeJ40BMU0FuozLGU26yq
qksjWQQ3cvMZGEqAyHrtk9EkOmy72JRXnDWinZQrq32JPAcYvUzKmtHivOXg
eJTRXCSMX+yUDjjJDgaVDy2knb9GU6wM9yoovXHbhd0vMVhFEhMnNdqSaJfR
4I6cXgI6n8UOOvX9SQFMiHfzLMKHgAjysvfP/B9CX+ipxS4zj+6usJ+Vs0XC
SUUsDXG1fpJOUa5bw7xDGQxcY8dD6obdhm/X0VLKTXC5HYfl17b7Y+Y7XORM
go0CXZsFX/vFTZtehM06Rcr5eI1CSq6pIE9V7xT5wdkFIoBRTI8EmBR4maV1
5jGGs2UWIIs7ixLO+7YqEmN4X937AsdNenpPVCwXBjvsdxDyPSAAKWFdiIsN
/G9IGX6dVTgqQJoA3kDUJTY7MxDReIdRkiuq5Dsz8s79pq4BcINjUslUavVk
JNDF+0uotnjjkCsO/+anrsEqqeL2jqzcJvc+3gala7YsMyideIbnr3Vr4QF6
qcVpid2IT7PQ40hj4H+3lvmnXWd+dyMYPC/q9Xm28tNvUyl8ab2/JPbziV0H
accmoKm1GHH4xHELNt0/bYutjiUWGTIZNqp+zTx1Ew+UegEYa/D/MKJc0h2A
6OTXWiI1pR5DQeUgldmuWLt/VGUa4DvkatPpRp9oCezjr1cPZ2UF5GnZjDxc
ZJkx6qGLQh9xWm5nFI4m1yAmQwWgraCU+Ozq3yIBR4UHak9zL6GsNY3wEBum
mRXqfLuyCz9NQ/jw3YJFhPyeXrbgRPyZF9rv0bCxvm03fLitAXBlPyHyGC2N
QHjUIUFvRs5uBnlYGFwUSY/6KjWjlvr1AwXT3kd+SyARUoCsrkOqbuPxM59S
FAS85MyULFc/CbzetcqBUVVbFi6nZpHN0DeSVo/vo9UCRd2saet6Doj++Gku
pVVhcnCaN0TeTtTeOVvqT+F7UdOE3VfoXVZ+hklCOl0GjXxQ7rMU2OGytSyN
+m/GiN71JJyX2Et/GjjB6D1b8V+DKp3hZ3wTC+Ptj/jJisd5dOjaDXXpSEsl
2hZfpiG6eal5MAfsTZOEBdwSxOZJbx61KxJlfYG9SceDJwuJexCH3NGcwxYV
RJ3fMuuDSMDebbca4h/JoqAbC20L1L8qatAGsDLLnFTSibT1J5mZrxf91PT2
t2gEtsEg3w1jq3In1Pl8aPQ827bHc2Hkzwl9a3wPgmMx8mPhVB2mJZSEsEjV
3exMhX9GaB3hVyQ0YpmzXUbtKgrsucNx8FqQPXkJx5PwGfpXRUM2L2Qc5iM4
BgvE8VPxK/NjNo5f8nvTwENPuD0YdsJPEXNsOhQfV66PVkjcWjrUGFWYkdOf
144DLbd+Z5WVGF3a7DHlPh1uzFrbaGLt2DKXBpsePGEA5IE2mBzGdXOhfMZQ
r3FV5Drq9RAtE/45qXkALzgGJecu31/yurkCtMf1zOIM7A9KdeqRl2+81j9x
eWEdGmfAMR37nDjEc5YinPQKejMBCvaMPAnQ0gpIsI3Wyz2rhuw7Y9zHIJBr
p377M6RZ3aebAVbmlzZhwwEnP3bnI/j54yaah4yql5QZL45KpzAvXGJdWZDk
6XvDNasZXcleRWmwi36DqBDgTY8dZdBRr5yz0kjYqLdra/PKip82pC5nv2n1
o7ACOYsM6hs3KNST7t8Li12Lx1d648qTlecFxtG5K+FydTe2BXc/pR4Pu1hy
zf1EM6k5oM7cIkbl9Pr15B1UPboT1lBKudFQ2N8toHdqqAE5sb3XmsfpnqqM
dpqd0EuL69CLZXww0/jLTtvJPW9EBPCspBUjwZ6L3gyES87eoXil/DxtIxNB
06RG0k5j7i17cQ1TJvYV8JwdaEva2nAtyB6ZuLvSuNzEfTxW5GdieEkyjsyQ
Maon8CC5CY2WMW6DEiJ3cc23/eOdtrHuGLQQPcyOojcD3A/cZkFgmObyqF2Q
zvafBNF6bX3f2u+oCwJ/6L7+g7NmtU4h2A4ShGImHYFhO9mBgW0pP+5BW49A
kYPCSYQq6nfbhilWBlmekFinKskhNY5z7/wf9cTUzgk0wn7vRaMcjWA66LSV
A+S2hEj6+F094yVT3PrtyvuFyNVZHaA0CxrfKhUgIxojZY573XMZPumc3I6R
hnIv5Xk5Zpoo1A5TtqUMV/LqG4+pf4aPXOna+8PHhBRC1JE/wZcjnJ1W7riO
5kvlYLySktLnoLfEHlmn8jZ1E/7uccYMLZEO/4oDnGGphXrqnklYdVuX2bZi
3zc3PIrTjZRW/OOq6c0SW7V9CDGe0lQQUSUs5uSgIRcQtss9lrqcbXQuhM62
9XOxIJawixyQKyJjwgsTiVpaMNlauquirN7fmfJWYURF3xY9ZXuJ96bU25nK
ZZb2w8Ueih6EgALKIffzM4lydVtsyieDQkFVY4f8wIde9g8k+6kIWSpEprZD
u23bJS1KGWJgha54blXhs5tepzhU1jE0rVa/o4OXKoVSNrsgf8R/qTsD2OYV
L/L4SuMpE/a3gAIvHdBX6szlVU0e0ZH64gn9SwvTGcLkvcQKkvxI8jp6i8pg
oSS+Nq0cwRVFBMKhMD2rNH5UENoEGaDA+ioSoEJnj+IuSX0YWb22qtIxopFy
svvGAKVWiSekuiWsRE5W9d3tv1h5PrebvB2TNY1cCnsukXxISc5ePigkU+So
QP6j+H55KLgKCthGf4thY9JfcN1LTT4Dh4u7sk746K+macoNHgG0s7P76kiT
U2FToTlkTyXYmht7+ow40ENvty5J9vfRJRGn7yZiq+IBC+unbd6scx9L5wY4
qekKcyzhQS/3TVnVePxlil8LvfH0okWHf94F5jrWOw0AVgwej0jSpcENbGLl
YK2BkZs1wAcI1qRGMV19O7UuweGt/XFPC39ZFhxNop9RMA7Ac0LV5c+1HFHg
PK7em6Y3RoXOaNZO5zozxNxIn+5yFl/NwrX8gcpTh4hdKocxKWdj/O8pUa1B
q81phjpAmX0VI7HyWpWXbSmxDuKSy8v8wdXY3Jil5ij2AkSEqPTU1L1/XZVn
7k9ReTslQztgtRp4T7dm8CIqMxO8XkCyFl98l+nPP+CW213pVVUr0DXtuSwv
n5p+UJxovhQqWWGRQmLs0j/YelaWBmmgRIedYnyhzd2/2RCQmMfX09ylxBDi
Qdzj9chAI7kaHby6uCDXJWMLvX3H0g9Qv3bCG/X5Nrfbdxo5PfyBMwBz2RGi
L7DtxVTsxn8fA5ZYZrP8o1hnlFahAfWJwcdPa1dQkUml7D9d5Iy5eTvC94eU
nSTrXZK4NNchTPUZ6q504g1diJuqKA+PkwYvDGIXoaPzqglsW9Wtsvf/3iHp
DbkiafRdGB2VrgB7PTUWa3KQL0US1Wj3axLTR8aA0ciZsWeRlmyzLXVeYQdO
G/F1IiQ/4XQpKKuHeqYAG1MOpC4n/3rehufo4zYkW5ZKbMEIfQ9hBl8QRevC
BzRhP1fPbRTbh1zu1eNjXmkFHOAkiA996xzTJc++xNt6uR9zWnTSSNoukoW6
ZRlPF2pBM9QHVGAicNeHjfI0I0xrN82v/9gjtvHA8UNBQ0RVlwHEEejpE99s
0iDrogSZVK7K2NEokYxdmJE2IVXa0RMdfhGRpjL2pIuTxmyQsEAjr62NwTVx
vfKchGBY7eo8/L9pmvOYxB9hTsQsXYWhf6EnwrgXxdpPhcTFxLwmMMJUlJsG
0Mx0nldG6zyDb/bDUyPhp5xfBKbVUlEasnDJM0eG9r1JqmzLZyzT6mvekCmf
V3xykw2S3d030Q3rvoNsCUoVagbB6rE7VcZfeWbcbSM+w0AhowC04JJztVfY
70g4XamJVoBWe8iM8wpz027qWbNFNTWxtCKw8RS8ScXfgKVXt/45rMSqptaO
BAWJh6GU6SHWigX4o+sf0diaQZDfWv7kE7RwwOh77ccwxG4DdC3Fq5o69VP0
CbPVvc9guEtN88+YzkkYaVoq76jRO/0qyc/iDpmS1Fz9fW8ksCXlyL6eUgHD
DjO17pkl/Bqo7OTYVOMIDpwshTrl4M9J51ERFXRKJ20GUW2YDi3r7HvQSF1G
5Oecwr1/BvkfRDKciPPs9LmlMY6XEz7exuHcba6Z7yeBCyY6vcgOuL32TWLy
2V8wftjI8I5G9pNeyaF1NR/w1/pSTL7evVl3YQ3/P/1TzdXpimWreV5weyZE
oSLdQ6TLcpdSbeWbXyFhrroM7IeKH5X6PNcEbfJJGj1c750xZuqPXpxZYLBE
a91rfkwUE0wNHcO9bbgOX07ZXAdRVYoUwikqp7gG4w7yx6lDj0iHof2kXT1y
nbdQKsvmK9XyZCnby78mneRbNAma47tcsZN2HBKdWuxrMIuZMWWhv2OPP4VZ
euibDH5R/8/R1cvMlH5DyF9E1BGZWdtJuVyx/J9tI1iehf6B25zqTrXbgfVL
U1fl1xOAf7J5WD7Pvt066E2sBh5gop2RnJOcsLh34iOOi7N2RWsgHLtFX3N8
dnjfENnBfgtGeJDAzPHO8i7m0sAlp2ZODayOptpBiBQHoMH35Pbz30TFreOF
PamFqU1E6h8Zhmhbq/94WdBwaTa8owl5zIr3ke1S8fAZO3nUZSxg9YNwmo4o
q/1ZKoJxMjJIwr8ZS+vQ6mXoPo6OOo4AQyf/ol107QO0atG32IttpVSC6L2G
MxSXdO1t25bcPjXEAToEKE3+Ta0SAZSk0NH97V9Ozp5PJqSutcag+NqCvdsV
9DpYQqq4/xJSLbn9FXE6usH3x2UsKA7NvfNLR5/+tzQaaZdjBEkL2VssNeP1
ZbB5mIl2gNIYKqQm3r+723CxIqooj160lA2ASMjtqb9pEpbGRiWEv8wQBhAd
El+NRlVcoyllQLf0vrBYpKg0DCCSM6maRlkiS3Wgu7XaFQd7VehFMXC7wee8
g9nUmMCWaZvMcjfZB71Zdau1DI5ez6948dMbpwMigT2Zjl8DlLXip5KX1d1g
yY/TMIce8N0181CFJBOGtHpKKlB88FN78CcwKhSXF587qMZ+jpQcAdNSf/CY
MajwAISxQnGavV21mxn/act53ZycVHymIv9cTHwpmrHfKC+QvVFlLj6Q/K0U
jk8iZh0wTWbBeJZhXJ8ln3SWqIBAkrUmpLvUiJMWJ8oXijzetQR5vdQ+XGEv
x3OS8p43gwVyFdcHPnz3nYd6v1goUyw651b21h+qq7aiR/V1cvXGPclHW69K
mKb+cfFxiZq1Ny9cx2cFrMdGPhp/tU9Qf/tJsn1cKt3bAoyLHPqttnX7DiVM
qJSFZYrzwIhA3N8PA9fB73cqfiCUxmB7/mNB8XcZQgaViUj48SnaWXIfVH+k
gsHLPnXm+hV+CcmfY04z+pnoNj4fE9MHTVyeDVsQkvfBHCmCtS0Cc46ebXwV
iIsHcr5pdsUPfi1/rmIP2ifOwhnpk4G6/rcLKLWmBgw6i41OiVx9Z2E0rBnp
kbSjonp2mgawh9dPXDfnupXA84edSZRgW4KxmDS/xP3mIhCDPKRlqQP9aDyu
kS2zWfjTYOi+PRAZfkNpM8RZS5Kbr39ACxGjMBNTGFvU07WnDMxmcxEND6P6
vuyxHmEmWv2gLeE3afIrbGxba4c3JOtnHU9aYswYKG+buwtcVCDdZkQAiFhg
CZHEHA5GcWofbgMmAw74duIbg2AYrAoXii/hYGEzZRquEVsK9uRG7ZBGa2e3
/jltclJsZvI/6HXnT+1NHJDfpKZ94rQiv6BOMNtdXDicjESeLir71Ljvvnjs
j10dJUSj0VV8khOEcOP+8JajOJMWaAUs+ZnxJprhOa5xXh23O/HoaaNeJvTv
bWTT+EOxHgS2MntLCjcywhwAr51rD3WClD7FlsgofeC1SOjZnYHAp8fjQkaC
2SWLdSGgHYJd2sNx+coaZBVvd3c/M1FaEZU6TBH4qCAweC+gFWo4sHYN6oqX
MS2UELapFXENVUsGODelruN7CdGDc78KvdxMM+6RYFoMbrMQkNYwaL7jvvTE
EM8k4AAWPGGyUZ65S6ooZDwjNItsdagTuanuWlOxEAT6fu7WhddCibUCrf00
7ZVKOcYjwLIAKbkol3/AuEilUruK0uKTO/tpKBGRjMMwEH1p1G+qyajQD8Ip
I2zwVvVNDqgNpPJeFZOhDziiKgNnxs5nfh3JbrPpFmJOWah75S0v9trx9XBU
QSADyEejrTRjVNMtCWqNDooU2TajjDGVfQOEn8ek0HOYZ5H/WjZ1QTWd7a+4
1BYC5V7RBKQH0Qg4/RhHZBEhkwY6zPrEMsAEoVOxOVecICQjFcg8Wn0Z6Ca+
YBE3Eq5Gt8pGvc6RF37u7kcYjnVXYZP8YqDIdO4rspvekFcKLEgItSo4MG3Q
UzPjaaIskxzJm+2DR7om3p2apZT2NbetKoLpg9O36q1RtuBgATsJEVEFaPdZ
eL2n7JYFHUgTuOtize5PVc6S8vMbcAza6btakVJeGRTZs/jr6iW5VV36S8LI
tqnVFx6NyFSw8WpSMTlFMl/QtXc+vt0FLqyelA1AOSpWU5175e69j5mxU3ZX
JBKb5ljUlTDcQp5SwNOBjv5cdGU5X/6altBLEoe9T9ljblL1FOXKHbqkVGws
3+OtriXvTicsy1iO1e0gZ5+GsOn7PpaGlPAeUVv5W96O7b6txySF0x/YX7p/
Z8HFruTOuFSmUM8U0naSgI9i1J8UZHsm74iepvftxjhAT/dUpQ//jHvXjzFD
NOjGm8HOV5exe6XRU3wnmkbsK/v6hVE/64qHXs7OaY/2aEkg6iWiVP19DaFi
fAWO4dHGa/kL5YGc5Wu6DckHQ2Z/UxGmSH5myYvEKIc0Ii2zeKYGKbGWxZGj
e1th6oV5PtOn3fub2evW8vctYeM5ShppDVr+Fp0tSYp13K6Y96zMuZzTAQ2J
4Np+1MwKMcoNTQ941zzb5LiFkynyTl842p4IXYIKKXNEMrJXr5V22oWIhg0q
6azJNxXq4CbbBRSaIocJr78e1k6QBVeVYB6n1W1ofWOYXoHo24Z0CScFAZg0
VpV9mUHAofKGAhwrBZ1p2QdRLolp/xwQN28Ei86ywHJxc1q+BiTbGAzpgarv
6KBWGMTcn3Ch68iKVbeK7mjdY4H7V0g+R+nw0mmdXNNoO7bjnuEnq9dVPX84
GoaLnRNO3nfMMfNMLtmH9iEAIkApy+nFIHnT6Gnh8fR25D16Ek+0DQ/Ru+Lw
y+VKz99EsK9sLaBanSI+bTzwN76S4+fmKwywzGZWyd446MI1ff+teiaTn2OY
uO0S1b/VbGQyX2MAi0ZXZgnHsu7UkF8ZnS9fmQ/m8LyF+SoIPPcClEBWmEfP
L2a4uYQ1OmSEvP9z3qspYjn94GEiLzt7On8YTTyj/zCbkRtdH1Bh8nb7uoRq
U/36xeONxAwNASp4oIyRDE4aspAfmPyLn0fYq1MzLuOwhfQpyggEWMviyjRi
IsuBj6y+t9lvqOLqQjdOMO4nhfbUUAuxrAJvG9zWrQAbtmuFOdgvz1yFAMP7
oJyb8UN7bAYgtwc3SwjUfoUEwh4rTN5UBm6mIb+VUAeVvBTEW88Rnp8Gssgq
gKDXvN2Tvl2bpja+lQrwVvBLFiyRbcmZzoHtXb0LZsOx0lA3WGYs3Xeo2b3J
+RjuoaCFoP/j+FuIVlSEaL+6DbBLmm4jTBYOJ2Pr5H4UycOJ0DAvAioier0W
bXZbd2tZsE9R7vz4aXegCXS3YrpO84OJ6FxxU77dYFnQrxZ+gNn/kQCO20IG
uEcKVlij79IeJKkGub8aa8wxpjMyMFFrdINOS71QTtlqa7GjanAkvYEJxzyF
3kNbnjyvM8wM5coHh1ub2XuqzbWHuwtqy5Usz4Hi5RH4rWVMJ6A0r3mifRlv
ewZindrhdr99dlgxVP99gJCddPPXgba35NVCnPI6qGhzzhaTJO4d+l0chRZ4
i5gBtj9nMAzQ1rp/jCQ9ulCZq2kxWqkJAEgHPRr7q8J3OGpJkjzoonTdFLiS
2fjVUTV8mCIP0lIdgkomqD42xx68uw81Yv1KyVeLO99WVa26GER5dhchHMhR
m+9I/Wvt7bYjNulo3mxQSGa0W6WpoHt31JVlBPr23eeyDKUkS0Oe9amD9uVA
biSVR4GNV+Kuj06LTrn1toxnHoqsnfwH42USHQDQ4BH+meu/xO8X2e3Dvzk7
DC4zIJVCdv7l4VvqrN1iNz8cmFf8nqMfwg0yPL40iWkgrvIOnMe8NdCKCM1p
5mzLWEipZFYjWPCimcx7JvXwlIAiPA4xUDklVOH1nmrdDz0fREB0EgW278X7
+ld4gVda8EDtx6I+SLkRq35UNDSR9kgdFycjGMeuxwggrpqDpjYx094Uut7J
D76LUUfk9OGXV9u2MZgThe2QQos3TnZa9Z3ycXFGeEiuC0nLEKIKei3NVwxx
atBsIgSX3Q0KnlUYY+D91VBPOCh5VCrAglnRHreBMZm2tb46GDSFQvng8lK9
hTqew1u+Itkw4aZSP1uzS5IfhJIBoaeUl6HL5ybhLFA8gMEuRBxkkg7Hnc4x
10wDKd7USX3y8mKedcWHSIX7Yv08S5N3QARNbDfwscG3si7MjP2x2o9kS/tm
kweZysrWk60kk4/QJsd52Z9lMyu2qJXoQ0dcAfT52POaug7Bq5sdPbrYCH4Y
x03uY65c4yh+RfOgfgquUg5kCOgc5sWKwRNvxb5TzpSHFjalrhS2JS1mPXI/
6HN2+Z3jxllfl1UPjjBAnqK4E4kQj1lP2gTBSC4vQfwtzGA5+I2hwTkAZx+d
dxF8RIiJEkDn929Lmg01OW5lQ9O0MhbDWGWTaHAGh0RR4V+uT3VZUtWLIT9M
i/Y4CUer5NDOErOL91vB89Fe3bA/TVlMifF0KWdg+woyukWatCQd7tOJ5Myb
PyYTetHbYXEmzc0wno7ZLVlGm6JB/amzwV9uaajO54zwkbBQtz5K/XPZA5zP
JjJH+IjTuxsxgvzZL8BRQKL9dAKsPWeXGYZR0JIkk1S3CwIaHCTfcjhfiC3R
BT1fOHm8DM9LZMeWPwAKROik9NnheM1596MO++umu2jIgLc0SwQeejbI5Ji2
NSJOqT07kwLNg35oxkVSIhQtu98swRW7oKA1syyXQEDo47aDROqB9Bik6aa4
ih9glrb2TI1Jh1ZcK3+qwymvAQE8GiixI7Ma2k8NHLwisfOgBmuZgkl3m1nL
X8qqv8lGeYI/ePqdZ8loW2m7V2jfh4Qn770pNkQZfrb9tdOMUXYjIfDPHk+W
+Ug/XkbMEVc8tXcm5khhFOpCG2aSJym3oOmSvzUW2WLdfsgKXlJLpWZOsKuV
YJ9xN64ndGs7tvbKSn9KGWw98DvOCA+Uh+4rir9IuSXaf8Ij64tMajXxuteD
n5QikQzhR/4GJf3URxjpuahALOphoyZIV5zcwVXPVXjp0JcQgih9bFOzdMSX
I8Da4dQ2+99qjgIVBWOlJaH9CqdUA39y8wQ4DTMPX+h/eKnsFNCjYk8c8qbv
cytJDaLpsKsDrk5+TJaMlVbXGECVVV1af2dDO30Re+tMWNA2vJ09gVHuAMWV
S48V4/8ZyN4VIkSHZf2jjNivyzKTu8H9UhU7VMvgtlpsDDxZMlTNzMc/L697
ce5XAuDmuzgNch6BOd+hEsie6y74R9jeVuRuUlTWSpf0wJzytm/G/yqWphfw
vFvP1WFmWpMWbInINlsgUcCFOpgaCKT9arvBJ+Y5bopGcV7i04Fa0WR09lDw
GhrYpDNNSzXKR7CPga7Nhxif8g9UpLYZcqhbeiXUUZTgzavd2zxMBTNZkkmi
pA9tKCxw8JXSXQ/aQs2EvHGL67g0wAYMiGRyt2f7HmHWTREU/JzLKPAiS69j
0e4Nm0BFwXDo7mi98Iw/9hsleQLRIPkILufnjQRWdacAgyOPa5HeoBg5N+jK
Vu/zWADcy6hY5CJ16nbRbjBM+RiiOMcAPbj6CSf/QRLcVdk9xy47h+yRRiCE
HXOFh91WN9fM6Com6gbHFHggmCHEYqoQYoorwHb5iN62mEpfxSRwgEWU+WHl
S1JiKFV3fN9tl4wsvlpT48nFwFg1GYPmqBz3gBr2b5JuUy0ODSd2+4d0/kPm
XLBYIbRS2wP/jfHcFCBePFckBRV1KX1mVwcydvypATXNbduDOP1DPH+aG09u
o6JhCFGG1HcMHb3susYtbRK6olaUrMOxuUqSI0y/n+P1eyZR92foIU2bofZz
Z8SUNxBCpDKrGZqXIstPz9mr/EpwqW1UZzPRHFbtKrDzS2fxJctF6qetT252
WZx5TtrHAX/h3Duj6EGJFvniZZM64vClz7HdYhZpPGEkWSahhJSaoFCJExQd
qfGV/IZmdyw7TKlk3LtZJ1glvPnv3vqg4Fsz1OWePC3C0zw957ECqXAlcy6V
E3hCAQbsd4ZS3F6S48XNYLq5NC/eYwvK1qKdC8/bOC3FKvkgi+M42zS/3uRw
YZzTkGry1JagGA5Mf7hb2euZ3V29QkUDy6mmFroDr/dmXJL/YXub7Mp6x2ga
hu3b5uwazTi20eEWnDdj0rwnKAeEqo2yBaXCRugVvnIDI1TdhrLxRpPBt8AR
NkTs15uI2nkJVqVmwHvZQ2/w8GMeITTO4JCxQ8ennp858486YmGRFdHPHQ3Y
jliPBhY89dWufzCx5zlq2Fz+uNBUGDjBNV8CZciHy50MCFbq0TbH2huu6KaG
YV2/Kp4NUfvymKXhBL1LMkWoU6Aod6IshAMap0/w7k6xw7r/U5nhU9gAhrS2
BiuMa1k+b0l6t3ntZQjX2GMkNzgZ4EbZvd58PDKLW+S0X6qk165E2+BicNAy
MNKM+EqsO5O6g1Jhw4AdjHSYNUKrcFxre8qB+nbIsaxibLYj7aC4F+uggfKT
MuT8UvHgvxaiG4F/IULLdlYcQem2qsJVOOuhGSq9i0j+pwiw7AUhJrgq6I7T
VHEVIIMZd3/aJkbI0r78Elps8rpKXZqz181Mjgsa1MjHV5kBJJ9Y7IitUWym
TpfproUhJavGvHGk8helIMmri85x9gqqCidEu+nOw9uQsCt4YgrfochiUmCe
EztevmmhW7HZQ5QIbb6O6t4ucQ13yfgtmYYvlZ2ynT/DfMWm6WbsK+2BpS+a
mk2tdyqe7Wn4LgZgMR0T9SW4AscTtl/zoyU8TNurCFDHBA476boJcBC3OeYG
8u34w85B4oEpZ/XBpQueQfgpXTb76RDjNqQLp0Fuz4U/TWAIPgg4qX8BKhO+
/w0nMWbLUBeQEgn1Oc/n2GWCCzEnUqI1B2+4W8hpm5qGTncPJEVdrDVFlXie
ahREDNjZh/jROJJ7eqzxsUvPza6Fyzja0csnVOOHGwoDlrv7c4spVoyiR4cW
MjiKL4poxBsZBgby8jQbAHAnGIeQ5xOZOCSn+WM8jqEemmFFE7e1iN+SjPLX
O7sUylubbl8JGdd3wVizqWJJAO9VQKvshOiZaXgtmnjUlTRhfk2JxUZfPmUo
8lo3DAsuFxvTPVLHbSEoGr6cv5R87dJVkbdGpzldSdEbNjkSzdYWQIZcewwX
VoJIjM118T8fs+vZ1iBAXyPMoIwTb+Fl/CQX0rK7ksqquAt98GgRUH18inxP
Ws8tZp0VzH+Yi9qyGHrfPw8tMgg+LhGm/o7XGmXzsL5iohsF0wFwzzGt7F22
zhKG0wwfVI7IAklIMPPydVkHtJc60XYSHLQqJONWhWAIdmiLX3LYkVk8se3g
wuGW7/8vUB1MO24qJDhrNByi0imltreiPCu0OR2WCIyBjzeWyjyExiJtfXJX
XImOf9j0+32wpb3KHbH4QTNWG9w9CGWaRjoMoP7ZATU6QQPNB16u4xtoBeBl
gPPvyU44qlp3oQfKbUylBe5bnQ9X6kITDXFxSdwtQX9eF85CB7WMHDk3QTLm
vongP1Rt1xk0auqe2x3R2NGvFhhpAPJL4yESEnB8R/KgmW6ZYhMKwOQdbBts
Ld+vqgf8yGEVdlWaYtMO4sHz6RO6ISASTL+aOd7xjiMUhshOHq5xY3OvQPQB
q8DT9S+BDtpIAseNKb+tG5FDJ3wpcnUNBNKzDBqY2iQpaVur9bK/KiYoVJ7q
kK/MeppoaaLDnFYg94RJTwjI9E9ra3Dhgy/7B8RM8QqcQlxJ8KpoePJTvpyy
VBLM7uvz/GJwB7lywe6IquS7Qb6UIPj4pvMNe4CPHzOxs0vzRqg7Af/14bm/
PQjVHMYgMf/oZBX2OURACUNA13dK5d/k8SuUrCXJqpLlXOoMo38iyVEiJRMe
T4PEoLbLBs3LQiIHzTtSIHVnktxOcM0nbYXruiGTCMRPXO8MHedkqoWeqGSZ
4BJe94CTOdnmn6N4EkMW0E/f3XuSGN1H3oluu+xB0c9frN94FKCgzwsUxI/7
uaD/qISjFsrM7uTynMpM3aOU7NcTDOKDZSgYA/NRSdeJgISLrRvRm4jfRaXD
5IPdsL0JNJa9UFO72GtoJVphWYKT2wG1qwrqnziuMp7ngoibZYjD9hAYcdh2
VAfAjM1Kcvwu/95PoTCDrmsB6RqAreGzeiDf93SAFbEKPPlc+UZZQkoeMdzm
6D0e9Z4TltKpUObkzjGuOdeMhxJ/KWbyUCxNFFAm86XASqLqmKFwotxaV20B
6iRmEAyUzPTmP6MffooCD1AfbTgzPKI73yrgoYpjXZUuh7f7pKma1Hp7vMqp
R7WknDIBYmHuYwfo9Pyo8QUAkX70h1HnrkqAWZamkLjsMam/tDd3Yd5hwMad
wSzbJcesL3D/wE5ZwY5neekQXtpG/4fcX9PpRQaZnKEio3+v/7CAGpffnhwz
Qn6lD3rKI0t+T4CW2NYOaXG7yt6CYCbPYeE5hEd+/ADw2mX5/XYii2bKusCT
o8Zn9NOw9tSR17ns06PrJrkcsroaBbtyWsBo6A2Xihon3zLzHg0cwaRmWJMQ
gsMw2mipuMjs0wUL4+JuJBC7SfzQiF2BXV3Xm2hpAYQlrcyC+QdCMyJIz2nl
FcVUStH2eey4IPPwWuC0d96PJidNsBSmHSlzUPN/q3rXJIYlb0ZCE8FoyNZE
7mfGl2KGUZkrEqavlAcPfLRTXlkXIPYJbhsLDbtH58Sybj17SvuSsV4Ye9RI
cBMHnRHycEzwyEupJ8pNZtNBCRHUouyp0xX8yKjE+8ejF9ax095OwSJB0G84
HstG19p070JrEr1ln+nwX0R5onV5aqDPOkeR5GUHF1Gk+U8tSBEKWcLUG5cf
bNonl7L2jAjK2XMZw+MZFK9zHJ2zWLkwkyMyNuoLFEOhdB18O3QQG9NyDeuH
OxxrA3nr/+C9Gf3xmIDb5xloQsGl7PzlSelKo3mKoahHLap33kssoVmv0Ku6
WTWrW68okjVZh6uBz/Ffr5qJszFcUhrGODTBiPXXaEQRcyJicxUeEKlEzVqe
1NGis2Iwb7PjL6ICAnroxE/O1rMGY6HgzNtwhnv3onXZFPjrQp0cxzf2fQT8
W1mrWVwHQCVZykRcFWvMbuEUIqU5nOSO3mKngt51losFC1fG0rBCg7SJwcre
9mdFlcGmHIvJprTX+p5ILJ7wbqWG734s6xP6ryMIqpjW8R3XONZAx0Lxqujw
8kvusaEG+mbFkQineQc3PSyL8MvguzrQKvIfP80uX/lfQ0+8NBYAnLEQauSb
pzywd5BiboUh3c1RxMzoHEO0yfqU2OVLNGfyt/wmbCQxAzn1A/wIehx57zFw
tPMMjIKnI1/BTfUHPkFna0K2ITbpg2Cprb4/PJCbMs9NwENCmJrdWUyD4Ao8
0SAWNSUp6SjwwPcj9n9IJULb9urhrhsOYEvGBhKv3RcpBSWvFeYW+wbLKjJ0
p36xKkkF/TkouHQOytpoBCG8F5qyxU719GPdiRFD9vl4U7QBcnWYShalykNW
fl5myz61G5ansuJAyl+QIPR3T1Z0iL7Q3R3hv1hnl57aCuSvt7HM7s0MmGsu
Lc8OQo0TdK3v2K7jI9P9ug6NRCw0kj7iPJ5XpXn3VBOxnM+1uNvZPF8sXcoi
6MiZLWXOGb1B/JqwvpTsCaTBW03r0N+xgpY9ChF9pY7IDPIYOHHx8GyIKAd8
c5wAyChSXz7rSaLIOR73AlnfRWRBRrqLGGIfUip1337p7ySlTOt0Fj36l/E/
duawYFUVLyvEX4AEs8me/ZO8Azk3pEWf7XvpsPalUvmZOp2BmG5DQzHZLH3Q
J2Mkj3lesAGVwtqDLJysxjMZpAgOJQiIRhkZUI2vUeXelI9g9UVshJEVGBQQ
eM1xFSORacnNypJkh3VWCfkQpf1fAp9reD4u7GM51EDWFAdtzdayvQ1zLO0N
JPsxE6O0YX1ce6hSlBakVG7bP8f5GdGmfvYjcGqXyuWzHhLi0afjj33dJ7sW
KhlxUn9mQzCuDoiXg13ok37d8E0EujFTQnJSW/nkgDkBII84QEI8NyTL0NH5
aQ/0CXdxsjAK1lex9IbWbe8jd2M7be37VkN4MGnYpJiKgX8pkda9/eeClE7h
4ywB0NhXCZPTRixZKkT2oF/0EtUa45dcIICFHQoPjUq8h4ThUUU8WX4hfwx/
YV44E32C33B9d9n9mdkseir4Rr4YlFn3PgF6jFBT/0RB6nZo32ezg8gKTLwZ
8bwD7zgX1lxMDn6O87GMEWrPl5uapVamx6nKnbUfOmXT+7/EV3lAbGtZpzco
Ie3CFfWyM2x3pMHxbMRNsWMGDWV9PddBm9eCcOoQbGQYFX3O0ojXvYgJw1KM
8xYVDb+KHN4VRhEi0mwIXQ0GVCyfB+xGdZ0fVUs6fZtJ9urhbwKheHXKTkTr
0nHnhO+hsSitE97EZNAoI8sQr4bGLgxDBdQm2TAyslRyMQ22gy6wYm86yBGm
31W9Fzg6963QOmsaBGbl6OyG6/+hJUBMmBLKU+449A3qscTLcoU0LpP1/fT7
CX4+WrI35y0evcEdi0GoDafbQAJ5yMkVcNiUnjG9nYkBM67vyi3bScFNyg0I
g7DK45DQrZu6Z73gZvnWBtuhfdoKRwizWmts1GKYghpw6qwna1mLU/OI41LX
fdgvUvOyUNlq4dLrqxfF1nsyBrzWvjIKcH5wicJwx0AuqcdV93qIm0rTRUjY
U9Y+PWOgdrIx9glM943CMbVkJoUe92fmAET1yIJ0zv+h/QRpjLEeykyDhwtV
A4eNGE/Fpn41eY+BQOOMRaLd6Usl+yJsI+vo6MF83N/rx6BoEPs6YKi4HOO2
N3OT+uLUAl1bjlIMjI/pZs0IIJKEljODcFIjhO3TfoS79V11wEqUQBYnEPpc
nRUT9NKgsdyqy61LsqsVN4pFskiftGUcXIltApKd6tvVqD90MyS+yDB/5xEK
M9+UxJzrRCavhOnf3tNqorwK+QqZEgvEkziM8C++yPPOXuMlAlloIgNYLbvP
YTFw8OnW2nyVrKgeVw/shr0JpEJSubreLW5/wKNaCK5k0BBP6US1EIhshrsR
EVgrf2QRK+ZXsivLYIBceSOfkNT9BB5GFhQEqzj6fjx54HSm5WTdh4zcnJMx
ymPL0cb7Cior7rULJAYuodof6ZgJYLtzr9IJsXOUKsAhCbq405BiwWHMQz4h
ezxlazr939oQ7i7v426o5gc/i8kj5vkTXi1ydIlq3zok4OJXK4QS6yGF/bem
ZtC0aOELmM0JJmgnspGDotvJJ/ydeS8/9t2tYq1eO//2HQrr343XpUb78btQ
JngWiMKq2BVBZMzc4nuo2QJ36SjQMAJjwW3NuHXpupwZK+mArjbZIv7WOlks
VpwhrNwARf45/FoRpGUvq6jsw9BHAnpQgjtTpTagh1qw9dKBFqfcii5ujmLi
zH67jmoiwaZlUrTL9++CVNUH/9LqXB18abUA1ZRjOg3odmrH4sXPNb71/QrU
CA2OMSiEnE49vZiPjj5RgFCgcLXzRmzuDIZLmV8RWM2eOZ3hA4R8zpBDDu70
Ww01vyuBoLBVwDVc8CFV9xFHRMCLtr6gOLL66k7z9CJOehLckBkL4dIfF/p0
87HuJtcKaJ1jkGwapIVzA7+NaYg0BLkQj88IUu29lGPBV0t5/0t/dUMwwKFI
ScxXvU0EJDDYlVvRVjVJiA+I8BkGMkM1Q0Q52Xi71B+Rb7J4cxa05R5UDCJU
361zRusnBVvX2jQ72Qo0IocqKFqW3RgbaLEkUhnAwMTugGFNI4n3axOS6qBm
D2NVVzidotFhU9qoPD5/DL7KCeF6TWrPKuFmSgqNNcIc/yro9pepxPE7Tm8u
Hktxy9y0QadZrmM8y3+2/k9IXD7a2G5IVHNXxIEKM7Z+RgS/h7fGhVro+4QY
WjMK6uZsPTXK18mAuRpnOiZhSr8FXzD04CohpF183dhW1R749QQPb0E0hFLm
h03ljEz8bL/m4dI9VozH95ABR/wdFL0rI8kFeUAenpUFwFrnJNRQNPrLGj5Z
FmXmDaUd+GHjilXQzX5BEAaQMLv1AOy6m1krG6zu5MUC1rTkDxQWpNwe+DBo
YiX/TJxhra+cz28gkEkcMZYYURqA+APcZPtF7B/bEBuhRW/xTnVoui+zAOgc
2GwAs/U2YrpCDNCm/aUDMv0x4byNCTO8y4wPPZFN/1icDgaVNEpqVXThKlRB
UGdnkyicO8KmgnsiOuib+4MHcARvlIZ8Pg7TYctYRMW9oaUIKDHFL7cr4GaJ
HZ/QBOO0990sMj8eqOpoletYfsfNlm0jWXWbWi7IKDsHsdCLf4MxahOzIeFR
Zy4DRO4OWsLGS5DDXA4v3qDeLSqBONsLOj3ivB0tuZ2jo42xxHJYnjISfM9e
hGqqhYYrifX1upPj/ovCrrgfQSwfUzRN+ig2qcPcLpK3TD9C9PXHoI41ixvM
4UzomlzCa4ysOWsGYaz4bqO1ZsaSjZkIfOpw1HvNr4gSWmUMYqgwDaKRiVtU
KSZ+SQKoTH8qmjR5upqOQoUopbTltzAykBgoZOu8oBPKbwsLa8zLGxyTLReC
5YJKOhg6X2GviR+Qp83x1AiiAbNYDeHs+Ybv15snAEPwRzi2pUvItxQ4R42s
XDZgr+nI5B4XCcR8oK035/Wxk8XE9KS7wLqgONhkwMX8FRXme48GtzeNDH4S
U6coBG4hwja/4PLqfdeEt8Kl4rM4BaB/tsjqRpkyjMeOjK6AgJhkdykEVCrd
EyVkqa0lxzWUZIjEDCfs3SA8dvMAhAm3ksY1UXUxBeTYM9NAbu6zHGfOWE1n
HPw2i+zuQt2sijeKJcUkdioYlG74NWzBOfbv74ggQOwiWFGkF48e2YBMVNbK
yYChDzBsQ3EbavDILVopOpbrOKWYCgvQ59dPfkCnOwc+lEeEo0vagt3LR8+b
phLe7A2OkHxfmV1LgL4Bd2h0+7Sss3kfPccFV3IZ01C14+Zpy2xwi1+xlxhX
vmlrQxdgccQRYIx8poiNKTTXPS3eVAdB3wRyvNTohY5h3BlSmOR7bCIafV1m
qW8tMcG6Y0wc3q3v/ciGuZkP6IUYxmgPsyaZFYabaJZ/apujFAndIrDI1xqW
fD2cXHDt73PmpcW5YYAUsqVFdq98X3j2b5OvYEkERNwDDE0j6+1NWWWOE+Sl
8g8IPmxyEUhw4GTHA1VGx/P+9+n8/FxbDCnXYXxQuzQbxQ0j7Vgk1d5kH+Yp
cWy2SRg9EnNoAWaoNO1/voAVV5UPx6SbgnX8qL3XqiFKidKyC1JksWdAp2z8
soPA54RqhKNZ8OKx4QVdjD/dQUfOro/Z+9eZA3Pm4X1hNj29KikgWGXFOC6Q
9CCS1FKqSSZgENJKKDprMgkX5LfK7tS5RkY2f2nktr6IAkTcg30BRGVVkRMx
qXPKL761f66vcwtXuTL3gVGGQLBPfACTHhCg1K4a8CuE2DpsRZzNvlEU67VV
9SLJM8Sy8P62VSjYOWq7lTzW/JX/k6uGX7fYSnguCkCs177ea2+gb9WK6OH7
K/m1L1otnHAx/UajVl/56ToUKfu+39I4ZmgZ/uSizgn0s2x7l32R9m8XKvL9
NfoJgY8N4e0Cv544C7B8THMNDK4Adcih1A0Yo4xkUOdWGgG53KugrK/DSp/d
v6yMmI/Y8IZM/3+gPaUVG3nfnBC2srSnjtV+eeK71Ogpl7v+rZjP5f+7NNzx
8jDGL6qqUjh1KgLvy0hXUIkSpbH+o4RdeJfqIMwwgfVqpTemM+dUz7A4EoQO
KCxYLwp2H02jIwAqq6W/hg/9J119oiPTqLhAemuKs3WOMhIO2+2xwhsp6ntc
665VP+fERM5KhxMNNtd6WVjrqydc2aU3RmSq6e8t9LhCvucRZe/YRni+YC6v
RZy/JZAsUQynl7FSUgm0jhArcH7Qr1l5kjPZiGw2+hn3RT2JAZEG2TNWA73k
R+qv1kp2uZwTHa6EFXKmLERj1xR+V125963wdoUfoMqqZNYmC2izaMyZei62
nh/8r7rQxmeUVjTatZdqZk4Va/w+MgZrjRbP5ZLgZYkEcClRO6CsWPzVX7XX
S3fU32pFMNskodPKyNvhAnIq/fovtdihsHwm2pcNAgFgahbQDuN8vwA7NBTE
YoMy1XlVAZvgNStGoIIBjoRkeWYWfcUaGB5EmLg8FzStE5s9FItZ3FbhOOHy
L5/Dc92Y07hcL4y+ERdUpjZtMlO6N3LMpVIZhv8S7SHF8rxVCk6RbHUQretc
P5ByIS/nh7THg5aQBJFxYOU1DISNV9gtzynMOiY6VPK5Y43ntLb8DQqDN+dx
0n7HFksFfp+XnIW0JDlgDU8wp306LWzhhcml5H6kkolnF1k8NimLdGMjMfGO
XP/O1g6yG/evS5q4K2Bbt2pn2i10jM0J7xDzEInL59QCXUv+xG/2hZv5jxbL
fI9dTPNHWk+Q+byucylFmw1VlZzIjbqbLLXugapLAIGsPbkhlg7FxlgtDshn
ojrst0FKbdDwEL6VvF641YqEyaqkbpfx8XpTfXKtJAONLfhseDBNXeGmj599
uI5A8bse2FNmtsfbpg8Km+kE49h7NDhj8MLTIYKNGGGsE6sEuntdtJiYbBye
TRdSb0A09us8pKLJsRl3fullDQ3z2pKin8b2YUMjLuYIyzlu+BE4BrcRn6hU
3V7Un+yxboVAaIFyf3DgU8gQoVzWeJKwz4i3YCRztqjGPhPRmObk8DHf8MEd
cinVtxMHMdgKeYViwYfA8+upEhw+BJd0SXARPAFINlbulqtiAO3yKXFi+u/O
rJS3YoNebuvGmBs2HqolnN0Qjd3bY4B4EOGSxrlk2Im4JXxYFgX2oWCXo0RS
tsKY8btjAdYRHPgQPnG1XhLRTJne7Qk6iLzaq4lCueH8wD5dogF1+d3nlbXQ
Uab+S5i9lpdUTNORVTLUfyIVH7xk0hbUE0UG5PdPgOIqXh86z3gd8jG7ZCt5
i4jh4GITlDcJ7aRz5aN5jIxjhr+ramBPONQoj9dg7RQ6YJbcxEMkNJYWqGzm
zH4AxfPzwrOGOLUNk28sBggC+eGbBYRuy1680P/IyXuGAmGbVEOgMvCKtYpv
dr6uLUlbWGeN8XZbEcckMH1/XFtodDdcXE18ZeSxCLZdontMuweQtOgnxnsE
vT9RhtQmXZ6C4X6Ax2Z6Z3VDt7Ei1W9D+PRZ0DUZ+xz4SJlVeDT7Dm5+n88Y
jMVLAmKgKIBy45vK/Ko3eL4QZ8VlFpqI31W7jIK3kMidluF5igxjCmRtPlY4
Aj7ZLaiMIOXEFiuV+g/wfBJDjLXq1MA4UMDtUfsRwtEuxHRQayoltH7J2iyi
a88Kb8zpRA+vweSMWUZQwPwlJEQWnHkYR2XWeMmZGNlcy3mklM2LV+B0lLyx
7L0gkwy+guRD7sZlai4vcQgVUGAsI3EpzUvg2yBt3C+2Rbaf49KMhGpC6E5r
EwxLp8yacBDtpStMFtECG/+cKurLOEJOqWVhgluTVtCuLwbopFvRHgBbbsiE
i55qScTiG6/0DSctGxC/rovollt0/fZHvHjONqsF7G2Bo+xApLwTTaxu/wiF
opCvczJO6LdBOd2FCxKUVABN5v5fsV7iH/xFGsGN0ciE3yd2cYQyI5Ns9z6y
pXsAxQMp1JVvmmBEpO/t610rubetsZeMZ7x2ru/bqeU1nu6xZ2JNTtbk0JJ6
GmQylH9y7hYGp9PNG2r10wRrI5sjkT0t2NWDHj0KGZJHt/tbHrGxk14yq/JY
FEDDuYAxnGCJ2b9hYI3pLmnpV+Dl3RvseE1sqxNAKQaR/o4VgyTNy0N+ZmnS
UuUQ92oi49/gx8TMDA8i/WOM/7rUOhzCF3TBVbwn0BzWNXEFwsvk07xqX+VN
ZnbzSqsKt6Fkuk1pdXOijJyPoyFNrB/LV/8ENbUIF8jtDJgGJXt+/GfIZfjs
NOwYzBPN00HcrMyVmCfpTRZmp9qarZ4rJ+y09f9pf0wysF/jGYE25ANQskZM
usVB7vX7TtarsGf+niBxfs55Qi06+bc4cAAgN1F0NP9/rj2HPFxEnnzzNKaR
fs7ZFILNZejlDbTBXl9MBgEKyhZTRwUybopgw5v3gV5SlV1MLMMqAI5U1Tse
vn6hvGi0wWMjo6SdRZW7TbuA69q4m/JHRG+og/Hmuq4Ol85CyCi/Ob4W8MAJ
wGoY3eB0lPWRPV8YyKcrF9fbJFOvLFyq49griXcCIDsDz4gMpdDup+7GdJbi
EY04wxE51mwPu4VFK/gUFVOWInGbAI7nT7see67CiBW5M0mS37/GkKmGwxp8
6PcD/c9PrYPLm0ufvobT/Aw0NjX+I1mxsGQfM42GX2YdtKUsXa4MUzmvvX5d
Pno0oUss5Jl6WTHn2R4XGpTJyuJDsGxlYNlHS39M3XK0BJ1Hz8iuPwLAuwIE
OoyjoeR1fa53W7KMM8z3JhV5IsL6/r2FtQnVTCpOmYgWu/syKJreZYW67T5p
Q+078EpkNiKglPS4Ihm6/7T7gp7D5aevKE7absCCOfx+0HdbDv84UKnNuVxy
OWarEc52T0rLiHmp+mRWsHwt6P11KamfkVjf+1/ujFegKvB/NTerwFBUXd9S
U6JzH2N8Pqjqd63LUjluFAhqofmnEOk8UoaaM7ZQ/JMeK2NHbTn5D403+KXe
QYz0w0fA7SNhtRvK56oVNBwDDpWDhyYZOIW616yLvN1NF9ajiimNVKmCCUiz
wNenyZ4e9gvf0AyE4OcXc1ljhrLhTXLwAZSEiWQTv947dxIghuZ8MRImMkZm
iuy+JYG5AiF3rnYhbfk5Ove8jsJgQCWr6W5H6eQ62UGFd7Vh/EsXRAFcL5j9
zzObqcTFS9g+Y+YoJ0GpawSj6wG/zUyNw2thJNGcFCrB0zAj7T1AN9QuCs27
dxqUl8ToTGmqtB0AlM+UIjJNsYlmNbN/AXt5KDL6qXnaX1fV0O6oDT9la5Ly
LfDkOXRzYX7ufLerP6z63YHJ8nsFDxlKv22raPeoFy/y8vdfE9nUIi4FD8vF
O5WQkzO65Ev9SvandNuA1xHn/cnmH4+rB2qb62iG/nfLrpZxt8mhS3Lrldty
pq1YjK0IiCuTQixSEAqF3gfThNmc7HgnQvfMjpeC2rPbvEG1kJrjq6SYUwiD
Qmuf/u9R7K3AvL+2dwHd4qzhWAnJUfqk5T+hOhhzGo85zY/mJVJV6/HjLXpo
tIxq4K0mmXeBTMgHEZzq0F5rNDzSXRy6SPLLogIiYTAC46lSV11XpMEc6zxM
qHpc7JXMJq5yx0GVzrs2qryWbCq3syMdOatRT1RX34GF06BWs4IZlIdgyPWw
Y5ny1LMxOK+UVzkN/NNqdao8EQduOzI9vi4wh6u+Ke9U/MtSYlWXeyNbDYl4
0ny1Nd+vc9/Ckn+qzhlXU54yMAfbPaCfvkENrYqGu3a+izWehKl6o19isv2P
WTaO0aH3SpjHR8ylSchgsGm+B31jHHWZxvQrgji7yRaAz9PPYYXcJZegaU44
MddWflz9aVevhlwVa2z5ZqJ8teIEiB2bYLqO4Aq2cXzW+zvA5KAXaF1Z3y8i
8xSaDf2qWf9k2Klzt+fMXfrTzuzRculxqCROfmbOiPcRXl2T/0NLumTbUzsq
Ie4d5C61H3aRMiz4UrO1rhiziTWvtRrTbP++3kyGNKq0Rx8VgK/IG50CJFSZ
8l3mxxwVyUTdijt5o55/Waj2RH6HLGHLQ2FqGE0RrMo7UDHGtmtre5XwtbJJ
GUVRJV+CmgYHvbjP3Aiu2B8G8n8RNTSqS2jvc3KhIzvNrQrct/5IVvrdkZsk
oagHgXQ9OXR93ufNhxV+Tnt2lJr8md/r/qeRLJwyPK8cMto7Rp2RqkYMFim1
x0vqEfqIgteLkG9peAp9hptYes2HMbXG6A8+yed/3IguMtoYTA4URw6BRpsA
z2g6TQ6qpbtYHXnVfVCCyEFfuMShnDOs+x2Kcfdt/4XnCidfI6C2CGAc5+LG
YA4jfN6dSn3PLPGlayuKiR9S67tM5GFHXHjEydsw1zoyfDLUcYXmXi6G6RKg
58g48cpW/an8dtVaG8JdWtwq+Xn8sPizDTF6F9x9bHFFbKUKtlRqIuAFtyGA
mYOq4cAtLJQcHtHf6Y2cbHe8WiMEIAyrMGrzVW6NU+n0vh40nb1AgMysdcip
oRPi+QOQyoyVVJ+aoAJ5kZ7NZ4Z4fJSaeJ7zFJ2cN7AD1a8GPQnyXJ0LxOTi
T/LiMVvVM7iBawBucI0v+OiGSF22zH3anYS6rRu7UcAhroedrG244iYj63Me
4MwaMe71tcqLNBNVDccKXeiKs2hDPrABRPiYxpyWVoJ57+QOXsfRPU9BNizf
5ETgV90ccrXMyTZ5jDr4EP31aWLErz4Ygekri2p0LEDvBbX0VOMwsUgCCAMF
itbaIaN7wpzq1y0GvZyGXp9p77mT5sdHeKj/gVdBBdSyTRzy94TommcSJ7ha
eeh/PmqiSjeYrVXlwXZrw5U8CEHT8cW77Qurj5mZl+n/mWb+/u8Nw52+ExKw
zHUf/I+oRh+/gQqSh2SDgoossXiLUrJUdx8hM+2l173l7EBL2u3/9ejjJJKN
2nmmd0An9qTz/gH7lB1giYVBq8eV/k4F2Z1+DhVVQ2lZPknVS4LrNOA5/8NM
WH0zmv2OWOHkx+IGR2YC9VEUSTvo6NrEdXJypi0TicMHHjaXFBpd5xerVM1a
n4PCACf5oE1sJFDeVD8/XvY1UCj/BpvIovMtFhLm2EmE26dzk21O9uh/e/WD
X1vBciv12jJETb2N9JIdgH+TX+qqgMdnVaniHBz2hNYunQmEoRd+IGXDBf81
vFSVOzz/55w5t8y6f6ZPVbpdN2g+nump9qJ46BdPzMYF2eGyOU6SE87HB7bW
8/nE6PsQCAbZxN+Zi0RY6GFBm3OElw1cWU8zl5FO5V08ro2RZ9lkba+lFJfB
deft1K6TQmUr7MeM8wZwGRa960bT1fnQPMFUoLUPd44yS1r6ZSTaPaR50bNz
ASu62iTlyOUfl58Iw+B8f9KUMMNkFuPWXG6ag86kf04gxVkcjZIPngChfKfh
qF6QOaMy0RIk0YyNqwhminFmhKqmyQzTHPWCQW3bbAmyPSP6DHDOZQRqsed+
8n4RHK2On6p9dA/WS01lTrTjYqC1q5jop4GGS8nts2JGIGFZmGUkltWChLp0
OuEMhFzl0sQSQLp6DaLtSYjvnmp9qROm4FzeQk+HlCyoqh2pxASrj0mbmN29
1qiHgGJgXSB40A+gKUsnjD8FgYDIrluMcatRW51cQKEzLB0rvYdLsebQQlpM
JQsV8a9uCpg+wJ2RFiJmRz/VsYqtiMvZQExFEbwJFCoQXsQL48UiTCmAeB6G
JfsJGrMOhcc2aJKy4BpTh8uMdh3GDoi2elnbVzgnsL2DjRRE7+dxR9dAhwHW
fHk7InTncu0b8fkcbt0s0SqtD2Nna782jz5XBFjWUf7w4rB2/QiD4qCUBKwG
J0MzL4sTocxOBWqb49eyGYHrq2TnYngxiB14nDW4jL5bktRNcJSlq0FOWg8d
VkkActYqOvAe2dCLGM4w4gNxj4XbdDGzfa346hum926fnUeO95LQYpAUIMgn
LAPt7Qc8TYN+aFFSvjqyiXaw+sVMvIKDR55agwDqdCo4mTTpAOSrGlTEn9IN
0hxKIgugaIzYNvwGQgNKw8TQnLjYzNA+NjW1XcfavpyXTh9iKhQ5XPbZZizf
pJuz9JBjxyZma1N3/xrkBLPn8PFdMlMxkXrQ/A9RAeri5kbPbrX8RiLbc7Dc
hIrDtpwGAZHv0I1568aH6qVmeHAe86yweSAew07IsBh6kZVaa1umOfDn95wV
VRnATAI8Xp88U49hP+hyPRfZnFuaXli7vLiWMkQvf1fo0vvWOmo+UFCfl59v
C8Qu6aSnuVemRPS7d+PTXpzM2yKlxDP1gLB3+3sYqeGMy43Um+K7OLwiO5jH
WoNmZ448djv0XfWAZxzKqeU1lyzuh4LOxRvjbYOeR38jXfE01L8wLYVXECFM
rjjXYv9I6wSwEK1s4ye2rPJu7oheAVLXZvxEjqjukEfKbqN1eLT7qjYUehMg
Nak84cGBkOh93IiqNmGL7PScH8/0wIwEmWGopD/g6lyhzI+G9wxrmUu5ey7E
uxii2pLp6pLD6BqyzR61DzTtKdfrg3kc+ncjfuQk91DJyEIHRIAOXKsKDz+5
+w/kisYJZfMagLa3MxD1hL8c8vPUll4XwbwJE+KfKi8LlaoVTSTqV6ibRQsn
zKGa3nXOphfoRt6VWcX9sBYHtb/Gy2KwD20xZwWW75n4lum8Vpt2UqRM/bar
C2wRMYCMkrWdPIrsywfQCceDHPijbXYvSQ5WhRf+fZ8PIhNhBaeMC0efHzP1
SdYaXttF260z04RIYVly+6pG5Rmz/GwxnGNUa/ozWykTmyHy/Tikvi/iXFOU
xjZQcj2IGVNqoZOV0BlBITkRSlxEe0GxtPYczFSGOlS9zYho16oNnpFFN734
tA/xQPyWbsnuytsjznwmac/nGLp2VDN8ZS/Hp14dea4Y6T0/1L+ZcnaAinGz
nbr3CxFkX0V5xwuppy/5SycEFNpmP25Rc9IniVytkHFE6ZxoVq7bX49jhV7W
pM5Wsz7itHYFCpuwgIXp0zojpKvD2ArtKPalhXMdg23KUHLaSkmTILr7OLUb
oB1kHp5Qk53a/UK8yL0NpfREnCAJh+KXIIDmuK0qFiXp1Za+tfBj9bq3lila
9601heUJIHBXTLn7RSKyVLAfLpR3eWuSQeqlUVz6xLmzaAck/erMkPHfL9mZ
Z3IeoCk6gHMRmPTWutzVTG2r0tV8WGJXe2u+RdEZlOCbOtlMPcvio4zRoD+D
iJf21yT3MuWeNWUhf4fT7NPHNFk9dmh2qQqg8ePRSRfHNrd38VtSzw1xmK4V
WiNqXarKHmUQUGubEXLzc+xmPJoMclZ/3ZPPrG98BAZ6C8mCX/S4LD5PoPAe
rSOckb+5ruGepdUGWicojOTihKc4UueMq4zpCa9n02Pa1a5QjvuxCc8qyIkD
a8QklfCFtzmIYD37DIl+O/pPz/LtVtHwCaqsFpTaPaTxFfslDru4aETwIOWh
nGy0HejMatPMzhNypdjUU/ebUokeCBO9RKVryirpGfTcBQdoD0I9to96YrGN
LHo2k57GxCRs0MezsBfCFIXtUHhOqCwOfsLufjotYnZyR3bL7qW9QHHe7T+O
9PIhaiUyGCvZdx2y6a6lUx1eGdwAl1HvuOGh05KgZdTKJ+QhGb/RK7xP9Fqk
Fvvkr6hcWYswHqkf0UB5JbI6ua6axAnim0c7ooY82zh5EgzZDdD1htmRBY93
KkbAbrpyAuk/BN32/fY01A87Yk/A/IVsc0GWnj7X+o0gV2lG9N1O0e8lwX5/
XS2g2DPmxk6XgwIHZl50LNARRsvUM7xL04ThoLPWKgHIe4N0fy5dZx6YtDVR
QaegrFPSr93H9SPd5tWqUhVjt/3fKlB7wN6y+rjCgOPWXxsQUmUzuk9MyPDB
EfobmyO5yfXaabpXJcX0pILv2EY5KXJ4bbOWxGglFWdcem73r+MspdAewnqq
8pcdYL7F9ujP54/rjqCk8EXkUtGgrkRlbbplWbYGhRFocTYW1r1jeApVVLq7
9EvVcayhOLoCq/sMfbfpPNBqIR36g2VSYAkhY5YDT/T6GYtY+X8V9+BxoNi3
VmCOLKDFIrWS769Cs5fD95luRDHYvpoCV/LNBYzOvs7uzrCpdaUQ54WIbnlX
Scqoiqa8Dq86yHkwzzN1k0LngxgFzHSu9HX86yUuTnLkfTqDa61hMoxlExj1
tjM7QRwunKV7unNE+l+ZZxTkXZ7+XQPf9hZG94OBiN3ygQvYnU9SG4jjl4bF
vpeNhTPSkkOol7ceG3IxCrE+blHSyN/uEG/+p2vxNWUNyeEcjM+iEHRz3Xe4
8A5QnkNukkTo58/HGnUThMeD3mETXGvMbUdRx1D3pJ2myAqWR9WK2LRKUpmr
s0JGgeNQxRA6h543UE6fpBjSXWJdVuJ3P+JvG4niOHYbMQHOCn4Q3nKsyWsA
bCIc3ow4ETtaqUBlyGb6oWTyY7SMNhxC5EHqzfmI9r3Ft1w/NVHChd5bJ7YC
FBMh0PUxxTp9nNxRzLof7y12D0AU7mAJX6lG+QN7xjLANz+FlXvrV99QtCj9
vBz5h2JGLe5UQrT4ZlviR1LSOCLq3Ea5hK5403u5T4Dhu7jtzQNSSKGy79TA
AYkBSwEhjg/prp54ARkiogIislHTykGzRnnVy6eOr9vekRoOZdFm3uwl3bDC
c9SjWYExBnMVZYIXWkHKEEqmLsP4sTYAzeUYUf4CYcyPd6TI+KROwUFAecZ7
TygRP7QXEVPhjXejKt/fxZ9fqaE997ieCGtu7V9bDKh2jTVyPWiR5d6aUPhc
k7oFw/gI8SvHLzjTSn4LkB5bg55O4VKtQr3IhwkLdWnaAttwD/s3Vh+1pfWl
XCH87K8mR55DaKiIEly9gqySgYy0eTxJlMvXetMUXSV91GA+ivLTEJiduX8e
3Q71XYJaiNieTLuZYLlZmt/7JFwWcXSp2PppYRW6ysczNkkHoaBhjCthvG3Z
HM3bHBQIyd+yrfMcFnycIt6uELynJsTd0ObAx4R/EhSJcf5/JS2XHP5BLqTj
Oqf+v43xwfVTMfemqymKRjidXzT5eFCn2XbZoPng5IbkLIPtCV0u//pvPlZn
qlz344peXimwuQsMneuckSueEfhF9gzm4PYEFxDoJhh0y+9rGeMYEg4394mj
PRCFoZCx3y5kmk0HFfXPR+O4a9lSs74uf19+XMYW/gmQfYmWUGB8DRA2ZYAo
sFWyE80ucSyPzV+n1hZGBrY2MnyR3wIe8QZmlEZebHwlES1iRdPPklX1WONd
wHNtPhg83u90R0dKdt765S2wrzYRPiCBM/Rq799GftHsIB014YTlucTekgvP
IGs+8KMmBprlUNJ2IlAZjwHCpNCb/yDmYWZlVgs546jvrinkFnOYSNobDoWm
bVrDbGDPAwhnBL7M9984igvBVqoGOMGPjjAR4qkgi3aK9JmhNjWl4WxJCewb
e9HHNYBYW+6CUgWzLPESvjkRN9v4m9yNlqCPxv/i8Uz3H9uBCg1fLUOPB6Tj
3Z17NEeco+iW2ptnCB2gp6a4t2by8wr2SkUH2quj3H0DQbkIbn43RfZZDapE
qyuHHWO659k7OKEWj6vgsnYJjpZNqE1GSAn9oAoYzenYtgiFLhG9NxkO6rrl
u8cufopmS7hDcU4oteCNYtW1Cbt+S4p6BzyMXoSODLeoI+anNVTWvUG378W1
5Afv55fKujPD4qgLMwlY4GvpXe8R/Yu07cVEWmJKRdNzgVv7XgsAViyRaXh4
Did1Wf+vsWbY2GbI92eXr/EmCkcfIYz9VpUFzb9SslFwPEtcBsTuDOgERGC7
XN7xOkq8opqFEBlrH3RlZxhGj3hIOfyJ7UsW+jbbCcmqmWNsEILhi1C2S1Ms
03uFJm7rmqxfUD7oqfvygAQ6oUoBmHT6/3MW/xoTdxZexdihslDKaL0Q7rJy
1Shh3+q5tJ4BBosuyIhVa3tYyBDln8bCoj8PmoPPxSmXnTrF47aAGZKB+ADa
k9EsewpBCtK1MFvk9ee2kA4YLMg+LetMvtoAlYPjZeNcsNKXSPwmQ9xxKBx+
RmcOUOj3+QI5Qm02VbdrqlxAsbXejBXftQ8WfWkRvi0BS/E7I7czjpjnBxDY
LBUnM5wb4896yVjaUyrMd60LZDgQcKVw3weYrnFQe8sM3y6jxh4je3pCQEJd
rPtCy2K68F/WbFxnrCoPO+vjcGt4JPb6u+oWA0APivuDyzh8Jp8AlT4bRH+Y
xENtgY12nnZwGF5PAsfMDwe+VTJo/KNpwHQRrumY8DFJYzPJgevG+NglpLdn
UPqfLVLCQXWvaNaEGNRMzhKx7M9NZ/SXZ3kgH0pwNjK8UU2HOA408Wcl9vea
imZGps+7VqSnPBqJfUDuIrURrj67opmL8TfWI6rpa/BULXe+u1awprL2n6pQ
Ah3/BGXcHkWndVv8nasGK/XvcEfKQAlOAkwPTn7Wx8OqppHKUI34AJOFqUjd
6p41EHkx+4g8opm7i+asIC41LexgzvN4i5h0emCUGzTC51GWqwNODwdzjU/s
0uLPQRE4FmRBV+rMIB0bdDf85WX/J5tUh1RQpohiS2YyFZDBBowFDDqIq2rZ
zFAexvOvzzGqPw3YxZ3DOJcOJNb/MdDZOaa/1BVwokxgXZ+a/N59UBISUEpA
mhRnreTmVrZCtngLbffNvNVKBPIA/7AAxBWE2qqB9YSN32ZRsGl8L6qYxjMV
iaiYcUtc/SaB+ZOncnrwLbi3xA2nGggTxrB+aebAZTbBrNB2kaCnGQ5+mg8b
6MjV25pXG+1y2P1bfldQdeMmBVe6Pw68LejQcot0Dx+khhuOnZx8tuRTbYk7
RROtISPPqJP+UvfA8kA786V9QyBgcyUm9sNgQ2La137ZymInL2NTx7gjOBMe
fwEaGClxdQeRziUu2cGZ8ePSHvmM0PaaCVdhUTwdYE63aSpDht+R9d1s4zDL
M4Y7C0xNLWLtflV0AQfUNq+YiDEGksxuixX4kFd3Wv0LRMMoAnGC80JESodP
Vab+p2anPW0vGmLwcTaRQIULjom83e19l9Trf4qutOtmX0xCY+ngBIt8tRpo
t2RzXxJ8EJkK8d0G5vwYvQyiTH9L5PlTmAi2Zat8tps80oD9tNqXswDyM1aj
fRuROtAc4NEYGiw399cpHWW7KHTVfLJ0YdoNzIzIFDT2XboWqtup7OueUB2O
bdRwUoTPvs2EySH6RQClNsaZe6DqPlDT/XcpR9/XyQ8Wczq6nsM3sAJX/ylj
A+kPypCgq/4ePyCauzmsN9Y1oLr+CedVD3ABKIgEThgoJWo7XBlX5p/fCjt2
vb/G0FPhDnavQAdy8u1y9dzh50SV/reJiBAHZWHeGPF+19OUpWoVKbF2VcFj
WcxB8u2Ak+WeCb46X2a0NDOGPvLWnOpvDYCcam0AmrakJlyDHEFQttpGdk/o
d2W/mao0YCOJOrW7DPL8jNZySyzuB3i+XLhOAcDcUgFraC13WreJM6gyEFqW
hYyz+HXnM4TDgzEvLQvJl/mLKVfHdAo7E8QvPJxaTaZ2RiNfQv6OxHGuH9AR
/1i4l9IXadwApeZVh1CYxFnCt12XyJfp+e5xAjHediE/2OwXhKkkwkbuWIYs
oE5vs3xsV7xtcdl764Z91nVVFbUuWFVeJu0tUe+x4kl6FxlPNwJAokvSVCxv
NwWsnHUTyOvy3NqyY5bJ0W/oCt7vrqDB4alMIF5bLkf00/AaP2UIfZBat3C6
6Xqw5tycVncyw/pcz3tfsYruwW294RPMu4/E3w13qP/rIqWc/cigAQFYMVVm
zfriE/cRvPjd2AQTfgUucB+6Rn8z+SfY8O2+QpmPJW0fmm7rg/Dn0e7b2xDM
V3NXe+fEVLqfu+wxOUtXv3/vr+M/5GBxAxwnDGDTJvqeNmnxGPzrozYWITu/
AfVIsV6fos3+JuJnQ5tH59F+mGVOR5RFt11Y9Q7pkIwj4Hny8ey8CGylAid8
bIWuO/0+csUqz/+t8tFSLyG4LXx5cl2dD8CJwHkL4hWCsxKmJw5AZRolo5O5
1siqK8qgCDalooxUdgRBDMX7PBe6RtwrvWN8lEotkwgZwzDb1pu/ObpBxhlt
z7zZz4NCduunDmIBGDQsrx3lTHXB60ZtYOQS02VaFFRvCrybmVaissJ4VkWF
tbY1AldEN7IseT7byV8viYWR6GG7Gvgqpr2bPD5wX7puWU9ZVKP4kQmkLXJF
mKjRvOTnkld6rMvbtfpBMRNe9+oAJt4zsLK1HlLe3CIW7pO1/87aGunB2uB8
gSGUKApisG4zFkDOEvPKE2b22rbmb7LorYl3HZZGF/XjE9QenisQiIvKFYx2
cvnKOa4XAGeb7PgJpIUKTbaAXqgHAAg9IHC4qFQJvDn4jFlT1+H6EJLylZZu
AzD1ycN6kbKBcdsKmMXB19ArLmlJCE0ufCMbbLj2tHUa40hSnm/SPNfTwh3c
ZieE/eMPB2yJPBDD7/xK+xzzMjRIyE2z9uoDEPUPPCueGwr5V4qFYsVQBMDo
VGkfzGISTQ5Uw73qTwBOxf+hR2Ifjr4GLqitpkwJpwBqoCOXjgc6uu5CFvml
Ny/AgkTrJQ4Z+6synLAEb/qz7Wz5KLC0ID0cRA3AXEXUFkyxmer+rI+MK7ZC
/Bk0vy+NqWOOamjFx41KXtxsjgijRKUQDHd0iwu0soQbDdRN/ewq/D4kQGJm
f5tW6goewGcSLc5EPlUwU2shek3s+jIxZu0pW+vCInLvYiAChUVv9TWVUKKg
aMUe53DVoDwoFXn3Bm97kfzIOY2WpW1nijb5z+ybnmr1PE/f2HddTRb+HYKv
5Cx7qD+KPimdW8k5VBHrOIPcOoo98uML5vYeG8EWv39rehz2rt6Hr7y5eogt
j09uAcT58HIfYhCN86ET+6oX4O1trS0Xqkl8MxUg9+Qyt9kSz7AW8FbVPXWs
8rn9Jiz+cdLtlHtALgQXJQ47OQYemG8AFptepS7a8Bt5ni9UVLYFHhT9VLrI
mR5n6ZsfVCxC6T0tr3RRwHUlzgPwbWqYuDKBimKAsBwhaEGB98/TcRBq/lND
dp8X6PQL2pb7cc18qkmKpjgbkjS2yvkbA+bj91XCR/prKEQnRtyCg2b4ooHp
hPg2wkDDYaodIrwKGVFYKao1LEySdeTIH7R+EZLb+KvUkK4maXltJgyVhyNu
ZGJ0pY7A+YZFAvIzgxMCIhCx7rdsn1Vhe0R6cD56paIeG1n/ZkbP7UzHw8R4
/dMFimkIEJQZnVuCLcCzrWa3RiklZOXWFDE6f/60w98e6vQgH03xV6Inb9gn
xvJihYiEa7VsDNJGgURxayjTb7Wz+iVQLff/rc7go2kUJ4wYAXNp+6OxMAk0
umD4XnDFnHlk1MgZspblPYFNbiT+iCdLn+Oy9YRtOn4S0YEqHbvkdH4cwtC6
gBaMzgm3HB0YfYRpehgIDIhqeBssOTVUD9pF27Z5EB7Tawpw1yh4DdowjtP0
yqyakSaidjHzTTk20yeEMSOY2ozCfLQArckUjxKqXRaEGr6czqnPg3FX6dUK
oSgWmrXNKpgucaaFI4VI2nNRbpvZJGxKU/x4N2Ux8IFnxltslxhrHK1/GOod
EMY0r5FPLSvmfgPWHm5Kmi67he7Ropubmk3XYesXan/5ZSZKummZCwaZCAkM
Z0qoynVu4wVpt2UJmYW4+w0UxxervHGkEz9uW9oB2fUWnJXSO/Gt6iMu4IeO
GI6/ejzeFWpKrhg9jtmVgvBtCG+1ptItG/ti31mK58LO3AgpB3U+9XSRmLhe
ai4oVj/Ai7juZBFvsdRVwr93UQ1y60G7gwEAjR+Y8nxqTvQCiplXnYtqQYX7
yQhpmINnUNEYccUZVpxXDQaAD20Ah6yp5wCYKawGV+txYWGFp7H9nfwt/rZ/
zV0KjK+fOlou9R1FP1DMMsiIiNvh6uw9G9lkEVds32lqpBcPUVg8F+w3BNI5
nNGHXa1QeBwL4CJ9v74NRRQS/qzWYzQTpoy7ID452sk/H7Au2K8I5KsWgMsI
6L3mrkenzeg0XIUa5f8+l3kuaSrlZJQwfkiFP2AVHtNXzmIVx+9kx3uB9Ku3
XE3nb2HDikzz2dMZURRznDPkxfeanftrNOGPGJ2vaRx+EcXGLCD2bTkYb8IV
btmHQvh4Cd2yyPKn8Q9AmCNr5HBNBalV7MFPCnXkZrvO6gziWunXVtqPMEqp
mb6Chk7w3RU3HobKnpnQXy5b/AGEyjBE9xcLtK03O4gHKjOSDjTBW9lH63DF
QBKGdxVcMlV5SWygnflf9ckjrY7f0rxdEx+qMoOzaS1vdIh3fK8qXJdW52vr
70MqtMg+ACnrVQUcmSVFcvrTS7UCV7noCmMclPP95HZLydJT/O4CX2KYTmTK
hPILigvqJD2gyu5mDdTP+84LQceTwOh5vzS9vR/2yAtY7asHGSKHmYghmK+H
w6/HodA1jxK728bv7BERxXEGm5bi9ehsIM4FSyuZGUC8lEhmzVhk5L5ht1Mj
NHN5cO8PYBitOb0NFa/bXHTwWyBamoVrSpzlt5YBOYprt5z4s/MLxBb1M+xb
yI5p5car+lRowgRjrlxPbxpIxYSxKXxpyQyqfzX5TSWlzubeb6MOKLADpKwC
et+KcHrM25IgrrtOWPXrLBFPtaUACk6MAu+VXlU8gX9Iw1u8RYMT4ZzJL0Le
8qg+rtgf2RucKNdizr9Ru32G44nW1VUMgJSTvWSBNajy2uf9sP+aGZkJv1Rp
POtwAVEIjBhSfeOswP/vHEA/716YpRdANTHME5glmuUdbvBT5T6aU9gQdTi0
kUDWF0XNPtBT66IfMVqFpdHTA63MhFTpY7kk+OFgTgWHoh3H8Np5K/0UGn4v
0vm1uxj3O5DTfvfFm/xxSJJNrhGd6rTnSYANRavFJJ8zG4/ThBoBgY/P65db
zIVpjyEN1s9qYyPAjXWyVUQgDOuQo8yf5QYn/ERuLJBk6PBV5SfotYvq7qBK
LUgJsE64RwWXZ2Zv+o0LwFmMydItDUBx1B34O5Kc/QeP6sLWSq9L+lfFywIy
wb7rdf7Jq5r2GGCx5LubUWNjEQjM23uI3iwbMDdKRIIzzbACoy4HSvB/shn2
WH1/yUJW4ZBRRNG45josdtrfJCUX+QdiVcz8upRiU3/Or1UDNJhcy9u7wK8S
Z3Y/lL1NnNzCp3GN27rcKWMGfRWwt52K6BWWoGh6TUpx+md99lmW9BvMFt93
yC3ttNx16PTjb3tHW3FbMvbRjAem9c2c9ALZmJy6HTZsrkNuRq96akA33sib
806d53VFLPlewaL1usGqL4ioXb3qb2pd+ulJKLipJnsaVffG7U6h0UC6A+R2
l7wbIxvYqXjImomqMOfXi2YBPdQMUBD8DdcwNPMK77Oays725dSTM0Zxk/DK
jitz1ybo9TaaMOx15OLZHpwIk62uPxfqA1LUHzgsIkHdvpc8cYMiNhMdBasr
S5xKOiwzMHuJ2t4t8tv4el4DPSydvFrqqbq7MZxVl6vqkgSdv6tVmRlKldOD
jkkKnjK6K01yq1WxQrNMLRsWivUwsdo1Fg9qkWKiSrzz8E85C3jTLJMWF7mo
UX/sb5bhNFuQEPXQ6df9SLA6rJFMfOswDk8O+hO75gnyRK1ufYiJ55DBf2D0
zpnwyFc/sDzJgKYiqhpof9I5XyPvGykxr6o4rVbRdgI2cBUXqq3Tvb1iTPtt
9O9yR89qHRtDTVqp2tO1SFM17yDGP8KoidKeIts/bZY/npzU20Wt9vPz6Qmj
HqZnSNfxv/jPQXXM7veh+MFFeXx5APxTTEoUaYeU3zK2L9U6mSCyCUveaFZH
6OlaA3bmmi2yKVHWPVqu7byR7PLICBcpSpj5jOE+quPr453ti2R8sC9r4gdP
Ovp/xy6JzyeWTWzBm5KbigOmx3G2uTnD7Pb0504LktgOcCNWE4NyVeigU8Np
rGgp8AoTP3FzlAklOqcogvw3BF2iFGBwcsI++vwPXxwcgk+f/7FQuHN7lhDF
x/9cto+m2k/FcaR+OU42Mt5ayaqHJ6lrzdL1N2GKxF3NIR3OvG6ARpAxFhuA
B3sqJOGmXZBi74RpKmmWndR/VWVRxE0SzPkxi6I8WDngwKM16krumoXVmRW9
+xhKo6NEbOEca/1RBODOq1mhqMMS+UQ4crBI+2plddu6ngweF8thCFrhK7Vg
KD+CjD7HIfrT0UxwZqYY18kAoVHEUd792qB0dr2iATfsyu0pG0dPVGuW50df
esb/Q2/Vtlr3vJdzG1okMv/N+u5tAWPV8IOQJceuZZArNqLqvBbFIX6JF+id
SOl6pZjxjUhnDx2m+EIMa7KP+GsG6QnhGbm0jasCzVolviKxCQ2Vn5FqdNYd
QgJxpeeHmD6Tjoi5FsdeULkW0GCCnR4S4WPym5QD9sRyi/uffA5KCU8yN6PN
fHcWkk/ov9E1YsRjBfqmrUz7Hrwdr3JZKwqqF/SVIt3J/80cr1+bE1Lb/dw4
cvSDAmEv5YN1Lo0ZF35h1x7KCaSB/e4EoARPAlMUPeGBarJxtu/PpHZ2LLj0
d28n8Cjz60BmEbr+TjxvMKgO1Df+H1Ie9/4F+4DjwC4hVwMA1jj3wRHaZdY2
ginTkZ1+LQxrG97dHBfju6qMc7tUTzWlqR5sC4gLQJG0trxLyMxzmVLUXvrZ
wlpi+kjoweLRvO6gutWhU5bckgliT8uXJCL60boo+Neu+COx52J8GcjNha1a
BmPuiYqLTM2pQgsw5kjOj6co+FfKFlEFrxfED/EhDrGkPe7dgqlYKNdkV+w8
leB3vOb6OhUU6bxY+ptrrwve+QhIcmPyliXDGVUAypBpLMtscwyJWmRbGPrB
XGGjAHRgEo/scQyMj86ej/hRCW498CUppaLBkQz52kLE1cuNWJbBjT92GZld
TkfeK1cJ6jAmrBEj4On6cuaDbeX5bQ2wzjMJfi0LUQQ+h3sfydSOuFl/nJix
5E+Bibn1TjtDhmj/rB19xTJ7fHB/3owY5zXkeMMAozfmK5VW3FHXjLbEhgEJ
YAKoD1PkOLI26phoPhe5N42f2puPFPUbR27EdQ0n8vx1MoCZui3qA4VMbDEo
Ac42ci/ShCMFomq0UIQFBlxn5NIZVrxO6hrY9UNM4NlWyY27trCX/k8XkEwS
KtseDGBn7FRTL9IHPZgHuF6qj/wGvz/W81SujKN74Y956BpErqnuP9CcvOSp
ED2f+AKpXuK5E6HXBs7czSNWLYRlAyz7uZQXUS+9yKE0Vknlu3VJQ3M1XNvn
eTj56yFsoc9xW2nz5cKyJMSr9tRQr/Hf20yx/93hoQfE6dOSYPfpwKaBrq3D
34g6q1k+F56uf/rhvuKw7tXztWMFuF/wX33Apbrrt+4TInUnPCi7uomsS8sE
o3szRYPCD6VllFYbrFdcY902HDQgtx0MXhdYBJsoT1bLMcZOYWZuPtpX6Dn8
JfAs/2T0cZ0U4vt3seTRLpcA5qrm6f2PCBVE/Suf0Jn+4vf1iS7AelXryBpB
yoIuoq4H+rvvmCRGeUBjGWB9cDa8J9xvlsmm+Dx7l0J1sfEVnjbsJBlhvYo6
fdlNcP1W6ao1q0sqK30uJD7f6We5zy2GCYoMltJOqIqvv68/81zWxmG6+Bwm
xebF7uSTHglGSflsSzt0De0NtUPFByjA2mc9DL852U08vWFtFJRDD+yJPQAm
XjMvsqk6gOdfvbWzldSNXC+n56A/qzNqrTaFdroNQctwJjVk5ZaZTOK0NbjN
edzUiqB7G4bzzennX/VUVXHxP2CqB0N914fRBPpilaza/d+gvyGw4v06jQXc
UgO8FB7rbjpLPe3tnPXh7cSHLCIWMbEwTKXsbqn3Sljgxk3z76FkUkomS4DZ
0CanZe1soK6vKufrxWN2XFfEUFPGu17QSqZOfkDBWvd67h7nU2Tta1Xrhzh9
fxEK+StHEOtVgeDFxj7RCP8WbmxQxep0wHRPHYLgMx0cY2r03RkCVVzuVEHp
BHk7JILnprLZKNNu1jO+bozUoVj8X9sCGD81xH6D6aZ4MhXvuc154QVWoUlJ
GPdoeT+RtcS0t2XupomAMvGXja1vrbiYIlhlri9t8M7NV/ItYsl5ZF+oC4gL
psBCNmKyFaP3ZQD+vQXFdOJhAiLfxeKpyxXHlo1Humdo+iaTBusO6BTAduDA
dhFQefRJd9s8CG6lbiXtwuNDTLUM16H7H6QBWfwp6DLvVsXNfDuvD1ALxP9Y
VpCiNjsp77f8V2fOfrVyhWM3gyQeU4tTQ5M49gl5nHjc7KF4r08iAG/fut9m
ZjCgR7V1miby5TQmHJhO3jd6kl6LYBiygiDr02OId/CdF++6fRv6NIo6E28D
JcLpoHBm/DYcCFVBjVLp4i+k6JV0sg4q7OD1GMc1XdGWxXwf9/fiZtfzcn1y
8F7ivULTSmVzIdg3GFuXqugoShN4TZeKG49O6qF0Hnf2QsCWM7tBKQK0HmES
GKwZU1iuASdP5gxEZjn0Hv2gz1LE08cHVoh5obRCyycSJUA14EfDwa/KHRnm
OKmuxRozjxTPgQiju/Pq8nJ/wNxDALOHMEzWMG9cmT6Dnd3B1/TWGu8xKPZH
E3NDCHBQ6AzWArWDIeGMnW1xlpaKHSj+KZtvlEj74IHkIqdvcTXPzIPlA1/D
fqdIkJVHWGRXbPe0FJpq6cixX99SoCjX2LS354ZZ297E7c2+aDhc5Lmrhbyo
0tJBeE4ZXzRMxgDXq5Q+HkT+B+A5lk3EGqfYRNtzymjZx3YeSEjWn9uhZQsh
tg44BVzFzkkQ2RtQiqSxCFHFd7J3rVx4Gh/kqfcLUxMfgRIp2ZzJq1JwJvjG
uD5LW4+BUQz/tpxnfuPT7+bXvqusttOtP/WqjP6JlePyBI6MT9Lt6ZuQrLi4
tWXbt6gJ/D3jm2kU6ftIFKl+9FjkVUCub5eG5sp4XusaG3iETh5v42iQjB3a
f3+vKYAJhA1BTTQc2XZ1T/6F3XFe4QHz2LeqwQn6fO1oSi4Gpc7q0vsM0vCh
ssGItrFgaSbEw2lPLBMIid7ENdxaYkpPNzDEhKZtrvbyfgGR668YK+r0zyAE
KF/eQRVC+H/rVkBFZDfkMnb7Hl9cnJtcvMs2YBbUOJS+b6ewkjN7B1Gm4PWz
084Xm5qnnn8ugRltReiJhnN/NF5ITlgB2ndclT2EwUYOhH8D1FabIGaM94X7
n9BRIq1C4RKyKQr20mLM65vcUH0p82k1FpHxY0xS+4N5PvomcUfRHNslz7sO
L0TCs4ZA76GRkc3xvMhiVOcaDrQZV7FwCJCfkY4qbx6E3UIfxkX4i1oTk4Ha
FpTYUVS3jDT6YK5laMORKrxoHUlYkGXJ7rO/K7ZOMu7hhl7N9pp63LZtCmVL
VEZkm/S8j69qzwgAmq9YB78ZedL1hRlcpXhOOoPNIQNRzuYLKJaayKh17Hd1
8MLoD2yHicjlpeEgwJcp+CK8w02TacaY1UzqjT+47XXXS7iq6+j5sqXlYTke
mQNPqBar9VBZTuQdYvUlH8K6tlnMMcNnaYVLeBms9PRUHwFnh+hup+4vS+qa
C7aU2Q+jJbsmLbIM70Bk+jR9w1udnw9iuvDQPYym2Xk5VuViFypX81L4RdN6
S46ImDP1kUYr7o/1FMUTydKuBf6IyDuXd3RxC6P5k2yNc6KrPTwY6E0uvCKq
SvRcXt7bEryNWnlcqJxq2XP8OuRkNR6Fl9AKkUJon+3saAnS2AQSRN2BczUS
LWq9lGf5y4pSjnmjqLQ61TTo8SsCKBusGgTyxVyMOVXMoWh44uQtsa3vSEPo
ytsfK2tCDus3fZ2CVRzFZF/rkfQ2gi8IOy2Oi7pr3n3UjGd/eo1TkHPKU86t
StOxXqJMDaqOOc+qvbB8Onf7cYM9ITQBH65z25NqpnGcVRCB1WYk2Cl1i+0D
iXTgbmkONA0+D62547croPkBIKmOlzxMCLg8ZamOhi9dkMldYzqsfKad5wi2
G+mAQzWF4eAHpcFl5s9meHs5R9Sb6Fsfj8QjOgTVKmFPrUhtpYdftRdZimBU
V3Z2CVJEjRspXNvAmlIiSv1qtP3vRb7NlYVtMRi3b63HOn6+pc2qVzQHBOdC
S1/PVtl59EgBIxPZ2043w1wf91v50bpXJ8+fMpTBe4o7fa4eozlEfEW83bNh
JYIR5mj4toUResIkl28aH6puF4CcAN0f5ZsnkGtK2H4CFfjGXn47xcBEbo1Q
n+2gxBJMTi93b+M+kVKMyZX6pP/7zxn/XLjIzLMpJxgdldYZLklFTvTMa/3J
dA7QCnmenMBscao4BFef8JyvYuP2VEfH003kTUukEv6jJM/4CBjDXMlo4h5W
ngRtYG+HhghhpDoPAeu0qApPMlwOOcWVpYxQRgnDgDYwSgeAyZtr3fiKVOVq
4PYaPgTUSTPm/6wNYR9v9sx2lSBNl00X3QnPluuhrIDwZaHhWo6p1iID1PHI
8y/EX5sW2QqiSiVxrXfrVsFhbzJ4PZhDtoFIlhsP7YVGdQBmLB22EGOaKs5g
ydkd26aKu4TbDQGN3N4G9wfFblqNbVhH7mPGijzk9knDC/bQAzuvn0DC4BnW
W+bjpCRtsE7gEwpuaVLhEybp7rT4ByUmK5NP4gGjQM3NlCjfCGyCaL0fhNk5
jeM7dM7MZRjZ+VtO6dNaxrX8mP16Tp+mScQ1dh6bMzjdLOSnGc2WdaLXNf+I
yCjHAzj/+Bn7Jrue9QXicoFqYyHucbDPPlVracGRMza4AFGPrEWVO/yL3NB6
UT2cXGT1A3UTKTbhShDGyHUED0OmdVSfQ56tacFvXJqgzC8je5ygt9TSiXDg
E+DWhmNtoD7iWWxCb1ARD6pM7CaFOirQt2G9L4j9CkPD4Ff8GtuLVEvGB66X
BGyjfXOxDL+qfsFnGC2PM3Cw+qFh/STHHt32F8TREhm4iTlU9W4Y/do951X+
NZc7eUvUhUv8Ub5CJ1JJYsmZJYZfm/g6oVbTtsNC9EPaJXtMm9K5EdSVM/VG
Y8lJ4hB+y56MRuVOsgPmw56evw4r2b+jGSnE8XjBaxYA5fjdlcyRwZC4PpsT
2rzLwn1xHVHiS4jNIiXAJ+NkBpqH/uCa1UNBy3OPszU1Y5eC+F6uy8PACWmV
MgPOh+9xj0CzvO0iSdvcuEy43FSTuYB2nSzRkuEI7O4nX5X/41PtER+CM+k4
qlNFhc7CTkfsIq1Ge3BbihJXVLcjHX4YwpeCOkzxNWye8vOTagt3rWjypB8a
uCOad/WvHji6pfdwObkehPJrhIfqZgRPwjombd6pUaGCgJGyme0gxTHSwOzl
3KOo0kX3unc679uXnHcR1ePvd3wREAfZzysNc2eFzC4ksHyZTzO+reeOWwjf
Gt0LCdtmDDUe+ZoZ5KEO5C4Du6aCNAchPeFC62SZxtn6Nhy0IWyDMBOdJ6Kx
ZOIxRkqEB8NCklUhpYIk6YFcn54Zx9dyDDLmg/tkuuVqvhdlWB3uBt81HpnD
U1ur09FcCSCC/j5x6shKr/z5vSj5fPg/pLl59NNHUNwFsVl1RXMjxmrp8w4J
cp3wclWxVoYIdTYJGZzTPL55QPxCwTUnu//N71ml67p8p0fdTTtz3SIont2b
MymLH6qzk4Mvx7fD6gDUxB0llfz+MzJeB5j2gxpmOEKEAiREXeHaCLtwAhX0
qRKB4YyE9psNEu9YtVjjWD2jNMPYlVSDeqZ39HTZjjjW0moADgdzBpXjnyM6
S8Zqqi8OCSw0og2gvkrqiSXO3z/qiXWkG+GlkIAJKIaMzjxs1OkRcGCueqxZ
udiswOeXtBeQ0Cn8ju98n67mA3bu+xfGvgrrV322Q1LqtuM2lI0MmmiF/Bdo
oLzSnRq3dKl9MTsmQ2a8UVcJHRMXmzRDZBXzJbr9PAwlatdTght5QTmLeqpv
4iMJdAM+cqAtgG/aBYb1gDkvfCIS7phpfwhCo9MlAbRmPh50Zlm61knj4VzV
A9tb04ZgF2O8DfacWjJ7qOu7uzsfy7hWFIVHiPNsnyl9xkJ1JgYeTmLqteq2
fX1+tWL2gupu6IBh1dmVRacHquK0dQinuX3JuRXizpYSbrVx9OTmKbtj4hRe
q23m2dbv/nB9WlFBv0nuvLjkicW/1ZHJd9hRHRZIDjK/UIoAkAB40SXw8yvC
hg1CmEIRcJWW9t62EpIyCLbukxxeQn5tkD72rzzWMhwfOJurPAPtLi5rCPYv
/ibPTArb/oet6XafSl4yCHy7CzwGeKrr5/U5AdZEZDxGYzjiqd/hoOBNILFZ
EefLWQAQbhg6dl/UIriq2bpLwyYX/btX+OP93n4isWJ/WP9t92XX/pkqskNY
CchGmTq99kJZSAVr867yS2gM5bop3dnaKoe/sBkWNK4bZ+yNoX2IEGZ5ekeq
NgHFDrBX49jtzQWnjO8Kg0QmKBf1ZK8fwNxZ+893Hheg+az8nBXVIY1fIoh7
dgnxOkA4+8PAxQfAXPfhWKQLzhmNgNoTSiTAf/BciS4ePg2kkrk1v1rjbX+o
/VBX93y6+bHcsDXcomOv/X27XOAKVvDj/rY/V02KJtB5a/7hcB4kWs64YvJV
V5K/phMR0CnCse18+1H/onJMHfebo2yxoUR832mpLodyNiuhSQH2YnPAsoSk
7HjNo2MbaEUUo4XR2WGAi2ZToNYnP2MCViqwKR0zkyGVh2o8G+u5pVH+VLfI
3ILIqPDQrw+67S11hm0iq31zIY45w2dwpiAsJ7UBZpZ3xmusCCE6EJF0/nvt
4tDClvoEbsSbw1UvDnFBoANjxAwzrsd3G8igGJlBtHT26R/01dJoh/QYmAHW
+2O0ZcQoTO+3zTZr2YsrVqroZ+zOCcZdcXDIInGeCTYEET2Giune4dZXVqC/
so4K/iyq421Z2keugQkj8HZGAm2pEXmG+K8bpiKrO5FKTbuEO8fc7cKbvJLC
1UlfrEbDE3KsRnY05jn9+NgLkAh7rGUn2IEobzne67P4c4jfyLO6X2SJOI9m
eLFKykaZZiTGIvjpkU7zPNNJrfYJzOx5W9J6m4WLb8WJCc0Lj32YY9FDwNqQ
BoWjn6UXCRqcXaarIHKoCngW4TApq/JQdC1YLcuri2IpMLqTK+EqlvjrBkcK
KdXs5JezhEzAy4H7qc+WbwVrdXHv0MzohNFSZVuW4PSjH89cypHDZuefJLFG
VD26f0XoU7Dp4tVvILPoZTaVxHLHUG9cfB/ZItINZMie2Mh4lb6lHpiwDc2W
pGkXhTEf/gxFzA8exDl/aS9txf0gIIoNbmVpx1Cq+Ge52XmUJtz86NhtvIDb
pl3u31Hsjl3LHg1MbAcfz0Ixb5tg3OadK0tv44yPfDc4zMXVw1XCQJDJl4zw
a+vqXJpghPOn5/5o7vUBi2r2i0vWO/fzFW0UhJ4pI0+D9Wev/9PwLyVpqnJH
SPqRahLE6+SOVkDv4uSnc8BSSj2IUyP5Wk/0oC+wlZbJZ4rm9JVCGLEmx4co
d2UgJCCHtvUXk93WPrZeFGu2z6WLoNC/V3agZc/HXeQ9GXNwETUbNt55wuNY
zoLnw3Q6N+pcvO50ozNHbeISd3RaGMsD+YU8UElk/KsGgjnzdEXSWvI6m0BL
VmY2DlZS1kqmfblzP+OaJbnrgIpal7GoS6hZRv0tM8eq87kh9E+TgX+Tz/tO
SL3RpO/rMdCw9vKYZIou6SLoSBhbf9ObvqowkOgjcXnErANiN7dA5g9nJRVJ
wBzb5Q4DvmMqcuBq4hdcGHOowdPqeApbgApvRdCx1kc0c2miMhqQxe3kAQPI
uUG7G5LiM/C+vKMXzMCHFWJydHR0t5LCJM+ol3Au9idKYjJbVg7UmOzowX45
kI2uScjIryRda51uWCg29VW0vnD6NXUKle7Ts0HOitKVKfBS+V19OLh91bcE
1Yy6i+e/RNW7fXYpfIVBlV4LR1NG2ZP6HV3UnyII7SBRx6qyaIl76W77EW4z
mS7R/30GjGD9B3Af24WE3EiQI05EG4Sotvp7sBhd4q7xb0mLzReWROz2r4w9
RhW/3I6pSQpbtb+roMxOMcc8eK7Wf7SGC34Nkw7kmxJjvC8Q1wJESXbPD7VP
CAbc+fMt1WCUvr86KOvvFSNhL9pcCXm4jtXSPPkavg5Wk4zWTvCtdFS8rUBZ
oftbvGDnTIt92bCc4oz9i1L3q+IYjsrNW6YlzlwxMkl5EB3g0MrGOAzcu8/e
JCBWCUxJr98JLZLgs1KkRkcg/05VVWgYIdlH57H+mrCSm2CSBBA/z/htEz1t
SrFXk7YVWPMHWhB9W9vuFbLxyqD224NApw/94DQasSPP3fWC+UqJzL0LvUwa
jOdfKoJd7P40HCPaKpWxMirWcs93C+7aWvtZ6sbN6j/l4UQX1XmnUJOY/uNn
JQSEuPOO1Gssb8jMg4VJiabk5zVotk6t/Mzu351wtXC/41iilCzoiTjK2Lyv
mpzZ6DbmJan2Rh7XA48iui/IuYCccZQmANNAww7302r1VHTnpCk/vbxVlGlO
hwdxLWuxauAHkzLib74bofhjubFTANO2aW4gSCW+Cfuu38b12Gc5iEJqvZxU
HtHS+PRCrm5gOcu1TKBRJ7nskoNla0Sk6kWz/sG3VUIX0qYP60J+3PansxSR
PuQeVc91G20RhdnSMfpnBIliRZ/TtBlKdaYnPYtp4Mu7TcXl1g0WCZIvw45F
p6LjWZ/7od19uETcfDfet+KZpvArAhyPl7/SFSwEyA1xZCjn3STsE3tTehHV
A94KrMUJ10uzNZBrkSq0iUaYsSY4dRxIoUDRIwPNf5ZLM5SYLRhM2V1867Aa
c/QSRA1SJpXKKRDoo6k6nU2pgHCabanU5gAGsBap+/MqFdmWcy2ye7AOEbb+
ZejJojJwZWbz1CGhH9bCSFzH77X1s7iec1zJAk/SLTqJsICytw5vemWgOnPj
zlOtmh6KEWZXBhAkpXYGw4asOw3tOfDS43gGVbE/OuyuYeyCfX9pMfjjPpae
dOi2R2TT550ob8Y1/L32ktpyxVofT8E+W9Km2Ba3QUh9evyVt1B74nwK8zHF
dWdO+TEFA9I4bxStNFiAzKcoCdxg7Zv2DsaW3+Sl49Ptz12ya2jwhIg7mMpX
idFE+kxkcVLDQ+TRGqO87lA+zOPQ1R/m7UprW87ITLejBdJGUx8GTjzThHMl
ZMN1/xp3rL35Zy2LpQRYSAg9O7QAblLfYBxEu73lZ7aw6WSFzRO0fl1wakI8
U0Hj7jAMvAKevpTNdmBCg6LXYRbO0IBsoI2ULkAYCmBM7SjOEIPCD4AoQhBi
75wn4UvSisKmctUEo/aafrU6/Uky+8syuq7UZRjZbyW6ZNgi03wRe0qi7Ojy
FzUqNwUExruv4QYESj8iw2e7nsCW+MG7H/6GebjcjjMfYuk2A4/qbXTmwImd
OYBQEznaXvDfxIfO7mOPC0X6m26u7AFClceyCvdKZ5uNf7udM7+TS14wr5BU
ohRirozX1fZD4iSHIOArxdB85HYTEjkKWqrNilYPsPP1FR7OS6V+a7cnM69I
v9H7Iqm1s1omtXdq0uL1d42U6k+HUxXupgwb44xHCKm/AMxznL7iuBYZGP5o
u4V+40HGJI7g7I7+C37RcrObr02B712xGYycM1b6o/dqJ2rQSy0ZzXtpu5iL
aDCxqw1ugkPbmpkFYRK/m+da67MUH49n79MWjC0vQjQyOUPJZvyipFh+VuJJ
W0wOaOKB3KXfA37mbn966AKkRGEz2x2L9GgUPrSlVJA1a5OBcxaPf0aR67ff
VHnRzLyQGam3flPOvMglQIZJbng95cfC1iWnFHrUQwA21F13aH8kvfFnPxOf
ecYvGwBlHb4sgKEigDFPgkcvmWdTv/4PEw1morN3Dy0JgZZrHcrrd9x60nPW
INMMVyP5zJK1KGedEpc1OLYDUD1Bea+m4bmyf2F6qKzqFjHIceqacmLKahQv
GZdu1qBoeoRSiV0vP8BrK9x6Ul879fVFfD4IC0zpOkwxdpkBwTOXAWknkaB2
nFQ5fXPb6XVnJT9aPf7Cc1Btp38VVCfqk8EqofPS+SMbYFYV0AFoR1aI5x9c
9YvJLmeWDmCHtzLqyJhX4VRJD9TKHmy3ill2RceG9eZIy3NlsMYuv5B7HBHL
ckkV690Kdp5mhVM37WhYlti3dWduMgjiBPgdrQRkYOIq+wSr8Nphwonpi4d4
KlB3F8Qzmr+QpLmn9Th242n/V2CrGlghUiEHFtv26B07orW7tpzbbrO/07LU
FMaVWunvfKCJ3E7EaviLsmKNd7QPYD5Np042PByfn+oylSsEOe9AkgkoOvkb
MYGnQWccrR3IFV44TfQ/rVUm5MxwBCc5PEASbnYrCUvS0hqNwnWbas47oVsc
hHOAbbEScpkW4UmgkHFEN4QfIG1ACzIBHqRQnvEe0TiFoMWHdPcSWqh7AAXV
4brGeGYcVCIJQfe5cbVvAhdzTlI0A4Ta6APELu4uihVsZPxZkjRcADwSn5+R
Jkn7nriZEQ1kkjDYNkCowshMxR6xPJZgTq16QSF9VPPrQlIGLPet/D6mMATF
mOkbSf3sul3h7BrbvoEhHJXPI1wAAAQ+vp1DgoJQbzA4TdivnJSdpE0awul7
EZPmk+oe9GJhfzaAAV8/yWwZTwz6f8vgxXiQKrXAqX9pjJDOV7amFl+oDnVD
aPv4N5C4UK7WBEmaFevbB/pKy4H2/P11AFS67aycRLygSiv8a8xNvU21A8sD
jc9OeTnKV2QYVSQUbWBY9aDd4XJWMLJe3yS010YFNWjPiTz/wU57AEZiQ0v3
yPfSBW2yGnPCN+LJKOrvc0DXGvnzCF9t091JHnR217rREN2gSGaLimpdvMBC
dCJooMwpMvT+RSUmDTk+3NrjPJ5LUMeiiiixTMN14MyXJlCuDOd6DP674XRg
EVCt46piw9Zqecmnz6XVCwX51FKBVHT8jOnLvCfHXaFrhJqFYx4mCXt+7I95
+zxEIgyY7HBjlu8sKKKEh/woxEtqycLF/B965oN3slonLF2GSZ0/m/9poaCp
rwpwkyee+XycTr1guaJ7+HgBYCk5yrGfylYq8gxF6EQqMfZAuFJjkdZrKylr
DouwJxpl3SGKyOQbTDXUkeGAq25/APFDUnG4ZdUvZfJBCe21VbXhm/2QDkL6
LLgObqB0H138WplbiFJkCVpZ6kdV4IxmskP2LKd9Xn9cKLrg/1ZkbJ6c0cxu
IE4jJ3Co33sx56bVley9m7MhQVGt9kxZGkNNy0hsNN6gW7PzK5TvxbG5lUQq
1V2NpeIvDOTt+2P3Sa0VctdfMHI3GJJg5wH1mEGYBiQu+hgJ+wQuGGA7XS3t
n+v+nZ8ogWaKaR1bZmpNVjS25gYMj6SLowYWLBWXz/bzwhDH5atWC1kcm9v4
zqoGkAJk3oEn3iPdUeK0MfQ05eEmdzCfVwo9CEAQw9pHoSo74EeimC/tBp3i
iOI4xu5ynr6ScnbEdS4pkPISF7V1upYsQkd5KfggtkLirdY+cTjA1BgM9SAr
Yy2wjZqEOPW75LkgaqP0zbjdbSQewNQ0n+5DAEQTg7duUnzEdK/suDu9jILa
sCEC1JOs4Y+K9NEVahJdHc8LqaDgBFH+gFDfJWVSCcWgkSPTSX6cpBmUJPrd
a17ydRLOFXowWOiQn+yUntAVC8dhaKZYMhcJFCq2r5JtR1cXXOSJDDLSS7MT
TGZNpqOuhDBB4MwubLAu3a6kwqj5Qe7c+WDWIdRJSaCvS56V8lj1iCO1hehJ
6XEPStFqDCDkkJqZNs0Gq+a1o46JZ0S6WV7uMxKAMxsLAtk66pvlOXAyOSyy
tO5wrtsYA2C5vPd8Ksk6dc/RSAT92HjsNKo/+JZHzT7RpTsXXUUfX/99crIx
DnwAzxoTUGh9BEEQhY2jSs3+BVVzzxMb7FOYcnmZuv2N1F6Y6pGdVJSDeVhN
LTWNB5jWZ3Gn5nXmhOHLPt3z1r2UtuO97IZyRFaL7i02/owxP5zbUhZMJz6r
EogEpQOOUwy7BtuY3mLD64LB2ib+ulj4sj/SK7yesaIur9b0ih5LKTEBzICs
5mZBTyswBBJF5H8JODCij2gn/31hTrtGhl/MIgObk4St3NUMCYu1aY5Nbc2s
0MEuS38Si4eZqWMHqXvFGDApT3hE7HCbYVHLurThr/Z0CYpf45qJUwnR9WBY
ilYyijt4rAgukxFQGH6smyD3yOPzMIK8ClH9AjEf9thFQOM4/Z2ftUYP+BkD
I9v/J4TA6IEf2cBd8e4XbJCvLXlPuq6I9BRJot7gr9O/9CdCHCUsgkp0aaeH
yYQ8FikbhiVGJsPczliQ558IWX7nol329K9LN4imuVV5N0PljHawVEe60joa
yCR8w5jiARv756VClqykp+3JMeohQsIP53/D6JMw0vBRl4rEUleVvoLlF9qI
H3i9rjuouL8FcFKksb9x6Fj95dehZJvh/t4iw6BTZwkZtSHEbuEMXZ6OHFoF
r5ziOaidEwogS2SdTvOnOe1i7MUIsUbsMsMzpyFR7giU9/n6zm3az3tP8wM9
DQecw5qxAv5BfzSL6xHGnYhvM6N8tu+nBnlLW4EGzAaDK16aDhPB56+Zb+ma
Yemhs5VVLEd7q2M//rXoTCFDebfPtolICLcQ/Gantj/rT3Sh27g+VAS3AhhV
LBUbj4eMGxLM/Jdr1Rz7ZucRjb/m2nt8KYCG8EoRWcifyQvBn8jdC8HVZMgY
eKj/k71fKzBfViYzhqaEan2yayAwefd53aT+fdwIM2kCtdlwRU3i0tSG22Qu
3wYw2vjQIZEUE6H/gRPZ+9DCj3t/Xt+VpEoUnMQwYinw0O7/jJyXfwh20XIn
4zLtcaA1biXK5tZA1u1S7xmR0dZtm26OytvnutPi8UF2gPaCmI/oPH7gZ7fj
OGz9S+x8A4Rc2bQJEj/Y822mS12lX0eZW2/XpSJHbTCuK8ZwLS4Q4+CtZRQH
jkM2XrgzWIefKdwa38Tt/pMVvoLwfMa5blt8FNJpF7uYxYuhjvJUFv6bPlwS
Kb13OGO97hwq70zV+J6jKlgtEre4v8KRD1Go1qSJoT7Z40f2NroasAOhOv7t
V5ypmynnXf+d+4aPAnDK0IrQeOeKzQk8xBza5v0p/h5Jcc2brzE5AoqcGkDG
czR6SZjV8kwo3oXn5RHCL655nR5ApoHQdZZIk8XzOl8izhDfYVkP/y5e8Z4b
1dHJT5hUDapjz63cFtmJBD23iUSrDAMJaPuodPI3MkgORxIOKuk2iMzyQFNd
ke4TXiUz0lqhFcCR4+o53ojTPDte/+UeMxiJcMuhkYTtOzsojmkkdYvXS4aj
VLJKOh6nNu+Qtmrhf3BcHAuyDj8EhLdeL11y9U/FV7B7n5Afnbk9u9tieES7
GhqeZ395PUfwYxKsr+PjY/qRHTKW0xcSC9Armq3HElqtFyXyj1MgNcVc2amA
KSQy3HZOcHVzb8ec+54m11rVXjaLbQe90ETE1sdhGJHIObEKX7HjUVVTG1xN
Dprm/hCq1czBOsy61zA4gz5kWf9kcbliTuMslxm29/4WJcWRHtBTvI1FNfvI
L6VHsSWoGq0zL+pTZ72iHCMNF0stA0QWUC3MXhSCzrVItBo6YWAEayHht0bJ
fMRr63eKziHx0hXb5u2STd+MT+v49/5w2c7/+gY0+JH0sJ1G0PvYN1TP42Pa
qyO/ocYu5lxpCirxRnP7TMZQrsSE3JFLvmkcsZlW0k6tBRJDCKtNvcH+9aci
DVV6rEwyg12Tosh02/raU7WpQHES/l/G//rtT03AQYKhox3r9x2dzqDLApta
pHPsU/3AO1pFN0L7T0njgJH4SAjEfvTJ71kbYXGlAGq/48VVv3MDRs5+001m
ZgcNI7ERpnwIj0HggdgZPBCw7frWKjWN6WaKKN5bw2UJjb2RHo3GLHSseUW+
imXjebxad7lv1Uxh1mcFFKF9D36e2rn0CEQ4h3fl4+ZWyFw1cydkIxT/6yb0
3rHXXiEEgqH1cbnVmTl53iBTHuKkVtzfriq8u2KdfJcKPCHC/1kjn4H/Bqni
7L8akfk5nXJaezU7ThoDkugB2gXY4x8mKmMvI9/Mh8bSBgo8T5Ffnu3PgZNO
ALo77c6mEjxp7YmXqFue8y53E7h5p1SFKYOEOvNsLhfaXgfJFAGvqeZpnHPX
RZORXb0U2zY/KnYIaewsRCVS3YFd/Db1u7rGVlgtPKdTph1iDjqi5Gn9BsLs
OaKL7gH0ZdHXLQOCUuJYOB7xn8QcGrzlFHmAOW2w0lcFIVu1OE3JUX6PGoyU
g6J2PCuJv4uhbCvEAusNGBup3WYvOPqCWY/zea/WLEXQX3XCgi4oUuvuwY7a
7Wq7mL6ip3YK1OOlAK1R9lsuY6dR/snpgwxnL9eyxbzCXl0ra+EEALMmKdU0
CohFS/8OJZfVqmzNlV2H9fq5pALR4WT7bddfohdz25FEZausU+aW6axY/gRL
6SawSJMtDXkgmDOfYOiIKW3d1KYncZfmLg0KAhbQBALOyN2ps3HqYsC++bkU
gsMvS1PFBh0PY0VTZlUdQoTbPv53yi/QLkyRG4NyCEdrtrdmW6Knqf+ZRkra
pfmNgPT2ifzvEqQWl3lJU2T1NmKPR3rGJnAOteHm7C1eW+o4K6XLJZ/ZGjWR
a8wgQ4+DeQal2/c1Ot5lev0SQDLxXH0qrnoYnElEy4tSITt2RgI4ixMf7H10
d6QuIUcpSos6vDgOMRJbputfaCkAzbYwvuO5yraYl2H65iwj5LT+pnZoUWy0
V3k7t98/YJqDISdEXUdamM468j0l/AnqbNY9hwwCz+ihyy4LDYqRaEh4EKxH
mx3FvfTj/xYZeKgmZfBdjl9Il0Gna1LZ0zrhkPg9YJcnNI5jTvdep0xZHhxK
w2JvxuTJ1ODEglT3Bg5Tr/AWHfP+mTNSzn5c8vvC8yR7UX9nFwZy9AYJRsGu
rxPawGkdFIDQVzAZXhXHhou2zv1d3xvN3IYUmlBBu8YBcc8WSkX9C/wE4oQV
xpe+F5vCQIr3i+k6p+n9

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpehXzIbd8EhsSdcosBsMDDmSfaJpaN7SK1ix2euYzgGkXtH+SwtI8DHK/fi40AlQXs2yUYHIwQEb0W9bg3T3WPA+/jxcYTpU2zIJsTT58Pd9UNZJ6HuS2LI92AEMrbtvsmAwSBCG8U7895mw82Lc+0SQiS6Xp3qWR44FmmjxVAuSoJaM3nq03m+z1RDZeaGfKkqoZGO9i5ZRLEKwW5/giMp7BPqwCyPNLdjUvRgNq6M9VzI4tcYmANkHgSdHqpa3/ndhXiAcSr8DzTBtv3QzyzmIcDf24Ijk2bAyoVbH10Dr4gz177UKrpqSB0+EZMBTgSuc9S1pKYwvBJAEJaiOfeo036cN3o7qUs4AKYXXIPMqOT1H3PUazuTwewwb3d0WvBcmywJ6iB06M1+RNH+ffKO2C9kZDjiFItnzpRXwBhZyk5NV1Wo3rulN5F4hFjJokoFI3krotmDiw6V9JVoYReiLjeOJl2PeYmBf9INuhp2pzRoOPAaL2FD1NRE1zzPlwe9iLzAYb/MX4qp3AAIwE+wtOBU2n1EiZmXbLWCSTpHdl00hbKekg5NaEqWu9c5g7WofWKuDW37J7Q9F70T7X3O50mYa7wAM0kGbwK4RFi/Z33rRYXk6SbjIS4Er/2UCtFL9gsEvRV6y5kGlaAZZkD0yBEOIg+ICqnbY/o5e8ejGnTy6QDu+WWsjgsBUiUSVBp4LQ8Qk90EIdoKUWePGj0NQie9t8xleOs+ZOmGquckmtGS264bHpRNdBK0FXSSVmcZAULDeYZSZAjTcu6ukrVza"
`endif