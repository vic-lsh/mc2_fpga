// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IzW2JmGYAIOXh+PR9wCV3nDXQYSfCw6PZXMF/CE6zq3VyvmjjDl3F/JloVgd
kyXsixg3tCe9z0/0x7BUG1A85Hr9nahCAeY09yEO82Z2JOjGCxJdRoGv4goZ
fV7GlGlxZK+t7pip6AkrAU74I0RqtwpZF9vVRqPDSU3iAmHbjyfznHG3v+GG
jD+t/PVTTAsOVhry8o4eit5Vo79jFjFjEdZPfycb5UmmpAju07gp5hi19epI
6RbBzrPs598GLnayDBgmGFSNTyZDh1v3NMtxxctOeakeKMMuv1f/TW9w1qMg
dXQqOKBhr9K3VyWZjOR2UR5bbaP9UZBC45IkcgiN2w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RrFmBLrhzuP8mGOCI9ftmvq9XpB+6wsajHldKTexzXPGaHTeReiICsDCdDrm
FikuaksE8nsXEulwwT2BIq2nnEgqa25bKAtjGsuoYTpZY5KVdkBX0NVTXxSQ
/a/Q7T20Z9DaKiRJNigLBNqaBfTqcROTGPxNFEwPR72d8V+b57xjmaHOgzlY
MqKbGnfU3WXYKJaNlZvtLVULeluDg/HiYlnCQrX5GDiXv+7u6o0595Cebw89
aYck5e7DxiH6f9unVMHjoyVcPfIO1SufQIjQq3nxJk9z5LcLB3V1oufDOnHG
JaUU5ToMYb7gK1TZB3OBMiyZKKD6UxEEykg6GvWBZA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FHGybF4znSQacyi78BJhrssdrbul1YT7IRCryQAx2h6s9JL61olZHm3pky7o
4z2i6HzHyP7Z0/wmLGSOMFCS/3GklQK3NPAGg891K0P5ihydaOUAqtFK66eH
QNIM4CwLLR9/SLX8eXkSIxeNEe/wuu72ep0sZDT0GmySRka1AxhefrLvTyOS
fRIQaXj9BaRo0O7ZeIDDe3DQazeZzmWnqSF2VG/mFiq2SmeePmlSAGjDhuH9
z1O3ym/A3yBYANo0+6qWvGn0dDTjdwKT3UUayYWkIEyU5fA7CArxkD10kwac
0MARgUkILF/9RjdIJRi1PGxFCeQ2SCcIsVF7R6DEUg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qmxOfrTz/5XeRSqzzoH3MJPLkqwxOA3VvLXgxt0Gw8hAqmKWjNAIm9bas/yG
7R3Jq84v5q0DMbrf9+fNdqQTI3fmJ4ldc4bC4795s6/ui8MoqqrJorlg0l6G
eP+7ip1yfq8xunoBB7knXqFBkwACXyJ13rcuLacIYZ4oiKVBEvLBsdD6y4nF
d5G6xMfp/EHZja0DCeaWiNRHM1eQqK7Jm46BkgXN+PYR1K+gcyF+20raGk/5
Dg57uSTJO4cCmtx4s6hSxpIRVfwksaZpTj1WqYmpe+nkRmlRXbUyJ8Gw4M36
1+OWp++vEqimYMnNNWqAs4sjGDWpSYThIG8VKM9fvg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OaiROnFNsppKn9uiU8M7gFEMfJb90Z+K5ciEQafyMV8vCn8MLnjj+aUnxHT3
2BZCw+mDjPTgMy07av6CTkEDR4Jz2VGqjDFVydMu9n/0qfXOibPLxJpmUYzc
4rO8GhPK8Wgf8qlGtDk2RiZ62aR6+lr4qrXGg+CX3aoSb01ATxQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oDVP9m75xgZM0cScwXBvJidR/msavsoVHa98gLQq/Lo+sJEsZWMVbaV5kT1H
VZzyjH8rBCTrMOixeGG219ajHmoN4KpcRxHK5NsdZMxGBe9Pn4Mah7T++je5
N0RVqME9FwKRtb+bDl62GtUXw0a6T7us792rVRlU6KAf6vyPuBVh21bEGX7A
PFrZoUAmvMQrtaVNoCOtczCis0o9o4yB/UsfsXTCh9WZi1c3qjpOQN3nn4Uz
cw4heNKiXkq0O5ywcSb4Y39JjQWDuOPkVD53lu+/K73t1Bges2a2fwPghYVa
G6Nk+bK3XmDaMyhEjZnsFQDxeS66XKEWEcs92clsSnLKgSYjZovwyXsI03u7
3kUQRbdvpDqlVttUTzz6ULwjupRVgoXiXZFvnmJBQI9IENIZSKY4VtwsP+wY
R0RSzqm3p5UQ5db2UHtlqGbtoYoKJudlCiKnMj2DWWz2UfM8Ek0nniYSxmGl
9Bc09zulM2yQlKsN3ibFydklnZ8FAyIf


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OYnLywOwNDKwKAri6ZUGO/2SHf0Rrw06ysUOXYiSTO/Ucgne2al07cfrBPRp
NYONy7TMPBpe9ERn7QD2bFUdkFSukqrUj0SozShT9mnu51IhsDgKgU6NCRvV
+sHx/Hc0Oi0YFrkStI9EIM/nsizLHmY8Lwf6sCqxxuL04f17GxM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fgoc6TT/aKDlQEdArnvmp4ezKbibSeCHvaEh4rlPMdBBCoSWwAUjkZokw5/2
azF4vXbughGOY4rjE8HZFjqyVXpcsjMlf46f0e9GObJkNcVM4ti8C2SdA8hM
uqFb1+yHNdtEJBmEVNkiG8SpOYimrgYFhi5VxORyPUtDOf5U7PA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 85568)
`pragma protect data_block
Y9Q2DtLCD3Evwn7f5utGROZE1u2mgyY7TCphdyNP+lUl/0JDkilRL5LRZTM6
/ivbTybEhEH5WhvSywQDJzWJIXXZkVgDEC6ZwFU0bWmq2Nrjz9KETqjG6Jdz
CmQN1MZu26f7xJ9B/9FZsByCLp0kwNl2WKjD0OFYzDx4E8u+LrgCFv5bRQP0
NElAajRebQYnQMOE19Fl2ML3PPGQPzBG64ytm1SFN63eHdm451WLXqLQPGGp
GOGus29dIsbMBZ5LsNWldXtDhpqVoYiwFyULUekBf4yZ9m77DKLnQoH63viY
KPj1LJXKDPXeMw90H2+LrEnC7pysWH9XneopPC2NfIeGnfYqNHmGtFIs54gb
9CHFJluQSWZTcgIjTHxcBBuYijFGOFjXuXy2NfKPjDPZbIbB3zHFgLmOA+ZC
9wEEd8t2w7YBhBEpOeVnCIxMyWpOxvaAmpfZPkCd+PylY2GxudWSyJIVceLg
F1m2YDkLyicWCp38bcIK2HunCC+5fAlekXzrBwz+rgeCLYauWdYxLGDt5xD0
2NYK/JgdtzJhZyFZmsAn7LZILH2gnmhLJUC9923+C6KddYcXtn4aVGAe8/M3
KWpWfl104IgdI/f0ZPi+xIoYr60AxeTDMrsFEDxKoOkLmKwR4KmeQQxT9ieI
idCIlrnoYZKLENhtRYS8rFdLg7opOF/Hy3KeE4sqTGZMqxDAyrUTNe361RF0
fCJ0mpyk2b2yQcHuU0tlkNnrUtHh/C9cLMXabGBcCiQFGSw0FgOdCx6XCbHz
g9eoZSJW2y7OjgYo/v4m/iXQ/gxqZmI5dxSd+T5zTtAtrOsdTujBrBFYVXUZ
6nYNE6YAqd6buOu7KUnT8/byEOIUhIXLxh2Ck+JXkJSB0ag7F+/6nZXJ7ig4
/HlVomj/cX1gTc7mYdJtkzxks8PHkpfaUK/fxK0IOhWWoCHV3oSVHPWX4wDX
iF5fohXljqMUO291ktsuKyJ8RR2L9+jDFspJxb66O+7dsnraF/4kyWHtZ29U
B62uTKanp4+qJgWluzI6hrtXJXvLXS1v6h8hyTbOGtaa90dmtc0obkxsZARe
yWLuLAzHyoZ460CgFU9VBXaPM1c5CetlzWh5H21DIYIQ5pXmGFX8ODV5Lw4d
BLd0cLahP/Jhjf5J2ucEnrI8qhkzSTeaRm5ymo6F3Ny2BwjazFNtN6fLpXQx
v6aon13bCuPPXrb2BjSXpLoPare9z51Kz1Xh4lEgyI3RKxoo+9CojXQsC3EI
vKnslXfdjqx3ds8WsUbegENdXz693ATvzb26y9Hs/1l7DpKyQiSg+BD0jeNy
58pLXOoWpZgW6Egy4JCX6np8C/KO94i7ydO2sGFcB5QkfxLCaL6UPDzhi5zV
naihuPWw4dXFGonkxj09QFrQ2XQfNrWcn53L+1zcFoTa0BuSlhaQROANOzU/
tidnX1RxhNXAExpdl9fuV77snYwTEKpLXmjsbSiRqruDsdwb58gM0rlKI1/S
84b202AtQJ7kr5mvl1b8fNTgkHAlWY15EZ3sSFzElMbjkQZul+YYj6ZbGbXa
V1am+Q+emoiX6A9dQ5I22uymHGsgqfs8Hzf7AGdj6j79lEsIP9piy9hAKi0z
q3AOP9V/8ErHlhZompZIdR9wh54mnxdeAcnpQYq41pEqI3Tv3EtU9d4cR52N
l70GTo1wkUKW1t9G1Dbqs+tt6ft1ZIGTxTQhBBbXqkGe3VkUqG2FrFTPVApy
oagaAVbuNmqqCA0dubJs3O23Hdjl9Ggat2abcLDgAvrake3R1HD4E937012J
lAz6FNzKUU+UmfQ3VGtMds5n7FZGpSscv8Vp57G49KMTDcxZZmsg5mvIo8hz
gUdiV+uaJZVcItBZ7lkMdGFkkbjP5zM4pgZeTaURvy8HcWWsc2Nz7zkMaiss
8Gxo5Elty36dRkMCOBqRaa4Y4dRYaaPK1KenAWDlg9fSLo0CmebwN9BOEUi2
KwIPFiKmszjv/kRauSnz0wvJdoykNx5qS7jy3yX9nnqB7zR1mBLZ2HtoP78y
uJwLECOta9fXbJVBJxQxzIYjmjmWSf0iUJ8x2qIKFt2ooQqeTVjyPwl+/BW1
nzpjlRISF3iY+XAhsXxM5le8lESB6EjiFxAebkaGrZXtZyfc5MvuI7fnzG9z
WtKUj0WXH9oGoDly7/PUSo4DwsyI5Rs6KtHTEuQMkl3upe57WsHZyeRZ/57G
1D5arLpYZlgCOz3Jf5mEvYULDeSLL23Yr57CvPLHhRNNbfpYv4LKNSa0kyLm
SogpJKqSurTZbfQKW/Zh+SwKk+PxR8EWO9eTxsh0327oDXvsnmbTUR9oeRxr
pZqwjOp1pPvBcJqswT5+C2vbmS3hoyXsb/XHVAlI8SbemxRlivH5KAl0UkR1
X3p1S+MhQC4kFCOf2AxQced701Pj5ksQ5VCvDpW6Kiz5ehUga9o9435nXGE0
DUBcludIEwS5tCN8hUiOfF+aX5oupuUwRUS5EgZO4S43pUfg8XUcmyTUNDxp
LAKxXDM9IMiJ9VWZLwomo2judeKdBO8yWPcmcregifkkKBQT02VNblc/wqRX
SYxt+ZBVGCuuHe1POFsQATvY+tLiUBkqH4X7Qt2Ew37FmmaD9r55mpAa+3ex
Dmop8ioH4Zn35Z86hZRXViPwZX4S5hlp5EN8zbu/PCOVBNMm8WKKPWyBDsTz
vOwJCWPI/TsqYxTlzTki3ez1TmzYQeJK/YMYaodzjpmrQXk/K5VV5/LHT58Y
uiqiD0J3lW83pmq+pEpKuWggwEVmDpnf2wH3laMPJlUc5eWzFBdKZXEn0WUF
5BbrNBxmX5+qE1BxEi2C86b99I0YgNXtu8AK5jaqazRptxz2CHgA90v/8sEs
u+hxobnoerBWG8j0RsJ/fhbYae7hpfoxpJUyT7KzcGmoQBfru2FXD/+TR3LC
Fh/h6XkCyZZdM9WjC60vsI948mTeRb4ylHAChZMVnPO5xlIL5VqDCCuWJnxm
7mlZMlDoP2uN1yurLMEYWMI+JGpyu5XRL8agAl8iEy6SihPLrhRPUr3+KtpK
Vy05xU2X6S38OXbMOckWA0q8VUwXU72LCf2RQdTOc/KXpj0WYwwdhVn+z+Os
59O7+v/qM3gAL3hin0/Fe0kQCxwD912UylHW4Xmcbwc6Ig1M2Zbp645tmcjS
0fAp5UznZGVKeRCuwbG9buIyiPrXCYIzRO7TRyFyjPhW5se9ChxajXGdK/UX
JJ6z8dupABLC74fVklNOEXvHJ88FEFRtgYJk6sBjixQNoz0n+z675b1Ly/Se
5/swYD/MNn+9dbJexdP5xHjAJckHKFmMiKw/zwkI1bfHgiLG4ESplR3PBAdZ
ZWksaCkU2DiSJWWgwIKnvjGbwgwAOBO93t1f2QT07Yg6f1CUBs4S2T4BrVcV
wf3iI4tBI3as6r37MDaPGVeG5DRQYUtXnlHijZLpJMa/XLIexX6KbYpElrbH
YtuoRVikpvVC0FJ2vZlLZSZiLP+qcze+lNTGhHCGIvJRjYetAyxlmY5aoJe+
Bi575GdIldn4f3/hKBHueL3DGmMz+0P/3r//19S2l5zwBdxpm9jpkNdd5uXG
by7Sc2zy6q1431z4elY2Ps/82iZHTOtJ5Psd6Pm4chf08KGpPX1/1eCcjJew
qHhcYJNaQw3VLoBRD7r8yoqz2T8VWdpoiSZY/J49GWFD0hXTawzb5TPZt9cX
8hxXVtApw/7ISoF16+QA6sj7bK/8CW7awLH77EU2DO0y0pU9TwYzuxSQGug6
Tff0SrZDdqBjZHVqjQ3NxqqhBs0ewP61PXSjcU5DK4vvkzv1/hyVauMyoFU+
4bO4SgO4zDbCkmt58+QRAE5RuRrCxMf5bMNrlWjzyGsytRsBa/zPBOEcGyei
3Rlr7l5EkE2RpUAqxQulaZbM6pZrlM7kq2WMZPGlSesuvXfmCfAx6dDWh0dF
rHQEIwNWFF97/1nEt69uKL3vs+37IdEAm/rJROTseLJzLKdVACpbQ7oUkq/Z
7TGkqREr9FLri4pxXrRsbI7qB7Dq6sDm9VSsQD5Wc2HxsaePXcjlwIPqoEDw
sGKz8ItNSi0m+Zf7rKilkCMM1hbAWhzdX5u7JDqbkXCTOfkx1yrNR4ik8wFN
X/0AzTRvAPq0BiMRdTkRRRfbuPoKjFW0oy5E/BLiX+k/Lmx6VercACRKv9Mi
OotDZ7juT0zPvtms3z0ARNw1CndnC/DovrD+tgjR/iMqXq4YV33I/sgqxkQW
2xmAc6wqN9txZiXkkoLFOWhiU3SjtX3f2DOK6OGkyKHgpgwf5pMuStALadl4
SgVGvsrZ5cKQE+WsvzxvL7J22NThsQhm1lcqLBuyEitVyqblxpib0mHB51WS
pmlXAJfs3GLkR1jokUQAKYl6zvTtEmsxZOYLfH22L7q36I/Er1pRwQAroTiz
SEpQ45pVioIF5+dIYHuzLsVn3aMY1mEbwwTwGfJBPeXVtc3BMf83Y0ZtmsL9
041paZgK98VeQxvJ+pJwQt7OTci+aHdH5bAuj4pGaA2ggq3FJBgWzx47FSQV
NhmJHXq8yEabbNHHxQFlwNUpXJ9rKFXBxCjj6QxYY+qvxI9IY9ZXY3j5yVuL
CBxjUAXb6Cnp1QuNErqZvza9ovOc2dtsFpgVy8jG4n8zD9gdrLTQoIZl1Zv6
1Nkf9z9xM1Nbi+uGt+Uz2/O3UFJkKLULafTyr2eg0kG1T8kXER8iSNQyP7K4
WCA/KpG4wFmfk8adNXwbYAyoG6jEq2B4Wpdu7/B8ZrYjgU62GNNHunMRt7kv
JIDtLpEe8HHLKsmTs5K6Zj0yMQ1M/xktzetIVby5oFzjYVWQbDin72ylBHug
HEgWZLseue3lJ+g/XpHT1pnv1CJafgSsKwV8VXcpDI249jgykn1hpOSP3VTz
k9aNf+qzBDUdBMvURryOViHnP50/W99By4GuRPFVaXjUeUrMku0Mo1qp4Ll/
Najw63nPSLfXsk34H4TB/IH6WAxDUSUF6ntWNmWQ1o/nzEgQLdrREwSEe35Y
Eymssj/PhAwswFBicqCOSRjmDz41uVjljLNp88ESvIjPyh6mHLNV+vVhR3SX
YXwJBS4XFb4506WkUpnBI0PkWEXyiktzFnTepkzTnbwX8da/e3u/dnQP6xqF
yYJn9DDB62ydIxuSI/xQS+Hb/SbYwGTg2YJFPmCYjB278dfspll6ZQ7fdtIX
xkCvsCr0BuMnwvtGrHy9L168rNf6GX97O4mWrTK6NNMZ7/v5dJrMb2zIWKFC
ZKmcTBgBw9GiJCKOoQwV1xOZQy9hlSgOF0mI2uYtZlr4K3zxlMG8eotkibWN
2SLaNh3yk4OjgNnuacmeirO3BRVQucVjfbq1hmmAqZtbgicmPR/mxvUx4yu7
0Sq+nxVO2bJsuDdY6flXdWPrsc4rHfw+ZVOiDiG/svuWTv4rpOKJpV09jGa2
8+4faC/B69v/GptCVYC96kzu1L+ZUL5roWRioCSbrFRDpJeSRng/4wOuP9zb
lDbT6cBT89Y3mGNw8SMkYKiVON5ybrx7JCFcigbrlgyemIRoU8uJBuX1oCN5
UxQcKa68JmGblp6abHBZNp0iHjGVjJVeEhFqxjs/1uyqYjWz48zSCgB96tV4
dN+A/Xvu9ZumPRzCM9X1zusKOAlyyY3CSCoAKvvYUwEVouAPm+CyffQDvaEf
tJaQBJOZybLkRid/OBpTtm36Tl20xwGn78GMFVQuw/qzIpTBIkvtejIC6lIj
h+QsEpkFolQp682iOITcEq1ER1t0Ixcgf3HwddL1jn74i6JC/LpE6zeL2hkt
Hze2VJ1ganG+5PtItjb8QtHD+UrdLrQ0cSlVmsMWceOeUI0a8iZVKjguGfbx
TaBVEYcQUp6LP3pGYHGASnz8eM9RXGBxi/XX5CMaQLFNRpHGzm45eHJJXcdq
rAtWixw3kx54vvRg+aHiQ+zQmEMLLPsUXybkKnmSBOgOObuhLP43Rwir0WRi
wRfPaxD+eQAWL8LcmbuG9OIyJ9+9R9MHoOtaUvaL0qtcOOSwK5G2ma6OrZqi
vMRnIeYbjSLDrTuOMYqgXgCFGLOOkkVZVRZAdjLBGPjMXLd7RPdeM+6CznCb
2k4e3AZPKU7k0w5xmj5AfiXXnGQX6ftAUpxiH/27RVZSW4Q6lD2kt1fbC+PL
+bfJzuRE5+ugYZVAbzQoyJo2covbDGM8fFGjOYmE4ICec738Yr2N31JHBivC
cRi14/V10AW+cscfEubFjrwzezxv/6GKXbpZrAusywE3arvz/7TZXAHbpUpv
9lC090C0+Iw6BESCwPm8+myL/s3EKk4lp9iaiJQK5U4Pt7fSkehPDmOmv3ap
FNKIa3bvL70ym88YCHsevKKny90AwMkaF2FN/Bz+8YkCnGR7p6pn5tmahpAC
UF+ZN0tYkufJRdlsXSqmngi9KraTnju+nNVpeV+MyBDO7CH58e6rAfvGDuhf
HeZ95XJYEcHx4nSk2QCc+KiFxgmeqwVYojG+eRibL2sABJ+qqxHj1prQE5sv
1purR+QF8gOuStgRsDKGb95FyLyDOcIgbgPyO7RMLELe0AFCAkdj37V63nyj
Kg5iz9HZUhWhcpQU+tYoGnoXLXI9ctxfdgn8g1oG3ezUTd4+aEkHATa4Gt7t
AccLksMjI3ru3NxCo8rzcP6jrYZqQI7tArcEzL5ODArtyjYNwGFqoJoybFvs
PTIxuLZS3Pz3XBvZD/iQhkqGSzKtSpTGWlDjvO3cWDGXQoD99AH8UyJALojf
8KuuBSgQe57rpYu9nKDotcwahVEW1edrXxuqiISbSJiuFwzUKsA6HGO4zsiU
B6Q3iO4T+IIN1RtrKkgQ6n9N+07OOI/pM6Akqj00Se1FpWIiqLU/IMEVNgn6
exHH2wivua5ztF/xCKVwkG+Tl0t3Kqeob9a3DlCJE9uJk5xeG9rzaiSLChCN
kvxWxb0R3jjXcvibfg2sLxmV9zioHrKlrHmw/Mx/9QJeGUlNHftfo9bnqHKm
03F0SXn3F0Hrsn30rsj1tKPkQSFZX5Qlx/bOlH4oTRX5YZ447BqVFzR96Nm6
9zdoGs2mey8a86QieXPK4+rfGx0eFpJsWxGUNGZj7JRCm5FFrqKsvushSEsO
nCPyIjnhCdEUuosBV8mbqZfv9d0eIeKNrjXPs2Qpy0W31SEmhzrYUkUKb5N8
LIz7BZM9teswQcOKRgRx9YRGPSvSvUCRpSKpiP9v8Qg/G+3HOBXDK3bvy9/s
HcqNqXZI5gQoWSWcgz+4yO264UviZfGU45z+8pr1336NFr0fChiPEDhmrhID
MceV821QUHMSb/4eHqWDyzOpa0mx8B7uPTBPy7Vlx/tFdixY+cjVBTAPkeey
dVTkHDzvR7e9j/D3Vgp9GDBSOMCOy4dHH6iwIA3k1aZE/C0SzvQAaxCyyz39
xZwaSNWnbB2SVe1ePDlBFxIaIgkYBwmzgNHgYlb6YF30B+uOQ23VqecOcol4
/vddWzIW1kcBnWkVpLcxNUJXdvA8w3S7N8tM/kyykTyXZYCXEqJVULIwozga
XmvPSaMnWeaXP9DwZvb4q+nxcCqjX8LtrSv5plVXcUF5fbnIwJ45WtdD1PD7
tAERutnFT6N7y9EXgkrZRLVvIoro3U04/APykyQ5rvD4tPVyNumcAXAdvvta
mE4SAiVww+5kwsf3kPk06T6W8m3k5cN72WA2uMXYV5c2DeNuKMlBao5XJkYq
p+rQFE+vbM+uxySUTh3gkpqhvIIHXNCJLgcBa0ryvIa+9Azu94g5oZU1dROh
qHVXCCEoZklHlGLAidv9OUpXsMWczTXrClgSBqSKP0T03yG4MifR9xLIYDH0
lkSp7ZnJ7w9asEFj3E/cEQzBnEVxwN20ih12VzyStXB/11clucMitDKoDNDV
a2B5lLbdxADThHO2B1cCCDRH63XwKXB6okTaU35tAXvluzli5adTcCN1/YSw
kMs8RdoQyjf0RgNPDNmZEN8JtUZA0Vu/lKPHuASjhNgj4TSll9TVJ73HmHfe
HHROumzpkfYfZnpOYPKcgJdDcM6S9m0iAXCg08i6h+LCxuH1e39oyIhp9mr6
7CBj3xqg3MFNe0NFMHOVpHytu+iuP9GwfsTfUHBX70OOa6J5IOkCQb9cvghj
mmm0XjR8/yPd8mvANEa5OX/2mC9aONYCdICKzOwcp4QvwJsQLAFO23KTv12H
4yZhi4lC60gLf/GpIGY+iiSS3NmQK5V3x9nTr7TQ0Ti/YAji5maHbN7YTy3j
MUT2DHJQ5LX3YQkzRmUFgYr7TDpcZmJhmtucD3K9TH9K8C8raVW19zJj3kMK
kwkeIKWtdgFEnNUsgivLTP8YKECZ2iJ5LiYcp0KlopIG6Zi9OZX1bKsyM/wK
oOpr4bgY9PsuqrDY+OJHAuS/zFGv1gYUMD7tib9Lj+YEVITjYZxkzEAuaoch
YDI9Hpkp6mPYvUPjNCkPVrAWYX1CQh8WTnh8FG4+NnfALN12IflsarFrJkAW
cDZnEWQ7W0sOJCTq5MCJwFOyvsFLBYqGNxvCVcXtsbQJlXwZ2AbRs2egKq8h
Z+xuMHq2HEgWBRj5rsQQJoDm/ej++peuKZoBhk3bthICTwPDhdvUL5vXTOs9
65+/kA0rqugOy8X6JD3+nRirBEZQ1+cwuQUkJ73DxO3RPDV/fhJQehopIPUX
/LPYu2rCnABoeDfLziSMG7NV7kpEaPQ+9dK+J7jornRI5gxLKUR8SNzLMKRW
d9k4G/RTq1Lyo7Ie8vFGkUKSZCHZIhWnhix3t//9iIoyxqIl8BRGbh2Prvos
kgc0orYq9G6M9LNfnW+S82sY4thTNo3HhdKIkFjqY7CQpxlFSoB80pFs9Wyb
mKxWcIBZQg2sfNwqb0o8plQLVB5hHmeTY+bbwDrdzi2sa2O9q8Wzk6abEaZy
tJ2f/DrF6ZjI7LilkIY7kSVodSEkspoOAWPXDaxkwu6BGDJNGruishaLCmao
dWz4dwnF3KxsQCbeSRHAjJGZgTvEFFCjE08ofA3k4cDNeK93x5TiHKHWmOTn
UplS9a2mcidjqxIweHoYE0aAL81BXMvQndiDlAUqdhR4KwVsRh1nr2uyPyZs
V58Lc21vwrjuLrXnrGaiRCSF2iBco1enL/blgcX+ioOAWMdbNOLnhVoqUUwM
xw58C4P9qXeEShz46002+x3/EYA28KVDDQS+dZlptSSjzeaFzq0hEeYqAkZf
ROV/QguSWgofxMAfRzhSVe0wDpZsJnc9C9FWoYz7IoOnJGAx04V5HCAo2Q1d
oCkFX3UqdQ9i7llp6IoTa29OI2l2MJnshHvOTJb7LdqkPt2v1QKRpWKa6bxT
DDF/9MlGOU4elikWZq/+XBa5azB2dF1vBzPWm8ANpaaLfD4Mbu5w9nUYG/5Z
kIa4YWWxbsIkNS0REjiBlky35jHbWeiCYn5ELCRVkQlwNrPzAEjn1WpbikiT
8tyltaeeck7fhSlCzC1Bsw5aHWCM63nCG2FE/UduX2VoeVf0cSjFCZmkkWjv
dFzsh+6l9aR517WKnued4tPUHalsyO9mx1MLkzO3ujfeG1R1VxX9gnLXvpTW
mwn0sU/FTOK8gACuuUt2O1/wQ81lSyfHbzMOv/zFYRDpCADc4TfUn0DVdTcr
O0To6cHB0GDOJz+H+EKl97y3cOa+YilKi8gs6CHsuMcFSH1tEfzMjEiUZEgA
6VsOVlldxJpMmu20RipMYX0Re9X60YiGs6zKsaLzs9hZZWD2AlxFIzhA8lJ9
vL9MlbOPCqa5yGmL3RsNkeT04OzwLjSeZB0mqjkHSv2hqCci7cf0ueb6w0e4
Mgfa01yt7PTGUjBGv0JoIOxRNi7kg4ycsPuMqrAwTgAXQ1HAXE78d6fKyy/h
ty7Zeg0QEfHMunV1EoS8iVYjiGf/L5fUwT6rTuzdQjq0BBqGQT6gj0NdMk1G
7XCS+NeMO7GABQK+Z9l2wevThxCS3fn/+EsdUEjytaKIKixqb7v7f4LkcamL
HtfucvUNMGYXk6xA2ZDW1NoRyH4T4wgcwx2vPICFurSIZ2kBxphXGvE/koMB
bZblPrqG7rLB4qrhJYBJoLp8hVwATSQvw+v53Y31yI6lWrrl8mi5Yit1deX6
HmtLNQPzoEMOqq1jiO8CmgaCjaiCo3xfkhhQbp4uoMKCl3eidTEfS2MiCJoL
iDw3L6zQzVAnKPK4/26KrDQgsofcGPqlo/hXg49Qlac/IwizWyNmrxV+Y2kp
oIITytxJDln367el5uToCc9BIdSeudIXVsRvLzgGX0Fp18VHB+w68PWAgbbI
ISl2rzAMrZORwAz5B4FNBzUv5Ez74q2GLHy5JXrGSptHQFnHJqT39Z+UIINX
1xVennm9nxxPAxuJcN1GCG43us+VFCVxMDM7X9XPJFBWhYA92nSyBRQmUaJG
AojgEzlGbesas7t7d1+ooeqZKyi5XsRlGI873eeaZ5pUkh3nC+o9/nTFuPy+
rTYK3sdgEOmg90Z98s0XEsyhnEXP9hVlopScc6gHMAwBBNnLYo0YcxlU+Kxt
K+g6VZ8eHkNa3GRVA2/29sMuS5PQEB4cvDMmS3bU3BwjhwV93GYjA40z+bNp
b8vWW2c1EV7ZmZEpEErR3jQgOAsWGCuZuQas6DTxmBcjPhsYo6NPlv+tlog3
oIR2ABcPtK4EeFIkJm5UZ1G4DmSxm3U+EdEIDBRdl5letuRsJRRmkAY+De8e
kvDiMi1BzkL0RdyqODgSYyggSJOzhGMqCntiYh6otJ3W+QgtvJP2IFFqseeW
OA1L/YidRxyZaSa/AdEY+6ijydOmWpfXCX55W3TBPc2agVUWmvQft3czK3HH
YOii6PNGnbLT0+ZRjYCdBnvNDJOdLYv+7NvV2OkCI94zzZzPivpEuZSViUZV
TvFAWWiysHZppRv40zXIOwLXsR/If0Uxy8dInYarIbNkBzSAJEJ0jvnX8lGn
qTan/MbV6FZcZKmBU2y5xTyggPqnr3+miPfc+p7ltZyk37txpTqHZpgNz+nX
fZbfG3Tk9hsUfgE4Bi7NUQg7PwQkOAaS1+jDnwaUUFmBA/OeVqWY4AwnCqsS
nrWiGeVGXHNZ4U3w933frch/9YSgxTzAmOZwe6bme3Rt8ezIffvqTkeDZH5F
CDVUi1jMN0G2dp7kD3dx641+3KLPwU+S48Ht/Foo2YYycjQBHzKxJGhGQ9gX
H94ro/zc9Bkv1kKLoKeIlkcdacF+D5cOEUZlfexbRnB7XXUELo9gkhwZk/oG
Fw4YV2qG6kx3W3F7YCbeDnsZAcvcbnkMMOevj5gO+rcsP8UY5nzRhwva8wUZ
hFwGdN0kU8a6ZnpXcso9xPuEG49qi6Hgw/R1A9Wf38IJ6VRX/pqrYemp30T7
sMggUOODezCwB6I9CKTZQyXvGi7Z4+oQLrYdhWh6lgkgXgwPCTSssWol0cTS
B80f4B/Yg3a2rk8Mur+sfi8l6QQ3dw63UsWrcabQPPhpi+cIbHVRNakNLIP/
0CihgTpKnezOy3Xx61cE1+2qTyycJg7XU8rf7uBDOnDy4WzMWyz3pdXj5nLR
J+PKBnENM7aq4OZx6x8HGqFp7ZNZwkHVeC61FUanYDl3DLpDPSUwszXNTaqw
SeZNzA0a7aYNWOjpcYVQwp2f1c5uZtHwApIxPVk8PTkAYvpzRwRhDxwH8RDk
0Im8FCPf7NMjxbBccDK3QYc/wmugH+kX4PDE511A2/0o853TLNu9R1b/VVhD
6iFATJNLoKRjqa+9z/AVAEk6EkOziI3OqmKQFrByKYVQNYu5wnzCaqsZdT3K
DzPVne6sPp0eOkPT+tl8MAR//kQva8bybN9IWf1+flQfOqHPBqSm/R8Mv7YF
FYP1xs8PZTer8P0MPI0WOOjt6kFOjS6qXEpC5SHSZjqgVAcLOMTqlVUFSC3k
WbEUyl7pbdFiL2gDGwAKM4wYCuaAwivW78OtjocROROCXUw1ylAEVQBAS+qq
wQEBDSFYR3LqG+G7yNmCBbqv+vVXUpeZTlVAXiNrNR2v29GVWoC2nL1NEPQy
tgerQ4q6dQon9J0WKvLPjYPOu2sIfF6ggsMsg8AEnyKEBWYIV0g7xO3e71DR
AbI+83MijC4RYfp1nE1yrXIoRpJe2L9LUeD0Qd08CK/0WJkHAdAHbxkkOUCC
FhSubX934rLfT4E0m2/L3724c1+ZzZwYjRbPhzmHYW74z0z/4tEtuepTQw5T
N6n4FiBRexjeuNVgn+aJ0G5nhbtLXcTU5R5eI+/StQEwXRWG86gMdMd29ET8
8VDLWEBU08DxedckCjV2sq19RQ2uqGkzjrSjgGDFCe/F13Ix2ghxffhr1bMA
bhEpBdNWbJcHK/MpVlZeZFTOA9XzoJaBIZWrmmbAaQxrf/0ww+1Rvgf7V2+G
DNxr/9Eu+Tm0x3PDf6VVDfdsfPf1L0ijodDd1kVnJA+uExm2+o5QQx/+a60b
ZPIIXFJLNb9CAwym9UMwqw6v0dFah1HHazifc34ReQEe1MAv3knL1uBvs2Pf
9K/eP3+aEkSmnu3/H1TPlSQlok7C6pAhOfHtsilOgxT1jptBsFuIOKVd/8Oc
KIrpq6dVemMFE3goxRzfH+ulJG/n6Lsltxk7MTA21Yq/lsvrHidqE6WZG70K
hRXMbOIWht4i4Lqv8/TQqm5GnR+dYqHTQ9sa/q8bABsu/YtqKrCWlIN2rnUb
qHvd3gdyfdzSXrsZTykLAnBTW67Q3VUWPSdou+U3wri8gDTJr/yRU5Elk5md
jKEGUDnOgP2f5gx429f/CFRvPmYHLAo4rMI/px4ccLan+rGBFEm4HZgPm/W3
86xZsoDdj8QONmYqc54yFCmo/v5FGG9NcRaC9xzGRRJJGsHL0dSsM5of2Ycq
qL/YsQtLbGYbyaYmW6qzidtPDUpgfQy6gIlvkZn4urW4iSneGYRPGWOc0dEQ
bTKqr0ZHBEl8zMzuXlnCh2F2sI9+ly1KuvIwFwgHH15pxJYmw4Sb1STpAPnT
Dg7Lh+lx0fh75Ue698g6Sj8Gq28WfqWRuAeQ12UtYySSg0ThPt40oP+fODjm
6u9hjARB57rEseYBZWnuAEsp4sJC0CivU9LKlF42qePpp6wZt8cxg1TqiA3B
VT4F0dhljvOBulthtCNzAw4ByLCDCh4Lk/Cxhenq5gkbiyiVyq2c+N7cvYm2
RuMv2fyGMZ/sALbh58SKc6GW53NHi1s6tamugBI2dUTteoFN2FwVFQ+Ozh/N
bDkCMeMyRmZjr91lJejvv7yqtxob5/7GPeKuULIHgjVI7cbhLuPtmHTad6AZ
H41UGkOF7O1WVddDNFsIx7IpTlqkIzabwv7hcu6tY+OHG2pWY12kpJCBl62b
UQkoIEsHJo9edvkfCzUHTW3Xmblk0JnbrcKExpe88HRGgZDymENKc+aj26Lf
/0jelN84uBITQWSQRsFEhNKxkA8HLuXiJcT1oX6m8fCTxu6vUgG63At98K70
IbZ8BdicwsmUTFoZ/usxt7yBMRw+24bzcemkS6ZEnBEiXfSh2ld0CISUeWck
m7wTcEwBtkIXySpwJUh129Hqcqz8pRf2f2TyRMdCGG9Zx84xRt3DUhNRYL4G
ZHSpXW/EVX2878MwAz/g6tD6XikuRi7ACMvvt7IIifeZCq9MtilSF6FZc+Yg
SCAfHujARG0sUcpS1Gfbrwgz0uohJnRFw2GNFB1vyuyANrpvW8eR6yf3IkFr
jWjq1MlfD5/WfJdbgTsfv+eVG2yG4kscFskMP1epDVXu9TY+z1EZyRjImyS/
WFY/9Nh8bgirNwJU0ZzuDJ4dDQiagIfDvjLmFNp9FN+wuOQauLL7P6tKSX93
6CbHX3cWzq9hRqR8QLh6TV72/S8DPbx0gcU5NhhF+GKPcoKF/Ra2QnBLjj5m
SJ9i28XlhhZCHX/1WdOjiR5Ub4boT2JaLTlb6xF+FPF6UA5+eJDUlkaUB3hS
M2uZkIMp5eJLUD5aZwtpUnLrprR+TPcaTdD/628/EypDLlEVmWoMTvoD5y8C
oH2k3NPsDjroAVQGT6M3hCXUQvJ7qeqnRik/qG0ernw+2uZikg/nYg/5NFt+
4OUILdHeQNM+HRPEZbz/hg1Rpoj6zajD73d6PM3GCd7tiHZOhsDuuQislPjM
aoHnKrFRnLLaMekMGqRf7/QA+wI1FXmEwS9rEo7HeVDLEBfb74+wnXDXjujO
MySTnGmV3IgE3o4KYg2llweeKNiDn1X8H9Wk3FCNpSoxbiwcaPPWwdSlQYbX
KdkLMjXkkzPQa6rIugiCIqYzAzzM/avrUzLZN6JUsnIGfxH8ieYff6me4KCM
FvvquBLZlgAEcU6xnuerVZbDC0wCCRew40MLFypQMnqhg3xvCB92S8EeiWZ/
4B0YSMOqmxyVBruNZS1R+zAuqHapBwaFRoMgW4t38uvTqjXkBbsUYmt2pWK+
yZnLh3ZJSPP2ZMfqRpxYlO04jnUegaUnnkuxPm7BkoOMWJygoKTAbfT4a74s
3RRf3vRZwlfvyux7lunrl8aVRYzGu9QMySjSG1kIkkl88Zofm2HjsNAVy5y4
HffJj1F5iW9pDxMFZXyt4PfGvgJA0pY9p58Gt0YY2kRXSv19KY9Xr4+cRWst
NvqIPIiEQGp638J+dhLnsDUMxlulx1YC8Ico6C1Yj/LlNbczNd4gHljpjoGK
SSI3GxfFdFm9Kd7ZufNykWcNJ9YQWbvOrxKJdcwD8hJgDBG+HsUzeadjdUBP
LZgpF1LqP8TGHUcNtVGgkd8tEdN83iwnk1xbZQBkHA7e8cn6EXfAYeGSc04q
RzQ3MkEOTf0ZqOd9py2BYYXih8/cn/BgAjNP/uUtMZC98ANacUnu8vAcFpDS
3YeU2XC52Wmd7bktRsQUKK7KhXrkxq0WLhKBFyxybQa4DsoFGyAHVCmVByuU
A2Nh/twSHcKCHKZdTPtFS7amr3pwU4s/3X6eo9ISXkQ//Te43ADUn09+ieDL
idFM51Xxb36VdOzZvhyH768K4us+g6krmE//bIrmncsy1EHjook/bjAUYKjn
YngcUcn+aTOHDoRftmkFuaiUdoFBWbqPZ2AII4qX8qbBP2YBN1LjLhdsU6lH
wj2J0hsrHxEzuaJ51HznIawigkrPaQYTMaq/dj3HgmC1UuciEsSZc7AoKsfS
36whNG4q8xlHiS89Om/wz9T0Fw8SECUlmaytcaf/CJnDuvzCnq1+Tm33+XY0
uFUk25XwD+MWRB/WADGUMWv8/fq0oUyI4xRDMBrCqVfCmJhoOcj9p9QEGQI2
ZcmCZaKUnktNMXrO9G7t9rw/m1sfed0Bsy3DIseDWKbUK7nWHJOJjrPbUawM
XHzvUQLW60WGVZcatp1fdu3jOG+aZ11ayNSQSZrd8JpKl4+M3UDyFFlNZU9w
KCZKde9Q0ExZ07p6I+m8Yx81GnNH/KReZ3PFwviWj0TNBVtu0aTlQc6nl2Pm
wLxAU1Hr25KpuxLCk6oakXXw/yOPt8tJEvzjovHXCNspwGWMhzePRkuS2YZ+
UFJJzUiIjVeOW5/ifLDjV/Pm7v+4xx08BweeOzshIWuFW0GdTbcAxh0Luxqg
i2gbXNVX7asPq5V1Mu1vGABpsJy1mKrIR4k5goFdA9C8YEJrK/q7dbhZmdWK
slD1QCAClzM7TCk+dH9fpVrT7+wjvND2w80Dv9UOA8JD4Uxy8yH2AvaIAF2I
k7Rj6ZgkDHsMyOirvW+2oPvtbzYNc3AW8PzNZyJOb7XLAjVKGxIAG/4AMHb1
ffTub0+yH8lJEX8A9DcwMtk+bf2I/nJjWeghB3uHecSHyLHQ+W1Mbp+AkbWE
zff40fjLAabV+JiNDsqmamm0KBWVNdSOXVsWVlZSFh4INEjKO+l5gwEHLaTT
+A94RdV9DMHI2hCzHfnR0ll5fBNXFHiY5LdV3JdkQ4i0kXgPuRYS25v+g3Ia
Ot0oduw5G/8B5pE9q9r2/FhjIueFnkyQlLKr1Pl+d1Q8sA6pyu6qM2agsGqQ
CJpn9VKXHNpKnEBM5l2+u0SdRhtMkzQ9vuEc68TxR9mWSYxyJbLmqXskrAvX
UICY7PqCK8/ehbIb52Uu8KcGVolvUAgA+NuKOavauyOl0Rk59ZGqWQbHSr0C
8TTLG7pBaUBs0GB81oHS424leWKZ6koZvzOLyck9iD9g+0HW0T55VEw2Pcqi
A6xDPG2k/14t6SvMnZjwHuoTCvCSu9yWM+JttpScjxRXfyE5+XS7hfDcqumr
gFn1R5HtTymV9UNXJlRq/S+eGoy0xuyiDGswl4CHAkraojXxevvw/qy8rmJW
ls5x81MDWYGSMMvojdDTh5P7uGLOrFSveXDLmrd9xQnXaYpuKf79XSoSIIIR
FjaLoK4aXWjN3NLSVfEiKVdhMIGXEiJQYNaM8X+cMIDQ50fMcEIpt6dZRK6t
cgDofpUvIqAgw7mxWl7TA3ae8EeMNh8RsOwaeUIopl/jIbuCQlM1OJ0+G0mX
QczLJJXWQCOdkhyVb7WLFldzRTQ9kI0Vv/Yyyc1gNg5fP1LTvgUooNKo6xeE
0sOw9+l+yZJPx7ht080WZqBWgyQv/svMzO8ArmStolPhFRNUp3gwnJOhAIr8
ionOXrQQeDQtBNh7oVEEVAetuUncWzlqY4Wmo3ScYuh2UQIbH6Dqj3Usrn4S
i91+7lvfaHyHx7M1CO++oP01a77RUrfLUsf9TNtLqhOSsp7pB9CJ4ncQ39+u
x9hR4YiUkPbg5a5vYKRlvSJkl7bscRV6O2rz2QkhnCHQodpAUdly5YwiEDYf
Sjpey04ZkSYktQa8mPTgYKHf8/mWAmpwIDSqwvzHg3sQu/koGJ+TNdsBeijE
M/L3oaa3lvSxQkgP5MzcnqDY1T4D+Bz+Q/Nsh4YlgAGiQEM77O9JalxLG2nA
O3XMPXJDDX8FC1URqI46YMV66BuZ2EN3G3M78w1Q1XLWNzgK8NUr8T071uuR
H8hAYiWbt4kGN9k3wjOJNi0LgX5uWfmIRsVFysZNEmrK8oLwr9qONy8OPzt9
3miea69ZZW4zVsfbYOdjr5SYTzA3dHNEYcjLZ2qqIfB/8MHbXIx49RSDFhTd
rv5Mwx30SN23lUGjflX6cYGOqOWG8Zt5PzRSCHcWfhbJu1Eo8M1in5QOxnyo
G953Yjtr3O61dotD8nI9Rk5m52efFKH202XbS5UFu9OAzc2lpSOXRFpkr+vB
c9SBae3bzYjVA+WFdEtgJqtmEct9MkDdZBOS63WfVzOoRVP/w11jQAZoWhmn
015mhpAR7/P6W2u7qYmqgu726Q6EUIvBL9Ee9Z7NZktV4GsRWkW16NN52oTR
uHr8EKGVB51fG5iEBZPpUtWtiSM0aNq2DGzrh1meFZfmbGKCN+HCK4tzNmu5
vD+sVYTeKSzKPri/j2CvKf49klc5Lf3+3KF56cpc3gF68m3g2pWZfrymbeRG
arBi7TigmFu77RfhvhZoi6dV7bqQ6x3oR2crroecWuw1IkmSoNbaZpeMULeb
SkOJv2i/adPzXUv+SzB9cr3Vjxio6W4bYc8f/r4Jwonhtv08LF9p5xdas/6Z
fHACmfu9hIpRoo5VYkPGgv9eNmuRz5eX7hqN+herY2MMBdhv2JR+Bwtg/zrb
epOh/d7KQQ5CP80R233xI7i08aHONh0Nrh8hqLbV1hYlmVGnbRMKQIX3L5yQ
CsbfGNVxDzbCJciGGZMXLZKKrgQG38QGyNjZybQJQ2xhMzJS3aavgZxZ53Xk
Egq2L6qKJIz1MaMnYmjl0csQo4VBZ0n/kbnny81U7L0jThG3+txB+mNuAt5R
b2JzZ6URZYwB1iIvbk3bN9PmoM39AFQdLMVRPifC7rjrBST3Sfpxq5Tf/AFo
v80UdDsxIO9yDqjkD6HGmx4Jh37PntzNZt43JLjamcAVMmFPMT+upqSAarlZ
cDk1T/kNHSBDU35KfDzrmi3HWI1m7owxh7laQ3s6a8v1PWmnrSy6ffvWJDoX
O/ckDWPtiFfIc8PuenmCdOHsiTd3XAnk/7DcglMC4CZ/cqEv9vDiQj+YJTyD
2VexbWhoH3mXDjifH1zKaLV5EcrldrwB5Xs/tKks62n5WrnMzWrmsapAMYLE
tTp7iHvyU5nzz7WbxC4hx6asZzBfX2VVOA5kIXI61a/7mo+Vk5uc6Z4G790Z
VRVtvP03JzFVXFgVu/4+eemX+vqqUiY1mr74yww+ieUx0Qm3hUR+xwRKHE+P
32YaujIqEWuOgVn/2uyD6v5tr8hzsuC9Bnpyi50cqA0GvZKFBW+kGdQ8glxJ
PlqkrVs8Oc8fcHrL5TIvuXCTW8dU/b0wlasWSvlpYRffOKP1C6xPQvgo55Ma
Sf6A3Jf12vkTNJAvQQ2YtmjaylI0Wx9MPkpJtR9AQx9PJETa6oKxamn/MGIC
IVgRB/g/XjYtWzX0EcEk3g2a7S5jvhMmYERshHL7RO65fZjjUNLPWCjqZ+Of
ASp0wEDgIt4cIPIybXdwUZBqWe9fT+bIWrdvNaiS6XsZPRtaeZXT/5oxOza7
52T7M/S5qucWfEeZZEi3J1eTUXhQMFd/Gm3pOzb6j02BsflbpFRjQAtoCysX
xl49uVpPSR9mWFm8n6E2mqCJbrV+s4qdFKmSTsGh1l281FMBFnahG5nAtfHV
W+EziQBGMOWDe3Bt9RPrqq7NuFPRegA0nyVuJ+4X0wYNbqGGduRUskxG5wgF
v1MW/iaA07IvBWuhG7GeersjOcj2l41B5ZcBsUxNIox73+8CdvxXuGozXrSt
a8P7NY7UY3mK0rojW+YbZL84sTEtnwVWZcfZBR8T+Q5JoqBvnnGi2KoUML2m
2NC3LipKl57YqAPTfMTKMOgegJrf2+NcA8xeg7Il4ocZpblSBTeQu25a0sXf
sE83vMAZHUpVvNo9+CmKWZq33kR9LcU7RNRH05Wul+sRCWg+464zLiqH81zw
Fpfj2L6hQRVchw2FyVXe8llZWgqTuqSZ+WiL+bfjkzZQyle87neqBs4hsmw3
5GJ3qLzdFtPoY/kZfYe/J1BgC8mO7vW2kwDfSqi+4fix+Z+JYzMJSLdfRY0/
7kxHgZ5lvbtsYvuafLjewDdM3/4PranDMtKWZCISsW2MhxZshY7S0yd+/TOX
+gNMdVQijBt1SiaqH+pga8Qzz4aehti2z90QafxVMc9rCnImGfSXCcy4Pukx
R5BNjLvrxauegapPdnMiZdrbvFHtwN0CkhAy60r0pNcjO+vE/uGkIK+X3lMT
m4JOogzW6UGiyCnKr+fmlZd8foxzVHQEItB65bWl7BHhQmALhxlkV/ITgiMY
+6SMwxHarkXUlwATbNFpBVQrYq5R4HntstS4OMtyYbbknQJoE5UQRD3rifOA
e57DzNrGA2N5/MSdPuqP9pIm1wK+Vh4ilbGPXsYQvBdlo8thU8lBBLH6abBI
2VGGPmyjr+llQwqQygadMJAEH4LrtBYLKIlx7biQSVKUe7N9rBluSrd7U1bW
T2OPtNTWmOojeVDWbJL6RfX3k3rWFZnPxqZ66jP3xyBo1D9dokDhlrzLrzmp
8nmCmUkJlDHoWyoWW4lpFwre5aJOiBDkU02LqlS+HrLQSR8/qwstb0/aZqKV
bOwoWCP0z7nQLhXkd+5jYSkMxSz9fSVSK6TIR4I/QVlMDX9HwpwT1SEI9wW5
7Ja2BuJiqFqscY7ACf8HbO8FHSJuFm445V3fIg8v7jRT8wXL6ISwZNT3F+wY
8HC5Hr+WY0YHQOuDjWMnPZa5g13JzdFTjbqhwU5m01qtMEycBlsrVvQ6oQQw
bKZtSYIj+/Tfos3uosCIp5HjodO507wYoDb53/fxcNRi09AfampoM7swljLA
9ybNFkGeGFwY0Ng/vN2kBOKbEM087L+ciYNhMxpkjYHLNQnZzEPK1rAGh2Y2
UoSxeEv2WLPZIAdluSKbmFswC5mIcolZ6nDP4LGvza1xsjgJxjFypXJvdzj6
CnhO3NDGvXx5rBZmKsY3Zt/dm7gR2M+G8SK9OwbYjYUK7PCHcT7z8JWyY0mn
pWSChndnngZDIBB4yo7scIY7dNMfAoNeppPD9MxOq+01asOf5awr87iqr1HO
m5fgAw/vVkwE49yIhTro6G/4Zi2Zu5FXw01QsU/0syg8LqX9O39ezAEePe4k
ag1/EFv54bo5JTYluSaNQjit1LPKughlSbi06XDzB3zQ8Y5bCCdtBf+pbqgt
4gflGrsBQXKeFMNA+8e+XNDwb25+kuRjzgLzHd7AeJze8g70Caf6cdvkIGB+
pHzDJrHSUF7nzX4nI4p1iOXKASbRkBZu2kB+92V24u9MIG+VVNLZnBZiepwR
33YeDaVPn84P/QBGSHDaFtq9NS5eGUqlHbi45nLCCHTPARi0KY41IHjrPHQ4
cr01ggWRd8fgBVO5P8muMWZaEMf08afviQthQzzJlMX6OlR+DF29aWpZmYmA
QY+P/52Lztb5iUJXovgJaJfIuT6YRX0DOQVJ1OpMoEyxM48uwdW4c+fNiZY3
vomAFlMd464NeLlZYgjuWZEgH19YbV0nYPIEVNevbkjaO77Fw3zld7DiRBm3
1mdasyGNzeRRVzZw+v8fDhamg9AgjDSQ9LQcU4Iii6CjcHfWS7StKmVstdz0
UIYnDxQsqHr9+jTOHq8u51eYglhyk/FJdlM6fxPxolHT/DLt3eTGi/E6QdfI
CZ1ORjyUUePWv1bbMR6eUT80QGCvw/ZujgI8LrPhJbm1B90qL2wkYPSnza9s
ENk0S/oZkBF5XKbGApNcqGaO51xhDE+9zFJ7EbGfKbKWeSTAHhMv5LgiKiE1
rwb72mpaXa3JMwFjcycvKdmcyagIRw2fexUeoDrLBsgLAEyusd/n/5PZGgCh
CILWyjupm753DVyRMBC6UROPh1PsgQijwYAJlm93XxGxTEDM8Iolqj04oYPI
UFmnsC4qrjFf+rzbr/tLL/E21ohMLXAI6RBTDd3ra7UG9jZpi8EVMuPIvhSc
I1R9Yb7XluOMOsC4rZinWjhkBsgVLZo5tjs/k5XGuoUUpnwesWEy8rvE1tFi
X1Kf+W63ZyiHoRgtlDePvPYPsaotxSDgAZnXTJs5zAjsENYVTifmVt3Rrtro
FY7FyH7R1w3WERADLHj/IqK6VdcCSmqEhF6wD8o3HuLIgDI7YB1KhzWKGQ23
/lv2KaMfgkL65YMsB6r/024fwqNxUM/vCvCJ/naoYWJWDRSAr82EzRNtSLiX
CduOF0l/6h9U9J5MfdlgnMPDPJipJ50e7YFH8maXCYbTFr8rGitsvnb3/o4W
aHxbYUI74DaULFAhA8lBWHYU/gQpJ6ofag+SQIC77UJbnFzWTLht9hWxr69R
ifhpMWxCEuRrBv4uh9MDt0lswPasBx9udlwpXb85p8bZAfcaJJ4IYstMIgs6
s/XW3CNhJlJo9c0R8/9ZDH3GKA8StfuiJonepxUOU7UC04TpoughSHkXUKxi
WCYbcNxwnnqqLnT5MLGTu5IS22sfLrYSbJ9jVwyBX8pI8li4nI+BKSJoOEpZ
ZvzPe0KOtjbtWcFl3X+SUcKzeHiwsbZR0rJFFjFCxMTBMv5g7LZb8eu4SvdO
6lSafPzjok+iVPP5iPIDpK+70DI+LXcvz/v62DkxtY1/BQeV7vEGUnr8Pftq
UX7q1dz0Hjk/9/6aaRi8zWbORnuHKt7J3eEwWVJa2YjlB7P4g0RGYe1MwxRm
0W11fikZ4BuKDaOcdZ8l0YkveZkBlUfHCgiLE/DS+YxEW0zFPrDkhGpY+Pyk
r74nBRGBGZ4Qx8lL4K8UlTnIycUFpObnwqqz/hyIw7Z4o1aJLHNDSkrpV740
f4qbx/SrfHyCeaKIP+rT/1/7HJSm/PE2jtG0DJMojLQ1JIeMP44+SrgPf8w4
PGJX+iuFMr7F+c8bRDlYzS9QUAe1wnPa9eiRrIQBHPajEVu3vAOuzix8q1Lp
nWJ0ntOEmfrtNpqX0vVSDI1u+ATkirGcrHqcJw2ZLk6i9Nn1x6rJ33LhKTh0
24AfqSefKxCLi19uUsIrM9n9c6KaPAb7FxVmGi/ELvGM3aiGOlzHvsKgJ8gb
PVwWk05nXcVX78L8RYyLA829pCpYBK/zDBFw5czYBAJ92X/LRVFxlzFyUJLw
U7dfRW8qN6EIQCCYX2Bmua8Xo/3kbajag6+GxdOYZcvCPfPBLMqPuWzt/YoV
Y6ibs+LMM+2oI9/j9eqqImr7i+9dJjk64fqs4cl7YVmryI7qpJ7AnBrzzm7X
9opVvUVWpvEXsmR/ZYgqSFI/Wk8b4ka5I8SyuI2yt4PmExS1JTHDlh14YpXu
pPiw1n6dErXRePK4cleIWErr27mJ3rEWh6KPnFbfHWrt0hJoy2PGoRTVoBTo
S8Ct267bozXeWCbaDDnipw0lxpLD4jq8KNDTMiJ3YpnJug6vGq7U0Ajc1Zs/
a1UpZfDMViAYQNiB4vhRVzZiE2nuTnCAIrFl8Sag0j0fEDW63E64grQSZr7M
l4y5k6qZIkVXoPxxo0x/ebVnEu1dnNcVvVbzid8U3n+SBJYFwJfUjVo2IwS4
7QjZCfx4J5HCG141uI3pJJcEsKV8KgyvLOOWQutB8g+L3Tl3iEL9lPbMi2y3
xWv2dkoBwjqbcLgKaSIEb7FUSrcGrTcwBBzthzAdAc8flLSBd8vyue2wIAgt
6k5Qefhf5vj0Tmxu2JWpLqboyikZ5xl7tDJRDL0zf9tkOIbmJCIt8GdEMsh5
O7rtUhL0LbB25xa4uE9WSpZAzU0bo6cHYl174l14Am6/VPqZgEbBM4HgfesM
cWPnAuecmYFcNY6LIPvqwl92BIznach3TF+186C0wEk1Qu4K3kcL+IfwAOKS
CJYcK2hrlhMX3fyTNfOUwRxVNxjUx0Xc6C+vSYaTsR6sTGbfdM+DFNHF2Crn
IR8NrM6EMNi5J0SCnY//zr8IRq2orUeGn6UpDZ98vnk7LgNAoFeDwu4tzj4G
mjHODYKuI5HvrL6IDxKKtYdBZTc6vnevxOPIp8UAqEbWo1cqtozP5drO9y4Q
Z4ReX9dJnyt72e4Xsg9MCe/NLfnIRCytjRcPUlrtFGbZxSJSnLrd/MJ7eJj7
w/+NbvgxzE24k9eY2710PKlGPlRnPDJ7ok9gQu4+LfEplD7ZaqSoRYRjPs6Y
i5VtpdYvecjU1zTcaLklN29kZcn0DIPHPek6I2QrgOrz9h0LcJP1ldlypJqk
DLZJ5CW7D9c2FwzALxnteQVL18fVfRoQo9hr4hsHWUjhEN+a54hkP7d2vD/y
Q/uAqXPdiAHyp2l9Z+z+GxC4q0ZFSUddI5uaEsUCLEHMyyOUAmOnZzwBDzeq
+mgYA1tfQVLEt3Td3sWB7eBxbqro4bmiEqCEiuEF8tfPXcNHPFhuezeutENG
HuhOcFJNWYyfz0nJJX9Iw31GcGY/DsYRlKRbmPzOWkjLgXeD3n0afLBodJcq
sRpwZZnGCOUyQg+tUtujpK0X1cBBDh+Vt4gFMsw0n9Gl5Q0GYT/+WSEqepiK
OJT0ujIY7/QNVRfYvXXTLVwOaer/6wfDbhPHfDwYtIc0WtTDec+A9YGi0KSD
5/qnyETbjF2AD8rgsAVJeDOUUVr28OwtZGk7z4vfmU5D3oAoLoi6P+IXG5+N
dx6RzX4g+NLG2aKs/RNUx+CnbUJRYcWkRODtG/oaXS9idD4Q/L7ZsDn3j43t
h7tuwEuPVS8OAueJgyL6dELdJoDjx7tJfgqypTxavI1oTZYjJ67/hv/eR3oJ
5qlQePIF0e64PmV3YBo0HqWsPogDjCMi2Lf9Pr2Sc8V71mX/5SC16Fz9yysg
zzg2/CWDn+gDqYl3+SAHlX8/5QrUP24p7KV7lcFefDR+veziPiU1E1jA0y93
Y2cUekqw1MRWG0lyc/ckEGLzLlqsm4oviRdTRZ2UVNrfLXNcldXcMR4Mlfao
RB5oTy8NGyAF3XGew1ORPyzfVWP/6xfNhQUiUVSTo74TwaXYY6pqCuOWISfB
9Z0l8VhCJya/QsHzLjNfy+WMApDzPml1UO8ZUXxMzqEQS5uFt761+w3kROGQ
z1ftVmZsegPOCF+Z4v0fFJ31Uf0Qnn6VImoiLhyEXW0oNpQhhiJSQ3BLVDsO
LSTNynApl3d+K0wQRlTKLNYV9aFcCHqQsfoDJwcqrJDe6f8vsyDa1cnvz/cH
FSVsX4a2uO/683RYNyDzP+1PVn1cEu0tuww4bLIdGWc6iwV6laGImeTWo1su
IHBPJZhJXciyesM0+Tk1tCFxRWyg2ZwBI99of0n16TQg6JJ6JHAvEmSpNeCl
Qrn1idDTUbbbSZSPPD/GUalksTr5OvW/Dv5Vb9KcFqcSTxPCmyzjSJXEu+9y
bkcqEUo4Kp7P7W8tCq0LyrmHIwos5twD4JzHSlKb53RY1oIdEu/1Eob2UXOP
GCK9CRj+Yt3r0mcDIY8V36UGKLVKQEd4PZyh/SQDnZkzJVkpWr1O23wWdnWR
jairXP2jldIciOayOCXHy6F9DlQtX2aVxH1WZPiPi0b8wH9tVLV4ronMaPtZ
WhtMs6HyGUPKwAwLPIcYQN2mPFqayKvgkllFD1sR41GmlRFEYcHIb+mK6THG
dF2LtJ9MovGoDKnA8896FfaoCd9TLPnaup9rinrwLBDFc+z4JtnPADITZhZ5
aShtrL01kLisyelrUvXWO2L0m+zfF4RsGRVVKbWP5uQbIKQpZU+zXdfCW1hG
z9ozKS8torgsPBmq1GzWavHdbG3+SKwraEa4ieH50yYDIAC3oigoB+psMcrc
cvRNN/qP0V6q1vciKX4U+sv80jXVKwICZICoBRFpSbNHAT7oWFjgqzX45jgb
49scFXYUv4wPBogMIl1LqxP+a14k7kmRBHr8B64B4NjTQEPoXLvtIcTag5Cy
tXe/ATuIu8SkbzDAdyWRGsqccWhxDGHfI4I81u1159zAyeag29D4p+VP75+X
7f8/+lPGI0s/5hwKkrxttq7bmDAmhYiafYTmy0sc6zV0IwTlvSbazbF2Qkle
WzYQ1sLU8uI1GZ7CBA5c/sFxL0BIx+OFmoclwCqXmgDwZ5B7pKRRdccdZ9eR
phtpXym3QH1WdFDg9E3GIy3fY8GhMCdRg98OWzvzjja40b5B5fe6W7iZK1Cp
hWbUpjZPYrsQJVVKZObCEcwU1yPeDwint8ssskGe6iLjN6Vh+cHkRVIFGuG8
TbzvX1eomgCS6EyvBWP98gPBuVJlOddGPIIfXo9+jadA0GDmoXzXti9fEPsa
UZ7jNDyCIbvnrfZeLKAY7QzmuLQ0/ja71aGPDoeoLhsTPTA5n+/51T/peTKI
aYLM3NVK0smPQZ32rti6vFFpIHJRVniWKeDYAxbxq9FpOF5wjX57422QADGY
MZ7r2AnEhnWJ8INIsEzCXUFmGgxGAes6WHxX/H4Oqj0sXzj7j8WnzLUiIbms
TNa6A4iXNNugnygiqMBd2C9dM2FDGj6cKGbXBHp76Twr2JzfoAG2rOXOvNw+
Wf/nxqOXGTnQWUUQyIIFOBmGQJVFwjtDrSM6ClQVsBfcFHJf1SyyadahqCWh
2jgon5QhEgR5kOEzq+1C2nRcoPfL88v8C3LOZ+MpkkeGZwepgGUhh2etyPw2
Fxta04wX93LYnheNjiucJzTIx+ufD6XlY872RahOJ7tLFGvfYQaT1C/Qo86D
MEDPu/Dw0nGG8lLnv8Gr08wvizQrnLffVOFDMb5QI2YrfzGgA2Ul9oilLXvN
Wuty+8saQ/PKq5DpnsKIvhcrDEGb4oSQUrXIQXS9ystAunLZpRTBvAd3vN3r
aoBD8ho1U1P5cneAU79fe5MytF891cxFCw7zJY93u9N6isBMPqOtfXMUyIBS
d0zNQ8Jy4y4kEiLHFypRsFUI0cQ8m88ChbvZwjy8SOJ1XLY4+VUJC1Xmztjz
h76lqEiGK8MvK+erCoRNrGyuAF2wpe4am3kHkh5Q33XQwhwmdfYgEkX4WEnY
gHDyel78iqFMtwQkFLbnCHjYSpi4flHgIzqHe7STX1IHKXC2IAryj0tNv/Gi
r5ijXJXMuI+rxrwm2zOFX6eSvZ6tW87nst/MuS+IKVWTczzPHJjgxJp4Y6eI
1pkxPWu76DJ6xcmq76qbhQcqNWkLVMrcx0kGiOnYz+l4LzXiQlcFXXq1I40K
W8RnlVunhDKL5O6tFVv7dzN9lB3JHJXnFMVPwqhceS78FEPho4bfRdj3A7j/
Ujp+t+x0grUAUv9zpX1+aonzqrkWpezCo+7LpXvnXEJn7UDpCOGtiumT5wAq
IJOGG/r/zn4mvYKlkKyVuSnw6bhs7buqBOOkXsa2azowFds6bUJiNk1LjbVP
s6ggq+lxTG07Yz64nRbQrtrRqmxI1S/NNC1O5IqHv/GrKiKOLhDtim8aBncJ
8ymNcHlHM9gGKc1g39NiA3gmZzWFaS6T18JNy4QiuXtuVZvCjyo1hTnAc5jZ
GytiTBiI3LFAqJrMPJwf11A1i6Fs1EQFP8UL3mJkbNDOySP4wU1HJejyaCZu
bZJyXaYYXGQHBGL7hXqKel2rU8iYXkRWixcaq8TNEueDUSTpVQ/n+KX++5V8
tQim1BJh7UVcxh1H2IyyHRw+jXYjO+X3z80N71G03nVOoRKG88hJwdVqSTzB
LcyNhAblI0x8SV6eArqnnzASA0un4R/oqKdfbTBay7hypAxVKFDk95sCu9tS
lCS73Et/BH5J7jA8VosOaY9aaoia/9cypHRn9I4WjWyrPrGkJRJirAVZ2bVh
Pve4MpM97gTqDsoxoWx4AAEDIvaHtkWbL71/tl+3RvSLFkx4XKCHsZ/6wLs4
GpraGulrOSk/n6D0z05wD8g8j0Ufd+07+ycCRmYq0TkEHgf4Eb1+ziXoJMtU
SoWFtcZm+fQHebtFGdWsUhrCF5XC5or7knUy5II622UmdThrxgDmPJ90Hd5Z
CA3p0k1pNC6AQYt7Ulpa6sMOBEMl68RESwNzHIe8TNTvF2WTMEzP0iJNEddl
N59sAC7CLU6SPNQ7FG+trwQoi1ocAzyRIVR1F+hozix53MxhXzq4XztEdvLz
Xz8PO7gbwwtL02Os9kRkN/gktdPvlNNXzhUVUoVnmG06vWIqCBcZvUAwR/mb
n3L+RB3221W/t6RAEX2IZAl1Z2UUfMiCDIekjnoGTfsotYMCgA1T0rr/hdDX
/DkQaqaqyKoDGWiQ5Eq4dPpfePsK9h/ps9ShtHWvtMJjDKvboWnLMIKjhv7F
zxxr35Wg6/Y6qEwb3CS7YgCqSwMw/cSouN08rjQUG9UCBolHH9qcb6MeIZ1d
UXUAxU8vyTN5h1iGvJhQOmt3PKUp6zBcyWPxQfubfyICrWgZ03ZgdhosZ370
DLJKcem8kWOSf0+ofKM+VSsByXCjKeAIp9McQq8I5GUxwJd8lUmxuXYwT7zO
L5Iho1ytIqrMLmK0Vg0kBvaNgfkeV/H8SD+QJtnMAuZbxTyw9tBB1W8aciv0
z2ySwx/aeT8xtpgPop1YCU8cnwkrJprMh5OREg1mhDDwgy1NlAyDbCl8XbJE
ozd8C7OgUh0yE0NydGT6TPiykLjmsqozkVdWTkfvJnQo2oaloWaR316U/Ae0
j1PZTjPzSBYxmm649IrpGhBGcRxgpDjR7aCIjNOeevcv8mvC8qgWVFpA2h6v
citVlu1UYxHJQ4GMLaUIiosNryMibkpb+XXi8UJbgIPBx7GOzuwwshta0QSy
3ALhZbh8JMO75JYpFmrOcJyWDdW1zJAuljno49Uby7H8T/I+sIGO1CGRkc01
ZMDWwBVBzkhrHd17be4P/4WejEhvqMnVy+hB6NVVKcqvXTIH3focbniHcfnF
mXkMb2xrd0yOX4+PCiTniYLnMSOyFQK4hU43BndWdV1+HAfTJ1PZDw6nxGT0
1W5GNtNOvnsoCzL82p6xfASVGLOwTWFXH8HUN8FXd2TnS+MbRpIZJOO0UvIQ
NPB0feoaU/1O+dkeoao2yyA1VRpXkR0DKxwM1naDaXtNGCH4qytaZsjtlAH1
4MZMaiZJK+cUhFqthVaG/6gZKKE3WmMMzrgyxcQZVeG9YiNbNqdA4Wdt7V7G
G9Q092B3MrZDqbsxPgXZRME6MOPeiiP5ES4TM9G/243oAM3eC7tFe2pWtUji
SqNU/HoJiP8LWp+thLEdTri8aYSkGCktkFNzqb+lEhOLfwq5V7vJIGWgJK/c
4wWVlgO0a2rzcdDDyyGI8KtdB4DtM4Z+qHQyGksbQ8NAKx7UqUK91Whisg0M
AJ8E5rmU9FPJh+g85X05ZOTky/T7LUqr2/SNorJBdKFawf9uUr6AEJja68ot
8c5uMfV56u7PndHLbsiPntkijipWKPf1Ikw8qp8lhAByytb7jeyniIJ1OMgb
BG32hGe3pgYx/j+JnzdKsWyv+i1sQjpErDDu8OHg1CTe/tfx5mLOiEgnF66m
qOqEchmd7jq6MHxeP8208EBvI6PWft9kvod6eV8Otq1UXprbG3K/x3Dx5/rP
i35it1d7aW2vgllLZvki5KoLP9MwkLghXtd4ox0/ZEgYhYe+yJ8gXXNvwZqz
MB8hEMkz399oAWX6Z1ppiFEBfn7KkIkJ7qjn75jcshJLgz+OzHHLZ2c3JGBK
wBByvPPJLcguP7+CIM1H0jTQgBTVvy/K2GLf3i/TYgAf3Hcns4IwFjy8nuYW
SgR6oa0PrWIViGpckTDNGe+Rz1iVj8iXkBRoKvA+Zw2czxMH931rebn3/nD4
p2tEQPhUDRItksSL0PBqm9eYspSidWWkhsjgoRqed+PxefR8BL9Lr2co4lNm
fJsB/5XWzHpsivUiZIpAPe79gMu22pt4FQcRlNR8b5ncaI6X+1XmmqDNqdMg
ER7g3jujNQsIMWkx5YnSiVLy5LcEQ76CprI72pGUBLXbrPprObfNqTAspT7m
4FqMGHunmuaD4Luin423gjAcqVEqARu3Tup/ulQyK4Zieo14WxrQlEMNn8Hj
4z5wfhMOPfPML2726sFx/gjxVV/94g1HNGvBQFzqqa6ZQe6KW5jtDCfWcl4T
Z+T3DFEnrKTAxi6YEmp8YUHwq7wZk+Jla3+VtETZCwHnWXcSVt5aYnmiWnMO
GzVz9sq5RiZnMdfosmJ3vW4vcgDmv2z1mF2wJBpW4A0WTh7g0FPrFWM3fKRK
dTK5qPOzjJcsh7blfh5FkoPG9lhx3w9o1sRtgTrS+JoxnHhwLol8vzod75Vn
kVn3Em76RKQvfWk7KjY9A1mW0OMfYN/6pl4fo9eQNiEpd3nXL1lfOQfgL4wo
iYkEE07kMf/KYFmc3uynBdQCr54dsdFDMR9V6e2XLeqZXSnDqUd9AGoZqTa+
m65R4qY21bRMWhJEKqistPE/UwcH3dfKCCIG1wLEYEeH5haS9wv16JVDCkAU
gZoeJWmKwM77dQVrs7PAKO/fCbDPjxk8RSbtvtbxuKU1odhuW+O3fLIR18pJ
AVoAsPlhYNbKp7NOiJ3gzFXuSiPG0mluo6PNQ1nVUd7Nyp7rgKFkW4s+rsGA
QX6k4IO+splzn5hNyVoNEciejYx+iOgDx33yBxbrVCb1x4+y6GLq8f4Jc1Xe
1oV2MRwtS1PiCAP0DWx0ynJp5JYBJ5A+J8mlpezCc6OluhGt/OCmT3h0Iuxy
UfM8+NPx1xDjM9AcrGPnOeaBQ0MCokEWDBJpqnv9Epmw6u8XQ8OxrpQfG06+
o3C09fHSteUuKJFc5xwJNgT6odQ/+htvLKzatCJ3p9yHXKgWMeTweXpwTGyF
Yq96PQe1I2P8Tsbc6y84HUmNgvB2z/7MoPsFRWeCtbHBf3Gw1DMwMZsuSUox
Fc8Il6E6wWSAom5SLdo+yAEmabfnnO4Wcl3pd6/2J4CIPIR/m6qCG1VIRWI3
3hvTSqEUOVTj+QTbYuu9nUPknRyGCllQbw9gLX1dDB3w8IOOEG5HWAgBWR7A
qa51sNnAWGaNvafYa6Zt040eUVeXQzqQIU7ofk+elR16Ik2Csx8oW2ee5T/I
ODsOOPYAmqEsBHx4vW6zsABUVv54PGStzD+FXdmYyAq0p6tLJgF2ZHpRBtWr
Dj62s/9k9AFIZmf3fYVJOkAYB1WocE95TcUQUxNWXLh0P79vOwsGK8XScsRk
s0lxYZbgvSYliRHAX2xvJ3q7S7zaJzi+5GcdJawgx1TrR8TToqGSl9Z05i19
Z+XCbsALLH+WZ752ivfbvsBXCILamyoMOYrZMqZ53eMG1QLfAk7evXVTYw8d
2SL7dFeTpUm35BBW/UyiBRQeZM8xZWVg8ejui1HBXpCsdxQjJiqvtWXu6JoE
PHe7rIEupYrGuvCo7VgUnGsBC7UjxdE3Lt6b90TnYS2VzI16Rhq8faKkPh7i
pLO7dbiPFrAmz6wsHZeeGq9vH0mw8cnbEcLBn8O1lXCrkukz7z9Cufzutda3
6dsOxpyAgZxEultzZQikaSmGw6co5fRJXn/vBpF2SE8tuGjE6vYvNhtV1IRc
IippDXpVlk4X3msTDtMWZGjKylFND3QcziLdnRvpYl3Cq4LmVKKIgfil0a3Y
tQ6aiQp/xdkQjMQMPhan6T/WDStRMb87K9kMRcQSeJzDOnPjOA6kW06UW6X/
X9M15GFWQhpMuEYEu42ik37GOLYqhpGFycTEAUQ3H6ygJQM+JjJBnp94BLwn
pu+xM6tYCdBVJyiZZELYyEKLcu9CW+mkdcHoLRtf2+KtKrikdJqTAlkWBSXG
ZuhpIGLfwkXix3D3LH7lcqiktPdJxGUvgbz10Oxe+LjQOLMjGW7i3zgaNjZx
V8zuk21endDrxvPOPBPN+1P5RipFwP9doCXWJ5jmpc9yLLvbzogpFPVIg7fa
EMu4BcrRjArdDAUan22oUA9FG4/xAIAqQVCONXuxA3J6dmOI2AXeUmQmem9g
5dKIImc9nN0RTATKFxY0YgTO3dBYwV/NE0BTjycvlUfhbPvdl92XTITzMpP0
YyMxeKC7FhdpAc7A1typ6p5l48eqOT/JHcPe0+jNedoVcIHl7sr9w7KNuZVU
yemIjDGeSD0uNx/JuzRh+++6E1GV75Sk0RNsmOX1TXQ4BijlKzOT+6aPhjab
fJpL3EALzUTceoJNZAd1FjVPZZ0ojr3pXqC/gX5FqHL0VtKfmvbsKZ0NW7aJ
nNvubZZeSKjEfa+p8Ep5pMpO1bvTkLLjZQw3EehzXn1r+CmEVPfgvLlKf1gN
Vd2oAJyFrOvnFV7o6VqEGnIJNcs1xPNnXimgWM1OfdCgjWlBVz8eWiOaFD+Q
Fczg6Ohwkb3c5Dc7XB4zM2wYTUI52ugyoXf4xyMqDRlXLbbstGhLwSM/FN56
UBltJBrtWs/2KUgp1T60EfF62DKVbbaGIks6WoCF1pSeN6bw6eBwdHvfjKhK
wjsCF7wn4VDeeJiyu8zdIZM6Z+Aa3SYcDTUyFg94x9qcC+WpG8yEo+xPEmUC
U3ds0WDrmnF0NtRmKyYbVU9hctKbRY5tDQ/KVMo7DQ4Zk2plyEjLnrJ8nxYu
cNRJpx1K2Lp5A+aCdtHxj9VvvIOXuMj4scsENDTRQqD2W3OLmLMxxDMqxr+w
I9xT9fdSyTzV+d76zRpGHfpfYEqLsyTjlBpFnpZq0onnT2zHU7fSUEVn17b8
qbjOF4SRpi8SGFk1jtdQYtfHJUiRGKMXMlQxCCrnXrjAK12OevO1uESu7o+7
Bql/XyYhZhTI3ufVZamPNa3reHxv6zBg96VNVNVOlFrSLxz7kseNOezD1+OM
qqT9SDpTFUGHapBIxSzLFWzk1Tk+Fx9kgqSwhM9wtfQvp52Ah59PxTUPV4NZ
jj6cX+bizSqmxCMqFCfNPwvJSDdX6+IoX8dopEUQ9G4bRpBzclG1bNxdRdpV
tux80+CdkazaENWgmVTWaACnIQixPKUwJ6e/k6lPlm7cEZf8JCDSB4M+9gV2
tt+s+0hknwipA4Q+1tV/SM/mz1Rbz7NYs3m+19mxDm4/qHTajTj5t1umCgy1
7+XxFxvSakCs2EGUPAl9jmjtkOALpucHh7GfDUtjtUFAgoGgZrhxl+WbwFYS
w09G+rAy11BVw3YRl9XPGwZtEpcbhQllT/fSOub+qAovmUgxP0RL2MNgkd9L
+INyGLXC3+0EFDSF08K4UobecUVkIZX0/x4EP/yblkUI4DtalvkNCwhWGKVi
gamr0IdbUwEo5MxECfJZ7dKB7npN3//mARKmPmZJ/i2+GUjVkkYXhrIRzfwc
7PEMT5qEPEvmAEcxCpmCx9wZTjZ2h1V+liv0W0vLjE78JGWRwSmEqPQXvDZs
hobyFQAN+n0uvo+15yLgctWO1ftVj2QWW181YNbLRwDQKKdOXUXIaT1OZ1KB
m1D/Uu+rD0Hr7oR4AvuILzv78dtJYv/LXXJcaQj0BO9woKVGgioL+TJGfjrD
3sDHuE61CGnCYTp2pLVDK9UbZHgcYJb3snBjSj1YFn7QAS0fXmbTOcl3Aqlz
9SndNGxfXh30Taq9pJn68VLHpFC0Wwt8cUNtNXVr6mH2BrXsW0iTFcTxzJEO
vkUTIqzlEvgetvJsjVEWMBWSy3Tt2FuP8PSdXZK62rAr8gvC24/AEBH8i4Wl
ONRBLF27vlEaZW+sz7AP5a1R3KNQCrC41cMLod99zhWo23qTWdsVmcJ/0OnN
o1Hag8flOLh/RqC1tBm6Cf81a3nOY9D5STZJIOVIgUCLpTK5f/xbCz7GUzVi
+Sn3WRzkgmwNOBzu1yUu7H1SSQqk0uU3ILAHxhK/ye3qDmQyPcx6qtWomIVi
vQAS+WLKrI0ouGZX9kGbuGkWHwIX5n7jkTIT/uzBdeArAiNXlHd7nOc9xcv1
usU5axIVxhnu+0NZNLJ0L+JN6vbrENKsK0DqntWjXQueBWDu81kLI7hPUfRe
jZaSHzX0xaSgallkiwZPv12+LK7CAGqQGVZKKVIYDDbOK1Tvh1pG/x+OjWP3
ZYwMhVNBV7aJuEt7g4ZpluvP6Fs8FfHaImuuWmKc7VdMJKonFL+z2+RFLZ95
sP68G+hQBJqGU3uaL+Z3tPm01+OxwIgdBydcA727Hdh75tNv3+JDyB4Gtc2P
z/R1r+lCIkdzbxmbUaLPLH1jqZXkVPXjQl3xrtxc3Mr2kaQJ+GBMd54Sl8uF
iU9uM8IQ3VwkMZr62SYBovwPEmJ+9dPYTJclzHRI5gMKOE2SSygzhECbuse5
H6/I51VlnaQ6IuVMBZkLzDaK/GVLeJ62aFZoiT7LOvqLp1g2knO6MCgJJCtZ
vTibAkY8Ff+crQEVmzP5Cx4Q2wtZGiBgs+3NPkGUm7woPm4RdPdMaQJH+lLc
fOrgbSNilPkg7q6cjsQtsG0vgxIcM0wLl4JHW7aRCTHf6MXxZngofMC1EUIA
BX44ndOzKSfCdLzLeFC7qWPyE6B3NTmSAhwraFNQXPrcbrF/umxxL0qLPaUp
oVOR39g9GaUfYjP7+yaXduTrLlwXLF6NXslMenDv6ChypE7kpUMgY0b2sEf6
vc2pb/iMUMApFE6a7WAbIXf6hHqgNqMYoIgiwP4pTnN9OUyxjK+1DiDj3TfO
mZ5XWKctogkvg2sk/9ezwr0gDD3yWKfac9gPQEJgBSjs5geu3Df9IhWBHKAc
2Fv8yXN23gIHcHzWyY+wuypKFCwv2scyZ/i8qpB59drV93txRslRFqzeFkO/
IEjGaag2/OfMzbcHfDxbaoDJUrSi7htpKpAQ5MBe3K+E+fTEWk+Qo2ADTIoF
n9UMhf+redjjiaoh/EnjOYizsOTYgQn8qwJnbMmztFzY7O4lTg886g8DavEC
exQwLlptyg1lz0VwULeQWLmy0mAHLKT5OlHjn91V4Gq6N/B09+DZEQSM8MrQ
z3gSaCC4BZxdDgn3JY8SnMdOvIGd61UPw37vOCBjz8LEdbMz7jwnTCaQ755e
K5Xffc4K2ieWjvkhIATB77Q7hQkA2Wfjtk2DJCenc5z07jcl4VGjSL6mxfJE
pqeNyphcR+HXc1C4GDDsborLp639f/zlM9l6ay5G36MVHIVcjQmM6fJE8UL2
gKKJ2h7YuBV6vJO46Mpcew092bFC3ZccXr1Er+ipKo0hCKWMqgpIvsAxhDSq
7+0rIHYP4Iz6l2fp+XGlnVaGQ8ykbl3mCYNoml/sEal/zQ+8qtusi1b1a5bT
QsT/LrT1iVcTdkMVeEeCdzvWL31GSMfuCJCFViIL0gitYSxfz6Ak5BAEhFhL
y57H/7E1QU7HYCzamZyIIdhMdFCz/mdeJSHH5jN2EU8qtBAhhvImGUeg5KOE
Mbur9OYZAaoCvLlRUvQLCz0zcZm0iiMNvzKUddkUSvQja9BiqyxhJCrV+J+w
3VxxvEXusa4pCVcN618maNUNKg7POeT7QbrnLpKG/IOgV3LuAshmikie4dIx
VnbuQyew2NIu2a53FyBhh6bokMfWaCFCXDc3zowEySJ5vvcYdClaMJhn9cvQ
ZxAHdg+rfAsYvCrjBtuCi6YlvXPZjkhCBMQiNunCSlNiq8lNzXhpggam+zNX
vHae4XtEz4ipBLQ2iGlWd3ys7LO+WZyAIcFeZOM71v6MMTgLFFANfNBQa5TX
DmbwT6I7nq4r0npDBgv0MFcy+TprxZ507NnWAVPgEzi/eGUfgXDW7cW8KS0U
pg65S9WdBRzQbkC8RVo16Ko9rYroWHk/jgfizCc2HvBHMGt49AezNGVEaCkj
dQgwqFYJleROGd+b06XvZUKfOuJuWGf3OtLAVs1xKFmvc4QULkOZg1uJue+L
3nJw/ocTuRyUjG3XM7XpeAxeAkQuD7YmWJllIEYQr7clnnR1YqHopLN+R+w2
myAZp3kFNBA38J1TiSzDtOV8UGhYTaask5p3k/Skd4aPhizEAQWC19x1rESf
yYB18QHvrBpWYmyaFLp6DrmM7PQvhc0f0TdtIGtJrQYjiBRF9SsXonhHRjpZ
IiKAXpA4OMgvjyiVdx/wWuIskb377LTDX+jO7s8cEFixPvoG3PAIrBvxOQTB
fRi0MI6rZxBlrr7Tgvei4UNv/q32qmlzRqGbLLTNHQrI+iFU/uE/gIetKAgm
Bjrh4ZmKQ5zVnVT0zuBi0NZrPLh8i2TIVib0j0/sgEskVmjkbMcGRqLbWXr4
nKBf03cNRid6kAAlrMunaHxR459XkSE9pqxQ5Irz9DTFpiEi/VF4UZIN5coY
V35Hx26A2LjKsta1HRPpAzFKHw/hByBqP5nZxylBo6BwyLC9hniIu5s9giBY
+5Ne4iQ0EUWj9hjWM7IUklpGw7efwNySLcROvaslqOPiLJYB8AVR/zShXaWS
aR11RwWy2XV4oHcquZ586aggh21Di+icU2VSHyGHw5CY0wmjekxIZbNsgvhb
ZJzXXSAHecRK1Y3JdSiP+wGqJ2K10Mf1sMG2Cngr//t1wqL2ohq+jgOUxyHn
ir0j/qOxv2dmDnHaOlHiMV8DZO0TCa35CN8SZ8VZpAoKN32q34n2YXC3QQVH
3BOQx8iKVjjzUmrQX1u5SWd6qvEIAfsM0u9BKR8l0qBeZWKxZRu61O1Jpgh/
D4fx9jAL/2y59PwR/mzPzbAsDcYw+oUjFtmN77IC90liDGQ0r0W32ukLak7x
btFAjQffRMgC9zBfVmswR4vD42ArbEV5oOFNLzUfpA/cH4fvC5hwE/QULzNf
k/I6dbo3qRIhoO2vXMc9/zW9r0OcgJwHF7WHNMt2bOMGZpWYLV/H7d20TYnw
c6D1ml/oFwV+5GxYY4lxo4Ys0HJox1jkCBCjJWFPmwGBAXMbOMf/QfCYlAfu
r82Bt+7Vufl/6pn3H/oAZP4VXkbc/SYYs/tBraka4+jnfZDHfhUksOOdem7A
M7hbCwQ+09yeXxjunVZUt8q5RDlveqt9aHmd4zmXL/KOaiGB4UJadb/PjmMV
MuvazvOi3FKMIhFoN5kLoAS7/6Pc0RBesslrnJWO4oyi+oBjWnLgJ6D7wudA
8DQbQhyGSu19xN4KiuJG1qK3O2LJk+5kLmsf49kodp/H4FptkGCnThkNZUC6
+u/TU8pfl2exKUW+Lh0Mx3ywWWIg1xva0mjR/BuaSUyR+tdQH3ump6HaZpya
n0Xy12jM1i7mTPpS6D1vwUM2UYEL2lvlV8peLIPqqVX1vQ3ZztAZQQNuXzbK
SQlpPs0FaugcxOdlKZGcmwt0ADb/ss1oQ+DyKnoeAe3EFZykNqVOz8s5jaCs
QOEionN+wQAMP4qIiBv0ESv/XoO2dGRTAJn2XRH1q2XXoZeqGBWHBtzbt2Tx
JHri9ixSiexns05lys6irFI/NZwfBTEH1/RkbCp5h0H7lv9yO3cV0xe56JbR
UUbe3kbPg3wGPGwRbR2fXH5z38xydMb18n53p7QZ0ZcQZT3/x9W8sORnojie
bADVMV1kwPCZ6lpa+vGwUv2st5fDg+SMJ5/gC9EuH1we8knkK79gHjifUBgg
j/kiOoRsrZSynAm1rQKD/Hrof9XK62jqjSwFnw9Eq3vyQror/VOC/InMpTI4
lnyzOhZjLHNynAMMAuMWs/0dmhhYVIUGxQzyd4oP4cZTQxCmJUxH48Pf4K8c
JpOx2KbyduQb1zxYqe4W5X/qK2RImocqeLCa/kOLSWE6o2iboPlRjfIjVUYw
z3JMDoZmGpmHnpBXOyENdTXudJqCy/yNoDttMwj1MHluk8279nJkcZ75dYD1
vTnnpdPfyG3QIZc9dg32HEDLzEJxsJrNVsGzoaaIVbC2zl81J9X4BVw4wYoQ
CkJ1tdwuA8B8nuxSIRv3zSelYhHWKCYkyxuAfOXD9ajCQ8eGFj1UVmY827ZV
0Im1LoQ9rhb3XDl0zUhsSfCAFOVf+1aLogUX3VpzwyTt8jQU/WBjz4aD3GDU
WM0xloHBXschJPbA9KIh1T4SExQnLGJuAn4ehC72zz10rbqlpvf2BWZBxzFx
huiE7YeHXog1Y41/N0iw581Eezf6T/FhFfLhufajZMToZ6S97C2sBPSLziXM
DnTTuvJWUXGwFNubplAq3OAS3VVL6aetBy4BCnkdmUyVbfESGasWcvQnoSyW
DQXwTEMPkQI7szNKOpGPE2LuJoAaTc5gpXbGKwCFYTMdkbBsv+W9eO9/SGGX
Jk2MPCKFJmsoj1AWwe99A22oIY2qriSfBGQETrOjq0uYDNdHFUeIqCleizmk
kfpCaIKeKVdf560EGkjRN/4poM6cAW4eXssnagvr5kTF+aAqrWsKzukustgI
oKyL0KOXS2yZv7leoWUBRTKTfa9E5pEP6ih8hxPhgsW4sabVMNl/B3ueBnzm
9HH/p39WeCet5jYJ4WrU55ipd+fgpy3wBg3lKBpgAqFg205nwkSGLDOp3bJs
YAKMqKiFiMnvsNOxWy1qRSh1C+I0qBqaRhCdBm9ofiLjNNrPxPty0iH+ZXrB
A+isyEGYb/AO9jDZorX2WVmmVlahVpxDB5Q+DqcR9j5LWLnEqzUb/vs2nHBh
KFzsT27B5fzzq0NsL5rTzWOmgjBtOt0lU8xO9K+VfEY7CM0DSmkGDfIkjU3h
G6btAXOcN0J11fgUzpjHdnzLo2lBiz0ExSHeZ+aswsaERZuvDsd4be5qBM8q
33sQ9mehOLDaOrFXjsTtA0Pgll/hirmPe0Q+OJBk9KA0u6XQrodAyqgQsFdU
cilf5t7NRk4bX2gmfJyGll3Y0LSUn1cjmf/OLvmQPXpX0FEWJe2fIZqx9xjZ
lyV0BTvPfG/QFGNphnE6unOzXpa84s7H3NGLa3oPxG3HaU51d18tHb1JmuJo
PTOPCAgXwOg5MxrseT8PvuZ0jzv2QMJ61lqI+cdFXNaIgJvL1RSJv7Ye7YVB
fxdgC0gyHJb3/gGRTyAXJ58yL80o6z1ZcbqvgKL5IeKXrt7wfIWsl4mSRQ01
DISCd8aYmfvMlChduYDF4Sh6awgrenBmLtZiu0uB4GAp2XP0Skh24NoaujgD
JAu8uc8GR0chxFMEpZyx8OJyhs1yhCwbunittqksKTSgBc+itLU6F9GO0nQJ
xv7aIfpOwemadwQQEqDBIstW8uNsH46ea+rlYAc2GIGCrBgfQNIIrOcoVvPV
DgxlTBQeRk6HIEvnY/oae8AD0AdwT1kmvCU7GV/OHsvHeNs9fYQdlA8471dj
9vmiBWcFYD5LqR/KvJ2i+p98nRYunrRfXU3KW7iO61L+UL0Bqj9a7ZbChGpb
2nf8/UGlyQ9jP9mDFgsnNza8uvxt/M+RHMbMzNszFVEWEkZdu2av5/T27W0N
i4MXzkUWPpe2tY+OqZKeEtI+2KfPv2wibuB6lhMylxH5NqP+WAi1IpWs9a1V
Huyz9WJPCywgiWf4CADu42a65EApK0ex1aU1+p/vaRbhKtPgvB5Py72YLe50
xINMKkl+55vrxGnIAeu+/yJyNtjNPGB9HcPAg5hay3AD/YmpIqQaONDUpNZ9
iscA6qz9GD3PkIZ+8wfQy05g6aGMyGOIh9ifouk+fbblxFGS7ytVcpHocG3i
K0f4ZSaFvfWt8oW0mCsej81K9xbhI8Rs8hQov0CaOXfQ6Wg4bDIvxH/B8v7p
VEBK4hEjWhqTO/ofNYPpR8Bod2J96KSUISEKqgkPbVGR1Ceom/0umnwxGzJS
haeoTax15zJ/2R5iky+p3GTMk2uQl7ZH6AxPpdaDL7+j6pEvLSJnw7lZmVw9
1FzAYQvjj9cNM9w6ZNLuE8om6pMSbAskIvH/cDi9rSDTrKGR6E6lOChHdiQp
2342QwfWswwXNbYfiRKHH8IcMk2eJ5SR2aWEQ6HGeSi0TjTGu1vRF3+XqF59
BhnOlFx6O4ol/3nV2T49gW79i9Vg3eyitKkeRiDp3RoLxz6+grW97LW1cLXU
o9m7IvRaPsrt5u7O4eCguUrf1rFYdLJu0mD/4HWSTToLPwm6ZxKyP02t8rKE
T9JyULWhNcPDh2AtYtsqQAY2z4aoSaeAQZJXiHgrxh6AWmiv5jWkVVDgbqwR
4Mv54NFIHEJloT7dQ2Ksrds2jpe5IMlqoupj58Be/tuicN0MkrBVmwziavqA
4NwTDKVBOjR+Dzoo/oVsADCUBA3Orgo3vS3MFbytMxIwNHe7lN4QOj2qcdq1
gvC2601e2Asa9uL7UseIDoJcrAB9k9JG8fY6U2vOk3mIhuyk1P+XtLAtHZyw
my437zAedaWN8UHJlITrHq7iREGHCoWJixB4bHvjgFexRaY0IyYj7ZQQcdA9
1tfoVGLaIXhqnsWWuVjzoOCKEmO+FB23lt72FSWFn05025/+jE3lo4+JkuMq
78UhJtFiq98HOHQlMRj1b+NV7h99cErvjwT8RseNz4wKzfk035XStzOCRjAX
yyxuvL4YA7IcuD2TAwYMVktPBEoOyg9pz1YW+Xy3LgcRXO2b0L0tqBJJUu4W
gDJqJD4dl6h3HMjFdHjRF8vU061ZjW5cTQeB5fEVJN2wt4lmhmviT/+0tyzM
VbQCwsjIyk17iJ0Re1P+UzpfYlrx772sE1qMraFz03MsRcqm1P3cUQZprnXK
UkNEXYFIEJGM5ig3CFNdNVcIeaTF+k10scM+Qyoibp5k4nyUfZnUZGJxq2ah
pfht0jIpWOOjDqlQR3qZ9I2kUutaYdWZ+rNuUxQFsNNHFfYsxRxjftTeZPvp
8HVHKPZ6N9Ir2RpZ8hpnZ3Ei6cwaUsf0qseO2wMbCbRIjt7wCbLIioJL0fxz
SRiw4kQ5x0bd8mJSSECqXosSmzeSnjA+ULzDrdNT938jMHLwKOnRx6u3nPw3
7PcCDoB5CnB45eL7FLOgfx0JCUvs9afboy1RU1UDV0N09YsT+LdyZoYKBo9C
7F/0TCRfhtWvIPzmzuLiZz7zGUO42mSvKux1zK1SDNAkJVX/IbUdMYr7VoU2
rAy1SnoPSQJ7CN+nRI8ye659TTNaKltkWM+s7W1oiyWFyuIaqRHzt63wVxqD
Fu55BXp2gMoV+zpK4AoM6iJX+eiz1SAuApHCtcGzy7QIoMcBgcW7h2sBfHKq
K/vOURABSh6CepohD6/Z5R7yTtVvaZRC9GUA2C1daf0EIC9cmsSBXwjl4V9/
MQk0vUOUX4TEfJlgKi9/uPTEMKhkq38CTnavhkYDZy41cs9tOJ2oJjgzrZ3d
MFjGVWQUCWoV55jTPsP7TU/MWmu0BCu20Y0777bIxjb69TlYFjRy12rKwUri
KSSAiFSN0r6r+NweMWDr+8bU+aF6sAioUBWIyTI9PpHenBH2wiEwpvx1V22I
TIso3Ed9amfWKUwpEEEokd7yq4xO43MqHGzbIiFOhl0Hzkd5VKkBUXIPPPUy
RjJ+5kSBmQTZ0k02TNOrcMv1UF8j4tKK2lBBPFzwrfudhNp+XV1yPNHKbNO5
gHOUOzNDmuXgxO1sm/+cj7IABz2jBMb+8zyJ+uI5gOUrVpEDhJEAtbs33Un6
0L7TOUx3EpvbOtbxNfvObSoOkaLiESJYETOLWx60gTzClte5f/C256A4k2NT
hrXpaRj9N07e+ynzWCqzlKtKWPJBEV9kf4t+LhTpFNYhQ5vAgp9hPYdGFM8W
H7Zuu7EOhZOPsmt/F0gcqHPg1ehqOqSYJm7CsOJRvtuYC+pxO41RbNWSQnxb
Z0zKWaNIWbncNbbDDZhvNLVar9nUTlP623j1hDrV6Coj7KW/q3D/KeSYJtVW
39Xh8CmZqGhO0FXkDl6J0r9QpezzN4xLVbEEHdRsTTGxgNZP4QGKNgveMp8s
3yey/6Lq1iMrZ3wviZ/+18308pUbh9ZbugqDcu1tKGK0Z+0yl0Fj+FORHlhP
D2WGSqWze2BMxyJacImaGqE4csf+4nSIhpI5kHHH5jSwpTR6B5037k9Z2P1+
W7qyQhdYVsIQB1O0hiHDgDnvMK6LckOdS3sXmSQaY1eSWbsMwKRK+Zch0eQW
DjzNuqV+8+WbJ76KRxjJ1Hmith3HfreATiryUBd0xbjHNeUxuOnMfUDsbt44
Avdr05IcDCNR3HQ7TXVyNJAjJx/MFiop/PCOahquH2vpNBWeddyyh722fT/X
QOlaVLuaDa9pXnOxfUsWuvCvP3QnhBr3sX8T2oE7USCP/V5sVI0A5z1j0vlt
q41v7KELUxvadebuY6jm8Vvw7Iv9/0kKBKi5q67oot+3LFhy2CMAMz3NfvCN
USyujp71HnQXi+3OkZX0VcrC5+8IndTr28v3QwIv4Q1uQMvJIpoFLT2Vip2J
7TAb0Vpfwx2+WfjZSMNHe8MNtsOHvBoJWRNww6xlQM47x211HRNdL6uvQrXw
EulpfcefudGYuwUOJYfLS2DNax+/M5wtbPH0vy1gO8NRFpXdqf6oTaVHH8IC
ex/qKdWBuEWr7K++B5PnqVmukE+ueSwP/DYBV5Pmsal6FNwz4N0jr7aMcDQ9
0FsqFE4UEcYArkeLNgDpRDnM8Zpthtoya+ctNywJ2xngdzIAcMqSj6HQjJ+l
ld5Dhcr/fAwcNGcr+39bepqs0pOOHSTf0qxBj7zfIOoS2yj4n0bO1O2/b4Fn
8JEdI5bDisgTzhoRBJQdESoGIGEnY5/7ucbvkzB0OvRw225OI/cZy1y5fwjz
KIoU4oWnXsflnxDDhUgD3JgDaBFraovhd3MNpvqr1++ffBUauBCWXPS4nCWW
MqsHFZIP57kg9iku1Ewyr3ag+ScpEMrohxuTEcRFOOjp342fx/S/6HhlRC5B
/ia/n/Zf7FzQgVpbzqgQVd19tsUIxM7lCsnUO9CgNdtLMOEvlm0HvlnTZIfm
zAJRVqT4Ml2I7VUfPK+s4/+7in//Ck0OUyjcA6lTcHz7L88OQsIWOq9hq2g6
JtHhrzIyqwSUqAObFzTPDrptOCG7TGuXoHGC5BzkQje/dB7loS1r5DDPXg1z
zInAsHp4eQkuSnfeWNje2GiycZCrc6EKBvFp44blduO09wTz/MbG2iYi/Jp0
1XVX5qMD1ucvIKVdfPbw/iqe1C6zX8ea1SP6slXAS1/EeBnWiqzOCAaGnEAq
bD5vo+ZqSL2Hr49jAOAg0cf/ZFQxMBmEVmhtUDXeOnMDcRuEfrimZ7wf52+n
lO8b6PUvtXWku6m5etTHKFW9KwZ3Mb5TDlWmwMrE4fkSAYsLKIvKA3wiJEtd
dBsYb5EVnILOXTlmJDFKM/mOV3sMlJVEqHOeYmClBuqmFn5uSyJR90i18jZG
fwJTmRUf7AgbGj6DFhUg0yzusACljlg+J9taBI77MOZj3yca2VUB7ZCnERoo
ngnekbfy4wCAG+DmHJo/5vQuMHRupso2sEJKSje35+UUvRr5XKkhAZnFR88o
LGexY08xAAEHZzUkKWp1a2i9tXLeH8qowUkr5JndDbq45tHJ0JMjXdWx2hPm
DB6DpIP0dqx8JjF7OMjuUUp8mSWUjWphpWm25MJjaCkE5r4bl/yuo08eQNLL
T77pR97UFSpyU5ZJwJja0r95ebyVeUIwqIdWRLZQ2bLgbmhkwNyN1wl7TQ+s
d3v3cGAS+U6gZ5B4AjKxCIH+dST+Yk1gyJscF5Gb9amLjksn6Aokb8nFr/oo
shmsRNI9J00QNP1X9j79J+uctIsyrJFisA/e26sYrO/FrJh41FrU12d6sk+D
2iluIdrFXo5TqOCksG4q9xrXwk3EGGtt0/1vd0+hfxMQj1PnI4+xw/tlgYMH
mtu+Js7JVStxhlNaaEd9MwbUnLK0BcAyAfDMb6K+t66jpkrqa4sjEmBou0l7
pbuSm8e7WrZVVUAKbOSAp89gaHyYnLSzbl5zcWZJ0otVSxenfZh2tfFbqgcg
X2hZxPAytkOeSPNVsqmnxvpzh4Cj/RyGmyB+MZZt68CRXo3A81kTBw6gJ0mP
3Y48C1G4rQbXlpLsLBzji68PW6Vg26F0nrbPsGdVTJNnumT9VxSTAYeJG9ZV
WwfSTqfFjEkreu0wyYWfM7AW+y/IRr3XrCbLM54lvZ0x9yjxJdIrQi6u6Zv8
ZUkUF1TfdiOZer+08GHaGFuirKHuTsObUToM8zCt3n+/KSyq8X3zDWCyL1Or
Ze4kGdutOsSsRCF5k+EOiEtOq4ckLBQl8Lvi1zBNAn+55lPU8uclA+BJSigv
bVu6yZGPZot2GhM/CnNrqHF89RpdFLaLvMzGUMkiPmonfWzDNwHcLNcyrZRI
1yTc4kL0RSag//UsrKH61kJcFsfYP7ZSKbb3St6ULpwB1s1ICTxhl5OIslDJ
WQEkgwDNim6ss/2YVdwLUkxMaDXwByLKrEK6ksurW8eauYhybo3FIda2TnKm
tTE8jaC0Th4dV9kE4erl/DQpGUGTHPBEyv8lEhktG9wOc++3cduLDOEmpg83
CWkpQGqGsSRHAPc6nM8wPCCG1CF8DvHR+mo9XswwmHDnOhwTbAGXy1+tH/H/
keQZLIDC9v3Vobtcfgiwz1mQhawzaKE3uTkMO9K9od+w5FDXYBzNjqY+3jDZ
mFQk8G32XTIqYYDAAvkWu/64CvEcY4awKG0E19VooyDLjryuuq9sf5KXWUNy
LaM9rEXB397EMkqAfxnWkpiKL9C8bGwjE9yyQxurti+Ro25HodLqdXVxWN7O
lzIgP/SvvQSRP5mGjSEW1tvN5ChO+YrdnN2urHtN8bX6RbeAaqLphNxVVopk
DC8u8bbFMPLV3qnYms7Sf+cKp5AyWNUeqTAZX+bB22rSvQ2jMrAIyQKPPZ7v
EMuOlQZkJxUoHKB5+LW9jTwqbW8JbdAIFQtpLvh7EhXnT8/B6wFr2pac4f1s
WVDSrq/wzRcGrKryrkTR9pEpejKzSjfmhkleMrDNaCj85EfVBGtFL0UNmYMs
yqFGVjTm2GFRwhsVAg8kQqEG7yXwyFMwiYG2Gu0tw/P7ap0LmfzSXZ5u+eVy
VKJgPJ8v7LVKNaZZDIHuNW45PIbWkk28oYuhVvQnyJzIW+aqtxvsihXyOgnR
hR9iQPH3G/2A/0FruMlpUZF12ZAEcjeLGTFIhqq0ekuhGEED/ZryrQU5V44L
gGviWbWGXaNxClbbkv3dZ5A6LEFVEO612KDLOy8+Z/hZVbE0oeNk/x7Hniqu
9cg/AVFJI5xn2aFQ1cY9HM822hU9/Ty53wN8QOe1xGJCMcb0vlnDm32IP/mn
PhLEh2IpCx7GDEHKATvKaU5oQDQALdvMwr0egTmEs42FqF2xAhNmEaf3q3M6
/ddxftxUCZzQBdBspKVpn+eCBN2o7h7n3lraUQyXQgWaoSRAvXbKypbUjlJU
ZtgrWOox2Svfh0Xj6LFtW8hsyvKrNEMD7jCmmf55VL+tEXt6AWMrJAOEmBYu
c8mKRTomv8jjCfxXs3Vs6rh3fOrCtxa0nu4XPdqZZHJTvxcL/3V8FL1oXkls
oNjQhbbLNrZy5ZIgWnGQ9SRuaY9KwsMxQV6h67zfe13AW7Kw8RS61oME02qr
GoMTndM1Dc11q/Uts/sktd0vccHlQ2fuC7Q8SCzfFR3zoPmAoexZtlI/lLx7
qEH+jPOvG44iHSCVxc6gzpi/RFUkrgwbQO3YwLar+DmEcqGb4UPb3cSoc8Gy
jh8uyRlikJu4FqjOAT3u0ag0f5n1p8G9XhGgNsaP8F4Ms0L1mnws9TGeLTTb
j0/vASNAis8xGfFzHb1iV3lij7Ng/nZrQQUm135PwyU4tIQluM8yOBKpjf54
izxivQpqDluhnV24y6/VSCZ7kDCsgGVA9OJ20Wv/mVucbX37bRCzVUY9mYGT
V5yZzgcAluMAzDGkA9pXzq6zS4RsqQefo2MztiYxERBXAUM6Py+9reF5vjDO
kCIbxLHThv6B/gWbZzDHOVGrVMZPzjE+ykfShpE6/KyBWsL/S10sIZ2m0SGO
CZdzoB9hQCIspt3wyjnfZzvnGrSydFcrA3Hh9ZfZUsTcbo39v4b8MB9ulTxT
DyT/UbtwO1nJ6JOFvvZ6LWpU+WrOipT5gJOdycvIe+PzhIHJEakgdd8igOkj
NEtTEmrCCp0CgmHi544lLM0fYKyExJNDWbepukn4YoUPVeJzao6LRWqaCQUR
wOGoecER57R/MYLuxVrsfHRFVit0T7FXJeH0L7qGRqIREIywdvKh5hqpeeTh
Mb+eB/JLryvWJX0HFQgroAbOMfIcJYWwAddpv843XGH3wtGd9k8yZScuJNhy
rnttM80ADjmxwX/0VCIQzSb4Axgk0zJmu5UBeMyfCZprDd4nucvoWLp+rsZX
v/ZVhpC+IVg9OvZddxd2PeInPOgRYyLqlR3rNuU3SCbMQs1NW00hNxAUo+YD
aeBVqmYQy75JXBad4fKSjJc6xPqTCkcKGXUQlv2Qx1AsceU7qBYjeVHbxvGf
erRzHQ6ZQRE/vCHVy7CGpCsJVwvgQcyLMVc7u8c6oINmcIcXpY7kTXppDkR7
zdIEDGR35UqmREljPTQFY3bnxIYyKKDgZestz+K9cELO+kt6SsWeOI0JQMpe
y0ZqIMN1LlIgQi62BcfCuNFYawhDY35I54Yz48nUtZ68gYvk7x51nPhW/u8B
nyPRj+IxEkibfVQXCRtwUbHXE/JMX+oVlKW2dxy19Tjm5T4ZuMo0om6hlF8z
l5aekOPZHmX1lvulKmkiwyIKJCKZuzysle5AZXBjKXYcxw9ddBA1C/wBoGPj
8RetFkwBH6ZnvlCJbdOtlGGM6h+M6L0vUrRSo3gZn9k0qyhy5MIOE3olQ8XD
GkZPLyGPqQJM+yjyRMKMnQbdnAYQ3FB5erRvbIDIoTPsK9gpusZjxpxMKhrW
RJBkyVhNCnEqoZO+JmNuHieKfitFXVqk3l7tARq5mYHU6oWIMjH80gQL9ca7
P9ReD2aeVWSUc7QCoFhst9MxGU19RLmssD2FJfA09mhyidOCo9FQ5CI3fr0Y
bHQVn6JkS5iLfTW2sbGiVrVEWaPQBR0rp9Z5p5bwqckSFCW54kURrZr2z87s
O8CQodMClp+Z865SmxmeKs+pwNENsBmOOWFRGAvGOMtw9INve9RGGYvyLmAn
4wzwec/34j9OujugPspLZlBXDWEdK0I6YZogim1LlMXUdLRPFQvcPpG3Tdfx
MzoqMTQKjmWzY7djq/GGH5af9KbRbii2Eve2b2qliuUyQAiPUNOWlsholrnc
+ijK4D8Zvbgo9e7beQGnSfUMAoCgpnAQAIRpu0a1j23t2Sh8BZV+2DXV0Zkx
zOTPEDLXu9Soy82u+29C3SfCac8O4iTs2/A9dVk9IOym7wdGlh+M8pOSupAc
XYdjMWv1qCuh+4cGMPfEB1WrhDaSo4enGX5dxMd6G3rRDyr/f/cGrNLMJfIS
8ZBju9VD7sLDg4AT7y/6zQVsaLw2QoHKqNgbD7i7uE11dz8VutW27+c79V1u
KfC0FEHEUHEyLQMabDtXjszbgVljfHMfYNHn0smqQkPqAES0eFP1A/JrMsZu
pe3k26wnBpe93TOZnzpfD0X50Kr0AAy4z3ZzKstCrQMD7YNLHzuqt3uECd0D
UgZ5dm2E5R1BoSKUG8D2IAGksoMRR4mIIl6SoQCkXFJDGMVLeNIQ2ZHXrtuV
kmIH/RXX8pQFNuluvi3RmV3Nayngf1C4cRtolkFB2jW1uNbHUPhkPJIPaevr
2nj7p2+dPCQVNprdCzr+RTMVL2FSRO9wHIce3R6FCXHdfYebaSNjTrKyvbDW
rj7Wor0eQ5/QPrwlXS6vKclV78C7/u5+ctwNqsEdnwSiiNigHNeRuI27wkuB
cbzppvaBOms9Tk+Yoypuw/g3k+MacN+Dvd3zvQb2CWMAvW/TcakLNEDJFeLs
xspRX0kssUVLAaDt2b0joSQj8pJEhJSEfZTrVT2l/Vs7+KZtno6SGsgFWMnJ
PJAZzTXU6wdVYXg8EB/YeLBMv1wF05QJZRdfkLORXcvoaDvfh1FZSvv3+eci
88xkJPJgzQXedVoodtrCPZ3aMTKTOvpUR/Jm173rtSNFJDxj2OrmdMAD3hN/
oKH4qD2woSmNJB8P+lgQmu6wl08FB4WApsTjadOHkCulbRln5+H2vqGMm++7
4t0XnmvqmLnujbsOOUGKvug6HXPKWflp7nnOKBQikLPYtZGd1ijkBsJcWNMi
A+4sXyGvFrZFsJs7x2XboS+8qAy+ggVWqfSRwYcvKQBKEF7JvzhrxxtPDlpO
Fac1EUph5NQwX4htxn4uHdUsX5y7oXM0yhwOEX3emtcp927eUEnO7epdY6ns
tsdu7vsHriPhd6L4O1oZsa0neknv63mB5OsSvCrOHBgjRaCypz9OAV81NnTk
XC9q4kJ3rehhkRdS6sEc84fDtIsVQVQkmbEgMfjps7H1sAE9W4EQ8un4Zsxz
VcrTPOUhZdvAP0TaPE/C0KKxiMtXFQDAZ9T4Pivm2kR2r6QdcxYfImXBNq99
TIXrTPTLGwtJ+spaldsWM0aLcnhb3SaXhctatZGOI30VnYv0EoDcrZ04bSNl
56YeXcZg9GbXv9+Orx+AzRdjG4fbV6SQVzlk27bDWqwbINBfnUIn+dihsNKm
zL+2V7y/sagwzBpEwguiDCho2DzVxmFmOvJJ2UunnlZS2qs2wogvafx+WyKt
/uM0ck5F+W/DCMhsZUTCrIDUZMdA1TBECETczjvLok8S9B//Wybw4fvyzRQ4
jpXXCIqMKnKIjbrk1A2HDY5UC3mGCnSH9lxUuUC6dTU+JjswqBz2sL1RbDr0
q6qOBAFAmrOwwXiOOJK3PLX9GkuPa6Gq9wR26HbonB6ajqLeI9u6gYJXozi3
OmFCwkvRoEsXyjoYGwB4KdDAHUQjUrNKl9IwfFk+brIOn4KkymARNV+En3pE
iOwlpkSv4uVb6SgD/AhJpozA4MNVprO1BFKk6wMieRPQAgeDU+ho0vMLZX29
uduC4btRocG9Gpad9yDgzIaCItvf4Bulh0uk6AeqkvrYvvKu1QmxdIFfDcSY
fwk0hJrAnCSsCSlQD5mrwLtTakJqj8hTBq0pI6Oxi8mTCSclByvjvQkD+FNv
ISyLRjCMpFtaYAv2r5OYgnzKkrxHB/NlAFoUPZDYKeJtiDj++VuuVOVAv8EE
ut6v1Dex0V4pKbt4Uw1iVDAN4xZHxf8f2h/y216YHf0Msb4i68qAKeq5VwXT
7RmtcOfwI99e5ZB3xZgjr2QttqdLan+Li+7shxGGbmHE6Ys75q589Dcb9fQh
QJAAAT4kQ+I5bIbDlXAWz4X6lGrs19LSDZadP+fedAGMzVyCxauPRbVLangI
42mE7oz/AIpKu9WmUXc5CGwh4opfFRAdi+XQNqkmHow4iwM4GNUwxYlCSAMc
m6qmKMnOafD1GQiT8vo1c21ANNh0ROXxZ5d+gX5aSqzH7cT/3giqPUB8FnrF
LFHvB7Dkki1vq1C2zXJ2OuPxVusppZgOHTbwaHlhdRfCvpCs0A2iwghEQ996
YO5Igrl5aSE/PkjwlTP3icO7YqDnc5MhF+/r2V76Fn6jmFKzpflWVrWUY73J
8MCuCi0cJS8SYubwZ5czLM1DHgiiTNQdUAh3ty5CIsnfgq0RPDClqO9Mec8b
MJEW2ghs+vWKPrb9btpm3m0v8N7iRFz44BivbPsVUkySl/f0X7Hla/q//POU
bI3gOmRmMeKitxYSweQUFibxNmTfxF3TvA5R+zA65XrRuhk+HOEHbQs1m+mf
aRTm3Obom5258JSFidVI+N5slpJSM3X1vt3TYw6SXcafp3Cbq8mRahQB7LC8
swVYk5j2Zu/eYaC1bAq69taqLBqt6AHlCvRHFdwWh4q10Wy9ItTDVJ2eSl2/
m8rlKaS7BdxDEQZWg/k2WAJBZP6VlTJ9LxXuk/H5NJiAFcU1RvqvxUr0s8XK
W9FLJnIo+UU2sZ4co2ShMb3oRygyry1U7LwwUkmyIvpPecGprXS9dhx4CITF
8tGHevFZtjqp5pQofO4zY/U9/Q6MPh9YhjVdplB6d70YseMsCK5nGDb7pf9h
GyrC7V6FoxTSZ8kNR+cSmnN0dN1A4UQRH6PnkIU3iLkBFQecXzTUZUEBGmav
8XB0ghKtZRXNhgbOCIwtMaDrPMYeWYkWlOKvakqbeWltgWegFZKN/0DQ+QXq
RaGQZcBwbudkWw5O2mIwCKgZTwEEY9mHNqa0UvusIPyQ51fz6gessgkES4gi
mX5mP6AgVbo5TjIdP3l/0ek8CG+YCofIpfrX7owyzm7WN8eerhxBpA6qfeP7
jX3BpJZtL1qvAm3LBB3Hnta1twr4FEjJoDo9KdZUEdoj186Ga9unNA9orcDA
6u+FU36pKAS1tz9tWE43STgtZwIuBM2hLCbkFUPqPHUJHR181b57T6ETicAC
+nMAEDRwop3AqV0YEEsbXBip+c/S2cOVtd71G+yITOFNNkrjwdU3YUqqlKmv
+VYGRT0srr498/3P2M7UIX9QHDC4kSD7dhB8GGa70tg2HFetFP8u+VshkIYR
giQ1H+2BNoaMPqrAlaCsVbML2TtHYxluk880p9wcfW0ypTI1qNrvgDliGp3n
8vBSDH4uKXerdrYc/ynevOdK13Pe9wd0lLAv7KCrMkQp/MGQIz69yWpWZ+LK
QSkWVq9oTOtKahf4cYqZelXyBJ2f161U0woZi1JJ/j+DAOc5zPRRmDe15Zt6
rS0tZFTBuhH2ApYzgALH6iIoiljL77I8umSxonihs2YUTrvyXjAuJlo7ocBw
jr5YVJ4ztpXafSRXTl/aea8kmzJY9EKD01Ad3DMr+zyWC9vQ+dltr3hS8dqb
6FEOkSOrUbmu/JwH9QP+TLBE69hRNtKxet0/Nk3Ux7Ed68V3fCfT7nSElRNw
onZEb3TCUn5Hdz/1KkFfUE+JGtYsv7B9m+lYRAY0H8U76WLuyZTpiZx5p9bw
vDTpkxDMtSRZfJ9fMU9gcZhXUtRU5dVILi1lHxF4iA/PMdNj2wRKZKQfolcg
dY5xwJ5MxJgVjbVY63kuNWOnUF1Y3loXE12ZBx/Y93/B0avxZfDMRBZqMjMb
oL4OVElylJEfMlU25Ef7StoUBqC6G1VaWnrTtwo6TnBmlcxBgc4ksRqyNhhk
mosYqz/MRiWUThvQmR1wDnobpEY6D3iaou83JaqyMW8+w3u7vR+RKz35hCt6
FwYXFeoQh24G6Dte1x2AipawX5VhztPobqU7alDzB0ZE+iHtIAzdeThd0IC6
EapX6CjrbtfCNgEhGqvgnMjNNEMA3vtPtcQBzdrQKUxVBFxueRz3ZVBxrHKf
uvv+vROMEh/O1qXnEsndScZP6OvekGIdZFLQ/799uHOSkDrDlq+ikxP3B1Nj
2PMRpdO42dS/bOa8BNeCnKOrt4a3IOi45c4cvqsf9seCMpLueSi2VD9PL2sO
FV2nB9j7xlmwOXICVqZHBc5nWXDhmR7g/mVIw+gM/Dw0Vtrdgl+OIX0iVkgN
o2MWvv0VZPr9UyXqqTI5OafLW3Dcledh9WAzkw2sOnvrbTlgdpn0yyPZzMKP
bACKQdM7VVSTfAzr0dNJidSdhrh5GypYn/B+qhbX5TdJQp63T/2kWvYffJjV
6OMeUdZQruV/Y4hnlwqf0NB/ArwIYPPBOViE4a4mFXQsiXcXZlMgayNfYu8n
vkxd/wsxiKYOOhSbcUB7qpiJQi63NKTV/3VsNQ5gcA0kpzstEbPEqsU+BDen
wEDLt7UbZGYLbTnYElEbu3PZuTz5U08z35VbNTBzxFlCfxQuImdK3XVXGzzH
B1SyNykteoAhxm4OY8NoDD0BY9z8sgen2SqRCurXi0gcZKmF5hz/olDqEkfD
fs/+k9Q+0TlcfdV0abT2KUHVBT2kH9/bt3uy/tGyjGd9vI9Z15ckXzBnDLQC
U8stnR4zLO1XrqAGsewF4HeH5uNw6eZqPHiipIL8uu3FZoodTIS7qnkSruK1
ejN6XBDzmyW3oED4UUQY2CmedXAFdjGV3WBVirBvjWgapTGPtX3qe5alIMl4
J6j9gwKq4W7Mmuo2Dqctpik111gjL2WQxvy4TM6Oyh8qgKMvLffb00+v4arP
9gQcfiyN9oxCkN0P5EJGc/WT1yaRAC1IhxbiHvoJgmWi5ivFyaQgnSody5LU
CG6mqBDeKI6n2VzHAdMrLmfNtXxfjBM3Ydj7RVA4kt45tLWjUPYrav9+ksts
r/S7qYJB5Oyth7LsaympjxjAGtoL4rfC+gwESNIoWBfBz7uboVpepstgSt/n
6r3lDmBTOnN0KmcG45bQEDIx0VC5sQLb5QF+LklyglW9f62Sa2gJ9Oy9dZgh
aAB4XNr5XYkNJA8nGEnJpxDbEbSzrnYK1Ai1TJ3Y2hvxauwyP4nLwiC0eI9S
kX1FoRJIzdzHuLAzXl9QdZPhxpOz8oRHmi2KBBclMKPvffpaqPl8QFyz1Oyn
wGMq5EkV+pMUDgbAmsubghzBNfHDDcYddYWAIdHiQwLdkygDkDE8U/ShVhsY
L61vAfwwX6lYptNC13e5eQA2zX5EJH6ZdO5iQbVAEg2oK+shK9HSiOvFqF00
mmxH9YvHpoGlWpVqC4Fch/idfpJ98oP3GMAikincMLthTno96hsMMiWOoRu+
eWpxuV0h3TLxYd6ZknU4lWTqf6DY0HNFMvDUDZ9MI+p+JtaTox7U/swipshT
fhbPrmoe8XVQyegStdg8isaackAWVjm7YXNjzsOQAN6lK4zntVI2Dp6efyVK
pWKbrs99D4WyCd0HkqYwZI4H0bns2VvwB+Xa2MbY2PvCZaTyrjFbrvpCF8Dz
gnS2m4OYIDvgmJHsxmNfbPEbxLSDdVZPacKJr3H2nnRY/7ZmGSPgt0FfQCFe
8PJxEuMgixWvO1kuiffIssVLMVfdGNOgwWp1e82BNwu/9qNjtvWqsySzTacw
EwDJ4Blhb6iE3oXUOzvFU9l7w1GE9CEdaflKbP2/y7RdfML27bluWS33F6qh
ILuFBkf+XUvE+B6xlT8B9wbztaL6H6tSxfV0RUust9qe++VjJA7DPTNjMx1X
aABYTlAzKY9CCpF9mCfJpE5CXqz1cj52BUeehI1v07d1o7ZMg05EmZaQmfPw
mNf+8usodWR4fT9TYKaQPTLYv/AScMRW/vZewdH3GRJXU4Q3A6NoIAm85jSe
6YhjCMu5qg7K/yOIoHX3Q9EYFbWGiEz7/ZWvr7k+tHgVi+Z/++A3/AdwZwdN
gmjMTD1NlEDzpprUcsRcKOUzyiC1CRo+IfutDg7q0bUf6noEBQ8Hsy4/Zg3J
cGOdfEAjBJStAuDffq4199WvYs8nyvOWJId9g1Bm1QWH6Fw1TnUYCVLywsht
IdurtTvQxEgX9FmXtKc4YAQXZpwrz77FbXIBiN3mkbp8rsxFUauSnvD4PVQw
tlcS2Kssjfxt2LA/YSgey2Jtgm3fEE2hbPd+iUID+4KaN+xNUcSy5uZNNJBz
pI8dqW2lKJJXrHt+8yXkKgk67Ei+JVmkXt/lQnVHT9uXxURQs1DrEncb/wo6
sH4y/kvCNgNFwxSRfl+Y3WDLNos/I8Y0vgBj5gDF0lmpb/clkFShrY1ihpr/
/2gV69n8ZlO2zWZJOcUrQ/tNSqbv16M0dpLjrGKBM/DZqwhFtylTq8jQZUOu
yILS3Z+oeWCRySyE6oaI4Ltw7UVNCHuK24QzFCidABYCg4sa2++4YQZzRBAP
c63+zyaFtGLAVM0X8seDEFYomU6nZ7v0GIPloZrAET18IN90lH+aZOYih9cj
m/mDrLfw4GwdOfOpU0zTv/iYwQ7KdMfbEQ8I+gnbodRusGfFvbvGNIJxL8Ci
0M1VoEARxmZ9CUa1AjBFLl55XOGTNThFHIwt4f+tOHLE0fmb9RY6K57D/zqa
OTN9r6L18PLdQY+7dGCuvYiLNF/DKX122rehsMQAGH04kZ1zPRQcW+oAYJLz
RuFmeS+ANlryCSFKoLB0fmCQWu9DpDU6hdxhlYNRcnj6KmBy7FQsqmRU1SQT
tM1uvX/FQDvyDqhdUT10gR5HEYlvG2LgQUyqRd3sNptTqfcLrQFHf54KiU2g
U1SPWvwqPpIKV9UnWxeMRzyU763CzI5tfg8vteJgEMNZRDPg5ibI6pnCXokk
VC4xZ4VlszR0DDo2QkNeZg4q4Q9SBK/PvkNpT0In2rOJGsX61QztTze/55L1
V2oWxCOAE/NrCREXTzUjLDdi69954IYmAeldpVx8s4dFbqhE2/vjr3OIGssZ
ryDPjyIiTRZ6j5n56qYUThgTPjLtLccwzdMOw16SSxj11iKVtmj+oS+70fCs
m3wQ2m1UldumRDxnBI1EyMNVpu9qcd3mj74yhf3fPMJwvf/l+yeFEm0znw7F
TbexLWt6qqDBTUOcdGKgSMinpRltoRtwMeg9MUtAbdqLxEJpndG1Q1+E3ks5
RY88iBtGKxMPstb6B3HRTywZCMzZy/zcqJLQgspun0H3rV4rpoWrsLcHNvLH
EABdW8CkghssDCHoCjr2me44QD0zZCDRhLoe1DMy97YCONq9q9YMvblYjB6/
8Xjxu94Gj/DUds4/lVXlUfY89e18KrWcm6KwF6VJszukmCBotgcCqCMLswRC
ASD0yMttXyXMeD038+39UGIynFvC55qsWXGjgT7i77zV3FsAV+/cfUr7pMlP
YUpS5Takhw20dVZFyyharofG9Eu2/kMjx5MGJmIkHiRM7oIit38O80ixEiPv
E1ygcMEDzdrBQ5A7JitfWcbwqTHV4o3/AbCAGVExKfoYV/MEJ9QnNup8bqWL
KJ9MU/B0vNAHEwSkntcNTWPwbIIaLXpWlIdHrDvCbGnSbquaRVyRjqj1I0li
kuvlDI9HA6MCgmAmdMrYGZu55LVOEqw1qcAWxwjdcCr0Po/83/iZLfiG8zn4
lKjH1/mBY+uBnNf8qFpBKfq5uA1oC40O2m5nHaKhhBL41GMtSK4tUAABIwmn
BFVpFTNq/8b3gIliIwDJEDCFm7yOcIxKfxWSm6BufCdojLhu2CmJMlRxWzuf
6bEIkp5GEa5LvvDG2MVoi6RtAILsgqXQH+geimJit+I3wC/KMu++TMEMaHks
LoV7QVkXOk7icUMT2ysSI4PXLBlQf/cGlfgH3uK3pXJQSemeeFCnunYidbXC
ub9WMzhc9csi9Vi7IP5Z80165AWaTBqnOi063jW18rJA39mf1jpjUiOoyZpc
xH0YhXhYaV1xiFUDpJF5nmhQKsRpRQ4hmk+31zvAWFt/nTxz1YOfJVU3ZLNz
2eOHEIUev1drxdHI4CX97Riqj+07yvQzFfKKjGt2gsLv0eLQ+eb1dSsYoi4D
OF1yIKmZa5qeX9rGshQ8exkwX/RvWqQgn9mSEW07FzA7QBSmJweC1arFpo1U
7SaBU2tMi8ODuQ24nKMDkFyyOp4NnfGTTE2u8wKDlsf6VYT0H3JydEYAqHI5
cR8Mx9oQ9LgIKQWjC6SecW0p5HkoWmOR/D+u+RLIA6QAAfB8KHCuE3G5nAUe
iE5enSP1+hKIl9G2Q9fAlPpsYSryvmlTdMEAfzdPGWxs5RIHyVdvtH4fpZpN
Lzun3U2NDEheooBI646OFi5PhLWVAjphvTl+CHpU9yDnRgt13la0SDr8wC9E
PC4ry1FPUy+leE+k+DZWgqtG7eRqOiDM4MQeEF3lAjPHMDwawmIB+vTTW6Bo
4rG+ELierMXVNJfAC9lhcofE7EbHuY4aKdYWdlUnjK15b0NTxIFpOC5CgUHP
FYNKbKMHx2uKzzQ8xA1dgT/gRA5qaF37f8YFRyROxi9CCa6kN3eC5HQUFzXz
q10bndcGK8eILSsRQFbRSYcf2IuQ70xZXaS84EWxpH/ue3UVYGH8byWjI7+q
MLl9oR01bfPGzAYIhru5GG6yNQNvb0bE+ilrCmeed9Wisoc9lX9E888E/pQI
zncEeA2J/sSccSzsBbBN/b0xdLhpp84JhTNCUtNctQ+lvCHzUYGT/Xa5LwqF
K3yJ0YF/nM5x79CnkccNhSbYWyL09x4dNQTOwptO2lZiTMGnO3hrzTw+ObCY
6Fa3xfKWlxFVlwV+OvDQ/n2wBX+PsAVBIAYNzmNxHBNy3xFNplTdJYY/y/c2
+a3xWFcrme0vXAOsoSU9tTFlX+22keh16e8/GiIzJzoly3FH+0OD/xKAQQQv
ubUTfqgWJh7CUij+vHoQClVY77YYwzkNvcWiRnwSXBLHOuUXWbvTrrQN4NFk
+AZQ/xzDsbqrCr/e0GdjswIAJ7AIAATKDFMQSEEzqwt6zn+WvZwb9teJOPmO
tAMMGDe4KnkFpdsbr9t7T01c8XOkCRKXDhiND3xXyPhyp1qb+12N6+q8rJdh
1ANEMI7UjPCARlHFzIuGK8f8I3jygnZed96z4ajuKlkskF1vfnNz5zPU7S7L
VuW/5o2d/rUJfMziGfiQqKarkjWTJvXHIPKbeY/qY1QHV8YD+uuG2MBEGR4U
fpvb2BM8OmGyL28Gx3oIfVEThtS6O/KxRfCjQOGDk2Qe4irXYnDXHmKF61J8
IDilIPTqc0AD5/8yyg6q3lr3OKbc/KGi7MFhzxA7+b1EHBInyvY7hsC0W8UY
A47nMONRCJHTX3Z+vhYqavhJcmkihCglUcB+MCPL1agk1n0CPMG2/9vzOaac
wOEd06qKbYraKt1DDwIg+kDX2pa30DcrYcKyZb+HJXZgEpV6XyhxgAO72xgZ
0ZlLMYhrM+Bdy+IBJYsRh4+ds4Fw9Shsz1lAkvoy5xvx4cgXCRhYgzxhCE0D
l5nG7S7dT0rSrvFQFHoavA/wS5WNkctuYIRUAFeJmPwW6cnI8eiVs2I7Uenc
CLwABJd1ArtqXJ7ehpmKxBmgkAlR/nBXTyd4NndUeRC7LwfJWCEX0W/mO+7j
Q+M5XWoQEdC+5ALftSFnroz5E1J2uYCH+IAYpTkoiU9d0SfuaFg0Gsj3f2Dp
dtzq1bPa9hQk2JZ/BJovd2RgMfGBQLrwr1K8m8SEeJDkm8Mgc3Qnp3mqKpyl
38swpTVVGGNNJTJW1IsOWZVsI1T7pQecRCZoaBOZNqZ/qKe7IzK7rFpD/o+v
DZv89iRg45KDiD5yILo95aQU+ddholilJH/k8X17LRnmfKQZMfDZ0EWLvkrl
GWAYIDQZAIl3Qu2G+FlY/hLe5C/jJ0tzFXDHv/Tl5YH5pLsNAE9ijuSSUd+r
BaV9HPJq2o8xOnyC6GN4Bw9CzhtF6zB0CQB8Fr9O3e2Vq4NJqLDuLhY0iP7W
nNXyx00hp307YN+6/P5mqPsowEHUH4iDsN3qHDmz0h745UitM9tTGn00F/vn
OwpLYS2vFfHCkd3SavXDsz/bVjXs+ojWUWWis89q8RG6iJnIuqC+BARGPkU2
oifeqPPSs0wf1LTQS8Covv42iucxlWBR+5hhLg1fQRetlz19+4tsocfmm0je
+Ti2OMXYB+Ty16PBwYXOpnYBYXfM34Ba6hSWcjPG5eTenogZfHytvzP1So7u
3hH9hXdDRqGWfjhbYlfu0ioDOw3ulZNgXT7ReL4ndNF5lMDoYgTBLA6qACh2
mXGs/y6K1+ksVgpTom26kgUKrk1936SmT8VRLqMLX63Khff1i7rKdCba745F
k5Q/e+d9nKM+jRM1GF0SHRJqG/e9/FDhoBnYvlZFmcDS39VaF9UV0mODOk32
5UMa3mCZTNOD3XYN02gKLQwqtqIIdQRPE/5k7zg9lO8mlasMCAGrWQp+BJr8
2hvhXdXm7mks73nGuf35YnyL2I78iu+23RYfjM/SS56GJAHiHOhuygY5m187
5Os7tGdncqfckxRFM2M2sR6ykIloXUHAMehSvO5MjkOpyXxhIiXM6dLVSBj+
FpUzwOY6XLf4lo5SEs7ajrH1e6CgDbmYh0Yj2u6tQYI/HIYFM1SJ1ZuxZxTR
u5cjX7il+VgqbZ8CdyF4Ia31Owbq1qoZ7NdzUZ5BnoaLrbLNhO/Sgzkn1VHu
sscOKHueIcvR1k66gWdn8jj75jtkMe6rZc2cUD0w4CfGvj/Qy++ERwarMJQq
2bwoIB1jfrSSEWwD3YW8/XqAhhPYcPsJsaG8DxPmeAnSRc01AnUN7J/qrpBW
y8hDoxHpH6hL4YSzniNqbBFA9FBDUYqkMXqpIdH09F7NzgDP6boFgkHFiQ/0
Xgediz74CiFx2trnK/ahN0TVCrLHtT5iXxo+XV6jqBBqdPP8zehtB4uc98w2
p0ZkEOBN8K4Xgv5Lenm+W0TqNZoXcfXQCo7s+yPp74K3XfeN5tIJQY3nfkf9
pa44CIc14VjfNLWmmH2vcFJS1ekJdhlpT2fHEkEtchxrGLTA3kb87DdWFTn8
SLH8ZYZhHDg+P++lYAesfiMUKxcIJ35PGNNaU55n624fJemeRlkBDNfPgUEH
5dnvLFiYi5WBda3K8aVtTmXOzlZtPNDoLhKpRc2mpTsAsAwQx+N8BfeCRiYb
AbE7GAraWybuP1bz33SGu9klXXXp3QnNgL1j12AIzMvT/uFC50mLLSjawbrt
dp/l8n59DSjO5CtOjpYKiu44883kVVq+53FWDyy/buVYtuOJk9QiGRkeQVVe
elZI9sYrmvB+BbN3kyLJ0ryjxMaO2+boryT3+v+Ge+9wlKJL96QRSl1ytYCP
aotn99bO+3AQIpo7REh885x3NRym2uEbMPYZ7ZtmCSpc1F0qHKSDgjBfuNsN
EfbR5DvIR+oGm0kr7nv0rlYz9WoydhrePET1Q9lAHx7OQliQxqyYJsnScKw8
wvBr58VIhZ/bceeeye7ITBhmRyhri9QTmPyMVom0zjNwDofJYj+HZXTaSa6W
zXFYc8diXPfiRNyiO7ZbJmd0fFn9M2wPgv//KIC7L6ytNmigVR3lGNYSjycm
7HdWZ+wQ6YEqhhDkODyO/SFX9yUeZV9QISIwEf5CMLRWkIQgBCCt8/+CN8A7
ZVvNPg0DXRJBf9g6vHBeb7dfeU40QC+A97apaVuubzjZW6Z6hl5bbb0YJebc
HxzsVmYaX6MlXgFCdFo9bhS2qv2En9M6bh++gUJJqHEhJUrEOjKlQTmjUBxs
cI9oROHuhXyNdfDoAJQ5+74mBSRFgb5AEbkiCnQ1x81KsJR5pL1SCBHaJq/2
xfWeHOmfMSSQWzRpk9n2I24M70ibLKpq7BfYlvvZoTX/4HMBbx9p+a5wRPAQ
jxIBr+sy4Hzi2vK87AyJyCATwUdTpLi1tFVLIbrkyqM49NC5LWSV33AiYQLS
ztmxoO2aEks49zv+uaH4GBc54C5tgZMQ1JovZUKqV+wdiVuAnoh+iskGXh+y
sExSPrGoEnkbhnDWWOYymRVc1HYi+XPmBRAoG9sGaffVOzX2Qs76qIUyQYcx
yRY9GHQG5IXcgdmPu767WgzG80tVWLZZeD6jmOKUkkdCDy6XihqEt5Ky/sIa
VK8MaYZJ3vQt3cnzyG3SCCqfo7RRwof3dUYH3+EaWFOMetjaiye120nqf3dV
nWHrwcPw8ySxDltzoEt4+zcx+nhW/u+B0U/s7/Ksa/HWmdRU3B612Gnax1Di
fbCBoM/J1hfALp3rOmVhPewIVCzrMcXsfeNtfxZ2rgCId1xsUixy7XQnCbqi
/GoLTTIPe4BdF6hyHvj/MWPtsV7qnoRdjNSHcKca+Y1ezocGQ4a80irIojhX
3ZFXyAmvua594tnQQEfCZbVhIF1IX/GL63+sZ55ICTiLhmpln2Mh/H9TLjzN
Bqs/IkbLrurE/8g9WE85J53kekd8qoXeINmCwoI69DR0cbtshQB0QdhAZvq0
UT7guNnL5a9hR+ZZnaLdWvfD88Jc0PAp+fRf0cbFqxtf4i7KlPWlRC2PPvJr
2cj3vu30b5xcSte1LecEsei0IIT3/WNBG2oVu2yKV99584XMr/dnvTPD9xuE
aHzNaxhw3QLEorF/cA7LGN5W48G201KRqI8GBogJvYXgBUj7oYgo3H1gcmMF
rtVUwD0GarGdFgg0lU6vlyvewzE57+heOitko1kDj3EwJDDMT8gsM5H86xRZ
s+DiHcYbL9/rzGcQZWSCOPnPAco+QYGYERUxigwxsad+seWwTKI+RFf2LKay
4YAzDuiU3fKrKCptqBK8zh/X5chqkHn1/AOBj/vTXdzt7HcbAlljFU8q5Na2
M1dlyWarKG9q988YNOJjRujtO8OIivpLbT0Xtgs0vefGdCQ+sekSzuItIiAl
kOxKK+fImAM79qgS2+C1nblEzldVrQ7RRTuJAIk2FqmJKALZnpcb5TuNwUpq
xSeP5L6UouV+enPrkRH7qrxBIjHVaJVlyr61r6X/HEzQl6L/aOReKCao2HZo
NOsxv/0kYX71PwOw6PJL8dY0rn61gD1AZ8Wown1u3WFH7Jvx4rHy/KGp4+y1
whMJT4dwEHQbGpcbKx06aYK+hCUd3psFvvLdNWkTJu8pt6ebi7c/VNHU7Ipv
kBmH/X7EopqZ1G+mQH2UniscbhHXTJszuSdnMElPP8ztrbg0wyhFYlgF1Q9A
/bkBnhp+6uus8KcB5CGwPh3B0NEoIrhST6cccL8v4Yzf4yFSAPCKF9f5Xlbv
wpxIh+P4PPu2tZQTYYbpBr8fBssGITwQZ/Ca3EZwjZyS9o4nK7Ft9cy6eBq3
lXrHTuxoiKy3l665GeRUP0ljnnOvSv700jdBzB4SmhF/TdIwn0mErpwl+68C
Mwo2cCUhgpZS9F/890RVBEzREbmWRWLJJNf2KG30LTuBfgEfbJqWlckhD6Bq
KduWxkFnaf1bV70t95RbE26uqTXltTMgAc9FuwbI/mtewU2TvbS3A3cJVPMg
l/35sfyBAj8GLeJOG7K3bZjspTfn3HNegu7HrNXo6v/UgO3hto/wqYfCljG+
5CKqZ3fWclYokvt27wMzughuhYzcvP6wisvORVemrRfBVXakq1NHrGi/0g1e
bU6rZlPGAc6TSXGt1VNJvbtQwcD1q0sA+qy09RmZ8wdq5Iy+0pNvi6ONby4z
AWvwXljUJkddbfIjx+GltLL4oqVxKHk3lcwVVrpQJE7Z4K2ee/rf+A+oRHaq
E792RG+AvyGaUiMsggyAQ6DyucwctOgiyZVj+mSSn+yUt9ILkBXDGGTxJQ5S
v6yboXPMIEqgRS34Dub8VJoZlAL7gCfGC3hPO3xbmqj6X7UWdb4Thf5d+bh3
6WhRGPJv3yoNQBrot2qRIKWyh3xHoyo0r+9llO6eoXW4Rb5N/9k6jBGXzelC
PuG7fRmJ1xdAjmbUO0eOv622nFxpROC8RKhLBINI1MuOIOMH1JMb+hCFCqAa
4TgX5NjJmgHJBFRvPCR+Wv3bokUc815DeXzNFJT71mHv2vWRS9Csy36W6prh
8Mb296hMwbmIXlOd6RDyiXIKbVXGcey6+n5xx1E8d1GX2DKHYmoL97vVV611
D/toe+aBU2bbpug14iRsDlNLEMOzmWojIbLIRlKJi3JGR9FHFRSbJKkkbSPD
G2A1J9dymqYxLWz7pDalrCFOiuwCA4lPdadkAq2+UcOygFWKS/5vn2DvmTnF
uuWNbLt9/zbJEuy1QtmWpnfdQTdzZIYUlWO30ghbfDeXwP5jqyMFqCLBD99n
2xmk3nrERYgXCmOpKgScgt9xaSWCqAAVt1toWjjIzyi98NgBmjTr0YaBgt8i
85ET6trbhGRs9sgtUu56zsLuuROBY03yJUOAo+2QRncPy5lQMpyvrpG6ucoo
JMwcFeAcYeUR9WboOIlZxzbrX5ejBeKNrE2Qrdi6x7CHl6jjnr0R+QaWvoBx
HVFxB3uXhyQH6WgaSSE2ob8MS+A9qMBzVXS1bjnuqxauBALRb5tjWfmINyUr
Q2uprKvUjGwcP3l7srJYyJ9lInnMWKiML4+DeMoOJNEVHo5VkBF+7meZyCAH
s8nD70itGIalTx5tLj91+p4/13BEBT7yRDpd+yEo5BhbNdcmm5gR69uIgCj2
fK8AJs6Sn+jNRoKecY4GlyzS5R2jEB1dcMSLIKsY1NbMndtMq8L2dOCy2UQI
+QTi+lOochxwFrmsughmcy6MN7d8ARAvp4hWaEMWhIbbMjexVzBBazhoUSri
xxe2eHyNeBEj3KpUE2cZUHTGAxUtuarMe41c20c/QVsreGbcMf2C4z3pL7/H
gGiM3ohlxAQQGOnO5fZEDBc9N1UdnzwN5Uz5mmn6N30K+Yqk9XePF6ZnItPL
bdp3RgHH/hC2m16D7vad/KQzcgLD7ZK9799gh/5+apwgrfByPzJduDQJeXWR
MYvxS/yND8VRZoV60RN7Yu/NBE9t0/+I1Rx4w0UyFTt+Ql2i+RrDAn0sq3uH
FlTqvV7nvuIH+gl6nGevpTTBAT6YGyVsHZiL9xeX/ERjo4KHG66yyZSYSOnz
+e3j2bKgU2yiyv17sSFqfURoGQXvPOV+4gNx6oQ146BvFSfBzPPfJqFFPBHh
bjqh46cZFUHNPmaRaurQyDq2BoJ+5gtHrqRLiZulzx6qvQqcb8mVeuyInlJA
yXQM8YFkFhAggflelZbkavZAl4oW64hTqiu2DJzqUYk4Ai1X1e5JSSNI89hP
QT02VzwdPzcuSRfk1InRD7PJAe9QwvreIMItmQvewdKEuarzdMWUQpashJXB
CdLBqm6dW7TXQ0iQY7QzH8V9VVxJW4b/TG6B+09G/J/Yv99Dh6XLzfIoeeFo
m/xS0cwNg39j4v8O/+XS8TVxtr/AJogdxtNcThv2EpFytl+AjCGH+j6/LBSZ
RhBUwUAtZf2J40KCpzNz3QiSe/0nPHJZ5F2PTQO0O1bwbHm9thmRijG1Hlyh
aowKckgScNC0bF91vtKtmzpj6yvFUtkM909LX+jBp4JMjpvHFoD9fVa9uGY3
E31qGEeRGRYjPA+9ZPXFkmsEyzv6dnsT7CV0NFjLOiCrpKQcO24zmU89uCki
GPh1cDn0MiQ4ZYtXJO+uVLH/PIbXQp/dP5edOoEWLvwJDRk40ZZKBDnyqvRc
f7NlSixVjJe5GAdHuiSb27nMZgJYSMg4zBkEkZ+6wh5MQkEWJf68DD/YDXUP
IZTshbODESjtFwjJifcEDJyK6bny2o+1Ca/B1XzmNjCd5H56MHUkO7mfT6lb
3iNBfZJmzhiDwSe0+ssJLBpxPTiR1itdtSIcneUdvVPQ+zB5ILQfORHUN3kj
g+kk7t9w5zgqC5w81x/a6+B6UIG0JJcJXE0b4xYDBS76nMDkU0Jsifnm/3rp
toD27xHBhTnPp6BOLxnEOsYzmOEo5gMn6Et9ViFU+w/A0MZcyWQaND77dmqj
qovriot+kAwp6tmmblTVzK3HVENzyzPT7rdVjQ/F22wJAQER8BUpoYwphjcV
EsNMr9ZcegXDHdpeLIv968AFb3/x/QkOLE3NOBQ0IukPu1HI1rbdfGvp7TDy
aEQxkibFaashyL7HPL9p8LS17oi3O/oAPeA1+VMgjbb31npLm7eV81jC0yOR
KKqAyhtETf7wVlpNrTqfA9e0mGnm8ivMOAYk6Cx5D/QhNClvRIMPZAaC72/y
0yE3c8j92//4oTN55vKegBBdZUoj1+9KZ8g427LNrAoYoscT4mI1FqLbla8D
dj2Cm1qfBj6oQxi5Ih0oODr7LaaCWlsiwd1WA6MlTkkuvpD3maNCqOBd0iMB
pBAXybDhPtUkGJQMDOVT+SIkjVMEzOQT4TtWEMjTdplDz3gWLSp47iIhABZd
puXuOP62SEXW7NBmFzij/KCCPJ3o7ykZR1g7INF40dxye3R+D0gkezNPT7Lr
scE+ULK5RL7kGEknK5y7IRCzMviRRicYqlG81U/RZEchT1D5EzgoFPKap5Dl
hKsmtwh2rpmumjUR5QAL8112cRQiKcKNK65d44tWB5boVanzmHgR0mGsz9U/
6sJrZb62M/siMhl+fC4tfD75DRjAyOnsRhX3R7DiuykL/XYQApBmkRWAcLPr
00VZLsD8m+rPfRlbbx8JmETSLwbFk4vMEAMMrNSiCIRqFlkAwS1adoD/c5Sf
HwnMLRg0XG8JsV16Q0bRqojaOX/gNzp9Y04y/rrv1iMvQfWI/4ntdUXemyyT
6chz0sDFwC+oydSZHxfO8SkpuXLyDpX1JOl27R/G1bVQn1FYEKq8mS2nAbnw
qIZ5qzfE5tACp+Dp6oRh0CwXtDss9JlFh12VLMGRqZJXyTqlXnsUgnf0yUxI
ticipz7ywqD6WeO460jw7hnONjQQjVEpi4HvDdPiPco09fGx5wFxqKZ0mf48
MucMdrFJGGTqHR5fnA7CAXRv7cMpIZgN00hax81UouXMrwP2BGRiXj7hES66
p8Y8wRbAb8ombzSnooJm7PodMJTxqDIFY/AcabxXj1PQ1qAiu9f8xSerOP0N
MBE2KkUpkDKbiolcGf8yc/N/18VcR/PUR1JAxZPJOCU1IYdot6gnhGj+YMu/
pWZ9NCWnmTLctealk0V+CcIpehCBDcK+pXRmFtghML3MfnVW6mH3FFDUycHY
vhlseUOGxksZ0Z0kKSqO9/i56/bprOyiIRytwKpBIZXpfHpmJv5sWBWKntRO
MiaVgnpDs6Ny48GwaQTpUfpjtdELfgcKNXtDrmCvTxpEp+6oNUhGtAi2nTvB
CEuB+eAEB3UanFyg/xkK0Op9vagIyaOUi7SUXhLA0AvI9QPVHE1YnHMS5Kdt
dr54bjJOby+YXCmCM25OTvAZ42lJX6FgFiLguRVGe8epa4XqMU81g8DRrnua
KT0/GwtBTZFzW0ODTwR690lN1XieKr282JOl818gRy9XW1gWQhNKHtTzBMd4
WAp9qOxH0Jtf5UkWFXD+attqLSkPThzFKhh9G602qXSX5wnJm+WZTavbXcFO
GBnj1b6RIH23Qu8+FcBxQdWc2lxvvEuHo5BRYPqL/O++DlY8h2oyREeYlR4G
Vwg1gXtA5Fn32VjTM7sk2dghAse6tpAqR/ij0iyFNm4jEKCN8yXq2xMDGNxC
19MPI3eFiCGMpPPvLI5rr4S7PefZfdEevwLftHyztKvye5+8fF+iOLLgiP2q
bkRWq69wVcFJi9FNPmj5hcYS42Ld2nAJpYmWmrdgiZGUBzk8ZHrZmDlms9V9
0A4HUQkBk/p/DQ5lkMK2v/9NUnOsVR2icnc/aF2GgeXPA7L9eeEszfedRstr
affNtlNxoSTYa9EODWpKabNjpUYFsFUjjMigyPMUcdNOBa5j65pIT8If1x4D
oFfMcfmsk7s/djet+RYuUCl+bAro3Lu0wLOEQWw1y8rIidh+Ogz0VXBn+o4t
Gf85vGE7gPw7wHuHEJw6LuAcbuEOwQFDrDOilattd1r4pZlL5xRK56eWkD1S
7bgV+3+X2QwEWQ22lD7hyXTcb5qPU/B027UgZtM0LHujsYdei2ajWWPpp5UY
Hxiicl1EjKaxSAUJmPvmkBfve3DKDIeJW14mBekY2iE4zqkPM6nyABBj58sU
Bgb2eFOku1iMXf+eS6KjrBZlyOyb7vZ3PoVuTBzL0tm5FBAZusOBH+13615i
10ITysZ9Eno8+hwzaQHrC4Le9LL62YAPPBLOPtca/OAeaKx3JVUPFX5XRGJx
vjwrnPXrd6VdF5vDYTQdi4w/adAI4nfIGdHV0i5LiseL7rXT8ylbLLzNqVNJ
veb22kGssksqRkLCDZZwFE6G/vi279TkHFmpd2GuU35NMO6VFrL/K5tYxg1s
3uKVEWkHKQWQXAhZaNbPvaJBzDmrLZSSJdh2JuNTVhDcKa+LlB5eqle7Ofbp
jzeIgwHjArMFfp2FmQiqTQGqnF+U9uQt2dvmNmp/Lqueq7xIxWiT+4O0TYb6
6FhQofUdjLplTrToAKEEFFryMVlxF86kD5J3iSBq65roRHQS5Zmkg/DRFIeS
ywd2b31kxqbrJ+CjLAhaUNWu8rCRkCRZP1sW5cgv9BUMcNX4VUatL+YIZE1y
JppUUVWPuyNY/j5QUXtL5TOkRC+pwRKeW82x/wEgZcT2ief0o7Pzn/k0NNj0
lj7IydtZzeGn8EL8a33PZRzFr8supT9CpJpgqBEGIpG3DHaxwJ+So6VNI00L
+yWmRVvd9J35aYl7LoLtg9y3IaE9iJ6/8OUNSxUMamSMz0l9Wct/yKLngzQ+
spdgg0LfJsutyRY6gsGQuMcCOzot30kLaazcKfMiq/TJ7hEumFzDCGw7nN96
Xv/tFmQQoXjOqMeuIJK1Gtaig+rEGDqt976M0U95EYxzcED1AYwIOY7bw9MQ
hei1hO+6QK7X3dhVNdOGis15MZLhWsxiXCTBG7kYGhwbqaVzUkEQoKSSQ7d5
M5gkodlBiARO1qoZvYrbjlaJE4i7iU3wLI/8CSKJFJZn1DUjH+DaogfrYiet
PU3a6eRZxN57N1lHwHN5pXVDPlYQPSYYrhBNZgY+OPygcDQGzismoXMr7OlJ
DP5Bq+6xaKiOA1dE4rqpgASi+l96os265QFZE2xJx6YmNgDPd7fQemmUnIEw
fDHCRUR6BwB+tgUffJ4zdlSsUTFgismPS4QAb5ojBXhJMc5m5D73DBTr0aZe
nnETPFkHqYTJ9SjHQrE15lGf3Ff2yuOxsDwJLlWmTSbaA/QksJD+9LTwNHw5
ZKOgIr4hy/TNBXRVdNjlZnft3JSB3Mx9yQE/rV9QR37spruS/dWFOw7/rhpJ
evC6LDDvRV4+2Y+nQS9TaNCQ4wdEBSk40yookn3QgRvHGa4GIWyQ6/TPxvO7
jQYchFGYVMwy8haHNSDAaK0bZgU7LjnMP9YTDM9wBFPeR4jtTzd/PxvHhDLa
ewq/g8PIzjIgQ7MSFVJ0gq7m2d6dXZKdiC1UeVpcMlU3fgTUGbNVwLBkPfGR
J8PLsbz6cK3Ru4p2/eVXgjxGVdvi3JHR2u3qzjJiL3fdbSJgMuJg0TPy/Apn
H3KKeha8+6DCU1R79mP2KKMBJIouGkS/8gM9ujUrFOwpGHA/cAeYrERk6RNd
JmD6LSePaTbOYlLcIBeye87Sa+O/CcWm+XqPXX/wQqkRB/RSDD9TPU7yCf0A
SZGZvqkv7L8rzXxDE6KKgs8wDKdq89I01+AAyrBj8wQga+VfLWnE0VO8pVtu
0xUVQgj9kzfrBbitxv0p7qfQehWzngIKriBAV2XzsTGTQ1I6dUCR+ixz4bGT
FOJeS8mhvwsfKfYLbpoYwTAkXh9VDDCUflLanUYJ3+4ETD90z25cgtNDGzlr
ZZwzWNW/kfKfeosVKaVgScg7pSbYiMsQC1AhkfL8rFnSlFy6oCZkPSH5+np1
gtzayL34sNBYTi+C9mLAfQboS67qzVI1ibKGCy2/0IjM0qZ9CkTVS5R5M7+C
yr9Bh16wrgpoHVRlEphPS1+z1Xz8iSoPej3en/ltFZ4lOR9VL7IKAdcuf0pD
ahPS+rMfMJR3SGHg27BqRkGvWIrr8sAqrZ1MPTeArc8tLrTsPnWPzA1psceO
+ca5oL9IFvlFqgGhMN+x+ce1TJQga32olf7Kqt7o+iJGtWkPlLJTOKgS0fag
k0wZSMUH6KA5mScFkOteQEibCMivOBR+JpFBUV+UrBzT15tqhLq9vgyxSmsu
a+c1tz2zSiGv6tskLCQ4Cx/41MlR5PurAmF/neGEXWoGkw834nQNp/UKyYrP
op1/YR886i4qVCiJFrWSdfz2hi5xNjXBruOazJI0bfQ8Nqig0+RYcJxTJ05c
jF1jEuVL8DYNGOTBwn2q0GRdiU7LUzHN2qxzmWpiTvBbunAWFYy8vqKExi1C
1ti460qqMJ7STtNxQQRZfa7V8VhrqtjmEbmHz1lM34w7h4owanonSmdK39OU
Tf+DmhhhXz+IZw6y7IUicX0IzdrKm0E7BSct/HNR7okdepPpRZ0QC5aKxps+
PRV4CUuky8AzSmRgznbEEjb2EtWce/O3CDuG6HalFo9tQXny8vSCut+1H2Tg
d1vQw0EN0YmT4jIPHDIcO9umV/faYF/od1jVDGyIMThLDk+LsOXwD/jN6y3l
qmpc+8jwc3bcrVS8UJVwL1Mm3elM8NJ/KAng4UYGUWsx8K5S29vXQi98crvP
/KWY/XuD1jUjuiBWHjZp8ZIvw08EVci+cvxhF3JspQfbSqUW3XiAiTrAdnTY
oQkNLU8mLzihrdOtWDruqELWcp9dhAObhRzQ2rHdc6vW+L/bKodcnL4VEstW
YZxZpb+7qUOvX8vM0NkNe5opo9xkpTsbZuAn+d65+2F2xg+dFwY5flk22dDK
BiTtb6LMKh7Dqq12rL+E/9gJBbMswCviBgqxbR0sdBDFiAs1ZJhcWp6v+BLk
QKwSWW3n2gO5wy+6Xt0Ex4XEbX3IEhSHEfZoYYnGh8T+yce9sYe04G3Q65wT
t3tRzGBDW8BOh5l9EIvdL3YaybY+hPhHVS+k9t2wQpVwRoTA/b7958OUTUN/
6XYCkQzeXVDxUKiBLZZ3t+/J/8HNZlF39ISGlwyu6/KL97ffETdpPgFnE1d1
u8Id3YFtB5G5TUdoSbHXnh7yH0RKkDoAOx07bqxiRuvc4AZRPMNR92K+tMMd
IKKWhlMFYug85XFDMlI7zowngdtzTtfmpGJCnbnus/6m5z0hHfLBTrpI2SFc
+52qpB6heRiEAIsacczGtjEHIwskO5cRBK4qj4JrikPNNfNfyGXWpYHP0Dt2
t8kVz0kq418lDyPpNwWqkgO3hfBRSvEqMj3RjAk6a7N3bBRwhiI59AzRWoIz
1LwIl+4Duw1tU3PZQyHgktHzN7tqB0CodJ53RsT7l8HvUC+/wRWlj15tdHYY
5RZZQ370+CD/nIkG1AXZu+7QpKwVjvGOYd1m3+oqcHBHBtva7koRebzjxxZo
x2dXW6Hmi9dswIgGH18e1nwlV06ekIkS0U9KWsE+CRPnb1wmGRblSG5vyffL
thsECYMXfaD6EEflAZLXZVSbyDCdlCgEpPNNoJxvBtySa9JXf34bWNw7FTf8
7LKNHmC/2tVi3TcA7xpZWQs1k0cEBgGtBdDxSPwb7jbt2kFViB2SafmFVetp
kHcabkwNyA8dIjFMgrlIhWjyOhIDC/4eqbUjTjCI7jee+QAdBbkvS9/uEo+8
CzOTKfLwFfe2KFQWmboNh5IOT16Mzs+AKO4pfWwdIOqx6c9Do0+31Nsra+cg
cAalIc+03YffegSFvqpM440i7qEsyOacma/4bRANi10ilq0kjlz69KTEsrt0
jJDpTYQZzp2lViPkFT5CXkK96xmR2kQ/rgvy0ZP3X+rB7Phy6zyysSLBhID7
Aj0IxwTAi8wX0KC+YLpmrhGJPB45+kL7DJUreXA5hQ+mgoCZphrnHZ6hfB2r
SDOphTbQvpTtQQc7yOAENG+keimPlgXZN0aLQuYSMcazCXq4pMzIxlM8zCoR
WZMOqwgjenu0ePGX0xiVXNK1iMkPdDsSnz7ZayqUEFKdNi48/7we6HIAtGIr
/1nnlxMiFvJ+t8T+0ny+TfqcjcsG/EBlz7bD6Rv7Xj4MKwipnm1sKes9ofCQ
/oj1PxcI3v5HkF1cc2btgrhe7hkrmtkBb8LUr5prdijEjfXVJiZ4owMZdqxa
JlRsXAonxycWN5cohH0lXnqdXsHYS3waPGDKsUElvsoFmwY0cKhUtrk2/8O3
cfwKNecqpInFOuJWJ2Ycjh0JhmxdZ2DmQ6RifZGpxNZoQCz4fFp8YEmYMX92
8rUjeAk+d9sijeQ9HleybaSijEurlPU2c5ok5K7sxy3HTh2GxXO52thrXyrx
/22KGWsXvw9n9WUqKGzjBbamQ+uc8NOYEvfN57Z25duA3yVKdqz6s433W9TA
Yv9LrqqsWzMNlWnWlFoDw1vpK/B65WwbKntMWr51cWRnfCmCnPjOz5PhOahR
nE2Pd6qrdDIM+Hpd67/cm42NgmQKN8jVf8sSWGpliuthRvAWmzrQXobYJTJZ
TVXlm/ZlcZuGzkVBuE57IuuvW8x4mpE8Ax9ErP35bkxehIB4tnULhw4Jg7Im
lOtYoMBfbAOyRshPQM3VDBpxQatXH+GbdsUHfsiYMUj2issRqYyZ/J4XqvCX
tsOMVZeg6X5nQVM162Yy8O7lgc7IxfUcN+RQhxn6gm3mVuVX6yIMb73aGpZv
7umthUMh/A81B3zN7Y+YxZOtdYjxaC1OqzZspVnavI0e9GiAf2pgrvR5Pu9e
iZ3EuwXUuJ2bNpMiWhCU+CtdOYBYFJ/rHG6Na84Q0JF3R+DcZ2tVJD8FXKmk
scIc8yaOVNBP4tflIeRQPr7AqhyxVJZBDvyQRfHAKGOGdoPGW51kpjTIWI/g
tKr0r5mLYDcO0lbR1Rlm/xf/whQo5oAaMqKvxL5HhapSUJMj98juaWnXcvd/
eJiRsnuxeaUnH4HCi0gEXwYAyYYq07JMwwVlT1cnkgXuMGd+ahkuksFGkqJz
ttTm/bwPOqWFY/YMqTIXIwv0YjVcHL2Skgo4lFk3RwReyxvN8DgNyDb/SJeH
c9gREvGIRmhmdqD9LTdGVYs1X13nJwf8j/if2BNU7qY+v4QLWfXE+sMqqkG4
3WMTmU7/Ta+j4mYG/fVTguGkZm51RIvL3O1sdlKLZgRAW1M3oR7avUDCxU5/
CcCJSXSq8Aog1XuDpVnpYGFTyKdfDsSz6uxn+skIfJb6abh1IUMWLNlHiEdY
6bRTdkp2BlOREDg6WeG71gEEFaGdCQtuwjXI77JqSUb0h//0JH3JadT+5rEN
FjV/kuri7rXbGhuAo53Tl2uoAkqD/xp2E/Vk78zJfc67fIJrtlZwkR5TsPwf
Ed+hNd2+2Q/FrHt4MYbDBlwREf0ykI624ssMUapuH7ZtUC4vK5bSJX/EKSmk
LIgctU1rTSo/rp+LmSTB+icOnpxzRMQM63WvKB36X9dpMMBQxQ/zFYeHrLww
mw3F8Aro1V4kRV+Rt+1awoYIxYtFJbJHQbHt1ntdkqsoWG9Fj4luR6oAzdCT
gaOZHS4pzU5qFTP/kI+IHuKc1WggP71ZKaJHnn69QKgzGnuqjiJvxAPPUFj2
TEbIoCYPoMZ07BOsMIF5DvtfWdrSyeuQ9Xy8ANiBoJMhLY9WUfIxmSkHkrPv
B92xeOyAxrUiuqCYe3u2eLVziHM2zncpZgu2PvEWr654+u7xRxF2zhJ48Ibl
5xYAwJbdemtdbo8VSS/HT4hV4uNHFfYDocCJ0/OzwUXnMGLcq84tyzkO8Bta
ToehRqOBMIE3l4JJcmcNijEDhgwmPBSVsBpE+OwL5PhOgM6K/T4DJF1LOz3N
HcJBz7BZUIOBPSeM+nv6s4HnFAQHt0bbWmh4CEwGFmW/6gLV7nbmr5gt+IVW
fP2CfrIs9qXU+WMIcOQah7/U0sCUP58fN5T7Zp55VDwtaQSRLjfjACaohQdg
UqfzkrG7CngH2t5hJBDCFtadh+3sr/7a2FzWn1cjwL9XGc45XBZxJZHw18Ue
Q7HEk6hw8QtIqzKZER+kTtmrZMb2tUgyUGbbjF0gSwhaosRP49qk5z8tQ/Xb
JRvtWEvrM4cVoX5oJxkh4/Vw90iy8VVFOK0/MRbwhYwvTchs6mKHeSmtHt63
jnUNQeBzKDEebwWmiHnKzL7Ja4F118PBDgDyrSAc/EWDoLt0lsTaJkiGPPGQ
fBCxDfp+pxFDlNlQJxalR8Cu2wWEh0+eNA5Je+BYMAzEsQF3af5HVjE91ua4
2sEzCuZyEYjBBEHVihpwod/TYHpw4nCLgEqeMsbdzzokwlz+6g1vGGOV4ori
F1GYLXlRJtelM0CYoCemgmKHpmJ1KciD11834hHNaU09tIu8W7b/QmKZO0tM
1tvmLvuJ4fe0Y/4M+UrKsO7sapt/cyrBPdvzEnfP3SN5rVK/kD0Tbi66DW1w
5XC7S6FwNjdZQSDYpJvErZ+X8g2F3ilieklMPifg7xovSxs//w8qJs+WSSG0
Ww/FE+TZsA/dVVTx+NOPnEcMuurflf1Le2KnKEDvXSEGG4sRL9tYH9+lfHrR
Qea/pkqUDHckaafVu2DcnefhVyGDNMsPgzNuNzLkxT/pH5Eh80RiNVZ173OB
gq5CoBFTKqASA7oRPQoTdyrXDGE00ZHC5uew2WjOmFVnjMK+1dWDJVNZo27F
SKbh8ctI1B9QnH/ZEHsLh3sSUb+KeBfHTQJGWZLXYyJejU6mw0+ZhaLTvwTP
q6RibBFpZ2bLPaRFMGSQd4460zJoHjwx1UtTSjulKrLLB0BK7odOFlOJcA0D
8521EeLHgZdkvbnKZzCHugtToJfoSjX4/0D+jGhmlB4tq67Accw/JewnU5Wr
89UGN/Z0OOqgq10esyyPGTZouRVGqCQvxw1dziShGEIIsVBwVIEHNEwPqRTp
aT0Dnz7WBTGQSg/XTNNQxUgHCfKtd1um8Hs4X1clYqrbRG3FyunZ2ULLhxjQ
CcTFXzF0oATZ0LeC3P86f5Ha9xpBofqGmErRdydaUNf0yaIB60GOGb2PO51M
q0o7GokuLQ6hUYDFdF5hHT9YRzD6cq+s3eLewthbL/5+zDi6Vf48i+HCjlPU
wOcrvwH/cmcFxtEnz5elY6ihiJ4KRE9rfnosLNwqR6U0ByPwwU8VUuaaL3lk
UaHk+R1vJ6TlAvID+K1VdzvwKa6bvMK4nUhPCUJZxA0g/BkmuolpCyZ6aAt7
cDm7kOO7QTP4D3/2Z7nn0nWeLzKYGiTCEMv3du7JSiL3amEYqkyq3bo+gv8L
u7ZuEbys/Y2VhPHOpKWqSao+f+urn8cW/78tMmT44Ko+YDg6vprIruzJLeXn
jkVQ1wt+aTimwJa7h+mumA0EUfzWe9PeQZDSJdsNJk7iJn97W1u0vwSOrGcM
ZDtiPmOjYgfUkeOFF3JUaDzsm09Gk6/JU1fejFIvWGMnXvNezADoFhrBnzgC
EY3zNJwPUyqrSPklJd/kXHtE37UH210ul5/8fFlR9tLnM2L6NNLIXT8qDwSg
s/sTWKazOpddRuSRkR/Cq6qXPQU8Ha50LmY1JCU0WJOXAfNH1AxpWorJy/pE
1srrFXzmTANCs/+c7zQ95luLDy8oJH+enZ8ecBFWQKm0AvIAAnsnlGHudYYu
yybxIepH0wQ2mWa9uSFc7k0nz8xGEYKbQJtlSNY6b42HeI1lYmLznZXK6PWv
nu8PSbAj3n5aKlL3DyXZMkCnsYKDScgdVVekdTUZA08dX8OO2qlUEVWhnqgC
xrFUqrMCHMwVG3kY+QdF54XwjpKC4XcsJelMJZRyeBRvoAEG7D2unsErr0rj
QeXfXaz5veRiYpBbrxeT6jxzhUmdPjvp5YZO0wchZvXFXS70qhYsbXnmJ2Vx
NT6HWOdPtGlaSZnjvmaYTJ4ni6rumfxwR/PrhrIc/qv3kAtf1Yn6e/+cw1lp
Wn4PYG29r8flzUyVM+q5qj3AN/1vVfHF0daY+5lMGeCcxFOexoj2c9RL+am9
J0ME/6N+eR51+tAzrEFdOVSC8TWGmB9PRG7aWv4m68TClFOj5zD56yfJCJMU
/gWbBg+D9JQ23aVwrT0rDYPZ91hTMt6OoY1M77s+AfptG+lOHql9yW6f00ea
pr/X8iJPl8S8+vlvRxNUJf+m0fW9Wyg8HNoTvkMljOA9O+iBZl46phH247VB
N0aD1tzSph8BUJjXYGBqIYSIxRn7YxHwTmdubrB/oVY3SO9tU/Y9XSG6HZRV
uoB3AXA5NtUkS+P4AIKzKfadNHXJ5wqi1AKG55x8hiRSV4EJUqbuVQlsL5+G
pjyokbgOtsWB9R23YHyJMyjx2hxLCYRQBznrBs+KDzvdd6/Qr7iBphzKvB/g
tx0rniqs1Ise3Tx2fpv9zWNWozSOlnliVd0tZdNmkKvb6oonZXAbD2fhmSHk
CPHT8pec+0EihRwWeqjr4aJQJyvwSO1zbgbQDsBk1Igv0hc0eEhhusx/lcUh
UPJAQ5J3q0QpB1Vl8heXlf38DOpXdWRpwiqQdnNUxCvJf9HKIz7lJqi2WRwn
SZIAKoyrHJrLtEC7SSK409IyqNjY4JkNlC34IJH3mzm0o4h9h8TUJpJUwFX6
IfJqCepPoenJ5fM9Ii8bStGhrXtiLdxJaXZ7FWNtzaZTcEZsMNdoTifX8nUW
ZVSDC/RYk/IwzGMhTn9j6HdhaB+Jyq7qaFxtyEEEEyXTNRyRKQI7W8bcnzNn
05nxN6AlgK7ngsCYu8iSAe1BwZ5B72jFwKuvqJbkyTUdGg0/MjCrOPTrKewI
Mm/lF5ENko58mvt8c8C6aDJ5EQyTdoJQbmjX0xEpLzJsb9XrYEDIYk3K/cnk
et0GjNCIZ16OfczERWO3geWxh8PmXP1i0ZGK8NZ2bNjglLw2nYXXF99AOe83
ZS12oe8Q5PdCLIbthI41Zt3YDMwijzHfWSiq2+oMFzCD4U+f/CiD/PwyEUsZ
1DFsbScqf8ALXYfLdqhCPOO6d7sbj3UZlpXoI4Pt2mxkkGD6U2zoS6+qAIh2
AmSDdcrBVQIzWXh4wV+z3aXGz8GBFUr/2V88RGV8tsI39exM/ZgAcDv3UbOA
VqC46wHuWNzULem3kmNMQLXbNyXN27c/0kXtWMOQbeC54LSCsKaCf2y9j9KD
KpHeZpWXOJ/co/iGfZg+IDbVrDafC/IznvQ9CQ/x8DnDT/P2d79VX6jYo99E
+FXsXHIfnVAE+6ZzU+FCrXZ4Kj46xojhQ8gpiw7Ew0y/STvfwUoIfPJvc6Yq
SDcswfvycEcHiTblEx2jyRk9TGfLandzmqsvdhIO9PQlE9ziiyfKPWEMIu2o
MUAzkyUj7xjuUn5PwTOEAA361ucKFUpIzl3BwnRcf/FUHo+QbKefw4NQshfD
wpwU7e0UVcBrhA/roKWyxrAsBFd/C2X/3ru45TxhksWuHGlG3HaLNdfwbtuL
M2dTCUJV3TWt6AryVsocMecIYHJk2DbFdBIVr/T5ikgbGQfPTsUpU+mbuskW
YjyNIg5qXpaAIEaVURRHUjCr3rSlQrl4HNiJJUTTrxW6XqBYd12uJKNc9gPW
1HXO0VfCjCXF6ieeju3gH3lWBSJOTee6ri336VzVZgJ7gfe3EN6ADSAPoH3m
wUrY6lJC+9LiGc+nasPQG39LKvGCJ9QLc3CbLVFFkeaZwqqYqBCFwIphUk2F
Eba/4spLEuYxuh2ev04DocJJpX+UPfG05Nkg6Vkps3ASEG6BHKE1oCcoFSyL
km2y0H92NPeiZSWxyyAxJhh9fHFv1Tt8XqpKQNIx4BLGgEHFqpGAV/fUpUjV
kCDfEVVjCBU2Vlof7XW4whzXSHqpR8/o/GCfvh4lSmekpfBBLWmVDIk6hyZ/
NcVPF4aWgnWd2BXO78pGXK/4ixRvobzUsQEPZi/d+2Q7lLGFv1/h82eLPCvf
aI+yHC4KTuLf+aWHMEdCtBsAJoWzD78+qpA1EPwekkIhIWcgJsxvmn0hwjdI
iKn6KApZXDJx8R4Ae8tET2/vDvw55mTYkUTNoGvP/HdngViXaSISjeCf5Dzo
+9/o7ruXS6Lvqx+FIXA7mtdRr45KC9tjolLjzsGPL/CIQaPyY1CmxC2PFs+T
bAcxkI3zLQeYcI/y/5E6D4xW9rpmIM6B4PQsyQ1mesOZU0d0Sq/Jfid4yzES
MVDNAN8mjgfEkTrLIYgR5/jKT2qmZCGCTaF393E8P1ebVagWkB6YL1zd+Fh3
3ZYVYRjkFLR/YNDCUuqT6yhtYDRFcC06rvfpA6YxcTTPgRozOrVg3l6YGsmm
5wsO/pkIMEwm1g0HbBk5Vr8aTGGi8hYD+jzWj4sQthFuTL5kjU+1LoNklffw
+MxxHISQs3oNSP4eyNwsjsFmE+uSfLfuCrDpcBsXEeuO+RE+vZ2kzdSZrbMk
UdtN4UIUzerIR4wyHjtjWxJ0IyTENzrLtcDm+r8RWL8h3ZajqiYOenJUMp0+
+i/E3w0MaPUGjJgjQ6K5bQuSlayRpnBwKDprssERZI+W2ffDi3ymfV+ZFu52
fwA1jkZeGXCE6A15gN6X+WSAeJPwo+/bX7Xc+Dpgt3Rvd5DDopJ24UqLKtVd
8oIIz06isG9FwUWs+GP0//5L9Uz/sMvk7BqvvTkzl1Cl2AVKbhnvktlX5DRz
ydCH8Kka10qC8VjIw0YP8RRXMYHsPWaAck0GJ0SoUvv2vG4sxOk7+ORosGpB
Fc6KbeA/SQhK77kpGKEmd0FGGK2WuvCAzdv1BxzWoOD3OFIA0th+3f5qkGS+
ZfRUAU1HNCXuW7kryVkllBs5WuV8Wq0ix4Oenm0tgg0V+pMG6UGzzkeKKPX+
B1rJtC0jQcxOsF4SP1IhO9S6lgYukgNTHnRrlhLKD+0GLnsbCUheg81OgePO
j5SbKwPSxfdmNY1sdvdBVK4lUG4R9hp6k1E7KVRfWjCNRdFj2L9+1EBWFODP
Sc0SJZUEPFQXDlpMAJG3kKIfFitgXCS88mh5JNWc3IKkfMTMKmUR4BuojDyG
z7tvXDLgJ1WljgIlmBdiJooHgQirEQ3zM4Z8n4vhgFyDrEy/i2q7hhfeDmfK
6Oe2RNT6/FlSIQ3Yuylu1w/VcDdvNp5GAIiAz4PpRVUk9WVn9B9Vv+qgF72X
R8Pk/+B7tiq24QM7M6c7VnSvEsYDY2Eam/eihLiUJH41HWkoyNZ8LIrfsVZi
lEvMAJMU+wBkvtZ8s0Ah7AeW/GYfVi81W7GMVd3xcFFED9ptqbCZ9B85V/Nm
1WK1ojaJEpQB7kuu0NjEFLO2/6cWRGZM1vFslTkL3YvS1g8NeuGaDh5NtOn4
el8bQkV9SINum2awraDLPIcnlFZUO9cuOhx4jUQZxsv9+3GXkvzgsnPpMLkW
EisgHDjJ0MNgyzo9+2gx2nWz217KoMEVbXXsTeg9jFx7BvUGzpMI32Cr/LZI
a/TUyIIsMX0+S58Tlq9hBm0aiKpUcpc+WzxH3BnsUASJIJyQHouSMd+z+WX7
yGTg4xU9bKaq3PlyGH0BCDmY7gAcdqNh4IzNlXWQBY7GF1TZ3NKpw4AcR3TF
rk3dO3H+k3mJCM5OSSDwXjEL7ScuC643iXQQ0ZEG8WnlttHlgDQ3Cq2dzkWi
Y0fUN4SDYliCXR4olmG+qU8FmxtJC/RrXz/KM+2KmMAJCR2g7mWBiVQX6XbY
0d60orIaaM7xO1/pVn8jYJo4EghwfC5dq77EdGs6+N2ypM5kocI/jfWNfWRR
xwJmZw+GT1fnsFjh4MCdKTFSUD5KMOg7G8+QXbgfKQEtk/TIVK6/POsvC+yw
IA5EpGVX8/ZnZbFpEvDewD+WXZe/qQop0YXLbjdpheKqQuas9ujwWF7pBlXH
wjt8kATFhOeemzSmKJ9qg/ig0O8NjipKrlE7r1ysSSFRWCwjDU6Eo4/HJqXJ
HrO7zXUzWBiwMvlWgCX3Cj5+xoL1efVke5jBfVr7Jmkkq127VbyZQ1CuIbFZ
+ntc9fYHQfbx/oEGL+acZPFCvkGRjZR6zP92A01U4jmyJp0mdRA12LxQmFmu
MBw1OlCHsj5132Wh8V7wL3aNZRpJekfnSa9Fjk9h6lmiUd8r0tNmYcm4NH7Y
/n1kZyzeRGZVjvNe+jIdpMkuS75V6qD95yOW5e5d/n14lUv3SWVh0apE7olD
b0kfQ8wfzDSnZLSM603cLomDmii8xOPJJ0uXcTS09dv8b8lcEwUuGnCLsKnL
ozs+3d7S7DwI1SxWB0160B78qBIbA5Cs8J3uFXOQG4YBD8RcPPl9gnURpzKl
xeVoMFsJomK+Os/2zwC9ySrwrKYMsPPaT0rKgBre5Dqxt5YVeWWkbhAcFDN2
eioSE9Y37UVVx32PUQgy5sGGz5olwmDD0LKhz3PadWwS/UOHkNhxkopB3QpU
Gy7ZeRkE83TES2NEdA8Jm3HNCdRoQ91hZW26jBBFo7lsGPD2srpWN9OU4e1t
Xg0oDYqGayuMnkvCwkvCilnH+aYl4PXG8oU64rvRAP8PEeY24FOh87TqUmh9
M9aTCkAz9/3zfbJOP+7ILsPov650Uz2v0HQjOosOBtL43klAxmJ1AqZGHHON
7X+8shh2I2MWukR8po4zxq3RotX6kxPxMXjA0B4whYp6BcjNq41xeigm9E87
zWmGbCIuTEy8phUj9VYyZcTed2SPJ//P8d5DU9/caiqM+7pA+J3AnLYsvQDR
1QOewYGe/yQh0or1hWF0FpJYQEzJcZD2+PbO9O5qYosy5xGD/UdOLuTF8WZ2
82bfEI6Gtk6f2cla1MVdRD1kLg6MZtgSbY2gBS+diPLI31p+OPLImvdk0hlU
86+HS8cuLd2ioa5H0JG/6SmLnB8BF2qo0zl6r05cn/hYMLWbFhI2bmKDCpVs
MieNdcviBBYCAuBfDTU06V8JLADE3gLa4LZ0MzK6DwgizZ+7EtZiwKffIKcf
dX/cOTyrm7kXtv8XRfcGRhNoFQmpliRmgFyn8JZ8sOp8L8s8hk5BjZsu3oP+
7CRB2uEZ6o+e3njbPKENYdCBv/klwQQgvONnEzRC2dAmoTyRWHJ7YIzz/FzT
ndbObsYkZHxriorYtGIylorZpkXpIpFaTqM8i8BtWkzkQMcKfGW9zXXnyTUm
b075MXmPipwXw3islesMebXGdm8gWJQaw9zpR+SDFv7SVUra872suocl3fM+
M3puPV2+EEVjElw20vBdye9OFKy56u5AIIQdlB6OmEsJsLyZviDvGaFyOksW
Hei/zcQafokUI1gyp66G4rcjDnOVrguHYkwEGoRWlrVqbYXiDFahaJjjZa2M
z9jBxgb06X516/HTOY2tDGysbfP8EYlNyUkGbOypI9Cy+mASLPchyxw66k9/
7MsG/ywNSmT93X/ScXNqVLOySQcIWdx+yuiUGuB/bncCx0U8mgw1RBYd+nUd
HGtUYy3r1YMyByaPEk7EuG7qxo9qR941FmQcm0sXkXg8dGsGN/T01+gmGgrm
3TFgKQfRZPl0yntJ49WiMapPB/qfQ9mi6bqRAFEsKTT4N+0jL4YfnW5ovFUb
RO3HkrGXqahYfUFTA7dQw3awTq8SUdOlE8VY5E4CpMafKK2S3YfGMUQWI5yr
G+2cssG/wV3uQcugn28agtY04C7VzBZKZEYn3pfk/Im+z0+rWzKvKNy5XLEN
9YUv2GzfvZmG1feAFekh6aJxoWoitF6mMqWZZDuf/zdtYDsmeMFrqUyrDsOl
u91cmxYCdl34p3ni+AuA8C0kpXasZf16/dLO27Zoy+A0AqPuoOff6DJMBd3d
11LSxu+UwxsrButBWKNrlecqCgPwgU3QEYHTw+tHtkc0JmE+FOQO7fD/DucT
xw+MNCJQJNw1BCngx6PKhTXWuqudfVUuhEu3oTMfP+IicJnFC6ZmjnNzcvYx
2DsTVFWyhkIku9vEbJh6/o22cE6+U+m+ldI1YUGdpqJgC/tJ2CcVtN8MFE5N
UectAXm4ZfVL4M2bwfBU8fJBHqYmy0AyHqNy/F7TMauB7fdHCzWYN1FZq0hR
c/Cczb7sbTTc4lhiJgJU2cEmw/zkAIm0TFeGc0GqLzG5PxpnGBWxiZqYA6U0
63VYGhvWKTNt7+ykg06RYMCqOFG8m0l1GkquVsFcGfNu2rB/LFB15tN4nwoa
sYytET5OZjUaaT+HrFNNRAda10wuTO3Jus06DY19+a/0rloIhcIYlu1p4lOO
mMyWKenzWOIFGMRP1bbtFGDbK5sSUudsH0c4gd5VNUq2hYbfhJOwAnA3R0bc
dXVeyYzmo9r5Az4LvjnvvdUk/ihlJV8FIxD917yUmn8iqyCZNPgOgD6HpplA
1dTuMJV2ZQpGNZlz5WNXFXYrg1f8Cyi2NEXhn0BkQw4sLVEsqxZZVl/IywGq
wuIEFrUnMmV0IBqWEzC/LAvI5NS+q8GjsMgLEr7WFgYTCRKjb7XfH4o/mrYg
xKCpn8GOuV5E8GxdWr6U7NtpQhuF8PeqQ+2+xQa3rvZeJnxQRykL4a9OwDSO
Fes0VhInm3Km3K6CIoiZY/55ekBWahUYmtH4YZFu4ynFnjAxjj5ntsmxsbYn
vlWUa6xaVRJWceuGp6MlelfwAWJX5TpQJuOgu4H/EVrgwe0kkqTbcFWqKN9l
X5pRl20OjDcIdDQecK+JCNLoGkne2HYgrnMt/Q2XGFLs4qgs2ItTh+DHvOQY
8hMENVuefqzQpZHipM2/6DbMBHir4ri/wbht1tKCTL7HguIVa1C0LyzpFrdG
/MwSBgsOd9XJnSm0ydMgtKbSZBeciPKP/EbYB0fAJcB27sRssFCHEmK//3RK
UAKNcCERvHrgBTjdneeg50FBYXodLGiR8dApzVEu1dGEuC8AhdJEcKX16pUy
M9IM0H0OG9ro91xUK5YkOQZvzcgkVxC1HGd/67r3XRBgd9RV4heuwX6MUrwQ
lpSQ8Yca1b7fJcsclpTMFfVAd+4hsWSNxzGwpVFUb9Tns+yKwKFM6q986W2K
moqv2hkwetPucbIDXLhuMLDaN38BP0Pp2i8ZwJSbdSH4UGhZhI+8Fh2frTQn
gomvm1wNayvo+y2+e+KBQu44ZjkmaqkXbJtD9OEM3rYYPRXFShM9Eqls8hRD
CUsaMLRv6bNLavRO8yia6iKNne4br3XV2FAs4HmUFdmbu6hPFGsb1BgnTH6+
ofR1UNQAMPzA8XWsXsXmQ1zN5FfTLorV/I9qipIDCY/L07Hd1TeMN+oOnsH+
3/gwJDUBTt6lTunX3u0gcEYPxKliBA9GCt5nbXHHsKcZO3PVbjk8kmq5c/Mp
CJHV9q/goAh4JQMtKh4welMKf0RYgWCjTBI8vb+Hpo6Ec/Nldxkp/Ad2gt1l
HnEMqNGQCQq2osXxN3gTLn69qFWUCCY7s067f5k2P6HetFoub1x8Q1uxra9v
3o7jUu1hAukfmd7oAsvl+OptOeZol+Y9XwDrqmOakRPqEYcvKeYAGrv+9BTU
iBm9J28CAMYZl6pBQ9UVGg5CQ9cTD6FjlRYzdpjiH/SPcx/lcQJmBfKWxWAA
4CPpY7rKPhV3I3C/QmkwfYA9BKcus/hok9ChpI1i/mS7D3OUj5pN8Rhnjuuu
EoaHYIWs0XvtvC/xR04PyZOZFWevefMdbP7WInimo7nH1oho/3Wt/rLyAX6w
3fTx4ovYW/GzpgE3i1/pubW9MeO9VD0KCSNg2paLYJ0wGp6NtsIIY1lBNGys
N8u6Yf5ANCnntIeUxwIPRMEEScdb00c2Hk2ZJhkaha6/+zqt+UdHYYCW5CSl
IFHsMPZtOqUJ3pJ+0u4QNKloqOBm5nykPfQgYlKg1thL7zxuNHGW5wvGVW9B
d+TeQMtN2L7e4DYw/6sQ8xXFxRQaETfYPzwjcq3WTp7NK+zHEd1V+gK4O0hO
eCFhY5jdSrgIgKrFKBOdHUt/dj15WGZYqJ12BK66/xkbWAy4xgR3Qq9OsjH+
KKxENg1eydsjkZ0xQIWIppJmPT8c8etn0D2H7rOiZiydxWo+yNF7owBHnJj/
9rd59eH/Nc24FVum0/MGPVH4Y7qk52o/sy8J2Swd3ct9uzT9439ZUvbI5Ery
qsdti5tviBJeXLYz2swdE+GD3tv7bpHktTn+rR+UE1wN+OKbTyRqI7Z8hmSu
4W1pHDQE5v26E6LUKjyYEQFVdtlyGaOBsHd+PqCIo/aOIrVyUGkf0W+18cBI
++eK+AB0yp0wUckzwiZgrvVZseO0AcEsLfpMLCpX2J31ZS35/mXqEnFfZdYP
VqM228Yjt1JE0CZuIxIPdV87mjQs4Zu0etFRrwQ+akm9GDNCI3o7U4slVTna
VqBPbnqY2Z+0llm0PcDqsrfpDFroofkG/X2UVLubD+PtQOQbguzsFbkfZF2v
uQJ6FSkLJfZ9iLopMmEclbaeDAUDaaJMG1BsDVRsdscDgskCOd879F/qnsR4
aXaWLiaB7MBTmDfcwy4gAtTHF+FkwVw6jUr8f/D6x7mcKn7mcHG0JZgmyzmB
DU5qD3Ukw51hPW2dHmwS/xO0212Ef1UtpL6QV6uAZW6/apVZCeAYWychqrC9
FG1sUsp6kOgWbN3yj9mhYpjvFrAw/zY5afwXgNoWHLrRN4pWmEacVoeUCdYt
u6RdoHczzA+BRNzUPiQVZg+vq+q1Z+bHpnxlE6+uCOMyFdN1tZoysRTsfbWU
KVMNRlKUXtcqhkC3G7KE7fqE5oLOqbxh+PKdf2A4Vr9ezo2dX2Wp0DdRYCu2
g96h6BZ2DJd3rrnKW/ic5EQykNOFJZUNRa6qVk7W4pP6W/dY/RaMYV1TE5cO
rCQBum1sJ/WhPDg11/DTkJxMSWsze9/imOcfLhyoJydYH94T2FjJfurGL/Et
PhWQt9gh7s3i+P1z3PAp8UX966TYvFjpjFlGmXxVReAxf/Hk2cOE0wYhx+pw
XmkPPr0Ov8vHOe/RxcwH0mPowlCaW500JlUMoawXJfcEM1tCjdBO0dRNM7EA
uoNB8DDzOSRa6YFeukD0wKYz7aAYfFHb+XbYWuLZAaTk6LLtk4Y72aMr9YoG
BEbVEEaDSBWDonMwzIy64Zj9xfaTiX9NQXWAZoX3JTYGaLbPmM873FeVojjA
DEzwCnESLOQ1TnLeSXYu3ddZ4j8MCPnJoMK4Vuu6tQpUZr9alax153j9OCQc
K2u2Nad1EyFx8eBNPJPtnvBhuU9aVIRGZRN3Ewlj2rS814hADTMTBV70V3b6
N6VzyyRWY6IvvYhgXirb5JWVZL2iSy/V3woZkioBcGgR6ODZproGOXBaeN2o
tTub1wdTWbvTq7MKyI3coP3RehY96W6ee/Jt1RHl1GA09uQ4ATsu+FYKYdto
r4jRjJvqwq2T5q3yA+byuW5lnttGsi2nAtu/VdnCc/s62RIAEc4Yyh1BmZib
NXvuM3m3l4sX6yU5eBbS70kkosCiOA93RFzypxli28bS++7ptS6tiA2XFO6m
LUIgb/9Ydi7AaOqjL/JDOaQu4fukYNhq/lp8O5bDgVJnGJGSZBaPmHrVJtLS
HIAInbO99DzbFq3B7wSL6es1nMKLDulYG+FuzUDzYyOe4K5z4tg4ZliFARba
4ZZikAzUMXMzJ8B6KUfA5uFlAeEOJIZ3jqnqMFg2AR2RfVhJE1QXJtPULtIT
M+LkvofbNaqiWOaqqQKZMvW1XYqSxlersB9G80FJLP+EcBWewHsGUWN95wdY
iMou/bLXzzw1f9YjQEQ8MdF9PV+tw0+kSc48cgCs91oKnq15z/sWOcKh8le5
B8jmQRb0Qx41nyR8x5sBiWiX7im38fIUCRgOi8TH2GJo0r4LbRkhP4CND2yw
Tih9FQXXnvMX/dxJ7YC1mSIjcsMaYEfV29w1aK1kTpldETieEPfXnoxEV6DM
VI8+NvDTa88rgvOXe/IO+Pt2TIiSWrkUrYCxyOzfp69FU+DM8v8kn9MCEN9V
GvYK8YlP6PAtiNJgsgsHSgjXtmGtXPQPm1FOo4fMuH/tbI6J7O5QmKO8jHdn
xcwKUuTEMyIcfEyhtkDgxxcXanMlQ6vkasPsPFe+hso7sIl/b4JcAmjVPBs+
fOr6VCAAQUhdROmRFc5oiPb/STrfy8n8obJZx21TZQhiU94Cx8I3S+sCYp/I
H0VemIqvjuWWLwndo7wzmYRfbfr3eTzQwJWrQ2cfhghE1ajsEM836R+Dbr4q
xwN7UVlHGe6wT1qLJ4HMfGXVTYBOQzVhWi7I1NIeV2vi4k1Vj0l8wKf0rhpX
z4eWqYimaF8QQH+VJJz5glVG0OeV/FenQZMpi8nI0oqdZf/QwNbDwUsaw0+U
9XFwDlzP23rKLhSvQ/mYHRGRtxJp47MqtJhUGp3R+geX2IUZP3QRCkuDPEEH
78TJQ1qKelMOElxHfGH8vToQqkwmZXe2tNfBJbmPb/SyMIMGWJ26BFUOUYLx
7SM6y0SnGn6owg7qgmP2osENsUomr+ffFL5RYdMBKivPeiSHeXUkvnmBNfOC
spjejlOjqucsYqbhsqJX9YZq2SFMx5+3VfK9rFmcx2mBX76x95FQG01ZLK4A
sGMVuZSTIY2P2GNRkJM+JV6RGLWYT1e0pAOKQiEbP9TC6VMJgiVFfjwz4r4D
rV5satGTwCUP026o8wIrbO7CtO5AgFwvq4uJ1k9/gxMTJ9FNydLoRaK9hj83
+JRcUxkEDpJvQoG5alxTkPjVQKrXqElGN8uQHfmmSxIpZQUY/qFylvJUq7pQ
/cN4So9RvUGoHmtTFepioKRny6VCchb2Hxzvh6OCfjb2RoUg6tuiLWdcikuD
nXmTl4VaT1J4f40H9w2fgkxYU/YDq/VueI8+CSfyX94BUZoC7n4oqyyW5a/1
vsOv70pXu9bjXUPGXJmjb1PQcpVq+c0dgQzVan7zqMM4qftSCIHGaZNAqI9N
9Wssb0LtM0a+NA0IFi6M2sR1OCSqI+pR5QqvMFqcUmXEJhwLpkAUcfobtKuP
jQf3WaB0hxYbwSuvHX3PI0T4R/jw+/ZJux4KXh4v9xFzyhkokyCCey91uo88
Tph6KDiv2c+qeyAfT+YfGyWIySJaacV0Tct7aC92UdQ2ZHP1Z756nd2jyGoO
V8z6LInRvKlXzADSKXNyMtxkqe6MWXgAAeFmuBb6JrxD3GHbxzAn4UG8n7z0
Jht/qQiIsyPFyu6vl5xUHR6IRhON4izFRFhvgJujX1ScwmKh8bos/Rqj+qIQ
83DNBMAsXKjls/Fe7qFAGHBTbTDHBtxeFqqB4KEPXjowrvdxjDPZegrLNPvF
wlkBKWJUrm7EySV7lYeS5n+z5CP2FQTdx2QRDzNqeZ0/gq0b3B1JHUgk6Gxd
M0nSygj2EHEv6+7ds8GgHI+inmsXZgbiPdPHXBX+m/8FWd0LMaSe7U8VHZnn
XHtaBgmFcLGU5WntiOfdu1vtbX0f2KYMxx/WuO6nxbd/RmKSz728gS4Usff8
I7utw66mkQPSJ+IcuWbR2MEy15TFaYYGabsotwG4jVto+zOVXJHdiR+9OvR1
6JN74nHW9gRHnQlddFNNmNJ8iUHzAfK3rO8FSaX3YDTKW7bJakXeggRtWeuP
MFStzvjNKUvG8Yx3BCilaB1bb4h5QVmVrptxUPMlL67Xlz96Isqg7Me7SP7u
x1JAUX4b2Yr9VzNkNX7U/jkaaGEkp4rVaqlSJC86RpRur2YB6iW36Sw/JEkX
/TwoBc39OMhmz31c+henri7TQOgYt5BnQ0fnE80KppOHQ9+2cROR8Loc+YAE
dp2VbbWxgE7F2ofRsTpYbw1FgJjjlpDU34vFQQGwcKiNoHCQCM/zyn1x8kx2
IZv/rfL1ESIASRNkUdxgT4pHM1hxFHlqbOVj39+nL+HKeAcE8roYZGxMkZfN
nd4vT6VCbYK58+2qG+vdrS+58sq+x6Ri3o78zWBFSvAMRbmgTLI8a8E3ytdZ
MzU/N9You6nzNPHZgJypk5NSXF5n6V3SD1rQfNOKYV8v8n037wR1MsH+URGw
3NsPZIey76TPmEwfpKr4vvO9IGqVpnFCsIiSDgOdKYwLsx1eecaJ0ucuTYz8
C/xAG2pImfOBIZJejAY0+CacU7S3wFzMChL4yx7AlJK7L3gXHzhEb5/cSLj2
hTg74UsZEN8pjIlnR4xv4yVMZj9n9f6fW7y5ODusZ8zabnktAU2YP9zdG7J9
HtrXS81wKASemP2kW3JC3Zi5SHRU4W/y+02tdJCfdIZllZzaTrnOmem38Rya
RWQ8itdUNKEvxqkAFDeKR3jXU+s6yBzhpNtNZvNK2dQb8MdJJH/llHsQ74rE
HC7SZ6gDS71YShmweaofPF3NnaEeNs+QDTNQc0UjzWc4w4gRtR5ggBCXVqP7
8WYFgIsM2frFoFR1Chu93EannT/6p0PBOjvlPbefS0WVYORi5bJdOMfe2fum
WfMhINlYofcW36w+vVp0YjcHkg0+nOfx24qDe+ECclHt25vaEcZGFrzpMPSL
oE0v7loJkaGPQK1JY3Uhq6D7k0AztdeTtJYDzxh6VFRMjHzQBKR+6nDUmxcS
4D6SAaYb3zdQIHj7FBqDyD2OJtjLIl5j8hwzVVXZbfKH+wuoZlUTzaaU7Sme
Lg2i7LDK6U6OshSe1Yv8Fw65k9j8exxNObUEd7y1pQVYc/NBzT/liFWJXtM6
oitNKvyk1ri7Lul+4ouUz5Y64sEC5NDR1wddfs8cln4wHINktroKdQmwuc/I
lIDq0cdKgNCZUgGyyBM02hDGf5Q+CFrKeRAEaOwprTGDOfjuTDuCs0A72tXz
u48YY+o/GYllhfIR38iGnv+McRh3qF0WByaUa+p29hg10E+5kQose+bVLSJf
4U27Q2XKmR2w798Za8GTsUYP7ph/j5Ps67ch4Spp5r2rOMDtaI69Vipn6pPG
I/tExmb6Gob7v7L93vE17CcHMnoayJA3a7dRwqzQBhpBbPfRo/xnwqP5KUaF
i7drdCxYRmmZYrQuvjaisn8RK+AoS6t0+6YqKNpZlOjipPvWmw9euBvrrSv9
VqiBF80toKya+aVHRGtW21IpDxw8C0yINQGRtsADEzbvxScaSOyl6QDhbMav
kql+SwQ7HUIHIbn3GxW0gwu1Nqpimo29N4d1rclr1rHfX5B8/2Csb9WnUFCL
rFBr/hwMrmr/u4rmWI7yllpIzu0BOpNqwNaaqE+zWJm87lGQtPbUIFDHTe5E
d0jJLYRqfSZ5e9lH/nLMp0Sm4hawS8m+kuEjzpzQ+sZ9F9zO8M0rsQvCxZFW
dPR1U7dj/o1bgrgwv5xWuJvCJZG4Wt1bt1jfEYsGKpuiGf9EHBXLngMGzcQd
sC3NJ9KPiWFQy1yQ7cwdRWOupGUaHf3d+mIWr325OlxGdtZWz+Vu6+VAJ92h
hI2DCjZXqIddtYjja8yyjkbbk3QVfruefcaAyg8TLgwmK6tpxJnc8EqPaK1T
5XzgUnV3G/z7YcNlP7kqlXW+J9e9ta5nInQ6+fcHPguBDYAzKSDinY+zFgIb
XJIR+5qnGuLf9kHhhJE7FuI1zaVFzDLOXsCjpb4AYHNrM8/kVkGqyNVY0s19
l+SSf1SnW08xMoFkDLITmSyyxLKGu5WP0orGQ/GUK7xXyANb+m4meE+3qPgs
+crZFbTji6D47gftyNqyMOUHh7zfTwra8sHBEEqtaS3Ag0Q2p2diuGYSoDss
AJzw7/y+VXChBR9pQQ8cHrdJ5a81l977DmqPsDx3gK29l025tyOJwivbohqq
GKrwgbbvXe31l5i8dJBuHrZZIDR0uob8DV7gIo/u8fjrJoHy+rtpki1DbzNI
unCZip+wLuExrx+n50nhTY7W0SCfMSAeQpv9nPFw8WaefAKfdHhEnqKqFJkt
b6qg8ti0xpRm8+Z6WD+ZY1jvD0vE2powZd3ZqXZTsSDdSdrousYUk30HTtzY
pbWp7Z8e2B7SIkw1KXFXSpB+LHGtFQfYViiYmxce5B2HPnyFgOyJs+TLYyHy
metbCzzs4dWg1t8gZA0zSGNg0t230g8p96BZhaNS5psakgpkkV3Ans4qoYSs
paK01FBP5D2HiBmdWcUSSqILI3/13d226cNXlQhSJHFjb9Sbu0GLlIcKvjjB
KEJVgMdh5vFv3xEIjbTLpKsl48PiLwTpQa3zcp9s+GQ8VSTjFOIcjtMlbwmL
jN9eEJnThJV2Co+6FcKb1l8/wagIXM1bX+BfacmhZlpuGV4gEIhQMG2KLO++
UXca2Dtui5PmCBK5eOzqHN9hXeORv7kWyat70vH68QqXbQ0OZ6dN6sUITo0Z
7kYymz61RMIgkx0AiwaN75h5tiwQWGxzChiS4jZjDTxXWqdV5KM2ftlE4rwf
Mn1l8ox98JG/5hqrT5SDW0vO9q/O0LcRI5tOn7o24+hoRLUpFEiYrsFvMkpx
PJ7IYYjLExvuFugglbKrB3PkiR9uKs7sAt9X1d5FwGhcKVEKMNqPU7lNCoX0
H6LBN+a2JhJvaSUepZEYqNNiS556S7i1kksoNotsOQu/+7CWoT4m1l2YWqXd
ZMZDQfu/COlFFltLQvtazINH/4+B7PxqW+GdL8006e3ULMWN+QUG/3NcDJib
5+RT6rL0AXcJqpdB4oVru/mcQgK4TIdnWpboikJpAW7dY7CMZPScIGKTwxBl
VLPL8GsMuDmAY+i7mPkg4poW4kjw5jkU9bviLcQ+R4rsy/sFkPlrF6E89/6f
VZ/H28xSUW8EkQQZZDfrxhSEtH4rOBbYyTRkYOJGPVHQswx87JakTZF8ETx4
KcDVmiaoiaqWkR2LrBKlwbeERApxtEAyM2RWmKvp7DOfFunuxaY4Nxxrcx6C
Vgg8Q6UgJwBbFtQO5RqMwUoY301/D0ICwe2cAvZhhfSdr5/ZNyNaM5YZSwHx
/It9QEl1ZybE5DbpT+i+n1DhIGRQvjGVUPxMMZXf+rh9DbvkpkTlzm0nRyM+
ohvZ/z0Fh85HWdvAtoLBecB73GYJxUnAyT4zyLVbv8CqTm6YetzgNv31KlXi
pCejYvXuPYYv1Rz/8KVinRzcAdJpDw+IqH4tZVYXKctD9XeB1pWrFo2TW6S6
fN/sMufJrSRFME45Zxs9E/UVdVCZ9udfb6iWTFLPnfamEfOXERJ68RX43ycT
dqScSwlCKW5Gji8l48SsFU1ypID+aPEEmXfZhiQlXX6uG2ghfJOSYww3lQmJ
CsbNnlhgGcjGlyYyo2iXI8+UKNjzy89LxUmHXabJQQz+kxKCxB8dq1H9zQbp
SP4f03jz2Ti3QwCdxwFRUZoDfXDl5qP01CrlUEGbOcpFdBh0Ntn+bye25K1h
OTDlSYOq7sP7QsZmkOvC+fLl+Q0nkTD7Wpd7Kf7VDsKzPnrSPK9WOz3qORsi
mfcU92CkPJVPV7CBR7WBc74/1NcpxHcvpMfuLPL1uLmJ9Z5XUzMn3nhTmlEP
CZLkq442TF9sNWkzktvQAJw/VyfguwHm+pXGZoWGAcg6X0WlQFbvqT0EIV+4
cJ62WplBmXKhu1ByM1xVTr03kA5dKlTDj7fARxZEupThCf+hdAOqUIgZ3LwZ
cpY4koA+Yvynl90sMszYatIv9v2EPm/qAjSpA23CbC5E0LlOmrptws6tTdoi
RR9etBvkhJ47rclirWXZGJhRYiDFR/e8jUBR6VnNor1qmFjTrWfc0zfKwSKY
usn23YeJeRkstVw7u/gEWnPEoaUsm0INBpVI9OTN42ymkVDdFdn8MknvV0sv
VCQZVaIfXuLaoPe9AdJ01x60Pbc9ub6oMT+kpjuJ3ipGB8zz3GbbHYWju8v/
qG/7EAr/uhjv9gElLlGbEXUykslWON2GH/vitZ14dtWeAWvdkCAIDMcZM/Q0
HIpH6TC6HP4Y8sYX+Lb563pa7nRJpVaWiCvRT5KAIAvy3k1GTGw8sts+0gh2
FzOJzVH5JY3eqPMPOVzka9+y49JI7GXyQGAx2THX34Wld+znMieN+A7seOox
Mqekl+9HV3+unUY1DhjbuggDHLQ4OYlfrN6rDeTepy6fRXtMnjelilcaWiuV
zisoYTfQBxQ6u1hQhER/K8irOU/vZfieIekphQpp2PyzV4kO3iW5rlzg/gjY
gvE1rs04p8yo0jk30kVO8U2+zdC+1rZOYligDZ4aZDFFGMuuvmutQDc4I905
GDNy14bRlftbecm5s0PICMs+ypbTN+Fo1R8Q4IEMIbvX5nbbAYNwScD1n2KL
Q52wGJSPWI/iCHYjAUiG7lKs4LmLXN55r0WwYbJo/O8wqeMhOyCVDXN9zjzu
5GDns8O5Ety6rlMe6cp3AwizoRW/qZpJv3pnjDpRDOu0ql55zPl/hyaHk7Yt
xKx1EKG+ptiCyK8bSgqyy0d3R5qMRK/wXr1wfTEF0V3igGw+tw20ghnl1e+T
I1XcXlZHrI/p3eIwJf/SDhhm9BN3ODaHGQBtAk+QwRveKVwSZ8JY6xM30Fl2
JutLlow/L+CCnMGLAlz5jhwtcCdHi4Sa33LgxQCm/+IL7K4qJAHhZto6R+jJ
WQ5468Cc27JIw7sy12VY6X7/AF7TdkcQneh6T7atYyBGuG58PVGD/cTUPi+r
HmxPL+UvCnJflBHqQ3m5pcTOFy25Z06MKNfGqbD8DEC5DSxMaPWE+fTEtKBt
Z3Gdcvtaf5bksj57k3skh45zi5O41NZgWg2xSi/2ZzxohMT29EPl0SroIBEk
+ZjXF/e3v4EeKrVJ4MJ8MlxUZSTPde5RW+r0KDmbTAF9SN5Gw0dCKo8sMsQy
COl++Q3bKlXc3WMNigA942cWYRGyrP1nj6UKMYKHjNwYM1YiVEbShKrPgDaX
DVb3g3QjMvUd8s3P03DpzT4xgsM2fVFUBtyHYeAZSDQXWEKKacF5Jy/rRv5C
ypQEdTriS1Tj0RJpzaLLZc1v5WxGFxkr8ko1qCzzMOr10fNbmVo0nUykuPz/
H7AdjlcobbT8bZRfP0zZGiTey58Yp+fjHmn/lM4YaSKRluc/OSg4DsXU4hp6
fMKNd+ijBfGevBQfO5/7mTvgt1VG/Al8OaTo2xgfHmlH8ZMZbzc4i14VAh2L
gydU9cSOHD/uBRJqtt005lxR2lUlV9AMa5AEkYTLsrF28SGvIzeRwkcKR0v+
dqyMPhx8rH3jM2HdQfmNJz8aYz6hq4cAwi9VlTVP28Fm+mKnXMC40zX/GcoY
zEM50Mrf6aSXR9qWqdTkpfjuA+qmN64POn0pbdKIb58bLywzb/EFsdkk3xRI
iE/rOaciDYYzeBMVM1kBZXjrErNZcC0VEXOyyJIEDD3WCc5es05uZFS4z8R3
Mk3ELOaCIyVGg83A0PLkv3HMCljYQddA9XtPtfmiYyx/qO6bXyc6/kd4wuVx
McLZVt9ny55BKoGkF2h2/eAQq7Zt0lA50ei68LaH6kQ4V9hfc0+tr5t1TptV
sqXQ+/v5h8kWznNsYI9nxr0DNzcYYVs7eFz8/UYhmkpFRKtJ1Ibju06+J0H/
Ajc/JqaZjICnScVL3XY2Ov7MgnW1zdlMugqtO6ZUzGauttFQebpXl8Jrfd8m
ZzxXao3TeAlDh6lFSQajq51FFoaOsuO8QaM0YWqk4MTealLw0WBA1Ri1kSOz
A1SNdz2RKmp9SBdH4yrd2+u9YN2L4ANr9NIE8a0etNu4FXHh+1PxyTDH/xi8
BR4xom7mzA7g5kZAn0q3qRIZMvchFUA5e7Zu5lMGsJ0u7ywNoQK/YAYv+B5G
Cvd48/O535AIzkpCxr+tnr0FxloJ1KSmVe4XcGAym0SSKw9K/5nS0xQsPZ4b
1XJ/uCtVMpxBMJRoqfiy7oCzJqA4QNsmVZwWAF4uG9OHT6BgyPqxAYVj1eZu
VkPOn+kjPgsA0EULNoqizYlNlyuAi2LM7gbE6Yf8AFR14nw7XxLezf2htmnK
OjnQ+/ovuJhYAZbCreN7SDG96hZSs9ABPbh4TnrPry956T6SictWVIxmGb+j
dsxK6tMY4exsSoYtEQw4Yb38x8QKyYvBecjir7LmyokyCF4Bg2Y0smt5phZh
uXVL3o2XxPNC+3ldVMWlrZEYragh+qS3LeCUqZ2uI9CvfDi4aXjyBOj47gQj
QNA5nysRMpy+2/M6dzCw5i3jIfz1+SS284Pfp4fIXn4KLrTjX/Siye5d/wz+
G/MBZDd25VgxuU4IgbP4fhbMSSB7QH9CaLk8CGWva0nmLoLRsRSICMCP5P6R
sVSTdIs0hVxuELdncVGct2cjBI7M/JAwdEsjGs2Sas/Ne4rx/QT4jMYo6pCq
fIhZRkBnr29vrnvDdpcls2BnOxAe2G8dk0uXTWyG38pvVWBkJMkCQCNgnRmw
rYn3AME1++p1MbHE+RBKd+YJ6L1wWlB6Gg/leV6nClCt9KByGt1Df1NMOYbg
jGehF++g9RL4jEZoq0n628P4pvcaO8En8NHhcXyW97eS/AQFTGU49RhudUxE
vuvuGnTJLxG/gnfk28AyESdGFQa+vfcBUZpaAEk/3d2MHe/EwDpWBTGDHlvn
1v3IhgQuLq1u+8wn6+mrDjyXTwU8TNTCJTeZpAlzeeWgpDxiLwWKPLX2BkB7
VRr/J1Vlbgd1qbu5v2oUGPkdrhB64lJSv0fKXZHCDVjCls8eZRWllu991B/l
4gjbOXMWr3/xxewE/RKR0pAUucwufBbYMzwPTqsv9sHMKJVuFQw3ZO1M+dA6
nzcSlLpsgDiZR/FdYxCy1oklaV9gltWaLQSABmiWUBGhtzGY08SDdx9nr2/8
FobjeM+i/21Yb824xvKYm8/R86QnQz59f2fH+6JXZ8z4+5boCS1tHsBRAKkz
OeNZsZfsi7gBsmp7pQfd4sErsfDlkhxX7GyR4Im4RS97JahSwZ8ZwFOyt9Nr
zxkHVgFWIHx7qJtITD/LtPXgOKUh3A0XkJL9gaF6jT8QBnHz9aorLdHoJ2m6
zDWrJ4UjjPtfof0nYw9CTIgNnLj7Me1rWRVFWxJFeavbbWgjNvE9QL4ysEny
jJ+GEtMpZkC42ylWUuTF2uZpt3pcEYqDYKqu5iixEQi11D4EAblc/1h/45ZU
WJx3WvusX3YuaekXs6PWvY1me59GfuthiOc5ZIecH/U5Bek4rThHf14elcri
FdWO9Pdl1S9YI7KPy2zaWMIjSyXYzAO+QqA2WpFRKZZ6Lg7XRADLGV2KnPST
GukAKsUACFJIG063z4UPp7bI5XQsp5UE3jvZQkSvb3hUjw5dVo0eFN/nE5YR
jkMG5/xapBwUGwgVl2/glRcXRKwRu7vu3ubyJt2go/xrBSZi3n9mbjm5usVz
QfanDt9LnEJ8/g6LmbRtu1L38xGGh5UivSyvuzwgs+cGu/L/zCBW2LguaHPp
yH7cxyL50+zE+2+qN7y88Om6kFWDLGu1cnnkZFUVKfES5R+LjUXS0O3cLTjd
Li0Ux+MUU7T1sq/uGWkWAPrNmS/dzDAhjKCXiE9fyauJpXL0FBOPkTw445rA
qcXBRQ2SyjO+g3qAKpSA8lT4Q78msK6nyuvATh4XAA5PS0Cg+tw0vtEWx16J
EVmbdqC5zfZcQB8vWdXQqjCWHIJn7SVO6qqWtoaMT42zThVUml4zASMT4CyG
oc8urDAlQxVEL3t9fJw6QfrurWmq+VRrsaBmetDNBqV2pV3CmS5rslUOW+aW
c84veLN7TIh7XyYHr5w4x4qO3mnSMbHiHSVqx0pzQqBVS9l2hHFfo9+Qtt3f
BqgheWQHy7IaDvIpDBqqltC07B/2DRvImm8MT5FW6nHu1jAY7r1bAooW0s57
/NlUkircLX8/WhdigS2Oyf98N1AVIhEB8mourTP+aRGIvO0AnjXyLjZl96u3
Uo6knHw15hh08sV/sg8A1sMdlMoUguVVLnNNZYKvckjB07GU+sBE6ZaO0GB5
OGFzsrEy4Z1nur/YxelVYS8w+hXUvjKiI0Y7TOKd8W0pFbMP8LRa8kJ+hiTt
lpJFpeDhXHi9czcPos1/jq9p2Yv4INKZd6wv+ZVWgs0t/NHS+5t76OWV9sUH
nZbluFYOXVPm5rpxme5Np5fi8UMJIwsLNEoDZYcv3f64EklIGBBuaOP6KVs1
rgS72O6f1fBQ4Fyrg52mjHd94O7Jd5WvNAeWGXMH/hLeDO89VFvjaUXTssCl
a6KHOyhJtNauUO38Ry0Q8cMDgtVbr198lzjcMEcAjhfKZi8k3D46E+BGJCh6
aGMH1oCo85Em+9D8q2ix97MNcL/E3p+T9mYqoJzcq6uscB5J0suV2m6ehvj+
ofAqEFVMxYxJMEi/P9058J//YEhxjsSiiP5yhjr/XXS4dW21OSCgFhzCjU3h
UUUOZksLx444WlKQ2IqyYrNCswY1pJxQbVqDKpp/e0kyUgWAUF1H/rzhxK5F
8e7xoG5JGu3H7KzmrjKpdqbqEU2Cndwet9rJpegx62TuJ6p09S6Zu778hF+P
7OqbDKaDt+8XFUOyQbb7zt55uC94inQXa5dzSioBzH03px+o3AdRYo3aDHI1
qFsJBrx7R8MQKvcJ4kRwoIDXwibz6KzmfXFLCX+/1hcTD6p9KJhL378NDn0H
bzdxB9twTnh/S35mRnDfCQsN2ORYBipW6mdHUIHrchqtBjJyOu5ZNmpm+HRJ
CAMlENWlcpCCiyuxj46ze5bXCqoJQ6POMRnOYp3mPvld2dxAEWJuNzSkQY6V
rgJSl2vdyq6xqxC3i6Rn+qCEZwE0shoDulwcg7BZvaQwFmiUzF1U/CRyVXaQ
tPmDn9RMkjOfyEW6f3Dtt44mxdRgkEtcux3AEUuuqmDCed2oRJnICtZlqoaM
FofgRbJTFleqxkT8nK8j/3u5+/MGZX61DdtY1UWQXnPQABH6O7eK+NnmZA0Y
C9/x/Kc0txMuXGw3pppzUeVAxzwSHLTeZ1ZqYSLDceTa301AoDnV3Ok9coPj
8I77V7jhzy05d7JaUwB0TFfzD6fdRsVic7z3HXodeR2IH2SjD/NPWsxHQr2C
SzndDPSA3iCo8C14Q00/9prbwpNIzBEmCpqZkRkf0717sQE8mba930O4buB7
NlYDutXMugImqNIcV1bj4K5hqVLuKueD/OsawJ/MWK6CGUh/mjnx2bYKSgqL
A1RZpxVqQXiSNCbH9HIi+6n/VFLg4V5j7KEARfejUEmfsRv75VOQPNfve+EI
/cLIo9z9r3wE0bFGZCX+91kn1rBC9zIkovKx8FkoOGmROToInRHZnFpXV97j
GPItwKyNWLkpizBTCjUwttkRYq7M/DluwtvLulze7Upq3dALuVLmeP/dY33b
ORD+JvCPVGqmv9G+Ohzm9ISPuPvHoJeTLgzLsxSa9NIOCyfk7EpocCsvTLLh
lsbykRQxnRq7LhalDA1S+OjntfX335/giTThPkJC7dI8DmOcXekZ3xUGFZb2
YuJWKibdf1q8DyHRGbf2jqabbCnEpKed0TertOWNNYazaW2lB875nfFEXqkq
5t8heJf1gtw68UhnaiWcVnjj0pWtvS5H3mmMP4jxDrxCvoYGBjTJq6735JZP
b2h+oyL1cmK0gEK71b9vIGyFNgFNfDNrQIL4IKpSEzccdePzmOq/QMHSXtcg
IuLOZs9FWQjcaEzi2ZiUXut3ze2yLkvECveyP1pUXeWm1eD+gW+RMvnNnf1h
JaJKH9umMXRjAPh7kezR+MxDJ+zMsG9KRPxVElHkxv9IyMluusnr6MjHdfNq
+XsdotdKPKzDcaa/ZuU7W2Q2nObOaJTs4VbAfyYWVmiLw7hDgFx77XU3bV82
1ZgVKO8GUcYgB3hIM32GNa51VUtw4bhhtJYOyltCgDTGAjaysXvhSsPVJpSZ
2iBcF8y1CB+k7FDZQhC44j+FcxEuJJBAoMnLs+KA8L1hkRY/IeGD+UGzwbI3
MU1Rcohwy8Sp9aMZ+zmVjSfWfC5PI2G3QOUNsLCZ1n7Ropd47XNDVkUBa/49
IuRwjk5/CVAy+iO94tlQQd1zqTtMMEEFswMN0S6/Ocr7GPFHixrkrC0l7My0
aLObVkyVtlgnIbhn4j17VQ+k1H3kXdQw6f61baNWreUdddQylUYj4JPeAG4D
B9rzZXMauvF7SU3PYYPhMvYtUkD4BtpgLtlTfz1YwgX6CdT3FhMkdrB49YQZ
V6UNH+71CKobHQgvugKsV0QDS/bYsW12RxUI/FOiaSylTuy0Od6zM5wpGg4s
1gZ93PIu21Wn7sCQN1IBmYYNNf7uFLjW9JFIh5FpcLAPQKc8+HQRKQI6qkrQ
fYcdc5DRWEcB5tYkxPMJHnmuk0fkXR/6LVBa+31lo3Zxk7DB8QJjCkTARrmm
NyrUXvEuF/oj6f31Gkmt/5Cjmpy/Od4KH6WawHcB2WHHWaAnez1GqwnBtXbD
luIQsfTi69BKyNuw0wkPrx12aQl2MA0F4fq+hcswqXnFe0GXM23KCPmmhSuL
WDrh8bfSREY4JojyFkSGjDSZKPDd7O34eG4ymaU8M2frnwTG6ABqqO6P8HCO
66ezaJfXHENPwjQO5UYUss4bP0z6lCKahtg7G3jQZAnSjVeAEDbYFmOgI9AX
wZXNv9enrwjBz0MJxQgELeIj5Wh+3L4+Aa+echpyFI5Jbx1tKY3RgEjtcbAL
q8hPgUwP6SjzQ18pH/LdKm1ED0cvlIuYVn3RoErCJj0LCGtsTIX/rF3wrb+u
qg0a6hdG1Au8Rby6svsx5Pj4yXmgVHgDBkoTMAhUKmg6s6es/WlFyqMLi6gf
//Ild/aL8FHh4nk9YXfe3KDaqzghHcnBBVmhWgRnPUstggIzUd87UY9gPbiw
U5E8kRxqxeVm5aaNqGQs861dDxIW52g2fl3Yu1vbO1QsvcCOXJYpfKCS0mLr
zoCVrCHz+w65eC5XZd0JhVDQkoEGCmPdiMXpxWgvSkGgV0GpRzzm3JzRhh7A
YxEbh61eVxHH/0VOpoFSPlPy8ZeFVFLl5gMdCI00ByRyU5bFap0TWhxMIAjN
uWA5qxCRs7XvFeLvMebn5H8Aru/XCPzFPozSknZH0QZyHvpPqeTB6rBj0vNV
ZyFA4WY3ah43c1KcbVxyAZQOfTjOGyrH3R/29WP1xKYfhDJOHu+sbYerNYhi
gpPjggvJE4wfn2obdwiyDcg11z5jPHFauFohNolDiuFjP1PldoY6GxUlYvzS
iyHGKcuT9rC1vx1y5Uo4Kk34GNZaxTWykZUSQeyh8pVmFxn8zAx2z1qmGlhD
974c9glInvA/EyRHzYtmU1Il+Yc/Fo/UVQ0ELIX316NffxizcmoD7Oftkjg8
V5LQrg9zvvP5nf14eAtG6B+RNKRK9T3OocwFTG1FTmuCy7fCZs9G9cfzhGJA
Mhy76GpramCo66nO+TVx03jXA7Cjd18o7v9oacsR3s0IlC6IOame6PXXC+K3
cK/Al4YHicMVBbPj8gsZHnKIKnZoTcKHSPsqyWdh6527WMlf6AB2XDV86di+
LAwulHmq2W6gvkwlmRAu5SZDUosh5N7ePgy7GGtjYXReth3OnoM1vgenzxjV
Rbv4qDPX92Ci4eiYQk82W2qjrn8yW7Zrws87+aAihf+sg1VMDZZR+pnlQvFY
mqg1ZBEQKfmKYFG5km1U5I64ksmQanAVyqg5XFwy7/MqfecJVAS/3MEK/szp
D/U4zcqNP7QrfH3hrIgRWK15k83Z6pGKGhE+aKFQsk6eJiZisz1wAyN1YT/f
GDgg5FTOlphaPVtj/+ZV/iMyoenyt9gmuKSkCCMddKuWUuy7LTUxM/3VNh5l
LxCjmYwl2q27awJayDGK4Oune6FxUXXrTUgv9wzFdm8kNPEgYJkxx4FSSUU5
P5R01IjwTwchq4ffuoJL48Qd+f4BGIjucf1b8e8qGOhwlopYdyxTsRGjjx3C
/3ki9NW32ZsvSVfebDJdsneaRukwKkbrpfKZuzwK4BTeHn6rYx0wdKLie+/C
ojfo4cZVdV13iDDd5GzHfd9jXVtU9/f6PLdMlaWElo2aV/3Nn7EaEcbJq1mn
aiuCIHvEph6XctZo6MutHai5cJyiItOELOujmy8L8xSp623UBTRHn7OvUxHO
07Dj2oQuqCEI8St90t0QaCulDsAexlvKKZmxTTRKP5k9bVNMQbqnc/iAL2K3
NrdMigSJAFEFXjyjZizEUp6lL8x8nREAaWnrw9aMFrecQuTN9JaeEUvRm8YZ
Nq5V4RBWH/+E6ghcSyduDLqSzj6lusa/nSh6dxMEx8AeEvf5QWb2nmCyddSv
qvrX0TMZYEvpjCWsHjcmX0s3vsD5v7uxlIE/kVKAMfHXj4kxRdZ4bxBAiwzO
eCFQaOJtrKwg8yb1l+K/ieVcopjuJAWyLWffiak9fmVbquvqP/xu45FuKDes
mun7Ke8XDqsY7+l0n0fsZVwhBklfWHejihzO740iXVjucKQb+UO8Ddbx2ZnO
JUJyiq+91ArsjvoRua9uye6/YjnVlcDkoTKsN6ziEvCAONzUnxv+/nKMaRQa
JaXN1PImwiqkNVl8tfw9nwBLSVWCJGbYfehNbuTBun+TexcjKBiKK500xtom
VKkKTQcDdZsNjAisWwz35VhIF33m3FKfqeudyOdhyuNWQK+Hg+PhZmW9Qsur
5BB4S1saZJtV3oCDPEY6qFD8K+GTFSdpA7nKtfWYYOYqFsyDgiKIQL5VZ//z
5sf8ex2Z6XAqIVsgd2STSWKUp200UsYXwFRPnLK81+rG/h/Cf0VgR3YhD87K
YEswNevLjQY+rXsPgccqsR2fVDTaGZJEHyy/imGQ6G9fHo154M5gffMguHk/
Fx0qoLFMt6WPHbqcg8CRd8owdu5TYLRUf+Xw3olhNubbic5PN3ZI9XHuVp4U
P1G6c1XYHRUpZjV22k5vvcfXBmlIzcAZh4/m+puwdTmcYwq9FgAOio40gdQH
R3jwci76G6pIyTBivIX7jTrRTN4gitCmMDcgQgynD5GRVNmpT8ay9ui+FRF5
ciYfX9WCmumbTU5BcwbPBPDg/nY7ehrRovV8HTZvUVHWhGGdl6sfM1AnIwbS
h/qxV5A7Swf3aWiAACaXE4RaRyKhfZWYopyMFqIJr2cLB0IdYM7F29aYeOPc
E8c5vtbtZPChsVklpvWUq7h/bpzcvYXEsj5LrbtV38dnxLKM3/0C0pyvb5oD
Cd4U6bBwEs1VR8m8nxSvR8IofknJIA6dIzc8Yn/6Ct0d1DkUsYvmhvdVKtOc
N502+Mfl2hzGU4i6gFnRCvPLx4PZr2L6wkq3pNzwn7NFz6EsjI50l23WXBhO
g+HGnhHOELDNcB5DCRK20TTY7vau2CHRmXsu8Z99cAYIb/uVN3aq/J5J3qiN
nNvQy2k0rv5bbUS8e4/imF7IWCIME2emr8dTCmjmh5KVnUxscaTjX77InY78
ACsE8w71ykFu1wXXHEif9WXJxtWYyRXUCl5Sx+VTjxgOvBihv095VoKH++dj
MCQU/bh/BZI9D6kPCpVKzqA1rK29aRSzGsif/JaqizHOohzBUn9QF26+QpYV
0lOB8QswVVxYBXRgvsum78QRlqNCcDcEnjOLn+nFg4+CyiT9bZqtNtbeuOEN
UYMBD4SmY6nd6g45RBA246lbWGGjkHjja+Tl+/aYG4tlIvqAriiBKJzRtd30
zuAVd6LaEvKdx7ttIjoXYtnPSfQWUxkpkfDQ/FnpO3jw9Xsc1Eb/6MVOUOtx
sWQ0n0++ByVko1R//Woepns/hFFtc9FMA5twSRAeCSAAdmhpOex3LFTQ5lyh
GGCYZpo4w6Q5sef+eQfH+OkM4ZRW8sULLgCJTqy5mjVeNaHtGpDv44UclYJo
uJ93UmAOF0ymG08FKUEXmNVwL/rD9orGNgUSK0nV9uHlr/LQ6s+0Ua83TFA3
SzcW3rda5/gAlS4lP57IeX3/x80+ct+ERM4ppUPe0UHkFbP+UUp5pm7ZaauA
SQGXMPzC3fBAQSmaNYLQbIg0K+7ighXATjRVmETUJSh/aBEiFbT3CG0BHc1D
dru31iHRQpdiLWyG2fYyj1jXNZxmCVldJmRO4edy5huVyUy/ftqVKfBJON7m
mgWqmzjB4Yi6RkJM7pQBC4IG6Ul+6dBPeBlVun9srEnLJmnHOLqdSU6DDGBC
QfZGTciNkkBr9E5l1p4vDr6ypv1wodp4LwY6ipADPoI57RyZVxASFVfMEZkg
Ps7ONgTjgG3luBmWZVfH5QzzG4ysYwMhrHvzJ2pV7kvXvszW7dEnrQIdq3sr
S3Q3WTQ/GQZyfxGc3wJKSB9TxMRn/4WUekjOXs0NWQSFKUWoMajf6l+lyBwz
kVccxGZg7ciYVKUWjQA641POIe6ir8WUzm9Ydnpaw/9q3tVRX1MYr1JFa2Hc
MmKOkVhs1VEp0yC7xnLzOMAEr3nMNu7w3IONh5ESC3k3GJEKY5jaMtLqlu6b
EAfEjs49eUi6xRzmzl2owHmMdQ+9AJxq484oAa/eaO7Wj2Jh/VXjNLF2cTaG
YzA8cZCLHKxFyapk+LnYxdlb9xMFZNazae4Qb4OWY4hmwrNqI0431wXMrcJ+
N36HkrowRj3SIzF6vx4puxlZ53ogzV2AMp3gMlu9UYPdL6XjPj7hVnfqQbch
Cf0weaNm7lAgvmGmrPp5Idp/FEAgW7PMfqogh2LfXdliQZPTafWhhGfM0FtK
xOu3TP/iSin56GhpMfv/6fcqSfSALTFccTz0pUnK99yMqml3dCUzYhNFEEmj
xuCc5owbvUO9MWLA4sZVXR5u2y/Br17uIaEovdSi0MBp7Vog4nbFAzqwya6+
AIKmbbR7RMiUb9qSb91ZHrlpS8RU1pHEaGjaO7h1E1C5iVuHgWO1VBMGyA2o
4Bg4Ac81NPSVTBubxYR5uMrOH9SMapGkPKLQqLHAiawWisGthWfDkHHKXooO
JesTsmX0lbuY6vFQHgib6qINfwcEv7fy1yWvgmX4JLxBdsoDog3x7yQLEgyq
SSHOeXWCaSBfySIf8NsqDW+A5pFQv0i6JIID+pRLrBTeIzF8F6KLR4xhSp3G
TBTBfsiNciyG3Q0tK8gYcK5tuQTomK0tH3ex8G9tOjWUJDrlxzBSoCX1zKn8
Dho31QnqToCeGuvhDg6smyP0ZPTK+pAFHlLl7oTeDi6HG8xIRHMYOS7ahXxL
xbqjr9mCaPbRw7hYdYeLJyQ2MT8561iAcrfWNohp354vOCobzvxBwQ8+DriW
LpQJNZ1uX3iHDvNhgIFTJTCYd5d5DkdxIifIj5m47B9kSEpBT7/3dPxCCFqI
AUb3gAoeSB1pkg3xPipRqaPWnsN6JN4UPA/ztoDnDg42C2C9E44l3rJLbVKD
xgIn/a17EOBdzUFB3rEBM2v2mcyPsSwM+p2BnBBqIMrQWLH8Q7gwaowxJWeR
w0fMjXDZT8iAZYUmglTrKLz+gNpDU6jgCGSXPFBDPV5FGZQh3rAEgqDKZceR
vEKqVXwLtxFuWV7sPGf1Hs+YOuHWcjwzSTOpHh14rcW4FaPAM4h9SCEGG1iu
O1Brer+LS7soBFU1Q05pBrudLDHtosLvdLjM5iKMXeX0SW+PlTgBBJXSszB9
NwX7Wh8p6sUfLyazoAsdYRenmWq+OixPJ2rrpGvc/9kx0yXSpFTBAJVBZO0u
cfWfjDIacGoelxeC29N7JPW2EOjzrFf//X2ihccO6pzL5zD/dc3EAHW9VpGN
d9qGlyYHkwHhkA+RtLZU9o03fNYqm5ELhZ9K66KnmIEH8lydC/xio/FKUW75
A5w3TLpTtiLg/2mVA/zvAIAvqh/YARtGiWKnEnmwOlLi4jwyq2sV70IhijYC
Sv/IGF1B501RjEKXyS24rJxv3bxYatmXY6OEs+c8SNEkqxGm69rcG9I++WCo
0OCpvz0aFOCiDnoxmb1jd1oGibymt6UK1z+O5z71hrW4Wb4fzRAtLr/oW6c/
Dl5D7220bCUSI4odEDIGy0J6+tW4nSKtKFE+MuBuoCQVoR7mg8DownSL3gqp
JfClSaf0zKoKl3r+2w+EkClYHx9kQ1BRh45ct0PBh4Mgl/XSw3lndUppp+iT
xBS8tCqF7/AeUDxJVsqKfaDx7JR9h7w5X5/NorHHoX0wsm/yaWOhbOQNe5jd
8i2sCWqKyB8JWFYRWAzVcsljHqVypzGwZOOjKXZkOWWzqPggTNsT5bReVhgY
Lk/1loM0FD2sVCXhX7r7oj8K4Pd55x/Tl78OSodsSvlFoDi+CFP4O1ne2TRh
KgahV5dNtPxCfX5A9cXzMfEaxn6EYb1pi4CgBjSLTy+PF3Y8hmdT3q6ELRuw
GGnnuV9dCMGwMRKArc/3gAhzCvLKOZ4z07O04CTScgRl7nZUksieg24AWZFp
SqA9B868ZYkv2Faz0elcpuRrsZOENvTc9+ph1o+6l6fYPSMq2s3yIrB52WYw
JxtlgxerS6gE4xT4nVqe++p9dDcKWKfnwfwx3L0/PxNnhoMpTArLqqZE0hBa
s9iOwPN7bfZ8dpCRSpqutRsUDRIrqc1Q8FAiHyTcohbG0o64SzAQFzuj2bM4
xS3RZBDMe+zCfXQsONo1bkkiEx12yCO7jVODdU1D8o6AtoQX/GcydGfc0T+1
bMzSqM255QkQR9+65Nxpi+Gkf5ZIixL9BTSlrgHXBSDA78I/hAvPH1S5YWVZ
wzFcZc8ujBxnZaDRwq/s7uCDtWRu1zDmcyQpD5Mp+CbgfoFGhNlGRysmMGs4
d0Ff8usHnEm4cbmJeFofpLkSgt6HwvIO0/nGSqvIaz8PI866k/i23NLzPNnF
0koIYkJ70PXScR1Wn8i2fXfX65DvCBgkVHEUNF+zDdxGVmwRdcyV9ne0nzeJ
SzSZq2Pcv71mChN+9r5fqV/FLdyl1besXK1KhqRaHlj+dVVYTGg/C2Na94iV
YTZxSWoR+I49fzpedLku1K3M3slfwcY03rdRK6a57OCdlfamCiIcpEUM4FVw
+w7C/at5FoFnX7z/prrKMFh6Iu2jf9kNFF6I7ilGpMMDB0hjg71ejrcKimWj
+ESFltUseBKrFN1WaIdHc5p3PR7S/Q3uRPTAGKgIC0VzhJBM4MG9PJaHhnKc
Wg4Gx/7A42iUgNxFc+5MxPlez/4noHI82eQXNZTGD2culSsUHLZuwkeZdyOI
iE/mwecUOv5yScRmSJuuNExw2zBW57NZjj8+KTaD1Nb0cMsepFuAW70D+8xV
glve8SMroginrpSZEiPvjcHWuU5fnYvWwuxVA1H90oMOl3QvI9UtCCr0Vrsf
xV1ioNEYTZ/WiDYA8WEQO/fMjNnf0/sDrE2tqhU1FXlQjldi8KxsqFlpVW6K
YEWqx7pS4blkR34ZD5t5qBzBIi13kbOX12T53+2AZ53+uj0ygshJLR1dgFjE
ZiWrqSHJQ6Aomra6JfImFlhUm7jPSQCi7nLtz8XYU1rh+pP0i+QrN1XfgQDE
35lTrPhJsvNaczpGZGuUw+mbYvMF30mZE5T88SCePfjtWZe7evGY11odFhgu
PnE0DEPW6W2lFI4qCXXUyZu9+kVIlJjJAc/fy27mcRpz+g3u+Fefgvk6F6jq
vfI5U+4IypQKPb3wFP4BOQdKvd8uri169Wy9AsAqiBRhsbfLxpmJA0H7HTHc
gA+ANtrqkl1wQIBe+fCPk2mTs+6XqVfk/7vH+1dX9ddwpEgiS/w5bTBJHNh5
J76D1S5o6b1O5UrlalREyGI8YtdOcs2BhAy1WC4S5CbrBHKHvwZFPbqSrQdZ
ilvbxrrAB5g7thPfcPmnoa1A+mTNk71jvimmSN5dtwj1gHzj+7MCwLRUKLQl
wd1xgaVg/RthxKY+2Xsf/FhwFrsSRzwsFOjVLXEZSHu4uZPZvY/RAKLn63DG
r0PaG3MfR95JUgqJxEGbnMpvr7JlaIdkZkOUbuKcVfFiG5rPzppj/l1Sg+LU
EaxItgSs17IniOuvpWzvrELwc/o88t38iC6PbVckYMGRs580/cS33bhkJ5LE
jlLC84Wr6cBG/+VWZmDygLnyEoujyso4Opq3edPGvNfYYSqEC2xTBfpAeOZ3
1gqtomaUy9vTDiojjyyRCQtFvMLUPSSxBKa+84Cku67pq5wK4RS7Dq3EZRyP
+UtaknySih0YZ+ozZ1xCjqWvVLITXbMpUEv0UXL/cpn/Tva7koLyCGoUGoKu
rtISah8RJHQbNDlTZXqIlGLAS/DbkerXiN2WRwphkcSU+IcU33S0NqVO2LLc
bi/jN2QMeqo5julK4QNm8ICSgpzotChRC4325y+FRX+uJpal8w7rpEv7R/9s
Xwutd6lXbvVuBkKB3OmAjppmlIUBj/lIZWkcpneh7z3oBJJ9vrR0lInh6Avs
5pWxkRkwva6SFLLQd85MFSt91ofDQMA2p120JQuDRl3H16mzCvo1RbZwoack
ZA/Q7xMCNsigDmtpkKWEDpDnqiscpih/c1SAHxVovGsTMh7itvbZYfv4zwvG
64pe9PQ00+rTa8QQkInAGZOSIYpSUF3qPUgiNbc+IaMNqqhQShqHFyjxOe0z
h12qs9R+o9c3m8PS0nudzl6QcWQmk3i3K14n6vTfXC/Gskx0KWXEfhQ+C+ry
1IXb1+cB2dzDpnSegTfNqIOks5bXSTkW+g6vQmzY2TMH6jv0JcdAVDf+WWoS
Pj+vI2VfsMZDbHTjSO1QdnwP+tgqU7vsQ0kR0JPNZdT+bVk56dBaa6ei/3Ex
GVMyz2DcPr2DHv1H4eRBLIS7DNeDp6b4sPBd4mzP/RaFteWkzjrAkk8d5WjQ
6msXoWivKluCEoh1Oe6VG7/rTG58Byxs/x501A+k4KLBnvhg10oQEQim7rEa
sGO7k/BavSXdVg2j3YBKnFLskrJV5l6SSCN9NS/DxSs6zCMg3yXzzaExeuAF
LXdWmygkqN+fSaOOb+QBya6AsJolvocidLWy9FSvY/VOjleboOfWejHbPMsv
p0hp14TpjuAqSKe8AWZOHW+zdGaib2IyxjI7CIZJsVmSq51zm3qzDL0ETr7W
Gt8SQ9WP3kMDAU6wuix8bn9Nl+9cU6m/dLpIlS3SCFg44tUrI95NtngW5TNN
UT4fhR206EnJPXmH80Lb2I8Mf62/kn7ULF1CiaLPeqwFLlAq3xGBM2DAAWfD
KhoiJ9lJYkU6KW4AWstSg2+FyJAmefofee16cWh5nG1p91BapKLUQcA3Jnc4
dBGuj45vx0uKlWKh6ltovxxE1zGYBaOvu71prYJzh7ohIsEhjg1VDteF5Xwy
cTQDSCT4Wp3ZMXi+tXpIe5EOhnsaqiamdL6Jk6TR5uSdbjkoNnlUiRjqLUMG
nq7qoo4+hEB6gG7sxVh5d7vqdYLHYk1b8N+66AbuLoaL07Ngr9Vjd506tLwL
mFugokuzQt0k3RFo9NWeQIOkSZJUPYCO2jeZQd5U9ikdp3utNgvRHf8q05bI
DryXqYSyfQhPmVvrOHpTyI6UhFqBOSNEpZdtjzYWaEo1XsWGqolbTJVZ51D0
72Frm/bdfL41gi43NS9bTrN3zQhpWrT783mimbgQT41RHLJe8gAb8rsDT8b1
vmBga8SGrac+b/k/zTAZA9P2Xu0Vw4biIpWEHFWReOKY+/qR9QEMvnMRqHeZ
NHbtDShvgQbbs3Z8SktorIPjUFFGyLihN6uIFdOYwmdDIDxUzsJh8LTgRe7p
hX5jQqgpRkXab00M4Ev3AH2Q2ZP30S/IOx5yubn8VVTIWBZuCmHhrz02bE69
cPLv+Dlzf1Z9HayWzVn5f7CW1rfmqUSz0ZQ1D6Fi5iNs35O6Hj1z6kcYuIfm
7kEBHWOnipi25EzHs6Z+0IKr/xlhRhdKVPGkua2bbyZVGU6xBb4qKrOqcBM0
5STSm+B7FJykEc8ldQiQUXAe2rKOZz8uMOgeRTwj2MBCyC4FvkeoDJp1HCJK
/sdzKfoTwWxmvZHVD7/fCOVNNMs6O95UlTBZx6pfWKPF8BJHl+VrMR37+IKD
jrl5qZDY487lUeDqm4/pZ+RugGxpjmztwBpAsiQuWqKoTWIrX2QOc5OJn6gz
LGAmF3poUgeSYeKGgvb4j9GZNDihCWjN8O9nkH51x3Lyg3mN1ys8HSOjIrs5
7vkDB6gsqCb+u++GcmiODHlhQdZZ77T6T8ypfvmplNnmAShiOMzBgSgAyPMt
6J/Exu7SU3a5yanbYJxmdviobUZxQC7A/uG6C7CwaclMPA0m+iahHA+Ddkrn
4hAEFiDSpB6OnGIkxKkTjfFWVC0KT6Z/PSvIXwlMkyscT/FSTxmBvZkGG27V
yObrNn84PBWaDlBYTNVqlg1HQ0bMfjK+hjmsOngDIyIozHWsE88AhDoO5rAJ
b4WAkiKeVynV1r+HMG1ltls77wboXsOOf4L2lifKJOwgzbNsVxMj9d1uAJ9E
JYUEMT03pjZFzgGBLnfE9SsAocmfca/Sp8D88L1T3L3PJ5AOdYb+gD/3yAFy
0alVu/RwKm0Fewp0Zbba/RAOtirk3b5T1IkaVly6aSx4ev/jiyF4thGmMtLa
/R9nRfTcA3jk9Ve4/P4QKDaH/3r/SaKbbc5ip6N/ngoBGBoNdUNW2vt+52B3
JMjJmDy5oCVgjDU2Sg7qGG/ureHqnIkuJ1oBS/wmjm1zcXU/am6v1YIPBsV3
FuNJO48WlP4OKNfYFcOBeL7/siOQsVgDI4tCpf3/+vSlq0bZD+3uJNTT2Y1W
y4BcPbp6M/c3FvLnYR34MlrHiA7XELMUfM1ci6oNjAGR60eB0m7Xgxay+Yjv
YLS3YrVbPR8tCNhBtIzYvivRcXjRaRLpqv38/3NGFI2HUj6RFi6w87muWX2b
4kgqLdddCzqtysFLwEFLbepTZ+KgIeXK4imdrCRXlXsHPW0oKFHzEVPP8r+8
OYOcmuabtds2ZVP7R/iRGj+huctZpzllGUJl8KIQmRFLfxVn2LJfAYtBLWdx
pIQ975X8PJpFcr9msb+gqqh14KJeXvxJ4DgKeQCFMAnhoTqz1lhyCk/sR41D
lL5oDsU1TPL77oOauLsM4B+7h+aUS8c6ZpFHoNodORKoljTWvnrG3KopKxlO
GFAHo0aCDRa9EYYs+O60Jh+qf65yiJYlIlrVmj16WUWutWXe9iv/pE3w/Egs
PyETY67AvO2u34GYz5u8gjWdjd207qVzK3wtQOVbVTViK+E6Ny71QD9OBxgS
shu+nOwqUt8Zg1WdwlZZEV4gRSgEJmXjjkRVBJwYSm/LmQaJU1wAOlCD7/xi
KH3acfIdLQYMlFXKdM+opEdOKNR3f+uXrI1hoWO0sG0NI9H5FuygR4/XEaUL
xPHOW5Nh9HZVw00rWpCGJFz4Vhqp/mCSMQfdzp7aqEqfUQQ/QEp4NwTg7lX5
tUylgZipGcRHWO/emPfPzEQe6HF8MG79VgI+nnYl8f62H3gDaysID8QiYEag
zd4X7ixMLoNQnlRe3jLMPyZ5D1F5R77nIgOj7H2GtSFr3rgMAo8MoKd2FtAb
biHSvpvqqVouCieEZofSupxHMRXBn+RFO5mH72MW6WlescKSIOQLas64b2y5
p8W/Yn+c9BRmmyGT5VsQWoHxaW/K8MYoHMmoZ61DlAUq2EJuwrLvDFShlDNS
YVd0KF2Ppo07hKK/Tydx0ZHcTXMao+q7kLIT/wa3QS995GR0tUl2EO5MwT50
3puWsZbt8G6Nvu8pSwRABWgowLzZ90YZy58rm+QqlAT21FCAKxLzykbB11Qh
Z545hH8WAsRWYZwqBySsnwiH/HywrYLBWO6CLgjOx7r321TeM7TWWOs0FLif
xQCMqumZ35ZXVdtn6OCjjXvomAcQwuOaUzb0klVn1pwfxUjPmz4Webg9CgCj
tB+IJwTrbaBkZNuZjA6XGp54MPAtl73hZF8Jp2945i6KdoSkaLLIEnRGJX9L
f/pvEHL86tua9Wgnpp13io/klU7rNw7jdifHM3+8PJEZ710Bu6ctAJO1O+0E
g8Uv376JGhumUW8zgIHHU0IWMjw7Z05vfEQTFmcnMD5bNriSKZJY6e2/Tif6
iUe05379s3VSYh54VsQiq0Z9XDGL3w9t8WKaJZTB4O4/bY2lyxyJBkrIvy6q
oYuZxDn6X1yvSlgUKRp4F+DpiwrArE0nUDHBRQBHydyFI26+w66Z/f0zjZv6
t+HllD9lu4/1+LPi3YZRHkyYmYLGhILsm1V86Z5k08sMls/HhaLFZU9iCzKy
XaalDmKfP9luWV47bzB/uZVoUVvoVpA1XykkPqI6IzZGBXSw1hJOvzxKOqWe
N2yYx35sCFa05eMSbqFkVwEsCS7dMPqWX7J6HYY1SDdZMGCMn1zUXC0vip/w
cCXo+Ach56/wxvwz/U5y93yMH8uuFkMkPWhlyIolqMvLAtrpL0SkQPIH8C1p
4e70gT6IC8ZaQD7PueTrzwwashJoAIG8Mx90tMmkIY1O6XQKdwFKoIzxszhG
4gccpgzjjn2QMQ6QMylYAleDAmOev7sxK9d8RYaaI6pxe2diT6UlxjRRzag/
zb6k4kYKcppVutuZuXhVkzWR/6YxBvyxDYEnzGAk7TXlecR1QUUuCH4xQX+A
WooGzi4OhOLxJPgKku5fl/UoBAuTafuAQrfD6zsc8f5PRcH77nfc7FhMpMO1
tOcBBbNZRe5/4iWs/+wIqlXGvZXNBLocYmUiesT5ndM2joNDrXWtL5GmgZtT
SbHLOhAcIXbYuRAYCulGhIwKlpr5BEU0rpm5YEhcabGjUM/9FDvbHUrxr/xn
Rt2MN20y9BwMxODILy32K32p972qkqdZHBrCQWAjx6JRbRGVbJBao5oTAuF1
+ygrYM/QEZ/CUDw3+sg4kyhnRIENEo7WmE/X9/i3rGQQsInV2h4W+32N8Iu6
R1EnvOyiiKJYXQlfRx4qr1EY+Nk77nGJzd3rjP3UiMgIQDZt650TTZg74xEV
5o3Y/3cRKRae+YU4YkIyLI7Zf5hTPfg1KPup+L3wRAkC7iXV7qiQWLxV0FCb
TOVD40LYnt152VAhHEzYsP9B3PljhYrQNG1y1fhwmsYlRq/Wu9TOFJ05zkqS
PE9wZMGxvC5/NidoHTZ1XUPRNySBLcOqCuHB//eXu1fJkSoiB+y5OdYcLax8
VYmkmYyYVufvToCo0hN0VVkLWR8EX/dvVCn+uEGY/dotxyFirokuBa7+3t8l
ncn3u50fRoM42gbTLkkYY54fCx+o2HIjLZRB9d8yj7JI1Sw8lEXUVFQmPUzA
AiH3RgySkspAIMG9iO69BbYJ5jgeJsl76aPpEP7yCTKMoabja3hKnv80xxyW
HEc/ewhucuob8sSXGaOKphQKUtTRtN/ffJiQC2dSB7mEWqqQibRj6wUQGF6j
d+Q0Mvx3tb7kFx2kmQg9YGk06izaSepsQLu584y9bliii123CshRvk+Of9No
VW7wHshzdNUUYhYcDFvwTYJSNx/QtZPnhunTHjloezIs1g1X/G3WYt1AZ/da
VaNlpF+Flm5m10irw5YHRDET4Y4CQp9w5wTLbLTb8RD0gbQSLtW8Pc2CfWPm
faXxMS9gBG0s3ADH1q6x9ghNKEdoPFewn0JmtA/leSdFQBOSvx/qA/OqzNt3
HxW6J28sGb+sGF3cRI72djyzzDxwbJ/RFV4OHUgrUW1U41HRaAOL03pNMYmT
BYlbbh/Uw6Adn0oWb0CX6dJWq3mJJh/hCjnNA4ruLmvF8LwnKJg99tGW/0md
QiDkyoevwF0+Pl98grVZe30eyKQEQfr29w/0yYPsJ7F4pt5KSX68x735v/xJ
21zUQw5Z9b8a6S/f+nYoYLGKS/WYnvfI88FQRVczHc4zg/+HUv9mDZTyzSH5
cNTnBT2Vr54oNJgJgJuHznNCePcjbJggVwLSvmfrJzCP47USBOtj1cbB9kf2
O+0ogA8WygKPDetgo5ZHsZTZmckMiC43ftq1bBcYDCNKPLCwSMBca8kUHyEi
ajDhlfgVFumLAAvrMI4fR59902gXnoTjC9CNxjZkOULtJHCm/lRFRA2OYH08
ub9skHKG59PrUk/e0XikL4Ce7RaeSxv0/LDdmmJVehvkeQRIEGrm8Hnyzejz
AqULN2pnn16p+cgCMGBfsn9AEsLVzAeeWzjXSPLLJcFt3kXLPXx2GW6Fcl+q
tmWahh0OQXq8U65YhBElE7ramreikwshWo12xDH6BkV0rkqM2mGtJ9OePHHa
Eu58uOru78nei/g9SSnjxlfV6kuX8SlERXeOShyfvZSxnUQRXdMSUjRjpN8k
83MDzy1y5rziPj9jZQZIHYZH7ZmU5avsmLDj+evlA++8gJ5TfWuzqGVQEqSN
4IJp/ke9qG485D9pQgjPch30wI+KoU1jA60H64uDHLb5i9pmjywokxcCjcQP
D8ARtBQbceoEAJa+VC9iQ3weNjmphWbTG9NrDNNuoQmjKHv02eUZz6vCOG72
VGhAqoVg5iLL7miBWEzWwvGpqA2m8XHBMktQNMZBuqo3edvg1FJVvT26eLGp
mTIFZ5Ax4NdLyjxQCGT6cneUcp79Fs3kX0lyv0oyXGrnUecnw6ede7te7oXC
TmKcj8PSfyT+JsAgr3lzwoKHug2vWtjrSD2w/gR4rOIOBsxBvnqq0/ABgs1i
yxsVn9L7C+d4Ux41M3w+QcgZf6E5COUdikUYlKMjHgVoPPlLtKFiLJomip8Z
q1tZHiS3LG2n0OAPmHSAq6hMnQsNjFPFKlqc2BFmfbTqkQYX4OfbiHsesAgh
AdzwucgoVbS/r5kDufyiqajbwC0FacHzviTOBw/f7IgMvtHQcnK1rS9mlnCw
ZPVU+avhjxLkW85F0If4aRBMS0TxfI2y7CHb1U5IeGYnHrSxFgYxTWaYGXAo
iesUXwKh3e6bSYUpovtsueSy1CxD7g9PVAmXIaK8AY4T1fNgdt9mwdajStpK
YmjLDD2orQjaYdA7TLZwBOwVVaMI4J/4GjXbxIKg/50o1ScUeMtc+25G5eTd
/xx9Z1Sopla85Fn6MpGDPOlSMcNwZ0Y7CZyk9drl0l84cw9f0vNC83D9voyk
wLViZFQNhyf4nR3FjMbQoTmy95zoGTWgtAA35LDxGD1bjm9l1FX/yH+OYi1Z
kmLD/yy9PIZRJDFLzK6Wob0qimAaP0iM1LoMS8YlmCHx/ShiyaUVeDThj9qf
AUnLFUkq1RN82tT6lMqud8RSjpx8SakaGA1p/HpGVSd2XXG0caDT3Bh8JgB4
peXxCj1psvtLqslmQ7fqGICkjb9s2vJ2YVWxTSVNi5rJ6e72SDA0oWN7GLws
2SOlyIxJ+76wTAoO8jpZsd4QaMdRN3sSKofxuqm6SrQFDTFXCiJFpSvtVBnr
sHhDzGxUOoJXImY7zqrp85JUEx9DNlu/6gWNr55L522+Lj0i47BJQbJZ7ZTF
eBO3svfH11E65nu004lJhHqhNl88twpT702H9t0q8wjxDsdp6bhFDAu+utKX
vtv6Aw1QqxDA3fHyS1wFZOLQVc/gnmiuvjx1fwSVtzuPAuf955bajbUugwTn
FUqsByxbS46FtzXnFBQi4KMyuBgZK03EBQiNHmlF892oiAjqX7CarVMlrYqD
M3gmBkekBXvKKY45BvkBVdNttgjtCB9AQ5y2Wn9P5IkKzYkoSOAp8QUjR9u0
DckfF088oLVENApquadsslG/R+NNH6GgLukB6MCjsrXZpeftu3kIPFbW4sSk
xHkV6kn3yFfNxOInMbKPtbpgi5aRvYIod32R+ejP9v6xXs2ZyscdCfiewxQT
LhXLvIpxmzNY1OqYBfxX3eJ5Adu6TO/fH9FYSNJbPtllAnVucrcgoqhmpZUs
Pp+b/oq6Mcza2AS4ZDzwtQ8QvV1tVkwifyDEgK2Mtbp/8pMvUuo7j+jhf2GP
FFp9jO5o2burtOU3+CzLqkrq+zyt+QLoqPxeKrub7Wdv919WRaypj3ZwNeXR
LtuGUSUzpFPinbndrv9o2YsZq6A2i2emdGq9w1fQ1L+1udDpSjtOWbG7NmrD
rmIf4/MnGlqveDDEszD6Gvz51AfbbCEU4VEi+RB/0Pj7iTs+VFU60tsF/JUd
yob246liVKC67XFAv1cvKzqkhg48g5OafqCcp0B0PbVs7ktE+ROwJvbVy7tZ
FG7plrPRXExuo9NuB8gchaCqVzseKhOrHbFwAR2G1TcLq1gA56ZgsjZwfVPs
LNGsnQrOIHdg3pMJ0SRv+Be/yLVjqfLY+ZvwgNFFQfN5kwoqzaSukYCTDF0C
EJ7M34ov1aoDCI3l/GUm3mHY9Wyth8TpIrwyV9prnvarIjmrOB3I22Qx0T28
3axzCh845ktnRDlGJ8ROjSNN9RHVapfVlDumDH6TZhR2YF8mzsvjN3Q7X4ka
xXI6QcQR6ulQ3MM0ePpUFT+YFrni4rzN0tJPg/EBoiRhC74zz5XCLzsHUaPO
97KXey3dt5bdT01bVK7+PGDdDHXy5Xa1xIJBvaMPiVXgUF1sOW/Gv5Geply8
aB7flpK7rEaYcN3/U/u0Dw129MU+HG5vDcrqzmra5D7s5VoNlal31x8HnaBX
fCq/O1ip7p3WG2OVcrfJ2WpRbRQQM14B8XWZKg3k8byI57pUmNfh3d4ZHvMv
GKUVjaTSxlIIgaujOSZV/ZHacGr7VC1xj8mnUgJSSXmqKSacoO0yzEtlkp5m
MMNtkNwoz7ZdFh0/hCcF+/3Ada5YX/hWYAHrqSBuHwzCqku+V3bBGX+wHVgl
WycNh20TOyzO0BXa4p/payHVTnr5uhhPlER2J5XSvJXTmdqjqA7EkmSM0Jsg
zU4KRNvCRzfjvsgsNQyZYRpEP8596EyshV8mOcC8NTf6yz23DIOzCTj/eYZl
4m9cb15UAIFUfuVFnFWawi+4rfcGjrCFJxYpICxx7ZfR9i2iuZnFPYSYF1BS
7kjejoQQYHT4Qb+8uSr7ooHop+MWIsBEgtoaDFOa9wjaIEQ3WDRJtao6hxrM
yViORkC3JqOvaAuDmC59TNd1KVxMBms2SV+nqlQT75y1HJlMGGwFy5IGgBpg
jvZMgxeJufBfK1EBFtu6mdWm6ZBFmMpavHZrY14bnea+2VJ3x8SEhMcV07r+
50ctkxNf9Q4cubgplR/cMinu8Se3VXt/Ve6XgRcChhKX9SaLBVxzSyG6Mngr
fy3ljZft+K+4l5Zy4AY+50kysN+XaftW/9oEX03YdrrN9nXJX2jWkN2DmIO/
XmOCyyMXsWy5Ssa4xFXrJ3HglE/rlll/LNGLOjDe3QtT6+gImmhIFCGMVJhX
PC/+HDlovk3vqfChudbGG7ltErG0pjB9SvYKKS4TW2f0irFguiLyZlLYHBSJ
uOS6o/3rGu3u0TdAW3R0DrircGmH+y6MLT4S0sspvzDf7VZO2pQR5MVxk+K7
HAcZxcZPDnXy0kKITH20zvZ4cL62ld/uT43Y8wOJFsOBft7NJW9FmoYZPGeM
amMRhuDXkKEyQYpiGXJ0uNgUikF/EZZtTwgHiZ0SomHJTU2nFGR9wuJ1pfMD
upxMbahye9DQW++UoS4d6GAh3vf2rxMQTkDP2wyNkrA/01vYCnsiJWyLT9iX
b8pOSR/AXDJh3fCHujYWbwGocFvl+a/5Cka0sN2/aDXvLDjzSFf4zfp74sCp
nQJaCU+AwkA4EYkVjt8A02kyMLlWc56aRGTYkWXfMuAWk4DxxfBzUv3MRheM
rrj8m76sf5koPqpFy5H6mDboRrsoqNCpp3uPmDpHUqS0mgU99QknMQ4gt3zg
N41unPzpJTE+sR5hs1kBA+DPpg8bAvEjnUxfgSukxC8GqkndMySDnKC+B+v7
peN5uOhGcWLQ98QxQfp4N7ldDyImH08vQydiAhn6No1VOrpdT2lqvpOgGsD7
WMn8xUWb6mUphNRUM9k2jBRUjRqEl4OIlaHjR322bhyXTroFlkgvnfagjmSD
vxhcGqjuesTwMSFzq1xlqPuygFdfG80LqjIL2Y5hRT37mAojsTk+XeclZYZ3
NEbZ8+J/fPeX/QdD2Td5cTGPh4MoM6gH6iKEm11lR4LS+7BmvijceKH/BVVa
X/7fh64UiWT7WkgfajfbPUrHwlC9R5H3n0e2ABn+KCEgqTYj5AFAMKy8mSGj
/Oj3aQov40SDAno4EweIHhDshLJgEBr1zm+p+YHe0DdyQ2wSkEANDSa0/hz8
wc5+oYMjKqy3lqLlTBW0YGgvl0hOYYpztQj0ZFtuijs2AxEtiknO8+kfF3Av
7Ah4bB2GoCTZtG2YK6pF48st0H6esSCibKJHX0VflU1p2QgLkgyPWQ0vQu87
AyDi0dhDOxt6O4DrSXnlaxAhDctUV6oJjs7pONPKTEOOAlHc54p9nLa4HnZ9
hmbx4q2MjLX/AhJNyBkbf3Ly/kLZmzuVfVjLb7W9z+YlwsNc6xMvyVIaOTgH
tN5yMkw2Hy3QvhPnv1smx0TZZ4HxKoP9WYm8obe4EmNJ7Ask7YGGH+FfO3qr
ro4BsPzricrtv3BWIpDj0hUCKaaBsMNQ2+BTcmu2NOpgsGhyQJ+2hBFEQ/xX
yrbYXNkfqJfvbmNw9NsQe8d0TutxNuSJkawV3qQptHSpKPeVYNgdet5wAKhI
I/zXP349pYzOvpDeS7XGWX4rTkFeztkbpYs2wWum7T4FxqyvxxNEeIWr19bH
02hHe9sLDGaEhoIUGVmqqSILyCBOSrrVzZuUNnJOmvDP6CVcvlT5a07VCgqX
Tgo72wK/H7weK1HS0QP52c1WHkrTPMd2Dm9GrswUS240wgcBOyVclAQtRRyH
VYOPhwAjbh5dudX/bv7HWAb0RALdbrazhLu/765EK4UTfSXP7nppStYvt0k9
VcrTg5Pp+oIM5C2LH87f01UcGuNQ5ujiIA+fL10cRtvBQJoN4x274fUwNL8Z
f3xFgUSH1bngWZWgC8zce6kQhJqgDwo+zC379t4mV2UxzIg365xv2oLyo+Ju
n/Bl9udKV7+3w4QyiN94RaEyZfXqvDuY01HU5AEyt0ZSUE2mNOel89J8kRV8
REFmofKjAKLd33A168+vkuRuhbYtxx3/gqVQGqVXlnZl5IBeGzRMYg2DYRgg
xf734uJg6V+a0QKtKtr+bPIu0oqO5Xk3i3G+kGjqPC596jnarizaZeKZEX3H
LXnvyEgmHvy7E6OohQ/QT5cOVzgnM3LtUmR6gyPXmosDuYSUK3k1WIb0GFZa
sHlAas162MKBaegCEY7GK++Cb1z9l5UY/ZeSfbcQ21pJi9N6Ih4Ki5F2OsMy
eEwKEa1AHB52T4yjtVU2VtgOvK1xFg8J07gORmP86dTtt7PVGBWnGCzV3wG+
oVh/pWTNLS4dLaUgsxIDGQL4+DBumKnpTkBda/9TTLb9bDPdrmUJYqVtfIcu
DFJi/Ez88Pl/v491G0l/2NxlHwEhd6OlfPT/K7fixtoaadaQ/yO1SpurfL1P
dA8RT6G0DnneX2CRjopktBc+UtBfQ+CX185zSzeUB7lXi9h2g+M8r7fOncM1
SGr2nCvqZMCFVP3BL/DlcX12wdyi9WgrpP87Z7XYkKTWsfeisaUOE8cXXZ4S
06w2L1gocJ+NSxpop8558+pESV+AxtEkSiD87/I9FT5mOYApVYOFDa6OaHIv
A1XLAj6Fb8UkhkJjdfiaQfWPQE65uYLFI5D4WgvydgA9tpnWog63X6wOmv5P
wvM0R+ghQ99ikwMemayVGkQiXXxKS115RBlyx8Gq1rbqNM9w/QL0czOkRsyl
/q/SbewKcBhqUPsyBwYJpkED/rGgfCvfIBOwdBSOwbB/W0S9Sm3Iy5R96FDL
LHQ/FTo4ak+ofL/L3m42y98ZBS2QwKzDg9CDYqjzBBCS1Vj1XEF1eiVY6WfQ
dEA+ISCGji0Fiz4pH9YYE5UAhdbfTSIwPVDhwXd+gRuPhj9p0Gv689Btgerx
/GRICwmvKw3VVFChR2TA78irJRWNqGNZEZkO3jBfeKG37xnj8TbNVuwY+ksi
6Xmi4/eZwTHJ/lXknTHumvat+ioP90MHGnbCz2YpeXSBCGive5G3xBN1kmh2
Pt5qrVjROk7Y6w2O1v/GVd4g2lgd8gnz0FzrgqGzYVkRdnYiUzBwrvl40968
qjDlVruwE8tLHnJv7BC7ZKPvAjf1l4336v09CffAueG2es1hDaLBiJBuJnUs
aM9GsQHzDqP43MJqU4Wlw3SPjqrugf8=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1L2GiZI9aKZo9PqIxadnGXzw+qT1M8uSgcTCZe74c+HuVzE3UzRmW2cWK5Saivlke7dOu6bi9NwUarMPRrHdl2OXqWedoY/xriSQfGv04jGodt8Rk3dm8Q0RUAqBCAOuph0RyN1SQdHrhbuN28lmDcEn9jmvurbzCcPd2GFiwaGNJ7Dyp1l2z5xzd8p9DioIMhbNE+Vl5A0E0hb1TDXeGDBtICgyLDbs9bk4YXqAT9NprHRsItUcx6eUtBTcgI9juhpahvWadXwy10Gr3kdNw4spYyuiFHMxGDvybj4v/JVOZdHLseCgXBNjhyPQuGXO4RujLqz3hEbnIh3Vbt1CFWl+ZCsTzRtNM/wXxcM+dUZ/mAk5893fm5A2etm/ImqPS+as4Lmdr2Ga7mSrkoSw0VEg2ocuWsqDtkmAIqLX4hRq++xnkyyFFXeemqDknB/JuiJmIG9XOoerM1tkmY4dVmTI4tCosh4FYqJhm+iPucNNiZeorCo6ma8DdYdEKsZX/dmL50zXzMUp2wvh5u+t0m+WVc0gsyvtAWZzL8wbcp2lPwjF+hiN2DWyJr2bPYOom3wdrx4qxChO7Zvjb74IjOjhwq+X9hSv1iv2Rvy8nKyb+3eXjQi99a2fjc2h+V8ouI8kphQOAY8NNokd9E1xooL8q5nrpnz5R4KN50I3QfRzgQXMQv4KnhRfJ4RScwEwA8deu2pAF7lgSrLLCLaxNV1nVcloJJlys3zF5SNtMzlDdCLrxC1wkVJ9c4WwFDbsD3nbVIClOa69m15huDlwTZD"
`endif