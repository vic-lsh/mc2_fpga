// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hFR+np1fwruQhVDJ6jRW0GToFhZJzy9URj9mTHrNIlbkHgMDIvqh7yxk2tev
Y2Ck3f78yHHT8eR6idFOekKFNXkO+bzeP2bw3TIcKaZV+4ZAo/P9Ji1V3Pei
6Zq0AWUppBYurRxQbF8VzhsnIMN2vVWXNUSwKAdTQseDeHz1ZdbZjnEsUdWn
DbsvfF6va5MtCuYomRsr78OJueUYRIH5yWf+Jaxi8XJVYFU7LsnSz+g5mcaj
dbGbfIDEDneF/13Kx+5rvGT52rPmdixifdSZoXfGK4PQtFgizIUAm+KmTNrL
f8eSeCvq7g0K1pF18Nc539H5GaH1FSNQ2vPTHzPYgw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iFdibzR9XOvYUxKj7k9M60b10oGtLjjuZpiB/9ZlvmXpv6LKwH5nOAIbpCnI
U4l0qM7AE6ttBGumHPtijt1Qg2WtTatWyYI2y1RyZva4oxgRYcIuPZJIKPll
zyUzUjNq+/iFKOltVTtAIsajmTG3IObiViYpFFBXKkJ5f2pej0rlCwioKlWr
cStOz9Dk3U6YbjkBnIMLDazXGW7HF5CrDfHWMS1QeIQL2aEg/fkRZCPXodUN
DfkpH+iTkAVUqo8SgrTC2mJcwtSQyaOYwRvkizu6glWfM/R9HQz/Y7ztneea
QrS8JfuHbkXZmoQm4curRCK4IAnuBSDU7ZUHMndQUw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ctqA94r4QFdT7Xk+fv8YMTVwRVyrwJ2mgLqIhGlcloo/yzWC0+c1PDS4I4yf
CCkI0/xz/ezxFOYz+EKfm5fxVA3uTDxJQRFNCNweH3iJDps9HxU1UMWCc6Fe
kHOTHFUcHNzjsiDjUgTAV8I7OltY962ZaI0yNPqKNc9jkxcyq7/AUwuv2kBk
ktL/0JDrL3AyWOHLWtmEnnnUljS345r4raTK3+qHAwu4wk/NcLgmaFp+l6J+
YWnbhg9XYxsqlMguW9xBuESPFXl6YN63rEWfdggnDA1MyHuvXo8qDI8ynof6
2L8dWhAsO596HyxJX3Tl1jCePFvo5eAoRTKluH1UnA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lugbhwXafSPL45hda4RUnN2agIQRwGDmSGdj++/SDmuZeANP/CxMUeAbeT9t
JU+ThLhEw1/2yqEmvbG809EtCJeOYs7r7tvrjekMSeu2lImDn59EKwUf9OcX
yBJCDZVX7DMNoF2Mtk/CRHGDNMItjcik8jwxlLUVTkhVHQh+bO78sVU5EY+q
QbUIN2NHvvYoaMgzZ7rhgV1E3ry8RxuaL2b1hW2EfFcaHdqQxlp/7ZtWeX87
uF8L7/eZoruWbmjyFg5vhnArKL+3e13bL0ap9UPGW+vT5FoPMGxR6JjA1JdK
mYPkRCNGqw21u/h34TRlVbd0/3igPmhSCbssRjcrvw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h6HPtWz690J/MHg6rVn2H43mQBungZH7XrFIxJAimBiJFw6kFi384Mo2nlhr
FjarSVkT9UbIEnoWqHt1QZGkrt8UDsKsNfTRHI0DwAOOTbpkJXzAqQg1xflw
DlAUSLySVtab2oixGlGRDcUKfawPCcxw4O/ylDHHvPFNyYDXtVs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DrDp9dv0dr/6JRObLqPIFALIKT17mM+cRtzeH2gP6BmmpZ80JLYI6OQDu6uL
ca0lNhTsCTG2mkDiQpgMH1AbPp/rpq9I3ZaOCJWGUm2JiovL18cZ0j5f00Ev
J37gj+FZt2SPG4U04DEzgfLFy2gWgtJTnVM0qo46jCZbmQrPxSAmp1jNPdGC
il38cgDa3lKoDK9Y9nEa2qmUiVuUgASomfGle79CphyOb+UklmHXUXTklyaj
mYn+kgru3Ns7Ai8Yqnkbrs5FBkWVGodWLGr1/hnZdj7+RIiYBbGOzSskargh
PJJzCsAGRg6XzOF0MCH/IaAY9FxVdKtrnxrN6n/MxV0wI/qZbgzVYM5Dp4CH
iinq6PjmDh7D8NYgxwnfTEL+Oc2rA6yWuR9T6FKQnEYQaRD6qGFUqZoueLaL
NMzXWyggQSfZKHWYmUdarM/Y3aDDohAsTYWM6ZYttDy3+fTd7thz4lcqY0Ir
Xbl7vRFduL5dCuASAIxU5i31uPZ8T1iT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MSvkG0ypcc0Bn78AKBn8iy7FYRA+0GnQH/0/gNrr+VJCI2TPHkXrgCKStHFm
Trdn0VJxuxE+ZVM2P63mNv+ES52MdE0WlO3fDzXl+HIIWEKdGYNddNikK6xu
MEtGr2mDNH2zNhH9Sn9Y3yAhUwsYxVl7D9U/d682uDP2Swcodn0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qZtC324lESmYauzGpP6+4SZIz31yazTKRTHsA/dUmQJzLU0EILUiwdXCIAYp
pJhTMHpmFMyBjxKbXA0M97maYUsmjsFZozOnVAlNyIqYaj/2apkpx7cO5YqJ
JmCET9si5eKTUlkMFm+kI9qwYtrjeWKWAsND7YozCQ3X+vVYKaI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4016)
`pragma protect data_block
PdUQWqseMeHoLeV/RjBC9pvssl/5seCcyIh7/+IoBl7vBNwhqP/FNezoYwf5
LAFzLeNtQkXhjYzEBuPKvuSWIpk4Ni/6k7hO9Ss2Rqx+6pJX7fAzZppAuTAB
kb93xCOUc0BQIfyqHtymeZk0ErNcX+IbU+c5B1HQGjrctonTcZtTBOKj5PkJ
LJBTDmKwDVGCYcVv1WXLwUCcxYehfS8/UWm2g8OFX7nJAO/BNYVzxGrx+WdK
9bLQyTtiV9pe4DGoPN6nr6bpO3woI/ALV1IZZzMDNwOc8UVLm8fipfIyXVjn
iLn/m8iw5nVnQWCxnuDyGu+fRTO7gLu0MPd7rGdDgJr87zIEklftoywC9RmK
Torf+QBh4wQ/5iKtuIFkguNwHs637/WJKKgmhE/N57/plnOsH5e2xRNAnb5W
03Tx3bM0Z18EOMiMkfFJ2hK55ufg6Jt2WUbrgsQ/cPmoBDnEmwz+pXMThYQo
Dw3+0mB9HaAO6S8YTgC0yI3eVlpEzv/G2v4wnd9cvF4oDnrp1DEgX7IhJYmb
EGKK6K53OtcRMPOcp/8nZLGXYkb3GD8MSMoLOTOo8gXouGj9sKHONKeefUkE
x3iyZxeXRrLPMeCfifWPwRGs6WqiIZu9l+R8AM35f+HUw1v5l29ibrbm7meV
5aDr2lytvrszTiuljn6dqtORhgXoDQpH7KkEFNGh6tOd/KT4Lqv8JNuxf7bc
QYJ4kxkhIkFGxi/qDq137L4tFvlz6MbjUBPXeeW/Az/bN3f+uyovUFM5TXMA
fJG4WGUir7Y4P2zwBI6MCXb6I2kivFTyaBqQZ5fEkcghNFqpY3melzE9+vpi
N1zUYka8SzPglIMpsQmqn8BJVA6yhBD7vjwfSeoVoDOyYXKkuhT+KhuUYinT
V+WR3tJslkq9qeOUvzF8GGSK0HIoWqUFIc4dOPQjP4YPci6SLngcixXgQJ9l
oHKw5x/y/LKKFpHE8FTnHGBG/NM1w+iUgoKr/jEumWk9BDsnyYutq9AVNSno
p/LPxlkpdvrzH0sJMhbzOQ2kcuyez4lodNXznuJ6sY/Jgl03evG9vPdHNr1E
iwYaSktzxI4gmjRnRDwI+GWN+bEYxuUp8BHc12dgbM7vYXxVTx/xnOpXe6uR
Oyz3hB0oM+Dv3DL+pDRb0cVyIuXLG72HCdxE9zjSz+4D2lM9upta3UyqzpoW
9Lepg1WT89+VsXYoRB5hHWUIWZi9+notCBYC6OknU5vk4Qt/G9hY5DmFoeT4
CD36X48cVf0f4Bho+r24xmCn3qIVafcXP8lAiei4oqYq8QVc6E3pGmSdngAL
cA81vAojwdc67Xg8EdSbgOZGgCgNeo7uwq4f+TLRfnIzkx+MruDehJ0al7lT
tVmZdb6zGKbb9+X03YouE2QNedHxreL0du+PRVI7K7d3y2enxSSkpUP6eiV1
TYlHTNgJuKIAnWjQmxqLNCIG1o8NGWnNZniWJjP3DTFQClFzmfVcYC5bpOFB
hyeY3KCf/FA8QBx5JhDW6nh47+G/p7nKLdhguonAW2xZTW2OUZaaqM7fj4jg
L8buROvTiMjYs4f97vxgeV3iNFA08ftSDBysgo1vCW6q6n25qcYrWGoIMN/y
UmNygbmWfHZBx7mqqucStwSLGP4iYVIf3iQKF545kmf2FGJXuB1Rx4mMn+8M
bSyOgtKmQDEIFTMc5YpVcCkRZzMI9+wJodIh2mO0ug2WrmUGrXSbXCx/CrRs
fNljL9cpiQCk/o2sK74g+y1DMNuY/K+Va1yEX0+X5qlYA4cz+Vd1ya1I9UuE
x88rS2hrOskR3ZjjHbWU8hRRtLvqCv3iKt8TYJThC3ljQse5QCKsl4YoNr1k
mJQ6Uldhg89AkZzksPgj5mZ/q8tnwtY0QeojaNsXEe1aFOvWasPDrx4p80rB
LZMtbgL8+sVUpk+btNt1HPaSRpc4hfPiFT9eJncL8MVirGMjOhRKeAbE3sV1
huMDoy4pJK+BJtJAZphzaePNOsCyi217ab8WgIFuTRLzBVxJdgmNGVtt8nx4
xiNxwjSYvggEA/XCJoTuqHmPOetRinPJGrgoZZzkq7Tx0g/0QO8yF81q8CWe
ItkAY3b/7pARzV12ZnLZV6hrqJoO9gcnIqx8PdJEGXfljXLRNOK6HJkEt0kx
eYTtfyQ/mZSzhzd6KeFKeNWOUp/vlGqMqtTU3nsuXcmfWtmIOvlpE4NfRwKd
V+8OBt7yFkF47iPrKkxJJXZZEJRJ+DR410tdfb1o4lSSLRLZSi0t8/9r/JPN
3/IB2njN4qpN4NPVgY3/qq0ITOC6FTslDfIHaeb3F8SclA/eE+TjHvTL4GDq
OQZJQSL13fLohRfYV0RHf24+hVsSZjPnLylhYp07oxYnoHCBhVnlVfL0DABm
U4j4jP+HlAtOnuA3jFU3FqvS4pD8AGYBiva70XOd9y4mx5+mMflHEjcaTJcX
NfR2J6VNtNOlHL1Lv4eUvQtax5JT9Qd28rTHy/zEwPKhFYShzzanDwh6zOyD
svj9tAv8uBZIU4e0zUoEU3hURs/2qSl0kZSCZtU32ALMYgnppqJnr2TjJWjf
WyCiltrWzIGyy9x2x+buJHQv9Mf6DVbGB6cQUmnzm+rEptWtmSfEgEvK1W1n
86xnYXch3LJDwYSy/0kLyn5grjtoNf+gG7ScD/ltEuuucxWfx5N+RC28Ok9y
P25+w4d5fgB2toBVO0kVHGrSXmz+aWqZfvcJKO7sjpRzrlhnvPh4OYpKR/fN
/GaQ89bfS186HRK+F/LCIwMLotxZ35HRLfDSmjMX3l0VjiK17CgdsedGR/d9
z8syVzj8rBW5Gb9+CwSAvXs/gCCCntyYXYvx95hLvG7gDTlTgKaMpW+YEWoy
o1d/5A2vUMoZzmFD6G6/Ezb7kw4erI8cPnEQeOmf+pdXWaBWo2e5BRfMTErO
05VFfOi+YJAKhtA0JAuiekmMDdmU5o/DgcOP2sjdCMg5XJADMeQdVsPkW+0x
D6mIMIt5qiPNbqvj7xEmIc7Z28fhRqB3j9TaSRRJfN5mSNdKIYGfLD5dAVqZ
C6csywj/L5yoCqteZURwybc7E8HvuW9WN00WynE6WCbjl1YBsq42nYUPRHlk
C3kuFtDjaeyEw96xf0FJEBpDC60FyoH/TqJbZxANgQ+9KKWMeIZVjGO5KSQ1
evfiPF9ZkKd1A+pv3dPFd7KV9f1HzWoFawinmLDyIVdQn2sR3LcZbGoB/5EY
itdpv56L2rDeU/b5rQUxTUW2MiIDSS5oksmiT9vtSIU1KZouKQMOZrM85iSB
6n42OFIUJMpvm2Jk20dc9OxsN5XzTzZstDK5EG1NxvvPoHT4j3kJ07qx/SEF
i0hQVDaV+tuENSaH4Xq3QAjAnKnWfSD+6xTFI2XOGNUIzTehx+n3LnRZNnKM
wP6qu7a92PQzQjmQEjMrhlCEFnVSNV0fmUx8zjh6Lz91LJ+zk2t1okzYsF3b
NB3P/AFZ32BemOruenNPdndEhB3TsRGX2ELVjHHuDwDbgc0cQN/7KRZHhPmO
nGfDt68B/81asoJLhT3C7eJfO0Lv141rgkONK2KuQ3Sw0/lOpq8B+OSUxW6c
2DE0IRSKgHslKuAdk8u5aQGUUNCV59+PB3uLHOg3XMQBnB+Sld4/KhlX31as
DO8l0tWWzcWr42uE8aMQ541ozOT1fd1PZUFUbs8tFViigzWaQrkv8Q2Gzdo8
bPVZaj96zugIfGxqZgMFrZ3tRe96OnXc66LQkjV2/xmHsFIDIo7FRQyItKng
Cbt9emjKsT02HDVui7pyjg9UbswYgQiMH/WNCgNY0AisgWWnhHq10jCq4LGm
/pmvasPDIGRvpkFWjxRidjp1nMA9NusfrNAs2iwKfTb2Jf1stmRP/JBXwJdr
Ijdvr6CyEWg2+wS3ACt6mmVHXxrGP4J9kUIZHUT5TbfV5rs2Pm9S3fWKojQ3
WdFZ3Zfi3VGHs76hb5+Una0Ecv0+/c/83JO6zxvm76TE2Lctsyt88UU7vkVS
Gj3P76/m7lcWjTOdZ8t2kZMcuOltJCK8/2j/SNTZfEGId7S2FyvOcrt3uJIM
Lo3ZAUX9CK2SausOgRT7CcZJpmJa2nkPCbQRTNzL9eWmIW2K34FwWNvZBMJ/
z81iImoy4bC8vJIAdq3S2AeI6q5QwyIQ55ZJ4FOcMOEW8A34VjKvEaw8PA9Y
VCrOLve1NZbfVl4TY31U4T4CHFnEIM16wLtm9QmUHEmi3B6SUwm86bvwA0e3
jR10IAZ9nSbaANRJEpeDVyeYRJQwDQiOMYldor8LPtoER1MFb/7hAWW+GY8v
hfdQbmcDxWXaQs+ZPUw3OhSkwf6KSNX6p9R1T58A5YqovnrTLpl8prFRoD6H
CyGrHeXvhVD8tGK/m52Nw9rtLbSmPiyvFwVVHO4oqn0dXd5Q/UOggOlgx9UM
FywtMXoanJPaS6su102jtUfs+tOGBZ1sdR05npD6KZNMliyCtZjapn/S9EC9
Yekjhwxr7CkI8lbx2ee2mKEhVUJYORxoPzY11ijHNauTMhkGRtx7Ow4RhLvG
bldaKLVkclrzv2rmJjnXk0DxXYCyYxotH4N2d+P+rpE8FNoIZNzk35ILWg+V
YpWOqxTXHBPZVSX9LdqWVhgSP9/GP1h41UTkxVUJdcyqu9e9njbW4gz/1V3r
Ny/TJN6v6RHCy3cM1t2A5cjlV0RpOFZGx4Yy1Aol5D5ZpTVNl/739cQytfeu
mfh3wMXsWdUilhU6bhcn2+qkE1m1LhCrwzTflG9dG0SKVB1TdczQ1fZA8YD6
KAv94BFVL/MdsMNOII8n5E6fKeesIIOkuUQOUlOQLpWB4uiGkhEgaKXHWioM
ZDPOAFAenEQyn7qukKlOl27xlDxlqEzn/CbVRIfysiOmafvWsMWK2MwTKQg7
/3/CjHxlQLTs6SDNBWiaYYeMv2MyU0V2NEkaSQRe79G8W7Si3pLwYcqr2bz0
DHxKiQ1scLxI7jvN08rI5bPGyKQmj5RbR6gucFw/zTOdIgZWrK1yMKr8LZ+C
h5nJeuAaBHe9C6PSBXnhuuSFgPaN2WE/RowMQLne0EAoswMFplF1Guo7vkuw
7PSoFsWjn+eJlfr+KxGrluurqooKa7qnKgTTrC6HsGp+Y8e6x5lQAxEMXIrU
Fp/NeJsq0/IAjbdOnvE650rx/FvG/Xm1rGrCrR5VIKV1dKxrkCsqawVS/D6d
reKgFzx5l5Iupcy9uzXYRT5f6WJdbT4k0issFyuDxpP0kmuh2y4mMsqZYVI9
2sBApsmtZ72aGjsgNZpH1zga/7q7DhE+rA6EoBJUFiOioVp5LBzuTn7qSxWi
LNkmLcLqF9eQ7v4=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wiW1foC8HHXdlsSNQUL/hOnqTLFM/mSMkPtzxUsoipnDBNi9CBmTDccvTZcuT/aZiLVIjZ7CR2dDYJRLXBY98vZUfVkwCGVbaDa87/lo/7F2L9M/Fc7VUOzT1WvYeLjJxjVJPW5OrVyBGbjTsbz/Ha0bBD3RIFHXSataT3ruBk85MtVlWi14KdT6UrZvIoWBJZHGdMbDxMIu0t57w4krobo6oTQ7v2qY47hY2ElJZ4hHkAxw/XGSd/t6JATC1SnyYGST/I05Dwz5QbIpUqko6LH3eAr75wzNnVvByFNceqV3pQAhAbF5VrrsenMrcghNeOS1KN0rIIeLuA8KY4tARCn1Y/xVLcoTg3AlSaOuTAutq6pFpA7ZvTYJASJeK1sZtbHTOVKVeG0PazC+Ckhyst1bm/CVirD6jvYH7Fr4zO68NF72Is5BC4IaSdBey4ucZ4LdSXUyHoU5FcY27004qEvn8MXlNgXzl1Quoua3MytNtSm/pV3KAnR75ltNs8/DqYjy6ApITd6JyRb5sMxLJ3a5E2R+Dxz7UY26bulGXygTyRxJHjaOFiuqSIQJnEN89nZuSlr/WrmaWkvCbRwpBSUkA1IDIwu4PuWXIWPMmbmj/jbqnHABazdwqzx7PIkVh38xOjNb0eMmekeLwnYpu0wd289tkFrUacEnTciZMQoYr5QEu85ztn/19YHYb3bjoB1VWzvorUoPTfe60ZTfSUusxYuS0yuuikYbpaOI8DivPhJj5OrsWhGnTKCKdPEu67OzmrFgbos7gIRMQi1U6hX"
`endif