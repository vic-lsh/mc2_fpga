// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
piJhNA46Jyvxv2RS/+dKAvYxl6YAdylTuEZESiQD12QJmX5IXT6O74+tSWUc
kM6bNnJ6zcPDLVB1uL8q1x4kLyRnud4UF3ektFoWPOc2Jy6Z3/Hc5qGf/Sg/
K8d0xg24esl1doj4ENezDFers8UsBvM+ZolhVwIgt4YklMc8GTpUkPt31qXA
WTOwb8cePHHj8HYKHMUGx0g1IeNFlqZzcdCik46bMyylaOG39/oissA6Y7AJ
brBJ9jQiGNSmNHvmEtvllKD1BUTLpnroOMO5D90sRnCzUAePjx1UOADKghWG
43Gu7ukFS43XCyVsdfqaNToL+nn9l3ne2Vt0hpxzJw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fOvsNqAEbVBTcl9eDaOIAofPdbbz9uOx7fHUxb67rXgUwPXEOisOZlJQjpF2
R8BRd8MAAuStEQNzBviKewwmYefjUQlBPNrq9yujn/vkBBfHn9xsD8lZWdB6
erEAXbzevRv5uob2BwKR95oL+742D7GvNHvkFFmXdeZSsjz/W2m+KmhPWu6B
SMalCJJX8SGLYi3qCux/uzdJrDebWTTE44ZxcbKFfwrLvYYDLS5svGyhMvao
wlXBvElNGldiW9QeuusLxqILihpAvkK10jpCryLivavYxB48zfa9NSIZFxs1
4nJfAuRI9fUHbwdxOvmM5nQuQ3wFQsbvkWzNouoqkQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bfa9AFQ+yJURRUpMpx9ZRmQj9c8dXZIYXHpSPxvuscEH2Tgp/bKOaCk0+XZo
gj4A9LWveKMZcLQNcVt5gLtHNWmXkVct40VrrApdgN7zPN0LtgCP88HK/eO+
Q/awFEoXXRDZDRyFQRqJCy7A/BXZYZqaBIToLNNmJwckR3Q+KJftyEIooeoO
JVqHje7+y3+ozKVL78e7QAyrpj7PInOMWs8cDnYXR5JdswI5K8R2EGMn/vNY
dY6Jhr3Obj/9MKnJ3q499dFdAAiMl5SQz1yv2eJgIhaVgsHyj2VhVG7nd4fo
ryaIKR6BOU7btKjqwOvPKaRuyoZMh2/xSMR76ZvLeA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jqZ3GRirkgOmB7R0uWoas3af+3dp49tzURAjAfymE5YIBGeiGiJLwSrInsKS
tums6NMDaiFTbbo8YArxEj8EE6Q07z7jy3+bbbwyJAOCB1Kwkpkp8f5G3jWx
CgyeT7oHHZ2uGfX6bfLXhtmK91C1JRqso9qy5D1Pk2sM3HMvpsFtaKEQjpYr
W+nkomCSydhQc6bzERUM8Pvz+nIm8rpN2iJgCMkA2oYCTQNQ41Mv7ruKsQ/o
xXsVH1byNhuUrAKx2RKEv05Sm5fphx/sju+nEy9uc5jeDwjoy6QHEA/wH6xo
DYGgDHnCKKR+C4eda2oua57yPLq1nwHWSuPyycXcnA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AtjJBTFh8Tv+ynW1t+4nMxgDlnIrkhrkFi610A33f+AI3zTbKsgnnyvqN0gV
/9jWli7ZZdZ81h2RSHl01X+Ddhsfi6YKOJNQdYLcaVwhxDOPetndMsABsZOc
W4SlOpOoLrynBxZ+vD1hR4j8DbkO93NNU62aRCRmNid8LoUsnAk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sekjDUvq0Y/BCntQXaRvCYBwAUlOfdcowpjWX35W35xgNJiErYHt0l2tuggm
mOETt5O9bxhbI7R0mAyPQgftKjZwLM5lrDepPPEe5oRkugDbuqPYoJudOM4Z
hH28R5aAeNT8EAJaHuwhISI8wrhXl+64ayXZyeYGM87MNBr1mP6kesF2GKBj
kJETQIND9c4sKFIWI453KfSCEM76QGd8BpzPM8XXxbs+425YFczAc0Ql1+Aw
aLrB8glhIY9Uyi83HcFUYV2OaN08TB9e8sbp8HqyPvvtmqHZXARmeefgT9FP
6lJuyEmerEYHontoaFOF98DXxpBNop/dd7+iaZyUzjLGuDhoASGsDcKSxIjK
I8pJIE+KjYXfgivG9UbSjqAMI7N7tb6boqaO6Qn49gqeTzCUt7UAwuxyGJsk
3QAMazom0JSC6QwOyPcQOcSxZ2j+tLg0rcsaGyaAyFXaxmDG8hwbq9xxDOnN
NbPiMqwCYL4DiHMBR4F8kMqytto71dnv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Cxz86lOoSt1S2xmCW4atCu1oTMFZqcR2f3+VCsY59TKCsNIJO/zK7ydfoxK4
64dVgJnDSNDG3ItoEXfslXnpQ2ZKY/KRpHlvd2JZNoTMVklrYftmGJpQXFlL
RJEDj7m4oBA7tQV9DKcgLf4EiwpFd2xwTOsjeAPgqBM8kZ+xv9Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ErBvDFcE+AbbuY1v8Tal0fJE/kj2pWFjPHurDoSkzafXJwSAp2CG7BxJeulH
hq4/NofYVwi7oYqaXIgTqctL1uNQEDlfsO/W4w/DnKT/Svvcczx2GlQefxzM
ytNlDgaqViFKpgquvXO0T4PLvB1BF4kTKgwOPsjR41HEyfyALPs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7872)
`pragma protect data_block
RAtACbHNJYZNmo3f3jyZaOwlTVfBfo2xHG5AJDluBSrzwKhsqiq9AOD8fjfS
tpsA3zPiq3iTTC7hQnDP65PG6zlBv89nOZhRxtFvJtF0kMUQUaXorX/nLAgN
rj0Bsz4UzgwUCFVmFZM9rtdZ8qyhREaZUUA2Xxhp8SK54pqPFRxLtJLtlrKe
B02mQ36hdhUPOlTdhxIX44LLrYEv6XoX7u2bZiCty0uct/v+YxmBWscIw90A
gCd8gnr79J9qLhZwXuU4aEfochQo4kcsrB7mLStGjdUVMOp7pZze6gSiV2Cb
Lo9xeJw7PlE9N6Txs0i7/fgdQj+epxlGo18W2anEk652GwP3+2c8xqBV6BbT
4/A/jln4ED8fUDV9qF4DEPcV12ImeeZjCJeLVqANi+pr0mkt0ytqE6IZVMcg
yZqzpf/O7U9WJmYDMFOUkr1NtF+r/Mc4gp9hvQ6tIAEPM3SGyp+zA3hVzQeG
qYQDMwf0E8lu/XMYzQwI4ffgVi9Jx86wK3JPnPVQYNguMSf+qPY1HTRMFxit
xzCft5n48KI8q0l94eT3hYC2N/U60m3yD31wUCZfBfoGlD/mNEVpUgW2gtgI
PpAL5riujLXaeGlnMvRygvuyEjy3x/I6uNoo++aeQ4zrT8wd4Zrie7SXG/HO
TipXdW4uJ+ORCv7tO8CvHmDNLQySzXGbE9JiBRl3wWhtSRmLe/NbsRVqbtNc
lTGgpTGG3swX7E/oy30YNWiHXTexNQA/ubErrV0d2FgKh7JfD23R+KQfJviw
NbVEKWf8rNzKyVjLYj57k4smYW3VXhuoM1AlnvvvQDWuUz/7g7b2QRlZkE5k
5R7W+KnDwZr70lC1R4QwEszzkl6EAJgbLO3GJWpKWoQltF+3DkUFgzbXYWwG
U0zdLGGTTozY+ZBojQ7kvQqzdQujS1u0Cqzp32HVnun6CUqAdgRhQUCWRbEO
uBnElj3/fkgVFgzCoa2gKjRuNnJlMCtgsTUqPbAv0AQNqe3oq0gu3R4cd7a9
uWMSL1a4zWzG77cBuq4U8dZST1tJ/J1GKU2wErGMJU5WxNMnt/I5sGswGq3A
3Rw9VIp5GkT+P68dkw7TPn4oszNd4qn837Q/eXy6rpjoynVXBLguejdGJaVm
o+OQc7JSNIGJ1Tdsl0Zx6xauNdcZ+qSoemXoPAJ9QoJRxxcx+ux2q8Ar/4dR
qOdmd2wvvoxLdfNAUGEK9lx1C0v4OoqyOFJqrRvCpOZG6T/yDUtZ2a/FoBwK
E8xX/5DlJRTZmbciLmjra5/nexHIdSxMxRYOWXdrJJ9zco/AeBRjjKP4PSDB
fajENu2pXbCvDnAFD+O9WwIGLYRY6ffDm9ME7mpyBTURVlVYgGeyuxX8jICD
/Kc795mtuXHrlvnty00udw6VlgM/etV8uJ8JBst/gGek0edYTMqSAblmURxM
aB6WNYppHnzTl5YXzrXG7Yi7oVwkF+gfhpHHu9uvkm3FVYYqz33U4pyhrVVW
4ZiEcdVHF2qLHBGQO4wUmNdVlpDrPBSl0vfj7QeZQgzii23aOog7i6Gv5QIH
bykk7rzgcJC3LjGe58/FUe8LCeWsspIV9Fo3zWAf+klUnsXWpihrZo5KYqoE
t533GliXfAQ/+GcJTQv+2Qb5NmliPkgOIJnS300Q0MxuAtM179RqfMF60g2T
uFqT3RLWT3il0JIMBvyI2z656r05zdwkBt7O/qNenQBY4DHlDyTkD0fsGEBP
U+Dty1oqoGMg5zwBBMsgalsT2XUXPhg1tt6qPNZuHd3Af01V4+Tinkz8nF5S
86ApAVqLuOD2aJHYhOpC0TR75juAB5rncfoKFnWCLmaqMrjULKv2OsRLb3hz
HUaF6RHk6HxMSaFYdtWRw2mUCs+XGKbwoAqCanHyIHQbqUnnsquAWJYaBRK4
NNeFNVC5bdyy2pHcR/Zvx8yHx8foIzbNyn42mKaruoNF0PPe3S63Y91E7QBG
3nCeD6VKcDrLhgP7qk8K1yAAi9F9yQt5trmF20Hyx5mF1YrmYOUH3uzg+WIB
2qT7KgRp4ADs8HnPflBSwPf1d+kn5IXnYajE15QhVT0HiQn3QVdf6FnKQBeG
7N8DZcs0iJkaVZq0CJKE3mOeNaveWnaLmSsshNsnIjh5C2rIDGR4EMx2DHp1
5v/u0kAzQjTP/IzlK+PihvkxoCcqWpDrT8/IY3PYjzHUbIfOOFJBq4cSjal3
nBRIylzt3vFMK9qGGqivOYP78Wh65Yj+SBQgIA9wm3B0ENgxqwCJxST83ug0
2X2ZqMMoVvkvYTZmWmIUW3NClU3Y/LRK3wVzAK6oUmYLQVYnrvteE6COpp/E
LYLyYIEma7djud2b9s9u6p3pU/03Jq4TC17c3aF+KrDzGDq/ooERQfcg03IP
5m/2FnXdNVHlZfJP87ibH80ojBgCwictd3TW8e58kDGeAqN518FHe86Np1Js
TBJhcvS4XUeEt3KpuLmorRGfMyZdmza0rdXZc3K1Bm+yfNqTuNDTvk3dTXwx
ZrBY2yl7kp7TyRVAPEV37Dkwj6ui1Q4LxymXJJx/B5VppbUE6Y3BuXri9B1V
a0WIxPSh0/oukNNRLsMvZGLfWxh3rHbR7+oStdSXtQJeFLrKg0YsClngA3ak
VaQw9h0Zwc2GM6ttc5oBCYT3B/FTQ1NqXvyxjnioqbF6RxNGKuHS6h5VRObb
IwpYOWdW6AHIu2g8gWF3RnsF6x8EZ7jykpU7g8WHoJVIWbKZqVL4JdCLhd9I
kV/KhDpnGiSEtncjZbgk/PT1wyptBOpOFITlqKl8uDAOghZO3LM/gF4m1GyM
nuQstJnbYtyAee0MaB+exXAYjWLvl4CpFx2S2cSCC1oe9kmneG89xwdBD9lj
FI76eIYj1myN2T4MdZ2PuD97BjIThFb2qdrQzmgHzHDwuXMcqxV0zRwP6xYN
g3b/vcuA8zju6xlboXYviWzWtOlAq1u8xkT6MARCGFwhm386FBs1vpJw3okS
ZG6VOdHtV8hxFcGkUeckIF4ly1vfmg1WaQAX1N8xf5Dklq1b2sWSs3kQ/4r3
OTbE69yCoSR8RBseVi2cauorHnWJS00jmZSYNYsDAyrmmxvMP0cVU3oljV4m
envfFPzhbiLQdrIY3UF9OWhz4PhkXlTs5BxeNaMY2PqaNIWIxNsI9OGpTn/V
5ab4pPonBDO3i1IOUcfbJNp6bCQ971UcLo3z/kM0SJF1G7yHsDIKWC6cV77R
disT1agMqQtVAr3KLncdpq/BmpY3WE2F7KSM3ZyT0XlwU9ie83Zm6pSoRAfE
kgq+Q+7qRogbFAZVHSM9H/W7/JVZlDh7UFz4Kte4i+PsWzvL7XW3TZapIkg1
RzuWFJ+b+ELjnznxN5N0IE3LdzFHmHEvxAS1u2h8SQyYbbwlaxfcrSBd9JOZ
MZDmvfgx9jrnMhlel5eCizCVbakbDLVQfZa+gJfhMno9H4BiLNCnJ/oiKfKr
WOlXRSYmEnLjRObmHbp04YwNhVK3NwZiq31bq52WNP8nH0BIDWpYb9P4cj+3
HpH+4pi/lHNQ4/6judSJmzt7Cx8+yfnmf2TU3WvUqOgGUA2R1aLTVZSCfpRD
90sNCYzp9+dExY2j4v7yDrUKHUk3jmD63oY8uQE/GR9p4l5+a/G7aAHfX5fD
lrkfbJI+gZoUwV0Whs4IJ+MZCZxopdUPzYtnfGLLrjUgV4rsTIt5/f1QAcFc
piAMgI/BmJT44uobPkPcjqX3hjJxMY2KpE2OBvf/4ZMielL6jrsYFTDLujaK
CQz/xaV1M4To1n/gbTCOxN7RQ+hxm9U+JusOllcFxHo+tDQAYLN1SzaHm+JQ
EPtGXM6P9TqsP5B0XiciPqZ8P4vlYAe65OZyN/un3hF69elMuSfZtUA43mL9
t8JcaWFT0J8lRx6qsUuRtLIkRHXYvBprSQMzS4c5urcUoIM8IEsN7qnDHBzh
ysh8/Y12YigtMCHiOEqRsOmU/jBbD3wsTtbUuLQomTxaipivJPn3S8gP0any
Yo/rQBV96mrVypkPbQ3IBbO8k5Oy1CGjjibj8ACHCj+zCdclRyuinI79+G5f
2XKUmiQWZpxc5cSAzmBXQWe/a3aJ9qtJRO+gQv9kZqvsiCPhcqQmkQ9toMST
Uoyih6qjSzLuU5y/3vy2T+X77I5caeg1dfoVMjUIrlzCE8nH+IrYeR8tK2G7
xNVq6O2cqXdOXlK5CKXtjyR3pgW0OtFubNNVaJHAymkqneun8sznouUpWOE1
tX+kqUwBfOm07TfRVgIxTCTZiJW5BOaOIpuv2TIFUb/H2ivDlvHD3N5b0dSt
CFYtvwPAZByFxUKRjz5a6Ati/oSNiGKacnn7J7+wD2Alb3OO3hj4qYEVz+1U
VJgLlnrGWOmT/fXiqEImIP9MFwliU4jGHhKlk6tmCKD8sczWonPj2H/MAwTV
KvYC4Ux5Av5z5XK3xVDd24tdFzjnS0qG/J20lpHswTEAcX1k4WPX61WBX2Ad
lt7C3FBKVO+ImFPtiDbGj9oyi3QHxCUWzmKjr2OVBvrgEiWaw+w6ItdqvEos
vVmBuMZmxmzVyJG3xp8OmFYVtVLeLoIgKakX2dDKlqtVP9Whh19MA7I/7yyY
5EaML9ZyWQ7MBWzUrDLBzQOvVlrxP2ob5zXoJiBSjw6/9NV2fp6gaPgk9v5W
Sfk7KJMJQZRasc4WkhC5a5jBL7DBnC2RifC8CWsYsyh2pKqSinM2AEnv/LWQ
4WUP/5tOJ/o66YnA0O7owPYW02/zN6DIXB7x7EsE7Ta8+vKQl/cDumLuaqjX
lHrMRiLj3MpS2ToIw4SgWgt7M+V8r2SLIBkP64bQk8YqxBJHxmQ+J1QVLh6D
wlT/AtcLAJLz4M1qGr6EbKKZM452e+4VRH2ApJuzmDOheMEZcYBK/Oj1pWkD
w6guHQmiO+AT3jcd2q09RNYygc9YrUUgEamc9bo/uj+ctrk17IINmkDXGvxo
u3fB2R6WkjPgmUKRodmXpFxdXr+MESyNsi1OupUdOtJaJwYvQSRjckMIIjZh
O2qRDz1bWOaXcLMFz9JOcnlSyqeTy5T0iJGVCwPu3rs+iwTRo/zLXs1GuHxd
0l4raFvcYQDjnV5fFA6JceuA+I41MiHDOC08qa0D+YTllIhzGrlbDNx724TS
dwQxZ7FVNwTaC3lOCqkORwaMtk780lP7muqjGDrRghA5J6ZV3gUUSqKm+Npn
lrwsOwVQ2JgjvevwYRjGS0ehzrByNRnG2udSI/VeZCD2/Spgpv0V7C7BBri3
7Sa9Uz0aVUloW5qRCMvqkwzuoXlRw948ScWTkjV4a2eSxAwQFqzJ88i9byuY
FqKQ9oALHn8x3FsYWI0ZBMcPAM/3kCtLp6Hov5xJeXkc4qTy2B/y5EF0VAdq
/720yQsaYklQjwp8RtRzFtFJWtgH9+/N9SGneepuAOlekRqdC4fAa/23UKmJ
aSrSamI9WsRG6EKCD+pbZYuSqin5m1bzkSDS8M4l7P+3Fw8hJQ+hixuuAnIs
20r5NR1oVeKmnwGGoLCzzfr46MuHQ+PLs2HMXGPd5zIEy5zD2O3ANWMG5eDa
B9h+5IAwjrVdEpGt3VmO1o0HgmQmWZkC5DXma8T3bYgWLeb8cKSViXYgiZR0
Afby5EGlynkdubwaLdIFps6x51LoX05sm93PVwcxZn9furDJDkqo7BoZC6+d
yCTYyVvbbv+bna969tNE2UE7imnynLZpAM/YODqlaLordoUsN4heAwsWiKT5
wfy/ziu97+wsxouIIdET45WtoxKLUWNDqttvsKSWGunAqbCmuLDBRdEw79Vd
7uJJgLpWcKIO5aDrPedE8L8i6xTv9ssX6/1bQ5/wNRkJZsxoV2eH9D2dtgdn
yppuLkr2LF0V37r4DV95tFt9YCAoQkULI2DN92VRWz/iqk6QdX+iB+dNDcAJ
dCNH/RK8NvtM2XKgqltSfAbJxYNic6NhprkSaMuCH4jkxK3rJMlM4DE1Ee5s
BBpO6zJxv5sXdiuDUkTZSOsVQoLDY85fdAOaazs6R4KTkuAjVc+zyq5p68XX
m+GkxQAeTr8pH4tF3bLpYPZyIDZecCcdJD9PIaW/Cg8uJ1PLx9qyNFzKK4UA
0c+K2iY/m1tY4yJIzVbjquU1moTQL7olNqy8F85eQ0yl7e8CWirIDDPcnlid
kVWxtzCXG5EB/aDhx4M5aot3v8SbZOUeclgdwMG0eGtHqEA1yJPIHIUu4p67
eEk3xLreqogYcjLoor/QxBSLSTvHA+u0/gBGL79vebj2HbinMqdoZ8RLoYn3
5s9kXeCkQCE1Tg3v6CYd//s003IZFdStDG635z6Fx7qEAgk6gv/jHu93Oi8p
lyLkcQfBw6jHdEf9GB+dZ/xkhfeG9UIl3G/CHlmr9kAhSLLqxzg2X1DyGtMi
1ozqIq2cVZLkbnIVU7msL8fiH0sJ2NIP2AXpSOMoyNqwLCxObSGCUikuHso8
cldmqIiKPQw0dbCvFBHopcmnRdgLEeBrysjcpavp7iJ3azhjyCLbX9lwPECL
5MCFyMvL6yCsIAgOSzvAdDtCQLUjHYlYSFyGntQ+QJq+E5LT09kp+xQo+T2N
6338CC+yL6ccZJfI6AbZ1RY7Xbte+0hylhgE7rniHWnbrC+fckoZSSY9ZAER
UkfvxETkvdRQ+iF4+vDCnc4DL7nfwTner0uP8G61KjD2usZuPvKSkt7UNxHt
M5LQIK/n6Ycsd5n79/viHhCva7gOrenEuClcCtF9WqtQW0AqZjLfG72IL8cz
lfSmn6A015xoU1ZV0vPYVEk3vUHEdp5VeaNVH/oOcqkqxwu7Ak/6GmLR73QQ
pPX5eclQZ8Pk2nJU1Md/NtojWTWkMZa9VxQLAJgMo4ZR1xKZlGNFn+RSwAMX
QeOglIS/uYl3IGvdVOH2N6jRMDGsHe2x5OQtfApqCAKkiQ2aTOp+Vl/8lvYS
GC6NyExja6hSl/Qycf3szJSZ3qa+g5gsRllafy5OrEYabxTXQv59VFpSTTys
P7WlzqkPEEU0azC9fNv0wGp5TUbF4quSS6Utp1ts365j/JtoVS8vlCDaNGQz
4NPKHGG95abNyt2m9Q5chjc092R24/j/mzktpXWp+dlzddlPcA2u36voeKP0
vEPUza5YzUgpKwU78mP9LWJNnQE/JXmHuku7L4Fes62s1UfUd5lCynWhxSP/
Kbo6TnBXQvLpxXR94U6rbu3xKuElRbqwFA4EltVbLbFcrc7C/k3keyeDTnqr
Wnm5vyjbDmBw8S2rhwLwkLwWUW5XGvGWbFPnjeDbmtbLrORr3qJKWp4hqSb+
kjvfyEkzA32WUtL+1wqjHNUKXhup42ta3w2bXGiXIHd6NqBrBMMBTzePC0uP
DtQaIcWYHujI7F9y9dpnyl6E41AHzk557qAb/7nYKypiow+5T+AGevhDkULU
ymGF2nKhIj8BZhxTxoA+RjCgQo7nKIYvgKSeOwjOMGKpIsiHx8wwTuYq7SI8
UAekCJzDTtXjg7uw/t8e/sxrd+wjcReMAapRQgjW/q6xGJ7wPcyBEhGrevK0
9B1s3e8TcS9Q5hneeF5/TB4lvaDSANeMF9jJpv+AozjqcaLLMug3yk+ioN/D
GFvNdNpR99rW4An8i819OWdJDd8gPaGuBGZ4imZ7HXkdjPFZFUCH27kl7db1
OhlITqNuOAIAoAcOs5KIoKBFUfYH63oNp/KNHrGk93IbHYXLaXMwuFARDcVF
FWpSyD+GtLL3rW+uO8LB0cb/wMxq4ic9keXgPH5twZWSMfFvFfyoGDwP6Nn5
q2cV099nTSDK8iAdUT9nqhJa6mTNsWYq26sAVZSPh+MPD05cvG3AkSUhpfr0
rpoOfHi/XBV/JPsn1TgjNgEjOYP5EOT4ExRLCynPTQZ439aqDEDvO8QIQfa9
yylBQHI7zzoYAtLGetphP7qYNGZOdV4VQPfhbvNBECOPYpbtKhnmhaPrmaH6
v4sk2V1JoKnsOB0azfNP6fLmPhsQxBVZQqtk5ajkIWODnqpfO1MCMz+XBFdt
kM2kS4p0XtJAmxnvqb7C0HFk8P8qVtqaI7F1CGAiFpOWU2AOhdMwmHQOkl40
f4tMgsn0cYUYqPjSyRrCjGf5R0QRA0SJyw0oumerZ9rV6hrdLGqhkfHcwKs6
kkegPnxyi8nFCO1NCpOtXot8yUAVU/zT5/7gomG1w39nNh0A51J+ca3nMsQ1
PQFqUb79K3mjz0gtkYe/960TjrNZs3AxVpkrAX7OUxyExxPY3iTmAfsHIK0f
KgTH8CXyJBNNMsaomB/mh2R5sjqRcJDkneWMfxgXjY20l9DAbjiSfyP9Nztw
1HJTajjfxuO4GxhugPU7x3qepdAMKUdZq1nkg73uRA1wEoOZOcSnKbcqyTX3
QxFbgpgCKtF1roi+jfehi6m1AbTatC9TZq3IcMt8+xKsyl1ceI23vEP/gd4V
ttsNsdRqhaYZbk+hbYHXLYdCeUxu+JjgsUW1o/BFzg5Y4B/5rqfG5A/kKAYs
0HpDNcxzvOKjhTHLuCPiWc1ek9uD5a2gHTxAdAw/IKh7uDUw9aOb/O8NfGTJ
1ViB1kJeALgWvE3MpYXo81bH+v1OLPLZhLyGMVGdzvdvqMJm7/5B87TcVkXH
n3XsaaU1OlzTWfHZ/c07xQv/NsWhz8KoudtpIBy3nIDzXnIC7/AdiRczPX6M
GR/mbQTToJm118r+Lpxk76dVcvEeIWWeTLaR5T3UvUocK0Hby+i15ESrT7zF
g9GOWErfuGZJVX5lrzAsAufj9osAzkCERKaF11rEQihwjDzuax9mH/O5oyNL
reqwFlIjb9ekw6lE46DtxTG+QmRDF7/wrCvXj0A7vAPk0/YwJOdU7DbwJTFE
XdfgqqirOwfCXtCVTbnYjGsEOiTor8Ppzn9ojxDKYNefYXbCZPNnBSqwMopi
VnQvDc3FDqM4NuNo25p8Gu3zk/nCqjax83YW0e6GJw7XwX3SJxTO1U6VULJ3
LptSXNy0od3q2KZBffukEhilzWdtopSW8EqLs6cw8ZGIyOOSEUjnvyOwdAuY
EapEf2hA2PZvkQ11XRoZwo+LlT5bs3Coj4EN4Ursk1xg0lNV//FalskW4LKY
Q1jlzOnVn8evAuqbT0J13pHDmdXBhx7uT/IDuV//ciOJFlkM0WIJhYh13VA+
XJH1oxfDHvzbnEylR/2hAlXL9C8hF8gyqx6k6DQvRxyRIObTvQQPKan31QCS
t+o1/PIaZVV5/QihvjGAl94aF2xahZYBIYmll/94TFgp+9Lh64usW5y8n/Dd
UaZeKokEoayRGLjFqxFM6qFFtcuqTglTGL3uWBiWaE1Uf0/mjZ9kQ56hsR7J
LB7PXvBm7vLLDYgrnEJ/dfw4jpINql20HI9MGNTF6QsNz5qDLX8zMrzZf2e2
2y7F0mL3aCam2fhRlu3QtY95RxtgJtGgXvKyZQsTRuDm7Cji54SqUN7wXlaD
wlcDHCByPiGkYaSJiVo0AN75vv1w/fbYP9xtNfkRhfLaa5ZSJ9ryucYPvmVa
7L0f303GSWuTzedNh/e9LybMrIw0DE5wTjxBXXOuspTTpnr9851hHAsb5HPy
ZulyQQJd+uRux6JpVYwmC7iD5IUR7FWTZkYFQ3f5AyDepDP2CyVYO2HZTPqc
ZeKetQHssfKY6RTtD8WuXbbWV0JAH8kBp2V8yRF7KLheJ0Ve3sxEmCM8jsph
Ggta3lAI++1RLKMk2Xy2eSvWYaLD+LAeCx9u+s3fGJrFcF/Pr+PQ3s6i/1iH
xhySDIDarIPeA06sw/Swuxdk/2C52H2QaEPnZ3nlCvZk7RvbRWWOnkL0jUb+
J70mkjSSmCe2eGVnlGCi8VsJYfI/y6iR6ZsEYjf7MbdqxzpUWNb+E/FzLxTH
uITX9ZCKF4yifeuotqGvUHWXZLZDe6n54PJBIna43atEE4LpickgvKwO2mi5
JtpwXaWu+g1BA/P4KAbAmiMPHFS1BuxbnW7WphQPTTUieGfhvwGoj7YCH8aN
3Lm97KUhcwF1Ng80jdjlEYHw5a2ln/Ka6EiH8dGQMAhhzyjwnFf0xTabPOGo
odz7hKWuQu1DXnMPWXiT4U2Z//+su15++lA8P/VFX3fGgJJycD7qO2Mxli26
ZCtBEaTK6h5P7KvWjknbkHcnkRETpbrXlC+uqYtF+jK0FquhaO3QyYepHaGA
RGo5CUpL/+/4sdLA7OfIG3ynG1uyAvwk+ml08tKusdfu8tjNYQ4LaJO0FK/8
IEAW6IW69zn8eiF17rpBbs+ByTMNWwCsXUYqjGg9qxgouI471KCpDziMWwTb
W+K2X1H/tLlsZTrCMzv5v10Zz4kJO7KWg6CvfTbjEx++abuoRR8t5oDaYXRZ
m1jT7hcvKKiyvcnOA1geI0Cj4hsynlC9W22PfOQQA2Es6/hMwy55BqOXhnwM
D6xp52zlO4mzdSuZJAn7Nw0FexjMD8Xu2XIal7Ogkr0MSJLJI8EJdBdk

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EqicD0WhRX6oizU7fsibWkFroQRgQDLybUG/pAg8eRmF6skaclUHKRFS5KukkK6jA44Eo9hAG8YF3dSFOFIaLUpn+9btxcIAuF5kvgqikT1RZv0GUzWXVyTqy2i6lv8tjvJieX8gfGCAEikEZM//WfBqoeGEMLIMxgPWAXVVx6pEHfDv16UNSzPUr4R0Ll1dNfA2QYSvLG0V+3JVEsTnzwIGOxKxBFYXVMziFM1SyW3jWIQ0akoDXHHmW/JuIC5ujnm+hRyo9yvdoUsDty5hmUZZ+TbHnGc4UQiQC997JrPKsvCXcQEKagKZ9Rd2WfeXJ5aROiIkJvfqZy1zX4OAhl8I/ah9tDQjekXr0t4TcWLMrA/FlDNIX+9zOMLp2lFtj8WprravNYQow3VW4IOB1UBaDQmp6Jkx3BKscLdHbnAUYonT7vLQE0B0v6XeRFOtsnyQhU7OMooJuvt0HumEyEjR4M+2MdCbRVuuRZCNOKgOsZotcnbUrzTEEY8uPLkdnHY8zx6paq614PX+vGKfxKRwYM0Z23SipVPeW4NCMU5brGTj6cRt0MocLZmzFcrb99ig3CA3+3nNO5gkjY88H0us1y5SWnI11mWYxjAmjLfmNzyqkLX2Gr1NeYMnWraUpm0nhsxUQd+mPkXcAzwsVBhr7VyVEQasPMow7KL7C636ia7KZUbtYlyIhEQK4uyqtBeIfO3IV2Dx+8Eu/xCUyuN9iYP5yoIEMslz9ixKuXBaVxtbMrJISFK74j+ISxvGovzPsfDth/C8se54CH6dLNH"
`endif