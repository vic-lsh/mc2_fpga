// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sWa+M5/q+vZtdqLSEOYqFy/7eYz4ZPQxHk2xNu+GTDAYt1W9gpPfdZTfPlvJ
JXBhs+/5XO0DXKsZw/E62USvXQ9aOxEmtXJxAc7iqGCpqAIOhN3AddaAdzb0
5XiyLma/OUPx4BAs35Yv2FLRuxoqJtSWxCeZu2BKK+8w7FzQo1as0OdRK6a+
vIQkJPkkm4VKX+k8KZ2f4maHwpc1gaGwDsPQsGBBcpSoF/jT8vImjXRnsDmD
o2pUjpcMFl+fnY3PJFZlS2jEocirlYwfEmlwOqZ+xf1Z4hUzRxhpoCPuhqVM
lH2slQERjm8D4tTbk2dbFjVpQ7hy2Icbi4eVt1vIiA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EN0gUypCOSzs6feMmOCqTLcRx+yZAJLah0Owh552FDVeOXwXPoh85Ud8Hb9N
wnmD1vYGW2hmLDYsIIjaONAWyahM9LZyQO1Pb/QfxTaFN2JV9+AwbrSjwa7J
KVLLyQuEt5xH8BS2fMhZ19KgJzeJ02hfu7GALzxR/DIiXGJ0WVyUD9URD3Ls
dRNWpaxvNwwf0Ie6kZ2JjTLu/T0P3o61NSWq9NQbySi338xzNkfOyhKGwrR2
xkMAmcGPtFv6BX4UOUdgFL7/Yuf0zZoX2eD6lF+llQBIZnJfFCGG0U5VVitD
uODt0kjH4JuNs3kHP4C0J7f0gQY+5xKnK/Xe6AhLYg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HeUqyZ3EJWZXVso2cvBh12QOpFucnEUfZ7VDaUsKuZmEjR9hxGB5fXSoizg0
yZsT3XWLLmxtalUC4U8uEXV5ePf45NvUYn0hw5RVbvZrGIalYUWndDmne8R6
fs1UqZMJgYbbbexVIEI1TtVL5AjRejMetD9MPWFxRYMxD0jzecK+lMIfpLgh
P9tN/sTja8xrbPSQx9YV2wfkO/n+uFQRW+nYUt9i15NXTxuDYW24vb4a45eD
ie/4d04NgKVoE0yD6AK/bCOcQ7m4zs8Nfz96lZZc04V4xV9t/BPGnVfrSeGv
g43zZaD+wO+36/BFmGOVaFl3ZY5ON6/qySHwTl7gCg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HvK08zx9ex2+jVEnOTT6aBwFym3yFaiFDfDMZhSjXVc1hmz+VuIfC1hN+H/T
BOyqfslOmHOVDE6dP5gSvmEIu8c2DKVRd8/iC2IXUzrHSMDRGnVovh+m6CVp
gVm67MOgNCoJ56hycwzkAolTqpSkojyZhe99Pk6JZoLZQdz607C20kH0c2vU
o5+Qo3tWhrVARcAV/sWiC6Y0kibC1KSfkWBNDpRfHxWTOrejhve3c8HSQISK
7G9MR8ndQzqlDc/B5YzYLB1oxfSfnPSAc1mE221OFADEt5W76gW4DzUEOpKT
VYb0xmuRekAUHoJW5cJjiG3jnHAnvlDgjlfCB6leKg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FzOf4N84u9Z/Ap8Q0fXy3EQJ55U4v+r+sasFbfp7ytrLVhkc5Mfy/CFtKmyF
ooCy3etsaXdnNr3Kh2CruExzFZepSeYyytn8skvf2CAyb0u8xmjB6JbwdeMm
/NY/xfzZLjg2Zd5Sr/VeDLNPLRi3tY42pYPpkLEmuQDNwi8AFG0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
swu/2T8JmvWL0ydEtnTqArWFsTS4cmtpm2Iu8TW6z6AMeOrL56chzLQpCo2B
xoS9zXxgSf76dDr5J56yvFouN95CMae++Vi4/E4v17AZ5ydliZUU7btQp5AR
n7h+IYvb4l6Xtr8AD1872g7Q7Qd+UY1N47S6O/vrGiGys4nv0MOaZ/2p/Duk
EUg8m456/O8JS+uOdHsEQ9wrxx28mr2VTDZCQI7L+nyjq8Z7c7aon77pRwYw
fUP7QdzZpGKPddy/paHSlwy1nMotNuxkJDQTtAkqgZYN53jFJ+DJhopDqD8o
OQFy59+ZEXoj1KbZn9HvQ5qNuAg+NBc3hUZnxgH86vvOWKdrBy3C/2r0Rvmy
fmxVf/Ba/l90F1M5E+HkOT+JtFV8a277cGydwtPiZi085dXB+N4bgdvLUEB3
ioegv5qfZXuaC2ZoEGdndR+FHWpt55glMQyxDj8yyU1BZd68laLahZHBIiP8
A7Mp8ns2UTZKdqxY8rzZczb6vXF7AjXw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hsqHaSquoJnMd85DGGo/AncA/xZaH3ryefyT5syKX4sMHjNse+MA+vJIpVgm
V7VOpA8xlIoNn1qpfD+7xi20ldaBSDJ0I9MsLkE+D6D3i8HaMHbYF1xEJZWD
vfpiSKrPvDqoS2ZTAD8G3MIp6rLfRgzGU0O3UKPfP7hhEvdIYY0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
stWGUQA7fw0tjElbUGbNgsr+51cNKJzfoomCjKBSAWbin+lj83xE715UL0vE
QQF1bbr5cCOWnCOs9DEwqOgb5ZyxCUaWR5EoPH/MfzkE0ec+MuJ6rNDTN2D0
b83TPLmR0s3EYd05XKNp3J2i2sk2lLAc5zKk4AWg9zIGnBhrAzA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 417232)
`pragma protect data_block
4qOfEmlocYuA9WN9Ps8nU6bKYp32V3SdmR0B0xr/WAo3IU+Vof/9bhqnVcXq
HfND/DTjmAym9za6WLQQGoDAkIr/wYYBd893HtDVRqXfuFVbpuOaaW97GhJl
xTd+WjybE5ezaZSeYXyeqkcY/if9WCAb9/C6UXSREfHldgRr+rPdP5jEsv+a
gg4HrSLPbMsv8uMiGGU8aAWtjp3yf7cYJ2U7bq3WTf9kEJ2rLDOP3rF7s7Oo
S7JFUffJ0Ga5pSveKy5Uyc0ywnwQkINdTLX5/iijJqlLYiowSO47GhjZydBS
9Cb2/vnLMVmu0xpFm4PSvuMgOYbpGc5RgeS1y93E6N8VWdMavDoEPfPSKcpW
UpL2x2XOGc3C6f/RjhBWRrP6Ziv0jiQaPIWhE+yD/XmT2n23ojnpgSjl6f9X
7KKkHo6RMcuzZ4NQApL7WavrYg2l3bvZ52KrBJmIaqIhub+uE8gs6kaypGqN
v06ZLJakjajFhOYTkWBBiMTpCOF1e44GVV+4UPOFhoJDcN5EKGVN4fOUWtta
kFlyS6tRJkqNClOfZg7VMFY0+kdoCw7SoXFaq1n1yNz8ntRYWl5PhN2m3SFF
zwiXJ2QSyE0DJdMElq2Fhqw1+/qNxcm3RK0Lf8ck4VR5QilZP7puPtiSIjrK
iFWV+20VRsdvhgtxpzkE7ZoZizp7RfP1AyMspFvWg47rOdnY1X0akuZT8QT6
zPppDztFfVbK0M1zEOtkf1cQVkFZlyZdzfRhbf4tu/Gaj77fhCXTFOKHypBx
4vNEdAU0I0MsD0bRTrP7s0XBmvefmrde3rXFme7lkrKY8S6SinByYn+Hy5Xx
iGor0SAiH2VhvORDWL6LbaWddo4dhUydExSAuqr5JWuwjL95V8/CphCtXVTE
sIUsNuw8Y6Wu6EvUkjyxvV5ZnKzIcnd8AiVvuz4IrKmyq+gCXKE0OTIeJm9H
Y5Ng3bM9nNPgn0rMoMeD8gKyNVoLkqek8/AmdgKFlDD/e4106VT1l9dgWv5S
X8yFtpM9laDD8ngR510RDZD4odHiXEycEI87xWmU5lW+l3BXcGHJo6ThHTwM
ltgu6DRTbBuw3xyzwaIXPmRgOwV0bcG7JqXFMEF/GDTQgm/1kE6qfWj0m1Kz
O3sTyYTNLjRo3z533gl3frR+H6sH2gxjSz901qFo4iYKgw7lS8HS/AE/22Iu
u9Wkc4YCXitC+XLpzxDdyR4W3cIa1Gjrhfr0SQcl1x0IerlpKVfIJ9UvbGTM
5PB5bRna6ONxmEGqFTN2TkpTkFAkblagCyJdZN4XIT0fbmc4Uy70g4VqlAxE
9sEscRm/TANF2ookkXDwRZcYIEAbOiZfVxVQArxTQsRHZKID1c34Cebk59fI
kXab5Dt6w25Z1vln7AKJ+Y1hgWzqCLdjZ9UQ279fs3gyGMKqFPxGNQrhXKnn
+3R92Eu/GnPgM/lMDVJp0c0U4RpfwJtTdhpiAxKKU2Y2BNq7Rguz+/Oag6+a
9+0LQ8w6HqD1oDoEa5sVoUtoKfoeUwAQNJXIRs61i54sLWSDMQKtErK1i3/y
cIczPLyQ474wOGYpfJquNAOZLIg0yB95dQdy8F1xOSEsox6Lw/9RIE6DxA2Y
Isq6zzj9ujzd/sivSoZKwaAw8p7nKtDQjuY08dYTP3lj5edFdjUtWFRpP5tV
cqSOMkIb6peih5vb/RICY70AH8CbtOfs/V2XMAUTmMo6gAB7PokedeEVPRdF
m8MR4zIYH4k06DP7hp/wliHS8+wJpoHIkbKRB3swU0A1amSDU2RWpXedcQz1
EWUZRInoyFSrHHqA+V9CHXXIqmkI0kyKjYa0gYg/phHSSgRS6lqmGnYNXlVF
vDrOSeGxkuatODJGDIYC7sPLmMxW0cuqgOLoJ6v8Q5SlMANj+hGQu56x2ISe
erDAiV1P3ayVxY+sbyROwHo/MTtN/ceRfnodRX2mMqxM4iMQ/2shVfzdlJIo
PiflIKYab2bSgRgc+YZm/cMcvY5SN2LLo+Uh0aZavb385SjkDAcGFF8z8bbb
OHtu2YYwCwC91PpPauKyh9Qhp7VDmIUzS4rnrb915nJbK5X7oCVtG3WZcmSp
p0GyRhvZPlJ8Uv4r5+pR0O8HWrE/WmNFxQEbqP1ZPs9oc4FL/IGA5Pf8BXe5
MXfYJy3ben1ZM5HNhVmB/EyMOW3wQfHiLQNQsa+Fg+p8m4nwVkwJ0LXLd5R9
4CDLn5692EmpiMK9y5fbMi4JK78CsnpaHXVcifZZGEVUUyRK/nfIjFurpblG
Xd2p19W3Up48E0qoM6pKJymVFDM/IjJAA1fL/yXFkb3T+xF3TiCgSVEQ4HQL
dkiO3e+cnSeRVbo3zHfmVftm45LrYxSmNBzIxXkGNrgsuKLvumYPbQ8nr2Xg
UGfEuUrWXG5a9NIbAMYByKKB8co9rHSMm1dW+DGKPd4BWiBmXUHLHSDU67tn
yQ1NVUjseCda3uhHEMMZerm3sgAKD5XtqR/BzW4XimSXgXUlr2P3K2zWr6pd
12ASWJXShDfrSDIymfc5KnGrTj7kNBu+uoD0SAnm8DEo3Fd2ACjGrQYj3Vzm
NnCwMKxnHCU5+9uBk6xAio5jCR9ZZg5tnXLT+o4KhedvxGX6hu5OEsVnIIPw
qLUL9mkFVD8IHYdXKBT2Rfh8zmoEZRRzGfIWv5BQbiOMsGaAXYbrcrTItctB
FFOE+rmWX9fFwt2vPy9snukEcEOcqdcigdRR4qakl50WW2KgUJpSQxDhB60T
8kjwWE6OcBvPqcoa++w6iAwztD+VZrAOogou7sPNEzqU5Od6ZxTf+Cb4ucPN
SPNFnxwb2EgNVivzbTEA85KZzNIQ1aQtO7IW2UPQbFAEtd9L6tkJLjoS4mGI
YgPMpW1VSEjpBk0iQtGEESFxGGp7t3Y7+JmlZyKos7ljCvbQTXCMf+KOARPW
Dw9UquG3D6r/mf1bf/C2jFxcpFFZafPE7GLldZw2Ez1uX65dL7i4GKcn3ewV
8i5glrzlFou96UxwsWZUHp4hT5TRi336X3iVYettidfnodCE8e/qjgGMh9f3
3bDpbt2CNhFf+yVipX3KirBZhHYfPtK40i0PZeE7yI3WlkL5gqPVzWU01klb
0iDTE/iHZtbUngs5b6wgR/mDJ65nhNJDofFh9nBwDDHkelp5fFt83beVXKtp
srzF273nERAjTRYuuFFq+RMTEcJulUGrQqJfBhaiW6ogoSdWobiiZeh6hxap
h47RJQMPwOCxNFRXJnrQI8F0IsCGMAZy8cLw/yNCCN7aQeJuEA4U5+F0gY4G
MoOD9W/2SHW7KXA267DxDYe1EUOkd9OlotOrFW6C76GjgDEWsUHwA00ghbjn
gyrkKRoR3CabASaDikEjwKrWy38/0lKCZ0Ss3DvOu4iIsgDRgfAEz8s+XYSB
o8qr5ACeSiZ0iIIZzmvmNVuRGG2ecsFocfaJliBU5vlOfYD4aYOl7ZXJVDZz
4ExuVn5dc+P2rCZoW43NgDl+DCbPddqpD9yaRJmFGEb0lhvggFQaqRYBQKYn
Wa/49/1GsK6oqP5q3FPDOa74uh9n/+Fp/VYlO4PWcdeEOjIrHm/NYDAc4QJX
sUbhrYtz6Bvyv5EtiwVdZb2jXTtscTcw5xW6MeqNye4beXlBv2X0kvb/V4Hr
wXuakOZprw1L+nTpvcmlpb0gH42XZxwUg2Pb4Tx+iTZZ524o5t50AljdgP7n
aKL1bLDs87q+W1e25NzxNknD85TtEwpfp+YbQZJ//esfiyzpjfSSV2Tcxci4
ab2q3DJ7jhhm4vWnM4BpvvdScvtMNdVFriPec3UX+OhSk9PlsIY9OXkF1sGN
IJB8bevEVWSLCBx+OZKPhMD7sK42vUNeW0UdMKQg3wjV+BETZDRKcz5fepRY
l5Ouht/mH2S/EA9beTYq7R1IG0m47TS4gQah0owxemSnxC6aJkVev8E4KgSO
gz5TM3XbM9AZpg15Owrf0xV4HN+pbdDk1NsTwUyBWOueJyfTTOVcv6WrkWKD
SjLW27VNypAJF6AgUKIx0hkNBRuGexVnyp0Cy37hbWthiUNoSVBoR9LJ+FwQ
DWotC/Ij0f7pdek9z1FSeA+YLbWFSKhThk9624jNWR9cmTaILOa43O2uhshg
XZbo6XpeEMIBYN8mcE4ErspPk2xSHiwbaEPrsMf5V8IYMilMp8DPWkZz6i3K
VbNPcEbXSfDYXQYI8i2a7Fmn+lzAyHv+0/SZFHeYBz8hEk/um/8D8yX2lY6s
A+NVHKdOcRGAMFu4AtWo0SYWMMxfyQC/N63xfDlk/tuuOQMEr6s483bQYSdx
CvRZsVFVqHudPxnKDBHX47xSz8HHuI2OfYTghsfEXGK+jYr8x07JHQeWm6ho
D9Dm0hGuNEn0jZTFQLbBb+Ny7nUbziqzy72ijkW5BuUdvlJdaQ/A2NbRTdvt
6AWuwv3MfWqO7QmExEGKKJ69OOmvpOI2mAuEyhrE6j104dPNnojS14f1bkl1
q6P/Al16Ir3IiGDSAXdL1+LtgMW3G5qaLWV+1oPzpyIJQ8V7XsNehqtx7Hg2
jN6U9LGcAhpk5rx7oMGWio2sS/6dCf4AHaau0ccs3IcAn+1l1pqFGKaFHoM0
d47j08G1f09Mq+c/LIReOJvol/5/mRHUF37MU/5euRbjN2C16kv+ecnDpms4
osSG2TAzBg95DfebF7If3iM2HD0W26v8aqG0BhjMlOioXkhirqcGajvsZ98c
x1ULw2VkBk5P9AmzztD9o040l9xRnBdZ0qA/dkbenTpu/KXt3G3MvdJ8YjcC
wroL6hmGBPcFueXsIO7zByYR/bawV5cLLSOOIsspmguoNGDZxJtrOqH3i2KT
49qyog5T1QBVGCsvfL+GyPtHp1cWu3JDNpNqnZnKcqhKBl+2whMoUiVJvhZ6
CVd3ktXSyAdII9Zy/KRJFND54rEQ4OWSKK0BOpv4MGEPqNQ5+TJXV0MNtaL3
pk8xLofmFeuKzRvRR1pifXA9beNAHFokY29ehBR6Sj7NGJZSwjf5wgiPIT9F
9AIUZjBv2Y5F4l1oivefkyz6kUkX5u2AnHOgrOYzyf6u4KvmfAR68j+XwSry
2TEAT3Fe4wdY3K0ZFPCNvEytSVlOWutbXBT440xtuIXt2jEV7Xg6+8hia72d
mffp3sAfhjTboKNmKPE3x9RLxKEllkrxZbDVg43SSVcrgqjdPm2XFfJ8C+Tq
3k+9aOMhf4AHxx9mwDdQ6m0kIzCPaDXeRUjXz2VkvU5sebYYEnaUCIDD/wiX
ZrrAGZvswocRoFP31Kmsi6MU/ilH25MyPdG+CiJEsfnMc6zTkqHvhL2jdob5
VxLrxrtEkb3qZG7pJMC27nV7UXobEs7XakwEAK75ke2XH5vjynaAwN5gyU+F
VDvmHSlN3u36p15GbhA41zqCNz5GwxBF6OksQKS61cwxXaKnogRYE5juwwRa
+zMUwMlJOryDYq692MC5JqODKT0O5DpDUUmRgPDinptxOksNKhsaEZHQyWna
mv7lGB+actU+hob+EXBzMAVsNElflhx9Q2fHHotDO0sLHOj1GktC+EK8/akL
jOqbPhM4XDeLTmDFuJOHZ/xWUiHnmBOCbNpDj5m5e0esVpIY+Mgqhj2Tgfk8
l3FgQQIXjolwWLfII40cjRP2Mhxkvs8buSDJZSXZf5RopmbkfIMEUWqha/lX
VsRisu4Efk+dLYY++rOCiAKcfUTzr9vR5VjXNflVEkb47q2zBJK2rIGeeUxr
Q9kTQo98IqSnrw6nhYj/mEaW7bx2gyPFTbahFEHHhaYE5IMa7bPsasUp7XW6
5eC1xsOv5SyKlYTIwwKbqNkOi1Q9KcqKzuv52iPQUI840n0RDLIc/SKHfC/t
cDW0+uIsR+FpOz4LzNDY4BtrEnGa3nnenHduUyvx4gh8TDnfXt5zQaqoX2Av
Q88bWAwNs3XSHDjAsbV91keRdRJrt8xuqdzbZ2h+VmdzqxkmqE/fyoJ8YUtP
tEv2eIsILnhnejol6Y1iR9S1wcuWQICVJvPvQM65QFaCpWZPH7nPc/5/lAeK
yzlUn60f1WWu5zE2W/YbUIeGFgtPlTR0zP7qAET46QGkynwZv8Sc5lm150z7
meIssAkRGdhnSo+EGsRiaQ853j1lyFW91/nMeMjkvt9mwv4UAsuGIhctbxm3
IfhkizYU5C7qmBytB00K0krqhdCajy6OwHmYKO9IxPs9siTC+xvlJ96+KYKu
tdCWSv/GL1dGSkAHgTOnwdaZf5d3fqWFh2J2AdN9ZMqtq48n93XVGdM8a8jB
c2ByUjjsUy3UQpxvWPbXtceywgnuQJfW7JpR79bJEyBGIh7P0TzH2YF9S5dy
wzIaAwnV2X1PGYHB9USYgKLoKU3n6c9f50NKxxdwaFrQ9jPNA/xhKWQNiVNn
eAk1X18p12xl5OHitrdnGX521C2n91tROMzFt7wFospJx/zd+7YZeYY9qJN8
YEJXjYl21EiSg2W/IBSWLDVRzAyR1TfSjg2a5r6fI7Y3PHwgwn6D068lXE8u
O+tDPAl8SMcoNAEmDeJYwTc+oJY14ddX/zLQjO+8ZbSXwPHTS+QkMiWsUEUp
UImqKLzYljS24VPHHpahonMP6eNGg90n3APokB2VDaXGjju65pymdcTJD3+n
ZnCT8xHqsgKMqyUku89Ycd7FefLuLMaqG5FPpkrPd3uGF4vJRSf6X9GJStQ7
cL8tImYQfQ9/VkaZ9FiNRv6jqYjyXA/bjylBevd0Jkg48SqhwlR1WdvbhQfx
LXD6G/dX3CMSeMLi6WWMn14AQ+VeSHSiyp7UUI/RsEl8pIOqi0vniWEKBKz8
8vTfPbJPCt5JIqKAwCGSRNGdhXxe/vV1bnU/DQQlpSly7MvFAGsl5mqnXISy
gLwAscrl1KIPbAY+a/q0Snh00c0e6sdlyGgpuZI9oWHYxRQ4WKOf7Ukt4Hte
ZBdZyKIvKpHqkNI3YKHVu6LTXaKfOTNMxBzR2jc9Pt/4Np8k5xlCOxNg2Y4x
L98xod2nYp3GFx+j3dtPOMWDDlwZ/DV7iytlzntwPtCEyevdRkSJVFvJgxXJ
E5izkGUEnSCCs/vc7ovkwkIFwD1OF5Mxo0huPfg946WGcs68ollDouZ5ECfk
Po7Ou78jrUlbStuxAebgp1sesTJ0dqlWgheUtxlMEzLqHYShV4OShsngxn87
JvSwnPixRQphzhDBbaZKFTkXHwLZ4vNLkXrELUqmVyaxCVf6HYfSHUVBOjkL
+AR6OphULcP2tz6qy9l2HMRk1KUhSJnfiMZ3mWoJm55264khNayXDwfTA5gg
1jrKlSD5Py/GkE+uD8jMlGCQ3981/nzr1BiuhC55FYhKBYnSOTnikF260upf
ffn7T+vjEAWBUAK82AU7ePnl/M+/p30leOfLfBr5jtg4HnQ1N+Z699FIjSv/
yrwgck1ipU5ofjEALf4w0/tdmEi1gSA3uHu6lH1qeHDkxPiE3mLJX71GfrAz
JPtCchSQyPGfszQI8e1YGQf1ygjpdjJKmjptZz+ncJDAKisJf8W1d3UqHKZk
BHfUl82DW2Z54dRYVgRltPgMS1B+HzY/lPNBysqkClX1JwxGGF7YPWyVVqdX
w1oN9RL+4VhNEiaMzIleVmZkL2hjkhEvwjL8v8fJlOM9tRRxPwAkwJrzXnU1
6Rgcb9wB+OHDz0XIKNEWMPdRfGPdPGtES99esMzC0g/PywoQbLw5z1nn3/5m
/pxvnc6Xhe0FelHA9EHF2ERngsPWm4HjfTorbDHs2Ufyl6Z5sJvomRoZGlam
5R6PPVIPtKR7Ea3o88cnkRr8aXPLhU3oQGS63Kq8CiVEGQN/iagveXOSvKil
yuog9aLJ3izplhZCFA1sRX8KLTi6w1fSDvcA34sR59GP61L8XzP8WBR7nn9p
1lyBW2DIGFCJY8x8sovSzP+pM2Y2QwwcEu/sUT97kabz8aCCpvtGXAF+KRRg
F9eLiO+3wI/6QqUQ1qOHsOGwA04bPxyTkNHWsi0ReNyhv6IHZpOezZYykoQT
vhnadtZgKml9HM3yZiVmfXIFO+HLcICfrnbkpAprFL/1VKKFAYW58kBeg7Kf
Ol7ha3LqGjlRAGt9TTxGTLysgHXTAwJkIyHZoyyJBR8wxSV017LW3dR0ponn
30E/Uk3tVVJObQqn/q3UxzukTlfmTwkQRG0qAKwGXGiwPgmqpVkgF5wcSIrL
zICoCN0mPltHTCPoUi5hzRPOg2MCBvlRwU/MeqfzirrBuIZsZq6PBAGl8+5w
yt3w9+nRKkudOZSrFvVsGwJaa1oxmRRm+JzoLISAHLkP9zOUPjKebIY5E5d0
VrAAEOvwt/l3vVlh5HZhAjteu3pvhvbvyRAKf+PNHxW1W22ZsJ6SQdc6y/OL
Xzgb49AWg4RXvn++cJroJKnx7zuSBNJWQTl4JRPwYfUhVyIT/6wJ+8asI/Pi
o1FOdypTWdLr6Fm6twj1DzDXie/l1Z3p0QF8FFoujTd2DFpA39Vt56zFUDNu
QjpYT7EPyA0RfIYwb6drKg27fX4bDvR8HCdvAl+pADXyWLODJ623MgDcGPN3
Jo8KBGagF1I+j7i5eF5vFnold14ZFdaLVsrLcKYVQQibHMFMk9ptdlfFUlQW
4Jp8Ch0+5AB3pL21grZ9zF81INrEkcv8c7/BSgJX28u2y6lLxnNRhPr1NfNJ
s7T+ybWvatZnjv5oUd75e3h9W2Py6GMd67ZfIxdGGkblHHzxt3T7pN3nwDub
RKlSMiVmSis32kL60rNB+wgGv0tAPavyWqD00JW61c2MRgV+e/k1mkuJd8fw
WoDbg83RZ/PzL4KyNuLSpuucGjFxe4wqmIhOwc0GwuTGO4eo/BE66XEusxA4
oqbcjInE/vIxGccB5KqgcYiaNVWAR+mb35WbHYQ0A09zBzvA/IldctRZVpqo
MwwbYvZtYzqNTTAIDbbtQUoRXSzJem+LNSoMq3aVBl3sAaNmAWOD5+NqHkK8
Hq4WiGEzkpwbIGhXOJECYKCYnpJf6IjGS8auSiUrspafy8KrjwK3fIlmAJPd
fVcY+NoltX+VLKqaDFnQ2wlebrvdzrNXaNW+vz68XATI5v8AeJ56QAFO5qcq
AstIeNJ1eY9WNc28CRYnDYsVplQpCTM/+XaKj7F4Vs8qmk+f3c117kcdlHbp
XIy7swMPH2dnClE9wQLmQTTcB2r00tKcUxp2kotMhhcpbQz0TmdAQrNhOmSm
Bv2CNi9Jue+zJ0I6/041GmdTMBUYs4EvAFke9Mr4m1AnajLkmAgOHa1Tbm8f
LksoheQoKEIVGqdAISMCGxocMQlvadTjm/5ofX9BIVjDfrx7S9hEK12ZGM6g
IUGnoqXyVx87B2tLybwCZzIv0mp95aKwqd8aqZ1ERnHAYAstKfVjmvmiBpAg
q5kF47mVY7eN4qyY7R3nTyM+F/3p3CnAji4OuJdBKiAVFb0x0N4SNbj0SInp
MyhlxCoYOesdt8bb8WYd6rmYXDsxxeR6ZWjyldi6o+7Ch1mq6yLZuZs0WgZl
wUReCG/L1PyevjC3exsaZPmTtH9ubVuHvawHLoxCm/9XUJYzwkqFMSx+HxBe
WLqUtiSGGLcq5WXGwSweggUQf90GIbBIVEQA9JRx8jodQNZa6HQPGAYq34en
nc5X6EQ9a0xS18n5+xx9QOUplQ3Ze7juVb+GkbZMEhsvcVhbRZGXwYtcI3qo
Dx1qH0P+2sGurjQgq2fva2uoXUciEL9nQhsvGBu2WyRYgMAzVr4JdAE3wwmT
GHfRvEDglrFm9NBCj81YAVJD0jcr45Md6M46FlmqeB3r+JfnuwCeEMOHFRTc
/VL5eD+BXf1RCbwRE3ftbWLLnWNHPbKDHUwJgmUlSlwfd8sniCFoW4l398+1
ZhQd+CoeqVasG3MmWOlA2BZDrOscN/QHKB55+zQRHd1DEVLuM3LI8/gWv+e5
a8f47uAf24TFd0mvih35WxM7CruR0B4qi05ydcM9KGew9uc/CQ+AVtMNxJfa
OwRmq89llESl8Od7e77bH0zwvTAsY4gp3VhHzmHB0CmsbPJklRTR20a8pWjl
okvETU1v8zt2N2EocMX2D8DZUi6VTPwWuaESNwBHGxNFNstUnlhkx0/p6Arf
hUl+mayhFK9txzYYMHQjGTshYFyUGRzhSXRaf6aetPhs5drYsXiZXhb8e8gB
y6ffs3oJd2Sltzc9pwiuiYldvhOS+vhAvhJM15FYi8fDcjYvGYyhQ8+tH6ix
iuJcnKKrfoHvIfVjbECqoOa1Y2gH9Hjh/F/JsajelXRNC84J4vTKH7KUzR+D
wW5AqrAdegHzv+Z17s+MjGoBG8KED0YWFgPU7gi/nRcHfZacXoQ/oaS6F8GL
2ktamn/oUKIvNBHhD3XtxEWwxnW85uxjZ+eC50nLsRxNzSJX6XJ7YdJ7y8HE
7kU8dVaVtgTOZd7ESbIWGM6xOh1fghJjRJQD8rdCluoo20x9s9emsmIQFZtG
crz8KAhHZUAl54bUmUa3ObUFM85ZJTYqWhdmnlRYMe+kHSJZAEE7R97G/nW8
AOiL/xJ04oatnioQ12FeTM50Yq3kI9YQCuFncvLaitabpTQcPEVGC/G9NHHT
rk0f8iOCONOD7VXs7lrKQRRYRuqwtHyasKOx/kfvA+xa/26oRD9Duby9pFlX
R50vRngMm5ZIHFP8a3lXBsR89CAmLLPx7w4RrnM+TnxwlAdmtxa0XVL8ZE9h
rcyWVfwxTz0LLYW0ho7X71pl6cGHzlwGdf9jQPfWj2aOeJ+vQGuve0cCqrX7
j4JACOuU3Q0sVau3OPQ7vBqwe82mGfUuFrvk4FPLxsQQaxnzj/rB3XdEcX5h
Sbp/+QpmMBevcrjXLZSz+85cX2cMoWVtvQsB1BOGMdATxFrW1RsSJTLHdgLu
pjueJNxppq1olkFVeQ6PxXY7GttG6IeCPpjprOPT+fGqPoZZi45bQXnb1yIo
aG3qCSfVnzdo1BHTE+Ik45A1kTuW5nBIClcW+BKRfhCBqN5x8JxAMV+6UQOF
IV5XH9hnnoLXISzqgPSwYLeHuWl2qt3vgZVZVXcfhgRvMCKk9sUhtWIaJGEQ
o2LaRxzv8fhtunk++GUCp4kFD5EuTKw9JsXXD1rWLcNZ0fIFyUgMEWvl4vM5
sTQbyCp7DCgQJESoSewxhpX9E8VqqtKaU94QlnvIbqTTHw2vappn7TDnNEyc
LvIgJ0cONCWl4/W0rnmNvWGWrk1H/QrFyXODyFr7OA8iAuX9jQfIcd45xUZG
HTi2v6zdCUxBiUXH5osoMLNWMRICJ4s6Es4HNdu5D31Bt2np4eSRvESfm7bO
a0LbXKP/45E63WKDPq53/pnxPMPqlfPcN3a1sUgVMJ5KX5EKvKc5Alcpk9Zy
3FtChhOcG4wEW4u27VuIu9JLaEs6OgdYQ/MZKcs/6O6zMEXQi8zHVKOJEvbC
swfjfHuEhCLHeoITSVh7HF3n3aFrB9hC/tKOPLi5GGbw1fAcZNolEf2lwia8
1Fn8DOgUPbuagcVV45Rlp+crGNfxw21T2iqxBw8mrMkNS2O/dV30He9mQ1nC
Brov1lIz2aY33uIbQpuGHzjpS0BXUyi6HxRTcvUUIW1rDWbrY6zJWYda0+Dg
ec4r20QKlA7Espk12vg7DWDitEgVr8ba9qZtxg8Os3X65sSPvgG5LWY/Wnwx
1J4BBKDlTfVbY5cEW3/MTphfT8xJSKbGDDkzDBDB/7zq2mNHDTpE4rlHUHOD
tz73j/LmaTXw2cJAHFZt5kgVZhZVL2b7i9cLUaiIr5rrY2LLn/GA6TW4POxc
mi0+vTUM+cbZhQMkIZ/xzicTGrOsM/gdAevDU3p9BOSmRDTtUu7ppbOY/oQD
4U+rvUsiU1cKYJ1u85gSIEaIlR5eiGfj+SBqCFSfN3PPuHyY7g4F8o5kDgaU
ub4Uu8iEstukD/AYTGFpe2d4Eqq3/L4ED5Y1G6PSVCA3rbJ5SKW3h0wKT0H4
gTiU4OqQH0+JR5rSTsLbw4tWhdSlMNed2UcP2G+govJjFj3qBplfnOpcVISw
WjWEd/AeydInq+DzeMayTNsfLhPaMwb2Cl2PaSePOGGbafwaD45VjPSvx7+9
z3Hq2LqrZjTFBr4IEiJASRRkKo6/kXyhg/8hXCIyjxLu1scazsQlqYEZf/8/
S/L9ZOp755l5XSf71Z0XygIbxQMAMZZ9FhckEpspizVr8/QRvVmSYnA2fx1X
cs9Vt73qysPQYe/L0Gu5Wj1zd6VU25gWo5VMK0rMJi5vENqQhs7GgD2NEn+d
dGdtm64wYfK+QcNFIXkkXYkIoqGwJM6LgpOYrWPZfkyCe1DRFvueoXwt75Iy
3YF0BeznqBhiH5l85X0xANQl3fpShXRy5qwu/PE5FsF6m4+OBAm1q4azIuqA
YaI5GUsi+P7JNt6CPTUKBCjczqHT/Ay0xgWUuWjuSH2G1B23fM2wHmt6t7CU
8X5/KEQjzpyTwMEs9JyQfd46SPoAl1kh7HPUpNhwjI3d9jbfsmpTKBzt5gF9
YtRggLzwOPuqxWYEPPJifpEegqAJH7+AgEUeySIIT3xEX/wQdxWxyThQSDW/
Q8/uFfJe7Khxfmp+rjiivrmjwg8wNhbBSpnxE7+UGlibiUCFxF/gd+Ue1Nkg
g2OyZvJ0ixJfw8aEkw7lp3xmlWsu8303amOB2gOTDTLm0WanG02sl8CH5iYg
RnU9/x3kSIP1dYfnAIUmcSGjI0kUeVZkrY+vlJEZFYCGNjt0BVPB44MFFH9f
+mvRpSc/yB4zV4KHi95SYuEYbIEYWCmbD0IX1rqmwTNJ5TmKhqjF/rTNqGTc
jaYiMYkFo2R/WanfuPT0JnXHkU+Y4vayObtD+mdiK7SmyEtNBu9w94MHapwK
kWdjopUXQxcJ2149V3b1JNnJ4PZU65CapejSEOKcw4y39KHMxG1wISkpZ17n
sJ7OwZGn2hftA7cHkIzYhZqRraJOjndishfIRuc016vwqPpX8vv7ttFMznQq
c/11p7xqsTLTA9tRUYxwafQz6JDT7ztJil9XYiT/sZbUyatyx6ToHyXzVKSy
RV1BLhwZzGZs0MQMfqLgm763hae0+dRfsLbz7T9KBP483rytIcx+z6pXGAny
ty7ql7mNMtpJwldmt6yQAeuixLlWPNddBFI7qmutarsWQ360vxZHhm57YUYo
olEXMAae7oA9wf41fW8wk3YqqiubZQ+6FbozbVlkAZ14Mn4OVxUqJjKwfK+G
X9buM9LDD68kMfJmsM1mt2Sp1GJZOKnrdZXbnE3rxRJitMxoNPOdCQBoRkHK
MIoQUKDAyFHwghtO2K7zYsr2BQuKvGxy1IXXvSsHRZUlLF9ZIGGdulNTM7uD
cnzYWVkqSEpR8gN66mAolYdDjHYMIoZC5Ov7Me01P3Uw83zGaMGSxXPemDB/
v1Wk/21tT0Dt9Qu1jcq0+U+ES/Ky1b6dfYcC5zbQ0NSx3FUxOBQ7Bnywjs+N
lloAlR2xDUTOL9Nt4ADbgMkZm0FcgKh2WiW/cuFLHwexXlZQCfKSbES+sgGi
6YfqZX+5khWcBnnTyEzy4Sy0nOP/gppUoB1GSc0kunMGXHZQjhafA6XJ1Xqf
F/XdTuve8YfJXjHSaRqkUXd/tF0pB35jd6r8g7bfPLY9ufjn8w//TpRTfJHv
XloAH/M8/XLFLj6m3DJHh9ObNX4TozVG+x/gopLAug6Hg7w1tvGIgiAfr5ja
2uTyubW6vF4JvyOrNbQx2PHERy3D5QecLCwFX5NJ1eaWapGr523PcIpOuoqU
cR5B2ldjRY0l/qx++cmqVj1C+1WV/4WfMfSZwGEC1M37D34FjmiIoOZoYTvC
6lL26/WGl3b+OxsU5ozZJb9XUDaAOM0fjJDHnnI482V5JKZ/Mlwe8eL25mb2
Ko2SOBN5MtXiHGHGalGKjyaI7ZgK0jPUVkWTCpUbdoQuln/0Y+Yqq7HNqAUe
6LfSJbIunWc9UcvrxnTYafIXzrrTo73TzQwdGbGF6NOWxFVcjMvybvAof7U4
cQaxYfnHS/b2CLXgr3x2XwIj0Qxr6h0wv9pEVZuGhLacK8gERudC0dP18zKN
2QA1oc+J5OPo/xCtQLoFpNqF04QK4Mf1QW0ORFFvfpg6rPZvRujLmKcAKF3C
0Div4wY74UYhu5ucRI/9SRFnfhqhefkCPxi0x2A76FOwyyl7tEDuoSuLtDN1
YdTGQTRtbhNZ/3DFJolNoXQHFcC1cS1frYTNU3dXzqGxEvLARe/5HkcPoOCe
XD+Rg647+ItA1++ikth4zBguuIR/oU/TkJI6QyWKaOQUVuAlazNoBBCMx4kM
J67gCrX/uy2/Hb2G2N5Qe5VJ/bOu94Vo0DOhjxUWDukJ5QE4n6mRb/TFSLvb
idXYhpqQMuCPKGyQhsBO3SuMgHUnrWe4SdtQA3fz1UJrgEkaF9OadLXltNrW
UsPCXhtXMxBy7GIgoGVrWYrQrSholGpJVjBVizCLKOHBAnkB7CkCAknmrlOs
a87AXl4w00pk3TjFH0azD5tmoyEyJoim30eY9I3Z7EhZp3UNic+IKpoFma2F
ih9czlH316AW7QAUAz1fITWBA1nX3uTUvIWmi/vNPfbZIQVW+6IBzWhiKcZD
a1+4uKUo6VgrU2XgsSZ0uzwbr44imt11NLZLDfKK6vV1XVmfWrbDLv+Hw0qX
Jm7KrpWFlf7at4GEBlw6gK9E4FsR1oyVCYT0ua85QfDgaOtS5ncMnZzRnxX4
UNWdtSWVQoOB0bElUlVvIS3HfZwLDCMztKgVk1aogCLOXknNGLslYAGpS5sy
z/043oh894koWeu284GMo2skZhcLSVcKR7ED+4SL50lgkP49wjvchdxOe867
DnvXsfhJHW7SUMQl7nfzs90NtIg+qQgNW900VvwhDjJgoAHE6sDZspUA6BNp
CzOXITpgAByFZF1mXW244r3I+mnVH5SnBEvPyWsrN+m9PfK1i19DliqgL9pt
KxNj+5OTIZ/BqpSMr4hM/8LQxuv5DXK8V+2XFN7of/mgLYzz+B0gvINvTWa6
6jGfBC+WZ+hMUF4lmQ9ZtLQB49fTBuZ+oR20n53y8ksEvWDHjKTTPpF7Wb9o
wx7Ooc0v1hhFYn0GWHSpVLkrU/Pt2hZ0RuMLJIfIaRKS0aKdSgYncsWsFHHm
SI3aT/Aw2IV0aO3LdfQ5immi/o1Yw1EDPey5XAQVbMuzjYmVyFxmYByWeXc5
qPfLnZ5sQkH356f0dPtYCGx1yAPtXMAPsY8nB6d7BkFi5CUdVSEYhRSfZUMG
tKZEMNmVMClVyDophMc6Pc9nkA2f3ivEAZhp00KvHNa/ciiT83W24lXhVkgR
M99frBNAQTipI0Yynx7Aa+/SiNsFxlzz4zj9Iztd+4dzlSqsyS028xtd9WEX
wU/r58UFMJQWAX0zrYr1zPCcqzmIg72sh0aFeCQN2/NAa5wPVgbCetz+wZ01
SKwm7WtRS3ilk0fvBkBrN8kkc0O+OfmMNA/mg7l6d3U2w9VIFfqivSvcDBDt
ztD7J0vyxCfGz6ngQ86GWPgjKfAy7d/lEfhHrC0bt7nD+HqYVItT/bP44/Nd
1DQauChatYqyBTlO1ptzNUllBlGnbXOxmcPzdgwLcGpJcgC7UpZhMJi3qNn3
/hUj2l1Xd2UMB0glzPbsDXUfcGkWmIftYX7w9cmgYyHje4TyEEM6Zk9ek9jE
KT6/Ji02Xk7eZpyNE4FmXrBB3FiL9WlxC0KjT1TyXCd4WjbpfY+DaLroGuL8
z4pMskn2EtECi6eo6ZQc5Xa5tYHzs4uGaA8M+dEC53Q6Mwy5AMNUGiVEt/x0
GkZSCF5cgGuBdF5szEkTaZKL2LxXToa35x3dQX5NJS4te/CYjJlt04w/pu3e
INQh52bhLEqOSc/jJXHbOkNPprBpds4NPmhlLZ4XWV4BwlYl9mnaC7wf3W0i
YIvX1VtuGAC2k71fnGAWDeRPTkLXuVZqJ+04IOimirJaMB72pgfTfWaeZL5Q
it/ogYEwrxAmD1ij4QMOKVVjZA9PiEDA80tVD+iLItbbonJDXlSzzztO0KFL
TIOMp6yYB+P19kZSrx69UMjl9wcBR7SsQmdDDqn2PNjJnz5tovhffmI6WQPF
2dSTaIo5AQVGupK95vCdenAvoiC4VbblqtIBZ+oqhDo8qvcrr0voasOAN2hH
0q0J+0JfYEhqiPVcxryVWc0Cx5SsACcUj8j17VpJmCV9vDesL1clxApkiMEf
1tEJJVq7Gp3rI7saxyfike9mALb1S7jyTbz1bymdIgUmSgpHPpWxDmzxBe30
wMNYrnED7OIhzQAo9qfvgXL1Da+oJW6xiuAFi4tJGpERR7cTKeAz/YEKrJrP
nNi703btmmuX4RkTrZh14kuAl0+X6fDD/08CY7ihE9+YP4yY44r/hRJSwmX2
GnxEPXZKROS85nnG5pxBXd+klLSSm36eUQ8UYfheBvmnG3TIN94qZ6nLdhER
WQ2s9YWgAnmV0u/Da5UUJ0vksY58OarcZcMk/tD62/Hxr6Wgo8pl1yBb2fY5
fKAVrPRyuT7AWWedou62BtikPmX6UX1qkCMSh5BQ7iUAzAeM6vmokAyKfOyV
J8GT1pKmFyMXtSQXUU78DwxPAQ1phfStQRleX26EKOTWNgZFcMBR8e3p8rWM
MezqyNugSUp0eTMzmMSzg0dlz4NgicUL9pnG/HnFqbFP+Lmt8245j96sR3qv
ZF8qIR6ND/1kuTFaF5j8F1DwogvpFS00KHdQPJ6wB1rE5Sy5SVqcGLVghBTx
OG4ISZYqMPYTht0garX9TBqSTJiS+WqhaSItc7MtY+vP/vIHpegp1SO7ZSc7
Nlbwitz73Fq36KPwhrpgRTRaWv4rUM1LI5aE3skQ6wnRh/o8oQTW5TF5kZq5
w2uTl2LMMkBxzDAU9kyMetXS8xCu7985mW2nmScWBFFqezG3ue2/PeoUUzcJ
4c2IdCUb1S7ZWdvXrrIDOVqWvxpFDI+fMq4ZjxHuRRJZRakqwZDpFPUxLg4R
Z6Ikpw8j3r2fCdFpIWAwHZ277pZIwVrv7WFVJjQBgLrvrJ8PfZjYMf+McCD1
FPDH2Opnf0hPFBpmk3FNj4bt5FcqGy/kdaO4L0mNRe5OoHIuhFlXs6rdjprm
USBa1U+LxyHZtZvb3uJLSIeFfmPvCYjXH+5haJp/mww+UKAb6iM20dx+w74x
dpj1RDTVQocafREr+qKmOi94tI70rpknzdnFCT96BXlYARYrRL1a/Zkd2+Xl
s2EDMsMkMLlisR9vGMcZYZLFjS8QVSVhbYERccLVq4lsKBb5SKX5EFhunLQq
dHy3nCFtH34E1ykdUNQ1QkD5h5ZtlfTI0yOdmvsWWem/gHtowwuqlTuwghDh
zlwPzFfGIgYDFkLTg0Ka83tNsExbDUg3g1bYn1FNa5v7arXn1lR/96Yl5liq
CyJBPQ1ULAPoiOzRCBZsptjUq4beM1gm0qFAuxe2zDPKEbt1uiRKiD5083kn
amEnHO/qPXApBU/QlhUwF8aVsziunPEn+9PYe6CZWJJNdSzoZ82jHjL9cKFg
yv0UcGBoi4ACZll9AK6jjqA/RTHD2ZvCNArt8LplCzkn0v77V57Tdb8Bum/D
6YihuaFChePKnQkSy5ERaHgEDtPZcGffsYEpg7DbFLuAKyCfuYIPAMKz+hb6
fAwxAhK5ibqJUOLbQPT3xA2n/MYJTaZRStCkybmRFHsGucp5Jnaq4s2jSi3P
9n/dn5ozV5yScJrd+bbRq6Dk+9JNWQGcw5T6CsTSOqLdUIUiBUsjvANztafs
1iQWNApK0BrZonVnPldr69ZGnHfWSdI7RvwdVLs575brfJwTP1/zhxRPDpg1
63h8FysBIGsApxZ6sxw4QnNZLTY5tmQH8GsokmUk7Zfp93MDL2B0dgXEK6rq
SwtOLDGuf045ziwUIG/Kq2bmULQIb1TfyilL8rx2AKuQAGu1RmouHppcp3T3
V2/A3DJ+liowqimVRD1BR0qAaYfsUH0D7KCR9IaIUhJBavYLBznnkE0Z4Pc4
yhqnCpS/fDhD9Q9kNQqqnVFR9jtTJSBn9ig0n/c7J8ESsddwebK17RsO/CNX
88j+3usCOpOXwMoaldOc1qSABhhyxF0aCYOMfJ3y7wa+pkzVT98RHndGjmNV
xZg8aakwVmXSF5mqyosNtwzu7RD1DbfCUAjmXCYmi58fjYOmbNNcKXjpAT1r
t6NLgp+FYndWspnCBWbBxNSRnW1QMcYjuOb5HVmqwOZ8ZSt+wxIu95jsxAx5
oKMv1OK2FMA0R5HRdKYMdRNsMTNalpNtNArEallOQxk+CMXABluOibUHjOJF
Yk7jApMyLGVap4941NdrJK0wP19YN4P92CWhJRcLxmvIWEURp/OLqXToGFeq
qPtn9hY453Btxh4pEFw475hXQfPB0his/LEncCr2Q7069unb9zgeH8p1ycj4
PQl1AyBdj+zseNRDPLhd7fasjMf8w/sImcYtOppAk0Yuq2IoYLlxOK6pAgA+
mVU0HcxeJQoYMoDw2f7rrbDhCbH9vir18/I0hCMofNG7ELu6+/LASdwUqcaO
tz5AI+TSHSoC4ePYCxjPQqEsFJfy1jwIz5xuNohM9txCg5pqLAYGz4EjwKlG
/6D+GEpTr7ELHNaMgdjrBM4/cnAEIGQcnwi8Jhxz8nl+ubuQW0Y0WwfFpLT/
xfovi1XHody4Mlm/lak3NHMgu0aKbNcf+M5FrnFa4s62xRFT/WV1I+R4XoFf
Qtu3DCrK2WYmqpTQtcVrYQhTw3GrGwvIBwDZUAxd3YnRdRq99BT6llTIuILA
VsHXSr+t43k5m1ur3xDoTjUz5ihTLWyv8Ki1dpfxwZxss3d9geCZiUlazXLw
ApNHdyL2w8LlmtBpxlLk3puZ5xLHlmHefDl3mVPILzW7QSksvzDPYAOyEJoP
XfhHhcwGOQNKdq69zhFHOwYN9Td3Hvu5OMGoFLdxwPlfs1l1utewfGW69Zn7
1Y7kvcuNrrMfHRYH5mMp+NaVP10dTuAeixG3mDksxcIn2bdI8y3Q7afeX8yC
pzebQbF2kDiXH+/VKOimzeyDfCiq/sVlzuEZJZjidzJjLu08QqT+QP8oiYAQ
qwvXKBuxR8DzxNVStZBIDesfuKLEtMlBjs3CAqfUtKjK9qgwKUlkSggZmoXi
0C2NQuyIQGfvF9MXL0au1WlOKTpemBPis0NY4HGSqcWfvqsaVADBsp9KXkyV
7ckWx9BO2wqIKedEmpyjc01EHnlmEUaUTMHShDEggDcifo7Pw/mG3Bla1i4d
VDBdWQpk0p9if71QZkAub8uPvi9BBx1+tfQMwBml6qQycVjQbqkZpQb2I8Fo
mJNU+M+CGY0m8bZc8GcktSyuzkpc7Pmh6mOBwWz9a9BW8ydVfL67Nm1UH+ys
bNAlENGuz8YrtCWR/L8Np27SYJDBCssP18jMrr0WEq/kz7GfHfQXelAitUTt
DUHoyqsF42rYL1Zr+WGLLwxNO0wiOTz6D/6ihCpfOyab5mSUFGXBceKVB+jZ
Di4tGH06OqK+FEDVoeCQxI2o3lAr4bIklTYov3v9HmIYuV+/tSMX/q0c0kAK
5CPcDMOaAqcgdqzQ7J24zm/lWToDEWEgOERbl8c4Q6k6D8Xlyl1TUwmC02ro
T5hbvt3ojzLwVWivOefvQq9Ouz1oT6c0XAc9fB+8b72wVIlfw3BCRvlTD/k+
qBz8kXSNT6BtSDFdB52IpxAG77qY61cXPoXpCoZ/ihQSGFlbihfOU0zS0dFB
mxUAWYcYR8Vcpkr5UPsNY50urewHIPUXu1tNzKt543ihMKF8CBg5MmEc26ow
G4+2V9v0n9UUh9TyT5fd9AurObE8sSeGX6Tvh9V9OgzCrQvQBYqfxJjkgVsY
h8JhECSjZdYuA38vBTP3PNkCWyrSpslV+H4UMIcsKRtIH81M/eMq3EUHgioL
o8yhcxaar6x6e/2V7RggLDpeszga518WLczBAgxaQjRq0LuuZX6AEYSOxYpA
5uP7dbNzS5eS+HZCWSwNxuRJAYVOUB8yTaf0INnnfcPq3tF5KchN8ruFHqFm
z3AHphBiq2OycOcJGB3CbJYC84NAIsQweX8WABlhducyHnt4mclhTqrdcEzS
Q12/pmMp5FWWcY+WstwaIyIWxT/ZWk8itNAmX04xZwHlSbQtz3lvW2oEsDK6
eMvjNR8hCPaZOt/4cLUH5UnXdowMWnFcsN6J7xA41Dg6nFc9iOvc+5RyjGYR
U3Amm4kr5iVpLLSBgrxa9qsi0A6n6La9Gv+Vzl1J+6j4DVNnxD2MR8bFB28d
uIlIFA7STjXfh+pa23XilQMhCaHph1UUwHqvob1jEk0BUw0tyZb6fK3NasSV
wGEqL/0J1Nu74nD5l6VDWvTVo6s5EHtcvxLrULZcib8CmPoW6qod9PfKQrES
AFq/aahPzTnKAZ23Bwk60BdxtyXlHoKDnvscprcFM0jkqxEF50oHk62ce6s9
DMtFS2U4UljtERjEhaQ9YP3OaHK6VT7j94teLS0ngMk/gqiFkT/LI3YxLKur
+bjDelZdZ7SFxav++6YECE6qKj7wuEtpaRV1hbX2XZ8BSi/ZKJtRjLH8esSw
A7hDNx2YbfGLKoLlnw7n/Vs/D9cCBM2Dc0bA3/Xfs/4ni6NnTodWqeWzHKIa
Lmr8FGF3Quknc4SQmkNa2+p+icDKychqk8YmB2yslHnzpHr9zSRqRUhS1FFk
spWxFbXHvwdW2x/WseGpl7lprpBEUjoIOp486KFiPQSli5Csh8dmggVPikeE
ds2rNujk+O+FEFKreHakK04TE2BGnHGM6d2QPu6Mb9/pR2DuUmuhEEQ+JOOT
bzV3gALKNd+250Fm84nl1tCe6AIDa71r23wgnow8AN+A4APWZyrLkVjMNDlC
U8WK8C5asMY9tomL7zab4mUh7XbTsqdLuoSgadlxdTnWfOIheyrHkjLzcmwB
F9NM27xZiooAtvFdAGnQJnBosNXBN86AwAtvvGYMjxgWfBrygPru9OR1HPBK
LM6MTLzuNv4ddt57AQOKAOCRxgj/YhfkRDmRJoNC3dgSZM/xumAj5MwiaYsS
zRmw7eNhA3rSw0W3ndy0umFQhnSe7FBdW+hngzIIqQWW4hrqg3CmJvMPepCs
OcCUOK0EpwkIl5dBOu4EwUJTiVbK0SibPCz22xvqvfuMCf4ayMeXptHzJuz3
sp9bXYICjqQ8Kljv/uOqYyCqm2TRKr0IkNFM3RT9JkDKMiMQ+s9CUbnIO+o+
L5D1q6FqWpXuH1u01pb8ljVZyrbcbh+YGsMTpYL5y08eW3G+x+Klil0XanTr
JZ92VvMh8FSXgceeEsz9nO6SVThzpfcZGQLL05dYcN2fmvF0SW0W4qqlsqpt
yZbRBmFnywiX1VJyj18KLLdh7OtEmPvOt4pr9OUftrLFRslQXN006TdsI5FL
1dMBXt9iL3GzMoTqMCIxtDFyJeXA55o11LftbQ9FJd/JgJU1v5GbCv/irCbY
DT926dWVxqN9DJcB6iVzErsfqCjxqSGnObZw0+hd1v3XWMpjRIjEeezFY6wj
BauZNyuDstk5cfapXYDdO3X8WQveFJaYxV2GZ6z34G8gujYpDeX3I3v/+kCb
qX9AmuNc92I3CTw5cWq6w5k8W7crVNE0gTNigjMbK7j628nj0Lau40/2eB7v
RrrB4h2stgpstaGJWApd6XHakhJRCYj8wfjvWMDD0YG9i9qiUjySbG+sWNlM
Yaq0+CBrMjafpBxofpq7BZv6X7W7tctyIw0HUJ59Fv4nQLpiGXEqezL/PNX6
ZGLbE3jPTz6KY/jo+tZytQT6Nba1a2gctCdm166nRijAnsG9BSz4LxqVbfsK
n/1KRBz2d9raIX4s6wVASPGf/ZwUIlv2F7BfSAZu/JSs9wiFU4wENs16Yuej
QsQ/OmF8RT58oHwesNI/B+wO59o/q5U1+KSnHr9/CGS5NDyiyQgLzKZQOX09
d/0zKC8HbT5Jb2v66vtaTMNilyIXJW1hOvQIkxBcIAAr9R0agzgt6eB2oU5u
kY8Tp9JRCql/12/RHEy6oVR7m1kHowszbUEh+PIuRuud3BG43dvjHXr0Jasj
IGAM5esVdteKO/cl7T7HMLkxtKaTtPSpoS3OLUHlHSpMboYNnOb5ajh20uuX
yoCyHXMUukI75tTZ/09A26M5789tCrbhAK56HF1WiizflFgtmyVcxeC8IMhJ
GSrZhaXEbszm2XDiE7Doa4fEStswT0FdWniGevNOk4+iN4dBFlFTWiTPVfSv
fq5VvzGcNud7JDxaoIOBQUTkbG7jl4595I0XG1LDCb/pbUYrvmaViSDiHoTY
NgZLCTwO60oFBlC1swRSC7t6D9xW/Bjq0ouuJZNDWDTaUcOqI040eLBLKQYI
rYV6CnKHrrSd4jX1IQhTEfP4yDetC+vHW+wquvkQ8mVZ4lRvSX1NGlBxgoH7
jH5BEUZWDLHtd0auEzGkAguPMN2i3d/cpGyBPbFAe2SATcCTIG3E5aQcfPoE
eyI3o3wc2r8Z5r0LddlZHbxE8kefEtQMariubdMe94gopkW4nkBlVOn/3Upd
Pr0svO9+3Nl/ibz0c5mEE22HI6CvzYLQ6ChGBpPcPiA4Nt1d+42KKkyJ8LxS
qaMlPKTT4MLPPc4OsqYduMWoLtNBr4ebQyih8Nw6vlGDOjFF6xmQwthqDAWb
Jq3XeQaEPKiOn6Zqv1Wvz9wfOhVTQO6UYbFkL5O9LHLQiNrIWwCrrGgxdKsr
TtKFOymFCS4F5IhLvhpCnLAta6QwAKEVD2NShs3SfyirpyGrUUskP7SNn1+7
ZakCOZMqPzlEiPQzbayy5DpgxTyH9w+JDE39/rxmcVd1V6i8ZFNO5EUvDOAg
Wg/wHerwX4i/PvOEMJlcq4jyPGfzMs/EQYVHYN6KyZtW+DbHTICSYvHMgf2d
5kEpqs/oq8YVXMj6QU9W3L+JA9TRReZM6k0KcSXlGnF3d/MMhCp3Aq8J80qj
0qDF0SipRc2ilNGoWU73U3qNhg1vfuplj6Us0WOLEpqLtM/xQkmDPB1AmgDG
UEHTzb3Hko9GsMEwege0eAMeCLY4gCFewXctSciv5sJSDwP6eyrS6rIINbau
2IpfmF1SIQgFZpwmUiyRTRYf/zLCiirshMKF1sKw+ZbsDisMZv1rHH0xaIWl
4RpIpcJIW9D82d/1EqEzmVzXq72enXFKYTjty7mQp9Dlcjvj0FUCJOG3dcrv
mh0AN5F5ddI7nvH92VKuonk6Y4ZsGMKwa2rHnRI3BaMS+0vyOjuJEwWI+2uC
IyXZGushRQ5EIZwFPU40qNkE3sMBk9N398PC+F8h1qzvnaUOUJclfqraw7M/
9MasoGdfkH9xFja5AH7PdsQWutK8+6vY04e52BjiFef+y40j5oCAt8EwrJIc
Y738OEDfYdQQmZ+L76fU/yDwWbOTffiof3+RrRjBipSFFMu9XT1NKyhtbjp4
nFNlStbkMAJGBknYBdDJ1KtmuCYlhQm5r7G5OAWGwCXfQnesQ6hRtI9kDz9b
/6mE6LjOOx3vpaMrdbklJR5O0WkzG1e804Ves3EQNXEuKemxPwZN0LoA+1BV
Ti1pO/Q5e+U1uJjfXdG5OOb7n2JfOFcdUb9si1Mxy4Jfomwpz3Un5s91Y4+/
gZ4sicohOw4SOYbyzs2chgXDpTw9zAtnYufrEXenGUq1nV2iYM1E6ItDD2IS
t68XVa1UQZRk3eC0wB8/qKCsQisH6R04JGgfWYaIK1MQK90Pm2I+aJgO5cOO
iRFvlLk9jWy/LYSWA6pX6yM4J/G31mcl2sgjavjVbQcXJQQUMv4wncdZFUH8
snCEQc9HpuisVFbmtMKzm7qErS6ygzA0dw7W/4I8ciea/G1hj5YLzhfKvzNG
hrPPe3LkbOJFxqhItH8cLxSruyKMSFW9x11Bed3OV1KhvNgYA3qrCHv8SR/H
rRxKuSVGlQeSLhSZtDAJe87g3pNjthQWQIVQHOk8BjmLCp5MxGcO+WjtwwmW
UetKUo8y+ieHeTe0/6/oZWK7uHfBYNqohitYf8ImBL/Cc6ZXJ4/dbAiTXvWo
F/82LT8YVLHSCiJ0XCrYwNyh8FYA/FbjHzUbgYLYjlpeJVyPVg5UXfDc44UL
3KuZuMU46exUg03arqLxiuQPPBtj+AT4J4b+Ro7hge3j5E17DRyh+qtn19CN
ASaLBnuzAaCwpBt/Yyp5TSQGE9RFRpOCVRNJVtGNIZVn4m7BqHzzCPZfqp+M
aCpv0XCfn0oZEFfLiwLzpNFA6ma6hQpiTFqKGZuAJsm1Wxex3tVeHjmctk1u
mZSTSloTWKP4zPILhDzO42Ty8x/OJwbb5TWMkpgAcbvHnURfynmEmHkRX27C
FWz7u/C3TijsS+QSkL3q5sBnxWKpwx46s71ETuJPPsE+w8sCvLkVgZHGnHX1
gAc4EMnHW1OS8SP4CyGP0DPuADl5xEf6K0XPXR76M0mP3s/4oUO/Om9PIDkd
t7LASPrKpOq1+MA1+9UqFKEDSg0GbeXsntCJoUKz4fuye9MlzX/AQhjukY2D
ZYO6/qpYc9oKaTK29XpNoY7wlIUsPQr1rrFTs5dEKqSULgdDe2hS82doIqG2
KQHbISPmcd7vyzbB9Qt/Je5D768BD/19WowsN03Bn6lkuDcw8oHmK2H/8bw+
LNK6npIYM8CenaIXz7QgXjsVIeUJYg4NwG3gO1wEgES+ujfIWWp1u9agjQe6
LdiYsJAUJ32dg4pe7PL/ycJx3yLnJa8JMORgUtaI/1z+TeHt9mABWfZ3xJlD
elWyAh3+0OfrT12qKsp+e/2SFc4OrJjFC0iiNLKYgLWlQgTQY2+vzQiGW/Ob
H4WcV9n1kAY30Usa4jxd6bEKjJVx4forfjOuWtmNNuOIMSQDtGjGIfwhYaR9
BtFtDRNlOa3Ag6XzJxP7OeLbU4bW0qCBvqSFaDT+az7SFgtlx7udrqzlHbKf
xpHBbawV5s+/I8PqVpVqwmLY3AzItZoPdpmft9gGRO4BF2GGMv3AJHMflmNE
uydMpCd4bxo2MPzwo3iKWr8bB/u0U/I5vYMRXGsASz+siKRKHkphfBATu4zw
llHIez1wv8xTFNEC2RyvFJeJqzhupfqoqdWvWeLeikGsUQPkCH2EhFSGEt+U
x4YO5bYr21jM05vCHrMfb8TzG8YNo4spWyplO7x00ObP13IbxDzlwqHqriMA
B/W23bsZBXvdOzbQYWx61AA8xuC7wOMOGAH9+bHa0oUNwlpyBT0NyAeSK8ma
Kqpv+2ki8QpNuWPDOIp17Yk5NdCdYZE+h1UxbF/2fEbE8WLAUJuAunoJBYU0
s7zqnnkz+btD7R0iOaVKB1+5WjWznlGNRGdQfQXESGXDDbH7647Uvh/cTjon
w1UXYozRxTtOErdWZpqXQe+EigvLXkd76fCYdKn85htXMRVe8OFfb6i54ijv
37U4X/znuUIkEHjsWjlvNkiyaQw5k9pX3+BCxXxgP+sMIY4D8UQowe+GhOMF
6yPGXrl/fKv/T4lyUffc59Vk8S0e5sQ1+tgwsVaqvxvC6/z5HwnP7u88Opmm
IcLlvKiwnOnyehZoyr25f3FpdeeiawN0GZCFkh8sic8VwwkWKtIeoDApf6pj
cySmWArQZ97CrO+Ch9fLWKP+xrTt837wiIsaURBxwwvokZJkygXZEdBs4din
kQhfW7vLQxskVenSw+t3lD0ZobC/7hwN/him3UYf2qpeayrw65B8cOLz+NUt
+47Jm8+EceGuSKocPIo+memYdSL6EHn6oLj/111dPicO83VoZ/IOQG+9TO6Z
zlTUsgRmna64TVIv9VoIUPjwgfLv/9TFdekAyQ/BVfXPKnBb2wrGgb2vB1Sj
qGvHG8sBHc7elXktx+jyf8+s9yl9Su+tC2iGep0xEBEiF4CY5tu6Mqg67X8D
bysJ06L72bjJukARQdGhP/xdEovOFmXZtohFhoYjL2qVYko6WZWlzV/ZOOB8
y8oB1EDtxe+sLcjPb+9GcFmQ2x/DcnkIZjpl4PrKensNGdJOaGRcc3AfL6N4
+6LPmHCA8xQtBklJACehKgADi4NAFTtpWY/rKxar1HLy/dgPyo66H/K44xbL
AHU9d4mAthdVNU4zWDs6c1Ep3YXEUY9Y1pWhHnd4INwdvmLt3SnGxFkJvUPB
chtjbn5MZYO4eZ1ZKd+oPuzVsIrlzEdwQZBGH5+Kt5EGvss7w5+q/yV7OfdL
+Yi0X6uru9wO+eA+qZ2bz8f/zK+ein6U75R6ohbnfOxUfZ2rMmJOsrEmK1kg
Be8LmpWFgkrnMjST1F6lIqGc9rqIjdnUp133NwY3rA8goJ9yCbuOvxHXmRi0
2JuQw9ThgQM6W+01JqO0ggbG8A7B01t8XvBJf2gqzCXpxBrmAc58Vht8icSH
4vhULOfJ/7BSViyO0F0xmwlz6LOMZ/LOiq/LSSdnge5w64zJ9JUQP1VAAC/5
bFVqpZNDH8EFJKs8kxPssFxDmPPAWYRjdJR2kToPmLLMkD16GahUXUXRDPrZ
IXnWk5MeQs6Jc+T1eEmwZDV36qaFjLR8ClVcYyDYjBCs0IOFzNLnb9M2Wdxd
T6n/l1tUYmAV4fP9hslWr2FT3JhXalXVoh9y69cHsB7cFYasTejSGbNSu8uu
DnVxxbs/xRLNck+3Jse0aqzn7wBKEOV3M3mefcHmuls1ejjBQiIRsq51qUXC
yOuZPhwUzxQV4T0GvwRaTmn5Pfm76MS7RKSHyqYU2l0K8sQX4fwOEZKsImWz
QFHI0BtuZnzJn3f8EW+AGAjPMVow8ESbvRLg8EWdjNWS1ai2G6UZ0ge74pW2
77NiCYXZnLKO1GATJz+zlOqbveU/hZkQQLuQ5oqIy/JRRgyb6CzHNMbvXwMw
97FO3eRwvsvIinsWdG9jl/5OAZqqmahv8HB1C+uu2iBGSVshvJfVWlkqpWVH
tY1bkJUH9DXsiG4oQqqw/OIwPmP3w9g+f0hvsQMvedbUsyAVqOv34aYvnuGU
QSUWde0tcRhAdnWv5/SwMNioivSb0XnbA+ESqHnCSwZDCszjSDRfU6QN9i9N
AtLyBqneYlKby7U8RQFtKtixktqpv6TRlrRXDO9+gSKc9995CvU2h+m5Go99
N/b71UZjnbCJnTQN4cStYT+XTl6Av7LZ1s9+kXv1r3TIxdE/LUzJzUvX8FhX
VCZe9fpzrPthsemeY4yM4o1s2FWATWRx0Aj2FJ/zq38v4MO5AKgYmO+O+hm2
36qFrhKIk7LdKJyV5sYQSzsCKaeDRfjw9QRQlhK3+d5qqznC9tzMSvULOai0
xYXBSXsS9si/WGrdpi811peauxf05CKCcnjPX2lS/8i7yWikPBX+VCwHRgAd
pp1m+T3mqLzse/kHleVjWeGUF1zaT4WEZzl+48/jGPUB1QBbufDwlmqXWe5v
AR81Fi4ujf4vc2xWLty6ABs3oIcUPNjfYQH6MNbFj/dH9kDfZuHq0KSxaSin
4qufTF7kRNg90okGJMiHpMdoxZWwML6ggNxVV+nc083LaUmgHLyS2208yNFu
OZKrbj4yUJ1c02Sf6cV2Ot+4+zIc62ywdgZq2ch3Lu47mxn2YNRIL8/Xf1pV
lzITyCztZ0drZ5dTXZsGtFe/9kQvK8umyZFrctioMbl9XSh5sSs8U9W9j3xk
VEQtFG7XT80c/aVODN/HXwW6blN6MWnJU9QkB+lmCeiUYBOnQhus9Csa1UXp
kTMV4sVKohJdDxP/71VUtMUS7gP5eMhDAkibI7I0tgHnJnFVFeSux2so2e/y
+bSlhbvjDfHyt3S6zhLYXfZkGHNHaT+dWPoGv4D8tYtr50xdRwOV8aZWcIr9
NrUyw3p5SId6Xz6D9oHN6fbCd1ffvl/FgBgTGeqs49/YPsm7hGmSXhXC51ai
fp3c87zuLob/AUqeNKMZTP4qxLkYS/LkIzkBhOa9mAM4uhjuU0ymcX0ba5sq
tqdVyXElfWsswlsIT1njFoUqqaeDcVBlHo2QQGdP8Loc5lqDUJQcZUW7jQQ4
Kn+qlIr8T7OZmau9HpbYnYPWcsRKYwx+oZlqULlqq5wfUnSxtOh/2kdptCG7
gZZtqiHe7su+XuQWAQc5oJ22j63OTaTLa1kWhq6W6yTb483npU29KNctRyPf
XiA9t/Qqu2GM+l9j6hSBx3afnTV2Ka60fWl3d95/r0CRUfYdwM42winolD4v
ueqYAMT/l3eQ+hmGO4ho8cS2ArNDPiAp9ITirNNyDG0+HahuSQ2wDrh46MMJ
kLGiG37UoI9/B3+JFYtNh5pDYtHKWhiJVgQO8ubLXm99/nVT4hHJ6N09ypHb
NFoJDW6GGI6Atf14g90YhpFYY92J/OHdgCRPaUauS0nT6URFTsARtjvm4gBe
vt8GT87OMRCX3O7dkb09t9pCJcpBQTrMXv06UZEZRSNK1pVrzPmbHlBMEj4v
PHnrcgRleopiT8EX2XiKywL+zF6RuAsLT7h8euM+QXCobWdXOAgLegWDIytY
tkbzBI3xaoYzi71/0ri0hz/1WTX9id1qnF6VAcTHY3PthUW/zhM6NLW+/c2A
UhigUYxYBVnD/KCo1bGqRRX5j+maRohf3ouJxIOxr23jqi4TKFPF2TYOZm3X
7kZHe6Y8xIrI5QwQ8epEWVWHGXkqAeu2b8hxhz/oN7GQZLlBuoVZNTsQ6+NI
DIFgQb5uYSxl1XF8WMrEFxB85xcLASzuytbRPw9Mg1phcwV7K/v2RsWt29cB
fp0FQdykJN877kRmU/bQqZxsq/1xYeGVqsjKYUtTMLaDwlQjA8gbaDUlgXvk
mKxUTKZjaXHN5z4zzLaTkalV48730FJgTPRIuzcwBmuf27kgTnWPynptgmwD
W6mebJOWfdq67RrwBizDO1Qm8Tjt0HPCSSXPI27EmoUb3mXXtCL5AjzKRJ84
XU8Nf7c7PYESpsvhxFiykzeMOPV6d+3KpJ0rQxf8kj8zh+FNEGSRt3+JD9qw
0H5c6x+2GEhKgqaJgHOZIgAkWffqR/DaZG6pax9Hpn9zQk4a9aQzF1Oz2XRN
sRGXtcSBT/Fdkjl3YLy7XRtBjIyTYKmcZAr0CL48a7lHxDcVz/RZeRhvcMVM
/3PYQB3i7V25+n8o2j8ltB0q7x1JiF6g/kF7iD3RFjELWvFNYItf958siEEa
ZpdTEeTdzoBF4XSqw8Cb1pazxKTHlmGaqKUOMDEm1Rs/s1Xz1J4F1IL5JNfP
ruunz0A/LQf9lVaug87d3VX7u7ik/+BPRRbSMOIqHvsPllsuKVd6s30O6WJj
Q1j9AQ3ENmCjEPmLiwg9wxX/mnUohu/evZyKD7QSK/cyQoGQewzDyqBILHEV
aN0gD+H8wlsmPoCtQp6TwtafwDG0RJ+gJqMjxi6J2x+fOaO6qtIkAFfu+qLr
wZF7zXfDOED9EzBPVHvxmV/FZ1oBj6fF5i7RGgylnwvxLvz4mCIpZt7QZUGf
6gTAv7UEdR3pZZ0WxPFW/aMn2pF+yxL8BdYPOr/1cPgzjZ6BDfm2gmiZI1w2
02Yw0+WuXdIJcPU3VDdZBgM2+5BcrjWXBC8fiDhfjthNVzZQGDIM4QIRDMdI
Vweyx8ceLGgqrz92GdJ1oi5NW9xReUZPZiKTX8TyST9CLM3UULyngGGjfn5B
xiw/amKc3i4QFSt06UM+2f+Cgw2z+slXUUwy1T4dQK2jyUOnremBC8GT+0az
158iiGeGV4qCwnXIT4KogZHtjy2429Sw9B6JLOSgH1Yon97RVOs9BvohZzoG
E9toHN+Linx6rBu/9kyJUIUYw/cWiny3/CWWfUffNf7A2ADTq+g1psjUUpKb
POJLK+LuNVP9Ycrq3xYCG1tYScoXyTAKogekTm9LmqegxRRT9+/DqwAqDwZ+
g8ZOSJLGeB9VG2TBFjLXKv10OHHFYjOWiJArtyySV8n9i+4AS8r8W3d1raop
N3Yojv/oytnTOy2MuVjfsvpbYyXA82sp1HSlHgBQiYmtJXbFutf4TUM/4luN
5cwzq4Sej1xv3REj4aVOKyihLk73XngI2f3vfGQV40UAYmju3UI7S2+iSWfV
IwSGSt/+Iv9rUTtoc+G8Tj2MrXAPEf5hJ44qhPl4xTKpCbae/00pm4xBKHwl
jCGjcQseg3oU+5rgzQI1DMLx1fdCN7vz5eeibwIDEDhpcfCclAMGQYbky22r
7hMvrpYlh7Jb57WCMY1rxT7MezJMLSnRxmMoi9KCTOX02+pR8A0erVfc9h9d
iAHu+yOrB1oUVLHiVbBxRKrLolQ0dDSUPIscsSgtKMJLEpQLjknuVn6+x/pI
duzV02d2Xg4iMwV++HBlHPdHscfsGYHfcslmEpXKrZCtMHYBL8OLXzOtx5t3
wJMNhEgvKzAobGL1/GMeQboZW2LlMU8hSVsby1CZkbG9yOV6EnLUZ4gA33br
r7qcpsFXwgeTbvrvZXr5fX6QFgQMtDbMrRRWazcdx8yyK0qkR39q+hHBD8Eg
2AsGx3LiyUqvwjTC4nOZf/a5NrQ+090kzGCiNJ8U5jpY5eRTViRqwwAhYMbk
9P/p5HmfGiKp5g2KUNz8uS2K4FJdb+u1emeYmaAB/tqhjtwekkCUv2IxumDC
KXGO9TcISDN46IW0ofcdpIM72HbRcTt7RENPWAXWLC3x+bhCoF0PxIX3l+QV
Kkk8/sjRTwCtSZNYhZkXUyR9E6EcWC9Q/2Ms5OylHAQbx9c4biQcLiuKGy27
EShyl3AbkmMP1SEU6u1gwp6ut+KLYa9BtCYwW6VPJ+tKFPh9taDx04smX0eq
mjLEQSvNgVjeG4Dk5Qt7a6JODgGX5B5J4PrGU1eoAQ4lR9aMImLUX8kWxqGH
r07V7M7TBXGzYmNnBOsjy+OJtVT2BaPCuaDPEoPqyvPobJi390MTBl0Piek+
bKItbCUSXOeBU1Gskjo/iLXGjwtubXQJ+f+GG/F9Ew9isPf5x3N3cuUiCz7K
lqJc/bkWSswV9fVojcXFOniutN1dZSokDGE3Ug9czZ0gGYBL4ZOWqOdNS5Zs
xf2rGc0p5gmdsSUBMFLC03zahrxuHrb4nF71TITdZGYFQGLpjCki6288Oflm
DsVjOnGUsPSoiTlGKOFsNU5eyyENhfgOQDTI9wjWRbkOYbDcgAZy4BMmTIqJ
1aCTLXhKbuRQSOizPumTR2qolBviQIQwf9b6Hax4eR/lHn3smEQ2LFCw++CX
BHrzh0PnnSQ3WbF91gFvfnA8f+4JOMS86gjO+NO2NuNZSza+PXtHfC96NNcR
6x1ICYs6oQxOSxwhOT3ifd8kDB3yo8GmLqjejSNeDZPa+/P+TE/QlDZpioFU
baGPXy4on4P4gmmGqd0j4GsZ4nT/mNVVGcbPV2/wXtrT7MQfrU6tqSvoouxi
AfvJVjcKHaTk/MKuSiBFiZJpmW5NM1ILSzabWK88/YJrCLNcNpdztu+U/x73
+aNMhOxSVzM/O5LHBxVSOWFUttGUUIWQxDg6Mj1PVd0XvnZo0t+WCbpOR2Px
3oWtofWnMYh51uZuuAwcxWowR4AOOQ88QLFQc8bDPJ/XqWa/riW2JjKbMSS4
nHqpSUJ9XfLhAvCxCcOhKfCoAQ3aAdbJwXdkYYfvCgwy8r01R9vdFWA7wTjk
+fF1pJVAW4QxGMtNvLxMy2Le0eP0q5nXcr006Cm0M0g+fTVSC0dJJmczUqc5
7N3uIbMLpNoYg5iHVGooO433dMKU1cV7kZ0t538UQys0FN00uK/vlYylSC5t
NrXonLWSngDP2M/fJ7e4Pte8XWXTCG1585kwr425yPKb1/dCO84sogyy+Dbh
Kaf1kvyhdEc7MtrXLZJAp9bj3RpLsMNN/lK3ebt06Tw8R6V+gI69veOJZiI6
E6xtrlUvPxQXFyJkT7qwq6wp0ESVNrDTueOv5MICnYv+lWgP7SlddI/B35O3
JeP7+5A+/2EOWWQpZvW3Z80Kq4kqFxFEr23XPI1qIEX8kCJSv4hKU2jqN3Bv
LZn5VKDNylJeN4piKSUHxnmDTj2hFZ3c6VPx0pjIR+BPhiDOEQElW4c/MabX
SAdJaoD5TQRaMg6fb1ux+TcAY1MjqUkB8zP0NFTdmOfod3BucuPUl8ZA8Qzz
lj1TE2Te0ZM1z7Dmi1kVsQpKUgNKImluwCUIFU0W7zrXUhO35CxkuaxrjcHs
MjqUKCjXX6yfgLE1tdy/liUkq2Tly10odJEgSZqNha3Fh3HSp7hS29yVyWSp
EZmtC8AX7cJxuH+SQEOdXkKmLj9A/wiTCdypG2i0gkuyZGHBT1QnO69O0DoF
CYpjS/VLzPcw5vefPdytvy0KQN+8xGjtDOPddqIS80hcKR2tlfjF4CAa8nsI
fmVl4ChZDNaYvLhMoVR4ol/niLb5ngC5wgznqV0UT/2ezAvRMO0Le7FpqxJg
mc1qAG5qosj3Hg1OefCkEfNfrymd38WvDiN70Lz6Otv1qp3xrIMl4Tmr0pqM
/7vsZ7xrD9LG6XAj/RWhzYGyeLFmv/bFo5PZxZWsdXYzCnMAMaBYJKQzxqnx
U277UBE2IsOCsSpEFl1+S44ZesBJJjyOGrpaI9mKHvM+d8MeyD7icSZtgn6v
33TDNocjAjz/Zv6G6FqjTi/4aR448Y5BdeSCzdzZcXHG6SQzI8KCz9aTSjvP
fhZUdXaItHTYi4maBdLnjvtKQzvmrANP2iNUWmeyKOrS00u6blB8oZ0XtGry
GT/5scPy/6nwaq9KKhV5/8LakxUFHFCX0QDYOejsFvHkaeQ7nppuUHSp+TCd
g5eNXUCKnjcBrZsgn0tyRXB2h6nw1ljeK6dNE7qfp6SeXZLh4q6JopGgMQEC
dM6eEf4WS783mwQk09RA141i2y34BHFQ2OFA0Ap0VB66DNT2NamSakjrrt/M
NjGFKisbvH/CUrum7gx876ODDvXHd8U4YOy5MptNlyqS13E8YlaPiYi1A2YI
Lj8T01qxYVR8+UDESlqqPdKUX8wEq28xlZ+LfqXNQgsfRtsf39xvC3QleUkz
Fs59edvP3ji6W3S4Q7TNpwAuCik1myNWs+mR2l5K+wpQX19SrhMksWhrz6CH
11puJjdgDyIs9dVlk7rbedniO3S43QHHsMuVFzs6eXAt4pTpmfVRhgEsSglT
+MeP873VDKlGkBUhYCXfz/LPXuA5o0p+wvGziOct1Q9hz/GopFw9RUmOtb5t
e28qAN0GYmO2ddZ8oU6EqvnIqYw8YDDnsYQd0K+YBqMAqdd8U4Q4nS4FFhER
Trd5WEGcOUlYWt6x1BOcLBMqjXDaggzmVwXbYSagSR6cHDJlE9Qtk28OUYgH
4fuIrbkSuzPjdA3mk7FUoFu6sZI/4uZk+uLdZVYeWSLx7rvi0/ZrIcfHK3rg
znsxqI4vsXaRlTfrT/sp9uB6ZmzCsEtcmBb74EVxSWb26ms1RJut0tC5ynQa
Z+77hS6+7IXBUmZaSFbUBZsz8nSEh+e9TdhjHOwyvE/wDSK3WVgrZKCzIc2r
Z64NgZ+iuzfEjPS73QuXxrMSskH9w8e5OqCbOIezVD6QCe88omnEhNjQwEGe
oX5F61/p6f1/BJ0msz8DvU7V2X6Z+JTIAdpd+QWyRmoluYFEgIQOuVA8E6Td
MSBo1TAjtPqD73tFZBuNy7pESw0u7r60NBjTVuSp+ZO4uMGNUeuRHszcTkKY
mSUp5ogHIGiC7oHSzh25NLO4VRrnvJHc4dHBJSNfCfzwpcqYFqwVCo1aFUc0
p9jDLthUeAqf3dgO4sn1fuuSS/zwbqZ1Bp456y+fm9Kg90qxIxrEYeO3Zq9/
t0+sB1SWAwyquZN9qiuTCsLdmbhJ3CqZ255vnPA4K9358WRplCtq1cUUyZnT
5fOQSTKp7oKc1bTG/oDCSWfHyxpatcbIi0THDtbeDQiCA7UYvT2ZJYmUqZEL
2y96uFx+9UctMAYvG03dj79aue7I+2X1nJ1JYZu9h/rtPQ9H396SZCuFrbcB
ipWON/nqEJhhnBv3lDrm5LH5JMuHTE666QtxVcoRHhhfXoIDySLRqfc8Bjfb
6Prh93zPhdvHrfsB2YUXNuIC5Yv7hAj1lhOtBSn4AZIV4BIcA5o//TIXeFQ1
XKIKcozV9mnbloBTuIAwzmjGP4k78ie1yh3TDHfmideNXCn08qxwV80jOAQM
SHloN3D5XhU+/QRqap+c89PKAECUNIsLWq6DgiOpUEokbxHGChps6BHmcRUj
QzRJ9a3jzsVJAMZs2LY7V09DFu8EYKrcA9W+I9Btox/YWVKkh7hA75neDRNT
PCt8CBbeBlGbi24z6YzgSUcvvysHR7FWbAM/jXEsZxtyz6S6zUshbcvstHxq
IpV/U8ekwhc0FX7NavPoltvxHC7PGzpGaMR7KOrnuVTEAvNlLWI9DR/X8faT
DgB8pcGi/G273gBCP4WeLC7rphs68B4IFCvCn98pdvFiCmK2TMIyy99NVYqZ
zhRyn47ewD200iEHa+C2DOkPfgBRGvtc83zJGpZoUJZMe7nnJ6uogdFAb4KH
I22xThJXpIK3DmA/OvkvmtC/+oRN/DVyBbg/tZcnyPyS69LaBU5HQ12T9JKZ
sukLmfkyBgQ9hYPsOXByGP6GDzl0YuJIjVODP5vtpauh0NZmSSPtg9LHEyM5
9Xw+B7hHOI3P5Wqu5CtfMd5NeyF+CfO+Y2DoVcfkPg0AZuLKFQf3G6OqvOMJ
4TC7E83xDsVuQbdT6NH5XnIVXtj3U78eSFXyFkuHUptCtyhUBYnUSOFI8C53
DY6avKYp21u2+evyN8ZtDGe/0uwv3xpbIEfA851MBJnV3LGnc82z31TbJvnf
Vp6xU5tC77V2o8qt1qBkjfjeX4iPaxQzuX3xO3R98lFmAUkQ4ixRyxdu0IZy
DwZc0oNSUWhN965y+05f3XBsPGMfe/EInXpMsWbUiB7ecSvCI0ZPXygsojLg
tL7BLD+IUWHExoQcUtEySyYhgIkD/w3f/GlPBTWHWr2CNB+K3qmVzBD/7pHs
rwMCYkpR0NGmPPSfJV7vRNdoX+xcEGiHmCWNEcdoQIl8KY4YSa5hmRckaKRB
CE+Yr+RYRaamCvQYlwKBD0B4XGVaDARNvsrHyE5ubfS8iHp6My5HnBo3zqQK
jfFa7qj35Olq7O9SWCHppleypGMk6mNZ5/WWuSNS8pSMvHQ3DhgOapLQdOTR
XFiadusph2uMjzVqDH/KJBgSlqcMkstwa+Svz3qgEZa8xOfeata10oa2Zfsp
2RMCUWq0SpAagPOhiZ/P5MXnTirZswCmfsQRhCZKaqIqVa+iDZNDbqnjKx4T
ZipJlebxYAy8WjuTafZeEZtYC4+3WJQ48GpaUrS6TL5GQ3irWnuUX13oMzyg
D3KeNJahlJF6RWousjKqjaIG4BVOwA7ZjrNhAtjXxU6FVZaGVhNk2vdadMvW
UhWTOxyZXQ0FPzfTFndmn6ADxl2tfJ0r/5FX17o7vkhQ/tlgBtLmGABWwNYL
D+MRIra0Q7cWHVk9Snp6X9co88ejS23Tj6LG34tqkylE7TsYwJkxUNhKtebX
4FRbe+pDb8qQmVLyrnxq4GqDEDYGZGBROmxEsY+8yE73BM0rxVHrax1njoEY
J+NgpJxp8d+Wifva31EzrzMiRMyOEK04u47NddCSKHgjiCitifhGDAfwLQ50
ztLWlEetZWQd8+Al9vCyFMQOmNStGNKwQQ8eUMVQSgvkBLMsOn0jyXgUIzix
qDXaez8PY9yLsK69kKv13Y3PKb5Dt6FVDdy6CKfloTwWYNBqkVWgAASg0jZR
ApaM4PfQbeKfCdR7jLSEI0MBHGpDhdxLvo2M3qlmRdG5S9sQj4KtIZBOCbVa
M2S4mqFF5v+iH6mZAu08aED1zVFmgmnvfwkJ19d9B+rPiKp+pawrKK94msRG
iyaiMIOMUCctWtIjY8SJDhu5q1SQakT/Adq+rof7lOJQl2I3eGGiJHDoidGL
MShfwWOjKMXHxl/s+wz2kwRHun9vUjrddsmE0L70yYAsNB9jdDmUnlsNroJz
OCP5Xl5lel08qjHoqKN88GRpDR51pnphvKwZW9ZwhoztdvyUug2TCJCjW/vD
WMbZfMKjgeoiVajr/Yg1KZn6sVFTs+hV0jsyZdBvOFrWxYxgkuQ1xAY4+kDg
H2oMwwJKrkGKVnN4THoPF26cPS9ETJ8tBcnb0qo2Bfcx5gBj6JCGTRcGNqfT
fwWTzdQgZC3CQ87blH8qjVLjQqrnHYCyP9lZYCAP+6TTtN2ZVA3Y4z2W+m/0
IGnoq/QXjX3Q2fiuNTiTMS6VAWgsAo017fNAdppZk9b4XjzTwi2JPnqsn3r9
NQgR0Bxvb9GvS8lNwX3BBwNbAPtcURZ/7aQRBKxy4xgBXVNY9RNzTCUG+A3j
kD+e+uAFdrKhl0PHZ1UgCAv/OsnAMIbBdfpGge02y/GnizKzQfsTnKaU9hq5
qQIKWe4S+/JiQ+Pyx7Apw75a94Za622qmvqK8T8qCbDLYbKHh49IO+hbeoHF
ApcQifuVLH+eYfjUl6PmcsvMJo51T2o5gwAdz9FEwyvSrA0/ijFcujOU2nA2
JwnlAJhFiF6YMIlvLHvIAfoUPbb/1yOfBygjRrpkQwjpe2y0DCMgsGew9Y3Z
hRLQoTQkmyzl8fZ0AB3u1npDteg81WKzfFFomyTl24auoTqqAPFfJ7ZnKlFj
ZfrMoAy1E4IgDaPCYxq71L0YPvyEUWqZieB4BbNRNfQmeCEElDYjWWSByyQi
NIGIz9QyX0q0H0FDhvK99ri/r+4c1aCD4BA/fAH9lgGGYV0AlAcfo2Hbs1mL
qgCHYM9bsvbWczFlxT6pFWdiUz8tKpp3N9CySiLvOzQCRWY9pr0ka9mRL5wI
2hRTfkVbTBe30oX0N7fjnkzJI1shVrUILm4ZySr5v8Hr3UcK/MkRkCWfzsXB
ddObEIMDb3fIIgBwGPcC8GZGyATf5Ydvazbg0Zo+GEUvohYhJCv/rDNPsv/8
2ush0ASk7D8eZLD3VsVugvvfSwsknUIddLqo9q1a9VKXhu+sETlQxGn5eflb
BOiVtdDoSFeK/XqZqT051BkYKWFrCRGAZrLXglceEuk5pzJIGXddhRdBa8JK
bl1JBTcZQmPsT4NiKGl5sFAPwisrmr9YE2fC1ox917LGEuzrsCRwqDhKqCzF
A+7vF/9oCtyM9zoWgsvXblrcUeafjHumnLkSn7x+HQVcV+p3VyBB30BnHoVX
5TckBSJcchSs2maByGB7gwcT1EUvtcf7Z1+YxzAPvXau2dSs4JKIwJgJ2lv8
T81COfuUxerbcwcsK0PpATvJJokLrLM/UbAiu0GolE5MIRaXKED7OOgeMuQU
YeEjhvhlnfNmD92+VluRClbnyZvHLN4WTyV0O9D0qF1xXUVAXusp1q3MhlVX
aKD02LNLRNcSWpWWkR5aavfztgnzQb/6ncYna+X9i4tUZ+NZy6QB0oxh/uLo
fH1esDY4LafE9LaVqWOU/M4YitjVkZ57Eqkx665umWNh92ndnD0xe/sr2Mtm
ZuCMwnrJXUWfWGBfabA1kmip8R88VbFkozkZpmMVavhdUFzChrfhlQ+vlxBk
/Jif6JBACs1md3Q1yE4aQdr9/Uw30xWD8M5im5hfjsdzY3ScxX1CblXkl6Br
b/sExMeqvda35NNo4aDxQNf/WV3TsdtxommyDW7vLY1vzoTdovuKQjDAaoXG
AH336nISNU/baejxR6wXnMAUyP8WpgtlByYE2vED0Ota9XsOqpnmRFLwjYiE
+1zlc/LikKKZaVdvCIAdzgXCFBfZvkKcgdNnoJ3sTwDOrTi/wYq74MoSP/KY
0oGg6N8FfZCnkfiw2KYq5/fzYtURUuiaoDfobIm/db7Wp3cmqtA3Hx09jAUp
aCw36cp30DptQdLgnUkESpKZMu2B4wOgo6v9zt8CDE3HilFpCpcumtVgiyqq
aps7JT++Qo353UtznjtsPhq7U3UBTIpIyJBcCwZ0pZuGlgO8tpUGi0JZPt0w
kCJw5+p1jB7b6OiAA87lnSVbGtoB/34Lp8/yJxGHfECxtFWCUl8uKkKg6Ly1
HgRUOWz49r2vClb1zynIZms9B2HsUxGMX1/wO+qIFQl9MBtHa4I9/G2Ebl3Z
H89sGc57x94dqNFbU5CAPKn/U2V7NRaitVLMxgzo8nvv+r9sP+OG1yqbX1u8
OnA77PKsglM1AcH90TGNqaMH0uSvsmYo0BS/cXEtYOCYtLTnGSj2JUl0OYmj
GVxD2diwt6oKGNyJ6Kf2TlF+LMFKIrnBCBapbt59L+/t5uMKfjNxsPUemekg
MVYeQaltX78NugLh6P9DPfxzUqPBIsyROk1qapXWzSQ67zXEdhpLrmG0MWTR
Uxz+Gs0BwY+I1u27wHSa/8vdUR/OP3oH/pLPRHzrB5DYNrhTY9VoXW/EWvaV
Hf+uLHAzFqapMq0o80NS0J4pNh00QL0CJZPT/ShbpkqnQb2jYOnc1RFxH8VK
GPQ79i4L92RojJX8cj4i02uUBXCJU6TK5Tcb0XepBrdd+F+p1n2OwyoVn6qM
XcGpBG1JI+DCUOxLUXPqwGhmAELOVOl/9bq8IwpjZBnLjoutzqmLo3jSO/yI
UBkiAlHVZUteALshEV24mkdLZNhlzp4Mc0cKWCeFusjKhNHxtuMRZ2xObtP2
jLToVgpONdyUvx5LSsnHXa0aFL7KgJnfHUUKoDY+BzdTcKgkyMj9Cfhj1qVR
cyNvVoDIqwdiEx9Y0r+It3fLR+TQmtQbKQ6Bk7LzesD6lpP5Z97UfCwB1M+S
ta2lNjs14Nml0QDrMyH3ht8ZC4MOFEK3C7CgFbvywcdyXl87yS0lyOuBldQl
w39GMqZ2Cdn7EypQtQJSAQr4YR331oX5BVkGh+FISKbSWD9dK3OaAiveT022
KzA+2NoIWKrGNkW5Uw7ZRZ+kdEPU8vEutc/nsZ78O/CO6FiclgqKpIo9kNvY
hEfJuSWosypQN8JrFmwOSwBnOpZNt3aMr3fMJ3JAkldjxkc7sFWk3z/3kiUX
Rzi+iYmeLHNsJCznLnIxTpDuHhGweldNYjOMHlq1hIrdz+3yUsYyRXUL8Dgt
HSU1f0ZD724Y2GE5AmibepM5BHzEqfZC3yYil4JeYc2Q8OBhH3C14cdF5txk
3/APy4f71Fy+sdlLOGFtjkOVFxiUULhTJvSbEVGrDqOi6nWc06wEgJKHl1HS
7xIiSufrcZWBO1m5USMS5aD6dxnkgsjsCAA+B+s6rl2w0vxomVojZyIVj9Ya
4D+ud90D2f7S9RRFoC1CJPh97KYZNPcNSMMGlh+Hb9zvHa3ohJElyjItKPzY
eMCDLMnxKZ9nWfVSuvV3JiVsDll030TgUCjvq9Lu8974GL0jVdEMdu/F6bjr
0PnN7oeYlJRhEkOszyyv2jXkGDk2XAEUtFHRD6VBsbCrunn85BwHuJnwGIE1
pSYkUnJW7qf5BeTOjyE+3Jgg6l4DQLR9jKv9gGwaIUXIgv99W9ysaPkMkEsJ
4AtU4eTxCYPjZZqSa0qIakMuvQMUrBWnfPXjiIMadnlxCLCy9B/zRb6ndmnd
knUOfMVSAvOAR8NtQtDwTuuE6AB5ZzCSVJWVMj5OmJx/dVjVc4i5wu8R4ywv
eksOjcqiMA/Ex4nqrwHntxxByUvFweQjtqlG1wxg3mHWGOQe3aEnzRuhvHtz
qU62N2+eLnJ8kCR006xIKqfsM7DQUD8YY76fadPm+hun1RXDtJlEGQdeFqTZ
9qZqS5cvkpR6fjfbqsTTzZzxJ/SfdnWl2B2x+i51XqFdlxScQvPYaiMNKch2
mFJ1i3xKW+y5DyNBOfhWg6oV0S0w9Kh40/FIDTwvZhmBt9xlOQHSCtvJM1u2
PBo5YNrKODYp3MaUWbLVsbXRFMN6IrIZokbuL/950iar7KnjB0o3mLYITbMi
mIyNPB6Nx0J9XuC0oT4feL/toTw1OOz7w6MBHEhmWk/5Q7Y0FlcpLhAzdYuv
Az+ameg+D+yJlj6YW5U5bGau2SYRnda7/z5wKjVT0oQ1oHQ0I1A1N5e0WBb/
iiVscs89kSgMKxyujOdVdQSryUSaAWqpHnMRBqS5ZKUx3zAEKMqQR0bQLiic
FNHMgaPEUWtvdSqcnpejxPdlaAJWRPjCIjf0mO1OF9lWqf4bC6ZOJLzkgBrN
/c5SS0axcJGrM2wxjgaWg2xZUMwGfMK0F49jrjsZuQDYq0nHUZs399z+nQof
IeuS6f7Wqciypxb4+JmjRejQRcKPNUshUS28EpgM3+YIu77CDCvNICzL4Ipb
W83czR49uMwb1dheRl4ibgPW+6Pto0ngBLjWyi4llObWST+7MXSXbkuivGdg
qc4ZO25s7vomrmypJEM42nFBze9obQeOsdA/gNc2CV9FDFr93RlIAcVVzKr2
c77mSFpjfPWkf9dh9JGUn+7Jsuse6Q7P5bZoJgTIsjJ2tWUbi1+jm/iJERiA
hbqONS95SHkNsJrcKQSC7a+8e0eIY4idhUTTyHETqnyRn/CWVO/jJFeuqR4R
0uvIoXfZrR1lHGFExFiWhAsQiZ0XgC4koTn8Tj2BRcgCLKTTLbjtcm2CF5z4
gexHp/rGzp2Xiq7TDmjJouDQOkSZsE7tGxP5jf1RYNlwW1e2WIH6ltnfv5lP
hKj4OpnD73KxkctE6/4Yrw/wDbJ2o1fxeP6pTB1NxnlQK68vlvyBj5RSRYeF
vx2GmTR/Th36Yldm8qtjFAi/emcQKkVVDG/xY0AmQNYmi1giVeZf4V5tUDpH
yl8fYPBLmy3K/kb4xFMB0SpAu+SZ6YBfKgTBOn7yVHGO1SjonZgZRgBgSGKQ
Alk8/hnCqJOSDbFiunxG+kZVBMdecW+twhf748VJ2J8TRuuUA0T6M9WzhgfZ
hsdTezvj9EdWAdLrXGYnzUKDzGXaAEiQBlyEGja75QoIpCQn4VBfJEokuYVn
/pi/LM95Eobtmq53/ZR2puamnD/HKbnZB/gTExc2x4Oa6RU8w9BfznSyQXwr
IT/f8kVtM7ad25xdRMPIaPfMrPYDxnFCvNzi7/6bCnHHoQuLNHabCy+p2dD0
zkCke8zQ1SX7e1FKkLxz79LxcWdmFsuqdWOOQ6T56wZ3+5/QNL0GW3P1/VjB
5osg5CZK1kpHN7UbGBeEfra0RKws3bRa7BdBuBxHWgR7a/BSvv1Vr2G+SpXp
p+4W76RpGT5R95Z6XxobEoHpAMNG+GaHXN/8MmsufZnQy/qWyBoGjBAFbpJK
H6WWDAqtzPB0iG8NfIzhRzfO+95fWRf6fnNU3ZHe7qLxjOvKPjoTZQJzTl/n
RA7Mducz5QZaYjL7m8xcDg4XN1T7Sy1Wf3pWLQAA/wT0j6TVIqjKvSDG0rO5
h3mXsEeAomrHFTsNZwrIvafhBSaiPQYaoyNPZ9FcBRLN+gdl6H971gCt+WnC
ltQVlzwCIW6iXFd/XsxOKpft5eaImATUEEA2liIfqqthTSg8wt64ShdloXQK
eSZRQnIXU8Hc2GBECKvhupLJ7Y5/9ln2p77Wrz7qLIGh5T0pjJEGRXRlASA6
Xa17NSWhMr9O/FMTNm7/8Vs7Ytfsk7jNJTWpG9MaiKrZcf4OGC0UpQGYLmFQ
lXTUO6QEWAO2v3/eAAtKeK55d8mBVoITlvBZRwfehOEnjOMAu2IpuiAN5Yuf
JpbYecVHj+NmRDSA/PY2fMohXTi+5/BRLlemSrSqyL1aE3quSSbmqQVb/b4V
EDa00eKNZ30xsCtCbTjvdabwA+yUNj8eR4SI7Q0SHAOBKr2GZi6FAWiVUAOo
fB5oi7FZN6LUWMJmEKtqg2E11X4ocjN3b0xLm/cAMRvc6MHr9tnsCgbWHNoy
Hk8RYvQ04Xr9GroOPhPNyDpTfwhgXNMaaCyjE9ut8n51bfyUy0gQw4MWvaxC
rwRvW2XWRnFeEs98+5wv3CJWFeVrL9d5MBvz5IJV2BflVPjUmbIMB5zeE97Y
yzvcGgOyIob8WNzRvtTOLaSK4bu4mhnwHtAuvnWqlOnm+nqhLEtX/wssGjvz
KsBRWWfmm+NiANLXVPW/4w2auPMjU0NnZFbnVv5Nq+LhluHhymJPIOFrTHhb
FhmghUPiYkkBZtS1Nuy/dyZzYoj8bjaTWli4IOj7RhmWNeK8YAXR4RaU8FlD
7bHErby9viErZa28WRdpiWT19unIjdCYtBPQqcvt1NEGzqcIwKiQpAR8LZ6Q
qvMz1yckBKyl/cObK4Al9FOjj7aa8cQKdGC3tLG2iBPHFquiXFs+PjB0iqQ5
iWe9c+6Gzf4We+phIriq7HKqHoaPOo/ixi31iIdWSxTEI/crJzW7Bq6jN2PM
aAdoh8GhbQKp4qx23w7qdMt9F7xilG9G0KG7BG/sRyMua/hUUGBNLhFNcozv
lMQkmbgvQjh2R1u5+0Mr19XEjoFM3mBwaOTw0WlAzWjA+6lcrim/9hl9U+2O
Q7O5QwnlFwBreonRHScbr6eT7HlI3znsNA+Bt3AavDSo+k45J0EShhNpYZkt
J5iJ1/JYg2owXc67BSDD8SaUME3FFJSFx2I6NMuiM3vU0K8sTHavHW53lVr+
1UdTmSXUOPOroKXCjB9RuCiK1uepWttJH8Fd0T6IPi41h9Fa2xX9u7Y0dMuu
2537p8hc6VIuZqUxWNfLkeldwum15s53TTmO6CoWnm3ybJfZ2pzxpSwnvLwo
Jo25C48fUeb4GTMRq/0Wpb7JvJrfJqpB2tlaT24mc/KhKxrVnivxiTC2WnAx
E6+blCCgy3S1r+N5r8DO3p7Sr500pCzaNaS0P6KtuM5hxzUnUKUvKWV/+OoN
OA7GbQWkMyF9wUzFh4OYBFXevBJFTbbm24w6QbPBrZv7ZPjdhtO5Zv8v/lP0
KXxgHiHPIcwOaO1fua3O8SkBcovn5iOeL3xSfL/9XhC0eLHacmciLOCBIB+T
h0kam9vAQAm0+5Fku2yFvEMuKMbDPII0mfEabuKISxC1POjvhDc6f6OFutg1
c+ZdkyLeWF/Gdy2rjr4BSnBQj0EU1Z6YvCCcmyB+OvQbRgIdHPHAc1Yy0yzh
xrjyC4k4kgBWALZhsdoZ4iRoSP4MC1UJPHR+5CBLvgPAYMJ/SwM1n05CwAjN
mKla0XaY6gsahkFUJ7ceYTvgrzDpEfySDHZXL1Ok8PCwVZ/BrzE/B0j/aA8o
iHCcZZP8M7R9bI2XrIO28wq8r9ZnR3/029nmhI+F96KruOWL06vMIYsyyzmg
kcwV0JWMeNYUBux701zF2UH46XJCnJX4hO1eQdVPXuvn6GbsPLK6JnmvF9/F
MxGbepoIZrgK6W28NhlyTUdCFm9aH9Q81NOWRjI4xabqMqbJS86dThA2uYpd
aSv7n0fWs9OwyehIXuwf5zaeoUWbIVeDh22eoUqceo7MX7e+zesHuPoN5wuq
4GcAr+1Gl8V0TzvtUxsZ3jy/bVUlceMTayTAF+VtN1mqKa1nFBLxEn4vixcc
N5bMfvgKLMM7C5VWAz/7zU+EtEGgiXix5doLEI+PxHw4//tMlu/pCeXEoRek
vMQpbwOJZOMPZ97b9EfzgwSMrSPb8uqnHuMUjKLsAa3GIdcHyn2t566asHC2
ntZIds8oGKGae9EepAGNZyDz22KQX9Aq9lqgjshXPJ66TxJNuN4ixLMZCYDe
3eGHYeVdGBroZGfmgevMXWHuWWEWIiFolTcbreNmGPidWbsJeNI5WO0rZGJD
WqcyU0yXhDzY+kx5ELTuCt579y142StDFF29E1QlP66OrFJCkGRbUt+wc3WO
3oZ73ChSds7Dt/yu0JZ1C1Hz4qIujDjNpXUEH/wsexgq53xrUEMfIpJDmJVO
vA107Hp9YWsBkKUP8R6hQhiiJOycS0FGD4d7yNbT5sc3cl3ogdQqcwfWxQye
gMc4QnrnXEYdXFLtRnplZ9A0QpsrENoUYiaXR7hOp9ZmWYz34hEBeBBaKgLw
jZcXItHiW0QAfwXLpWUMwGBbsGuKCxMzt9cA8bTVkscCvcVX67KY5sa6KDAP
qjI713N3psIMmUxQt5tJ6geu0ArSLpOHFjc02T7DOm53Khntx84kTQJuUrLc
xBUx2vkDVPzmwXA+UesY/pN76CooKWZxZ8xWuSo7Vl/FmEoV63ql4sYFBl3b
Xl8hDvYnAGGc7CbRFNZEgTyMbh5g4twqQLeFZUM6YJBY4+gndnaFBuWLxpi8
cCl59CBDk8armEDT4nC8BDYII+beITV9GJfHgK1b+dNQw22egLcMtipZyt8o
//coL3gx4a4kFkn4kLYKOAQ6hZdL7RNC2CAHxGGufLb8Z8Bw7HeeR6M0O3kC
uTuVAIPE/E45+K86z3rpc5Ie5eXtmsASH79dulvGjIegaF8RMXXDuuXyFe+x
WfKDLvsGsiczJtKln10bhtXXrqnx4ZNNOcck1CNIf6qYnGZYQ5/+7zqUOiXQ
vNPyGsDGOlTvtbNcJqGsUmZ/8pnt1eWSMK3Vi+/EHGOhDSKto58WAiJOw6Jf
/NvntgtBG4xWxURyiFvVdG9V9tpZHJv5KvbJ1EqfE3+fTDOHAieWSmZcExzl
Gkt2rHoymm/MhlCZPaol4qOK0jc4HmhXIGYzHnlLAoEJyMqAL4zAAsmR5EAS
8vGDIajxm8SHW3O7bzQc0kWufdzMZzarJPiV6igtDylja2c8W6tFUwlQBhxP
8dYKrobqbqfPB/lv0DMzqeVBquO9cvz/BO+O2huvreF/GTZ5eOanxN6myVB6
GC007YuVn/IQm55yHmmdSbguPqmoeA2JoNMMgtWH9m6phOCXyXjvcGquj/vQ
BnG/30BoPM6R8CTOYfxPAeqFm18IyVrD2PKwUyF9y54gas38LGpRh9ZPakvv
JBu/ZyEDGl7bupG3lpHG0JBdvaHorZXNkCAiHFJQL8drEIDZGw7KwLPxx8dv
1G2XYNUztDpfs9g/dBuRViNHBYaxDvN2R2HEZr74+Rw8L6p1GRQNaRTokoov
Jl8ewtsJDMBKPlI9CY0YKFGFVzvo+itFpmm2VACoKbA0kiCJJCwLoU+5fFCP
4ulnZs0uzFaCbIwRboYb2Lr2rs3qR5ebuMBdvrW/mb0TxbO4GXNQxjz3PoXF
uDM6LzwVEnJQ84svvDVw1U9hULmshYCwoWZBoUEOaHdblgaIdQO2CsB2Th1b
f0MP3ZdNYVAlAAJ0Pm/8J0c2UjT0otf6EVWfnynzU1eDmekyPHKSPczmAGiT
Vh126Iwtm6PjHGS88DKU01j/VgelYNwElMEKxqraRKoIa1KSugFoL8cUuG1G
/JpJWCUF0KtUcDEB54Mueay4KIY4BXyUAcCgzH6UJCRroiCmGst3Y9tS0OSv
yxZ/ati481MRJD7vG+qawMW2ReLD2agBIqMsFyW8TaBA1ASaFUvz8KH2uIhU
gF0thn3B1ulpcVPQNClC7Hs6jE4sOb/SVSsYukjTuPZg6VtxkFdlapgAcxqM
inKG1hrJ4TxEwC9v2QapuZHJGSyNrxzWy0Evkg1AkBT25yCQXByMCmhMN02s
QBmfu6oLZM4KcuIAKkZ6QVh0JTAjh0Zqz/13bhIW0e5APx7M7I8Jtrqb3MUm
2wySWIQOcnsFsdwaGmDBLm5Eh80ewFHuzCQyOid/ARzENGbyMfdpjnd5icrl
751k3IbZxQzlwdjcaScTa1z/2MID//RGiZaKhnDrSnRqZiJZdDIz9amwd3XS
QGdNOFN5c5KpjEzNoPePP1Zjkv9pPGel1tSJKlxiJAygMoaUhYtlECMyhsNs
KK79alAW/24DL6+MN2hYJHHOWM53OuFGQC8UUZupsMXFzcjEBTrduJdjmrmu
uNhwTI/MUaZFWf9GLdWBwcjWYhd0mCxya2Z2J6xY0ieySxA4w4acHxR7we2H
5R5IX14/QUD6xB273+4hnWSEmASk/buGWzA0Ll8lWmvPetEqVTQccfvih31F
o+pNLaXHh4cb6E4X6F8TSTUbWOrZco14DHILukLLJ/Lj6lHi9BleIaiVfpoM
hL9eCRqIT4XtJiL7X+Q9zpZNeGuUm5S5SmHgYuMLpN91QXb4qJkpwnZnQUfC
siz4+rCC50gRBIo9tJoeivzm6qsqxtSXoTrHkqBPspWaCoPAiObHG2+wd6vQ
jVL8C+E074f1NmH5XJA94RkcYnjDBmHjR7CwnwlIM9DxU9pqF61jjqGkn1cd
5z9y/T4WJlrJ0Uq5M+eEUkh6fALM5ZYPBbbGO9/Af8LOkq+DNGLTyXMIoZu0
LhA0OK7+iwJPOtjEmrvLvqa9wMc0FxyI7NbJyHcd3VcHZgK3AEfavzo4i6Lf
RGEp9W1XLXchpt+8/xIc7Nq91h+yJdrbWNobckIamMN2VY1R5eXcve5hpRdk
rnJDgzdtOY5bKpe0pgISRxpNiGbg33aMYiDlrI5mvDniQ5SqvMUUyLnfGmbV
YgJmOnE/0vRAlBnHcwP7OMgjJ/CR+6tUqAyJ2EayC4lN3Yoko7G25luC3Wtd
DMjwNLz/ijMhFID204mzwF+tyuSE3w1biCXp/r5R3o2iUfw6yVYN7k9Wfx+8
NHgglH8fnC31itspSEUD/nA+vW3ykZSuGgQ7x3KO2UfC/KSLo/ybdj3xGslT
RBGoJod8PMXhs+Avz9zKF573KOOFkOyXxcLxi9MPrBkT72NgkzShbvC7G54E
t7ucjpvVWo9BvQMxaKMzMkDd7cL12UBBXoxxZT2nkqg+bzOIuDPulov2Nw+z
11gYrnlJtaF1orRYdCgH2IQeIJ9f9ZHs4lypfcaDb5QRqT09uN7tfbp1hz+0
AUfzcyVoeFjRvx3vGeC+gixLvIMZFAc9xFH7aE8Yt8JzMJ1tuL5bHDLhCZik
60y7aTJRvPuufQRwodmkCgwauxntCi2mbfSuTGwGIOpztltERf+v40fZbyNc
YQrWCnXLiV12syHRW1bngFg1xljEb7fLAuc7sH3E7SEkcVZHrmzoeE1FY5Rv
hEZoaFmCyRipwi3NgtmoKhzGNCd5OlFl5l5x5glHiuihnrhYNQY6AIKlkqGv
Y3hAufwgT+NwPP03C2ZlqNE45U4AE88zvANOAhqTMnjocrISDBdY6KOM2iJ/
qTWBuse9QlWQ2Ar8Se5AqJ+vLUjrM9CSMH8ISQ1egs8oBuzJhiR50P23rh4j
nIRvbYqpHly2qBKh5+tgVCdt2WNWQptmVvLOG4ltntBmAWP6+eVImb0vAlym
X/kaOz5z4ntohF8mLM4yhaMQnso9ZkGNO+XN/0poNI+9sSMvPyM6Pz2vwP3N
z2HfB88e+XFA9OAIX8TypTXxfxo5Wjp4qYtDCvxEzW3/Kx13hoLhbdNlpVHL
zu5bEzKX8zbX617QQQ7xchKAmqh/Lf1umhwQmxrxh1J6eT9GcCsr5THJE4LC
aYMta95sVqN1TD8wnJ8SY9ghTjYGEre/v0o8UEWs4W4nTn3uf+t5YIKD0qJY
w7oDuvcEURgzbfaQ4EUkySczMhQbq0ro7KFXnQ8lNAoIn/6XWoldr5x8SCvm
Mt/3zQc1feeliXojs3Q7Fi/QyoVhm3agxxO61Nx6ek9h04xMv/NvfBEurxIs
e1twL2TaVuhDmpn4XfcGv/CU0S9/AJuIA2xnPE5fPoymZnRcXRp9VLioj53/
uMXX+wDSGQhy+HlCni/MNeEexYFH4OykV7eJoQaKpWMB+8p/O11K2QkJYZWH
jWuClVCEw0dLAMuXEApAQJHqibQeevZBp1BibVrACqt1GPPyc6VkS9sJeKYg
HdvaGQUlYJyr+7JfqvuFWgbGbuI8nOC1hh7TNwE3552w0VsD8cbFtuypLZU0
W3f5Yq9otXmxl0NcrfNb/6MnDaSQnHRD7nT7bQLa/1cWfI84hBgqRraABU6t
b0fo98nbB6eyec4A8PB6kGg+8+V2FE9sA6R7CM9mQG3a5fa3dbiy6gMZbST3
CM/F4a9UdjFgklv6xPflI28oe/Ojohotu3q3+9QaAdTHSmIx0cECgUZiKkAB
CdoTziSWZ2Tgg+IfkTwkNt+cJB9cxZlCjTK1GPdElQObG7pc0CGXQLiJyQCI
bVXKEq8MbHApQYzVBEt1ufCYKPGCWMbvRz4g5ZjFkw6bzGVFKM7+hC9yuHqi
FcaUQh7T08U2CWyGycbwn9B2a6cNW55koJaXdKQOTRQu535Z43on1lQrDh3w
WM6D77UqqNsTNGq1p9oGiWG4KluV5FpSjkt22IvbMKGGRcrro7gdy40V4xTc
L+v7Rznc6u7Yu4XsMPHqxA78qMZjD3r5ChNgJG7wYUQxqneHsnaPPzhFVlFE
qpbDQ1f/lcfi1r7pKxqkkJdW5US78+R+PrjUBxNKMRuuKq5MUiUdfbRnJgB/
vz7ywpkhsnfaK9hTQouQqIZCRs71I4jOjreEB+avC25fTDMzlADzoyxxsC1m
VwlFoYF7raXyMz2dJxBneF3I7YG2e617wrwLv1X+efy7PwYCuPCjANuwvi7w
4luflu51Xt0VokNjIYaKIjQgMmYbcb3S2NarXhArZJGUG8UJWv45hOluRr3h
8cLSh4MhcYXk+APHbVnFY0cywcXelLotLxGEZWNO75joMl0dV1ycG1Becj08
/8ljAAeMhmp681Nva35WmPdEkzuv0KeotFTf77mBOLykntNpKHb4iFtF28zp
OzJbiv77ADrLWs4vrOiAvcrTd2wXcwvYvRnWjWUN7QGbehuZTnHJZobvL3Hj
aEDs21PcEjyl9N/t1QrmLRFVdrWDNkvRGA9Hb6RiCvgwDgJ6TTg6txl2ve0R
Wtr3ylSN9i7UMvGUOm8ZVrH7SCqVryV5p4G+q3QObSAfj2EImNSqI3x+qtwz
5Ar4tOnQkGywy5N7gVZ5dvm9IwhDp/jGCx3lUS7Y6g+PZgpvkn8R/uc0oO0+
XMluB/rPmt/v4VhOxh1Dt/CV3FP3vdfs+lHJ153ubUeWwyCR3QHbOxACCnjC
lLfMTVxs3AwKYYNMuE3DjJWCblC6o/1FHK8oraClko7/Jm0kCpu4pHNSV610
RAdbBQSREKrKR0qPV6hNVv5sYt+RdmEg1guiVtpfX/HHNM/N5G5U+9lzQQPl
5Oeuwp3Py24yjS70mexkq3h9ZIimjaGmBcDVLGcQ8me3NHU14F/TWw1aGFaj
z9tINesPLyOuSx2Mvvhwo/O5dtdXDReqynoImWJYrBNz3EeBIEn2ZMuGLqAo
/MVzLoCx+lCbvl6ihk5QX2I+EOtN+LJzVWVH9+50Rd5qWTC6BcITquNYeP9N
tjnjYkyvQjErYvIXrMcEN35aDhHPm0xKhpe1jPLFuKtRMV8eQ8eieuAQ/q/P
KCTUDTEl+2X+sjVk8gDwfY1GDOAThPPi6DPmLCmZd+B2fzs+QAV3EK//TDyr
ZiUBSsulbAg6BOuvwzjDw1FN3Z+xWjN2RtDL1ERBGQtUiS+wbdfnvxFX7Sn3
dF5ZPxHp4XP6FPIV+4mJ7SYk6AkBG8PEzpT4KfolpaBf4LEIZAnquYPnqWBy
zthRXJgQRyrArFMQ6g9kVhlewsCSLQi0C70Vzs6rtIQWA1gPTf5y4HoCQBaA
tarCTW7Mm0pR3tcU2YwSs/mNAGQnMK1YGh7GSa5UIM7RN7SOjOBY/LVx3lGJ
TELf+4mG0YPUw0n6TMtnwoZdpG8l8Jhv82Xr6occHr0ezvEZ0APQLaPuXxoI
NQsyW6eoy9z1KY+CUkztIyOwOjDotAQ1RGjH+BHB39NycrWp3dTEGxJGu8v6
dx1+RDztwl/MhLA14rzgJruF3aPqrRQrcr0kMUPKmhxLV62G8SGl7SI017fY
RIXSFw3ikAK721iyuW8BAz4cgT80U+BMAr2B63A4z26RS4rlwGvA9m1NttBF
DGs93lLROJ8WILP0b10sFriP0uO+Xbv9s4PzydNspA00Q4jvVblCw7+Q4ww0
m5VRqtgpHUHNnuk5BODJ2P+ayzoo4tJeNDqB/RsOz7LflnB9TGaXeud9pJD4
G97Bo53eepHMed9Z8zu/boX8QjQdZHrMy3DUeDRgfoRQVW4gmWdvA9tvDuY6
ayCOJOoh8wiEYXZOc65WnG0pSDLhjODROMvXvqGlxoBMBKutHP6LnX+RqK6C
V2zku3A7PDwfko2oSWwXK0qIBEM6t+zECaX9nUL3lHe2Hy0uOieKMlhvndh8
gbJ7otaFcfSClsg+wobBVL+KoRkm+WLqgzrCb6Uk4qIyK29euQtOQi0Wngkp
CwzRk5q3g2+/s5vekAVW/0nIeJT4+J7e8fC/K87W63BlNQNs9mFPxrEA0kCl
4Pv9R6XfAh+hOZP/oo7ZpBCu04puIDb61Ph8oMXJct9byGrzXsfNYDzYJ/Hj
QrjQhxblzVzprzZgxL5oEcwdM6Lk+d+R9ZLBbrjcYN1TRA6ORok9FPj4prUC
5bQPgtDxT3CEkvrceGn3q2Lnx2MYFl1QcOdFloixGuwu7sOE5Cxt3QVG8fYW
TzCD9T3ifAFwFeVKNSF+O47NQmjhOM6UrF38llo7kPLM6nf1PxJhOJBm0fkg
oHjzJl/7DWY+NaPMOE4MFd1EyUsdD4a8HxoVyTdkBUW4+KIGsZkgyWB/H+82
scyCq2MlMWbxZC8hvjYm6eNWHzQMkVWEO3wPqA5t4naNHYO5ZJbvz3obbgHv
HP1pCgey7Pcd884Zi1k42U4TF3FaphpXLTPLdEQfssW4g3dVCxHvR+KPqmY8
6jJ8NP+uu63mwRBgczdsnshFzWLqC/3kjJoVTkmKs/E4Xwz/SPqCHZ0F0BIB
B/m64ToWiSnmdIt2pT5Z4RyCl2KF8bAEQuUMva5Ih1oD0xFwqyTDHlEz01yI
XbzBEqFDEIjDn2KuugJMNZ6CwNwRzV0S17+LIUd8TJTSu4QuJWE6nnZWAdoM
/XisHWzBxihNOTKVkvzWdCxPPt8W0z19NKUHNPaVKAPwBBpOZPpOehf8gmX0
g+qphz2MGpB09QdysBEVqvHXEPIBX44rNRF6Ot6MlVhlEbtIi03h9TxUEF2t
gReOmKzaKb+/rb5dp8eicoBKRyx96oGvWRo+fIpRcTki4ZEfup5dK3TjVz7i
MVjuc/APtFezIo1kBxhO4mlB9SIZNkR8ZBu63D0JO4H4QWAZvh8XDzinCLfa
tiKwgukL3a3KkmWw8mEzX82cRWjIF+Y3zPY+zvBuYyaSeYeOeaMOCBnMG4rb
ih3+/VY+xbKx8Yfp0+yHvi9EpNQ0IPihc5GyNa5vA/E/IlImrG6O/fLoHDFs
S5jE3NEBDuhfPSOg54vLOZjtpm/vr9yM0fCJLya+hqGr8ScHc2vb22OR7sVD
+wmjKOm5puRhThnMYjCzniFBBpjET3Gwn8aE6lglQvmKvZr9Zpew4FDBpbG7
OVjuZAtOxmuJG0HmL0u+xac1bJo3SuMkfsSbyOeXopfmijdfwXHnfJKMjSAX
RxF3FA8lB1ECeIehyE+odQUvUDnu+ecbpNP8tqW/XFLCGQ4fyJ30nkIpIG+T
jgwp5bSQonCbvP8dHFFict8no7YIPKCDL3pJT01UxCeuqRU0nAwpdohRVDDs
eOW4mBqFXmW675q2WJxIinGwfuH+muYX1pEgByUNNPUOg4zbgV4Uk1Q5hREx
4A6yKTFDHbCfKSv7m4IpAj0vt+YxiBfoN3QPDo9LwqRT4CcyX8JW469zUvsT
bv6R775R3f+hoVIqH8JpqFZxia+ijX/DZG9CwsBrNayjbDqtrIa8Rcf6TtxX
u9XzaB0ZxnZGjxwNDvrjofrRlEfy5UF011RoudObnalewB+dvD2OrKNiG8fM
VuDNil+Sf6F90gD7neOgP3mE/DuNLuHWg0Uhq0S7wj6llRSPWpGA/YvIA65Q
yTS9Sb9JrrXfGJHgd679v1lt4oMXlUHbQpHnxaQRq6UDqO63UpIHzqmjxq18
i2NnF7hEgsTkEhUCUoht38afU1a1+Gw6WRvkVkXUfFV2ZlRhNOLFR94JBuQU
wT/3My4XCPfqTu5J7++2yTovCEaBM3p5CrMUQi7qIRC4zeBqZ3RAg2eLwlUA
SLfPK3FWMgJDnE0D9IBioFc/tF0EoUEKUp/KlSsjbvvonLBEC7/E71I9cHHH
Z0U0K2qPngtJEwA4n3gWQ8Scqf37Zxed6O52MsfMlus607f3wTTHJR9cwI4W
tDy6hsA5jB+bUAJnv6/pB87Tkei7Ubq/FDA8qqOmpHHIw/atFdaV7IyWVJmU
dmRtitSWF9fYOxBA1tdnn8WLUwxEQnzGFOLD9Tc89r97xBQIXoRakTYiwyXb
fznX8wEpK7xTEDCLgmdZpshXpC8253bwqK8sjAXXs5weVV73jVltZe6Z9LS8
bxdW25TberSg9xfag8R9ODzvYoiXOzJ3tqCAGLUcRablELOwmFMpPr3UsE15
TmDTuSfGeKQjm5MRsFBmWYDPF9ypIj3CvY894NUbsQYKr5G7mdObmbuxXZJ0
aySfU2im5gPnizzkaioRI7Ch2G9x02xngN4Z9jbuUPXCmOGTcaOX+fdpikQs
OuVeNymUAep/4/grxX63VEiZISHiaGeFmK1gLXKYtW7QH7Y9tVc35DW4Xarx
V3yGcs1f0+8GUORaNimgEgKFxa7Fjt+61NH5r4rzQWiCkChVPQLj1KUaG08v
U0v6CV5nU3ZbYxYrpBZ2dT13fO3AruZLRA4ImDIk2smm07rvXx0AlF4wlHP5
5OMMNdEZz6c1KeeCcOEnClE/XBUjy0jdvynrrZcmzDsb3BgoPpHX1uVw94tB
45r0FaONrDuY4BVpGedZDjeXNDwPafvk8cjDx5DDxkcJBdiRSmjUiARCXuVF
iflmzKLcnwU9nO+OT1G5yhFgIzzvFG+vPQqoniYLrHMbE9AtszUuzisVPuS4
3MR3l6dMlReqnH/W0wDA6WnUKiLtVzoATqby+IrJPkH2VVV6e7X4T8a6r2Hx
tdR93oMu7hDNRIZO/Oq22FoPMUC0lwLjS0FNLozpEOW5UAU3COYgHvRH6Ae5
6ym45v66xQoctJRQzC0QUsxzq5vQNcG3tZBvUbjODv7isGn8dM3XI55ld9ys
uCjDDkARBeBaVeYahRlHorPeIXgkR1uDZPwjwvEDIfM1i4WnQKry4JkbaQIc
2tK+gQ+yBkJa+7td8UhQEHYKoSOyiLr+aPANmABGXbTolzrc8n8i16hPQyvr
Z0Td3uUh6H8OXDiOyJXNs7jyhPsXDdt368+FI/Ah5rc1oKCl5VL/VuGglqG5
mpWM/SSyPXQr5C1Sg352iRACJSJH9cwJP9RJf//QGmOAnvx2NHuUVp4tIWhE
vTa13Ua8i8Zu682hbQOpl5q7uBApGVwW+8PQeqRmbd3qNhw/y8QoXTkK5zjr
goXfS9137aiS/PJIUncipfsS29pEln0GrxGa+aDLygkhvMjYT/vjSXcpzVqm
B9iP2isSQP1JP5VMBOeCfuBalwxdUSKZX+dktZD6oDA0RejzeBXZt6K3GT5W
4gGC+8mDcAOxmm7X3q9rvXdt2ZTi4f7Hmdx1aplkYph//HXb+6i0j5pURt/q
qa+OLxRXvXegP5c++aLZ6689EC7RLeKrqSp7fJTRMl2msliB4PADaetwTgh4
stZ6MR2JsUx1L2gT3K0Op9G8Cw6qzlyeLfM1UPmE3UJT7eb27QzFiCXbdKZp
w/eNLzvjmSe43YdXuvZBcKaRsqbbBYbDLTlVrbl89bWXCRGnTpvHC1PqJUbv
1755gVL604wPS91LvbH4/PoMqSvIg5+rGiRUJ5k/k+i1EcsmMSTr/XlGvfHu
F4ETZzbMmAapOTS4VaklBdMGiWv5HKWCgS4QYGp84JwUUZ14UgY7EBi9Q2GT
1HsiythqLODbGkr23a1MxssM3/02rCcEe3W2Yxr4lmtKzuXNTSfUZYpSYG8G
RnJmJsp5x5wBHwVtq8A8MxvbCGqsUobAit21e+l/79WHLcaKqvQgK/VWQYci
SLcAs5mujLNr/360yJ2YJu5EVVD02ODiVJeYZztkrcrwUuutmcIlGo9IFiLl
MMvoWuE+EckPHnQJggXZ8eAwsa23y26CzrBOAVspCY58s43sGlYivUDJ1HQP
Tm2bj6WYh+SXm9wUfLjY0G/lhS/dtZVq+9GyuVO/+jJKLWbVgLahBt5AV9GQ
0zNd1LY04hMJCdYFHZgiN08Pz9H/vwpfNKslVulMwGjaa0i1d/JPY+JfBf4m
5NWsoHFvPNNpQ99zQQyDb55W/paQIXcpIvKZJTX8Xep9DAAIX/QJspNiEl0U
ryc1nQdmmiusE+4M9Y/sZ4eXQ/SJc0W9mP4nV8Ol2nt82BMmwE1MCQ+msU5F
0ZPI++7lDjNNvP2kEeioyAmSSXC17jjv1585LY/A2+74Yq5IjYjoTlZhfWxq
5ziDOcQnw6b78DelpUJ43oxE6iiXLOSyBIdSQPlyGD7BACushUruI4n5LWGc
M0VaT9vYHGoIuNQ00sJ5r0WmWfkt46QYevFxeofLR4H2zaSZv3DGRkjMqUyH
JCilbuiVGvD5DRKU3Tb6dSSsW4oJIFU/sOflXMzixHcCj3Lru4d53D4byFQd
8ziLnlAvDCrV2XG3WLAD4NI2yd9UTpD1pA+7YDdITXGJtAYFayG/kTsugtQh
6TTSVQOvo6DM3GZz0fv9CdWQ4M9fWosIowSsVf2yLevu4DTtoD3NNq65+H2u
zHsexXTXttLylLB6VbeKV1vHhUJYBcgDV1DUqXp4QDC8RhIjZWWad151C+Xp
T+i9V3g0pM6fLajmrTfoGqRKIn1mpb1S0XfYJWGhJ1aokCkuFLSg/WGCaY2t
OdRyp7dPJ7wjGJJmG8i1btY/7kxF/zkXtxQv0u1ldGahhLSSS2JZynwHbdjh
w0Kxm8tadUtVzEJPZsp36cbyJYE3ZXc8NcKlHV2StlEBGM+HW5g57GxiC4cB
FrsNSd89Yto0ZNDa8sraZypis0Y3OVQ/xc9VWIwGCFSoFIMSzOwGdg6amZtX
AGmyq3u7nhIyORfDAxt9J8aQIToDpWTBSm7Wcdad4+61S5aQhZ2sVX/zWlve
Di3yCVgd8AgpmYrZpnARQeW6UHZ41lLMjllkYtQd3yhs4HVJJthGznrX7oTK
Be+RWuz58tCJkmh8YZXx6pFbSc8IvL35vmXuJzgwyFSQef72kycLrFYWriXP
GYjEoBxBV8+R4pc6mPGRreVRe1sSUipPDnkBOzXzr8qX2N0TVxPHVoSvpqUT
D+bz3y4hCQsmRyCbhFIbqiDzycZ9WRRbURp8BbGrCG/K6byXHpII7128ql/n
828jhNftJMGdqGbUZ0SiQnWPxeO2c00XJ8n+hlugvWIG1U9ALq0S+dsEqXaL
5tqJtMq9FqIM2FUtqEhkIZaeRLnDEFSZGMGj+nrM0pubSrlsmXH4scYb70s7
A0RQMGsZTYoKbK3XhyFu401LpOc0fFT5uwOuK5YJhuyQ1N8/fReN06OpRhRM
KkbIX5ePnvd3HH0feKaeb3NegOZ5oRfQfwee9OPSKuorgd0jU1IOUg+YORFR
2kSyDDU9x3TF6DnVaOIK1GaPrg76RkIcmpIcYFjjVoZLTYhNr4AIm9Om4NgN
9VmRdHkr9xynbH0bIdY20mInxk8QBksQJCSapLqM1D0ImqkKdNqGzSDuCQOr
fcZClnKy33IHBhRRiB5LBmte7j990a+S1o88EHwmy44cvJwwA388DvrTRV5z
/wbZn9yvjTqOLmC/xnG5277i9ga/iFfSK7OyA8JuqujmnNijfjQPRgO2TMg8
OLiQ8dTGGAyRaPmTYN2eJt32FAGOvM1UDZbV3/BCBIwcgTevYGnZ4lC6gnqO
5o++4Dgv39vItnqgMZXyrZvATjULqNnY7dNWYNzdYLV6BDLbE0PUvuCkbcfI
44XwFw0/E8lMbPNNQrsAxtBtuNkzvWVGTBOJVXAld5ZXO+3sbehjv2aUzSe1
xeabvGEQVlR06lrwqHLFS4GoqrsQnTeDwxb2MEFnoXNW7+xRFFpJs8wAgEQ/
Ock+a5PUbdnTUYLBJvZe25gd3cbGaz49Kbicf6WUHZ/Zc9HvuWALIR8RC4K4
mV+BaTerpGeUO6e0vikhwo6px1cIlTUSilNo1o6FU7M1guOlW9kBGoroPeg3
ZCSgr6qXZadUr/lbzk+c6pzqKUzTVPTImXInUN98Q31VsPFdqkRwMNsjIqXc
G4Jr4VvnZ0akun4ENGAJEpLmw0PRcFNtyQ/XbJjhFgTuYTaT15WZS7Yh84Zu
c/Nekd7lIVGNrSPBph5jhFiS1E32H1llD4Z1M+iTWzCMXNDwAdnUJDnUZkVv
TKb2B+4rOLUaB4OXi5vwNb61hBHyGx8luotG2s02VPtq9vdNFCZlacDM6DC9
IIJb/dGOCm9AWG+I1II3RAcdf5oHv2DZyHfXCzz93HgtyWI6Gx47DF2WbvdM
Xa/YXxt0idfpnmpWPtICn7AsArLWMhbTUzk7Jk3E5vftwOfUlTIX5Db/Xyrd
XENZQc+oixuN5yytU5f+QaMHr9b8zmyPZp2TGb65teklrDBF2+4YdjiPZqXE
emyrdZAJPxOseBcsnyj2R5L1Nm5X0Zc6c5zr74K3tvZ+KTb1SgROsZO8OXey
P/wdVcfv1hKTmiwPgF3ygaZ9e74ePl6sN0VP9mb7Pi9IP2slyIeZTjVIdGBp
nZDFN616v7QKpCi0chLt5XCVI+CA45Tf/nIIBcEisr0S1mZmR/MSqVMvDjwk
PCPB1TgGfoDaI+DNB6GS3ISkSRwo+Fp0fRktppwu8REEuR7SlfQsyMcjoyIp
z7QIErP66XBAk+phWRKwFvRx1qTJAga12HmPosQ+EVJkGZp+AQNQlWSisxUp
88xuZDihysS91Kc1MydfoBsLdei/LVl/cjA86Yoims2Jk3Y/cvl63S1p1OAI
uSiHUvww1QQZhJKZQAO7iAE74ZJWHMdNvs14/aLwN9aSzveLARbo827krwLu
gRZ1UHthhE+yPVyKNihAuSQtOjeJB21nDf14q7cl0i0pg9DVOfjq4iETEfrS
/G9ZCgvIyIdgjRKFpKxfW8puLWeP5Kuuj6YRwWknmTZ/Y+wlX9rylLge8GUS
L5n8Fd2lwzmAsVUVDxwylMXuluM3+3a2R0bttkq803chRmJCB9CVV+X7DTcQ
85lhQrH4qdwFuYnLFvs5qI259gSSM4YHcB0vqtKpTz6khilxo22bPLPUvhk7
ay9PGkwBT/t8VSMXX+S92on1tcFux98ln9LCxqYElT/0TSZCDqeWK5A56psi
mitxva8wQ3+k3pxI0xUcktwGBuPsEgl9eu5Kl/TwIGi1GvIo3JsevXl8pGdq
HRh08fmx0NWfH0VNSSWDaJBw7KD13e8aW5KdKureuxT5hl7hwuxrllvGzMuA
UKyBMdJldHwdb/4aEpCzALGANLNSIIZaLj+TzZAwW3Dl0tbBI6tR9Mhqcez/
3qVvcZ18Uoamg4oNi3Pawy4p7BSyf1JNiwec7QTmCjOATB6YaTb8eFXBNb3S
GJ4uak8f2zW6kK2Ji2J8BORiJyweFk71PwTPc65mABHra0trn85CFdICydGP
/wTA3HOz1XQvyeEhgpemrHnHiXIUQGvNFIscIH7BkoRPNIYn/gJ9vbGxo15+
OrdBQP8uZKSU3ucsEgfJxu91uvw0L7tDBdUPEk0t4dK3qiUx1LmNoEZIGz4M
hvDSGRH1EDTZHKCn3DfNKjhT6VO/mHKiwUGExLrWUUVYplWv31LfktZDoZcq
XSiWUqV/FWcr39gdMlwE7JS7ioq34CCB2Ig8QlWJUeec/j/UwxlJVcMltgE3
3OY0TsUl2ObSaHv6NnCv/dKYnxsZ6w9yI8hs4tUWK2ZFkVEb/8M7cXUuqDag
w+P/IJ2IZXBTieC0I/Ix5UPbxTg34SEKa932jT8g+9/9yLcNeL46g5j9PZ8+
f9gm8hLYh+T+136y9mEjCaO6BCrKoWVS5xlgHgc9XuM240kHHCoXJXUiOuXQ
aS4yUEI0kmYWhXoZVQ1SZ9K5dZemahvDwjhZe7pNlmZW2IWwZmD12EZ8kwYs
aseGvQ5O9thRvVaD5wQRq5lrPXrArKVnFNjMJJtV/HgSGL+vA+zLDtxxf7+R
iRQeXNHK6y9nHNL32giWUrOdM17cN0AQ1ekxtKEPae0skdPkAWYG0C4ngAcn
yB9WMjHQ+NwnCBk/YAGNK9Q7njmXQUbHux/7y+IazsPDCuGtrqticpUMS/ov
dHlEvj8RRIJsshDCNy8EeAV6vXe1aNy/MhUtydPbhMoHn/+gQWQ6nA9wbahy
vyipVPPWJd/eEBG9LRg6THwjA7hkjo28l4dNONid5agb4RWH+OsMDAUEHJHK
TjecPM8HKrL5dzWd++RzykRcHTJmmqWzwg4DZncilPxM5l/W4W2InVVn2EN/
tZ57+ObU2gYAuPF6yLzcF662CYJ0Mi4pt22Rn7HxB7FTMU/8UfSZU/rokQ/W
oqbWdvN0UCLL4ZOhUv9+0dw9Iyp8JXLGnocJAyrRvy/0bV46yekSzOhtw06G
QOWeAOcu3u/sBm04o4Ndpeofp4cb7UIB6+NHSNu5pnhiSxwZIU1Wq72FIVHN
YQ/iFkYBpZ3/aouIFyPkzyMG7JHiDEQtf4Sez05XiGExACCdzkcTKjETuzYB
3F3TvcV4UG49eQTdrxBLC2Ot+XTbuSEgOknqr2dHbvp7cvmDW2iwZYz11A1Z
2Rycs2p40/LrdFzcZAJ70rFxFsttrvebABftLsbDd3PrCterlrp4hgDfB3uY
ChpTIm0hg1IolGv76dW2SqBmnvhsyy03wS7bD5AeyFWJqEGrqRatPtG+bs1Y
dzSns7/QmAk1Ret/Sa3qINOfjFtCcbVwNO3/rYuadqpCteuykLMv92RaWl47
OhDTKuEuL66dWZvYZuirQkVQirh0lCbt4bINW/1MTHf63ovgF23NA66hHG+4
Bua/skD94RkFlxs8ROD5krk58VesPKTB4LEULWDN1OPRgNUufe4QjWhwQJjb
O0lXBy5G2O1ilQDqP7rd1QZl5MQp0NL3JbhBnZsvhDqZN8hP3iOh6rjJwMWb
nXryxPS+hkNMlLRDUIei4gAXVuC/Rl5SlBQusIrHR4xqyRnRf3HD4JEYbyQ9
bYbqbngc/EGSMOiNfXIDu7PKbkYCoutnaohI91Thqe3PjSAnZJ83YrLUI22h
fB7ryHzYakfh/WGND7rXThSbWeQ+DRDHazREPQBHxlrnmrdtsTTl+MbSW9yN
Tj9KcEvGnq+6Th+bkB2JAh1ZCbtwhNpJQ3J5lHO7L7FiSJUsusF77iI8weU4
rudD9gsIM5Up4VxjaSQiloVrX6sTyvS7UpBLluQlfWnQieNGIfAlPrmrjvYM
XYUfSmWykK957kThagIzGJBn43VgHs/3JZif/8IPvnyoyVHBFuxUtFmp4lEF
spG4GzPbFSOQcJ1XvonfRTUOoe4DeitGq3ESjCgKnF2oTpP4UAV1U2hPeE1f
YW68DtP+CLeor2kDDWeJgpW7CIxleNjzcZX5qCuSW8DL1c/wk+iszxu1CMMy
PTtnwD2Hq/6UFut/s5ya3BhZ4fb8s0zOOShpcM2lCIZcrqEopdm72sBYL0Z0
kmpOpRNkwPAqSDodW9uKUFp4wqaUucAe/LsTk0jLFyrh7YgZwruOkDGEUfrg
kmB3jGrkedIfReTDoB4Q4e5Tg46WS/Byu2y4fZQO7NREVMgjwYbxpUbBcIK4
d5h8My6ZdhUTSHQOg1nycaGL++rMqBtuYABhKl+sGmja3HDdMjPCW0JFjL+Y
2JtrPlRwIiRq8zfs2x4osRPUx4qML4N1jpj0j7mgBUBMwoUjyZbd/IG6fI2D
H5TLyKqq+1jmuqtC6JOSXdyVSdJb06PSUXlyHHwiSCs4THM088L+PoSS+YSx
jr92JU8qHsq9jB+gCaaNjJPDX41UmPsfLtEdlfAFnAIKVPv97eXNE85VZZPS
bUmeHXBlrxPxuFOwUCO1slB9M5iOdsW0TXEH2oPOrNR6L4OwcbW0jiKaJQs5
9I7ew8X/7cllBYTGy4VlcoZpTn6OsZi7jUt9/X0bHUaWSu9d4Ma359EsAG9k
+Z+l5PXcMPyeryMjCwVCp48vi/Qa55eMhsXcyWaHXYXddsAsthuFHdZUxozx
gVLQXckQrnNNEPV1LA4E+nQKwPyO5jLR+bE9igOz9x9KIU/xo3SClSG4Gz9G
qJXa/9mqdhU09ttkL9KhQHUTiN/EBywE2u4X2gI1qg5btztZahZ2k1Uc06M3
Ss9AZprSkVjlqjltuqipbkBsLJsKJJYi6hw69LmzaIasQX1PgsCFwmIhuKQI
Vg0N7Yp9O0GfA9IBkHv86FeVALiEnIkJU70LTKzz6FU7AV24Ocppfn2xSXQM
Y5xw7L/79k+Axc9PQpcPcOav7jwfAk24VZUWzG+Rmxw7k4LF9fx0GQ+Rs385
Yuj5U9ooXXYzr8SaSAAd942eXt3/qWLPJUMBag8384nOtj9FB4cbbo4jcTl/
1woaEGITD07O10TGayfVi2ETwCmJolnpFS3Dtc1kwpdEs9Ao4z93nZHgpAhI
nCjNmbVI9PoRiEM+2NQAipSbcnV8Ez4cMNn5TEoKioGxyfKzJl0DFCa0lo8v
vtUDaziYIZY0K+/V9IaTmO8MEHeEayKcb6plbgyqzcopE0OXBwxODpV2I32k
fT5A+/DAjWWuaXScLqjtghQxKW22GnQuWq6P4SWeBJcInJgSHbehveaEgT7e
3ldNjIecwweUmuPThEC8WCFmUoza7t5+pjTMfuQHNS8ul8X5WbBnV44y4rmU
V34k6xPQxZEyucigWcwcLMAMfrKgSeejU9lgB7x3fs/i9fQDbomTcySemui4
kWeq6SYIWZm7I8cVzfquigq2WF/SbM25XjpoCAmtYZLkjaB+S0VkLcrBGYIU
+8r1hOY2m/j6210nN5thDf54I4hK+zQsoqLenpC4MWYIiG3gC41MM5UAgmut
bJi2btfNOqmtAsaAi/2eQQkRauA+8EBVd69depBLQY1Mj+CvyKVboXRRzvkT
ZFzlNYpr9fW3cn2grj+z4YWt9Sx2h9StllXolDt5rbqbbbRm2U8m5AIOU6JR
Y/1eKUGSCBZVs2WV+iVi3YZFHjheoac4unIrce3VSrH2LH93arqmwifxxYGO
VM5lT0wcRXA4w37/mmUKZb5gYJHwRchvfJt88eoACSZBOAQIwcznJp/t2RC8
0sGi81TZ0eImOMt7SNpt6Xgs08/ZTemsE/9Cs6Pwo6F4P7lyBRTnji+f8YGY
ZKEA4oOJR/oZmWVRGrsKtjbXDBMgpt+geR3m3rWYMNqnijC89bxqoT1780Kj
S4AXSb8N4p8kMVU/Ixshfch/3VBpyEMbjm3iQcFEDBo8Yhz9cH2U7uy2H88U
0Ew1g5IYLE0r8LLb2cxz4gqHGDKp0rfmMlIUGQwZJB9Y3liuMCvjmnVmAHTb
H++Ck+5AfFdfzP+6xeDfsarvMj9+eGUPOrmNLcm37shxBqXKjFCRFIYxM41v
hMefiUCvcjULqQtv8thIPwZ2daw2SUe9LTSl0pJgVO8hdXG7wG+EYYuzSZGX
W+2ggESQSIxZPe+Az5xs8osp4ZAjeIGy0h1O7jSNR7TyC5Fj6hNVF7G28YG/
+jo3Vyr/o+tRBR0zndasDJIOzYoU2mZhfXhizE4uCOd8dR6BR1jmR8ekqdni
hD4VcFB5pfXN26iLRBzQCz+k1JsZcIJUXMfVw8HsiUSjhnJ4qdhl7zu6pfTA
zoTlJJTvHU9wjYxX/4prXPnN8Izp6YHscA/h7X6LA4JidPQ3uzcxi5yjp9tq
WCGAOEj92eMoTTpAeC98q/LAExaCNu7dyaEk0gYmpRVgjV7RsMooSaFzAMNE
wH8vHh9sWKg6hwRizFm/cy6LpaYz5yjNCXSCzyMzkq+Jj9a3VV/gfMY80pdY
tcvIW2wPajs6pXDwaLwQEy3Fk5o07A0bDFiIDyRhnDn5E+J2lDgIlvJAlgON
7Up/+In1H802noGBbHIWU0qx4PzKy4s2mitr3AwRoCUb8xYCtsKOLZwzfmx0
PUGoNw487Q3UYrTehVtgSlRtEOalkhSBAL2KGU1q0ayLJCQ6pL+WV9XnysEv
i0yIBXcsGk3aEKj9zkOb4yJ5TuYSOx64piTHXBb7SkIILBgLpq54UWKZgqko
nL0thzsxZGceFqO3845XsXHi+2oXBsnjRfoC+2TtSwICgv/xgmOJSLZRXGN8
9HeCObbkUoRLbD6HcP74Z5TFxn9imeuvfLfpnWcjEAqzXuNufxbACaVNCKSP
v0kySbb5e77HNPn0HTS0J0hvuROdsoTM+KiO0HFqlJbo1fg2vMpktHXf9I6x
mNCjQHKvP8Z8uM4FqEQsscdTNtkBF1vH6aB/KgBEfjiRz6rRyqlrwrolMq1W
v2PPaIQ/aaqg3QnHMd9KFyakF+zd+gcxk24CV5crF9FJcGg42lxfTQ/IAgDf
RFakT8113xUOYb7X0JnOlEOx7pIfnrHpfgTLTLOUHlyIXtyQfPD3aPsEPcoc
prJTg4ZzGrPUsog+aKBpKkJj7h/KigN/5z7O8QC0lunKfrop034zg7qZW8jC
/3Opcv9jSx3DBvo0yHUXrYfPeRMEG5B5lztC9aYJC/ogs8Mp6PTcLcq8RVLy
rQsf6HGLdVH4GC0QE/74bJ55vv02RNaLdHTcu1ea1yHFVyiEcmZHS+Xo5KPM
Mrx5ZScFnnttJB2xS2wrl7WBMtzHlpSS7JkldgOXsAyD0GyqCvD+0dEsGmbz
z7MQm6Bb/pWXhmwo2z6SnUL3QSrIVQ85Dq1gpafYAZ0Hp19fXNsv/fSsH3tP
OlBwOIXwOpqdbrGIG5L3o5FVxd3f+DdqfhXzQWukDinYjfrkHQ+QNxBdbMuF
KO25EqIewmzbSBJCBOoOAFz3qa6Ay2q4ANtu2+AxZtfDcZ6P0GdUqEWDeRGw
ReEOvDzpms3e4ZuA9i7ygguHEDmzopnS6Oj93peBkKyTAU6R49L+51EpWJth
g0IamS/gmhDk/UdWrCeyuhr11B9RVcWmP5h5yLQzUkIbTBNbc3bNCXngFstk
9Ta+juwSPTJX7A5cAhTj8szs6udj3R8gllM/K5bgwadUNbVvD6/x0u/U9TRJ
EPwsdXKZI/OVuWV/zd67Q8kBBh9F4mbAmqs9D1+dJOJFRAp+6esqaYPagZv2
j/iO4E0QvE6R4xlUmkkb7zFnhxcU4j9xBUXx0ID5toNgEebtwnzHuVLdqh/Z
/7zCsxIo8czo7SOqNWiMi8oG7RTnlwnFUNd9XIxXy8h2BlwdfXA1niUdDdDr
L3cA+2T6seXxihb5hWxuul4FfBzzlkHN/E6Ul4tIO2Ol3CFJeIRk4VV2kmEH
8SCDgmaNGoBD0ht/mIS8zEtxZtGA+gLnmOkkMm1NvRlmHrNPoKfE8ygaeKKv
nf+V1bCdKHM2mjS2y/pMRdgnYO/izm7nnoz1uQlOjowF3C0noS15Ia7TeYho
M6/lw/KsC6x7LDZypMRTO9pBwesbseDc+cfbtjmduCc86eLMHnPybQhTdBEJ
egWg1EkYNJF7k4+C0zTPCLVSxJwHk0ZEffctcDDoHfhhYGbQ27CjiFhK+Z4s
zndn7FsoSoUm4xQVzwJafMZGCJATxckPKkB3XobKcACnxfzPu3j5hHoiYvxO
hw4dZ4u97V2Vz99kOBrVwFkov3Gd1CH3MOR8oc+GhY0QEXZt5W2tXI+rBezu
o7mhDWCldqHriV01h6ny+kwd75zbRJXmT6jXC+meWXms+yOLC+jX/rJwh5by
zlW+/dN5Rm42zCBfOEYadD/1yE4pBxjDHgUZmN0rKOyTQA/l2QD4Byrk1DPa
sC0XvYm26YdW+9lknijA/N41YBwSSDNvfV39H5nZH4Nu1k9E/Bk9gAIlcPnY
SoVuod8TEoghA5eH+zL5vnuGjwPcvh0gJK1ToZhR8vbfoeCHWcG3D1s8u7HH
Zt40H9fT7RNuxO7t/rYyGFdgrZzlB4L5rC04x7vefBlouJsDbItWeAZsmSME
oG3sjHLcI2OaGkJS9KVl7fIGAXDYFSRD/VJ0NXfg3p1RRM1Zpg1oPXO1N9ln
sL9/jJrkIF1VPl1i7nj3OBQT7Zu7Ywne+yo9CP7cH8rN0z7jrrNogl8W845i
ViVl7gzQgJpMhWnkbSi0w6VNY18ajKCauV3oQpAA7MZvkAbrPBu/dBI6xUUx
IT/HG+tWNREpTrJbLOglAtOu6gOYEZDorlc9O2wafbyevv1FswwEyRtEMOgE
UhhI4hkmaFnpSHzc5kiJ0rd8sv7F9ZUCDJYKF4YGgfAmJEmgdYhaLznrvhdR
U00xpaAO1V9I4H7s54qd1VCqRsiy7KRZNStQysceCYdfJSJCvtXJSaOwRblv
dprXxmthHK30V5S27TGkz6OE5i3eVndWbz+aBzGHUQ1rz1QUjIdfqReAtbGF
eEbC5I78/nYYP8q2TWuczlYGZgRYzAqpAH7V0GDnd3pk8u2mkzdZOLVH6l84
UoD60fMRBm7eBl6yFvXWIKqmpcl3ex3R7ytz//Xo+8JSYp97PVIDKfGHUNAf
Ddj4V6+87vFmqxANm8du9jqNRkzP71SlKH+w5cQ2naRSrQtWSLfK42wUxK4A
AKY7fBto5ctyIOet885TEymXpU/ubEb3E8ceDBaGcRdV1+RyGYvbJHa499iL
EM9nUVhDS82999THG3BEOfd2pLEaVTnX4B6XyF+zhIXGUf80TvVubATJA4Zk
ZbnWqlRSV6v3TsgwNyqnZ9ZFb3PK7uu7o8eFn8FVmMFI7V2yBHO+/NlCBXqf
v4ZNUmqzSogUocOnI588Wo9wEvHx1dDjaIizd+mgzwwTn8EcoQREOuFRFrRg
BoGvCgBf9bjGPZHUTgB54vK092muXSl4wBO9RveiSPxwKYyEt1dEjTEwOjps
2NhFcLWTQ4N9iuY61AuLuyHaJlVwE5HyHB82XKBE2E1TuO12yOeOBlNBR6Sw
tH9007IdBp8HYuB4Ng//F+TyXA9wDLRLt8dMaKp5W7kEJ96f0H6U9EOgIjv6
awPu5ZJu08r9TeDcfKllQ8TBOETwHxRSDCqn+Iv56tz7kL0kK94KTKuj59CF
bdKBYiMAbOHfYCXgjw7gLZOmvC2yXRbPXPtvJA9mlQQ7jaT9y6D9xCjn8zES
adCl5cJlmy7N7TZ4wimI9c6c8kCKT62tiCQGkcCcjIiFiAlR0owcB3yESXlb
+0UMe6p/UWdSLU49IMvskm6WP++AQHhsSzjc1TrXARn8+N9cjmJBIuAPmooO
yMuEd/3jNs9XXcP2ABobBkJGg31aQPl6dG2s/TMxx/hFkfKfOQKfao/FS6KN
cD/pjoiCareUfchHMDk1zl7xGtqNvyLvnNidLW2ScZMEW36Gq6+1sSybE68n
4gDpk4n7I5T1mhNeEPxbbqYtBFZAv97xTwvDLO1Oil0b1YGvFmt+5sVTCOnD
3eHDEjDIPtJCZB3axEiwQtklgbgvnAy47Nk067xVo0Lq/VfqxXOhiS9b80tD
TYKj+fGbhxZdfkpGPFi2r6OjJ+OVf2oqMKrHukKgY1ovQucvgiRWNTD4tBWi
/4xmG7GtpZ8QcsaWbyW3V3kWGJ48+nFb3VxIXpKDnWlwM7hmmT2r6i882yzX
Zfbd7AGy2zJNv4fAHECblZ5SRzQFfa5YHlxuRmdkQjqgN+TMrILHerAXvCnY
SDJyO5+i5c0jbZfB+yGRDB20MNdYpELE/tWXOcquMW6B0WvufFcxHZmt0vH6
XY/nOx5jmHPNzSURw804lVWnzXmygfnqMN0wAXZJIvPodLbtBuEC5gAa7Nqa
e8Yqk6ONIZlVBVi75etnwpJ828U6zAMTYXQKIedco7pyHFnspj3CeTIReTep
6Kaax057ybHUf3aiyNwPLOKMmQkZ2xODpvtrNFA7UvIGnfEG/ucqSZr3RZTP
KIyvyPXLsW/+C1uNfOraf89J2YcfROVTbUtyTaV/h/frnF4jBpCMoetd5SLO
E3o02FWLcT65BDPDydBzTDQRg9lPNdhbPZzRFCXTiqNaN79Y5OAYBpTY2wOp
ZHqJ5D6yDQDT9GP3k387cGVi9xnIHdEp25wpk5WmQL/dpUTIYdI/rOK2Jtve
GPjwhfCeMqYZ0tvXi15o2BBG2L9i82/VpwvhuUtxyLBSeKIbi08wp+alxjcS
V5eCYtUQsr5bj69bNQ91PnImIUznNT8YJkcxLWKmiaTqqETJ7mriC/f+hFmm
AMmcEHicjeg5zl98WxobZTvrM6pNJ6G4JkmODO+7JSnfMVI4vpxXWY3lfbW6
DsPyVGhkXaTuDsRdfQfvCx6KuWsxMR+pPZ6gGwh/0ANcVPX0U3UBopUQxEkD
U/AfmMVt1z2qqUhDxoY+Fk3kYHgYgr21AG4ATaZlPMpA5w3RGpTqWO6j9vfl
FTAk1wPwtu1NHLAqc4IF7hnsjEgm+D+rssivok2x0jRy2CLMjtD517tVG+AH
Nd/4TiE6tm/hMjMmR3JOMyWCrIRLWPyeuyiReKpXt4cc3Esv1BThTRVxcPTB
B5UrE9x/+a6+CuqGDZ4b2iITQgSvk8u9Ku8YaJs+9X0xDEhVPavnqPK2AKpy
/KAlGZ1gGNDqZlfZ7w6P+qkYv1JlWg904GUvoo7oaRneM/jI+JU6eNTZQtlA
I3O1K8Pkmr+N2eYjC4DvyYbL3f+XeavfCcw7/lewmeoQFk4T4LDnbBPZhdA7
ApvAhkGH2IpBqY2FR0Nry8VXjVbJI5J3WcqONCNu7/1NEfR7Tyq1klOwfQ6L
mHfEgrnZPYvHZH1y7bkC+a9SS6kXJEu5098DLHnjQ1JWlXqIwNDQMEb/kc8B
A/ClWHCITxN5CPzwvlFAufgVDmvPy6UR1dcjI0VShSZFPvTVU2w2MpojO86Y
RKaFbHN/zDIFpfoFO4MxOo3vcq1BmQo19b84nVu9MddaXZF9Hus90MUMV8+f
Uqz1TXYNnsQGmzIAYGX0bnWX99B687UBDFcKRJP6AHcDg61hPGKdL7aflSQo
2v0gEIwTldg/a8ZUw4JRXs01IoKya0WA/Ce0Aq9jKJsugPEWD4CvDuZqnGwK
NvoqAwhjDrh8i1BQEcGmObLPduyi6p7F2x9yREahIl5CfYfWpuySaV2ecXZd
VIt6zi2QCaKJDt/wlJ2gIGSVduVlBGG7C7osEJZxRPU5GVZEBSMSYZPfaTds
khi/05egLtjSPGNKp5ALUoCgLWRAfnW2jV6Jr4NNs5KAXLLfQsu1F72KZMRI
f5FYHgwnrh/LIh4nV34QFXJbd0IfXaHW4hzQjerXfcZEEaBfB3D7K1ztTaAB
hSxxTEvSdjqSsNXYRjDsRTVX1EfHrUsaeLFt23eX4XJSWJEi4KzHq3/HJSCr
clB7up0ha+Kjw9B1UBD35BRdyc1RYtJG/xG8aOsUWT4f6UPF/5ubClmet4vG
93Qycai6z/rTo6mo2sE+dTHxi5ctJTtNKYFxlNQNf+NWqBljldIXh6RSD7Oz
LK5IprVDr1dEHGH8f59ufbRVa1f9Fq1nmJKTsMceBsdrs9UwZG9XeNCT72kp
nHOWte3Sjv2ZBXSxcYZhnla47DptmsMgUPcNIca9fzWKon5rDjhqV546w8Gb
MVCSQ4AuPCAQXxGSBoJu82yEIIwjog3EkM+GHqdvnpmc0sdnAs/lCI7IwZWT
3bKK1j71qgxw+Qqv47B1jRwobnX0AyO5JmzgCnvwNJTogqzYhIkGwh6mDSe3
UsriSuUycg0HSdFzkKE+6vuvSts71ESFhOf4LPOWdHNTsOzUoxrndTr9YyiD
WErUokaqu9Fj4hgy/yXmT2LGQ2tce9yipDTTYSNKtgZmOaBx1GYuAvrBshVv
W88I33NTnQgLM7dJZ0S3OiNMB41n1C4hk0FSuYWzRMAOJ+5Ihtrtyghao7o3
FVXihlGCXJCxAOnWwYsxWx9bTN9xkJaxDLss/fZIeFRezex7f4GodfwmE0Rm
OtUZjoBh2X00MJHptOrA0TyYQGdmAg+o71297ZjKDPdEV0mLDX+6+1pf+8WC
kfcdcNFYSGH4NCf6ugduzTAt/VT8kVGTIdstD33wtmP7HP4UwPw4JW5v0ut8
w3TJZ8gCnzxtAMnMKAItLVOSBsToMPIIY7BGTCjCXx4//OptE0+rN1JF7TO9
GGa4E9HII5hdKX5bGWEf4whuBP5hRdhcsX+6YMmVjWQk89EkjrSOPtz2VKxT
iGRsfRZuLH+TZAehgh8C4ucSovgJEU6iDMHM7G3wInDdFnwvNRORQ+ZWs8A4
DhpRyjE0nHUhNJDO+KbNDw1jxUR9xIYyN+mZaIuYC9YB9vBd0s91FyMbUrUQ
gBRJvgobf1x5calhmuo5KjABuunGbPk4jcMgwA5+oPGDixxZAOhLAqHbQ9/t
zNsKQGqBJMdOVs6aXgXrE0Kb2fgL0eS5bWaGMTTHF8tCVq62DbRQQ7yLiYbK
rYe4QCE+qk7LJcPV9PaxzbuCMqHXard08ZwHBY2iiWUJZ7uqeYEjMArMCLCx
YGPlLO+TLjm4s65/3PEyS6j8DeyjPRCMCGYzfhWgjLGx3mhCl9J8UGnKSbeJ
o0r9vdQ8slBWYPRsxBE40Kc7E43hhVRgPQyPeUoKA3UBxbfJwZy5wjmbCVo4
2djAuPW+tAvB3jCRgf1SZdLKqR0K5dCDmZoyhuGzZFcixAPscwyT2I319mNk
PSm7r5wVo6FduRkbQlqQmmu5g7HVigMlwkICeotrJNOxNkx7+svQOmc19E76
gPMoVFJS1mHyUoRgR/uimljX0OiDl6YRCERWVLZTf2aJ6+nR6qdSwleHwM9h
3Qk0MWrwmXwZjiihRwUsG0DpXJdaVignXHaesKhMrKtgxyeTV2jXkPCNFKWe
dXa1JwUHZ8aBsKr4mkGvCVB708DKNSGWIoZ0RDk/tzQ0Kw7XEDmiLqtoVOF6
GeedmrOf8+afg/GVSZVHuf3bBkHkvADnpyN/KKe6KKWXuzTnPvcKS8Jgi+sy
BmzRjFHxtgqYLF1+N2pbYgx7wcqWoMFDZ6YeLErFA57au9uJLx/qVKwEShqb
lqVrSTssCj4tzSwkfZDt2elsl8++r5evsisX5IgplAhPipERGNhol0E2LtqJ
K6JndLZFAKL9i6E4LaMhCdINUc3C3u3Rwuey6JqcuoPlEKWLCwcsPgafDEjm
20dTx2HHzzGulZgcVy2gpWIdqNyMYgGbcvenizW0eeA7LU7PJZRCqwK0Oht9
Mhcfr3/RwQm1OXG3G3SV+EbxZmZskoEUPu51NXrEy6z9uqSRQHqQJ34kDoJf
QHIpu8NLhnlUnG3iGqeRA1qnz4AdG0+6dDYpam0ml0zSY0VHstOjOthiNaVr
3+lOtNAPmb5FK7UkhslJCCB66DX1M1vGMOJCXxdsGuvYeZ/SeLpMyO50Csl6
f2mfMEYvwf8U8rOYmQB9e7yladTZ1ZAsrNJNkfK+3jbTdWdq0gmJ65hDDxBc
LbeUvExEGPnRLAneErsL2xkOSLx3JyTXwa0lghfX7uJChVgWDK7GE/e5hRzr
XeNpSwYBFTs2P6a5yaGqWStNtHBvTr6RwGG6SO/idOrwm4xMsCYWXcPxNsoz
0kjZkbuzM0wSTSCd9MlhJskFLrZ+UWVRSZirvsrr98AcYWpks4cNgiZ8xyV8
aQJFq0WYrAXTVsMhGyXoS3UpIIxNsLAUil9kuAZ2zdxWjT8yenvw2fRscFaN
c0o9VWg6p1yl7MQO58fcxLRgGtoVylY54dyoQewRMUiMz2+KeXC3kcu+ErdH
G8QRVWnOVyIHcdDtsTs8pOyedpdN3270LuWmib5KF4g8RCj4ys5aGCJ+mKyq
Nuot18/JlG0IJmRwAIa0YfYqDX9mlP30ljJQNUQ0JXBiy2DS+ivo6GFDCcXM
5wzR0v08QCMZ2vNiMj7Jbqx71mMU6eK6FQkjkGDqztKgwpOypHPJhVm51AQT
irHqTePHhf4irOBokAt+10iZvkSl0AX023cYfh5XwYbTtCwHKHf18aF7mToQ
6Vt7girejoMCF0S3P5N37DLORkofz3+fqBm17MrmUrO2AXFZFJzJXgY27Wa1
yBbO/pSwFTlEET8QjFzn8EdaSrG9r+iwHrQ1COHF9Gt1KRUvYOSkzbYYFE6c
DdNOZhB6Vbk/K+Vb7qxIO9MfMKK4ABsXYK4xvArjvNznPxmMGqrM6O+tECf3
+Jf+JP70jdy78+STqPaiUM/1KP0AXKMFgE7kmGoVruKbQIsDdrkSJRVCbz9D
xyxmSj6fz5uPp62c5P6moM2QhuE+vDowzlHD7LPbKnG9pPllKRD7ONCwOpup
S2Bq1HtJKPHZ00t3hIVWjnJiZiHK8EC3wwE+DcwdcRhd5yGlMrzKLJhrvo+w
4214psMjxrg0dgIAGdAu++n56e7MndUUGNTPGbFzFJ9t7gr9X/Oh1bDygZyi
O1l8BngDINSV+ssC5psE7Wk+4F3b8DhvyjPOEKVJsf4/FYXtOZnVm4g4Z0AB
YrsZDGbsacGqlyweY3UGBKpUZM6USfk+OdIhHRqJqv5nLREUSNw+fbCcKDfY
lFCq1f5QJaYRI8t+o6YdCWkagigvzqNlUKO974ZNEdB/jLaYJuRwSC/JpRGt
QyLio9HRGsDaIaTL3gfTalEcjocWk7CXnmumZRa8liFSpEaWv+pQ/2wIDWnd
hAkmJEdU54tTMdg0kG6/W02loLWAHenbk/gx5oB66Rp6Tt3LVO3lmyleC3Vt
UzAlrNSmzI22ZYGobbkNmBvpm2rJeuG0GRqKewegfeih4j1xDWVA+Bkl4/mJ
Khl0Y8WE4GsSMnVual3NueAON+fCo0bkqeESiMx1kCUKi22pvzCKr0foYbnv
xylSz25PxXtN5AWqfF0vYZ+fS+vyOXJ3DldC/VUKfTm4/Npelsb3LySyOcGe
rTjZU7aPzzBq3O/3Va/2KIes153744B8FhW3noNuZmdhFrFeI5aA9c6Gcn0Y
IAMRPZlcIq75y5JOEzMbaCXR9uR1eaqGA/gziQv+U/uOONnT17OxBWA6iQKx
z2uqxsUKPzyfL/HGfojb4u06/dWsOImYjCeM+pM8/fRh/n3B0HITBuPzubGz
OdTVicVhtsMTf0rhCo0A7mCfGa8nHmcwjETKCLSKRNBC6y4E1fFkZgG471AQ
D+Bv5pmsauyrKR0+kRP+vT2vX3Ilu+ZeoT7/9JON/4EW8s1rTdf7yIGu6v+H
mH4H9mbYAlzzK1gDf6YyHQO98W8FEmaJ46AWTCtgotOPumx/nJrfSjEORIWU
OAmdzy4BP30m8LTZRQ6dV08rVX2Vqp5DMAYIWlhTuTI5cKqFfXYvoXr1MsPV
1R5RNuhZcyZ/YNfoprhbj5NvdEgERKsUcfSKRvDxoEYETi2+1MCWZE0Ev3ql
sGSU+DGV2O9gTALWBds+ie/q03qSpOrvlX+wVZA85B6R63tPe5zZYZuXsFDw
rS6hq+2un/II4dlLymq0sr1TKCcdMrVRILQp42o8KIN2U1WcnSjeasKv8ZRW
RjNlumO6aW2R2P+gVBcjJhL5x3QgIwudHfELHcUK2tAo40dBwvkqRc6QoTtW
1Ug8+VMerFAjGKbeF9PPfwNoV7ybQlQVo0yp5ebP2FO/D4IZ4wAf8G9FVSi6
gtPgyu1AlgU7FK8s9LEtXLhrF4xX1bgrBCbMV7Fnedd7ed1CSPyrSvuFwe1R
xk3283JyuYKDyXs+NO1iVFQHfhDCi4SqnbBrJUFXi0ASMwj6V9I0nQfZk0CU
Z6LM2XKvEcoODHY7jLYgZF7l7mcOcT0VIhDsVPyZtp7u658IwmBz/Do0xSjs
c6KkkVChz/aUsy0OCkdv2yQQWc8P1/qBrp+CM/ZkO8sqy2Tz+fZrimDgIAjt
K3G1yMogLPDoRq20EaKnXfQsqmIaL5zgHZT0Sf8fYcDgSLbPJ0sW+0W6T3M+
+8bIvtpounPNaAHbF47s1lBRx75IsAQ3zBh4xDXkFths/4ACTy+gmtXnbRxh
CBmxRAc5MMyU4jQYiQqo0v3EwMwry1OWF9TkB35u6OAP1pO90Gsh7rtUe/bV
l/Rv4Yjj9G6DRljf4ExUVuiWHpXh9/fg/2UuVSDWSlJWcNStBE55eO2Owr7Q
fgC0eTcDsnQKs/87r5hid668fNq90+cb3sfujqqDouLUBksBxYMz0R+oAFLx
s9xfv36utrLTlGn5EL69QUgcuD7H+RhtUPnww2g4eCdvRxcUYGood/rS3CbJ
yWGmsHLqDUEEGX5PU/i6VgUmlv8QMSGVL3NF3tHA5MXUCNg7CsgX2M8pNtNX
YjIVr0v6j4LP4lW8PGxhCabOzcr7ArM/mSvwGWbKwOABEjJIwOLDND9DHH3I
ilFaT94LuzUaRmoXKivywPrDZUyCLWxWLHOCiEoMQp7Mbgt4O1vmhppJ3yfS
cBpWsxLIy0LgA9SUtnfTtpQEmHkTdhl17AeboASv+4/efAXKwFLZI/vO9av+
9uteNudkvmTQvrZJeZLFmsIl9n6pstfbQj1/dgeVtIuLV0y5pwSIEaUw4jM4
629OJ5wKx2xVLNGa05Lws1ni550iPUjFEATXAFjq4a1eq3XTJwPglunpoim6
8x4+iqk84N0vZEYnz/joek+WE7cxJQSdkUCMDQItFeozdyVH8X+yWfmjfbLQ
yQUnbo4u/8SMxX0mxyWSK3TcafG2kMLMTQ8bb6r9vBzdS70H+I7sxiGA8E6W
8w8IV10JXyWH23+DcKJi7V0ToJrORlLKb8c0Jv+D2o6d1matMY4JKvfZgMaS
sKuVextxZ/HvRYnqaCHDHzn7/ToD4OYH+bT429D8M8vEq+phAR2FiezQ/Wuu
ioxP+nCox+M80RqZjRgzUaZ14cvU8aGHVmTn5XOyPlSXCfHkR3yfDDtBIeTE
iMjskemSKaSwWcBqqGi2Wu7IAqaW4EEuI3Xhdy6pLQ3CVHC1GOpI/oR4d13S
zslvpZ7BUcMVTb5Rhq2fCL4Tly2B0FQ2uIo38NmEVMlNiDcvDcuCP38fl4ck
zRMLi0hFyHpyx3ESh8+h9VxSNHJXlBXlnlkRjTPy83IhWrN08+xMq/djOrl6
fzfCpxTegGMTyl0hX9A+8lSkPRFFZ1U6SNN+N2HLhMRiBZzz2WOBBLMrGLut
5piIYEeDaPUe+Z6r5ECNJpT6tgAVkNLFxiXtzoZ5l3edU7FjJYpCvPSKwAyS
/ANPEUgN+ZIQURtdIZxxmn/XSsYrtK3g9Y3gqS+ICLq+IwBESSWON9b+zqeU
GQbnC+alI0xG2mDcQBjYPGsBoPMCcu0AoDbCWpJpzbVkr2j7NoCRXU6J/N8A
uhzIjnY3oREhNHWcxg3Gc6mcZY7YPQZuSWf5IfRySjMVg3QVxCDlOQvaqSLh
gOV7EenlaCDe6sYD2ZSOB4WFqf+UYgxL50YJ+eVGpmFXLSgua639tSP5UvtI
7xMgQqRih511n+ouyg9WBhIyu2l9SGXLlOdIcWXPRjYdL8jBdpIj03ZtrqLj
jD3jhD410i46PCKgKPvCLwlK2R3XjAWRWTVc//cDWvgY6mYLFSjq7YKCi62q
ZTSns4pN4ho6w/jLDMvYsxuGHf9oumAAD2DKTxUwnCrDv/SM2hYsA5LCiPhE
iWrPqYd/RdVLtRkEMeRWU/Et3n4273vX4GhIyhcgn52wJC8H+9IFlYiLnYMG
oPIiyQSHNytn/eN7cLNcuKtWtQcZw0HHmDBf6+rdJ2NjbV/H6qXh9lh2naHT
T8BmvK03iiyfLP6ShCn31eQ3pG9mehKEDnbWstqmJJQHhR47FsniKCbES0SQ
agXMzVK5qys9A9dRKu9XVvD+VH7Iu41YxO/TiLo8H5Gdebze16tUR5lZm30b
XUx/WDYv6GeLiPji1mBjF8jPKOe0sPY0iZ9JpFSyoh2FrGroC66SjGi+4GKf
DMR+bdqaejRfr50px+tPYBduyE46ti00lYvmecnvO3lRt2ZiLIzccjaTWAkM
EyNKAtOFEek6RwnPwWwDsu63tfdO2FIUe/qV5pYMv4qo1uvraCdbH+iHfKIk
47mL1aTmjHlFB1r8eSfjewdkc84YaenGpFGkyhk3jFj5lQsjKqIO5atGkPNd
Pol8kVg08IH7xUaHf1tubrANz8zkuD2sKtyb7ZuIEc0UGwlKR5S7osx1lPXF
ugmGKboZY84v7HQ3qO4Z2b1Xv7LDUztydZQqkqtN3lt/i2O6Vs3sBWyRbiXL
YcgnR37OXZE+OV7K7hY4n9EKoQ4pq7deyHIL/zIjDwKHqo1f5hDpr5SOR6Bt
bdsmidsz1fkMyX2KfOQSyPQegeghBD+2KaOfSG3+eArfb9pXSP27c7Lo+VYF
uUjXi7zuw5hkC6RMK7UU1VSmNJaTlSu1PZUsOpbMNOoZXqEmcg6BIWhJ3p/q
I6y06vZFWLgpCzAwIH6mmAZ9sF7m92egjSAoyxJjSsdKs0J9iKg4h9E157Bk
48h3ukBbwVVqentbNh0nUkKOda3RGPJmNGAIljVRLsmuZPy8AsD0toIP9CLR
0etWFOMIUCkWKbkA95wKxzQU1Vl5RB1vPId2EhSYfDdEVsURDTBFXFFQQOkS
AJxjqJvsJex+LvddOxAnr+SsDXDU+ups8Rmt0vgBtVGimjH37F/PYeuQ9ASs
wQLkgvo7+pkKZGQICL+cPf+Lu0nmHhoqQlOp37Ph2UGfz3Owok4p/y2xyA0B
KFme6OiI8LiqdHE38NcW/5Lt7217ACnvS6s081BT81JS1RZ0KNKCRwgLe5Kc
j/2jZaA2LAthRR4UpuY4N5iDBSt2NblESAG++fD8aP0aPyIEVGzJlNHKcgTu
s7vjTUjWfg5O5PRMzpEiFzUxsn8Z9Mb2KJpZzMAIDZb/zIO9tZvLJXcX9Jxo
YZL+0Ev5tUC9mSxInkMW8fnQYIVlBMh0WNkLONPwv+or6zO8fHvZMV0D4+JP
OEyWH024Tsbr9ntSHpZ4pubAOs0EmuQQst4m0tLJSalp0BIH8H4t4APL6l9G
mjljULswXw3yx2XLxjoSEZmTQomJKSdCL06qXSYAHffCPYXGYdEYHWV0DvyW
7Pakm7AlPV9BfoxG/wClDYtytljOPO2JJFlYHpg8nmHF99GhyJlkLBhVAp0z
gnb6URtNZz58Ml4Tyoz/J6UqSLqSTz5Nz5+hiRP5CtS422YShFwCPWjcYdwZ
bV7XnL3pdvGU+CifaG0/ePUcrQQHmfRYNyvBjOMawonZvPpg0RO5bmjzZpbh
EtNEiGMTTxomvdXk+h1Cnuy3nQNKmmPpOI3LVyLJi4AqyNllXIlRuu5mFCbh
k/bfUm4BL+Tgf1afDAAky+4AjEeI9n38cOOGd5RkEhWc0rfCNwoiToCl9ljy
VKUMAuKEKHUTD+d65BOj/a6k+GZyMFZZdHNB9hQuhrg3mkXeSbevglz70sjF
1rU5AN9zvNOnwaQKZxBbmwCdfk2kBDRDOk6i9joq8FVdjcHCkpeJCa8tfB0W
sLyoCjfnQYZkdqBG6V9+9uyuu+zvi+pXQLNik8YOupgAYOmp0yTkGK+WO6IG
rhhstohzXJ9d4MdGa2JgqIOJzfc6lP1W3hMSrRlgjRaHCJOQPr6tGppjRPqY
sdkyARM0hV1lXr8H+X92+TVGmQ1+MSmhJ+xqijr7WKAyM0hrrb1t+POMR2Ib
OQjYHHWWC62nLQriYTFsWUTPHISouh+mfLnyDAIWbzYbhMJnziSTmD1LevIc
b8d+UmBnsSsrYqCc/XDrRDkkKJ+UG9kzcpByVKv8/VZCDeKo3H82zSa+zRll
2dD4lO6SMMq9IaESzuAOPRm5nQOCBjtOL3xnLMT9BcryE7yhBG+2ljGkk73+
3HyJ58gNBS1ds13loIBSXzpDbX4TC0RD6kiLfONRODHOlGet3aJ+WnxY+Sip
Xn8sJtuPNCuMw8PHNKpC7ZfBPi6st1ppB8f/9mIjgaoga2PkxwJgB8W8qu2P
wIJM+3oPKdq4rTIdy7c7fFh3zAtwUt23f4xp3VeUsoXBeVJNUtKhWCwI/wX2
muEtciXGosyVKbhT5T/hZDMhxww8Yim6GoMFUoSlVW7joDQLU/s5MzD6wkcI
4FILUf7RY3wU9whmL60da5ivWZ6kxu0yRUSWhAiswcH88QtVidufyb+jXruA
seBz23YIke/VjQC1QjGtvUAOKOsEmRVoZCjKi1gVty1c5ehvJPVBwLqnA+v9
1S3W6nUrNKDYV/EcgbcWajUdGYeoXKoJRgTqWFbKG081ed59lDJCy67/SlZo
jJqgj46yj+eMcaoZtQyfb35YVP33g5cbE6GQC2CE52bpKw18YFBn1HFa0Crl
Hk2peVBr8t1RxIS6ZqT0V/0nkoDPjIIYXBppnrmZJ7Bighk+RrZ9nym369aR
qaqN01Q6JPI3VmAiSH60V0NpbTl8j2NoREfToBVGsPOfh6eG9eauzDfdXglc
99o9pIMgrYzpETCgFhhWRoHfEe1V4gCJju9/0PbdCSdDgTuLHaJOTkHf/SrO
Vs0+o1uydMWDZuNQyVNpKD0j56K+SdPihZbJzy1dBsaLrNGDZNWZCR4GnlyT
hbeXQ0+7K7h0WrxKLyUDSBL+EbLQ1G0dFUvPsc2A+Hdfqfj4DrnhoH23pEej
94hvx6q9yw3+5ISgT+lGVrbnM/Bi0B0w7wQLOJ7EDdKUo1ZV40g/i3aGFDtH
4McQMNd3GnRzODM9MLiCZ12Rba0larXTlTGbXBSLpYXgrjjE9ygS4BD+/Cqd
KNKjGoP3OQlGi5RPE/Q3qQxFBsay6YJc35jhvZlCD87NNb+XdI8x/GlenwVW
+iboE4wKvJ0WICVQNzy6KMYqgV8+Cv3XczVT9uaFex5SCsoU87OtIpGb/N//
T0rKCZeNvmlLAYUA8dIXbUgHwWM8pLiEBE/uL+LsFCafxlFgqKawILWDlsWM
43UKK+eeXM/UsP4FdZTXb7ALMofzezvmILfZDCJ5f5ZtUUoyLEmj6jbtZ9mC
65lMjrVqsjGhJTVIIw9+4gGIBapNtRdVUnJ51DafiqSv5F8vS9XCu5zl7xJy
F+IDYqXHowX9/C+uurs13Q9iWFPlw2/Tl0t15sPwhWfd0TvrtcHOk2ET/XR4
WzTPpcPLR/5zVIlM0j3mhAF5pcGFpzcYFPZswSlnPM3nXTW+dfptAaL/CkT2
EMikFqCygVg4VArvy7HhFhbAWva5CvyAdXT4FXf8jhNT1O4a7gtoN/PvZvvr
dx/Yo9wHwnbCCDgUeGRIrJ2FpJ9wl94ilABHODUKLWf+BC7uv+w2H/f6sJwu
vDPHa+PWyuvhmZwgbcEhqDWQaU52RVgsENBfdJdWivDlsxAhxBZFBsPXK7cZ
vjBs0l/A2yErm9GjR9GpmQlE14akNjk6MPluQZiWcJajG5Mz3btjGxaHRNHP
dMA9zrQ8HQFgMIjcRmo4k5TZS1ydNPhVYUDGpJr0UI5LWgc1lIiH+o7Zmqpg
pEdO2/l5g+hPQv4CCMs6IHwlQliwQsKoASdWcDPUL21JuOyjggvJKwsElljg
KzSq6ZpUeGney0yY4EXDajkGC8vMiU++PvAho8uttkux6HuJa/eLxndqxsGB
2vRT806fByxqnv4zopQoUclorlM+py1RY+KMwGPXgGjB0zlTwBkLoKIv8tIQ
1y4lkRhGlxXATcIjNBH5PYZ0M+3U7NZOXCFrqD+ssyxagyhG4F7GpYXcgBMt
GwjbOjCnMvrqG1dsLmvN0+uI0HqFbE9VDjGA9uqYtlH/pMAb9KqavOaK/E+z
XrGv/IQklDco0r3rDJAmg3i+vLijWG+f7twf8LslrGqHSc+qAqkSOp2+X9xQ
J21UK/CNCmUiVFGn383ZvrCAHlOgK4d93uqm/h1xABn8HF5K+nZdgwm4GZS8
O0b8oRanXpdWn+7s51O34CG29A8LoTWGSyxDRPsfhdbKE6QqAt0wz8IZMtV5
Y17s+lcwKGfjQtTMZm5gCui+xewfvcqYO4pYI+GkZCQaum6wbZ6W/wOeJLi+
UEd6l3RdapIi2ZoQmqOBZ75+MZB3zu/m1ehA1st6lQkaV3jLX1VPA/aAXKfG
j7W/U5tAC7/XbF2w7TuhWYghGnu4C3ey6VmOmYDyn8816m+IxuRnzfdAIe8G
tFYE2dTIZsrBi1B/RQQtvzfKpfJa5P9oprYd/cTwQwbn2kYKD1LQURAx1SyY
0iIJ+3VQUNxszR+zW8T4DKbwaad0uaTqE/KaF2oQlst5arGlKHEt/Yc/KjXh
y+7OwWlgX1uRdkb/s7bfKWINBvX4KfqigUNJkTvyE5e/f2UWyG5aqLjLeXUs
pFzAINs+FBiSHQVlZPmSifRTgprO/ic+V+43+ErUfrtqKPTUyxxG5h2jrw4c
AjdnmdK8RsBbadDevi8fV3U6k1MoAqHiRXx5MDFt+/1gUsX9xm7QVN3PnIcB
pmINSecc+xqawRAp52jA8pEjLaSQRCr5bA5Q8EtwA2l2ST+iq7v3CE1Fzm0v
hrJHBvNp+EBLiUvA3++ApSaomLML2POVOqTs9004HqwbszKj0xQDaVcHSXos
rNRZ9Zzf8u4yZO/dJjx37n7Py7g4y7LcH5jbTm67GoQqRiTD44NDWY9t8JTh
khY2QcbK+zO/F+22RnJ8oj8GZWUzT/wFM0lnhIrqG4HikcFB8P3tjEak0Pld
P0eEQNcj8oY8Xmv0rSFYUXJAu+H0y/GVI1wvU/EkZLzz63dFC2E7BFVHAsLv
Ec6DspuHYGSvCL/4Yky9+2d3cXgsV+SdYLHaD775/9bt2PGdi6pOxYN7FUi9
T9ph807LpdOKQdwonXNuk1kwg97REuK8QJDj+M7j1JqzOHAtU1NRnwVtcupH
g7o4HwrgalQI5HXUkNu3PnKTi3PacfTfkGl7vGJWdMPaJuGY07BFIjekFe4x
SpiVlLvvSJLPOZ3BE6bRbLS2/3tI1XGGq9YpH9/dMZmDAPz8iOVGAN8gOKMS
b5zjGSh6X47EchkMJaL0lgRbsF2+3sseVWk5fmiZoILlgw1P50Z5DQEBUczI
VelEO3KIPyENspJ3gxvrrld1+SXOvTsXMJgA+GflFr7dRDbd4ecGUfcz8K53
uFaOFubdtFYTTvQU0qD5WjlLmw/3hrSlRBub5lYj7tLU5UC2UbErKmL3+a7j
BPiWfyhLop5EkXoSdFcSbQFM3mnQDw7ZjAyCoHTT79bt6URqYYnfERRofM6O
dtQ0EY6FhpXN4rcory19obuUZIrHb97Dlbx31Qc2QliEd4jQgS4lNkYy/1Pf
ux+iH+LDa1V75yechN/siDL25+FOtgLsO1YpjB+a/4yigvJvenZoi+FD+Wrl
BEeQoSn/xDSYn4fLnn2ZNhjkcrLYYKeX4asnlicAFE9PLBvmanlwFPkakyh3
cprtRpf0eUI6M+4Fq1UC20FuBUPX6BG0U2w+CfTGpeWeg+jN35vKikBg3ps5
KWLynD8I/ir6HDPibpbCqC6EDQw6YRuQ92ZBNN450P98Q6RP+stNFbhedLvr
oFkDJ5XsobcSp+ucwrkdZwZSFLvWMmaLYdyapU+FZQWaLSvvryoeEhXDVnxn
TPCoAeESpOur3mKyT6cq+tWQHJshi+zdHSe6YVvs4XKxyVRVov5m5EAzIin4
ZASPOvOTRNgkLpj2gJ4D7RzOCOEu9s7xTENPRJHJqqp437FBH5T+t+h97j+c
FjrfzYFw5CCyIwKm7y7SQPZXZlUTL39pWuBVx3BsgYHc9495eIR0EQKm+OVw
ki1lWo9gazA1alK1uqDLcNykLav8qqW+ja8QWYM7uBYFHt/VK/2Mh8sslIfC
voo+4Yi/CyQk4oxjTvxXpKUIxf961RZyQdwfJ8TPVP0gcDmI77AKwvGKqXer
jkszPT2oGpzht3fgWgE7n2b2vcGIgN3kdEpJpAG7F0Vo38E6NObiH6N8adNX
0dnEzk4BMWUlaxdem+/XbCzKbUcdKCmT7i8ERQdfSTZdwcA3xIg6RtBxRROx
txCrsUbMbzk/kCBL8BD33Tmcso0u6dYNEdaSyaeND1i5R27JyvZeg0R0KIJE
iP+2TGG4avGF8QatyewQ+xkTDQkgi8nP0gtlgxk1fp/b5XSrmm0wK4k4WuvH
AHEV+0NH3NQFkwDZ0kwnlLrolAGLW3OpWRmyn+jbqc7miUVAinKOW33Q+221
VBVQtxzJ/AXlHnWMQ3qz+vBllb88YNfWIR+Nu4ounhyLw/s2M0nCu89dYiUy
GERW5NFJoAST4fzkl38+GZyLuMEERLBjUajAEuNi9pszNZjU7SwAP1ry7Mtj
UbDjjDLfVFdi2c9FHxqB6IpQTrZvYwfVIhXCynD1VtRA0RRnr5ERTaTvpwwl
HGm4B5RefRux0AHLN+eZy1BrJB8C32pywa2aoUj6To7qvJpQCXJztYqNbpr7
97OAH5vtbtqwGVmGyTCxl6dZieQD97SBw1JDHC5Yn61wNzzeuDli3UwIQ00l
0g3Grm0zrSTZ/Xtgn1jgyN0qBfXDn7CKkEcTJH+ZnKLTp9+VfK4andJueKVA
PUWSzkPQp0NbmUFKGGQoXUv/AfXpZQzMFOv9M7TIWitC+5F9ADK54eDsNtCy
vcrrGI18+8ctcauXwXgO6P8AKyYvakr0R0KaT8Nz64g1riTOB+1Dwj497o17
JdouJyPHNtkJK809wwZX3cBpZ87G8q6yXUcNQYPSK74jEO1eAjJ+Qans68wY
na/L1Q+mKbD7rvYcX3XuzSan0dK7JL6avTj7P0aZnVSoaxkxjeGMBIh/pY7y
GLUFEcilrykAkpKbxbfvgEprOQMQJW7/XPYk0p6uzni8GNfKPZmCOqNuKJrD
3loK1n5c3Jb4LBlLYPZ9YQeGs4kuUmTuztNcILqCOWq56xfvGKPZoqmsbwB+
LOqqr4RT1elqQ6zzso/i2aoVzEwRbc3ecFJppaZCFZuYcnj09MuNiGMzUps9
IVne0HKZbko9OVjXoOzOiV7FqHUDcB9F2OVW4Dp496AfMRHECegx9myNv4O3
E0lPdCOq5IcBWFSUbJJeNDurgVGWiK9HFd3J2Lg20GPU53DPx6U/1jG3KLfA
PwIEmkA7veI/5okTaqGJPIOtfuYMoZFSY8IgqWNCT/K3jW0jvxF16Zas1gxU
ZqJolTBfEN3NmblTQ3Dla8ue9RjeEzQXv14ngrMPZXjgzVsSiPh86qLNIBlL
rsV1dgxLTip7VHCWTiwn7+FWoAbjONC14OkpPHZVESME27se2Y9h3rAMMiF9
9yaBO0K5p35R3gW5NMRJTXWaeYiOrHg8EdN3oQyucko3m6NOQ2hLde5yGtB5
tagqs81PwPuAHi8HyJExQMqUaMnSr4Ke9+ex9dbbVlC0Fj6+CS1rxtPzlhUQ
GMHOf9PqedehgRsXu1wl8LWnaz4iKpY4j+RAeRlCmZfjpGxU3yKzVC0NQQwV
E5pSKmNgCakWmto6/aLSrp7O6QJsT2lcdsstR0Fdnlv37f0R9gLdDCqYT5oC
N4naohEKEUG1hs7cx47XLb5oRm6771QLg/35k1vtz6JtzkmFQ3htr59pWVSu
uAMX91zsw8zN5ZUnBIz0aRIYK2sTrWcxS2He40ja7fFHt1lhHCwDTObOo1ER
IvAMfuKih41ZfJc/xi45g3M8DZ9jqvfyukNtYh9QJCCKciFOSEfFEupnyjOj
upa1rfvDjU+L0806iYz88vbzrexYPtOcdb2BPLoSHU3R06rmztyWE9B5dh0r
tj+yfIW9cPuAN/VDRxzKz1hYhtWr9j2DVMgFU6VWd7a5YbrR6SfQYsufCZKT
hgL6QjuojR35hoFPkonxH2+p3C7uD//oJJo1P3Ssh2wEkhnWZLhwzrpiCKfW
zaN7uvRmwkKf7DAUpYWUZlbGQVvtYKydtM2OdcfwK6VEg/L2bEEwmWvOLjhq
4RUuKpZki9r89quJSfAnCxi5+ly3A/4YMxT3M9vLphiTuapknY08JkekERgo
qT7/eztkrdB1HurX/EOEQZ4lsshVBA+lbNXxPx5vN35cFm+K7gA2NBQp3tmh
AcP0bQTsp1kKjR72Wmy+bNI1AekKJ/MqNXyxMuaI1I2FsPOQowsPU/bb8nO+
aJT46HeJdpxds9c5gWhPr7KLJxXnf4Z/OnKB4vnwysICQU325CRW9n5L8kEB
e6WYlMi2qvRk5hEELWVcIpZdPXbFlkwmtPgLotlZTnYFzILcPoPuiyCgIwqG
lH0rjtyXmfRyp+ulJGSzSnnNqbFLlUd+mxLDBQxsxTC3/sCtWuYhFpUFD5K4
OQDEhKXvD9cvj63+7sCQSNBK+H+B3ujcdcgnxictOXqQqZlRxoC+ZYrnx0eA
XTbo+ELjklVxGvsHIGUuCvsula5GMW1guYmO40tVgbwCG/slRcFZ6pDXbawa
iLfIctqCrYZcu1ftHsS7hzkCD+IBdS7RoMsZ71ULw50lp4Na0Dom3D/mFmiW
IgyHtR+VYZQLsuBO9/MF4EsIS+/pF0YWz0QP5MVf19cfbB4DEyIC2YxTdGmP
CTmP4fubrLqS5aPOi6G74PO91KHIZJclcQEB/5gz03AdK4/lwnoHNRFHJScP
qBi7s0j5JxWeqWFTnItnpaOkxaHbGyWMm0c59nsTrvhG7ftL+4qdLDjoR23P
Wsxb8fzuNTDhwVUHC/BRnTP+dL01NqHqYIr/LbMgh3W1ukLS3Ht9OIY8dfDq
DaAULC6lKRO+F7KRC9W1CrhNvMHtt4R0ES3OKoY3EKTRgmrb1hLDiTNJkgdc
hCYs39iU47NHof3TdBt/IaEKbzYLXIA2gcIJbEQ2DSiSCghDJ9e8HU5kFrp9
0gZLN8DBT89K6VKAyNfwlIxEa5OpGNEM1YJybOUPrmR+S+2Bjgv1wtDgywp5
LjuXpLCvZnlJdzKGU7g934CKQz4g47Z1S6alyhxhsLuAaag+IAYElPbjgu9p
cLjG9ucIDbESNAVrbdcVKxmczgQwYe++xog5F99QAp8mz/Q2Z0O2/wmRawm8
v8Duyu2m0ZzgcJBLwKJtYsVYPOEVW6D8N0u5JZQ66jJQ8El6J2+Bkd1yMkxY
/yJD9Z7bbvWx/a0x89Jgh+5uO0tNgY8vAPlcZypPpXGFVfkDbktitQ5UTPA6
IuxqOtTTNLa7WSGxoTV60AF3nROBneJ+lLW7WtqVLhYDtQaW+9/zp3vcXMJP
Rg94rgGCDGDNYD9qI+GGPaSTkrK6FNdM06KJF294OCsWqsmtx3u5ypSKOIwY
aZP30Pxa9RN1bL097LxG8qwD4b62DwM/ytmDvcm7lDhyZS4gHYvVpU3V16GO
pIYEqCYwEtLvhBufv3tPoriPVPLjLJtD5zPxfx3vY8iy5KkW8+cv2E7leroS
AP5JD84/jPur/WpWko7V4Y4nXQUAnicNiqOv4NnyF5mXjiO//lu3S97SJiyK
BPt3qXQ742MLHreB/5fExCR0KqMIR51GfDHGUBd22tTpKkIOHmUfDqr1ZFAw
9fgzrJOHd2Z6DWVm47gZSYbeFn0FWd/rYqMcJ5wPc3XMODMU+sQzye/6mrJE
L0UFV1gKmMQhDDq1ha31SrmrR9xah2+yDz7Gu4zqrQLdpC3k1KZpXuTtH1O+
PzD6ubFwusezRSYeoVa+YhHBTw9tUvJu8BScAlTg10h6eWxh3CQUQjB8nsIh
NRYfY1cYWDcAExsFXHWRKp2o14ukQoEBVHRQe3veu5wU9So9XxHmiJmbNohs
t8T88tUUVZWee9MGJ0fz5a7sf+01G+TSeNv0Z5abZy3rAwOZJpHCIGgayuY/
q6nDGW2lI9vbe5xGLeGXcNB9eKf6U0uvkcBu5wJRxdAYAKqCMh2kZtGmhYpQ
l5Y+545vMZdbPcyro/hX29t35gMBMFKBqkduEzpkOt9NJB7yvbstpfhBVqgn
uT2fh+wwOYkQ2Q2b/sF7L5q+Q/7TzkJrdo/v1AX/xPm82N+HTF32reB+gqjB
WaET1SjfD/diQWZzyvJS0f8bXyV028pWvEqIVVutGuzA69uMGAFYtBpXPQea
QP8R9ayITB67C8kBe1TzcyQ9pDd3sS3G1TzawRJWnz2SZOFv4AqJswpei/rv
xHK/ChyBsEVwbo/uESsOxFxwrsWL/yHBS3T/fKKjbD6W8jWfrI9LtYvn+Wrs
cIsLP3tv4OCBMYXyRtGcp8Jj4duuYnlUZb8YbhYhDfirY3Gx3YarGzWTDJji
Gw2Naph7l2c1Fu7XKzxOD0QMfxzrUGeWDpEDKwcN4xWgPMSH0ZM8XtaZgcZJ
J4x00nbZRBLgE24I8pXBBHj+fN3s2UPYp47u1GjbCvGsyDVyYqNOp+LGISVF
no6YcbZ1indRFc36zxgdrnfrgT7octGs0WFeTBRuJfqjKliiP6w55ylOCF2t
E/Q8LFcuaf0uR6H76TNirGYQmkHKbxw45w6HCReChTuFlk07ii5jszEu0aL5
VhwG23WyEa8LCLDNpdTS28NFbkXtNykYuWMkObq9E/6QYwZMhbZbxR9vCEWT
3fUpBmXb1st7j85Le5ofMm1KVzxSW/qIkYNu2gWu8MjIm7n9cL7NzR5GA5YY
8Pi36ek3qCL4oXJd77/PHlvURnQfCqZPajwM1EmxZKE8Jm/6HmQbWtouHW0K
PCcaUIVJrg/WXKLO9AS0gbwf651JIppDMT/hNEdpukmepkLX9BMlHAO1lN9Q
KLhcTU5+fVRlMpEevogcDyt0DxMqXlAfTy+1ennaFjNnESuyHfMy5CSIlrA9
Vn2Yo6ntuMdNtVoD4p7aSU5oSt8ZsLF+zHSkyh/g4xpq53BlnMJu18EBavol
7plXQewXXiLjQRGfCFlrs2sXAu3Y1K+EijltRtkUrmZopBdepp4rRrgH1fbN
Li1tDdk46wTohYsylAsr2XqS8VIAJsbcy7Ghxku/xTkK/D4MLfMSyMB9X67Q
rQxVUKdKPmfJF0H5MsfnlRWLEc8bU70mopd3TwYN0H6v+0iDV+0oCDG4MeuM
vAIQX3BNGdL8heZMWe71t4iLAbxCykPoNE40TcukOGaqVt3yUO200cPLVmIU
Is/h7baPdngiOiON5b9vGzPB6v2YM+zhHyylcui6cF7gxtXBtOo7kkix52KA
r88jXzMn7ZMd0ShoEB28SXwmDvOkxgkfNA/QztMs6bmE+jMBJ/r8iXfZ9ijm
XpzqJZFaRq3GcWSlg5+WUGSJClicg4T+iaXyBhJ+BbermE2x3d18QovJQwwy
Q2c/qHEBEXxbjt3zIE9ifgepd0f3DPaKVK/dxujKT3HwSJ4+QquA/6HZe28v
Nu+wBaDtwNIPYhW7wJvn7jIzgdF8jrn0S0QF9sCV5HKu3AG7fo6IsOI3XjeP
rBoP6hzpVzJtqbXAnS0otPT5MiodJmF/P5ewaw3tJHN4bdfapt2uKWXKWF8N
6V2DwLS3+r2jaXsWIUbBIxcfrOcWKmr2qkaXrwdPZSgGyNz9P4s6ZH/1K07O
T5W/CcpZQd8fW8cmtAgJ8WuPkLljZlwUcexovYM3/jZDMc/RO/Xd8ZaIF2KB
NAKtd8mcehPABltgKfEHqUnvyCDgi3pRFbF9c6JBWg2+26T+2WSrVCSICeVb
VWfaGnejHEahf1T84MGsF8sdLKQkye5WICkXtc2/tyTzsd7iYzAF5j/NMnfP
4kP+v11mwlaubomA+Ks1ogPxgI75ZkYJltLqX/xalIbGJ1yfZuZJnS3QkSHi
RWaemn+wI1DGjA0yyH0C10UFqLhMboHGrkoySigsHcuTsk3GPJ6FEhpL2HmN
QKhzK5qSEqkvlAZgmvqh3Mz+H7OVLt7RXDTvRXVFM22H+mCHeDCBplW5EnBi
/STUXXBhwPLl9bzri85kl5W1tKm45sHf6lSoUWqDZfHZu62R4g+D983Zi4lB
uS0GTvNW6wqZm2iOMzX3+O+lo6Gnzv5dysu7uYbaRxR/hqkumeo010QhKw2Z
aAUhE7zAMrjRkXusUYUG65hSllKIyJFslu67oGF/RRUKu1bMhyX0GE/vDa0X
FZ/8322Zo2I9VdwZPcR8VRU8sAQroQp1DDHj4Pt7ohXM57/+F5Ej8tL85r93
N9heaNjUXXcf5wohFj5xBz61R2By2TyRBb3TQmP35gJSW/ssLVzBUAwF70dt
6UvwA/GjnYaWDy4RSjjQ5Jcpsy42ZFM8ZKn37cYJiWt3DAxq0lk0WQPYKsiX
sZerNFe37Ei/TAhK6OY6xcp0qQZlnYnxubEOeN3BL/PQzCNOVTpIaV2fJs10
W1XQZhFBZJw81XRsxOdCGTQ1Y/jxDjqVatp7d58Sn8mmRLlcWrNJDsA+vS84
DwYx6qdELFRGFt8OThyuW2vGY8sv65X+QqkdZOEBA9TH91rPhZZdCpv9O7f5
6hip5b8TLJBn8XAoxPekhPcOvvhp7u/PcjW3HH9SnMRkGSHV0QhJTE5Xspga
tYpscxnM/vsNJ8oSHNzwgsJ9f0dPPtAf1LBk9lwwi5O8EfdH2CjAwJiRZVAH
G0WAp1Vg88BOpjLfqcFsSBqmrP5D8Cuv2M8DH1a1m+JWbWy8Bu/o4lyyatfD
uECMErnsa2/Q7Tx5EiipszoziEZ5vdRY1KgT3/cywyNpKx3ZkBGBMNAKbtPt
Mjgn9gSuDV2vbvghjeHPzFNTjnRejj91Z6TSXQdbH9xYq6ymzExoW6w6XqWD
gR3a9Eyx9/l5uWKnx/gWBH+wEgHPUqf2kIuJ7hTUusp4z04W5qRhcVBzEiZm
CpNlHM2iibywgCvWld1rWmUBR7835Fs7kVfsa7xeTc3+JTiD4CzBjDFn0VNL
a1i7u+xJIwZFTcd/sl+x/GFd5dAjVtlvBVwZejfdPqigpCqGGhhW+nZBESkg
L299x4MF9j4/Q8Z3wTU75K1LO1Ds6eD11rwhr89MdvD7mfwmiYSPk62zUzTA
BBLuAFHa3gjYAXZp5rf5NEGvo5j+p4VPYSazJd1s3SrRvFQAe0uJPhm0EFVb
jt//rcvNRpgA2JyTOlRk5v39kkupiemFBM7GkNG1HObHuhgpLLaIpDvOTUaQ
6Zjmg7x8sepa4zpdmLz4NReJo6NoQOCa1OBq9Lc2txhxIJ10O/8nkVcE8oBK
kOZwUKXqEhUucAz8RSCJFlqf5bcxLaFBoSPuOFbzsPE2hWPsInOrsPTPAmpI
Z5MBxrF9MSApah/ePe2FLMi+t3pe03F4QUkCOfoZVVgVcl68kF/y8868fGeh
fkOq91OUndfb1c8Ag6ZOJ+KWlDvybHSzmsxOjQ89GaIQlqPwHb4mU/NCjetV
ZKEgxkzu/jibKPSpZrbBXCtB+oLE8pwtBciWHT7q5DJBfs68WqWvUWeRFPeC
y9qtz9vknxtkw4QYyVZLvy9y+xY74FH0nHAIHaBFzjtHt4LVTvZ5DlR4+t6j
l307Ln2HKfiSn07jH0fxXAty1HrzlyUGSHvrO0XLEgDZZAHUfDUjCXERB+9L
2wlIGNwsvuH1hni6nY6EE3dymW59DA+BVPCvAHEWhV95Lfg5y6uJAUoK26EM
mtoiuZX6t27fKjPri+hJ4VESKt3mEdQjFi2lHBnoK2KhN9kTo5HEtfFXBBaL
9dMl5q5IJXvhR1bbfuNM03d8URciCASayCd4a4FLLpXjEU2rsjIkvrc2kcM0
YFAeEJMX6pgQobBGN/5i/6HkC2A5FCI8/KAgkxaDA3LqR01XKd2t/VDW5vyw
ODfiUZoW7s4rTvv9WGDjOfzB1lvc57aLKMmS98MmWpoSolR5KkKyhlLu+ivw
LnDDl6LPyO/m91UGLoy9p7/dtDfQAodRaB7vIqoevtnubViOr0fg+ZvFAVTi
hHBVoK7m0YqUUFBChTykNOMDulFj+4gqpvqff31cTbaCmhnvhrfvGRAW2GBM
mQfZ+ZNd+OZW9J5RpasZW1DA0Synvr1AgHMm0mLqhcRgh+n6FYxME7ourDYS
iJj9c+6cc0s06y8UJL/yisADo8eM1NQxXw17j8cZrW5OeyKokCAxO0USp50o
ya9GsBzKQrIaRBHmcQZF8J4tJCj2RuRSnSiNpStCGUAateg8w1xJ/sYq+M4N
SDOSBlixVO2MTUGOHMY54TMHJA6IsBcQeQKTljsRxNXNQqAFaBAQWWpqiK21
UkbjTAnSeiBocjwuiInl8A2zfEwCI+rm5qLHv8ixKROsvmBKVTaKYd4z8zxe
Icu8hvi2gDySfOPHvMVpUvho0/6GfcCueXffplmZ5UuHtbDhlYNQpZE+QsK9
VH/oFIk9CHlhmpClOBbbXShbNvMT1D03w/oW6N78PrwTVnWhTBEJMR49p3tM
jKIQROPMieUOTTkT98aQbFB5xurbEwQkCD0UCwT7waJaE34p20OBlekrtVph
aqAy91LqBATzq/fSBdKXgwQkhG7oRD5VgkWAcJOe+rNpfjYRA5DC+oFMTZkc
5tVv5cd1RdMPAMFTn52A8dpt0pxY8PbTDS5rMoCMKL7P3xWiqzMzClrQuY0G
7AAwk8hY53tpiyVOcwP5hDNpXdu5D+95bZrSHS4g4xXSZ1girIaP8tTXEeIJ
UT7VCW7kC7YwtdYmCbxcuOxwvyfTx8lR2q86TelAbmUaSxUZ1MF9tdl33uf7
TlQCEo+5yRBn/S55zx9kCHWG6Rd8mwA08nzCHPgDz2Ti/zwOH/Uw5H+83UV6
T0mdbYC63xtu5pwCSdVtKnsj4jComq+lETJ5erPw8M1R6ndIeGV1YLfdB1VI
B5LoskFBgCYUSzK92eGy9Ts5qmtbfFZDksgFf7wyBkMfYCpuNpIaH6c2+zPd
iSBVFMVs34NZyQER/eB4vFjqS18pAiLHnNbayfHNtM7WdB1cqFmWLfMe5eoL
vsy/yuqGDWWMzffkYogpbAJeEOVoCM6FRC6rDQjr+2TQSPXii5BZRsoGA8g6
GmcWIl5ufsGI9sYZykT6d0me3Iw32Vdp5emFPyFq4N9lOCP6XPUZn+FkJOaf
lzoDJy1QNhsej1m4c1TzThnZSe3vFNMH93h+PPfIXNcnQENUVKqmjSF8gzJO
EphSZEjVcbRnB+wL0BnZdSnjZcchlokHYdoZ0R0zCHryiSX5iayD3HlOUN/r
R2NJcmk07+4a+VIwWMgnb8MDRSMnGlykX0kMnyczCY2ST4bEc1ZJRlJmD/s6
2H4SRWdzsoQ4UXmm4GQenNZVGtvQDYdZZLFom1FhEDNsWhT97zVoxJ2ugAOK
v67V8iGZPEce9PNWJ0YyWTkPz3c8AQHAnsSURJHR+op7g3ZtYVfmo7tHSwpf
2vRA4sLbiImTX3jI07J0bKIwqiHBQeXgyVDbJF0WKJFWxO4L4QtFC7iiiuJi
LKxjbxlWI2iWlrJe7NKclZkJEBGfOi1As4+81qHG6tM/797fNmVe6lM6WPae
Rwe9P4cjtkIz/a/4CEWv9NyK9tIt4kSgNr1/4j9fmi/8QuieGDFrAOT23FDb
nhBD04RTkZG8tzRwpktYFvzV3ADxlw9qMWqiwmwpN67g3US31CvVCKdN7Z6C
2LBt+rbcy71aMJukv3ixitXzhhF943HiB/mZB1HxIwY7RkPXjxbbHIVo1XGA
b1lZPq2XvCScnFSir9fKGTO1TS3GKfe+AuRShzB0XOlazaSVmS5Gpbo6XUxa
8BWwCMfe2DOLIM0AXgaVmrl4j2LgB9FNXOpWGYRxkWg6u2PpGNaUui7dEZb7
JsDQCAN6rQVDJRp/LJuM0mmRYPLdjcbCdRfPzuGVfrtLMIX+cLldG8d69Vl+
AsW/Xf4ZS3gZvpCYhQDTf+f1CCPkmXPBK2o8NvhYSe4WDioSpvroMF4ji5Y/
mGKmsQOCNn656b8zKYVEuaj8zn5zZwSEEb6hehhcyzotscRkWOfNM5zy0fvo
wl/V0af3k6pg48vHnxrUq2cL92Ssu9JBT5ZFQsR5SogwaiV3Nb1ZB8e2UfhB
pBb6tTIq0Vz7Ucmi0m6ZkPROJNpdE0ACNPm3/EC2nxXO7nxfPB0IqSEzdxvf
Qyo9NLhNANJf8HnNhf+2zDEUzIyLGIjCJTVJL2cnpfFQ1t24T2mHuY+rxPgH
/TbPHEubL7caz2oSMZIyPwYDNfNh7MuTKruMW80232e+bdMQWuTiwvPpcs7V
N4cwrDP3tW3/tA2K8SMXxgyQeHFBgBYLagFUR4HxgPEAcCo3rjA3c22WKzpu
VvCFDKMcbYd4Vr++Kfb5/yNjgoRrE5MkaS0I13rn2LVT2JfAy/Sy1dliZYYu
z+tGWUSXYEQYy2BRrjMCFys9N6P6AkPYstBZ0cGAlc3gSQg/UgljdTDY1crN
4XtoyVLd5QN9wxPjWGr7CIRPrEZWk7iYbbaklf1gKRyPyjIiqpnKZ9lXXWrQ
vUYqz0d5RbHe4QSGQGB7ywfnq1pq/xJijv1NYX//FwYXQEp5f10LT3CE7CQF
iWbj7m5xmGYe8mMHTQwdWzhjfFS/bO/ROgUY1l0cIL0AEeoA/6GGff1PWzaK
fTmNrAU+JEI1DbIDdL7s1EniKvKGqrbitRRe73FxVdCFcCVLpMQHGafZD2TP
KSIQXpz61X7qiqLvMFunr6QWOOjJPPUepDznFo9AbdvfuvXbg+803WV7Z1IO
Jxuw7EQKraP+18L2YkPP3vTbG6EZXWiyTdkVZjJbR3R0bjLAPdTTyqBRd7xb
cGZtU0RnkTi7ahfgfmtCkEErAKg1R6h8PxoOBWio5cliOyt5CWYjtBIIgLti
KPSsRISoludfBCjXZGkhlZgutLkVT0GZdPTfUVWIfNLdUqqRtZKMg5udJlM1
VyHtGeKhqgJos5DgBuOpQ21p1LKDhj2zWB6fJF4W1KsP7Xd9Qwnmc8+fyaKM
/C2hqJs7F4d7Cf0lLyWKCnJqtTBiOBmitLyPaKnOmKIQ6ymIYatQAfNaBlcB
uQOEdi1m7AV9rSjB1I4vk9Nr2iq1AbgXlTG3gMXwpYd8tcEp38a+uXDsEavx
NCvo1njyybpKHFZkUqasdTfWDMnA+eGtvNXMm8ry69BHGYjMbvKoHUFUUinH
GdXqgFLbeDeBY6njFhsSIV/1lG5yyUare+OmRg8rXHI5jb6IToTF6NVSEUC5
mHQnQU9KLPe4hVd9XxAT+rXH1r3IwhtwOqmkmO0k6osevbx1S/JNTaz+Mnts
/yM2mMNBwz1Wzud3bG4TqD91TCa0Tu1FxITfo7RRCDDuEl2C6vmB1E4a1uky
sJODJx/0KXYRpB1fYW+ATd0JgVENXLDgpRUHA1QFlHd90vVcpKFF9PmVl451
BQDO3QRXUIVrLYr8KHg4Wz0gAaOXKUMzp2Da6aLW6ANi3oIg87WB6I/RXgxo
5QPRF9v4XeYzYZxkidQRLLvorcijrtBCiHrj73P9yM0RoMB8fp7XfeA579Gd
pJHypqkr5xsQLy3VyR7fMhKNeKH9tSZG4kreEXF8jVp/WlDMpacd2AlGIxxf
yq6xX8zsRRgHxoojIZ0YprG8sxMd6rVv25ozj7G4Q25pnG22/EYKluH57s4J
A/JQJobO0yd3UHvlbRyogNi1S2gYpjtg3p3AxMMOcJw08LQMA/UWsds3J0mn
apEi5lO21nQ4RW7D2eC/Dy1yIqhN+OUJkY26mIxYUlTwj9JQb0rfbrw30QzK
B48midgevCP2mueF89/JSVRrTgrfRsh+0eq7ZCkk9g9diDx5y8jtCJtTCd4t
zPmjNcja+hgpvt38Fesla/G2D5ngmU0qNsQliVUjPiZ1fKWFhGXSDa5jlGWy
/VTTHktsoGDA7KChcIsWLC3VIZNDmBck3D+Wn+LDkCPVQLscuKyYAfKmwNKi
4kGpMXhyvBJ3izTktpsBouCgcqFqmBDo8/LPaKBZ9G2BDOBYuPU5rdw7+nHr
Yuilb4VBNeLAV4tRLifkhBtmZc58ES+ouR4Anqn9eCXiPxb9oVDP+NBRqION
iiAId09ZhqretyntqHMp8lynG22ThKXZ4FadtG/hOV2jBzhsyl5zFjm5k06+
vcAw/+jHpv1vAmfLSNvqPVtRFlCe/U1GmX9fwnIvdSQpfuSXg4T9MyXoV+xa
2yoHzhK+KhelTF/9+DgjccCa78B7kD82LZzUujPT1gdhJxWEcbJYvQbwGoRI
kbZXWa0WVcoDZ6CavfblrcDmby5w6qVf8o66fght8RO+tOVfSwn239r7rBKU
WOud9SFeOAj2A/iIzaIJbAN1mmT5SASltJyoucBlz8IyfA9z/ifiNSQC3zdJ
pSmPU9/1Vt+mVplMCZipvxItkJRg7+N3FEiX5zS2WHXKsBxL2InmtM7XA8AM
ATpS8a0qKPzwXIBg7HTSXA1uT+m8a6H5qSFD2QSsRKNr2kl1bYy6AWKGkthf
MQI3WBXjOOy2yZlzZC5TpVrrR5GMMUSiHw1sqBvyNGCoWOav4u6o/5I1T9Lk
l9htDggDZcBBz7tZa7i9t2gjEJO91DjoxvAVPZYFE01H6Hu256fHvm/YoGj8
zyYWfRMuK+gnlEGgBo+deKKn7dPuMddKYSVDpfLcL9lF3yUMN5aa5Rk83Hje
qdq1cq8q+wbsbHQiAvw+0Rc6rLPOCeiMWZ7UR45+iGNa8FhNtGAQabn4SAyl
CfCKgaBkAM5kGNB836HoCmTOUc+3BgeqyvozFUrGsa9iucr9i4tsL+o4UdSA
Y9wnC+A/eeBCAng7PDoryuZA0M9zWP38IJeYR1LHeflJ2rXFcjWHBcRjiZRH
rXdm9UZcOQArLw0BgpdG1x+tQcEvzQVR2t9LWwy6SrVxLhNELiCGQ5b1gOMM
iD/7P+85XyvNpnL75i+ii1LxfL9Tyvr5xBZ6Dbynks6dZIRVj7hLPM4LNilJ
gXexPcrCAr93Ug4saNaurz8q7k8V6mn2CGb2Gq3t8dCkBG6NI6N3bHUkwsfs
N2FaBK2I8hgUsFJoXN/SNW9BzPFVkPhh/wP8eaq5UCotfHz0lFrMBuf53tcK
k2GaVepA6PFzrUxn87BRXtTmgnS+QxeWqoUPc4IuH5Dm2qJIkvjxdF7hjsSi
pZDbhuYKqi21/QLWvEVh6JwdXQBi9FeF0ji2wUyrQhVQKAh7SSA94lt3LGKm
ONSK+YRQ8DzHgtSqVQ+qNOJ27+1XcW+iOHwqCplkpa+Os+mIcjvPhYR6lHDN
eyS9siu2fcY9vz19iWUXiprs3hhCvMztW7n/VBAqon+L9CQLMJaZuwNF7jy7
Wj2bMuOMQB6ux0cgrxODcw2Cp7wOYD7Fk/HCBs7K4LC3uIZF366oqWQIIv9w
sVPV3uJbfqXcDMKNubZGplwlLZbnAS7ljwtJhXCsNm+NzyIESRu5uJpio1lu
uNFaNl8TSvjd1sS6iMFSEQRuIW6H4JOe4I8fEWSn2QHmSaGN9xMSDXeLIFXo
lFhUOg6g9yHQViny3EnDuKnQpEdCCIEJgn6eYpVRKPzId31vyo6T2P7bAdoU
6SJA3DzTKECPVFrHJTs8xkWw/D2KpGwxlqilAGbEYnpYj1ssDUGwFiwmbmoq
GOlEbC4BT1NhwsnlnzzZ+GQ81kvZ6VR4AKs2dA6j+BsZ9rBOtB2HxCOBui0Y
5oy+9+Bsb3BfC1qU/XBC9W40BcBSLhY7iYD968V1W0R6Si9VyivEwNc2FHYn
ds41Q4/W2envplSGsIEZk5bbudT3yd9lYaT7d6vgRC8ttOkGExl2K1tktFns
Gc3d0B9vKvmC8ncvPzE7vZJ/5mglYMVTOcQHQze0nUxzEqxhm/4TWsT2vtuQ
mNqO+Nxy8Q7ARjiP5Fy/NOpaz0ZGxFxLepRpn6SlXoCcP54r9293A8ElpKHJ
sb+4D1NG1O4+Q2hv4TXByRAIGW222QV88GPpAUQhl3CbCE69lDskg2JIGIpG
ECofV1qkvH85a2cniwEVgC78/W5Qaea8J/FjrRPUfYMCf9gR50ssO2/s5vQI
4sTB9LkIXKbe+9Mcpgs+XqbABErutXwWa/XD6ItBvHzZM01UkYU1KNBOrZaZ
8FgKzrE9YYVjJVNe6iitxCzar36PKVZgNOSqpuj/6nWm5t7sWlh6f0AiN47X
ajOLgUPdtvdPsSMDxZOMZfcJxG6lh6lqWyjwr3zAvcjmNhCdwuZWVXDUGk/J
mIqkPr6P6xufImD1nWtftlrtbqTYT2j3n5FSOYnQPp/M25Ej3mYZWHBLdnip
94VSp0vVkVuYrmkkEP6XH/alQ29Dn350Zmeh74Ccv/M8qt5bqym1NPUqctdg
Hmk4b2XdSgTh85HYwtFYTeVkCYSNmfMBL+WoBiV+zxUDHz/McHDbIo5U+4u0
jDKwvjrd7n462/bKtANaXWpmbpj+Td3IF1bn/CzGhigO8vUlJYMYozTqI1g4
+uDm/QiCdfmsGbfGa/lVz26DIaij76Lk3STw/2fXMb/uio9KdEFuq3Cbv24+
4+ophdRv+3fGN3puS4Bw3J0hGzsPSDLVnx6mOecvb1MbHsFcTGIcKOzAc1Ly
rR5+lYhABtAPdCuQXUPhIHruX2bNk2MTj2WtGB2WujFUNkzg1+ULgqjCpUYQ
2etQhx0+BpcdaaajGekfG3xzcv0xsXAF6hf5S92FEh+C5nbSTkbmkUNXVHYa
V9k/bqu3KEEdpZ85u35Kgu75erhQZGzZWzmwT2EaH4Apqx8WTLoeIv3tAm5N
Ae/3GAJD/KWxW6yQGtP5n3Cuy3wtzL218IjEZE60rSjCY8AnFC0WNr6dPr6X
tRgihL9PIQ6z23afITzv6wLCoFhzgiL48np6KcqdQR1IkT4fzIZhCk77sLMU
Q89YsW4RoH0obSajzhZBwm7g2WmM205zlrtC5hhFdzAkA0Fx11djnJVfYahB
+ahCwdZpOqL6or7y/bmB8F3gkJFeZsogTmHh9bIt5w5p71x9KrvprpONA65M
SoQEiQWicsd4coS8HFggag8kiweTTelpuO52CN6M5UyrZ7hbLMcBS8D0scBo
BynHbRyOPMIGDKz2CTUaoOaMipD6yC7Agd3ZMYyTnl0t2WOzb/GqvjOcP1eW
1C4ALWMiL0QBkAXnTyBovKyaPFpuapDnQ4FdqcnxLTSExvkJeEKJFoIFPgqb
d5hxtIRpL+hrWgKYRE5ZutkVwb4Ro/v2YvRsxeQ2eoHIWnJRbBE1SL+3tlz5
40QDiUbeVGFF8bhIjJQL+OMQb+mTkMOHvilA6Hb3xnGJ1omwG2tDuqayIGhH
AFfbBSFWL+YIs0geEu2Lh7qNHr/+kBmeOrzLow5uAtef5im+xMF9gQjrRR7A
rpQ/tmecur8jaK4KrdMZONg2kzjUAdxohSsRdwKqOsT3pWrmg/hxj2NXavxk
jL/zHZxnXGkfI3J8Tss3TnslZbmrknfuAjU1WqlcTjXNABpzDHrTJe0JQRXv
GVfOKNrXwV4SNbtqvZUNSdxdIJ44wmJ/a95aUl8zT9yIvXUep/R5L4FUYei/
/tWP1CmfT8290jJDGVDMzK1j5bo9Jmwk948XjTBcJ+l8qqy5EhOQHI2YJMzG
JVCZLPKWCvrKnGhlCuF+4O8+z1wJTfrpmy4IOIla6cXC8gmdNH+3RazhflsD
HHeB8ccPjcBNi84Pf06AUa0j3/rfRqI3lB8EM+0GO+namobuHXIPH0CQKSzY
btE52pgNpWm5xquYR9B6OLKeTUC8Mn2AQhInC71A5WX+Lz/axW5j+MRmRgo8
G67rbv6NXMUofVHUuTgPtI4x0llhBFfWE61A3KRWCgRPP760TkDN1tE8Zg3l
6zrTvNJJxpZ29xAEgHQT51NTB1Wcjk9iQiaid6Dn/xdVNYCjNnlIFandG0Yn
AIleSG7niWoAyu1l3vSPxvLATb/sg86brfACleLCfyYFbeVn9D3FgPsBYPRl
o4NFXQSc7EefaN8cRfPYQREZYA6hB/EGA/1SHpTqMIfo09YiewLKjz8fyBmV
kdSOAm34PPLO8Mq6pQt+3fcTQU5hEt32Dgia2N8APZdBAiBWB1ASfCwVgoWd
EsJE3KDpFi8yAiwij0EfjqCbii4r5nuAvzmGaZ5Trgmx8Yf3vV1AQMQ21/Le
qjDx1QOsOMVRXjXFuSornic7Dt0PdzhXkkJCRTfLHmKl02h3NU2grnArZjDZ
P6v9TNtfg/uxX/uDfTltIKFut8ZA3ZxdgzCK25MjawFYvoGkMTG9pjkQT61x
OiwMUtgrQgfixIpZD7kTCJXX1lB6TqeCxi+F3rj+fG0TxiYxfaNQE3l86MkQ
dxgarnCEoqy167hdLwTkE5Ce3Nnqeo8WLBU8+wcrz8CM9HJvZ+kNSRVAoWnG
1r7y5WlnsR5Qe9AT3v0UzEg5x+kfb7CQ1tiPk799VJq8JbxN09+vuQirv1ky
Dzh+m8Xuw4AyiramrgEshK1EZlieRkN5PlCjW6onkwllsLJ6qwcTddzrf5+f
Z8aKBcbDAA6EzvWiNrARSvWEux/UcT/ck9rGWkGt6nAF8co2wca75D8AUCQl
Mwc6B91cSaiRn8np1HovGk176YbUj3HdCaO+Q6mvCbE1jDxnx/s1E0X4V/Vm
6W1zfrNPGH3lu52RtuWcxNQbIIE8yqZACPTKO24W7SkGltcbPII6liVMZD+p
tkzUkpVLXNk5fG+JpAFqW9S6Az6+tYYqGh6qgVememHLz4IqSzn//qggTUd1
McAW1hYO+QGkk5alK2vQkCPl5m3LqoC/2EpOqBgtj9244R5fNUY3zZSxG8Rr
u2JCAdA2f3at8KZxumfPIUI2xSDoaY/J1i4azjHFt3KDE1RC8u1VsCC5crGx
EVJDTg2LWwCt3rTCzr4b804ZCzvlCL0LYL2AqmpTqWWQ0rZ+PClm+rqcOvTR
iEkaucjsHk2bH6MW9d+pguCG0IdJmcmQyo4+g+2B7B3FDhMMPR2PztcXHSgg
uD5PL6J+UkrN+2USVC+jFjt/YdFcVmFTSDbS+NPK/hQLuAnNu9Xtw2Z/BVX9
UdQODYdWer39yBHltBPfYtNGxHBhrl1dvd7s4oyUL2cT5jLFg/BhQZ3gy0m6
Va+S/1YhnDOS9fT6RIOS2tgw3P5OiOwbQgpdBp+8GsgzE+7NhEttZNeY2074
ZvTUWqp181ztV9be1wdntsXd1f3zTP76bdPzgYdk+WP5opsmWMChEKma9q6q
12zKWbMZh3ujtEKjQB9PFQs15MoZ+MwOmhMRtFZBDeqlEPAP05hM4NMlgfOQ
fVRhdONSV5ifCxxfEPIyxf3oXi4lyGuHhxDe128WUtDWzO74rDOgeWNQOYHZ
iak4tGbTrOJKzbRN+NnUI/Ww0MH/I55oOWBIPH4lv5+iSxJI3+rL4fd+wiqC
Mt1mhIFBszUuQOYnlRbUPnQGLempylBGnOsD8Q5vc3wb7CedU7iadEILaJPX
QEb85AQB6Vwv3IS/g7n0fWnIYTxcp+umSzryvRr1DzcHNRJuDqTVte05pSt0
BmMyp8BQKn4gyJ3uiCswTU6n9vA8aFvODEvwaSD99VyIam4wjyb/8s63RoB5
njIpKM7iNGUXaAJp+bk1lXjqPdDT87ZZqtMm2rQTRgNnT2wtU9KyHGTp0K/Z
8aiVMCXdP7rmKWRdpSgmW4965qFr0WwbiiWE4EPpU3baLDf2kZDTESJDZc1o
T7Xfa95cI8e6SwBMIUbjS7/LP+PzAz6ypR2mtHgXXZtPG7qY4kq6Mpv4cCb3
1fQhZaKQJsSiNPS8SojE5W5rmTOiWcaP11LVga0QfoVn9ko6xGT01OXIdeGE
a0EBOT1L4hU75L2ShIn4RyKr6IGX2jGeS1mFoT/fWTMzcLSa0qG73YP3TLmS
/Vs+nSJZSsNYD1yufSq9E49xQ0v6YJIPEKcEZMuayZCabn/Z+N5nvQFQpc67
PgvnR8mHl4ksXopGLmMe5I9iZc436ZDwc0rydo8/GV055jPOFT3zBV/38GtI
1BQLuyHGdctaWaWK1V00Zf0a9pGoxr1fe3X0FakcrFESQ9YhNnMhn2N474IJ
VMkVCHRzzmLtjZoLU5ah7RnYQod+vBlLiXQeOwzWKNWem/vFpNVpUVggRGfR
td2shwJwfkAJUfU57IZ1HWjjOk2OvbmJp/Jk381aKp3w0qhHC/FhFk6onDyf
HXrLQcRCPyaI6eQlLaVrxcm+iD1FBsbfZaM3PcAE+8gHMreOAOFsOKoACeqD
xiRnKCbDudp+p0I1zfvLk1VxTDiWzJJO4+1TgVoCctF+J+MCHxLbevHvdRTW
gck3/MwGY/TmUSqiXe6jBDo/dkTv4hCk6AA4T9J79bpW3yMq/aFwlUDCoZ6w
Nbn/z1mQ0VlxHP52CsUf3Id93gbJCNEAT39hjk6hXTcHT/X2QQTw5KJUs/94
OVo6YkZ6tzvAUoPyLxY6PmIe05Yh3Mo5RLVxcaSTS6Qw9ro24cWReqqdB9XX
/9HbpNQ+9SToNgt7O7GkK5BgJHJPwvtydUz82kDhn4KaTd8FybxwWHh5hWU6
5EnZv4+mtsbapQZOx/ksMNEOwGCzf0+or4EkZPhVLN1rpdx52qd9aRpjjD7G
KPnAF1ayXqySDreFUE19trAfENprPXQUEG03SYs0ELyzf4ExC13IdvCeZGFh
D+n0015MYopwoaeqPpMv9g/WCTwwqsIZtsU/AwUdLfpeynWIuhz3kQMAdTW1
rG2xhHX1jpgq7o7JrwoOWJjfI5Bf868wUcEfmKTsuabjuZUH7CdAZAnctwAK
5CmR32grIytar7cu1265e5OxIe8jgJIjuz01Ea9f+mm5JwoI/LSV+T6ERWD4
sY/A0mdUYSsqPoN5nk4aGpaQ2AgRxMRnx/b6aXJkPIxDzoWVU0Z5NBkuj3pD
nJ/Sxkgespv+5+DnbjVLbXsUbxh/9U8VbaBBMpeu3RcsSszJjvqg7zPpzW8m
L+wHnHrN+TKNgE9+aGXAKY4RRyhAH2sHW4T/CQzseZT7UgP04qhxKM9jMyc8
gtDY40v5g2d8/HSYvaLciRIlebtQKMWH871fYoBRInU/5CO2I/bS59YynJgU
uUSAcKK4m+q9xBA6i+yZrUu8l55Rt9agfQ6uB+aQFYyQRleAa3otnSJjrAAj
N6nogdtrqx7CuBIaz94Iq/UVvaIGKHju1lbXOpJoj5KmpBzMoHk7DWLj+zwb
IyHnouhpoavGUDeiMgMv1rV0xaGYlPL/SlRBXHUfBMYvzOSUXsB18OXxOBH4
hGtsdb9DpYEVmRSq5yNRgIdLlETUQZpGMllxprMaoLT1HXRpkYC7qaq8sjlv
zTyIK9ASXE1w5t9Y+lFNvCRlvsQZ9QwPQvFQqu7XWDyucESz4JTZXlzHGkNQ
qk9Q9kTvk4okZ4x3wLLDE2Wmv9xhRH6dIFDF9tqsPmf8j8oNCcN9NdLVKSUT
zAsVYJEPUv+dLexnWloTPwLc4P8TRh9oWrHS4mQaKI2OfCNHZKGDr2Z5y3/e
HGhvfaG2ZzSJKPGE+oQwph5311Rm8Lt6AVQLu2pGPLhNdg++GteQGQjR2dMx
q90hnJWkTRUUHq3Vn3H1Gm9SyEY7jZGaqEB4B8N/g9o+Stw1XwAaeiNFVsRT
VDo3Uf9CAWJ41NH65pizfFNBT/SJmpL9ToE6qDu27AFYtzI7gW2eeyUsm20P
VkXeZ3FO7Ejnl0ReRnPrmwxpI8NpJ2+nu34y3Sa/jfbCJW7oO/R1l4bnA4bI
Bzq6GiMyCAMjjhAZQ6EcbJZVyn6THLzwR3wa76hdlpHLl5E0kf4moE6tunNo
kymDJVMlUS+q26GTg4VDALx8uNamgjERABIuhSsB2KetHWKrepXemE9F7xco
jUoJTQd9JNlwdXH5dkPgg3kKea4bb9c7vL3Z8lX9VuRfEHxrIDrJwwDXdD4K
WrfsaIV2zizOt9twFAl725zhsRKndttfJ9mnRrS04Y/pP5RGifradOMoz62R
S+WjWGOHhaWRz5ZjmRveMNrJLJ13bYjw1ADQcvlpNxQdVo70/N2GR0rky+n1
u+mYvex4QsrTnCu8K1XC+1PL3syZwvIME0LQcJURRqK5K32uSTd6qUIC9SHc
p1UTIBuqWtmMVYK94PDheCksvdOI3IBBn85sFigzsCn2XUcSNbKt9II6bCBB
2UeQBZQYJRXrjl8+zUTr5iqjLrK4OZAJXQVbvbH+x/pHK0kRWeQQ1UNrdAU9
KPUKdBSI/Y7znF0209Vgi53K0irq4hSqGHNOsSXQznp9qBKq1LKtS1WwkuNR
j9y0g/wK7GrUJ3eZJAjLai5cEQejYMinrW93j/ztTB9AsTTyBvGGIL639nRO
dhUmkaoFh+Pz5T4Ypgg3kRf9C6UG5YQS53cK23OlbUlRC+RqghnBPxDWyRmO
Ie18wgG5Ol7FhyqoKQuGIIdL2qavgaBJ/AT5bURALQFrFq57qKtbu+7Vpuvi
0rZ8qD+b1OcyDJVZx7+YVWguZ9oOkPFoDO0SGaGEtrV6INwFymN5li9YsXG2
ERglGYIzIzcvusRW6zJjo5Y4IXKNVXaxxpxrkN5yeHlC5Fx+7MUcQrMEv1n8
vGm/IFGW7MT2WoKTcbik8RgZRZGm0J8VcdY06dcWMhS/ukSkkUwCIq3WdABo
g4Mm1AQuDbv9hXp17zItFh7aQRkKCoYCaTbl3kNOdzrzahw8MvYkiVYdGih1
1MbNSgU18PNYTreOo5xEiG6S2na8j5c3z0Ac7p7TyB8rZIOfNMULJli87V6+
Pznv5O35ne5oQeCu7g4hZpBvcEGl2Zjt0RPRNyguvZ4y7s+vcKFwMO5EzGnh
RVMeCEVm1hPrOZeS+sQ81u1FJRy7HMDK3b5pKWLvEYldhOCtIGcuqOL0Dbln
lc/MGTcQBTJgQojY20xgrxfbpqziiDuRiTc4ULsKgbhVNzpznCirJITQBZbI
dESBUdbc7CdvbG5FUM1ijsYnushWMvwluIlbH12kExRtedwWU/MkIILw7/CW
2OFONvf/4LHU1ZcS3gJ+yRPA5VulHXXPMQ12jwt7ziewi4Tn5Z0IBslbdq9M
Rxn7utO5fNxLiva2w5QUq1JuK+sfUWw13bXJR6KSTPjxYP/7Y1Pdsyvxrh+b
h82AUDBqHD918Wea1nmXKa7lyNwZsmaCJcRIM9OpXIAHmK0nzNKi56VrNCQt
AiqwNdQcOmu7JyWXPbQEDT0mkQt7EG1ErfdK7QRmV99onH0d1yVzAzqjx6W1
SZrSf+cR3W4YTXU0VC5KDIqidU30SHNc1QohpyNjI4vgu3LcHInEsIWtwnZK
2XYw+IbOrqeA1obm5OsuRFESow6GsE6pt6iKs4K5q3ax+W2OTfvEgt8QkUg/
G8bKo2y1yxv4HJidwv6+i7hHexsIiL/3X866BaS4skNxPq+w+XqJVZNuY0wh
H60aqrhuOQPP6WcKTym6jC8krnwi0qWP0Jf2OkFMCa2+OxaI6rwmC7iGXVP1
oPPUKO+snHkcd2Sjd18zinhgXtg8WAG3Y0eXemuN6xjx1T26yvgIPW88cTwb
vrLh54Q6/RPXWbF9ecaF8pEEv70RcxLpyCEu/yjKHnvmrbceRNhBrqLfxMuF
CkKBjIBJ5p5eZxIcSUEkV3UzNsROaWPFB/Ro7blVOVQSfD6WQrV8au9hse+6
BnZIXnw7A3noMlZv4VEZubkCk7HwSc3iHvB9GJRq8pbdJ8//slgJW9EAzIwk
B4ba0ZREaE19SYsNJ2asoERoZ4YCYHkmNYdsZITvR07vFXvKY1MusFCQ+quC
l+0kRZVNA400pNZIDnuBTfwiLRUtNSCMA/9Hy7Lw8atXfubWgOVkNwMDBvs+
MSuzW4XnrYUdfmAhHo0gigpppbQ1uuH3xd5OxRRI72akoLcjZ5PjCx+k2Fme
Keuhr4zDMYQ3R+E2uhoRp/7sh4Zao8KbXjJqYRlKepmnflDip6bdtgBTOWma
iT4YyywVbGAAIoBeN88UBjG7nxqn6smNamYVaOq024p6vhRIhJzFV8qTIFEY
vhmyDtDObKH7PWKpZqyT7mbuz1xezlPgDROh0Wf8g2gHneimgSMrNLA33ve/
GMUjGxmnMef1PFx5+cbxBA4hLYpW1B9JaXjSh2J0h9ovckNMepj54BLOhHN/
ldPCCAjybHSZt945rgVAkf+ikWZQG2YcCuIDadBgg86oCwlE9IbYIGoqxcFE
4yRonxrHRdsWUAILIjqAQICgAzzqDb/gkDkptYiRF09T1pR9/7LNsKhjZyvv
8KlS/HlVJFqsaT926R0zO1XdgyVElmZiYR7JOtGRyJkjDL/yg4nFMFQYO7Og
RpQ6sdSQCmcN0pD7N2u4cHPUaK7IsLRZSYMZLQ7aqMF/3VJyiMmaCdsGpN8d
GATi603clPtkzzpliLK16j1+qrcDXr9X1VxhEdt89FGz5TbO2zgjgO4RcYEV
noHjiXBu2VdvlAFV7t4rl5dwVwwPkE9VAD6fgzHemujXiQ2iNk53t3DvRzF5
xK7briRQilhG8Y2aW91nLCHLMAuRXiPhSxfzBhMDN4RAEDSXoDoPSsHX4IUL
l13msypOJ4kVppyLjgUTl9lZax1GzeUTJi84MqjURmA3ZRnXlAXAocfV1qVq
CtOPUoWKL3iTcIkO08nax5myoqBuJT58oGxOXB2XhWtsoGQsva9BgkOdSEFu
1eoCzRqBWqHRbjjwVL+WJkmHrU1ImNnahXsYMfeMseLHtdIHVF6PTEtv+H7l
9tJcD0jviOljgNXa/UpNLO9+gNjzazpKGMLwvuyopHLAHrTHOUzJ/MMtkL2n
sY6f5bMNl43UQk15po5ygfnJYgUCAEE4TKHJNPElrjWV2Na7OTnHsxUkwl4d
KRtLytya2OUbaGMbmElcGr3JMbdhyWtan75qJUf9fTR0ocWbmyIqdQE00TLE
eE2PoxcGBodv5K71nyH+Yc6+GB7NpzUaf7rFZRdYTmBIV5qPmd+eCDb9a4kW
vrFpHkam7nJO2taHDT3MCx8SPaO0Jm85+KwvHuODpryULxvVJRCG6M/b3UOp
Dobz9Iqes7x33mcCccI65IRCxInnnoShAMUSp3MKWE9m9e3IxGcLXAitYbBU
6b07KIh/iGaiTSH+EjoCklvsN95K6O8lU4mr//+Btc9EpEp+Q+6Mw/cgew8b
b2z8RJkroeDW02YvNBW94Kev+AC657/LLWHGILuQxGVpc8mOkKqJvgGg5W41
jGcm9tgcWj85PyATxc4koL93i9TzZf/k1WxmBimjoPq5qPjd/YCCscze5usF
Pv71WcTYUzEBSg4TV0RWrbVOk1vtJjeI6SBaGV0Ruo8qyx0f5Nst8XBGcbQy
b7Sg3ck5PsQ//gJXu1ALhiqATalqalkvOBO2dMAKu+KQV5xfmLUCKkqiH9jN
O9lqlG18fp85NzuDIqEs9EZSPpPLxViC9OPftyTQh7ch+FHiBI9d01sqnJRt
JwgP2Xeq70LZlub3DK/byi/nptXNDXXcAz151AcAbabkA6Vb05saOY7qHaL+
QIEsyKzBilEEmjs+2PR2DcymWanrNtoswFnAApppXlh1kNHOrsuLC2jLNH3O
xssQS5akD5ojkQxG4ljTsM/4vhNsdgMYtV8nnLZ43xopUeOOx23PzYBdKAfR
2a2gaGAp8wqMgr0tLltGZSeffTCZP8Eakvo30+uaqpuxH+k9VRvCJaSyXFqW
Fo3EGsAHK18dOLGVbwoVzQMVfCDR/abRO58clN6XZcl+ugEfrBvuhZk5leFY
0xUW++l0pwsQZlwpgDN+ELznLvEDraIGH7wZoDizHcRfGn8loV9dQF+PHCBK
AWxWzYWDi9htPicx3ddpAdWK8tH3R4junRQnnkdpKh6KUE2ZtblAHEF6goCp
VensIXe8KlOUz3VGNGYHctGjCsv2qYUPLDkQ3qxIxfcS+3MAcTJiCpB5R7QT
ZHx2SrayWitx0iE4lEeNuhmAC6+VyiiU4fstB8nKi8fUpIWlM9gPBbjM9k8u
W5Cg+ubc/hOqlJJz/utuuVjPwjKo9Hi+FyWq9MhMqp6WftgIlDp+HX5inn+E
lU3xzUlX3JQSBuR+gUNLMiHJ56bpOrJMl02A9Ws81abf1BDr2RqXHu7E32Ph
3B5WNomTAL64s2LRUiEVciyERFN541E5f9DumP9Du5qmUR3X3i4jSh2QawqB
Ff5HdX/nSWpocqmGFppJk8/HqV13qvxJAkJKwQMTNEg+Y9G2XnuoHNgvBc0Z
hcds7WuvkpqiTm94F4JWs8LGYnxycHNNRoZVKvjhEDEMnkfmTXCko7TO3F2G
8tsTWWxN4gsqsyLN0zk6mP6U1EHrIKO09ekvBByzStUo5yCHlFyivc9TCYVo
QxRXaxRZg+xpntSgvPFB4+WyRJ1UjBG0wxZQ7ey/58srkoAe438+m8po2+zN
L/gA85Ey3FCGypoVN5MssvRetArB1jZiWk7CbtafjvXEyJkTU3/d1h6TYikn
1OcDGx9om1MprjCqG4raljV8BQOT847tEfx3TPw1byrXG+ISLa2rSn5qN9Bb
S1t2iKk07cgmHdLw9Yrp/N/Oycv9cOhlt4rEL+KxQeUk5F15DcQNKF9MvtoA
8PIZKGtZ0AgbDvAEbGUivM2MobQgAU7e6LvM1ymzdOIzip2hBWWwInfRFfeT
J7qeJW4/krjvpxcn1XAHQbGwbzj5698h/YCPGMfSoUy/okqBtz0IjcePqbd1
YA7HQ802mO20/90iQc2joUKuGyIish+zWx/iLYWgv/6VOk22TK9f1ELgs1hU
6YGgVSGsPB+UOsNPOfbh0kBbi2paG3c9kCG565kBs7qH9qx5ydK7VGJ1nAJs
Grx8IMVR0033bbSgXWyHz6ohqvkgvI1R6TAccLCuzxHnkcqtsBmyJDlC8e49
JquhNQ7UtrozXzUrnbqMMZXdEJQ4rMrUID3XyxfpsSA0MjMZYk/W9gr94ur1
cmY4YdtcS/EayCBdfPKOexmJm10xUtGoFmisE+c6TJtn4unxgGd0WF9dvBSh
YHKVoChJdeA3FhsSC3umbYE7G/wSRR0y6KYCgH7raiiQfE+KT4UPbljPadNS
PIim66z02a37L6j3KriYvEoXdSDWbn/D6QjOhf9BBtYpSTc7r7hcBnrRQsQ5
G3lWj/wx9Dp6aAy3QLfV3DnwGmCKCeHBPN0ElODWHCOIcnLJ8qHMOJJyifUx
t3ySYfAVK9VN7puuI/l2N9+amzAL38mM96V/0/nOcdY9ADdjNtwHDpMgMoqw
Jlc7YC+gWeHWzCxb7tYjmlhvckUS9t0f27kF5lPnHQh2osMDHg7yqUf9GLVj
7O2xwAyDZzmx5073bKgsCs1/cfv1uZZsDrrhqnFQgFH2do1ioS68dGQbtKxt
/sNv1omga16VX0/0DdsMs/OTIBkwNMo00r9LpqTM4GQ027zZH0hJSFcxV2tk
FW/ylSes6NKpukmc6cYliYPVky/ptaS12TuXMdfMTwg5sduVxN1wnXEUfRve
OF/0Mi8ZOCvwPFP0a6cwCMFb2TIKQKG7wljs+EYTexGp8ywJXypRb0ctaw/v
Prjz86AMBjJRkwquJIB06ngo4N5NBwmLauKWPlUEagFIf5vL9SKO47m6HOHk
KfG0wxBngDhRnOX8ZLIapHt3Dtplz3NCHWq/OowjG+IfwUs+4MRXEJSAKMrR
o/6HWCSFJJeZAGLY+sgk4af0yUGp0zIl5kpBE+MEdVCPBrEHQiiVjCv0PKYc
5V+cSj9B2VklQoM3wYQ25HJBfUnSrG/m5UEbLo7Y1c6SeYIjvdJvCUGdYF+q
85R5z2Sex5ZR0BSm4zOxcAG1MZk/i16kMMqAy93jjKG/4gJMsX7NTKKvpSQv
T8pXDtXDYhutPN5iCliACQSIYF7/3JCr6lXlVgPO5t6xqF+SBX+IMu2CVkqP
TofZfi8sx1UNOfYauyrxGm+b64Q/ReQEMZb/jDTrtz5XlgDNY66wvmrFenFs
UFRxDK3hO/xWnUTyMm9+xQuRh5kaJxS10t+XubZ12JNvMHvz0LO1i2YuHMUr
/WAaWA2YZOSiWFphCBjq6n25J2H2k5mW6hET/5uyEUIpQn9VANLRcqoua2Ba
hMx5sfFGv4e0Ze5sRcHPaVOPYSb9u69pMHC5S7ZR2AP6raz9SJww4YlNxH8E
pny1N+ipSczkqiKDVID7l5zd0k89lTvVfu2SQvJvenLTAhGi6FZfB3p4cQwV
86N73+sJYHQy8WR2rP6o6crgo8mjsDsUS+KfQHE9rA0JYEDxTZEVogkXZFo6
lVEjoaLFUQKVozIOwfJVZkJMgGtQwhvV0cnvdD1b2JEurQ2zptUbvBTXO4Iw
ujl+b20bROeeM4rdWEE0aMIXs2CaUnCjknTPts37AnowLXNqAK7UNw+NaNaU
RkAhHfzSRwH9EsuLlLyaB6HU3/zKsVRxWDPNt1JnPhqXoKzxW4KYa9+gX1Pl
InAfhzagbQ+fj6Sedag7PVflHyfDXip2+Os/ROg2MP8t0y22LrbeMl+7Cf6D
leYn816As822R6rTLrOP8uARB9w2qVW0rXtMEHEtJX3uULkCBl2VLGWBBgDk
4sKRXF2YH+bXzpK3ldMUfI54gT6tUCI6vdDSrqtOo3c5cyDa3vZk4Xs/abS4
BUNWWab1Tf4J4qCyt8pUyj6zqMwlNB4cCdwIKXJFAk1A5+W06wXv6O69krpX
55ar7LJpEyV32vE+/+CWyECpyPIkKq20XAKo+n3eugaq7TmuMZY1IzcQpaik
FwQyVE5FhtYnawLU2h+FBffjGXlVNdgNlz0lrvF0op9orGkug9XhfNaTn154
Uehd/HHNlmuJI7bTjCEO2AOe6RxdlMGCiIXVQ0LDb8eCx1r3YvAcKlQTn2Sw
x0vZGrmrvB46kgxBinDYxD9WapAr71BwepwRglmMAaXHPFnNyUuww4ADQBpr
dezBOdS00oud2CsnXt87gGwDfI8sBieVHC/rhRAcMzAcChPWZhnyiaGsKP2p
NRq0b9VTDwz2rDMT5YFEI6srtIifG0g539rHLyqmRrzYFCMW1S1jBTnKeXqX
LLP18izP1PbYWZajiXKiyDMG/UgjtovgB5yT8Qa3BYUvLkrRw/tzbsXUbJ0B
c62wJgl/efjtnUsDCBcQ6gm2Vi7aVFNyxyskqPq+o8i5PhXVRj/BpilNCvF0
JX+w66QGqukoLJ3DMhrQK6jAtGYRlD3X5m49g9khojqF9aWxk2WXAvtm6h7A
SyZiuhXaWoaV7PCwpwXYSIhrTtnHLuycDDSmHPPHP3O6zx2zVH97JHC1R22U
rb1ux5oBR5+kffZ6MU8iv38r+TVIwCo7Zm/VEIOOPxKdv4ke2onPhrxKy3Bx
S5HKuWPCMW6+FEhVQfhaQTUBj1JQ26Gn0oG1sGU3/n5K9BMYqM5KO+Mf/RCY
7sHjahIdoPrnKhZuESTbhtQJawjrq9egmm9oxpGnc8+NeqGfY506eKZsMaSR
P21XMEYgegJXt1eIB+UBwAp9nwbUteojBj7f0nRC2FZl4LGibQN99y+OlV6D
ICRvqEw1rtTq3g8ezv2vNc6s8xT85Lx0UCUcndqrArA2rHP2zIlKFlMTacaJ
91UliPzuit0smw0iRWHZwbyx8LuXSOdm9asdUopq2BasQEMW6cwNFH5Azs7c
nWcEDBCzymN/b5FWsq+7MVeyEaeRWYrJM2LIE1vQkh/nPb6+xk0mpGpSklAH
89crmxTcRUrf8fPZsIfB8T5HvZKDoZWZG6UJsq5kaGkxJhMuRjyZ8SBnWe7k
mvoVSANDyevJ7ELpJYfXi23M72jIdz2DqHpWHd/5qPJ5f2Z6JbJXGkUUJK53
7834FLW5NsWZX9ppyACZcFPcSIXuasg6WiIdQPGgghjuZs4YM1XLyghJbsqR
V9t25ElMWRYDNyeVGhFoSGTafWHTJhZS46KrMM9GIym0mg5BTRIdiLBzOVc+
0/s7ne/qgG1B/CFfCYfFH5tgvFnmU/iLzxPbO9vfuShXT7NCZl45XMBnAbSn
L02YqR3ibzCNA5xPZHvwwc4jqJXzbukimi1v91K5LDB0b+xo+2oqClC3MxBs
RDGcogDfufzTEuKkHPjHegmlm69J912KSHaLPL+4wBAfC0KDIKS2PKJ3nYLS
CQYSGUt2t1xrXIJHLLfbqL8stKkSKH+wa4LnPNlmGQcv+BV9juJKUYrSIB7o
dJdK4D++m28zTb7r/yMVTLI3Ow7Ixhj8sNv4W5yVTjAGu6pWU5onWQqoYlPi
1wzkVrFQp4loUrcocYwEa30XOiWn3550YUdeJn7vCTNvCHvhjxNeSne/d7hQ
ZEZ0tQjoPXiI0uSU9FpFzCYi/c33deMMm5RSG9+blMvtl02gGfRs1u+QlFC+
nx/Q80Q5/iQ8ynQ97MyBuqBLFaziC3QWenpXW3Mclv8Fq0Ze6fDGT0VkqmRa
NOE9ozCTZnYpJLqy81pFuzOqm6DjSLmpQ2qbA9GIq32Z6Xm/vBQUbBPk9T+z
8MZUTajThj4uk0SPD26+6xz9/5tu/lcDdRMNAdMO4vcyb/OC8O0zZy91zvyd
wEICMpgyDWGqUv3v3culurDU/uNYd/HaNZ2TzjlKkxLrSMRwplVFBtBSAgbX
Osm2skK7v5SM6ACoHX6mCDF8WzaSLkz4JoWfPgh5vUvX42DuUqGCJHJfOblD
9T8pqvIEBxl5xzgVEh/J3C9gd7Qd/C2L8jjag2R+w55ZfpiyzC75c9nntUJm
FH1EJSIHgrHVObRXeJvSIQzS1A9Uq9Xqir8xM8kgxclOQ/dRXLSo67Mvi0RQ
i74POmFRbMclg1YK3FxieRsat7sWCa3pOE7kO0B9bClbEeO3qElP8rPtPoCD
m3dhC2y1cL5FWMaWFvfchBdyToJX0XqgrbPOPIcZshb3dYOWjkhQ2bVEekMH
nsW5ZvNoZ6RpT0DQI8OTU14ObDfsivdZNGKiglQad6hLMPhFRZnH+nggnWms
NajI++sbTJAOuv2AbdyNAOPp5Nif0mhyNGZKIiB3bXVA6PZ8Rnj7IxeaU6FE
vFu/NGsqGqomRQSeWdp01mysBE74X30yJ9HxPCJExNyKTilj3VA5jGwuebY/
iyfU0kIQo/QmI/PEvOynSLV7G3eFl8XZ/gogBOcPJumwXGm21YEncfRixqPO
bAtQgWiDw2qa46rpE1P3AtTDjReSg+0A011GIBugqCJlcX5WPk2rctxXB59z
2rQu3cgn57MEJ2WBFJ2s2wph6YqVHgHASuCg8/5bNu0ALpKS82iJ6f4ELH4T
ajRxibUVty+bHih4EAgHceiivgDC+J0Tk7/RSbUKN+Xc7SvXlw1aOQ+Ab5Aj
vIpv3Uwya7Ytyh0wweb9iyX4kk0bAXKZzY/12BQCBLJSEV460/7S07J06W8b
CG9ro+wOI3O3XxraGu36lKXlHYQ55SrrFACimjuGidbNUDyNNX8s4mkm7aT3
LLFYxFBFMAmFhhPL3mG+14rgSaWdvbsRznJz51nsKpMYLo2QnM9Sr/GE6APs
ubPn1iTf9mcrXnNBHeg9O0EPpAlW8z3jvbRMRPwwDRysTDCIJAopCc7eexUw
nEFsDmj5D+s4OFXqmIBRjtTXjrelPTw7IzBc0u11z0xxg/2pQKpE8qpVVWFQ
FPu+Vsed305vFF72b2x/ZMV7ehGf8zrmqkBOmVwmbzBifEYGRj9wa8CkVITO
ROtV4+Y5RL98byJ26RtloukIIuZz2lKDGSIvVXaeXvp0ftkwz+XTcA69b1OA
gDekGJd3nM9yrG6uOL9S1A7lLOPFnMXxK1IIiCMbrSm1L1rEA3n3UjkfEIX8
oM1tXpWO8ELJnquKLbUvS4a6l3b/4Uuk2oYAHxQ4vtuMWfQBirsw0zG0xg5v
xk1vSc2dImzWszoIaLcGTar537+KnTL3tTgkv3rGnOdRS05tljlQJbWBGnp3
6bJgQFBBeqLD408jze2LkwN15n2bzJzWJtln5FkAPiqgDTHR5WtBXoVy6taf
NBmZEhu09duKbw8/V/CnXlQWFjxXOeP28n48m+MX5c+YBGQ7SbFbF7lhiMft
3O0VLQC0f0jycGiGeqHB66BBBYKZzmqGbbnS/8ZRN8K4w904prg+xTupi0VL
+gAwe5Jq+/XvaFnSFhZ0L0V/7665vNmEHlRwjNxV3ofsqbtWLuJzwuYYww7J
Yz7QnkZqaqJqK5rxwPwe8boyU8+WN+UmyenG0XkJOjha8smrLeO0a7iJxCJD
OXh3ygCD95gFG5dwWhjeORxFOQcS+7SzyRDGMs4tz99TBzDZenBFldQd/0qR
7VB8jK/qT/6QCFjjUgOkNYl/kt+/HvSfDHRHeBLOWre5FiGER82v8l1AYJx/
uKk9fJwiSNRIhSrTiS+MHyvZ81AQHC3r+5WhJesNyh8da1gB4fF5fgIJWVHT
S4AQSgjWEMTAuALjFZxiJRmObQAsFwta7IKgoStKN8Nr6gn3rs+B8kQWHaQB
xNNbvunpAtf92Vt8ocypuwFtreumvPF4QwBsya7eUJ0NiPh+JpGun8ceN/ib
6//tMmrUKWAOu9UbmNbED7TBZBWTjlEObrP4rbnUIBEPVKMktp14RcCZGgRK
ZNbhFHE50IMkRgw2R08GQDxL7/1fZtqMcaSjTr7WnWDoY+l1x53MdnuEFINc
6hsftr33PPcpN1anblFw+eA4FFWtFxWlOGQtJnOjB3+BX/hdu7JezFyFY8uK
TD2bm6CJpe8VQc8xb5iWlSmHIVtTzh9nHZ8r2sOL063bIQUCfglS9R/hgmlx
8FLAuC+NwMGyRLZikMpXAtOLdx43aegbXOuRqx67kfO8AKN3JwbMF2lLkX2M
TzSTClMmlsynNE5NuiWuNN2Ic/DbF7FVGTvF0iGzlzkhNtY3EfJUZ3tm1Jt8
EiXjWaESJ3ybfpOd9MUXt2jrt3hwBgWygqtKLRERtRBr7ZQbde5TmMLQs8tY
35UyqrIt+avThEjzadP4j82H1y8jW1fTTkAP+3jyp63BkORTx3po2a+uWHb+
CB5XYBEiJJfIKsx2yOjNUwyglMmpULY0ujmngUAH1McT1IvKYqE+lX7dTf5+
8RuPaBVzdaAHKEYLan+K/6CtA0LI741GTb/wE8syJH0Zm0FWgDId8aEonc0C
9Hjcx25dT7kJhIDbcZhKZtMhPUO9Hj14eAkydQKyseWiB6IKE5+Fu9gHKyA1
8I1KYpq6QrU9T4YhxVy0Mygq19MFW3tXS9rOpttRgvAwV1R1dwQljvZ7j90f
thEtN6hwV45HpDM7RtONMZls1p755P7QR7HQ4wA258p7kuDPCRGnmfbfmGUi
4X8sSl/l0jrZFEM2iix2K0mCWjyg/2hVDRrifBX7A3nhiT2ti1fGIu7mk7/w
1/bwRUie/Rm+EJuDCFhpyhOiYz6XUH7Bmm3KXEVrkh5O9x2LJvUYP2RVdB0n
aNrmrFtQ1V6aNJSOEej8il8v/O5ZdWJC+56tE4KIox9w0UzrR99db0wnopqK
why+2V8N9HYHXW4clPZGt5x76djO08IJ6KEBK8tGKqfJGCut95VsqYRyiQHz
uXg1P6vtZ+mhqiW7RsK3imMW78VncS5oh14Cv4NUuRiedLYJqHCQzXOzAOzn
1xx/pWahKRKdwHdiCymSVkid9ASVsOIFSgZqW+y5dBYexpuWej4kzFJSW8U2
biN55NN+vK++62WzwA6T5aGloOtzhB/EQn+W0eo4rmH2FLeT+nWR97TDkKi6
cZmiTxQ3ptwT4+nb5Ql6BuPxTDoxkLQkTMN5EJDwxn7C5MV0RAl/x0mdWEnX
NfLHSF92ofL85TKj7jCXRWFd/bdLhGwjDSpz4M23o0kaJXf1WQMUthrL61Sm
zvCwYW3waOwXbiCFF5n5zl9GeT4IGk4tVtKjtpPaqqxuL+AEfE5Te5Z4V5c2
QO98Bd6XkNGIzz7CEhXaT3ZZ2fr7s2Kx19FP2dx0MhbgwCqT9Nkl3hYsEaxN
1WrhMpcN4gAYJKQWvjX/5ujxPaNATzRvhZG4L9pcIk/ARyVgb04QTnBSpFSY
OtEc38beFj1Ww9dL8t+pWDqxHLZvtEum1M2SfKh2re08CfC5IjhSaA1LmS0F
IZKdqEqIpk2v/nhhP+VfWMF/wO4vkDQyGHLaOvrxkvve+RkZqv5QD+/XDD+q
6B3j5icgyzlKL7RZSB6Riz9YZEuqH3s2WnU9dh70Vd3A/aI4ojaDwfsfdf1s
wbRD31QvZtw48lq0drNTlt+jYINCG9J3DaYC8DaBYk1R2Dpw6bhnK3Plck6w
y94Zm1OgYfH73K5+FrFdUxDiFRJ/rQb91Co1OyCHwEPdMlrJ5Jt/z///Jxlf
MMmzFWuYPvCDBF898C0DArIXEbWb2AByxu63+eF+J+SA56qTbodG8+dP/hHc
3NKZxCx2/TpBES10PCcBqUcRum67OIglzPYkWFGnvrsQLm1nJR7wwULV/Iii
ac4HvcO1Mikyj32sKrIm92/pd9i4Xw1zUjH3XABZokZ17HmJj/X100s6KFCt
5B6exKXXUvj6MAlPH1XAiHHeGUsJM6d6PGkpoU3qatsMANQNwqIb68cbrj13
5O5mYVE7o5bY0l32ZzEYjFkLvlkgqN/sZIds1zP4zYxvB8idg1M7YIXCJmWZ
HkvGEBVHsWAixzpdRLVTH8bSMI5jSyo28o+QVVY/m3bwZYPYF5c7jwM7xIXi
lhu+ZDD9CkhQb6ujs0xvPH/+jTmo1JZA/WFDqD/owmZFicZ6WIQ4lXDdMWsu
V/uKH7J+i8E4cdmqDzRk59iRuEH07jcUnjBaZK5cbheielcN1lInxYvGAQDK
rZKeijYkzuS+8zksdUCRBIbdrGN+zhqbyQ7OiF82EqF/izzWlvVJSRv8F+XI
jlpaLkAwMBJb+tHGLrjerZNFD2VW30kr1m9oPI6E2urF3HUvbgvb+U+U0D6U
a5sMQNsLj4W3S+0GFJbGWq84IuXUe4o3ebudxPJxG8t6j10zrIBmW+Y/vwgh
gteguLTbyPS1DpsAZTEmETTnUCIf8ghID0JHYVrYIJFf+0OKSUU5N6NtxJ6H
Qv/y50XWpV8FW5RNgRQ3FtAIPErd86LXqWsyXG7tzx2n4V5wrorT0E+b5yne
VYho/Z7fceINIu6ECmVX23xN2LmrcTQBrhOq4Oc6ahbfO1XCrdNTEXbCD2Ln
aY09AAk5bLVjQtXDwjP65Ufzd+EeVt3MwtS1AcTpoW2VcHDNyPvmaBz+ahRP
JNCv0Iyzvd1Vi0eNcvfP7o0cBsCj4Mzw7smw9r8d7leaZb7pTty+jzXEdr0c
15FRaPH869oefEUx9JTrpmYUbHyaYf1mjD40QABqqz4icjOdTMr/LEZQP1pS
/zvvDuVlkwACAto8q5LsfRbBQQ3MMyFySuWmLTM0OL4u9tC1sjLu45Ce8nyr
tywFgM4jAge0fehymVIcokuaAC3CAkBMl9u+fQHjt7pYbXFvSUilNgfqcFPU
KaqlSOsE64Ok4qOBBAwx0Ef7FycoNowXP82D9wt1GqnLjCssHRXmNQ4WP3np
HX90UmAFTeEotAwtZrZ4QGvjRQmvFdX0PY1lha28IQUOTg2/MHk9roRepSJy
tsqOKm2VR3K8SREgoTvxKN4aZENFHm0Jp+FY/NSqRTHR8HkCYuIcpzyO9Kiv
9RFNfL87quc4dPbok61d9IyoBwJXCQ55toY2q0X2QkajNe9pZOBYaIR0Tt5N
3S+kO0GihhY08DYqTtelrkqgjxSholXt7qYZQO+sVjE+PkAmdA1a00WLIGxZ
h2sls9ySZOfD5aldc95Fivw9WHNPuyWOfQUOfeDmSt3dd4vUQnXUS6tZALkj
uwdqeRxCkuY3U9XB9hGot6FukOGEFM47xVRQqdTKFYVd0eaAID7M1waNqzmv
BIrM5G7McC8AwucKG8rc3Rj9N3jZsfohAPm6wHfGZhnxvACYdKGN5LEig28G
mkPLAovphEHBLj3mVAHBxTmO5/8VJuN9YxveklMdayKTV8zHjwFLbmW44O6W
9RjR/8VmUwj2L4mSIwylxCW3u6R2zAeCNI//AvjNHgFL9sHqMSCtSteFg2rJ
aOA4bHJc5tnGkw+JSWsDlPKe4SvIj8nLx6hhZtJmjHroKqfN6qjI+IcGYhzw
auvMkwGMMKWKcVYun4FzxVMmBl1cqx5ZNh19nkznWZzRN2UeNWXt0wiqQ6EW
W5ElmhIlSUlq6jgJC4V6KzkIRAJVbcyaTT/O+tynGbplAMO+0RSSqVg+7JsG
GPPgpFQgU+FS5h9I84Yf8ZlRPZwNuagJTOLTJ37yW5CO6ZqOd0n5gCP6hmXi
Tk/vId509CRURUFIIpdHiV12DpJ0lNGNZG3kghbhLPxY8ZMHq11Ms2gUC4rK
LAvG8uTX3b84JGD1zWY8UB/HVqmBn59oFhn6+f+HqyQbG7slOC7sIPHNeLaJ
zJFam8yp9VR77l+G0n+Jt57RXQuPisTHQvBvkcIa5FLp+s+QtowGtRmtBum5
LKnCkZh6e/RDt34P6cPvaTuzDdCcun8hrw7Vsm4t+tgd+XpYfqmWGdQ/1Ke+
ARbvE1W8l+gSi86sqj5Dy8BUU3dB2FFr7k67g5QpD2km0IdW5fYl3iJb2Cl7
US7pHA7qOAd58Jn1v7ASfBj2frn2QY02tzFnrzRmpLpK/zwrOn99ZsQDDnOT
DXwvQowJD/eiapinmpcUAGM7FHV9niSmpaNxpC//RvWjCxNwpjYmwwL5J/nx
6HhLGKvvF9OtkB/MPfJzSvn6pULXa/9zTtTK+kq+SlMjoc1do/HyWMVr/deV
7XzW+SjVA8I8280CP0A3pFkiuKf2m4ebs81yW3uGJXEGRjblYoaD6jlAeC0X
NqaBoZL19prfLcwNKUhYu0BchPx6ttA0usU4VctU1vseGlNcef8A0Ogzo5oM
OrJj4+dDOGsB5bsLl0ZLhCmFgEjewQiQ5dUZmSTspRWVOnUc6V5MsX2kJhIp
fDk+6iJSaEFm55aCmgqAqO0b530T3D6O/TwXx/LD+rJziepHjXOZ4IOMslUe
w5c11naxcKK0ueWl/kxJzaJO0CNe5kbtxnZX+hx100TXGk6HdL3w65rkEigl
h5PunqeAka3PKaPDZrZPSizPdXx6Y0IhvuBXjlpwRYjiKza076oWhx2REpml
5a4Xi/s4xBXjSdo8lx6wavBYpRlb4YzNB44Nr9yRYNDMzupsumbZn4tutMxQ
GkhUYVu/Qe04GcahdUq5q6EbaF3KLV5GpsBPRblbTgOF1ivt0wZkGMvfdY8i
lP96BE14ijMIQJI05zmroLZTyNA7jsIYdJPgccr3QSSkcQm07ld5LtIVtxEG
LIQOLj28G09mFEs/IXiLWZ3gmY1TFj1iiDfhUFhq3uQP+lHHbn+WbGQ4HQz+
VfCSqkronMMIiJsahINw/cY/h669luyZMiXtt0HC1lIh/RcxkgQtfz2Ewmh4
TIx7CnIFCxxxR+ZA3ETW4MkfVvvAveJohYXxNbgj17oTd98eX9fKeZnelNqq
LQf7wPldXeNGrsZLVIMLMCJyxPIVPnlHXdnfFWDVYKOPU4YEMpjRCImHAFVf
3UDfbk+owwsrBy/P94JFBCu8kwo3O6XkjiDQ1ohhEVK08MK+EXkYGGoiJWwL
EDzY3oy8P4R4d0KE4Nt7axeDl08fqyVaULtaIbXVBwDRNV4TVb0UfZdfiUeT
WvSzklRj2uSVn4tXQ/n57/nAMHoTo9unCTH17LwVA9Ei6AKdJ9P7lu+51RZz
6kAONsZEVxhGkPaAX4h05w9hi46tZsJq08E3PeEZI6Bs0e6AspPKQ8RHdkLt
UFn/dHXJUhbWO12mcyqcVZU5IfIud6DDh35gSdGeFxe+jW3KF7uDQLcya4o8
XuLRoORAr+mmE6BI/AK3Cblz5aR6Mibgbnj/L/tuUR2EnVa37HV4Yt+Z6V52
hEHnydCeZSQ+inrwKe6xFF8zCLdi2NzLvDVX17WKsqSl4GifF+RLg3S0vM+s
VhslUyTZalupCO/aL9i7OldqqT2d3hRvTyMwUL5xk0k1O0nyRoRVxNcj22SC
1cl/kKro5SiiOuNgj01XF6hFjXUQ4i36HXCrW4a+DfdmyctBpqlA7PDTPfvU
/xRIxog/m8mLfSfO4fgmU8gnZYE6vax9DUdq/kwvyCVg5ltxjd5zVoYK4nZt
4WCharRqg/AeliaWtJIvg4OjICK6knxTUixUazug2CyQrGehpIzvd8GmmkCR
Fre9TleuD+9CWSz2IfXv1kgEnchkUK3Nn+aR1pqHHCU44f1EjqbC5zwULOKp
RmFQtruyRGK4IqoJUCeyaDkHhBuJmT+geqcDcHcrV5wOsiI1ZQgo5j6qxXJ0
EddnGvV2ewEymIqLUDom2QmdRnohXfuXXCzzo8pPe8ui+JvcAtWwE9SnHIiU
ZYAbudGlISrxw5cCSo7hYJKOpmG2DGayTG5iVeXA4lxjP5KARMT4WcZLLR6d
ffIwG00UsIAiY7181kQhQ8+U06oZ3WvhXR8miBSIG6n80cHEfSgHlJ6/TI7k
kMaFhfnwPtZ6iDcntTM47SAfr2+M5ejnZc0LW/TtKSoGKyA2BL/pMQ+78ZtR
MqwpabXdC0Ie9pTD2jz1QaWAsnNGmSkP5BgTIh4/pHZjKxhEsGTt5WVQdyo5
lrMoxcxzW6RnSS9nAxtcY9y6DDd9u+HV1hYthVyY38GEygpUWskEVG/Hxeyq
r9UOPg+c83sQJ7Z1DtFoYW0bzXOGLNgIX+ayNvXo6CFRIxrY8G9a5zHlzEvp
dkkP6rlz9gZdaimBKqqjvGvc0Nr/BHEoEQBUTpsJb10k83HGbxIa7YWMGBVc
ya6UQW0f0vh0QkRfyHLgjhg2PO8wTLJNz0SL6jMIqzaVSCAvYm34ESnMA1lT
Lxld11zXLiqnlmyZpwqN1aNR5DUyhaRZxWSZW0tZ9xlCJ2wrSio4fkE2eILE
1uYjjJPHYn9O9poUr8Qf33C0iFntvo4cTCOHfApj7K3Nbvwg/cP1GtJR3gFe
HA2H+Svytc3qLuH+tPYUX/hlzpePd4A1xeO8peVqRoRI5k4zQaxHefkNbJSY
SU8WpX6Thub5h7/CNrZdx648LOm04VKU5ZWNl0dSkM7RU+2/wcILltp5FF7i
x+K8R6RLEokSiccVbvxs0Ij0JYYKoBWO/ZGCumD9Q6TqALMHjIAUxfU22vvI
PkyJABnDaUXvqaLW+X/4j1ucAhJdtw1d8oC0STJrx4Pl7E0zW9VCeSMQggcI
3kqMAoysybs26KDr9+lGpgcG7CWlTNjaDhstwHqkwdMvN6nh2LWz6Y7kYi2S
tFMFZkZjyVxVBvRzJY+b4PVcvxG33U0dTdHtIrRDrY71mciktwIIcHnYIlBb
fLWQU6S23r3lYGSBU5ELekMDIj69ErKii4sMx3ZdMp1JnV2ishoozAjR1+aX
fZ3QYglH/AY9DkbBextNT2gn59s4ohJEQ8mD+cxYFp2wNzVjyqjBOkrSZHeA
c3EUweEAhxZG1pmkVN46e1HrMmsaKwYqeEMi/wn9l1Lckjj/sCT+gCCvvR0G
wh76tuFLreL5b1hrD06H4t1DKtmw6PzeJ+G2a4Rfgkh8GjAU6s8oVYXqMI1C
A+uaAGR/erSu/fcLStks0D01zjdPxL99ALjpyQhzU925WqhTdCHNFiFJg0/F
rAtK3fJ4eplSDc3MWmd16elxP8mDmWo/b5duPdhJBpgRSCRnWUuLxNxJVHEO
gjW8isaWAbO4/eV52lC3VbRaLLv4gB5TRFiM5HOLNn9GgAq9AtJcAnC2GgYg
h+5zUlGf1MWG+qQov8Frlxo/XB1da+o9D3KxFPgwvy6D50teshPpfyD1Dn1c
4Wrpz7aOGeSbBbqcL7tqhn6U2AAEaRcnHV3x1PE8HnNu2KB0yx/a6lbaZxdD
R7Mm2QWiepw26JATwQsonjaw7PRFjqe+fXErqeu1T6v+r+qBh2BSjpzt4z4I
oIP+4Q4oeM9AqZ41lDXJ+zH9/itPIp4ML28BQBH02+skR00CLEfBpiB+LaA9
/SwRF4NV8ZQOY5IbnO6Xafq4Ecs4kBtOlPRLFK8UFlJRBVCwzWmJVZwoz+Xu
rGD/LtTzXQN/yl29SAPIb1UsLHvDCdjRn4p1XCAe9XyuIJKZomdIyxdfwjZy
KxMM8h9Hmq5YqZOPhFsM+feESJFrulR3il7fTA6PYTxTXdi0WIl+tSa7QxDg
hS3DC4T/1Juik925vNNgHlfL0mx3F7dglAtInqdEyfv/aCiqmDQuJykDOEv2
AbMXQDAysKttFEEImAGdkuv+4vWUrCqg57FAWEMlg3m6HqMOquLlbYaEAiV+
fh8I1GwYaXjhUd0hYnA1/Kmd2HSAHbCWPk4K9NbameB4+VReh9qaVD8Hyn5V
3ay2L5CZw47tSVvPB5ZrS4CcesT2c2amoBoVvxMdY0TV1PF+xpkcZZoRNqxt
+/YvZHvKNDUudn63bnk8wuQVIJuQYe3MUE9xcNkTPqyo+zmqNyUeWP0bbqi0
IT1x3MBkXg8WjjRQ4cK0qLzAkPDEkaZ0BTqcwhx1adtJTCs7lDxnR5BSby31
+hufNZzFlYg2Sk8INxDEPH8vGevMYe805x9+Efd4oVoZNSdvDP/x3bPZ/b4L
y5XlkDV5cJRhu+tzmqXoqm3NUlfb2dHyZLe84JZLAqHAv0Yp7YKbsoYR86d+
KETjuNLP29Q24ZF06PuMkrRNls4yZ79iHhHlxd7l1P2ijhh/tlQvRLPPH1lC
cprr8HlMLmPTXDbVNTUOq06uZ6OWT2rundTJYZXeFfQnJ46JecDfl8w6gBlM
37fClN723ZL1OyvskI0azJ/99/y0AEW9TLiZDGYlFld6HLa8eSHi77M2seIJ
U26eENF0w0y6zvk+l8V8OAU/GrwcPw6BIEQF2sHQSRZXqNgEctndXzJ0JJe9
kQEtr2NNK7wT6syYoHeNfh1Es2o43dDVLBPGc64fUGV0ABdl7l1JvGep2VQX
xXa+MQtW8cZQ10b9EjFVIR9kWwC/r12nQ+RfEt0K+1jnFvuDXmhQWwDNGCK0
A3HJdWyg5bV30t+4YiYPw/gVS7ILAPI0TWHTVaY3+ziUieg5BTRnBhj51uGE
i5y5nujPGMAIRiyGnsEMLUOgMnjpHikQfpk6gqRSZjuE+EZiyTR2qG+L6XN2
TXH2lvzovfvjWHNsL0v9rHH0Ci/Knk81EEmNC20ZvCe+EKtgrHxQ0LlAzTEu
d3PBaAgYVEMt6cnacpblvfDLvVp11jpVcYTdU97Sm8yluAjWSXhvoYVMk0Jc
8sbmyaeU7kjwjxviomOgWq2dNKAtRYPHIR+JVWksaWS87ePvDZdt070/pRGD
3/8/S+wa4i9pjF5352YMjfdc3NOvF7TIczsXpKj+5Gf0GVvhLiM3wvz2k+Wd
7YzZu+I/dO+FipqVvQGXrcQzHKEk6A/Uxor8XnuXUDe0tOn3/h63y5k99ncQ
cGQfiIy+dWxBwcBjl9zbhW5j5V+lTWa0ZV3tkxSakkSfYtz3CuQAytBzjbNq
nNSEi00GZsGLuQV/JRKtf5agghV6iF0QL1jVaTrzP3O/uaqborSjNH9Q20Lr
AspmqcL/PyTfMft4rMV5PL+zN3M0ogIE18Zi+AbXmQvy2CnQgz5ADAZQHCTe
RMBK8KlcwZxMscBObnTom1czsKEbfoNj2ZBCI9cTTFXdDbLMuhrfUr6e5+IT
+Cs+q7jrRKSPFnJIelZQL8OiC6NM8J40nEFMaaYiHiLaOXuhu98ON6cKDdkA
ufCEmlEy9uXzVM5aJMZ1h5UtrAPYtz3GSorgeYnwkQP6nLI4v1R+PKdWbIdv
Fs8UG+A6SbCYA3Gktwv2kIRfj118MnbOPxZgr3fYq162c2A3dCCTNubBGEv/
chfaDjWwvGkMWYuf+a8wnVHCotQCKrJLO2tU8LHxL0WG1Kui6ugUvi+rk3R3
lbuP1SCSa96DOz/HOWKAddDYvuXkWGU0oFwTw3Pcpy+ideYxuyEEpCPkAFhs
VLxTk57o/87mzH7zm5es9hQ0Fho8fQVOpeupUySBRimf8rbPCxSlDbs73UHt
D4p2Nxz1r3vnCY5W4hLujZvmJ6ya1td4alYCn18tXgDZUxoNIQSICpBxmgwI
+ldpUTmSAvVaNappnLNsqgvx4CqDHezR2Y1uI/FO771+LbsRoTeKDWPZdRrF
5ivPKAqgmWQEvVX6/jC6ST0DbsXwhzsXvnhe1Mx8LgSQ5G5X+abh7uTtMo8W
sdkPytrpfJuxqYYwrtfWTe9U//VbCAaz60jSxII+/jv6KMKaCjgPEYefcm3z
gke3CPJUydk6ynwQVNZu8jnz1F5BjjQWEWThSgA0yKUueMOCxCMBRYUyH9tg
iAtUFPpv/MH5kZXC2d6w6rxDHfZaedDZi4whQR+Hj3XFdE4Y0bZXZiWnjJxt
chJwkB0jfnW3z4XGQayMPq/DS0Y8+CelmLi6yYWQcaeAZOMpie41JIsBnNwH
zsT5Bvb4oUEcLEdnR3ZOVHe0IvL37qnG3lGsPdSYnPlOyNQe5WKWFBbMa3D+
8AcwCfaoeZlbylMv/TWsl/kvGZ/ECCOWd0vHjjJyXcOYyDLToGG3Qg746GXt
NL0MpVvqfIQivwDVGt8/zeJrnlKcyFUYvQpyjRB+wMer6/gztHRivR5Gebxc
W3NVoTJNk2+iIiXUIlJ0E7voV95A/9D+iEiEaZjF/Ondr+KWkfQ+vvhmFvk9
vcAt/TRXxghq39fMGfNLzNL8MrF0Of6Z3ygytHRcQcIfYNueU2dX0ra/D/FH
QrpVEIzNGamxS94iSp1Adjq/TyOoPTg+J0sHo5ZtI9urF0qmHS7926mLXWdM
/w6dXGbz9V49NjHNI+O06/JiCtLo4lcTIZPu8ZqjRoodAb5ftuyr/bE5Xh2e
ayHvPhp6Ck9yvAVRNB9ze6/u8yrefLr9abPC/wSGw5QgF2GHEJesdXaJaOJv
YwAKeYg0Vl1HYewtbXyJQzTiFOoSCAg5c3GG9xJ41jaZf8JcJU9pQbghmXhV
aORVpC+mNxMliLKPZhVa8lwpGF13pkiP+mooUSZasKU4gkxzNZbLEjK0A0If
FfAoUUF3Nx0enj/SyGxoB/cpTc75hsZtfK/z/Kf3n1kPdAJDIKD/xkw/+ZSt
Ere1I67hAGQtZcVdtUfl99S7ogFt5K9ARnlrEPvMG757Ls77kiWLRHq78df9
/zYgBAqculalqPeVqYZ+orcLv8I/uw0RSYwbArXVNZ3PYhClNiHGHNzThu8+
r4d9tzX8tIYzLlfaTRptKqulw8GxzC8tXBVjPlEyHTbBZGsP8i4oK+HHUmSo
4Y2mz2gYIvxV4ac5iZoXzkHqttbz69g95sIFHmvHZ//Xjk8x2NHHD5qNBGDL
weGGyji6nN4vJU6JFBq+4/CCW2S5IK0XCUiTjFLS5newOAbdoVGDcujsMjyv
Ambldmzi9Bq6HiaqPA0R3exdDCGbExLVbljUqMlnZWoOLDSIM6o0Fde/rlPi
icZqanP1he3HNy9kfLEOlGKYJbPrwk08I4dvRbI5YqlYocEBgxx6B8Enj5yU
emcGf/dXf7w7AD75QgjpgiIZVOwO7CB45brvFq+deEnuVpAX+Pdx9AxE/juP
EacRhwJgdu9s3iYe0wbH9lnT5BL0tI2oqpZEphkUc+bkhuaFCHMSK06owc9b
cPyObvtZcnc4P2siAL2EBz22FTJV+YyckF5I8Q09EtzkuHj4L/l/Pjopmpwm
QMPqbIjPUAlg2EqTx60cq2qFxzPJV1AH2Fsfxx1QuCslpViCHSRSB08mvF9O
ZKlqN5ZKDWFzgK8FTiX1KxDDw/sv78GmeCAK2228DbbDiX7TSGy0aSeYtBIB
SXZslbkzFgT13wKUIzFbwWOHBZJ9/CIcQGD52gIDhZVuhosXro+1lOfbC5tH
AKgnRvH4r8keJm6Ba351Kze7ocKvcwQj/JJ2Lzbt4Hm0/B2HriA7/ndM5xtT
gq+2+rVIUTjpo1auBHMugxom1Ed6QvezkGxMwdOJW3afgOAc01tJMKDDFlq+
hOO2cRpNSEZvQSRcQ++6jPXbIlggJd+ayl9EQnL5fB+tn6yozk+n9pqSIokW
z5hwQiEDBOQUT/kdLlzZ47rGzLkPo86ywj/dwE/wc4pZk3hV3Nx7nvSJ15sD
G+4jGLVXpWu3LxtxheQcakwq2xbKixfxE0T3GFRocqqxwPpcp8IKHEZz3rWb
ci4yvKrQ9cFlLH0BUZc7qOfqG1lfXndbySAP8Wd7qcwyz8vxQDuWnNdanWrI
2pEoFczKL+LY+t8xtr3hAvh3gJwx8xBEhmrXFSzyRi1eKmWlftTrQ5o2FG7T
Vwvr6LEDmjhml7YFjoz91nokhft2tHUrgtABr77mjr69XXBcyegVr1zS/Yxe
xm+PWT9vYgMc1ZWsTl+ReoMuatv05pegImWx6zp6Zl15bq6YkbyiRJ5sge1+
uzhX2J9FyE2tNp+/XMsMs+9CRSHjx760237Esqz+RAsCWt87qChFRuA+pL+c
izVXZiSNdDUZjBp1j1RGPXuNr2ALDsQvnZZjD2J3B4ngPItcLpap/6g2o0ux
ojDecQgHbKK7Q0UB9fYs0GT4G86V8UY9ZZ38PkOA3yaFviG3UfbWAqRKt7ef
CBCs5O+9V5jDfO4t4/nEVH08lyNvKnbn6noG6s/XrRlHHhlvojZ9cogwId+q
ygF13AfmG9vPTxNHZpSqJWC3ZTnAN9l9K9IuAZEAejKw6dAUBW9//5xz7O9m
pgoHMgLXUlklVpfqHvT3s5cAyZimgMyy4CcIvIsbLNJ9o3TpsOJ/w9i9PT3V
B0OQG0hoJ8wtQVXttW2548XAgn05ZH/S2ldRe97Xy4eKiuJ8rCx0YtgUwmCK
IPcgZwAVE0hiLukpEiZX2s/7UEbpk2P3LUyLy2eFPtx/IQGqtXQfQtSnAbdO
9dnHsgxVvR0GkBI0xAbh8Rv3zqMD1cCq33x8dcV2JKjAesgEDHCDqkNTIy6o
hCPKNe8DvcBAloXa0ABsMTxzOGhlNvtx1VQW19m1IY2O6QisMbIZzp4SgQJM
KTCTqM+pEokGhT/hZIVXRHV8/FyjnGkuZJhXv8wvWntCP/x6A1N5qJ2KQ3/Q
9HCQi0CDDsUXivmrKq7v29bJDkdj+boGz4OhiDcKe8seKqOEFjssEG0eSGmm
YguGjU45UK6rQ03ga96NQ8XjsHNyWhPQ/1ljTaPg/rmomPQgJtJTR58vRPc2
tL5ZcQ9L4bU1NwJho9FZQyKUZKBFAwLz1Lrw7xrrLlSg5x8lIyejv/7jGg7t
1Lbs2EKXxcqpdOfYqHS85ntsiDYRlMumKvF6ym/4GU8U2hjQ1gUPbSDIM0au
NOzKt1Ip0GUzNEu6Ey56rF6mghAd8yHfa7oVrqXOEQIxNMtFnvGGndD+Qyag
ZCAfK+YX7iTNyU6ATXeu93vbD8dOSIIlavxOElOSvrggi048gbTYtNEXJvZD
OWHDPcBm4+cASOgnyGadCL3d68lrwBmeQY+8Z8NjKThjOw/GCD8I6RfB9as9
Xs1uhO6Atjnj132/041+MyYnIxmvgKprJCWVTN+9bsfxJsnZSEDJc/5TAuf6
WFibdsWobFgz57qJbxZgY2iKvu8HexddSn7LHBuKZm4RpvaBK7zoixMG6W4l
qvgKN134BpRbCIeFw2fdxWgKdsbGWHGozLA90X+w0zGSUFpF+ggTdfVioH5v
XPwLLVek8UjmmQU34jfoN+vQZQD/kNWWTW/D6YIh5aq6pr2RMgTFsvF2PBel
X+1NLjRj8jQM8uxjE+IT+11RkZPm3G32OgMlLAWr7ku34u4PnJ48ZCZMsupo
K0rEK+HbCTlptnMr/xDPcf7dY0lMglibDKnt/b7BhIPcaYGmaxTlCYvmC2ab
VGjyVrB7wroGFrYwC/hoDarv3mGI1nhZNwArK74GzWBisPVxj/bGKMOVPDMs
Fp3FpisCwfJLUKuZ/cOo0MH5lzp/yDEfPyV015Uy6WRirAUML5VrENZIgn3W
1e1XUGsEWcjPIg03t4C/7+vUIgwnEYlwnuLrWyR06GK5N6CB3Xe2Ewpojr64
gVUZg9tmp+BQ6G6aVBecocMNFWUgsqtlpSUiEpKm8etBeE7rt6CVkeeOPZqG
FrA5sBR1VUaXWzFtyl6ab+4UByUCNO0jDPBuCVsP1oVcEdybNTUc6y3kd/JK
n7Oj3r/VJCwoKzYwCj/X5ssIfXIfQ/lneKlU8J2dgUHrrX+E3mne52yUsvE5
/KnSW6MNIJHOBjyQmx5hpQCDOrKRbr2C6KsUdM1U0UaX6np95/+SeJ1A3v0u
Ze4/90l48okrdxjw6gRCLIsC+h+ebgi4VZoE5vQGkqbjCFwBIwxMhfNCGiuh
3JlgXqZo02ulmRLtYyakuO3lR2az/bmQrSF3G+HG6Ftz0/1yqIwPdz0P+Lrp
q5nHFOZfU06GA+M5519QPiMHe7CyCoAGRK1GhuuiIxTQgIj92jpkSnBD3Gve
i3J3ZU1uhUlDxn3t4HCGTLlZZoHj1b39OpfAckgHbfnuFtkYbrAtbVQ87OFB
zMH4h+nVh929N85/aTYKdmRufbbqDP5zRaJQ4uDl4+uNK3ehYccw9szfpJUi
jqT4u2VKPT9+h782daY9Gp7r2CIsMp+q2UndExgnLULzoXIJcZwuA8cr0zIM
sabKYuXm5LtYY0k14fg+PcQ7Yh8OBFdleKlsUk4/8cVoLnY0HI6OY7JdWGqV
6Ur6XYLFKJBTDbsPaMzdb7NVqzLbSwhZ7VA9wJidULybmf4Z2TlF/Hqttubz
B0/OnkO++86KwV5CaSHam1S80yE3I6rzI7S+8TTjE+4oFbkohHImjqDkpMze
VZW1fIwwQ/I6T1RfLVJ+ZmrUAzseuj2doRKZy3gFTuiqOcGxB/mrieAFuNIw
x7NE8+lYQcjfm2Bi73XNKE+sycSWFzG6ZpZ1hr9/wPLXwFFMsU0Hh7ik8RA6
Ijf4V4eBohpZW/dWIiJZJi3GBdV+AhAKIq6msaUlmcDFxYIWfgUfuEkfSvUG
e/VsUkcpcSL3WM5dv7NEuE03qUfH2O7YV9omRaHnwrxML+LbKcK0EQXGA+57
jHirHT3CY/vSClWNvfE0io9rk80k2vobOJC3fi6m3yll2bY8Wqgj4c2dYXa4
baLg6qsZR2Bvne8SZE5cAokQGLfnk94tmqKtKQkdu/DTCHRfrjebbZrpQxDm
zeo+ulXFFBKH8BiI1Npn1HA7c5dqQ7ptooZlkk2+WxAV62oZ43IxrJfPFxno
Wc37areK7y4qtNjC7+GeYN5LPQ/IDr66yi4LPRodAo/cGefWwsiRRpIro38T
CBhpRJCack3yN3F3hFcDrOK32vMDI/0+DL5kTv3QPNMoKD2YfyrGTark81JM
mBkPK7Ehl/B81RID/FyVeGEF0Wu/aaSgBIHVYgQ7cFJtuHlD2awoxRbBCJ8z
jeIyIKW42QmcGbIgqv+jEVDs/EO+GXNO4BI5sPallCnm3WKwE1HMu1ymuavk
3+ZMVw5QMHJU9/rJLiLoo9H9D6O4PcoQ35LjpKtjld+qbugJBFCT0fTubW0f
gyurfpWUcapve5+9OTHVs1RrmvwHkhIPdcWGtgvZeL9362Vd4YIZ27AQNtP5
XmsXLPIn/vpXD7H5JvRaOc7oAbWQ1/5xmZlHF4wqd3YeUhUpFe+AcVfZW3h/
tvTLAyjX0myXgWLrl3VnZ/FrUQLP6glzxOMeaI3vIA81m+SjxoziZj6Vktar
1lvWAwDb7mwTlfDr7X7YDlDUW9rZRHy6NrWc04K+Q0DTsxt5bmieBiPXtqPv
yhKCHEGsak4PYGsMns/EJy1vR3SdKbyuT3OzGIbq5gRwM6DJstjGj7+4w1hB
uBzfd3gjCCuiTVgn79T7TJh+jGs9HMKjNP48kRhbQ3MqUG94/9oj6r1BPNFa
Va1jBQ8vZ8Ob8wD3M5w9dmwLG64LauG0tu80FCWr2wKo3gOp64u7Gdx3dalb
VKN3hQ7lWf+oRFRK0Bh3J6E8gMgGaSLk9X7nrpEMELdAbk0mfkDkjxR8ZxHf
E2HpnzXmgzpLX5FGEMMsPBxwoJjY1DjaZpMDCYS3J9wLYvTII824MVu87Xmw
VxKUOcI4Y7toCn3kIXTkRedQFqYagLP44nb8uc3oBSLLqQL/uUPvr/2HKs9y
Ulqaj6xU09jlxePub8q1TUO816z8DUB61qeM7UdZiVBQZGmNHBH75D8MoDPr
fUmfUJZkdnsp/v8pptYkyLY6zp8544+reqJP8Rxmv1e+G/MxqvJ5wlfJ3EfF
tdGgL9f8PyKuTchtZuBHVvHl3vEnGORCl6piL6kH0ohUS5P2zexYswRujafd
3kB3/N3nP91QbStmPpYrvS4tQ8jiHVUDTh+4W/hbKfWz1UfVg/hfLZh4w0P6
FGf1ZSSrdvuQIBOSEOvBFVgduxvj77scm9+Mo1wUiPsmjDu0mL9wdXlIg0vW
9/93Zfe5B/2RQ5IAv2sTuMT+Hu1qJB6SfKVtRkaR0FRmPw6sHKrQJ6u+IQJB
5X7Z/7jt2t5v9SaMFYeLgrvkRl+6uL9e305Bt+XCGjO9m5Zt+mIduAdDsqfI
W29zACxyKA/oCT0rHi0LiWvUHSiT5HLeI7fMvphBqCq2RI3yjHycI2TZuBeA
AW9B8aHgxLR2eskBsMJq6Bnb8ILiTCy9p2zrl8hIEIUabV8SPNAjNoG1bEBO
P57PwqL63UF+9Yu0EVjN5jLQ2L11Fq76n5CtvI+adiCvTqmVbKKybggAJ8XW
HRYYCJepcv5kXXDD9d1zdswgtHAYM5jgYtVX3yrq3XFEaKyDsgVTf0TYDBKx
ri02ZFeJIhEZ7YbpnAT91zeQzLDfko8Hbk0N3N1vDiwJYKWOS75x+GNYsZnQ
k5dD0X11HhvLtioU5U2ONBiMz/g0ErR2+YgvPFPJBQz9Jx8GQjEgbdYkQQwN
4KqW1QnA/5f0LnnkBAHL9HWcEl1ct9SKvgDMG/dGUyN7+LttAWGkHqG6Wo+Z
9T8JxV7CT3KQi5cXViUsY4PWy0TwPtwwPk8Mbe3zOb6F8Ld56B/9WMitQIDi
bgIrED6/r9u7q2vm38JSOmpXscfMzHAWzlPVqJCGPRZnr3RyHKn/CTcms4fQ
YLJNQYUbTQCk2ChxMk1KDRG3vLtsQ/J5GmLxOf/e9oqIvOg1GOfN/kN3bYE3
eGhIF9jgJEHuF3y0dJByevaeoA6O1ZqD+MxWWpQU6pvuQR5FjzTZS7p1BDvD
O4tIbayByqkQlV2teHkJUij1vYKhsp/SpMnpV8sOm4mkKQFlKT1scUl/kVMG
VmR07XZUIujtBIXFRK6I6cYNsxvEkP/P+rRqsMZ1QOegeTuTs7cp3Bsdanlt
eg3kXHW/VLh+xiFRLTQBQHthlG+IjttuECONkyAHJ8qQKL7qQiZnl/QoA3gN
PRXqrN2aIa8vnYs5X+6jnwXsvUnw0RItP1LEr4qrbxON0Zdd5IaDFU6ISB4n
U/TrNyAkrIA6nyXRs+jXKAYCZvkf12j2CmCYf5C3k6lMmxJIiV86amFP7leu
AsjIgTLwCHzt4xSUPrcLGskizgxrYcJhBdWU+rClQUMeb/zjIhjZtxh/HyJE
FPbzSMnD0S+yPly38o38uskLkOk9h+sw0fLKUR87yf5NggbN9mcIhL/g/e31
w8fdfVqwsEqQtTCqHJBA4Y5fN5tQnDIaTUUOfMcZfLRnomM3aVM/EBlQCWKn
o9rE3vj2JRWoE21BR1HcBCt2nBDguMQhSRuqIjIN9K/4A63cSksu7mxvvAIA
CKB4nn7CVQIYIZ+HPVcjXyKTSt3obrbeM1nhdJmBr6jMFPHjHR2mqlhx2HvI
e2q8VSSqQL62EGA2iHs6E+ftqtHv/n423wCMLpmNUGFqM8xapPaYUwK7PBsI
5J1KVrs/CSjmQu40j+68xRRKhTaowJkR7E0XCu14yCkjE6uFtjH5FTC2T0fe
BCy9aUTfM3ZGj1EQd0XvwVWB7IrK2TyWED2mqcQ7boqZ2Roh6F6m7nvkaVtm
m66fkqzhdvlApgQZJNgh5cmQTQT+/4cfMgh7z4TJU9vWhws233KUDeDF7XBu
OtzRbc24GDoiWUzQGURyrKlIMiYDJyHGKQWkSwo+7l+J2qX1kJuLkeC1a6Pz
58VVF6gsZOm5Bg4K9N7YCqP2yoFvyjwljidJ8NEA4JMPT+lkCiaWu1A3qEr+
UG10Esogs/v1ZIlfxPjFtdHN2gyQGssUONfL1KgDxuhnMbixwX92W9He7aPE
lTYeNG1Iu4A1KBlsGAwyh1OxbPGB1/DqhV6qCiCy82clQP48ViMlT+RQMbbB
1MmD1Acf3gHX3443GFLvruCiJvayOFAh3L7/3x8nzMGPjNzzlAMlg9F06h5P
gbA+lquGi4Hnd4hJD1GngWxRo7VxfA3PzYleCH9YGGw1BR9UhKAC61jc1OU6
pDJeSBtPNHaywpEBfrtCUqeBIPO/KNZtuQjoHiZ1UeR5AdmzSaV+tkUXOi2L
Tb3gCOJImYl48v3zD5K1KD/I0WwnoE+tkpciPtUU8XMnQf1gEEOJUQmrj3L1
ZqX2SrtoLRIk0GTytsAuaf9OhJ3iFLGc1abug72rrqF/qg7zhvDL3Wyp6i6n
Kfh2Omm5/inD26hK6cX9nZkCUmwzYhbnIdlAjaC8ypLeF3zrDQ7xPy8NPqXv
c+8pBoVEBrvj/2uoc1nfaj/TUjqAFJ1Tyto/YF3CmLB72SknbO2B8m5+ex1V
crBSakSduG9qOpNlUJdFnFeacQYCegXjTETal/+pboaVMtI4qhwogEDMqyC/
I6RnwALoBGViXGwe3yPkrcCbCOLtZBr3NWBn1oAz2lu7wWzp2gyEElYfWNNo
sOFLwHYNfoKh4V5YJIkYjAFp8xB+GVN8wWt4wAJWvwGeC2PgfRztU0uubUaa
gEKira8iUzAjmoEPZo1nyxsTF8mSGuSVH7ajr8Du9SmE07mmpmerc6wnphVD
la0oMKkRG24TvUKioivQsS6QXpU1CaLw31GjVaPtA7CyWRr79qjsRQ8Lhqe9
sGqCun/yAd0uIY15w3pdTrS1FfJurU6mPw/3wj1V+cu1p2pvPlzCSdpy/rqY
tEez8FNBthwVCwykg6RgKy2Sn/Nz1fTe8cPtyb/ufn0wgwtdbyH8Ceq1pnlg
lgPPcJsHKv2ijwyGmR56il4ERhCS2aJDt5VqHj12FHNts7+LR8spTghvrXbN
S8w20kpNsoK3+oRtob9W7cjsPBU2ac7USNed1vj08GK7tPiW9IQDfHrXr9UQ
Is994HrJk/H7ZPad9Ie6Gh26/QSW/l4o1kHmosszDYx51AdH8hh5a4kWzaqs
LEAgPTAIRZ1SNX4dT5QVQhGiD1P86oEJPjOR8AQ7EcIzBXJYqAHkpUQ+L8+P
h3C/BHjhDZsFVLqFLCLzRT3PClRFdVsR4Lva5SmTYhivb0p9aLivRm8fCYSR
ePC7nH2MvO9BD31+nsPZSmjMUkMXBMa5M0RumQLcrqh8CHCXHWFdkY/2I37o
74N7SXLt3JnYYdeoe9Q18+x8D2d4RZWfWXsMGJg41OcxVI8wAHOGD3oxIfR/
EM6HEouemdUhdv/4AvlEjq6i/38WRAfDDeQSYT+da8Hdukj72IHmbult7RPA
u+k9VmeqzQXHwS3J/nYL0f3cXTXU964voM3LQbndlu/ZY9KDt6EEO5VNvIpo
1wdLe6PgCpzWbw2gxqzaRl3mad69fkqh6lC7+6kXssLBYd3VMpwygjyzuqnD
8RyWZ6kv/+LhgNc5+SI6ngUrW0ba7wMxxmBhYXnl5w2UAjO6LaNUdvEGVqho
phztrdWH5nUZlQPbc5bKZYONjwPcrbUOGpJbJCPX9cry7RSHC3+sqB/J+aVa
Z8+2ghfa4qE4WfwJHWc9WVu+O7fMAvBsbMPjP9whv/QN0hxomCMUXLFBcq+q
4N1ftZbBcmQw0hW0So7Q0JVSO4hgkJnKz6xq3rWHpkBoZPSyyl+o+USaquqh
6rN/DDkeetWuoIGNGJOy7L5vF1inZKhXIV1/SySpKksw90skpPzSBlwVrx1r
Jo6f8E/qQOx3Y7uYXfTUcLOu5E6FON1/3JBiJsLZL6eLra351hwKMvuve3H5
01gelOa2YPSFG7wbYbhKAn2OfvyRmtvNuBSVdTTLpRcGAV6os0TdEGiifcdN
MTd/+xviheLWJpW5260B4Hp8OfJlyT4WertMXq6HULFsmYDJy96Gyscrr4hF
HvwK7ymh4ki1MkjdkhtcFFiH1aka40cJWurOrrBPz6JTUYSMzJfMw5Fw8OSy
YPcyqnOJqUMi7T5ZjDrC9ono8y0H0UTy+QYqPeleeT1mVVV+dDrcHipCA8NN
2hIiCHGL5ZZeOkjqtgt/uuMHsysfEKIwAo0wjppnRSn0BKBfkxIK35Gwk/Xy
1WTwv6cSWCDbSDnYXcBbQvNTNWYNJgTAALxi6gQvMc2sLUDm3mSH3K/ZxBam
H4V5j98I6fboDQPgCoBMFCZ/59NX13qcucTEOMMbLnE7iFkgP5aI1BM2kFGg
B+5wQsWFfFfXL574KHmF8ScHSah9v38jaLNbRP8dxDV98OrPeuCiWyIqk14A
radmm3oOJv+pIYZlZvGnW2i4Z00h2qDCKMqbZT7wBBy7etGvAAdAdSOyiIJA
2/sZHi7ktSaNq9teNPZFQq1fPwvADMn1u2WH/0y4C38enPzlTPkpevRPebJG
b3aQ7s7rVUpBqfDNFTBqmNmcRD6Ul+tQoWcM/ILhG5GFF20Q+blarZ77BjzM
DjOYvhL4etpv5vsX3p9qy1+0IxYXTZce6mx/DMQ/Z2yQQt+14J+bldj5QdoD
tXGhOmJzWdvbkj7G+IXNryFnrbAq05x5IqdglfiQoNK6+d1rof+5+i0WQbRM
omvuEtgEjm6PgHERBkg4Usrvt2Pwl9A23wIBvjPuuDtlIpMzhAc5cDbv54rD
ymbyXhIM7UhM1fdMiL1105/WbgJk6cvEi8Mu7UTOO9XqTSSHDVDaXM4xrDFc
BN4etuef8cb6rvTRd/G0xrvMgN3zDUq4cXYaOjKHM+WW7V5ia92pVzI0QOVR
rv/jrUcgAdOqF0OB7AASSdrPPq+hLDz5phhsVPh4unFOiJVY3EwyEDW9qB01
tIipMn3q5XO+R6osmavy1Z3KK9GXih7G+1/giQdweKoROFFOYH4JVUrh+nuA
szg/FdDOqfHaFndcBqsEBBjS1pvUVucMWYfZvpiRUGevc2kXNGSN5xGmoy8t
T4erAVnlMBxWuVbe6+2beUk9epFEn2L9Xooa3V8lFVT0Nvs0MQcyw0GWZu6t
XLhPIE1/OPOrSz+5AzF2c5VlhdAjHo1thzpS68C7nccxl8qG4X1PBjF2RQmT
merfpPVoKrDoHZRvSzuN5OvCscM63aQ5B1qS/uKry/sQTNuck3Hm1CLtdRi0
KjSFl6oHfq+bk+9ZHEE0RmATuQmVFIjrou6cQ7sPRQfNzIGdgCph2aMRM6w6
E4McEvJSPEAc/kyS6yGT6S6PeHgbAxKzN9pzMWSLehkFchStwyDNit/WBVIZ
3VCG9g24tcPt28k7MlTVhaB2idUsfSPn37+s2pv/opjmuqswatj5IU/ghPrN
bPTO7uyr2ButsHQQMTgWMjMoUOgEdCwPcOZZiB8i5Gy9ZvgQEfF2Fuplt0GO
ot+0LYTJmh98JAO9JM2xM8J/JntEpw0oQl17ivB8P/XLSCIdKsr0aYNtHc3O
nq+M08xM5bglqFYAmt9nCoyVM9A0Oy5FckK3p2h4wahCxxtuXnq6EepcYCVU
7Yn4R59/lCBnrtbNX60onXD14uNh3DlNCUqfcPH70E+wXGP/pdkZoU1NbDhQ
LmA4qgYiNoHkCmTbbs6NXMc7LK7FTx6NrV6dTq8hQpq3h/ilwoqgJeYUVu93
xSUlvZ5Zzv9F5QImxF2dJ+ZUHgcFFoqqdYjegk80QkdxVFeoNFduFSSpwVe5
K+F7ZrotpEyzM2JqmqvYPjIHBA9s3jcbOn1vIeYkTBbx7WNujUXDz7sHBPWt
heRHmfx+RWSC45Jlan2+0581kqjRGtrg0ipY1LwIYl4UDFQ5xKdQliKzXKrH
FZARjg6Lu528YdRTl0/13/3SEas+HQjla6JcgZL7N/TVlQ73lv75jWp89Jm+
TfARO7FDsRHT3s4bJeUHCH2jwNTy2MxzhL0YOK6QQ09ubqigiP6YDARvvZE5
b/hR/3/12I+0j9m+dTSc6D1RjZkbzvv5m52aM0AZooc5+egVb7/1X1Ntf8/y
H+dAy5PS27cw9wUUsXv67pBgbe30hUKJcbBU5UUqQ43PlfpGqGpwWcddF128
tMl6KjExXpGNCW7PNHXgRRPVHka08wczC+UdQtX2AorhDbZ1A1wzkULTLYZR
KHjMYv2uDvlzrVX1e/ocq9hcvxe2ZJgy8DEk7vDFUBCbcoSB7TPbjN9ZV0ql
Wk3YLpd/d9LFUXz48N84NR9XPHkxdeecf8GYf7yyeGlwcMwTgkfVbihEmKqS
Fttx6PlY5GEFBM52GxXhACrDLjtFeyV6+04II2rbi3PU0SbMxyC7FX0YP1m7
5zAab7yMOHr+tSldz9m2+Fx7XFxidMqDDk9xBAUycpWfiLk9wY/eJU8tMN7Q
2CQZwYQaCJc8jPfwNgRgmdE4AYSSoWUEw6/Aar8WtdDRDaoSS3ri4cXczZCP
r0pdOV+Iy+waN2qpmGUx+vmpK00CxMXAEVpwxS05wzy5Uj5Eiy/ul4Nst/C7
LhF5sh27KlArCEm3IRz3thYK367fkgXyoQAswqMg3O0M8LP7zXt+QlcMg9TM
OOH6VD3qolkr4kuYAsuBCfQj35eMIm4eZeUWNrjcdy8bbpqnigJsRtyMDrm4
VV59cHqdXewqbTQaKGa8SXkYrlo5Tmdfsd8GpbgIzbPU+PHlDicm33CbmFlI
3q+P4jggZhpThfL5qxIYIM5j9Rhqemc0cIyG3fqWEAI9z0aETWE6emS+9Mf9
aZNL1rcdpMcif3TyeNXX5Nn3PVnAKeWNadn6U9cvtWF4V3DOO7OQ+/1ICI9y
zs/1zQbqFn9o483SuDwz8vV3nJs9zZNO3rZvoAxdKbh3J3dj+QSGOEuznGDb
QHvFfegiZQN6TtE7bWPVHOMyqVsv6D2Pv4g/EIcTozhjHfqJOCizGV8m4IfU
XdNW8I+3pMrJteVx2kgoj6yyJqFhzr957JX99a4rdhRBLGVDRsYmJhiDF8ko
gyGEyVPkfIwKA4JAxZamJrkPTUdgjw/S7bQTlyGayRMjl0VYHGHKH6GNacQs
VQOKAweRinbbsQh6vVi9NZXDLfjCKGaYmJFWkW7RPBn0LdxcBVePBkxkqDrX
HF0mJzBsOEPEsTdaUSa+RYZap1YWCe3Ah9ANZISylI0HywIEjm4KsyUOELYi
oOKcsHgVHyuHlkMTx86nvg3oWrW4vfHE5MiF29yNroQ9h25hwCPKN5wvKOFk
tQrErZ8C58/n6d5kV3vCBBcu2WnhESIiilyS4xXzXfUUqBd6OfWb3SGddTS7
iNJnmrBmv7aIqv55RgdBX2EnMRvkszOhhwek0Acq388zx17Hggka2Q4qm2Vq
yhX+FrFdLKjYcHFsjsbPPEN/xfM+8a8XALno7iWXXcvMWkqmHu31z1LmwTxC
jQJK6vE8R4eaiv38plsdkKkCT+m4THzstvCzf4azNArKHOZoHM/TDZt4vlDv
RO8zqXroPSxKlZt8sbBV7QU1m0/3ZbcvG8NuVxtFNb7O8EGX8RNOdcKMn9vP
5wQ9gsBBaVEGtudaFRXU0Pqrj1zs1TQmMtlMidz+ahzWjipPEXskyM19wt17
+vJKcN2ju8zUbhqlfeULDgf8Fnv3b5QsJ4vdDFqL1rLVs58l1/sQNUOPnhW6
97yTU75YTLWzBi50uN/Mw1sK1tgR2aTpaBCxYFoF8RTvaRxrCYB+ZN3cUbJz
/HYXWbD9WhOYZdMhLkZnus5KvwtOtUgaeFYF213wOFK3PAXna84dA5r4BmeW
rZz1hpS1olyFiBCFM/NTIQQItqpwYEc1mijU0X8b8pvh8FQUk/hSdwgmg6q/
sUWctTWX4rahYeitR6zEA8xNYm3P//ndT48czldz3ijc43Dr3jxiNtRcEL92
isY3Nx45oQjy/M59WukJtOFKEiwZvbeRMbyLPcbRFcf8QWZ/hjWbtXwopG39
137FJlkqMZssMeXd9n5kDogIPmvIAgwNA4fwezgn0dB+7bCDKl5lHg4SxC27
94qakqN+9BP9+uMsgOZ5/0j+mOn9k13LJIDKInlTjsx9qr8Zx/Dpvbb0wSzH
1KZjaWZOHEq708loruwBLYZJfDkzKeUDCspepyOkonzaQKScb1OG+ZUzQJkT
gg1u966N9qDSy64iHTVOVAbOYkEGUDdoOEJP6dvxJZBrzcwxehp8WHBcPMV3
kiU6P8wSYbon9END5j/FmdXqiksq/eqJLimVsoTndMIXjWSuIKRmZ7f3pz+G
KKDMtDP8vczKGS/7VJ5K+3RjmPF/cfJmQFXzk9zKQbeDTXyldlCOXCX79S1I
kzDhzrxaxwL60amxNPjI4zr+IJ5cF9XdM0ngca9l9qqDlspRJymUsjX3XsF2
wLCKW79vdpiszD+LcVstDj3DKL75b+gWFAsNCA7CD6PKbfTUXiQ51WCrENGu
gXXWO6rVv45lUKWeyQlUjFziihQpnyELGoi+7jxHfjzPMJCZ8D6hZrDNJAlt
zA0p8q70IYrc8RGyIZH9rv0fnRy/lLvR6fIg0+BR+FKhBYc6nK60B4YHlp5D
rRVFoM7k/HWc7kDASRDcgON0H7qoEe/Et8KE6MBJawkKQTD+PilARuTMCtp/
cAT1Uw5gGVZLSn0TazH0+iUaDZznkC1WwVxpNkCggfMX8mUVAO+fBB7KiFwu
442PR3nlM0STnNRKJ+c/zrfGvnEfigzkxowscOSMABkzps6plugpKJfAOWFh
2myK5hIl2g2OqDSdg0W9VPZgaGNrOdNxKBnK674CXOaSv/uD46TpXeULsHYg
NpbK7H+KI71+fJktGT3/KZvUDbF3djakjPZaTBtTyTiATCFVh5iPREKteInH
iY6cpBECYiPuR8vc+DVDfvFObrHEUwsA7s5uoBRzjObURvN0peUzqpVCH10R
ECaPh0O36aOMlxH0Tuyyk2XYKD1bX8KQqUui2hr2cxmuieyHC8+qeR1WXr3X
tbxZ4XPwmhTV2gR4qIeIddutNS128mb1xDJ1hqPjsDtBap0dtCLmTL73Dt1K
3wSz9YLb4iALY+zD0ErStZL8dTOh8xLwn5W4YnMMKVD27Yh5piLQNgb2m4vC
La8fH5SBlxoOCSAmPZUdcPd9RVUEs4i2aPLcq0YExG2onykTOr0m2NbP1p7g
4Eq9P5m5u0ZYJ17YPXWGFHNVHWcEIOO98jdNHxxpMLXji3oIygj1kih8B7+T
aI3KsVUY1ygDdI2zoT7NYMIZm1arWssOV9yuMEpOyA5NMQ0OClH1PmLac+hm
KaAYndQv4qJep8mMMG3gqWa5wf0e7aIoV20jUyi7i9q3njJP+9jMhBmrUp6d
1iKxl3hfMSgFcAX98jsuOby5MQ2J2z2/6vRrc46IJrQvF4mSZ+h3AWuxxBhY
0O3gBBGMxkdGwkAPnKjzSjdmfN2/bFuh51aFJ1fjrVvuFeUerTn/BJXW9G3P
PR6pyKsyjAnFj0yy2hK3Bp4fKjtflXABfb1ah/suorL/vnUlEuq20gFvXG6N
9WcJ/wtD7I1TFxVHy6GT+jxNUlONgj+ID6FCxnlTq2l5ztnqRmAFAJHJo6KZ
KYB5BV4w0prHIhjkwcUpCt7TiTZDV7SsqxC7SjFxajk7sIO/kkY/wOXWOVUv
t07KYXqnaYcC+gJV2ev7nI1+fxBWwvwNN98/JGXinDmIx041ZmkxvVKTqN5z
FStQFp/Xl++phUHoKAj9+T1EbF/9b07Sw9UFtOfiQB6BBZxsMuGpgZOJGhQG
tfDi6vdoxglCEzNwnIJgcDkWBQ8qxEsHzvZQeO8YtxUtYW5SPd/FwXJX5Vhc
kaCk8w/KT0NskJbOiiTMSU+X+rjNTwwKZia+cForbkJQ7xZEJ6NqTN9TlLxm
i7GFiZ5wBsHfm3/D6SZ07V3hMu0vx6pb28Ni8bJhWiwd0g/8RyHny9QXd0jO
43peExAhsxnYsXTO5pheM2erkzrnq/mYbdB3RmscEZyECgAHTACqQUbncDyT
UOSvUN8WEe7X0TOyfk0uVYsMAyeNz3Nv/AcwLvkc0Kd0lbZLwjMchYtyORlD
R50KFn+X2eS3Sjk5qm6KLkJ7fHOpguCxUlB6xdj/+HWjvP5kmGGRAKqUV5R8
xu5APYIGwdNqLfDLfmLiWrzq1wgZrmLRMdMxxsjqBuWQMq0YbwYJXfmVOh1X
cjmMfdWwQdSSl09SC91K1lV9OoLIXnsMc378FO9mc14TI54t01XC9GJhQakH
HZxni/O/53jiXILUJj+9rtsk1grhO/fWvDmLF+KwU8AlGbzyk5A92l2Jj5Ap
umi+j6H8BY/2Dp4MKHNDK1hjB8YG3w49is/f1n4hX22eqbQNUHqmX4GxT95C
N15Lwu+2BIBeJDGAYyJyPs5aMAfOMVxbP/f9oS6ZKSTozFf+qA20eq7WujD2
9j2oW1f9RxNV4WPDaafYjvxc9Uy36nq9u171+5SAYfP1avp2gwNnIRThkdbj
iajc6hmRTV9UL1+6BPsURTL8l68mxgG5HpZDSHh+qqVV/8KnyWvZhooUf4kA
GC/fSk/RREIFYBEDVCLHBQbomYntcAJcIGNyXQpCxSOmkohkY7cZvvPEJWSO
fAs4/rcSNvGBg5xJhXeE8nva5judPA+LiipJ6QkCZl1pKV1eKg+0hmTXvkp1
566amQRDDhRGfDJtPN9eYx9XFB8q8u6M1dxmp14VJhTsy4hUEVDc3l487AbX
EWiV+iVyVyt8yij9QuLIFEOOoe6l7mebSdZq9WBhEiwi7lvDYPvtjzExD1Ec
4K4oe76nyKq9bO8EjfjBczYmEYdFTOZH5KU0nTPLXA5CX4yrM/wTyEyBjBJc
T0r5xAzKX4Fj8RE7E18kqY///oLHOstgjGNAb7BiU86UJ/kvTDkuTfSYD3xs
us/GZCiEVBKjP8C7iSeD8dHcMuyQoj5zNq/rbxHXstNiZHm4N0Al+WiCcbhV
3RUMVNOZOIIEP3fosF61XmuBBTQ4Z+6JNJuanRiNlBbTjldTRprZ+nk8Elt2
yIouXCapLeuUdmFEIl68ggAPMkDhnTiqn3hdG7puVNFwUED5p2AuFNF2++Xi
7z35sBaio/d9x8zpO/jhBjOTHmXDqb7uoko97d3DLTLad46wgo878/PadA3T
sbeNCzxx2HAj+qGBRV/9ZNnwiRyqRFTrV8eQibLZgJyE7UcKCm8yxT7pLmDv
yl9epQJcxPaiSlAdv917GZ36ZMiIZ2S5fYycFI8Kvc2b4nk5RmxrMP9ogM06
gKV9SrNMobqwpjvjurSMHxtYIAqpsgEqFVNjc456bSBHnSYRlj+touM64QBU
en1z2RtEWCG1MKtBwF2/1No2j4hb9Wxg/roywyF8m7QyM7vl+2XEogj63372
PAYopCXXIJVSv9DUqTj+SD8YreIe+R3mp3J/+np0cg3iJUgSi7RSwmaO/2Rh
1KigKcLccZ7Qm5IH2uWBH87dLDc/o+FOqr/yykM06ToXEKgPTZQqHxlmZktE
plP2EiGhwZ5RRpm+ML80t0FdhzKbpR6FE9Pkld0+UUSUnko4hTiZxeTN3E3D
QFnwaOKz9HZxHl4xeWyBJD4eJHR36gwjsg625wrn54Zbnt/xwCbn94kk6yed
hANZz/hAKm/Ya3FkWMWZR+6GkRgxNsYAikLLIWfD8SiYotocT7JoYob9ShMU
kBhik0wzQlJ313G7nyf7WgXc6+9M4JvfZzVa2QVVX31brl96+bI8we2vXs/B
VOFMsexfbRT4jHTNWD9zSLGfHO/y+ztFs97OKmk9vLAqXD7IffYnT32gZZm3
FMTj5irmnxCnViRBSSj/M2yTazoovlLr+Msx/+Luq1D+mAgnPA92XIA1yeMJ
u1zcrPHsXkctNri5gQgIkk6wZ2IHXmzQSRJQIA1Tjj3JFv7L4yFpMYitUZG+
mZJLm7oy4AfTeZZZHakE5Ecc+Y2Q0RIdy6eL6zaravb796BBPk7TlbEaherR
Er5xB1VFNdxNd2Untq3QJtQwdKcShOLcWsv/4WviuoNcXGn03XtxCVQh6QjJ
R/1qz/6Pq5hAevO9H4Bt1ssXxiJhSQ7MrxtJI5BzYt0WYgygOjQY3Bulz2aU
GQtVawKhSeMSTkcDSbiR2m8V+pGbYt668F0JVuKOQLZHEChpA4TZuMuRGhWy
EzL6fe3nIkXcxUT9hjsiDxvWKYTHaY21OKMkqtkN2nKVrJmCK2yoIgceP3PC
+NlPTHPTTwFZvRP0rU/neMd050al/v6QgWC7tyNvfR6gvETnYYUCcgMu78Ks
ct4aspe+DlrSekALp2hBmeuQXoh/kUmCplKeAPn0dY9e+edJbV8kmNF8Mc4r
UOzesPTENrebuqi/CID6oJtn7Ti2dcQJJoLq+dXKdTcXahtv0iAmct/HlY6Z
T6rKj1hg5j0EaOkHypFiGtx3OvNlpzI7aMMIZYhyGppA/yKIGWxcaiLEVUpB
yw+kU7b4kGnCPLG21wF2lRIj66IUXnFrg4AKj8P1IPedwj1yKqRp4fDzxwc2
X3ZRoVwSc4ER/+I3ZfbeneZTHYW1k+tZyEl5CPU4rtQukn/Rq7U15xR3/EKV
YaQidkZDhaRciRRab4Q5mr8nAoeG9C6747wbexUUxpPSBHyKj3Zb0by0aBcp
8qrJx98qPfbNJovMgKXZoiDbetY0ICTex6rLCXrPtCdrEObV+FSMj0GJ8y72
ZtQoowqX87q0UA8Rdh8VTp+sS0JtsHl7KSJOXcF0YCYmH4Y1yW9bRK7EDH8q
GfSFEe+HEu8hx/84z/GNHM93fIoVomw67eaK+15EozQ2NbRmkFh31JPJvWiS
KFhaYso0Bufj5bu69TnhxcFjkt/Be9NdcsfWWy/iP/dME4qq64yJmfx2BaLK
cflsZKNz5P66ze5+4mRzDyWecAHfg05PuP8+8PwpozQceLtOriHTyv4rSMp7
po/hySIDDHhClO5jShgfotmwbBIB/iYPhtcPMY5TK+bquXJXipgN7YQqtYPu
bOveXGCg2YNoOgMP6lUzoWVFeFXHvwRY9mLS9yOedK3Y+hu3Ykfn/DDT85PK
ZvsgjJrJcvw0acGjA2KSooSgN9r3HqSTpHKdI7URjFm8n9Uk8cHDXZ3PjxKY
o/40MsXHQ43PruyfWz/fg7rmljWOO7IYiAdZ8HZxR0Sb0Tw06ga1Ccwhh04P
NQqnW8jrj30wkyApkO2utMD/pBhdvfs8wj311Adz5hNtPcD547vxYeGp3VbZ
nm2YOYh6MBoR2FbYA4mQjKH0KHmaRJLAJOOm8tNmaty3/uvQuLKBfPKU7Dlz
8++X7A5YR51gwZ9ZMCGa4NP55U6YJ6vFDdlUq+BmPXdvTGCXuWE2EUaUEmCO
3b1K6nGYQf0xbDNZmXldgalDi8oKzdfmK9FEFLKyqMnGSf91ACaDwtWxjFN7
E270m+H9ibxFuFZ1L2FUUtX3ZQ/BYRqiuPJZDju9BZ8OAeCCRmNaCerZdyWd
tux29HpTB1edy6ACtVapQ8FV7Wi1VLtbKFOqNij7Gb13z2fwRyQpulXXIsZj
my9pL/gTaVap1UQmeZrp1pE1SXJwmxNxscwf4E23TaholXn9DXjePhg/cHh7
ZMiiWc7AHE1sExlETIdhiBnD/NKBA5sY8hvF0KixNAzfLjXtoRJWh4wOmN+9
jXkRai/kflFqJSBIGZw5GjpRvvxWTffQl7JADqYzeZtc5AaqeSz4a2dqjE8Y
aX4qNOE7yBXM5CzRYLbndXfNw8pE6Pedtnfaf9IcqQzeaM1+/WM57UE4dvoV
31GT2PDCRDaDn41S4niymtgyLBoT7fiQQaINGhSXuO8d6Vxp0cf8zBJq00si
ol3GG4zaGhDgasksnPZ47MUe6Msaq7rtI3yANeE9SitOlKMuKBSkJ8GDhglx
NFSyH43jWl1h4b6NP8nWTCYM75MBAx5KUGpYCw5fqdjct/hYDRE2oq9S4QxK
B01eCzk+Mcexjb/ZI8ksmc8oggvXAcRDI49bgxaOxkdICFr/oDxaZ/RiBpOr
tlbmh7tofwOupcwJrK3LgW/pl+2Y7NVmDhxKTl8xXGkfeudGjcxJmmNvIjTu
kRvWNIkgIlK5q2yYR9bGOl8lojl8/KfrHN8lOrOIh+o9eX3bapubrkawy04X
cZF5PkH3mKqBbIxWShkrMhFf+Z9VQpPluveCJpvyDdfJ3nbga8+VZrCdC3Ly
LNMnh94MYYtlDVZUDwtJ4GPfHjbSyyrNCBK6Jgk5Sd3fFjGjAne+Axw8HCP0
qGdmYylYbUUaNtpLki50EPCfd1VH/9La7xGwZHy47enSuW3UT7PLnbYtGOlk
nP1N4VzC7NXtgZ/k90sxxPNTOq0GfDGbaXgNIHgTbLpfVcKOla4sKwx+Wf3U
u0HeacIwLb6LfoiOqJjKTRH2bVHE26rAQWkJ7u/J2z4UDyURSc/qHZs4pARg
5h26migd/lFwo9qsFos66QXzUeHpo0d/PL1b+1yngHOgRFzhfW5+XZLheaa+
lGnF2I3nIhis3O2SDYvCIQIMTPZZQfHBoQTzMYmB8xvA+2GPtzHhU3VV1uNS
OrVaUFaO0zReyrqHEm/Es5leWB+BLOxiJiSyhXbVHyoeHlUKaCYjd5h4vU4H
14i/PQQ/euvL9gC41VdZzGsKb1zIEgqqKnp7izg1x3a+MyDJIlaXRfciTIBc
NI41K68OD2Gukb7XJv7U4un0cCFVEtdRx7FZMf3Ir1SUhUfjbZNOnnyTdING
Fia3TdSZLnLhmyE9NtJuThuZ6/ooikBKGF2pV4zTpZMRaLhZ5gwxA47CULaV
JemImlyh0bGMLslE6LH4l9sWaw5plumoQTnoYwFIBiIPJJ5pAE9BYhIHRiA2
xNsG0MXu9L+L2E04tCni2s7PatB8IrqPTPXh1PHORy5AFBS/via4pJEx7Qis
aoZQePhyYSkCGEYepzrg0zSArULPmd2tEvffs361eLjBAp2QWXCnkEtCLj5W
Dv4vN9i1LD+m66NR1wruQXX/sl/1dswhynt/vEe48oku7o7lodOz59SElj7c
VMKCHlX5i1k7dvGQVIW1hjjtCwn0rI/A5nNSDMgB60g5q3jQdkdxQDq7sIIm
2qifunbO4IdlEChUhmY2Ufz2pYAx5vAJ5JUmDxc7K/h3FRkA1UTxFGLwRgu/
R/o0p2WSo8loreX108IvBQv+7rCzKzCA8VdiP0Gv3BxP3X1D6hTnhZFhv6AI
Pt1O5cN2yjNnAw9BCUUDFUUQLWXTm/nUlAkroK/CZYAlLsLvbLsh8yMjhydf
v+jWc6stGj6t5dAYjBD4Vb8NfIXtEW2VBxsig173YF+PRH+QcC0Vlxij9kdH
y36El/MUAjqEWncZjdrme1iH9Y8d/tnsujbBp9phXga6hPJ2gE0WkBuN0eFg
rXoWqWghobR/eHtWKBHur0M4Cb8MkkSxGza2Qri5XWGNbC+CF92PHu4KNpER
4p4yROqHYr8dovh7horZjEr4McOPC1ZuTPOuXXmiYJSrFfRpi1aP+brxO5zg
sKlS9OzTrI98/tgYHfTrnjIw120VeIC4Gbb1iVGnXMnOckN8M+FjZLliwF9/
VlvM5/QKfdG59rgAHWsu6vZ8QQaaaLcdPAsUslrFpJg3p5z0W4faQ4gfH7gg
XB+2CTSYOEUDWSvoVYh73ztKdYYCK3tO9Wc313/8JF74pdsRuYRPpMKFw0DV
jwUSizRRZuNRb9smZ60iOR5ryNgd1iczLvwm2ZNjjufpiWtf1YpZ1jxCOMB3
l/8q3fNpQ5q5BGg190G4FyvE6VetpgYNMK3SbCST6uD/xp88Cqwr+PaCxrLP
reiP6p2GMLDQxmKkvKWkF+tbEYmvVZM5bwHaIErpd47usp6On7Q4vWrmOJeT
vWMoiFQjE1RdG1jU0gzxgjGdS9CAxNWsOp9MxnVG2OflOo2wMnzcZ3U7UPzY
az0nMBs4253/kqAKjE1a6MJCO6/zt9S+4LAywS+wwd1cc07nNwV2boov11Wb
CfT8XWt+SdLhczkApXhM9TVvKRKHoFlVJvfqbLjTwWMUewnE3WJgDSMWbrDn
kMEUpBWdiLbMjOwabWr6q3JIuEnR+mWeCQ0ZJYVB0Sd02ZRhQCsseDxzU7QR
qNDZYo5r1KhYbCqQ2B679Dm1IQmnztZrWv8EpSKwSCP7FhuMcrqh5DVmMdOB
Ga7DdGdGthaQDK8ZEnDpueMRJKgVzI/YjAAnp9OtlY+OutoHEljrgBG5wYQM
FdzEn7t/5NSlCdYbMEY7exwS5cZJfWMNySjdaaLKOoOrLKa6oIAHxFb8Snt4
aXkhyBsMsLhwdxzfH6+X44Hzb6zH4QG0FVGwMgozygzUDEKt8TISgeG6uHIl
mdxENPWtEznKUnqCIa2yut8U9KX2v0zw94yA9fBsV5lvgrj/AjkS+uVpcUN+
dNtsXAZVYdmhTRbqlPE4TCl8Ish5I6eQ0R1dpat6yDiw5BoW++WMhqLE5lAv
FXxvmO6m0c6qy/2lpOmEKEQaZiupVsioPzqqYXLcAkZGS1LDQ4VXqP/oJ9hu
xAzUC9YCv0PkV0vYYsiEP1dtFURljWJYjjrLZzpFM4pfejS9RnSHQatjSBrw
cpkfRKtL5ImD5TPfd+kvNeb29eDP+1zV6UxL37wPc9natH2sXwCtNjhmGNsb
46GG157R3U+Q++0gWInAocuRbA5461HHJOxGZBtuJ1Ufce4WTFltt5oPYd7C
eY5cYxl38rNDdDaaZq2B0Et83wyYHvCiIvpSWlavDf+SkKtsI/YEA99J5NkT
0R49XiGFsp58vp/ZmAYzcb5I4uveLHPFxm+qrYe0xzXN1gnfkOD6UwgcsKCK
x8rmDtKY9lzrYlO331nNuhKKw8yFyCX3aWa3B9uh9KrM3Aqhkejk0Wsld3wn
9/U8L17O0kceO4T/XtdJmUDCGsGLuu/i6FQIGwPjEF7B2eGo02tBvcP+N5vN
OG/Fy5D8k2WWUkr+6HEwg4K1Xnd9rRrxasoNXIkxr9kr8DWb1XeV+Xf8KAkN
A3yuCk1raHXMV38rfN5G+L/j2K5k1mgGHqvMfXClC6ULoufbv/jT+KqahhPS
WseFeNKBHw1AsKw89RVycsIIccW0LvRiI5Rs6Gdv5HKhoHgdE5Upgb5JN++v
NpG9b050vbgoRvUbOa3TKNM/LebVjRx1PufxanbTKXGOJTc36Ijh8/MptyBC
ju4c4LGfJWCc19JbrwMsg4GuxdmvFIkJyto7RLb7hFmQSt+cP71UU8eftaXq
ovts7cKMpwlPdNVgGEIGs/rDPqm2r0ZwnJR6VtkFoxNQjjF0O3axhOtEMTFy
bBKfRUHeN28ZbpqAc9Wlek7S+IGBiSYhVFQ8z1MrSlZJ69NcjeNaS0tJAf4w
tQRpxo38it1dPOh4g5MXUgW4YZdvY4fRqVcH0JoxQB/mXsOO4d48Hxm7Q4ti
2ylsEQm9vO+djWdPmcVF6HiGJHFA+B03pOC9VXoMnsHRdFFQzwKrks0rMoSS
kIJIhmGxgBXCUZvJzNVR6XQGZROwnDQ7bK98BEuV5sA8oOJGPGJTWgAXLaq/
LQwxH4rPAij3MXelwUwPbeUNgWC0gyVq/0vZFV1AW8LZb0dPbLh/IwtTESj2
mfhkoZ6PEGBwUNLa1fdF8EixnZiT+xT6esYzROvgzcoxNN1oJQ3HeN1cyog+
OqMZtFxkjBY3tCH5uu6Bt7gzhufY8f8w2oEOX2GiB4dIQiCztShOY+rxIIYT
w8pRZHLX2rVONKV/ciHrN4ELLKzr54rglXj4JjATawyEl3ZyAD/EwB++r1MQ
/kC0liI1o+CCMLpLxC5v+8uyTHdpGyQQ/yoEy6IhioesnClMiNmLWhwiMXtI
yF0y1R5b9mSnlzrHyjgGEjQpnRNx/+o4s3pNKPd9qTsN2bFnThMcFdE0IJMo
TfdPhCmH251xxIF0Z2wciMLN2kbVUrQD96C4lAxJ3p+iGvoI5c/hifFCqrJf
Kljo/bRzcwraublgcFwJtOo5pvO26wRZM5q/T1PbAerVBnZ8EFma9k9Z0CFG
XV8LeUiOeUZf+Pny+XPExkAJICZBSKN8hu/QZi8L89tQuRaMnX7pNpsk7dD2
tfmxrifsmz4skfSzyH44Xv23THqIqXhenrfPvdcrDX19ZGHhVjsiccR266sw
JqSxQJ1icoHkhHCFQbi6NN/7fnvgxuqvJz9yp1MUZa03AF1GAoWr/DoRY4Dn
FipTYsS4QcXklv6lDyP/B7e2pnA7vrX9qjlkp3Z3BIterU2aLsRT61rJ8qYH
J13YrJaS3p7ySf+QTmBLCmUsbGtPT8gd74IeVQP/nzSRVzOygUnXsrEuBi9t
+mNRGqHJfXIT7imQ1RL7VUy+aSFy69vATS314YoS0Cl/3fZ1ynoAXbuOfxhI
6xaI19gfGblojV8CRMNZANTOjnDaqmfKvX0sOCshBydcerwFJKqDcu9cEv8R
ENL20IGFWAcyKdmiBijKGtHbOqYgV5LjoWkBjV5e/KLjj88HxTTRuNwhhk9l
bVZlQ6l8e+0P4Xvs49tpX049uAR74KR8mXQJO/e5c1c0naj4PCTkqYs8qtI9
IjgIYnVAqpfKEjCHZR4loA+FCsHG+/CQ4Y/hks3/TGZGamarEnHKtJjPmEKK
kX1J88eaS3LerSQuFwF7Ob3IQg6xyTcEg6BwvH87bxAxtHrKKCZhbrU69lmR
6q7AXOZbNLtWQ1cz7UdgKgMgRhHIq+twlj3gvaiQvaxXlEbilbgoFCr+16u2
lPqYR1wkIPbtdSWResSNQqkGezHJo3Y3b2CqlU6Nvz13r2cWrNTNpY8dlbrJ
V3kK1XV+z2OS18oswVJx+s/oVFGuXPYTPz9QjCHpU8AhHyNQiySMDpu/JZ87
NWHshsPxVqxHhNh49iI5JapxGxKQ9HQyV2DrWBR3p+f7kE5SGogCHaXzXC8v
wK3rOclaIi3/AenmcW+DqJkrZEoJ3zKB0mxIvNV2zZNBYXen2Iq1RXIb2YRB
QQCVteOlsH0SbIgyXkGxtIPhxaubnpN19HJabIs+EjW0QwSRkyb9DyhzKIOm
zTniXJStEnyA9y6qz1mNUxqsXvRu3T3fIuBTQWMMoGbwGmM97Uylethm8cF3
4LCINJI0C4OD0Bs3EUCJamBY6lL2pb8zVh+0SIY1rLfsEV8sT6VJtjCVogF1
ydeHhc7yzmGzhwqef13iSjUR9Qana64iexIH/HFOmEs1Qt41YHkBjdW22gWu
gythSZXiCiVdBtCW+Rq1AXgOSIxSlw1MdzVk0CPn5tPOAHwjFnzgMTwoZuSe
Cwo3Inh+62U5XWv1HLYBOW6hJpq7CmdXqfUkCZKUMqqAVdVvkMEhsJdZwnUz
CDf4dF1gtGSooWSs+Qd6CF/KxfLNG0ovE7oXjxnBdbZHPhKI1iQWHR38/LOS
PhXazPwkKm/D4feaFjKK2buKPjbLJrA/uFzFheZe3qSTDCQfUfePElDOw410
lv7AxPeCxq/tdkzDB5IztZ1QsYXDmCPXnSG0fGwDPMnAc3+d8seH38P3fkgY
oomklHNunjgNSH+0TaZiNNLbYbilqH7Pq1MPap6oDS7117j1eKl1JfcySVxK
i75o1uQj+fuusWRVjsBXVoMs8Nc93ihwoujS45U2JAK8E810Tt2JmwLAPb+O
A2NIELgJqK4lSa+AoTgAqG3S7lagbpA0WEQJej3T14RvCUWT6RZH2R6yvtqW
0cc6Gblxk0Yu95U1bCrlKlqf1UNnbJqG6BjbPwo9+79F2mxQCT1SexELos/2
78wQghlwtYxU/1jtFtA/Nr5OEia24uzWA5opgv1305zenRJEzPhLWVi64JkD
MMZ9ueRtLj/1WIS+tpqjpNdjsDZ5jCjVQ7vMsO5blEBtnmcbP6WQgs4CisXk
1jAkY/vOcE6QZMaJep8FY5DNqbTltimxA64GFRh7QeOrUNa6e7hCx7YO6Rye
AmtUwyzaHPl1rTPVufechQi/ZzkdcodCTs+S0+XhM462io4nnFJFde3RvWVf
+0MbphG2H8hg/Svf/vBAIKZ+YTfV8YTYyY8+AHxwc2H/pg0Kmtfgd9xZjDV0
j9duKNMVVI0UCewtTsbZpjuQ7syxcCplTPEMmHKpYupJto/2fAh3dZWjNQTO
YLLtBOP7rzIUvnOVZoj7M0e7ZSysl3VGDQc6Qil4RcuJ2JndxVV+Uukh6wSQ
NaPRJ13ivNGQ4xCRm+KndEPRqYXnp3WCyFud7kdNnbKQH1NYWuBZgNZDG2CA
BXmzz6Cb4Xgifx4JvDTLCRmmwkxlxJIP3PWEObOa6VruINpvOG6bVNMh0gNv
ldK2P6hRDBxj7gceehOrxA82R9tqK5SpCFa6W31vVax1svv6QLMsY73ojzQd
yEjkfV+AwKVTu2HWd4onDX35R8EZ1wvyXGvHEfZqmX597yjSVsQnzXPLazxo
rD6uLYeLSwsYVNrHhZA9ZbcX8NYBkHC5y3lZkUya6NjKXrXaklc2UwgPXiW7
iCNYFg+tPFGLlFZ1KoCiLf7tXZ1i0kcdtQaVu10+wySqnVk8udx9mwA/qvM8
zxKtVoTX2J59IYvUDVDoRw3hYK/9/jBhu/GTZbyWuaGkTNbntKRdbtFCNjyZ
ddb2RhFlIDUjdr9mf0/L5RSGIgaZsdKj141UiPegUDei9yOVbo001mfKl5z5
Kc8kpkAuE1F2cmV+d99vZLstKUuTalxa1wwpVcsDAEj08xAQyI+q6LbpNwEA
10yfYLIWFS6nqrv+q0hfeg1AIhrFkSOYKGQ6C18n0cPeIHB0JBswCGs0Ku6j
omOjf6QlQ4CClcsX8L5j8uA3T0P5Smus2CGhYxnYZNzEwyBSU+DKbn1aOlD0
3h+TVC4THbZm3WdOFHfXGbvGflDPiGqrVLxR4ncdf9Mfzf6eXaCW5yhy0rYY
Y/WCX1LjZMsA1IF2jDmrnWIQkM9ugbmvGfvJY6GrAQd7yT2s9xOEXTfKXxNo
kuUuntFJ4tZIgo5Rib+KaRu6FOILiu1Y+ZsO/BrLeY/zezxZtYLM6wBiO/jd
yKvEAougIXg8D/o1sauFFci/dm6puPMW8sj3EG6XinQHWdxbUJfamjD3K/R0
SPf67bw9MGr9oUZ61+kQU2Wzl2GE6OaFm6mdB7qYzO0iTzaSrWW+zglDfL0m
LxyQ2plHynaYB4x8QzzLKGxX9cjb/59t3ksxBh2aN0JoGhKazVf9g31AMwuk
OR9sicC1FhzJQqcv+Zocr2J3SqZ6f3eRor8O/qaLfEeiC7nnVICfmQjOJYK4
7AlJWiHAjLOlilVL/ME1sLYqOTNBjlxXEUCDunr0MUc3Y7zVPVpI1nfjW3qN
Oc0JeUtw7mD+PNMaN89hBIIYFd6t7mW+5sYomj0ow6VBiE92JYQvjkkJVf4q
Cw48vkhpAWvKzBwP3zlIlLGE3KHIGkHfb9h3d0nFXFnQKiMMy2QmyG2gJTk8
7fFGmPT1vwgaWzcpEQONXLrQ50VX4s5kuwBYaNWCXgSvc/BJgSvSsnddxw+m
o3OqV/6dtshVAUkF1jym9quBD67/iVNzjd0YyHXfxVx1zoZpvkvFuNr0qNXS
DMcygBwEwsOzkudrbsFko1QAFQoeoNJZWroaeLu/blY+mBDCZsNHC5LAYNw9
3ICpO0fMcjxDzpi0cAe/AaknKExBDcYv3uZyuUCaOouAbYMK7lRX4olYTAIi
RAD+Qtlp/v6B2Cz7uMw4oZMVYbP9myyy7o4Q3lwsdYSpGyTesUujRfibUKlf
3ny1nbA3RwPC50XLNFl1c5X+fGtib8RrptMiresEHG9ZBMjkgF364vtuQwsU
x+HU2Ne+RYKYB2JRMawrBld7igHKGRrBieeGYuuoNG3I9SSxc2vFFEysUi90
kfaU2t+v5Si8KpbDYt2DG2SBA2tKEzZo/epwBV/lX5IlIb70vw5LUUGSYbJp
9ly2z0YyrbnhD5fWAmt23qiwVkwLrm3dyRpXuNy6ihNbeXjQUKEI99q8Kn/f
86jMSZHEIRYqyuqUZk+fTGAzQ/WKkVjowpF8E2Kod0qVOKyDHsjwE/M9AwNK
EK7AbNpXPXo112ghL3/p5TQjm4RpsZkF9jQb1gJNLXJE9j0Q/Q1MjYVEb9d0
MpmaVrEpBPvXgjSJz/ILTNvpXv8lyxDCZWqBZvUHN1g5BoMpNNi74DZ7/tfp
8n6q/IOm6SVufEjUn8492pJBzwIAsmDZdiSy/KpdzdYDem1BXuzISlzd/jFd
IGc41rvt425DLMvkRdM71KYxI3qgx1ElfL0vAv1leX3+Mytbcq8pXc7l8y5r
Gb2azrfMEMqwH+tS6cTeBzPG5QOErId4/gaxzFZv5y+/LM23fh7fW7kKRepA
Xdm8adav2QKvyepr2ajnkxtKkQVhpITFTbCoRYeyBeSepm0c0V7bBUS0pYhr
FKM/GAEUEOS5e8ZAX2shIXK5ecmp2lmT4TMioYvm52h1VtOcotbGe7GsBYQw
IX8aDoM1rx9uMsQ5E4aLHpIpsFbrjRk9/cPaLbrKuS3ARMRJIm4QJFyrVu+m
VrthnPlF/RvFsLcOD9x8hU9gTj0WJ7fEkuvgJHYCEDiic8guaiPKSTOsVVnT
u1MraP+Jzr8lZyB365zgvg7CT12bqcIDqAyi9giEaIGX3gQ2gDW+4lFA6t8x
B5bozYDdcKHbdAIDIVUc8KzFvKYaV432YOiJ6A/V+aBDNFMlLKxFtrcmGmYZ
piDgTgTxp56Bma4e3rJbYOCNP/SWIwVYKz3uOi/hYSJTal/MMtLcKFvGwCOp
vQ0J6M4C7ZsZs9otGzEExKH1STdwIlmHyCsf2fm/eLUudRZl9e/0x6bkTIgz
6WGHJeolBG/Lpgc2c8cxXRF09Of2dKMJvJyK1aTG6ixLaIIPd3TmanHoWmIv
o588dQ0oU7gtAnIHLzggIvq8XeWYZXeYL/vG0xkToINxzAhJ2DPUl1x7SXnx
UGrgsYw/bhEjTZEOTW2vlo0HrlgyK1c9pmv236zMbBYYlfbN5hYANdsYUvJN
4Dwhv9qggOEK3jGVvgI0cFvBiCup48ulP8iob6+zjSJwgyfg3krdWtQGpij0
JyeAhh4Sn6du/sld2DWpNsmLR5DhmNiIG233tKlEVa71NtAbYtYkNq4/6fKO
p915JAH+w/jmEGVk2x8cY7qHdBl48fesBuvCg7vGPHgCKs8ukiimFhqwnp4L
li7e1BnHASd8vjA6P0C6qxBVd/8nUy9I+XDqvCg0QJASM2IcDxULBL+d8BwH
tLBW5LUmBwTo3hq7D7elHrhGPNFzX8N4qeb+EwNWFOExOR3+WfEPnqgLKZ2J
0FsnrverMUJ9rQk9wzWQDFvb3i29g19yknxkLlHlTsy3blTjeMa94f4jA9jk
XhewTTEGeUwbfHRT3P48t108OTyiF8G8LuD4T/4uIFkKcqaIDCniXrlejiTE
HCvgwVXK51aSRpw27+8AIkidMFT0NxmN0XietIPK3PvCRxtBLYZ9yZp2xuH1
uSs8z3ucvhkPiJXrGFXjC+fuP4fOUVIF3nN2phdgAKGU68qGKBuu2vIZh31m
KWQ5A/gBGhIQ9ToH7iRVHPPHuPBrobTH7e65NJAR1FQ9x5mFdyTbolbdtomn
CB9keDZhRxZbHrYWeaYfVYRkrx5GeFDB2SAUNA3yF6Pa/QfAJfGRz77ngR8a
PoXB4UTXifZArzG3hZ9nQVog5GVK6J7/ERpQS00CXfBzplHxmb35HNLMBrJl
+CqWZTmOTvHgw2AAbL0xvwLJ9nR1waLDiXLcEbdI+oGXZqU/jiVSBqbEseFR
NrMrHcr7QK6WiY6PpyVprEi3C0fP6jtazZgy11VgsYwSvhZoBLH+sEFhhqN2
F9hCFKSgVcG0S6F24MfwfYTOgyd5YqrzPJZs/ihX8V6VEAIuz9WHNsfHhkSg
4mkjeFKmYamKmKUIa1JBtWHkfj990pjXI5PsuG7Aqy8/rCl7+3emOqivNDgp
cGN2PTrpibVhvbBtYPTX033zBTdjJxWKvxPBbGKANZtVbjG3Y+Ebj/YADGo1
6xKtxOVlBFreicoG3bfJJd2l3VopSNP0AXUY+64ZC4fb9M8RWv7V8llayWk4
ZbTyk9Ttzh6BKMM0+CRfLIk3C33TqoOmCMWodg6ZwDl7Pylwq1xX5fbsnZbr
2bWsqhBeup8Cpc/GzTZ3/XXSA/46K1FC98C4cdsPf7KSmpRPZgjSo1JOgQhB
qNIDfJisiTwgWEncZAr16i1NUOVdROodJocZ/wp8G3ArAJPOp9hTRRvWxri/
3nozy7yPX04yOajZ8pL5+W+pNSWVWsNrG2l2PTaIogncXGZ9Q2H4V/oEySDy
7B4JuZKWMutvek4G7qMnhalnp3CYysSbzcl2oZBU1obRrxNFTDIA4kb3P/2I
iW1yQ/82nLid+IJaybGqSO82p8Vj7YRwnJRCFqGIViUrt+kuOUbAMUwYSgL8
5SMg2TImNh8379tNa2qRBtqE2JL4Mu2EXwKkG80Yqrj2751LSAJ0oZqHkXgn
2gVTnThNP4juoYrFrlW4ps8BJnx5oPpmI+EcozzncmZ+HRtTgVnLJMSBDgAl
D5OZUbf+Q9OIAg+41gG3jsR8AXrA2m7PB6S/eYPgSk9DyyYgu4WnpPVl+gnN
PXpF2jp3hJyByEfPARIYh/hzpJYdtIXD6mzHYLCus/7Kvoqvf6YSRsedWBKH
kdQF5/uLtg3n0LHu6KZxp7QrABOVt8DAExaYO015eoLUFq4HIOc8SQOgK+Ft
UWtXclvwphxnYJ87zC1T84Md94HnHtNEPO0vAyNLoG7b9Bu09hfcdziRAky2
SY5wMyhvpoV+rHXr3a5SgMdYcvYV76/x4X2qKGpTGP0SpVbDywMM2OKSYCLZ
gIDI4gCUB9LFT/23cugggr4LdCC/k90EPvBM8WB0znZoy7lJcMPI8M+/qG1y
QzGC2DHSwGqr+bsMll6qPt4/D9m9Gp1KlfpsxoP2P6AY+Ns2oKqhnVRF01e8
12+Xd7Ic6zNGPISxm4g3J/RfDMHJG7q/qP9E+TyBElZsWiJst8dnKK0yk7QZ
i8MJw4rk+Ar72lwSdnp8vLWDWu97WQUx/PYi1bvy2cwbMPV5LLbdXoZ6PPON
fTHpE6qNpca7s/12K+aXD8pmoljr5zbQWFPz0nxpdT+fIQ6n+5ECRh6bRqLw
gBW6TepxavyZV1EeyL9CY2ScZ8MQJy2M45+IgD3UfQ8u3HDS+srQg/vZJNBQ
e/KGhk//SZQHTTLUs6SetWzENOOYFyE6uGF3MBbLC4i9bq9G4i3/+vu4iwtf
OpMfG1ha+123t/9m5ySFVoDgicRfBMfuqtX0prk2HU4m2kU0DPW55nvx9jXA
zdWH9CtrnYMW/qgFEyT+tmqUknl9Gzt1NJiOxaGro6mvqQDhSuBEQvG44FT7
np+jILJkkDkZaNJU3CZrSAZM6T+UBKRhoGnLdIdFy42RhMNX8TXKarcBI9yk
4mD8Dl47yIRPWyNowfxyPlWw9v8dRlYUTIpEJnw91RlYMj2SXA/4w5wWjevJ
ayOwH2PBibHYXthDbjYXxo5abQn3Qi47NKqWRZaHLCDIXJsDkj62EEnQjxgr
7xhPw0478MQtLcTrwcAKbxrH1T4SBkkYvA5uDEukxqEO7euAxQE5sKRqUARy
KjPFZNl9vdRzqzFW70npVUMMIn1axMXthWbobbLvXtUZwX4bdCwWt1NmJj5K
+iHTdFBSeGI6cY4ngsYAoPQUHvAtMYz173F1QAj5W86f6IqTm7DiQhH8LNGd
5fGWG6XiBvPGFvgLY7Ylxs+m/kySPQArtPLA1xXXQ2JdYyg7ilgf/GqJVNLv
djIgKvU5tujP/foHZ9DiRglBrgj9PV+dftI7a6tfMlphAvkXFCG0cuOjTkSA
GtyW9feiTeakLw6wvSagadc7tnxABsfT+otPnfGryMknvfh9rbRj4Qlj6uG6
q4bvZKAxuDmy4MMyDbKdYROCFSao80DoaY7hrOm7cx4Tyffl9nlYtt3KCNkS
++lNd08CiFJ7UVpo7PThoEabaw459Wc8MJr/f5ykt4PocjzEI8kKyJ41jfLM
6uz80QmlV5mE6/GMaXPxjqTrCisnueApY78NOX/ZshfA5K5VaFLdAyVTrk9e
vRCzVJ+Y9Onpr//61tCrCOOk21f0+TuLaA8NNVGIJesJA0ZSMZLoDHEw7tBv
OZ6ZSDDVXM1dpt5KkhfCiG8EnLF97v8GqK83NNDdTWx4RTCGrOZ7TR5vrFoD
EBwEFuHUUr3oAOZi2bxso+WjEWZoK81daZHL3Mq8QBFdIMhjNRcdrpyrYAIK
KAnoxWrOJQa+Q1pYvkl4iYaWomIQidKIOdgLlINumvzzYsaF5NjGLikN4QLB
HQ7dDALyqmKajq9vCD/ug3Uila22fEzejF5y31v2EEKkXYee/y+dRkHZXZdn
diO/c9bG11jbEUEZufLyxkcEKUQku0F+m1t5Lwi+n21vj9LF3FmEPrgYfyci
hi3YIwuxFUQ4JipTcOgC3ZBzVMv5N+47EIX906nBjRVJWU+agzSSqe/qMQwq
uUIyna9aeamhHvCUnUP4fUt4/uyxvjyv7tyD1R4RAUW/I7DtoubqjIPpCPf0
pkBEtOBD/zId2uApnJrD38HsfvDa16ZjTeynJe6lNzh1NN9amNHqwuW+VdDo
zsKvY+JXl05ohWzQm300p1tJjTVsc+7+ufbPBGxOBSghMdzJ9gvV6QsbV7J7
C981787rt+32jr/yzVcAK0hTAx0Q1T2YGCsu/MBomS612TStKi9S+7jEPg8z
n2n+/NBLE/FCILm3LCKN0nd3cSCxJ1PEmn2ytLK/S8Vh8raM+4d2Otk6I0cP
UGtQSzx+rStkxveYk54Yyn4OgWEKuq6FW6eg5hDeT9uFR5YjrsL5o+LEAgaS
O1S8nmOBcfUUrF/aPL9G2joFOiwfp1Iq1tR92aWbs1tcKr58tule6a/YV0F4
s8aj3m27uhkbhRZEB/CgxQmofGzAhehbByIt0nAggbwppmQFvvt91uDSIlcx
r62BVwuzu0d3BszdCKgiZ585zlDWg7oFfBcHoiBhE4l0edPaKqxNzZoVNcH0
k36l+wplPqXRe0HPaK27TOW1Bwmad6WDkMxuzjug+YANkU4sdF0TyyLFxPKK
iViScRVV1Usuyjs5Y79ppGqjudRjyxnprYmSX+V52ShzZifxaWHnKifQPVmD
eXswKP4TPwb+bFl8vF7DFtNB4OI/mWrhoYq28cv1I9t0ol7wynRPXrM+Bns/
gtaKseIRbwu3zYZgn6jC3cL4mCSJcnNx0L7ma6YJAJz38eNEFeHcUFha6Jy5
ZWHZzBk/DpEdMZFyxiLe8lvjJN8FPA748uTekDKvt2igB7JQArXVZ33SQgMi
TDEuwaoJ+Pk/A7/MnZwDojv+A/nEyvkI7XVNtjVkwZQsn4yECRnkDM8e6zhn
1Wv1yaljJnUEwLgjJUM7Ukax0tFVxiEsc+NV3kIjjKvQh5ym5te3pOwWN4Ku
xg6Rv9d1s7htb+/ws5+Ght7WLjdE4MUK1LHf1UofFuQg6olbagMG2Gce0bpa
S89SQImQ7a0P9xxM5j9ymdcN8MWKkE/YEioYWcsarZhRFSgSAyMulump7GeP
KZLeRiCgi6EfyY506VMNWbjsa9UFyOuUYjmMSJxfJH+9sR6khS5nKyXtYdtQ
JzyOGj4dCggRQ/TfxTFZuykTnbPkbJLATI7jzdSCi/Saxx67fACVHmQ+kvPB
vad82FS3uGZRoklSaKrtfOTWsukW4FWVE+cel5BCKtxC8bhjPRmYBjmb5CiH
PNyL4S1GqwZlJWk3H+sXkQmHGeqiwncCq1kwf+UaW7o0N0z2HehOzVQI9h2r
yRTPuyZ/maRPHe4V6zVEp1gG7r2GAu5YdqKMmQdy7oA+441pN7UrtPOpGGuC
cQ0BgOdd3hGqREeMw14xEX/SRpbTfD+SLs5F/h4tWfAIb5lIsRnzJLhy15eO
i6udi36/fWTTBjWvewIDEiYmf6Uy4i/1ZBC2Ef8dXwecAz3vutxKmczRV0F2
H8zwhaaAEEErBZX3NlcF6W56FF+ox6DMYiVjvNZwdby4AxylleI0HqwPW+wp
DRrycRDdippe8UXbcqfr3E9FjQuHFACtQ2TC7f+9W/F3hEJ0G0PVsd51YR2T
T4U91kMhIB9jcztCBy81Ui4c03yhoMF4hG5xO64rL7FtBf1G2505lrSo7SeX
W3omu0c1MyGLuGjPW16kEAWPc+iiIUq2huxRdvuRz1EcFaimXxwe1yRkcJVR
kNQFEylrabCF7P1WrUgL0O0SMjgCVZr50NzN6LtkHuU6QGnzR6x099/42qbE
G/VaN4nfekiW7jEHW15evsTBrPKO88M2NIl/g7GbAtqlFSnlULpKF2R4/zAd
6YX+b9Pwp2Hw7trfzSWdLUvWWKjM0R55h/6Hjn3qLJzvvYSE2IJb7k0mLdc9
hLVLThiiyOAeWS1s7GFoPhuZz6yYHZGUoduxCBPt897ruDOLudJcr+NOG1KS
Wf4GfkLv5fVA2g8JJ3mZ6QwFNMHKHusZJmEDGq6d874Z1axSrZziYUZ1J2Hg
HJlFzIwZM3i0HjAowpooIcIdDs+Xp6oCFm/OKbEvltXWZIurWbxsKteQhpkY
FY6qcd2x3SjaNLonREa80wQPWIq9imDroBerjUAMHAx3TTRYjLvOEgl/SXXy
uiHI4EXFr4Bl8LpDlq8PQm7EDMEhL+vXthYgr2HflamHVk/2ot1MKASEtzQn
6VNAkYPafjtJUfqo8TaJJCpPr4SAGTl89OfpQpsOq3tieUA8CaUH0DATG+Iw
xb3RBTN9lLabvHKVB1VXox+DZ7Y1an+oMsWLt1iFt2CWLjmf4FYFF4pROOFs
1e5nLi/Vs+Ab1+R4omTC76r87IFOE/Vy+xEzW0nCz10iWBY08JX3+qkd/YyI
sWbyTMQnTZU3hogrn+LxNqVHp7gAmTs7XmpKxJD0AcbZ1KczoquEI4SOjPXK
vQWKcm6ji0HbYQJtkSoCK8DbFfw37GMjGN3BfFf5zeBhFaCgM58C3vH1s1ik
mdXy5DPHwbIAjiyyg74enL8+V1yObK2cWoKBFv8BuLcW64tfpN6x4P/w0g1d
jSr5s3kE8F0ywp8Zt1JhAapq9+ZQ38NKNl9gXVl8P5zjXFMblBOfJwj8Lzi7
gmhMGThuHETVx7a7SXocXjWiu4ZTUez71BknTqIQ/L9v5HFjvyjxo4+nWQ0T
g4W6uZ04/STL1T8rgxvSfSLc9Ly0ejuyuADP90UR+W/UrnKwVHak3TaItpfG
H2yPrwpeZmJ1z5FMZq/hZ8K3/7GAugDskCXrzUkxPddIbEEAs+/ctLjV4WdF
nvMYBkoGy5XAs8m3qJt6+l8La5hTebDA2t5YS3N5M11vH/qUe/AXdZLhs2O4
0CGbyCreA2H/lnNQmqDhO8D3hEG1MOFvcHIPrhAVB90y/3XlVNbIBeapW5kn
wjTBE8asq6JaHTzq4ZA9OdJdY3MCyJjFJSNqSrSWTmj8NMqqY8VCQvPWBYIE
IHdALnOmyrPlFxBGFD26/aCC+q2r8eGNTgseCxVqDRDCho+ebZgglbb788jb
aN8+zOvc28GuCOBIdf34Dn8XafvbT46T+R9uxm52y+6zPTWw2NXNasfm95Tk
9r8kAq0XXB/1zLdWkxGbmoygOnBII3x4c04CnkzlnTgKkgmUic/ybrQvYZwP
V8yLwFqvLcURJxlynMn9AX8GfZBQ/LrQBiqiZ7BG65qjB66SXoOZoEWQCkdN
towBlYkH+XykYAi7UpopvKf5A+ZySumSwaykkHoLezmYnaeedowwd3+hJQDF
yiPEv7Qvuy4PbqNFYDBTILUHgwWoyvK0ac7LfFigLM6LVjxfwNO7Pm+gj5Hw
9CRYFWxcIcA6Vl98GzaV6Q4q4tcaP9N4EbtnH+yS1gwhBLJk+LjZdKcbX3gL
YVH8INgTbdEGToQJVytFw98SnO7l0iif3g++Lf5JNMbaRKba3B2vUNw/03Ko
yf7gDg76AVrc0PaxQTyycKS2JHnYYXBDqlrgB18kGaMMUAssSv1ShcZDUon2
4dxONQ9fwxbpRM5TbMJD7fEBK1ao3d8kG4CQgPWEBH3+so0Cg1iK3YXxzPVr
1dYWXpkbR3HVAqtgJUaSCnSTz4aXjlvtFQ/zCY7H/GnQLb0t6hJ9wP2mYWGW
VUo3hbcebOCcJz3LhceaU93vvjJ19RO+j1U7Thz4Q2w7D96zgMGWhLRIl2Fv
PO4okEoYUwbcSZSxBwIk13e+Mn7cmw+87Xi0AcQkPdqPDIJCsEtBwm3TR1Ar
/Hm9lSK7vuhTyndT45QWouGz9yJkvHGbxNkPQ98kQbnd4QuYTBgAhjaeWPBh
IbW5oFcsPNbVZW0gDJM2tUx9UlNV+WZAp2DN1R2vpFhSiluWKq11Vlfd7zwy
bfz2lBz7snl6mS8xXDjmWgQAj8SGcdEvOHfdObwKqITSen9mLp4GzKTuAt3E
phylAr7oZuJe9XK2imeuedw/cbpU5nCtM0JwyaTdGYscvV7XNkSePD+AP/co
Td/435D9fN5g6TXLS/1uMsIg7fpwFuUtLgFiiFfxeUHEX9c07wlcCy15//UA
b5WvNR1f99UhpVuZE/i6YCZ+nXaUEqcaUUVw99JN7KnIrdpusYNAIADdWsb3
I0gpN6rTCZx3MI3LpdlvTbWQN/Fw0PKkcsouVkkpfpB4uGkBDDETFbgYAJ0o
BJMi9/oF0dXtqEhskapYlQSv1Sw4toRSe7utz2dkInPKQRKqN7c6ruZAXg66
M7QGXhOli0N/DTzZFksEHbdLENhCG2jOcoMOV19tP91VzV+Jpq9v4fMatZF5
nrVXLNtu7urs+tRjOQR2CEgjNIXGDsklCWK/IMxIDnAY9SQ5OvyeVy0vbyHf
L+pxaDgCw/01tUVB0iZZBWq3tk1Hw6waMaT9/7iu+D2G1YCIqng7h4j1BYiy
oqTXaoXKajipCfaf1E1EWHmoN2uPJ7dzFG4C1KMOoUWycn7kCMFLoRc2F5k0
rsCgGRXUrxC8a51HuSX+PviHv9RoWgyCCu+9GVzk73tRj9ZiyUQCRzc4xTTP
+A8aVZVbWLzpyPOHb9CPilU5Ps27n2p3SMPVhoNcPaVShUs+GUkCkoUfz+cq
ZL961h+oetj1l9yESYOhV6zm15nWkVf8kPL3AnkAJjBwZRkRBFHPKykYrtvE
+BzP6whE3dRbgB//HlZP0lbT7OG5579Grl/9uvhSVbFp6eRHWh5+uyIIWR0t
6S9aLJ+ntV+F+4smqLHu2/pcj5qC9c7kCYD7itfznDWuS/W8yyzo73YppZ2M
vTn5jWv68sggv1WQ4+Xx8YnFKgiMbFs1uFf7pdbX/wyiOuu7io+k710APk7d
3Bopaa2eDDaSa66HXqUb0dAt60kiJJlBEsolhPkqYyLymhG5n2sh7NUh4T0e
y/2m+UsnyCZRhe6ZC08qrmCs7asAS1RCrgMhmDDotUiZVQMKKLEzPNZz5oSw
VMXYHa+mm7dds+qgSF1VMpcWjYPPqSVO/SSoN7u2vQhNeD/ZI/PijEoyKiuP
I7uPYARicQzk52WEa2JYp9f5FPOVjPDBsdd+n10+t9kEHZyRr++GxWHN+BgU
ccJC9k8Mq44fic0PAwXNWeqO6DcqOrQEXMcBxriWFtcd/WiVVxbT7DLnBw0U
IJzgl54kq3xpuCDmK2vUxqJ9zr8+3wT8NHiQL5UaJTC3GqD010ngIHAlCHVe
QlrS51/c0Gz5jR4VkhL5elJU74QHRDC8mhourMXqxFpUVHpG4+f0WTXMkeF/
sufnNOV7cDS1wPFyIoWa7TQiSiEjeJNSJ/9M4JcQD0mgrXXKQ33R5soWaYsb
j0HEn+scqMNMvMGEnuFqVas5MqBYtmCOmM7cyruxV0WNhp7JzWsscilOVhC8
moM5oJRXu0TKZzuyGfXWs/RGIBxLb83N+F3nJNFAQGmRZ0kF2YJkeB1roeuS
XVH11Q5XLVljMjQ7Eg4rrSjoHuiRqc4FFdqkVJ5r7dlwb250Pru9APAm4Mze
7hpTiRcKwS0jH7m0Rj7iTsTAg+nHVQav1Pe+JYrdflRen0XRl2MsYXbA6V4/
5zOvz6eZz1/X2pH8FWqVVKEu70QDPTwDjbWg+qBpxKhyDWM1hQzKf89RaAnh
VNeoC09QfRDnGtVXD1RFF4Icw0lotalR3g+PF1D9wHG/7lPgf//L1KphfRmd
k4Wj0kzVnpAYZ6OthYk99I9ki4OcRcuxZQt2BHghaw+zn1Qz4fGP0abNTtVY
ABhqtJHjqY6Wox8+PeeJWvqB+iPxTWkYa1mVs5/HpqFEd1yPqXwgLNzwYIzY
WUgaopyFbwReXICogmYR1SflgqC2IJrkBNRSpnst6r0RAmcG3zY7ZDTe9LJV
BY9AWDhjxU090wcl/IouKItG2x5ZHdT4kCnj0BoBu/AUo/QercEIF35lmk4M
d3zrITmbQIt/2g0MpmyqcEHuy3xYaBBL9Cq7EJ2oQ824w9zHh5k/bOhr7eF2
sDkPA2lgs4d61L9viZUJy4emglOZoAGBW/3KN3f4OB7dn2C794tALMMnOZjd
hZ4YBSI3LJ+HyrPcAhdKlSBjmCWrq9znajOi94FzNNLsbstVEN0elgelbFbI
8+sR1MyZqjJHmZWp5HNaIcDrV36+1XiXreNwo1z2GX/Npv71hJGzUk2+H8nu
tzX0V6aWOiS/tt9G0+4UoiRypgjf6JFSqore6Aity53YV05AZ11Tbbw/xVl4
WFZbKIhNZeM9BQ+tTT84Mz94E/1UcHlRoFC8HkuETodq4d8oFIvs+aSNS3t6
GX9SyLTv9o3TMDQ54SqEfG9zqdjrwdXk4QsdAcZ4URHNutVIKmEDElBt1NS5
4B8HDWTPATw92kR+/iaTEvscI9aLt8sDawQWIgsBu1BfN05M7em8yePP4cE/
24YCEvNAYXkQV5B6vsMS8v//B42GzYfaTkjca5Brars0HmqoDnExKSV2SivK
BLUtR6qFUigJCDhuUGpro4r79nSSkoSGfUgpSGDkHjwhOBqvdHbXHsw6oxg0
GHQ9LSaQPpyPAEw0iAIUP5xTrFT/gy2nmYIr+toMicCYuh91DT1qUEgSAKbx
7rQUH7FdyLmLi20eDB1Lx1Oz3UFfD8fETiY7YLkErKw3QTe/P+yixvh3Qajf
8loU4CjradQ9RhrQ9W7i7zlFw63JL0H1B9i6na/nsGyucvj5y93bQ2R7VMXw
MuQ1KvwHYNkrIt97C89+SUG8hyVX+cgctDx72cDvaIH2BYHsaaJyKeFriEBG
1dZzx3Fyv646mqJSioW0sh8Nzn8N+WT4G0H6WwEdsxscgxD6tiaVSumSdu3q
aQtNpok7zydG48PPa1tNpL69S39/Gxn/o1h3Xcq81RZJwBEMhaIEhTK3m7WJ
4HFyTLjXjTbNOXDbOib+FEN2aEM31oO4atSlURUNVYdxC10Tj/BIqrIb/cdb
ALUCW0r58SMb12tHyI/lo4v9XQHymij4c/DYITK8BndJ0GHktxPbSIf/sP/6
wx9kPffhZlq7Ic/JhHDyl0HCCPZakogX1Yj09fTvkUHaC+ElR+6+y//zt4Ea
quTHuURDieI6K711+Kk/3wUYhC78mfVLSW1eL+jTSNtjvRG2AF8YNBKRgMbA
8pwmw1Gj8nsRBsKeAP268BIJZ/GU7YmE42wlaNkwEgc3rAURr2M4zX97mJjB
lVtZtjnLBkqcE5+PxYPVXFzTfi0tmiRry2zsHuj55+YWYAhuYQ8J3Iq1xCYa
DrSN+ixZQqfXpXa5q1W8mCdXrvkaAJ03z5Whr7Xx4lM/8UBOry4OALmrWlge
p6N9XS9G3N5t5shst4DgJDd90Ri7fjlJcaY51mE1dXdnIN3yl7ORPAE9U+xq
oH6Lc5PLSZUz50cReVToe6zNmkOMAg3YCB4k5sDzjiaRcyCx4q/f20vKGlus
6kZlVxmMihDdtzHIbfXMyFo8TWHw5LfZ+KHTFl7AllQVwJG87B0rJsVS1MCR
aPbg4t4m4BieRuoRWX127wopEZogjApokQ5E3rwkNaCqV7KC+skM2W8LaJlD
kr+PXZdul05TsFq2LjrsC0NHgK/2sEayT56CBiQRoHvizHLOLT8HbFUrykDZ
UNrJuhbDQHnIZpKqhW+4Gv3+czbjAejTUenI5X9RCvZmwTn5tCBiW8opcYVE
1l6IKK8ptWB/f+qZ+8++Z1ODcw1Zopl38zCWcSTWOsaa+/rK0w7rlToUHijA
vb5HYVr9yu8IeK/lrgLQmzkLJ1osL5A87SbQ25uFac4Rihy/sMa1w7ez05AB
B8R6nwM73adXJQuwZbfnwzyj9dJZ5+Lw4KOrWq6F7W+LjA3DzhpkKsyQOSil
SGCkRhJxTkKGNDmh+qDE9LKq2st8C1F7tCzgkqC6GYLzA/LQ4w7O9IAGIee2
UskcDEWqyDFUpYCqhxqugoje93bBsv1OagqGYHFa31sRD+62vvMr0X90dA+6
MAHvo0MKQN4F8nKhNtOkn1Z+Qn6FClRrEHp66kUIqC3krH0h4XvJZ0tx29Mt
DRyY2DXL+/Xr3gTCPVdBjsnW+7+dCElDxNtTUJGrxRiSQD/tn7N3mKogmyTI
bREgp+vBFp4P6d6FAxFkEH13ryicQKoXyikGZ2b34hynJHw+H5/DqLSOzcKY
IiRPxNCUHrUz3sJRk2qe3qmp+JwFzw1XOzXiprWOPxIk19C+F16MyyMmRfhh
Aqf84JycLK6q1B9Rhx0f/2RWtqnYO7Tt+W8dsh6nL8FZFzFsDC9ArIDJ6TZ8
7+f6iMh7f6hQPa03WK+stimg8ANurFaVKZUfkvJ61aI+uS7I1/t1PdjtcDLr
JOnVoQ+7AWOMnaqYIlczDnb3Pb87VzNrDzcUVEGejEzzEJyr6kkvmnq3VNwE
fLLWzGNki6/kZEB5lFmVSZQ2vCdzdFYwuRSbQJi/v6uIsWTwF46+VTb6nfPj
L+99sVm3zTO5+liufQ5MZt3iuCuw/I6E30OuVmzoLL4iSfm2P31zD/LSSNKI
GkiN771nl3Su9IkkmtOogpG1pDkvPx5dTktuJUh3y/vF0MjrUtzmwUYT9Hpc
SLYRmmBcdSdujEzaRQW/4NqW3JbO7F7H0MC2rDa3VvhmxPTGgxp0agQEHWlh
MeodSxvj3tcPrRszfDD0BuJ3aQuvcRVlPGXLkSJoXol90eqFbi4EgkiPYfJj
HAkJOVNCWB4btwBhjKQw9nhpha4ADCbl/qA7mkMR7WM8m9LSbJT3s9h1tVCG
auBlVG+Su8YUHSEVKZCs3/+cY8qcafleH7uhvr28mGj0BqTUmG9SfmsoZL98
Rd23EgCu95D1knkQzeLzKQriJT4sUA2YWHGntjdeP0LoQnF5HNH/kycDVBT3
cp88ZbTVIdC1uZoTEE7RjJ8xvwHPlSZ3bu0kXzu0xgFGMbKSRBt04HSMIqW8
loeUTYGto1a1wnQAvORsES0XZi7PRRWTMM8zABF1dfvSrpOJ7jaTO6vUPB10
Xv1+5Ay3cpOV64jlYy2Dwlr4EVEX4Tq4Xj9szjAnXohu+fJteMqjcwCxAbqq
W9dzmCPA8u051jw+czZ+jGAr4KoTkc50iUnglZh/iEA1New8eb15CzP3TwXl
fuCYrYb4dYWp+YhcI8gyRZy0ZfVPEUe6MaAuuH8hmcCIr9NmJUpWGihaapMs
ILm+gux16xPEoRwLx6avtM+Xkwa/gZlKi8XGNeJ2FEDig8obWnvxEqXzyk/N
232qUo6eJY+lsFwHuKba/LqVvjVggduvN6mUe0XMESoToYOPy/Vu1tZ9Miuf
whhJqkpD1Uz/lWK5RHpdkI3aHKLOUSdC/jjOq09f07wtJB0Ge49z4491Tr9z
iKpT1BqG8iCts51z4P54dLO6pAJ3XFpYFLJuHDFfDuUaPgcxgRjZ3y/0P+lU
QjY332DUZxxjoke21ymjUl1RTAQZZp6EzyohWRD9pIzIABOyMuKcRdwYM3j4
IuEc1qg7jUrnN3kYTat60svSWfLBQaZKb7czk6Vx+tmI0dC3BKxLpQN0bAxC
ORaAND2SKzZO27II00B3yPxORfnMgVxw/aV6cn80BhzIRNS9paiKAhtgMPvl
tJdz0LgztiDZ5BcNpsXrZRaXOFk5sNgRBjh28EDa9tk0hijSbC4HfQeGATvJ
UGrp1+fAUCFy9rIA8ISP7Oy0iT0kPRCUSDErkQz1XukMxGze6WIPKCo83oJV
i7VS+QdPnbk5yE6y8AT/Yo9aJNMHh7i5ReMrCqYiIWw+MdD+OAaOCJpeCewH
Rw6vk9w94RtAplHbzVO0hFRMAVP7f9/n6kR1eRM801RY5lFOgJvUhsxCILcC
/6ARsxX6Nbiu7tr+hsDTL+Fse5qQ2HAfgI3Q4dkwF426EhKZFeMKcsXtyl5g
+VIm2SUyjZcDUA+PjcLf6U8VHQBRTRGPoPXVAXM2nhTKJGMoDHAWicNGiIkx
lI+K6a4CZr6qD4uEq35VP4CFM4WMAkQ6nsrzjUHS37lIvY3+Or0C+5HqeoJ1
xhUuCHj1Onru6WMP5Bt5lwpYisrQ/zYPpn7v0KfBbgyr0nP5JGkqix0Tcw8/
m1jGyQOXi4pXfx7tWgYSHjmte0GBdDFSk+KSILGUT44TIvGrXjGxNspFBQo1
DrBGHGNPLl0l0Dq81TQTI9ds7zpIiuM/Y4qrSeeOnbrcUFQzRSno0ugIGahD
G7xwc5gUU4o0yvtUf/DkuWWgqQkkZrMofMs9ZtRXLzXkdFL8Emdg00jXvNDs
mZBxiwbW09i1MhB+/tLkloUMLSPVRt9o+T+HMnVfq8jS7jrUl1Z887exh2xk
ymL/ubPHtvv7GuK5b5uFrUs/aGtYQcjf7DiFqzAGDtL9Am7RXPzgy1pnXSpQ
1OhX+vSsujOI8R9xtR+Yfc8tYQqW+/1wu/hS/km/vUfDatMvdk7p2eMA5b3j
w+ZE7hpAH44coExTIfGjTf+afZtDqAzEYfHBXEj3WbueLIun96sMXJFrL/br
82VKN2vg00lBLaaJiVAG7trzbwVXeO1yB3OoMGv2/Ey2cezvd5UwyvQuV3Y2
VXhkZ6dNSF4iTnpmL2YiyE6+l5jnPuKHPrQkoUQ3+l5/PtVn7wVdbCsCMgdL
FFvyytY7lqot+kiPibewUHLE4wpXwhRRkYWsqd10Wecro2Cc0gC3Yx1IhKoZ
/Xq9NfIS9nCFeP6sq5nM7/KOQ1U2jUIQnZLYY1oZQbmCZtsJr5okmJbJCBKn
b0Idr2B8v5kA+PS6EVzdu5MWYctsj8S5Jj+Dm+++8BvTAvlXR8ku55xnw5Z3
Trxcw+ES8ykksA4KLCO3TBexWVDq2M9tIBmggb8u/DEUs+MNcQEUo5mkfr83
ay2yZuN6qUIrk+Dn1n5wSsffd1WtiZFZbDzL7S/TT/iS8Mz9joQRhM6Us4aI
BtRks5CQu0zUvektWsM2XR2IgOxAocadteCnQolwfhV2YNAaUzc74V/dzMAP
TmKD+DxIRmVxc41hqKK0baC6Jhqq5KSIeHMwpzLRkzrPWoH/ZDIaNWuDaTEy
DyLV5fQUa1XZ2AMqCmhTZmaDL6lbICPrC44XK3PGqCFzJTtiCddhqi7HAlS+
vk1T4k7v5Gkkcs2XrR+0m75ft2wle0YHdJYlnzZBbSOEY5Ml9j6qJWUGfgUe
ZGEnjRDwgeqUMJr8PI7lX93hmsHXXnTkFXRYMvU4Fvm4NbNi0TnCJA4FDbnc
inh1AMfEApDq2V1n0kKVWrGkQF3i8Ohv90N1On/jcwP5tGuItlGYfx3c5b8z
vdGCLcWnmFYmte+NQwxtSF3trP4BEWwB4md22iC7GBPb8wFcz85jY7onOIo3
S6XOV/tF4W3K7TlPZrLTJCxRE6PJXuRyTihB4n5EVRWk9h4H5a+qnFb3ZeqQ
TZ5tSmzkZzdNEuZHowC/5YZp7CvjL9xzWJemWQhK1RYHV06igokKN5cKofeH
KGuQJQ3iuAwyKVTmc1HC2TrW70ULAh9VxE3SnYuOMh6uol5tQqtb8MhKlr1k
5OkRfYavjRqlLp2BqodehgYoPOmRz2/SsW/mt3VUY5fPfeY5MzhSt11KUNXt
VdFv1CVnCjenn6R/+t2JYD4aVlC3qTVvrhLFixYFyc4lb4mbnX15ClKH25nU
xHA7hZyHBpnSfDA9/wrVMIWm3LSi3aBcIpzBgf4xqeAXL8wDo4wB8bnJNuRR
8UMLe4J1GDOLjAW2BYxvVWfGozTVevIDuRVx7qiApYwd5+4eKHK3jSxA+Syr
PzLefwiWMB+Gs0AXemVVXov/GXQd/mWXsFwPTJ8Y9/JVUcQTeoVA1M4TeoUb
IK34REt7ny0WvKDSiv8Z02BCM2o4NpK0kTvkRS1Gs0hIWItdhRb8HaKQLQuL
baSM3LdAF3lfi+FtUVCm4VXLbJqzjWuyFU5ixcpBn4bizNNDaIvalFf/arDD
YBgiApROOChTvs/LhQOqkfx23Ch83+WENe1nAV+UAlhO/vIfuOwj0LBHCCPz
zHTn0lh3DYgq7oPJAw8JsnE9DYbHZSaoY3ml3zP/iwT6PHX5VyvEUAOxVZhE
Zfl+RnPAy8eyTUahPIWoU8/NWyWLd1H5KHe8yBnHVK/HBtt7ZKv/DHiPVuPR
jPoDdcOfxukC6p4xgs0DGNu5SBtCse3QOC3eNjh8gLMVlq7LE0SZlxWVx60I
PF+XZyAwyRURt9hdxyTDfTsOtB7q3bXyOGH3bdvDEQm6OrQ4ze3BuP+kr3mL
XlEVfkDojob6WXzMo/Xqgn/0hHJ5rwx4hADsF610x4wz8Y1O+XSLj+9En/7B
dMLLdRJJ9e3OY9YWYlDSA1A7gD9rD8EeQ7VeLnusLpiDrsxOaS1QETjEkU70
41rzps/MCAXR5IhMo+tYY1VTHOFV17DOe8iNVHT4sT2aqY1RlGhnMvarpGy9
43ySGyLzvmJPS/GSskbyztM0T4FbjmimQer7lkENryry4QbGowgD6WoSyG30
9Mxy+PJ5ycnXIRHI4XoeFLobUPt9YmnY3LOmNoQ/j39hTuWUZHVQqQt8/lO9
CwQwWsQKqQqAKvQD78V7rNPtr4reD2uec1GeWryrvPCFnKTno+hCHTTpWoqg
aGJ5m5ySDZaa7FEKp80d11dpDF2ZZ/gO52qFWOAYgBtc9QP1mOn1zvdW02wx
f50rRTmv0281p416ExeL9IiOM/eh0tp41enDsrWWQY22T87cr6xjrtGaIk19
dmY728yPmrJ61FxLjtkmwuOJcvZlVCzklGC4gX7rttFgmEWFDtMjeMh6QtyQ
KENFIO0DTYFTdiyh92V2t/3V6Fhv/yuPWwg4NX7F+giA7j92iUxGzG2PiDCI
qze2R3DPCAfXo5tlL6HNGT9OhjN6Qj2sZlSUL8zArIvm7tlpXBSE/R/4fSwA
pPMahalEy49sCp1M1jilFsCYMmtWuuV7bRqjNgZfzmY309UPy7yDdMpKkhUq
nPVt21YyiBJG0/GFBxjlXm5dS94E5GfDqHy/pOcf/D+1miC3XK97LlZ0Ybng
7S+j3wF9IAKMiGE7xU7k2wu/3R0rSwdnwgaqNT0n0u4hFjSiPPMPv/VUpbza
ByEytIE5cnm0nDI1k7QDDysy6oMHNAiyxC9JeHqax86NcZXuq3gL1UR1NfDG
yHLzDAaQnmrbBE40dgpLDG37t0hCotntPXMPxUoFRxliNZ9LyxY0aE0JOSJW
fz0aIt0JYg0mrpV2A1/w3AB0w50viZ/SYQFsbZe7iRacdml/7K5CDeejrcnC
9/kq/e4VvwpAq4IMmM2UAp5uYfAHRwiEuKnfSa0MCTeY918jGh+45BI6MKA8
cV5tloBaumV8vQZdYl39fGg4E9q843n9GtQhhR+CH8Q7filcfgiAtc9sYgHK
YpaxYt9yPwMJwjXiioyTD0jHrCyvwX0ug1L2WYLLOr4vkBMpevg/N4cZ20+z
4ed7tIvj2Ok9HF+R2RRPznpd8UPKPn5Tobarrqr53owsPbODof9UVsBlDL4L
uZjwJtA8uGLVXqMgHoL165Vnhd/h68iDfXmsIA1IzoKSINvMTAADgw/F6rCc
s5SGP7gntpTqpOf+RmpGEknYgD8IaOfYcwuYCQWUNiza7bDVVnoR5LwP7kDp
LsSoDvXuJlxGaniltuiSx3Y0/M1oU0+/c8IiUpS3lhmYt8apCwhnhXZZs7i/
j64jVOMZGXXjekrslDNOEb5K0IDuhHaM5BKeo7d359FlndACtnOXHc4ZyZMc
A2J+6ByUUGqCrqcSwKjIqTscaZAieTFAeZySOKpmTuTS2fsC/0CSbJdRSsz8
rAlrM27rhGGggYMreOuuwXTemmgeXiK8KC6/aThkxS1vEv9SEBCdWfCk/2h2
7mZDef7MaDUyirBlMSCODkmCiUudbhL2haQ41UfBF8AmeqLSMtJwbsacA6y7
t1K68TyWEE0vbeyfRbVJUS+fr4e41U3k39OqFkcTbfEvik2VOSzknAOJS8h9
a0RtUm7glMPeLp++VrAt1qzPWOt/gY/WD9vJfzCi3AqOikqLXT1k1aEi/cJ4
VPllH7OyLQ9b796uzsMCIMpmwoQNnKddp2dgY73yJ6r84p16He8P8pSOPjhB
lyXMfgtFvMJiEooZJc+Y6DFsSL0JW1e91CjjxHVs55sVOuguGDx38wmg+Rdr
V7umprDmOZYxHy6FbEX7TZCbLfFEw7vM1wpM38KgpWgWvY2SCAReke9d9Vi6
WiOpTY4hOCJj0idPg4Aggs/p6kD5zAJlmruD2qkowX2UqzXp6mdagWCiwPw0
SWb6gbthL1F3mjdHGc2Hd41ugpUeeZj6zDtqvNNnOynHpYrsh2e+w0jab/8r
iZ8rbZS2Y7Ucpdpec2I5KUUesrvDc5InVpqKLkyz/qRJ7G1HoPBW/9H6zKzT
V8xLHf2v/zTstvyYM69V/SJdVD58mB9g63F8AS22LIyd1RV2umUmiaG8Jnyv
yOcQuQyVn+/y1SaIGlpTgg3D03dRSzRH9bPYzxZZOtrYNqhfmxDEUOh0X9iJ
9qLKmNNQ0dzk+6WyrsxO9UBFiQ4eHKPE/53Tkvxh6VESfVtDc50LEERlk0cH
EMfAnUemMxj/jpnvGlJ8MdTgbXppstw8e0+bHbSs8luISwfSDdfpOB4Z7fh2
UEMqNccH1JUUpKIdPpBp/so9KcM1pZbzRQR0X0mE7lfsYVcuMHl1PYVFLoeQ
9kdfeAcMjaQNYw1Ozw+cN09T+1XCIqAXNRQgBELI/g82B8t0v1nS8qO0dzzv
Hr2/l4oxF7dwsCJAcQpBZeVqzH/5SjbxQ71kxFkxSFDJVH+Rtj6aPKx5vKYg
smyuPZ+9t3otH3TZNQG3wXiPzTu/lDneHJ66iLiNO+xfplCUCO39e5YlzfCb
2ZiVcPcdkYLdD0MSYK+RABHjmptokO50507DRs3AhS5eyMG5dZ5Y8eHLQyhs
qPH5R5cqge3ZSweI0NXMcOkCVYpyc35QL3seyUF2H+s/rjubj6QUJIL9DgyH
rkhWLBqq5YjAF+WIBpr7ENWxVgCVJtKCx+KJAmnz6I663fQVGPObekLfQU0T
m2cq1RepIOS5FQZGKyLEQlIN70dWBnIxxI0BAXI9doMaTGOnfxZFyAqLRrWL
LGj3CNzL8acqbDghd9Y6V3sUNAPNosetxRatfxyZKFnGYiNfDjn3eMeQ0bkF
a0qMsmZ1eZkBMdhSDGrFX+nhG1LkA5hPDArao+J7aNU6bfsLlLSkNBDQ8c7X
JwLqmmpfkZJTpbgS55G6TpqpsDRRptlqvZtkGcge/hi7G1C54WepRD+oXTVf
UyXEn8lsdQfJQAA0FB+bEGv+rC/U+7tn29netTikAFHdFJY89jTzh95HCRLO
eBAlj7SlA3CeQOhwvFwIt2BmeK5Yxhdn+D4YFk6D0fRIgtBtSEif9iP2W0bo
tVddfveSKrAfIUcXaIJ+hw1W/gMoQHiYljXso3t0g49gPKBHx+wzy+lc0gfy
rQDUZW9gjGPo8JSdUlw9A107WYj1TMFs9ZMNQzZG7RFikg2W3m8e4x0JC3EH
I+y0C/sAApnyeBC0IpbTEZmkFBI5rEt8L+/iLwK3O/YbuBd0PreaCWWn4JBy
zcwnShZoNfeNpXxhbHLR/MzbwuEIOtxzPhvKUoPHwzYr5YMlnGBcnYHyVEjG
2YPbTL8N4b3B6VdS7G0PmS26KneCrVPhP2bv6OqLiOwQYF/LJrMEzrVwm7ei
hoME2BXvRp+ReXwwY/ps8b0tydvVvpXAHyGXISivcZsRw5hocLL2UcO5aHF5
cGjga0eeQEi6HBBg6Xi4p7aUGcYjQEU5NJoQiAr9nUOhotGN5MCt+QWtW46D
5janR7l7c3hJGfxLHFu02av/Q+GHCA8yHnQUJN2Sp8Gr3qsP53UjTBCM9nhf
Pi8s4ROrDVctQXy9fuMbAyYpc2LxvdE44vFLEujxERNge4cVMF/uMCu0DrXO
HxlrJIf8htupz2xe09mDGCe5zEXvzvYj7/n/s9E/010ZtTt8sRpUXsqu7pj9
0LVnK4GUuNW9Zg29KrPNuh5ZpUpDgPdHaXGi8p4HyeLpJQYuUUQ6UYv7aIHn
f7HGzmlkVMvFBaPr4xxcv/iNtbi0IpZKQ5XgkJ+W9Zgl3PvE47aLAtwJej+M
c0pl3GyJkk+pF1Ci8vSAiTxCvu1eYMcidcPNpVzP+n9dKUNKjuxd7zKSMa8J
v9L2vqohDa4lKSjl/6T3RN8OW0fufNRYHxTmy8+1TiwVvDNn/skvygVrFIiB
ljrxj1gs07ERQYh9TZ6G+PSzwNQGm2bvfceD4ovLXxp1o3v0B9DcAMl09FsK
Ep5wkpQYQs/0YSs7/uwyPS+HgsFSZEjAT3NCD7eDutvnOitBF7zljctied57
WoF56ukk5LxCPjc7eBCp4qsWSQdv7rKHi1iuMIHK5mNODOWBJ3WbtoHllSgD
6uyxrQc83d1FArPuuH6QwgJTbvM3rtRoB28nywp/hrgXq0n9Xrt4ABWe1684
sOX7RFVaAEHcRDk/4HMHQQZyOpIpLNJZMsFPejkPW31ydFXdvKIB6QO1oZr7
ntfzQ2l6R0gYkmlIbGqFJFuSlffQceSro9m4+icr+x8gPjgYU/IWB8QmWNMr
irbFOaGPKSCCPKRgWryS7dgLpN64ngx7B1mZcFGMDas0pWJtyFc/XqzC+f2s
0Ey1tcRwormCuwJNB4dZ1PPdjYVW19fZN00L1wIg/nJ9EZMNecOJ4CkE3c5S
/i5M57foJd7N/vjS9LK2R5hkFWWN/rEepx0EZOWJjRab8nx0cLBKoa5fKiKM
57oMcDkRyoWhkYDY/P3N4TV41WP+vR41JHE+l4KAbJZUNqM4VHg14g+z4gyD
4vPuczp9vQRUo+9yrAV6RUf/NsVS5F2KkCLPldNFdpLRFphvooEC+p+cYvzW
oMcSRFV8pgZT1C2TE3dNPCtyFwuy2oAnE2AfcMVSVO8fgZf/nnVBWeYADQe0
PzOvyKoU+U9dLYjDcKz26GcyNNeSHe8bKxSad8+S5Di5A+zh5zF+P9lr4ja0
G60nmxEVIx/50QlFWtJIh6M03wA1ol00BS7z8gG2jjZo+82nd3EtEgqwssja
3Q1113aLlzKnGXXpPJHxn708oMqN12h0KnzOVWwL3eSgUQpsHR2EE01n3nF6
VpxkjFBK+/iAUlhnteJN2yOLobCj9R7YMMywldgGU+DA+eZfYqjKri2+7MhM
V1yVc+VK/PNzQoi898TSZ3Icb9GSz5jCOgzUtFIrMVlcEl+GlIEL0RUpUIkB
soqiEFLou4PRMG03aSSQTiaSJ/JFJ+XY3F9CMAo/xqsRXw72jPgg66Ny4ou7
/WfrZZC0esdXP1eXsFTH+9ZSymh43IFH62C1TG06q7lZXglxiN7xXy9MSugk
ocGnAEHW8fDuFJZnJNIKhCOgsWuzaeZaUGqNgiOPcb3LgQHg9tEe8KZGUrTM
248z1h5CDpGUpsAKwox6MrhxzQpWbfZTc7sEzN2E8V2CNtSrx0aoZDxOti5K
7Wbqmk1lYpGGWGJ0Bf/t96c9mQdbYgHIDf4pauSfLe6fNyIsstM0FjHGn2RL
6jaxC6PJYcnWt7M62edg9dQ6aTVaY0Hmgbzty1Au3iGbSb5C58G1R2v088Dg
hklzGAskh2mfRGSM7uSkz3S8/ZOWaiavFGLyulChQa/Pdb8ZSM5angpTBwWb
lnc9UEwtLwn/3E0/QjI+xQ9luNjUA0lRT8PKkHnWI6SN1VwDdSWecNbcdWEM
0YmPzG0lDLyRA9VqC1vZN/vkpp5aJdTQXX0tWXC7CMnwCpKH3KXix8kxNbSW
Z9/ZNEaI+wppnYRjDb2jZT8grYOxKaQPdl2ADOYDbf9uEYoJ3y8W4c8XlEYo
gLEHYWbSdvpNWAbqCPpU0Mz2U4TkvY1IyHR6BUWIyIJPd6glYMJeBg2MDYBq
rCE874ATIzWK2Daq6WPsfCZ5d9aq5eh4Aak8hI0dhv10BwYpLS7njx7dGREH
YbOXFEwWzb3Ki+chIroLsbA5K9oBxgK/ROw77aAxD9eyAgSGWQaGODkNDNaj
9GtIzKBDxddLfe2bn8ql6B5R0tk3H+U6CsO0IwJTCLyPJ+nybhulyz+JP6jx
0nMZO1SnTZlgLKl9htEdLzkjc7UmUdxnXRfcrZ7bGSMj2PuOQYYdApYk9D5q
jyvik/4niP9vC7j9otgLeu7qVQpmq+jbHwAaDiqBcGYbop5R6bZkFj23UonR
ez3tu9iZhrudHZ7mF+FrMpdJBK5AofrGnWr8m80uVZ9cVWep3aN3Z+S2J+LJ
Ri+6jt2/5VGrCgDteUGoRDoKMmExSvI4XvZRPCXuTNdxY4TjDhVJ1WZ6h8mL
07th6TTXYE+c/gSALYVRYjc+pHypvxrNZd9k4+sfGLPhSZy9RNz711bBJP04
s24W70LQfQtQkNoNAriiRkzdIBV/ROwevpLC1JzMA5d2A1AijMdMfZfCsat0
ed/S/Y+KjSRAD57qCu9/QSmMFZM2F9x+Eu44DiqWzpKmCDAiMVFU2Tdp74DH
JWW37BEfQUIkILeEGeIj/0M9vB51w4feobZagBZv0RVe1irgM/tbSBJ4vEi0
cJg+0A0LYX67k+EmzVrqIfEu7ZS3Xet/2xAlHErQSQ2JTNhVobQ6HbCRCmPL
PXIvng52bRyF3Ao8mBxmJCQuroTBGovbRSJ9w8EmIBjFT5uJwFYd1azigVJZ
VJQg7TWBO3YHyJKgdudHOeArode3FVO+9XV2fJrmkhTIOZgW++mSdGYQGGQe
yMyNol4OHC8evoU5HogU2b3WukOZqLHrT2qTVugbXnYufDvgbs3d1OlRLssa
dRHCiISXqxfDDhT74YAz7py0bTFaRVviykduPbZxUhyaij9u5wYz50ZGTUsQ
JmX+he7t5P5bM88OzTlxbwd/xk33RXUlrtqWiO2uNxCHMD5PtFB17EB0JXU4
p8qsudjGOz+8S72PyIXO17ZLpAQ4zQy3zml08U2F7C0z4SwV5UzwNr28jL7h
lsqhPzv39hZVtq1CbgvYNfJtE3pKTfyMXUF7htUjy2zle2Pz3wK3sTpt6/He
xza9qfzXFnxWASLj7UNjlGTd35hbNS9lA8oH/DBWCE9kQr+TmmMvc7iV83nO
CgUte21R0Wi2KdIlX/kyhugRYG8Fq3Huk1Er+i9sZFlN3me3LMn1SF7D57C6
qe4tc9BeCe5ygzKqWV47X0daH+AOKrFT+gLYTuylSu1WlYjrG4tsN4uyl3Zb
+gtsJl8qw5mc05J09u4GiW1nxCseIB3hC6SrFFlIF7Wbr5ACfR6H3/iGvpgB
NkqWvcItH+mb4jM1BuPC2j/0gR9ACjd3UWBd4FR+Ck6dDdPpToyYEtwOEOGi
rIZ6bjSvLZIsxARgYeq+8GY4bhn78MdXNDOZGml38ygR110isaw9TRt6BRBs
UEPwZOmve+Hbdq/tG1ibJry7+DzZ9YJAYVeqfk65pdo2G4NSR7Z17i54v7/E
UJsoSeFLGDB+dEau4WIBzuqk9hIQrII3o1HiZ99dz0e8diU1qThoAYA6UZdT
YFaNztXKUfojPxn2ok3eJ6qUxxd/lFl7r8k+1A3H4f1RFn98Zk7qoU1+W2JC
MiBvRnr+LVzcJPI3j324ZAXyZiYvTJWWZbI0mUOxGkEwUCf4chsGxbrMXYXV
Roezn/vXXc9czC3698wf9447Uv1Ab44cz90HU0j71Hs84tOgue/2IXJ30KI2
kRdKjLCxUBrv9BrMZbr8s98Iqd/Q3q1W+2hP4A9AR/dk01YGh0GB2iOyg7Hf
DLONU2sKEuEIvVslrIrJLyJ5W4M/F3rYxNHD81qCZyuGH12yBARXClC8BffF
LSCFnspWjSDeJMpTbTlkTXaMHDPh5aXYJWILOdRPenBovu1BJMRNhJVaMsDd
MR03qiz2Z6BU6PoZpsENC+E1qahKZJSgZYoXVgn53kRn97Jwxma9fe6nKhrv
tWhOGBdZ4fkMgRHGKITMiEkbbnPjIRBkI+ukUROiDxI9KAm9DOiycd5loHhZ
ZzWiFr6chWZm5UUD//HVRee9+M34gpoal1CiygqvGa167s8Mmz+gxP80t++O
faASdVOZ8ug1rNn+AKclsG8k2ekYhMbtDoCw8t0I3EEF219HEjyZ4bVBD8FB
UtH0klqfo4o5wpG5GYczTKO7zHlrKOd3FOKmumWFpcBN8v2Rnv9+KgfqBBSK
4jLTMr6n4Eq2TLx+ytSEfI5eoxaY7+0rhgElS4uuSmGo9atovXvpvii1HnZq
CLz7nfrn99DskMUVWJkuXHcyouXlnijqJWIwr0dSxzMibIswLrOwdccJxE+a
Avpo/pj5Atn9mBSCiA4r6qF1CPjAXs1bBhY78DGXRHGnSGZHGSQ29DLP32so
kkreUsKiYWBBrfQJtz84OVzBcdUaEYhSfGoNCCDUsY9jEpyRAhOK+VnNh7tk
wPdo8iRLn+hB3alfoiL373xtuw5z6Jboa9g98rdD2Luloc4tpjW0XS+puGih
y35kIEO9HKjeQQi09bOhXWMaVvY/rZ787ZKEZgk2KMLBxQZ/XK2Yl93obSet
O75WaFRCDxm33bNy8oRXjMBlrupZQwBXa9jJCwlUUBYyX65oARnOTF2rmitl
rYdYWB6d3x1cj4vIDjr0FGOmaTsQ2ST43gmJ8wJts47jK/Nka3cwMIl77qyF
8Y67RM9OYHOp+2ADAg44UQQPZTcJMe+We5mbk9K6mGVXOhSB4R3KVf7LcYj2
zjEwXkROa39TyJte7YkN4gq/hQehmDne5uQg4FFsBIsIMj8BsxSORuUHgKWo
MJJuymkyHsGAiAZ0Ze/yKwJG6NcvCOaU+L2Db4vIU4Z0DkmSuMe6blMumawI
ynWq++znVAttRXFDl/5GHxnUprzRELIXrH7oP4Z1jWCWx1S9JyWTvOUOtVjQ
bqWjwF26DiLgzKTue8B+PxXCTl/EmBpKCOPNmeQVjxIdobXF8kkiMGhQCQgs
EA5FEYFW5Hm2u406mFBikASvVp5VZhG1AZC7G3OOafLzbddmMsKovpGM6sXq
Pdea4XnuNon6BTAeGmJ4iX/SPR/1wBOmaKr0W7jEt+XQ0Wn84BAfRjmAQGRT
8T2dIUByjKpviqAQksnBWWX2BJ40wwu8PVSOXl/b+t80pjpZtFCLRG1PfhIk
+UGBmcbJGzvso0lKYX28PwMmpUsDyzeSY61wl6iwCEmE6vWP4MkdpUlszR5p
whMn3HlPx5W79E48CedSfDVcu09wEMLPFNGezQue6BDIAmezwz7S2kfa0WIz
wH4VlvvJz3VETyNIUn6/F5MO0J2xWpri3zKL/9mYEIbjP0aBgwAhALM4zqcJ
nwjb+re+pb/WRLXx6v94BUwr62seVkvjOcajWlttrcm1vFNVDR/QYBdfLRAK
7blM27ne8fT/vnCi7yLla0rd9YOkGXM32/Z/8FUPmpwEeuxwwf1UJMRYl3jD
yF+7LWIvBWDOs7rJqPR0IC0aWtkKomfvI5t/mCjXVLzEZC1MkXInSxb1UGbZ
zO5qQPj/69HzWnYDkLMAiJmgyL+B60WUijzkyedxcWv0dwfBwRFSXNHqVcZz
kUeWVIOsQ4vVbSm1NBSxc6xu01OtmWnwl+ywsuyYYaT4FqeBuvObn4rnVRNs
pLz/JNUbiE9wgGHIRMu+IFuQLsP62FOJyfV7odVjF7bvXlIr0SGGa6zkING/
xKUSoUZ2vEigU4647ZTElAyaLg0i/NgugZkoKONpMMmNxmTcVtMLrdAhBGj0
n54f7Ss9q151FZl9NHb74D5Dkgb6iFwbIsj4q/TzVB0AooKNqgtbRW7L1by1
14D2WyCxajmuQ5GF1IafKhUMSfRTRsvwFaY0+8JBf2KuXGYR/hcH34it+bNq
sRH2Qd79Sc2yG8JrqpRezYQRe+b9B+ZXOiph1RysErXelRvtBe8oWVqBQ64w
II5eDWeIRw5iBZqjCOZdDgOcs+aPDQ//9Au6TDD/YxLn4CHrx2xiip99tBM4
hyjFfqWrewpjljCYY2aXgoylV7SllDYYXwdPG7gMsrsLit1Z65XhYgYciPVV
v/42wRyR2ggFsaWRTCQHs9YdlDZ67vxLdMa8F7vvNgNDldzkL689EolcEuit
onmwfqPMVQ7nfC0U1mg4RXx8UxRxrYbX86ae3BapCcap502tR6mik+od39Hs
m4bFBsoTvx1HoRPyT8fneGXtIe5Fd3XxngdkUD7+h/2NpMTQ9x7NzPi+sMu2
Wk0R8uquF7IWoYOuJFHkiKpx0vKK0cE6gwaL2kMfLlMSG3j1hgfPfnMLY3j5
HSBqNCaFyxEu77NIqblLKpeBWaKEfqaYDrkTtzm0qd5e2kyXRLqBxdeIUFEh
8ACm2jvW1WlpUNsaj+S2fP7s3cjigKT8/n0RSwkiu15M4QMURdyaOI84KSWi
kZGlrM4YZbzL9f6pH552QherOlV2yjCV0byDVT8Cif0mpk/ePyaxnKOzrIqr
G1zIIU4uR3c794EDQ5VWR1os2jhvvVMhYuubOaJQxEt+cjFF7oB8w/nLjx0h
U4hc7XZrpTBYRh/3lsjgxMec7HX2COVKX4p7+WOy0ci2u4jTv7e7D+Dl+cU9
NBWdbqVEVZSm/5+odMmUMW2VIOby8eLHQaT78dRxn8dnYLTUOTF07AI53FEP
bniL+1JLnmA9aeTeyM2vIpvX2h6fODJb+aFk62rsl7OFMZvNHBrYBJZdneJm
Wo/vgFZuFZ0RoWsyZUipVN7PrSw6REgXT1Z4wpDRBV5ocVKpu6lZg8lznxfq
mykwPD+1u7TDM7UM7x53KoAJ3U5HtZjrwtwTUbuSk6EBXiUsW07Bhbw+dUPF
SQvdBVTKZg260K5Tixb6NLxGwxAQZFT2V6gVMOYDYdGgFNwzbbQYnAfpBlL6
knci0i8J7v1qUqzUO9g1hWtAz9IlZpYpbX71kpRJfZDahW+ZKOuJJRUWAi5P
CvvRXY/1/OyykQRdBtQgWgrlgCsa1t6pjOd1axJU9INEzHo6bmzdMDWcKNFU
dbzkbwEr2fAd5W3VxelVf39XNCgmdEAYZurF3LKILcU1zuGpjcmkk7LBT2T0
vj+HpQmVy6iYRqnS5TcQITdQjhKdW8my4vXwPVAP4e6P/nDBRTk9/xZ2Rxl3
tRidD2U6v55+6k1qBoiS/iYxnezR8KvHz62nHD6uLCPa1g/oW34gwphWjgda
4RS7NID1nx7e2cQS/BhDQ5abmpcIclB8VEvDBV1g5CZ4jngZ2RJSF/vYynQj
IQEcVYdYd5VAqWMF8dBYZDSXZdZoqrDydZovGdJh98Z+7iTVC9qLEDFu2oLC
9+ohzb8UIt+QrUcZPwQS3Mu5sO1j4mmbnKiTujkBH7kHqlQdD9SRw/h14EqB
xF0FC1M4r9vs9YBxVsbpLjWm8zci1d00I69s9PafCCKEUOn//gOZBK5bzHZO
zK+pNgdyo75ZiUB0fI64VwHTD6f6VcdJHksbxzA1upNu7vsZeNGxRW3IU3AO
UpWHPCghG09ErWeEHfyC0aT6uzoup+rX8BFWLSviJ8vSI/8eUpHtUW1/a1yO
GHUfxw9zdRtubti+Ao0uP8Mvu0h+gogsxYN3kMuLIodX8jUOx+NTioNPvzsT
RrqcPMibouRjWWYOIOs1pdvbLg+GrqGR5N8L2/twpRuYhsBomH+QODIwmbuu
CNlNFwQ3IM83tjmkDPVpUWyjiVR8ftvBAUaVT7GLE9pgda1VaSzYpZ6U2I5R
xP0zpV+LrJ28FBzi42wLSLOjhhmjRDFvBSjyj98MtnL1KYMvyjgWnEZ35UOk
LAdQv9iXu0QW47CpHq0ZJbRgDu1LUABwlazc1rAALx9nPzrg1E2gHzcwkzGp
vzZUvaHPM0xoVTHEBS+8egC8y2HJZ2Sgpr7ZEDmQPCwbLuL0yx/bDmkvxP31
Zy5kbH1KjXkc+a8nNARv7Rg/O8tCLTw/CW5uJClm/cHTUlpcuCcKtPTkUPws
AVydBkFYRtrRHtQ2VKneDqElW7zRXssfi0GW5MqbFZtYvYXoajyieyLkJ5PZ
UIk+0WK9rGvtGpTNVto/0c+YeM3adetzr0nEKAX9mAbRVTvB1DwOdvBsPmCs
YJw+HPuKq/cgTgVVjp9WEc9nwhnAyZRn4dOyaXM+ZGWSeKFKirEHJYqgFU0N
sh7pbVLXOosHYItatTHPHpUO/OEY6445INpTKntx+ULqLYvMbDm1qFK/Iplf
8XeyaB9UbuMfv13IKu34Ygs9bFq6F1dFPuncNxorTATAB0zCS1eLWxncJ5ox
/R4+gbClLSVgc6L59iPCDuQ4/QLBF7dJGi4N9kKjAoiDhpm8YxWHZA/yertF
mTO2ilV4HqThNdb5aOLjmGF/8HtNOJlVsZgPIqSGbFcccN73HWEDEU8r9gON
IBNEEy+jQ4mIC+EMAZLUAxm7gLcvhGN1pqE7VMiQMLb1FipMw2NQgnxJtLTC
z8CjPoQFyaNDJFX9pOSLejnaC38tbtxFgBwshjPWU6UGxBXVEna526K04oZP
bE9te/K+XOfhKuEqcVqKfcOcSsDJA0QIqz++y40VXAAOHrmFils5GzGpmDnf
OeRPuk2H4YM6UTbRO5z/A5Ecs4H31ZxY4ffsnjs5V6TQwD0UWOME6ArQQtz9
lbMcgVaH/NvY/R4ueA37wOba8bcfPXHV21E2pI9rVPlxMyp7UjbFUeyAnzdt
rab9Mobg28c462jiPZe0pYPZXKNFit4On1QOEhtbgAV1t0RxFGyChB8BuBbL
9rYLLvvMOKOLs1Ly5sp6XMPzYZyj5aDjcT1B/wvXdcA+5dwMaQYbv2Rpeyxw
vbQD7FKM3udWadCguWgK82F/otR5gUZxqWQxj5KnV656Z8z1tFtHolm3czd1
hPHMRdiQrc46azB0nb4YNx/iFI+iJ7HtlMtuFj9bEMsieTQWhitW4uOu/EEt
m8PF3dK3gLZDYsNYsBZ9bYKOKzaxeqhYhRFyUkYGz5tioBGg+9jaJr2wtG2+
16qp6Ej9qlpu6EVTv5ykXPrUVPigzojmHjtp4Ww+MdD+j+Kpgt4XTMZQLxEH
jVoYb4n+/iqUffLFxL2jjQnYYCtp3wDFz37kWl8Qq3BAFWZFHHeqBLcEmH68
vAnQdVHPpQOwi2w+LZ0hbHPrxUILU1Ck9bkEc1Ep2mQ0VQjapnCKR1krSLTq
VL+qKAO9eK5p6t+stNBfTNBUzIj+ntYlvD0A1eB+Uy317jnOK2RWM2rim89F
n39VNtv6C7sCSzXUzLrUVpyVnfrd3NOL8mG0F4/EBpllli1lygcAbAJ0TUDj
TOh1LUOhVVCwj8k5h4dYKA6GYLsQviYXQn6AzLgfTDB5ynPbwCkQGo90tTvX
UywzzElYXAALUs/NouMnaeotL6ClOMIUlUIqG7uN++JBLY//XRObVjUuNzX/
RitO9QJqeJ+DugoEL3ryZ/Yqv5ms7rce/bsx9ksMV/Gida+YwrMON6VevtLd
Xzug9X/K10BBMU3imD1uHMwdovUtdY83Y3+Wk1iFeY8WeMTjYykUOWQnfMWf
KgRO9lLi9z00eX4H1HpXlmpksI1r4gQC7y7BOQV6WqTZ2pZY0DOGit0V5lE2
M9ryxKVp/SmUp4NdX9ZCHuiPh+JVTqJJd2CyXU2PMzymX5uziNZBKDJ5v7P8
i0iwM/IJw+CWRjZMT2O+vsjMqT4luJOM99cXlUyjlSco0ySLS72NbXJysKOS
l2/woyjNpC/B4zA4agjE3fE2KZYPDNheYdOSe8TclYlBTskiZ7JB+qFraZfR
F4hFtTzvoZ0Dz5jkKRgeUhQ4SH7ORDRsuGPyADlUSbMFyRMcvoEuL3z+yXud
V0SUrLHYxJ+rKMF0A2DJjWOJtxQyILIuoeClWRScJfzzak2ETXg0ac1gcBCV
NKLP+0zffRfQ7CLcZ8Fk64WGi1DU7IOLuZ+MVe7L+vCn6I7KisD9mqBIvHQe
M8lN9mkdMz6gc+rGZE+JjnFHzHx8gaP8HOcZb6B79ToYi4FxTV3e1aVQMdXr
lZP6JT0bKMuIq45eswsaCP/1+rS4cFsThWjhBfaPwocqiQ5KOntN48BLvw6x
Npu2cU5djE4xm2aaf8Yjd0rjh7Y6kyKmCF6UUM3xsI16szNAZ3kLmwRZOElK
oVpRVTt6d1iGKC8EfBpV1gEO9VirUiAuuRw40x5HkyC55aHAVQtbM3UKq54n
3ojvsGhG4qC61bgVqj16OeNDOFxbxmVniPceIhX9tZY+iKIBUv6kyNKlBPsl
K2QziCX7dKPURy1VEHNNjnnO+ujp9sSAbbVfhP54I+TFhwMSTa7OzN2Nj8K0
4b6tmR5/v5gbyVT8hUh6ZaHa8YrgOhIJlERMaWl9EaaD08IunUOfJXU2U0hy
tttluybQrbwDNrEy6LyPYJ3meHGLoNHqycVEbSLlg1wNEDn5rB3i9bKMAU5N
WlBD6iSWoD2px9H7mA5U+BsMFQVijADshOsPJTM1r79n3hJvCC73aHZ9CK4+
tifktPJuS8rnTYm4O80qqSGJNGpIzuosk5nuqldPkbv/5Vh/BQoyZIoLaerW
KNtQud5ndVTxQzMaafj8xQY9X4EkwutkYS+hlMddQ6wOwd3OCOUYqF3Oo0AY
CflPjoOsa+dofHBu6TH8QWYb1OuUs/FFA5nlIsDSLQRsZ2VCiZuLdLoXJOtd
Gy1zbqr5m0yvpog07OhAaKfV8Nv9k2JnqqJpBf0B77E1nPMP9XUj2a80Or2i
P1R3sZRkZBEfF3/DNxe3MV7Y9e6s6V/013oK0asRmApYAyr5V4kGEqOSj4Ik
aY9FHcBCPOOUVZ1vgDoQw0LL56PeWGR0zvB6mmgOR4E0apSerZngqqZT2SpP
yofgItFHXZaCdGJ9AyJFQGC808lueQRZamVJytyCo97sFc7zvbUhqogKMIYW
bJNkaPl+ps5KGFWjLvJZ9/OpX0XoSqmZk8E4dw2UXv+J4IRvrcSgUJ4DrOr7
z5n8+zm0QYcqJj62xmYfEj7BgZsVHzlva2MFixsDU7WRF7g2kehBBRjg8NiP
/HvBgXwGMLyisXaqdXbc0ialNz5WDatj3wndBTO2T+RViuiCpheIDYwGBzcO
cmYzAVAGE4WuEA86VB5G9I6ATrHqk7RlKHFSUo5WipVgnfbvX7+At44nKA1N
LEj81mzYR5rGOUY5M+9HssAS8/L//gkLaMK1kcaOzhkayXnW08jfq1NBT/HK
cbqFEuKwF3LLc5oSd8SpKjGEwLrSutldnBk27WsCdISrPQ8SZ/aay8RdDZaU
zSYV4iM97+STVs43P7NQb5Li/r2D2npQudYuiQ3vsDh8T88zolVy8CUJ76ml
OyBnTLbLMqDQMM33vgbMFBiDIKpRPjfnmMdDXiGdkxH9MtbHEoFPyn/YhS+m
vWREkdg7EwC6f/cmv/Jn98Si8VwZCfo/2uUzzHSFamkHqqVE65PRyvDiL0bd
w3P8pqh9e+Onnbm4qKZnSe2U4ZVOTz0CFGEwi+C9O5LQ8JVlZSZNeWEQvoAT
KwMUEIWiiJq+VixEIpyGJeAWRGpxX++jnFp8XxDFvNmpBNA5TNMTbWpaNBU7
NsXNdvtJ8znDL/y88yPnP+yu4egF5bPoLAKMUCw3zTYp3tergacOJ8t6jfdX
3u6om/E5HJTUYYu4Aoj/+TVhMCbM1RnlVPtuEaXWwMbyYi9aq0aFnY5cg47x
1yDggxEAZKNCkrlwh/7N8ijxk2DP1507+dr6JvN1jg17rVoynyuU6i54mMhs
Zyg7eoE8whXu18r1ozVdsm92SY/FjnRsn61JRmopGL0h1cyU8ZEY3LIzWeyN
sfyUBqTvfKVkHCkVQ6SV+IM+7pb1VKOyOGpPY3Qu1kCJ4/qweBziIiBk3mph
y5DqHhOXiC8vpQlOO1tQFQ4C8b6KwhduZUlhRjvNkwa/r5N/HUcPKpAGLfbC
G17IR4MEWcv167lmJj9H+/TQIreSr8jIniICwif18EuSBr0149ZVk97/2Czt
DO0GKB2TAp+wqSjpAYaOS3DRSXKywdHsfLDGyuIdfnU5+QX6CcDNs8dnZ+u1
U8sZHgZjULL9xerf2G+C4UJJEAdQDGaZd7Yru+zZ/6suSAYiCcYS7tnK087U
0VXFHEqgozWA6wKFfDLIdQh533PaadabUhKxWyfTr65Ou/V/cUfNOpG1h1rB
2bF8MBIwgW52mqGRmpuHKoczJr9irWSUQ/M61M295CaRcvQG20OS4CUw9os0
JHCftC+yElghFDRBDudAaaRa3wygpv1KM6m3BPDpwWNWXCdTrFpYERfUTSuV
E30lz87MhPL+T94cEA8rTxkpBOIdBhoL4w2XYq1XQrDuiOocoy9OoXRpyaad
ZetL/nNifh+phCfXSujQm9rG6M6+YeoeUVpnp1V7g+sM6pNF2cW9S93C6aF1
WQED3RiF6aYb9hu/L8zTBC4VwxogKrKwSojtWcGjlYdhkY5hmGZ3vc9QTrrW
R3/snx0KVNj8MiXMo0izPhGDveztyPYZ7HwM7uws7IYThFOvNEKaoRR+4GyN
479mlB55HStSnDrYagej3UUmVE5+V56FPgiNqhlOL/zLshngo9s5Ydk8ec4u
bvJxKA8COT1GTUj82DcAAvCG0wd73P5zoAJRLcU6z8AkN/mib0plUIMBA/jb
gFeVUEOOyqxvFITMw6KEq5SaEupjP1XqI9+ssKnGfhNFPceKUK14bVAowQSF
a/Ysrdp6hmaI8SuYcw7SJeGPCjbRoPf/hWuvU1n+Z0a/EONp2I5yx4SzCmMx
npw7A59Wx+r1DejsD9VeioU0uLLifNyoJJ/eBFYYtn1JoCzNz1adz0isIPTp
Im7B+yvBm7xlugLd5OoqFlNSlXLiDRibH40flrVRvU+PSL6X154O8o9UTAva
AN26ozBb/SQAyACMX9KFpYe/9tnkc5YPTrTx6lR70XhkAEncTnWNBQUPVSBr
J5F7OqELhk0Jp5QB8t87/PYCyDFNEIjeG6wE9hoTqD8h/kgpKtyhzhHxce2F
bu+nVWqq0Km7WFw+eYEpIf+ghEzhlzAjy/vD+p850LTDewzU8SuK3tp6I+l9
2r+KvITONxpTuRIJKukOuei36JdM/ETlsgzQ9eJuro9LCVnlqXANxQmA9Cxp
WOMr08j+JKx7Zu7sFg1r+z03m8yHq27Wyb5Esk8RqT91lD58i6tIycmVd3Xu
mEmOyDexD+QJLBhfHBgYHQbb5ZGDDYSmJQcAICwVlZBXmTfZvuqb5eqZQGvT
iiXCSurrmlBygXXkxq4tDPHRTxWPwNKdiWUlvKf1e1QAJu8JdxuNsd05NAU/
LA3JzAz9mWpQy2ZpM5fD1hKYA110n7QaCGOreLv96ZJaZ+pW3jWJ27DBTIXK
eKYfIxIRsOPFmmpWHxGG+b+iaFjkhOFztQnDr2Hs5goXUTiVRdQna0CDo2oR
w+mPFgrSaBK9YEnF3BbIjEuiDnvPeFVc9mA0H1aVa5pEPsgJ1KY3PcuifTUy
+XdHFniVL0v0upqA7q/DVS+DwjJc9QdsqPv9nw2ug5VjZFhhgFJ1yPqEbz/Z
CPEfXEOEPZY12ff7+YL28HMuvQ0jCKOCk02yBhuDzUK0F92gn/X75NppygQ6
dloM/sHSqeTl25w950EVqS620wXXzISDXt1jvORk0goRHxzq/qZsQaMbZb6d
HSF8BB/4VlRVSuSX926zqvysgw9mz0fiUMU+pDd58nUOEUDu4PmHzIFlxhOz
Uy/yxGTht4VQlJbItb5GyBmE1nLFLBDsfSwDOr7M3eD1U9UuvKf8YzL85BR4
CCle4AgUdyoCAkuKyuEpfkmLJkKaBdI6PLPLc9lEwR6i3O1+pJq3w+Rh0O2T
5EmJqpEJUsxz/ngODiRr5eDudBBlMNTSWau4nrbdAKTaa6qWiAfHxl0hzO3s
SgB7s+TqXITV/npCGSvnjFH8jRm04IipahaRYE3980fe8N2MAYC+kF+L2zlS
f4tQDfAZz43mAKNM6edVhSDezhcKU2AGT950wLQmje2Y/iiYi6n8WW6qp4ml
Cp4s99b3qymTkGMX3RrYocmVg1VpXBTIpReYdC4SxkiHtFMIFtScwZsX8lfH
Crfp4gn/+65EYJmnX5KBIBNDfWOWhF6HRgaeUvKGE87TFG9toBOSF2apXs/o
DIX9Oqq+RDC6y9Z+O6TJ0EuKBas2S+6O/+SRdHJcmjd7DceB3K6/6wOhnGKX
0AeebBqN8OPgTpPT0DEjUXDaE6V/z8phD4/dJAjXJHI4hht+88jOqISNSWTE
JIAFPLInApkF0hLW5H8u+OCZzZrlVfs72f+DqAYlp3YAB7Dpad3GjicX2MUd
7sOd4wrD7zRsekgYcmYaafUd8gzYP3OuM0tb28EEOOWpdclYbVKArAJywfy0
qaOSkji5STzEmSoWRvbTWxbq3Q8sdhy+bh85XzwehgTXFQJPtM06J6vw+dz/
dP8EMY8rPXFQkzg+rvamS2bQ9LQjjfFGiV4sTOh8G5LnvSYZV7lBX6lDGIeo
+5tH2jHVuJXq17/fF1C4PWDuHBNqoTZPKgFSXfXIdzOBd7+0mMGHC1YattxW
ZfWKtFdbxjuLbv7Xiz5Dn5D0x9VPS3Tlmv/ID0pizAs88i8jEcmG4MMFGdgR
DeOuZQx6vQyKAmEd5INPjuKd9/6f++S1hZWO48sVfQvThdYZXCmPCy/QtjIW
IzQrsJjy1VGAmKrFLNzPUHBzvU/qg6hk6lyXVZen1wW+drvJDQwHc7neAe5a
iHy0aqUE7l9KBaLlYfkni2mfJQp8SBIdpVY9C/R/ejn3cC+N1KA/ygj08nhB
mp6ROuz6aLTeMPmKID+9hgEyjl3jcYyrtjmWZfMXVovAeCi1myxwhtyq4ejV
960BMdqZAoG1fggjYiUV/PCRbc1YFuhuBjP09cIbYU2bsZOGLSr78+q6fZ1q
wPe/wccMuueRlBRmGS1r3T6v25ICqacSTowxzHox5MwDZ4n3pFX+CRcroVO6
7DGDCXFlOEMBlEw9KfnxFe9t5Gx2mPaqNtrBfFBe1FU5Y3tPbtAXOozoXimI
060da3L5YbsJbL3suo0iVIHOH/OVOTa4OzvJW8+JIaCbJRfL2+8ws8RM12ar
suXCpTkpN+aihPoCAHqquYyDp5DPn3C5kl8MbAErrHXm+bayQ3ncVnWgzJe5
23vI0SA9iWfkiC5fTXy9ShiNZ6Sx/toMmbPC0FjVJQrb8XF6wrl4rv/jD6Zi
Nt4glAhmbzVcki9HyOrLxrD4Jocbm2RcI2kH+Ei4cM+hPl7aH2agl0iGMeph
jwB86CXP6FYnJbCkSYpwDDy+2jzKynVerhx2p32hIkBTtGIRAE7QfrClJrPT
4KUi3ofHAds3hNRoOOufwzObdr9QVMXI+wfvNLqfVU6mD3HXhBtnRj030gLv
4L0FXJkIlgOWGo0GZYrgNV3ZAAjfKQfowQ+Ch5QFFlkxvjbmNHQ0NgoQsaHH
vqZQQLUdTEvuSVTQmBUFcd/McyloI99DhRVY/TmZOGDLpvuZfn0mGTnTVVWw
9p5a+t6VJjFH2T96RTW25qDt2JBOyept4L94mSLk659YD8rOYOwxy3YPa9Gm
h/1MszjlMIyPz9/p11ZfI8ZUUYAVg8AeKZvHgIw9HIVceQVpGwKH85paMaFO
KLYMC3zy8Hs0LTxOiB999DEaG4bUdMzA5Kjq0dycgHN2x8Wb/RvGmLRVvGqO
FLTX8X8KfNQflmZcVXgCrjD9XGIzVGkb5dv8dUhuGIXeQ9+ElQt9Yww2ZFmm
fbRCpUTJXr45vWc+8MHm4Exwdkctk+VRyNqfzsfF4lpeTLa2vfF5s4RwBkfp
ISnSqAHunfkjLnHf2t0eA13Lyxw+8/88QSGO5/lNTaJPBlnV0Lnb7d1k5OHj
XLZmNrgLAiuH9DZa/jsrV/DsChfUV3RUPbREk5Cs2wsVKAfd3BqEReShNvvE
R9GZAJ3PttgcCj7PmUsu2coESXb1ygNC0atOsdVkUY0o9/z+NX5VDWD6EF0U
XLwLEI/6aqLjZopfUvgGswvh84vt0iUiKiir+T7S1CniLsX9BExjz0BszRw9
+6ENlAL4Hcygm1JJd1Stab7vKi/bOHc39ZgyV77vRQpryekkzlAfWgjW5itt
b/cOtodfRQ0/cndlMXKtJRgbsxCTx4D+MBoaf/WTDqmtxDx7rn9MoTkYDBck
95RDMr52YNAK3Z5MEIP3uRDDWliNj6CNAuFR8XBKcEwIvmZVRmgQK8vQNBXK
ro6gbkGMxgTffgXh/1nuw4uDdXT8Tw1xFal42E9WImxIDnXsVDVTf2t2eTwP
BZczxHUIomuDsxRv8H1bawIbirEOj5lUT7/aUpX6oAiN5GrdEda76Z2lWIm1
nMHDn3bjvtbqA3e8dnUw7eM1TyC4c5y397YLDFROz+R4TnIg+GeEeyEvjO9T
6O9XFo/zteFTdBrikxUZK93yGdmyFwJQwAZ0+8ZHnofW/gaRd17Snqylqm4T
zeq54Wr5MnByQnpES3MpkuDQRb036nQe8Qqp45CZG45ipyb24/Jy68R+uiT3
y0y9efq4gEpGRDHxRtm1EVupJ4HpUgVNvWePAVD2PvpOiKykJMVqqFikfh91
OD/3nEL8yRl4tQEEIDSJAUizgFtVfzfIooSrDIkDLkSKqoQoTPk89T0ytrw6
/fACLa01GrGqTx6uvN5vHT8nUQJh/sTLBawglD3Qmsf++CQ8PEZHBTAi/N5E
M5Y1OjggaH3ZysWVumAF7oEM/VxdMAnGrflRfkc6XNlPOw78aVz8+rl2atez
xDYVrcc7UrJh3JEHKQEJ6YnOzX2LkB3le7IOXhjmA1TLWnMorNP5U6kd6eEY
18VnKYixDevcFTYk7flC6zk451IIkt27ZNmTMwVUrrN+48MzxX4PFosFLgy0
c11YW3UaqBmIjoh+82u1cOcTwEoKe2R25q+30S9IL85XOWgd0aGbODziGVbI
M09lrDoda6bCD33zYI0r0o0upwYbXbxR0mlHyawUi9D0Q7lI1LkKfh+L3cn0
SYbMKTzTXxu6gTGDmV4XTCH9M5wvQaE+5R1WvwKrYNQe419OSPjcaSpgh6am
esmS34aeQIOZt3CcYiFTjklyzxSbwp/fC6XW5DuDfz1GFGL/1qNZtqDQQeTJ
kP1TgiHlzPnMoFp3+3N2pDDlGPOeaOIyrEVtjYfkZGpmQORXyLG8H4Cyhfac
fKlAeJs77XfDNDjQjLgH9OFw9V2TkbYwAPTQp0Fqt/PHpv22FHpw/FF2+JuZ
rC4vIHcQV4JEYLf3IPafBfQuQ/S1I8R+Z3zLr3mVizacZRL5kgUC3cwgS9WT
QtXg/klQ9BuOc55wvUh1SYHPi+5be2QF6P51pJ9BEeuaRKMT/7sYjSTHzRI3
FNEwI/QUHVUxr40ikg/C/MfAGd2tGYKbyswxsYFYLvXE2YkyMkAqODmN+9Z5
/gtFR8hPRKjFlowgH0voHXPwMt2Ey3zRqWNTrNcUfugUUFHyBsafd97EAQEu
XC1OOdBbXu226RSeXnUv2h+Aky6e/nMdF4lhFpF/TVNzpm+o1QQxmsEIRZzE
5HRfQjFpZKY8DjCbr0rVWspsagkBG6TBBSsVeBTTG4XttjgfMiynjkMsCBBl
O5xaM4P8lzPHRJJYZ2gx5W3iB/Ntz/eB24BjblTkIS5QXzaAOxmHlOuxsFfp
k2S/6/yMzF6dWwJzi3PEoZz7tivXfbbrV+0BjwhlNvEpClucdX50U9Q6VCx5
syDbpDYqRR0pNa2isyec3G4vA/r+Jl8hQUu5lgpfI/bdXWwxbj0MWfhllyHB
LO5dsg6ttuGyy8mVO+ywEIXIz8GyiKS4W7yePT6QMOrPXpdFPMXA9y3cKdXY
HAp50SK9kZ3IwCtmwDN85v67PbH74C9uMv59s1qv3mSCNv+4RTLXH5Vz/DAG
w1o0xPAE35g11CODQs7v3NaRYzxRFQVP+Wdrvsqlwaz+Xd56G2w3CYsngyrB
qlkB6qVrp4KIeevlywl+x8d7HdHV7bdCH9i+G65+8etQrxG9V1QaBo4AP/T5
4noHSd64oVsBdm0TS4fJBwcWDyelGawWnuZWVgIYkRt72SdWmnXdqjKdQFDt
3C8eDrkrUESL1OVc6VPZlonP1FuTydGsWhmSSdNZ0Vf0E7Xh9PDHqXfE8Std
FhGEjDSGhF0zEzvZ2ZokgBiqXu3UPOfBdJcUIM5Lub2r/JruJeI0Ro5zIlGn
S0shnCeW6GNXckNX0yiTU9WHkHkdc0E/VaN261Ld6B2G6GTBDKUNFJkKpSZY
gvtMiYbrbpVs1A/t1QmeeeDyxaXTd4MIuqmhmeRUnhZXvG3QbX5ISFtCyZ24
8jXGQmu7OjLwgKP7fAxDD8MYsU/k4XwRd9e1gcNQGfp+eUeY8dobsOV0hkR2
G5DNaiewrPkirKPooYmsP1F0bIebsdJiJ3ysX7xu1YcxcWIHO25OYMTG7MH7
Un7jQJmC/c3EnBGdddHbRM6j0LR/Sfc5cuGEJeHF8AcEsoc4F/U+H75naJCk
reeZbrulEaWOEKBeB8pS6/23TzHy/++hnpgsTZkI43/FG5Mbe2rbrK+hX2+I
n9AMZQrDvrUUhYMo4jwKhcFrtn/8KnrZfr+NRDsf+fkk1KCkaHXRPLQLVsNW
L2An5yOMncIG3ouZBdx+6ME7Z0oR8kx5XelsJekRRuaoi+l/A0CFYTNZVNiK
ygZoLMeXouttA8Cy0BJo/9U9ID0dlS8oyXvPg/Ejc0bhJJpgkDB0YZMDyWDH
YjrNy4tsr5hCBH0Yj/EZrGH7Vtb/+NFIG/FErsQmJSTT38qHm6ubgQzCcqBv
kg51rz3kefNqNIZGIZx2GgOxJuuCdPD/LBCz/szHWbm8HnLvFlFK9zqzQ8Jm
WhraFLwgwDFTXwSqnP78Ld9pb6Ryxz3rYaYSiSMBlHrDceGxqQtBKil8ZCQT
/69qKrAcSIhIdGxMbjk1y+BmLbpNMeNGW+yIKhD1NsYivOmyCa+EjdGG/zCU
OAaVBsiPztY1EP7zkVaaNZ4mFAS4H8UPjJt1h5HAW717+yzck61w/CisHOhx
dk80ZmrWoKE9Pa89v2ERW9YMn/BdfVZsOgTcpuTVB3dN3wg4XB8fvlYxCLvX
FiFjS+EW4ENdmVV1OivxMw0KQdjZedCSDAqciq+61HnrOpY6+x+ZZqWMFqAL
Sk6Ixbsba8w1eQk89bFmG/tMuItcAxOk2udQNtwKQsHyashPRmm4iSkkQabm
RUiDxaRRRhHoahTWxO8uarPVnmsDZdzDwLHZsuDz04dlQypNvfK6f1Zr7ZlO
0dX6JYILcFizllu4WeFRhaZ0TQSxKsuAiOsVHJJ2C2KHi/XBfDuFWprLjKp0
bFp7wx4rL29YaZNyLr5IrxalLaBJbEkHK5WIQeNI7byMSTl848E87PO6Jn/S
t4OCkMC4DcY7X9FnUP4KC2AbPWvNT0tTDKu4fe/3H+uh7yvMn4l3vNnBhB2r
la1V5+H7HoBLRdH50JX0n5EMOWZnAzvPEx4L9eBFbOcSz3UouP5mm5TOThWv
lsst0O6Yg5c4zdBIU/HWsaE9oDg9FZzYyqYRHqeI+8iLQiCnSk84llUwfWsO
j08d5H1JBP0qmDXPvcSSN9zjBfdp0YKqwP7MHkIqwXo+GhZqZ41WNHomOclD
POolHum+Rb0y9cuAHi+Mz9BrlScqN+iO9Ka9gQpOtvI08BPGil5d392kRX6b
iAlgmfGZXWpaIzyS/psr2WmDsNheEYRnZlIXwKiNeaVI0DP6CEmx1/hJYgF4
XVOlFO4LbX0WOdL6yy+VK1FtAKnKAWYu4sPg9nKXkZ6stRk4081jOKr2JLtD
r6FfzyH9jvrSXQmBpv3jXOmrJ/eafYqgdYV3tgD7QibDkQILZ3KkOW+dHSAz
J8bcvuIJ1BUrO4b8QTqQgHoiigqeLi3LEkKRdQjeLMmMgBH8F8g69qFxaXZD
MTMNBxSP+lZ5n8ozaRC4h+l5jWnoN3KbzV2on2FjUsHN4cfu60a1veioN0qO
lkU+51c/dMzRK8/3i9bs9XRN/YMEu+zhJfLCecZ5Nhl5PZurxrm9IPfAauz/
lEh0WIRrZC7ohNYWgqBGZotNLQnbbRzn7NPblnqP8ZR3B6C/9c10zwI6Cv5+
omTvR9keoV6SFo6RZ6a4hYTyTYTe/uBMG0Xj5HOLepATj8Myj2enqbZKwc+6
VicNZ12V8L56j+kk0YeAxbBxEDqEwVBFfMMYjo7EVYmWJRunkN3PJQBAMTmr
Tgc8O0munAW14WS5MBF6QOl1lDa9Y6lS35o1caRtD53XQGK/Q+A7iHqCL/ey
DSTdT5akRSq4oufpMhSEAfAMjnuhISe2e/V65WtbD8uLayni7IfeCs4Py0mJ
BPPe55oE060MX0oMhtUhLhfb2GeiLZECFSNHvWemxKnRJ1LQk5C/TSszFKMp
JRegns7yZVFOaAq++T6wpR65PAreKTeZzUgB0zENc32G0Nsglk0BnPfCeFrf
r6UxVUcS89HLLconnfSjCRnJ5lIxqnM7iDTHKY3ABpTauq3KdD6VsIHrS7EA
BQ4avhJmfehdiOwMIe77Gjzsr+0dhCKrK+edsVNmhT+qQf1dvpaefXiCYRot
O8mY+EK0llF+qAP17rX1QX/Kq+riHHv0JUSrIRvpcC2z0krmlgtcXafvJhrf
8PiLZWLPDnBiNTO2OVbCTHPRKU2lvyapcp9NYnA2c8Q3AkH2wHsp4VuSxj5K
PLk30yVjSZOEl4yAQIEABwxbsPfHiaZ6QcF0t8GvCRQzm92ykB62iFydWCIF
ncZFEfZLwbhuSqq9KPSMK1BBInJ0ILjMC43j5LKR/Z+b1MyIy1KwKmy4bfTZ
evbr1ik3BMCv705y4CBLUvzvxm3iUAmQZHwxIMXcEpnYsooQGzkBIVxAsNZD
1J+UvtKzaM2sFLsQOZGv2kYgemd3HpCkPQUDnLblaXr8dOlaubsuhHGQn60V
TX9IMCfk+F4B9x0HrspN49NIegtCyVMye2EwJmSP8NFlNuj+ZL+u0TXOcxqp
Rkx+oQYGwzDoG6qkxOYJ4xYh3moF3YRfPGVcSkVklUjIJgRA3YJGUq5A+jj7
2u+RkEhAFHDJfKPFDYDZl5wtqts/nyW0IagTXHoV3TrnqESgkf8vuUCfFNOe
dHVa2oXBsn7Wqkmf6WAWxacsY84Xs/fqfkBPLErQ7yAs/uU2iX+CasexOov1
Kp73TUM9TgWS6DqA/v9Pu28uL1cQpH/b1yFTRA0bVWZy3f965RFQJZ0yE0gB
fDbIpvSt/XQEfooXUApSawrddw0afiQLf99rcU3HTMS3nDQ1Tei2SduZRZNL
LM645qWStx8zl0jHWQzLusN8Pa3tNfl9pU0PVsftXw9q9adTfvnotZKq6Pow
F+xmo99uJRRpvUwzh0K50xkEJy7PmLXSyoWFRfIbu6K3nNgJ3KfnTJXiWigG
RbR8Hvp8YhCEPErGTXKaR4snLqesFeftZ4gEJctmO3BXOuJth2iOEGTiK7gA
WfTJA5qmHuPzvk5AGhu/gPJtoX6bpI9OF3l1DogtGouZrFBPPGWnc0Jfy2Ym
ZjPkNIGWbVemvVzpoxWqU0+VfQbXoki3CvOC6zDH7ZJJJThyYkbrbyhnzmWD
KFom4aN66GXiTOmoqX0dBaNse5/g9cbFNopJ1nkTB5V81V0TAnAZn8LOg9oe
nTM/ckIgLWlHx54d+IaLiYywjj9rDby0Bbg+lfSSlYILFA4A8twe3jTlV3bY
PCLOQkMRRbhQCiJRYsoM4JDEPpol/+YbgnKw4jmc47GSTaqsq0/l3HUwdFGw
Xn7qhqvo3qRYqv5q6A4P10glzHvCCc18dQPwZ4t5o8k7M7w7bmTrfnjMCVSa
lUa+PhmwY2zTcYAP+5+QqXUaw/hj+vN913w4pnlbz28XMP+sYBQhuX5qmVCr
eN4mYZfv6vzaQJonhTFqoqcIEt+Tj6E6L+QJa5bEGmnzZSo4sy3VkFNGX2mB
5nxzHH5fTxa09z2YfMfCwYk5xpeW8G9HuEB7q+YigZa/dlEjO+MHQ77Ds8In
Q5QRWaZTeRyYIoxAT9/XdI1bRDQ++R0M112BGw1XwTjC3lWqEbdqSKU3eu/y
R7yDg/NTalFud4GETmWJXgqd8fqAl+Qwb4t1nwIDGLoXX4fYwbk2EWa4eWPr
TZTBYcwAnwL2MbfLbFzbx5x2Mlr/U3mxjUUHAo2JYDZr1k3Bw0tugiK4W92V
efOgpAp0KvzfTtaXjybxUyE7rBzdV/XEEP7/dhFGepapk0ToRiNT7X9OH1Qa
PLTetuPzYsIZwPc8ZgrIj2s9DZK0Fw+iKEUTdBxzIfC4KcwBeoBncHige4bk
2bELw2dK6cYBnmoYB8TQgvnfmJLs4TvV0b210TNu7mu4Gg40lNkkLZZZ8DJc
DY2NsoRky88uoj+cTyB3JaLjHZnNZ28OCrir0BRWtDKlMuaWspvsCYLIHK9O
IsFaO7W5/t+tDE8FgcCCHC7p3VZwn44I7FGTj+opMW+LRZ9gzh6cbP5lTi4V
GlbkwIIp6pMseyuDc2Jw4HxDLSpmjjxyK94wsLirB5z39bZzPUUghuC2OXr6
2H/9wBqvvrz1WCM5y8tr8p98Cm2ALsKz32zELaeH6qwYVntQQJuii2HBsgqt
LjQNEu/gC0RsWNROvAbFKp81rYFzwZFmR7yPKXjo0dJBzb6x7ZzWKrBUCIBJ
p4/dJVGV1mW+Le4+DMAwv0GK5vANfWJR92IVrH81+TEMewLx3W/uilxfpLj+
wVlVPp+OiPBm+zwRT6GgRyqgRMJFbESR76a9M4V7MRoHX13/YjUgwFHPOUnU
IBTU9EbzqbM0XKTLMZ4KEBgxLhZT43JZlkrdkcXDHVr2Kyu1Z8WtY/2mQ69R
GsG9GD0oeqxwlHJKR2wJpQrJ5gb5hByZKxXnRqKGJWgxDzOPDmFYf5yU/FtG
LIscB715UCjpiCkK3BRzlifimAuws7s2CSICDqXQHul8iGWRPcpw6Tj17gNl
3up1kHF82jqsBAy8lLpAgPUIYBh16IQi+DVKF1h10DQD53eb5WpK3pAU2xIB
vOuDQjhenkuV6MfoCZjyUPN2u92jPWpp2/YRl6K5hZ/j2i1USy2URkjqW3Iq
TBe6zGYD59lFUI42kMiqLoI0Nf9T2L50ETxpdg+RYViApSz9Bwmn4PIQdsnr
FVE7v/ajmZx9+fkl1wC4g9xRMQ5LeE1JtCncasKJSUyF3/0MnvLXvrMNibWd
FICTvW7DjD98VRStpaD5ud9RSZuM3So9qSx5jHQLng2eAz8oKt2b+14kGnIq
lJJjJMPx9jBhf/4XmhCmZwUUEwNCQ/YgE0yAHF77Iec0jJSOCGf/Ffv0mG4H
8dAxnQ2qJO2exbZbGVl7HPVOb1gOW/fxzcur0zs+nnA7Fqlbfs2VnO//h1+H
CBxO8p8k49TCPpytAxTkDzR8EK/I/sAi75e1v+25Ml/aePkkO1QBr6qrojRI
7kSvQyRKLQJGCCXHKwbIE2kq1BmtnPDkFT/PeLRh08ax9FFp08scCdHc6IT7
LNalIz2N3OA/zqbJ7E+26qxXCCQj++VgZKxzD0Vt66kJg2VGBxxjRsvnAqw1
91/TPQiG8R0VbmOU1QTLxHkdBz+RYCeBpQs1MYBez0sHveSZijfOV4I+Mby8
d/IgX1kgL1dekbKrLUxbIzAoGJ8M5kiKkflItgelxAXN8U0QWxXWFtrJJGx0
x7z0O3yAGQfc555d/oJDo5CGfsH2dAwl1o6013VOpFxcDfRGZKyvT31frfGt
UolsVAXiXgecXo4/wOc92k1ANnlRZPYb3SjmgjpJW9pndaYo/RqtuClOY8iI
4FBBWbhGMGWv8zZCtF5FFZgLB3C2l8zBe+qCziirAdsCGpT3LjZM+5LBCesB
cd2yUXw7t+uJiUsd2ROEVNIYckFXaa9ETkROvKN/zA1eTBURffjF2GBc9QIT
iaU/MdO2r0jI9DNuwLzy23bf46Cy8OBtpsRimxGcFkUT4dkWcbH2bCjUNs1e
7QfR3O92X+0m21Pk+Ks59WQ/+vhj4vsq3OL9/SrxU0IYw0MDK8a89OJyET9Y
/F8mUtzvoBksp7pX8ypVi17ErWDignfO3un12P8el1H4sI6ZLE4beD98MHyS
BCC8+JnQRX9jC/9ro1QZpI+eR8tlX0GlAWJ8JS6VE2d/iKXM93fSaU6N+jUO
c1o82P3uGlFqE6VQdlHOezlexoX2cpBiDugOxp5B7cwUAp/mS1c+Q9Oj7q2B
HPCBOUeQ63Duyygd/hZPZruxJUCXMWGy9SsJGlYvTT5rIFxabVhs/fh6WutW
ab3qAuJC4c45KXPPEZ44+Smn4LRe+4EjSYRW1Sibl88aKiMQ8tx0e3gygwGL
7tXAqbpLFwA+IwKKAAFGkv/s3FqokgeZS+ZNr/r5SasSxMrXP83+TFL0xZFq
NzIcWn9YUjaMT3lyTZkC3zOghER94w2ikF5NANkBcQ7bvHu6bzwh7m7NcCmt
kWAivvyRdIBDdzyjWEWmDe2RM+79fK2SAebO6dOEidJk3fciqgkwfWNWUeHW
3PIc3rYKK2IhyGEV1yMvEdNATX1pQTVc9e+jzdkq0CpDyJfxmSkRqta3NWDS
xBpIYDSEwaxAYdohUnHfYujwmQGe4yoClHCyqdWyITWepkWpVohq9Uv1H0jD
GhAGX8AbwBdzGDCmKD4LgOhVtc4Hs2vwYXIGvY/Ev3RA+4Lj5ELtp7NJhDBY
WxjtWomkHkQwH7Ayejrmc8YvVaPUK9fxBjLfGVMBPXv22SYNg/6dp43lhZBi
AIbxjuhCJB/B7lcW2TIMcLu5k70l8cd3B2YLcSuByGzAlspRR+vdPi2KAKQ3
Mjodl6ztZg5w62KXzoM4WmgBbtq6Axx3V+b0JBfcPHKIWCD2SahS3hqtwe1+
doMmfftSnVTs4Yuvi095A9JtMgsXtAP5HbV5eXic1HXjvxZ+uL8iMojUkZbD
N6ATk6w5Kmxizj17qbfoDTA1pQ3kmMD0iAHLuEe7p2IqsKsly/K8qWRqozQN
lAxi+fBmNZLLn9oYI4yqaVf63Tcoiz7nmwGF8dCH+O/39Ao3Ndtd3G9yp9jg
WBBSTZnI7oPmRXqXj3avZQQOVUsJG4TF/OhDLN7bbuKjV4Sm3nq51bBnG4Zl
iIi7NlGGc8ue/30WMgTMjaItUBHSHvOf0epjYCNXCAx7VYpELv1aPHkDNfOE
ob/rRgDdRSR2cR051ikXkB41XlkZP1W55pfWD+ubQSyKRBYIlKjW25N9BY8I
BL9iw25lvcZx0UKxVKm5Ur2jaUwVW8n0uLX6vPeQKe8XzoJbmmBjDSd8KX3u
bfltKhC8/o3LTZq4Hw5T3iWaeaVYk8LWaoO9yez0voyLeyMIYkO7/i7XnIxA
eRXXv/Er5PS/zEZTT1OHKKo4LkdNpNg2NF4KyM/7w3NZ+V9Ycao6DuIqO14o
0P0cYBXeYCRR+SGjyujbbnGiR0Vg52b1Q0h7TIHJ3LymZfopQbszeHGs2fEg
24cpqPskoMURDQ5Q5D7Vb0jyAKjhMMNQRVXmNeC4GeD+mV+zE6hMjeUJ2Aun
giX4s3KQTxHyhX141GCTxL3CcPZOnJef4VPh6HEKpiy22mO/39f/RaNIChAZ
EbR4xeURqgj4n/YOs1uLXVphSozZzyfqzsbaBVeZzILJW2ir5C+5QjBzoziB
mw5pzFhai+VFnQKFYLgnDhn6Gl4WABaerx5jEJBIufKvALzY1mot9+FEMBTL
q6Rriz9g8m7ntuqGd77Z/RaMNp5Ywj05qRYkYKCk48QZoOd2/hHs6gT/Z62o
BzgXX+PNtYjuDiXT25gWlyC4tvSV/sY62t/cU7uc/KB4BW3eRn7zn0S0fGyV
rrUr+m64Kh0/CYjx7dpi6kFf8whd7UyVdlCsXzHmVT0qvRma9WFkECo8w6qj
KXYhTeJjlF7Wh0k9knR93Voo7XoGznLQ62QKWaTidUwVhd9oI0BVpSIdkQCi
soHlzf/kNoFtjLayDMmsrWFO5wS1g/3v27ge3wlp4tAC8UlKRbvoqC1d7tbP
JjTeTx6BAW0jYmmGsvaw9UEio+CRmfTZhmuyANQgE4wK3skzBXm0nrdfUYb+
PavvcE7ylbzuxZxAN1o6UhHS5CRiNhv6qouCVuis3fGkVUVUaPhxPbWjz0y6
aIQo8b8SmaMwf3pPCQwO8wm+hjPWFNsV1oEjLF08dkvIvyxTu+UTbjoAONt5
YKODD+9eaArbqcIlP239QLesS6rwJHbepyjMflX2UjWvV1MduuAAOAj1GEG3
37lPSEajFtxeoWsAXTT9wyI9ZkSz7K5R8iQfzvz7H/gE22lsA8WMycO+OTZ1
GkjOiTF+RQKs1RzFXnJGQFfkjgs7CoJ11TVeTRabcdVwNbnYFCQ76XJSCIjt
1EYEqFnhuX53qIi6KhDZgK+WtjSo6XYA/oZfB8/hb28cgve+8t/eCSGFRtfg
gnqQoQ/c7hMDOOmy5NXFqx1hRhMteE6PPRjKvRhC2k4RP1SGQI6Vqj0uIJz+
7u+AsTX/HZOKpyuqDqY27RITTCYIjRX4FdfSaSPwA0ub4eZnTWdMRYbePmU0
KkXnMMgngDZ/yfLowr9s4qMWxctANJYKCWs9XFVIDsF871B/kfxyl30UHjIZ
TElVsIMwvMxgAOrMPiKsIDOJpUke97Dfq2YKXiDRyvY1GCr7ZtjJbL8bWpOY
UABvfC4EFat85LqFZe5YNZCz55x7MxGTDUCpP8uifsAtlMP8Zk1CT526mizO
VGbYd/T4Tnjuhk5oJhaFgO3jMMFStr/jjvz7aicGG++FJbVnBpod1ibTKQYv
uSjBtcDY0cAge5IAbCVmDdHw89ZBTsW1/n79Ql5qpGdkBFaqqc4sQhZfSmkC
IZjEMV7orEBNEi84FrsG9oEGTLQ2eBerJi7kgLQpmGwPZ8+fK25QecEkfOJS
YeR25qBCy8PRI9V9ms7/4+vroNqwNRq+SiAZIQNckvVh218DlnNWuz62ASsK
tizK1VySFyQ2iXEjlnXIzlcXVnFfmDtmYdKo5GHdyVEFq0ezcaUyyKAeUtO0
WpvtUp90QwLXTqBN7UaX1b5b/q1co82oQcoZCphgA5SYeY8m454Yt+ZcMuBt
ZQmiy5OP4iykJdYSLLIykM/z9B0GQp9grXb7mW2Nsvd4xxcyu4LW41U1Z/BH
c1TwDLjJZ86UpA/RzNhRryNjiG4SVKpO+RVCkU0Dai8fub2xpPMLkTRFyo24
R5R6sKlvFnnn7ORrkOMpvjOwerVP/GejANg55p5+tqhwjnI2tWUmp9r4UkD3
6Q3w6rRhQqrToeeFEV+ZAoND3pEjAxnyjsXOoBdhbTe/gAFBbUIMXZ38c64s
KMdF/IGYyUn4rI3lEtJ1M/n/67+J5qae3YUHr+Fh1ioPTRto61VOnnrTATCT
QWJT3C639HuEtvPV55mEbQLBdYS+wPUYveIb+5K/ci6Rv7M0dYKKSfKUvQBu
Gvs2JVmKqeCejOPa6lYi8e2PHb1LgEl+gLeEpY6RoTQ6uRE656xCwl+Yksas
3o75/s7Dhl55BUcQRpKyGGQCdlkjGD5d4gGxifaUydfiPYcFZ3XnFy/HVqsE
/sbsMnXENcoUHGp98J4/5/O72OdyFjDK0LBFVQzKNkeGFicFMZUfmpOp3YhP
mboos6EBAwXVtQ9UnVbBwTf4Q4+DhaigPK0DQD/IE9LnS5BKTL1GffncXUFy
4jYuVeNUbXjDC7GGX5T2l5bm7dukVxnSx6hzACC5nRBwJoTwwnRB5/jrGicd
vKkr3XUu+aIpWGhmu6fk6bXXolemjdtzmljjaB2LyI8wBono7qIOwzc8KSPp
oEQ9yGZzIfskSZzvUVudgwsMYYJ/LHtkpEl/EceIxkzv87ULs3rjTBRfRips
RQh77II2kejUZzMefejzV5f8qLYN5h3e9d2iNTZ7752S6+zQ6mC5FCn1UhQm
AMO8b7LD0w3MB3ONK8ly+CvZY8Fn/temrXuWTc/7+sPP8fpcQphRinsIFzI/
hqf+68MctSD+f2xynVdOrBSqHYgUJLV+na0lTKR965BKHOrdFJTf6ajQpL2m
CThZ4MZWEMo1Nh6qNqlxPKqwJHRgpHHZXz0VrfjA8DD79JNiU/theOzyrnZO
2Vb4AHbTbVn6ByD/n16EVnuoCZYBJdaSQsSLYhKPWy3OWIa9kYvv5nmOZt23
EKwei1DF1DSLlDAfZ/ExWF8F3J/yGQ5lqIm+uLdVyw1KAn4+T/D6vN8WwCRW
eD7mVR4OpikaVbbPQkK0akAD8YCtT4kHTA9sqzkkzBO3Qb86QCtXn/fKoEdl
pvMhiJB/WBcGjwjId9I1PhHXBLfoSJUPpjVAKUpwmXS4JgOry+1XQ78Rht5o
7rcb5j5c3wc/CFrqr/JIJ/23S9Ng/g7kaPpZPXX9Jyl1oBIk81v5qqRI+KBp
wMrN9UjRMZb01xDune2096bUmXL9ZdePGUaMjkMPltZyZQ1HMy9yeAgNXxnr
VqatEznNNwnojtOC5CHMy26WNcG6uSJgqibKbzb+n/dtC82DV+7SDzMe7zKY
atzxWSHOPJxkcN3ffivEo283xpz5m1Co7OzHxbzG+THm1vC0kXxqruUR58HR
XPRX6urWTGWy0q5uMb3eeCgYrKwpWXrluIg8FfjpI7PH7yxV5Gb5nFY7nnP3
fBszsVwhaLdVhQ9V06JMd0NUQdtMzpHVvwqFPA0j5FsSMHYuJPkbSwTzMHkp
f3e2I8pX0yvUaqc16g2R0Deys4RkzydDfDuprmd8fDOOgkVSzbb5CEcoNPD2
tWY6HiH3ziqKckg7VppgecYN4+kx9pAo1pxUJYQCq5XdPTnOmzL9+hwIUZsc
aOHIWkvPYO97Jl8JlyCmumzVj+wVoqlTljQcK3wj+6FzAIkPcPV8UFLHNwgj
DS2Pi1CrVdFPD7JYvKvoaLXiFru+ETUZ6u7CPUvi7OTi03USuvAnEk8jWsI5
aKpn5MsnE4ChE2C+Ao45MO7rZnkivQv40xIxGMc1R1ey+remDIwfQAaBnNyO
waOqZTpddKP93/WvlRUZz67FGUmgRzbWlGuZ2puIqYR8aYcczqjWbzpEllb/
PMc0VG1GiSryjROopRn0UnUnaZWJgO57q+RYEclFEHAZMpByo1xXzubF7Fqp
QHxAoVijrZuucrOeO1qg12e7wONSiX6p2u+/Z9ABMnEFzuAKHUAVizX+I4f7
2YTTsd9K2zCIj9HxHUvlAPZjnUA2NGKUIO99MMu1fexQcsoGLInfrBHsNV/T
O4uQrFVX/kfWZoYb5uXE8fi7eoWC+hZ8yKYA3dGGJhr8kva2d0aODsFwpzEn
DxfCZ4BjMUjHhMIhxobWjYUzzrLrWmQBLrb1vCbdhZoCnGhb4pC4oR3uZmwv
dvQ6X+p+OdkkU7C/HzAu4CogepPnxEGcrHYCg68BrF3YF9UlHnUCjk/6wUXs
BiiNW0RTAzpqo98CxSSFmuK+GjOnC40GveavExjwJrQdOPSrNMsUykeS7aCy
bNWxgodHa94rejyzlo+SF7L8UtSZqlwOPmw1DOKec4GTK/9quD67LJxK30p+
xqZOiqaOwUz6UNMB1VjKvfayGyd3RNjIVl5KnwjlKgLTzR77xwFvyeDEyBTA
rGweca98JKEnre5qaqdct99GAAj8Ob4XT/m8f0lCnLZvTevQ0BFGf0hGe3Vc
QpVgCTfzmL1kfHv+JRMn6re3hwV7Mjkup46yYg718qF1UboNrc5vZrSqWtz/
vZsCMHdMjyP+ezPVDDt7hUAbC0dVs1AZodlQfW6SGzrsx/z7BIJe6+E7mvyP
wllfV6FjUfGBVI85yDVWFJtK6Jx32/pASdi3m9rQNQ6x+Dlj0LZpOQuaJXAi
ESBBXIf7UCJfgzQirpTquw5i5HwfF+MJkeRKBxxuzfpgzv1tpcRlo7C6MtWs
ezSe1q7TZfCYEcHcgvWU6DVNSn8bNSJUItFLOhX11PCiql/6eGqt+kE9SELx
MckSxksKEOr1l+LXGM+cHoqt8NrgusDfyqDwp0bIQk17qvL23fK2HHw2yZI0
YRmnNss13K1KRmOp2KVEix4hn1fZG5DavGIMYRl+21/IGquejp/fYTqaZgFd
Fa4NyNXwSm2kcxiNcHqZQvPrSFehVTIr/g5iZ5QJR4OmQzr0t7vW/EsRxrkQ
dR5ST9TZ1sFpTgeWVxqqpn7+cx48me7IIIiDWhav5oqB/7BhJIFAmOj7/6W2
oGxh1XJqNEboqUTTLrNXrfesK3VWN0v1pLpXwfb6Jv4VcDwwiCk29aGZl10O
yHV8ttifXbTe3cdCTi2S2aMep0lvcYX49JmiQ0J6Z/0rDqsYQt+NMvQEk0Rh
5AWUb2FOFpv0pnjxDSEVsQr3ilMjsgmuZDZmHkSf2dN64M5Drp+F90Zayd/q
ESwNNkJAtD7btAfLyomC1X+y666w+s5NcD+F2kiBL8ZuM4wQXfTwI77i+gEl
xzjBnEW/Yi6J0+xxKHr8tM6nn5vVxHCNQ1jLrEn+sHQI7KAx64LCr7qlDL4U
u5mJR5zWhRJaYC9zcZPuJh3slFx1biv0cRcck3MerYiHOJ6kAqvbUOrGFF59
7mCJYpMH8dAYwQhEl4BTYubES4mGDWropk8sPU27JIlo/dAMEYMCu7qRKMgD
AcYS/7/MqhZzmMJ757MNtJURKpnfnG1AvTdMWoxoS7gAu1I2EFQktKki09AF
TyPpTs4KQCqeARkJBUMyIiWrf105L4BCTOQhkJUR+eHjyd4THbae2dIsO9WU
B8h/6+ll90HwtgsqEYqakgIAXE7OnVlibP1aAgLOw/A7CygjHVsa9yhfhkC/
d85CTIXpmqHLHH+31bsd8YReRqVgZb/dgdZ7eJzBTye6r5+UUIebjWFyfJWu
AjDmGH8ua/tCnNEn22+0HCeJ6soUpJMwmPPpj5Sbq9WSZoykjyxpEcRGh83Y
EKcndC6Hoel3xu2IkH1pd3SBOpqE0R3i4OCRTCz/kJ0/nsQjanchivPjvziT
LTXlNDNTgoG2YsuSYfDwXgnny27Ibnefm0OSMriJO9b4QTw+TnWsElz07wXx
NJxBto9lejsreqTQ2/EaBiOUxnQFaZGd/EV+NrSXoraopJmMkGcRrxyLyUvu
U+Yt/ckzTVPESg0aIfKiIBgEUTxLdFw8jlArRt/AfUYOhJq7Cep62X2/7XT/
Vvf+kziI1NYolNTEgRv+C2QOTXvNvFmpzng+P+Sd4LwUMnTK/UqJm7wJC68n
CJx9AjHM6lEP5/m2TVJabC4Bv5A0lzx9Rdcvfko9vf51X+QhCPJ4ghEfK/I4
ym/X8en7uuRsvlu6L1CMMDIZb7C+RlapyDHVKgigzUJkSbI+iVCvLDz5Mljj
+IWinG3EIMX8E2Jl3fQPNSAa6LzkrlGMKhIRrcqPDMEtDnvdDjHjUZoJKUSX
RE46/60Cc1EN7bYoD1zA1dIEMSUnJUH4HtzWY341IHy/WJmfdCPiBs5kTAn8
nLlipoByovFBbtjgdKtFjJOTn//3abXnS37PPcoh7JHsoKVv+HpMw+O+VOIZ
OTS74IW2ku1+P7vG4JV8M8PY1+eWxljko9HkeXQGPWMfz92SyZqWcJTGQwTB
+3UiaXwHqF4qgqncOra+eQrOBHbSMCodI1h8T19soDq1Kh4IvsKqQWqzGkGY
YtodVPWuuQdv46gYKOwT27SLixYj22kmerOmOxcQpqPm3eES8zBVBHFQjVwV
CP/hM5TE6VLsHbkts/129UGd2YriEzc4c4FWv3VWRC5eHW/omcspG7e1rMta
R9wmrNWbJMpRxxRYsV1sBAx8l4+sTVlQ30BsbxTkBa5hXjXTRpiBE1v2QFXm
S2QTqgdfHfk1wAOy6YBCxchldKFVMYpp7ciSt6/q6/KeQEuoOSo55xImnNJx
fJabxwL34QoFoY5qcMzOvB82ERgOyUEGvjRPWRhXzuog1cZpR5RV4LxWeeSq
U8uWrqGQ8ZflzUb7dzFtwSc9PZxZqLM6bQ9Yb5r0Y/57L/E2iVf46uVoyI8b
tvRZV8VPVFf77TtFkPF9lMvtDMqbQ5i5aGjfltjCt7KarZv6QtzSu9eE/VNw
YOnSAVxFiWLH//n6pcff6lcdIDfUCKmB/lY2tmtoJ7pqMdzGf/zs0B3gClWO
KxEI3kizgDX2Ma36Znfm6N6Yq0aCXVXrNoysKZ/ZnVDr5a2/dxQQ1BCluFDA
I+PB3L2UVgX4Hh3pDx5Mqc8aHQh6Pu/qbSmGtvrVwO5mwsW454GgJyPKQOi/
K6r+Pl8TXEr0GTn2ozyX3CpXNtJ+cDGRk7owZ+fMgw5ERD4Tk5n0od5h7bx5
pVvL1A3MWPudJlkiADqdx4MuFiyU6ITSvwjCWiUr+2YJmahaahhIZkjDn0Ki
1XMKO5raXeLLYXy0OmgsXZRTAQpoVhRCIjoMBsPb33xh5Ahqo4fOXX6U4ow+
0rlDTBzfe9ptYbXhWpoaJJMwya+VgI2Dgb7n7fVxvATVL5MSFhpkj2/cYuwk
xoFIsOCNzT6U1lHG9fEco0H7ufFnNBNI4y+dS/OwY4OYPah0dj4Jo6ETvb1j
282WSTnlcc5V/gEMMQO2sZy5LElpC+K6Cv6Aw3vaRZlsmc3Lbv/S9zMQ/T/F
Ov/v8GZ7mCiNL+Z/kprkS9nyTP/TXWpg2vSD8Vcft7eouSroiAKEXsJm8ixk
BoqQTKn2iiXscuu2rGhnOrqlVxQqP5d1nbMbFKnx+uiUYKaOcNUSiQ2KApJW
auOqvvVzkZn0kcVvDr7KN+GfeoZTKDC/gs4ev7ugqJcN8/bCyKhI+MaOCy8c
LOTVKdSEH4mcB0xD1MuZz4V7HkDfr2OkU7062jJrITSeiRTNiCGb5GUow/JT
I03tTeSj7tw+/BU7XSEAK5m67NGavEsNDXKPo4xdAvrwbIS5YsxcfxhRWljJ
igbKCpuyAvUUzbR2TAr6g6AeGqhBv+5zIInup+vjRpn9QV8DNaDPJhS8NHza
W89LpAt1yRohQ0T8x8pdcskBbVdP3sBJkfcW8hc1nRSzyvKE+qUme1MTlkGN
tkpU0hCwgedyt3AQu4XtQRiw15rKYzu8V2YH/S9WULUVoDJlcQV7xoLwr9se
fM2xE20gRB2tXXKTwm6sJqvOa23Ps7SrVQ0+iTHawvM2Gp0oJjkiDCS41Mie
BUyXe2xNcIo9nefjxUGyKdJjaxbVs76NGWWJ5g2rxZqNoOOgJGt2y3F2LZ2/
Yi8pn2VLmiExkMDa7Q9bHBoexhR8LYsniLzjXlpyZwKRSs2LApQyCY5n+lfb
lGXtMrhWPOE38uKVYRCpOiLMluV3PZcha49qa+R1ilsIP8ziv/MrFAw5yBY0
DaMGqIGBnYSNQspYDTt5j2ph8tYX1eq4Xr8/sh4W5ZNxdYJNGnBUTQfamnfg
XILt1xsFzqV28G/21EzttMwFC1nL83b4lXQKMuY3Wlfdyh9STEvZs4bHhex8
JqCFS8ECMgWfhuVnQhF9f1p7u/yuNy+SnleUq0NuCYTrmm4+OrPI4W/6ddwR
HFck15FOcOTGFGhED3CG0p82idDlS+c8V50iP6buTb5uFHAa2Mx5QZx0aNLU
P+SbCtvyV+y2YFr1WX/Y44dVvqf9DL8YI5Zf7gfO/GC3/SEid3olimDblNTY
s+v8R95s4XmdWY5Qd2MnGSi43xqyMSqIPIHgcNBbE2xLQSQU/mgrkdCiOLfu
lapUGrmlTxtIzqBgTQM7a6N2+F0vFnB1fD/7yCaYzg/7aS5yEGP7Ld9jrwM8
wcwlrpArIA4jK71V4od4yQ5Hsp62ag+aXO0jzVqjuZsIESQQgkzgmTpn4CPN
MZ2MlX+aDHWufz/l12zAIfw81ynvkKDQ8pv0x8qTE5dgGToGwuZMihJSZkrX
/25c81uKN+JLWNbLl9EIVcu83kVtWgJjsiVbcfaZpKFmP2MHpmGb201jVL/x
v2cWNRAf9vMXpDvofl3H0Myu5ZUBNEKZs0MJy3hN45VRaCwgQp4FbulCYCPO
AFRDFESnfxP7QIdmrIxxAzmGDWoSYvN1fDZxde9YApWHZGmiV9UcvZLwoMxN
5aTubKvab13meNkiihc4nunSOFlM2GYTgF5OhZnFPNBUyR6TEodQX5SBc6Mx
mN2Ou62jgn12lmkp0vG19oiYfgCvUaR1ZDGy/O9iSKB4ShRfL5soNc/KeSUU
SGuO1MyUBcNA1vs9fJowFdfHcw97jDio6amSRZeMjqS7bTl2OCgQptX3jZrx
gol802ybKEkKKGQojMJKwW4SU3Dd+I6nHbqKMdI0dOwmF8r4UFITg3fW6rwp
kflQJf/5AFmaCRqr5aOlym+6hzqnn4JM3nhQoniXjcwMdpuFqOSPgvcxFZ8h
6jcRrbFXG27rdSkG/lGPC01YX2bsCd9wRKhGu0UeHXfUrnCctN/iKnkZ76pi
dw+t6aWie8PIJWom5+US31KrelZyeVh0SpR6TuwMQ85UvJlN/XGXZtvsz1mi
uPdXhsL3Z3Ie7RDdx0M7RqF7JvGmT/lAaqyd6X9erN4t1CkLo3CBKBiS9Gon
dZihe+elgumMrsD+xx9pc0DxYphhhhXRMc/gVFUHVjSqoi+Gn7ZtAUe4wng8
AZzBGyVvNHOmJveyoLSXPcehBWKB5yTjPvLyiUa88luUkTS31YyD/8+sJaIM
qlj47lE4BpMRng0zwKyOzfyVU1v38ZOVReHrVJG8O8tZUobsEkg8IG/0yhXJ
6anGJglxK9TsM+xVyaD0h5GG9XcQWL0EbevztN7wzW8o+wUuyFT1sDWfad/O
9GSyIZxkmP2xUCAULVM24sas7cRxo9BekZXgOSl7vw3URPts5a2E6gxc+Ah/
+1pfQnNjeTekRG22H/aY5+iYV7ocRaRnW2YbvRB3GcqfNXXkEUAq2WJQlime
Z5eiU1bB3y72iwQ4jo/suAtRqaEdzda8g0IoN602Cbm0RDHjbhnVzBYq+1xa
z5sEEbMCe/kkTloGWezYFS0d6WpwZ6pJ8V5504UgLEHrZ0n66/oHN3DQExVk
dsS6pbxc/Z2TZiRcuN9xrWvF/iGA47z5VniGnjisWfSR1EB0Kt4Jon2Q7Y/B
9SNNtqzcD0m7jXAiY8l0LTDB7cTwXjT3Ex3T38RP7uiQ4dsLN4AjhQWts7Ae
NE0Sda5tCCUa+3vvM+Wq/rWIcbWkJVeobw6j5GyZzPUUu1LVUU9kPKuoFXVK
x3qWSQEMGNTev7u2VItvdBDB2CwBevLSJK46JdKpajsFcUh5PbkJCH3BwxBc
Fg6d5xKwNn0W25I3p8SpblL7Y+dZcXKZ3LnRkfqS0YarbjcHseToVBbtTBhy
CgFDzmLIBCPalBT6gXJdA1OMNhBVWc9SJFKSsHa9WBrWAWUimwotoe3lTMZh
Z10d+jBRYog35Bzqjvo3mluMdLDzzCjR3UoSXgRVrvT4Z3RthIYoHvMv3+nx
flKScHLwoQZvzZukPrLdtsD4hoMCJgyd59ohrsKRsbPnrJiTJJOtZHXqiTV7
4P72F6zFkmgAPXWzWycMR74our+YEZiljHE9J61Pdty1xhNyBlVplNKAAp6m
OS4jqk5zXCXQKNLaiFa2cptzg/M2plBgv54O3K34czddlNGpVc+tVC9MwC72
W5lsmZgGY9ZbZSr3FVAM40rzqM3dzEPC1QMlTXat37V/NKV4Em/Crzot/AZy
pX0JmrgJDJOzKKSPfD5JacPQrNqBEwBsyCkVVod1oI044xKixV0xkB/ny6IN
eM3M2QoBFfHXd+8d8QuNO1LtbOydXrKas4IXy4ZswRb620rlipGwQIp96mg9
lNdHAtrAQ54PBmoJ+RXXUqRbAV38yBLaQC6AhhLLXz11TGUnoAF5s4y9S0pU
PMz6m4zsarzr0ExG/AptjsWBXMFI4Ja75Lb0Q7t5JsteH3cKZBPOqvnCO4nY
z2PxT1J1LFVIOdry8f5rR7NTldh9z+GRAZzQk12RQRvwb/0kq9KDXeHRjaTs
VPMBZZPzQfHIHxu5D/NeUVtzaukpCFW+bBePGgHG4GTUfjHTRmAVokVzAnFs
+LfQEPhBSD/USyxS/5A1TeMxAo8UAHWBRABP+lQhLs29utF/gD/LkSK96T3z
Qtwpme0WP2WtjtDuv91eKl4Thi/P8uoENfslj1zWG9HNZrPPqfB1MWJgsA+c
TxBeVPepW1JiBEJHowMH76AY0tAyOSrUx36oSPuHbpoZsMM+DKDzbxl3n7Al
qocDELLiaYzWG7x/GDEF3KpieePyKdqZkrJ1Y/+/p3oFCjiIsaKQMHj+DjfJ
qsucUUulAUBzlYbBFHht7imxtjSQOt0IVH0q7wtN7npmcjF3OAVcO/jVll+r
rlN5AbMXP6spAIz/2xY1zGIDmH3MxQcI/1BCKsKoqWh9/IbIYOaHz8cZ6s6F
YCgmEqgcpGpY9dMf2np51mvppgA70cQVuYyj48s5bDkLJ9ZWn13twt3MEFI9
qN02935h/3M+zbT07t6EpQRlPnrMJWX2QtASmiKfmTiimrFh7R5GhZtSkE6M
q1fvb483xMuThKKlFtGc1p5MrCAQ727tqjto+gU6I0vJWtm8s9I6BYI4nhUh
vJXZ9fHYDOTzu46Xtv/V5prLpKgwD1CYKmQSGNxiLRjzDMd5vxHxN6rIn3Jl
h32jy5ZKYKHQyzytBw/6hx6wtGIp1oHwi4NtIHVDzS29XOD6FcOrmYLqL1nj
7YRI16UD3G4LUsctIL6FLmfwiwFYNtqPreYzESKvT7k+6I7N4pWA7OqmXArQ
FKX8BtjEFqrTrEW04xgqP3TlGYm+fU7bowCTBBKEHWSV90rUk5FDvQoY2vRG
GGDgB4eOLhhbjFQGOSxjSaalNn9y8yL7bw8gyHp+DiBWeMSWObGCN786lStq
SsIq+SjVmC4uu7VL6gBStuSDKFmIZ3rKg+zvHoz8joIKZ0oCSy5kAwhf9qjv
TbXz5uwatElfYxqE2MvKRKg2c/Y4HMlC9m+0voxzMK52AyXLBj3PEZhOBcVN
aTZIEhjSBpW/+buJORnsiGcIZA9obTzSONgG3QkUEZMVrblNbHYJKcYapR7K
x5SZcLzab8cyePjt067ygCyHWIxBFhxqGeXPphT7iqM/hGAspG7saqEsCxiP
Z/hwxsZhoUBcNUsUcbRPWkRZgZMgA40XwsRBbT5GliVoVf1gN0QNO2G2K3J7
HNaVbyqHeyHwEcWWaLjtKoZqWTMB/Zbd+z0rzFeyEo5AJzuDshFURl8K4Y0o
nYR/JbEqpwuxw413HNYkEGQzHIAKv24cNWHpk6/uTFKg6obkWNpH5IpYcaQY
Aq23Q2N/HrTwTaMgP/QoqdV2LiRl/sMEKlPYS/uELdb5a11gSapSmJ4PVRoB
7JHiALZ96t3ANfiWKJPEXVI5GdUiAyUBuiENBkBf1qCscnxypGkYyh0/JtpO
HHEqqfQZlkOoHAjQSqxQ8ZK4699FgwTxkztVVnyY8jb0Yrt0PwWLfKUvnVVC
g4GNlBF9ChMP+PDL4Bh1ORbPhCg5XNDys3bIiSmPCU/its+BaFSWXptKYQqr
QO+5fTX4MHHuxhLEVd3757zx1vxAIN/I7Zl8lePwlAhbW2/sTejE87zQqfel
FNqww2P21iCoc9HPZpj0FvowklxCuaKjfAcHkqBG40Ltpol2zRWx+H0Fw+kX
oOa81Drznou7V0ZucnQZ2B1J4vLW9M6uBRjLxZsCg3YB1sOt/ff62jq3tSzU
tt3TMoGk8GYwJtdA8xvLQSxNLpx2vISeX+Sx7ElX0L0Oi4ZD5sSE1rfvYjL8
FntjrhxvjRElx7N1JjpF4cFdJ9mhTzAxQ2MozuAVcLQQGNM2dSxpyJYWHd1r
GH1qvlBoRGbJqs3N9Vg4RBAly3Xi2rj7JTlBszZ+aePzLRmVCGvHhco1MCvy
Zr/ZTK0f700H35MTBSR/gF2VAYuhMdzt4+/KvN69JHmTtkt14Wt3L2+U2Ail
L9LPp4uor1NvcR/SfbSvq36DMUjtb2Rbqkz5CWMAhOATMpRGOOJMThoJ1nqn
GNSrtRqYPATgEhb5xicRWOKzWdOk6lfAYiDRP/lp2+YFF71z/66Iv8B80wsf
ZjjDMi4xfirQffjMEljwR1bFl66lkvmS6XrnvtOfv84q/MS7o/YrZThHI26F
ah3oLoVCsaflC6gQDOIu2cY1KknU1kHpJD8lsSKfKBPyTfhply0Qj4iCJVrR
W3o4ANbC4QuzdBoUYmWoSvqQauJ8owL4HcAbMdAGTTfSKMYcxLHTcCuZHbaq
6TUpTo7EI1ygCCB8k9ykxAj8+nahVTiV9+/B410SRW9UGq1jfA7gNqTDQFxc
vWcqyopABJO+lbhWQOceLKQd/aE9hnpxStl/+T2kEXq3smDW/LLjSHNt2ddK
4D1O730Tkv+21hl5boxnIj9/s9h4Qa3W2rFJjizxZonFB7bn2shRRVpNQarD
5kA346S4HsiOQoyJIIC8kvyKiy6QU+U6s0MItZ31VUV+VVcdTC9/AE+RPXRu
hjnsH8SQT7V2u8Yiq9myq5/SfI5zI6pz9r68gUTalLr70qF/a0gb56pJFBYx
KvFUbGa1iwYIUlO4BfSZzlLdwQQWdqcttS6aPbOzuDLJGO7MSopBbo738itY
U/anPbxA+vRxr7OgJE5stdGHjgwCTsT0vUH7bLyYAdOD8TcYkN03IVUH+teS
osW+T6axvNOj/1IhJzD2yQpD6a46Xt1HmMvi3+Y3l9tr7+yiVCrscHPftfvN
WJOzm8bFFMPDxOiYW1CKzGWWYDRuVwO4NIhLCp3deZsG6/H2gW2UhKZq5Zv4
yKk0qeRq4cWMbf7kHqlelEfttSWJ3QKI4cmYcf4KPmPPFCeSnc0GhjVAYyg9
FlodzMJAWPkka+aVGIV27GuDkLnSBTxefSML2p9hFDswPQjiEz3pwl3umQOF
YgbMzK+3mKYLYXPqPTFtvOXRPXe4am/m0IdP+dq1Ue80GJyHrpYWoNlcoXT8
tXICJxKxwUR9r0RMUOvNPVGgcDmXGVWYu0HgomjqFzSkbOwt2S9I4272aUkI
fmFwkazbz6sArdW9T4mukas9NSqPMfXXlPBUlB98wtQgoyZcYO3eYK+9+mN1
SkFWDGIn7U2w6rKhrqPBI03Jyrqb0z//6VqdmQ/5BOP4IM+D3vNTQ4l9Lj1i
GpHuEr0WROSoXRqEO156FylbIcAyawppGXG/C6/eigmPeQFglraN8KRtPaMm
aQM2bXQDhYAbGd8O+tUnRF5kjtsiLnstJ7RbePIC3x39z6tW/QFCYgh2FN6W
31ujmnahUfSxX3w6fyTEAI9u2a5J0YYqe2Re9aIWy6H3P5ULTchy5pLrtkHw
cuaBFOaPP11qjbjGowLy7/kNkrzwv3V6vYGMouJ6ZxrG/UD30jlS5VeoLztW
DbYWoPiKb+cIxI9tPL+7H2RgzXkcWj0KeokEvgfC0Ip572BjvdlpUdeYqPcM
+MkmbmVKSG7P40+kbUeCfGGSnCsm3jo9ua2rmOs6CR5665rQILFB4mOJIvlN
qf5wbN/OqcXIKyta5ocxv2AGTU9xt+ufVUQhA0/Xu2DRMwcKcaQmgyiPjk6B
eEao3fXg58aRmhATGCgLclTAN2A07+IxD9rNX1G5c/Yg+lQtPb6UtlnkXmCW
MDhvBalVMfpinFOGNqjjrM6vfXOQNs0FhT9L/qyZ3Kp2UtLv7B/7fkSCTZM3
JyeZypiFcZJCEN/B4Dvr6kPuzg4cJr+pZ40hsPfmPfNHZ76HHKetb45spEKl
/TAs4MB7GG6jgbwenWwMcx6d8pf75mhrhmbq1/Oyc9geXxUslFLUxdj0kfwp
VMUptGVHeqxBPJ79SVkl8X/7U71+trW4rHpJsITiQQ5ne4VjfAyXcOQh0BnT
3eO8LCvtTHEH89sEGPiptu5vUCpiKvYlsGsBivRf8R5a5Fu7dYGzWGp7Tfx/
A0ih/kOgWvr12/u14BKMspQ4eFfMXw3I+yUfM0U4PrLk5T4ekoHsqTZaAjCB
KNppeznbOnDvjwot2aoM61A/Xq4dLjT1bm5jlC48S340EQtSl9Qb8Xe5SGq/
TiWzUzKEAMGIT/T9Mu6h1mHR1Mvt0JNfs6WlXQWWW63yQ2im1AomgQlyJhqU
+Bc1wSWnd0rkbUVkPcUfAFP77cVivmRnWZKfsWI+4GtGlUJDqUyo1TUAZjby
3hS1BsRaV/rr2Dnq3T1Oohu24TKz/rousyg1JXThB1oxROGp5WT960/w8DRX
34+j+WysgcgYHouaCTMEwa0nyDdQuxnZsIfbr3vCB0M0W7L/JUG//D0QyMCG
wUczHuYBXOBJ5+rwaOE7harAJvi7hfPGhIauVluGhP029NOx4GiaP/0nCG8m
YRCoU+sekYEdGUaavPQOT4LzelEWmVZdKEwQF3lVpgQov0DePwr3VWDeg5WN
S3kC8foyZF9MNvRz2yMMHACj0KT0Z2JIR9gygb4kyhyyWWlGDqP7SZuwJf7+
k3QED35M/BzGR4+jtQMecK7c99aCOFOhNPpVMpJViNybKPumCb1HMjQLoTeA
3TZn7nim2LL7116R3101MoNg/Y2VD7pT1gz8JMj6dW6F8SKSgmq8XOjMD58Y
zXpRUMOQ8zF/SPpilxVMpnhdQ9mxQ6oOK0pqzXmQaS2zyKKumUgbXFCBkGw9
QFl1sTh38AgyATi3LB3/fH2Zu/W4rcVjbHRYFsSOfY+4FHArvnFJ14rmLYHz
N1Dvk70Cdf58dde71fPIbIYBiGPY8I84JMv1DQjb1BAQ6KjEEvPUmQGPIvuW
B+AiAb3Jy7Ouc+sZQL5aAd9PFQXO2Qx6eIcZ12g3naj+dB8ZqGK2XRbOb7Nl
3+1VNewLxNbq9Mh7gS2pgZCbWL5e5hDNkRCwibRIES8C8sZHUIUA6oO4Otm3
OZoZtkku7mPm6F7/ZIidudkFhdTvxCMOCArrCWyYtprYJRp/vcds80TmEcC6
i5QLkJccjliD7rBEk4u+Kmp2VcVZk3GVInDKmRx3gHQu2vi8gZfqleGypNVK
SkGIN9AGk6NRt77qT4jULMyBPEWwCz2KpLpy//RMlWExTJn6DcGDIQFCjYoJ
1r8p/wOSPcIOvpJ+OGSZRc+FaR0X1u1liil7yOmEBdCjC0cl3OJVBLBEeW+Y
CkfAK8UPuKdW0cdhxrKYEsTVnsz4md4MRWeiPDQuiGecC5JYYq5Y2vHEvAey
nHcdwbEF2v6VwoDAT6uk43LI3t4Dnjp1iaj9gtfzLleRyekdqWF9VFZSp067
8v9wP+XhLtCn2MUS5+Ih4BjWXTVPl5LDXGtZCk99cWcsZZx63Rr9QTE/nBNh
q0+IZXBJDJtXi4CTqCo8d0hVkGeVBUXRUVro7nzHNbXWM+Rajob+vXfSKpmZ
lHUby0ZYZm9s5oNKKJ2BZIHoVjQugq7cm5Zmg38rFNH5MMVy7pcMiZVb19tm
Uqa6nBeFdMMzXLKAauXdk0l3ZxeroXaltN4sbD+/2bP0M0GLdPcbc2N5EYW5
qyf0sIeJESZ6csiAxZpcTElIk5PzV1hcqLdwlBDLDMsRHeiwXvodPmxVuzZ/
URhMI/Yvga+ZNKwlkUvAvZTZgjpKrejHSgASk0RUyZ+L7Ng3abhTjtxsvCyu
t2MNL7bJgpOya4PfVe+UXlwkJBR3BD1bi9jFwD/zqILP893CmQFgVXRp4glT
cPygiSbpVTohSCWm+rQQbe3bIqJcvWIXT/x5H//4VWK/rnOeT2z4VLApawTZ
H04FwrXdNa6Cm1IBGgiJigBzlO8HZqcf7CSB1613sF+O9QCRQsIxxHn2PO1n
JGKYjaKrafbHe9ePW6OsRpxl2I7nmmcx/hl6dl+CsesjqwwvHq8AHZQWjknm
eeDfMG/mH9bzkrYYMGAdoS5Ksw21RaEiOKhHpDXdbckhIfiGPzYHmbQgs0k2
WjWzL9C6ZDGi2LrXvY+U6B8w3CDEkJFOyVGf9AqVnfuZqadBsnz2sOA3gg4J
Hj5QJ+rRwBwLHFzW63CIHCr/u7evIW9C80HOzszjgOvw9q18puACMrqvRxQs
8UF4xIaJaqeJv6P1Li8R4Lf+lvhDzGapc2Bt+MF3oe7RWs2B5MUKcC7VHnPW
B5wQMXYaa0Je1qLKyYLhi7DntYcJQg172fsuSCNujoVldGUmap9MdKvTTJl6
jPqA/1WXvXUxGPxoweVWA/WmJBYOktm1HdxJ4YjJr2ArJFv/PJsSYQJAXvow
bKGrtQC46LjxknxxNKuysSU2tqz3Znec9S7bOrVMu1h8HUQ7lkWIlXjxvWDS
0028lria2C6BGCoTGgPprkbktLxO4UBwSXfP91VpQ9gdKoCb4A4Da4SmK85F
YXBJLGy8uo6NM0KgzHScuB44PCbCQyeTB9L7oyfD1SrH9F8q9E9Y6tAQz017
YZiijUWzOtiGv8j5335D/iBVp/fWkS6+Fs7QwOl0pXUqQq+xkWmS9WF5czk6
2b5S8QXfCOQh9Q9hM3I/UliXqETAN2OACydJ0pmtk6ATBgeSPyXoc260ywx0
8NiWxf7q+ltWwm3wr4NCcvBkMCtZSNCp+Ndt84HREHes9FRrX9YmGfOQ2wPF
+UckPmrly1Ip7U7DnSqx1Tjy/F7n2IsI+Is0BJ4wx7RVfnjuPpjp/aRe14gS
xAwS1Kp+nFCVu2t6ExWc0AbNKbncQKodTWH1GVlr2v5r3x4pdbW6QqrlxsIY
zylIJgzAHKkRZZCixjxP1nms/IuoK33Na5TZ1KxJqgowV0vK7f1lXuJxwCPW
vEr1776APM2CCZruIcjmm7G2V5F3gz0nj3FAe8QOe0oKCBKmkTn83xbdV31X
AUvW0jYhRZhPoupEUr7z/mb7c3s12StCuXQgowFo/vqGYNnFdWdKNEAY6f66
ewp4ZZ72oUJUzocw2yO0q38C4sPTnhw1EvwOaL1WMePNx5I4BUiNGHeQxxVZ
rnaucHguGW8hXlOuOiy/a+MSmU1gcnxlWhNO5posZA0svRobiIbuRQUxjiC4
+LmW0uC9JpxAmrI6xsg3m20cnsYIXnyb8UQiG5GV/+VboAyQ+6HlYNRk03Np
t/RouJfMxUAa/HRsE3hPcosKbTCQ0ZzwPafeFQ8d7Y9f5n3JOnEX55zWKvaK
IHQQSy5tZ2Rcfcnlv2qq8HjqT8H8HA8jrlZinmMk/Zz1GKdtPCrBMhhdqKbt
yY9bZtI+IOlbhglum/T8TXsSof46CNV/RgHbtpPW8SPovi77Ucb5SqN4YSsq
j4okCJ5tPGPYtkkW1bYF5ACQfkBpfLgRg+AMjQj5awYMnh2a9oAdg93195gl
iQ/t6BN8pt7P5+2TG1PjsZq3Vw6pEw0OO35ceFcID6yUdLbdCz4qhwcsSJQN
0vwOWyjANik2hqd3eFx3B7qgs8cgBA5YrgCdpgkjlxhk9gJnBD9ScCxfYyeL
38IF8M14E7/KSUKjvzFHmmeNOC3wbfoIQuQjc7Os4Be9KSjPWC6XvaiBQAl4
pOJ6Bn00T8DLk867mwB/tNM2uBu2t+gOq9Mlx8/xhoicdtn6vRb76CbpLaCD
ui8OTGhzSMtn2r/HOu55hvcgaFgwfZW0UAGS85JIyywHEnGRcTahW8tHUZ2j
TZNopaYHTNWo6ChgdXgmdDW4CuK5t+6xwNRh6UYhgrrq8GNFIpFZLVYlI4ED
RMy0tfdL3JNKeT7KhXQ47YjsJwgCP/5AGgoDSzidlPLMATO45iW8cexlUH4T
cn45xF9vaoyGbocNmchitgJJXF5f6DKguErMcpAUXBaAPoOilVgkx7/hr6VE
zooQMuvVB5Aot/ScsbsJc8lypOXYRMAESvPXuXyCZ+zeIRYJcypjcAdH1d5O
NGWjYWOoMP4NVkWpWDKwQozzXi+rbzJTgp5tRw2GJKVEUNidu5OjAz3+/+tf
X1reLN10VJSYkaTPbQL+Oxco5J1mkaymQWJwrQcPIepxHNrzcRq+Ib6D4QZt
3PpeUvyr/0ZvuxbBwJiSO8e98zj8EAFkAyef8KaQ66IUNcyvFRMPAGEkKWtA
MaJx/zgPW3exViJGA50PD18wC0x9pCCqBviLUnQLdec8X7zLrtAJorTFLKuG
6wu5RMKVk92wV6YEBEduj/gwnJBu6uECJPbZAvijlwsv9VyiaZqNtD68vXvL
ET2Z3qFIRblOqa1gymoCWKWpLQvx0gMe/j4l1ZJVDYQArLoDbavWcD4XaHzg
g/cTECQ1V4iFUjwQAuWnRtVpW7cG0y02FQfjzaE+Thm/B76NuXHXDtWqNKa3
FJbDjXeRvLNP4p9OpYXwbDX2xwyQpAqYV14v3xtdZ1JJtdOejPT9fKZ0I70N
P4OtVeFIWs4z9yQ1hfwlCjQkcxthqw+ukVIrxlmJuE64rIOsQT7o3WK8eO60
S7hE/6UBwqd5dXUYdViGqelON0Yk1K2PlGjUCkh54tuQ5x/iB/kSI674gB2m
MbajjF2b5Qs8X/V7oSUDMcbs3e6CcAWQZSY+kXnE6Lo2PJfHTax1OrUTnUUl
nJwz3rIrxLgnjo57QG2KuAJ9P6ZdMGqED3fMIieVs5m34+ZiSWVQpt0VbslD
znnvkIKLdO5YIu9rVhS6njGTxnyzh3tIIwbnoxoE1CkosX6Y3uSswbL++O+M
WNPBov8h14EieYnEGYActOX84qz9JD/PGIBeNbhEMTMN/D1Efm5dyeTdS5vX
Sx6tP08pl4zxOPCYAblFh13qxpcKngdjaceq5QsOqPq1Oo7vtl5hHZ4fdAqa
3xpWJgMSXNLqQ8g2ic9WREVlCQSQhCW6XWXg1A/mJ4b9HXc03fUH1vvKQKd5
d5hZWaYbrEWciRjFf3X1gvsI9wc7XAMkVrp/pA6d3+iiCcPyVp/W1jczJyUl
O1BsdmmdMpEhUny2kF1/63nddoBqTkwof3UHWWBgf/nlTtp7VEc60nmpcbqJ
P3rrbwIog/EUW8eto+OXzVuf9LwJHDzuNKVy7Rh5gtp9yDb6XpyIhEyaJfR1
JJaiqq3QL+pV5A0uwFAVu2ZREgiGFWfToZBL74wOyE0dSU/pWvdZOGWiNCnE
JzWE8/TfZN9JgqGQZ/wv+u/2vclfF7MsHI3lM2olYMMi/bNyZ+lbUE/FaN2R
tY5iKirrgYF2hIdEvFnbKNKmOT9EJ++uXOFUQVX6zMwH8d5Nu9szFiei6iWV
7QwqOameKV6DqL/GQKnDpsaEbh0qEVDFq1dsG+6Mr+k02lXO7YhKPdPf9GFL
zAyGuuvuTe9k2D1VqvfEpscP3Ca01C8wz1H5J91I7dGkNyFnY5al3lmfMS6u
Nvh/Nxk9xcRGLTN8mizYgxpfSXk3fhIJHtY1IwkOsL34c/R+89sle6nNRnpP
Sh64SOj57JSiQz2GD/w3j2s751SuKAw2CveDajhVOnokxnc7LjxVAwqf31aG
pxxYPgcsN0vqFTZLSanNTB/GSHUmNBhp0eg+33Td6MEPmpk5cQuXmdMKVZ2s
RaDIbiNI9C9JLVf0IiLoVDFFGXeCM39jqsCdkq/0NmnRrRb2UWveyB45D6uO
rRMl7o8NYxP2SE1u2VufTTqEmQgOjgUplxBKQ30E+N7r8DZfNDYhU9LmLzOB
bD0xkCYyO2UQUfUHgHbCYxc8dqFcLAb3iQh4daBIC8QIUhLSUxppzGf1MaXc
iwtNb+B9rIt0oK0a6SRNCoefnCrU4mheTQArdkkmwJIROdptZdWEh2IQ6bLR
3Q8lqJnbEncI4GkBMftNwRGuWsegk+4HrMn0HKqUSXsHftzVxBxFOxSG90nw
GjL9wBVXBrulAqMV944UFim8nyoOLvEhAPIfTrerv8gNM9mtkHbZ2s2oHBoB
/nVS72lI6VM95ahaFuRGVYpMaCSw8VKatUYpMWHGQ5CTVAmAMLZl3urYMbaR
NHF9TDMlS3xUYJ7Cinf9eMD9cjgFNpnQX7C1i1s2plgMALRzO+S+z598jOtu
Mh13wbsk04F7Iu49GKxqwggfljm2rujCRjnvHJYNxhVzEgnjJE7boyYTXlyS
PT91H7nZlrasxKwcYZY+ru1rkcbghQgFeYwdGoH5hGmKZZTKjFiljD+ib7Mx
WlxblRlS318mZY9mK4macflN7PHqfUzk3kF6xt/mF1VNfyjjT71VKSEx4hiy
+jukrLIF5EmgP0Cf0WR0I4N3FNwGJkoDDwYgh/B1j/Csk7V4gtZMbqMRQMEG
cApGNn6kWkq4FsU0WcsiWsWdxhUj9bxinvS60XOZWZhMvhw+rDUzKNlrC+oF
v9RuyKGTFLcFaxDtKggTsa8CDhm9hUjYHxZXCgwA02UWt+giLDZXdaWSLrg8
0EQ4tzKCYL6E7oR9++FYbXpMiNMWf4PyfzH1d4FNOg6pKllBnEcDPmA9ZA29
RSZ19Y78fA74+6AphnpHpEG4ouCZ7wZ5ZX5Zz/3qN3VGANxAPmdwlkJK1BrA
j/zkKTEU+2lKo0VUWuA+ZcmDfuM+lWQuCBhKb5h7KbqnjBbeLFggghLOz6JW
iy6ClgxLU/Nv05rNIMu+ygnurSAWoylU3X4RWD6UUzez8Yir8nbyBqYTsdOV
QYbrP9Z1Jf9eKNhMIfmyBsWwDNpXHzhVdyqzWPqU77l9dNVCch4txiL4w7vU
dCyHZ2sQT3/hdlxKXAYg6vrTFZZXd53VZmsWziXAPfRWgUOMRikBESanqxNN
TczM6eb3DXNr6+p95qeZpzcsQ0NlK5Xgd8vGxeP9t6wtquZyKjQQeOir1GmI
9nNWL4PakSZ8fuRJHAcnKZqHpZN1F18+OGs2CeNYp3djmqR6FkmHYm7aBZlL
Z5ya2eei/kdpN+jBSLUMigI/y8IgMmm4mbTZ/2r1ElgwhAQte82tAu/pkRnt
KWlRaVgrmpCC13HNENtXDbLDZ4YrmyYE7x0WMTbNDkbx0OeQG7WzCi+g1v+z
wufAGSvXiAH6q4oGR7pTzprKnOZlyL+foYCpspg1qLSIQMKHViScVvFGyu0M
9Di0PxVgaQCCoZYJT4WOxJiiZZINT4PFPXh6rF4zbUy3sNoS9T1nrj4sqs66
8agb0rSjb4ozgvw3gONvH7aCttZAyRhVaNMd26eVlHN66xcp4kRByTVY1DEB
EUwtySNE16pIfS1PTVaDK6Jues2d9m27Q2fU/SYgEjXPx8uBWxVMpbxFCpL2
9KhTkD2tCzGArSnAK92EFGV7FtDv6SCihfiiI8EA9iCajeYK7wTbwNb1VHxz
8+wNwAvB+bgpPVEACyaBA+qTIremtXwHCQC9Ri2s2FnXlElY+/xBzdNn2bTS
zCIFbHrlMpFubyQQ1D3CvCQWQJ8CtfyeCH+5r8hYKMg2+NXV9rLSulWL2oDj
Ksicxc1Tym12L8XkDYhD3sjZYswcEmkPss7q/0NPdtiPAoX50RPtnRGlOV38
Ffyrtv9p6mI33JgjDc11tOBB3F+vktMGFpTaSLxP93ck+W79pkNdFPBVeK1z
Abl+JY0dA+hUMgM7gzeqhXT7NJM+GjAQ27Taul1RedU9kFtpnfvmAaevI8cw
Urfjls4qb7FOPjpIZ7SVNHbAl5Gr0eBX0UAqR1Vx8i9J31ctU8HMJ5EPZf/c
sLF3pGuiUzXfJwulNTFVHbLVu4e8b+ctjjQOeX+QyZX5qJIu57/a7XycGnuc
qvDedrTw5emLjDGB7QSv6erQ/hMXvKeCybWxo0/WwhmxGLQn7BjMgMR5NCgG
SgGXp9zaANhxhKdv148rxFFkC8EuWHt1wLiFM5nir+qs7/0pnIlFCWvnc/Fg
4OfnSULLntiu4/54M8bs4/tZxnjSLf/4exhx74R1hHkMPOLONDIfhbQ49lf3
3OD0ExqNcAJAKDL3vNa8jhSRPUOt5FEt+J0HyD2NBeq/nVqVbIoEyEJV9//J
jC2EqnH+l2WFhUpMxSb6v8/FophXM4n5frlHSNh1dD3Mqo5ZyxXLAhJL7qe2
JYMt+nDv/0WkOzh8rhD/sx+rhdhqZadWZm1DRF53HRImIqbQc5a3tVIfyxuJ
flC5k6QOMmiPNg0Fq1vNyI7L6CMcwZMnSpHQEaNp0mxmNkWndWNYZYeHO2fk
r3wc+ih3P5YihqdrIjHr7HI+sy1R8zNhExj+X+KRuK0WVAwU89lZw8yamm1J
hk//WQXn7tLBeLkwDLr88yOB5Q8MPERz8JLepA3qwx+sZDR5XnoH5jCVCSNv
tMZbNIayEXqGzOVsHFb1olBMDRzauTmaYw+k4Tc+Pymqm/YpjnAjjEglokVf
RojBM/w4llzh+VT7h/vRhQjO4su0Mnio1KVaGq1FIoPNqwaT2Biu0XILUM/Y
BhpG0PnpcZUpZHa22gMP93rHgG+UMZS96VE5NVqPPDizYQpLV27E4Jev0KZG
wfHBys0c3nLdgzALxDPdBLBxxsQ/0KMdgjHRNVmiQ8cupCEs8W0R5ysk/oB+
HiJYQDZc9TVZVQglkMNP5lmtnTD29WTANpL2Anp2T+N2wSEDjKVv+Hx5O4v8
vjUyjYtwxUNDKLU/Db5EC/rNGEUt50Xor4BTpHE4+26fszg5H+NVcROWgBh3
DdDxEWcs21Gb/RzJjDvTxClU1lH7bYeJcj9EqFl8jlTC68kLOXZH17yYL6EO
byLt/9KFKiQvd7U5E63eDs/BiYYk1t9/8By/U5p/X5OMkTMGB8tDe2Q7tnmn
JJNiN47Xu8pwRrkCC1m1xcuyJ8zn5KQXtjjQwt3q49YLUfrORjbDFjuRnYtG
Hep1SLBGkIQ0z7wG+CRU3LLOcAwlbcDkN0YSu94fnkdG20KhpY0AtuX1kmwI
zayP7PdfpQcqa7Vev203RRiM1C8QrJxayPVpn4aNB1vx8iuwP4909z3Y3N8G
FLKj93h9eWQKLHMUIcKzK+uwhh18HJ0ZkCdDV7mTlUgZI+5QFbFO/QhggKA6
4TJfJw3vn2OSzcwGO14SVxAuClkhc553d85XgyBZdjZ253HevSlAurIr5eEU
i0uNW5J4yUrUYiupLcvlpYSwzPIC4nSgh8JzP8IXlA2XFBO/xWpeOnIMxe4h
FgQBci2JVBRtlctbTCITmbRDZeFByH/jOeyVaYOLx2VpBJYuf72wtzGzNuvP
F+9+2Jvs0bN+EC+QWdSGi+g+Nw+l9aO3NrXUleJrkmBB0n25RJ0QeJiyhFKP
SBL4nfUJdgbyxER1w7v9LIGANQQTAgaDwv20sJ980uN8imZRY5VSQ2shc165
NRykLr31DtFbkLU06E+Znq15QpdAL0+pJnucr370jn3jwc5So68ULMWzfpIe
Fc6lYYffLDIqaAjZDecAL9a4bmowklfSwk55blhsOj5W09zYIuECEGszcNw/
7404mrWpzpa6uAE7sVNjJkf93k7jAFDLJ/NY+IsXwGzHw5JLG3UhVXfHBdco
OYe1mlyKAjA0cfIxmG1R9nF+LjINDHZ79zOZuwnyFabMTeS7NbVzHk8QquGa
8Wb1VvSRFKU+xf8FzJltGzgxpFoMVI2Lqe3P2SidazK71PgUJVbgJ7rqoZ6n
nNXy5HQq8pJuRP8eIjR1YF9YGaLRa+a8nQA2YTnn/JPXqUmozGSuzP2T+HZM
o6/pqID4k7Qa0YqnSB46qlHG9ZJrAO69On8svbNWTe9jVHz/r6TsgfXXJQFp
6H7z10Ofs61Ex37njdyShUcM2jMwx+xoUPwvT3WlPDOFmGV3paufRdab+u7e
ejfnLUqwsrgSZ/Rq4jduPmB6c66d8f58yboTolGKxP1Oe04+yGFhAVF4m5Kb
G4dBPBAFWJhjUh4qTwvui+YuVmmmyph3793KRBD3kW1ejWFKPJDmTpndkpLE
sH1VKD0PMEkX2Op91c7bpL85Nltj/KUpRMGBrzux9EHKWsZ0PPDy19jQLJFB
fKWSDSfMkkY5JhgtW3OnSrJ/V+agE+6vTLkf2kbRsiUiPPYdUnW6l6k1PlOD
jYk6UY7VD/rcbzCIAYPZUJyUUOJ6mUOyYpW85AhbzsNeoBdisxYb9FpVeSMd
kbLWLdCfBSc55zva+RTodPS66gjeGSIWU66EoMnbAhMdwiIVpdmnxEGgqO1d
o7MD1VaQYZblUCujOwpnHwPX5Sd3r0cFlhFZbTvPwOn+m+Abqxk4eDTeFp/V
CX78c3Dh9J43k3MF9E822JyfnitYRP5qjydmThfdEakVMfef8y6Y2ge3/xAl
s/ZH33fFBIIv60GCI4jO1lB4g30e5IWuF2FddvRVyNewKN+5aqKmyU5ceJSn
LylJcn5+obbZD7er9Qkz2OTYmUEwXLsVha8xfYukEQq5+myt82IpSNQcuRHu
5d6bft7M1GpCmwp+dxs3tH71NgDlMLhNDwgu48QuQ5xvTXDCUoVilbr3h+va
Ju5iVcOAoSYcVGXd/yTbREV2u5yxv8K/WHpCyZl4X5NUij076rqqvwdMdu3a
D2OakvvAg6eDObntkHyEitog4yUeRIBUoqjZ9vOxMnvnkXJ6QQAdPNJ1DOQQ
gxG/4R+1YbjOjWRX9N7D5u8PjhKfFSPI4FUOVXODLdhTmmN/CGwof8Ht3TmI
4EZg+8AJtpFH99OIrQo8Gngwh/GLqLorS+9qOF8dPCToO0ffjJVM/DQylpV/
RKQpgH15zKm0D788MUAfgsa52EjFt23AapcU3rh+g8lkSZpfpUADifr47DBj
Bja4FhMlZwlKDd0dY8QZYSdy08sPUP+FLJ/pB/Y96Ph3Jtx4fQ70k7B2L4It
90Z+n++hxnjnInBOCbVQ/M3t4h16Xm0gj+swPMyugzQhV3lUAr41njydMaRF
2M8UNdqqHAXCKbBOQkVU5r/ezkqtxxrwAV2D0AlBS2h8FiiIwIJlEp2gW9LJ
rMugZunMZm1x9TCz6zc1tvSsIzLVIuIgOfTwwuoTebMIITOQ4r7B+o36KhYl
7WT9bDcnAS/2Remz63lyn7Y+UqqIShLeS4gk8nX2Egb5Qz+/N2QRJBaPnkT+
vv36vj79Gg5/iyMLfA0hTTosGTRk0ueLa9lWJy2neuePlqs5BiJuOsgL0doJ
Xg0uA5cijRQdgQtq9RRcDiW9uFN8jriGnJP4w5LMgB4Rhf/HoFord6UFlobQ
3u3hpPt8fUurcRvOYRcgBLdVtbox+CPM2AWdRFJ+rUBJ5uMcrFwzzqKDtlBb
5P6ci2NGPohk0RJVoWLFERnr0nRfr1RHsOFDHyZz3KTn6xVo0BTbCLGV/FAv
ERA0usM3NkGzy4C44Wg3iXm96s6d5nfxEOmle2Bmmy/8jcyMeOKQA+gahpUe
hU2edjy79u+Zw9LWYlFQA9c2A8cBU9c6yu/1Xwk5rRYMorgkjXD4R7zjZzA2
ZPXhgEKVmlqDb5puOqxya5Rh48IWUgiC3RpXvRx2C1WK8S6eyJm7Agbx8K3c
Db+kVGa405J0iQIYK0p6DrzPpDrnkkv+sVT25v/4NcJkGjhhNQeBduoeJHin
PWF1c58bYUMzd3iF0Wcu8IzY7d+yp4ynuZLfWLpnjuR+tqNw5XPW4rYuE8RQ
EzW736wNyjykwsICQFQbNWSs8jpoKPIZBNSMU+QYPfan5OssLH4oC/p+NKz/
wK1eKcNz9PoIfTmv7T6XoD/5wqZ47CeQ9yEgbfyKuoYg89iD6MKuc+iYq2Ux
FslT651FRR/Nce1fxqJRK2+QJVvlnCfLp4YFqwsTcayFmuiqlBEKEyvQdV6g
KAxiz09yGRwjSbRNSXTAKY7L8+EDzj1JTcaJAz6eqKpB7rjB3FtEu5wzPYTt
m2s+8YGycJMRgbHCedVbe8iajLlyh8FpuMD7Ql1WpoZYCSit312bw+1EbxPl
6EI4XOm9j2TwFddK9BeezvQ+LDKvmCLLxxmFHJ7bYh51edK7eShe56NkTStK
eFcdx5n4LUNkU850TB2RltnZ3nheVs1M1Ng3E9MIeX3jI9+Ax2/2Fu5Jp17H
BUHRrVp6chdpsVDjMs9J7tI6ISi8CaCvZuBHSasuvnZxK4YI5cXvaOatkRjL
eKlCUuXXfvqYFcNozXni4fWn2BjpmCQ8P+ch4nILpDVZKPi6Ng5cDOXZNKVF
TQG0kg7bMYegWVRcb/QlyXB7WC32/EO80vgO+UA7dIxR/Gw/7VfuXNGxVxzp
Tf1lbYvvbbt4QmI2OCiE/5KjnUkU1EKIkaao/ZAKdpvD85JIXh/1971IQYr+
DX1snixwAlYkeqSrgwnJDkHYo/H/8YfJGDnkOTjROre1m+D/9hPSIedM9Q+o
un/Swb1J+QG1WguNa5yBDqU/fLDtT50RL91aN07+0ItTnMdAnvvkzQSQs0Ke
6QiUf+ZVF1xTC61XQFuiiPKpc5FVwbDBir3/WN/EVknQC8/R/gjgxIklWCJH
vr3M8rYZA0cHiVfg2YlT72e0BH4aAsFNL5nfAGVwGS/dV1ZfpTGBTEf7WZXC
KoGAjmeN+CXecCPIVx9bJ9WGDsfEdFtiSPvN3Gs3fI0plLq6QvB+JnyH9Gb/
7ECh3V+r+qrJpnc/dXAzM/uAijbP/Y3x7kJBLdg4GsDobodb6bO6AQZc31ny
Hy56WPMvuFz06Whb+GDpBf4Tr+F+iGdmW5i5BNwXLPCLh31b6xdvdei2O4Qu
3XYEsPzOVft8zdlBXPbSEEnRrHgctU0eS5E3Pv297MFdj5E24VFp/HEJos5M
w7iyIRCHvBCqxvt42Evv2z+vGax1+BG1zLZGk1uF0GChiTYErhGjVo4ovJ8s
1ILym+cGCW81776N58sQQIzsMBTQzTae73NZjDXmVw0/zEewB41WlCH5p9hX
emIhlDK783lG2iDwPG1zkF5MbHghwBvPG5zShDbKcEeaFzRq8/YpFcgh968t
K7/fORpC2s4q5pTgHfqjban7+ALR4ZNw3EZTk+zUsYiLJWmt0KDrfSQToC+x
GFzAMNfg3lZ47Si7wAxzLwMNhUUH3MaqjPNOSt5OSRXQ48HGryBQWNmMB6Am
Ah/HKLFU8cXjJ14UUez9eBu6ZZhDF3inwHvlVrpFJt2vCyfYsKiMZaZyT4au
WG4hbItCiEmGAAPgZnByXHCPAAGLgHDvKUKUf8YfxHKlQx4qAtp54OghGN8B
2cSLiBFIpP5Sd8szR0ay8Cw59ArhOfkcdQ2fo6V2xZuGKEfvCYcrQLPPF1Zl
t2FAH71U/GPcOrJ7XLKYaGK0ouEaAqUYLTgFaBSNI7L2qF53IQLjtifkYYbK
OwEIg9LpyiP/hybZeBPQf2tZcfsGGVYzC4HydMQbTCRGdxvyxuhkHH4Bxo42
42FYQoez6mS87NESVg5ujp/OdgFO+YPRH7l5CeHdLHb9Z7QS1cxIzXB5DJGw
QR1QSHBO8FerML/bOGUuB6iPhUSiuljBOcuFIRYyzXJiMvBuOLwHCvf1MIXu
zcVHZBcyaj0VehdJ71faoH+XX2JG7pF1DJmzotFAnqqsPwCbW4TV+b/TguXT
m3+fkPRvQuydkaKTu/w6wMD1HmpCbgM5TD1RxDZ6xacDFNp9jQMQknPe/nBn
UcuLPVrO7sgtv5ZD9BPLPe3fIRWyg07MzplFicndOyqI5MqzO0KqMs3wtNjA
J2ctDiM+HIf9XL7C+LC3ezZ9CI3vQUEi8Upy4nx/kLo3y9JIt4FVq+5zxFyS
AFJuM24cTdB8z5M8gLY1pD45w5wL9UEDE46HFvKvo801OficW+xQDWk6oMEo
WPZhvGNGjS0xkAqhUnEYw8GvKW5kNwYNqLaiTjKKVL2DVoociUxC12XOSirc
2rI3502NQTPnMfrl9ZbNUpgkKEuW01EipCE2fBwzeehmzvvmxsV+xuSFGbh1
qBquVi8/7RbawF8cBgsz1/+M7F0DuCc70qXOy+R7kCm4iiLahf1vRmzK3v5e
hJGYrpv8ZCUm+Zhu6KuOrI/gopo486LSsfPNLT4FQK21ta2YpKvmn1to5Xkf
ritb79osQOQVnSxICVoLKAdOQ9HoPxAheBMSc2jLcwvYnERZauZW1XsSK9od
DpLHpHGXQ2txzRZtuhXvevCmcomB1u0ya+BJ+OKWtY7wMzWtA75KD8S5gA7Z
tNAlMCVS2+vWKl5Ym+Ch8z81ix88XeENbkkBitojJmfqvv/V9xxLvx7ZpyBT
Mkv9NsCBOFtYC20UkUfOLLgovo3Guv3MgQhln8l18eIc00VMVC1otu1xKWEI
ZP9rGiTlH+nlN9Xsq3pJhHq5JocXoJnz23aUdAFZR1SH3cghUFY84wUtxdkv
pYjIU7yCl2lMemYbkrszzJ9EauAeZgT1ZqAolMjz5n07tcALNNBMzoFyFFOf
Wz3lFCM9ITnSJ4Lm+7NPzbDCHBVxG8hkNtPLB6jPSCa6WfHHocHQ7mvu8d5Y
l6rNJQrBCHg9czLcdubW4gVuxSFwG5CM2Wt2B+kpsnQAc588Pde+CKMe0FY4
ucJh5OsFkXyuFaZj6W+PrTYdIIvc8nF6g9y+9hG61RhipZcI0cKZ4eSbqoWf
2Y5hqENHl+eQ/bdh3uluJ/jXb+cZ9u5/KAePRkqkKbsMEaRIs1n+juwOaK7C
ATrei63JhNpsS1CvthzqV5IcfrNO4YHr9NocltntR9eDvdBkSOj4XjsceTzN
whY3eRqX0b/WopgQ7AFciLdHJ2Foo3d5hUxoVyquSNnkXbcSDeki8kO8rZG5
KbTi1F4g5118Ve0NDFUAyxtaQgKkkKfztCSFe/NTGerzBOV0hz8epE4JfteP
4fJpCvjYLrf6DTpar8qtNnlQonXWlhEr6XrWjneRrHFYXZ42KJdaXhiVxAVI
mWOvKDyDDyAKrwN4RC6xho+nT18v04y1BqU0cUSgtGpeCvYYNjR0o2Gw6TWV
DtvSKk0fj7pI8835Gh53yTOr6yZhjCwX2W51u891x+CwTbLW8PRgT4QsOxp8
rwEYsxyz1HPgKadP/dEGVbWcq+Ms0NxyF5lJ9oYZNHbs0IlcGdpFBbaqf1Tv
xVg55A2a+4/Uovf5TScYAnqtmXH/MU2So0slJwfxxL19vhiHvmH2nDYY8qfa
qKLzbxJq3FxYOTfrvuu7bz8E/bpXDu+hCwBwYVzzOc5KYb0Sikp6NkfECYFn
WzGZlC7+h70HwbgwFlNZNtxRQ9hP6+eMYgGXCGhCu9A3L1joJZpMaSY5E6Nz
u8N8lswSN3vdDxCX4LJADisuYLNscsTOVsQY3x7qYQ1aVCUpouLog66fGHmx
6BKpXwExxDlcvlGysfQz4nmosFT6z5fmI80uhPUn5lPd2hbXLyIO9x3MKCJD
24H/dkwQuwCaGYRIN91sLkjQ9FZ9qpZVGg6oCjnpiLBAbdmsuXHrpten+N4d
Zn24URCmQVrHSc8hKBpkK/oJ2e/TsJ/LjrOYJW+t3MV57mm89Ja5xiVHd9V7
9mVUdH9XfAIPVUagcFDsAStBOcQxFxbSEmUrXYXuaP7CkfMO+fK5LepmFr7d
50WqJFAYzEn8lnLvHMS3h0IvNlrTujpgyzEhJpDYlbaCy5Kk0mTtNo4Rtvmu
NKb6XjXEINV/N1Ceogdgmbj+XCxlknCGbozoPhhjTioC/YnEm7wjYBsUSlj3
SQzXKapMtnx5EEJJKtyYD8pHwXAbJH1cJ+hBe5xQNkv0MeTekwvmc3fK5Ro4
Uku0QL30mnHrDUY7myV0HcefBkWhNceoE2Ix10ok4dRUBHuax4TTMWEXAgrT
eOZkitf2LO/TwVrV0hn6Qd1PR0651GMvDsagJqyEot7iLUNfS/pHRpvJ9M1V
LG2vKKPT/oOyDES1T6sY3uEHv3fQxaI7JnHLhnzf7c8m+8S9Jxk+vkltyeAe
uK3YjkaAwzTd8CcAdaLMgoAflCcuGhql0FipHxQYxfBcsegzxIrTYG1CwtTc
PchIBN/UOFLjgfMrC+4kL/MpBHqxmnoJWuBvPGDjvl6T5ZkDwHdp2jmdXANc
2D5t4BvWSPnFgqxV/LvYz0VEKOuZxSj6ZkE7oYajxtfhR2xSUx5U7OISlSye
7ldAnGoDVtDenKqJzKG1NqNpZIdrNzvUbkr/C3S0cDl0CPzlSEp3uKHYGNkf
9AvzHwmnQpPNj3V01lVq0hr5Z5r8eIfojJBeMfDfLgFEPKTtvVxAz6G/FtxI
B4pyDmM+Mc1ShZwKCFjEw6SlwDZ9SSV7DCG7RIjcdbTrnv/qCdS5ksjAufyQ
bJ6Jzkb3c4su2wxcrHiAygHjBENWHmbXq2zge7uNQlUKgqTIyFVQKiYfDApZ
AKHF6470f6q+mLE8eM2uWe2XqlRtWS7SZSbjudE5Abc08hAjOpXmDuuBmG/Y
H6HXyozHGIgEbLsVWLJ5UwTM78cBT7PRL9B5snMm+bB8OmIn/TahuGBq33PO
hSAsAG2pFZ2fie0xIqGTFtufYOXkw2iZEPcu+lPZCXC7/PDnC7Bym4Ez8jzm
GAvwz7AfQVVjMYN2OT50Mu8r7j/sZ2xV2Ob68w2uVjCQbWSVKS51elsvjo6X
7vQ/cnLHuD2dYo/APRWRVoM97VMVCsMUK9XpcohKUP2rQ8IchSFYKfSrpDkj
jhHxVM1jnM3SBXxSwd5HGskxG9Y9ZLN0DhFVi7kt7gdzlDQu9w8FtS76Qs5e
hGJ1nDpf7YxTAQXLYIF0uLzMwk3nA/iUcxXoY7DbnNNwun9VxZSyvdbIszwl
VWicXnpUFa63y0/cR/LXqrJf5+vaD8fJiUQ0TT1N7v8nq64SloG2gUm0HSZw
UfcFNqUfrmSIVpZO0HnwDd3IWgS2ZwDaEF52n5CaDuXSzRabPOA8u1OgETy6
IJv+fuuN9mpwY8K3zvcbIpd15mZOt+lA6KaXX7ZxEJa8rQsHl+n3smyKh135
8e/5OD5rlhU+4j7DDjHIxlIA6OL/uIfnZ8meAnd93W57zmcx1CO+o8dcsKtz
iriedZFdTo7DSH7c8x2aSsaawNgjBy1r5PuuPyDH1Pe0v5BR5m4taYXml2Qo
TpUASyto4xAWXUbhhJcuP5bNN7YaWGWOCDMaSHjn72t7dQ9NR3icCuh1c1+L
wF3SBoASwna9Ah7ggr0WlSZ5vQodSc0rinJyN2ej0QqMZstH0dr55LKMc2hO
hrjy+xtFgm4PfDEbPh75GQlSjHSCVeh6rUXrv8pbGkEWaHlWcb8iJK8CxvSe
aFIZA1JKFQNPnEJWmYu7VjtaPe6E+0yQiHHfusRxnmTf0Xl/e+VkJUemJ/EO
E4nIGvltnYDEr+qHNKXDZ52ybH+/luBAZFdKtOsGp2Smdzj/vmL7X6Y31xNs
PbI3V+on4QT60I9EpVkYzEgs5IVganEMF2qzaYT5D5ogUsssI67QHQw19RXG
5fY9ei+FgxtI5LHqlKneJpZCwePd1Ao/91oeWYy0yaUHNa21Kv+jHlds7doM
wnBm1SzDY5LD7xxUUfDF5eM0mp+2oEwYLblOXMSY7JJcrQ79ytxexkgBcwfX
Mzf+ydCE0ofmgelgLCNmO8lDy1CmEnDo4ZL6kd0nOMi0R+t0jmIqJX9EgBXX
uDmuj5aL7qXoIJDCdjoyTWuLF8tz9JdM4NCc/Xbc1jh7bVgxgGmZyLh/EA3H
LXuk9Q4s9haH2R8d0n8kgWLPUurrBYsys+F5rlaVOjjPgzhyNte63m5wNOzZ
A5r8POEAVoEvL7A4A9TnfmbrUEEbqcZEzVUspOD5/GE04fj4BRsbZgOwjV9i
UcjLmG2B1p0eogfnUJLTrZGvJvvEPCKMqDs3lXInaGPYu9MNFKLyfNpLqBQk
8KhRxDNneqAjymbLuabzAkXTIHHcrATvSfblQJWc21TLo5lt8pVQX1UeAiO3
j4KEVQcfw+XcV3VOc3pQP/Z1Ap1uq4W+mV6hJzjbWezgfDTXq8xHR72ZlhzC
pAQptHXZOepentVjx4xt3zE6PTsf7GTET4IZ4/I0eujJlUSrHXMnyI+aF3jr
wip808dR7oFiPoPNlVuDnwgLoqbzbsP79pDaJ9QlwuhdQDVXB52ubxqIvqP7
pTVIckL/FRXnTY0DqMirmQ1vC8UoB4yiIoTRfSRgDBX98jWe3C3GiGiBntEA
Oycd2q2Sozxs0xm5QMbPsiVdzCM/Ow8duE1/197gsy4/CBnW9Zcqtqdb9o2l
R2o8TJj8tDnUJkiUh/GlvNZFGg6Rj2oSTfAivnSbI6/Lk9ZXUvp0P3FIxf6j
EyNzuXQek10JJBqZaj5+MO9OfY/yrg+iItryfSnJHmtoZR4rYXb7UjLBb8HT
dFoJHyK/xQyVlas4ioVWnQFpwF5sA1J9FjiFeyjxuUxPVu6iqWSI2skRVvPJ
v+nSie6ZJZ5jn7TKw/3SfkoSpmlsn5nRWC+wSvNdoXFHXh2nJtVFQDOqxhpb
5V63rbdjuPLeVD1xTEl2EIRFWI18vyhVRR3PIPE3tzD4ABX9WvekiZkDLh9l
CCr5rM877MhkOlR0V5NBimGkNN/1nNM/XdnYVVlXFdRPE58erC5gpLHaqc0/
UkjvpFqQJ3CosV6MfyJOh6ZNJU2QVuCMoT62VUrrTAYMR5oMMuUNnLduXvLD
wD/x+IXr1gmj/mrP/cEgQEEPRYRGOEH1yqO6q3KMkBvvWTqeIn8PE5ootCd5
BoCYVqn59fKm9kFvKSFZ7n3O/YBpxehkqxXiAuuylxjYfP9ZTLHJtZMSMjVy
CFP9Oh8/LKpCnPgrnOzGU4JuN8B79KFZeZYB1i206IGioyNxTJ25rsZZRuL6
regxJZPFu9EH2+sXUXEG8G2cy7nSKbeIohel4h0mFmtIduI84QRVql/b1/rB
wl6NH2kbvX1JmqCjMIpUE4rvaHeAbAMS7ezZMuZX0+RuAmJ37a0AKGMuU+oE
mxy2TzIJmJU+oJ+Yg4QbZkHOQt4tkbW12ttldB8paqDslqkCXNYb1DcBQpb5
jXu+fVfvyGNdci6Sth3G0dT9Ku4kpyz+JIWXc/WY1TGRN91KV9/RaieqrDmF
iVWWmQzCYEYCkOZvRG2RUCm8Nj2DNx4/mwi74eo6gf4so7KFJW3jsmZHVIBm
b8ClQ9wy3yQL6xvnQf/83fWcaBBIQzpgHvX25+U8wR2b8hnmRafskz5WOYaS
jsaroMeUEROMsfMqm9Y19JIaW9sWwyq6tEeCJxO81TPLyZOaj5GfVR6BF5gE
CLra6mLMHYzMCq/Vf/9tDcQFIbjXPeVXVvwnL6gJu1dIFXDrY1kNSO14VF97
0KuAhrTCuEjP0j6YLbGzv5Ap1/96Kex+LNQCqXMLBZLR1WVrg3iR2KVpYZmj
SwijGBPLoOqTpG/KmB5FF7wgK6UL16vG6VUtimhnXq7BDcB/9BzJpOTrerRU
wxaG39EdSiFO0FEwF0xhLuZj+A4sFFyqj9346/Mh/onZyszx5iS/wQOsoXCd
SmHG+M5zzdPJ1MNcrdZ+FXUSCQ9M7gMpIsKwNIKPIcqKw9NOtvOCQck+7GXz
pZyZIn6maf0Me8l/hwphYyFrx/kgFyDJu9alkz4vUcv2t46OK3ozNZxuq9UW
xgUbQYFz+WJ5W1J9wEL6YcU5AZGjvjcchpSRKVlffyfsxO02nPGEsI/uLOlY
Ill0q+obiHAfJ86Tkyo1DhvQG3NaL5kVkzmV8383LG3rjUCw9WQQNK+5domo
i+crNOfZkZnBRrruz5fwsHwFbBhp9nO0KqJQyqQ/Le06r5PYn+YeZ4iWnAwH
GhlIfxzW+aw4Pddf3bg7K7ii7J7y2Hb8BVPHS7KUhzlt3FI3066KfudJZJWs
6QkuVVyFCcuRpA1zKMgrSDa5Ie9Gwb/m3y9PEcFvr977IOAVKhSnNqdy1lM3
qAxjkji4HihlRR9m63FcZWzyuxxTypGuj+m/gyft5nACH60GL55vLq8mYK/i
p+JtCDzNnMFgv1z+Oupylib9E5vY3ksC0EKjycZsjddYGuDV7ihsizR6ghXU
T5ZSh58pDbBKVZR1Hghr4ECl9OO9/F8XL0mSGMrVhDKc6QatoyGm/9Qpb45A
BuVkqGV3414ct+p2G1aOIPF3fywXkp123RGguGrtEGAXCWLvN2BChd5Bh3AV
9NcnH3FzVoDYBXEkrKVfRY+11iA5arRy1OKxnNCfUtNjiXIUMw8v3tBAwax2
v0qdEs8keZpslZ17nuFF5hAsgaj+UIH+dKIefTIXvDN29fD3FkMbt7bAgMGC
6UlSN0dluO9wPyq/A19DavW0J3Y5YbWwGYH5sNwSbq4FJ1ny4CLcWsPW//5h
euuqtUxiBkv9u7lTbRSRC6ECoEBDeRoeTRO5X8EVMKS4Zx6Zm4byjggDBSMJ
svcCy8+nY9iLV4UR+aEAvMYsprV7QY3NyZu0VaJTb7xWrkW+3vFD6JJWmGw1
LzHy91rASupOUxuyDLg3Sk2Fnkke55xLPfxeybmFjn+y/DOP/X/+xvsFpPOs
8B+FwKtVZlqW8oJNHh6yOEPLP7I4Jn2OWVip/njpTYw3jo6ZWhHZ1x62r5dV
hIhyO9y7wWk578hdKuu9BaOoLdNWfpS9Aqdev9tBqjvqgBBKgn/45l5o7poj
5t1BeOcqjeYIfrEzfnymSE5t5T+bm1wYLvi1ioEp6luzCbNMPFfOoLSAbrZm
ECDe2E891lDON6HNBBCx0U2Wen97r/AOQvY/OYk/ZQcCSNgYLt/lGEjbnR1E
4BF//LAakDVQvnPAPjJ/6hJypAV52cBSPM5MORyUL7WuzJN194IGspdrJ5Ri
P83LVmhn1gzuecGn4jYhuUKm17qzFBs0L/GJVvv3KN95T2vdKHNaI/qObQhx
o0a1d1MOgpDyx8jeiv3IeTITgzaHh3LuJ9PVCASpMIS5LoFJ2UcvOJDeITS+
oRDVWK2KaESBmvNkbEUAV8JSpynyTGQj3vLnQgY4KhbSgNOJe5/aR4SvfBVP
CDovUq/DZ/6Ee3scaCv4okrZiQomGT/PwO/jpH7Qd2TKOG1+3eWi9M7isEK8
htwXesd1LCZrFQvkW1nsXLer/BiHd2rTYLFf0p267y3SCj24aO2zfdPeKaVa
gDUkvXcCnq9FA8Si3cpPVOviWkaWn3u0euxv+E0mhFiPGKl+892H6FlAWxgW
Oq3b0UD44XrJzedEsiE20J2E2BZzGVYIIqih0lWXv7tT5uhWa0mbpt22H4nJ
YA6JJ6pvxr5DkX2W+KWLO/vklVXbPd7ZnxjHSk2Ld+fScV2p1Yr5vCeuDTI9
WIoS9vUhKJorRUmcFOIN1Y/Oae2urYFgGE+PXyCUb0NUUEE7i+gbtJ7fir2p
OV73+Uzo6G+gdUXFE3tG1eFtMaTs2vYZWNYhFLib5xsw+InKi4POYJ7naxKG
DNUAbBnmE+aqY2MSFFgothq9CbpdsBXg9+DPGP3QSjGjWpL57pwGt5mn5q9i
LI3sTOw0P/q44EFBsaIUefrWNEJOOMA8fQA0tMxODl/fQJjFVqFubCkaq+ik
CYC1O/DGhcLogwKyHI8NnYlbQjAYIIVp77jpwgUQZsNrWyYdL5Icfv3Xe2He
jLbTozE36qgcdgLAdOwWot0VW1xLg8miZuUe1ueh2OkQ0FyyNizAmi6TqtAv
jt8VNlJK4Jk+zEtJkuT/zx5eB338VvP3Y0KNnDPUsohGt8IODKQQB5Om3GdW
R+/4GbSBal4cFeNCj9GFWxZApePcVO+FDprDYR/ULprqkyT2SrwmN97ptd+Q
PvUfLez3WOUVc1M5mvY5m0UQMXs3tJRkvDWLQdNPqFcEzG+b+jGVQFDsBW5i
QQwWCDiepnmQNOcWUpLbbiZVk4h66SEe7FjLdZHEyQmlP+5UK1LIKu7vx9/3
kJJMk1CHO/NYDpAlr1GXvWvB1OZegn0o764laEqZHThQTjf32S+owtZx343d
tl1A+/J7SR1vQz1fnbhVLQwOMXiA4gCVjTZv3T7m1xCB+DwaEOYe6n8bZlCQ
0pngzoiZlpSv1MOgoaHiJQThirO9NV0oGJTfsPOPVvIzscO+SzFp3rC2qUqG
JzFYLfHfolqQxjwNBsne57E5JWnj5eZlAI4m1LZZpza0FJLrEE9/mUobSGJh
8J1RRW1yjo17qgsvnJtKpXBWC/1Yd0xXjpUCtasNEA6ILoX/azBrO26IpDFC
HFO5nlyS8JPR1Sh8hrlvXJwLEXNNTNwVuEY+Bnn3298Z4EU42luPaRCTja0D
rteG1YdXR7P0wNfW59BCCupVm8cAEFNoAHODyg9Mkm/BMvTNZKt3lV6qKzTW
L/KP1f98jVl4m4EGAQUXC8GFScHyVwPOCUbhQs4MJBwZLqGRFOy6J8VulUey
IA5dQCt5fBXcjcODiRWtity4yw1K1uYsuQfIKvqubPEx1kFrMv82gF2JOiLx
LfLIYFSU9zGOYvvBG3H9ntuZHXr1Uimf+TjjtNht/b9Y+mTnlYr+UcbkENRa
DpiMeLcmy/ccjxX5Yq/xcNoVCfkJLlbQ/4EMS8IARHE2rPi2Mk3wLY8P1Ha9
ibK90LUNo1v1zBsytDDqkss8Mu7FeTNCeTluWLrQyhH+OMdzMsaau00aNV+3
qqKZuCJjnclhrSodI/B7oZzF014qYruS6kYDx3OmOFFDyLZ0pMKRhzT7zf+f
q9HyikQCrHy1NJMk4ELXmcF+B56XDw9qa85azXeL8Jt4lRxWJruAurv697Bp
ygYjpFt0nerNn4LY+1bKM3M7UG3fmDg4MdBRwcDwkjECbIhLXCHTEwSq+OLw
T40rUcfT+dxDGpNrVOVFpMR5cZk2Ay0YhQkHlnObI66VYiASIM3BvrXROOB+
6/m7miArJAixRH4MHAlNqf5l9/rClCE8Klrx45ldD4MkM4jPVaYkzG9s0iIY
uggk/JB2eytPtIuF/x500hdZKMF/VrhJhCm5fqSftl1wUnrnhbZ12JWJVmer
xYiaOu1inEh51CnO/JrAUXFHYlJh4LMfDpZKoAS56OzVucZNysBpxaSLT79Q
Vx6LAZ3lAMWjVWpPPsH5uvahm2UA8xiJxzGHCjSkxDZD6uo6bdkT3ndSMoiQ
EPuHGvrvGifdNrNMmxjgVM6nehiMWsyFJbZRTCBwEUWpytQL0tffMs7fcJRv
+6J59H09W5iPV//eJ/UQqp0UiO0eAXq9asIg0GippRh+HiavedO9CdUZpWGT
X9s5qkrJt7oGVqXzR/aRB7V0RF2MJRZ2lmzHjgHkT8tqcF5byDDEgYgUFaAo
Vl/O7VyVZNpSSe1ia/rmU7r6X282K+cW0wahKEwKymlkYtBmsUSguWzCv9t2
wRPu2rwRAIzgJWlbsvLbKx0W39iCo2WEBaXQ7Wz2YRj/GSRc6XJ1Iy9DMIfr
joJ2t5jp7gyYFLmF3uU5rG2wlkvWWyGOSjALpsac8PjqydVa817REZ7T2RfP
E5zEWySDHfIguSfCpTxsDnmFLejVhAmqdvi47HCUGAc0qE+xMw7tx0yT5uk4
UQFKX/VINob1PmxyK+nVCGLd7iYCDIi/NY0SllRVQElKvNQSoX23K/YmdeFt
1y7n6TX8H0tQxdpyxTgnvmOZF3Bry1w1mbQnPcMRBDi/yyKK4VcDzmGhCO4i
9jZjgjXD94KsS7IVy+nHxaB/FbzwSykgtjXb9eciUKUxsiNS3vuh6qSCX206
H6mYG85hYK8fzrd3YVpJ4E1QVtvKPiq1Okd8wesserTGv901dELuuQ3V23kC
qd7RoKDNvD1Fc3bC7REm9wbnU+kO/axG6cbS/7Z9HP0YBn5uOO5R8+UW59w4
twhQzxf/oEpmnr2XHcJzAGe3d7vKGA5/ngC5CLRBVKGAm96MgXi1rHH6HUDG
JwBvZugtpjbxEUt53Cwen+Mdf9KG0IEO73VVfI8HIoWCADPWHw80tvsl6Y1X
8vsIrRLa552tFctJilsT7lzBCl93f3BWy/Bw3ynNH2hqRUkpBAVtuNS4ZivR
rnKGV56GLYQR9bwjukCDAIw+i8emZe8649YR5JoOg0PwmAbe2I//HoptXfi0
SoUFwFsUzKG1MeKK15BRMSRJCuyZNvqq7vkEC2BHRsbx/f2taQ38k7ae/6Ok
2Q8Il4fLIczWgdlZTt/udGV+iZ5yOiwjmIwnJZrwi2pU7nPLd4rxNXvTQieQ
6qp76U6HmngVWBhKZcvUlgN9/muFAZHuiAtK96UxxxI5R7bKkEMhhjmYIAfx
A/iexcxzC3dmERKiSL1qg/7jxBdNetAw38iBPnIvdiu8N207yZCk8M4x2vEn
sbSHYcw2I5ldMeQVQ/CYW3G/1OhHq6P0Hh9sCmN0bcJCjBXbOgb8c9L9TsTX
W51GveCGD/CT5nLrOEgJ+q3otE1fX19ssqudgKqjpqnFNggB36jnUWu3jEE9
TldLqCzrVn/eGRTnDPe0sHnPZrhOkxeuz/BYoPuH7aywj6XUxc6yryDDMmLI
IPvYpKbPcOrOcLE/bKgixHmtr+11emBF6damXvRVwAQKm2PFgac4+gSmivM4
dO5ErZtEnLLpS08OXWsPWAPQUM4U8AenAECh/DQ38H+oadpg75pFRnWwPjFy
N95/ei0gfIsRCJPlVCHzzxnWl1aNjpOucEKT9B4ayMZ6z1kyBCvqxT0+ZEv2
4pmhdGdCw742wC1N2wcbE2rbHh+OyD33IK0hljqhmUjqJCvI3+Ig8K/xKcbs
E3fPqROZarw5fHvxXBGK4/QvCuhQ52jgtWHxgHHtJ5mUL0MFwd24zhMJIdVf
3lDfuHRg20GqNXXEK88rxBBrdu1MRSfdp8c4WSbDepgrDgl5l2SRmGnhfL6B
rcCueP2hfMgDtlzK2/F0CaFdyhtYWvkFk3HAGRjmxo7R8Hxt17baw9o/qYP2
dOx2lK8mPDwfQWFENGATmvZa29ZYRlI3y5T097SlYNGbtTXTMlUo61pspGXS
tkeomkOoeOkE4I9bPKpCnJPNKiehubCdjtds1RYqE9LTCGdfKNp8oYdIApiK
fZrJnsnY2LNk+2zNAOIW9LD0vaRonLgbGcvwrwYsC2AtUN1Nw6mrmpv0a6+W
YG3QmEJ6i8F9SmirRzRmIv4c/t+ADcUqu6NlLl3eogkuZUsgEXRX/WlKHtxG
qMEgdXzmSi2uD8/6nw5ZlX2Rre7zgSXIr0+2RKcqknPyGnqdBB7jo8PwB2Wz
wkETszXCC+X9ikLkW5Ez9M5/X8eFv6bo5kaTDMSb/R44hKKMMFOOXqL+tFOY
IkJED8bTCD6+FAuy3sAZ5kDFb1Ijgx9aAQGsAWQhVuWIVFmRuGigGdjgCHjK
1fyxXJfD/apfcIRRVs1sJfMn/lDj7Jx3GQL4mlmSke8NwI7FWWxS/IFfGKn/
SVVekqqRL17glvAEbFSL33uxyP+jOvQAJvkSHTT/hay/2bcXEp7OQ+JkJGz8
6r0/Aa0R/YVQWbGAz42suP8J/e8V1PrIsaoEG1f5F34ZNizTipWBwrdTddcB
0jeLVa+NZhPY1KX2w7TgKhBlBThxZNCz454u8Uoqzl6KRjWUmJk6zLLcublH
Gw+SDs2bEr3FKBt8kJtXwWlr17uqQFXgWnkGvn1x78jBC6FolYpFiCo4oc8r
7dOj89hgHuga14R9Z4I63KAlrINAmTJsgz7XlThIwtXKYEWPsPULIcQ6VmNd
TwdptIMZk8c3/Di00VwyitnKkYJpt9Yl6t4AGfDyeC4t91CYIU85ZJ24dARi
hqBgvjsHSF2CRRmULsbJnfrS5nHFwG9kcmoVBcT+NyYZk/4Xf5o79VHkkJca
VJRvRFyhyPWF8lN55Zvbjgq1R98yPD0A1DW1EHsSmL2z6AyOHZGzQSLD4dl1
x4XYrETx5qWVlELk9tjavPS3AujMZCV6VHajcatmbRk08BaJ/LfRW1vaZ7SW
0lR9BMqbYYYNkttTZtZt7aknxSAFG8qrvxXvKKcyz20VEVCeQL+WrRljs//A
yiq7cF354ENWWIuLv3vIxxyqyYn6guJQ5ktzBT++drHxSE2Qq3mKlr25WQWr
CZCcBVQdHcDaYcW5fqEWuPchJscXLiPNljDitWnBKRHDGnFuR0e2eXkOnckO
/tLnlRPcn+pp/riVa6YoYUUegd+H9+V1IkoXh+eQU8WsOSvHoFW6XaZ8ngRg
DMhWUBUlHk+flmHALgdDMalW5jkLaIajVrMKIK4BObh0rYSkWbuxZlzhtiPy
BzAp8udvUVFI14DzL2jusoYP/lmppXkKpmiNfn/wxSLy4CcHZ+dsouOsFh1/
+yRg/5p/L3hK1oW8ilBjOL9UpkwRZrRPFaSM0iQOHWYr0NX1sta5Sl/cN90U
BLgnMZkCVAYqBaxMiNKb7kEpHIrj/ns7epOCDJrbpHKIpavnrfQ9pJXKfcxq
JAqAUS94Hgx+jyIK5SojV+N+UDUYZCSCs3oV4uu4oHRdPjwk1AdbIkkvPB5Q
A8S6oiiQ4leJfU7VHiTU5hesS0P+6DPvCZdN//2y/NJ0XWl7g7ubXDIpUww2
uUELBC2QSfbsRvsEcAudsHFLpgJkiATlqkMmjuwmcTP3bbgvW4zOrNJF4GWz
hZLUXXvGmuniA87hzbXwZLhtF+7yZXh6MCSX++HkKUyfwlcQOxWVTuIsols/
ffiPA44VjJJl+8D6EQre3fSUB6uR9rGQnDtY16y9O5zJJUPsq5HLeGVmf7PO
IeNvWxRdDZ6D8ev1fn4lavVcCpOfKpyG969Gz+qZuCSdVhAWyvfFi96C3l9q
b85yjm649wD6yoCsBuwH85zxigczPCjm34ATZN8p5VZei2Q7QVVDmtAiWAoD
RgFFRZhCTK7PJ5mUs0Kt6SXVWOti45z4eXeSextHvgcMqE/n+Me1scvBJyt/
p1JMiLwRNJRORLo/QqeXnMM09vdBhqmgVPY8RZ1HdoXE+9cGbfLL8cN+QKDr
BpFnToOL3+XBKVg1XX86wiiBWK/nuySd13neVvwpUmZvEDkpKscabmkHZnYF
XSAKZuvpkAPHWE0FPK//04j7udG5yc6eWE/Y3XkPyNTRzO/nZ1C78ry8Mb0G
FKR9I3UWGOwEfwtLQ5TIrwuZAEQC9WIR/D4ROiRVsS0CCQmQVP3G/1cYNdQJ
gnrLLW0Guy0lmwHtaD8G1pImMWag5L2qFvUkyLibMR/xmNvz1itLRbbsAseQ
wp9zdr5l8FdibKmB6sfU0hQdHqRB1CchQUBCxH4HV+kfQWV9h1UH67LqgC+p
zzzads9XkzV+QHrWqd8xcLMFu9kqsj1WDIr6Z9jK+sFffmiLGVscpesuvptb
LCjt51Hs646gzZxJC+5uHR6C6yNtIVES476iGwYWuuTcFG7wKjTo8rSBMH4h
vNSOVD7vVmsbduz4Jd95szr7Pxn0gJzExxlT1cm246KXhr81eTf0PbYXYghA
dsVg4JgsRrJZM3X/6SgoKHs/jQJeXJbqh6u135z8CTdUST+JqsstLHQyQvix
tnfpCuWDK/PUzjlRotykcV6b8EBnWDg/O8VfOiiFwzAoz9mSiKpCJH2F+FJp
GBxLaVZX48oBH0PeexzPSxRm6nJXszgoKeu3kE1szFAa1z+u3qvMShsvA2MI
vbj8jsYTmDq2b7Vw8aQidEgAPk4ixb5Hh3x3iCD8YL+Uza1oTE7YCBjjmyCt
oLkD4Z92LbniypKaT68SYaL+VE17UvpdUnT5T3Yx8VlsGVpbzyqCT9vNQ6hV
QKj4KwI5mWyWaFaW1zMc36/rTWFLV1XwZmiQVihB5SeJqfBh+ymY7XiwyNmd
BQzLtFX249InqkID1/O3LS1Rf5jXfZd7W1a0oq6/GOKqZ3hmdlYTrC6ngiRE
P8icYnuaOJ7M3w1pQujU2VH9miq0Q/48DNSE64+QHpECogtW4Vnbrbnl9afe
3ojcpIQz1Oe+OouymPjOyk2qqwViONcRXrUA5ISUQ7nklEpYKYoK11HlDCYw
vSZHCQ0cIyvpD86aE93IvlyKCZl5TRKvZVD0g6rxevQGdW2lxHLYrSL/fSlt
AEifiWuRU6xKeFYYfMTe/DekeOUF9uvX608jqVi97gcuSy9NVd3F/vKXLE9v
MTxQXA60j0QBGq0NGZyDld51kxghekfIC8snIjDWHkoYz6zQ/M6rrAEwkY5D
74ceRRd5+noQw1GrBvk9mM7clW5Ldy/PlN8CfBqndUlzGJtpQK0+OovEPxlz
hH6KUZpYlWnOQw7MYpgPtphv/2T7XMIZ646H2q6em13X/BPMX0RSXlP1xEAk
81fxi3/BArf9UcGbq92kf9tSjViG5viZI0zHrYCKk/VCJw+obZRZiquEumSc
sbCL6oW8elTiv3+SkwFZLU0MGgiKxXQ8M/inv3OfqOecZPBgeYUxU13MoF8E
rhKoXAqE/na/hbCv8SFW8kvgFNv6nHcy7a9kx5Q689udmLtJLVjc5q7B7NCc
8q6oES298b9TFvJHdhsOG0EqWSgyVF6DjpchQH++rhHYgq9rPoftKEj52bsY
jmVokKnVS7FF/m+4ireyztX5QPjVtqEBfi2Fqhg7BqmWhB9sxzF9EKjLR+IQ
BWF7rObWexMIuEgN8jdMAPp0lHtaonGszFXqqojXdmUmfcVWlo+NU5sXL+Ef
42Q+vjf6b3tD3dvj0FYSIvTrAw5xGKA6VUb9u/WFnUsygiwCscVGXdrSEnOK
zYBQKlEjavDGE+7Oe1z9lEd2hWj188JFlnu6ZHirlOAIbVw3JeXlTufZ2w0K
YjF74GkKPm4XE5Cj8mDQMkVWOMMukxpPLpEeJMYjulrxGEGMq8XVkt0PrJe6
GbFHkt/8oDQ+sAEEJWA/KBDRSfRu+qxoPJdJVbTHF8ayhqCquUMP6kdvYfrD
kuI5gx0tqhe2CYUw0oEdFpAfGF6cjTUe3HiYg0hSfe91o58ZI1l5uXG0X7TS
0sGcOjHH6Le/qI6maf6NN0YShMkx+D3iPB+ttMpzqerjjjSP9QZZ+YROMkLh
uwwpTPVmJ8taUyhp2B5bpf/iUMXh2es/HKBSc4Zh0uicrhUU4mGMmNsDvh1E
6wHRL7cOvHNrryaNwTfs5oQY34UX9WWThrRwWWHb2eCSTLGasvRC7VizoVye
mmsSS0tX7cFAGXh2fsWMFJD5fR9L7xPPJnr6Q7kOqLBVrF/LSLNmLQFAUF+y
7IPj2QzdbeXAk8ytOjTzAyf5pRpysHWrLGtLNs/yqHrgmPah11oIAknvCONc
i212CWewoOtAzHH0PPA68EImltgsJ7reipTEeM2T5dZhyp6xtdfzF+/UM1Qs
/A2A6aODL9hOjscn9ogOho7IL4tpuqSE4zrXJI9zfJh478BHJBeeDNu83xse
x8NQONYJNlT+aMzpSvxbOL7Yau3t1PrtQGaQfMENgfF397xJDq2QcH5Eiiu2
UGU3QIsjwDKpW5eUReRVeoot2N35ddQnnURfH/+RMWjM+DD7gqINsxR4TrMX
7agFMHOA1UIcgb/eeBtUx6PJ7ivPNuBr6TSKhwka4tBs61J7/T3HsJvLfl9w
09HGI2b0mABWHwLBSYa/POpK5sMUD8NfTfNkUWAA9eJX+241NrbyC0p6Gu4S
tEwmUp169i7+5s54/a4a07mFloa3B4CNCoypKRTF61NYDnJRP37XTEEso9cv
tBYJ86kxVwvr4+EUlWzci0z7Svx4iqgdEFCW9vfVe9JZUQJuLK9bdOXu0wDZ
N3/VLm0n/Q++x4LLVk1WYWJB01W4xYvX9E2APmL7crdgHWARW2OjY1xMw/al
I0PSR39nRpnLZ0qaZpSyw+GAsX/gNcEQ5D3b6NLNIvorbSAxctefwtA2dlJE
Bn2Xc49fudOxWTGq1GtBFufUhZ+N3c27GKHTL3Lml5+uo2cOBEojPtxmHGfM
a4UN8wXVL/Uz/mTqfO+NF4MCi/dQ8bsG4HyeV0nAhsTWbYWXDtSQh6uJupsv
aFPqmW9IhnSAjgvQqSf74gOJyDV7Gr1pgEcI+UAVmBL5Q8Kyo1EubVqjQK/U
+W1CXYnl0u2MXXxkLACW+VGgrY80OjF/eIJQrJPpYB6FO5k/YelPjbaa/JLN
XGiG6FDKYPWTIW7FysBMsSyKAexv5F33s6zSfVV3VoGcrh6pF75/eF6SCLuJ
n3Px74OPwtqDIUoL9YIFJ+xiV+v6O/jH6YfQ9XpIYSRvZby2hyNngG0cuVKY
CW6nOOzq8GGaXPs5eapp5dbj0QsCFCqZnhBzRCphyJ9eSOC7QbkLR8GBIEN0
CYsyzVbSNOjPwnvujfRfqnBWui2jlfYMg5H/si9zmndNGDCtvVt39QPk75ih
iye3gyT2UtGrzVNrnkYbY7LU9AdYyTSnff/ZkOYHd01dW3+q0o1YIZJfgz9P
fRp+Lx45EluJDz9VRukS46bQyZuV7ke4cA8Mf9F+HyU92yRveESAMkrbP8Tr
xP2E3UoW6Fvhz2XdGcByQY16Y2/N0dNWC6GmmYuAUNkRtlFtLUV5wOEJKw+N
pyCL7QyaYKeS0oho6O7Nk5hE760NYp3YmUfWeebyTjz4jlo64HWurohVIJ/M
SdqMGvVfnsZZW0rJdfrCmidBst4q0nfD1el4GN0psOZv668MiY1y4PPQo64q
RpE3mWgVN65Xkd/rhoFrAUc30NvyI2R5k5ZbNo5CEkAgbFOvZSTWFkiS7kFf
hoLOcwS0wPWvVV/wftrt0CcOdirXh/Jkmt4cxYLixt2dVnRnWr5Ho9U1GJ+1
DHZehbvs2jLEpfFlmpWWcyW2oj+4wl8iNLA4Sx7Zr0KJTUGiX9dCLlQDCS0i
7hqOjeMoYmW+6F6DNGx0IdzsM93P2+/euDvF47pNuoM1RPFCQucPaHfDx61O
e1YK+VhLftkeaF5EwYkq8IvF8EGa1J3pRfvAtG+soa+no4YGwhAeUW1yBIaj
po7I3aBz/IwMez1nkKAInOQJwjsdDOTdb8huj+heVe3LVqlvQtss/IOKHb5J
VsVsiFtj7px8NeVu+EJUFUpdIRY2GIzx/mtwwjoxR3usVOgveSsJD/nMJT/N
WIR67FcfvMAQhzcmy+edSliYWUBZzW181n1jkSrFwfqJlL3jPl32qvgb0EW3
fjlMpmt/6JnSCn7TKkK+oIvLYZh67PmJOVEGTAtnFR/EwRNzsQOokmzOPq/K
avR4qMP+OA+Mk5ymbV1BUhYFBIT1NCHoiLlVW5JBfI0hNqRpFx4krvVlly01
iR5l2BpFW27AIjv8F9yb3W3YOsbuw9XxFNr/zxKW0p0wPUPly1dq1VXfI53v
cQASQSjSmMPaBHejV3Jb3QAwRfZPw2d6fczRx03iYxD24DofH1gsJ+QKS1C8
BJZvwg+47Qtskg7YCaWLYcFBDA4FZBerfAbkg7J7OPcs2vd5u9t9gq/4dJJB
Aqh6p51q+XuTXo1Ty5o1JV6gMfbQLdHzQC3mEKQownPmM3HcZuDdF+QSHc3Y
D3MFxS1prFmZ80G27BQgfLTiHaoEM/WmfHAGlGKzjzIhIJ0XoGeX4iha5r3f
nwkJzOXYM3gHfhRrAjmmhihcvliXRPx2FJgd+003hhZZd8zUoYGJVk8yCVoi
91qcdDx6cyTz2CiOV07aNTJZw7GYc35F64XvhxY9QLKt0D/eaAsZeKvp51/v
p2ssuH0BfMKecuNFcLj+Sr5fiLOtrIvRghd27bKmSKjlzzsIgiLtS0lxEhZu
Zqv10jO+wr9/cSis8iPTwGBYV06DDgpOniQnExnHymYK7NUkYkp3rHSYCOz+
RdGoTbcDuMhsT90dnALQUfZNZZeBJzOgeXhmwJ92ZaQIbzhjuOx7yrtoBK8Y
KFtPpm1qCl6m+ZTntv/x/iS4p3Hcz1xHNBVIzCQs2zFCSCzeg+ZXF+KRhIkq
bSTCVsdL8DB5RR653upiNNe4bMDvlKlMYccuzafuRwiOeOjUyj4kreLIGHvP
0AzUZHp1+ZrU+hX9fP7Rqyru7+2uwJdjKSJiwma89BLdQxV3X+qcGinqalCk
r11RCWeqQsiuB+BUkH87W9hc4xqskeajiXZtYMq0P7y6bWynx0T2Yy/2z3su
svUWUfs4c3BWFGW6ocvJUPwVutp08idXYQqjYdye53UbFNC+0huou2aJ6cjp
k4uBWP61IWiPw8dIbfee6amz/UdQnq2kV3WPAaEYTTd1Z8vqJFf1Ep8XqeEm
z5RUyL/ztk78C5Gihr+h1rNPUowpGyAfuL2h3UaxvOwPPrZgOBJ3bnduv9cT
Gk4i3XwTDiF0rPRM/n3EH+EO6sRmTPmBDMr8d9ztf/lPjX7ZC7QB4Tyt15Q7
CAvLQsyQRVb958pNngxDpUXNTI4G2Hp24rj7gC2mHRRNLQYC4IXwW+fUbFZr
XRuPQrEkyT+bh3V12phZyJrP9DJMboUaqE41GCkdpV3wJPqmrjJXAXzfSV4r
G6SYhnJJrrNzTpwteywa94KIq+QP3WEbzK5jkpVC3lsxidpC2nhYjktxB6RK
UknFot2p5l/jyO6qs17wJ2OyAI3hY8DJyVimJz5KngK1epVe6M9bRsw8WGPN
Fxcif3/sjSgMaxUX5QAa+rZiomd9M5paf0MmXTfMCVBx1lcVA9EUjFby7CM6
03sHXf4Ta0XX1q4c4Fj71CC7dJHFAuehCZaXXMHQ+/5KydiBOm3Zuc8A7Jhd
QEiXhqpkKiwqxiD9bDZDqAs3t/Kxy27xUH2TgmIhKUWWAb92m/ircnRmpQH6
sA3fI+HVU4+QCmKL7u39UdWMJYm/0Pc7UReqFh412Yq1431851Q5xb9/+KyL
OHlIhfwvqwnCbc/a2mI8GohMWxJwQsCyBypITBCPZmxXqvX8aWz3/uf3F5Dk
JF7HKTZcpjdLgok1GarfQFKvXTU/v5aUwc1q5Ag0V5s85hbl6Ldh8qG6t+hG
ctU7LiNFAt+BHIH7ELYQulmuavmnVTF2yjMH9o2YIQg4r1XNbrhYcuTmFeUN
WJ/72GXXxuGApxlUWJ/duDlYzK8v972W2+i9w32pWaTVWk+Cmg9TooM7I23A
eoeRCCbzCQ/jos+bN6SDWTtYQ3elmu4lDG6uu2KFBfCSHJhw+rjrWKsqHNQi
9BHvMicI0hXZS2TT1HSByzjBpSPzsX4/Uff+7hAa5HroJrBVKwBT59R3Woj/
ip7YhhtaCIc0Mmpj8Ej6Yez19PMkYATwkZOxueew0q7dxaiy9oh3eioCWiB4
WTEhq3LPOmNgJOD/bexy+zdgY1LbgJjcI8IgdabwMba6zDFPGLueZKdii55G
4aTtS/EP4Pk3rnTj/um9Z1cNppJRlg9pbDQi3WqX6UOlPpu78WJfCUiFH1cT
1zq0Rd8N/QxXmm89mEMobhLvg7VJA1db5jguy3qa+XI3DHNyI7ETKk88KInF
kyFTWvAFl0OpXIxB/gATP1fMAMCRz3xdl7ClMoEjILxqOU0XEpJ8jAQCQ6mo
gcA20XS9U2k0ySRykOGGUHKKI7nOoIYU5EInPlQzTXM9HPIm0cIadNxcVx73
fwsdPPeXxj6Kw5JHI834WMwRFx8fjd+Uhjo+N5hEyyo2mY309E0wA1F8ecLM
qGFzocV4FvP5HEqqt3oeFWBenp/Sdcj51usCIFTrmJ7uqTaoLHwDLMrOu+/c
rLdislfaR5LZ6fxPesqoypJLN+DqWKxA3s4V9kD7c4a1IVaFaGWrNuK9nrUk
5gejOJwzjIZWAjklHscMBQYjUTHop/8hG3DzlG+948oreTU164Rji/lvTLHm
Wz8Y8OrM5m+YASihUNkwRqocObDiIQlTiHK6Q3JV/hzLtTZBB9aUPnvO7atg
Kcj2WEe3HeQjFdiDsuOVX98Mmz9AE0tnSnPlw1v+CpRJ1bsFCdg3rU6aNx4F
J1r2ldNjTd6wiO6NwSi1zeQtx7BMRNZfb4S7GGivqQsA6TN6jKZzcCQx4dcN
c/JXQgBvzGjnsvutQRAiqa2zYgr8j/eat69w2Ta+aVKs3ceX0iUNCMVmx6jF
fnJoCIvQSfrgD4pNJ+jgDlMYrW2UARhGWIk9AfmxaG8vVQ8QPVwYtsjUX+JD
lSjdyFBTB27s0psyzlgkWirOhPpqEQmDBEvnxDP3gb07b74XUNrcBQbURhEh
QzOonw2h9oujPPO++Cohrr7ajrtLdq4GOGhDu/Nk4P7mh2uiT+Ji4aCQvrHN
uuXAAwu741wD3oRHJQcOijuelKDTyvjJONhnU026hzmPDJmgJm5M8kDfZGE3
uT4hkLI5pN6UundYlec8IxFM5BakC8LhYaWipEm+03sjBx8y4fmGxnUSH0Xm
/SaEKptc3cFIfD43Rs3eb+N5pInKt5bfdTVtM4qXVKiu3374JbG/AHRyG/qg
bzqjpN+acilRvuzA6w1DsDew84yyUm6qR5zEQydWMALmJ11YiV6gWBwRSNC0
x0jFrGQ2ar4rVOEIz6RBhy1irR/H0myPbGv5I3teF4eNryqHiK1wKiTI6cQg
oqAi8zVuPaCN7Vu1frc7KriVBkGnS+ljdiu4G+gucUBKUy7E46MiMqetgFvQ
YOAc0bKvTgdXVOPALMb+MceaJlt3IIVx2tdaT7WI3AQwBdec9Dx85ds1MXwH
XzxxV6ImCbBAqgRdXl43uyqD30T0G5QWk3Ofo/LPYPGsmgxy1E7STlCS3uUC
zXfzzZ7Cs82jlDCIaKeO7iTrMjHj1+K0iiFAE4v9AZ0WfyvRhiu4dDRXsnY7
VhHWoGWWNyQDNjrZC/fJnMFQYgWKthKf6O/cbJ5lAr2+YJ7XPJeumzZ5ZfQb
dmlgFBXg8+q7L2oWmE94j+4MCYJ6aDRAebmrzGh3rKa2ExzXizoRhuKXHxWo
Ar9qOc6YSPLAqiyXK8TgHAmbWDPfMbdjXCnZH2DjxrlMZxxmUM0Nek0AVEMk
hWltbqfhLsVOABHV2DZwnCEjrGRcUknbatR3qxshDO/cm9HXUGtclxrceUF8
cfpLX9vBY6xku05OMYZnSIppgstSoHvoPayGM4Wu/xawNC6SEaBgcdi8fOZB
4r6JtGCQuqwLBQBN6bcMk7vA5qxX+qRVPho0hKgoh9sTWe8e3ALOMQuiyEC3
DELbxhTePuxoTQpWt3qOtbIS4uGeGpjcC4zRGx3FfTh55KpPiiIIeMBmHUHE
5vxTrpS1RXKGkxOBYBv7ZhTDa2jzul0Z+2CXS5ufL8JM9aVCGnKi739S4n0c
TK2ZjxJEm6igPjdh0CSYwXfeT5Bcm2eohpPZMEd9kVWl/lIeeio/IUSHDXP4
kZb4EsAHaITotuuZ4YSnJaRFacm61l1vdgHd/7bOMcnPZmmlXBbmyQr5WPPP
Ka4LkWcO9AeNDz+r6feNdLXemfterelXy/KjxEPKd/17s7An2YkoC7uSJYlG
1y4IVmaxmFuA+rekztryuctLwzNM3OAysIwZ6mN5Vj+NSBxneqCPkSc2gEf+
gwIXlPHOvHmr5rRmjK6y+17lloJ5Kzgvf4iVvKMHOeBXwHH1uVZLA6ulvP3a
gc68/4HhjwdcgfU3Xd8hgb/rgIvNnntnTID7I3+cDMl1LtA9ixrhE/HtAPjj
1mMvmpSo1YgGSyM6WDNwYnulE/HRLpFU0YQOQqyQi5sRT6wAkPe9b7PX7d6O
xJDMA7M66jf8UxgCogBeJS6eCVJyPoF+shR4XGqaUuq03gPa1rDpVOiYcC6T
I0QY+8BCnpsSZbfTS5qGpgqgmSL/pJueG6GpVRFpw6R3rlCn5eWsiED+biC7
OT1YvB/7YCTAMsARg6rvX/ZBCuXJ61Foj3MmtFpzCouvkKn7sJcveyMX4g+z
Kz0FL9tpXRs3sZZNyE/8KcHWsuAXbHLazMphCw3vwwAXVKiJOWZaJbVajdSD
CDmTs0VG3GzjH0NtzV9CyKW7EpTCAKC3s8Chg5c1BQQZPdGBjDlB1Pi4l4q1
ZlEK3+R28PgPuLWXWuPJkXjCnwY8eYLWps2igAfUOLV+W7x/XBIJ5xi5qWPT
xTJePR+aXkq9yiKZm6lk8TcbPe2prHeqxDSR7XKEM7+oISxXx02zqEnZyWuM
H336AFwEcQhEqRXOzY0se8FnWeRybFd5ZRZXLhKD+E8+hGuQ/+4emF5ZqsUU
oWFg94ehFqLoULQUU6lyt5zcDtUG0fr0Bd8zlE7vC+GERQ1wCvM/C2RQNCnb
pz24+JKV0LV+t+dRToTF1Dy/4j3ziJNFyQIcHUrI9iTp7rx/nNV6iKkmKitz
XKE+CqjlroR0LDoNGC5LSZ5zPP6W/QhFJpzoxztj2MiEQj3FmgcIcl3dsPPC
Z1fRzDXfnLpDwmj6Kj+E2+4lqmBlAcGNlBfnBbthua/99lHq+89VyyCcUh9p
L3aRzr2zblL4+CHCUl0YDnasI7/BmLenvOVsimO84CNkWuYgH0CLaIdziJMG
FUtKRNAQq2rdfYsI5YipPgbsF/nazVxx9vkZq3jGDX3zB4ohJ9vqrTcmIO7w
DDEO4PdzHGlYGbh8RfgTirKWlF6w1NJbMnoOxK0Q/9svtnrytvkK889nA/b8
7xLfp3CmQPjjH6oO5klR8Nv/rvXeRH6P8p/EqO8vhv4Ej+yRTsmUpVmY8Y1/
CyQhrwK439ypLdkxnpdAcLrbmecwUZyAO0rUvwXtQdsvf34wCNT5UrHatV1B
LGbdHVTscyV61NMGEn8CnmAUFl9/J5XVPmbThbbMoZKVzB/FC7PUhmG7vRxc
E799/RxCMWXbdoFVScI6XDDFSuP3L8mSbEn5qTLoba/y7LYVuXoI73wC1Vt/
bDMzluHzNMuscNYEYqnVQJs69KwuQrqUlTn/gMLjFN0ltLglrcWT4klyLJsy
ULYwcdTV68IVRpg7xP6z2eIdmikrAh5xlbJOoi9BP6YtvKT1XX3kKDjSAkI6
DmkpUUiFiINPi/e15WXMAvwmw+4Tti3Um5OvqwK/pkfbbrqf3MOpoBUXhkSi
jOBnYxFkyTE9pJeK5ddO/rIsiBqll0kE8Tb3DT8XaMaCGxQtpdSrIBB9lHSA
w36cLDTAQ4lSkNYy9M0HgBUds1fM2ljtt873NlNr10mHTQ+IlbVQlC4yN27k
+TikH1Q87CutX+yjyGNtwN9VnfuLq4CRtMaEX6kNcAKyYMhk4bwcFLjlzAjr
qPtFA0YxpAoTN6ZBaVDaVPVwm6l7IyordK54y+p0JnYqbdpx6Qy1I1SMr47n
Vyk7WVmqd41w3vqjXnaMHSgrLYNslFKwz3uVK/KZJdlD+IwuEbRufjg24n5V
BHRwdKgufo0O/NeuHiRRJXN9pyZdgYytlmBPlDwouFsihVcYuOzhwKZoobKU
yKZyHJ6J65nSzLYKsNvHWWjwMtQPIAgMRviF1NH4NP7T9tFZMep/9+Rstyng
uH/PjVJnoHFyoZhTOF5+9cGZhTb/yCkKpcJLlr4YNp51vqqv15VAlovNwWVy
Cbu4d5Xd3ySUNInUjtcRHkOzNMWynVPl4F8YGV7BzmauUa3iHyhzEf++mO3d
tu8SR3tCs6g0CPF2HpucwhUi7w477NiDcSAjsFw2TGlutmdQVMCvi9MdiljV
htTU4QNsRvJp5DLwn3WXqu5iXGgBjrbdvWN4z7oys+yAvo9x2cVf0mxMX47B
jI52ed+CIH/lKl9CFWdnItyqWTEof/IIChC9UeLw9nc6VLZ6sKbnewghJAu5
pnlhP6IwvlZiln3H0eODyqu6JXyDS5nO+S+FURnzf4rLZjXy1EYsJTE+EwcZ
OMfTmhD+DImGydcbv3kcz+nRs37euhjRhm5NMNPFuRTlg1Pa5+o01X/0OsVN
nBMaELQJomut6BViD1felYdPY1rwTcmPrrVt6gfmbcr6Hv7JBasqGOqZJaYx
YUdnAmYGzoqAP62Wf5Nw+7/aotWQ3yLPvtWszpP5xIShxo6rM2+FRYnyvzli
R9eU4gCXvqQSP8Lx097hNaQ4S/SfLMvL5ehutJInh8UjWlpJu3a3zrtUypyh
ek+slfTA7PN4U4IMqbtnDqFSMBFTw3Kf/wjW+YgeOnatiTCiVm2SofOhG0jX
6VVi1Rr7kckJWQI9culkfHLF7kCLx7FbC+fGUyH7WECWyEpY9WQzA1caL2ZV
MuLSeimED4L9l5Qu4nPWtNWxM9oJY17MDZZhwdZRAboa9Vt6w6DTCxzpFS/y
isn3CyXZdiimUIYLMjOVmAOPZbZMUEhiRrfxlIin8V0KwQrvPReNilE6/+BT
yEESM5BijtoJhaOOG+gTSa3N1z8DHwWSTIyEWDNfS4sOW0pTaWXmilI9cK28
JEm1mFo3ZLK92l6pnZqwk13wSkz6XS4KIWAC7EXZZ+Z8NSzIyDZ+S5AjxuQI
zs68rZqlLCC63PchhvOzTEddPWHE5UW07TNBbULnDBqeua3rQk5R9tRdj7fb
Zg52RljhQVs2UygtiGsCuqZPFlqWCUfZ8Kqu52z7E6gE+HNWiB4YGqgJwItt
WJuoaFAFxir/xfpUDHhTYRMktiS3cafg6iRiH0ga5epadYl4hWN9dEZNwDO5
B5Rjy9RdzFXEFTYk4WaOh/aI5m9zHg58qiQtJsixZgLhYlcitqdei8ZrwVTP
o5XtOxrYQPwCT6Y2eonoaL596lXZVa9Su+zjWoIrsKc+9TTu0eGtOdb0Vrgo
mf+s0IYdizjr7VS2ZVrWpPcOtw9GhLp6Om96wDMuldOM7TcDtGaLjUuP7dvE
bM4LH8htMU3Nk7rNVtBVdvbzjzjdTTGkyzI0c4AzKB7IkBOObH6QHA8x7Av0
RNNe9tQpNe0Fy0d4fqnM7Pkl039R8KpESX28b2gouRDxvtKbAfSeGFlcVwGe
hsPehv1OM+pcg/sJUMCTymASGEgihABmgjyb3177mC1TEEHDiV9WeLl60eYm
q1PqqMISCgJJuSf9pnVB+st+aoFbB3N/Wab7A+d3gxdD+UKzCd4xFvtLHfKM
XHBq0t1O8QGQm7UQ9TnNey6pa3oND68noO36d4vke3fk9/0gW091QhwURYjC
vH9MbKnIzyfM7Aw56W1D3X4OGpJdoXaXDah9YlTe3A8RBnnCTy0Eh1tKwGzU
ulz3ewYpV42vLxLTEZTUCJzz3wuabwSyDProKFR3VR9IR5oEIFOzC283eATz
SKJGP9bkzxoEDr6aswP/m1jE0fhzUR5TUU1QXu6tvTXAtWvoxujmDapZTUSr
PCMywdVVSt0nnb8Y/PeX/eYALUDM42Z38pZwELpUSrAVD9XiRw0rgqhyfO0A
31DUspTQyLKiCl3Y/m04KEivCBnmBFZK4rJCrSre78Js5bu+ws9QifT6sT5e
22j8yasaqW+qgkCC7eLu4xA0YoiKbtB3zvz6+mfnCvAspMEg+J6yIV0h+e3w
KOt7KTK0IxJ52QDl46YhlShUjQGCWSub/zmxjEal15tFik+tJIFAwf93Iuw5
VQMgPpdDHLp4DvsCbFcuHGK/GEtpx3lsnOT7sglbRszG0dOjpWyl0sL5yzpI
gW8eUG5BIlQJ/azgfXQ1XlWj+/xU+OrijOudRG1rXF8Hc9VmU5j5vVgoWod6
O6JOwiv6QJG+0SgThcdTEshqeZFgcyXX6g5md2fyiFF5mpeyS+gBM19Rb958
Ac95UnkYOFuVy8jkmWaNv9pD8p28etuSzWBXv9MG7pjiP2z48pqWwzglHXJx
61hV2nKGvxTYziZ1idbOIR9ORgzOIrwJDm7k62Z5SSgRgS49OyisSdwhql65
NYTjuXT1VfsryeLhBcNo/hvWQgLHm4mIqyAJZlYT3059xkLBTi/3Y5IDsVGs
J/ZUTch/WVHTlrxV8ZlEUJM6xGJ7oByDm/jQ3etuiZXRY/YYN4EhxAsi3Gij
aKwNGHhCN2fRdKTqxywKz5ZNgV+1XDjbrnCLmzWdenuJAjli7seqelCtduDi
Hm/RnZv4qWZL2rIdpNwMOofVrABqThqo7y5YAhfhUpFP0iYJ8cg/136BgeQU
sC3GPIoQHWirgJbl0df9P7BEwk7hrIC/DXJk6dyTmbDmlOPDeHvyME7rUmr9
rzmTMqydKm2rnxxzRLpv8imy456S2Rce2cxoglUXg10Am1Q/Z1AblpKy0JUX
3knfZ7ikPQowW3cm9DARfElu0jvQqE0w4NxlKzv7rW/7B54Gc1ZGfTJuuB2Q
HxdbUd7aCRhrjnj45oBj1hsasj8xJbojvzL5ntp44wTaR7FvXrXthJ96jUp0
503NVAZyac6I4y/C6QSYarFF3KKnAi6R1z/NLMVLn/hQTNGqa/8wbPJ8mkMr
rPJdIa5n6FEyPwZzcFRffx6OMc/Z6mGxSgtxsSGHFJRWhpW3d1XREep56BUI
7OgF8I7mOywIb2OKyZdnzBz4gQM9AoOjiiOL0eRV762K2AtAMj3+Jd3j+RbY
J8ErY8KKBYvQBuzNrmaUt8oqJM20RueEcI8x2v+rBgg41XPlkGYeItoYiGzm
XONbz8JjXUSrfUCbA5+SaalMccRtrtsyKDnqBN57xRvuKt9w46Z1yNpLX3eR
ZsUS3TfsphpXzg/6MUZGOHeDkvX8vYY6G95awECdi4ljaDMB/f4/12UHg5e+
R5Zm4+ui7lqQl8CurVcV34X7L8QNWb3pVvIk3ug8k08l3l8jDcWEIYBxBEtF
L0pPNX7ozFcXFwlo3ATx8YiUN8gHs82OrL1bbkavK6Va65qHIvzS4dES6VB3
RhwktqiSS/4tX6TM2kA6D5H+Uh3f8FEPgT4wBQLR5aYuKU5MZ/0dXAO5bNNq
FhqXtg3KQvNn0GL8F+Dl6T4cggvdxnNN9zAAffOHmC0gogmusVjK1LGp3lmW
ijIXC8A1kvFLJAL4yfDCckhq+WIuoakEQGixKFgCWbxZWZzj2T4Z7IiDEhDH
AZgpzk3PGd3a3ypWu9bQrk2pST9dWrwZ5CXtbY060EV4t7AnB1oVMCkvIgY/
wXj8xMgaqJScWhOOXdk2jgoMw2l9zSFJBRk/FJeW8plaQYU3oC8kkIwdj9Rj
RDgyYXBS18d+ddpRaeq6oTmRDQNy9fA/j62KIe0KdgOqX0aDypj5UE10lcjh
MK0DOlDUeTc8CVRf1e0u+acRfD4q9EyylHcJ2BXQwSdD1TXikmz+J+hx2zjR
sVeJwaX9KZWSbhLIm+PSrJFOXEKkQmkeyjZiHxUxBaIxftLCOuDdh1DIFAZB
vsZClnTdg7P42KNGqSLW337NPLO3LFaz9BuQgIQKehk2NZFDeJbRD3AiIpvX
xcUjcOIz+9v6/YzJPZV94A9EjRV9VmpIYnbFH6RtVbgWGUZ88zf2TnimStWX
M7rTv/XrEzhWEniNmFuzc8aQ/CaSeuXI9dA4jKd1az0XWp6Flhg2L4+xCJT3
9clEbvoPM+RhdDsQsAEELV6pUECWv4bS8Z35BdOw/cJw6vTU+DVQkHY4BA7z
UPNjcnHaxG9/gGpgkUIcsy/4vKx/Wyv+U5H8MCKfCukWQ5BTWVeB0nGDXIKI
GFabZZbNeP8eTrwXy15MrcJwzl0CzYdwNOZnIXsN/lYpge7Zv5MMvKU5M9y1
/4hD/0Y5lDInyXQku4g7qo27AYkxX56JPfRncFq16jQ8OdbNGfRpvznomNms
z/qMsIAwSiFjq9AjvtmDPjn1TKPeaKEht/MICwex3tD46JlQdFc2O8P5IROF
LNaepwx0/cHelRitea1Qzgbzj0UMlgApXPwEoMqKl5Hg2xPIn52pBGBpm4Yb
L45ju0FrTipzzE8tlKnQI3atxOteu7Ere1Z6ceexonxR7qDdg6FOtgEdaTXC
cAUaMmJTkuKQNIodVZ2OV2hMaU4O7bvhtJ1OpnsbV4sPEpFG1DUZM3C01jBA
VCaBb3ISjPthhp44RPqRouiOcwU0ne3Z65+f8thHFApqscDTKzYJ5Np9Yc1l
YPfgMl65Zl/Ui9vMCLW6yH3pKMrATuW5lAEGcJKk+OXHkiuieCzty71w+qGj
u8buTsIgbm7vF6D4QYdgU21YuVnnodMhVOxO0TFPQR3WD4BI74cbMsjJ3ARd
8op+6HfuwDeaDnlYRs+I4gCfp7mRkxe/t8OAoaTl7UqrF0xM+URNTRXhykyL
06WncP3EiAeY/7mpRvMNKMFZ1vOAkVZK0qFjwjgrpYGn034LwbJosfwUT+gA
mUYg8q2Q5seZ+eK40B7rcZFm02Qh2kzZD6deE5ZROLa21fQUIw+pcUL/jCW5
InwepLLtE6hrxNGsGBhzwpmerOHpd8/y38QoMxFfq9S2PctWQUegA3DGXnoO
usVKNZoI2yQJOCcbb4jlqrhn5mZIYxEYrFPGqnnedH6LH71RAmBLqCKyxUu5
frBDM41XHlC6Z3wcytf+RwDDUufz9BeiF5O/ltNp8IjM5SE9TBtTOzt2U+4P
CL72EFNfWE5IJzHUkgrr8k6IY4T1hUrcwqYpeG/uMESwiHSjyv1lnj6wAOWr
7nJKhdhTQre3bRS0danU8nHJd5mSRkwP/edhWAh8179uXhDmjToTUMc2uNLL
Wqx9RznlhRKPdzIeyUw1OGw6uxUOqZgh63Z3EA5I2zUMwtmUkv+dlq4k5yNA
OMxV/3dkF4xwAW+S4Bc+tVzWZnJ48ucbsWvSiGffUpuwxaxCZD5Cs19IV6/z
qa/rqVIhc0JxQP1ree1lPUxhIlzwd4gqh02FGOKSjRhzdvzMU9ZYsq1czlS9
fkSNHFGlFdcojbDeIT8jZQisgAxRheqzAexPGglz6zqwFC8ly2VsIxBWTbX2
QWTlXhWsGM/FiAZe39jFHqemH6SBIYMjS5UmRWrP+L2Q5Ms83KPsPiuwbL9i
G2i8o30OsQH5AQEiIXe2sZgkflMVtsPlahx04pYl9Q+RGzlRZusLRj889ETy
hV0k4q3V+A59PENWN86shtkfy+bjvaVf11+QXYMKKmRqSxCCmNtAcJn50Wbo
n7xV6gi47aZNgJWlUd2H1BrFYys/uxHKl/mJeI3fRZai+gvQk+leI1JlemlO
LD03ZpuPmpxj1bAci7msONOymgL+dGady9mgxWzjUhZAdZ1UCsGwpAKjW6tL
zQiCD23FmrAYEJfpRdexdWORHak7PgZkq0dhfN7S/1x1rD1v7VCpd16SjqBF
XNRuw0kLbfqgem09N0ED6W+3icUuQ7e/pBMRDZ6GBJfKBjfDgwh3oWpqpiOM
Hj3lsd7fAIT/kFQokYBIotG0z+19SvvmmboCD3+SqbXq921wRG9UFQ7ICijK
KfjH/xye2Yiv5rWt56ySvjsJAvNE6smMtKqk1JN3PKbaCGmkgzvn/+0fv1qE
TTxQTCod5z/AYhPIQ5YccMpyx1G4Cz0vgRS6TVnW3XILhvvLnut6KpAE8Kdk
fDC5gzIfUyrExpLwcWWbMEESFFjB7+54c9ZhXaXCCdiipzQTA8sy1S4ln5xR
f0CLlx9HHZeWMStPH4wk6zneZ4qSJZ/4ZO0m7RZ++tFxvCZt2+3KB8W/sYpm
dj95qS68aSoOvDpxTe5YiczAuE5b4rPc9JxIbAzsrH+Ob0XPsjURmQEdV1y8
0O2VDiIJVFKG2iG3mlfTmzbAs1iQGdsqhHCeZS9vH1izjN/YzGxYOCJcfcr0
xzPNk/eeHTxmYlqD9xz/AYHg9NP5247zvBw+nRwAgG0bK5lRvOHc2WBWuAjX
4JcCtyWp3N56j3nfDqxKiloa3L7tG4jYqDhf16jt9yRzrlzLeN4leFm2vMj2
nn7n6eXozjneC0DBg1xldxdT2bnEUfIYEgkhvlTlkUTcE9QQlnoJRquH6aL/
VZxtOWM4NJ9raGsdEAuBRqiG4yeMifuFYbHqZRtx3OOFLs1ZqQ74WjEbv1PE
mbdyut9COy27eQTcxO0bVo15IywZp5S5FlBWR32J17eybigu2vfhDv782BEM
ErYN077prhruoBZD0eqNwcgasaLOlgVApPfkXK3MsFkNrSHSJFamgtM6/t1u
t8j6IYwk3BpSz79lQUAKvaeolMTVa3vKers2+0PQeYUFNcpMcTtR99qdCMw8
+j5V71FwUgJ2Ke3Rb910WhOK0fuJ1/Mc5axQdxUL1L8a68ya8/OeFSw0OiTT
sXe/7jgfmNjlfd5gfPDlfj9VOYfZ2+TvyEZQYNHqo0acqf9NjQEl9ujVKSXn
a5ZHiiwyA3jzhio1/Qwdnrrt8+tdUnptwqfarl34zpHHiyiyn1VjnYgE0Qn5
j2O3mlda1dyr6j5hrw5DtaQpItda26OHXXPOKgU+0xVb8T1wTZLR3Wyob3/S
zoK/QLVU8rEFha/KyP6WUGVfREUpElP8Uf6fFMS8SVf2006taM0my5D5XXzf
muRKMUmFE2tMmgMtO+AqkjZF1TezDBxpAaS4LI5H7zy3hh9yvvzBfOUWOIIT
i3nGWg7WZAN0DmoAqCWNXXyeHexvAt5LXLkrqenMnb9WXh1mS3uKd4VHmrb9
zH5CQqvLJEXl1ROHMCDGsejCoFMwVs6OblULpPPtvjOgLiE3EA9lL1qlQhpI
BtwKhVwu8MgVPXV/GlGw5zFg6bpO+uRWoSX/qQNKtIfh68P294rs/5+KvBma
h+PZaJIiKYqeAlWDZwmhUmLKz49roxVpcbSSiMc2UTUsgFQnoXNkVgKCYqYK
gyt2c1REbUQVYlqoT+sUOW8lSpqkdAfiMNCgHXgHm7jspgSUhr0jYCjQOPAW
fGAGTzgBjiJ1juhYqjuTzC3KQfT3kEc9Ch8N5aEsOI3noz3Rmk14XQ5wgvol
C9Cq1hlzBqfwV9PK9rC0vlAWRLXoSACee+vpbhNyxL2g92V44MomRsOucyXa
u53TZsiXa3W7zeAYvAgqLZgqzZLovYPeyGlHwrgjO2OM2lRhK2m4fe7CfSZO
4ffDaB3tkMp7b2n5skDciysLlupVNW4U9Lav8UJ4BsQjdsxzWFVf29HDjnGd
JqkQt5jp2IY725VhCQqRQsnCjK+j7TXzt7/NrXv11WdFz6p1YIaEk1v8/3hL
3X+3eLO2bvdcANlZoqs/Y2GRryNPYzpPyAVhnDnUUFKRJUoAJfcl47ynEi2p
Go2C4GJSV7eZTiNJKS7TkMJox32PZbro93vaQC+ucPvjntzwRtt6wZuU11Lw
7amGbK9OOClwkfC7utjS80xdafN1AqzkwT0xW2+pVJvdcU7j06k8lDembooy
rMeUeK7YW5GS3dr9sstAss34I4vtGb+xMraK89WcZXvjqxQgeAbo1lyRA6+X
yX8tBkWKlBu2tvT+An5YrFKWLcfZtAu2cBwiic+bP+mh3ukJf7Sk+UOQnJdz
PcjJlw09XncTuEeLYrivX81cVwYKVdvuXMdT3CqGraQKHqsv787tImbXQCqh
Zlf/eQ2Vc/SYk83mn9opDZHAPRDmfRstONQu1lvKhHgkoNyLoMmjTIsZFu3V
Ju9/zmQGmh/etQC7X6o2+JsUUfGNbr/E/lsb2F27RWBKTI8DRloxIaUEyeZj
N/CCJ5vHdQY7B0QNriEPuAXJ0RvQNoN0eaDP8ew257XZPXo50VG1wAWem3Eo
Hb/vYWO1Dh+uFZ+UypZZftpp1MCNyVRPvoRhBpmpUtJ9Z/I0PjseSURNHgFN
OYFqXsW4+xpCtVqeCQ5vpb7bG0qq1o/1yCfFx1In6EPvKLiN1lEyYchFv2nT
AexpS7KzsRkkr4yDu7bLK82UvJH4luaLzHK6EdY59wwYOtGWGGtLP6A1GSDB
PjLuo/0S9uboX/gdxXIM8h2m/1nPdTsnyw2jZypPNddQeIK5V5O413Y8VK6k
lLgmT07wpbsyEUkCdYR1hkRIBlVWSdbgeMkD3jDYhSroYQQyS9SP/CZThPQd
JPaxSn8OqwaG+CoIfW4wZ5m+I4VZ2+FFMMIkXhC9Ot93x/1Z2a37AtNX83+Z
i8BojUVfwMoRdPGjF6PvIpArphMH9ly3YWLeLxr3V0XHZSldv+s7Fd9gQS9D
sqCV5f5LNrPRaLAW4b4tUBy+pehAXhYF173IDEJppGxUAhqRMfs80UK15HHg
WeTuyIX9rxJMA2R6NTbrFTrEgKMO7sfGl+BcuXS3q+4pkzllkvALumd5W3Zx
U/onHJmWdHbb8QsJ47zGRxZbOfiyiG+vuZnk34Vgc/yJZPJs2WwVg+aoyWIK
+6CazjxsdGT57MUk8VDRtWQ9W5P44zplfeVwmuSNqsf0QVbY4d8R3rh+BFaE
GH+kHCjj9KSNB3GhJYe45y2U7lOH0yQIFiu2KGjG91+F0suIZH0Rex1LEBZY
HVNNmsOZTD8kBAbcOKitut8I/NZFMqf3fyMmyFw2euZDpSza/zCya5a/j7+j
Xf+Y1dcO4AEHi7xJjK1rTO3DsaZCLbrQE7iXs4EqXt2tqB1gCZ4IyuYlqwDf
uGjFCtxfiloJqW1Ke9LDJY5hyZxM+KxX33F1b0tgDRq/5jsp3mbJ40yKh5xR
7bJR2zOruM1hsKtX8Q56onr8DsJY9ZT0l57blA6gRCeSQYxbwqMH97CY+mTU
FRegDf9U+V4POusMkh3V8FI5cUAKDo1w+ybxuK6FnGkx7gn7Waiv/9TQlT42
B2RQR1YlISYf5NzN+Nst5+Lykk7kfThK3pSRr3RD1ECRdKHET/vT4mwPBGlL
YDPW7e4n5grT9k1aN+Op02RzEEZnSe2jjRaYLO+EOktp8skimnxPFGcJzM2i
gQ/R405O7y/CJmm5/uYcICWfJQGedu6Ho6Sfb96fmvSMrDw84NRqNZu4uabZ
8Kxk4Sbv5bQqyVXpWwWLd7XGHaTn3hSyVKqNRk+3zExEOhFMbDtIQyqe9rAt
/N27CsAlx0kpcvqGduj0goGA7h3d8UWJxGAml2aP6OkphUGoaawP+3a0VACE
qBnhmsbVi+nTNiSZwGgCOAMLxCrm8LYSEHSlTGVC9Qd8oeRrYZqxROb65/iN
Yex32VBYhtLGX09LBEgsD6nAcRVPticKjSM0efWEyXuTFjOo3jaqeQBli9mA
nlKKYsdoN9Ej4Tfs4hsKU1A85PblJs//tLMygfsBjS+WrhSKh8S8qZNb8f+9
MJXDgaUb5OgOfwjuO2QIc6Nccp5e8Nn/vjNCCWcY5rydb0bSeloY1D1Tj0go
bu+Y+vm3s6a5wtaLHpf8foKF7Q/FreKJOsdAy47FdR/nlkNDSP2mK3AjqSqT
Ybv6fugHSqUsphxBXRj+wgYPXP/cVyNB3D7udV4E3Q5FHZEq0x2njPXfAS69
s9yVKm0us/5pz5fW1mvcyqhI52fZW4+ls5jAU3YNhZVTiPJWL5NpDQHaKqcu
VtaYlmHxquNf/MWNgMA0DP80I7sL/2zWCD21mmba1ury9qYYRo8r1ht/7J9N
5ow4TpREJIdenA5P0y7BRTzvP1dbDa61Xlv5W0yAX1tvY5CuI6yXcDbGRmu8
HX03ZZziHBT7aC2VvzQWXtWRkqLZZjQD4VYC2eqH+8Fbt+S/OSAc7OMQu5MN
z2Acy71ZvZ7+ODPwwqGRFl5eRXNrZWk+a/LllJ50F7p1pyqN/x+i9wzW3Grs
bNju3GI1GTM0sVprvR7R44UelBxSiEVqffOIUtMOA/g1bOYuR/S6Vgu9cjZp
SpMsV47AEXyq1gC2kcHifSOCJQZoWIgXixU16wq/TclHz75mf76oP9x69HGD
fS1wF8fBQT85fkIdZ+sVx5QJ0NQ70x/r87uJZoSZq4/tgsgPJXe4UYizF5h5
1Xsm8ucB9wXBxGOoOU6wJSx83TJr1xv7W+DRYdTw0LCiFWbpiQvmFhwMwenB
2ApQgpLH5M55XvwasGiXeqrwbYxeqsMLJgUfIc+7jXDGsyUMshT6VTX8Eagn
b5yMeywk9kQQsOwUPJd67/cD+hfoX9NnZ7B7dZ8xTj7NEOu5k8Th5gwXtGsu
ECNvbtAoaqwxpId71bnjh05hLIGyObnT6t2Lox4NhqGjx1mzgELoMgdIYFHl
8cNfHZnj3AB/tvcAjYShWNi8q/RXQE7oAOJxxe8ZpzqkOv+noKALwBIUp/6e
gjOaQ1w4PyjYErjxmWNjkZz6OiRJ9bA7Nxg5/NVmUb+1VWG4kyoxWcFPytS3
D8mkMHxb85Q5sljYm2Zloj+brZ0QNoXQRsOWeaTcxywVi8Rx+cUDqLXPBGmN
zyTE7XnBosO4DVrKxIwRNYfRHOHqW2YD33fJV0YoGvjjYt5xfT8+HNDrDT3C
LvMLO4J9iwVD2pbZ+vkZrH31dciLqdqNfOHQ8m9yiwYIx8eRjV1cmeryhupA
0UcrZiyvE1duQkiYsw1yQWzYBkG+k5HrTfh+CBwt9QR2bwnHPbasBe9RbvuP
OXwp6Q0Dd81eQffrxzPGqfwYyb7rYzTNVp6963bHaSqVJgMMaZR0rpBkVN41
LDFnTFqivTQwqVMf4B+ry61sJnG6gS7F+8KSWLvzbr16Q7SSsGHn9twU85GU
zOTq6MRf++BXrWNQOG4+c1g7cha2tL5VLGfeSVJH6c8cI+eWUZllUUFtB86a
X6cBBHu7ikALwZi7kfN7nMr5CxHnWJrrANF/J3B3FFO59kjHb7HCGb2unP9X
LKt4YojediMGk3eYyGBoNblsodh8XbGFtNx4XokCw46iZB5DwbPbh1rFUXFK
7F2FK5hvVuXdHI4NSLNJK/KeMzOsBV+h9k5WxuigZhMcYat1cBSWW2CL5Kx4
gQkpCKHVXL+cVe7v5B+eIw+R1BY7tpBlc6QubJrFq8myy5h0CllFArgRljwF
QRhr1CjyeQmcbwY2YU1GUf8juBVxKAdyuNRS7TiBFvAlfN8KeH/h4VybIw7b
HrXG666YlEElLgqjoL7gx04TwdlU/YKVYKoHc/UAG4jF/jHyxAUpiye+AQyx
gW6XIkw6t/18pNOKhqpE4sjL/mPajqghm+6Is5J6qmtfA+yBCRh58u8pyrnQ
ad5yiEz+Z45ecUHJijU/WjXrhzw/kih/j2VcL8vTQ3SQ139iRE49PiFNmQXC
G1njILEN2dn1Ro24NqAZuZV6JvFNcHuUPkzPpQAs6D1CA6IqOOO24g6VbJFW
pPDnuDHIO0OQqBUvMOzbu4T+YE8sXi5RR1AeSBTcda3lEduH71xol9aW8Ung
y5f3IfS5lK0xqM8vNl208SLQParU9ngD2YjgZ+dR7f3w9TYPusVn5SfGNAnm
1vMxqhTB9uk2H2das0ljo+J9/y+lBIey54zkCX5drhcKihboHYHk4hGABqN9
nPJYrpesdC5wcfd2qsmNuojSKExF5YTalcvzenGXZQIeaOxH70IqX1dpqqPT
DRO56JG5rqH1s58coWxBUY9ckHC2jKDuOtlTy9GJSTjdnEqDNBJrSiYZW+Dd
0eKuqzgANc6hQcpUhHMoE25NdCus7RKxq0vfFHpagaC4pjMSuPw+wtZOQ7CD
dX9C7L/LTR/Ofr2sBWgy1DUZlxXXDkroecleeRZvkxHPaq+L1jxj0qsz7SXB
Bh334MCNAFvfyNRsLehQZqRWOI8w17UOB5EUqLzoqe975pfrUbhTpRYrD6pF
71Q+l4vhXI6bgMDIY4QLBaS8MpNMPPH7PUhx7i5nc+jBzDnltx5q2769GRbJ
8IKIMF2H+sy02nnIfy5CCg4zpsqGtaAup1N0dMv3bPMLqaHvf/RXrR+4EUPr
SFw3CpCGjQ7fpYZ9L6tL+65zltvg8VtNi893sONvxoydgU4L6+DQaXAlGMin
Gcs9w2uWsebPs7idFkGrVA9bvnh4hOAYMekgvXpxOJJMRgcFRZABQ0OCWmyU
4SMPo9iGirkCli2i1QZCvBUX1XxHcEMmRLx6sr/0Wl/SkDKGCGs0wrHX3V8t
CN0fatN/0mTTt44h5uQjDQSOR3jBZEtSkKgrNtuiDAEBiq/+h03Q3oWGz+6y
rjhoQt4SFzH84CMjR3r+T3pICAGzEiZLfR08hBYMubxzyqYbtuUfaWVcx8Pt
HaB3yN+GbbXbuVGB038GcO1PQUebNkIFNBN2WEGXMU6YaQ1+F9tzSb1V1BrB
a6I7cHQbwCOrdFJIg2hjiNilsWCdQNWcmWrDrZmwU1FJfi/qvZZk1zRrVwcl
gMGW/2SntqbBh2bZ77w01S1HDv+JI1CjR2XzX31MlZyTUI5VVN3KUYXN2v6C
O4tuPwtdoZupdxrofbIn7ShG6OPO0gqsQCxR3CokvgkXHEMt69HdBnuhBy0j
ymIakDgf3LIS68QgG52muoxFAWeHn77EVOJMnjhDNcTVOPo2THIMTjpzD3BD
fyQiCmxBXOIQSziDuTk+iWr7VV1E4RZDQWi0PeXFWouK820cpFgPi1qGqttu
YyzAVrhDlpwaMNqX5b5rJO2Kvx3Bk5gVFxhC9SAIdPW8E7E9zCM0P+oJ5RWD
cLQigv1PyGDLHaq99lLLIUFRHDrCo952zXbwaZBoB0oSdceWopLOi8v280p9
IbRHfn9DKKYY7t9I0F6iRVp8xK3kFkP66APlg3JPDDPlFW1LRYtVkDd2pfwq
EgyGMoHKwTBaxwde3YSzNV0eoFfZ65kd559tJC8QwZ3AtTFP7TbSdDsjt3Uk
X7qn1WNd8UgF20E6vk5nVCehBYFlk7X+/XIIWzuMLcNbrkgpsW0oUIwnHQzJ
AO31/GRKruQaBIpTqwdmCuz0HUx8Inzm6zsJNYiDcV3P3TML7WqVTFI/Jk/P
u6wSBKTj/qqcveCj035ilnUxjFzZctYIrGx9v0W7L27/YIZtkldUyqOB5r55
rYQyZ0zuoX9idKBlH+1CzxnVB4n1TEf/z2KG2kqUX1cy5rSJADlNXx9bRyjI
pEAR+z7y4ZDP7jliSkdKp6luGqRGgMolMfsbGNqGI/T8AbbIwHNLbNZi/Hfy
SzVMkB0kdFbBLqt1C+1I4C6pgBcBemWIr32tqO4gsoWOdxWZchjJaJitQJxt
XXFvc6vLG/MjRiqUkVY60M/7rTyEpvxPKFcaRB39RFUQ2NpoD8HA5vGe1MOu
xvhz9j3eUnsO5TsMulF/aQ3/oO51KWszn8tz1zK7SU0b2SBt+dx2NuXIl5t3
mbjhG3Elibz092W3bLx8jcYhwQd24agd5j3afH2MSudZg4Wco2eoMpy/Fb4D
cAYM72Vx+aZ6JdeKY/RiCcLY5HqygSus2rvx25Ex0pN4Ydl9THq7vrIAwq8F
LrJV38Qd4wGWA8Z8SbjgtqqvQonlgclnSIwremEbYqT/q/fVG3i9QiZzzmxo
ARSjdA+1Co3d5zVLqjYeiCrK6Hr4jZlAl3HrZd87dhMOe8sSSnVexMC3sIyK
Q9rVeWKj6b11BaEHVZhkI/W/2ohHnOFy8mLtLGBaSRz085Sv2c/6vbGe0CQ+
+FVQoX5gIICER9j5tVwG/mer/pEq8SQvk64Wiu9ZtBRTwBZzEGD1mzywwDUH
IecXzZLfV3g9s6LXhQn9pnZDxG0nbBkNp9zpbKE1vGPXfOx3OXpNbLF7ZsH8
s2xuQR+n3SlHojTd/zZZ0aOaBP6KwUxrTwjousEt3o4OVKorogI5F+f7FoPc
+JUrW7EpCfXp0AoXO2LVSpkncpmJK37dKJzk6dymw+l2oy+CrgiGDsN+r37e
SGuuz7jcf/xgWmy55T+sXv9GWNsmCkmSx4fhSKYvpSxL4qNlxdYFQ1y9K9eA
EWgTBCskgbFdq/dNxsLWPyagQN/75TENi13W7lndMhLasnFDyVJwpUkFtbMs
ePFyWOtQWqcjNJPWWe7g2sFcpJ+Ecfpcav3ZYJxuYI2neuAhZ0+YtdRakN7l
+JXYcFAklRKHKCfGe9FrcK6w4k0+9T3wvk4m518nSF+ae41DTAcpQB6xYnN6
PJYClibVVSYGclQFCq5U4h0FOZAiQyJpZZrWzyhMjCRvvSoki27Q0uF2xMEd
2+P46Y+QIuRbaCwwAk1EdvvzhbX6CGi7hrJQ7TqWUJKfWnSilCpQSsglASnG
exrRfT/WBPVlBYUhUaKH0Ka+nMqrXC0/xkAhDAi5X9b1xX+qIGe1IkpgATdC
b2enOrnalYynDBqvf6jCnsXqr883YhJsR2pBn0csy9X/HQL48VoJHqr2yfzm
wDsNlcSWEbzUCZ+RPg08imbhdPPGuasCXJ8y78edu+eTX4xvh0kLo5KsDQ1t
mMRS+/TphEJ3jP7pCXFmehlwbEh34q2oAnRr54X8dt+ZWgbVg6zIem2+rBWv
Oixo9hZUHyD+mfpJW57pDcQhTiHPQINnFETQ03Kmtbl1g0x4AomF1iwxA2xr
Dl5T8uAAw/MGUtpJvk5LwDpEyC50Ap9HSLhai47D7er93vF7AtIuQlKcT4hN
gXv4jF8TJYHdqFKO8XU4kwbqIG5btYhWrOlVh3ua4TQbUuNETUO4WmhBncU7
j39pHRx3GzzgGDYvSu8ADtti9RO8StHY/kRwr5LwGpRDyno/+6ocOnnyPuy+
9ODL3hsl71uQeeecltDnVoN+v9bsPmPGc+GZ5iJYaSAng+GvQN9Ia/Ddy6dg
yIUTo5fY5DXH+kDRWnnLII1qPLU+aF1XPsIXuqilWCfCFod7yS778p0UACeU
FNDRijy71rJckaOGD55/yYMrfoNhR0fuGYy9tBrmFXf/1RIHV5yHX/6Y13mu
8Av2CSzVZ+LTWHtyUfhzcmtGze9SRCi3mpYqxuQO+F698JpbMT/y3wyPygTp
cQJCFDhddv8pBLP6+ol09cSntlXiGntYrtV5qlL1KgBcuVn1JFsfDRbnKAxp
2EMK4Rs6MSaYxDaUlhjIPX+Uhsz760MgfhxOhYwwek/nwILIXHoj/SbiQIal
DBNPWdFTcfPh+3LtmAEwtzGZl2KdElupMuKvwjYPSPgLlWRBP+B2+kdR6OO6
yP9tITj/Oqps4iyRdkiLDwlAROW6MWaDDZftaN/YKLjIWNV6awc1Al9CaBE2
eVljvWOuec64ramCdDIm1cTXSez9yVJuVLGzxYLgT+2WFdMsTDl4xJjM2XbE
0XxcpR4Z3ItC4vyHuuYcrVENzPv8u++wYiNyGQQPiT4RXIq6jM9DbBiPuDHh
N5CBz4jjWZ3+dZoFyo3k97Ada6DySW7J8ImFuFwmbk/yaI2E5Yh2iR8rAURJ
zmfWU/3OR25Mnvlyaf1alf7qoCw+kkCPr+1ArEGl/wt1E56JeeK1hlg+1C7O
/ORKuWxRHwvdtFekE32GmOIAAYBq2pvAwp7czNAdbRSJA0XoigB4ZiK71E31
niguexMR0XXKGOOJiQ7zzhJ2L06NIX3LkVPaK1tYHQNJ9btzK5BRClLHpuIl
D/en8/UJMH9KszibxaY3Rq+7MdiV5siCMQLcKlkafA8kzJ1aZmQXv1Cxrwjy
b92meSB40iQXL5yc9zIlFTxN2ohiHKLWOeKUaKbKqBNShUAFcGKysEFqR5mX
V58UbzXFcLGfVMG7u3JWylqYCuHjv97xG/D0RsWcj66OXwYmaPNIJAzh6ubI
cPnByaUWH5/F93QssDZyYXLLFPnWIWvPIAaeL7eeGgw+J5LlizrnCp/r8guT
y6PeRKD38JJmwqxUpa++LvfC3TPbai9hfOl1z1kxyERz7DqFp5DaqYzha5yZ
upG+PoeQcndJXPtLscBr0p1bknRqJHD8bQ3moozbjEZ3ReN8Vj8iuSv7x/Pi
u3d9jZxyW9LIjxA9qjsVMdDBn9avtCjnCon9V4pSYN28abQV05L3t9UMuCc+
2a9p13UQhJxgLJd9cSET7I/Mh9gwFM1nD6/KrpSAklsh/cBncmeaNryarzD5
Uvx42MUI2W4kyTAnC9E2aUK/2/nUvsrvoUI20hiXv6XXkMrbIHrWpF7tiRSE
fwfwhnbRCgMgDIJGJbcDmHgM8aMq9vWOjOCudkhUKizyBnurbPxD4XdQYOzt
DYa8o/jQq0Y+MSI8H62RmNwuDM8GP3MNlyxUVpbPiVfcbd2V1802a0b0+0pw
poNlB3znF/goaEkoObOV+xKFFRi4MYCh7S2TzP3t1pbeadMCktaW3kj5Bt3Y
hzOpd4kvAswIIEry3JQYLsWZkbhMk9fCFmH9CeTkuDo2B+4uvgIGoS0G7f/s
kfwmhHdci9Aua9EKtOAOqZZg/oa89aDhZoACeEBvvELezHplGrtGfLvON4h5
02i23f12VNfVJqZNikItZHskMqw5xrmVqJvFFEh3PoJD9rjLFL/H6ertz6nF
hFnpZs+Px4PjoWmwR9mrcA5wBWKHe9RYbna3tFvZANluEUtkDxJIj81N+jMl
stGR2a4COzfSBC3wH3Dw90EvSjcPmm7a0VRJBxj9CL9N6Pi7ZJg4dYQGvwnl
UQLiaWEb591TezubL8Qfr1/LY0Xbmr305L7XjPLD6kuvRpB9JKNJtdZwW6pM
Wpb6hFOfS9rXILW8n9oQrsjPcsVfALVwqHseusnNl5cat2lDXYO1EZ4We3GQ
gJ8OSaWdKz8Uq0uCh1tc5CROPSNo2VLAmucetDN9qQcPDOeFBeNmXCjY64mc
y60dNPFzjlztjGe7qydzpeeez03U/6OwaTEFb0nCjaxdFqj1hxv1eFFWl7Dw
bCQe0b1ZtOdF+box8BwJklkYei2pzFGxqV2d3st2MzxMQCBFWGIIDRnT0hEz
teIv2tw+ha4XzV9P4LEU5P9OaOMPLSOPySH2myNA3kHD2AOiwf815FdxPhtH
khRAK3xaDZ/21wBrkPG+eexWe8FQ4s1Dca/yhNOufVEHTKAd9GVimMxWbjTT
U0I1TTD8yVggH2wQbiUHflQfCcNC86h4z66ZIfyWVnfJj4XQcf7g5uOtOFGZ
j247RnRO0iGFEBalnSVn7giMrG7AkpdvemVSHVCSmq5svkQTgA1Y30PgJhQU
G2Sl348hs4pSjl8RZuMHpiIpjH1Ur3zcNwlzwzoRUKhQivMxoPByxcyyGVC4
IS09EY9O6/WrYBsdFa9QNJpZb7Q/QNiRCxKINcKWygLFBMI0nDlTeaSWTj6q
J7qIbbXy3DS97x3ZRgYtZUrMzSn1Ew+gzZa7N4IC40F0Rqy52xpNoO343D7g
V+SDJ9xsDWTuZz3eJDAnu5BmvhKeDeW0rdrCdhOm5I1ttK3HQxVVQwoHHguS
yH8YPC4gLijRD4P0Eh+WqAAFnJVdFFjXfeskzdWIfhzf3o3n/nYJWMIgelKX
GJBjSq0jR5kn6PIiJ8zXJw0iuPf/E975LakIpaR+857xVsCm3t/h9M483xJ4
/ZE4fnunQM1zqHqBG9yQ/8iP7LtUgQPhFmFX9KztOfOB8ETBjEuYj6BZ5ET8
VQAv3HKhiv9/SqVWhMYU1GtRE3NZ2vDHztm8nK3CD1ITepKEgwq9n1cjJ8yE
o957eFV+0TMZEazGDqS9KC+RDgyHi8vXbC2URlS3pp1v5GmOR7SR4aw7sTqZ
RDzRZ+9bsANJXnWOEnlhluWAReGi3BJKMW3L2mpxUModNKOzdbdedqfHE77y
ZQ2E8tZHEXDXoTirCvxnuHzWK+OcFr7ncP9rRIqxc6wMFbRZYa0qhPexHNy0
DKQsjFR+PMoGJ0FrXP66PrxJ2M8aQyiIMIgh1htVb57Er1EK+bduGlZxhrtp
BwM34FJJsB3WtJhoCjCqpH5McaRdR4UfIlgY3A7UDxqIIEQnofOx3prd6WNq
p+LC+x2Fz835+6XNI2FHW9B9mJf41Plc2SKYN53TBLO0wMV+/xuuSodL3zWS
FXJJPMDDTea+SEhYnUEGNsQU+jvz1GyGPHht+PgLBtPKk1kdf5tdcOGt6aLL
sqcN9UguCAEBOKoYWgfA90lVWlQoLr3f/Kvhwfz9iIhP44z6YthjDZEmayhf
ssQuNhO7mT/cUIGVH4uE2V60eil2B/bEyVsxmyGBN3E72ply6lPcEAeTb92p
uuEx5UF5AjAWzPBm1hRSPjgTDqurqdFYSRZ4mAt046+aJTRUvfbQ39WF1cCP
llsqSOk9tjfX0Vf254KPAF8EYptQ6ebRhchkDM/DqG3TtVsKQRiKKUw/CYd9
ssCe/ymtzWjbY+2bOArEismKpMCPhTg2/KdDApDyZAuLCHJMGF29GM/zrcr+
gZEpyI0sIaSaTEzGZ02xPZ5wT9wtF3+imx81qNa4abx2fwlBIkc2UOznnRNS
rTodItVB2TAt6KPrfCZSveV3lZa3n23rTBBre8JzTgrNsjlxIyhs63eVNIVo
Pun4p7vZ+KRRkKsOz8ULKge0CJ5vr23LUVVugZ1WKW+nvszr0NQyGi6Z8egz
6fbgTW7RKusAGi570r02qkmzaaGeFz02uuEd5OXvi0Fgdsvbu9+GSxWGl2f3
CrDJg50GTTAC51N7Q336qkplfubx+gEgQdvh0N/GjtJu2maKRBHAC8S5BMWz
f3Z5E1eG7uVUeBIacGEqDKU2IdbzwXGgezeAh2H34efD6wRWLT4L84+QkRtq
d3fqUFo+oDlpJGzJV5ACn85ew1qzMRlEe2nrN0Ou41S9WRVhL7duhWQXfO16
hSe465qMCuQ7Dkz223G8uAV7vOFhHeZ6TDIDEg/CSsagXiqTtTeiUKmyYWSB
1+6mYQ1DAhQWr6N+RlKlyzQkRiG9e2x/Q9oHip8S9udYXKIvHHShDEm32m5r
7qR6ABk51AsgEDVn95uy2vZJP1OM78/Cw13j0wGUvzRsR4I+ItpdkZ9z+6GS
Bn+S2kb4vW4Oh/F+9zme3X6FlVpReMg2jOpiecj17WtMMxQIMvVIx+309iLe
yb0EyEKH6t7jug+Oke5OiMuXNSLkzGFlC8pc6122H+/uua6fdMb9z84UDEcY
52bCqkjYnifLQdDmIl1o2DL47aJMR+5k/UrihkFZpdqB8eAvOubPZhJqHJi5
XySvmNcuC3HJCYK7T67Sdpe1UzQhiHjdplAsZHb8mNxGX7iWupFt7bPncCuD
YurWsTOP4kgQ9uNHIzL0pDQnCgZKcMBT6zv32zZFDISkuF37w0THLP5TECqD
QWJJma85NBdfnkVANEyeJ6cJzr60M1JmFcavjL2lR+v7raPjm4wu5Z9FGgJ+
a0Oxt7bzSv3tcqVHG6nK2H879Forj/Q28LLgyr3I4ryzQSkL5qQHKckxtiIc
afqNp8sW54AD7n+Ml6ZjNqzlchcuIEk60Vh0TPPvsa0FdB+QFnXhJB4lG6Nn
rcJDaw9AHnVF+d9F4i5N4TOG7EFJie4N4O8aJ4gaoWFu9tPuEQbOdUsxLbk+
LONR93HpkqlYp5AA8Mc2zkCGterQ6IntlP+GttlK6QOFrKRrCIPYU2rF9j0g
2Kx3SMApcDHUTwnGsMf0Pr/w36ghUHwKRUoE5/R0d+/t71JcI/zOnUzfWStz
FCHxr0sybxd7J8W5sE6leH7I2Ro+azZyhzj0tCpW44fulwROXpdwIokFqg/A
ICAp1ciXKSDN1nVYeSMysU04QGeCTY/3vZ8nLkkk/yDdQr7p0V2/zFlINbiU
Dw47FFzxAfz5erbT1cjvrVYc+rKPEvm8Jl6iN6GuIVBy0IXEJvIZoZlFEoqh
ZIbHb420p5uBiGIW4DpU885U3mNBfzs8rycA/6V1SchajxrTD+CsQzCsCWii
PGC36qZy2Tuf9Jejeg6aMNsgFHzJ17ZrKJX7IQEXHM1ESrrmRQ9iZKb4vSGQ
DrWiOvKArQ0ITGD4jMJ6ZaHnlLIv3gCEOyW+JWihSwuHAVLnyik9q11p5wLr
YI+9meVazq3rqwi0X/EqZ4aBjvC1bIs3qdjo7Xpf0Fj+ZXNadUphhAcxHUyY
crGLmHsDmpw9HBgUUIlXcauWi2G8FEuDykX0iMyURQFUWONhs/vn5gwYxIoQ
jB8YKcDjnhXT2LTG5wDLBYw8ItJdKilwg8VKM/ad/IO0t3ZFaep3IfbwBJAY
c9lsuGqITx1NuQ9rg8Dpw2URJRecWbI9smpilBS9xyA9jqStF49U34RgWtuy
hoMtZfoMwRfSmG+xRz5UCXRK9ZzqZeEGC/kTQ+HcQco7Kbv1DM95iNJr5pyo
nlcVL6cxxakRx9NyxIwszNL3nwmNMcMChzcPMvMSOrEWCGPh8/OUIsXRhrhS
zD5v5QLtqnB306nJnut6QZL3iTEaL9wBNCt2netSV9fPbzWWx36kpRDB+wxB
MvT0aJGDm1deROoqMurw7ushkYPC7zQrEbFFOaVbYq1uzn+YGYcPTnvdP5UY
GxR338JInmwlb3cIFCUfMAVi2Eu/k4Mo29X87bsFgxqTdVcbx7C6d5i8A+1l
/asr4dGDqd3eXTjs9NrIbbI2wzvg3R+/Bnyd0lMWsskX+aVjHU/nF/3vlJ2X
sKrkhBgLhkbbhrlmU6XhqcrjUEdsdD4fGAfjxMcJbML6juNLao4Z9bTy56qT
JAx7fcpHCDJEvSKGcD2JeU+Fyq1XFuQxbwjLe6XgAv9mpVCOzxCtUnbS/aGN
kpNmGdX4ZwUBmaKk+SPHrPsiEZ50haGTv1JDj1Xi6wnruC688zsF1qStkLQ1
mMN0f2Q/qFdHvlF7L5ie8/lnPdPrEbQzmS2QKNR9GAwon5knoAlEjeeosKJ+
96Rs546EcgYRR6j+3/wM+staxI9qXneI4ZQqlQ2Kno9wpXUdoMbK/jjzLbdn
njb6r5P8NeGZuu1yVIZmW6XEhYrqg29J1a6flpZVsQ888R4wFb+RPz6V9C6d
uQcEtzjUxGIv5MZFWcrdupEjT+ZlfTGlW/XOAsuH0j72UidtJZsH83NXtoL9
x/cQbcv+5/u3i+T1Evk6w6LYNWobAM30M7GB0IzmNV7q2baZiDkQcLsCba/Q
GsfF8BogdIwd2uIb3lKYUSROvTMyeJZ5MrYBGDKpsmLrOK8WYfaqrgMb63La
8QnxLnvMoNycdXcmHDuGj1JxdavrfwomaYWrsvunXcjATYKlSgJbJPCWS9hg
fJuiJCoYZrg5OVAqvsN8RpQriGQa7hQbHXBAaKVN2UoNoZDuyRp76PJrFRSA
07BwV41Ss4Q6wl77fuHjHQrO3gRV9Jiy14HBvTpo/6CA6T9MNssdUYmYg5yi
vkTtLEJw3eRdLDtVRdZ34SDEEFWKYiXLp2q/GYtQZ+OT9t+f6rLRY4sLTlNy
v9fCyYXUGXbWBiXYZeDCdjQxXQ4k3nWxcZVeraZ17jKKpY1SAXUINjr+voNk
RoANCHiyFCUZZnmrABkr92uTjBRsjBqNElcHgzheNDSJM4t3OrJs8csFgGeN
vr1Rjf58wq6/DjLvFU5vRUaeF0u4dsK3l3kLw4kbArQIsKJ9cSJlGSTmIwIk
fJOhb5h7qh+ixPKuIyBaayP5X6kEGWLTz5sfXtOjHYDzujFbjcr1OhBKPrvk
kfA6xTpQvF3teX52pX4BVm9vP54IFPe6XySkfqYLPKAKXWtQfcyDSaW+k1NK
ccfKgizSnjSqQ1bVhPSE9WbbuCz3Fmb8+GH+4oViGfx2VN4KRBaOlnzsbXQ1
5GwSbVjCq9F37dYdIclkIYvEgxKrLsWt+08nECM7rHKrxyq99+TDKfe2JIDU
PxMV2dOuKiDU6NGKMp0uu9N7DvCCPRW9y2uN41q+BtLkWNY3SEkLjBrSkNpI
fM+umNZE7HdNA7gmbrOkPbmFe32PlG6EQ3FxUERvwQrxPYNPP1w3uRcSHkDI
ZWOmYPbePFIBj8UN5cZi1FvEBRlD8f7I0tvHNMuK67ycy2XCMEZwefdeTCKs
4/sEfaOBz0hHB0IFiCagoGjvO32y1zNon/pcJJNKWlAgzQ7hqzkLH4LAKnU8
4nnU1OrmrwccnuzlYOvF57RhcYDmjBUds25qA2DYDbMy+FfdMYH/KVKbzG+1
m17MHQ4pMRKBIz5YNPyRE4OUA1XqktkhanZ5M3Ii5uvdu6fCWnVtdXyyn7nH
5QbsGB4nBhksiKDtJHlnw9IVM/l4UwA8pIkVZuq7KnPsS2d1+AGGYLPGKLLZ
Tq55O7lVG79vEbPVR31DpFRz/ykiOPFqJS1SH7Wcqwg+rqVtXbnPaQppJeCI
zyQVXX+vZNmcCqR7ysSX4VwkFGc/4/z2Q1if3lU5SHkWqsJfibxFF29fgz60
DuPKVkev9BVgXKzzdvDJiP63dk3UT5QV9nQ/xLNz0K8swbjOMp9OXHO7Fk2g
Dkt/hJNu4FfCjWO4XO8EnJ2PrsE93SstieUk5Rs1+WN/8/0nX0LfZIU/jPOu
/KYiM4O3B3Atn8k2wzaSVL9umXD3IwPPAraLinYf9GsYePPo8JZDuy1gsbbE
iTd3HnPJM5jVYrrlQkzdPfkWFVC1z3cBirve44odT8AZI/cV3GIIu5KwNt58
PRrvWW2biH5+brtRZyAgvDTG2Auf8Iz5gWBp1JX73NhS2zcls3wGyLz9AXJY
S91YQS85GDWh52WwdRREN/6Gs8YjHoawDjluAKwB4ZQ/QQAo/YZ3cqhpmnYQ
bFRoV41g8sTUl2XSZLxUO/EHyEJsKAfmo8nVD+HQ8DjS1++WKDf33KgkHg+W
QZnx9pSM5rf6jS2dQCJU0VB1ZRNeI25qr7l2fk0XbKbzLBIIvDHG+8TBE+CY
aIdoX9n0jjctLvNLGXZg/L4dnlrya44vITLZqt6owRnaOC8W7I1IJJNnvbxn
3Yy3Z8vod8DSam3xIxpX1aJhRzSmQLIWo/2JdRRfZck1xo1oH1VJ7SLJc1Bc
X47LS9bmxxlv6O85gStMrZMJwjDSt2P/JZ+qh+DJB2uRCN9GbRq+Y79G48Kj
C1f7PpPp/0oSjPwiVg+HGSAUCr1JcGC5Jx8pa5Abb3Wpjd09SH62MCh5q4Tc
Z5AZTue+/2sSJ+n0KzsqIlYJvsaJCJ0hJ8AwDj8ZGZjg8+xeptK8n93qfzVe
w2B7e/ua7aoy6YGNAtQcS46oXpIN3wdIVUbEmkVP4oIb6mpKEU1c7dC9dxPw
wKUDUQtBkU2uwODdfZpNOH0in9LUXyZr9UbH7lRQFYydOv1nILc+ktxYBpJ6
eblYr3qcLBlE/U+9fsFfz+4UUrOFtKGBIqcvWj2fF/qm5noqYfF9JGlApEan
S+XuDDTnCHAbvSV0aXt6bE84T0moBzIR9GtRCMwdMhYgEg8ziR+eqmxIsAWv
1nWix8eGMdh+8R9IQCC24kV4TxR0JeKrOT/nhrdGr7EaY0TknmwUi8AdMTzC
xrvL4CafnZtD69Zb/2g0TvxSuV2YQzMQpMwlPfqogKpDmOA1WoEZayUwvR9T
fqmt978BJ8dTABfE52sOox40UOEGjaAng5duouoDEcQy5aV7/OyfjzNH8za7
xK3lTTgXOj6M42z+wOxk5Msle9iYF8bdX11fKdhqiyWf9GAsp5UmGi47uo79
7o6UxThcI5JCI6xMf1aQVGZd+l332ltNJ08XiOVwwKzgcTpclaRA6p0euAXD
tHU5T9Y2BPPwcTbRsKwuGROqYGUkIGeXf3n1Sm0V4XEKKyaMhZI53iPk3xDa
SjXA2tfdIFYNrVYbZR/eMOAn2ijI4jsg1N4/wLmAnUZymhcwOCjWVmpWyjqG
t93zMQT9UrPRyq0SLXyT3HU4+9LoaQGO4JZiR0Cpxj/U56P75udJNu2tl4QU
EhS1LqLpPJ4PiNCd6SAoM2zdSGNug24zZM5fneJ3MbTEnhQcT0Z9fADDC8SD
guohQ8cabwmkz1jkm4IYCbq/aOgAm3Xb4DhljCLOcln39/xkT/dVLKuMrFFn
145hEXdtk507hLxmZVhyOL3pvjB6wy+hHr2aIXicdk6T25yK6bLNybmsu6pn
OoR74jk4ZhqlLRVIdM2muMdZLPnkyT2l0AhNv4CMJYHkNN5MxgDwd4NWcJi8
F4NwM8diryDQMGb7D01LjrT0J0DZPRVJbHrbWmh2TjfCgdkd7RNVdXwGTFp4
FyjfnjMkA2tlmeJJgLuAnYRvUfVYcDlq80vSgfl3nZDTXxjWC1T3xb7pe4Q+
AOHM1DuqWYTmNzDPLR6JdmW3Ya5ql04XvPQp8hJMVyC/zEZUXArlNdG+MwZF
kItxQdzCZo6r2EEVI+3FVAZEAWR/P/HWR2MQqi6jMIH/thwuFLPF1skfftuC
D1dNB+7c4GoIBastK/8YxMId8VNMPyniMKnOjCCvRpW7ptlGKHdfuyaJ61Z+
rxJUtI3K6JoNkUcb1vRLH8DXBXhIf/bJTZjkDIcMegl7DXWW6bQpgA8O4qva
WXrwnuW5XGVZlmYjegBKhV6IYtpwuHWA0C6j4X45UlXbjUFSdseuuQWSoX4M
eKU46/O4nj4paR+bahWdtbJRwbPTWlQYdds0Xz/xxkp+i2orQOINDDWe1eEs
MqmzqDKWC+sisdet7KtfKsruziUKrGFEOSUSELM5wSMCxMoy/elWeyRzXsAA
7T4QIDVrri6W0hKtuius1BW601UdYvUUIBcZKptiSZMlLV5AcLs1XKkVCe6j
XUEtoT2VJ6+gcmTmIYfnMVFOYO5g2LUHAlPqyF/7mxLQW5b9fmenMAJCYikU
NbfFm3GcqBYOoX4oau88ED+YgRDNq3O0tFEqgfLU3YpeQpepMjil0om1xgZg
CemrjW+tEK6drqS526Ga12qVI3wa7hCAmQFV48QbTNHLCu4/cNEz74ZYk+xu
gxRuE8Lm4mAW9xNdyCNrtq8nDgQoRDhmxQmvtxFyRpp+TgDzuJr54C/5FRpM
LFP2hwtgfDOvGAK1cq1oah/9gDEqT0mfFvw6J3ZKXXtsXMDg7UuHsk+ox/if
CVczX/yMcTURa+bE6cnzA/v3AKTE8McdleTWYOEVioTEN+vzjTRkpgi5MS7i
sBvE5+H4dRwSjqCkD58ARQ7ImYSiU/pJAocvQnw2mwg1LC4Ejvp094myylmV
94n3+uVNFUZ/FKZ7G1cTcE7xPuE6QzJ8iccIGMKWw68YxQeBfj0JzWmBoLvL
EpQ/lNAhMs5W8r5TVuWYYsK0M0teiIMMoPzGiLhxVlUXXn9OjdiXk5tt4dro
21ZY75cyN0nTI5/7RhZlVzuERaAo6a83vfBQ0x894usequ4qzOT/rJHZSOIW
OGv2n3GN1yvL6w1RRLzSyr8dwJwsdNw1O2+/uqwye9wGR4QNCmtakTCWtOnA
JCABizF3WNwzthfPkqZjdS3Ra2xMTuCYHJHu2XkD9+90pauOoLPDGeLCM/bQ
Cv5jGXXP/UYeVlZMh6JaTMYU+9O3fBikL9hzYWsCFIMwM66DKBGmPe/SUrDO
1i1YcdCku8uvWfS2TdTvyVULKqbdqWGnz6105rkUEYItc5fKqWPNr3NEy2D+
+ySFHXgzJ0Bn59GQHGZO7iz8+SJ9lVWn4Cb0LTQZw9dKpQXtlqSUtZPbUxvJ
I49En8zHWAoA5wi5Q+F49gjsEmbiP4XwLhHEIP307IAk0PE53bd3DpDtnXQ3
sGXSAt831CUksGjGGPWQWEIUFrkEaAZL3gh51edvo6sJlGzxeAijp3NZJEsm
QFUd9/p9cGCLXhboo+xmtFCF4Yl/gjl0+YtmjPimkckWhVxEtL/yHKxaK3Sf
ru31l3TXaCr3EJtNVxCHPtjtdh0CrELG+scVJcWtAHmzCFEpjnyBY3VgscEZ
0i7Ag5q9/XqK4bg+M3/gzZfXZ547fZRIKFSnvZorKtdqwhxv8l0TUKCYZ2e/
VXWaOsGpVDAVOG0MRwA7m6eegGSkURVs4WmCiHGU4a1WLPwCN6Pi1O/xD3J0
/HRqH8GyorlOS9/TG78IHiU/X2xJ1z7ME4B13Ju/MVHFKI/7jiKwwlyZXXyP
6W+kXaM3EsD+Fm8vPLj3NAfY6GXUqqcb4JNuEA8DbM9A76aMFMLQnGmB8vP8
anlMT1xjTg+VYz+xy2xLyFPGh34lB/Tl/zGiQe6K+e15afupW10DXfo1uJNO
phWt6pLJSDCVsw3YSbPnT5no5kvczoth08EVC1KxHPfMuEN/uFe2EersJ+c3
CuGJsKOHs6goFQ7cQpnIK8IfP1PyaoVgpQygbfqaeZi5gkrrOCmu/Rsc0QtM
sEWtOyDszu369Mb2d+bwV5fX0qgbVOOVw6/CNrcM0+7WSEmoRoRaG9UJatt9
ZPvhK0DQm8rVvT1qr/4SF9evcAtr02Euvh9EXtP5BFvrBj6/5/g+ZS16B2e4
uWh0sqZD7jiXuo5luHOgyowvlCcvMNmei2DaUW2tuKSKc0S5EZTAv4n4GlVr
DPazrcYTIUXWUQ13/rwn4G+vWFuK34jK04tP9nKfprTKTVpSFoUfKU44BZ48
7257I5sOV6p8PIWxT4X7io1NgAKJmyhRc5v61/KR8LGB/WPEJ819KnjPAsnD
6zLmXmCsKBuGG4t+i3GE7GemY2qdwiXsmXBsc2A0jP+2bqcpCID8dis/q286
8klbZjoWMh1wb07+UVhIqqPx2ObbWhGjVzhZ5FiDnb0JX2JNEowMz5Y69iau
vYsfDenAAxc9AelaxQp/pl+YpjSMCMN7R4Jj3YPOP7Tot5baoMaBG8oFt8rg
2RHRXdZB5lL7il4b1gX3A0eFIbTW8AEcjLww/hODcH9gGHioz9dFv8QBtpZV
LVV+e3G0uDCq3A22V0+BawzTSzwm+Itu5PJVR8d95VWD0YcbddOlNaglQUSe
6LVr2rTRy0tPsGGA9bBWNdFqQ2zIsjeLoEwPHuES20NgMvt51v+FBc17+gVx
Vug59E7yjXmGizYsaAlkDWy4KBRhHUCCLUm8HTOweDUIjbOea0DROB3eEzYN
FWq+5KP/sZvezSk8lh4nQehB38CegEX8aQFlwi6WRvDKxQAxMGly7Aif4q/k
bGqr01T45P4vh7mLNI7l2Kza+NUJw0M/w1eYts51lGyu9TQG8QlGbkILp5YM
O++j7LuaENXIyB0alrQ70808Ohrdbbz8Y6ourndL90F0s8YXcxi1O6e7nnKk
d2jtSWfdHvgtWI1ApvCMo9dbcid3ElXiyd3Qj2nnjdO2561wYNmP0RwIhmPH
ickNVJWvxy7deka26dxF+eTccT8duSPMO6sogvm2BSlGceoWQI4f/9UWMl1j
yUZXnObG975Z7dQd7v3kDvO53MHsuFDuicLhCzI8Gb6Ro41Ypf3nXHqamq+D
r8the36Y7z2YgM904j9NqKBQnuzhwP7MiZZHcT4KGeQu9smJ7cGwOpXausv4
kuidZyxntD7m/jLfGO0LwEl7b2SE4goe8tR9iHV2XWl9x21kFWNJn1Vgjpdu
Mq7LSDvEqOTJbRMBIyOr2fNQLL8hJoG+mOdUuF/afyveMKQFk4/hDYq0OfjQ
0PD2uP+ctRzaUfCnZIdhmXSHhTM3OPltkQHA1Enc2hVpnWHgRuTTKouhxSG5
Av5eGWvw57NbQ7xtWLA2vevRIRpu59p1F5E7SnTMO31NJjMiPv1USDTUTgLy
2h+9x3+AY8P7n+M/6aR5SL059tPxaHf+LvG5U1WTpkmwAWNrRTgoGuJJjOvR
HTCYfqbaw5Qv9nf/wFt+WkIzoZziESqYd493GBPbX+inP3RvOCCrOJX7ZDw2
uEta2fBnzn/vBnMjsHqh/ykgoaPq30qHH0u7kaXX71DCdEd1nDOB2opvpVRP
Si75YZ/3L8hXoJ46PE3YTNL0QXO8FM9+uLX4xwOMhzMw8667KqehifG8e2Wp
E8ypxS+J4T56qPvLGvPBc9rQhohs6p24FWthuCYfrKVK38p6VqVCIgxASIHr
nreDPft56WS88XrTj3qqCiebSvrFvlh0659yzUpcwDXGTKHcNEMHIj3pLakQ
dIP678g4Tp+X6iha1y9M2cC1Su3evMd9RQjeHpQm92aeQvmt9gL0Bd68CHQN
asIAwXy00y81V1EoDeT4wkltlwpNulYG2Psr7764SnNt6JZBFjnl5hnG/r1w
5s/0DoSbdJDepuIMcdSvhqU3Xynazuqn2x12nJeaSaSKjgPtvansW0hSImDj
RXrMgsAFYgXRKSMtHlbZoAFDupegEEdfw8BRl6qL3efyk+wJNgjTkgkDJXwD
kBebtRXlNFaacn+7vwoakwlC63lEkFyFZ3EAgXjTSX+jS2OMTx27wqY1yLEC
PXbbrd4M/gDeFNSYvmm/bl0grbAT1HL9wEmCtEdugJ48RzY0Byld0/90dVQb
LlajaTPIuwKJEaF8hRbHNrCnM6OKwZcnFRYi/uzXSF7IE+1qTfjS+jNUQLS8
6jbeoO2GIPE78HT7T0ICeMwA556uBSN+F4Kdfs1lCeYt5TTfzepTTPVnyJVn
0RuHJdL2KNH5z/mk0rr+SmbaiNoyqHU6a8YvBasb5D+KRM/vrR5/t1GGvCcT
504GwgJm0sVXUGYJnvXskOz9nKWmXlyqREZlee+iFjB4UT6mniDSyXsvqBMZ
9PQpESljlA9WFytuHgftHrGua0izGZTNDV+x7xyRklYJufR6AHHQSTeg9m3X
igc2bTmpdfDuBNY/bNBI1i8cOxImNC+GdILqICsTYz/pdA6TZOZ8FA0Z36Wx
el5BUbWhCMsepXzqQ1fT6S20aaQLf+1seiC7uiCZXEv7yvGOwI0sjvp+dC9w
C+Dat2D/BymaE2FyAH/YPCANcDQ1hxGDCCbob7WISGXoBtCoc/RQwljVGptp
k/BUjGhIiADijtDoynjst4U5vP5so/qnir4Q9Z3QKAd31JLmn/LX3mOOCKIA
UwMOWi46CAuWBGAM6jbE2ZXwJnhiEDGTEoI7xGqI7iq/cBw5fciSiqmJN1Qs
349o5yq2OWoEEOfreVXXib/dQEP1/ekQNKJKGKsCCIxmlIMVJUSQNyczG/ND
gdknezpjag5VVyMQ+nv9Q1KVNhShnY5xYE6wlkfgp1i+EoUS6RiruaOiQIr7
3bNFKE9WNaOKQi9Ljfsp1jbf1l51esXz4DKxjQIWOilF8sZ8hmbCJWp/gdH/
3hTeSKAEV9K+I4qQ3TOUI2gZM+j3G+KRcetIZVZvrl3CUGFSx+pt6AlBGenW
1bW1D1YG4IVCZs5ZSg7RryfZbxJL6G/aFW+nnE9uszyoHh8YgRIM3VR8qwg5
IgpPxFLeyiHWJj4NN5RkOqQn9uli5KF/Eu3/iBNngGytB1EfzLdGH6cExS1J
X6CoOLS2Vdp6lDf/01nyckZAXIMRMfmjKYC43UaYM8UDIyk95nPt2hct4LUU
YmdbJjhYytksi46r/xFbRFBWI8OLflEJFFh3kQA2U8rsKxvAhL4etbYPU6eB
UEq5NhvCT2cVY14Uog12EumuaaMUU58YTmNGeQvksRWgBQTTBgVZIUG0WtIl
sXiXIHrCPd2+1IKBTVWwJ2006T5aQ5d2ZQXFVSiz+LsDYcLiQwUVqU584Bbn
KzA9Q3huAw11YgWBMCWRv0zRzbKBDF0nDF5JDX0OttzdpHVd56SmzKtsj+Bs
uBnO3fHUmAW7ZhQV8a+2HYsn0g5sRZlqz9SsKEgpPWBxdyka0QB7IyIfahMy
z8YQEj5QDOad8c6CtB5fJ++Heu4u2FM/MGRuwHzIeC1sTDJDtrQ/9XKgA9IV
Rbsdmm3A5sJSckcQLFJlr5UrcrAZ/BB0L+ymChTcNdAiR6xwDZkEt5tQVuQr
OiKRowbO9Cb/BoRSd23MePu9f+TZZAkmpHQpIdYt9lcs+/3KsVGzDQj1BSIU
6X0bWL4bF6/kjvN5I39EjccOsubmqw2igPjjcuDjeMWnvUWJcKngOpaxJM4f
6qJZxmGVIii393muHk7lgXK6zbqpDsLiV/zVlEH7VV8uPaai6ZcZE5UpCdqb
ZA0gX0aXmqEcOMgUKh0xd+olfNZRmfunXeFAuyuuryVjslhvqsNMODhzmVuR
BRzywmuM99ldtWZPZJj7dNP64SKSeDkSeja2erp+HvT1EdWUMT+xmaQjcjlC
7EhUczBaLagrQkhPJ0DhD1MvhE8hgQQQ6cf14CEl96r/bu1syLYQch4cgGE5
LQMqi34KhgHzUAh3VE51UU49RvVARtmM3qIr10eeKN+j19EoD9XBeUBaRCWc
1rcXh4wYgTMZ7tA+zgzHYuOXYTQghzVXMybQK3TuG326h3Sa1TmhRDYFv9kH
AGJ19njdkRTKPc2u5UP6g+XJrd8uQ0/bcthevZCFQxzUdmWRMKtWeMs49IEA
XWCA4ONTpQaQ0VKV6mSaopxRBdvbTA1TcS8iPzRsGBzWEHA1aKyEPV5G9UsL
fzD/zvYoFAbonza1xWyGlpzsubFFUS3h9GGFk1gWxXju2xl8NYaaVOZwg3cX
S2T+W7qFBpkDJ0BjsgKaakOgxTvrutjl02x7KSWCbxRNYwCmjzgHmhDehzHV
bO6MaXuT/vZBalzHBwyjpt/YBg/Rnfrbzic60zlpe6ZCbpac+AOx+4VCjfg+
uTrIwvGMV9fsvvsR3mIR0bUW/P8i2w8zwbw9nm4FCoRTxdY+zexS0p5pnR7/
Zpqo3CLqG7TAw0gCLoi/R/mVgV+2Gf1yzHirqyZcRS6BYq1hdldAT9HImzuJ
Lplp+N/GmpVCEDQ2hHAyCFiSDXJj0BKZD80oHmG67Ai7Pa6SkdkNVsAqN3z2
Rcy5RgP6noiZMmdTeMTHrfTz06nooAx3MxQ8voOwD0zB0QiMdMhgY7tCXPwy
klxTyfxt8P/aSjbBNDxjBpJXNyBKq26wsg/5k2vSMeqInGjSj4erZ23NZ+a5
b292qC8eyariOndIpp2jOrl6VgxCQXxgzf/knVAjYO9eWAUm3QOV9sLttcA+
skBIvI+J3wrVw+FFky6Oh32cR0ZveJ000eKBGBrbLM1P6q3mMoI87YbNHumF
6+ImSQnND1WSCshbvF9wAV93/UsPNS98KkLHpJ0xOuJZefHhfOOuniMfc63v
b/Z4i7GxR4VleeOaS+916AGJEIY9zRSXyqnM5+ea+vKTPzA7qC+/gs7ESwrd
5Fekpv+RHyq9OkCm5wyZeJm5ONbRNWdFkZg0d6Z4UoKcJ21WLKYUD+ASbgjN
qCHqjrc8/PsFaRlBuoWamZtfXEx9hChXV/+gPkcHptqcDiKEUNKuWdu2qYsf
AXMyUfcGg0KzleYFypGUpdesK2s7arh64kkuzx9ZWmY/RttThsFehDXdeG2a
oxkLrvCGHWPunf+09eq9sQrtWpUZKEypXMq8E1SyhMB3OdLsAhO5lHLR3QH8
wBAl/Va7rw1MF+OmQB0Bo2pd1hqsCplt9iZmytXDlzCqjgKqRi+gTMiskC+A
Ld2W+BWI1xO7Tlf4X4RSFmLmz/zHqyjtRK5fjFgG4VlwUmfUgjVz8V0FCOsG
lmqJHctEG8FBrsM/OqguhzEOSWKB2L5Q5v3n4Jk5RH9K7midRn+ZL/v2rHCL
Qs4tjBrdY1o8ckTSlRUk5CGsveGfENaFxcFcoIY3tmwdV9rE4C/I291nFb2e
9UwskdVttPS/wIEnBC733DzJjpg6sOW8Adh4GHIpfjcQqNLSjn53bP/IzE7Y
CMbCVLK1GNbz12uWALfaC2VGX1wxh8xD0hc7TTHa61wq5bWrSViu0L8+QQ/k
ICD2em3Z/XF8RvMCRHl4IHyhK3DatJarjePO93Q8WjbcJM/3HrPm2YBCEZU8
kPzhSLF8pcsd9C2/je8L8Ol30qYB1zk9d7nU9JzclZiqYuiFG9NxyEGW3dwS
bq7BeiAt3Vahl9YUjpzN9jD4gpyQ/fAkYBcYHr1++hlqld5xmkz39tnNv802
eJ6vrB+q6jscbeDsLYu7sO2R1ovIo4lUMr5HE3Zv+IddWeifiIgbntxtMvKC
d/uq9o8yNsY7eLI7/wqyqbup0F4FH5IPa7VgPIDRCfxmfdYH4jdnskt7lcBK
fxmGLNz8ycbHxXehhUsogv/GELT2fJykTV5EoFO1VJo7SQra2ZzMdKrmyt32
Xo3x5cmGzrgDE0U6a0OFbZJ20qiH8DSNvf3hmQGh4WBGSZ06DR+pvwsTWxSZ
6l9OW6juAlmCmBm7dAOxmUJBhQSE3tfjtEWzG9x7fTq9NDDXQJBhmzAfw/U4
EH9uIJeN2nQlOw90xzqDh3CIJKnXucER97QMi6oXBO6uAfQUHPrhsOGTacTH
QxYM658ycbMiuVoihbRCjJKBYboTIhAvdBCSSFoIiRQ47mEFdAFDBEAqQ8+w
yBHIVRnGokaKq6FQvGReSS17J8ObplYuOVzXhNNEO2UJY1xjNfP77kgQk+ut
qCVi0O/eTHrTABzPs/ebZHDFZs303AZJwbkfnEKmj22vU7CTySZBTJr3+4Wy
oLUd69pygZJgQZ2kuGH9Plgjs049QruPR54tqnZA3yuyYKZjh7zWSqaaenyz
x+4RRAy4+L4r/Uc+A/oPUzBPh5884DR0lBbrgXBRWh/BILwzOKXxgEueT4Oe
QxOhI8Sy9cgxVSuLFmMunvOmKMwAxRmiJwUDN1+1YBU/Va6M+tH4z3ukcWD+
7aBJMe97+xUAPTKJfZSokxJXn3YFGEaeu8BLSabn78L3bV9I4SxBUUaUYTSx
hZxD4bQp9l1I8FbDzZzakeubkhpQbTEbrveyny5YFkmjh4iiWK7A7DqiyrMR
1j9+m8/zWMOs1lHhAd3lnHT83TSnEN4+Kus/Tmv1w69JcNCe/dn6OZFZj0bO
00waHss7IUJc5ltmnYy3XzWxudu02Yk/Vsgji/qjltdFHQwhWOhWiQPSMsgR
v7RTqE96pMpANqxiaF9/2uKhC1iUjj2dI68sOaPc4m0Kf+83g4206iqPZneQ
juF+bdRTFt3v4EZVOjX0TVgFIQz3cEQ1jTnZDYXdIJ3RhQKuFTiFEY7ckynq
E4wPuvsYAPAMGc4bT+hzGq/8YMz9xQwM3mfn+0woK616rnyHgP7ZAI9KZAbD
BIq5aWLAko7tmN6JuXKQZybGOoxGwHUBaoVDNE8tqcEBpeJQFFsvFsVuos3a
uO7eFnam8oK7PLfJmncjdw7CnkifH8fLC9KUJVlXO4iMnCgYbF0AYHriNDK3
bsypGXP0MJoD1dUBzQTJvWKONQDH/MLT8Tnc49yEEOlfIMONqPUnHyFNUdqp
UV+BtcV+y5dMsCnsN4UDvCNXYXI5vSeE7iu8cPa/3YuosQEmf520B4rrEsJ9
kmswwXMPJxCsa3qKiRGCaNKE1y2ZTB757o6355ZjK1Gi2eNo5aBU2HC3q5OH
oCoYChsbGqgYkNShY2zyDkv6wH0hwcIhbRHC6Qas8KNSivqhQmO0eH+VIDMb
YILzvz3jAuNzM7hZYweDqHg0/8pSeAO7rNnk8ArQfXxhyUFNFP9xrtAiBY/s
z8KFnkb5gKHHipBz4EQtACNI9hktyLWt2w9Ft7azIpOYN6cDtXZYjNCFuSoU
yjyBmD7PrmeWX4UypIHpii2h1fVyV5dpBi0row/MpIh4FrCJf/gCWn41f5Ss
LIas11u3WD48fkm9jkn4zkvhXFtoc2Yt0Hxph2NCY1t06QiBEZBlvlyg06Wl
EMJUdrmnEmsNd9DnOrpakSdRgSOLrlBZPyvm1iWvu1ENLTMK+jPGNwxJV40R
o5tmQNGF+JwGX1q4XjIT7ZljTqssexb0eh+zt81CudawcYnRodf9CdbnImlu
AZRLLRNFM2Bh6F6DsH97uad77nX98L83gPY7ssNdNfvGq/xtPRRVK8QWiXw5
WQe5i1QlTzLXTDXcA+qT7J+po0zzinad+rehCv+HwFsGfpMF7n/IZjoJ0+rJ
/L6h4SKhoQPu92okvwWq7MhpsRz6as1vsFFS2V8AnszIODNg+3JfeRvC60//
tXN6ZONVtdYbp8xWPJEWxzX+DovAon0shmvUOmnMcohAt150EP7Bnow8nIRl
AxaUHECf7+obNXV4Tacp5LIwUSUvNwl0YPV7QNFRf4olqMTT/K4N9w4V7Ebc
O+CG9KaVyWRdL5BD+khvOjXv5zNsJPRh2t8H8ewYMLkSpSJs3w3t8YqgGHDz
hLGZh6SnzxqT0Vg9Q4ZnI8n9WpOxa1mqF0Wa/3520UBK51AbqRfl28btZk9k
8dxsnVV76sUU6H5VF8TO3BT4Z5NG4jBvSYonXaeAo7abPOXsmJZTKoxMREMg
H/DeJ1b/0fXPzScPN6jPGruSOs4KY6rNH6NE5j4rr54AJ8vJqiJNbp5z0ELa
e11ZRvjp2Q3tEi2Z0pqsSNpRuNwoB9Na8ncFzZV88CCIR8q5JvKh2KEcgyVV
Im+O4YEV1o9A6R6jc0zhbY0QJvgW+QUTsT6zn9EsZE8PcSePloKVLkfHugxY
Rxr3ngAGNVvHsvW7FBBerfXqrrBPGHJyGgYlv+s99DuWG4fp2/T+eFcULDAl
rslH3gtJK8igSvudm/XBO9mNlocUnlmdAWAgUru5rRpmKUbidro2f1He6/0a
eLzzhok/zKAnYewJgYlDmFOKICRFcsCcoBIi/sYqqClw+GSIpbDtdHSwSVcr
vcYlRxtKlNV0i8lvJ7Hs3Xz/RBr+b/tkcFmFA/wuNqJ6SqA90vCfPBvIOHq7
RvdfJOifhQ69E1ISONzk94u84dUpKfJemjowRzn2ILdP+XVLjHNQgbig7ffR
y26QanCCqttj3HdbhT53QiTHyIxXbjH49IBB7cWd7rQkRNlT+5kl449YHi6L
KAJGMjHeOG20mbCrrDTf4p5J4tyKaNg4/ZnugCNXXg10uv6BHeb1I+5MYl4l
Kn77xpnQNwTd50fukU4gCpYKBoWGX72VjjP0ihw9VasL+4S25b8XwxO8d5DR
qqLyfjnIQEz8fO8sVRYVLboqo8jodFHc1+7hSeRRjDEBITn373r9TbLbJ/zc
vmRpzvEcM0NuvJKzjlUab6Fnpbp1Xvt8wDxhVorT2LaQ0SZLxTEhphJEc2YG
o1iTNdeeMn6pHoAIT/vx/0EEux6qow0Bl/jL77aTSZJsYr1WmDiybOR35X6V
+klFHTnOSio/1MiB0rTHW1UyLZYkiPkwSToE9rDf1Mrf1e6ykOIw6Ie8j4xE
dnrZZtkArjdawgp5FOXaliwATSw92uYgzbeqHkLQqKNJMOM03gKdjintN1jt
AQqZEzzpC4GYuyRQzLUOY/VhSqRKfyPiNh/7xcrgzUAzLoeUygnP8xjvt8Yb
bZYR7Sz8S4q4kIL78JDsy+XTcV0aS7/MngOlC1ED4/oPBBWoZo6j7cRzIQP/
I0UdEIvhd9frAren1UB/DemzK+lv8SyLjG8KTo6uPIS7oS6ifLiwMfUYziPG
GZTJoeTRwzrO0/K8lOAkjJTcAsOHRsRrEatpX+uuI0ZAqUpJcjV+K/4CpAjk
umnCxySKjyNqC8+5Bvs/k5sTkN0/fNqROYPXu4wc/ByaPJVIvzxDzkHQjkZe
BCPz9UL5FEPpnjqBRMp+ZN78l11AxQjORZByo05oGJnWJ1+IqkpTM/f3IKpa
dJfFwNuG4GxgG62DfU1iVZ49xs5rN275YfADOox8O96K2Rz0GVJXCQHkc9XR
F0oeP+YxOCboiVDJqCtBVjAhK3dZg5jGjdBfzWnVxJx2U/rugbt/Z4Q7Ragz
eAuJ/rjhGPaXUGtsXntE7lvg2GJrbUUlC5y7N5lDOesyPOhaYs+EIGoaqXLE
aGhmu6ZKpyDLxJQPnyy6/ks9vePdqrMxyf5xuOOadsrtw6qAUCeWa6XoO+wa
pSF+lkFir5RHBL1PTYGIa41L444NJJkW1L95aiB5jcVoXwu35lL4g0Ku69Bm
Ssi5cRqj8Hh4GT0m2mzmwymhHwNHSXg8NTn9XtNlBDS7l/6W2KEXbBSs1SIU
yK8g9hYLXhQw8WKsODZS1Gy04l3tP9u0EZG+myNGkmKCgdVYSVOCHGgY1Iqg
5srHU6a2MvyDfzF9vIkl8WH4p3OgO7oT9aKDLjRMUmJwFz0ULfr0wjoeBS49
zQmHC2TL4nPgw0qf3G5EScRayxWq33TahgYbU1mKQVhtBhc79TvvCuqrDja/
i0MATEv8QnKcDinY0WO5pktJU8OVlaRG4wo9HRcL28sMIYubdYwE2b7DM6mt
c+ZP9TxguUb9POzjEHyfYl3i1i4bIlRWUmI2YlWFwV8U6lKD9eEK0EYLZYTn
BWJhdWi2aOsmbV23knnnjq7eEwf5bRyQ13wvgqjETaVkPszZHN26ulTWRaB+
C65mROp2ibNrnfW/gTRlWyVZYD97OonOpG14hyqwe4Cjvsxfb1GQ77qQpDxu
5UKiBSvS80oOvAXe63xIISBjXK7fzXUAtGKvJ65/Tfv+hQvrtPdi/RI20AUr
oa3fG5r3fHgV+jJ88vYZyXhKlmwk34vXElx5pI0A0bhRjaombfR3LmQRpaH/
CbfHH2zIpFyy9dNeNriznYAIuJWxYGTXSSjoQo9C2uQGf9fM2JKj+1kJVaYk
I/c1UzXQMkfMoGpo6HOyk1oHFpVXN/i3/eJkAGzPm9AwOsGlSsBNlESH9PNW
YHQk5j7cSDMsdOVIgyxXiB+eKFsnwp4zvCCsQtkxX4vcs9SRa97+QUM/TMpd
wiSjAXCwsI2QozPVAhO96+kD4/QgO7nsk4U00+HUZ0fjosQSTPu+Fc5VUEMD
zmcF0VUGR0Pw/ZDeqri+hzB2Op5LiPE0nZwxMjACAQbLdSpu0iYWTF7BOkvH
hHkvQLQav2udin/dLRD9Cv0/xiHZpP2W8gZ/o1ueJTpbGDkdCxX0lL6d8Y39
LnxHOr8HVj4KKfYyPiKGSzOVKQ14ZKJJczsZ2F4hwOH980WVDQjtXHeF3wTC
Z4b4B6GfiZlW5OWWLXRlCT5Dd/NBHolwaaeBVMnDAIZqWJ46LdtbmUT1JcDd
cwhgdg9Qnv2+O5TRSXz2PacNuPEsCvyEMa4HM4lZtR1AXp3dWAOmX0sTjdMa
gtkmI2RRBY71VrrIfMpuLF/MJV0RkO9b4tJoBB2GeORu0DKdnu5jNDcgAYA9
Y/HoJ3Yuhu09DqOX8/Ox1kUjgAdB3sQ3/F53l2Y6+hZvb9wsqXIbNPcHLbz7
IHIsa4Am84fM0S8mwideF5/2wU8cqUZnrDQQD8oWommcIdGxGdca7ZYtNO21
tAGPRkLz3BGOSB66EfuB1FeMl9Z0zUcZP0EHR/Bdy5gcg9evArz/dsXWq8Ji
XRHZc9hpNo1Gh8mYj6CAb3B2zkoxTump3yI98ybZxXxMQJqnhAlP0XOYX1N0
mR0LsruF9iC7aiu/ZZGgjzOpI37brwmrrG2GnMmu7QUeJgW0YsmhZog5isNb
AqvvaNDEoSWJVHN3OjujLN7GEuRhuVXpycHCzqgeehZ6amJXMuNWQRC1UG4g
RkH1eploB4UeLN059UpnL2UWTLv2jxHcNnN9SiXdJ2vzFDMmbKlXkOX5q2YV
X3xoLo7cTraTMNd8OFkzHK0K3b8xUV7dfv9laxGGoxarJ9XdT82JQdLv/XtP
4jdRFTf0/0RnAcGj/8CouJNWISzWbKShlTWGW2FqlZGnhkcoo0wPqdAMTsiM
JKNlLsmWGN6MlM4xGpncmMYXJOpgk6h7/WCb0Qg5Gr2dnn28qBKAdY0hVJ9e
097PyJQaqQTC+73QQX3hR2p67enkJ6ZZyNnuKUtGHlGcsG3ZpFSqz25nHAIy
We4YjD1dv6dBUHpQRm8gLaPgOF3GZTidWOSi7qXQHqUfgSXPbkC0blD9OsPW
4ZH70beEV6dsfF1VrEOOYRslun4dJkC4Q6zc7cN3mwraduWM+YmHJya4kx3V
h07SYC59AXrW5FAt8xkUDXJlvWtUM6iaze09TTOc1hxrNsrf3yIWY7eZ8L9e
ilf+9ONkiQp4I+5q2JTkLKLaz1ZQ0tOswBTut6nzp2zq2dTG6ihi0aSDu3ju
+GO07wVgAO0V9kzX/j6mDVbAY4D0ihujF5rE+yme5DFaoui8Prh0V/i4rQfE
/OkMcgUDFXQjzRz/hTOGMa1MKWO6TFmY7Bba1yCNR2Yd8AyU2wLT8ZwhLFtP
lZ9Zxwu/lHNPo61eYCe1+TVyQYVKJ+9/sN3P/3QXUlPFdpB9NWpBjsqpvHhS
IdG/uWscsXjoxJ5XDLAeLQbqVPaUbojaG0GyYou+eB5kR6TVk9sjZRW5WMxX
/4HINlMpYbKsqbBcnGGnJGBe3ZVVExDJvDE/AX9BcC4mFY8ikv1r95z42i6p
htizLF71tpxN2+tQ77jBQcOJsL3IPF6+F+jPOMMgkbiMQml1nUz5IRhKrrG8
Cerjj87l6boXb4W1rYV2WdTD1YgEY6Q5qMW8KePV+xw5M+Qt7M6t7eMyGWwu
k99ZAuXYRq0W03rJ6G3Rgh1RQjOj7ftyLCMgG2ws+22mp21Q7ZnMYtn27g/N
8afssPAq9dK73ish8SJa87WR7rWPWmq2nZARJ7gbqcTNDLzQOsF1BO7gOl+H
lFG4WWmXVd7pilZJgYKNN8xncKMb3T1wXUwUkiG4sdqMW6mp6zX2uqV/4d2U
txiszD9DCaFBw8fwzcHMOCCkWtlNh7XQwimP8patOWYzqxwp+1NwomyxwK/G
Vvo+GeC4QPMLR3IaTXzY47CoNGxim+TnrvcAkIgPW+JfUnkHg8e/mYON9A0G
DJ5DH5SP9Y95Ve4R4j+wI1dAEgYVnBADBrOzhFJ+juSaqQB2WuynyruNZYpb
jIUjd0zIio6s6Su0EQPCxrJq3n13bhIMFLBBzr/WpcWe3r3DYI2Brq77H+JR
iVHUD4hel8mTh7CZJEVd4NznhR2O3W0viiKxQWElRqUb8ZWNxeDZIw/0Noyc
6MtELqlEBzNhAhJ9d672Kz5FM/8pSOcJ5TkDCO25qrRhp3KXzboSoBpuhBNo
RL8DaolgZ2HlGFSU57j7euWP2kalB7rOyD98ZjPvFHzdSiHznlW5g985T0vw
bf/mEAWJ4/8PauWh+VgWjhCEYnGkBscDIePPSqN4zhkP8fuWTgp+HT7y1zi3
yDZlxeVIbw5/go/uqEqheY84VE5UZ+Cd/MyS0snSQa7phpTjrDS9Fko0Rrqg
Hnpblp1tyz6oSAUInsfEdvEXkokYW6x4A4SzZgo8TvjTbBhWCLuA2BqB22vO
Xztkxh/cj3LW/0npKy2BDTZ+x3EzcAbp92tzr4PEkIPHxYPjIahwVhC0ZlNb
7TA2SM3R6/IRfKGz9mBr/7efS6KnY7zz8Zh6RCw21jH8taOoOhkqr0rFwYio
+wYO15/VREVTxGL/x6vvgAMLGZsCRkaolbeCDI1QSvCmmTFJFY7qHTOnnddm
7bqAGtKKQsCg4t4gEE4U7juC2LBg6a1N6uNjcl7eAL8q/iykBcc1pPL+d0TO
0B9v7lt48WGXcCEea0VFik5R3kGL0BI2OzdTXyKxOzcwys+qEFvQpzveBrhJ
RhyY6DQ5sRqkli2EkgQnnJXUDwk+6VqP5PzKPWg3FwvGhCJ52lWBxVJcRWTH
yvxdvUVhHFWcM/bMNQy/bYoWNvW9rDxOcWQYcJfjLxJt8sdkfEyyii7JVDsM
mT++AI9zP2+UmjLGIMVGoTWOCv8xf7NAjrW5iRridJCatUZMukuMdv6aaJaA
bNaW2gLrDHJh+/vlNi5sfb70FAgi5SJyQUQfe59mgNfiGB5ckjHw6yb0tQro
QY9d9XZh7k5edQu9aUHze5lDsErTkJA0hnQf7jCX+bnzhbQ9grE94ILEMMvB
TWJ7rNfXINyFkSOaP0PNtNZRsDzneUH8IWOAuOAUrzPwWiQSQNjcij1vY2C6
n6EX/jk+gEC05t1o22/aXFwXQGCkAzH5Av/57LvTI5A87kY0sbZQHPWeTW+I
K1l94Z5sCCGm/oixkbUWUNbvHi1WVgWysNTA+qnBkfqsqUi5e2eNSBCOlmuU
MK5ol5Iq+yngzamg4+nsuMoW83+fVKJ9V3r3v5knyE8XQ6f/eGYQOuEw6nVu
c33kr/b/MeY9iVCdEmcZpO6u13PpIaT4guXxnPhub/0tjhJ1Da2mo4/gWtTs
QL9CqhxIgl+lWiAYXq7LYU7tzr3ZME5m/53XpTJGhr+6eBC+hLjv1mpqJGd4
jqFno22JRtWt4qPLfyG2KtNm0TsSWy3XsmWAiLYbp7bBaBsQYnsYOoNQqrT+
DA4+ImPXABnNhGrfPLLOtmE37JJNk73KlVWU+cHCE8ogQj2xGputzk+bK2Q8
UA2XAwWmC5Cg7D5rnZhi8FLXA0xRNUc7bKvQAuBlrLgtL2AEKarnbLMrjaq8
mHBw4KSM0m0Z3MBztzpwLWLJsDpHbnb72GEROpt5nFAroMlUF7PC7pLA+K9x
YT2sncLSA9zyszUti+t6waCPbjBNHtyPClWPYnsYiURZapO5pE685ZfxGoY9
xjjPL/v4Ls3vr+I+SCzx77wUI3aaxSTbzgIRSl4b4TmsbNtKTtw4Q5er8F7n
g9nnfeaQzJISc2En2bVDz1OWqEVpVomyzHFnjeEi61lFEoBqzIfR64ViHcCu
zJ6LZAlRKMxHMwF3dgW90j014KuH7Zs1+LScp4ZT4BhdZ6zwjIcz/6mgpv9m
4aSIQUj6DdH5ZvFmB/kA8tEmtQOUncSbLYDtHkT4cHKs/8uhDEEL2zcPWIVa
xuJD1OjI9IKFxrUMK3ftEn6f0S+eeQx0sZOUE58ONJ2uIPEYoOmu7nBM39Tg
PAKpu8i71nqrTo7odJYDMqujzfRZtyxGpyeQYyZsZmrnyq/S/+9Wx/EAld9g
TskIJdRsMtGwRto8Aij28hjHfvscIvaCmDP8KmUBnnZtYhef+vMGujfx+glB
L/ey2G+sm2MloaDmK+52yD3RXXlwss/f8rbGG6hS0HYHK8scqTiLUHGpOgW7
UWCnJ9HrIj/NgdcShfWR5sq105g9SZOTl4ABgSPtAnbhtbtVhxuWfN9TX4RJ
On+K5sSwEOiOdl14O0N07EyH+BiMDu5VPPMlo7868L08HEhwLYwlqDYVzDuA
3Zy5JuCP+6m2vDDhhTMChRkznzWUbJ5WcjSJGG/j3JYqnT+j2hcWHtUKJ3M9
WP6hkDWA/Focm7ohv0NeFh2PEqE+poatYONihMsU82gcFXXozWVg5WYpaNMl
BKLbOEVE4Dryjjv/K2xAs0D0Lwfl/CtLj8CaKKa05VPoDGWFrkleuzR9yPQG
K9wkThK/MOrAwGYiNBrWv5G2Hc3R1J5GoaLBWTBqFsMO7VHTjz961vthWnGJ
OjXc1XvRM6/NXisgBveW2LVLezCACzxgaaJir+xqN33VDPekR+HPKSLHCp7l
RdT6CbMmtmwlPFJePKK6hJw7QvCk0rP537fd+DscjAaOkntcTMCxUj74uybS
ZlojoBH2p+ggGrC4h+Yc912vu2J3rc22jCw5iRcspI6Kdv5OcXqvUrlGsNNA
XV64IBivFShNFUxKk5mPaDPWU/xU02glte7/dyctXJ4OosnaTnBsPtMpiqUr
2LOMM/39rRe0chfPOpdvQoswCuiJpPZ9SwZVOHv8X4+Hn4SBh4Bvk0XLLTpE
6okZeuy6QbXFpqaFU+Dns4fjGsI57RCMoEu8N3dqRVIlq94ZNIviDUiv4Ixt
X/klcR13TDngyl0OW/lvyy8yIy8IxhvKC6oeOtGmRiESZfN904mVYhyPJ4HV
22jqYzXpzRMzSZsW4BdZbMxr2bPsrKAMQ4QD4h73jaLt7iPnSiu8Kiw61M8+
Iud+PZD0hcZ8ElrnIOzqfwARxpXy9ua5t3btFTrfCAZWzurUly+YSRrS/m/s
c2wABMPhsXfgHQduwFPhl5ar1zwBKGBJmmA7rPSwzqcPXZALmB5a4k5JXw1Z
zoIrUrdJ5s5Z0Zceywb63NgLE4rK29A25Z8sPSuvfj4/uExh8lNKP2XKSfnB
IDUhUw8zZLCDCN5guKIPhUjb7eS6N1GVs3sxZOOIY5Flmgj3kBvZ22j/S2uZ
ol8yFZNSb1UQCvSH10gXGLo7KhZJnCWFDmi3dVRupnQenU2E+ized1hZkyQQ
XMKY3e1puBnw4cWo5zkFBJ/FszzblceJ9l4RIEmrTpkLmc8mp2MLWPcEuVrr
kYnDzNA+GACQDMbCWjnZ55mNpeOc4jRU4AJM2KnHaHuFhF2ccZYA6tR72L+Y
jEKIDTqACotZYkbiqQneAQlThEEsLqwGEFV2vqPPFdhnnsVsdcIHt1blZktc
GrOF+TiOsrQAOw6UTg1R59Vv7M0/a1Jo7dZgrI4jN1I0hvu85EPaGyAoowot
XvlyJ77H3JwijwUm1V3WGoZizcDSHoSt7FmP6OxpKvnqTtflW+FFLdbPa2Wf
K7R2dykn1yxgzEyb31JTizR9CgJqwivqg9G0Ps4QDYzqe24qeRn3jtQBHIB+
4NJ5Z60td1RfTlBwWZeuoPz2UaetAjGI4iwmnM6zanPYyBUqu9wLsNOA0RBq
KOpBzotqW7pEVBJE0fWA7TGkSbJ8c0O4094CxORWpM75YRgcX2ePRZO9Gdic
ZxVF0Jls71r8RhHbMKhRoJZUDBSNX6HUGrzj3EiMAq3mNNIRrhjuSQbhh+63
RfVKScgB96tsfXdP39+kOwrvHqvxfx75L4e/ZXkQ5UGF9QuIiRoNQCnA9WFl
PIDFGAV2qKT+jG26vK6uQT33YNsj1Tkg91aW0L20pjXK3I3IwhIJ2ScaoaUl
lL6kHAENyXW76RhyJeR/o62069r4zQMiBblu4DheJdKttlBgk88SpiKkL9+x
w8DysiyWIOZGZWBzWbOfMM1JsbJp/eoQ2meulfxyt1sBE5/KOmGus+QyM6gT
VY6QNlogPdIrAdEWK9QKiYFkzaFfmoNBCXwOVJQ1n/t0VtFq9NJzs6RKyXIZ
ntjhMNbt8sB6HEjhE0sUIlTlSkk90PFH4D5e6BbJBGjoYAvSKF1D/lNmlhpd
z/ijWLt6pHMBT/aVyR940l8njQktcKkMJGjQ0Hk661Y2UaKaIzU3IlxNNtdB
mhLseEo7eBFf5uOX5BDUvpn5EaGBWFaI7FcAEAmbFa8j3tPHTSuHrptX4lAP
VcgqynrgCtOpXtzcmhwSmVPAFti1/0W5iLFof9AaoemT8GhmIRdNYHfRCfen
/v6UCNdmbxbh5EmcspGssLwgyB8CwVJUIadqrhJ+C+AvxOaCe+MzENvTY9jX
t05JDpMIFGgpvsY2u2uHTx8Kwww/4/LcrBKyf7JngtvePnGhEytaG4/VHXOQ
2C06bQK7iC30wCPD1IAo6Omc9h6BN/actM2Efx2c73ZI+qZmlPwpjhagHVIg
TWmeGLJo/UMxke0xQ8D7zrmsIgwxGW0zVo32zkLzBL5tIHd9BG3IL7SW8rqi
B2tCCYoHxZ/UdWjhCeQlPGGcGxSOLamW3DeHfqZN1zDiqDgXt7WGbc8t8ZLn
xaODzSD/nE4ZvcE5zj5OkCj1w0Qt9MaxHdpmwxn5Pxk6u6xMPuG6OOYJw7st
dk5HqJ9GmimRyaiAyd591+swxFbWMQY1nsRskj8ard9TlvSJoldqFKmQJguU
+J+F7bDG0Jtmzh/kzMKWstUap4t/S0EO+iMs7HnK4LyF9xJL6C5qrJ3u5sI6
SOUoMzrEKMxaotDIjgI95uF0iLDEU7pRJBztqCBXZfqDqhmV9Haaa56aZNAt
I1AUHaLY/DIWMFrC/kO+5tWHiiPMu58o8deuEoFO6FI0wsGkoLqh1pByZqez
p9vJB+uDfplCnXC7oncSBe0cJVZaPmJGTK/3Wu7I48n/17MZ/Fvr6kxTOBOc
dk+RDZZ1Xylw4vaw/FrPZIWhbWwwleaeij0Ky0iGqpHoFBsO/Rz49xcxQMfX
zYgwdHx9jtPPBTsDUJk3pS05CHaeQxUlLTSvtD441sVFapujzSLgkzqR5H8t
YC2mwoPe4hZIwKlYpyhLvqo6I1unCKbUPxoCeCMeyDVoFxdC+uS6xkxeAemW
dO4mEjmHaS6jEpWml548iirMacIkdiEcRWJLTAH+6PQcWVcOT6sOhKo2jLwC
3lpZep9dfpLV/bfsUGquV/5vzZPb4AGAo3T9q3pE9YbqkU0b29J1vL06sCBG
5xZ6thHW5Rn4PJdwi7yOTSNglBV3eyBrcLq672fJPE4whdH46ztr6GCzfEHf
UnF+G1ydqmg9eyKx5IhPU0OXC4SjPJAwVwPq+Uin/BhBmOQ3HGRQoc4wp0zd
hwy6md6JjpFB/WSFV/q/lBO3xY4HPnMsanbjYXWkL2WjqhqGknOAWu960Jap
cNSrvBp4ogR/Zc6Mw6HESZ5DBJk69VDd+LvJA2lq//3f77oDUfVHxTOByLWS
mlbiD7x0b6vZ0yhvgPwAUXGOh27jA1A2/TwG5ZVF7bMPcKpYdwJel0pYNprF
GOQLdqUV39mGc6hwQx+OgzN/VbnuR6UGvCaNPW+MT5ddAZP1vjE97P7g6Y9O
sPOT8lRLOBfycQNv/JG6kwrbYjkQaIrpJgje2n7lGO0bxDLfOO21tnhPtzO5
foHs3W6mEYe4rro70Vd68F8W+EQTvYc54eAmfdB3yOOHZMh9wQYdcTO4O6QK
4xdF+WUkVucESxqqlsM6vC2HqfSCAXDw49X1KMpSwtff75xdDxA9hdUUAMfe
ca5XqegsFN9JWiuNIcy2V6gDezqnqUapq5bsSvlkRCe0zB07Au8Y7CgQRniV
xWtKtl8zQ0at5NxXa4rrbwPZF4ynIrxqsWtkwoX2XKVjv9bkXZ7rH+POS0ga
iX3wRpjg7KxlTyw2CxeEbYfSipcVHDvq5egT9zOT2IFtYeiVn6lVX2/yMY5u
8ZUkcl5K61C3y3jYCFFVjSLTek9xGjeUoKi9mj2lzXezbpJe12bcMh57ZXrL
Nq4qotQEzE3bT3xqpaekCx2QpL6ceBOHXNhOL09TllY0E5z+OdtNmUaRaLyB
bzB8uL+henDt4U87KFuvnchHG4cLw1PNxbFI3hiR71tfg1JYragyi/nYOKth
cO1+mSyJQn7B/O5OvyRGDKCJZX+6IT5iK/DuJ8N3kU/804jGK9FCny3tA3gT
YZUcfgv7VciZHWBj2f5cu2eow/65srAPj593rsvI7LMsO2aELV0PlwDXgXHv
Rm4AwhAeTU08KCp+DuP4E/hB78tHoRvK3rJiGGpHEpPaBx6RNdpDf0tPERiG
dA1UGn9sejk2icBFGPxMYj7EO1HM+UpvpUdAk5xX9fLs5oCf8FHhr+7GML/Q
w5hWFyIHAcShhMHb2DbE99HHuCb/9XowaO5vFDAugwPSxtKUc7vq4T41EcIz
RuCXumntTEQP5n4MtdB3SuslWQAGKHsMD9nbY6wmN6RiJrdi44krhM9RQ69U
i2ZHXw4+9edwrvGXHpj6nSiDjwVgb1csSO8gNHWimw/VvnnvBrGD9vAzbF9L
y6i/wZ5/3Lsr4SOEB/ihUlikv6TdMGCzHB/8C3+sK1dJQpf2SYjSHR1AiBis
GwhpypR23qmqIQqeGaVfqPvpTxk0OxjGYpVMe3ST5J/rDQSl2xevHjG4yRQz
HuQeEL2QmJLCJsC+LyZ6IepxIpJgpJznhgV5+TVbBJOnFDHobWtlDGUI6BOW
uI6lBJuAhxmp50nS2Gfft+p0XtA7RR4L3FQC6rmU9L3lllLg1SCMW1lCHgpR
KHCTd5ML5oVCeo8a1CE4FoQa1N90LxYHgT+Qsc8Cp/RtJh7soDhpRPovWPr0
YQ8CuBY6/cGu4eT+OFynk4dnw4T+LMdsOPWQXmZ4PtP4hQyPONr6tlb/EY/v
H3/zKV/A5PFBNjtnvsoWULcrhYkYrdunkX7EqNpdRxLCt7EuP0ZYnZXDzogn
BMvI8JpOWoH0k/JTNMo2cvbfaS1JbAlPy5btQ7aGIh6+rk9tvw4lU4s8O+FC
sHbIVNnKhkjaS/AkHSG6TMJ+9D2Os1bay1Bl8SSqLuBthkQ82+NiA7SHFgbT
tCh/rUSlLj93eEz/Uck9Mau5EjJntA5e4JL4U34MHlYMHAM9d7gs400MPjcg
MPLA1ULphZx/lXRzrDqDIp81p0HpqtWSaqPYdkThmvtdyTmoIOCNVibEPY/b
Bq7SUkFbTg2DnCxSOtYYuFbCEtKHuhiCXGXfZjAmZqxydL+sbpl6vmbVzxJW
vT9be0Dwc5Quj3CjW6GmZmISKCC+S1C8rIPC9XLI6TZXY0mcQJsBybtj1nKw
UUM0fbSguu0u2Z6LiK/Avt31ieHgiKbzgBwaRRjWPhyNI6ZrDub7G45mjzE/
GdOx3CIxvUgC3xaChhljXaAfwbXSjW6mlCv6RGZu3xxA8EpTOnf68sUXmyPh
3LvV5qz7BMo9BzL5ZdMfmVcKg3KXdiY7W4hYcS+Y0Z/e50UREQL7NN8VwFzV
lTDDiNu9A2djPa0X1syJlcC5CNoHVp1D0gdrdh/OZIVyzUd7Xlqu8OvfgtSL
JmaiOhf5GdGRGvPIRIBXXRwhBCEF3mCchvFCwX5jRbi6ulS7seL9dwmfStnV
M3K4RIdcckTbtRgwMrOxz21QK3hf0jI2nlRYTwZ4lyJDmE9w0XpmHJ7OSsnW
+b3v05UtakqdJ2Pu9I7XYOE9Bpvlqf8glP7pFFjq7AvNvxA/IqYdkdIGrrbF
jn0fSt9wWTbQcSn2Y6XFpQvay16UChBJUhy1Ly06zsoSesoEEj6ii8h8XVAh
mP2xa+jq+UfGsOaYBWqwrBGUoYN2oYC5kjNLH0nD7T7MV9qgg2sRq7edN5jF
vLFak01mlDB4uOEnKLR20PWIvg52KS8VNG/kEMqfEnca7ttFYwmbk9REzkFX
hk+bU+eQAFLclgyYkF2QpxGvvhxIbyJWF95RPMC5ndL6Cw5feeb2ypMZz4RG
moY/EY6McsRV9cYeNpPz1P9TT9lDQ680oCj47NHyzxqIa3x9JIhaB7yyO8CY
4VriWkIKa9qAMy0XTQv6s2VrsdcxuJ5RoW4CiA4Bf845MYncBsj4z5xFHXkD
CxwjfpdyD+pmiSW5Ho1E5rVbBd2YYSLZ+koj0bI/ili2qsF7zhdn/vPILmth
gtAZqvlV9q6h1rxVaA08EoMbvYBNY77wbRSYD5puDXIWKvTPz8s6m7ZkIc1S
nh5Lly6Cgq6MZIGSlZfIUU+PJNn7DKu42f/PAboNIltJIkZ0B5N5oxaDZsA/
ExSP1+OB2uruSG3UtVk5Gt27OmnO+aSbFeoBZ9FTZ9PUYBPd9XqdnPdg5TTa
yK6eCWev9ifBuVCS3Jxy0GqZq2dUZye+eqEcElbEY6ftAEZO6Hhdy25LhrRG
pPknw1wj215NRIxVOtBg7qO2SJkC5lkDsyVWoLKR6fI+dZIFoIETtfKGASdh
ouwsFZAHGO8a2UgbxEihIhRkjJ2ZoPzBAeWvi7qrIpplFUSfMU4UPTy+81bh
+Ucf+/FzrLGc+1N9TdC51x1+pYc0YAPMTF/iApkeuNa+r2LmpIltjKWyrMOL
sFHKu2/yOxbUoUHOr+aFciSb9DBnu/zyyxXwwirk6YhoVvhcrweKBFud8yUw
XorGHmpo3ojfRidf63MIU8dXz+0ew0rriiXo2emEXg1Y1qFmSZyocmWGcu8F
ypOljkUmcMoFon2xFi8y/SUWWiv2CgVX1aoOjBWF8Zr4TrThicz1p5L8qtnc
3Aac9IcYKfwBQRR8ZCK3bTTNPqr5sUiKFDkFAUw6xGM3TDMtF5IYG4Vb6+dq
cyVV6bap09a9B5T171p8KJ8KZ0Ub9QhKrsIb5uGIs4Nk7BPzexZsuTHnUF2s
rmPL2zWJ6TFJbu4vKPddHHfbJMGbDFi/Zb9780JWLU2tmFSf0d+wi5akbABF
OJ10gSdpGfQtZk76j8UP9XHC82764Ay92OSZwc2Tq+4Yx+bMvdi4zMyrKx2B
KZGW8Th8BBWET353vwWX7nPayXeF8xdN2oes3jMS4CUHshJmS9bDZD1sUFkr
yFwhIPvEgqCIO3DR6QErYO2ba+tL9T1aHjYZ8xEEHXOrd0gK4StiombvsYV2
1w2U0DWXqZm0lggJT9ffHN8RFXfK+YTntzBWjcJiEtrPb22MJvGsmJCwE8pC
f0KEYmxc/iOf9GlHEnbX+BT7Rxjdiw4v0SJunvx6cCfcqnhnkoehnpEbC0X0
y41PBJvt/49aZS3fSnHtt0LZWJC6pHxoRGH8SL9tFNHE3o4dTPczb0yppOe1
NSp5ffyMWRTd9tZTOWWtfr2mD9p7Ajyj7BCE2QFtrGAr99C76RRTeyvEKV09
gz6Hdt+/tBnPrzhA6A2M1Nx0CYcjt/yqd8QLfNBUOQm6Jx71+Ok2MyCH5uVM
GwxUFzX+pkLwQtjglg0gMvWWAiKOccLBIhjoyLjIS2MhtywRTKmRFHPErINq
EsOnZ42g7dle2EX7VZtcvWpxdYuz79/UtV4xu/M/IXVuF9AGPha3Bl0PpQ3s
fs18FLGjnXrU/4uyHWI1SbNGTH91M5LhtSSrghIGAqo6uPjK8EJ8gnZP6mSv
SgNzJB8+2vyca/ffbghj4CVCJ3fnCmIhHegD92bR11609LqGyZAtykBiCmax
D5nU9ReSk/n7c+3Et4BLAkcZZeWCGEV/hi/ynXnWOu4zFZvcSdSeTLi6Ojxt
zdBNcyWtKvgKUF9KKRCJpSVu83OJ74LMnQKctSrOF4fR7o0ovAZpE7W6jthb
zGmRVJWGHXGfX45l6JjxNLrbNkckr9qLvoaEqu4I4mDQWnWt+LKVj5mje1Ih
FcbONmFMOq2NYDZNU9iDV2kfTWYoMHt7rZDoXiDVqGchOJJlstDKtFpPUU2x
Bm4mugQgK7HaQsf3nUltg15odaIctV/W27z4nJx3I9pwDq76+sd9ErurCwHl
oie06D0GVfkCIMBfyltsE+jyOk+JODkM3oxhHBXXFZ2ybr4wD8EPnXh9ZX3q
Fq98lpW7MuBCin0+BFgeBvJA0Up7IYcxkuTfRz2ghhSwnYnX9QzVEv8zLzgu
XeEUw0/nl4TcHKaqGt4Q9ecxzSQTm8EeLSFEczFMjCh/WlS9aPWw9hOrBUre
9M4YDfA6A7bMs/2gH0XjL7cSYachHz8sl3KlpOv9U4a0vficMJJriXjBDVkS
1WOuiuY/edjtEyOBaRwMEPcZ9PjTzTWI2QGK3KKYBZItiS5veTFySSRepker
65LsEQU8PJlpTXMudEQVF59tTPnJXaZZPVJaS+2MwxbeU8iAVWsiQ23CpBF0
iy+WmTqbxHkdvZCoGwTIViyN4BdzX1f8S/G6V8IzYTYg0LI1AQuiI55jYKx5
G0c7Zdcn/UbUGR8QG84t0egDOVZrgyEUtcFGk2V+eUx441tmOOgAFuboqM4t
IgU8XcL1CWfDUZPPMfSkC5bK26UVnFDGxwhV2wge2KwTK+2vjkCBkl5DcaMp
2jvQ/EZtxhU3jkKMjvkJue5aQNeRd0Y6jGASwmJ4VqUZZ/GeKzDI51D/T69E
B124baNUlrktS6d5eQh4TNDCrKsGmicPyhmq2lWF1D1TM79pIkXpZcGzZBTO
2wsA1WDzz0cwLoTSV3otSYg9ZncTyKY+INR2YxMfmrFj8Egq1476xszVM4cy
5gkvlM4iEkiVg3rAnVogt6U2fDiTNwqDun6V9FJm4u7Lpiu7G7PwcT8or2rV
j1yiWnsZyMhh+ElI2Y9cJ+ZzKzCeLz6McV/Dh4xzBYK7xEJBiYMKvjyRHCMZ
ox/IPzcJuNaOd89KIpzMqkiyy4BVCMAZ1vn7qV6gXEg9IKgY853SM4WbkWDm
3zzVZy/gN6IEY8MJ2s5fy0yV4TVinyLwd3A+RZdGyCQpZLCXx7RLQyGQ4cI9
2t3Iqh5yUTXU16/ezDs7gQWUOzj+ZiYpx/iH75t31uNF8yH/71N3N5F1Io2P
s4oy86wfcxjh1/rPBIqh6BhoquKdgRiYH6rWgY4DmzVkdB0u2NwBvnxyKzrf
rZ1CCpBz8r8o3iexZ2/pNIpNZMwK8Wt3ByE4vsWs1kF3x8H7CMuvQupvF/YS
HK/sqKF9YYg/BEZ4crz9l0MVhR3naeP4sAKgJh/nZt5VPOeHaPLe//PF4jKA
uQHP82IYTZ5FajszX2btXukqDz3uPjlOTtZT7gq30q4noKOfRuhV4ma23gz4
EiJ6pi8purEbVOfJGygMMM19mY9ffEMjjenWQl49jXdm2kCmF7a6L4IU5SeM
9dowB7erQLFPnulJr+dG2IYVnyhKmwDFOzC9YOSiH33pGxk+BrAkBUN6l6bS
MBIXTCdh9vpmba3K1E8AvKx3x7VKqhAQsGnMkHe4gBJxkihmFII3++25kW6Z
N3Im6YhjZdJOZTUpsHvh+GojOycMwKFTaoKkGiZyI3R/4knrr+Yjtjt1EgNd
66zNHEODVs8ph6coPQhZhoYV2FyQH9MFSrgxFIXZ/StCpo/yz5AuElEUG5P4
6pfLtvQmtnCBa7PuNGFj7qA9WD5byPhajcRubR5Ef/6vxvMtbUeD/YnuIHlX
qM+w102BmfZKUfWM8bhKUD223TGjJ+T6YEdWZ8YLPYQVG4GqtS1rQTETVZYM
uP/MIXveP/gQfuxB0dngGpyTsk6Q4T9m2QMYRGT9Iaz9mOkY5mxZAFfHN5Af
NhBgOMQfi4yTIFRCC8VKUMZOVcycfrWTl3f9KNNBt5az3d7hqfLTjnPAvPUA
S0QSWn6eAlHeDTqYDTFB5CBJAM7XSXA8uA209uKjulghVbC2MiLkMzOSOoqp
d/8Df3uYrA6o1/KgoWlcPNNubr2NK8iNTwcPfc973K66hPw0BADEFZZuqFvl
/xtCKHMK6l+xHuJvcmE3eg6U3yTwkxuTLvt1UpAcSGu5HUkZ5OlETE2w69EE
uFWshRRrL/EcxhEJt2Wb1vy5NTRN0TcefT8vuwhQPgU0zwPg3VFk4TG+1scy
AHIIu6Dg0J6k6YeihH6R9H6Bg/EzIGIFFJ399CO00CZ5Nll72B6HEIubsKwd
iPOqnFqlrFX6TBKAbKxCP+AIJG/Xng9h4cPy3OROklqWNKB1r6ianIK95afs
f5R3MtS8QcmmsfDR+NKIlBAZREcNTOiAO0MOs+XOrjYnd1hPZApnrOB/Vsc+
npfEQVLHHw+WMQk6JDrzf4brOWXzh/edYR/jBVt8tLnp9o5UUfhteelxaR5X
/xyl7Isf/X/FOgw3AwYct1K7cXAoWKHmppQpCSXyQOkgUjrAUOZKvnXT9TV+
eH+v5X06VxPj8VeE+wBfUDu9hWg8BjQCKKJjNnM+s6By9biowPiY8NZI8H8+
bRT/UdQY/7/ZzK1HSLU1Y8nfOSG5NwtkWI/yYf/bKmbity9x9RXzx+ro1dql
x/A0EUVx1k8RKf8yaznztOuFjk1TnfJHipKBBplv6D6z85V+67/ISP22f3lk
wIw2CFglwnP5DJmPR/gdHTs6C8PBv8A01GLq9cXbFN3u7MPf4sXwopGOryx3
5uIPO5GlBHHfroWlXCrUCF5PUYx6m4CbSHUohcqFNAPsPUs/Gv/LNx0G3bXU
L/LFsrznTQKE83EeVRyo88xhbMPLHyLbhbToajCtC5fFaVL+yUP75uETAflw
rGcRUnWrT4Lk6b+ZD5pXczQoks9tU1+S5wh5orx1cKe3fdBY0CG5yg/38wvf
WjSB0Anp8lcuzhe6pVJwERSFU5dETDAODfWPGvB37tl7mlBA5oN/yHXjzrqc
Xe0SxNK8ZtOknJuucyQaR9V7qud6F0nJcdfzlCH+LNzJ1rZXxaNCkt7zxsyd
Z7XYkjFywnfU5rPTXlbdFIJrqvS5ZKiINbAsTy5DbRIH82fOiNIQ5uhheYuE
j5ikxPYGarGU06QJw/o/sZygFyb0KUbQKcZLSDkqtkdDDWyf3uC2vAinkpcI
UOVkvrZbTOhSpIDlmef+J1/jPbZaZCcuqAzy4+Hz2lhVixLS+GOarkqSNX4e
5YW3RC75+xbVHZgdAgYgw8iHH4/Igq8fhFCkSCDKBYe3YIuwCjtwCeEMcaJs
LbZjVe8NVL6rWkrXVv7kep6YMkJ+lhirxUq0yf1QnMdsSlWjqPGMPTBJLFwH
jHYSzg+sqAsYwYGO10nhn3nSG7T2rrHCZw6EBOk3w+CSh58rGc+WKLwr1DFZ
u8rIgXzLt3rqZw5GG3ud/DlFDvMu55ZPsuAAzF6m5KYezFK74uzIiqYmcBXs
0lO44ji5ryOb3ahGRQCDObhxDxujIR9UHiQH2ZJPUjGAc19/X98FjEqAor38
r3QO5XXg8xLZl7j5GDZEdpVgBmThVO3uliiDVi/WA8RDD9e07Pqzr47DJXxu
M+Kx7ZADDj4SwVkgJvOWiZAJXukzejWRE3HLjPoqD4zJYUz/ygH8H8b5CKvz
4daMArqF9qcb5TjfeVhICQvgI0Vd8yBWnVtYh8JYuBsgDD5wzWXa7/FxduBD
DrfIspyu1dvJzK3sp9LJjtytczpuWyyRkSu4GmxV3HTmyOdG06WCZz/pS0h5
Qy/+KssMI3QrTKR9IGrMlZHyY5ZqsPcgfCfvaUN9Q2GN4HOXlAWDscVdXoWV
fmpSuE0YJTaHv1nOqN+X+6+c9/BftlT1lowMmcd14eUTR57HIJ5pldVmXLgb
jgxEddJdX9Z0L8knMPBQYlTszYosTRdisVXL0VTBdA1NYmLKeExmqkORKxUm
ootte4HFg9C0kbJYJ2irxVwQU0iTRz5zanW2MHteY3WaVlmyhn3T9CYhJ9Em
fYvK/cgjsOWSRJ1AP6saLQT+VK2N64CQJA+j4JGofVH2eD0NGhcLoChcXqSg
CcxSpGpyp4R2RjPCloVlH4e9ncJsq9kbtIT+6ht0UUbMeAs4XCEQ5nc0edPQ
8Pf6js7KZ6dz0jV38zTr7uFffeDECwec0sDJH6eIH2uKwrsr6HnnRGEpIjO6
P5kNWkEoK8LnS3QUdfeANffuqHr45AgQ+vHLdW3G0Ln4IW+rk9hpmJXaXXrq
tVA8fOteThKC2+q4YjTDw2tUDMDogDJgn/04aRUEsp8Nx+vvhnigVbRzq50S
9GMqZxj81oNZjJelDnHe9Krg4X22aQM1+Cw69mASw7I7pD4m3V3Q4aPF3F53
OCGTB/zKl3V/Q/5NNRKSBKkCOc3U1qEnQ97+8vS5Bd4difrwvCzKp+mebP6S
36sjEIzFRTn+F2rx/S9LcRwohYjvK0AZ7haiLgsUz1eTgHB771sKT/LdCuvC
b7FpLAfOIGGhma/Za4Ug5GLIv1a46F/xPJm8hVT0ya3WsENJR6+ddCDCuF6J
aCbPtdfYLkj9ez4soXYurZcn34/RGKxDspq791EG5jr7I6yNgmuyQwCZ4XDS
rf7H7IdWnGNpELjQU6LAPi/JirRgW3DCNB6pkvO9bjamG/E/wVLKBc6k0/C3
dz/SW2bepON9AJd63DtMs1xtsH9LSe9pKIfS5iebhLdCrUOzxtkvLJ7gvEBv
VbIC6votYGO9qdso6AJlTOA2vDY2mUMknHGCTzIerbef164E96M9947qW5Ql
URk/jy0rwGwKzXWf3uN8gGI/7lgRok08rqD3Xr2BAhPFoOINPjWa0cXBytIc
U+WUFU9XGp8aw32sUgnxuHcBhsG3/PtM4hzYgNYtroWsBItG8K+WXuVG1zXX
fZIJ5mJb71zda04eplbWyq7n6MqPNvFhf1TkDojCyx6TczxVIoXkifrD1bO4
jieW8vSwTDVG0nhaRZA+mLr7nnsylqOfixsPvaiQ2Uz4VcIMc/FIXvE9i1vO
fCjob6oyEWti7HFC81HLs4oV3Gtv7seKgCuE0o2ZGH2ZKCDl8Hc5PeM4oz5q
dPPqlU7LIvTUb8aSSH6qjw/NigQYhW4maAD2MOta5JN3DUl6ZAEnhHOeQUkP
3w/IVrMizrK+OQaN9euTlBXO1H4+DOIkxTd26uUcaVoOLSNMuN9HLCln+3eJ
MOUPyRQF77mbs9VzMlb0je0WK0RgjXkx2xv63SF2bDPiVN+zMTZsjfOia4qK
3WKbgBHH16zePZeBGElllujpZfFyyWeUD5hUf/zuSXxWBG0184BpAogO+F/l
BdHtMZa9Gb7cEn4NMxWKECZYMGSY3o6OicjEpVAEmJh1Hecyl6MQl9JEkBd+
BHftNPkOPVIXEclDzrAqqU5+CWrN0JrpuP7UzQ3aq7B0xwKLsxc6XFq5mJVN
2s85GVRYErH6sQK6zzKYRo2da0zPYDDwET41wCxfYyt7F1xVkXVeJMNmiaXS
0SFm1BuGH0fk6XNNbSpRcbhRajgEPpeQyZ0zCSM3Th9oqhbgGyYwk6QV+lfx
g8MoFiZ+H8D9a9Y83WYubS48R5+8O89EmgSptvaJKs6MoHY8FnToGT4OetiI
TrCH6Y8G/y0CWHXT8ILLNsWUU/ElNnMXs/Uz95Vco8aUES0TPXwiKxUa6N0F
YZ7uuv/UrFRP1w/FS0cSHHvxVaqvWwVCH1QwoBxOFDpxACMBRwDTj7sssJXT
7hlPEhldTHNfU0/elAb1ODt9mC0s09nXghW+GibE5DZUifUWrxeomBF/y2+0
Uw0UgzIuKXheJ3qhZQ5EAFVqt/qLtN5wXoxWwQLL2Cly7gZgRGYIfZWAlMHP
mBuSx44rXC6eyv3C0WmqOgtg2ghkOANoHLvq+9bv2r6NFdkRTd7H5rg2DSbP
rsfKbyOrDXXaw7hY2lN0SEWEb/seeVMKMwhNbNwEu3WXNKDYiqU68Z4kUYpV
2DTXcMXBaCpVAxw+iPcmvWM+MNv5lWEIbQIR8mm2HbvbxTsD59uMgRQGb9sO
/cMg/WC+fEvXjGQ8yE7ApGczBAQmbSUd5JgBEsWU+Mg0fJtglyxwekuWwuNN
0JggEkFYXAR07AKRHmoWYXwCwQQ9gEye+Mffh2FmwI/GPH7xttS2QYTHNd7f
FOu4i8yGcWAzD7xedqlCojUMuEcao/peiX2T8u8EIjoulnEdrCz+fjxzx/ab
cdxSBC9zDTzuOvAcrNjIiLg5+Er1Cu4TIYzzmBDkriYdhcayR4VT9EgF5jFM
qXUfOH/ozp4nsLaKtrypzi9KvW+Pkoc9mXdBgPp8c/RfMsxVvL232cZxxmTT
GfbXplupMLGV0FBqSFcbpY5Sj39DdjpqEeIAeOBPMe6CAmZ6hmp7Vm5W0MfV
FDjeRIVeSLCdtDhDy4cbIOJYGy7+ieWcG16Q1L3HN0cH/QETvI8nC6Lf0fBn
Rb+x7AxyVndY5qAQtUT+qZBMwnNVr1k6HjI3yDwgskbMlPIdarfrwD6ygISg
ukBHaWGLyurJtMTX0bcFB3Wq++ujEopPQ/wC2D52UGkyr/nvmr8S+5piJ7xu
auU7DubLPIBJFWlSUkOHzh51rm3UmpsUZgeoFlmpSsog78/O6fx+vkBxkBBy
DIb828H5pXMeWKMVyH3QfJ7NevtbCMi/fwIXGrtYSQ98kwKEOOeQGjWccW1r
6uVX9KTTLS0uJaand1S+AqwUZqh7rkkv0qZAWfUJA7/A/6dMqdyknqSXRaVV
Q/1qRPWfl+Rwc/35ZD/skKhGzPSAog/egHEKJMjp/Lgr5Llgvg28yhw0Yewy
+yTen+qUBpPoTkjgK/0/qDf1yHZ4kTuoZwnUORALuABruAsBA0/27p08x4vs
xKdU+/MuabjZLeuBIfjhLF8YDJDBdYk46DVo7oPsSPsVhbU56u+Jdr5XPCLj
Nkvq4NS01eRf+CKLLi3ulPem5IU518aNC7I/mqoi0y43Fh/Gb6q18f9RPYJ1
sejmM0nySeT98bpEGfzY6UIQNU7X0NoVFg/MPQuoueiJnuW3iTuFDQ0G9ff+
NLoTr54FvHWIxQ6RatsyJiLuPxNUq0dlgFQDLJtynPwuVQ/VvQSBrFwINA3x
bTwM/EO7xzadTEXnd3tFNptGJAA5gd8qFfl5s+KVvMr6llj6QAARuqxhdya7
RMOzaiVOVt+Qf7NhJHJXKAQu5GT/us+Vk/FHmozcViJOg0b0m6DhvQgLI1tk
V9XGJMC90LP2bzGPxR+px2rnu3sxIfi/1vY+agPZdjAIk6iuz7oJI5wOrEeA
vYpqgOX4U/my0S88JpKOazDSGuWeCvvww3J5CtyaOjYTbK6hkf1KRps6SNee
2zZCkKPd9Gem7uSLmKp0W+qUxGHHB2YuP/LhCUWvbctID3XIuHdfNCvjoYzC
ILxHe7Md09wZWFK+HKU5J6RmQcIfM/OynFmvBfzxDqkUzsBazPEUYDvy+Ol+
6nhWsRq7ksDNSz4PSdcV/+bkcCFoySCWVyfXCxi1Jb9niQTNF5ulAyMPla/R
3saavBDlnSWOXlqYqXARyJpS9R47Q36SBE+fi7eT+Bb5Ggf05oeJ1KsDzqCK
ch9L/MIxfD6XImyxOlsJSNvYTnIKiMwG1sFbQxp12CY3t7p9T9vKnx9TP2cu
dNiBCnecQb81yOrN2V1nf8vp7Cvv5huK5RhfUHMupD1fF+4OjDkElRIc0Gbn
LmXe0vXmm0v3aD4xNK3iCDfB3qXKVKd5jKw0k3PjH5WHP19OO4OAc3sJbzc3
fkLhFK2Na5dOoPA5YQGU3J3GRsXoY6h19FN0tP0pFM3g6fqjLh3atKCBZcud
vmYbNm2nTM1LRtGdADZGZ8I4MXRag69ryE+a6ZNwp/DOfcxMCdDgKHrb5Ukh
S8vj+SlbisteUuMwyT/cCMkJKGoRgIUys5WkKrW1uS+EjPpExHBldgpHVQrt
eD40Rrx9PV6rxMsnlpq2F9aIAM7p3PmsscCUAWQ8RD3ZwFswrYYrIk0ZkGiJ
F6xTdRldCsDScL/4AONyURMSFi5bF9DPQI/MqKN/SwSbzp2mIPzrV/Zkfmxf
67Rm+2gaK2MMAGcYzyZZ2O/iRgQrAQClP7Gr/3N4EjfvHcuWFt6leOAscuzm
WWl5RbA9UJHzVYV8w06Q45GPfQZ9qLsVnA8DTP6V+5dlkifnmxewshyMuRZF
j0xtLG8RVOjKGP2Tw1jRTLWV9l525XdDNbN8h/oFmeN2ELcQGdNFqY1U+V9P
GOrErzTJ6n6OnDpDJsBhryj8KqvVdesIfPReXbYk9/USK2OKhbcx9+330BtJ
vWkkkORd2erByWodEZFucTmYcL/KChILEVcU9nFqmOerLrk9I/49Ita0Ttvc
jN2uftRP0pyj/5aJJOShjdd8tcb9joQgZ8kqHCJvT0ScBpMJ2lDWyo+/DJ4n
2mO73Fbj1TkBgBOE2aUUDVTQPBvsfCqGzWBEL2Gh/Bc2yRopOGyONvEPaGbh
2fujwX0oergohALnRs2W6Vs4BtmrdpLHVqqE/Hh3q35KOsF9zcywhArFZkFX
fTJ/wKECOesPMpsu5lYou9qewTJK9fWSsZtMzJ8euHDojAIdFmrkBfhhL+BZ
0M8M2GC5K0AtSmxfnATeftL4e0uSshRPp3UU4r6v2oHcYI2CjTscANXGr5HI
oc9P46eft1kXQPNl/0HRhE2fknJKEyHN6LZglc+2g2hlGKj+ig3l6QiiBaZM
Jt/gJdTBsSh+8XAdVOyIlVq9EirbZxwl+AnR4jkhR+aqLr14n4lB0ayf7Yoc
Y+NN782vUUSam7hnfde2+HkReSKhOWEXVqwWrdbhUB8aMjVOGhuMOsvTdwhD
GmgC71AnmxakY7zlq+wHMQ7fqPJDkEribnk5pso9jbF3d0L73BPbRGhLXVQa
DBlBUsVOzK5QQA1ikHe1oA2weOAqfqqK18nv/NRvv9wzFJdc8R72H1G5nN++
qYIvhPaNWPhht3jUpAxKEB8FzuPwT3LVpyl2vegAvJFkSxxhE6w1Mg0ziJeL
SelhD68VQeIdDEUtfm/EGyk5rH0G5RnK1etqMM2gGO/sT1CNS6RvEbrICV9l
VzxOJVM1g3NAV9n/k07StHUMSPs69wwg03FE7tsaUraacLflRH6J7/votGTd
y/2/pWfY/fvpuvJi/do9dgXni86um2xnZBHr9S1S6CRiDqIBL4bLi/Amezkt
hByTfiqXfwOMJjdhErhOpPaHV15bktya1KgtxAn1meVAKOgvwFc8yIkp7G+q
7ljw8Q3RzKbxGuinkC1AKB+XBsU3e/6SIdIacn1hhWBT9zQncKPKgfJh3GAR
ZM+Uc5M1LGaDchfjeECxM44BgLmAfPS+EkKRSkpjFhRA8bziVS/D+p1NmBJC
S4Mq+EeO9qcicrBU/cUIKfsLZ/p0KsLD3VPRGkAHbJWICe51//krHhCGYjQX
sHyPWTfUCkdJa/RSllTh95ARn26BkhBadkkx/c889NVxi3lOPoODXOEWD0CM
Pmy9VBhRDniNyuu2jTorqmH0HL+PYemBlbR6xE3rqO7HO1ePNhk6GTMXbI37
ZmPX6tm90cbQbGNl8MO68JOFLYSTb7xQnTYXkl9TskfjcDSVtcek3G6XDpPN
SLPDsVLi9mf7vyBdYg0HaVoXhj1CYQUSqflyOz7lGGyNcvS02ONuSHTXHTNS
Q2iwc23G3Z92te7iJQsxb3MKmMaG/GglCVNMuiB3I1xTZu+QxNYXZWrTBJZl
i5PkJeuAM7aOFYH6MfA+okt/9c95Mhv7tge2+zNmDev7W2/CnqBEH/kVVDCO
bRAXDpIrwiUushv/Qckz6Imoqrq+gzf2m6dr2ZrIsUG6EDmelYSlubw2QF2a
df95wFjZUmaQA6DJn5VrZBAsvOgwAhNiShVZRRI/0UOXPmi6CwH5/wmO/fuF
A7Fsethojfgr3cu+3hQF8IisEAvQ8UKqiQA6qwzn8zPGUJH2xYgcTyYE0xt8
XWKwJSG+NT+xnZH0v2K7r/Z9XlTdVntdBNNXMOWYrXP+xJUpL9fh2yGyQtmp
faefk+zyYuElQHKuuIoTT3sCrpAHFnwBtaQdklUCl5pNZAh39rlWXzK3PuT2
wU7cTLhVJYSAwe8D40i6sQeRfozgFiCx4LLuO9O8rOmjEizs1SZkNhi15IkM
2SYyJnBrZ5EmVFWl49GvCLf7cW5VODBQFS6QheARFig4KHaYPWKhv+g1aw/p
nypvZRW+yRr153nU5RhPbEURWKN/LSh2VBL0aqNRgEp7kqunWlH8Y7OTXmaD
AexsclkOf9BmOvZ+Jn42+g3G/UtHw3DfABhhDakcUzmnJL3rzs1prPgbmFWE
ND5n5zohOR1UVWO7cmhInE8IU0cU+Iaiuf8iF1+3JX2H+p45ztAAx5l68WN5
fVybibmpyKQDhj6VNjbMKawZFsVIkWjAZd687UE5SzWjZh7hEqtEKbuWvgWS
mFtEXql8VIIu5EIjgsO4r1lGqqO4ei2x0xRgnX5SC4/xRoXIlPiQqSdHFiOn
kPxgMyg/IkS8jsYPnnQk2PggEjrCrCvX5YWczhBMvujMbE4lo167XA+VI6Y3
9uJxiz6oEVYso7JajOD+EntWbCENnm3nx1djhtL0Kx/J9KKCYJtf6SD+s9n3
HcKBF2z3GLuY7h3ZDbyOo0hjrnMBD0fGmHiO6jZ/tQG73Ha7QTAHqJ/0lCP3
KkCqmEatwZC4WZG/7oMD+5uZHrLgM+W00QBP8zkIIj75F2M+JMDpW3dVIrm9
U12tOvylFwNJT+54V8AnSe8JoZFN+oPRJSDIzeFigKRwfhAY5PVNOulcw/89
nnUNl/2f2ErbIQSarZq2S07II+x+BEG+ftJlf7wXDEC5bIdXOZTo2Cvp4Dxa
zRTx2uiVoWFaG+fNJUB557Q1ETJXveS1fUYaIzFBPc/tnfAEpDyB906mrl1j
HIIftxIa/tjRIRol/t3oNWmwmLJgdrDkoUVtKRrW/vMMzswnDX3Ha50B87YU
r8lIyFO49pYTRqOo/G83KOkr0qAmKFI7xR470++qY2XWNQyOc5s7MyeqgE/q
l2lSkkKrsUdPWpGqD7WXeIa3Y3J0gMW2PaIRO2bycne7ktNDwLbQTX9bTsTg
SjOcapJ1EtQoiwk/pyZ6H0/AzgKwgyBRwgC0pAFBcILvS3MznU4Xd0prRXwP
rtyfNq+bZzTpYauAndJmNJ6i6CdtKV9zBOjt3PUgQizCqwAkICwXFz5vWUVc
YEPRZFMjmmgGWkujOmGNLe2YDlKlXuFqzgphGrUAz2F+Not1/kIMN9EI4dwb
VmuCKt+ikqhN1hazoM6i2O5qlIf8LbcrjPTELhp5Fp3BfqsXegjCVN5yd5Uw
vVMQtyultDFCqiBvYjSeyFAx9jWKjuP+TKWzvxxWHCNooloMBUZR60pFzmf3
Tw8vQqFJ/SH49Ob7e3ahWQdCF/RaYKRpV+OkUrpQtke5OLB7GY7Iwx9T1s8X
4+5bKI5ARHUi5RfeZ/e3jyS/VbNnim7kNVsII7XvFLbTeSEhmkd5bJ/znwBz
TzC4jIGAx063RFCgs2Wgg4myvvJfI19HnKwp144MdwbV9oAze0V2LMWYWSPI
9MV+5m5L36qK5rwsZ47mCw2wWt2SbCXxuQGu1jOPiohuxOjEB7dMZ9Fi+wFv
myKaQUIih6UhemW5yGx9niTb5Jwr5SFAScJZ4NL1Mq6E0ORfNDZKFrAmIp+P
72ag1tIW7mqrGDINRJ6rDEvAfNB8o7f3E8I54gea08zxLQYApbUEmuFvhjup
x5EilqIFA6PooAFfKbOP1Rb6oxAlVgvIdIccwr0luW4blVQYKG2Vcp6tmz6f
gC0FtTb0Vp8hBGN5KOF37lsHs020/aTDau5C4ZJNzaIKup5S8R4F/mvsx8eg
Hz50Ck2XE4z75CJzW1R1YIwDXq/99rxLiaxoesvNK4Dkmwg/4WlwlpdnNSfE
zb9emrFxJmO5mYKAHWCLuLY2Hp/8XtRMw6N1b2M8KqnadxRzpIqnEv9qFAH6
ZDgXtTrse91gjei7kg1vZGvE21hAs2WgvKgjQdoSZ08s9Ue8YckjtwY7Iawi
KVyGtouDk2c/c2Z8OvcDdNFfdhv+rev+jOI1ghpKMSHPFZJJxmGSTB/pMVey
syWRmifcLusEcfuMAw2xojMPEraZFmY74lPloouq9U3yt4w6YjxmwleIg8Fh
/q/vGD0hOTY1Fsbbu96sc6FLkrsngY4GJ2VhmxZafGoDwLXq32SlzIUWPJs5
gQltKQ3QNMQ7cRx10zgolehI81mtTGtJONjdwoRkxKcwwCkTOru7F0qQfAgT
9q0gOWeAFVwF3XxHDzGlbZ5oGFqFNfte9MiBnImsZxEDzU5tMVbizMXnROkP
eEI+PLxcG6OH5Ke0aTlu8/mr3ZHueVSv4+IYOExwfgpQlXkZAE4k4aecyeIp
W7c788DHELv7X7NYV6f6ZCQsbJ2ZS0plMdB6OUcU/21lNzEpreqI+9vxyl4l
q7OtsCk+WZC3XF/SjsjPo7IxHHBJz8BeOu2fCjItfJ1hIrpV7ZY8LTj/fb4U
fTMQqTZ/EnPLMr1TpOxOnPoAcOYd4eRB6wiqV56CQRWEJCeJULkNvo+U3bau
f64cNX5bXtLxMnaejI8ozkEK/fyLB1kgYW8ds5bEtlMn+DIxGyUr6HSnSSiD
AiK3jGdcrttFHrP7AQhZL35iGMnJnfGXtvDcfCxDkzi5IMultRz5sk9rBF01
jOsCHkYEnMS/0YUUblcuuHDlv3T8fDg0G4/HzoKvt+UtNY+QJgDWSPcQNqmB
KUUu0cnvcic1bQeVfE+6pKPllwgdJImisCiO343EKXcaUmBwPX3zwzKzTH47
iiV0TZaLq1wL+nYgfq9mJF+iP2pVbdK0en2bHzY+GvN0s4gOCcMloz9+8wed
ZHVMKvpOcpHhlPeW6jUfLGvLs0q8NAx/cVvt1PVc4Y08WQt7Vo1Q2XCj/QNe
PQ7c8LBlOhYuOnMt4fmbE+UQRi5eyfDmigte6XUen87TQ/ZIySktcI+mtVdn
vj/yWeq07/4j/FS2IzVKTSplJdBwxAMz/7BIE/Q61xAsOiwUn2+Va22FKSmi
2Y0tqyQfb9sieG1gF1U7rz3vatVumqBVQRqQk1G+GIoCL2GXJ/6h/HMLN0WX
mIADcmwGbp7ta/n4Lu/okOYnwnrq8NH3hsar+KV/9X+S7bWyqC8xkDRSt61r
AkRXb5CjKXOzTknh2LqBul2lCNmGP+bqw2xWBJZ4kPQaKOmyxDysVIZy/LfL
/EQNdtxjl3vyprJLTOiWo7y4CL7SzU+Ub9S3yAd20mi45P63cdUWg8nD6i5k
8sbkPXxsyDkxdtYPWeaZFPHe/6Ye6Xdmw1w4f5E03wYDelyIwk3AJLSdtwEA
D40wTV4xulbJ+zk/xntvGnx5d6N3dtIs4KUNaM1XKbkQZqzy1c5Th3R0BGpv
rzmuhlxCJyfze+ePa19UBLZ/V8TOWFIgyC2+CLcylmJ2iZKjry46juC4WCVu
FPmc3F09F/iaMy4ytFyGmprT/RNb9vCBMpBvMnsGnFy/0ARecAArwguI50Tm
wpQ0xiVs7PWysL+menv5D8y0GmOQ7XbzvprztttXj5y9zv7TJM/dIKV1dbnH
uK5Q+3LvoP4iYHUrqeoQkop7TiDr29d/fOO4Y6xxzMmCnKZWjL9S/GlZ23AY
MmxLYPb/Heqq4xsrtk1Xeng7EqtaBqH29ed6uYzgNr9TCrbbaMjXRJVgfHe4
VZCxAGePaV0zSMUD8+nLucgMqf/9F927NfnElZxz4iMxnsMYhrTVOoMENPHU
QDjQ7AnXzmvEkS0efoYNVpNUaJUHTehJJzELaG6Y31aMJhsVa+3dlwqYp2Z1
pzSEZ5x6pKs9ucA8G3nC0a2Tzr0TC7y6rUnYw8RiWcHXP7CejPnkaOygRiRK
XzvL2J1PVAT70neqtOALCxivz8CpaoTd83yJr21It6HW+ahiH04io5ioIz22
qS7IvWbJRJodcu667BJbCREvU3ur6faiL0AdydLiCEser4+AYoM1OMpwiaFP
+EL6ZKWX1RxmQHs2f2BVMEIcyoSAB0e+EpeR91QIlDDlPwIRCWRF945NqjAM
LtdfXLke1GI/cIeSY4KR//+IHP3vfXDcIhUgY7k5qeGhLKd0N9DL+i86ZXVA
Lx1kkQ1eU4/OP3AlIM9J1RQX1a84eVO+HnILwVL3+IzIZhOuSpDjGVq3lLS6
xzVSGmqkkbeTaOt8K1FkaD6FwBwd/cRRTLgk9+Xa8GggPceEA4qvb2FPjP/c
TyAwNPv3EKffNj485EHHIPRkbYLj4QOf/ug7U/c1S/cfOdYNIvoNc/elmGov
6pFIbZR94sr8bfaEQ0ML4pwPc8PozghsffOIJ97f5IGjhw8ncEhy0yXSCyMO
Z6MFtSnKOVVbURcX+ySFpRpMcFH8BflJtHNxwZ8Aa/jwuMdjGkRcoSGsreJM
t9j5yDU12V9Yba1H8jrkmle51X3WXmN0kV8boGnPOtYf0YVVH4q6gblvwJo3
KeOjpicyMcp5XT3KYXGyxIeA4yhjYOvqjyzJ/QLSg7jkZuV63cz5M1RST0WS
yOycfWXXibcMTiCeyu5yKBzT47oT0KrUEQLeRxpQWWKYC6PRRnSyFvts/Ss5
pU4QTc+yXasUU+yHAuCROT1T+5mbpw9ib0P0kcYY6PQtpdu1NOZnNnXMjW+0
65LcNnhF3r4/CB+yWdnaR1hXMD7dXJKGpQP0Hs8z6zO63RTXYRyL47v3LVxN
YTrdWeiJbAwU7Dld+gOB937CreQUMnO4mPG0ysTyjuFoL7esK4deK2w3Q+9E
P1xIqLfPD4zwE64XE+MeNBpIY8Hit5aFgZ1wR9W8Oe1qpIiO6bs7kMJgyQ6C
EeIebsAJbcviWf58XZcqGZjs/0RCBoRyDTiIRO69g/9CZXZZGn3leQfekkac
+rj8YUZJ8L5M+zUUV+P9K5X7DRBudgio+iP2WW7blZRCdM0bdK7lFQw5bus+
fXdJeQ25vIoc9VVpY+pl+nEfpR3jQBGftCkfuGVW3zhob9TiH7izJUItVgyy
IhXPY1b+PePpV6Y4f7L4cdFif8BqoXpYMDzoOe+kCZd/gnxLvry78qfNCgBn
uORjzfCxHKy/KmPV7TLps5sokwQfl4pob7ii62J8AWNdPenKFPzHduKxJfYW
ALB4TGR86+pGlbY8TrgHh50NSmbQ2y4n6Du2scMvzYluNEdpnn6lzDxECJOb
GtokZClAxK/5dz+8NNCkHQnFwTskn612UB2oCBKY4AjO4d+GQYSw0QgFJgBK
+EyMdMCmvcz+5wToX/vM7u5QXcWHBCFYvLw9+7XSzr1eVEGfatOaXWK9eXeE
CDUjAtzuvsg3Vj/fh8rBQPbtg3zSRuJgVs6eXM2KdkRG75vy7Cm3gvQCL8CF
/eu6QJgcQUXECRKfzIShfmaYf8htkGXdmzvB/OqumPU6GUsTFVr8hDHUWgh2
8gW1Uc+1oz/GypsWYv+NZicmgXHXNklmOewGXGj2b7EAiVsNmfOm1k9fBONy
1y/CxonAjXZ1qcAf8pnhWwtKaRufAwZc5b2zIDZfliTs2X52yP7H/jphhGGi
V+n0dD4AA38Dk6K+e3Ie8HcMX5akV/RWiLCxgfTLfUzpkNkeZ+BwgRs4V1h+
sX+SQpKpdIQB8gnt1K4SmhjzISnq7/OtpY+756DKd3zAdpFD8Rwe2twyEFRD
vHQP+OqlRgoryrJTvt1GYYMBNp4yd6d5i/3Ve2U2IdRzK/s3/ppruvoUeZQt
Rf5+f4fOVlc/VCn3MyVNVbfp9L0BhmRJugnCj0NTX2FXQkmYIin84+JO4cQx
HMwr9I8lC7zTM8Mhk9bux9nb34q8/7Tj2+Ayxsm/NsD+YuokSFUlfIoTw9ir
BGUQS2oce5JSQ/wlWJJj/1mWwN193gJNuNdxaFYxjwXcHMWs5dW5GZBlnIL+
5ciyZNm5YvqOc2+L7tjJmGZ9B1RY1kil4E6PLqMfPLMYqL+XI3GajCiq4t4A
PqyDzNczjSkOYLj1NlLk4biOfrvnIUGK9RxZOx5YBTbH8lrQ3t54meMKxHlI
ExqpCz4DWsmQJh904G8BFKGI0Wo+rX0Vsth2p6dfXwtMWYQfIqhUHi7E4ZM9
ljSmBJ6Ls8O5ZkVruDocakZ1yqmbSEudk8tBACjuI9+aCVMX9PDxAAcRCOLr
iWPxRroakuFOMIceNFIK6UFGs1wzYoVY6WuijfjMQG2g6dXppDQrPQzfzUiP
TSnptxlAt0Q6xotwMZLSU79EKLrKSnJ7eNw9rlZvNwDP1DFX2sIz4l/BkRzi
4kT7lTCkK4bNq/J8RrAUHBrEqQ3X8/P59z6OOlBTybElOf1OB4rsfyH9+vWi
e/R3/9dORykoAMuuY+xwlp3/mMl48aSQjvicXCjGnUQLevqFXLgdsRPBbCjR
8yOt5whMu4ecFQ6zCtw7U/NvZ++5nv6VTgzjddzvr6daNAwPgs5Wyd2mIr/Q
zCQ5JI9QUalV/GxV+rRnphGRSa4vCRq7UbXjkwp0Y80sCh3wlIaObQw+IKfT
rvRdQpbiUxnZIc7IKsPvG9yy7h3OBPZmObi/WNODCbXbr9BSLNdHKUCJ1IYX
HqfjmgZc9Zu7+Gf6OPduZUqbL+fTnX3VrTiJUgwITHstf1h808e4Qk1OMFw+
rCD8NfB4e1moVPeUgMfJCJFsQsQLw4n2v7kDSfMQdkHEME2ZM1M5kyC9cL3B
GN+BN9SISJrA1EBOlAlyKTlgePkc7KJBdyyI4SggyLV7WE7powlX6EjEczFu
FWD1/wPqmLn2QGcRD4UV1DGuXMpNI671R6SXT3VgMR4CT80RdNtCpQi8+Vew
xhtqK14o4isiyvNNM93MWZs10Sr8vJva/biI3Qxw1jvILyRdG2vZie95MPq7
L2/cl5NLb1XFXZu+dVH45cQiACl+UviFD0fIPwkIMISSBjCtXwT0ti2ZPtOR
XVaGr3IZqWsiPeh0DEcLP1kJ7A8vT5iS3JPbhhvrotRmFMMq7ZcDJHqrdl/T
3dlY00SXWlgNPjZ1/BfCVLQPZOFXja9KuYHSzv9OJE4kFpru74p2HTqa9ToA
OKW07ItOgd7vkLtRMKCA7h7oThcw+2vnOgMJreavF19yK214fP77S7GCd/73
LKKulymBc6QIWVhNrRwqxW5btrvmwhcMJa8cB4ZJQEtoif9n5XVWR5b0Xeo1
3OZ1edjHPPc/A931MSWT4EI4JgTrOadgXK7+hjmdoANrZkltqi69DsU/0lnL
qlxWOAq1QIaWA+LPYtVkt3xoZUqbmVQITqO1CHQZaKXjw7lrLlckPWYurC16
bo4HVi5bPuG2WMm3bV7zrEBygvt46p7iFeAeQCqGXQuxQqFBdP3+AjKm2DVD
CD9BXxOQ8oi0mvNy6gWINk6z8UBlJ+QxtLI6nC0S9E9WK54MOb1F2uj5gZi/
VhGqiifPLeLztcN0KyZcCjS3Rc/NkGS/f7WovsgmBFKyMOzszzK1A2zduxi2
5/2Gh9bGKbu3UJnc1E8f6DJM7poC/39AByU/MO99hJr61qrAEngFlEvNaRHH
JPa7kkyTmU7QyzGIoYxPzgSXLi5W3RrBQIA24C927AZj2qR0yk1PTdPmkwXF
IQdDNOwFBJzdE4wcFJ+fhgNrwkw5sC++acfmZkMddZOmK5LnMvjdCdffYEs5
qJ20JVZ34ou8RdM9IS7x0bH64sHoTXjnYyTOzsIM7t73I/7Okeu1PzcEL1yO
R64avIatqAlx9uDbeua9d/jkhKHVVSOAHXlOtu98gC2hFy7fHVcFYZCgljsK
rFhbwdfXNVZk/jG3V2KBEo9cul+wJmQclBToiXhxhQ8GfS9ZJn9x5/RXVPvJ
hmFgdQizoL/mWN2qcMi49ug+h/XKtCfx2Wvjl/wFvwh/nc8ENzq6V4DXALQ1
6hjcJgx5BZJuaORfUJZzF3wJ4StiCVcnJUYRHG93yiZygQmMr7gm1M4wMeLg
hFDLye87pWiM54aB+j1/szPlILyFVAsD2CP8Sh2HsJXOAUpT5PCYnYVIF0Sp
7TaO8BEesKa74XtahjsQZWEft52TFx65MGjHbPtpcoRnMsNANTJLffJwxSXB
mby1VXQlLb1AujLqB+dfCJEbkNMIyihHGwwRUvXRKcY4y43k2r0515QbXzt8
1MjZBU7i3BjogdiuprpdHxY932+hc9f7uboRAOaSiwpE5NTCnqfm8UAwVyVx
8alw4yYx7Vops59VzxTgSk5XHsdcuSYIiITasJKmJDTQUXvFsqQwWXB66VDI
N+4k6bMkJLp6wCRKQGctedR6tHjq/9p+eEhyzLWvgNSPILYXm+X6o9E0n2KB
OI1hRixFRNojugmI23nwgOO+5S7NHUNOTdBwRcwPuZhhwXsAJiNn3mXwCAL4
YiNfDEqnljIgl+aN83ITiq/E2ul9+THQQkeneFmJ2hSJUw+jLOv1U5XKBhiG
gCPzbbXZbP98FJrkyqRmyo63bVEjv4O4CSOIPy/tMGGYz37vPt4akhZQyDJm
hHJYFN6+PRLfZ1uruLKoenYNJvv8aVDXM73JHgGLE/ouUdpsz5fKDTGooueN
n4/uZ5PRd8sh6KaHCa8amJg/qchHF/zgag6a6+rFFGaEinIzGU2z0PDrbWAu
jx+ipxX5S/+CAJiuZkHJd65xW4Zde89lc2cKHtOF6OVRL2CQS2ftXT0KV0mV
iMgJzoYVusILShzbOgJubCn6i0zJ5qoAnrf7ZT34fafovMRD94BK1VRHYwdR
fy5N533PPZXpUK5TNXbd8girStt8tGClLC7f1CprNQtm5YqkrN4h4Ex6fN1M
dvbhVn+JMLMgn9gt31loQxu8l2j1XvTG5M3tyGXuC3uU33l3s70zeHO8lsKy
6nGgMBDagXa6xpPtx9FYxbmyG5cdPgu9YdCWk9sSbGs9Kzroi/2oZavgxbNT
R10j5ltYmcrDGj/yf4QBYbUkBFzAgsX6DduqNXnRxNFiuMOPeDPbAfYaz1TP
SFwZ9uljBBMc8cnminxKTrd+3YKNCQQ2qUWF9a9b7rZBzCH7EHzH9cxlASID
Cx+Db7KrQ8aQ4p8zgjCuWLwdCVBYwdwXrctEshZiGNOOWZdCO7pgjGac1p+G
Ec1/LUynfk0icncQogShplRscyvZ0JTfw1GmAXtsPC4oBwijphpmj5JswdMU
KXK/AKMf8teHiheuKb6hEtroJpQhBLuG38UXXY7Uc8l5KSNiZ9n2hodceXCe
HLx29fXU6QcAsNjUT6yNfpleqzTfAvM47yXe8SHsUcQm/fpVAhxCdh7I+VB1
edyfPrDwiyl6dV7+g6PObOF4kM3h3V0eIB8O0BG931NvnhiY5+zzdIEos1fn
VFLzNip1UJkfQ4lNokGXv6M1UVbKHyOtTmULUTThyAzdNQid+pDyEuWtbzaW
E3Pg5O8e47d5mXy4PzVfBmaaDkW1zTBg08YiohZzg8J1iisesfWT4AO3DOOn
zg3bPrfKaZ0lS0pYVxBGa6tfi5Hfh7S5baIr7CvFQXjRvufpRi9qrv0yyVie
ZrNhxhGLe7EJsq0Y8zpKwen1399MG3Gvo5OL0+BtnUz5+WGdXkYBLB9fSy5p
jQESlKMj0XZy617VUUzSQ+Ar2wdrGEj00Cg+BBGJEWeJeFrFi/kRzC97DnyW
vWZkuvD2NNY539xMXBQHuTyinZYGZ4YlptSEW48jqlvDhft7B4KzwDRLOhB0
8x54WZEp3R6NWEP17FEkjBJKY5PRXBI02aGFC5EgbtOmUyBH/t99SL1dlWNu
fcJ470+yujOmW6CdEdGdyG+HqYoa6HR+7GOX4th5YOnUgWTqdgnGMDEWrjLo
sBPZIzqIuB+OphpJj+hTDlVcYDmR44VgDJIT88DuXVdR771lqCdtAoA74xDv
zzkEytIwUG+pUTVpqtrnu38FRnigEqiWcjWy/XolR7PLLQjbdzzyt1r0SDJg
eKsZ19jORV74agYk7LzaBzk6K9UKhYQNVR8XUgiq6XyL+atKITYLNwP2NoxW
CbRmm1f9M0WRK4jrMs0twbFSYiLw4b6BjdnOvtZpiYjXg54/3uHDGlnM9sfC
yzvBvzcxbH6ER6nHDdjRiVSCS38sNIwcF6LEgQLW4gcDPt8R3f06MB90LaJu
0ousCa2ZGeUY/IH3b/r6VXB/VaYAF+QClo14kSBh/f1LzWugK2MNmFzx92cj
67ts39u4SuqGVVooJceU1g09QVk/cHhvpYgTJrCMY8hvxHYFqS2rkQNVX/wR
YX78uSY/IYj7d0z447y+a+oR42tubU+HOVTrQqwThWNuy14xw/fu0BuEBWsD
9ija6r6cHcpp02aVOS0MPx9fhp0z/j7SFZFYks5T1O1nniBI6daJ2PKFw+mQ
fGV5KVUMxfHEQFkyDjN9xc3ufNn2B2PiXmKRbHfCYOMhfuxRNgy9LArzwhhF
KltFi1LeQxJ25hjb2rwHFYp11MiSCZ5jdoMo/XTJjJWIawiwpGq0Y+mn2NJ+
2CnKms007/1fhcrBJN5W8tP0y4BLULvEBaF4gs+UYFAjxjMpBgUrbPSn7BTK
cC2K/p1ZJlPrDPdbkVyQY3MdN+K72+X+5wOW9xuAw3cqZGQuVSOB+g/xoOCL
nOK08yRcFafSFbbTfWjwpQhs3tO2X3sXdFo7ps8sFMUQ+NUoefYNiXynsepU
5aKt4IwnxjCIW4+GCNS6NKSVyVSY+qFqLZtJJV4MnDGE4CgijYVcQumhhI2t
Sj8NUxv7SY7DzUNCHPDt0PoJwlAb2oSwha7v1QEHyLEJbaE1+eslold40m0h
2cHXFPOk/eC0kTAG2Gryr4L9esdIe8YRgc6vxzlgsvuUj8dhOAJnNZTd864l
SYp/sdpyXPnrf1LUAqQuDxNwGng79w0a44hbYiMmonU68kEoEpWxmD66UChz
Skateoapov885kJkyJgZSiyJZkl5avAcSYcNXycIQlGNGah5P0riSLIANFqG
4Knl1UDVzCeN6sw3PYyA4/I1h3ei4SK3ttgPRpaVzMKZKe5d+nE+Tzc8TZfX
vXd6m0Qda8q3R04XAC1wIEtidxzzLBeLoOPptOZXgcFokW9rYciUYVh2DfZy
kLKu5rZM9TEC6i4xWGU9tDSNzl5XlTEHOzKyPenzSydBQYzbyh+/HfQ5aqC1
La8Ta5Pedt7jjenekxzzHCVmJVneVeGwsI/gmTknj4zdb/qi6x88441q1GdU
hoWq2cz/3kR9OFftv4EGEgBkSr6MsRPFx1flOH6UlkkN1mz70zEwb46yb0MC
lCIvnAkCNX7TV1dRyvk+5jkGOHCtf3HAy1fsC7Bhb75nBpEPXhZOFJ+F97ku
m93/q/VeDIzX3pNiQ570M3LZF4ZZSCDa8V5aeDgR2RF5/Zof/ke2/Ob6B52t
n5n0UtKmN95WeWJWMwZKRLcXnT+K679nFKfcBW8/yu3hrOIRnLKM0mdCJs60
JFQzgVVbVVPPYpJAjMb3+xs9KqCF+UtQvIlyqEVhHWYwkMYn/mgzPysaguOi
PusedgZvV2xaAqX8y+xJbiTaFqFs8iujhYgNyZwy4o0/1mSjN4HZccjasHWA
ocaOu4TZ6RYIFbWX1WiHrWMQRiXolKkZnAH2IA9yHHIchJjcst8htybYfpfc
07XSDzw+vyprZnAKThY0KZbzOb37bC6vmE6VAcH++3F/0UPpyWECLOQKvQ7H
bYmOpVRsY42WjL4mHLD4h+pvW9EeW9IYE7kKxWdM7ABlklft40QabcfZkzGS
M7yXfuO7JhZv8hFcnBd5dg6Txc7QJdWbjRksljEs8fRv00nW421fWOqODrv7
oUg9B/3wFuViA9wHjjuI/VGJgkEe5OoyO2DehpKYh+A/Wx6YMaomcs+dhdOy
amjS+Eq2qD8dgPa7Ef2WFL5J9osQrdI0ubllcMdORTO1I9lEvAryV1YUYLcc
PFLwpq55wutHrz3PICdmT3yubO0XzBYjrFHSNegFvenijL6ElCpBo00KN60S
T4c3CoNC0tYk/35ZlQP4XWY3VlQmjz6ljzJMFV2MER+gmf3KaM5He4UdBRE2
LjomOb/uLhCuYTwsaYy3BaoKNLigMHyLxZLmuvbbkQ5+RrV3xGW7hpb4JHqQ
Q+vZ3S/60qhLgHCAlK0IpvA03jyWq0ZB6lZx/K/NZKU0kMfroY/jlOx5u6vX
cmfc/bwLF/Ws0zL/+FaK7VUxOpqO9YY7oH7gIU0LOj7kLiwgrTff5g1rHxQB
fCCKlowMgAiV1SNzU6CZbZKOI/W1lFl4FPEqQeo20C4LuNiA6kIROToDVIFP
buq8YOJFW7aeuPV9Xsb+JQzD2IyQnEgBo0vukUbtVSg0fjR2IZ6qS/eTnrCo
W90gdateKXP6Erb/NAX2A8Why1k5ITtHgBbGbQiPwAYxarHj2Qr/bbbSrvxl
lU3PJ+doL6E2iclboUwD5ekGEeBBXdvGeg9KOeEOC8qzQYWr+Uotk+38pDtm
B4wBEwtBfMv5z1vMX/Ahkd49jXFfCFXhx4Kv2kxgpa9OcOIejQUriDAAbkjW
SmIjCXc56ZOC13x3ToNDua/B3ndQwdi/IsNZrOUXmCt4j0wsfAkIJXBbfUl2
jCMcSpa0iliu/u8pSgurdiaq2FqbCEbJo40jXrsd38Sp9dFddLwVtcjoRNe1
7PIET7nIt9idVoy7PzNDCtXH9xTx3642DxyMUV9ODaqlTSvAvb9qUrvZJsY5
CuOZLF8mK+gbUmA2bqHr9uaJNO2ry8MKezEbkYDStsYVn0XMmrV2fJZVZpNm
FSDxaVc2pSkEIxDMHgK9jjuG9k1GYAuIgVIEntUG9RijlUw+XEpHNTMBRkJn
dotRcqFmiDdhKwT5sFHUgKgdSfGbEdtyyZ1VhHA9NSl58U1ZDcioMiQIH0Kz
Isk92C8I8Ju88Le2vrIcDjScw2aYNVeUrhmK0Zdpgc0OpimaPvXgK65jA/9m
KoVFChHIiJkHqW6kcHmYaHTNV2QiokCeL+EQCo3iXRzbk4quKGsCEttowpNQ
NQj/Kn3oDwX5fayidWmXto/r7kp9xN+XV9qFzfy9f8bbXYvkvf9DTkYyeUnm
I06odI6G2p/XrrGtidoO4WztEawLLDLmuYPj+o3klU6JFiQVs7qgy8jK+9qo
stwbNHn91FKwfWK7A5y6MMme2IMFa4yyOY3HwEtnKJ8zl/IBLzO9EVh7qFEr
DqkdFXKtn7wO6fi6v6ESQ1LEUiK0zbTFDWen1qxnBurFwhHpxOBgKVyXD6/X
/DTaUQ56fE4PzNluE2C5PgLJLPQhuSo39/XB3evHS4TcU5HAda2dNx7S7mhE
Oo3ubmiUNmbM97cxuLRRtF75jM3wujUKjS4cnFjUtJk6OQguqtDqGd9u59Y0
X0+LnaP3p6wJxbIzBOB+vn0pU3lQY8wk1LTY5Gda64lKgdDTAvctfIJN8/xK
R6L9guR+oWve8vFsTqCDm+ahzxQZpkqudQmKq2P6/Nt9FVkWMrb+gGokB9PX
X9EdHiB9hUhY27zpWVb4sggo/QdkoUVrQK3CMvoTBFpfRDTin2Q3Xl7dw95D
xdHKKGnvHQCB3+Bzgejg4vL5fCUE/C/jVRQwuE8RhhkY4u3fgJlZWVUScscZ
eYtQhphh2yNAwuW3W3M0nROwcFse3Ws7VYPfrx90IP7v55iXUTWqv3wf05Ny
6B4INyJEjB33t7OOE1gE1BBL+kv8cl1JfSp7JmsL+0MgaGqzf3Pf2UtIsWL/
PvgsHndGD3auhLlCtVhtGsMPgdut2Ub9EwB3+rgz+AzBFfLrfWBvkZzkBS9Y
6PAK+9FeBIY29jd0m9KBKEQcKRp306xmtrziW23lcKFoeMsGkeyaqUBBdBQI
Q0pw1SKgzH2YuV1OhRnG2qSuNmlqSuf5Z7r0HAc0MmotzDezHciX7OVv2MKF
HO8eVf+YAQiBNyYGsT4oyynq/zZtvsYC41oVw40gtsZHUWpysBwDo9WA0MhC
uscDrU0gyhwOcn9qVhIEr+S7OQCOHjyroZzIlcdjVA+Sc0/B9oJiVziW936E
KP1qVGUpOC5qPgPNwQXmkkqt/QI0+vTapnGgJ1ViBGt4WlOTciAPNf0GrYMW
JHFxZMv4a/l2Ir10+MVmQDrVRaBB8Gi3MzNKSD2BtK++gD7gSAvA+ipZ0J2m
GLTop5wgL0cMMfNgT5pFlNwc4tgRq1GcQPyL6TMX44QdNAYRRS41q2RC9id0
sGg80ax2+/Ezp1j5PNHBIcCxfXlid22nNLMb9BDei9gDE27TMwl8C2V6idgP
eApS3iZriCACvPcc9DhtKsbKnbqf4CEGj3ig6AzzrN9cNVzSePYcrSzib2bc
K3bQcbTukgyBgQ1gRBO7I88XDucE5yOEJke30H99bG8X6fLseCQKBlESuQA3
ZW4H5szxtwS2tyMuLff65c3JwKm4mj29tWbHDrq1maojzMc61cQMOxYvohhZ
LEF4zyBu/zNrLmsW9GLr2ggyUjw+MbSb4ZvZ1Us0jQoXQLvvTqIWWrQQJEQI
rbfYWwag7bRp5OWC1OSFoENOLSgb4yN3JsCR/0WTBELTGLED9TsdmWdQOUX5
wmuTmx5HhidjJiy/Mj48QsmOquSOzXWKKSvfgIR352V6cTB3uYIkw8IqY71k
uLmB6FzYXef7hLDqtd4GhfXnRjfw29kU9gHnqgiuCpm/Mgcw+5TGJNSg4I7m
e1YXzsX/rnkfqe2yAl+ic+pmY+0NnwaqYVXU1mTXJTZ1MitdQJBqOTiDXcXr
iQqZ8smvYPvxCF8vvn711UlZlF0ytLJl9ErT69MyURoxxBhmvsVcViAATv9v
B9bFZ4K459nRsvwd8v1o4eGeZ/bZ2ZZvhPR0ia2bSbdCxNwLpS96jxWMGR/X
JgFwNyDZtwUhomKgqdbvwGIOEz7Dpdg8Q3Iuxquc/WHeuOm63ssNn4bnUmpL
R5XT5ct3ew10U1gKgEX8Uoh9iSzSreCY/SdaeAm4Jli6BJNDhsNb1XTjEznb
XMe811MHOpVywVCdQXZTNBiOfX0XSfs1aN3LPt/K2LteRsXFlrwECwWbg/hW
BEk+BGBx+gQiXoyjzM+DzsdAR8V+SBRav6ABd213ajPNi3jf+es0zwBpCz01
66y0bI0gOb4/lIWZbpG95sUfHkwszv8iUyyLIVAE9ci1+N6AbfyQpgj2h0GL
3MPKQ7gZMEXHOutc7syjPZzYjqmOkZsdHTuzP+tplbhCoWz70Po1ckIyw2Jq
g3hF8MFlgl/5GcuilgvdJ8jHWZqedU+3EWamoipOoK8BE2e2RH6fbI8uplrM
gXsrWbciLDVMxIbruuTLCKIR2yqxRW+xGmG34WXXKbb8c/JERrzoEgYB1Tvo
FJpw2UeYg2lwH+vRFsuQchRiBZ7qifbAaIYIAA0YVAgZemAFerXAft7OrdZN
T5PwqKbm3CehEpEZwHiaTSr5OxWxhsobS5McndlT5DP3fGwZV6XQ4BJ4fWbI
fhQ1JTWP0avqKAPrnbNPV31AEeVV1O2yxJQ//T/En/CttjlxodLI+mjjtlC5
E5Eohf5OmZHzRiEjksHVfIv0ieka0u/xzpMUh0xHgGOuOnZvLTHHLF2xj2qs
+1Ca/5eLKOf1rlU5BACl1PwBP6PFYCfk4Sozj1qiG+xIWI3Harhotk2yTt0s
oDBJVHMdzEnT0wXbpVedYl3zpT2ICVtI3jkpjQcYEJCLh2f2728y9OjC8vQ0
0VhYpOGzengYPl9MBE2ggu/BK5ET76G/0IDY77SHfy53MKhpJw+tETeGsWVz
geDjVOua7yf6CpJYJXVxI4Q1QJrcoRisEcldryaVsaAgm7fRH3VglJ320c+j
lKKgkNumNh9odFQsouugTOsWxLPdKxIw7c9uIwOoMmWBwiCfa0e0igRwgLYv
WjtpvZgmpvdU9iWEC0DCFegfuNL3vWgG0iRc5oceSlMfs/yNw/+SUsqsGDL4
xVWUvLiHtecPKvMgyo4uuQludJz1J5cyh1Pyo6abiL1zOVPqR+YcOqonASu5
gDAF5QxDp7sbZadENSBFLfiSDsjtKsN19+ieda4MPy+gpKO01AHjMk5rAJri
VojlIOXZRhVcn0aKNJFkM/l7kDl4luRBMB7yngamSIptK/MGVL9Ga3OwafFl
luXWIoBHCJEBtp5fX7jbPWffdxTwr9YPtJ7kU++upnuOjlhIsWwA0V5QHBEo
EK1xPtpJ6deox3KrwEWhN1K9Bg5UfPogOHx2/e82YKtX0484yDAXONoullVa
Rur9JcIJ9rd2yrWkTs1VNirla2nquO3loqBF42CsqavlNE2Qp2tLqS1m3OJ1
6qislIihATkXEBvURYkBrI7vnPvxAcjQ8pwtEqp1kcl59bMdvnnM/e8qlHpG
HS/4TgJTGjTvqgGDyg7lvab24+faoQcCU+A5S2JqkRWVtaqCfIi0iptI8vQI
NpK8ghpwEGeVLySPa513YUgvqxfU80+ZGGPbF50i1XqTs7aaPoiCDdnUxULF
wEbd/MKm+aRUrhvZAXs/vzzQYDbiU5NXsl+wf4RwMZ4Amzjsyr9xfItL8IoB
lsKHSv4/OCgL9M4vQVgl6NKGKpB3nhA73QdPNnmADRp/S+gG9FuCMAzgDtkW
wdIkcpAxecaehBLt1+UDjkJcK9TcnBfDKvvGjOoW+wjyF+03AgQ9qIw8nDIc
L6vA4inkNqyzsnSfyuwXP4igwJ31xLcQpQfGLoPEj3i7Pf7zWVYV5wC4mDgn
bHWYaoolJE0I5MjIYZClc7Ys0/IH7N8jCdl29iRZB32wTu7ZGrkIz6CwNCHr
uNWMC3mYgod60fQzjVth9gFKautotsXvDR3rHoPyXmNQ2N/i0kbzk33ZWNiR
zExnKVJI2z5DVwp/3c0wJ5SLpIZcSB1FFAWQhHSOHgib6rZhI4k9TQiYyORz
oa6kimBBzv5iT95aWr2g0uVDubYqxhxHDG6Iy1GPjzPGgmK7pZgkmSZLntdn
raW3ezHOFqV7Nj/A0WYoSTO9ZIxtxcg9NZmrOllJJ3nPZKXNzndgCIZSuIZE
KUlucNWI5GykR4u8PtuRlDbU63RVynCdrm1oCUE5eeAoQh0tAOQnP2a7QbJQ
w6nR3uxaY9NT2nF3dOW2+p7lk7lpnJ+3iyU5zQwcwyxH0r1vTPLLNalf7jX0
H1iBpx1rCD6kNnfux+UNYwb+RbF3rJH5To/5LbFYeojBA5OWMUlnUKsgIVWo
Nqcdn/08qZ8FDTdZSlK4q31EWGSTJzBmcJhcT6BX1rMROYY34593irWLibAy
fDeWz5vinMBwmlqmpE20CD7jxJmY9hXM2q8HJhN5RO2ZvXYFBHY1PZxujeoX
VHLt+eKbziMnU0G7fkSnFLTvSDFQMJMBV+/oy3O0jpCf06fSZ18NkNAu6Qee
DP4gu+Ba7t7Fn2pymvoOP/NBB0EI4FP9gXO8SHKaVBGst6hUjXu8nBuJA1pW
pX3Ux3lkAH1n9wQDg4vrOvyvxZQuRUCSZ5/ERhY0KYhxTaCd2eGxG57h8kxY
/12gJngHnb0/zvWzOSA5Ay1Q9Wz8m6t9Ryk23+JQ/BCm1c9iZyr/+kdrLO0N
0PCl/l2c5OxRGdkfMnBtW4uPQFi9ujmN8e8pVjVjxjlsGPdU81MCEeaxuYik
+zPfNB6Nu8rAErsrvU3xkCgxkJUg1Xdfe6Mx2UEbgWr9eCm3PlfrzpPMoFns
a7Rof12A+0P3AA+cLyen/CDIKmSRW7+8Y4xCFuG2BZk5uMMYPeCW4Aq+Fzq1
KzXJQ2rq/jJzEdubWNMQ7Jm3WAKNxJO1Qx/0ha1tLlNjZ361KD3/tYuspUrv
o/QK3IC2nibme1fX2SiGQTRld85YrTJADGicvudDWdiAqM6Y7FQaSu/Ba5NJ
pA1odAhFfFBwDa/O0kG65I7pqjaNjEub0caCC6XQUf9flGIRtoa1nYOSEKA0
r2YjDw+7M0Cgfc95Ngrxf7Ow+wTngkwL5dAfLKcEU6ecpV9OtUXzfvRLmyWp
S7xVA1U+0qenrs6Y7exIU4mDVHFYIUTwHOwC4vzqLZDE/tbjbUQXZR1cim6h
xLm3IPih1Og3vty0JWy1oxPJ6LpAlnrFgMed1ugf7BTexCDpSMyxTuBGZB2Z
vCnIkwuahmlV2QNtiisjOaRnVPNeAP358zfaF5QZphSgeO0aAfrtY5D37wqC
NcIWxwuPwNOAs/oroGrNz9/GKDnUMTcqilUmqwfkpShuDMqyqb9VmzacfnkY
75Ie6ZXFYQovzMo+7l5DjMHCsKstRdyAA7w+1eMVFku6wLiI16ROer78zegE
D9QXHyBSbO289NbHkOxd/ya6n3zBzxDFJKm9SaZoTv75xxswv8D+BFnMusLn
SVNPka3uLPICG3NXYdUQ4UopYtt/+XD9HGYx1x4XMqOtlCHNwj9C3LPI9Frw
Yptk/BNPrNx91SuqcoJubWW6sGZdpfDsifi7FH6xuaHOJ40MclawwOWgiM4m
ezLs+B2j9Q7CXNib3PUIpMedYhLJFoTvdEU/JULTvZfpayUnqmKBKFYGvVur
hf2E/h8rVnJs2yaCTpXng7HRcCiE/UV+Xel34BhjYvf6dAI4jFfVvdV03Bio
Y87RFjEs/bl8d9nGYnY5BrKPl4RvMFG5Q5sdv/6RydhzIiDMKrOSug+3rQC9
kkvg466j1jD0+xtrA2dq8tDUQKnvWOa5TzwcxGVxN9AC1IX6oZN/T3ICd9ie
bvOsueuQA/pZnyWAuS4nasgTjPMaAaY7mcYd4FtM6YdfICHQI9y0y0tSzufX
bIEF5hHaSSpx7bdSFqjYhtPrquiJDNdYvLIikBZWBspcPK0L0rtBH1tJtf+c
teTW06FyfaeIhaIZ/4hcaedXAu+Cc7QM93Q6mrPbTFfpmMwEhHLBSWCkZE9I
QXCp1dFjF74cv0Q6IDYQnPht4LPb01oYcNvtwTxltwA+2LDhklNuZRokVopA
B2YhedwH5u0p0n8NReTqDgldMMP+h5Q3BK3qBZPBbdShCYgoUj3FzJ/yH5iC
8V9ls70E1GrxIdZ2cz0A4cI9KsBKl4ixd8ADvTBlORu4nLJQjZdaiLmmg2IJ
w6G7U/wg6K48xvvjxq3pzhz5D22SIrX29RJ6t0KGMF+ablxPpEn9oPWL6B6X
nm9LyJ9NCu0cxKRfJEFUIYhMNgT+bqslVumyq/Rg+zXGo3tzTHc+EMtIzQfB
Cjne6erVMhwVpPoOKTU+XAKbFYIV9gDeaqtTyhdNhicggiKJLZS+HND3UDIZ
i2UuhMMCMLtr+0rwpNfJ+zpi1JynsM+gFFQA/9VmV87DwDe8IXINkLSpRa9X
j4fkMQynn9bAgbdetHEAc1+ob47n2kuvOZTAlG5Trle7XXBprrGgMmjnWFol
TUzzMaCTyohROmcGLzPeC+lEI2QDhJ7Co5IpDJaJ4KuuJUz0NiG8EQ2tIB6e
Q5Hzp8w24XpqfMMIMlSH3XZ1OX7/tDKay5GUIGwSJ/wxo0Bdlx0Anm6qE3i3
srHWByYH8s0QFADSc4y+KMl5FPcmnjHSdAgmCf9Zu1CdLN5If2D8hbnMR8Kb
qXSpdCas9BqGPde4Dke3C4hzosC37b6l+RNXKd3BUwEm1HiM/eMSK5EPPkOH
2qRK9j57kzwwUTA5BrbjmTrWmWNt1gC4sZBvU5FfnawU7qv9QRmnd8A6wG0H
ceJwpIPhStBdaA3H4ZHl8yTOZuALdDFlGXBO4TIHTNNzqQAeaL/Kjbt5ASR9
hhxM3tbcLddXO6s+bsuPZcwV62h6hE+pfs5FJLa70so/cVCxLt5oRmrQDoz1
3gKk/lK5ZeJfTviTmlIILuEKoCkcX0ap6n7fDqrBRtAiMZbO6AxHE/O6rZuq
FXb7wNTAUZqKomrCTBERUlNpvoL9Q8/EMbex3sOONdgS7uZBliSIsOpF7ANo
7Sz6dOUV/Z6+zGOtM28XSiM9e/DbXokg0L8xhMv6lcUL7BKbeDxAXl6/NUpd
jWbQq4zMerzCW4ak3RgmXPrJ/j3PYUL4lckKnnFjkHKjUGmFCzN3gvWEH0Cy
b7MnzIpbSNe9rO/W4pwQxEKb1NXiHZzxH0HrKxson7Byr2WHGavoZ2wAo233
t92iHaXDZyf8VsecYp8o87mYrdGVDNkr0yJ9dEIcVJtOji8aOI6X3SfqgRUM
FSpqnHt1pRM67IiwThDQUYOyo2TK+nTWMApHIf9KaYK21FBaxnkQEHToExqE
LP18evQTBZoyXUE2iR4B71z+HCSomY6y9IbmK6apHJzU5sXPg2Or0PosebEf
wLTB2ZOCt/IaYZOIrp4HUkR169Zd7gYae4AVY8AFu49R3+bMEHyyk0t9X8Oc
N2vRgJdtQt8kE09RCnbkhlYnRfH7BaUaiekWYmbk4b6GoCU8MXSghX8Cb+yr
Oo0c3olbRbZ7vQIv4nmk+RFmxeYywrcPZn/mTSEHfYyG2qkHjQYG2IdxTuiC
21kdM+SA/DQX2Pwt5zNPwADroJXJKqjg1jKPKWSmw6vOiypE1VU4RyJjDqAq
SVWWcDtDsz/L+oaF0O7Ou+4NQprWqSAcQsmFuM8C/G6CF5yfjyXrZqKAkWKM
uCo8TbRotRIt6FWx836lFB08Khplk65tZYOdzZv3yM/1jjCsULGDU17wZQI8
4QtcDHKtQ4WEYOs7+gU1Kc4BYpte42fKnqEYLIiOPXWgDLiNpHBeo5PIMS7B
g/K26FFTPW0B1Bq/0VZfB6+OCO+bcvcKu3nw3cn7ri1RbU3gqm8LVkmKHmR9
059yY7Enz60iyFhqjgTPFx43KNO/fXECPqz02A+Lknqm2UruC1pTWPg3Z8l8
6aTe1riZsnVnkl8LmepooO7sPYt7USflXKDnzf2+jxxdanPmSLqLoOAbnqkB
9HI984d1D++aWoyaCC3bPKMJLyHFwYKLi32bGjjs36wxIjHk1zcZ54JYxsld
A9UmJNvirwNVDtxd/dluqRcxdx4xvy4uWXzgBZouGaBF6k8aybzRQiSt8Oko
M72sd0nOjn9kc31lzpvPnzN3Xy81U6S3CFkqj0mE4T1fidjsAu6bwbmzYMGd
nj3bkhf3+afdCTp2kSTNNhbvHaNTjuN+6knJR4+3YXEPhOfwK5e9w095rJ6j
AFA7IcRI/aZTBiWlQwOavp3iG48yYg878qunVjLQ0amgn//VnI2CMWJ4rJtl
6nZcTyFxlp8ed30wwLkyHWSa/1fbkEOWd4ADN6Tso1AYCMwxjhwk8MW2U9/S
+u26lFGjQmPRMd19XnEt4vLDxEj1Rfnuz1q1nyxpSY11SKGRa/ChJGVa/qV9
fnHEzma5jZUM6S+t4lTw4Uil5iIgZkyvv05yFi7wKY4v2MD8FJ3MbX8ul3Co
cJlLh4voNi549IDs+hcIdrnHkCb5qsy2+9+S8GI65HKqg8zEQnUl1h/jloFq
8NBlUC6JQvsnd97reXBL089odQ0mpAVKcWYlIhDQ+8YF7QezcLh+LsvVKYOT
TQ11d7zwo2XIgL4Se2mSgp6SJgZJQaE1HjxxoOO1QpcJw6hlUC/5dovUqmF2
I+WOHGZWOWf+YBQPsLap8PL3MLqm5RZ1mUWEiYdMeYnrakIOsPl11JRScnmO
Mw8KTPgnrvNhQFK21+slPPWaJ6h6XOxXnp6RRbuPJoih0sVSQjL0oSg2VpHZ
tPJDGvA8HHV595HTW1FgSNKYnxtuVIxNULvWX0qOYyWl5sza1fufIu1bhq2k
O4KTC8j4UfdaeNmNzztnpNlshUSbtwMa+mr/ESxnCWIjr/1VgQ6q7cstt+xb
pXQ8Iuyqa3xuRouUUAHRl8FeHZxoyGW+bHmaTytMTKL0+Fr3QHZsiNd+p4z9
3/nMDt+nQ/C833cTQLdieqy5+obJgqeeQGgDGxLBsHnMt5ksWKbo8jc576c4
0mONu70EHDUL8E8ViPQqxz09VJf9zrFkFqjZsJZU1C5T1BtF+5OjHCcR881M
tBuPNs4MsQjJx7B/D4jbnjZYZ9T9gZjGDyTdv0L8PZXIjt/BWhywPuzstMfh
cyMW4tgErmk4rteRjp/bxodOM7kpRe12/339vNh3guBI4FbxyCxkT4KCOd9r
9QJMuYDTFPU6SKXb0zsPSIgoUELRXlg6XHo1QCnjUnylzHDUsBGNkgbO+3Vk
9f9ovs3Bx1OBDFQU8envCSwAkZdj0TC1c98kQX+BsekCD0+LzouCOxXu9g/5
Fm5e8xN+o60Bsamf9vjBaUk978a4UDBcYTNLDVwH0gcphd9rRyDf77uMHbIc
mB18EyvmAA/BBvkhF90Bh+5KsYZEs7lbCzUYIFFq4WPv5IQxSxya84LNZYrC
3lF5Y0XPNbkE0xdUokx/c3oCHtOdB/vHzDiXTfqklRvhnrTFVSCm63R9smU3
33eDxsYzOfDVGm1T55TXwz+G9zsxJalTbHi+VKJaprKXHoTLBNiI7HDF5Wa2
dZ98EC0MpKzGAFYtdRBVVYJszTQgHMosSq4MZrOmeOHfPqTUTNK2PLFGtBYZ
K99CTJv10P6MlmyB0mI2UjfpIVbZBoUL1nvGjVQzNGTHiGgvdqcuSLvqEhey
qPSO9mCaEcaIJcAHg5SkcxuidX7xkqp+1ekqxjtK+DtLeURMaqC7qze6TreQ
EmrOYSb6MEwMv7VWwKW+DPAJfaVWZs5mqRGnOxKNYxFfeGw+Mav0GRbR0QBl
+rb9/UI53KOHS8v9KBxOYucg/BjliHsC+9FYCKoFBDF5kqNn8iC3XZQ6GhDR
8V0iTZovGZw6CorxymU/LBnahcCr1HzdYwj41j1zTiPdZ7o+XbdCM3Xs3GSI
aDO/GZKqN5TJpEImQPjGCqr8YSejrDVNPnGb1gV9I5LqqBBEw2DvgbCHeqnp
gz9KLctidlwwEH5sfexNjtshoKMB8dEIt7ZLbNdlskJz46yH5Y30K/ZSJ6vT
8+HnaqAZXUw7s/Dsq0psknuv1isuxlGKmgUInpG0XgI3Bm/jDbO7U/YUGsdf
je1fFe8vVPUNdfZcEN6JlB7UX4f16MNNqb44kVrIpYp8WizVNVxuCZ7vDU1R
MHrebVLtDaYZaxeVMUlyNtKW609dbwORrmYIqwnh1ZDhF55JFA1AKmojChzK
/CKxtdegPkG9CECpMG5bdbkAY7FSu0MdjShUzQjF67mDN+HoD2ZpBl+TRfHV
VWPvj7VSeft0G1ZlqR0/PrIYwH4Y//i52OnH93FRD79cnmogtV9zjG/uyd47
vFDgBwEb1inRBplSbWFvXoKrI6qKWbgeXub6YgvtT/pdnZM2tDvthxunFhK3
VBNSLrhLRTWG81V65Wbw603DCC9zI0HN1KMJJQhxR/Eo9dohcfCz7LKlBt3K
ipfKD2IQfgliE7KBw5NK0HCY4jbAn2ep2gyyo6GVRtlyneuDL/oE5cTq6AQv
1cCQ76CXyjOL9hE8xfjsNKYCuYkxDHs7JsiH2k75aHJB7m2682KpFTQyGPSM
9DpON0YPdKeQcLtWGVtG55zmY45/5LZEQTR9U3LtT49G+5ofP/zm9fm6LefG
zf31NxeT3PyI2DyaruSVGt7mV5m4BaQXuS3eXDlLPaVmMmOngXAa3juPvow4
e/9EM2jSzc0rvGRrk+Ibm8L/++26EkQpGxrbgQ8Ot+ABJ01X6rxM/xlSTGCH
LYMbyAscmJ+5lIz58YwQ0fPPci/CebPnsr0auXCS+k78G2GhcG9gyP3Dg0SN
z3yphCEFa7Rq5lvEftr0h/In1JWCmdLA66i67CU4aRdBfxgm5kybm2WHsIk0
kCn19per1KMJ90RNE1oNBKzQFDt2Q3DlZGk/ZThdUuN3gzOwaQhaOjnyzP5j
6VSdl6iU8ZUUNep7mmi/ZSqSFFrJZOUaJD3Fn+7FCCy9wdolaOiGJov8D3m6
H37yR0HdIUkv1G93OLbrYDclbH7yabdTl7dZmXg8yQk3FFWgSH1YYrw+xtyJ
lQMDuAdRe8ozlJGoupEu5mvMoCIQIRoLD4D+rkE2tHZzc+zXO+VubVGL7SHk
HzOb/7wLpSn3T57SF3Cvj8qLubQBPWlsTPmWOYguiUqPDVtjARjIDoICLbQf
8Ka1apWNrexku1f5I6v1pxQzaDsM5cUHGEahBF0NHEEuXjNolQzMk1H5cIzP
5itpcAZbxIULXCeXlyeVKmVLDWSlYurCn9HSrXbx8DT0w9APxotlvGIXp+FJ
M2pXlPudamJgFc1J5WBB9L4N1xIUAcFaSgTZAwDhE4/q/owDMdVSSW71t6dS
jekH5mmb21YZkNhwvOdxesKsoy84LVJn7mq+htZdMO0s9w+Ag1+s+vmOXdJ2
aQOuAkpFKcaRt1Pm5cRlBbPzafliyPT3h67TMb9oz7gf4gHRFKqwbRTd1y0n
j3VqLrVCTL/u197XWbEf+XKrPNIThX/G9/YZT5dFQRT+XFsXkC8XrFbNjlmM
HfdKjTBRQt/rune02r6lytApBvgarZU3vp6fri2r/6hL+sFXHNargwHQLCsP
OPzwUTOylG5b+6zlGjS6/CJAtVBnc7qi2mJiG5Cpm9E0Fz/vExFYErCut0tR
uDba7zX8kA3Euv8eYgeVzttx2adJDwvJh2XVMxZ7a6KbPEUcBwfeUiYdobCL
H88WIxREKdr/VbAQe4dT6zYsCy2qpMh36/m6YapnWiXX8BKXcy8A5bT8dzsU
nwGns+7dsG+UZkGCbNRZLiXuLsE2oDFKRmVjmLOCJmzPYF/c1ZC1a6ik5oT2
3tdVt6qBKxQRtQAq5dqSYV6oK0o+iA2T+ZhbGKzqxdiSc3biAQnhJQpZL4O6
ZcfXX2GuOZJawJzgcZg8D5L/KaPwJUvZYqjfHYuUOHZs57lIW2tGS79xNEKo
0q4YIRFxKJU6+VvKJhzuukWiILIety5IO6EkIwP4/PaDWoG5P+3IYdeiEfYd
8RVKI6nZ+MM0QRGwPT8PLl5lOCa5pwVbzeIJov3wQVX2OeB578sf5D0q6PtR
FeFtl1hwp+aAev7+nnTIV883h3ADMGgRO9J8a/VDmh806ly+Z/uc2Afph1+6
ttiDcoLBllyVKfkwNVnIB3K62us8qm6tB559nE6jyVo8QfLV9Bo9FuhdJhXX
+azSVP8Rq4YBDVnbM9dEED4FCMCXtb00vMm7o0IiuJ8KDoKRY8zaVbAwBmUD
L5KiTyPbLkF9qGlxw0fupGep4Z7ZdOvZ9WtWU8u1lfiLx1yrS3skR1AUwUs2
ld00NepphrYEga57ikuaQx4ZTo9BO4W5womWVU3UdfzckaoC18hu1TUwCM6S
FiTejiIFbJEeEi7yaYEx71I436yvsl5t+NGvCFgqw/K5ozq6SZuZaUQZYhhp
Hlan6AwY2bHvQeP8KazkmoBaWV+3K2GoG4lYAcMh6xje0tJWiRZup/XOs/13
jRpWVmW/gFUHr126D/gD523bizUUEjutL5mcYUsPRmDXT+ApwOOVfgqZK8Cb
E998se2NymU2Law3l+sPdEoTUAoQc7jaOr55Zl4oGXELejojH1fwI2erUJID
r5KwQ+Dji1syqUxB12qxsBeDxI+NNdMjfSwbGT+zKhJDUKArx6ma2h5VhF7K
MD6za7Rx3zJMLd2gGaJdUHJEWA5AkMkXH/LdR/cciBQD9JyAyfsSmrTRy8+d
RE/wx3sK6rTrr8kiUsQwq9wQ3Sd1kAGzxGO4AbC4iWRysQKYtYZN6s2LqgUE
kgMWGz8WaMhtjHio2EMYumuwOGMvRJDZTMRw7OmxK46pdjlx3f4IYKWslqbz
msCA5V2o6D2fIPtyNSbS8zvHxPyXo7ZS9volAwKBFI2AfaaZb14ZG0HTsEcM
0214TmJio8CUD/3vdfFXveQyI2TObHCUjW4iZDM3pjkioAMEpK0UleHM7d6r
kZo9jSewGe+y5sNwx/MwC35j6euO4NmW1Z89eI0VSr4Dgbn379T+C6HezTMC
pRqT6OiKew3ysBslS8g5BHxRSnbGg+U0YYX2JdUSNhFtASqB+WwIXw8xIP8N
+Q2r1PhZPCSNCcLz45ahgODjITG3rxbEUhbsk1gFndvrvNWtOGlZjOglq7/0
wXGMYgLTkne96RgIx+tnAKuYwwKOBdND2VvJ0WeyCmvLQ342YaSCkL2euZrC
oEu/AbtQzS3MMfNMjucrG2JPlMyQLVRgvNvgH0U8WkZwWVlPf6MZjzmRPkiU
euabyR5J9DK68NTtXlUc5OtSNGLqZj0ojqfLnoOkmpr/MZJ+zp54n5Fx23MP
0VLQ0MS/TkuqADJEJfoSGGStXiiQICpv4PWd2nwGa+eLkOv2ylIEfZ+1l5e7
Er6RCLxFHf8FENOV68bikrx2ParD9foR+02hEv52f5NIPjCmgJDheWEgHLoC
VtcMNgtyNGKeWneVTgydQlCpf/t7QbIlkH7wODqymHObApBgQokWahwtko5l
aCU7xBzgD1Hp9Fx9mhDmxLCdOAVt/YDxnGQ17ibqtAkxkXr8JY43LOgeYkO1
79MGuxJJoWYSCHTzaV7A5/lQXUEY5GOLO0/90EyxhuT7qw0FTdfXuZeR5MsM
Le//pg2gbbb6a2CVJ9mE7pmODwSG+9o2feHxuebTU8575GwEhkbI3vL2YOa5
y54s665IgHawfJf0Pj5JMPJYEN23U5SiuiojsOPtm9jTUxBZp+2y8/T1R2BI
1pa01j98noczRjRkV9p06OkTfnTBL3yyk/HFETxSz14IURr9TBk6UVIOiZXI
VjulIuFM+ZNGe5Ik0CD7hJCTjaQBhbwSMqKdO8BU/bMbgzlS1pbb0ZAnSOmR
cFMR7JbV3r4ZtbnutTBOixkZZoazF1oZgU9fW7yssjAxEC+NBSDm/RbtTPCS
pS7bebbQzpRBCJTIlJ2bF2IhwJltlgiI1PqcFQ94IpwzLJ93e5/0rNU7byXY
RJJthiW765xOMn6E57EABo8S3hcU/Klu7Ujr18qUiHVVUPRWicPUlybn2Y6o
rxMSRg+/s8wVf37Etoffw52VDZHwIX0t7GpxreFpd32+jbdE57qR393AChsX
JtnK95GCm9kRMXMriPV5+Fpx8RsTy19Dk3SIytG4p3yndqYzSElbopS1DniL
dbdBQNJG68GFOHtbHFhFgAFlciwjyvOIvpfN0a4jgWSHAjclr6wMzWBv3WIP
LFzame0ZQjSmqaCYbMeHy5hl63OvlUDeQBxACXh1pLe02vZ+8eeqo7LORwXq
i9OhPdhmWF5RikT2V6BnRVMM0Y5FZKiwT5fOoR8WmCf8/tx7SbexmWoQIyeR
Y7nqnCI2v6WowN2usuHCluaSIR1r7YiTz2+LUUuyTG4sa9tUfXckz5r77n82
7ZjFwAm/omJgif24Fvc4BEpnnPK2L/CpUWpU5F1RF6ktmsyNXtu5nnuUJg86
U5wsNnyvjrGVKrV8WxU5Ly0axbdhgRDhRE0kiGv0p2tCCOyfJUW/ls7zPgDw
5qYTqbyu/3JOQ3QaO88KAPkEcjUsRYBPSfYyY/Cy+HDMqophIURy1dR7w67A
3qyKv7CMrrXWbC91BRs1xDI7KNiaa93D1LyRVnJRj7b01IGo8JDDJpuA/rKv
i+Sp93Fr8jA8ZtwD7dDSNH5qw+5JAZ7IxJKW778kDDkKs6CNiREInHmJguts
/7MCzaBbGSQJ9+vG3VuZ9ZlOmTnfZf6TRQ7ry4HN9S60bpmtpuJdJrlqkrgi
ZnpCM673OLLDXXi6HSjpVUrS+5xxkrapP2qF6F+xHmKu4GWqwDafCIO8e73K
mNC9La75aW9Idckxg8Tyb2gQqaXk5r8vgNPT9lRedv2knkdiVxsSxVyTOEr4
GgjkKQ+rxKUDsycg2lHA+anrRaQL8djf4q5G0WmlZTpejkzLeEWZHHuN7MS1
oE2DYpnyYPJNylVQ6WJOEUzr3E0HL3uuBBbnUKOjZaGBD1hel1/+SQIjmwzz
ZLFF6KHpn0hegDLKsazWZLiJ/2Dj05HU5zRcQn4i4f2r8zzmpB3f+V3dfazr
cdI7OwY3BUU71m/GGkiVmHBPpblVMDWvY3EciqcMuBWpBf8wzzGyurD3+bzq
yOBoG/TBIB7uJTY8wSiT6wHqIF2RoHlJPr9nLuVFZ3lVCnU3Plx8lNk5akcg
+TgrO8PvgXIr72wYvn2aEVIUt7wct+0ik59hndPbvWmgjMoNpphKi7nUwubz
8uMZn5ajs/eM8fGfRg6Ua2hewKauHj/AL3O5z8K4duToZqw1RUN62QI0rMOi
fFLpyDCXtV7bWazdTfES2/pSPPTEfycmev8FBDAQotpw1846txf5ypzgMqsK
UMsyDHC1dAnBI8Pf6RzAWu2DXYPeOkYUY/vx4ZZOpsVfX7cJuN1zCaqWHJbG
s8PXIBn8rogq2Whdw57ULr9/UN9ATnd8xtDOqpJPR9GvKa6sjgkq2U3CEayZ
40uA8kRhlN8NHQAJyTqYPUGUAR8wVTgTdXLhQlPUV+ZNmbaHo6q7mpxyZwiu
LYO8RA9gwvBwK9ScBeMvvMUC2V6XwtGfqo5Ta4vXTp42Pj/Xk34Qvv6x3yAN
5rRwcB0u5Unr81/wccYajempTBA8Zmij5mSCXZbTg/mZvapc9vjfHB93Nruq
SX92NzbdFkimSqcl7ULiTdhWQbp6kc7vc7nbeq8KzDtMemRN19XDUfA/z9tZ
giZsh891i0Mb+SBO4soR8gC5WywTI+ck/2+wBgEVoNXjUtSlzhuTiDFBAUfl
/LqXYfqEsgSAXJmG0c2sHIGKTJ032BPYdATeq4mg2qoYAP2xpsdcRCDURDB9
HJ+i/CQQhbHE80KRhMElDiNRaYG4UfYSaAz7hmnUHaZ70xdxI8e2KddRfYiI
2YsrPSU+yCLWKxBDxOP5ZLuxydXUt3bSvSy76uoFpBs2RNhq5PKnJ/bzD0NA
3RkWyvMvtA9TqMWv5MhpK/sd/yyhRy92pzyZ1/JsjDnNJVVt5UGF45PpD+5O
r/CHtdVzjlacmFaeMTfclZadol2DA9D2V57F9VYlVWnNpa4u5f6lMu5v6WHB
78HGrp0JGjyg7Nz+rs/MEt5+B1L2xszztGAnT03Ts53ohi1NbQrLhXrEWNnM
igCktvRJricEpFlFmlLk7nVfIehYsXV9VDuZ4lZDpyXsGnQeucydvGHgIhCJ
SWFNbzK1+d94kbVPIADk2rC/wjdSlsjuykyf799UwiE6F9FbG109U4Hg4gTK
B1Kh6EDiLrASucPiZRyYZqWGzUN+wUD1ZGIBMWnor1YVY9sis0JiKK8woyqy
A/rqnKhCoZpNJX1BCZej2qT6AIeGx1ohx983LGfJpzc4Z5T+eVYkQuwsriQ+
8jLnqSc+th4SDQcxB3wI8JD5lgqy2xTU9BU4S4smjhzsaWfJZV4StfhjugTW
bPXDl8d+R5fQL6qjGbdWFz2hGF9oaAGbqonpi0zI1G4J+Tr4bFRxmk5adzqc
OaDSsCxu7IjBM8YOS2R1C5CWdasJnvK9cVlY7KEnUqW6oaG2n+pdl0bRCjwk
olhm2LNwCliob1J+L4wUW3CoMnGANscPh9T+QWoRFFoO00Vb+W3CSbWBpejq
TdwF61t7D2bNVEteRinqCntIM7MP5mIkQRGSbKnLb+xfUZ8Q8eU3brJL3CBx
e8zk+Zd/UR+ODKftJLytCsLgz7pzYSn8n0YUjmxfWBPmI7kBEYylR03E+EpW
D1y0Z65H4uHXbE7PEN9ymV7/dHrBGctK8QTFpnX2CLNwfUvv4KfSmHVu7sDn
nQTch5yDOED52zrmlx8xnsKnjBpJjW6Dv+eguAnb7VRuUKXd3e7MXr4brG5W
KAlUawFU62JNVGN9dsl6IxWar8AKYQhdCEMZUUtHg1S6hULj3bnJgamMvldf
PM0u9jmT5r+9VK3Pkz5TYgEnv5KTuiaVzCi9wdoYpL5l5JWBzpH2U1dx55/y
2pBOjt6sZLWoDdIou6mOk7sQxSZxFvzTPrDVXShU2Jw0tLKgc0qF3XuLRifv
314kv0ZguVVm3++mBdTyZLlsvYSnQImGuD8DCGIQJVG3u/MoY0uhVw0Pgh/N
XKeEC0sYF0jz/9XFLcDaBea0WEOjPFJAXseyFc+pfMhirCz9YCv84OelUU9I
xrJ2dP5YaLZja5yMqn4UOblmOPvvHRM0ZdN6ZP9GdH5mYDozkH9NLpxX+cSA
s3eXAPeciulaUVebhPR5q+4SOy+XSP8vh8LvDJr66E75E6RLCWXAUy9wjRSw
kaYsG0cZHw0dl+2FyORFTyCaSKAl6JBliI+CjKjWx7E0+h8OfwWOl981PVnn
v1Qsqx7fxk8/cYPcqvwPqco/T2Qo5ot7EYZSEDDxZeeHTIWPi0QSefKryHd4
vKjlgVDrHJIgnlQV1koSOuUZVK70awlszZ/vfDNuLHstdtArvpDHSvJKac6m
qXDbDDhsU6x0BynjxotrqvUpRH1PXE+2ikrCstPE+QbuddNM2l0A+gOuPa/y
clWD423bkGkS4Q8GO5nJQQP3NLmEWKt6CgA4LWiyS04oM7Cl4a8ewTUrf7I0
90TCVFtrMKNG8XEyMm62fttLrQtJJGOxhiythilkG9x/NxydGmtfrv1HYNVJ
V52MZ0dMnYTH7HRHZ1IZd3ktBGnUMBZ7yS6WbHpwFNM90R/nAJ3h2nRCtpf9
mFUa14mRFrppMY/ff/UitFfR5LC2uTVmRyE1lkJMYFZy6t5Q2crtEHKLPNbV
GD+ZB90H0WLYoDDcqWQ4VdZcGWZlRCUyyYc4wF9wwoSEgNA8Zf3LlcF4Z1CH
rbXKAV6BBIzixlISsgdhtMPs8tcy7E7OsADKnk1Otxof/3d7tFmRsscrAV2y
anUyyHdvHL5jTCXWS5IEStjuuhylDvAZvPKID/9WvBlLMBpCGxSXG/o4smK0
WyormEyaiyCJKawXcONZBqA37yHV99lRbr7xJvZl4jaxcImOl3yBCCI2djR4
RK+4O/HoUMjGuC6OFkKeaK+a+gnJy2LlAkMDeNUR2JpULV94uRo8KufxGA8Y
XYOHRMNokKuu19MjjcCWB19e/HGOxLzqWQXGHEAFXipKh3NkvIxioCuJNQVG
SNlXuJ/KPiJIVEB/SAkrkinxR0GC+dB5wHkEe3XZnMeu3/NQENHZlPpFvann
4i3t+h+vgdqlKBRHsxommTY6tUyVlKANPx60UODoGWFT4QGm223EH6ulOHQX
0U7M+aNprWoxXspHjqaVII3WOoQv3KQ1mlZ8gi+g6bawunVfuOoYEzjMrMrp
s8jgiz/dr4dawlJ1zA8bJKwrDDQwFOdq4TJ3RedLZA/7REKEHmOoIFUmQ5kg
0dvJil3/xchHGjec/4yuOKE8NKbrskwwEZgxOn1l6xpdwR4eay8UcpFFQbl8
wz/rjYcq5DoQ2ct1SQ/KXxetJEJu12YM6hsZiDkyNUYBjzgX4NynRgDDeepa
8Evw2evla3JSI6hICVv8tSeTvMGiOh2ckrnl8wAbaaWdjl6jJv76AEEjVY5e
dgkoJq6pmhpVrGpbp1NYKUfx7+ixlw6P6qHldUiCUz9TaQgoslG5vT6aBodY
BjvPkxwo+wIxTwNXr1YfNAgmPb5vGngEPEbcoHguDXeZcwSWu6PRV91vG/nR
Ks02F/JfYdnV7TtDfgdiVMb/KmDCAwIhHX5kYOf75MPQ9+IPJAGTz3P5n9v5
/M3vVki3s1EtNoBd6YmIjP5w3WDrrFqI+b3O2ajwzfI6KdswoS26ahcoNrRP
3B3oeq1aWveJgmTj8BusSxzKickGGBlKub1NV3+rRhm48orSgNztsAHzyLuv
OhYR9jj0nMZcQSE4QWiCEvTMo3vs+PgtS4DW/p3IbVyngoyJ9cwCdj6Kl+pk
jUbicUqMewyCKXlw8/A8vRC2hMI1CE9ymKwUaavexKmPAGTRqG6NwQXmCXNg
1xn4sO+eX7ObRuLHUw6EUFbjw96jLkyix8N2XAIkBEuzakZbFenmLG1QFaqd
31MXbRxlvue/9BtESaJgALWUifiZMcuvEU8RltwSjZ1VjQw98Ig/7g2bL7Bs
tF1s+8UgloH6Ve0tC+wYTnWpXhujWhY7/RK/8jFGGjez01mg6zRWBCmprfWT
Ati7IM5dUj6C0NUgBjqnJQ4UMbNmj8wCWjcxA7BmFcbPxh7E66Nw4BMONBk1
vXNONXBVk0aY8dMjrRuvMQh0J3lil2YgMZhFPTWLKDTKHQyGT11hgMhOOl80
+8gwyOiWYzPvREoJBpMrAMFPDU4KbRAwEuHlreCMBZkKRaLI27g23UG0GJly
c5oO87aMtt293+DKNgvFxcvu5nWm/gGz4jt9Bo1m3cTl6GUORuM1o94BL/lI
Atu6ZdZI7227ABhiCTThGV3L0NOxJEB7F+EwIZDmjD7V/IQzWlPRHUv3QIdQ
3tPO7cEp2n0vmIWfEQfFwE494vxGfJX6RkAx/DSS77If5lOxTBuSo5cQU/7s
nmPwgyS8vE8A+l8hWQ91P5J0h9tMdFy/ftvs6uc/cs/c4Bt1YrmjSy58jkEr
npt7SWvxAxiPV4whm5lWj43T2txA49jjpahq0q9pyo4Zna0pxe+TC8ls3y02
Ptcxi4yDJ/G0dJkqCHVc67cY/oXdOCAf3RGaBsxGeVmHmXX/HAqR2GwNbmD1
PjviWM2yfT5CtKGXwbTwxMIy1IynV5pvTYaXCKg8JRUTORBHQBfzKcMXoJhd
MiDtGRn5MFH0VU5I0jTL/0e1j1K3XUtNIXnQTluZ8zmXlsoGzbtWyfExC2P2
u94jOD28+qXw6Hm7MJFs8bv2s2YHbUVfXywW1Shq3/aDS0+hWaBmuDO6gXC3
cnDEkARpNlD1QFss+ups1x0Pd4pEql1Pvhh7BJiUmec6+NR7TMsn+dIFMIUX
wWwsCuucGYi21FgIfKoiR7GyAnBSxum+48iJ7gsrdEb5NiJZywUXfc3okS0W
CXtd3FGw/C4Y3wI9MLnZZTpV7fwz0ZEV/ozbBki7+kwmmd6PMw3rP+YT7g1n
NAnwmFjh4DfEQz6TBYN9LHEhL11bNqmnZ1SFnFv0qphd2QIU+9UCIL1Y6pcl
3C5nk6aN8yEtC0uly3ds96PC8rF0SJbejcJJItnLXfJfVxeA22WNsRRV9O1H
U2JTjWD3Ch+fmlIovPIEfQ4uHC6VqSoJ1V9zwOUI1S9MXPOCtVdBCsscNlT0
NLtWKBXeoNDorcx+QCNLKHJ9V9S/CrTDVSanvzvFUh+U8H7EKY3NXqkU6icP
pqd+lJyWzN/BCj/4wgFhGIWJ7atx/3ZflnGdMZyLXJClYRiyhQWPVfs9x2Xj
ObsS4r8+mWUdJUz+zRn+DkI6CwwrLUxxy5/z8YGQyNpcN7ZzmRXF/3yGY/nS
GFDH/yE2Eq3S0SsrOluN3MvY7a3NM9M8aronfjH8yoBBgTMreR13eVYnq70G
s5jzle3KFUqVTOtHMuGLzUTXUMwm3oHnc4iQ6F+C5X+tvxb7Vs0/zo9Prt+6
r49A6pVYRGYTDygYHql3LsTgBVMBLjUXSKqv0pPr7ApDIDepIMyIhpDraH2d
fP2OyLo5lEgDT3AbwQwNUn/PEE/J7bj6vXwFGVZRJCzoliHap5EFt6Uk8I+3
exfwtGiQbyaGjU5fYcW3BKquh0VJNZgfByLEd0rrLCyjuvxANhPmaueDEHGU
hIJr/OhqoUxr/8uAB/bSkPrLC7jboMewWOZd0ygn4smDg3CKriG5w/QMFlrP
bfbnEQ1g4jibt615e30vCNUoGY9/UAXjSnYHF+UzSULG2LlY4BrOu5OnWXHi
5oDCIRfEooxNS9JXbANlyg/vZqwnpM0qrgyIqHjKwIXpDQkiiU+VCOBZXSJk
0L9bc8zJoqa4tSuWDAjbwK/8fmXgX8o/+I6XU+La8/BmhtqWh83KWxJmUMYI
MWD8gTZ5bG1bKjHsT0zsFxdZXfNJOK8V/7rndbvPnU7DL3bOTlJWFq2vy2TQ
LjkV5a++nuDejuaY7g6hKujwltF2t7AwAXhvO2Ys6l7mylbsNWDmLN88Fiax
4GNDgL9KIMduJN3Myjf/c0BhZMcg5VneIrGuLj+mgKTmz8mhhtpql4oZMU89
mSZfcn7jMVLU+LC6yIEjpxdYDDWoI37RU+BtFS2nrXWQ3jg7FfnIHGLv+QBi
HC5ktGmQAZPTfB6L6xmdT2c8S/DKPnssWsw9Zvg7toeQpwv3Kwx/cQk+mS60
a5uWCIWt3PdiT+cXLLb3240KKfG+43ErwRqnevy2YEFQWQhf/XBgZuKE1rt7
tFMPv5Ub/4oUHH5CZiQNWabfyupbeZG9ImOPb/T0qOY/2hKIYG8Ey4a8QxWg
RVDijkBFB7/Hs9HNIiIH1YLasfyH/J6ax0ARwPoRt4cHAggfKGrbl9orwUlL
o01K0mCIsxbb6my9lul+dVhbaM1Ic2rEHkUl+xPKZ6To9ira2yZQ3SNjct68
zBZMZ3zIEydm/kdNRsRQAa2wV5pvQoL+MeUnV33VnOL0yt98SDmsVkkKTiF5
ZEv9MYxWawhipMNEUkR4YJ0ibrpiEkcTslQfknxCx56LuZ+HpDk5thes0fGr
oFnyVRyoi1mvOa5B8+zO4JUB0Q1OaLAiiAwLtvo7qZSvVoA1ZWAqCsZpaFbL
DZPDI8wxZ6/23ph8VoHtOoCOpT+gmUQN/4r4bYcjn8NOmtkNayGTusTnzBTk
B8wD9YrJWd0q45RblT6fPkiCGIBAN7SHdGGvAiEJ7p875G2pfYDxurB8Q9/B
MZ2Gl/SNUIInVO+wlzNC0XkqoItBRWH0cV7qE7FJtnIXwQKtwCL/a4aleN1a
aSDk37qazwO/KlwUoJjbWBztfGbN9PgnxGq8BCE6ZcH59vXkcuhqXk9aDPhj
P7pFoFJr1AfJknSMGV9IYCsQ0xWmdv6yQRpSpWi+lf3hF8byeC0asLeMPlMI
3Yp+SBZx2boc6lZdTkRkJvQVeQqueW6VoGj0y8Njelo3naGCqNr7cYVKbsaU
tc0IrHUopIsNkFjBujCvWCSLlpfDxk5tIIRNqNof0AeMVDTHCOzqxUSOqpeu
6dHhCMz/AEp6gXQ8STveEoy/Tcj20T0xgqDv7Bje8VbC7J5tlzSGilQgHRJh
DYQqL0DGZ76ljVXBi//pplFyNwLslU8M9gVKXOiFV8RZplQBozOfxbdnkM5h
XVawCBHwydnuvxBnMpfZLkgLBR9WrZpFdIHkSt1zVTru11aSb00DKsfAc71/
q8JXFTaowgE1UxBRsicm6RHLhvJ5nB/WNCx1l8YTZs29o2hhhoXykXRKP/Vg
tgXd6GUQot6cGacYM/02PTKbtUrcIhH5p3mBFcJ2IxsElN6rI2Ud2GdFFVlI
QTgsLkl3vhP7vwxMnX03D1R1W1HGm4Z7ZjWxuf/l0tTLwGV7fzTqJzAupcSX
8Gk9/VC+Wg1RzSpcP6euoEEtdR7Ithu5yuwN0WH0pMxhGTm1cLSRqxW51kaM
OVpMxMADo6wl8BpcJ7fgTpL7sUSUthJeuZoXYa2/U3+zl75vHh+//nzZ3mJR
YUt5umfEkK+rNfGpQuWbG//bpK/SghpArekh+rcqdf9xUN4fA2daz7wG3xG9
WQwdVlUOfm+lrArFil9IjdG34g9pKSyTbaf+7vXD8HIanpSpqNAWOFZdYVBP
6YE0qOMc8dOi+KJY8MVKu2nPKEeKxtEG3m9jZaJDTNc2w9Rf+Hhog8STt6vz
G+MwOUCILTtoTqLDIoiNXwOJqqv9dx/3ku5ke6Mjh/79HW5EdOszcm676t9n
zx6DJ6VSyrqPQPwZeEiUyqbsTxROi+GdHuC72NieBgrJ7Pi3oOgCIFBM7Wvc
PuVPuv0MKLY/sy5tTccjEXXiY5FAeU+2ZLKR/6W+WkOHpOoru9NxlXgVjJj9
AAs3VOec1o8GmrBawRH4uKx7tUCn18eJNZv/44QOk7KDRhKKmI1MifUVXR8g
2tiUjD2dkZnddxKr19wVVjE/qfgCZyNFDxQvuKNhz9F3gaqNHTAhqukb1WKX
Ap/7rpNpzRtkkdH2qPFO/qHdy7aJaKSUpzmlbTNAORFIQ1tO7h7MNLkwd4+b
Ywq3nW6G23TwYstoHRpOnrP+dzsbfEj+Wgiqasgjy38MbTxDHgYsMeAfHVqP
rBnIjImueCJT9K0zx1gtmzAszvzUtby7F1CU+uad9VPehDa+y1S2qGJg7J4P
x7Rpz6/DXsrikW01EHNbVkE071rU+7UW4yFLz3OQmkM8QHwafrvRhSl7IVJq
cv91oGMuVvjExrEvA0aQ17GIW8wsZ6yBytXRcfxpozd03DFykXcn7L3U4PzE
AvGyl31UUQIbOKATiR/ZW3Jy0zudHmgyhIVJ3goX8FaqbxICUTPLFxzCMFbX
Db6jZTBn1v6xuG/EcfB5Ui8nXLGT9YCCZZSbLKiirWNsuE4SvV+Q0mdVbRUt
+0m9Ud0+28761ITHhMo6wrwcrbyewy5AaKtAbScBuMxkClg/6F9fULSbSWXg
1MgI44RzW1J/6w/HiJOLcArapKrWqyXkXT4OySKQWTVeZDGSUJQGTT1jcy9M
Y+Bbd/AUZvz+TtDCjyKZMKOXAXLxixt4j0ev4q6CLtifjNQwNEcLL6w1VsYe
7fEl+k20U+eDZQhOut5vFwAEbguUGaP/BNKsgR9K9JYf0nQccHdix8iP08WM
l9XhqA9NpPN289iRLx9Jfjnf/SewlIFOD/DVezBgyy4by+tz49sBHHScMn8w
ftEvyi9KvLAYfk2dwz1mTkWFOjrGY1fsfHscE2WmH4glPEFHK0shXtqfZtpB
Dt0VZ4AOyoq/zcOTuPq3pgp72ubQyrIxMTi98Ipu3OdRSIvJU0mCW/sI+bLH
v7EOsQgO5mt0PQir5OXfAC0ncopu3jpL9EwEaCc0wMQAS/EB+CA4X/eRuyVq
1IyLqncXKWiPunRN01vO393lhFKEgOB3Ez+iRAKae7Hr7XFfiMCOPZgm7JfG
m7j9Sc4+L7uJvDNHomX5gLY2B3o3hMydFpEk3rVRJqAUsoOWCo+3xEqYjbpd
VtZnn4zWc2XhtLEaMJ14HI3Z7u9VjMvfBLaxNA2qQ7/11GkCXUPX0WjIBpWx
+fsynZOz7IaFoivTUIMQrAac5yZLZZC9kispe40iW/CA1Q38LWXM1dZ0r6bA
/chqdoxtOGaRyRVR2kmcmgZTe4xKS5/F5WVArEE9CJ3gdGioV7XARpXPzI84
GFsMRkefqDQ1mCx5kYCi70/fst87T2KFq34v/9H4oqfDAt5OU0QK5b8Vg6eo
XXDuPnfTl7GU5ynGawMnn4rFxmpLTL6qGn9bEnfqF1DRqHNLgA4jDIQN4TnT
6UjjO48k06kboTIhMG5LAesZ5VKPd7LZr0zAahJbAL82HzFJvyiAQTlxGgUf
uyWF94IPF8xARnW9gIJhZ+wj6ef29vHSxgI0+vVWlEHmYlM+faeFD6CQFSW6
gIlFh3PGdgaDX/S4CWJElFu8fM89vI4F1e6zivT/gf5alyvftJwYdz4gjrOu
hd+xcairBU235PeK6t+ZRhVKbjiLB35wWg1rq9oUFPoZnjRBAnBLrZlgWqjL
meJcq0fVEB0Tx13etjdnR5dn/PB0t8T5AoBDpUw7QOBjTbFhQS0N507E9m5F
PMDIw9ZgQrDMzkAGMJAA9QTPREPaHgl0EZ2T7MYRCNUxzITZEUw4cWmWpQQo
L7zoGDrCAEfjIMo3U5zKUzxTdQIx2yjbv2XaeZAwcsWL1zc+GgAj4WzJWcQF
983WS6IWg6K52a0Jrq+B7gMBMv8CAMcADYZJb6GJs9jZTNPoXBGcSTS9bQcn
tyGgcNVBLauM31OTrgVXu8ZYCXdDsBYYuTzjyzlb40avxycTOorEPYccBVPA
6zWu8AcKZB+jsCdP+EyTutfKTA8HET2VKC0uZF3OLEjEo4FjpkqyfRo+Ei2h
P0sNe/29oAI41SLzLgh1aAXE+rZGUkacR+A2bdVcVGvwYvTKyAd9SmWsT9vm
3DVRJ88Y9DmB/XD7pIMqN6u9lYxe2MpPZtliqaeIOt0sRPNPQKg6asFvqcP0
4GN7RjgdAOlTjXcwVBRUwFYOE6+TpvvFt7kBhnnLhLBBeWVCdqYkHUhOZjJO
CzoQLWEwaCO6SVuRNQAfEEvMXlp1Sx+/fbX/a1MTDC4K5oXmKwwIDEW2dMwt
T+yD+7jEpsbLB6P8VoGboOmXX5FQe3w2qc9MrFstfZfMPBrj+9X+yk/RsTdL
uX89W17aQoFWeuJQxMev1eD3H28ymMSZJZv4uw6Zz4X7Axb21vDkDY2OPCdW
fdUDBUe9UXfxcs84ry7ROCdIKWRtUxSXzlx9kXS007MgiXPmDkBSFyGmXsRd
VN0b7PyLASKoYjyGPXzZ/D3q8L6UP/T8cRdwSeme0t0CNKvW56kIA4h0qGIG
3uNZTz8jgMZxW4W4OVlnSC2ab/abSQtT7zXL3z+ZtZ2+7qSEYcBFwfKJvw6X
R2EsNkYj6PwK6MRIcDBHdisdJJvZesStDm10Aqaey9GNpdFcgpgCMFfmrMoV
afKG5Y/ju+7J5Bu2gqwHD3gbmsrwHkxPWJOceVgCRHJW8youMFbnY8Hbn3ZC
YBzIUi9oTrq/kqdOFip9gMYgWmyMmW3Tv01CaD9BsNr0eguti5K+dHbd1Bv3
NSxZKhMuX0opwMRvX6oG1hoG8YKKJ16RkVT/eKbfgD4bsP8ObwR3lAi8p6QI
ZUyf+rcSw/kPsHgK7tGg5GRrmqKGQr1/UGTiOnyBdkMe1r4Z8YzPc7FDwqnQ
A6d3Ko2He02dxCY/F+sDJRcWVlYAr7B0ZAnxI4FTNk6lGhPOS9xKQ8ZL4j0T
IB4EUUp+6ajuFYHOPTYRQtE/KNsuolcwgS6HusPtBMq18x21cQOhTb0RKIrk
LA/cKPpSMs1abYxdos8KjQyacXfOdvnkcbLmX2jdKrbYEsTJS2m9tmv4/mWe
ImbfVQT7wZqtQBFBrZAJYVPf4p79TomZMhTf3dw6tPZjkXxum5hOupwLOg6a
d64+H+1ZVw4den+DFVAcw1GKLBCK44Y8Vz8PNV87hv8Ngg0OjmQpnsSZyhcW
61llkaHJqf1q/qsvZpJ2f5b5wvnYjK9WCs63BIEW7hKqOmq/MGQCQdNtee6E
PJUugWBwR7Oft+c9xlDb6nj3KXL0IHfHFoMz8ZzB308seDwoBhKCLbwwncXl
ubDKHPKm4TS2w+wNidnV+5TS8LnK6prnvIVajL/80hqIWVBRBB+tMGUDe3EW
NRp5ko/Pg61ofj4Y+RdcU6O5ZSEvXXrfl5MbaTLOOjKWTYPprSD8OpO7xxH/
ajfjeC0xh+v2Wlf61ZAEF/0J7eLe6d79q+l0429eHevEjcs9RU6TC8P2WWTp
G7UlahunEmhpNQHsLBVXEClYu45SRHNYcRZ2TwrY7ehccDMMZYs2B3QFRGW6
3Hso4YniENFH6gDsMPhEUDyWGrzux0TLvYurJhduKEhiUahKc8fj4OREdSaR
xv+fV8N+uTFRSOzFQUfdZmaxb19fRISqw7GpGBX6N4DtD3cBry0k3dFb8iyi
HPLVoLkP55QnY1BAj4xG+QWNzANfxVblywNTDy4bwZS4umAP3WVnhHiF2grf
bEWQWqiujhknnu80cu19mgSD6nE/VE65NTsAOoNOA/TDvZq0mtYD8HOqZU3w
lBDDDU+aFfZh6ywgvfdANxsKrfn4whlkTGesp8CEHH83SHy+KZCY78VPi1bU
7TW3X9Px46qqnIi559UftgTHF2BvNvIvjY+uxFTELvWI4iLLPGljk65FNsOd
lHg+ZAybLdOjcILwC4ZU0HxwrRLx4eGh/Ka/QqtXOvQTsqHjdawS4QLh9wGZ
522uzighp25+3d/h63oKGh4eLKwbkewO4Lt6BfDWmSN16MtTKglZmdJVwLNM
G+ea5HKVWL7Hih4dl3BSxu8zu6aITeIAw8M5eJnDvEyEHP1ooQnsb40kvwN6
zTfoYZfB4MjPlsaJQF3uN+/iJsUGrznkmSWL/bhS2IMdDNgJlUWbW3v5v/40
9pEhK4mkQRFVBZR23RoHXeYjTCiYr0pM0UVW0h7luEKjMpM4PQJlj6QSn349
hKOoWFd2c9vOA8sT6ccnahQQwURGIw1hiEVkftyKSYDF64IZ9FPwPrC9t+nk
lOscHfWY/EBWgNMmgtoykRMIlLBNsroRxIMBVm3N8LHX2js7F7IqInSoSD5C
HrnuKXEpkNNiXHS9AhWt8BWOkt5ejORwvpHiQs2cphF9f1NhuGxcaYyJ4Dcf
7/4mivF3gLoc1RgivgkkjiQWF6bMafO9PeKCmlBxlzKvdsL+/0C4otOI+2nA
FkBheZKyiVH1mdX6MbRENR8TC+VagGCOCqCMKkWEZ9cZCSnw3fZ39XXPR9Gn
NgSNnNzw+QH6/YMUEirrS708gaXYZ4Zo6UATQxHzdivIVdvSNwNkSip9DGmX
1+2jDxngcLCDZbMyMrlcpf6EmOxbjHghvjdfp4nTx9/XLTboipvYNoQGw2TK
81HyIXvJTzV7F8Fvzdc59h+rouCHdWYLrdsbEna9OFGBKWgVIXQmgggmwtB7
/MUYRNAhymFq1eGyA4HCaRIltYk7BNrPwgk96mIDsJa+QtxyTm2jqSaalA0S
GApvm2Ajhs2bSIpjUrIBDPEpwkiY+JEX3nUDQ03ZexWMo+R/R87YFVUPSox+
ntw1MGFYy0WQNXHLDGKQQt2FGzAkYAZTgR2ubaforzA+SkZUMCfDxlVT/U6B
3Idk6Fvh2e9OT3wYKpK2uzlUoPJlgY0gvjqAlDfc2ibgtwNsC7rSDfhhCVMR
HWKnpNiIMocKZKysvMDHiKgzW8WgTPwg32oknkjehlzQ+5wsoAg/fID2BaoD
LWpbAbtgnNuOWDasUQsoX6TCrfY5fwgi/wEBXFgxXVYuNxr98EaiuNI5UgxW
pzdwgpOOEK/prTZdyfmx81S9OLEGDeTWfkqnA0fNL4gF340vB+k2wEMslGZG
daZ/IUONAlfHIzGdUYyR8yK76nPwnnc0vgyb4jQUxjvWwVN4c+gQD7Q8lLqm
D16W/8jCIX6giYvAUe21T/gHAHKkmHERFtBYIw1Gea+9e8n7zY9FSAEfv8j1
ybcANBGdo6D1FYe8PyNt+C32l/Lbew/VAEqNr9cuexM1o3h7QA2fUH/W5OiS
bMjWesPqPSVKCC1u6EQy9Qh2nYLq1JhhDpo8HZkadOEtpsBE6Rwz1YQKVrMk
FBwLCZRHavgIkQSYhSFfp+xaccJHV/w9zIGrj1JkW0wTFdzazNlPZbeIlC9E
UFg5GyCfAlF7mS7MwWZ5ABIX28hV/EiK0M311vYaL5z5lvGA95DbzPAOxQyv
4UIg8bJUZ62lz4tT+aWoIhOzQK8xf2uRUtYSSyfeJt85DBmhja9L0SJI1hZJ
735hMN9fEcMj32i9cEOGsyHKlIYg5qN/g5oVXvv7/S0o299FTWfR6+86jBXq
OvxlJcpTqG79AvdhWn7zQTfYpm39cHM+r5TXkLUZa0qn1qfH2QIGnMP0IaQi
aa99nUTlrh1EuLf6PgUDrIGZ27WKNaxu7+R01WTBjdmJkiDjJCgLIq0amkF6
JsLAZnUBE1s7Sdzs3rYPyPiB5hpyiS/DzBht3iygmVR7E4N9F4n1I44sU1dX
w31yL/cAklyuXAj5Olh8uXsn8oXTXFdT46dmlfEuFpipY15uMY4FHkjPeT5x
w7cuKunfa2NvMbKkipBR/MX4Dg+jzcltJtSi7bpBEVBuKTrmht/iVJy8O9zt
ZYxpKfCdEWI+gTqokF7XNRfitc96iemMgRRPqVUhakW/puoqGxdn2sRbSEp+
WeUgSaa72A+MGuSz7tsyuFr4mJzgz+bxMx/IrEvdbVluiqetYfXhMwzSJBuU
Xmp64w5xixohW4npjhLlosf2CZxGEuwTA+BhoyiYT1ir6dVq3Uhingr5dFpy
YlmDHZ3Lkpb6f+twKtZTfNG2ujroZiWx0cjx1FDyhhvXjARjhadCHr1D9mKX
A4fwaaCfw3hst3MKQK8V9oo/g4tds+JNca9oST8m94ftyy08J6n+qRPX2Rxl
ruPT1C2JMOUE/Alhy8AbRAVfDlj3NUWtEYNHbT/o6z9C3UpqDM+iU+1NmqHR
LagW/sOSTsJf9LKKYgKgGdABr/mWPoXnn8PFi5UXIyVOAZIOqBJPNCsZ0Zu1
cSybMpqWWSQ/5xY3zkT1yN6RrMirSA1In0apW4476WYTudAA1FtNy0D56j3c
Nz8hoTV0BTaXIkHdwuOHgXmYBiydTkduqNVvK72zBwoI8xapuafLeqQuzx78
waZdB9UA755TRgkk1dpLgFW9BX+jRjzP9oVi52fLKaixGc/bUN03GsNowOCM
J65m03rVZrPTJehzHzzdepbASXn6kz6MNb/4teHtt17N5rdSWhlp941VnQ91
dL2qEO2dvVH+ilXA7kO8fqSZpnmJdXzWHRg/TyrHoHsxF+kQR/mPNiSPEChA
f5R5yKPAyfxUdOsNyKHFd9hu7grcd4msM2IxSZFLxCnARFatD1+oprpZnD5C
rxjDyyC6I03l6NfO5JWqwxCBBUaPNHGE3IhTUJSUKtDmkX7QnJbbFSQH+sb2
dIG/yG1bE7l6KzILE4OA7Rl4d17Lv4osIesF1rMNnKcqe4siGrZwelRin2Vv
Q2CmB676gCWb8OvyosG+U4E/1uuXddvxSERpu0x4A5ti9Pg0K0aXe9Ob5JlT
RnwK+zLn+uAf90GQC0t8LO+Fu07v+/CU5qzwCfoMtUmM7nqkmbi0JxzCGZ/g
Wqn4SIyd19So6tEmzrP3+9kLB7sSuImtCHsMTlvFBmEZGoXNaBfAnbuobcTY
unjLzK0crsExS8I62eHhhjU0DLxJW6fkA++j2qlob212pUFLVmeGvAX/51Bm
lJ5dB5p8QZOQDTzaoGeQknAuDLd+e3g8iftuuuyGg9NSfrRVbtM936SDFK2/
wKvMzEHc6v0O/zch48NQBC/K0AW3Ahab2CUf395OiEpHnxOT8DAM+Z426/n0
GnL1NH8NlxaQG9evJ6mFv7GJ+JfdUMaPUBHPaDLXQooL1VmqkRVpVPyLWdEy
WZHtLAyqC6/0i2DDKKWSIJUNUCgaoT3yMM/269HIy2w5rmIvsBZ3G7fzaSbh
sptxHlr+4B2Rk7Kay/J0NOGKWlLA/trxyJ2Yv9ZA62sM6OeJyJbFwZdN7r7s
C6ZszUJ3Oo2HhFm94FN/4wUhwKUCWQ9p591tJE+jepCB2OttJW2rNCofDtnP
rv1MPuapF2r6F8DYVyeIQe/0HTIWU2VGrMkWeaq7pgkcAvI6b92p/0Db3kUC
Rg0IRX5x9HI6CifBMvf1uR9slAErEpepBM6mVctNvBQ+SGrritTybLOFtelS
CjCbtT+pxICYF5GRcM8+R0fRHDdO6vIvBcyACJVtXB8QdTfgjsu5HMo031dt
nFbNhvy3oaGKVwpWN2OBjss8MPdCW2zdRHko+3MwFg4qrynujDY+eFG+SIot
j3Mdp5xGoNEI2bxSwh+M3cf+yA/BzwFMf/9FyXy59oNOHXbpSc6SAOnWsA6N
oHQHcDSMVfVQnRtRoZYi1TAcJGXosFSiYAFL9guQk1Q4epANQEepZordwGQx
vKc5DV5Oq0G8KlmY8vP6q7f68wLuJhruFiSGPiWPB2c7k2RsG6mfAwQwkURF
5VVkkgwyF7QFQ5lu10qaSsquyH6GX2eZCZX7ZQY3hhToFZSjcNXI3shXP4T0
RTXRY7Rk2l4+HGZjpnaa+g7Gqu3yWOH5NviGisqzT6WmCT7oyyfyx5u2ofIa
lEPbra4YgGMpT99WytAGiaCtOBIyh3Kq8Alx/jLK3IfbE+ioK/u7hT0AGQF0
cEYJXFMRE/CUYDLOfqCHPUWu2NZDbqyW23o9xvs4ic5FCharomfDLK7GozJt
VT/UMtcWV7GJtmqlzdllkOA0ffz71rS0VE/JJGbDQh/VcF0yvS//jjArIZxR
MMkF8NMDqYcg5tpmQTe2ZAM178j3tAkYhAgSvXlx9kkZKWRxMcoEFIa/QckW
nutkX9LpqVQ66Hlg62T7JQy0hkDbQGM55xxMRSOu5VcFFev2mn/isFymSQHb
fa4HT8AvBIbMTh/s7Rec9DSkyAdi+LmKa0M1hkvcbGsrddKRg7vjikPeyYur
egMremm8dwkIhnWPfWZpHy+FAJFwsMWOYw8jfeWZlWhq80HLll3Ow5ZjZjsX
WYLHyAQizdmg8C7lw95LMn4tEehXHIwYioQrLU5E1KRJfDPUkbEq5+iCLbhn
kSNDN143UDs5BOfah0BQsNGidAlNDrYuDMRi0tUqEX07JQYbmtkfkI5gqWWn
Q7ywP7sKxY0Dy+CvLOJlDXTKwyQJZTEE8bGLfdyvGGUu0tsgiQmPJ1CzD1aO
2lgCz157uX5uEX9LBZhiH7kn+D4TgVoTPR8BiZL5sXTu7sYaZmRzXT2V3M47
8onHn+KJnixTnetyx0dfzolkp7xaG+0xfCpd7gB4iT/F5hHqSJL+/FDQ05Za
eajfw+YZGH+6kW8pCpap8cgVNZCwqsOBJdd+FR5fdoJQtxUA+TMQtXT9+CJQ
yHFPdFPE8WeWZaFq8SUJ07BMThUjIB2ZDwQrlzYZgddEAQdN8P/C6lAFuuSR
qEOuRvCfBj2e4U9G3gPjiP2bMmF/ny4hZ7XeX9txd2Y2CDcKMQuTIabhQrzV
KU0R7vnnt9VIe7ZpuoVlr/oLwrHutClZ2zcetN/ZSFMb3l/Lx8SKBxmdkTIt
Wx3q01/9700e7qmBYx9NT7jMz5ro8kX6n7lW5kceIzLs1rLDclJLyontkWKa
Gie/yik3+gzazATOSTJjIKyj46HNnUro+AS3FPFVzTHXfAzsAcbWREahQflr
LCkVMOq4b06Y0pThu+Qyj3kJCLGauRK4fGr0yJ4cb+bml5y5CvvOZ5Vswo+8
gaBF547a03Ls12tY8wHO8SSvhYAChimbiypgB5CapNA4FTJ0nUL+ow8Nxk2D
QByGMFKXNipB2y0GhD+2mQmIhbPwQmAd+zBciFXq4RGTp+B1netJDLmNbE7W
SVrBZu+RMsDBXnmtd6jQZLGh/5BtuvGkhZYTG3mwv37osoagL51V3MCqW3/C
YYuzV2gXMAEpuRj5cgdfe4x4ULxWvIHQF9aqezhQXItJRyYRfBWI1W71tuOZ
f2bs+C9hYvL/+WHrTmziH3b8nqiTj1kspS+QFhIma1WKbabteRt456HWqd+q
4l8FuvRpuPPzA5X7wvuZ1eqCwgSmXeEM4vACa820KoletarnmQTOSxNpQzhP
dT5kj4u3dQWwRZG2ZZ45Xhhw2FAWb3QMLSOaWQLvmT+VmdJuehEUTUVMWjCy
4h/TxOOQcgsNlaKYP5sMCM63MZIbrF7CVwSHLiVfG7i7aqXEPLRgTyrlzGb3
AupC9caREh9q/rA08oanF26Uqh5HfDfgSorr43QsFUD/zkw3+GGc/qmqPhAs
oN+DL8JEsAkXBU8qhmHUOd5C51CGeETHyDtID4MfbHZNzCG7fOnzHMajmu/Q
xBigT1wQQlOyf1lWZlDDbZKNMl8qa30Lfz1GikHLHtw10G0OKKfuJ7sEcUTs
lmTtA4XRUu3H108JIhD2vukBD+sPfvxmm/4KV0HVy3PPasuIfm7jRcSY4Drn
PBsdcQz2K58lEypw/6qC+AwFL5iVh1MBg4oSWVkGwZiBGhkDg1bwvypHTts8
zMqkwovGVo9rxuWIFFM/uaMtzabezKiqYK6Sz75AdIMp+JCKsJn7Kek+XQfK
lhFGMLnsFk1lA6ugk+EahX3yK7ne+Q1xSmujDMAa8p3lNdlBLqN7BljTIZwb
tTzd+LVRXVw6JN67dhMdtpwJYx4wRdzn7BKPLPcitjHZZMkD1rulhrJ6DkWO
2E9oX8JrFiEM3Hci94l9Vu093/iqsKd1bUwIsaqtMnz27DpHYSuIzwdnAH8M
Ay0uWySC1e0ftbyfad8XbODQyew49nyJoDBM806RRn4AV9V+MDepmDh9BWHa
AyqOXTYhhETEbe5sh4G116rxJnuaUInfeq12BnqM4zTK9LG2VQiLKnhRzlDq
jVICsD+xSamRbehHFm5L5Qsv6ai6GHLP4ew3RNOmbS8ep5Ud2+RVl+xBhxT4
JrEbDA7IdFQgSMsS66ZpLdBR8ArEjFJxAZLSPpac6H2m1UO+QW8R09W5xlxg
gEf2GRr6LgSf5LNlIrBB3ZKEPSxMSq7iWHvvC3zJESygdDKm5P9ZgZF1FTVW
ow9dL541vbcGb6xNueh/rV/8N/jLoUnY0b/iWkckxvdYzozL6lOuN3LqQyRY
v1u10+Kx3UekA+QpwT2OC6nwcxKPHAHsiEyGu/fYSEu3vW+9CwcDTORWVEqn
iTizNPtihxjNIvklvmwl6srjhRDqAdSwVHCqVFsEQ2PKuR3mb1k8Cp0y7UJx
nTEOZy0pR/HKyO5SVbLIQ54RPyTgqWt/s+toR3514DlgfX02ccLjbIUy1nCe
2e1F6l1igYyxp8MrDskCWsRsPef8Jv4G+uhN+lKtYsMtbMcet3drp5P4AMnG
1cOpQC+rq5bDZ2pPOHpMRwKSI+W3ju3gPQIpADgXnZL1EaOOPC5tZrLp4QY8
+OnI0CNoRuKOcrBRDdjYOjQwQeoKdJbkxdsBsX5jsHPm7u+aHcvKq5uEXpn1
RH5Kw6hFjLQVM8m4svICzfYt7w5i6NLd2gx1YdBjG3H/ojWlPvxV1OWTDGlk
qmhwwcErE3vMM+ZE02NFFlSyKbY9qoFbV5iWoK9+Sx0AxuZnG/MyNGc5gqNC
WIMcK47J/dIAgTmoUy6sGwG5aPkuIWCH6BFDlp1+qIqICu540GmCUtTAbcmE
bDop10k/jYZrBAX5dAuts3Yj6frU09rjVsohi84h4hL8J4dMothTyWMCLVDp
nA3qeI+pQ4H0icuLKibPTGGHsEg5MaSdnCG6c3e8W5Dbum5DmYjo0Bl23HW1
H2PDgS/qTbpmb0Qpx8BccZAy5zRWCp/fw73eYCGNvirMMK6/9srgbtD9ZY/s
uXAVUowEto4VUPy641PDsiH04Klj6C08fELJWvPlV9doG9pQsBIw8PteSx3e
WRbAs70hZ8pqdCfH9StxWqIxzjgPHpQQFdA7m9UvT6gKMbgCA2f/GwuSJvp0
re4jBvTpERG424+xNgI75I0XFl+rddRyjU9WtDcoy8ZWSS+7AXma+S3+D2r0
ei+tY/5Jn8HS2Dw1R29aWtoeVmvO4pXwlgVcENbISiH4//1bdcleMym6mkbw
wdcxwg1l/ee0pctA/S07HW0o1mU5KVMqJaPCQsjxRnkCbxql7fsjakT0XEMK
FvF7Yo8dXiJlDEaXbJ37VeHJ2QKc9jYqzdIvMun7GVbwpHVq7gCRHRi9sxrM
bW5tu+m8wMssnUirPCnomEHXni9DfiMhKDW9FlWy/GdiuiJmYzfAIPUU59RJ
xmQr4H+0+JOPCm/Vgq57CIooRnV42JjSJLYQ2x/3pwLToZJP1KHADpLS+3UC
tOiwhLshop2fJx2BIKw7mckhAJ6EAgxNMm6brGeASieT8Du73How7sqRNR2V
fZHXWpcXLGvTfdd9YFrmPY/tFrf/XFAVA7/8qOTZ8jwX/ukR+cnCn8Sl5qi5
wXIL5+iWZ5QkZ5kUfEHL8WHFTAa03rgkR5lQu0kfZRB/DMWoKpKK3QtdKrps
5Pu/5i5HyoKCRwxpz8Md97Y15cyM/qk6juzKZKOHiw4VvBarhxKZSdYPq/cH
XnALeXqfgUKThPRnTRGfpOQdTWIFX4IC5MWiq99zzdpktdRKX0KNAmhdkOiM
K0NEV5OvE7VSJ1EvOLKn0yVVJr4j0dw2wA/Cs9yVUgIJa0xweA/pWIBE49pS
C51xFwh8uyg2VYC5RWMaROkhJnuIDrZDcGaEIJ4ea4b77fkb/M1j2quI2ZTV
AHEhu+de0jqBGkdcpZ56j2Aeu5VOIFPYHnBkkmMGtSISOJBIsW0UYkHETUQ7
ThXdMNj7GpSqu1TirjYQ0XJZygW3p34m1OhIPhCHvPKeaEYdSho818bs2rmB
jCAmwhe7hobiIwsA47ZX35zefINIcJ55V555AnsgXK//gQp1UMlslSNCHkIX
Va+pMem/oSy2OJqmtYw4YQqhJ9JGLAHZxO1ge7Ei6ow07xPj8aafjL0HEvRz
lJBLJmqRjAy1cAEyATBMEzPg3Iu6sxV29olLmBGj51NyIDn93VZjneFVEgBy
M5qFWpm/XRRFlh0pUFYqAq15/k+bsfQZtwG8SsXN2ig4tBHk2u7L0u35qkJL
EEFGF4GCCVYFqQJOhjo7QFCYICJfHY5MH2YOzFkBqKnRzbs3iZP8xZJDumnB
PphXBSbxntuLjhysFf6uEYn6jm6UifUZ7ymgDCL0xA8Rx9u6zvvX2rdpInm0
TBlfmJWj2iya+KpnXFh/thCIZTyuiNat1Ks84/iEXgKl4LVzvmsghgfACz17
lDCkEJ/bYyncH1eTsikYN8lx7nakm7ot4nob1ZdGddeeU3epppjU4IMyGuul
5liC1iggWdkxITSpeh8OxAbyMwQjRb+40PfMMUzn17jzedwMVsWLhC3bN7rF
aVE56OrlMdc3GThTdMcEjJ21KaSSKwmbZbOEsjsqnr/qLmU4g8CFG4sy6z3N
Ba2++OwJ3/dQAqKKyIGQMofGl+PKGQ8KRX+kqx4Cg1zP/i7Gllcca0o8EP+b
EcsxKDAZ6ltjiZZRaz4E67QDaqJIfUHzezi4b7NKVESESPbQlLXHDS9i+WVO
PKyJqBVlizY5MASDOs6nSisv0I5i35lwv3cFMoR0da55PRe1coZVpzpdopAs
2crn5/ihO8tU1rij+3FrkN/k3HkpJwEFVWbL2uAjIsLP4/SR15udL8m1aMmO
alLkrzrbsk1WjuKMdCkuRUEeTuvPnUVz9+vJdE2Xc72q5tGHpvK4QMQWlk0G
WhgtW7hiz9hfQfIZUkQGEXZlF2J08Qll/eNElwRMBM8/wdMkAw6dR0GE4jWb
VWNKQkis74suQR8xXAen0fFCmTCnwSti6H8ZsQEZCjkd4KVkOiEUfQepRpcX
uYFUpDlAkbAybd+JN61ZWGX4OWxA/apll3xJAeXEYy5lDBIxxhtF1r+Ltonj
NJpWaI7hXS8ieMWPkCdGCyznWFZD+xzFb0ROCfgsVt9GUXsK4DH+bK9H01gu
2g9YeNM4hoqkBvV4rX7Ep6cl9y9YJTCnNz1+bqSbKcZKfNKSGNJPRSIxrvQg
msd26oiyfyf8r7+nGy/R4DERzXbNnOk2ob6vV/C8Clwct6Pn5ckfOQSCmCSs
fi+A0Ewswj5Zasu6uMExit0r0Sh9E3tymjhLdknVlUGcO+wr2nSvv2xCWKII
QL3kC8LFR/txSozptsPpouBL/iL3UCnbE8tvc6ow5GUcjtWfbKdFNPaEJ6TY
giHc7wtzAK/+hcNL/hXSXV2kURx8qNGBgft1khitCbV2oRQpSdgle40zWAfJ
e4QmwEcS75b2zbODQv/TnFkMlzyLFXA2dv/qntcGVdX+bnk5S9C3bYjHBWd5
w+y0Qi9D/oDM2A92vu+Ug1ieeLENECMITZ5v3u9cfIwKqK7ytNVL1mJV7txH
cz0tt9SjWR48KZMoknVW6Bx+FO1gDBUyH1BtWxPy+8LPU5uLoqqnyc5Vnz3K
iqcSDV7T3VzRDgv0OI++tft+B13XrbJlG9OK6pBMzvZtHP8k2D/pRkXrALTy
uPL2k23HTJ9QzKOx4tDFB1r8/r3MOaGDv7sRZoXlhGpTGcoEtSv9AR7zVZE2
mBWLsba1n8X/JHE2uGxrWiM43YB0pPeMXF2q7rc7tUwgxpedTNsVCrMsJA6V
s8mok4JQG6pXYbWyVEGpCPjDTnd2efgxq6VtRNfEik1LfXPXBBem+s7Ns2kM
7WJKe8HZSjpzwjrVxop/w+DLLyh1WgS7NPCqXm8T/5XepTtUNOgVF3mL5oD2
P+kIqOy1tv20i6bp2xYalZ6G4vftiCI9lvjm0Cpwzrhjf2l8nNxDpd6mAgmr
HWxH3I5qq7FBhG9kGOCLIdZHdagOcYhyosIaK1a5w7jFV9iRx/nVoB0melud
yZDVEsKs7d3xnnYVqH3HT5r8K5LhIwqvbeO+8ZcDuMk7qOy0ezbOPlsKYwBm
AbPxW3XQg/+oayM/flV91LFlRyBPkuV2iekEuc7hGfTnw/nCxGDRDZzMXsdO
ShWDXiV56AIFGQ0toV9l9QYHoz6trsfWD53xVGiDeZ8EMJt+2vFSBawBd9CP
QF/VfbW1B6e9X6M+GVlLIRR/JJs6WTvOGZuHrmArHYNR3d0HmHJZkfWRD6FR
35x+RRjrBpg8YEIHaHIrcOReAwjvSpMhIlCogTmr0nHGjY8V8zJAuPIjmNS/
JvRKd8NvyGm7m08fXzXQ1eFzsb4obYxc5gyH+NN8nc4//WTaQv4cxoMwwEFQ
EKV0g30GhdMGlvaTAFOmFWksWu+zpC8P7ZhrtRi6aOOsceIhtDKeNssW/x8w
X7v1yvvOW0ku+F5TOZCDnU/Y+e+Fxypzc5A7giuDb+7zkuQy66hhLhVV7/EZ
9IkklO63mJhr4UVn0e7AwPtV0w3Gw3okOYmN0omLfAo3ys0ToLfZKSicSovy
p42XPEgNyZmhoxVAj+Envxl6R3a/ujE2zUGj4to77ZeAojbOxqk1Dk1msB/d
WKRNO1Bffqj57XXOq2l2GjPq/hPlKtzLe2WvEUUgNYjvAlN8R0enHjRhnbJn
EzSf+9ulrWKbdi0S1t2X/fT40UOakl20oFHD6o6XOVObjjReLAI3Ua1xkDVQ
FvifwE+tZ7V4JcKXiaXYjXECV7BNNe6ZliKsLGtlXvBf3YeKszxoLznxxUPf
mWIsycRtnKEmUISZNdzZENte9wmjUBVASY6V9n8Gf4k3C+oplsOtWo2xI/Xf
Awt0z4q8EQgDXAnfYRYwx9gQ9tIWAvN2ud0wnzCm32uWmBKB7HjQ+DIypeJI
Ga4OU3Af35t8Vn/ACp+3tSSWsxdFh99QTzlQca1mYzDhVwfaYgI3hh3GPPtQ
vkpZe4Vb1KJ3oWm9LRCjS2h6Smu5O6Sdx7mOUUnp/9XeLBQ9EnppjSsuOsoh
XeSfL/r3dAQzSL94vnTsasH7QDTW5xF5SAeuEovjA25iz8zvaMyMjkXSBayN
uFvIUtO7ZkQqMdTpSx5pY4d9A6ANHR+LDk7TcrtG3z2ilvJx6swXaOXt1lTd
PbhF2+ZZRxHdIkpypMddnjA4xiGDpPFffYSvTkxS8X/loPq23qM0gtos4z0y
OM8gBH81zXNAgByJReweD1dmtoC9wV+hs1aqzVuhwiodAAPK4copZRnOqggu
pgDUAtbT8e/hB/k+Gp4gOo75h071OiGxvl8AzoayIofsCZJx/amUqIgdOoq9
+XGdyfkLAb3odxyjUqKu/VdM00dV6bOZIf2MfzFChlDoZ51eUHMMoE6jUH8U
tg3Bt2ttSfy8pBc0kvi+YOBq+CFKI8CBvyaxxtpAxC48MYjZKeW99Jx36YwX
Ma/pF7RobafMsS5vaAFwbnceluV8RWcT0QLi73SMgkYPk0Lgo6U5Mz6hZryY
B+2kqxNcGaEl8AxBhQB678N1dhe6I2tuUEsoLJyQhf3O/aQqqrw0l2eJrUWI
Q8ww8G/cVDLvvQoakd+TPizWGdAx9oOJb+uV7fPAkLViVL35QlC2CiiMS81w
CrRhH2D+eFMpi4dVNL66Kfx+v9IczZ98QokJxBhkVZEV3yUcsvDA04XcSfNc
7JKVggNBkLNbYSzNfCnuIhPmaoCAFghWqS751LAQFOhlj5twTmuIX8kBN9g0
/5XbtaIkXmbWnj2qnTcfOS590LCyqIUpmgDeiJwMhaBIofcTkUh+TIbeMig6
InVuCahYOkA2XFsAVLCNoXQ2OU11hYvQLuf9Oz2ishhx8HSc486/10bUiXrz
6BC7L7Zg6zvCnjpUd7sO2PEK1LGDfDIt1OvBatNV5DVqArmPxjVZ3YD4Px3t
qLF4Yaw6gKPY5PPFKEusXnpkEYSnpNav1t6ECZcKZbgHdRlrjZVgF3S781Qv
pL51PmwM5in3GQH5d6ORAaQ5TdTVns5t9zf+qrRn6KWhX/VdyaAetzKNCtTb
5FvMGIEjnV+ojEN9YTleFPEDBRVQcVdXbepGNqvRycuuQVYa3BtzEnc+FG+E
pP6wOTG61bUIozeRycJp5wEjth8H3IY0kYC8S9crYMhQzvSVwpmJI+qep4P0
WseHQOs78KKtD3pZ1fI6YonyCNINBL1YFtYRUbKsqQ+/dxvxM0RqRDMJHBKg
J1sT2lNjN6iFiiuT7M3O1SFTVfZ+MTYx4JzeUxA+QIYowtOCjmkjBENL2nqP
IFZnYXhddwvp9urFJaZXFjoLwGy3UVrLo0Sjv4pP3jen1tMYHusfiT6H80CC
5SZQO5Pq6XZceADARlOIFH12ieroek9m8fSXnevcqIN0lascn3QOTLexsqru
+Bc0wsRWeOSYIPziu3eULujJXPPTMjcJQMiMWDu7Xjt5ft2ZebfiaI3aiOnr
C9+yFBz/zLqqgl0dnvWb5abVWG52Jsx27ZgZRMwCz9zaYnhwy7M9hLeKjxv8
x4RP3lpAfOhTdAPl680alXHzNq86+B0qtn9gtLYyl7eENkJ4BkdeJRRXHUH4
FALOojJ/zhYnJTntCmIDEfaC+5l8DCVQGxDOpcOSYsnhi95xSOtvsstsDcCN
s/wOpt1TJ3SGQStEjlE6jigPRFBkhhc2dT3DS0T2YiVEhFCLJ5Jba84Vb6dN
v/+GmFmF1x6fx83HLFW8dgXMp6GXZ1mYDdIbpWXv70jrzvAf/vN5KiFEIVQc
uMJW3tU/C+AAoAMJxwjNQxT8L2q2uWxdi5EUY6TWfOSSB6d6D5oc+4yyG9c0
fPJZx2tw3dpam0k8DO46w+s2Vfpxuhkv6u7YFR0QqOlQOQM9ErfASbRseoZz
WFQcmb0VswEOo2Sd+BYRkjwkW5tz9fOLNDzHF+7MMt5CT+Ide1NJPbrHLpMs
gcbKx7qXKCzTp00mbq32n9PCBr9tOJeBYjZ7m9jJ5jHKGZ6nONOnQ3wGRUbr
S4yqmZl2cXLngKRrZJ7XLumWXNBrNtT2FM/wMsW8to0/4XdsX+ewp01o59gZ
P4BhqOcKvh0ltaB5/XJApW+W+yEJArt1sWF756rr56qHPiI0e4SLqb87IFlp
VCiSCb8awIFRWGdP+bOzJLrCeA1/5X/6kMBCJ6OVcvnWHE6/xInb+xWUz3dw
uqr9HovLglh/RamlJMj/yNxWbnS8881JoU7Uc4bPfug2U0MGUM59okL8g1bs
4Gs7df177VvBEfVAu+F5vbUqCjFSxnQHchaNR/JSNuncx6kN1oIc1fOt65HZ
R1930MzWO8i74NpbQYp64NGQz93a8JR8M3oMNpF5LO3K04nd7DwxgEanzhJx
gnz/stYyQ/ISHaPZrp4k/2PywQAhFvEwQKFu5o1QFfEsOKwQBxpcf0B0pAEb
0eED+191/Zyj0+cEdPRZ5F7OLuNsdluCN1Gr12b3SelFoSyfQAk80TYf1knG
5lDyvRYB/0RKmDeHKHSxbcDINowuY3cSNJt9TJxKNc7qQhOWtw/iVeZqnMdc
jPcOq+nv1O4kq4fDjx4YZ/M0AZacddUS/GuOisD25Nli3HZMLzQf63DQNzUL
ajCeQPPh1CgQJpaTYRBXQ/mf6mvHMMdCMdYWVo2Dv/U1ntEd87D6YKjKmqJm
fd38aE4256mzTs+9yUXgcfn1Zkel7sE8C88CRZ887H3cd/FK6jL2+vsO8ayd
2sgB/WdVbQz0IDQJbvbi3yv7a62y9FNK4kdmZGEeKvRHLZ9BgPd0jAid4w80
KKzwNVGp4MRNPX0IlNi2wukWoWwwTwTGMCSUc8PHEK4Mp1HyIT1RMFbJ9Amh
ko7FW5oVt84Gqm6bYfPZQldLklYx51Lc0QGXEgWYL1mZZSFTvaaXFHQGp+Jx
wJqgaytCV+0sj/gJ6MdKbktOUOn8bczkSsnCFOZH5OlacEtX/4DGJDdxzTFD
YD/M8EDGCM3WBV7p110IbLw3e+kwbN3qNTp1gWuHAJRva5/pD6Va3FkhVZhs
xHxv3BpI16xhH/d45MtGEswzawdIFc8a1KTgsOmvhmyIphrfcdX2HWm0iXox
BOL6l0MheTmPZcWAyN66L3NatcAUygHkg8qo0jwu7DsXsFko1uqJm7xVGIMn
DXouL0JT+S8M6EIN6hxZvM5ci2auMOtOP/NO53LMw7JTONSUjmSjOYcxngBC
9sALIiDNyhGN5QGRojC8cIkjXKDs/9t96QM0EkEF66VtLbcDm1ME1iXQjvfy
i2OG/Ev9RdJ/xgW5lk7ruHUOsVdICsKkRs9V1l2jyszpazJ9oURIV14zjBWo
m8yr5Fipm8AjFiaei/fvwhJ26zyEnTvfs/4a9qw0zVSwcU2a4017is63sv/n
EIzfVYI60Nsc5BQeVyTwQ6QwCbQzB4u9zO7wOOKqXC/rNPgmPtoVgJwSscj4
iR+ev1/P3A+VeRbjk57cf5EcsZaeH+xcHN/vZ7fwCLc2574ayzU5bRAHzhfH
+QRBweYZhq9guI/xPp94Kv5/8mX88JYLrkTUxenTnoFq9i559ZDKNGD2RbIL
AcAScNNVmAugEmX2h1AzNcVDHWuySWcX8KzPO0AaUgaN9Xxe5xQKiCLhZuUK
tTUfmNlUbLol3bl4ssU3BSJx1lOiMiLBj3sb5nWzY3muH/hwRbPdejTgJEVr
X9a0R2db6UzEtqeBAD7+N3aLEvaSZlZoBw9nMuNUClw/cuVxPNVmDzFG0Xe7
Lohr7kEyS3Ofm3/oDEcFic3p/dt3cKRLbqic//sN1Vzs4EyF9hbhT+i3vgzT
mzrqKzJ1rXFPfgUZgBOpvi6243t2p8GkPJWVhXsAsZ3ZrrCJqDVENADs0UpE
j6fPoNCociFzp6HKjqkz3JCHo0Ih+K4nv8A6J0Syg1PDDFwZJYaSHU46Qig+
kmi9LO7rbw9LF+r9Y0TqF+k8YywvkHFTSDyLpVd7TA4bZiE8/6+GTzBmJKYy
qtNgITjSkLH2hFMjdn3ud4y2ghMMhNSkfdgc6+rEXOhTz0ENLYQ7QBbzHeX7
oQ/G84g0MXY6zqnlPQPk7aW+hrp78CBBuocPxD74AUgDDidgbKbNz6D5/gtm
QLSGzENOXPi/gmjCDEHSH43szdDdUauiuAf2cxwzcqfjSQcC/41+plSkZdlQ
KF/RB+ohHUtJWigyficUJ8w1Upa5G8/3VmF6xS0o+gUzjLM1/ADHNiTwJIq3
wqr1yPM7A9g0Mu3T87SKK4k1+sLbseDl6osgHbD8+vSg+GvjVuNqwnjlULE8
6hDuOw2xxuHFY93uBGYt5ulYut3wveUQVDWCegVWc2pjHdCX8UjlzaraBkL1
j7bqBMxaZsNP76BYsVW3OB9JOQwNF1d7IbEecJ9iPM9znWxC/CVaI4LVRYUm
HqXLdbcLLgXddtszNHsR0MO4x1FIRFV4HRAa646EX2jKG5a1MbKNCo5Frzmd
s1OfeTmCfe8c0NOS+YFdSSJSrnr6QylGPGtmWZLEkpb0rjCO2+xsJcyxueGg
Vsl2imkcvMAg1N2qZEGFVP21aqMeQiFsSgjfoBG9MxQx5WK3et43RFBx7ShW
g4SuiOmQNVXrBaB5184e4+qhsOXiEUT6fmGaGFC4wDkZjQGgpYTzrvQccOLX
2gjcWJjQUoVI+VjIQ0yaXwof/KOzu4IE9Jtf/k4Ncbkgw/KLSVqc6yw++i5M
wiBDfkfcx73j351uZevBYCQ5u1KcNWBZ7ieTsYYqBGv6gWwmM6IygWPcULKf
HU2HSVomfnMJBm4tr52o7YklocWksuwnkDCIfeoPhJ1lbLlDT9TKqrgaCT2Q
Qii0ElHPU3tCGh6sJOfRCVFIPTZ2GGDTnULtuERZruxXwEtWEXByRDI+/7eu
HTLxzmyXQuV0628KFvDGM2eK7yIP1PfjOFwgpj0CYL2bh6LqXOmprxCggc7J
3JakugG49Agoydj4ceAebUVElkoSiChsS6L7MXLCJVeOVsrUSAqexvsZmT7z
9+12VZI/Zl82l+9XC8z5JBYHUy3VArPwuCMpZ/UlrqfLs3G1FlmoDDaWYPL4
XHAlD71WbGAf4T8E4SSOfyI1Mij7ivNiNDafnkhaU7D9idzslneesLlOat0H
lB9vUAXWXRlqvodXR8rXGGV0fRz0Fer9YWFfDE+h3tHnAJ1ExXi9n+wbKb26
wBwr999bUTsYXAUQ3D8jBBkDwQDJoxN1S+ygkd2GwmPomS7o8MWcsF110DZk
QwTc0yb1M/detM5dPxuVFkOHxWxG7s8Tl3aSiqfR8wtK3XO+MB/a5JuPLmEw
BW7nabm8ZOU94M7efVJSxayXMdKgO4+aHFIM7YMdpOqPhzZPxiRkLpl2mG/f
7/t5AjwQl+dHAzwK3VOmtAK0UEUKavucY5Tp8zpCrs1mFoN2q400jh4Fi09M
HHZH7+wH0wJBCs4OVAQAHi+YwZ71jUi7wnHuf9WSB0poXmVVFrRiuQ5p0oN3
uRNFPyoNMRFwOAasFeQbFyT7AtWJEus1nqHkpV041XF7/EaZ9hMM2gjE1wLq
lnlUcmCR/Y2RiK/+XFjhWMZhzSfw2lY62oWV2B2IjSTP9QO4U2YDv7r3hnEj
ExOBYyo4OqRmaNzaeIuaKYMjuZiIF3iEQ44BEZ/2sftsXTcVf94Jfhx5Ra7v
kQ65FB4R9s0D64RGAJVGbMwRsidhUl7Ekjr6mT4oh30/pVA+p/G6KX+bjpaD
ovgu5g3EK1zHgY5s+c5CDJ0CXd1Zzz1lVYZnzFlZwLypqBiYJAKA3qTdOxo/
TzZ7QzlH0cX36qpuORDHd5VhhVm+2E/Rts08+Ryo8HYhOngco55M/WiyD9LP
OPhG3GiahezGg7OJysWIXfE0W4hxEiMuQyCslE5M13bkb2DexPF3fjlhaLM5
5tqNPt+C84oTmANEuSgbEi6wfJdv6eA0H+C2VOYnLeJ3Rf5Xxlf4cEYOdifW
RPC+TGcLzlAodBOChIG2QC39ly/cQMeUyIDbEjxlukdpEZpZK/LaXzM0QTzn
BLR1d6YvvOrwcKWgrroehFUTvNqa0DBZCQV31fKdC5xb1tpUIg53DIxxy0QG
BwZrmG41OHFZN3igdytdi7W0SkwVMlGtC2M7nIoFeNNQgdnvKQgzn0LZ9xXn
kSCFdkx+lzuvZKrQ7xIJb0Kd1b+G5lhaVIcP1ykSTjO3G2TMwtp9N+tRassq
UzJUJMPdJrDqocO2NBQ/6XlL2TMCF7ipg7k4wgp6yDHhQBA/dFJK2qvlBfEX
HcY9rnveyM8iUBqbIk34b6CKrX5WOK+cIOXmsMRM4nLtrkuMG9DX6B67j10j
/4VoEp60sVs3s5xMMou79vOT/gb5hhd0EqoKGf4RvKIR4HuvcjZASLG/qCZh
odxQQ1i6dxCGZSSI9gozXht85dpW715pihS3NOhWer+XWEXzU1gZs7+Aozvr
ctD0+iImvud4ZWJ6A16/x/LyAnMjl1qagUcl9Ih+ha39ZAffv6c6JXP1dfNa
G0PCcZjAfmfZxr2JsKmVpewkVy+ywIAsUGgtlhNYpzozhteo8IQL67FENJJN
a89WkKn/0FI8JK0IsrdYiTRTrOpW0Q52EqFqWHlMGmh7Hqm3I234IOWquh5x
4PSxSl+RBkZ1UCiZNOGgGePOBg9G41KRrGQQYOCZDiLsShvv222JfIccXlN7
j7t2eK2hb+dN5u2aStv+goeh/5NrCBckYTOEbB+mqjUUXE/Km6Fcmx2Pzppb
WwWRxB+2LvOb05sbi07m1znMhuOIgsZIlj0aIZcuogliIUzQ+gqvMQVv1T6b
qYC5w9Jf6jtxz0Q1xhXM31x2ZYJHB/h6EaLJYWAwOYjP9fu1iAhTWVx1niM8
3KVMCbHj7b5iuZzO0beyXzlOsEJFwfM85zauyolz67+ipKp+ZiUIPGfuMDDY
EEKmHUm6Rw8W1DP4XwF3oeIYckASXuUmtl7u5imXLJIzB3l3UMX0ijAcsj0W
pWGfUrPaWLjrvFx9E0HPg6mnwh2zj0eiGMI3zQsOMpRiGJTld8MY1E7N1hB7
2INKc8A/AfVtuUVo9ClHyhNgIoGo9jH+iscKAFwDzpI6LdCa4kDdHtrV2zMr
BeCr6JiT9dTdS2vnTAbGCqzBBYPItbJlFrDxhtOz0d18q1I4I+kbSGYb9dCe
hp1sDaE7b6x/tj5dJuf0rlpjcDnFf9uJ+Sxe0Dxt0ERv9MuIuA0o1y/o1olT
oNLu+t1QPxbfueK+h7p2HC8I5RAHbn8ZcRo+OJ7wtk7lII8g4SJUZqRC79MI
3Xgc/9FMoEgX6pds5k9eBOcucAWeJuAl/cKPxDYXbBRWupIBJ/wyJ5MIFaMl
/m6h8tyeIcqpn+9xvE2XfDKQH9dmEjDG+W+msJ1Z9Vi9mXpqEzJqCmW3j/9p
ZuXrGGRqqO4xyJICUs2xfrYoJmS1eCqVFL5GxRYhmn1WbDv0bZOMLOR3pW19
7k+5yktwSz+D3lpDzfvjuSzarU/+7/2TyONrEhVLq0AHh44sMhvrXj9fx/k4
9pvbp50ITt9S8kcUJ9aQzGCZC7XCIFns9u+uygBxd5i5gRmfZkGES/0LTHxt
A8ctgMJdQmb5ZeJ3hjDcKb4glQMgwH8C418cwY7H+Ay+URn4jwJ5k38Ut4Qz
pyc2JVbJsINrw2Y3igBNFt50m+1G7m1OhmV7GorahSz6ynSARfxPqiGUTici
T4T5r4S39as/w2Zi7iAB6tGeR79oF8r0qynoXymQ1sRUpa/pwGq98rIq9rq5
yB/GXi6mUERNtoaAjyjQfyZa3iyEAJ0f24xs9jQ5/PJSjXRtxczer5uOaiLH
XDzjMmaKV7IVFhLh0i+6M2VTErw38Ek6ytqnEzZHVU4vxBvQ0WTpE3BPzISV
7xnuI4aCRnApoXaNny1fTfwhSeLudIzNeigWdxz5iSytdLBQWmzSTHR8xQe+
kX8XQJIwGlbtrHPZedioJAldO3KcCNMwgbp/vPxX6OLqfTgHQRLQJgVbMB1B
oH1X5ObIfRmDW02oJBfXXZZYW2eYDa7wTPERSHh998v9zwq2E/i7Nh5pOnkz
+ITzY5ClwPTiXvBkclR2a3RLt6wa9Q5R6kSvpe9Sm4qBjeI08OE9D+OVqAx6
teJnKYErG0Z751X8kKUohqVoElMZrk6ww8tOTviuDa5KJgSrZtM+6dLBW2be
hjtWx9unWTjtQTqIrqYik3nSrgO09YGTmduNbgOPQA8U5gDQa4VQuKQENLCS
VIQ1wgkEJG4DM0hN3IRDzMOzf2JJ5FqV0frv3k0ejeI3SPLiQpYZZ/tHFYwh
1mL8BPujnlUJ51N1D0na4fkIigHPltkRFOR0evCpcL+Ngd6lu9sYb32rYoJI
PMi5tNW0DpW9Eh5qQUT/CplyqyRHpAGxfodbBVvHd9Ur9LWQf8VFuk8ukA/d
NLgvkjohsNSSwtO9zaQmDw1l7CTl196a1hbqJY3HMf7JlADrMp0x/nDGlYeA
1FsGgnKbSysmeJhOeaCjKimMd0/1LGaQl3Tw4/Ymh2/QBtDOaW7QONnJJd8/
1dTTZ87NkhZSnzYhb84KUEh38fQhP1fHFYn8PYWyhK44wsCWXaZkGnCoJJd0
ZbEicU5IYYvvctpBaOnjtYkl8tk0tXU+Hz2wyE1FxWupE4vnnmwqPMNXd2dE
2SBZsNQAzcKI/AputVGphet8xMkTmEQnRQ7/N/JRBKRqtq8Epb9k0Q4Geo/p
+XzDcF3d3cauw3muKD5F7XkL+ls+lNnROJNeAXCDavXjaC2d0A9epdF/zwTt
mDqtPEclpnnXetdlCKDMib1Y0E28F6fEEAcz9ijcCCj99s5zR0JC/Zrp3tBM
0B6Fo1DvXVGH6LDosgHFqCLn69PP2wE1kJW/NZbezz/a1J6/U/RMQDwoJq6+
SCagowGW3ZjglpgD56JzGi5ocK+Edbk60ofTHNuu3Ok5zfcJdgCgYSfZ4rG6
fQ3kBGYin4HQllhRWC6WrZtL63ziHjSo1FwVHNpTnYWWshN2xnMDC1w3vuev
2GgfM0e9BOY4ajDJsu763mdXkWo5N1KtlKdYdKCB2gY4ejTb2YfdUq/a/JQ4
EZMnNJpokB3KLdGk350J4B2X6E3kchyL5nXveUiX737YIyqkoU+v/B/n7VEZ
J51VYAvnz06/Wpdsg2LfyfzXyOmuuWbhW4jRTJ0qUzJBP19uFe9mFnuu7wny
sdkYYrJ2x82KL+aQPQ7d2e5tLak/ehHXRHS7V+ndXlEiJd05cGPFuxhF7F8t
m0bV5YAcmUw1WgfXcSOrkbF5o8tlh4ox8wBXYI3K3Xo/ee8DbbY4vy0nRg7V
PvtFmPW9TKsUb36NLYIKkpRgqB9AU6vexD69UD0+x0lsFRFwSoNt88FBdHoj
2OZFOFz2o/lh1pU/v3KxlG89x7Dw9iaymtM2i6iHws6ZqPqX1x+8Wh4M6luF
psTkozpNohtZGZ9SPh6N3rfVtLm/DX2dZ1HYe9heBOBugGNqlYw11wwk4I/s
J/rFLrVx2Y4re2nW5iKoJdTbUyhu5auMbpnEPOm6NySxu4VsRVwUzPfiQfjI
DlHK2Q8S/tcEZvDQnipOhVaHAGCN+ZFRJGurwPoK6cZnQ7ojk/3roW/2JUe0
PTB71ucGhQO7V7barDUe6X9cSiHe3f2BozCvsSu8Dwomjs2TRgANqJswp/Vr
FXuQ1LHK9ffrH12ke0nYKGifrKwEosbs4NCcq9aE5vRvnHXjxDZzCWDP4gdb
Y6ipJu/XyZAH2d1x5rHGnUPgKwz7TJNQerwGaAsueGN313hHqWGM/wm/GXGu
HoIZRbyCgFHbUHEdUrJxq/F8d//KfCBLNEwEkgOq2HtqgFxPYCSDxxppXl/8
UNaMClqdLCV0F0RJSBUqhMjSGBZ3+AmTVdeJJ4WLCkYKL/9fZZSHpQi46BID
dFbZvZFXNXslqC/Vu3JEipC7TlLvpGN4pwizGZPG2W5kSmwQKaN4/7uKDGKu
ubqU4uxLBts+7+e6mK0+3CD4yIWzMALU+1V4NZk62cEpG+ho0TB2V9//BLvt
MZeTVaDxkuOOLQNzTe6f/gqCPrV3WO4uZYdZdHVqNmZgBTYj0TjoV8qolWCC
ieHnhE8HtdJPVeZYFFmjR606TuAuFDuke55EpPRUb1b2lhbBU1C7YxY4/DLq
RUuBiBQ8JA8EFpQ06Uyvej635bMmCNmtii090NnTES3unveBB9zuDnuUh0ZG
KtW6pGhecEjX8R4oIe+QTjM2YbNB0TXuk852XHwZbmTCz8agd/Wd8fnQAaqz
Ov6Uo4YYvG89Ipc+MaOacwWBtCLOVWzfaJ4hVUCoBjD+YSDUUuRh0IkWYLlR
plH7+pjU+BC16kFiwR0BkkL8mMxXf1YZ5X8xHR57wEHL/DUsqRdIvrv/Izdd
/uEhb5YXzKRSY/hwZIB23VXlAMOQzdyDIf+sW7rbv5daLeXR2R+VNMT1swXM
nJS4L6VSuBo1A/9YpsES5hhr9M64t9UedvsQmSs5o/y2jEsQEkaNWu/GBq9h
LoltRWRpd5z3j3ElQdsf73lMCXD/RWU1AyDUnFx3LjmO1KIxgOLGQK1ByEYu
hvmLsil4nRfscIND68s5Z/MNaHqUNrNt8dFnJ9JLSOAMLH7qmQlqANBmtX/M
BzJsewC/oXWnwvjQJOtMvqIQtZO/2Idjc1mhyS7yuKpqgfwMdoUip0W24zXd
59nNQQxx1795kg/0fhaFB1aScdDN7txyxKhQM064jYSrVbjdYZPYiOAoJesW
/Bw9NjZHCMg3G9CoWGiJ1S0gwP75F/ueqhz30TXcPVL0t/0DDLj/yt4ih45t
rYJh/s7MvrsggWSk/iiZWtHhuKhgD7FtFeLhASeQQNBtZEzNVzVZz7NBApUf
mOsby2VuaNTtbzYjkG+8k0d6knoprL3d1bwd2b974HnWIzDtIpmhNrMm/hRH
RhEOEOpsj12g6oTfjUZeeIErFjElYVWxzXtW28ytOQ9HQqDiJF/JqonvYENs
xh09v6gyavlQwiKhkvRaVtOr1W8qKJguslJ7HUEEsQkypcGhM4v8E2OCAAuy
Szqz9JbPMU/Sf8xpZE+GgKKz/ugMcwpXYtsidle13ZKTJERKHWuwmg00OQGO
zVCl8e6IrUxF4Lt97DnaeROW0w33i30gxsslKBsn4mzrtDkaN5szaYMdWsFX
q+M6yvg+0bMSLWH4vsIkPjBwm3ZkL1rkTqvQ7eMqfgS4norH93vu8/4+h7WU
Ju9CVWb+aIfWA860hkrZ6xIAuP9wzBnQmDwjjkGxnbtxBf9hBVStJpmv1OOE
ZNG1dVK/iLEg7QlZfGYdt43X0ZZtDSud1ggQRAgBsPpmB4ZRx6mrjxZPxugp
o+EZe1KMfP2K6blt2BbHBe3MgRkE/uCQ943ogkHOqBfPMR0zH1yXgKb7qvLb
UrT1OKsz1Whpkf8y7EFkJGFf0iifsXrQ5zm+U8Jav2KdT+lrBZ1PREE+TtgE
5fMX3wVDUDWe6OlrSvzx8mPUy402uUC0Gb9a1/3BeuX84x+zFG1Gy2HrUD7M
d0Zsd0ETiorfaLBnScYJRc/ysE1e7olElOwV1g7ogkPfrVlarX+cxk5RVUiD
4TpAGgQWcQOisFVJkg7tg7GOQjOOgV0SN/af0umbKHr4nokhVTCA14SW86Kz
6LzQ00xZjH+Z/grLdNyfwo6ACNfcq8OszUdBcvZnTMFopygjFqPnoYKthlOg
901DlaA4+l0VLeTEidatohz1HEmclX/0WOug60MKCI1k7AoneUc/Npztur5r
LAS7/JEaFDPQrgLnvFNliqJvd0us0Go/b5XWWkRD/OXPuHNOltf1xhj1qzsi
PKoFE9ROOft1dDUw0H0r81N4I8oVaftoC9p2fCeK6wkQcLM6JBtKYbT1//2n
XsAW2/mU54i+pvScPRFhChh0NUhHjJU+BVeNmEyc09IXRlhBFwe0QkpkXpv+
P5uE0cJZM+X6JgWBiO82lBV4IJEZ5WrmfL4ba8V1Je7VdxPv8+eO8GHHGVcv
HAk8lmKNYc3s4wgLfTj3C86+0tAoAjKp4D4XZQXWv1WWb9td7wCRdlNxx5WZ
9R6axzClyhq6a1tPOk9H9bSq00ZaCpjwkHkCpjxTBPgYP0DNLijIqws95GQc
3wHuXRMPNSSgPrvZdIyWOLop+StrWRkKqLsOAh4MGQZanyw4sBt4NnxRxGXM
P9rgBiQQS5GkbwEfGaoyFhVBlakDMQFj3wyek6HnP30DP/516jMD04kqyoze
PU9UTHOy1N27PoZLNpco3qClQsVcx7gSkvEt9FgkL1WuSRDlZTm8RQFH4s6L
tO2K6UhRkIfAlIA5Mj3xTckE/oPpX9VowZ2qM8KpMFULWxajNm0YLuEjIfsS
pINXmFuU/0bt4tQC+Dlg7tN390SqiNtDKDO38WTWmeKPKlf1PD87IYWinYNm
c/xLbcKQ7Zlu2VFdUWDUEGf9FisKdLonqeY9sjGbSMyZme+9UFCoGTxqUgJI
EcBOe0feZIITLYklmKsOefC9sqdtNoPujWQtxdKqot6Yu2xYCi1ZEhSVPP1W
lVbMzDVUxOXpBMA8ftdEbJZqPBK4ADPzYAYNyUZOqpQyujKmi+ouNwMvHD6m
4tNNkorNnt9zKqNINF/EIt7N5K1k6W9PstZyQgvuEXBWp+Q8/SYMzkrqyqqE
Xn1CDk9gPYyunfZpnINBu07mEfbEwMkksiQs25KU5kI0iTTXDMe3+T/m/1Ez
mCHTB78Xa/PuyPVCt/zcHYxw62cRH2Vw5rWS9FViH8tdHUACS7r/y39QtHsr
bpI91QrubbaRfETogkPYznSifEKIA9AdFq3n0uRNnNmttxtFA2+8Omlexrfz
W8Y42JtnX5g4E7YptRiqSKqT1orTXrtUw67SrCO42bKkiQXZFaJFfSUcVtSI
iNr8pGDgmU3Ci2Y08YLBdjJ4opmOH2eYkVd4oVg+b5FKqZ13wuuzykmQh4L8
3JT32F8Vsg5ndYI7CC4qEHWFTxZluEIHeN8nymGDF+pXpyu+WAtL48I8EPk/
6H3SO+QGSx+Lki6NGXO9nUGu7egi+8u4hGUmVJ07bs7MbLEmWpRFDQih8S0l
nonhyy71LYaGz5vrHpJsbGzjfCQehQoiVTszD2SDno3XGpusHy0Y/om7G1iC
ebORo1xzeM46GRkHXr0SsRtrgGrWuzZH/i7oKYM/mELELRddT5JrFi1SODA6
l6u4+9bxFlE5l7eGBY9O/6L/+MFDdAQ4j6mHsO5eCipimPyleAVrD0gqfJBl
IxW4Inax75glSfjkDy+/LwVCvjMIVG4pidjwWxI1fF94L5r+ZmEfNO6JRrNR
C08Lw0sh1HS5OF8ib8zVQJUHeXwLk/MvxrtSlOhkP7PAbQBhu3kioXfNkN7V
YS2l3Fe7FP7wMLw1m3g/leWsCKXztmxjC/dkMXY1NuKugRWvjlwKgMPBkuXM
sZyovMcgVVmXT4gNvXvv3lDBsPZGpfB1Z1uQ/j2c38pM+8ipCuYiPk8QtYi6
b+OZHcwBnETECnfdtOjWu1POp8SIZhleclkROnFgQWODId2PR5QdINUhCimZ
2/S1r6KpVzPpGfMhAlNeRPkRyicygCsrDUo/lkU8c1UDIvlOfPlpM2q9Hlsc
SKsxeqRjdjh6tgoy5ETKIVNrDeB0sfRLFIhk+O9qRmPbL9gyRyK8/NmFtB5e
FHy07xRaCK/aRR7h1sVy4t5AFhYwhBnA0K5LJ7dOaOyl3Oc/HnHd4qKm6Qfb
kqjZNUGoiDFUvtYHm5lRXKLtiZeaaHttH8Rsx+qtwygJC6Lv7r2KNVvuL5pl
4S8GE5PlrAWioNd/ubstx6nlIDIRw8/PwBxDDdlJ83IACH/xuzAS6ZN2iHAr
4SwIwgAJN+3jQcco1Bkz1LO7NDMtNHgUgqnmL271Xel5E6ai8SuZZ4lNppGR
NJCFs73QmLMSSZ5jr21xnXAOBjgJISNqp1InpoVdFd30+EulYOjZPT4zDz87
MBv6lCKvqvYG4htea9bEND0oH4Qiti5SVNwvebdWj96HoE+/z1faw5g0Acbp
x0j/hA71r4T5pxtqWdpCsjUMaJotW9ti0OZVRFsHbxajK1xxkt3Zw2YQLWQG
iI6y9EWlqAOOVej44P56IF+c/zKLiJDC6N0I4sqW1014YERS9QB4z06JLcHa
WQDFEHE1s6/DrUsc31x/oc5X/DL/cFSLoF9iYWfRirEJ2Lou7mgD9Ptgu7nH
ejgkf9QuOaolPKh39R7VgNbUJil8SEFAatmkWHiMnX6BgL4UUs8RasBY9XW2
GsOjUN2Ss2EsNxx7vNfkzgR4IDi4zRHX/hXmfhoWVay6IN7blNzh1MwTmQEO
PpaFINlimVaIU8uyz0h+Jy+TwG3O//wZjFhGv57fnDgc0JM6yS2Bo9b0msKx
WKgC6wZRtUWdBM7EyxCD1QUB0sNJOAJSqUuOHx4OoHkfLIMj03PeAyo+FXyR
VWawrCpLgG9AJ2se53QtseMhythQRQU8Ra7PaNE0qMdQ7ciJsEXy+xNONBnL
app100S2jyXWyLlJyayY7lVcCyAKdODsfg4i//Fw/4oV0QTcekfcC0yS19ck
FbV7ZNhwymyi7k9SZFZ7v72gyIw8ZAAlDgmqJSjKwD0Sj7t3PI0fD7OOYa1y
CAAAqt6hdbYpMpsfIjE2LR+9xTp7eR4dMuMsgI4lepCdfoTiHQMFjJcjkRr4
GFlWcHndjf8v/FOWAt8kgG8NUo95DcoKzNdKhR4K5pwPCc9jfY7yHJL653Sd
u8X4bhxPJFGaQkpylIRxlxmNB4swOF9Fswl7CYdAid5J+QOowoO+DTjmi05+
g0aYyUky6trti1bXoINKtV4QHUD0TxRF9cq3nE4ovBe+IUtbgW2JcHIswbCQ
Y6Sh+njGE+oGvXx22KhUUm67PFG8lNvBN1lmYabsqnUHvup2CBmTCrZdgKfa
fUatEBLJq8x3iCZcPwajXWEyGxTOOrbB4gyqmSImNgpglpcs++NWMr/VfQrr
yLQpNNLPA38E91k2+IRxkEEcpQ5ySmK4rYGJN3RUmNw0rnFZDFUP7JJPQ1XF
3JigG6przTszuj+Sk/ZwXchOWVlycuhyY5Wx3AwIpRksZeWN09CVlFORS1Ch
rL3Ib/Ft8FYihZDmSkdZKqhZLSboWqkbQ1xtxg2AkVldfBxroDtIYvZnbYw3
OugwmpuHYwqIf/296p5h0qA4WnHkIDxgSnrHUduoSvFG888CFlnkcMLuePZQ
0apFwS6fQGKTL7FB9cJ7P8MRah5wpLJN7gJbHhnhggco+kum3jkTdIKrJAf1
9NMeX2NAeUlJ1icSVxlIFhzi/XZurRbVTOVnAILoNuvfYGhm3jzizbW8G1SH
5V5cwcstrz0DRgQPUkhydU55QtE82sDttNcNLgfz4mvEXRh97YAc/6T8Gq81
ND+wMmxRvdbvd/XIgTz7kN0nzCe1wYfryuQOfOp4MroVpm9Yec2vUHWSZwE6
kBw6n7+DFALqJk8uuZDjYXe9KiZuHF+z+scm8/N8PBu9ZnNBFrJTaDKjHLXZ
6Kco0m9yQBX8egnTyfSjPtqK17i3bQioj0XkAF55+/kiWgtK/OtU3c75ma4Z
TXNnvkbpzY9P5gSOpap17kpmFvHB6DMmE7U2uvLKFGJMTRzamxyIJ7GSw1dd
eCWInjfQ6ypAcZv/d/X0lq0TS+yk7lKSkBvlWm13asvMjKMLyL+TGlr9Oi53
SI8tVNbiSfeZIcJ8hU+F7lodz0cGyLFF+ukJgoQqjeLIVaan5gWS6jnDunFG
6dE/FlhHeQChn0RV2JUpsPCM9ZTxW2SIm6cvMdUH1dZqf8znf2G2LzNG/mjG
aS5iATNG0HsNle4EkkphHAiMLREVky1iBaRHpVCWkAAMCwCtS1tQp8Cyiy74
dWw/gqFV4qdNljn33m4+b2DAkQnLjFntBgYsC0tDkwPBHinaruiG567GV2r4
+PCwGaRVVmPiok0FIJjdu5qKrKRhT4K7Q+0+osgZG5Fe1DSG/1sZnEMHXPi8
9snftvAJbeWrY8V+VLq3rSBggXlqowQ5A6jKmcJixrnXPS5gV4qKZEMA1MWP
3k5S6dnx2Ezk5hdYCQiLDsPw4a5Ab5Bf0tEm1zdBH1+rVKy7wQ6aimckQneh
r7yucVkEeTtZ48et9kWcFn8St8PdUpkLNzqCS+QgSBm/9N2nfEwqjYPNeP55
AFeGbWJ4x8jerrlefMYEsSC/m50wTX0fW1AiGq5vcOnaoRoXFL7Iq7R8y7cn
lMSL4rFxnWts3afojrQeok+rSjmOfJWUuahU9uZAN7UprbC2nD3rFruiaEF5
rg7q6RJ8f+IPpjptZWJ+7xoG3vi+dW6aRgFz0yUwjFgmoVYTcZVxK0reodOM
WlRX1DQVULVxych3UYFBFjM+kxvdMPjnb1GbwK5wivRpw0yxoJQ4lr6UH/or
9eqXD4738Z3bhn7hH3oiDfUXATosj8YSjBy6GNHs2eYs4ELynHOGf1yyzJNk
mq7TrMQY7RZKp5PUhsgRZz2TuB1nRmlqdlDAshYDOBHF0E14oRuiI/NNbRpL
3hbGG7towBygpP21ZMd+pcdOAVTMLm3q3G1FknVhxd5ftIy0hM4/bbNK3zYC
8RNbaVHBEvhFypN/o1J8/QSpA0jZ8PwC2L3O53s+EOfcyFpS870nZsZvylmj
rNzo0DcWq0+NV0opylcSi8ZY6DlB4YepFayNlDa7TmIEq6fU60b7FK672s0k
L0Tow73tC1WQa3DITnnZGfp1dbTzXAImyR9H6YR2NXveucCXpBnEFDCc3B0S
Gr1HpZjPfQz9HL0QUyF7PdxjYyOBY1h/pevVTP35ntbBsgjWw7SkL6mQcxjA
PreVOVyzdFc/bQvbgG0ZFBR2zD2AzzoTK86bYwZz+kSgjQvWSd4quctGpkv3
Xe+WeoNuRtOLNflOsxqHerO8+BG9H7PQfPv1BpLjzWSVEICv2qMM1IQ2lslp
EOGhXrbgabMVaN+T6F4Cje/U6/3o5NdsuvpPW87jIFkkjdhfLFwLSkw/0GdO
Iivg/FOeKnr1vJfDDLnIRgnzjXJ3MlGz5cKBXPQS7cXqn+/wIo7jeGn3caEl
G0R2/Vv0XdTuIh51tWs43t4qN0QVHTSpewLRfOf+qjqwtLLv5vWZrsEZNK5X
hEujB9cu/06smlsLz5r2PuICJrESGb6pkHaUb4R7aQbRBXbLG2iIGZHizb3k
YlK1J1K4UItOq7s9L2lAR28lu/4VTnuh8DCtVgjuwJ2AZNdRyKGcCUHx8EAD
Mw/iWUmc+o+LPsK1n6K1ZTfDc8OBqLs/depxQ5eOuXL2VzFAae3uVFTPFGl+
+IUBIfksw0yczBxUuXckEeHD/Ftb4Hjj47GBk9RjHaZQKz8YThqAB/XfOZ6E
sDVOpT/bEbOuLChK0L2rn6A/zf0vhbjgRD/AC4MGcwRbDXRXBlb1bjP5cVXV
fUu3bDY+aMJBcDADe49j8vdP6/56hu8E/xhNccQvmdIxs79R7atVccpXdubr
2VpynqDNQ507ty0Nb5xQP2CCFcIg6pTYXb9RP/qY0Fprcmg03K8hHrpC8KuI
xMPo8RiiJT2ZQ8oO7XTIDMtcv8GHH7waiygmSVBJeho+ht2zU14E/roroTpy
2js0BifqvOpNGVAuLKqmmml2MJ4k8hmGy0TNSVHQuQZYTO1spgz0vVoSuyVA
pEesIOrip1tRQrjzjgx5ts+q3PQMAFs6MdLIlcQTHFJ18Q4YmYMkqGSZlZi6
NgXtuiXj3iDuwn/zaP0OlMK1dqNNl4FIZmxuVCXihkZ9cvhtFSK4l3622+ZZ
xKXiLwGjXZt96sWN2S8i/KBOsa8Y7YgA0tzA6BmbNxC5foQF/bd55NAUziC1
xH8FILtEt4iCcf1ZBwRWD1t7iGJhNePptUqjHRFHAiNpjIm7WALhnovHiuUQ
pfFdLZEnuS5zuaTnTIA0c/TxI1rMPufqhPmtg/ZT0vywhOs+Eyy4W/kZs8hY
1iZUKHf3tOT+v85wOfnu7YJPm8Z2CG7FNYlzJmQEZSCRyxDxqituKOmw0OEc
M1e9MYPsQ94jfRrUwnkp2SbfSg3o9KJylNQYayh/iloNJbgLTy/sYAWnNt84
ktkC85UJ5HUPcOj62+3gq0NlzeNhNsxsNkysfJMbTQrHrOT75L6d0HFFu1ML
dMCTAgeD6M4zvCo3hz9y5T50F1RhkVd+v5J79CCsjja1QeFSq72hjpyfNfWm
KMuAMbCaPZ8+L4S4eqX+5jF5A5yBwXKvU9DM2Z9q6+7YfM9PXOokkA/NaBp6
SA4WYjid7vbaKggOl+laXa/V8cRRKGC7WkAyQgEzFL8Q21nXhczZIXAfFFa6
tNqYiaI/+xKpK2SIVW7/SlGcU4/eLQGmt1OhSn6VqX3Xide/Xtkj1XqQyKP4
JOYhM6cWQY6jPNlnyl8MkoGvsqDIUk72JV1UfvH85ORLwxUkgjsPShRoID0y
joo+h8lUGBggEYmuwtThSoo7udNfFSXhynj7Eqki7uMXeB742z4sjRkLhmTY
9+35HWitssnPlYxv5Ys48Nejdw/e7kIqppFWVLg9d1jw/j7nqnxskk34iau9
V89F9FT8w2wzrVcy+tsHvgbBFIB5UY6YovuoeKOTvfNiI9TZm2mo6ELZ5pUU
mgKxc7REWA8wWmtw7xjkIvKzBP+g49MKTWwd/ClRNc72n0Ge7eDi4pPpu/hP
OX7ovlmZP6pbgZUSHqv/b5kDIcUHgyuPlQjNjyDOmKUSCcjmwlwgBOaJpKdr
aEuX/kwr1A9hoO+kRg1pmAfMI+ShK0RLu+4OHiSzUQYnTYdr2At7PU0Ch8A+
P72W6kPtuoUFmBqhBqUBLc7o3e5Zd2C/93OqSY3pvF5f3H++Y1C9wBVJjjxO
rb6J2cLa9Rmg7zwSyXXQs9qtH6TCWzHAmzcBjrbaoDx8irlv+GdBz/v5YHQ7
1wY/G6YCCW/FmkBeYAILuqvgo52Z5TxN75MB0X7vVNkQXGuUWM5Y+z3hdwUB
b2vTzX8TjyVT06U8DcaPY8gJIwokx2k9jWjSKobS2yuWrzpG+wXtaMoGlI4N
zT235jUcve4a//qrc8C3pwlADJoiHLkVkZRsvnhF7C3gI/e9BT+Jgw6mj6/V
Rv04v+nGHFaX7S3PXfFaADeG3V7SjQqgPQmyYTxa30FbsW3JJboJrfwn26ar
OnWFYn9Sh3fyn7dX0n8nOUu2PejzWtPXbBat/5nmi2pVk0UG1UdXC0F00D+T
hCfN3P+lEpkt0Yy41I9ViinbdoEc75TgGbMy0MsIy4U5/V4y2ihWRNuN+Jm2
WquxxzwhJqlkkeytdRD7lh0BC6j4qKG8At8Cnshys3nt7GsdbVMYZe1PEmUI
zgUdbXiB8h6FZZdqRpiv/wAQNwId5Cxfm5rByjFYrysSjla0h7rL5bJ4AD6b
JUlPNgvj05YBAcoNKdudISqxBpHyASGL+rDWJ0XFQWd8uSPi+LmxG+fzj7ma
nLTERxx3fRieLdMUf7rSunmDsd3ql2YgjVkM+D9Kl3iZL9m+HSCx7xRq0II8
gIxxf2mNRn+pGnPVHDP+Rj/RKJnz30gb+v63n8yKOO2aYQL6TROZ4vbqCSNH
6k8YpCuUaBj/gYd/CE2233LuCQp9YYoPb5MKj51rY95dkK05L2TU0Dy1PZRm
4tWEyvH//2BLuz/8qy9b5DG2vNbBDwjTC8vYVlE1K08kcUavuBwaGnJaVwFI
VIu6yPmYQWFDr4G6yho6nBO6A7vHwHn9UGlu1pW3tn5INNvJZmQxjahw1abn
CR1sTUsF/qPk62mdJA1vj8AZXh52MZcbTND0B6KcYcQvjkqIC9yxsrEdMXqe
Qs4yEc5Qc3GQbfpqOP0EwRj1Ll70XIRFLJ1S+f6phbCSCDA8fh4+Seb4/gGY
F/p+a+IX+FbCRGk49vd7iLZAQpWhpw/Bqh6TN7809BSDyqN/PKrBW38yVH5b
Q34mK2z33zH7sS3CXdZjNgIZjFpppi/2oifewsomBjetafE8vaXesRgDX3Zy
WOV82hkHeFPfXi4O+y5HLuYsDyXlLc6vfidyLKxAf3snqpkAMjqgqNIIm/8b
LBTK+s119oNoE5WOahXgLm7cNyVqJj4gNV0LP3Yje0K5WMOJfbD0ryCGcJRq
re58ziNkfRrk6cbwDbtZCPdSQ5adaPh/g2qu/2rJtVkEscGbZmvEN781qRSW
K3H5T03YCTOvNnrJAtLnfq2qqxsJArm2VLIfloqCK1O6awGJtCz0JCFFywPU
ZMbYQDGkFVu36H4whUm6FbK45tlfGONSYT8d1hRbpw0QRgWHlFxVVdb4Fv5V
oIbUdSnZfw8CjxB/Mka+pdKY5DNYiupVBl+HOzzd+M+K7nVXTWr0XrBP5xTC
2nbLJPi9Au0+NPtouvEKB9Zo1STmwzTtNp58ukB1wpnCLqqY85lcpbSo9hQL
IrpCPcUbwnUsg/cub/vfVCp6vDylLQ5Pm2I8SfSig9Dllqjd9rANHfJj/QU9
R9o7qxL+qes44avUjW6JJcV2CryOQDgPG8ROzfVp2E3VoTwlrJDMdG4CN5kN
qTped0waJqAqXQZrahbzY5xnQVXwaqAVKh5msc77A1oxn9dN6rWSnuDjX4cw
yPfOORhGrk+WCiZ/Y9QeS7Pb0ncRtgT6yQn0buJYBkBL3d/iUM07AbvAX+or
wmbhCfRgaxo0Gx1uYaB0c+hbsvqFL9DjEt+XcA2Hw5BVp0FtL2Rj0LE4k5oh
KAAf6QPgjUV810pjB8p5H2fm+/mJ31uhePoskiT2tIFpy4C5uYIuSAw6I0vQ
vcn3xKsuyhz8MGndjD5wR9AAebbqjMHDOZjgNBXpHpB7S9TQQqI6zGOsXwPF
8NdxO0vZqdew0S2pXhvhKyew2nCdRSkst5eUxEiljvGWE21qlTV8ACku06I3
cBUVwTOZZsHVfRcB/K/M6xGbn1BJDtWZJlJR4FncbNbp9afyScU/OkGdlSi5
eAP5KcV7oAlj/Yuy2eZ5zcrRTsKyiSJlp/Rm0a4cZjggaTIW/jrzMabxjmgw
eJWrGz9yOOr99K/J9qCK8Uj4tuRIz1mZbBFL3bmr7T9B8qY87+VHaft4GGJv
CuuYwJzCTKxUe9JfANlbM5oOoP2r8DwGteNxTxLWYaQRHrEfv/Dkc5ei4TJ9
wf4I6vPK/4pFmqtfoOXwborAyLDcZdeFJN9YaEtJUroXYW6d6mOUks/7U6oj
0G+AHw9HJjUnoPICCcRIOaHhg757DvY06L305ES5cml0UIiWPRW6FhXRRqtO
CNg6EZbvqOEMKqnvSOgmoJKFCtihkehh+aQZTDoStJ8qNmk+DNrRuhunJknk
utm/BVcerPsdjyFJngpYfVWrd/SkhNdQ8GWw4F2Ohfo2w4AIwh1EGJ0kevcI
cXPEH3ZCK5n4WUerRjrvBkwqXL9Kv+lqoH2E7FtIEsgE/oH13edgeREfmDTY
B8D6E3x2mh6TT0tTJtjgmLoQqx6H1tAXnxKB81pyWEjOSfl/BwbDlkiuMgXE
PqV+ohb/wncq/VcXrLwLenZ7KO0wHJmzG9ScA/IPq/A4IAG+7nSoXVZ5xgdz
5DsE9/CC1s0PBOKSrx7RU4ug0QcsH9GvN/7eOM/CP6OKIexBRswWZ0O1qcfj
FyUW/UT6LySqIulqJwkVrmDVTUKgkOpIs+D2JGoaBQVgJBF/b0+jlCMnuUaO
FCluA1SL9bNaIEWd0RhZLXNEAByi4ZUJp+JETBYO+77TJQhOSdJgWFTmXq0u
bNwBTBTEkRoJKVNf7a4/HEU1JbfQ+6RQqDqDs1DE6gxB+iJrRCW8PWfJonvU
Sei9+vwvuYkeQ5Ik45qNeDR2Z16TYsK7Axkjtb7F2rZW1ix+QQSw/6cJ0Xiq
ooI2FYmqcpTsZkqvcK46/3+0a7YAudUP20u42+FB/s8WhGPBx877DT28Uq8P
4vK0B6c+bE5usqyb0T7CFrlbVDudRgLMNdWXaDB9iBymrgMrx2Jg6qV/a0Qy
OChAeOXxWee+uyJXPLnpx/OmLnkuNu//ZYIhm/8gNFYFzdW55D5oo26pclWG
u89RibFSW1BVLl/NuaQbKUlp/PA6+2F1JzfFrA79hr/KSJZfrUYymM4KTYf4
rZygZ0K3jwUS/Fmm0txcBla0Gt8Ah6JOOa+uz5QgjehdPvBm7F+LJdER/7//
MA1atos5aJhzrYDrY+lxm3zp1w+nUpPOq21UE+DDqv6JKAqxlnBLcp3l2f+r
DBf6WNONVSFLIibHztlmOJi+aH4Bzi/hY1qAm1GXFBe0C4vLaUOIM5bkdOkA
hXaYE2KoVOYbmRdc/KbllAKe9ukRWhIzKgDSebDb5TKOiJCTh5+JwMHQJkY5
B9IY486Ibk/42fhtaeqSAT2ZxmUZJjQIgLKEX+OzPkaHz1KglIsmX3EtRPWp
e9MjkWlO1qXo6UTBdB/JkD+gQOoTJP9ZY0yqcxlXj+rL5RPmluiFPbv5y4L1
JbVJAouIuTvnqIKEYYfsmEONp1ajkysdSnOZz/f+VKq+Hf79eU7t/xvyY3lD
Tz3YnwYmEwdL7Pd6rMvchQo8Ka9wQv8VjctcdH2TLEiTYXAsTVqD0VRlvW3e
2lZ5C4z0ZmWSxHg+rdqdYMnmQBa1tTp8is09m6CWBBKJc45+Jh4sgIe6TOlp
BV8IRue79tcnntpNuog/kDFiE2FRq1cDNRtorNzLjFpUV3xjNoVvcBRnNDZr
6eKqhf0/6JIaWEiF9eFdAHnnQoD3VL+lbceRr8034bvrkEz6N9HO+sEyLjWG
TK151WJBRSEKbU8rqrS10VPX7tUw2Uw/+04TikS4PVUcz6BVyMqWWVRXDjML
3xpxy91hVD+BpK8VcGRL87yo3U2gMnNvhW1YPEO3p1bLpQygPypqxl/Cdei2
oR0uftBX+Px9pOhbEnUrGGY2YhIn87vLXxSk8tJXmaeUl6Mxmskaq8aF7HyH
9WR5EMr5Ea+51OZ02aitrJHogfr5FsTy4+VNPeMzPcskgsUGyhwOPIuCKJtu
xWTRv9epjUvCrHbeYyamWR2cK7rpyEdmAtsmKeSLkL9L7SGKR/QeX2gzXpEv
UjCBE7TEfdQgREmfeWVtxmCHGJGivRc0mIkz3D7yYGezEtV9E3fD58lrzmmG
/RGInYXK9ifD2/mbC5gTQBgEM5LS+b0Qv98aVKgn9uESWcV+wwzpULq5BgXK
sGsEg3/5ewM8rlrEFA4YTz91fr5jCuLg5hjBGiF9ZzNErMBDl61OwYRwPvsQ
aqxtUaooYXlj9DXALWlPa3DHjYFDJ6cBE8Vjjz8fdJtpo2HDFCltsWGZ4YtD
KCoAcVzRzV2/BIHcwbZLjo9TW69tpjzRlDLvn6NxcKEWav+1/H16PcvpY80L
oaAJ8uINicGVCRLxd5MXsFzu/jaWrpHzIz8VqEhsWMcxpEdRpefIO1EhQKNq
SkyT0hbhCLlEDj/8qYu9HJMSvjCYDs+VmzN+vXE9RkDepa6J1AyU1lfwFwcG
jjYpBUpateI7BQ64uA9/rO2SWt34tTy5xmWxNf/AKqoS8ceaKPXmd7MXRX3Z
yI1m8aPHHGEQSqfVHrKjJUjQru0N54CCv/fU8HayG4RSrGRoTphysrbsLomv
oLm3T1/ZosKQyqaoRysUQK7m93M7FaK1X9gFjEy7Ey2hdsnoKXGbe1RVtYlf
7XTIsyOzSWUT7JCWd9nBwRzk8KT+SKsBoJGvKtNs1g8frpaywHpCN+K2O8yG
p7YN3OMSfFm01nuHBIFJIrOyiNzvmItxVhyhh/wogEJBHP5UkBITg0RHKpJ+
nxgABWmVHJpPwLA/6NinvnpX+3eeWN0kIIfTfJ+IqDrGN86sJNiCRXSz9J7M
AH/goyjJitY8OGe6qPoUNMB4+YHHInVUOuRioUdDpcDhv/AoyaFAiqXV5oq9
FB41yY7XDdETVSxwrZWdwRnAiS7YDCEFc5mP6dKe5Yj3JfP5QD4RvKneoAdr
R+PqwQpcz4B8tPiOoRga8+9Zlvgv4SrT7cDFv/6tvmtm6qezGz1mpc0U0lrw
dlv3olQlhR2RryssR35EbnT8FoUyz+0XxIR4D/tiibBTZAICN4zn5RvKRp21
mk3obpVuN060I3JXyJE9GxzxJbs1L0sN3W5+pijsR6i0/5yw4E3KeMJNkRLD
uRGRKV8r0e72zmgnmTGr5M4i91BWQETJSeGoLTJZAb4KzAhKzb0N+J9bi+K7
rGlN8pY8KDkz9VLublDyOQzG6AFrK6qDPBEGW6XL87uSxD0LnFNCx7aIi/3y
LQpHvLG/JzZoPpmyJstjnCOMCTt0pLjQUtFTDLRxJgM4IXyYo7f+d6FBc1CG
rMF/mX6KZOhw0ed6q7MqacQ1FOMgVrLDGsStzsPPGiaV31BdIawYnLIv2RYg
LJU5BKkE6PngfKnHm/yY05FkkOR/+0JfFW/3ppV8y2MwpmZFXLW2j1kF+/Di
7DFKz8sBWey7rWbjfTdULI7MkQ6na0uBll5QkWz18I03SL3oRiEtLuvaU94v
xf5uPAihrqrlJxYFm/afr4dJD27ajuwGItw6MNv6uNsu4E+MTg1w8NRdL9NM
mfJNl5NKNw/2yWvB98IfSbXlTvSgFAxHNmjEGgaRlEs3cNk6K2mKnZyhvqrc
vhZqSZDXLcp/2/a7RcB8feljiW6KUjOscVE+Q1HZm3vO5cvTma7/SQ5b3XpN
furTpaYAfgQWWh7oLygODvGcO+GctyycXJ+yw4/ZEXGlnFYB0TDotKjbPZI3
KGzl/gPWxIgHrxMgjfkka0nu5y7EQV3sUhWumkBSeDQt0zA/aZUs9n98tN+n
j81rhyTvLJuM/rIySlYq9kHwGRHDkEEvw6SRz4uEkk2/RgkMVilz0aHDtUZ1
BCqwJIEiK5W9n0uPJoR12OZRsf0tq3Edfdvs32YgOGUwT7fW+vE699pjbRvY
goiB0QM2Xwx/6waxaBKjUp3/dz9m4obcXOdh8Jhq+BHsPiy/K8TtVMvtlSSw
KDBSi0JkFPRbVdcEOm/EvaiXfiUB06XLev2ZObMWvZxgRI57pWvbsQf0m51n
fAY9g70OUcC4c/uzv40WYBQtGhWtJ9e8lYvj4uNtoG3mcbjJwLdiH3cXSTfQ
cC5tihLhuVgTqBRf5Pc/4t7LHk788Wx0bUwQkgkjcbOVV3Yqw5c7SLq/LOBn
prVrFp0XrFmw11iRS1R1ouA23afbHhsVXoJ6MvL/YRXbZf8AIhXhGLVpvqX9
VYJObQXkhYTog/MBodCPE94mykltcgxgQTp4IM1UF8MGHWBfoQ5VsaljB0o4
mF5cWxTyTtWjT/k5kpYoRFwjKgkBUe3DGEKQ+o7H9cwfTxgHJPC4EqRPY1gA
Dx2OrhDMmWhflAUMrYJVgWz5QdKxAvHGUjr/9on96cI00Cptdfhgz+iZoEGi
AwLRncshkLi/J6R3Ug9F+Wo34og0arfu76Q5PxS6yXpdlKpsGZxaI/pkac7P
V9DfunhOerijkiYLXy5PES/yUXbwjKOTihXN9bDJVuELM6IOmpG8UflgsuDZ
Gy2DpVIPsptCqOKvHlyamPvDUEDO8sbA81CVceIgUKq8WL1au8zgWyaObcqW
YXw/OayzL4Bp//cslgdqollxutJU4WlKDWM+0Tl0Biyw87othlRylfBOt+hp
PJ1x3gQZQs+c9HYFvyyZpiC9Gw/bfWuF/tuzcJMifKPjmqyXZeUeUuBcym17
BiqFwE0qAi8wz3hd/PTJf4sqcn7ZN9K6T46HHTHZ4xONrzaX8DMibjeGpac5
S8Mb6Utvh4KQQm8RtDmxmkYWpDk53sYVb2dz7zcTzNgIeZcpVma/lxvF2FbE
88at4e6eYjioeLd2JXdPmTInvoEPBFVpBPBnV1Kq5qw9m7cqCQHIjZuE7IS5
N6avGG1LS9sLAd7Vy1zHsyUyriiyxJVitxDhtHcEE48Txx8s7EwzDnauhPIT
32ekRk0goFUJpnLdD0AwmYCZh8kJud49K/tJKny+lWsCD1dpoV44e65eUFd0
UYo1Cc6KCwCqWz9rbiAjiA1XM8y3BGMQgHELgIGCUjOHmt6iOMIx+ubUW0Wp
S/LnVYLgKfTrYGgtqB0w+FgmItigJ+7gYEQ/BmhWcRp7re87Wayr975ic/E/
XJsjpK9VA1GlcWUXvWiMMtDfbKCkDXFhnh/clnFxiW/6Hf4NnV/RqtPUSAzI
jLsYBn7fCyU8zx58ohz66KxhzraMKHQ7lDGQ6CFVWQl39vIfsKsDrpSS9mcm
CKhxJvpUOcY0XuRU2Moh7FG2TSPBa8haf5PU9pj8WZQL9uMztBgrkreDH1j9
/tgSUmmWJcTlZzR3hGqb8bJinAD+68cOw+QVVbI74JwxKW8ywab+GAMME7TV
HHL3UdVHYHai443Sq+ybNUqsa42G0ecWp4kALbt+OopYMhsRpYrdqnDEvkt9
IiJct1eydeGuzT7sGjZzLlyiA9miRI3bvfpgFn3Pe+gaYslXzmDaUBUUZXKB
EypBo3piLO4lsXACh/PeNzodnpsOaBYlDKcdZXp/+tRSRa08TFrwzAj5dtXO
xsEoQ9PBuuP1rp2LldsxvDV0QMrO3PMARQTYVBl8Xj246FYTZDe/90HcviI+
UdfxjHVFhUpNcpRyaanPRCURRdfOR0mW227NVSBVN1T2p8ZFx1gZO/XBJVhp
OzUQ5BfPmA2xLb4as2CfxmT9p8PxeNx6V688RCuGc96cI//p27ZXOwU0UPif
N0wOoYccP5d73lM/4J1au33aJOhxWvqZ1Yf9YSGotuV7MeAzFdK6yXBRvGTC
8SMCL2fxDoADhXnO0FSsYnpj3ppY2/mUJ+pLSczk8E2GdaPeEb8jBCe5xtyp
s2Sq5kTN3BpeJS6LyoUH1Z/XVyr2p7KYQelCwimivpsciPgSQOmPF4IZIfGN
ytTuPf6DvIzdOKOpd5qK87rUObd+MT+QilTeRA5jv5e3KuSJaljbEGHwx2FR
pvHbDCO8V4wS1DQ6LwyVB3l0oRk3Kfds6NjgdSh91JZlBoZpukn6U0Sokjk7
pIlHe2hUdiHtGoIW3lnaGPlBFGaXTSJd6yMaLdqrC9/KLota7SyfthmvLpnX
AryxbHsFZc6M9n5uf08Ezqo7zJBCxBTYwMPP/oclpaBC4+lNY3ZqkzcHBGfX
5GGKDLMfp9nR8X7ifBcqSqXs9drbMJZYiVmeypYnihBBh7Stnipjiww7Irt6
mUUAv7VlG6phRfjzY4yE43gPUbpsbRYSu/iEcpqg34gVUPC3Yoez4Ca7++h/
KwTcK9b2NfmjJstlCZsvRS9ZiS6mm3+ufqODlHiy6t5vebGyBGMQ57uLEt9j
GmMvNulP/viHVCPww9BqJ2a/Bbz8dtxWfWPW/hzBQf/eSLd9mWiQ5s0evmwU
wUKdxqZhodMUD42QzLilk1ntvc0BtecbW7ndMVYHek4w96SbBqZwugE0E++5
FiulTosiE1kbmS4yo6sTV3HU1JPIwLiOPbwt8BMECOl0Sz7PRLfSlV8oN0Iy
40sKnjER+JK2zFYcrRNnG3I83bK6cB6fF0bUXatNU4VseK+Efi4nT1u26XmM
5isHJEwWim1MnjE2uULTZL+8m9vvmHj372tiZ9iGnlKxcAYYgtSqTAU52aHN
uvsUvM557yv6VSC00bTokU8xsBrQj78jrnVMk013Fn3+pnXlJHgLKWOoS6V+
QJKG+d3mMZlHF/ybLN3LSiZjJTJxv9oVp0d0XrUtsZAYLuUCBCS1kjDkdQln
qf7IHXXUWcP8ubURRlVLwsmgUbRlri1nauvmn/zKD0TgbUepnuQONK+Q93gy
cNj4qlCGP8v5MVjj8YLIGFdawVjpnrqO2c9yHwYH2yAJdgb1ohB9uW5bp/yV
pszqjEki47hT2b8OpjGp6layHFE5/UVgXCP/dl9y4nvN4VvTUM5fw3SlMkJC
HLLUg/7E6Kcl2LZuIxy2sn0RhYxfs5Ukmh8v6zeULekvw4sLkQW0EkKkb5ll
jODl63hX5haIfft1TWfBWEoN6iH/Nxp7L3+b/h5UhCIx4Zg4Kn3VXTZvr+4H
miEKoL+pH5VuderO4tF6Zqt7WwI5yX/NDT0Oa/T7FaXkU1Y8ElppiUAMZfDZ
F7MTNo5i5KnGGhBeDQnj8egA7sxMorUOHdcK62PlJmfv8cc4lehkty4K8Fej
BGRtAG3X9KZZ5KmIYC6zCm9XKafQALqVwECxWjeqnvrCpBhF/n2WsSQ67l1f
UV1tUXggKN7snNPBU/ei3Eaqqi0v047alnMbCIediRBNwuzvPdcW1LyCz5ep
bNLm0O3QZQ4Ohw8y9kGYFLyMbVdGA9aO9PmFEIWA4IFcNpRMWi8ZGg/B1a+q
IGWdkkmuATnI4DzRn5lW8wumdDi5wGaSGt49qoDPmVkH+7DzAgVoK5eKwqQ7
HXVfFMSEVysx3uF4wAQ5IeclUJ2EDTYSQcExcY88MiZ0ZrF7nBpLTiPOp8as
lBsRcE5ZWo6GsrdCunRAZ6571zbNJAJcoNGdICP6nysp+nbsP5io/jp96VC/
HyPqK37iH9cGrAQ9du3kNU+WUjDAzsUUjW7Ak6e1mYb0qZTCKxRjX0ZAwaeL
71iLDgHjRunMNAM1sHbPJBXLXabNzItrLN0ngCm2zq/GL6yvTuub30VzgSyK
nY0vG+IxBjL1/xUlo6L7IXvKnkv++gEo1KJ62rmhs4URGAdoAH1yZJECg7ur
9tziv4Fdr7wxDmiOSAuZdvudlkHlaSU5Ll/3/ssFEzoaTE2R0O8uIdf/gqAf
GUV9dmQs1ex4i79+vMbQVCpEUXqSY7LziXS9UmJ86TefNSZQZfEZtbN0GCTm
1nWkvKfREcqZgM1zAxnd9BcZH9uRJ+Dc95/Q1M2J0H/JIW4nM6lQnqEieCAs
uIabPYvytZmDMeYCVDRXbzNZQfp3/uoVCvMQODsQkvRtqedzGZn8kGRc2pzt
4ZMjNgfSJAkaGIYHC73m4KgVQn8sFw8IDHcCQbFKYn+wYTeJQjvvX+3IEzSb
MXn2jVi0TxRYwiPScvLR6bf3gKfIheAkG4dIcH8uJaQsYucsgOsvma/zQ+gd
8VnACLEBgcmuyDjsfLwaCwb0i8Xrcw9MTg/ew4hZ1S0NI+DpFmcmI5lKJndF
TFCCYaG260mDnKBOF2hgOiyuz48izNnqFOx6GSueaErLSsxpGRomKF9TliOe
NK43w/cURHFLXLogh48XqmE+7Wo5NBb5A0NnSfCJ7AaylSyHE8STnqMBHMv0
DtXXqz5ghDdIuxUmQTyK67td6mUzkIV++MYLfhwpU3z9Atmf4PyBeUW1TofU
i8RU9V3y91MDOZ7VY170vvCGh0aOpJvGTkmNtsCS0UnZIGqNwUcSSiMcvDIq
JsDf5iwz6G/ojSsxYH2cQTtSVljAWFWVp9/Z+Qj/ihiU2RtrT51G3mupkdai
/4ovV1IIrMDcKs1U2+aCbAGLZkXPOf3fpfKKB4lFZBq5amBByAGcvPOHr8xW
HDoEupOiF9ALOnxODxz2701maUH4GcyzmAo99VH0RDZ2wQeS97TqjCH285J8
9HAv7v+byrpjgnLXmGFFI8l5qaCBA/f8ETGq6Nm/iAKEi9LAR8b+P+z+kvkl
CLZhPGdsJymJpRFNPqQLbnbdntrLrosAA26vnRp1UK+VaTDo+Hu17d/se2P5
d6zhawZPVcX926f1V0AAzDaYYQjN2Uyko6Uvv/pAHRNhjl1Q5nDpRkw5RUZX
S8KW1qnu8dt8IwviXp1yO5om7TuJPnY0geM1dfY5go/3bxa5dP8g7QKJmSfQ
s8kxKF5METQuTA8gQsVwytxkJajy9Bqz1dhkI8nD+dG9YxxPGgwiNKRlj37z
wthmFvp166Uc1Ly1yRfNbYcx+ZoXatpR2vhNlE9s+DJL62Czm9qwJt/v/kBr
ZkNKIgDgKcA2UqHzot51xb41V+FwelX4CV8M6bJymjabuTmZg4jt0LlU2E7E
CUEVvyyyp+gQyXO6UVIOT2HHY+sllt1oKAUM1TBn8WzP4ZHYxYqAPsPbr796
pYSHAeUfssFSYLpGH8YF7POmTvjiMLL+80BwAjc4AfVC2NZUVSe0cTPx8jRj
ZXbHkY1JOaJlmkvbhpKrkvke0Ywjl/agaPrUspSDw2QJtJKqqXUWG3qFlfqg
CCHFK/qFpQ2if3LulmvxMdI4yykdoYdBvbjB4RvF/4uLDGaPcjKIYpdILlcx
I+/mlGl6HdSIBWXtz+fq3s+nS9j0As7g5tsc5rnQCXB/y1lTzTmsSo8bsLkM
brml9L/WO6v1MzMxDO3vOoARVcoQ6Br2MBqN/XTEXSocbkt9lMgdCleXIEFt
RwE5kzPzzCC79sGexCd855wZZ7Dx5TAnE23n82L0o9kfeZIdgKukW5Ukkqkh
TILOW13dEqgv+SHSc9jfSlsxuJeW42rPj4nuatN1BsIPrIbyjicc1NUmbN59
cQy3gTnuYe/0/xIG/qwRl3X+rfIPv2c91RtG7Fc5XBYsswN+YL/OesurRnrl
e7b48BNlC42eNUh6ZZC27an/d/E+h6X5Vx/d/U/xP9N0cTip4Xf2AZ0SVXgg
IMr4gpTGu0GSYZI8rFZL5N2bn27zG/z4DY0qNCkMlgV3CAJGZUVARC8iQiJR
RtgEnQ/CnYf08aIgTcWN4vnDIjtJB/7n7PO7grMneErOemXfbKFXmjZm1N+U
df0hZRdjgVWjhmYWnFi2gPfO/8g/jImd6Mwv0GPyLgpRnzJXuWthZRV2IduQ
vPLGOw9M0nuelowqP+RYCLyDngoDRKJqqEJKAtv+W2se/4JkT949QvEJSUuW
c1uYo/kLHk8/I9WtqFmsvbTptEyJCVfl9TF301+08Th9oFa95qyPP++Dao/Y
QhaX9lMwFFbsrSHj8kNyqGPjfIKuJ2xrtMlkwDhcj/Gver8Q8HBONVIpnh/i
JsweguknDFZGQTOchd0AeB/Wgmz8jieCx8txE4g4Hs8nTdL0rDBvjS1DdW6h
FP+Lw3QWPKCc5SCVbRLk4iGkdaURRvFDdyi8jKpib78zKt3sUPky8U3vYwey
PVQNznqU/N1yQIFPK4Jwyohb0W0ZENd2f3FbPhKDWx6ug4HA15968L5PCndx
1R9df9FqdUCKYg1moxUmJ5fXOTi2hbILzWsPaPAuafuMlNd8/pu/q3zky6Dq
Hwrwdx4VZiwVxbhzv0IeosF+Ske1VeVFVyqac7WKGRxH7xKvc/rNOPw1LRVi
u2Tv8rlPqN0N9eWx8F8wmrE4OxOyi8IXsRPJJnobWku4wlJKMX3g9MNuS4dx
YOZNDqrCciWXm33noOa23G5KBpclDZyqAKtlbwAyVKI57i7WADxww2AEjpKt
udUCgKKH5QHaVfvgfhihjfvahH7eHd98jmtesXXgP3fs1sJzW8iqy5Mxaiw6
I6JaL9vrFM9uhQoCGld0LlsniTg/5E2eyhv9HwN48M0fG6QsMZcYb4MRdUpy
LOhgULlPtNKoYovuShnBycKEvoLWEw3Rnk+P3YVA9BmsoFhw8m4n9k+ZhcBh
cxN5MESS4LLDDKj3nq004seAeT5xHyxQ+aQTPo+TGnBHcmvHQdGmrRJnSTV6
aIr2ad9eVtUT2AsaLAgEUwyAUetO4KfP1jdHT71DZzWP8dwLPFcAfRmOoYBo
aKuuGlG4Ece86Upa1mLmNDxhbJLlF5qkC+TbgRVGIwC0oNBbuDuMoLk2saNt
0SMN0PNzoBLXGloDfDV2c9aSeL3BRHyboXNKcIkMBsJUfXKTOd/IqSJSMtZL
YSlNgMbOm+xy7xVWgiHz192BRj8u370qZ1TVXGotZStOgjlJ/wVZXoYYCFg/
Ax++cg79nNCcmccHREfBDNCUGBcVfp2aBOpA/y6xmmjC9zB57yDDzrpn0RUo
ClffAxL0ijcl5+yTYtsqzTEjXorzztYGrdLvkQyZMevD5gQuRlWcdSt9UCJk
qdGQXOF14S8BQ56dkOOGrp7kcVOqM8R4woK4hrsYVImPOoLjIyKe6MQ3cQrC
ZmQw9V5/ief+Io1XUytTFi8bUjU4i1+xXCKm3Vb2TzZqcM3CLtXsyjobWYrp
VogXlCI0azfrc3RMuNbhs0sauiTZH4aGezVm7/n4OiIeQAp3Ncb/erHthYpU
HT7V324FZOOaxX1pR5l3f+yPh0GoiHbwBk9X2GkJ20k0FvHpvCm8FdOmSRnZ
JP52IOsMhb+xtl+fNituNoQaZP0PoOYfW7IhlWZUDpXB/Z+JGPauZwfVGjt+
GFRFkW3lR42XDDf43fBicT5CFGEskr1y54WICs4jgFQFcZOZgxYMl4NYzYl3
bQeyXcvZ/qIrR/YU+A4ECQq5pNPutF76/nAJhhaY5tA6dmNpivrP4gku1QAb
dGsik9VLVNjpc60TMb/tQX1Lmdsbz0LBT/2Kobh6bRf9FwO0UVg5U4nnMMyW
8fm3L1VxwOyOe6QIJPnCUdLEHm+y8oNYVKT7oNSE7oogZ1NmZTlQKSYljj67
86xDL71Arhha8/ehvjvY06S1eVSTOP+S2r6IjbtFXhny+29T3o+Y0ZnKTFWw
gBTd2+bfydkqUC5hEtPb74kqeU/5DWChiGIlbTa6cfE3ltkHrP+YsIzdpoCi
8glkilo8PPRAegNT0SQRusSVu7iK+ix6v9hj6EYROFUJzwVgpV2Dcsno/jDW
shhWlnya64zVhmVrFpu7VwEpOenhhEI4EEEz75aQPdvFYhZuOGK9LX49+uNU
AMEvK5hVGtCVJBvi3uopOD1NTGPD5fQr2iZBwDreoXa/VmOz9isXLHtH50Dl
Ogg1Y5AvNH3obpA9hPpNDPW5xvw8KmDcqvuY/UW9JK5q3WkORaUAdCd6Ngj4
C5qZQkEfYMZtz5NfcIMqWPovqKKCZEPwYLQGO0kzqoy/U1rS6kIzbqiYl2Jm
orXz5XZG56JTt79Dsdm/xvxcsPYKquNxzX0Fya/v5R33PmbGkrBgtFUQfsgn
TkgSmNUw4lsTbttH57t/NjrFDJEj/eLAQ9eo0CJsBT0BKmB/b614V08SZyUp
z3kFzAdFNd1ZYib8MEfCgS8RlGr/oF/lQPBGEQQJy4S86tHMyRUm+2mwq2jL
iR7bqKZQEj1kSPLnqL9wUSBg/KzuY3phoCrIHQLgqngpjueeHoWcvxd7hQZG
yagzyhFkJmMUoLkcWEOXVmQzGI6f2lgwPqcWVsssWsVMtHuLbl2Ca669Q9Ie
WwnipHyOjH0sJCPjYH+gc3ReXbI64Wck3rs0LOMDZk67BrhN5kLsC9sWHQB7
X613U2lWBjv/PnLKxbsbP7DC8VlL2SPW96NIQBCv7/iI+y+sY/G/++39J3iF
l2vwomLM3oVazP1qWVrXDNJyP42cfLharg5IHn2KESWimunBCedJGDs6ozri
ZjYY2gHJftr46cIx4nJVeatoEYAfYhqiXP0zYtN5jaoyI4mrhsMrDtTxelmG
2yBH5FsG9ZWeM6l7eExIYkGhdLrLQ3Mtrn6ttQSi9Tlr9H9oUPqaOQVhesoW
gvcnhO7iSZ1AvlbTMSPcJ6skYD/DGey5VsoUgVJ4uCIV7jz2wxuXiT/XEKnk
gYzLuErmdmFKu7wqfUsb0GJYd6SJbH6eQt5we96MZTNJtcDybbn0N+U+W/hj
Ou1cJgenwtdZzOtIDMeC7zw4yip8Dg6IR8yRnecAAp+YyIJMXK162FumnoBi
Zx1vdiO/tmsZebeftDZyRg+Ri8F3k7ZEufQW2yCGnq9XQGeMUOLCtitxDf2r
BlI01pQgIrf3ZwDmREA7uPD0WKMTXd7XaEHwVZyLEB4t1tUgOR2ncsc/3zkU
g8B/WzUggqD7tLI3TSJFcR8wUFKojHLj+dCQG69YdiVwfCBsEwE3RAXt53Qx
TC4xMmbyf5WbleHZJ7+Az/PKuOmyupUPOohefQ/tICVaIB7qpTWwpBS5qpDe
vvuZJTZ2AnrCGwDPpBGtTcBJ++wk/zT3E0AbrB5B+F8auF0DqrUe+JX/3SHl
zdRwqcuQz9P6LKBWc5EciCFGDD+5hIfwvyA92SPjRWF3/JR0qNotbhIcuNYR
6YneTuF3izZl8tNzq8+KRrCxCAPVdic9GHez//2n6bj+UADzcGPwp0iaWfxK
Pqo1YxDzN334kmdsI+Fl4/tIr79JMswFEeqXr+h0sTFHSZboou4ql/+I8uO7
uLn3UI/7KcbnkZ9dqcN3cwctKSXHjxwdiZ5VLg2Ay0BF3lf7cAveetlRsJav
npuJHti0/qChkfgjLjYesMlBPPuvyZeVJYFstwHKC5S/bFBwXA31v/rUHReT
FXKDHImxtSMpCKpqa2GWNrRs61ttydobYY1VU9Hld/76t7nf7m5mLrSKftK6
tsyydKiuPj6MTslxN8pOylKDGtAnAWx7BYun9/odsl3NsEPJeYeCF6q0JGsv
7N9DIYf8sO+y8hSbTT01cLOrU8KGguJYSuUWQHtmegOpciVwYa4mVxhw31MP
Gyf1RKkpSn1muuFdORFtq9LPGRlMlLfwtpAp91rizEIUC3ZEWiwB/Sa3dmX1
w2EU56gYhQAuh8CxPfkX69W0MQZ7xygzMNsdf1oUIzPIw0jlVDHVo93qgmUC
HjtDaSQOcUhxj4qVtvbFr+5dRVEtgUwrUb69vdM921iimbAiXUZwwJbB2gok
noEyAk1aTxL0J6h+OCX+q5g1qz65oZgeHrVum4ri+xV/FZveFo3oQuXz9e7f
rStuM3NhdAyWSw5zbMaJlcfPu9nTq2DDNepeqxvVbrkWavkIO1brJT7mEDiX
dGUVbFiofUOmebcjgrmm3yB2VUgXP3E4Q+6tSIpO9Cytz6Z7aWJYlrlU4yg1
lWg+RZiKNOXH4JRlUysWSSohJlTxx0TxXGqgnKMtoWennouFydHEC+dMCP6y
7dvXFl3JRrEvf+FODThj8d4eGQP6DPjB28YfCn6x8VsVUz0yUQf+haFSc4n3
I+AKnUAn3isF0dDAnPHktuYuJ48mfEMafwxmYt/4rUSU6VuWZ6sjYfPrriVe
H+Rx6uRS9qNCQR45zCvgeLt87TbTkBuS1qTSeLK7pbqqAKtDrtXTfO7yiDJq
G6gkQjRlK7V6fIwyvL0FXSH0cfKlrUBftWC652n1XjIKlvc2OvWmDtqsg5zq
afdUTmO0RfJRcZkEQsMr0aOa/vEH9r4Ld9w7fPn40MmQ3ebTi5YEXDeusOL+
1XB8+1lw8eL1TeA9rhAmoUJfnGbZ8baVKym7Q2oCaqOpHjDgMqpjxnuRhOrE
DUBnsyUEVZJBilQj+2FxO7MwUONxLfTLo4jRhMRk8fx38DP+6YkyTRkjoFcB
HvafZF1hh3bC68QVW7ivlCWIUEGp3wtau8tjiCV7+0Q9HMIJg1zULyV0qboT
ARogT1d5mqMvC3uezh3yxlzt5RdyMioopid2Z/33zHCN6BXrsA8stjrrHZhm
h5zrHCTm+L0lNPFzSjt/i9h72GdaalfSgxmWTmIvX2Yk6OUMfxqvdiggWYFI
2GldYU3LT5q0GdO3SvPJvlnbmpSjsl3bExUyJG3SEXQDqCLOdwNTkQxZFklL
tWHcsRof4w+YG92M02Igquh1lU8rl5i5fNT9VI7fan/6Lyed0ph1Vpp4vr0F
5xVCJVUQVsHWL94uktsa77olWBPcd8VLWMczu767oZRwc2mzgCW+h3ANQ85/
45yJK3gT91WUZNDT3cNMzSfyJBm03rTS1DUHVtzLcZHTrb8A6K/Lq2VSwZYT
DoS7nYzGBM0bDcbcOz751fjl3vJURU4Yn7yOsVnmte2fXow4+NELDTRtz4de
N95uBTosZP9bVrXfoXB05Um6fFjg20H/4UoufSug7ilL8kskXgNqhslfxyki
bNbU8Y8AXEl/JOj9UrdFbFv97m+OaP1u5BeXq7fATbL93eIqcMue2LQTBjJa
baN6tcjbbe/IrJbl2pgphstnHPpYeC99C5OorHrg4YmhoGWpgemD5ZzCKJXW
6yVqvjiurwLdFZHwJK7nN1GQ7EIcDO3Mrh5GdIvGQqPn75VZnAtx9QAHiH1u
LmRsKtphnqcAUL6Xv2gNPbegMQK7vsA3T92da36f4kcpKqA1Ao4oXqQ/jF1a
Aak7TiH6yrB78MRM/7iUbKe5ZCshZwCmif2wAFEY+hCVbpARRGA0BiQ0sCGn
pPa3KU4BNSON8Wp5epzp3N9FJOsAq4hjSJfpdM014nERkeXea4umFlg5sNDJ
YyOn2Xx1CnHlsUAUKgqTYBfZt5awycK8i9L1/OAgy44afpb1nYZeIZQnIV0l
Sn9Y9gsKa5NqTalkALUhxbuelXfhipOl9IYp4SRvRmh+TYiypfySUC6ALMxr
VV8P8lNfY0wk6+A6kp3bC0htO6cogcGxpKLDXS05vUSa5PEmaxlZ1eVjd3DZ
0niGPbhfEqdFvl/whyKmOLh6qET6GXWfVP8iaDEa3ifkn6Drax+Tn4JuLkjj
tPiCVBkAHssMczkjWZrgji/Vyuva1p9YUecCHUzq0TLryNHp1dYDkr6ogtBJ
NMH3XVVEZCG8DeHr9VygkSEpNW+5HCBoiwpNf3z6S1+LJlEyaigpGHYlYGVc
5PkQrJjTZxWgwcX0IIpwCutbD4bJNKOzNLRX77uXXlqwz1Yu5WhZq3HmtiAj
r0PwbLpYCFznwNBWc4Donto9ePLFrPM/Uq5PetbTuxDcLp8UybXCKcdy3lGZ
Pe6SI0usIkMq2Gfax/yUsBd5rXx/yInp0hBzcYTiv0AlDLoRUP6PvfhOyvXk
3gmXbcfeBxiHNCtdZmk+ogsHNu2InifLW1ZizkDgbVgt0YB7MKsy/96by17v
ucYx5kwqr15VEr5xfAPEC+amkiVXCTcipFL3EBUxRXAaMp+GPTIHxC130F7V
yoY6f/b2COM3h9QzbnBGKgOqBruDJlTah+f4LAw+XgjJFIuHRFwZubvWKF2X
f0CM7Pe0Z34i8nOyxszU/WLF0VL/YHTkwZo/0jte3pJFem6WbMAC1BSS5LhK
2hJoaMSwdz4KdwRZwxv3QxXyr0CCkTy7idQjrEEvEIpKX10QDx7hDll9LiCp
+u3ud4PZs+VeXWXKobcY/BXYgGzLJGZ5oRRaWgDXZsz3PmAOTjoGmEoYPjed
Xze/O/ZH7Y3m860djT8ktlqE+pH4H4UcrTCIvwKmgDKH62n42ygbI63DIv/z
4GzHfeFdjDT19DC/raOh1dveti/2MK3DbIz0XAUSwv+WGiDEpU4rWqxS3P8l
k3+PKPf+kKlQsKST0KNQdN5oyVIbhuqLF+FcpNQwF+ph+oGJwVhBXWh9Rkib
YNht57aBtoMnwKwy/Er40ot2Iu/0ktWT5DSVzY1zb29GexW5mM00ymfkyZEf
frDM48W4ROQ63l71GeSv/2B2A8IxISHd8PpFETPrs1kJ6Wp1GDerElFjDUyy
7krsqETCNdeJdpJF/H5EbZfoEbWaQIqSDuJFAE1vOQVnKBzVdlZHSJEgn0qb
Q7wnFnAhRyQnpxWWDbi/VxvyeUWH/d84lV2NaTe3ktRa33NuQKCLjrqI9daw
rVhButdx/aAUCkmiAUmfeMxAqO5nBhwxdsN8Xl4c46AlE02w9nJiXPkeNEPF
tTaMR9cmvT9hmnmMQ+n7dc0JsSCLYQZ3Eq6P51RaeKlZbSlx66Y8SNLQRknu
GKpHDPrnyyYaRLRWNwwseGqX/LIYkeUopEKMNQ4RNCsbbcIRboV2N4a2PxHP
HIra9c+xUQsvnyBKx5alszDI5PYsZ9u3zjvJaek9UuzglpHiDFO0GmMDY1oF
8bYHML6WW1j1hhBrzU1M8myf2Bt48k5AW5kaikYNr8IZbn21Kol9dVdz3ryv
aPYf9EKaJZy8phS7h2DCavsx2/Bvissz4oCPT8eMKziCGM4+8HtYoBl/5W1q
kjstyAO0+zwL4g8jfCMgphkdDasTtUSEsfE2dV3j98WG3sm4o5hEroOc1yso
PKKV3+SkVFoW06U+E9ygA6yrxT5X7XpfIWJwqz5X54mkRvMjPjfvyyJUBOre
8vjmcUh5jejJCHqxms7vADC2sPV8OqIe9q0+Ak7lPJDj4/5RriKzvMmmNLyH
3hOoXVOHdV8MLVoVdOgcBe07YyDmPNC3zjaSMjrM6WcZQd61N0bTFY7klgqJ
U4rYpmTtUgu86/5FpZ2/gDwd2suuTAHy6CMbXijj/6rkzbYp/HtnydPJW4Lr
UokEsYpsTr3XAIllIEITDAmDjuYigyNtjStBugXVsJaGZSOFlLzyQtRcJ76s
J5Qp57SUTZxgHrgtIYnPc9S0PUS8sN87w9uBxYuI4m5TeY/d5Mrp/HWB5ffS
9R5IR8D5mhMS1R9w/oWZ8GvB/xrp3EdiWQWaKv5CAETmoLpIVS6CxvpTEwhn
vx1AXfqSkkMQYgL88uve+PBWOxWFAz5eD8zevg7H13sRyzIMbA2OUsA4xUmJ
3wK1fQ1WA9jfNx6u6uxS1VYMYFiKUkiOeMuH/zYcunkullddyR4Nzjhb9Zws
jR2thDVOA1icyjFYOnPRmkvnW7M17LQbio5ztNuUZDdFtVW/Igf/6bylUYZ/
X+KbCeu7jtsPGHffYlvH0PRjGQDRk1cgtCSmqkcdhyvlcJrWYizTEjirnAk6
6QLU6+Wkqpqjf2qAwfabVS+6mq8NxmHzuubcXayDvtFNux8y1H5gacKe+Kif
uplBdYHjjd8DGvVggNI32oNTFR3eOKn0ZP2EvEje3eJpeys/IojjMTT8DG5I
Z8LAzRVWONNRewiqrl4/+kWAegfw88sKY96Bd9dIRMHdnsR+CXHoLO3pUgFb
nib7PMNNTnppMQBNwC+HYBMErlG7sIWo4Q+uti1DWeEn8RmOFxtwr0YSqlxE
UhgMnMwutJhWyg3IZyt4Glp163r/605Ez8qMc8VFdmfnoLZsUVIjTTckhEab
Ri0nKkPh73XQiG43Qu1twy8Igt5TQaVENUs3G6wrHNOu/nNiELF2u0KSXKf9
KwFscC5APppu5trKixGQljS0Gh7RQhYnRQ/ByVyY1OXSYOAZE2hJq9t34Ovv
4gaZQB0443ti74urBINCbToB4ixKGOPwL/4HiF0/MCq7s21q+aseW0AQrJe/
O2lLjmgVlsxGLt/ZopTEDtZAGl6bs6cWZ6G/iiWKKn/k5uMf35qoy8MVB0GJ
nWXRnXlmWYxH7p2/ITxNSf3tk9RTVEeIK5VEeTgKAXYEHrt2xsbc4+lxyH5b
cvYW3JCOy53c62EzRjofIn9cWN8I4U4iklT6sGCaNcyQcn7KnE8eS9qMpBC+
Hh25+FG5l93Bq4qMezPD8hz+shL7xlMiDoB+lx2eT5pekJufVQFFCT/fOxuZ
lO48qB02r+Mkp1+EHtHCTucUw3/qe1kRUymT/YfeLf4LqUKHSzZVDkSuvdfX
7Fj93opt2Fp395CKqh/OLRPqkRFHSezIO59JSA9ellPQDTNRSZOUvZID9vww
O/Oo6JQvY2bikbHiszw6nc2G6tzYLrbcCIAO3BZeSO/g+nvauBc2TlEJjCz/
diq/taI/3s037VbBDfVSGKGsKgYl3c49WcrMPpU4fi8izR+fT2pb/dzVEhGl
TevIu4PP8cIHpCCLVr/zPH9b44Yu9ghn6ll5scwaQBjjpprou5eQg1t0XgCA
CKa5nleUl1zeiNe7yms38HO66/39H9rApBJVcJv5PeuNH2ga/rF8dSXkDDF/
HDcC/sufm3B4OSL2XrVj/X6JoT5tH8XWPnqOAvyLbJO8SdZO0JqXefQ9Ivsa
pkan//gxZEUsD8uSTwIOS8wr6yflyikdsn+AENSr+HbHC4jM33oQ3LuoJ+En
mpz+cjXIP0HvFo0S5Jj44Sjc/YPS3zgPruYzTU0FP5wvoPenwAno7acGbZp4
mFBkAIj9u4iMCUAshgpu9Wbz7hQInQX5lmXEzKiIED82C1UPAfe88Y1luL9W
vCgU009AjJLBRnbw0x4IW8oxgqpTlG/AqiR4AinnZ+h4pUIIpg4eZwj6I9jn
dNR2RKrgoayExGYVddp0qqe4Ye3MQYZ6jmsBmQyb/RcST56Lc7M48NYfd55L
9YG9GqB4w8w8uZBBUvqvFGduZmGaGjsCROBwXqRyAz3fahqd9uyUb6CYIWR9
M+uhqKwuQKecG1EVAktfpQtkEiE91P30k+Q2/xTv85lX5M3B/AsQaEomRkd+
9lxVdjP8aXc0Eecf6D0ovQ/x3xQOv0WMsgPmM6wlqlwbhGKdczR5eRlieQko
9BqHsF1KII0Hs6JpeZwM3eB6WCyLzRQHE8cBT16cqU2zWf+HXwZ/5S51rZaM
X+vv/nNNHFChZgtJdBBnQuknoRQ+GI2c9EHgntoh5WFGneunCiCW2nc7od0n
KA/xvapYWPi6a+mnWcSJq3l4C/Dt/jzsd6ivoZTu5UHmmaIoPWP6NuDt2aM3
mkz/yUna4GDADxoY53n2e0RTvQ1tcSgfctMnEXeVwQVSZtakVG+GdfpuNtx8
r+PuuYWZ7QGich+OV9XSE0mQ+KLor5dmfXPMJr7jDN583CeHLkt9bDWxgzTV
Dx/KcfGH158NFAjR/m7pq/4rZcSKGOB+c6vmJ08EeMtRfuBpye8I9styhc2X
/wwQLobUfw3nTLe+xwtV0Pez/gykLWBhIADCeONSVpoE1KUSgCtF/B4S35cp
ttNAYD5rU6xh2nLaHJTDtvkZiT9L1MmqJqTB6qzfh1U0/tu6VJWCeYqW4V0h
ChNRrToh68Mj83ajHxiYjYHwAmSqrm1npQOO1cSTOHQ6ajKgqwv59OOffx02
mH/yZwKmQ4/w9sF6T0iOtDrz4QicOCrtizMlhMR9kn4L5po6NYQ3ZAaec/Dl
NS0z2A3qlsQE63zyH1N9JfPed6toW9E85qMyTU+QeYuwBHt6SbVelkhfDMm+
jzcMA9VYsnc+Ia9dpcMaVTrhIzvcN0cqdkosZ0M4sP0795O+86kPFGIRqKcK
gPtu3CUP+YHhlVsDZSJ91R/MajHUTJNSaq13IPJRYHKhq0OkLuImjpMTmROa
3GwRevkpxbQ/1clBiq3v+eHPcPTMbt8UTsoDzwh85kiGYm1XwJgdUohX/UKO
uKIaumGeddLkpG16zOg2MGdAwc8gDkTLcmCgAhXUExy2rS/REvnz2TOXlGnf
8aNTamfMekglUIJ76/OgYhfsdRef23zILaBoCUdR6xtkpx0I65JxTzpsBOZs
+sG1Y850aHkW1DA/x3FpQ5XEPYs557vlBZTNvpQKQezpN5MUcu3UiJK47ve7
DvyhIw0dukD2Sz9CiQZR1YWZ0CZt35TVlFnWJJOYBAXS+DlmSca0PjcqOyQH
+17KU7UkC5oTr7kQRxZKKXyP7hRdc5c1X3V5a6dU4OeRbrNW+6++NFYRKzez
8mO03BcSzqwFnyw9DSlm/R/lAbfMKm+CgYdH/FjindHhFANw6Xh68MMhmoUn
/me909j0KsDEff7UBIuey7b81f9yGwM5mqscHGRXWzmOrTIj7sYekd/BVGdR
HB7sd7N1Ij0/9+xc07CoCnCb/j589CvMIKk02Rv2AJOi4EJj2YMeQO+S6xoB
qd2OSvNheOatQ/4L1jihq7UuAuPGCgYaxIBAyhmlTh/ufjrwc6xFx+mAOJQs
dRj3i5Z1glfcahdsHybuDArT3azssknOiDl3qs/bJUFGowH4TUc+o0wj00o4
+i7/exX18d2/N6AfuIrfHrhiHi7nHnBoAkjCukEehuPZRR3mnsGZldeOlipF
Uq7x/PlARf3ILYuJjiaXLmmfZW72Q/0LTImR69ugHuI9NmjiEPd5xAGs2tP0
QgypsYjPJghboJpKe/HZTfnSa6pJqMaBk01ChEhmXifb/nzfuYxLUIzCQIiP
2uZTVpkln9o5lna7lS9tfnIDXfFYcf4cnUYmFc0PqeFWDCvF+GkDdwTe6KvK
lJWh0smnyrhrp+jXkDJRuXozAPMyY7+kYyn7zg3MXFgVh6s3KoRJwo83H64n
lLFAtD1tv0phaIbwj+JZ1sMZMtJp2B4g/OfSBy9YV27igqJSt2wwFTbxsv+1
D8Hargicn6hFkiw8579YMPBzmnVzyE8gxx+w3ZHyEZNwUyv+D8KX1dBrtM+L
08NRwCiDhcwQhL4HAdBRxHqTPRt+gWlH1jJNGW5/E9Oev5rTVDU+D49iX7ds
naKzl9bSO9GKaEw+QcYDGIlmJjL0hfzTs70vSRQ8nwXOIhmZYXeCWNk/f/Kd
Wm6kvz1DW2GSQKE39uNjYGDF0Mv4AEaEsfzabkIQDUK3Wnl8HfVN8h9DP5YL
R7iIdhQRUoWphq1itmuvtg0HlfI3AOCTacWcNcaugG86yw8MLdMl6QorDq7n
g39NRRbDzKYepDVBO8ee1ywGsbbmLkcvXBmXjSDCGmI/zsVbh7x60KlZmC/j
HXKgiacIEh1rHVCl8q0dCE8y4h2B6373pDxyHi2HsbpK2x/oRCgZsI3kfHl1
sCqcmJxoij1ghiN5RMOunjVsT2vBtV39Ku3X2WRExoOiSXkZMpph4Y80OHDD
Mh1DjCbytdeIpk1lxmUyDnBpQyM8QFebONkpuk7IIg30M+0r1t4l5jreeI0/
BnC/TDgkmbEw557aWbm6BAvK6sSJNmC+n9XeKqjoZ/GlVxr+InOw4NR4LN+K
BIz5VMK0EiUaqV1NLD/VpdOZsTxbdJbPQ7EA2nDCSoTxN4nz+nx9uhSbjPAC
bTSskTqe+t3/7Yxuo0dy2Cp6ed8I94xOo0ULROSy/cDDJcyJC8jcLGVDnt4S
zFWJBjvGU8U7nMcNHO7x1M8HhcbmB8j1nntMLn4tIJ7g+LgMfvH/lxzZ0Qhu
uhMeERVzMwfXD5d01qAvrF0x8LR4byG3jnkCZsLMIprTnDs5k1Cssh+uqkEv
rC9wa32CERdxcRdFo5fsJuw78v++vMECJ6IFWCiVtrTetrfo+SR3olJGFdFC
spdjHTzVUzM5BHEonIt8iMnVihFgiJUvD4Dy53Cvx12KMQbzhy/gsYH7z5sj
TBaUT6W1uyXZygIRiC3jIDBE/zMePLnJWFywClMBXvnEQl4bgAFh3nZ63PyA
0vlNnLOlPHF1HD6txjFh72wpukoo30LRPiWMQ4G/eLZiqtKZtIFunWa4kROn
YpMjoWZTn9WXWTa4nVhM4od51GAoSdbd7lMF5dypWn+pcRubZ2bQa1vqprY9
AcWh5phtsqRP7fYrTXJY4IRhbbXx7eGl8OBx/TBx7bRaAb8FrWSyjFbyfYW8
LwwZ3tk2z4UjyQPRUDNmRera6tL0yNgV9nj6qQeKp/aTydVu8ogWlidilO5z
kYvX0V/f/jLdYHCngcrGacSqPiYcsu0GLrTdVBRCTPsPJyDJzmCTkxw6W9tN
LJpergEg2Sw0o85hFHSnY0cCrQYN+NYEG2hBBddjcwWuNMHatv6YJvuQ5NrZ
LvfC+2jtzXIQw3I9odLYz2EUco4g2OWgaKyGCkN/aoPbcoIFUrtFIkZ3bfho
OerT5kfYendVzubLu0r7FaeGtHpwd0kp8sJR0geubYe4Pe8Xsw9/9/ms9TeQ
DULPPPgl9U9zpr78HMiw1Uf/NOlN3mTn372wAX2GEtxuCfPA7+4xGVelWOGH
SCA/hZ/coXL11Be2egYmchlRxyr0VWK5J3uNqz2XWFTlMc2ysXI7NHCT9Jkh
ILMcq7sNn+ay+IE33nbBn1kDKReybvz0h0Fz1Hy90xrTpXT/8AXYbVhpssW8
105jz5Tx7xDOjUQRo0YZ3t35LW/HQI8OiiznNp/I3IPRTJTvsAGW2SdToioO
qeXdztWhyJb/+zUXWD94iQW3JnJ46HIo4aU/P9Pxzn0+wtGfDbEQ0Pk13lzb
HAg8vgB4pf944U7DtENSMD54M2zJyYyMoeifFJgFpsvHsqjtVYNhsGu+s7mq
urcgThMRBLCMHe81g1ERmaC6+nhCVpTjkIMskiT02ocjM8rh4qaC2Ak8h7MH
+Gc+MrS2csEv8Qzwdxed2F7+5vgtnvyVrf7YbfYDVpjr8MEMr6yWFYBJJ9Sy
Bbc1nEKXdglMpR0n5ek2GekcEjfcJN3Vy4qz2Vu6QAk2uuM9595vjj3vYsva
8V9TBFnBraPurUMByh+ry2bZtEt9iCJQ2z7gQ6tkNUextzTrh0F/jmXA/vVO
gqKuY85Y5c55tYfUAYU7TSeYMlCQwMqcR4QfLZeTT1hWpRFcFogXoVh1Q1AV
uvVc2mV+6RnBVhsYlaLS80iScT5Qwu+ZIcXtWOxIItfteKfoiUvLXQjmM1jh
ZNeOLucpiyZZxI8IrDUNme9st33peMWpyzvL4CgALEnVs9iB++p/RJvr6eew
mB78VwT4kWVxcv4Ft5VISxy+mL5RNRG4+xUmj/05zw1mRNFfcVTiIPK7ENpH
NMrcmO+zkWbqXw/V2k3rBwyoSRylC21Vnk51lqmZ2WB+CunVVJ1Ip59bl03Q
fApIhm/i1p1LPCNytmdQiRx5GUD9xGg1xDjdxCCI3BU0FgwhKDxpaHVv8cBm
1XmRbpssuw40hBv82s0Fh6xRNlZh8ShdB3KU8rOxekqBBIHqsG/ge8AcCKwH
8xbld9G3C9WUM5zO3UVH8hWb293f0pHj/PT0VikMmuPFibhHrILBqYN5lKau
suFzxDVL/mPhDsq5OZBw0J/44z6oegrsxDNbDMkwSxxNJJLr4ljHUfnTGR+y
UHyLWuyapWPTUG2qdtS9hiDl+mWZgdccbdLELP7bYUCnYzWSlwKAFQk72oy9
XN++LtYlXk98IfEn3Vk3++7CCFgmJH4jFx/H5W1OQE+KB11L8HSsNQjSp/fo
1YimOomIJpLRCruOp6Ut+g7K3p+hTOKzw7HOfSX9ovaBzPIYhy7b1T2nklY9
/zOf2AWT3+3EcO61NQL5IscC8B/64KgdglsRlzIgRZN7ioVDiEL6ubX7uIAR
oxHikwRrQrDVvqkCE8/ue75K0RHMiX11cCiOfKOeVbSwheGrrdrGkdMuOSdd
YqO8k7hAk5XB6qH1SNJfmotEnhayvn9q93cVss0QFZMm5zm8mr+7ADkgb28v
W9VdeMG9Q4Cm3ztR2ILxR3h8jbAgzWHsFxnRUGcyMfqlJH7Y+sQh5QvgjUVL
Uq5vgnisD9i2E9qHWLXsleEbeloed6lzFD+HZRMf5k80R+nk9LSGu+ibhnaV
1s5IBj173pDFodXXA5mtFTVcDolnb283/pn7lDfXxTjskn/2B4hNS4R2e5Vd
bXyf8w/UIATN7yGnqBxDPV9sDppQIH/19lUIyA0kyxf5Z2uJmM56Cpvw7zkQ
iFh9IynpIQyTauD6G6r4UMVN8AiQLVUJXA25dfd5NQUG3Rt6qu20YCgAjKmH
98pXYrwT6p9KgQ7jMDonvGNG7XzuJN6A4ksXx22i+2T07soK9NKwzj2SWf98
yBq7gzw2mAeOwkBr5DD+Y5GUsCSUSBW6JFXs74nE6MM0URlkkaXorUt5qlqE
d4qOkRoOiXnhZqOq7IBgIQpISo/SzDs+yxcmN0QTAbnW2V7CrFNxAS2KzthA
7EM+9zXOf0XdRmCQZfadVg4Cp64VmGBHRtdigyyZNDNY8gIAQboVIL5dwd0E
TBhTJaZZ3k54lgu/h6qyXl2mWGkhSlxm8xqsE41sJrtk5JQNBp2FeyHRJF0C
URfH6I1XZFAprn8xccBzSYf6wHU6jO/vAp72/iqIKb4PzThiBHlGHJfwsgWC
FODW5MDIhnWoqXfGeFtSVzBXMByr/n0gE6eIbYlZtqswvTJ+8L7BswOQs+Fb
v/RcamvvC1YxUJ9jpfRYIK2qMwnsE+gBlXMPrp5po1Q8Q3pLdZmYiL6Dp6OJ
HgpJCJY2gY6XfymmJ/9CDL9g3O3r5Pe9VE4CZyVZa8dlaD5U7V6jBknE4wzk
KMFpRQYfKU10tZrkjwonJMrdHYIm75EFKxCYxUk8LL9QpD/+is3KNb2FNzA9
mic9V1vhTlFrrCVwhatmBaFcsPCuUBdKTOGRD30K5J2+pINQhdyJislY5Ncc
8WESUB4mSHtPPcyksCYg3v6UhgLfUyCHZ5NMikBQMdbq3k4iuKgpws5UzNuV
vtZvgjFrrhu2A3TKGP3xjrWeZH0Nj8F8y5gEOURfG7wYQe6EU2Ab/gT4c1Fa
OAQlzTfmAw28dBoHS0pYmp43CdCIo6fkA38iQmTDtXSe3Y8Uc/K6V9wr3WSd
83xlgGxkClmQBbgqjD/ntzxDAH4DLWK5HDVACd5Ucta74kBBO7IDFOEikdC/
JED90VutuJFD69+EtRG5fMa09i3SpCNcxsa6W4vDE5EKoXzZ9OAnlNMCjEZ+
cpU+3dzPbIVx7yOtnXpM+mXhmloXg/pU6jT+jY4BcuEoFhqc12ZdDiM+wi1m
zkKpSao8EmDcvoi4B2Z7GupattyyoMksKOTf1b1W0zq4AE8bvFouYUaZwY2r
STycEhB3gNhPbuBbHtu9NkVPkO0mgdPwZmS94sSmfdyBAEGkqx+eOTqoJ8pM
O+yTpn2bkOK4ShVXBQMrLwhTJxr7Xj2nHG2qKEaZ1/KHzr5oHopoEV+6+Hol
efG4skBw+KwFrw5tDoJLkR2sSE3U5rH1yuFDzJ/it7JmtpDurn5G0lNydio+
Taet5r97bNbhMDNFXKsMstck59eB2h4plzqrHlFJbytizREUdlaCY7o0i2yn
hd9yXt/9Gv7Va82wF0bg8dsiAHw3sjxmUUZ25rEwuIqV8lELGVoCJufIkrLk
iL2jxer1K8aOSSptwS3vOKOEOnA5zSp5y1an+isSJ2/YCpnI0fo0r6FJn4wC
d5xyRXR2+7aIEYnR5Rtua9C2CnDOGlZLZdr2M6vYA2LCoHnjBY6Y9+ipwgO3
UspQAHDe+VA0SUVd6TDO+qVp332sCvq2OuSg45WSUVj3xpf4tWz+QoAzZOEY
10Zh/dv3r/ZDwV/X8ZpQxLcN0dL3pH7msITHFds+YJYIZoIgMxpiG9lJM/VR
4Tk+4785iSML29cIz06YEZogrbshLjuOtrdpX0DKyiDL2CgzpfruSSbTubjQ
vJI1epBqQ/brao4/ZgjCc05StBwyydiPc5mrX4tnWf0sZ97W2rluKO+DJYZa
43C9owzT/6T5JrC6AgzC6blJgXozjcJxl7Yl3XOYeCuuBKxh824/7441voQs
Viq4PfufcSY550wkR+50mseIMwipJryizXjj0EiBwxJiRlb7XJC6eJQbc1ZO
5QdAX1vPwf6R/1tLyiHt/mVtOI2rhuresa0ALRRY/8w/4fX5KGyS5SsaYYmn
kknWwQ/PnU8tTKv2PhqEoB/s6P8Iv0bW01sAD74rWBo1iupmGNAwB+qI5+5q
GyRVdNxG4n1F050HxFQAWnkZDK7beRoxi5G2QFW+S8tWq0eRj6/sEUJkXMxs
x9AsjOBA1X8VyvpyaZUCt/gNPOsS1XI6t2H+ArdWwvPAjwBuxht7nvXPR6ZY
B2KwnMMfTcEWbv6lqqllgSR3xbG/Js5QP2IP8Iu+zthQ0Y5ZBMqaUFH233Oy
KiPmRNoikfvD/KOCVLreWdtO7XQFDsho9QBEu1oG0VPFqwUQHAu3Y8ERy695
CKwqtfy/fdPWz66DfCmwKQNNJoTu+f9FpzXBxzD1Kyw4JZqDXC2acy1PuTyJ
Mhvo/5d5DeIjKtVsLhesZV7OgyELHTSQDIEmAvie3JEHb4a7RL8qvbW5H3MX
WCw/3i/H8gElYYOfX0MyQPFPLMaSllj6qidcu8ckCf1hgezEgWDvYA8gPmmN
SY1w+0qHdowKgvixaBAWS3tTs+LkTCg4nHHknQCuotr7CrLn4VnFzRTWVhz+
GiI7CA6Uo7rAEZdU3YUYnWBo1ldenrTjDBr6XRFUYayvJqbSUuw0flKmPIFc
Ehh5u25E/++bfDqohgzKWlYx0cE6xaBK2XD3LlwQidFZG31fpTa00g09Ty4S
ehdLdiQlACVGt2q2wnp6tdc8eDfhRS6RWJoDlSZdjEOAnF3VFkhJWugHaFcS
6ZM116B5EOuw5mN5tb8x7liTdWH0flcAqueh6TwrL9WvWcF48k+ag586X0Nv
tDLsUogYWMeZbmSCrcwIFNDTQD0Z5tkuIyCDuo9KjVM9bBGIeRgmpj1lCA3y
d2QRL7rS9JgAP6pZxb6ye4OC5fLN9XT/V2LuPakfVN6Ijq7V3ZXek6h9dVqO
Lb6OYKrygX9i2b1OSulIWEqGPXriDwqw/Aki7bJIK494HK0otf6nQ4wLfhMP
ojGSdxsnKwLDzGIsyJ5L93AMgA0LK7EGADy1e0N1TuRfIe0UOI27Wrea8ucz
5jCnkvoqqWVqP3h2CYXVHkrg5+H/qYOTqVlOJqW1c937KpLhBeFFOjCIF1fk
51quXNmcA5xuKLUN2iOVZv3jC6Ncb0hTAqb1VfFBLMI1ezRncAN5j7gyPRMK
wcWXxHKVWhXkpPlEra0RR+3tTmTalIugOz0tm9qWepliYlE06aqiCingZARo
4MS/NBI/c3SzYBmha4+s4MDLNJLnOmKFdLYYBjeOIehGNRaIfEwi+/shEq3v
WZ6mO7eyXTJ18uEgz2g9JGFLo15ZhLxrjEKL811uZ6jYh+G/GmZ3/6Zcm2VR
m1xUjwgycwnr8nWmKZwZ4d0aY+3UGWKU8dAjPRCHZ7l7OZF3Lh4sgigduF/o
3a6gfo4EMOaW1RW8ethqA4Jb/FsunZ+8pqCY0NXpaZ6qnw/5iaV5kH2rxQ59
/HKgy9Lq5V/SwmvxmX35zno6IuPBv3Ue03sRnqYvankvej0bvmNsf3nzplr/
6TFoNLvUVYHODafF3FYMKdIO7qWX1ubAxntiYRDEiMNFdsLDmCt3ZiBxxDvQ
ZH/cUCIypvHojVE9Cvn/5QrU56M1/OUswfTmauzgS1PghAGaDhBqItApqzh3
LIdOfpRZBLdzAYDNzKglMxpRbrOUUEna9go+THW53o+xmW1Dhw0ooOTb+jMJ
ZiMzYRBdy4JQynye97xoVF5Idg2ImlHOp9QXW/6VlUVjCdZEcEM9vNhZqjsd
gzjAkDWjeaP1rvbuqFkoqc3lqSFvxurguBMxikEWTDAn5kj1D4Tqu8NOfAJH
UqSbyjb84dgrhIXyWtLu4a53sPJgL4JGZzvPUbidxxRLbZGNpcOrjlx6r8gZ
gvJWIA3zp2l4mHef0URsYnCMHlVPmkLpu6ANtTTNWEeXvAusiQVqrVCG/Nr2
nNrkd6PXOxF13r8ddZUdlOpG0GXhFAxRybflYiq89OpgQ5TDq4S7kDIOk2FU
n90aHswQDaWOnKmnjP+eSySBtMINgMl/85Y5nORH5Z9quIEze9gnftcS5/sv
ZcHQjDAvQRK8HYEKoFUyeWn7ycj5bdfFoknqhpvMYoYQQBikgMeKbpVfp0Bj
yoGcMcMDahu31z5Co02e4Zc9yiPcRDrnMpkrsBPwXPufYvJhUQeHsADKCkxm
nXXlyafK6KpMTc5qVgUSMKM/fVEih29KpjZ8FHpQ7F3ddoZDCI6n2mv56IP7
XS6tTdKA0mK/s49G8XfjDQvJEjEAJcspJm49xTLnLHjK0+K1M6xgcc2oRoSb
GRgVvSJvhrEWpkPh0sHYjFbWmBJe5nkpgYQ48o8hQeO+xPyLpt6nh/DSCU5Y
KQ4E3jDpDrti5HwQXEg1hLdsTtXz6Z882IRtwn7cOBgVTwuDVk+HAGZCBdBD
vFaXRtqVp2ozf4Mhvpl5xJWzGHzKOPvJFDeMPEOjE0pFpO7jjH18omuUiCNv
NcuIqdbVCTc6oYOlEsYin0eVCveFonkVlyyDn8LfkchjIA+K9o37J4ZCenye
GYWYh4/gpQiRkydDxiTlzBrYgl5rtdbec4sEUNnijcdRMGD95RvmEaN8+JP/
o2ui/HZvn3ss2VpaCW1ogoR9/9vGQwqRokfGB06Grs6kNFtQu0axk4X584qF
46n19tsQLSjWTPXnC2zaCd8qz7SPe88GnVYC5yGvygWA3KDesTFCn5qYYdwX
SNVOdqRqagecNAQuLlyZZfAApQtztvPTDaqXOg/KYSiaEh/QL3m/ZfawAQLV
mjqi8u5kPOb7146KXqjrhepLVG6oW5JiI5x2qBm7nlDIhqGMz3/j83UAEUJS
gfcIlDWPRqwSajiUuDJduPgagIySwSjNQqQbkBrw1pBrIi7eEfKlqJyNqJh4
HGSJQr5bSoSTgHSGAPXgxjWyPsIfV/Y6MGE0yQoZsAxh481d6UgHO88crRt6
Op9uQUOCjJPwwcHxaGl0LFhYM6lGP4mtxADB9IBswedpo+Pdjp60EAyaUObS
VqxDFm/89eC86+Pzbs4PfIbof9IvXUjK/z9sifhygT4Uc5C2PEjhwYQ1xCtP
T+ihhBS/wflowkrUIQKulz0tM/SfUyNoKTPVzirNtTyA3sRff/Ht6Z/+FldT
700uG4vSNP04k1ZhD5qO10dVKYv9ZE2Hz0Yng5uKTbQtV/LSLYolJkLlK6iu
6ZZdFnH4uyQ/W6CWGjuMWjgBv5/AxIw5sYvbdxSaEtl+uIe7CISSk8EPS5iC
8kTijJiXVKwGs+0fwqdfmLhs+6/VV1gS4AAUKFDtvvZP5a3Gj7MfCnWvXhP3
eZXXx+5TXadECkNwiTS5r/dNSijC+0l99zT8KuSBeBglkK8OiScvONTh45fR
4oUjzxepyetR4cw4XbJSLpFjruV/v+KytwjpEC9vxtTdUeOh87PK2jWDCUwU
9Htc2G+y/I1Denf7IKRy5xT+QahPPC+bj2EHZpQdZaR2JwX7yjdO+aivLgz6
oT/w06eLPBnYEhMAY9Md651EGFNNOLgA0B/FSXZMkg3pauUvySVDG2UZ7aBG
0b2gKUv0hBjvRsaOFVNeoME4u8nWurqm6vkh9wB/BCcPbrv1jwp/EapvoYLy
oRFha4sZfwKNf7m3WWNH2qbYl6xwW13TMwemrh7ZqAl+qCgJMFdy7gJUU59S
plmIaom7bTNEFY9cojhHvzXKVsBBe/w0GJnN416ehEOgkFR5MhhV5T76SdtA
OmZSUPFgo2XRThKkNhGBjUJxk8V0NYUZHgWLqP/L6uUI037/KqwMgtm0pfY6
VItlU9XU5VW3URQB4KDZSUS7945S9LTsYyXIUGGtp5/1e6mb1o+E+F1lWHms
VTxtA6iHaYJDDipCBCeLmAKo79r/e8UQaNj4Btze0QAFbOtqVvW2qscTNPuQ
p8m3JlNI89tpK5Pce2nYh1Wn6GgokeSqVmhy7BjicImRb8JIWiE4tnMaEEWt
dLT8LIUt4FX14kvACFIBk0Hr4kf6zZd6aRs3WPcG6u7TjsWhmrr4GzGvlLLI
to+WjBWRG9BbLZjOZWnztI1u/TbIewTVFEAOLe3IjppuNIEou7z5gfi08rbt
hfPyIRhnvAnKEdwv/UMvjp5K6XhunW7ZUyeXFcWmn9drcEdIQejX1PdyEA1u
yrL4SBUXD41ER9fjBqswrtdOMT4TXCrCyzsURmiN+8a3rFPATUAo2QRnOJOu
11ttOndjIvzNjUd7IvjwvnpT8F/wOplWaDs6rAAnh5P0tPtAMycrms59Zf72
fKpOW0pUVl+p7uaxdQVSvG+7QkVAHWkdPmkl7vyx6kJ6HYd52uolwFIGS0bG
UUoOT2HZnzVm48PhiqI+OEY+qhC9wGIUUXUViUG2YLrrtm17XcjMbbjAYxj2
bLtLuvNZQ9KVBjlri7CcBMxWP1cwj/DVnXetyDlECZ+PqViu05309kprT3k0
sQhXUiBhH2Meu7CAdBMTPo+EGXoO+i6Ex+Gvc50qOZVJELxHRSbRTDDP9KKz
uZZ/K0+jG9KayT4QWshkABqn0jrzaySJ3Azr4I8X//oaKiK1zEulrhMpLDPY
ZSkRxmGJQfJGlh2R/94spigK3vECNaH30sePmvMtffJ3hDI7yQsvnpoXb8B+
6ojGrQy3eU3eDT1gzmMk08PAN9Ksq+A0rzIAocKH+q70jV3a7DdwfsagsOzA
T1qGmomJVOMlvdSosiXFDPxx6f9qBnQFpO9kXMy+lMKSnTlt44E9DWKTc8U1
HiEqjBReJpYNnU4Kl7f6li1X7ql4Ppj8Sqln5eILDwXnILyjpIvUmU5CT09l
Q7aUEtU7KwhBF3BzNqYO4Vmrvtjl9O6zQ7vKGRMDHr4avPiL7wRqfU9tlduH
sVlSrMeZRU+NDQOw4pY4U6Vnis839KGy8Mu7d56UvJl1jWGKKMrMqUZWmW04
FfzD2u28loHdS2mSikTdrKm/qZChkviKrv5ZtAuNDibqJBK5mcoXyQTuPzjn
kYBPSfVhjEz9W9j+q0hacVnlEt2a6/YrBlNNkbgsRji7hobeneGkxGQsdJSc
XlBvATuSOyn2KxVwToMTRna7xvySdjKpng44NTY+R0jmfg+8DSGhf0MPbu5U
zv+wJOYaR11IYKqnEZRspwSUqNu5lOV2KFYSoDDg9aVsdFHx8WBroJb5xUHB
veXULftpwNrWlOH5AUBxJ7U2p61BMQdfL5LG43JjE0k9mY0OMRRAbeqzjnxm
nGvUzHzctinTmFjxta+iShfPBwgtjfX2RhDsVmG1T35aw2J2o/anv71H97Xw
0duZPPClR0zoXJUhBq9yFpSHPVWY0i+u45p1IVFGgYKsZ8ESiNLEKBCRUw4r
1JNOXe+KaU6C8zroBv4o7zLnV3U0qcclwN8UN1hpHq/SF0hwD5Tm4JT2KXLf
UvkmeW18n+UhUKwbx7ILnBSP6hSNmYi/QG+apPh3f3pce5pMLMxoH6jovvD0
eUpDOyKLDwFEYJPmo+CiYMHcXONeSnSCatqsISk8ZqxAnyyFNHEB+LkvL6Gw
zvF1n7UJN9NKWpDIwCX+FlGSq9IvCfoeUvSgF3GY5XoB0Ir36ycdkcofHiIV
HOKmjgR9rDyPgdQ6vDA6umP7halDwGQPNygCgWlvkPf/ZHG77IIz9Kh3+Jmi
AJKfpGhYo8jYo/wty9MMIBwadH2bZZxldtDTNb9+1Tf4Y6Ty/VYSazelFQLL
CWaTL6AeIwJRDvUgmqb58moAolYY4+ZHl7+8eyiGvb6ZhG5V2hLQwW9JwM5S
xzGs5Sn/mKZZ0xQu1cEZS62h9MLUKJgwWMrBIbVYaGz055Uloa/ohL+YFePV
KCDPhwE9W4oCNaf1azZmxq94X0Xm/16APZIvgjXfHZKOyXHLs43UwfWbmUxR
nvhuEo3XTuXusQaIznN988lEBGVRMU+oDpOhr/36W+FJj43IFA74xFyB4Kzl
Tj+BU2m0RU4I+S6VA1jtk4NpstMTWJHI2rJtTYfK6j7igUTFt17pNEIb6Azu
Gdqjaut1WvnSsw+SfZK81hAzDm94Z8wdF4TC1Yx/rDKiqArLFYKlAsJk5Jem
1NWqfwUXELDwV38IGOLs+rdDLj3W4r65UZxoFQi9OMVmxSI/r+3p6FCVwJgO
/93PXtKBioar407FTbw90CEnzENWAv7hh5HXjUix/W9wbqg8VenCFfnXLfv3
1qzrHej1lM2CyqDE94JA304rLf0obgkRADECK1f981ZUzFoH3EKw0Pc8FWys
DJZWcv9yht9HWvsp4vpRVNRbl4gbAVPmfoZHVPIrwO/TpPNAzD6V/wjpSAcM
LZz6nEjbEMMtMQW51LfwAPwETn643AkOSc+dvE5Tgd0wiCFuikUXNI4TgnVR
Jwj54fdpN6QhMsCAgYocXCo50hJyD1e6RO17E1twtXJTgOMhXzw2TqhXVaHp
mK0JiSPFb6qHKqPhCMgS5QMB5eJ3HvXhNld2yom4sm23f3qXJlk2xlDhblhk
5zZ+uLlW1rzkhpc7ylbQ10xllXXjMRbm+o+UiZtFfbK//wtWCJKRw929vd/9
CYblITjWrChrgltc7+pyvxYIDmZFBnDhvd1iFE+NNoCsgIYnyu22wTWLflf9
HkBum9OQMBhkcj9UOqa9gCwNEFSAPIvv4BGBpdkCldPPXnmzMJgaXT0KR1Qf
Umb8QUnNnyNgvZbwnR2TnQVwTLhV1RKKCyo59OVBLQtZKRe9J7oZj1I2dVxN
OTcSHOjCQqGfhTYiRtNfKELVkWMoydesGw828wxf2AUrqtQlXeG8wL7mDt5y
ePBPhXdsAar4avGSSs5c/yMa7p91oVf0xnYPOM9Yrmj+SHTCCCnF+pPay8UR
XtC82Z9SggxFwZeVqs1vWts1h3zUtZ6xB38VXvx4p8xoXeYgNCPiMg9Ih8Ra
wKyub2u8I9V1MoGoSUrc43cpX2zW6dmze3qbxb+wGjlXQ5AY0zDOYNnv+xl6
opp8u5hgTT0gbgqJT+YGpSsFkNba9jD1iCqFgVaB67dh18a6Q5nOjv5YxuEf
WJTZ5nP9+zTR6dWEarPRfvxNUh4UQjg56HbL8iMbjHLPqCuBFL1kcrCtMt0T
TImEKvjPvecr1cFgI35Gtx1wpLVJQnukmyTSh0nM13iCmo+L27GwoQk/lv1o
Nmx0Xz3zpsiLWDllMSM0IjMqsQnREBfyiOOc3VX05FQgjbchNkZBl0K5hf8a
wGjSawjKPjXIbjqoXQu1RGASRD1NnkOUC/+C2Ugyt9Mq0/t3ulc7e3ctER3R
2/hGwYkq2lzQ9qf9406kw9b39Eh75e/411qifuloMWlvb86s2hwcVdFXKZQv
j9M4WFnbAydFTWCgvksUH3/5Kx3IX5JH3uQXQFVzfH2RShRBIZTUvLk3Hko0
B4jkrwWRolMcppgASWUbutEPsG4001NajBE5BRVJi27QAv2MDh6PDqEEEDQ9
CfbKBMm1lujYBbCorCaYig+00NWasvSU6CriGrk898cWmDFWhOdRfCHYktTP
IwLRHSTiJWWMNa8BsYGxaayhSOGV3SWmQTyGhVBmL24eHGzI1GowJPUwzChm
tTbh2RcYhw7Oe8dgWt7tDazuJnF2Z0eTv+j+Zi9K53DFmM1FNfLOCYxtVwTf
POu9aPnnWDR3jZnbN7htkcADhYxPjMFzyFNEVWSz/tSEXwGfwwZPWxS+JYBb
qSAsAO09TD4ksiWqKnLGDCf07H3qNqzTCSMsdqoXPjhcyCIlXOvdFRPC74Jh
6oKZpDTCcUkkIf7Zj312YqASoAWXTEcxqdCdaJliaAc6IAexsyaZd0nP0uOs
F0fRsIZEOY/rBR0EFs4hSUlXJaUzVxcmJWQn39/Mj8SgbPO+Yy4w601BugXw
PMTYtmEZQhqceNJsEibW0L6O8gyg+eYu6cWeqDtbXQjcth+/3oUrieYnXQ/X
zTE6BcQEECpVFPW5OkaqfMGFv6UqcemVzx8UgyeXyL7cV10taFZ8rE2SsCqe
Pji6nUs5XnYJBvsNaKRMLNN/2gPXQzQ/J24zRrjCkJV/d3iw7xyRWHUWrlNY
0qHo+rEXsY82kMCUnIJN31bWo7ExvGBakVegTicod3I8Vfdfc5WFlU9w1BbN
4w6UFdAWrmo99GHj5/+7lUw98evsw29WKx0+lfZyLWzAFUkLnBluQ3pAjPDM
6rbexuNcOwQsfIBpkQZcCwSjBVN7dD3XcDpnLu8OodT7oYvDzXf/BSSz0G5p
FcKa9Ornq4D8PiSa6mOCIhxViU4gAmQPYFCcfDjZZNUxmTMQO+2CZLFqFVrn
pb7EWt2vXBsFlEaNFDk0k6I4BndFS72nF9YkZIcDw/KLqn25XQnjdShfMRB4
WF12NdWSdxHWv9fCbJ1oiAtj24ujivVLsr09AqytLHrnxxriQxFP/2yqC3Qj
Dm6ELkuZQrnT7su3P8lhpRP2686JGAOGTCaVbY1SgTfcNA448FcbVZnAKrtP
i4mO3cXJj3yGFMn3iHjiR+DjuGguiXykzcgv0PuH4OMSLCvx8PWJZ1RIkBi/
Lw1Kb6F14Xo2T8YG9Abe07M8iusEwg8XbjnAqqjUaMvbdex1jPMbiQ86Yy2X
u7jc2PaajvlWsoCqlfPPnV//OyOtU6sTKRGwyefTasAKEO1ZLd3UrUvb715J
TGxR8wWliZ5n0Ll/vteIezFKCyTXQX6Y998P7/O6obbnCBehJywYKFFMOSov
Pc5K/knXkFUz1Cte0St0kTYPkGj7LbR/bOoKZdW6mEiFGFSdWIezUcAt8lgm
zG7EvvPdf2Vyam0yILgbOU6f7boToEUAeOljpGSGlC4hjltqqrfcFAvb4Vtk
VYuQUFd0nQeNRlcOKjTG2BmblN/S8bFYDxiFofWgUEg6th3xn94nx1iwJ5MG
hADcNakfJd724OMryBklxG3YzKmzN/VMBnU8tn3h5pmDht2bG8zgG7lZgXGE
mxU3NFTeUU9wZVdYC1o0In7dW2muQ4uvQslyblCAUccXvoOQO9D5nZ2LkGc8
Fw8uhHUt1swUapP+ri6H3Y5qIBV5ZP4cDezjXdGZHnezXurwg6hLN/a5KI8u
l9A2ot98FLBG0+Ocp8GJzgPvzW7VnuS75psO1DZy+Vq70mnPJWbBWZ/+mq8b
XrA1R4nMff6Duf4g9uyx9HDjuzC1d+QlPWr6JaW+gZ7FtnfVjfXkWQmTf6jb
c1cZTutWixa+Qc2K0LRYl6hgcwh+wmFTl+yiiXPD0Uav+RbcH+ctlLau4GTs
g6Y4mSyOMWSDZpFuqPYzpMP3fNov6BriBV07EZx3uIjH8f0WcSEJvOj7K5Zv
sgp8nB9UGvNNUq3ZuojvmeVD7ogNL7Tbnq7oEbmNT/IurL2D65SZL0qZqUlq
IZFqrQg73NVCfUBLEirKp+6ZaihQq+2qo7GU01JI5kNtVXP/u+4YnwdR0KC0
VoLzPpP67ybwKakLCZlLenmA7XwPv3ngwqf3yC9UUncpwzYikalIwEMgidbC
SvIQ0Z/wkv3TNsqnbGsRIN1G81KzftgE7Jct6Zn4XmBLvxagcranQAiKFiPY
+TApXHXyiw+xDbtSsD6YfoFwcL59nKGMUeCSEzZqzZ2PODVxCxIcfmA7Eqas
OY4Q4FVrohObkriw+wqJpEp+36xXRfwK7p2O/Tnb3lzVYNMwUjyA3ZjCCjHT
CwYOj4tAwN5vCWPr03zM4K/vCGVjGt726XqFSk7HvXjIa9GMsOMBg/lt31VH
xRJPgmdU5kIeSD4962PArmDUlCKwd/S674V8CsnbhiSNcBHkzSrU4NKG7wdK
3j2diFYvd10aRAChMZUzV0a8HVit0rqkjVxGaT7TjdmQ/4RuZw8WB8UfcVfG
djn8H11T2FcXqxo2y8obBmvQuW6Zd1A7pl+7ittJq6UtLrIym+AzVxyvKuas
2aKvSuErMz1ztGJHIu/RX4mcGzcSvVlqf/IH5Tqfa1zeP0C3r1OmA3dnCGrM
WnuYPxLbmrLeKVLrNAxoboa08NCwjJQq3watjBq7MmEioxCNOZz7NVBFuC/I
/BW/1u0fYCrLJnoc5SJsW767La0LHoGJsJxkNsCeP7PlOWcEK6O/xr1Y2XZ7
nBV0uCa4JLbN8ddY9YHWOgicn+II7IrAVZUVVsQZ/xDwrYtxwDkQPscCU6HU
4+Mqym5Sj1mxtXjpYI8WliSB2pFPcm0bszfkdTbe/mYVShdolHMdSwwTtFpI
BkdW3I0UkCfZ+5OOmuBl58JfnpHdXv+f9oIA1pQn+x3j0xKU229tbi392rpl
TDK04MT0gpetPC4BoGNOBTuZE+B/EhefAfPbjYQMCrRCrOQALQQxLjeTOe4l
c2p+k6phQ+J+6oLg7HIpKYaKzbIsxaSFVJXkGeBk6g9NRYpVcV9IFI3FDhyG
x85S94XWNAueuMtHtyDGDPxGy2N4rVjXVzMoR0ZBAXk0YV+/YNDeh70N7ykz
rdvS/qpM9xfL1VAaPfaG2p8ZYWl9HeVFuqEaxe64SWY8I2zVECGhpSHVc3WO
iJtX5E/8Xk/V5KxbsC49Yx2rNGyEqaXHvLPLYFfxQ2PZrpcG1xK9VvdxhmnT
N7D/0XypNLh7t5xPxCFTleWpd6SjKly/QSBVk+mwlTqyA9EIldgd1gi7PCJQ
9O29CH42p30el8k8L9v8X8+Tbu10kN1xOvcHW6Z76xycwlaFTNKQZEvq41W/
b7ShrVreEezucxK6EyA6DUmOAYVbPT2fzrKYeKiKmfOUU9Dbn97NhFZZqJRQ
iLpAuHhcVQu2kd42eL6MjTxuEMZLAyVcqD9i72k0xQfz8LXEtctkunjX/UCY
RrPIt5tREmcLlN53hdqKPTfcrr+N585o0ZYZEIWRfbfjDLmG1u05OkD4holg
K/jBFooFueoLtWtCUmQcGKEruMxEAGeKn+v8JaFDgRCp5VVbJGYDt89RKRNl
IHpo0Qa+tRKHeQeJwpWP1pAW62gbWGq6frIhI7aNwI12gsf8nEoHKQrDPmWe
9t6A/n7eUkVfGgep4JLWebnRIwjAPVSHkAkpvebVh+sqL6HTz/ViZCmDTmhq
EsDMrzDW0ygRLzFabbnN3V27dMcJbjUya5XR8AaeSCetLhBZMr1mvWexzIRy
u6yefH5lgJsVIYtLn12YBQxtl/8xKKMWuw8p0h2OS17q29w8Tk5sN5LJsycm
WQ8Gygwc3jT+MjTXDdRS+ceDLIkVB5gCSM808Nk9YnQK91IG0vW2AAW7GrRH
TnfijULKi7Uv6/3a4l5+u2uuTs0n/8fi3UwbpZaX05R0xIsejP7q289nlWo+
ZfAWoFM1dKQDPkAhIkWKMNJA0VhawrWEskw9DGeeNkFHW4L4mLKBkbOURc6A
ZDCD65GHUN5Sy3TITbfrJPFadVGyYMovbO/vpMhTrtyYu1V1/SMV3vu40vLg
QJk/ExDqafzbieO1Z1A4JjhYgnb4xmM/RjpphobPKW5TtZBRp3ADhtJXANXZ
tOp0T29ZNIpgktdtxfnhHC1Is+NGgp/JTzThZjWLt4sI7aefXf+lI4tya9x/
hmRye9ZTx6FEGPLqRxCpRq0/2DDXoK7A6YvLl6LDghPa+8jsohCcsR6N6IKw
Bj75pFQ/lZHKqcNkHHiXCTrGFL17qjMfCz7g3SlL9bWMk9Snm9AdA1gfKAPG
0OiKXJn4DJM4L/2KznTGE5DGrtwBOIF13qdJT/ArjdGZek48yuFQg0nWy3lQ
ZfI+S18xA/JZYvtbrJbB6cxmlRJP/4D45000/x3r6rjDy+hbxuhMIS2Benvo
dgGnSQ+WO3BaIRxyRx95kYTPOJSO85579cUOQY4zOZRJrQl8lul5C5vhWDuk
yjF6nUQvYmxtrGTqz9WXdhy3dsd2oiN6MVOiynn/Bu01ajkpafPqSGKFnOIv
4HYKIm1+tt/Lddvbx7TMBzRWjp0Jyb2c44zTwolJYYy/pG6m5hCwjFxWKIwJ
SSvyjh7vXH8JUdEE97O7P6mZot/5KYltcK7xtoTXT1F4FInoyCvMf9/GoTB5
a2doB2Jgwz94ApojR+LnOiATsKCeXSt5zfoL1mc/bnH5x8W7S8ZySycIykKO
18aoBU3qpXYE6uLV8+NQdmmdfVZnTM1Yup0Zo0ZD/TRyh9/PRQ21Hfqzf5dg
9QuC63oNyMmHYlmGtqaxUNq45ckGbym5ee8fH53Mh2EoMIrILM7d2WxQsRfu
r5pOdm5ZntNF3hVMBSSfd6PJ5r9mTN++X4gTsOqFAwABkfOhxmMKYL/A+p1S
wMs1KtyGfIe7t0tHdPjsHKW/mDWJKavVwrKCTRjF5DNwjQsNzOF4P9YJ3+pw
hxo/6CT2PeXf6D9PAXEbyPMwpPAQIMgiYSU3gg93nXZme4gz6B1StWFCH/XZ
LxF+t1La6FDwJo3rSf3Yean9ghkACPeG2+mF7ZfdWgi0k4aI53mqBtcMpVjZ
8v61mw1wj/16FNsrwPHiPu5YzhQctws1sQr9CIbiLWtMNsIjfiYvYm6gjHv9
Pz7wNhcUavBN+ob/bFYrEUaOrkyglPvQB7WwG23HJOHDbFi4Q2tFoQt0po8O
dXJa9ocAkToqIU4uwhbIkoVCGVhREbe91BJTnl/FdrWNM5bQuHDnpda0Lt2c
1Fk4RJEVo7+4Uj2aTBvoMeQ0+ajqOm1kBVLxclRWG54oHFVjajqNzZ6c/kO/
vvQFgslcJ0MfZuBhoFMqPKrrB4aL8/m5RRgwLZYEJLsRsBifXc9CbgBR3Aov
WX1LHhHJWJl9BG6JE8Skx7mhRHcbDvF4TrR5rkB11PdI3yC/QD/iK2gWIEdZ
u0Bea5XOqT507pMAEtIG6LpFCNMuFRMJfDOLAuGgpCk9ez4N+xXM4UjVqO9Q
mT7HT6FJgVy94kr/OJiFvbxzV05fSQBXZm/WgIyCrT4gS0ZPfzHxHmfyp4uN
025qkxdcx0zJV7VjmKrMZ0pN/cTO4zKjlUbN2fqWFok2ul+99mXXUjbNu33n
LZ40r5hleecEyLZgn51CAZtKb7WEWCePkk96sZxsLL1N3zoKa7K6cGIZQO5U
ZVjzOU8j4X1X4mfn0fyHWyTBQiI8mk7PAQzkb/cpbkB8SnszLo9FbnIx4K3c
6eHaG1Dco5HhOhS5j0WOpLEHNQPTRzsblNtnjOAshnNTjYfYB/7JmCG89S6X
aXqwc/20fe8Hd8qa/M6J0WuoGc0T7kw72izixK7mr/A7QPM5RhAjFax1yzfw
+vqcIu1QEdgMUvIw+E2KNThZsV8qqFYjgLa4UHplMJOJrqfAPcy63CjtfUpX
hgLccByL/SNvd1/Ec7HWd6/SwwJXQx/CsbKNzjWsQYLhzkYd4DnTjK03MWg1
oMolcJCFcaWStBq+t+P2cNwWI4K64pViVHK8bj/BFKBRy0YUvvwWP/Z8FAYH
ZdjhO5VBPmkNH6+SSdZhgEbK2vflV27XksQLyhd6gPurtGSUOoKR+83jVwy/
OAIHA6uwS9OX40V7So9E9zYSg5z8Kthu6R49ggFNJbDHP3l3Qpo1EFUw0lzC
iKmEqUcbH25OBHVkuPgV85ocuWZpSlMRxSBfbCPVWdfh+WYgBBOX8MgEuPRV
F1u/afD4wu5sKOxURZLh2LgoCcOBUTDChGfirLFkyf0F1Gr2+GgyFS4kqFHH
5PADnoNcT0LwKKYdl8SeGXjbv9pcXLwACSpsbseuJNhNLG0LHvEwXwqRaaLN
CloDeTfbyqrWyZVz4t6qXCdqEJn7nyHE2n5HNUDVmyfu2kVeqP7pftfDMb3Y
PStNacBKz/s1Est7fib9Qp5y5UNsSrkVUVJ/ecYrz/VQKWXicN6bnV7VaXsz
o8Fl+5/9KH7u/NHejDW+yQRVce9ylwrf1VOHgq7BApmtMSfTmCMIOOi7mBv2
5SKwUcTN282SxB8BeyzYKDmvYoohFe+fo7Z+HptBcYxLMAFvprh0Y51PSFxn
r5kF1Li3DG0ZouuFIrf8IAr7clJPb+geTJjpVYMbHEFoMHdMGcZHk9DH1/MZ
AA5QS8kfsOYUhQaIskDexHldL1QZc21BxzxtRD7JNfcwTFsfbeRk6ouhE3ZN
xIAJ2wwSlAAM2lG1Sc9F3InLlpXUgwKIHrcHO39HrR55l2CikY0e/heTyTwR
6t3EzZtCiKdbHN6PrLoKe8O6ZIFg3hrhj1PyjaPCJsQjUrhwQ+afNlJ2WhL+
pZWy4wEIxVg0HD9t5sXG7UDxaot5n+9Q8Uzu3X9X1YzGOT/zYONIiUxbKH2L
g/agjTfUTRBMOywiholLNKzSzz4wGjNiVlkCQbuKUaAfsMfx3mwxI/EUrua8
n0ZJ5IEqgqr72vk4tuzgKecvw/VKqIBDXBWevkuty+14qQAImyYux3QxbCzF
QUljO66gtsSoOhXpxR3OTv3H2QFIJN3XCcjLhuCrtjy1sADWfxl/mCLstuSI
2hs4wGqcArF8cpiL5Cjza7TigHO77nB+bMM7ioKdCDfG3AvM17d2GpO1+LAC
CDGDKeAzI8kIFGzNNgtAuRjxRFmP3b5590rLkgihWjFNt7CiEMUbf/ZUNdIF
l7R/bv26Mq2jq5Hkop6Cdg2y8kDdqNvok+APr8euuuW4yFrnZGcE9uJy9WTG
gVgFrb2cx6vgSpmmTIIx/ifZirfXfFB/5B5SnH1AkfdGyQS0Ww5K5xOGmaW/
iMHOoizamdatkhmU2iFSbR/ts7PmqUChEgtsR6U3KxdesbwMRwTItPvhtPZK
fArSqrUWB+hhCV0gBmyICM/r/92Xp95T+59q02GgLZx9IoMaDgHufnydmDNY
9gnYMf1brPdrYWkdRi6TFDbDQSukKTfX26lrINucZHsMFBUwexvXVHT/xoDF
vTzXVF5ZymMA3RWXYNkZvn/TqujZkZtpxc9froqaqSxzkoknaGPe9Ar24El/
hcZ+gfAgkw2HE74MjYvQsbRqvl0JSYTj6snK3CJZqxl35n+reGIM3dWFkuW2
fatH/nLggbHGr4kOt6NCVqlqcRWxnZMOay1r4Y8y4CShFqWBN/ETbNv3+18x
46yVaQUqEo6zx+BrYHKW3RLQuJY8GHu+/PoKo3fVoWcB9E7S4FrC2cL96L0x
F9zhRvWStahMK7As1z42vHV09N7NgO8pLlJc4hVimVJQcQefzk9l44HtZBIR
3BKbSOCF5zmNo4PCsyPj0bkVv4VY014mOQ21oh0N1gMFilnOQ4VAMlnPULbg
RW0nZXZKbKu7LU0/bSncCAJmfIjMmeIa2sXC1+iQIF5ac9YcEh1fWOreug29
QPc7/tAxVyxsJNYYLR1YRwphXmIcrDLWiuwVpJbx5igZ1deMk7FI+roxKWlQ
OmE5wv9BzRymlj6BWtCpw45CQq9sgtY4bV9NPVZyqsoXL47JkpzK7m4Z0oOG
uxdkhua1qzdOH7slonNH14LUphN8q3o+EhOtw2/0w+2nfMgP97+aDW5ROMCo
y9vBrbfqmbeQpOzmvm2HBvGI/JTTaSv/bWlVuS8xz3WKC+wKAgVZNm7pZ3/V
x6WkrmO/mcHX6QyVzVm6NUFPpKe6pLzvqQ5YZK7erihRb0pZXWV7TmVEqSXy
GMAX7FoaKjmqdyvwdqAOMR2XlnnwGLpUIXiUeBZB19N98kFI2gd4SpkMX3Nh
TyEBjGc1NDBorRcpOgltA8dYRVHyQ1VfslyBRm3pv/f5cAbFk5LLo68Gk0bA
jxUeFbamXkVNUn1kmePQ9AxOlaPXDb1I4vfnRE6HPWCrMcYZtXZus5LJSRxK
jZoqozSiYrjDvWdKzsZjJer2jYdijkG4Wo+P+NMjwmspEJl0kRIlhn+Ee/48
U15/dBJsVnbDBVmfBE6KiD1E2eQrtSakI/1nj76YijnG5AGu68i8iJ3QZ8zQ
KcsrTnIaY0vpaiBn1g+ZLxwUjr11L3+IsV5QTNgU9lpnZKUagOS45nltrF9f
0koMlg5QspyU2SR6agUaUvoIURmSXmySEl5JiUeYqKet9q/7hjqg7D7Ty5Fs
IzwcCt0aWLYgoPvwzKrOLRfnQrKIdqeyQlz4FbTZ3WjDqiDDDw0+2RqQJonT
9UrV23WrEJI15OfvsZVoKI2xR/09Y2gZwqyRFJnDz703b9CW8KsnzsvTZiAv
pfTkWQoqcO5/9NGgtT2yX/pEFFaW85X0bWub7bsDjqgjFaWZIm3f00jBmMPe
10zYwklkx+kS1kplJlcHVrd/UIHo9poMnYLp/41rh1JBIkYHYy7+L37c4vj4
MscQ2jCz6+Flc693c6bT/6wkqybkOQa9NExZp08BK4MzRK95jj4oWKfJBlI8
nN+tsYF8pbwMVZ8awJHSRdAz7ZFHfuahPxS8Fsw7fOSE5be3UhlydOxFK3bu
JobC/Vh+41YRt7Vu4i1rg/3307ZjldGofCfvXgBDu8/BNSCN8eYy4d9cyA9o
ipv+Q0TaFDZQftxPfGq6B2Q9s1QaY7QqRkpuKZWVvKBfGygQJ5UibvX81E2R
BhjQJHA75Ta29iQ0Nsje52vZUG8OiI5/BdC3vNme4H/PJt6TyHytsbuZFxpU
wLBoi60Kp+OnetpNvuVFbjE9ee28k6QQs6Q8VMHyMDLFRPGOXItE6q3LHUWO
71ohZ/W2f2Kn08yTebAx/xNibSaz0kHhfLq+JSwKWu0qMbKdv6d7+H5pqiXf
XYU89H2tSKuxRFY7pjXO6KN3vgjkBVEcFSSDIgayaKvju7FnPfjzi9KStluV
Ny9p3QtO802NVqNVjnMxMO5OSU9T3NNRq/UTb5hmItx+LFDEaYOM7PngpEwo
YmXxZnrM/wXlObmxjFwrET0bI65goSFpJNHpnrHtoQv6JpLgsdOfZDIAvQW4
OhvghMUBjm6yOeez5KhIE9pfXXXIllXef4Y4WhdnwyxpgSPQXMbQcp20ZWOn
pcZfaG+g33bgrJ44fsJMsOKJYczA0VcPdU8wm2U71/+vNRCFJTrQfOCeAEpP
jcoM5w5OXvkvAkOKIHM1Ou0iMcuf9ynFGCoi7TIIrOTzJ8+I9+NSk+WmT4s+
WrjhIPU5lFFVcxxkSy9LwEvjBupfGDsb4ubujh1jCSEOf/4pkISlyztdDDAZ
xXLZHk6WYQMDI89lvXkUlr4y/xdYn9gGMJFb9HraRSqISBlcPr0/x1jdX8Sw
IJFIBLc1rxj/int6KpYycA353vJJw8kApCj20NpOtHl8y9jNjIAFs/4deigW
PjiHHfLziqPsfHxE4WqiQ9nUlFLUl5kCCP5Lx0tjUimOL1jF8yzsyCcvc45Q
PFvOmQywRp/F9as+nykrnkZgqLx80dQ8HHBots9u/LP++gfcV+2PfchnWcoQ
VuknlM6GDJPocThjsbfveX0dOY3NFt+eU0M5Lkz4x+N45cpG+1g9Qu720+m5
6kcGUJgqghbH4PkrhWmnOOc+WvZ2/MJDYIZ2LU74DVllo8p2w7uCw+cTdGMf
OYpQrYlDHkTLb7MTqn1CBM7atMBjOj45+v4TQ8XSgbGHgCFTLW/YCouO8lvf
J5NR1k8rSy2jmWi3tOEQyoMl4L3M0xVp+KL2YCgjk2jCzLYvdbHfDUn0vaEl
X+96V8OjsKC2OhYVTsg4W+nFeCwe5ag2nxCaTf6VcSxdBPCVxL75nCqCdjbi
DJuJbLAgzahtRhOlyp0rVckhU99oMvvstdBy11Ly+rAnbhcG/Ic+7Vb/kCKP
HEU3g24T1/kmNoi6DGUAcJJSGBhFsWkqm0lDXKf3A/cl2wvM6TW6D5M3K+Uh
JDsmlY5aWHYQHFDf47USFUmfPZ3Kn/VCS66MnikemdIpR2G+y5GoLgOugMm8
+yQkfJXJXxpcnvPYJEPTsqP6Vt5RA1fYtCDGhmYAw81lGj4SLfYJxcVo/Tco
DaA8sqQKC4mc8XiBswg6hv/HssPNKoONK8M/F57rtIheH/9CO1I/uBIpmfpl
teuZBYlLEglk0ajhlqdXGL71a/XzaHka6MJj51tSgtNnSy7vZUb6vVWhXT1A
Z777GhdWdTeoQ3r/1jjilCMWcjUK8SsYZUuSCpWuy6lSy7UD05ZDcI2nbrQf
Q1YCzlZ5RH04VbfZXQCKaqOYX/OBKx2QtFpkD4n6myy+q9qsylXeEsOXNXhH
e1EliW6Zj4tWRUdn5Oss64QcoUCMvtodry4vgDv3F1IXFc3h04yGuTb+44h1
XLQ9V3J/lOAFIrhtBrfjHrfYS+eEhTDNwlTOdVFprJXEok3/ydhCx+D6hHyd
YTGcq1VuJWDA4B85ExbVtMPweeasuPclHodKJzDq+zD6/3cEfU3mgwpxusb4
B7kp1AHfBgoXhcwrzhb9hg7IbJIeYwZn8kXVZigi5jyXiKyNsyb1DrRe9vyu
Qic4aHAmOpeT4VjJGawiZEgRg8BKezTQM4MI2QDZG44XgbsrOtqsS8g7wvgq
evuaFXzQqYq8Ibwqhbv+OfxsSIAGtVmqpBX8iJ4RG7c7GRCXuxcl2MYdy7ru
vQ3CcCNVSgx3B8vWjHGvvANuNpMg0ESshXqXV1UZilHvXmQWEcKcSZ5ZCWOI
akAQOMXXuYNtmYsyEBOXLcVa1K1v2e983szQDiXSA7GPR/TNKI1jBzQ+8Z1m
E2V8hz/xMp0wTlIoj2SCGLI5sdnP1VufB30RpFmSZFaU9mEKe/8N7+3q2vid
DWAJRtFMuPhTZwW5zxti7ZiSq1msZ08mRb1hdDY3i8lkmgjHVwEv5b50lK8/
1x40RNo1IIb0+I6w8V31D4bBQd9ytxIi40wr0c7vCLKv49h+6wRWUkEgG9/d
9qjfb2MFEaB3o/1QCa424mAqjyBXMpRQkNXAaP43s+heqgSLeyE5NSRD8mIO
6F7/VjwNUv/ls3e45P3nT70hUfgP+XRTbJt3K44m7TVoEAjPDFPyR654ovEO
7sBHF+BcTQi6v/eR04h6s9s2xZEzA1zm4D7jfUUo9UUneTDkbf+ewxeQFxvg
UFSvqYwGjs30fWYgJ+GEHNm31bJ60DYujUmBvaxxa+uusl9NYG5Yj0+hAzti
wWbojwFUbfoQtQjMG4asbAUZ6c1s1jouCX0rx1x4n63bQxcNSiYtxE1jOAQv
FLf2nLO2Fb8YItLcusrXPwS1+qWka/J3H8ZpBHca0nUJOJe1jtrVei70MJF0
QdYsNXX2Yx/rxZjFy0JLgMsh8t+CUwjYi+zzHZ9BRA8sebjc9QlMkAdJxcxi
2X+o/zeytNFLZTQxPLRYtKAZHReZzMZD7ENMSxPVC6P9KyIrP4gaaOoOjXLe
8dwsNdLXiR+OxsvYyYp+AhyMsANg4FLyNF2ogjmhYWzeQ9Lw0qGoRplO1Gxf
YLcQuPD5r/WAaxCUBL0KyAaiiRke7rqjiQlq0xd4sB5eb55Y3XtITbVZko/8
WJsey/zDcA50pbgFKdLHHwudlw4354RTHPEaJRuL/YE7YS8en0skHM3T5esf
PKgxcdq1ML5xgLud0EGZ7pJNPdrl3iay2D3hhPBxUN9ltOKw/GClNeKnV/Rr
QDTRrVrUpIBi+aelvy3Czi6oyiWLaNWKyOLHZQf9kx15urbf17CDN3IE4hy7
jpx3L/GW+b5Ru4voEBF72ApnNJUv9d0PLA7aeeVf6FSiY2asCarLMrJukLgi
bF/cviMu+3RM1m+9p7jkDs/cHQ9nK4bn+hV0yZRsomizNkEFG7Y3bWGF3rBK
t5zYsY8MXeRLtEaptKU4ja69WW1xUctU1tNrN6WNQVyzTM+UT3gVpdGZg7F8
w+65UiRXaomROfhsWkpKMXo/vfXX/oeahOLl6fwNY+yyjud3pUBWw/vzGjyJ
/LxixM+ZeEXWdWQhvHAW5PJKjkJKdvOPB6gpyvlmU9nEtwOfFepCQGyoK/Fq
dqkLZZkWhV85uWqPdvqtStneZ0sbvh4QsYt2Nanu4N9LHCTUcXOulmr1Ij2D
c76kssoHhXwaJOS9lAE+/0AxSEHS79XtzxqgNZXOvYUCtxP7Wlu0Dmv2Wn/j
I+up8yb/ZOw8/eEyo3MT7UGn3kgRGPgG2fqlWABWUX09CH+LJIr3lH+3DJvI
z+qmgV8wr6/kh2WoSmZf5c8j/uqjkHfArfmWxYcvFqDrdg/e/h2leaJRgWGl
9ujNOLqyXC7RQNpVqM2Qs58z9dhJ0vTC3ZyUAygIwralxbrO9l1V+LadoBLI
CKZ3gXgFQ6wKdqefT/+cLQJ6fCecRdYWGS7ntUUf9lZ0BmHxDffZGywhdcqo
/Zs0L+ijwArvtIASgaeDVTvn6/+/MhpPnnrFI+wa3U7zKpmAFpUGQJxC0ox1
ef9fojtupOTqdlq6htPQ1OZ5Z51S/vafqypM67hVjhcMeuqhVPaIcQIOLX10
TEuUSMEcrDbnGtXNZn2ymapsovIhhumBiUYANDXeWd8vYP+kD5PBAyK6km7P
Unl6/i2IvQLNZfdhMWt/tdjunhVCgbAtriDBFvLABXtFGwFCF5nLS4eMoym7
E4nozYySDahXbVx9G2tlaUMjTumILy/cF/DN5RVebXTeWUBQ48D0wpjuAUAk
l6AYcSLRiXcDTc5/Ot8Kas0FoBn/baDcIrghVyTCDX8Wg04UXYaQv+mD0LC9
qyVXfFhtNHPJfVtNIH2QDNgxjGCU/flg3z4spBgXaoSIPz39LwO3T0SHpn6s
grXOZLxNfI35U+Z91FTiePWUm02fPd1wXBsyYcooSGSe4qBuKSmlrVdyzwnd
OSG3OvTi23KmQRUHgTcSIV8oXeJOl/eimmL0jm+eiESnzCEDBQmnM7Tlwv1c
FzSpZPNjk2bE5/vEh//6Xf390LZr36Bg5CAwRVGFio6G9lpMUFOyWBNWp6KY
g5sG1qFsEoJZ7E3VG5OlmyKanuRGnY0tjot2hjuHIr3qy2AGQzYNJOCk0l/3
meoSiYG67xTe/pQjnVYedpunMwSQBADfqEf1e2G9EEfpl/ziCjbQJP+Sr2Ti
4y2HFHtli4eqWTFusd4xzqidBfYLAvTGfH7DXYAsR74fCuG+GfXzBc6QndBU
JlMkC3jTDYpWj4rjL6sm+jq1A+zyN+eUzMKfDfXJCKbUDYw4SkOB4xd9OrN0
t/ZMUiaFDuaKYaj8gci/QfxWQ03iLzqAq3sAmKEfTYbWS5NcgtWR6gXg8gwf
gvovUSHF+I8AU5x+OpMsSA5lKH8GrQIA+7TB8mILz5ziNQUxeHY2zBm68Bc1
BNo10E+gbcd4CM9qZW1Uxth0xLhjfrc3UcGtoD0eH/IvaJL6TAsluldbFewI
p9unDdYSHcUAbttKf3BZtpaHmJYNBdCbtScvI9rQar+3imQvt7kU8AE5MTlb
ok5fjra7cMheDD5+XFufYIT9YEidl+ErA3S2rGoD7tYKCuasuEB2GYdq/12d
2aCfl8o7q4jcF759pNTvw2rbKry3/VQ9RPKeqFaDik/cutBndoLBkl06bahn
N+WMHbNa9C5Z3zfx0/j2gzYXUPPmN7xANsCyioBIqqtcKG5sFQY98zDXTfIu
AKF3+y76KeuAlZzA+e/KiVZ+PHGVWwk3Y1ajGn312eUbvpQ1KFgm+TwjpT3I
m364sw0W8um7FQQNV2OT7glQcXxRhDw3OrhcuYWj6ZmXqDNX90Ngk4dyqN+1
kPxuCVB+fzH8t7ID2xJztjqBajgLu2h+a0iezEqQIwxFm4qTSe5+61iEAxqO
UVPGNEXrTMey6xbNTWO4igHkEYtyr/KL8ZezlRmT7zvDH3Re/cHXl+Zu7NZj
BoYDFrJ+VngLm6propD9a78kknn89kzJVsSiU34iOjAhtQCywhycuBl65nTU
xMy3PEmZlltqU6ZE4KOKB+ucnMVX34WuiUOkOKyvI9w1WeVAJRA+P/7wA89v
wO2N56C+hfLVRnDTcUFyCy90oL/OEwOTccC/QK8Qf5r3q+apTLO9Ab8Z7AQr
0Go5PN2kOsZ4zO82yMftSwVv0YzT7MIZTM37TDKhdDksFDYvOQnisvv31E/n
KdJB9w37cka15YiIr4eJ+hdtlJGWfhTR77sceTKO+w6emOxNlh6bqBq4FzOC
aZLLGnEhtYfN8n6U0q+aXOtAx0hNGCSq8idvOm51p/OMHXN8J1SQqJ1BLG2P
HUWgL4jCJSOUY4Vlv+KBC7IlOOsXealBnn6iKiq08ZFYXIFsxOSooTFIRxKK
QwX3EvSrRxvCSrzcNm1gt9Qgcpjv6MldfNZtqK7Sjnz4qvvM6KGPXpXA0xQ1
rfCnW6eOKOR/mAdLJzbV4jD8K345eYAHIoKZyZDORONB0kGjaFFzOzpdBOl+
w3iRvAVIAHWczk58vTtMR0Pt6GioOIAH6k9TR3MefUlVZ9TpKs6PYupvwTdl
4lVcivTWGDvR0MjELI4H3SHEf+NRgutqHlN06dKU+B7Ux5cop+ZWRLYc9jar
7/P3yun4aJqnrIaEQhZf5sHJlwrAbLbXHl0UKBjQr90b3YYOiffsqbabNvEp
+fdWs1vynKrpYWsPR43CeA5qdbQ5pj1rGEHBrDpOkPLp3P/IKW2BXuQ9roDW
0ugnYlQaHKWWa/epLE+VhgQFZN6YZ84JMcTJnQW6unXyKTid16+5oWLEsTGz
XmSo8L4RKwDlYslQ710vc31BZUzeEShl9qcGHZ1ZkdFyLJhgG6utwXZ6dTzi
uyyhSRtbKtqp9ygmr5JSPpS0/2OjO7Btnu41frsI3RLbPwthS8p5/jTbPp8X
XQW9CkDpat/NNxmBa+hj4Oe3gEAekbBhymn/VCsymVdgjC3jvjYMCn2iILWn
UV5Uge/Mg/IyGcCUugOMldCNn3t3aZZ2B7Vvo8y3OSNqRdE3+o4f6wuEcRoW
68Hr42//x8mjtNfXvMxdy513DqjeSpzD5mPDApxe0GyhvE5njRE5fd+TVQdN
RPl4wyaFl6U63cjm2YbiW76+aFFSIZxEXxBJhkTiIwMk5qOrN9H3rZLZYw7o
ckOMveYOyG3HooAWeKXA/hJEWFM3orOtQYXCh39audU6OdBNer4eLV4JLtxV
BdnENyTRVazSLNOb/EEt6HEeQtmFIItqxMW4J1mvH/ghCxym5dk6kniFZw9k
5+BBDzwIc7n6R51GLKZ3gou44dvHTBg9vvpyPkHDrUa4xicavGR8E+fxAamu
/7GD21ZLoKoPsmCAs4lgy04yK0g4BJhBrUA1wd47pdfCyCY4xviY5j1UPMbT
JjCbEQlDkVVOfp0BDptYuM46xh9Z10BWi/JNYSK9aFszS2QQY3zHZe7fY8Ek
4CYxJNU9YyFRutRcBZ/rrx8WP/vXDqvxWPqDia+29OEF2DUeLb8PO2Ui39NC
p/83gCKFeewfMgSOSuCnt2sqxKIOBzhbBVfG8qOzHZ/uC6fBHx4C5p/N6gfY
KKLZIOvRAXtRGxMEqWx9Sfbana0Wx2DUNJ8FhJ5u9kj9tuplLmvRCfX9inWY
dyM+TWsdegs3THhG7hTnu1V8rlDqviKSDqbVMAqHiBPBWzshSRwZgxzBU5hG
9kE8VKUnhJNEdacBaschOvsjuQPqp/OcvlUose/WQuZRBh0fu0B/w8yj/jLJ
k5MOgaBFE7zVW4yWeMZXKflEOx8rifFGvYsThg/4UvC2CnjA0YwtHJoZuwvW
Ka5YZr33r74uArwZSEzBH53wGFgs8uzOcFv1qezw4bs9w3aT6ZbVZJMJEVbX
WQm4ddnmr+8Jy2XNSq47vLOhZfoJaU3sL+gbO8jr3WU1W9dyrZG7+qal5F9I
4lQcXkx80JjQ+po+EA2nV6K8LHcMRtkd+X9WIOZlld0x51elSDH5nOXz8txZ
vhAwEVQhSG02YIDQoJVN6TCPiP620WihNy0rClJJGLtfQYdnaVj1e4im5YYu
5mOLI900ujZxZkiwURvyj3dMQE+Wdpuz5FMBXlM/ywXnuElIwN2imHf6Pk5d
M0Ol903nw5dfIcbTYAM8klSfaaxNKvPYV5fcN7/2xV8oRjv574unwOr395Lw
+vWbT+/PcqRKcJJcywA1SYqNDJxtbpEThratyiyLwkQ6DY9tXzXjx8l9984U
Tu+e09pBm7I6WUD966lZ9TZUuq1crBK+32cHYfFe46bjeGMimaL6+FY4OYM2
Qb0VjKgHKfGjlqs4hy89lozX2e0qQNtc+Yt6X99SSDnw2jeHLOPXZFWetX07
mzg3u9s0hn0OqICrnetmHxpKrA7F457fMEn29pEKkxOveQm1V9caCRBw4Wa4
o3TbWCSSA7XfbUbjfrRw3ReKPGDXVhTRDcl6Qe2SlFXbn0gaeA34QHo87WMB
gr5mRkyycWhQ9zIOkvM+m5phi1CLMK7dy/Vk1UF/qyk/Qv+2vXohwL5OAEbY
TUVDF/flmg2hNnwqqBDZgPqzte87S8ckXdgGMgzYFOHBc+FSyLXdywjTJRby
0eh7U1xk6MboNxk9Opjcr4rsAU0VTr3bYG7bDWz+1am7EKwgjTdStSob2ZhH
QbtfX9EK+S5bcWB8lpmeyAh2QbIf2klebhf53+TqN/ddo9QbAlJdmI2iwuer
OyzBaisNM9cpozmcSr5RRT4xt4H33QDklHD+rQAemkbW31J3LeRmLlmVVfCP
YL+PtCn45j8/g/31bBIF3D/RI52L849Sr7dwgBXj6/XOlDk2inZ06EXkTBuz
B5iBXF0ypjGtz+87jQKoVRg8w5nUUvX7C3l7xemB1KxzspkMiORnVTNsRFB3
JCyK6YAARXEIlFuOHHo1rKrlQQIZIMBIHpBnwn+6llUPdmYHzCIiP/WvVyfW
EjX67tS2NNAy/B3kizOmAYRx/1igGcQMZUZLTWJrz4iadmpKES7G9ZaTPCV8
+MZ95d4EMZhESLkhm5Wt+RK993yeqiNyPh3OjdI5TGJDWKZ0Q9Zu4/26dlDn
2xRiOD9SCNBcV0ZUn/C7X7T9E/yeqkjuRigdVf7wLbiyio77S9HSFEMa4nwq
ZPBeDuhiRgbQNEdkKlEP7BFb4MqRn1lnBw7rKbDwdphPcfB34MUKGjlW69du
cmyGbODK0g7Ou3GL5AZbwKx4+NXKY1r/ht7YEkiG79RbUErNJ2X7dG5my0sJ
iUunKLfokRzMTs6grmy0OAutmr/20b2yjIZh5ps0lolfGpn4IODPicLPMskc
JLvBasneI7QMihtDT5ELsp49AqTdaA90h/I6io5ZUHpN96CQkC4eWfjTxM5X
dVsizXtewZ0Jfwf46HotiyzJsfxbCw9sV2TWPhmduMm3JNP6uVQosIrrGnte
70IrkPRNCCTinPgUWMxmab2xwUxh9olEPVTKZ+cXXt/K3cvxoVsFndi6iofx
nA13BAWkF8Iw+frblphPaYoNY6u3l34z+7AIrF5RBeD7nkOzaN4WeKpoRvv6
e3zHRNth/X4vlwEjbD/IMtX9dvnkVNCEXhna2Rmf4mAma2rUFKeUoIxsOWep
QW3g2Gpp8XZ753SXQBVchzsRx+LcDXNLwo30oqEz0R+o6VQS3/FnFywStCF7
vj2H5iZOJ3W70iFa9IjGuaPnN6X8tbO4ha8zWN2baQ2HDSBVEss1AXB1D2XY
ANAFUQI5d+yOvQMHT5IQTvaZq8jUpvt81sVkewD4fmMqUGgQk8KeLRYW/u/s
ILYWG3YaFwomGSNmetzJ7JD9NgcAkbo75G8qttESU5a9ExquZcNgAJn81ccQ
R27potcG6uT2bEkeZKY6bUrldzimxAFIiAW73Krs75CIN0xLnrpvDfMfCPV1
nEo7UfT/4EOvdufQe2aPrA/4gbVQq8Z/CgzNJ3NEv9figSFIcrN18Wi2mtFy
NCSURo4DSNiLAxZY6b9kQYq8lXsQ4FAbjPuY1JOo0rY1y/gC2J4XEpl6bCDW
sYWhoImTkt94D6a6BSxQjOaTwqM3DM9QW+fu/4NPTIIOVcwPMbRzeI5qgy1w
nqkPY6PmECS2H+wz1KdIVT3S9oCIBZtjU8V47hCbptcE1oLMP49CU7+9fmbw
a5iL1MMsOqguDfcjUtzQtLYvuHhWmBbNY5Gre4ONbIHt2EKgW7d2LH/vts5S
2WkLdQPxaoNhyxLYJTTLXt53EDY+p5joWJkincdcYRPXBcj3xnkv6RHS4P76
X3abMhtnC1mPDVAwvK3u74B0n0V992z3425R2IG1lcYe+7z6tsK9uTwuqsRI
t+KawENukKYAPMQ+EaM48ancwaF/fgxt5aTxn8KTn9JRZvtbfbyE9UArUENx
8jX2kqlhK8TSfr6RVwadHd8LzW4MuxkazOtSBpV53haOqA+F6nq1EsjSJgXF
FhVubbNp+nQtLKeNdKpctOzBpBhEnUXrC2LvESIlBap1qUEhyBLf17B71bIV
osOFRfn8+pjIO+rTo0JlyDKw+as9Zcxz7mhYqyUO9dRp43Q+J7CeqqAkZEtd
ALfpNZl17maeCDGYnpQGkRdsV4ZZEs42w3GUYue2Rurr6wIKf/MPhw75S+wI
lOm6DdgjMY/gU55C/Wrge/+GvLfCvbllVqd+9PdtUOJo3aHRLDMTgdcWY+qP
T9ZdGuxQBZF3/p+rlH/DkbBDVefR2Hj8rKLb0cHjFA2+rBfvYbUkSVdsrGFe
aSNp4AkqtUcSqS77hAPhg5rG1/01Hvqt/G0Iu2/4sb5niTfhrzzsQDITrx5x
Z7DZ/S6cg8ZikougpHlgC3XyXLUmcc9rMK6NgybuXs7SrcBR9FyIPVxd0fkS
odxWcbM/7YnG5biqZuT2dMOlYpD4UDCblUwPQmWnjAbEfdDUmgvWs7TnAYkP
hIR7YiW+RjCzpd784kW0U/4QNlkP4KKr5QBv5XkOKdXFSLMVQLHv8KhJlcMy
4Zod6mK29gqTaD0OIh34NY27XlL57AW5ZYB6JWMshsRSR4i+AzRf+uRpxLKo
7GS6RnHtT7WU+41B6pqkDNPRhDTW17EdC45m8nEc9L2khKe8+RjY+nFxghcZ
nr60yLJgRe2XwEO6oUeB7Ze7hCYaq/e8G0n8jrGPrhm0DkC4pTRqsx3o6EtH
ykD55ju0EKaXC2ATeDp6ZQ7hnO7ugSSVMweM7m+dpj0KhxbZIHCreZTQo0rD
fAtoYB0Mmqtar5fghkL5cNX24ijMGVpAG+BHnmFv+oKYqc706pa0LjVslYNS
ZOf6CHNm7AG78qpZtIg1kDm184z5i6J7eR3X+OqMpXOv2sc2Rk4M10b8yhkW
EQU5iQCq0NyJbFXOE8ix554ZVkMPkwPbmy5IGM38JdWgcU4Tt19tzKzG7Ogu
LEM4K2LEh0Gh43CuM92I5E18Z/YNNZILYQeW6v7LypYRgR/ZXtZKo9sdELdV
wFCR2m52+ark46RXnPk99TCAeHfK2h8zYMf5dCvNJXgUbpaGzKar+L+eMjqW
gdEu3OVb2cYsj2/8vak0rwPaV7SynkRD7cjdEDsPA8c3vPBXsYXfGbOCOdXn
cIenF3qHxEVYblkPT8qAmuFi6JK78NLfenc8gAaHmXGidw6ZREDdVdU9b34z
QtOq/aY3zUdIGnclB4qap5J23Jjr1nXJG+cRcqeu0Cv7NXSLECFWK4gzmW6k
wxR/qCGpGTDD5NL0xiV9gkIuE4a57o+7P1ZhXLtN5zi86Urxt9LOg2ml6jDh
KgC+OfjlVgQJifjRyyJH7dFZHa4ILANtQwbr681r+MH7DY/CMYDlgFE59fsx
k4NTxkc1hwcPJsK4tWkvISur1HLihuLOXi2zW0DgqzL0hxMle0Ix1mQDSxRh
ly0ntCXdM0z/7M9c0FaVSdw1ToKlOo1KNGrSPZTNvLX99Af8aZOXnd5rVXjj
8bhGroobjHxm0TaOucddy+gPqlsf5EV4Aom64+EFgwxWj/yyEMVPghKODwlh
yn6AiEezGeQqUsU1rg5GaOkESRp0v8LfFjRtidHizrOAKFsPU/KxQyEZ4IUc
erBSzs2RqhdTC24GS1iTTtSLzQ6dacobI+UJik+bx7Ku0l4lLeRHHSF1z3B9
Bd29BxmltpIDTS4X39+ALob1KDjwKzUQR6ZjOIKqON9OWgSbwXutRt6IVxuj
6Pyc2ueQNwUIW1vZtKE61kt4cSdb57gwvbcD+jFtubjp+O7e3R8CDjrtd+yD
KiSPygnQnRcWKWm4l9pi3NqRCPa2l3iB4dmkPpndD7y3IPWlXBjn1iQ1MhEY
uP/IAfFXJ9csSqhz1bMgij99oXCUYqVsGsMb/GXvyn7ZMrGebRJYsv1cJMzE
VNGWMH1N1jqszd2xVYDfSmXjoUonBe8Yryw/30EdT4wb00Q2dZSDE2K/NZbb
SFNc9vWJ9Psfn0taJEyvLUw47xkv/uLf2CqBf2Ex1YLm1i3kEkMMK0jldHzv
iMNx6rVfzhtZ0DPnYGtWsgcnATP4M1rfszx+xClisEMNyzNmVho4skyACvrf
31tYKvDJQzgoYf9xEzyHs60N/FtiYNaNWs4oOjkNtopIqR0TpBIjSaFkvU6o
uDr/zQYtfbaOu2yjvCRJgHu3d3Voi6dHiLigN6OU7woSWxzjT1ucpQsHCyr9
7H7cjwgk+wZ5u84/2zGPwNjjUzDNeWfJ5Kc/BQUbhtWsoxQRXhuT7UDvVP7g
6fRSYIQdDI6gIzucZ0v2WxTHIwtW/lLu1Dnr3d4P0MI3RKnlKtJbPf/2oEko
2m09bArPTrNrITI2fCx0H2zW1Ag2PLghiEsRfR1ZFNKwgmecA2hXmTb/isa5
xbyhOlTWIygbCpZOEn/wA5McWwTesaG0eZvyoVh+QZijiyGF6Pit1eavjiEy
xJqxD2ZKOPNu2ryOohbX+qhrcTFSCrrzvguZatdF3dCKDfEj+hK4f9pMhE+T
XPa1y+q3XUrT70Dts2hfw+vuBJqBlpvi7FF/tcn399KPyv0EGYcvEJ4qn/UF
RKG34I/lFTalDln5DHRWRLUCYBPdscU83jZS0ISk/ui28UzawHYY4H0fFWiB
N+oyKjmgXaXqQCwsWR5j5/qihRwJxu7FX3jVEZxyX59eJcESHH4PWwyAzy42
BdbIYjog1Q4kdUApmKnZIgfUX3Q1w9BdfRlip2FT5PK/1nERE8kQhCwFx6xa
8DQxwFGfdaM1rApI44JsOaNYZDsuzKKCvs5ZZdlyrSZbKqESrWJ7RRjHrVQ5
kjJDc67s6pJPZJgacMPCNHZvycmmFo+R5dCmIPcUXpbO0XYpdtbS3Ch17kaa
W9pMfzXTG8rg9nsg6ZiwIZsONpMDtwmhl+BhFWxCa20ZWNqAVqhLX/jjTQ0E
Ee9MKOKpEuhlk0V8/oaQNulGPdQ9MIdvs/1BhAEc37XxwRLfkDR116tGLrz3
BDwzj2TYMP5pAYr1gfxpfnbl2UBtgPJObL84Np5toWXLMnXuJ7+Xw6lsuC5r
iF2z+RPbsu9xwIMIua8ll+rhV0bqw3VQuToHxL7ZHvB0hFiQa3/wmtjPr727
zfAuyGGX1BvW5Uvs3SIu2tsvqHiSxO7bRxGjK2m5TKp8ZDbhcxThLSw6/hzU
BVd1cZqGhZue5pC+fnoxHPEx52j2mUnu862d4AJ3ZLZa99roQt9C/rYE9IQI
Gg5LOIQSIeOj+IvilrMRFBDzjDY99NKjvY+tpmNcQSC+gUEwKR3XvwG9Feak
YfjearoNG1HBxw8YtPhOwd10R4ROyKoQKE1WKBvqxK7zo4Qt7AXM8eVJ9Q0I
aBZXrTx+ryjlDGtvDdif5ZxvtjyZwzQHqM31GZMzC3mg2uVCptWagUWhCRPb
UHxPFzS5bP0fdq9dD+pVkXGtactd147fJRl1Unqjcx6LNnojpDUUmxK1OJPT
0O6hDDxoOq/Jz7AWhZiaRTET2V9mwFzICc1cuOssguuq101Mg4bi+X6YOl2t
qB2TQ1lAgTwdjO44iYhCbT0estY5Q6vByPvGWXZIUitL+xB/7SxhKJGlTCMp
7UjMJ317szBwgprpH4f6WofyMvVO2NjVD3zebOGVHtgefWa8S7DMlUkJIwBl
NmRgOTmnOVWyv9FTbLaRELkWPopELpahETvAlAqSbaqI0oiUV0wfhI0g/6Ry
gRG5CdNDxdLse3VtyHVh2mTuWEYPkYFx10kFc1+PzHYJxSS5zDuMNUT9fPe6
sg726/xn6AKelP6RowDge/7t3rvsbsDp+vyHBzfGsahwYQdBUZvtGinDqX4/
BtyC5xIZHspTSujGYnv6dISOVwIYQm03rzj6S5LOONl6sbRuMZObAwuaNsfJ
LTRw2sh/4CQLSqaLd3mGgEuYaaqGLMkHPax+NyKeqAAANp5o7z6LoOm4YDgC
faRk+cklyzqQfc5ySavJhjBWjVaRUP8KWw0D1Y0hWdDrJFTmL8F7mxHb7vcJ
Y7uV6ITUvziYczjGYh3NssvzCpylY67rxzoClT/RyzHkocze5mRQuBVEXDuu
BjQwkAaGcpTdahUzhLuFO1lb6xquu1p2yd8QjwPZb95c4VVRYdkmfPYDkdi1
Qure2B1b2lSyR2/d87OQnc/ayphagieTAi3v1Pv/H9q52MX1S8kSPd2izVrP
t20SCXLchFz6PgcWvmiI3G90S31S/93wEk4nN2tVMk3/ZwDamprTwmGMO3hD
CT0zK161HXKM/imkI1zHgpxLyPpUyOWI6hstSJ42pjHG5WW0eJsKfeYyjVRb
SmeMEVdqi2J1O/A/hWnZDon+GLXWBd/1YHrnxm1vBgBqQobNUhBVGy2b+v3W
qzJAjeQTIENaHvUfYpyXX/VBQDLmAuu30xNP83Fam0IUUmBDAs2vc3LAG5XZ
pwXgdJaLRHFEQm+QqDROdSQlqlPT+f1f8BWFY0PTmsDDtJgj8gG+hohz9Oy8
Fz02Q+08LiOj+nCqaTsnV6TPkEluTOBKx+lVZjNbIEMteYTLgryOiVQoxZ5i
jlYezBku2xoy+zxTihi1n4qBBXGPee9gMYMCMt7UseF8fW3r5C2z6bgDdAni
fiDNCT1rM0emMLs9a8PNy+LxhmXNxjYQTqtSB6/PJU24GCAIKfOG1/jEcxxV
AdUCl3L13E+ppDf7tOyPgfAtUSiKChtD+uc8uX1su38qRNUAORCxm141OOFf
gN2VR3XuBltFm2q0tSLfavomEBm+pzi0Z+H3KO5mZPLVjaL/mj3LxWLGvm2+
pNjIa9Mkwpzi31QDBtEgVFDRe5o1ywNTI5tjg9ab1+IpxFDAfb6cx/xyOLI2
W0m7MA6VOHit/+hqG0mktr/5mOQDIqO7StFgm056SDjEFStGr4H7ROUd3Dh7
qw2jXNIrStjCFX6qwUXDfbkEbraJwcGEE53ZyeeCOZOlJfstOFpQG0ZQNQ3j
avHTxsEsXJr2TciXWFGSfUfbYtWRGZsxVmadLOqhKbd4sXaMG2NtIiSFGaZd
KSOSyeYv5FkJvDrA+qAWmH5SkO4pEyjdnbbp9GSpo7SXXV9s07PXCpZ/PdWz
toVGDt2WsUOTlGE6EUREbtCXQjOlnhCUwsKAfB1TEBfdKf+0wKG0lHdifxmg
M0bS/bDSkqkWMhpo7pucro4bt76dxWjT3RQ0rfaEF1fz+h5ObpfSI/RTn1Xf
6ZSSQiDDZ4LVznPxxpHYafZQRyh7lPqffQMwuKWxvB+PniccbVaQBfS8gFTi
R2bnTCMgH6YheyOKDA1GPEb5K/zgbO8jX2+a2ORMgheQIU8ESOrb+6g17o5J
9jpQD+agZJ/V5sftl5SHwrcwRjn9m81mmJFFkatl9qvyGfy2PTV1EgLIl+Zv
gCq/KugSv8VYzJdlJpOO782eJDyuWVVq+y0SLybrvaa9dwk3/uRJR8SpOcya
puVaYQMBumeVZRJx3fe4RY7Bkdl11zLx1/OaeeMErN0vkp9HmQSmxaEwvZVg
eejS9trwVFa+l3H6iOP2jNYRYQMTVyoSFXkfaHq6KadQDm2c1pe2UZYMXYVr
1/ZYPlawc+PZhbvcmQ0s9l3qmWftFjjCt+ivxJffGbwa6rn3I/XACGCk9k8/
XJZB4fiawzcu/AF8OTu17ACACSuX3xPP0gYWaMxpgaTQ73FGMHN0LmYIAOOT
s1XZD6jNRKKG3ygn1fIl/Mj7TIzCSS4/M4CH59E7zc8DflkUBG1s/xA0Yl6H
x423MqUi+dJQvHlpyV+BEWz8SKFZbchmOn3qGI9Tn/+wR/ZnMwvxMm8gHM6c
8l4CgTKsNBjohwI22DjhpsFLpqzo405zovBIHwah4Y9HuuJEq3wjksGsXHDJ
UnNEqdyG7rUqx+Yx3C9s4cfLTdiXBmBWsgtaSJrX/4+syo8e6M0MVG9pHWya
MfVxqpnJgYKwlhVHGGUrNKqGSARiDW3ZIZwRedjFLryQ6X6pcTkWTS5unyyn
mk4ySmYdJy8TPe6YoJzQsqMIZZb3/AfE0fwmLr847zZY/zmd1AOAsJbij4HH
nIkOCXOmH7OI8Y3lSLGD+Y1yCtEY53CAWeOX6+GKtiuM/H4gSLs+/JQwUBoP
pcQ3qIdgbRzHQ6POMQs/RX9P3xBHP7Kt+JA76jBd7ebnM9F5AITch7wNU0Cb
ZjdK/97QtSGzrsmpV85yqB+KSfLxRxxDkQ4Adzbcxce6NHLmP90ZZlZJh+RE
zoAwfOB+/DkB3ycBo+GzzpDfb6xm0EeuB7MPeMcbCdaAkXMTFK7xZZf/Ew2x
xDlTbpyK5uxt+l0YH/UQKPoz7UINLxLcGbYFl0nnM5g1gNxfE6Wm+FzBTAq8
19NKjgmnnsnE4S6s3m4C39VMYSTVvumYvcr/t3HnWQxm6/G7FTOncU7lcAOt
B+32R51xUASYdym2kNZHLJK/Ysout2tWmXp2gdBb1O7fHKJJzbM9iGEIc5Xd
Z3Eja7oLMjkUK103sSOiSrQOre93VfrV92vldar3xlwN8j1iG+WQ6Jgr4op9
OcZ1BZH7vp4tvWk0Y6PNfIF9p3gEqgBd/yarNJKIuwuEg3Bs3u6upk3b21wl
eVkORQW8Bh+NeYZEf3tx2FKX0K5cfIu2YYMjXPmr1B+SVAasA1K/5N176AHt
XLDy7aZO/AiFt7/Q17w+Pi9Cs7JtYxeV72s6gMN5FqZ427G/0PU+0DP3qdLR
A2PyVQzqX2pF6l8uw3gb6+ZwxenwOd5N+nFHHAUzzkr/q0RDswgUtghoyz1N
DePcahj29l6eG4/iPRmuUrtMxITUrvvpN13yRLr88EB+k0XJGjPooTVt1gUD
RYc6VQRTz7f0b/uzZFJiRBOF1s00Km+zMST9glbqB4lONVDYiQB+siVY2eEm
5InEJGfywfodjWJ2lMEmkOGhQubRUqNYHvMPZw5MxFA9n7NkRwOqxeYTUAGv
ZeOxUhjZ17zHScrhqoWPZWtL+foiugWeKWoIoAzqgQa+18Zc2oWm5Kv5EiDY
FSvxsWhyfe25PnGY7GNQXqU1Q7V3brPbQ8BSOWQNyDtKlJEj5oIMqNzIibgh
kbk5kPX8gaNHmYDLQRB/BXgCn+/82eIKIVjqqx23SSWLWXc2T9MJhvV1szJP
cjy3gjxN9ZL1x4oDsVDfStZ9QXuDowg/8Buz/5fEEMctfrGwPdrMeVEIbMfw
0AFoS/NIV1yb9Etcv8Cj+nsjNpQGVoU80HQVMKfhLZrtQMvEuJH8qWRIwD4b
Y+XycFusDpxP9NK5hMVUDRsn5zVTm5dVyIZnNs3oJndlK0MNSX72ciATbZdg
3GI3IIYAKgJhUsNXpwLNyr4/q7iHZbpaGn0QMzCFFEt29K1LbtLD+xJCewWH
Ng+BOYvR9pXujc2RpcsBDff+rz2dXqldxOh4vWb0aq/SLMj3DHMceEQfo7qd
z2juBGJVJ2jv/sRGfWXdufgPP6KW5YIVsT4wP7h8ze+Ly8gCwd50V8yq8fTR
3Js5TPNy6WspTzXMu7gT6jS/KWrRQtPn/yQ6EEt717NQWmtddRdL/rvWsFuz
gHvRwvKD6d0bbFsYBBxRX6ErMSfh8d9CM42uKONvcKia+4AMM3Of9TkaTEAP
6ZDqvyRD0GvoeGXxKFKPbgxb2ujNKZt5EWXPn90kMi2+/45tDui1bM974dco
sMmkjSPFZ6YEWC8JaToY0jkEal5HsBWv8OSVN9gBk2HNCkWr2a6sSMOalwx4
/iDtBkskt45S/PprLGXnd14SQIIu4QlqgYEOHYSvp826WbdKjHeyNMxU+vV1
07jLL9wUh2fuRLO2GUhuFMSZtsjfWg3Ci5k0rzekTBA2/PWALIdtrBaBalvX
FttF8Wk0m/AvvMaqYFLX4HsamNqbYXlZKQQdVU/NoO6p5ToR67dCDhInW6GM
Qs4zV+KyhIZDpNzovkQBQFzQo8LLlL+VEBhMA3z1Fa9W8tf7YrYKmPO+3PEK
IVxIFuy5KKqaWVHNyPLXJEym+rlWfBXbBY/S3smqPz8Gmv/5Ih4YRa3vxOel
oueCL7H5lgLprHvuoUBSzuqZVJecgDvLrMOHB/YqHNykCvUudIjRu6Zyv3pK
ftBgrwts3+dc6StBIiU6omFpKnB7oNCjZl9RUWohAFIG6kfWoLkiyiRZVKlP
zeA06+ccYyc4mGq7tvijeM8tGRRP7lLp9fQ/Rz8zi7DQfOqeBGek4UJFooUh
xBaMW7Y4/cu/AiQraDxkjmSdpDVQ3/BPeC/bHKwKyJYUei3PdYmM7xVDJV4a
vTDb68bvCP1YKxdPSJb+J8duk6EaI/usgHqNBH0TOLBH5vD0qdSvJRlKSBFX
hEiuursmgkRqMFNYmxbtz6Fd+WkijPIg3jIdiD1qT42lTkijDH9Lj3Hd0aX4
ZKz50jS91XwcrldIswGySuD07JoUxTrhQAk/yryGbwiNmwgrgKReSStA1BOq
pyK8ajp3PKIIWyTBY4xue5+2rEbyVEpj4Bl+EaBEJzNFBAJnJBWNXuaPpcO5
eTwR9C4sUygIL86wgOSxygFAKjrvHIv4qrWdPjiOKLGx2hG89ElIFdan/D5m
7By3QL2f+CnH3xVXv8tnSRVj9KmGqoppO8HZXG/AxtH7q8jxiZLzmJh789gX
9oDL4EfLcdEDdNKx7/zweobfgX/dv1hj7hfRaZtVeUkJkI+ZFw279H2eIJng
rMg3jGgdRwIRtvBG2oJr/uU/huYWMImN2ZweGeqmBRSpo8UEzhi0u1knDdvm
qXL8uiUVPAl01d+3EFD5S6kOU2dTBub3ZUVAmBHiUSwuiH5SPkoK2t9oXA1+
gVAXwi5rfi1epNEbQoXI/U+WsVhYUUUUJ/M4tr3VpgrHSrzlabwtrAnX0Umm
11yH0fuejPqZl2QSDegx9UIxGJM3Vix5eu07kRlbYEtxfUqTPtuXPZcagQHQ
9WqZo9NLfFwqv7jOkgzcPhVPZAEYLc8cxD0LejBetwv85LFonWhQxNySDCUl
O1o4ziQ/r6qad3eRR3PnjlxKQLB10aCAdESKiI7jK1b5hpkCtHhZZfVOkib+
UsYm3ul75QtsWgSHRGxMvISXI+QFJObStqcNh0HXuXIJaJw8JfGqAmWGAgLK
zTwHEw+jnH7/tu/Vf6rjdWNYblmXn1LBCc8lm6rtRU8iiQ0ZAtqSeTwfIT0q
wAlriNn/nQcHaIcY3uA2mKfzQuyUrFVVBxwseq65Qt++UyjlSD7RQF9Nxel8
okZ50IgKqF/6Sy3jJqolTmbll4XUwrBfXNiUVKMkFHuTXXAOQ115MvH+mBYJ
KONUKKL5yGnY9L69O4lbdq/0dA4aU9eb+8JdCmhlK3imfBxPn5K4DfH7SEJr
9vRTvdC1B4zJ2V0NdUZ60YSKPH4hJ4HhttHOOfBzvKkiIaUR3JT/KGv7JqK3
0WYEnEDzn1zx1wzPqdI9iVOsfoEi65hoKp/B/3B1xyRFmVJ98WeBMHDnBZZq
yJ1gvF2Rpq0RY4mf8SnGQf4UsdFkot9nY65zwLk2O0Px//7/WwB09Wy+M8bo
hQb2GxvTOIbNBRlAQNbOZkJF757CmUvxx9Z+ieBQrf1kMqdPeClagj71ElB9
9sTv9Zlp1T6972MUp0iSQr1COqi2E0ftFhs6QBCAdictau6omuwA+FrPsn36
H3dmbnm9hn8UFdgllYux1ox7ks94MFEEAVfpEUT3tzRVJKkf5MY0oj9mMq8j
xszCzfqhSY5DZLUun5/DWZ0q9m4xQrMFRB8RQMvZ+AYnQnlUXHLaEemzXCax
AfBkofG82nPN3J/xJ/Xxdqy6AcRCvNsuFiTamR3TuwlU/ATqK4tvvLO9Es4a
9le9fjRHna38nfOWqzTFL1C6VSUjuySLSUV1GyzFl1Nu9YNCU4em3UcSDjcn
VRaTMEUDBTWS9q8ngFfXYqlfanjQfTFnpJN8JOyf5ODnrduX7hDwpMAxG7ol
0C5mrYkyUE78tUGHtbsFiUz6LG1IFsKOQrSuBa7text7CYd6uoSQI9o8blE1
/gF/xwi2aVUinkXXWswLCKwlPMJIZtYj+JGrQCdgLeJJ9++Yz9m7dhfdtoRq
1fJIUonTWsQ/MIB0BbW6LDtlSpRuqfWsTO2U50PHUEfBqT8nvi4gAL5OX1GT
4bNWQZM9iwkJ+GxA8YBijUn9/2eBP0HkTZXHB4IyzbIzCOTsuHHY+QmYqHLY
cRBuUdjQgF80GIikmnpjBSoGc6BaPsWMx60qBqUifozEMjJj78FE+IC2p5lY
b4E9RxHtOVQLw7zLhFgO1boyFgO1h/fE0pR6ENFhYP8FDpAcDXu/Vd6hEKse
8/xYLYaEgbV9lHqmaebahlS14sNCdusz5/GvWvqvD79uWhNVwl0GvLOisTAp
uEM0na2qX4wtdQLZQPKQW+OCqn3NL0Q+Ys2jix1XMaQZRsoTjnXZGvpjgln1
7t/X25/qBbTfweNYil3Zv3eSzBqC9lHNbTt79qMeWY5byD1i0wMxJ5oKA3hD
MSYEB3aSRNxuuH9wNUlJMU7OdEe4nhdO6tmp0osCm1RpkcXp61tvTwqki/Gr
L4mDFn1gf5LBSxT/KvqTnWA2ASSm0Txom+j+OgCkDYUpmdaxQJb1HHBQFLC1
6XuQZPGBl/WPEI6QRiyT0fEtKZxjY3oPF6CXB+tMtsDFP3aSWFkitzXOclaj
D+duQhldryR8yYdWU7xDr9B2HiVGtJ2rZLw7vCf+9jqF3eIYiJyHMNgYFXQd
F7l3mUWT/p5zhGSxv85OiKDW5Oi8kx/U61n42jXtcZiHwYtbJPSND3zKoKzw
WipaWWJb4Aq8zIhLcZS7TlskmtHP1xGYAeHDOsD2cUXOyiP3T+JL7Qs8xbDs
f3CwXUFGXk156XcbWNr3B8F3RF94GaIaYBdTP5E+WkENJmzLaaT9QXhOBcwI
6XheULreaUSff70BGTknonTlOu2DNrK0q1l7x3fp9/n3oTdet99fzPbRUHIr
gVIm96+smIRuaAhFr30UBK2eAav/DXbEgM4+VNHX0IsWlLI1LXeooVDY3hNG
pHK9cjDgE2eQr2PekSfKkgoq8QFqZFNh85qr00dofrB/ITBPB9O4XIoxmgUT
E2wrx/onPmyXSZqJLfzq9+FELpbPUBLNpxyO1pQ6HiEtxrA1XVkycuxh/yaW
4KmmautCMTvQGFzJRzt7pzCLzlLkmBt4vxJx6oikCYOWKX6BqG7JdPQZnm6+
YsUiqRGd7reFCenIy4TE9A5aaxvFyQw7mTqTu2cJlbVmndJ/BMfuSGnUOaJH
iMXRzxmogHtrOYYM+c0tEK7Y5+G2SBdiVABrkQP24O3z82AcOk/SJWmYWqgA
dS2+Dk9ON8NH+I/USttyC1JkxB9imMCeJZddymGFocy6NxHXg94HY5Jg6zPe
PLrA/7zundurjGsHThiahdGX/8v9oyMfLzN/yrd6LvBYUoMqTjY7q/+3A1yx
OPkjxqgkUU6BJA6vjs2JEwUFZUGMDKtYcw4M2lZV9s5ff2z/Xo8nGdNyT9Lz
zfliow6teWHdVijf19CWZITPFpSPFxk2ag+Clg/HWUvLjjd+nrlkkB2GcuZL
S/WJWaWF0fVDq92rOY2Yxd6AB42NaVx0cR7dfIusw92H/tglPey3ZhGymVLG
92XMU5tnzSaPi4PhraGhxcjzkk/zBatt6zHsV1b1wMiLeak98PNrI0KEG65d
dNDcTJUb92wfKwsibWUu9L7Ab9Vm6RZByxuVZKUz8zZuMYhpGqNIHV7qaGFL
t0zTkAtHIMcsVwgsFTTsbwygWMhVVt0SkpHAot01SDlJiPSui58lCMvOB/gg
uC50VUbfJ5TCZDAZrbM+TmlpYnflDh02wlYp9Z6t2v0pPaVV/BWzNBKhCQC5
F6UD6vJDKGFNUAmKOnZoidR9p86+UQgFC+n+/mJxbzDi2+2Rn1MI4C4QM+GH
EBZjlQdR00P+lYNZvgWAOB3IiY/YaE+JAN2O+IfCKnRJuCUCywBRcL+Uu9qE
6W3o395jolYIEuBmsy41YOoaH+yTzw+3LGw5Uc1u8/Niu5WPnFCFdFesnZ7B
vuxLdJ3xUih/Dx51veGFpBH7mOAeEXDYZ8lPYxTx5Hqcv/nx1mjT70piIzdC
vvKBWUnjit11RkuvwsB+WyrpzE2OO9mitf476W2VUn2zsJ3il+mLEX7r/PE2
7CLo9aLJ5zzuTGuXIvdcQ+ariV/8yqVqzmgr2gdHFnQUV90kflltaxwtWgyc
pwH+cgDnH9xht6Y+PPPKVrISlNLSjJl+igREgNB8DLI32c3IHcJjE4qSDzHh
jE6bqN/wzTHihBxPq0ObrFjKd0y/M2C7zzrtaJqGLopNlCAW91dzbINdLODM
J9rwdID6gteAnP+onxpeeh9+fWzNdW3kUUoAa1FGzHXpVZ17n+4CsLsF7wEY
xutdQUnc5g2yoSWvimnjEwbz053TBOhESPHKeFzC1Y7ehNjRePDq/DMc+8M5
ggVkGOr9igWjksmFRT5+BXJk0vMpFVN6YfejxyZdgQFc+vX3LUJfJu+/s3Lo
x6aOD4UA+d+winYo1nrBiJwi3SJ+L4l5E/uE4M4q42ju3oTd7NJTIzgVskZZ
vcMQYIa6qRfjoliDIezrLX2QVqYw9Dz9U8eoFhbctwSC+nyZjuM5vvyX45SM
62xkkpb4Cyt+lCkfuWbjp9qU5ST8q5BAVHOz7HpgAK46n9WHrR+QLX1y/B7o
vOWtGm44GvERx5PXoQ3XUXip7NopZF21BN+k5WhfddaYphxPR9ArjOKmsJhL
F0iGGvqJia1DMauOKwvWomtHiN9Tf8PI7aghpNDReIX814e2oq3KE+2Ud3lR
I3T6v/gvHSwk/GJKS8uHh/WVaDDLCkCUH28JMJ9PYVvUQf1s8yaUvtQrGlhk
yg3v8JXI7CAtoyno83laOsKZkhYijoCcQveNrGdKTIlNPZwbjxPVoPQdBO0x
WStLvOtgp1oPfv3NcWDygH1LoEJUkgF7bPKkh7a5aEP6rZHwA1rOcwr/6+2a
aboRwhypRbP9R+pTZjuTqnrbNjwM9VghmX9IeasL8gJEZ7b4oJhrD3qztpPq
1U5dW8W7XTLV7mgI7xa3e+UmcCMlenJ/KkVrOlL6sweuAq376TF+6/sQGnum
wLcv34lAsKlRAkKB+gU+tB8HEVOUjtZUCXeKDKEAcY+/PPHqSP8LeZqDNy2I
EDYKJF+hiIWkWpj/hWjH0aZAASZ+IFu+RBJwiDz53FcnxjkiLoSbVw3MdQut
Yxk91v8yZFL5fYMghP9Q+EqFADILY5PxOwskpSZz+QGvxMccA0ObG2qTLnZH
ucgAmQpFpVdegm8su2igYesDPC5vPvxGaj38VZauXfp/J9hyKC4rd0fh5zZi
m1qkGJgHeyenQ+2UGGBM2cyHGKPBcIoMZhPGAo2EuWnXxXuYlxUEkErAnxlI
KYq6PJ6Ocw7da3v7BZwWgt6XjPoE0Nz7pokt9bx9CReV16GZKLD+T5ej3OEh
70Z9xNBaYIFUCGHvAo4DIT5OflNLI6z9CnnjsFo7+XGvmvYVYaaKv6tvyMFx
nB+RrIZSwW+0uRYxMZeyCGhpIyAyDM4gl3YMxfKhurP3T5f9QQM5vNnOij4r
zMasTg22MZUK0gDfYsq/yl4nugW3Ew0P7xls2u4mCWHjqeEfeLj8FHYPcv5x
4RJ6D9Db0NOHQC4rn7IVrPk1opxIVG8Wh848LRJjsfp0toDbAJ3J/lxGmtAa
lrykWljFqNygsxKI1R66xgmfAbGJIpVuo2k7v6dYaNHw7H68Gfft+g55iZvF
8dEoFEykEPKzkQOklvhbIcL6ISToQgfWSKXSzpSm6HBZdzk/AV+P39TxWTyB
BX+7uNNjiL0W/7X7ndqenMudtlopm5160jGh2xNhlaeZmhJC3ZDxo3bRs1Xj
DE1tjMz1TO7g1BoG6y0KQcid8Xj8UyfLiTJHApBArRSVJAVDsDf9azOqWunk
L0J0RtIkdLSuHo4mFTgTj4LrHeMk4JR5oJktaK5zRClz9fG235EmYUQCS1nG
z7CsVmgN22TtuSCSWNa/n3pYCn2y4TVyYLw00agAoj59QkbwPg6As/tz38BK
VgyJXL82SECDBSVn2uL2U04ahz0PiaoXXbzUVJ/hSC9yk2tUI6B0P07M1o6f
HCRprrRtxaL65nGOHB+wMZ5c/1ZrBA+Jx6uc6dvZtRyxVUWaNNR7LUyUOQVy
FjoRKY+Xa85FrBMXxKUFHzKCJazich6kccCrP5WFLo8nSayQRdTLFe5lBFi0
iE6fib0wJIK8jhhzSs9ObTvUg0EZlJeD8jxtAR3cqP85oTZlpjhXx6q/BnrD
Q693IEvtemFKTxprK2l5l/E8YBAXwJaTndaLClSx97NoOQR4rQMjBqtXaIus
LlfA5TGirBsYZoKClmTZ0BQhbV1uQqyrGPN4QJyYWqVg+ZHeQq+NSERYchQK
VbPnKsb5f3RIdABv/FyX7y/oComkpMSKHNeaeF9AN9cVtYKXfC5y+barNSUW
c9D9tWnZdg72o9ibJ7OLjcJapkChOflAwCEj3+AKhF6AaHb0B1lUH7efg3cv
6RmEBqDwMqq5ZS0hq0oAwo8AtAekzLUT4jUK174JSpkHrYUvNu969AfdVyii
STs+9PkwOoA6bYKMP9z9JDvq2RH6uB2LEGMjJ/pesiaPa01f234j5u31seQ4
mBlprbc5VnbaD/zm66H4EgFUc83UWmeRjE9XL3QWmcAwKGi6CDBMVH01YsVp
qwZWQjkwRSIcSWn+am47sFozMxp5EixmvBC88r3OGJGCngsMeDuZ67lIid9q
lTrd86R9uuXGwTfle7Za2S5HBRNah37p9zmDG3k/KT+u574R/qlMhAliQOyV
1Lisa4+ch8qenE5RZGuk4uQH3zhWMMN9M0vGZyUkwEYzibGZrFNpckm3L/Ya
GVENlNBDexd0alTQtzc6AHY9ih/QozrXI+yV32pe5Rvd9oIl7cqPjPt5viyc
arvnOXi468SUx/2pmDuXBxw5XPCb9s9wTeNeXH5Ipo2I2Dkg02cjaHnbI/ih
4wdLKMowi66oQwUJzaoBDb7VtXL40gyaSjGhn4gI6Ny5DrpGcinJPBlDDzT9
Ss5O4QKQjRkjH5kbd9Za2zla5QZ/xEf/4D8DViXOxg7pTqljP2KnlXdq5tbC
9ULF6rzp/u9U2JzFk0Qje0RCVzYOZejS2mFDsM1IMkZDz+LGFUeUQ+3gMnAp
pllVssowd1RxypxLRir73P1A0B6Z2fNWd+q/o5YLZTMo65oD5KFhZ3PVfwJl
gXZrq2tXoLIiUtbvad7cnnjkhfEahR2Ccy4yllb8PIMQfljFUUQ9uzqiGCmb
pqMdkGOrcpuEW4oO2Tyd4CV2gdLYifnt6DX+fXYk3bXzTH7HJJBp61A7AGWm
yes4R5ZDa/zLrmTmuu32hMPGphogDZZHh6QAZlmjHJTo6Q6+Enq/6hunTeC2
bfbQ04kyfe9704oJl7qWXf+QqF/szUo/WGynwzLtuY5gGjR+YxaZxua4Xevq
b+NkWOvplB1Kl9qcP92TRg/rHUvKku5+9cd2tWAwqnNdIUW8iLeInGZY+QAr
J45FRJlV7sn3EYxwKeJe8ZId8nDDX05AHMNGlB520I5LV/yoKy6gD5Hf55+3
GeDlXU6Z7nAuGs2mb2k5fEktQsPsZeeq5F5iPpwkMzz4jJkXBkRv1BaVLNF7
ooAM0KnsbTcYWFt17cFMMZdmNq0DNha5I/7Pk3nh7jwUiFB0Gm/EvCOkWl0h
BhcUY5+n4JGMaj0/lww/NGw6AyhrR3/WKUw9q7ZuLq6tJqiEXm8UkO1eskT1
ENZ1fli2BRQtC4Mw1omZB49XsUAUimjcJHoZHQmcD1cyEAkxmafFxkOLVxwW
cXfUH8SMlnnum3QjHiCOp9+W/Oe6NOAqfrFFJaslbkAksN2M+4ohNDaAoOjj
+rVGrBX9fgicZ/0TVj9r9t7i/ASbWOMhI486jR+VQGC+NRMMmRkjcn0m+6eR
OO7X5Tp1ADi/WH+u6S/FhSxKkbf82kkeER6sXq3BRHFamWWVwsN37m5Z1IVX
keUTHVpPOqGBBu81dp9ereNc6CsCDmGWy3NYzlvEVm6N4JjIO2f9psK7FsR+
0LdKKfEeMkcwgHCKToxMGSwDSr7ZxOcP4UpTjbndLofPYPq2s2pBpnYf0eEI
GUUShRyZV8U+fetxdGrXieCEzEhNcaVoEQok5B/mHtMtujBFBYskwOTDjl/l
xKUtnqokuzMjFgAfsT4EtuB7o2ujzbYTH6DmAhxrX83p4WQzqj33UZIQWhuR
NLL/7J6LGz8rjQ14muxkevp10qkJ0dcrbGYjQu6m8jWJhZzVxqNJFTBGf+1L
KuMbcP6IzD0r93eBx29mukadhnRcCRZr5fK2toVDh3eEiChRMXBcxM+ivtKi
byv5xW+lEWoGamrzuhdv9OnOXt15V2CoklMPKOO3cHhD5JrR8UypzSFdOMkP
H1UdeYcxX9Vb5h8altefUQuHtZc4Dy+gl5O2QrM199hrW01/GZlSVqAQQuZZ
NnfYmfmEK0STm9FApI++3tu+5ZyV3glnAc5hjK9S5gu40qzJKIxGddx0WYIq
i6G2VP4sAMkM+THpBimR9omRiLXm9W63y65Yi/nNfr7IHTbw+8ZsZJdqCO+j
WMAefg+ba+v62z3/Glp7tO1J/r9QNho/k1fc2whavIvPxi6t7fe1mBw7IZH7
aMMFlXxZ5aFz27lBjWkOpP2wQB3UssUva3MneMJiFYaDIc2VRmWiGsWpNaYT
Q2WwnLHFP4Ta2aSnpoaRgaAWV/+UECGPiFJdQho5YZc9RCSwOI8nEJOBtChG
jbr58EJH2CzgyCY9ifSWN6CLWDPPgFUiHsVvp1d2xuFAxL7ah5FTnVJWQ/2Z
BfkpRXwvXTXnaZdVCZmVPDgmv5a2/QFBnfs9bADMcht+yruTKFF8YmWacbQt
RghupXj/8/hhWMMiDJh4Yu2RNFiJXF2U46BfResFCkSMidgU0QNQ77jaM6I6
/NUObaHKash8V2ph+ODuY2SoBrO+vgL62xGP8hkm2mmnnUf5FqzMsQEAHggG
RMCad46i+NHmp9vEnnUJ+7i/P0s4C6TJnZRhI9XcDMXLYWd0V7PN0nph7x+x
u4Su6tKVxaA1oGIQj46nVNVeUARaJpm7EcVvFGCF7W4rfnH3HKgdV5fe2Qrx
mUPsyYyJ9+W8ZO1Vjb/29zQGUPjVOn8MUmNfENPPoLHqvf9UaeNXzg3Jl9gB
dCmOw/gK9PbdZ9inTAjeR25Ct7nCcGaoK4oSjSZQ/2jGe15jpUUwm9X+V4MT
7cZFUChPO11eQi4BcrxXbbrPH+SamSh1TSg6vJRes9U10FfS4+91uJFJSjui
CHpM/mu8A2uzym93arB95Ph6Tdhj4vYXf9LEK0+ddfgbCHRWo6DtkBZPjWNa
YfuS6IBZUs77FJg3ocmLhTAQh7IpIKh9UKPVJyLRZLNvXHRDgiZAepx/WUm8
FikFvE+iluyRyJdfcYiM4kpNzRf6H+b00YzlifgUyU7TB45hEJ8pb9HqiPuC
nSkewLXrmRZ/A+IaFGOc3dJ8E03ynhhubHC+nFUfmQbuTlQ1bZDhjmxVv/9p
OG0qALJas921DBGsM2HMD0ksCl1eM7GQRvN0pSRoN3sQfo+YNU+w/0xjwjl+
hwbh15KxVW/2d3SDH1B8EkWIWawxp61Q1y3dSinubpwDyF0CCiJP08O/obC3
sz24cg9AOLLcADHI03TUcOJ+I4932dCPcH8gJzYm4Pc4OjMc2WUtoYh0I/m7
2Njq1B8XXIhPyoghqzBc1DqoeTqSv8zsFaXVNCS8Kim+c2hLsaNOMruAfGoe
inSQD1Z2cv/VHXnu0PWTcgNGVu/wFmh9YUO6pjmo4tPpJfskv+7j5JF1HiaW
N0absCn1d4+aLR8TJUCiwDjH7Z5sM+cXttitt252RC6ZhyQn9ROBfZ1CwCTD
tOphhMmWflLswivfq7smAaBYflS+ezHUsHbMfCIy9F8WNqgvbBv0PNCpK4ww
n2wGFPSOyYi0PSb6FnfcGm7MW29/jYVHbNvhHH+hmb9p4Hjuz/HJkJA2FEmn
cYnP+R6E3WdA4eeklBl5TVuLi/AOsT4RSXbZN2gpFvPVrLV6ACGwesPLccpB
pAEHWc+PGnbvejqhohCJyNO+xRdZ6mprbwD1aL3HWAdE+D1ybbAO2rin/6lH
GeJbmWgA4gm/jpm0jbEf8vo7nuBnxT0hiw8LYq/0KJQ0esno78wknqjLcJcW
iEoXPN3jQBC3uK8ECZZwPow1bGrgcoP33SWu9iEo5lxrKmetMVdQQcz4uOQM
nNDQwaduLC3inPbqAy2G1jpamImEWKQ5dRsbyWreYDCOe3ZOnkQCfW5LWFnK
gEZgOZV1qMOyxnkagZKjGLlzyt6DSY15SJtEBNQcCQ7kbFLjLAsxobyCnVT4
uMzmGSMXWYXhBJipvEan3+WNtLqoozv6TsOoNkBZysxJHEyiOa+HtcZdF1D7
v5Z7A/Y4XPGkayhrKcii9nf600n+P1uNkY65LsrPsr1FUR99Xhh09AHDj3gv
TqFizqd1vV9pYzRtZnB4mnEhxikU2dmDRLF2gt/gT4YN8qGO4ca+x2sPtBxZ
O0B02wCtRQavX8rbstctDik/ylr3BrP6IpqteKjf9SwZS12RaEBn4ufjpdkx
3uowmiaZeeomCmTMNfpr02oC6t1OQl9PVD/YQPH11eHVh2Me4OspNYTnPPBE
JvLLyJbj9ao52GlECghSEktPH2h/1d9Siu3LwHEcqz0m2JUmY+SmYjl7CzIv
wJs01a3AC7ZD/rjtFWQB4UrsEJgW4WJuy9E6fFX2qvv65F+WeuXhDxRFXIjo
1dxMiDXfUjNvRC1OarMXlS78vzOo1VZgmofpCyCPm4X12AF8xZ2vq4IVS3f6
wuxe0eOnNW0d4Ae40bPR7tnO4w8ZA255bg4dJWiwbEXS2hfH2/d/paiak0sL
pRT9ImjvR1eXpkDzuLHJzqyGvS61L1h29TH6sL9LS3kzDxB7KiCN+D95/RJQ
9CxL9uwyZNwKSffmnbJTWVY0D62nEmeOblNUCaOJIi1c9rLv5Nroo1MO8nKD
e7wAwHtvoQfRVb+2TzoX6X0y5eivWEQjoQNehtFz23APdR8iItswlzevCpmN
aGwxtrFlu+7ZDVL+NRG5SHJWvmLYC3GNxun0oWOZoNsNRBstHOBZSvmm9k3j
3GEyuLhjiAdKxRBGCHXTxY2hxWqEo2+w37D8/KzjkvXe0WKJuiu5Dn3pUHxQ
vUvAB3DWzCf1TzlH0dlQPRLikgUgLN8hqEK2LzKs/DrN8pDS8JlOcI4g1RTq
32Ata7NO5IHBnNX3XSscttG7OZ8GKCctliTvHFXhsL1I5KzuvdnFBOCwn/Oe
OewN4FcaNXtnbeI4nWGZFAkBiOMD84UfiXv2jg0oN2dwX27F78Bg3YWh/O2H
uE05bpBoNq8g89L0B5/VlRLBu3R/2mXpWtCHYl2V3WEnrhnYi/J7/89fMaPI
ss+GCYX6wwgzGN8x8UQSIYxJc/TqZ/MoDIPljmZ7zzYqvShruS5eJQYxUW3y
5CLIDDd45Q9Ti0UjWZITSjpFgUkqZhXnv2I/uOvRRO3ixZxzgvHg1loiqQ/j
YIaknhGWcWM7CnZVkLX54GVVighlg3i61IlQ93L+RMrACD8v4FAtQAZjhmgb
ldmlN7m46BcSECW2RIteNY6J48MbMRzM/5VN49m/Y08JAPy2XnuTIE4bIEzW
PNbiUR7Udvl3B1p4mnyjM2NjNTXUJ2JJrgolLi9JIbmueBxb6gaVFjaYD8dH
vx/x5bubIgkVfAHO5tZ8Ll1izLeOjecc1Q8bQwHMmEdQM1unEdHSZ7c2Ji+a
H6fcrG2DhjUjAwwLBSDYd0i+BN0+ZgSyjigrDmueOYhDmPeNSWsWBHtTHdtE
fr3KfltCtb49ZKtdfU/lFbu1E8+Y0he/J+I3PrJSToI8xBg9Np88CI+4F7XK
RUcHNCc86y66TiToX9flWKfWujWKk2JWmciE2OUIKRWEt+UARMFX8x2gldxR
4Ah/UDZwpEoMN7QI3aM9m/7+VszfIoObH7pubjA/4mj1DZef0rginYlOR0wf
dpXZ+2WZeSep/ON424/KC24CuOsZJfCL/xxE08WvhxzA7V3sPYOXuyKErw3K
U/DFnTYQmAaiAM2seaCg5q4OH2J3dWCIhQaKa3PGzyiTGkX61YU6PN9/tCG7
4invprINNnVdTToqgLmD+oI7ol9rJNadYdWau7L7+WJGWKurMb36rb78461n
M3jXcdohMX2F3dXgyQkKc2LuxGHrvQ4SO9HL8YJDTRJbqj3fX9Pg4uwzZzlV
YFcmnzuJEprEoTrYYoIFWBckn+a1H3Twa1TBH3+cHiWZeUE4mitHNPGVrjaw
2XoMgGP6k8Ss8N3eBpuwRRP2WFbcExk87w+qa7LHBPflHbyo1RFVk6k7nfnr
pRCNPDZUOJw2J5Sd3E5AJHkPpM+MIqXyaRfqPdUYvK4tdgEsywro4JJvAJIr
JpBICNUAoUVjcZNumO4k46ZmM5+kWRce2D2iaKsE0Qh0Aj7NzQScfbcwB6j4
q345FjFuvETWP1ar4yCg1iqN5Jq8iWB6kyEc/Syi4tomKeUNcOjWGCjvN4Gu
4oJjvL/a9Pu6LrjALsrCWNysIGqw8V2URAh11DSIGp7+Bg1tGlQh6ybTchRN
/UUDOn6WKrBF5anUzh5hUXzKDktXJ0D+0SDeebDhIKdD/rC8N0AaCHVlz8Nz
N6gHnKIB4dXedrfNDD36muPtLDMFffIjD/iKFCNrDeHA69lTM/oqk2JlO96Z
o6khC5zh1nb9yP4G3/z3AQRwWrcZRJY7iO48vzXaVcnq/h3CW/cF6BmdUF2Y
wobGJEm4iLlL2JkBX2zobCvH42Crj5GHNCV4ARVF7urrhXNNNcJ43QkYqCz5
K8yFjEtU53Siy42EDV6g3gDX4Ff+aWXPxT6HRLc+34NaDHDb8UIc/tjhsCQq
yWH2leuaomaHEgFZV8ge9YhiSOvLhJiUKYu19Lc6T6nARKyVDYkgwQ9a4cX1
txjFbiUSoFxPMQyDtczSeMA4mzp7k7agAGLPP7vppXzTaRf50aAvgJoDzIG3
DSOYBfzwu+JyoSwcFg50vjy4/0UWotDTnPLomSHKYTrkgGzUEFq9SmGeAmZc
FajESCyPNM+xiDEyD62C8lS1pg/4ug+GKDyykVfaRDKr8gwz4CybM5ZOjC6i
aGHZoMAR8Odq12JiHNRB787/CH0FP/Q1ZQbRKCtHczhH7oF7oZTubqdPBZjW
PqPQ9H6wbmz7KHuITLVcA7g6YE+2gzkqsTGogdq2v2vgVJFPTBMxw0GJEuIs
5GBY/CBhy1ht1JR79zVzoHHg5K5nGYOak2TqsNhBiQ4L8LuVIpkGQPgeIAUT
rdWuAVbcHpNmWRiWiH8sSaObaAWNBzF3g7AxLrBFSTcUoAkN62fX/nVtDP2+
e/P6278e8l5YDnWom7Qq4kRMyodbcXSIRejkqqxgsnYK1T+0ZU+VePeGDtjG
763lQF1T0r19eTGZtO3tqG+qrjCM1h2CdFNDXVuGry36BSYMbdiJKY74OruT
16iSIsxOyma+kBPBWlU8i7ZsVi/Ty9rhjCqub747NL8v5IKQ4V5lLNZCAeUE
H0Tw/VSdlRWhsQg776vnuEFVuKMH7+tbNkM3O/U9klMSo6UWSeRml/CiC78m
ksuTq87cDRaImE0hpkgwe9wnqNDh7UGl/+QLUMWMuWUmp0Vj4gz/tai0u9fk
fALZ3k8PNWLcOCeJLS1zPoKguAUQlrFKic1uqaXgak0eJBoa99B97NSRQd75
K9LcDQtb6FtZJpHoIoHoj35/OCKIfc5J3EGCB+5de5XEseYhSVToxI4cTb0z
zK6/H/25PuOeUSmM0kdPevBSt0y/IorfyMudpiQQTfCpT/vXLf7firdGzkZy
SH/kiVu7VnLuZnrVTwcxEi5/V/NulA+0lX48HiuqI7rVE/5rCcNQE3es+WYm
b0YYaxbeVxdfj9zAPxvmwNruIhKNxJ9uYcR3CO6LlThY+eZkSl69GDKPYEg2
DCN1HWoaYIoKkpbam7y1QTv4m+ye2MCYUNdpi2P9J/GZ8KqVtCU1NWjTv+Nk
R5ZY9/qRtSWu+jKKWhhfhP0hKmbmYVxa5iw6F/manwBNKjCarg39GIPuMlvu
fB/Ibs3DDLuppx7UUfBzDIWQQ5YTCvCXoWg4zLXzuyO3HO7LoiAGNYr71ILe
Pv++yViihdotWEv09KuHuHApYY18M3AsfxoeqXz7NNoXx+d8zdU3KZstot16
1TOTU8Zd6yWioCacI9SefMhEqFrrYE6hIqosqycKEW+8QndfyiBnyPgXtBIk
EUS8C5n8lDTFnrvtkCFcmxll07jGC0M4n9WE/5XgxSPT2p5877k1d2FkgMsD
vOBmYvPyOy2i/KUL8/gTP9kZ4cuIjK31bcQwl2QdTb85CfvpJe2eUJqiZTCy
uNvNSjGj2+bIqJSL8iHkbij++juUjgdunCt4z0GUV3XBHW+xkxfIKCp9T/F/
iCzalRZy47uURH9RBbrZl4HHdqNy8bZzAu0CHOb44aFjBylVoC94/EDa+qsV
fTTKf9y+q9/RaJIbOpPYfh4FY499CMdC5d4FhK1022XEdVuCRiRY0PZnOaif
rjla3ZmekXmYqO8cIRfEb7ySjxceBHob+JeD7Zi4n7e7/cQDBBhWLHg6nSN+
E2lnmgcE/7JPgqg0RapwmvczRqesHOnxFsbhoLCBR824E2tlRUIO6KsFtbm2
Wq5pTKMjo0thjsS6FcgxNfBZvazxo9/PmIs6nJ3/Ok50RM0aW0/HorUaVQ+i
RYsqsF7s/6iBeyHu6nYCk8bsn4WqgGLeE8YUI4OwiiU9LSf6Q40OA1BB+Eza
cQDjNzbxdsLuRYimEYVj1C29VFXkl9GaJFXXlDo8drKFoffxKkTh6N4IeEVV
fYJQJ5HiwDHU42pVS5KHe08Xl5hbs8J2t33ykWR8qFX4WTqMX4706wwienWU
d89EBgUeBWnhQqjLNI+DcWNV3JVatr9Ux3Kd+cdjPlGPUvmRldOmhZxhqFVn
ruFOWArX2xTW/Or+bHJ1VlnuZT7yvzRjcWOShhx0HlB9SzsieJNCKJ5PZlkk
h3mfFXQCYftxSkBVhG93FIjXerz0IFpcO+SKAznleJx6Cmsxa8wYOqM94exn
xffPofidMVewAHyVf6MV3QGTn70Vj+Bl8IfETBC77dA6IKm0HhxocxlQuTTb
S7VS/g8WFwPKkvz8jqc8xKewN1lpeuQc+8xqhYda3qQKbLgpixf8qvfhkhpN
bhppHnt6MPhGmtWulAGlTKwIpSmONhge0Y7o0AKHnmGwAxoy/UdYYtpKvnUW
0T1YpLMHcBz6sAA72s26iPCrexg/wEnJHwdrszbXj1ZC/VR62uEiO4oJSMOD
wS37o4rqbwHeliqi5m79BAl+xnFacZYatrQR0xRQQqO0SbMdjMC5DKlXzuit
7GzHRPQOJf8IfiLcv2i2t9xc0JFaTT/qA2yiGjhP5CsMzU+RCdkEGY6T3bso
wfM6eHkQgtxlmoAaqR0KJoLudR3T2qlq/X4hTbu4JgU/GrlzyjWzVF6+F6hL
Dt/JyG5YwyEV1gaf4CAj9UukmIzDUx89VRpVCvWMqUaCreJEH/KeIVQ0SOrN
9hiBQpFqj97c04Dq/2HJcKYnc8xJOQcw52wIyl4DoMAkZuNrKBPRAL0fuhXL
s2XRaQLn4BPTkxCxPjHkC0Fr8B1tW9iW/vJGTkVpvTU+nG/gYX74t18LkkZ3
WQCd3Zzn6K+y4wCQNNunHVoYzHtT0J0k2GQpXCKqlhjivx+IP1lRrM0rrx4y
dwYWg77ntVrSSrIpFJpO0DIs/6DCvjsn3TM9qnTJDlDsTBxJ9imPPslT0dbr
MDeX2chLQ88dPIp9lQwQ5aa4xAhHtNF+Jytv68YnDjFU/0jM3p0eGDS+727N
nWXl0JpFS7MxoZyzFBO3P9rP6k+c5qvc7beUAMubs6ETpGw7OOl9A/uNra0l
zII9nvA+7U7HbPBAEbEq3NPVcrs6WkrkAfWUUrirnD8gVai2hJZdpe24deZp
nnS0bN26ckemGqSal1xKGAPCnO8X74KPwzyuK4YEg/Yzb8h2gxS/Nnj+yoXU
8wnMO2qTVQvb3Wq0QeBcC3XdnzocLMyVXzQTCJSKYhIlmpVTjuDHz1AFRMbZ
gp2VCiTkPAnY62CwZ9JwMTocTw7IiMTbwqFXqtWBIxzv2Qpc1dFKBNVWFqEc
8NqI+0cS1jylWKnBOvEK/cCV3JREm3vMdQ85zLmY/bf1DL1jJL2HxtG7CFVb
L++fFkc6z1nGgJ8agBLda5cfxk+Oyz5K5Kz/EXdSl/kKpbyO3ISrNL1xu4MY
ZArq3FP7XsYIp3A2QucbYZ3bqk9RCHwCyJ7AFuggIyqGgZc2pYkz/xVvoIYM
P/6KWUxiY2929BeB56pFDYhcj64ZPbqMzCXQtbnBhv0zDMe2CVQxnEan/44k
5HU5g/t5znII1POMHQC9ZPwHxejqP3GYFuyYevkeS0GUmcvJ5egvwQbqwt8Y
fnmzjFTMaXILzVlX20CTY6jKrnd+4GwIaKPeHGYufuup9NEM3OBVKzjVUb7I
zrGy9d6s0c9fl5vFBIIghqBBvI2h+UrJ/DPS4xN1jahw1jlT+nFe/6Q0Gw8y
wW9y2wvbuiQPXEDG574Whdg6W58iwBm0+Ew3E0ZFu/3izc9e0JHE4BlcjP5C
kYDCSt2LHxkIv4cYuYw9OlP9uL7hl2mRFnqgNE9pTEkVCB1rdiLrvNf+jd8+
rXPH5T51MRxo/xf76VrmlxY4YUKAyoMQt+uci/3XHtT+fjr5XdYDEJa5507f
1JfiLIze58BCzf3nZTlXi0wyx8GnylRArWAO8AdS5KMYmCKFgtsnpYF47rXr
hmnr14wx56namutTIqILBWfF7blamEiGHVXYoWlWV5QBFIpBgRGVZ0rD5ftR
GQ9tgEx8Zvb+3UZaN9ichJuFU6ydP/p9/OrDhq0ojL9YdoD5TdofUpndhzEw
SUFxcW5Zd8JHTaV7ZvFrrmFBbD1+pDGftz9sxD4eqOIIAwbXVCbw7waghKwk
0cdfInKbk3fjUnIEPrKeeqF8mBEiBQQmkJCJRs2oaWXFIDGZY2a8cMTqcClv
/e5Kxjr0TsME82LIHqRYR+uX1J+3KFmRttvzsfdlIiVNUhDNDb/BiyRhRFMn
G+LObiKyMJVNRcnIzgigtOAaG00NPLKQJ9JYrtMwdvttKsqDvBP6eUNmKK0H
rzxZjQVNIpJffKg42n8xNmR2TBzR2Ppv2kGeCVmcrUIBkgC/YMkqGGGly5Hq
8INBnFLlsiZm2UxjIAUlsm3ZUU6FiukI7VWGd40QKIG5daCcg+F0SMUC1v4f
qplhUYpujL/7uYN+I9UN/YTARwfcDrYFdBipVEWHLchRKXbYcsyymkeSrjC0
6WvxloibmazmbR9lBtz3t7EH0Bt3yncIv8Lttf6I11rKaYc5ZWV61BA7LAmA
sWq+Uu7aHVQTA1GahaTBGaioN88AbBj+5+x5ZHACH7x6xmBSy54Y4+pEv1Rz
DTAuX3abRkkiCgDwr7QHgBCuzRk0xcq2ihPklYPusmRUwagDcQXqJ5a+YhgT
NMNZQkZSntjsWcL/ULwn685jmp1pYz9O4LI+Afj4Un1E/E5VAS+yG9KxSJX8
dge0VkQzQYoNgVoyzdutYwct+nCrK4k+VZBxZc14QNFpPNWK8qD8GUi1FgjH
pz3+AQS1UlSKYL6IGhdqw1jnc9KMpUrIUtDz/3SL6mq11CMqKU0ncorZVUwU
aGy1FjL5/FyNW3Iy+wRwJw3QeSNkQyP3D1Ag0CPRfdVvt2eE1Dr2IfPLvYsT
/mBVizptCBjxDy0J46cBMmd5QY1gcEdfNXfMYDiLajrosWVIQW6gDJMl+yLf
S2TzEINp8tvuO07sNpLXI/hUzITqdSvMqnn2ZcRy39liWudfCVp0OBhLI6F0
KyYnB29zt+QIpZTzSRS+izZQHgSYbkq+72bhepZwDxeXjZe3q2Fi/ggw07Lv
ID4jwnzCxmmqpvNC3skT9TTakljfOnmb4FP/D1uJU1As2t3FJJLpAFEirusG
wfwg3uU3ttO8GEyMKLLhyJ4y8bFozkHzPdbZCMCiyJvxLjrbw/C9Qa9t6eGG
N9k/dZQt6iLUmIaHrBLzua2TbSVzI+5TMlZ0CAFbC4Pd7sFoAwJ0/MpHEPus
HfmcVQ1ZlZmQ2fXczmPRrVGLAj0rtBcC3P1Dw195G/QodoD5dybhDEURa1z9
VOzj8nzGVA+1NrtZOn3f0JEfRTkiOsIo3jriHCrdYr2zTFBCj8VHYTrt1zbn
eHNfap3DsPGrcJ4/Dwj6oJtukOPmB0PG6kSrpFyQ7R0xtQ4dHhu2sUGc0xSh
FTkWCHc9FXYG3RR9gD652ahPgBrDD0Wv6f57Ij/nyYoHt7oC6ybYuH3gp8h2
/EnZYNII+aQ2NFPuj3yjMmAAovZtMKgfFVgziWYaWXY+coK2dt69gDSbbUO7
BBDCQ+Jfmt5ZBj/h9lk06WT9IoMhe1U4kqU9nw5v2/ZDP67MCBzmdL+x8v9+
0Grimk54zL96U+C04vuhi4lLryX1oEbMo791ZbV+/7rqcNAs85kHlH11kTd9
W7cK76LF6igb9UHEwjZGoKwCiEnMMINzEuPq1vMLepH/x7oe6AVEzbnLTWi/
rfDaI+QLAgKndPfjudAxCRF7qk6h6BqqX1N+TxUZgTUC1khh6JN6QMAIltZ9
k8vNkS69+xgXUXE0Zc8JEHMMCsNFeLPQeYy+6zRF0OfU5VDCBR+Kx3Y2Xrbw
O9Om3UL/g1YnCFpq+XpQO8WozWqIhMeHj/04OjDd5IeFNhrH1JK9f7vIjPGK
t/MSij7gcTOe4ba/b2YMdaDQW7PWFKj2lT/2FLu+gdgMlePblRmtgq3Axwkp
nGRrDKZYooPGrbUvqlHdTA6fmLr2IihXLKL7RBF5n7rkuPdzG78kEWsPAlks
cNXb/NQB/PLHKEgr8+PgLFDXuUeADlj80HQKaqyFdd+kD8g9vqBNTIDleVnl
nwuevA7UTLpGXnFAWbqJhZseffJATcB8GOmSA4bqX4YUanXO6EGEm0WomW/H
/McHFs3FppRMfCTKqmtUHLbLtaPuHk/4W8a/68iDKLI7BHWoWrV2olb+oU2U
ARw+KPdSgqfzfVbGhs8cV3UtQ++/MOtk74DMZO4t2uHd10DvgxHqMyCBaxfR
2W2yRiLv0+sYXdj5qmEnAvQE3NTa+mBr24B34BVSRLlQtOkNd5deKw0rU4vF
xcIX/YjPkjPoINWo2DXoYOLfzMTK8V3yPWltfjaGw9LH2vacVb32D4FGBceP
lPtrmu4Fx8A8mdaFFwQtQmSchIWdwVUdkr57jY0JNi9dUT373vE8xzPIsIR7
rxp01Ne6Y7veLhd2C+eEimuSajWKzRiTA+tK5eXDd1p+dmC/DLJ4q5b4qsuc
x0p16yfHTv5rnbhJa+69MiRRpwoULMdUZ0aPqjUR1g1Q7pbXFxxpdJa24XnW
Zo4vwQSWFXppBCAKBxIW/i/yv+O0J1ke0QVqAJ/4qelgAECaprJIyvoO/mwW
TNLkBcy7M5Ze3vXMSOYnDSpR4Z6R71JScB9mOqEtajvXk6OtOEoD266FwWwq
i/oU5cQMnsuQ2kTBYWf9j0mier5Z143XbWGbsiT6Mzm02Zfdugr6s1sWhMa/
5nwLrt3nEP2JYfN2KqcIFKwxBeaNT36pZABN2MgMR82JnNgsPsvOO9Q+L/Kf
N7NP68t0jRtiOrIyQxyh2AFlUoMqbHJFwhBh+3HiPSfe+N5TqOftP2ybKj0B
7HcjbyYxFXGxEsFZ1VjqikbG9DJeZhadxFDMO2ILE/RtjXUmn/no0Hfd4U37
lCQlKRnS+gJwraNwVIlWk1v1JKUpzmMF90hHk7A1iURciaVcGf97ihO2xus9
eCwlsayhxzu/74bbgDVqq48EsCitaCFL3UytRLyhIwrF8yv4mCX8CtyQoW36
Ynn7tVsWxzwYmqPX3zZ44756ai0RMDuCn7anzLYBDwkiUiA+1BCkQhHtjD9G
l7cPZ4SnLlXdBYxFtN7noXGCbVRNwNJc9Rrde99CRYNP/OCATMCwppwkJirM
JrslnRD3eqFVVRm37Su5uLdKg25sMBxecj4bv6zpWPQptBGAisZLqFws4pYA
JZzzhU1p3RSSEBJMR7k5i8/ZdcgFNHBLPgg8BoX+P23bydbfL16S0tW3luJC
c7Q1y3TdQpVq+K+tGD+lVvCpSRk3INg4355kcCdpXgme3hgdNivC+SadkT8j
gUpE989lwBLvgz1WN8nRHVCu1D8yjl4+gayw7kcvF45pP0NTEsaN/Sie4ywk
XW6JjHvRurHeR3bI6kxVnrRD/SaFcpe+oj1Ri4p+b7xIGYEv8WRni5eXU3DI
Oj7I8tbklgxsgf5l0MvkE3c6gMmzmDWQW2ouHhM+1RPHLsZPx/BeMR6ps5+E
34juY4vINt/j5mKS8n9NTxoDSkItHOhpFaH/2qY9EaGNj6RcggbpZBqnlugv
e3rgRxQFB2CUr8bjfRGd4E3MjHjzB6MQ29ANp3RmO6vecGVhgh0E6W+HCEaO
i0QlGSZcddP4CydVDU2d3IkmRZG9Mn+2wcRx5bHGZSTX33mNBGG64ekPHADz
pYMHbTlR9mz5zuoLTZGngIM6XIneUNBlQzDEsvoisahnIC8/8XPG2zHD/kkw
3G/3DEPJft/lphBWjQO5EYRDT1uFdmmnhUtCsi0egR2BpSyHgvpsZ9LGpiKZ
HWd53BD0EHrfes82Zq8wuP5eSUrhkLzRusTAvOt9AunQe/jiE4OIW7nZs87R
EVFCzstUvvzT7cAo+eD8/QvwxVT3xLx72CN32nh9W13pl+biWi4EbepylVHk
R0G6wTiBE+DCIBTz4EHY/V6v5FfA6ISTIzR8XuhmH+QijqZjwG15BUBrDP0l
AsIyTIUP3k0LPIbz3SLzHg1ey8U80FEejKidjvczj/m7jXHaGjQLtm/VoBAy
QEZRd9DricJeHKHbrq6wam/enqkaWWXmbPZBbcgQ0b/jgBteqITkAG21LxJZ
81c2kPu6uqTH3IwDTgOSVCFnL/jpj4E/FUK41b3/GRZM94KcDiv0GtOAK6W+
4tyX7D1XIfqQYofnIL+7tsGzznO8YsadApTs42n2XkYrva7BEuiUmAwOHwTi
D0mpox2rQhj71BlMxyXH+iP4Lgp1NvaQZu3d/+/mU7FChAw7Fr4nWCux2jSC
l0zdYS9BplPkkGa4Coans+eIvKNajriemtOus+Q+ZcWPSynJr9+pwf7+7ARz
aYuqH0xPVaPvs4Gi4ytd+h2rkCls9rPLij5ZrZuaoehnr3MyPSWsVjczugQT
ifu/tu3MTUpF/D1zVDFXL4CPFMELb/Ozec9idH5fwsoKrXbgWVltApjWLLQB
UYr15EdfaPsn2Ii0eAKwKLI7+Ue4yaJFOvTdS7ALLH+7BmY3d4xSMvaKSx+U
RtdRMMLwu///wm7FGEmOYkyux3oF5WwtweQNs1IE9/I96bi0vMuruGQAUbBk
UxqYry1rVrcp+Sm65sbT2FTf63nQ5TDnA1mJjSHMkXi00CarsYKSeFXL3z/C
DmxNrP6aUNC4fxoF7FEAhYIyW1CUSMmBIsShzwSaBmPqPuB93B2CY/WsxY63
GVbCcXh3Mose0n323YUZpm/joAKDgYa314Vowo6BVu0VG5HlzalKtW7fGrCl
ojc0XgMaCyroQh32VR40q5aZJwGgcrZvvPzTG0sUQ816HW+3F7qo2UdFV09v
NcVVky2ykyPc5dyIhDqCmmQ+04u54ROGR9W2DeDQ2P/PdArrL+IukaM+qL5Z
s8JVvZXTFf3z/RtO7ywcEFrx9lEELW+uEeKnzZBQ3N02Yq19a5kZRgHbMgNt
yi8nfmDb17/aIC23a3xYZbcov1LSs6DsBA+r9tkG9U4hzr2zb3BEKQ1zK/K3
hDs/+TvzLsH917/PVCx868kMDqIclmWvMui9ZAMT5uezcrU2gpHj2pNL43D0
wMscFL2u1iJQmKyIxTm8oHogcgrXekucko3sb/RCQDxdj/814m2g0Psuk0RY
LOFALOdkfQfGpdo2YBCD8b7CoqMPOuO+Rvct4ly2aX1Hli/cYvzwJDM/mFV/
QoIoyyAIYJqplV4mDtDqcff17f9T5OrS9c6wXnYO8QOwYFGjzxknjDmOmYe9
69YZvLqzBYgdSzpzuQqdGY/qYwaTM7qU/Nzr/Ko2MVY4gv33tvHsF2LncbuE
kUF5JbhMywLp64tm5YJAbL5cm8sHPUgx3cDn0t5E45s4/xGonNlHh0nNUnt8
qRdxlL870hsP/4/6wEeiajq0NzMXOtehqISAAb8NrhYUhMDkpkiT9fX6xzkc
aJ97iAUEd0BvEwi8irm4a1BIBoc3ZDuN1HM85BvIvFDLdoTK/xjAFPCxX5yZ
NwYT7XyGK6L6LcFn60NiYw63Jvcw4hW+fJLk81vlE2k51o0tZUPHLafwEAX3
1DFV2Wp3RQRIi7r/ouOxKz901s6y/0hUCFOipkGkwrQToVaCBASNb81BgB5g
5yeoqevLCaO7uS42/QzCIdGcmcIfljkYzf+5Kzk4pyCPYGlghCDhQNqSYXdT
51zDwbQkrEeDbdZdzqmKLgNzMqHUqbJRzYhbQymsMzgp7hQT4TlAL6gl7nOK
eMoTmE7FBCGyY+sltu5VsiRufOg5/RIx8+LjSyYTELPNBTljZ20bNw0jAmVJ
peGQZH7xmp5f5az28P1xB7RvCFZfr7CCzbVKWY9PGt4Qr2U2hfvPG6cbLiDb
q3WiHzS3YS51LvHXFaAqzrdOqvsyOzeeWVSpo5+ftSWYgldT36BQRgCNm+uC
9KyymuoaAKfnxeHz/QQl4BQScLcLOl+2a1oZ00LhfHIszvEdQgUSnqDpS9bv
HuWdP2oiPcFIb88OYU4wnV4HeDq366PPWhhntfpnbwO1QWV0pMIgWQfCgYVK
Msk2YA1XZr3EwmXrSc4T4ohbVI5k3OcojmPtqsnI9i6rNU8xjDN6t7mBErlB
gmUm9rUyS6H8GS3fJUQLs92AxmXm+rrRIuo5nqcM4dgPhQoeQ3VQzzNCjOf5
SMxYN5ZhunRxAP47Ezk43O7zzN9jlvhoHnxJARat/bJS8Zf0mm5GlTRrDK0/
6h4dMKhDJD0kW7NiEWc2L4YP/yn52qk/ntf1Do5nfNGlkom6RkR2hcX+3QfQ
nNCaCZwgDDLfYrUE/q01cJlKQXxcppgFU3VqWIENaBgPY1I405i9JI0wYdLX
BxqLQnEEcQ9Xu+KvAXOV1y3Nd0wELD5JRVodNMqbYUKDovgXuhbUqAVRkyTi
CgssKU5/nRKXZFgUH2Ff1Wxim7PqqpVpWitUvpPnGMNzaFOG25Yz9cRt6jC7
VCfEFJJ90gzcS8pugYwqgSLby/07dVODwtmRRVKOVvj9XCUxKXglzFw/GkoQ
1wY+nuVCsoqOGlfKo471q96owhwu6gDaGwzaBwDjr54h3tgZai6JIN3GvYYN
L0/BdCGHvNFo1F+tyMRFR3NaMgoKBQw2dPLyuuQb6IYFJfxaLHiPyQ4Hdp6c
M4o03DIMegoqx6SkP4f41pPtwmrj+A/643ZIx59hUoasLgqbcAyUlp6ovalz
9ThVr+9i+62s0qmJQlfmDOtdK8kpVki2YySSy8ieOlYx/sL+nq/YDK5aAXqQ
G8aP3L4ODS29l7uCS3oe42sLuEJX2ZSBtWCueVQVCTbOuOui4Avw8m+h+Gqn
jl1eA3BI4ytgPFVD8wdoVhcS0A9zpDdXa7exzd9Z4QDyFe7w3Ic2gsfP6HEd
7XpSK6aaGGYFkA43j1hRbm0llS6XmcFtmae24zgHGqdHkGRIF5bGNf3uxzX8
KIV5YkvTqJPKJCLaOokhRSx7ybN61FQqN3qDgV7FvX+fVOSNDoUPQx9BiI/R
pKI/WlfoSRajMW1MFOBIlCrrBlX1CgQMQLxdf9MGRukEJbGsZsTgppYaAxGH
RwPmq0fnQVH7wt/REGa/DTuG66zPlkQIV2mWkP3ilufrBjFPetpWZVBXs1ha
1/HgfJkYfvTn0C5Ng1xTduD7Ft4X2vSrSTBWZkwO38jUf0M2oHmjeZjQI3ss
PHjs7vh8+tC0NMDjRiRyWCmk+MxTRyF18p9fDI75SSi815sP/+vseD02VGbg
wqBNv8UdTkjzduG+RzmkXMF1VybKN6N7SoPH5XbaTHpyiDWiPx0VloYOaaU4
78KxNoApVn/REtyDuJI9D1vm5iroNy1+8S21grmVo8r8Xz1/h9T0zRMZHAEg
ob1tq/lXlMOw43BvVhQbv6u10fGcMAwtJDfdQpqw0CeuFGhjVgEcDM/DgbF4
cLSvnamWY4XV9Yu6+4GEsMxJJdoFE8FzBZrNPE4HWfY2bqPOjmwjJLBgaZnM
GhZrKolnRvUwYX8OHL1nAfK1sR4Vu7XQc7LvcAuGQr4eW1bmin4Gag0Z9zu8
COLoRknojmQvAINPFRdVKhk0sOE52dUX+a5i/lRFqbcMIZJfimK41hfCXEJJ
D1a48wEgNt2oCHgOY3dchytydVjd0/27kZ8u4u2wnCeZRidfgGFv3NitHe3r
gf7XvLb9eMRpD4BU69tNymldFSit7pc55POVh2xYxyy0kNcODMRRpcgvaipZ
zqLI0mQhBugDRiFWf+QbcztjtxfuUiCvnlocu/l2C9ciXQBri7oVW4JyeyeZ
dzZRpVo9CdyAEW9NMTLO6/PLEH6lsz5A1KZcbm/AaFcMHF+OJLhu+kpwlKZ1
wUZFcFpD4i7hCPhEZOWHPk7OXOXFxO3/Sxs6ypVeM9Ji5gk8H0D+cgwMc2Sg
Lcs7ZaPWlhawG4Byaq3UqMW5hLc2YQgewOuZ0Ho9wcEl5qnqezUEEDJdMlOx
Ei2/vuVvhqtiUdsjxi3L/r1DPTtWkggZcK6mKHyAXG7fzgtYu+bPW3pW4euo
5kfRO4Qofu1VpV9C+Eb7jPADu/vsVWp5d34YdV9C3MuY8OD2e9UliartKcU7
UewM8n92BJKfduxZWZd5m3xqSaA2Ou7yNaih3BHq4bvNEF6PzMMdpBsuc6QI
QQmXLpOZL55TA2UJ2QqWiPW8OMVImRNJTDDCmsIfPNvIbXrvA+LnWLD4jGLF
qaZNuL7NtOkhGMUlCw6RuTKKooPlGfxDnYgTqVJiZLgq6CJWKl4nIt4/EVk+
FVf9Nw7ECeE5OxjErDHV2b1Dtcvcffa1AuZDmAiwr89h1Bs1QiN21derWl04
TnSFdmBZBaqxfTNUXfeTypDFo8GbN13cNQJP7ZKaFa3Gq39BVAsUc7Ae65az
RvA0+a27bi18y+qftAwOG8DWch2YFrczIKOcpP8Mg7m6u3rOcGagpak4gOsX
PbwiLq9kfUrmBKEjKQD1w8h5ARKxD+ROAFsBWZZCRRA2VNfE6qfNa4qOsuG8
DXXwI4/k7feSz8rs9jtYGAgvM99VHAxUtr1VuMS7Fy/GlUclaLHeoABGrav3
BI1Sxai7wa+VBH3Ah3PeNTrMf1E42+OcJ13MpC2M0fC2sMyfhEAi2ksSdiTG
cxYcH8DLjbDSh8sC2fWWfyYlsuvJgEdeMHZcbqRWt43YKv3MEdeGM9JjW/vd
9p2EATrsVIyqcP6KKU8YPSkfuryTQ06bLtFXdUhmCEaHW+8jEL7L7RSaVFdD
qCeBlwvoXLO5JT/C5xUSgvgevs+tINvNXnshuWrXXh4PvNXXkipESlQ8T+A8
QNlPwm/iYg6FYLh39UnjcJFCqjALdooC4YI4ctOA1Wgbh/v0VVUkNjevCprZ
W0Av068TLYQPomLNz0kvVDjfMKnqPeTQr8i16Uz2liJ63FyQSO8Qv/MhCbOZ
yQIHkqBCPDeZqesTrhGeDrkgHZP69fzICY60J92OwfYZaBrD2NpOjmkUkzaj
JlFHVsdGu/cKEGNbhJ9D46v1o5AE8mUZAS6TPwf82MVJxhbPAvruBM8g2T8v
LtfpUIvwDN0L4/lpkzmC82WRMLpr8VP1NFMp0Wjtq8Kte0ITlLC0Khn4rAch
50woUTQZxoTa9taXZG5KNYnED9MBsQICbjjHY1h8qcGN1B8pMXbAMr0N55Ys
QWyepKKF35kHtwQE0j2+N9XCNcbZXxRM6/pwiFJN4VlcIMq7qE1GLr0hc5/g
VrlEK1aRZ9M+Xdxicn14DesKnbZERqOgU2xVDbLLFkX9LPK7VJsuyHumHaRq
lho56w41PtzK7VpbGmMIVsAjmyzWaC3xGfdooyQ6QUVAmY8Z0G78BwXfybRk
LOQa9yyaj0FyJ8ghiBbVlxWD78MHkwx3cyjIY4bejuk08ziegCjGqmYgi21w
nsKkKuN13HKqCVfNsjyMNvnTJd2kLgwRS0cw9ZjZxcmS0798TOPX83e7TunL
eFjv4YqWYzzJDD5/zygMJC0uOtDwl+v9cj/BpP5VzlJLKWgbJcNwIopbeXn9
IK3o4qFnD4sznybs94XFKpQFp5P8XWuVJjdoGGA9Fb6zlR+QZPE/Gfo4vU8d
Fs8Chj/zdTXgNuUbEx4JQUgvKHTRny4cNq7hRXXDIKQD2b48Uk3Mmt3amRAb
xNSUpBdnnjiihz1n+TbAJ/qPhfjFyT1MkXcI0LBoi2y1UjGs7LHI5L59+qNy
YYkXP3cgB9zxVKZtlyURKGazL3+bawNln7hU9jBH3J36/JMicjpxQPtV4YTQ
9CeZo+NBtcyN2GxNwOqyU2mkE2XMz6Hg3k5Xs+bfzC4z6RTeIBOtgLDCth3G
+GcthkYjMDC/d94uL5Avme9vnI99tPM3xitzYJVML0tkob26IEqJmKEPeT3c
ZH5dUwnBRfOtGY1rS50FpdbV/jMCWXd7pA3h0w7Sq1lKsFcU8gfsb+U03U4E
QkBwJZ6gaU5VW8nVVZyieOU13xXN6xsVRnvHW7te7TW5V7g+DtHVBPOSSGId
PNdPaMvLiU0QeSE8U3WiUlzEOoesPWP5gv6ciS35U0MwbUOWpZby2BBrsFWz
k9hqCPV+dGCycijeQKByBJcsDvdbpSVildVWm0P7SMx4DeW2MGSlMRDR5gXQ
VxDhE3ert61+vqUAcbJxBSkg2ig/cn9Fx/3CJoarh8TCzNE83eRjzkv/ZyL3
+kOh0FSzIBOEZAb/+4VCCrPkVg04FsjrpaUtd5jcKA1wGm0rGQNWYK2Pcqh8
jIMzShjMVmgaeBkU4pAKD9RGnfqJftu3bJlky8YdpYsaWYLYrW/fAKAOwUdB
bnp0Oi6hxzzCN2tOkpwhd+NgeMIi3GSwKL8mU0/3t8579WQZKDwXJ5XEvGYJ
izVeRkpr78TBfLJLzXevvdvlS6Qdl8sU5W1zkSQiupAn0mwR3eP8p/leNn6k
8UPwcAYacViaogZ2aiG4Hc2VlMv/+quLhwppSnFlEV12LrnzLoKqFTOMqmTR
5o1cex9G2sdCVlWf4s4KL1Ykg+6Hu50s52SlFl6tCA0vmQ6be0QHAWZXhMLC
zzIkBd/tmp/GXBbTdJjwtkSXjGwVHFbOUXyziwvYnQESH0ly9fTVxQFOHSq/
BMshRC9UXc0CcNhPOyFrVoazg0fDjQmnPxLuwrGFX4cH7iPvR584m8utlGGN
xBAdBKi8IdN5ys1ENE8z48LyGj1ciDo1xp1wUWMkZQli7KqySCVtrSJ1r462
fS7TUeEmKqxRTqAGKRHMO81TWzW/wmrjJmPY3LNneNXtOTpl58wRguzzKHnX
JscDW1GgG5SpuEk7wb2AH4kqT33oU0bVkuCvTC44glDTfMzMaNQb1NJDkNxX
LDbENrGIQhuZO3erMUQUCjiHPh6dDPJPLk0wAQUzff4KQ3t9RvzeOz1fTKWd
mKfeejQu+oWByqm7nW45G7SuUrOyVj5zPsFq26uIdHsYm6juYYSi1KH/U3Ei
yFDAtGNClZ5tUQ4G4dNwul8Bnl9LkGOOeDN20HXjTExu6N+F5rJcj0ZjfDGE
f1+6/zI3g5w/21IYD4Kj0O1M1hYXLh8r9toSjSbUBi5wYtAsfJb1Vv5n4Jyy
GtkhVLimzkE/+qwUPtKmOqTQ4ERA4OgQcfkpzG/gjCKbtdxS/KjrPgALnMsQ
7utrY34vY+S5AJh2L7bZ8tu3b/tCdd8IOXFhIZJJGmJnH5izVo+CuXCe2xaZ
H3zfujhsahfooPhHz33nTilxNWBDk0MZRw5UMqxNrbNnsaAUAURy76o3uL24
dAVDtyYoSYCu7BDBJVBVJsVdrE/hsdUBPviyqENfCwGtSZIXQQMX070I7NCu
B/Cvv9nCZ8hDTynuv2gpqFPNu90iWsMifLRdZq+BKRR0Rp5jxU3qEmieON+G
JJFj/ApNavVZR3YOakDO5NdfIC6Lv47zLydCicmSC/Xdy2fa5zS62hK34KXe
aVFfo1L1nhLF6fO49P7KRc6etOHGKYHO4KpHo9m0p4PnNts5IdFqHUhOEqks
KgIV6vER1DO2RElCwFyT60MNsbQIO6dwXgBvs7F5MtBm2DXVFXI69O0LbFsz
nACJXglqw0jHXU0AjQ81Xr6vUu+iJYoDwDS+6++OkRFH385QJARQ3nOYVXv4
7gA61Lgl2x06x6ysUBcOMfsYOnqYySP7vZs1fDJWqZCAVPovcrTHaAYJlHzf
2mwAVPEtc6qywTThxsNzm0TJQUr1U++gjKVGPvWtmWv7AIu1Y120d9DAswDU
gAV8VlWp/gx4w4rsIkEeaMIlLCMjl8Kbkdy/mEIUgCc+5Au5vnhZdtflfgr1
DHLLnwqe28eeY6JveUsyVb3SZiLcPstw51e5XqykFmWewGXwL8SqKn3Xna7w
U0x8pyRHXvpiGfzyqI+VrbWGToJu7LrqEiaOL8KFx6Pva4OKSCs/BiXXSJGm
B+eMEmCMhNbQkLedYewXadOCA7RKougbbgrMnxjLyL1k2lnDSoQuP3rF4dcF
1fXOQGJXWfh55aav16LJm9njgly+n6rkvSGy2iiGjZqdsNuL/T5+cfEB779P
QWJmsxSKE27vzMqbL8M8EVic7iYVFcBbbMKFZqjLc2/mblk20g2JINX/g2V4
tie0wjaCNNbad4+WeQLRjGGd7Ty/1j5msrzoCHNBu9aq7tGdiyn6oqABYlct
NPVXl5d+iBd1p0Bl1NRNQr5lGL4sZaODMtI3PifKiikNGIab0YVMRt9uooBG
6FRXGtCBHlDkt60ScypviramEnW/3Jssb2AH4WFb/aD2+qk9oVYoiHSD4Ul1
xDa7JomPlrx19TxDfPIYD1YXyMceJsu3n3STm+bDAzZNmDBdiwuoEg/El/9n
SUPSbpDyyjRWIg9lgerUOn6z8sFYDjsU5JEsDRcoTmU9U2htiW9Fa2XZZNC3
mYIxy9b+7gnFSXzqYMnzvkRelnZUGj0C1YoGShYClTXkHThOFK/4X2PLJth4
Jf3czEznGKmSx8CLnZzzRUc5VLFKM7b2itPEfLzJzBOM2WLLMWoGuPfm9Gbl
FcSsvyyUDgy9aUoUhTVuwin6bJCMLnNn/WhsnrU5xB4oR5x7PQv5HIGTeghy
EsvL6WTYIZh5uc0tmgx9jhP+bdNuQog+ONU9ldAt3n8lYcJidO+K6gLLte9a
21GrJougI38d4+zQpUqBAR+nqFaRlRLAsiCX9SWO58cprEzBI3JVBBujIuGw
HKQEUQb3lXsfP0gWenqtrumxffwSaKXcPBYR2dCn9Q9b21q28qLg8b4ChOKw
4JI5CkFD5EiseGrdR1XdeIcFmmusUC4p+xHXb3T0/XAX+yjcHtHFx3Md/iWM
HE3+vBza2W3/wT9VlDMQCYhy/5GUpHsMopq4obk5zhJ9F1DoVBBmXZdqDVIN
ThbxOB7oyUcQx7VLkh4KK6pFjnayFg3tFUqCaMuXJvhieuBRA/j9aClNw5hv
yjRVK6LPN+OR+HFPCJyo0yAxA/WSkOzd5EJG4gJwHcZ9dWFpSrKOSA2El+EW
BAyP1eJCIR177F9JSntp8H0dcA90Nv55PJYOF5cbnks2bjKW2wsG9a0gJj5B
WKgUxmsVeEhqimWhvA7ZR8VCkzrRB1XfwVvLW7Lof0XjD5Erfv4T3dtyfmNj
sl9zOhQ3e1kAHcK+ynqatLZoSuCOBwX3hYbXJprh5vpiXNPEwCvJ14EhMVwd
WE/awLn13gHKVE2V3Uar7a9HjLOgDPe7ZIErOJPn1/cAUTizly5n11L2Xcvb
DIJM9HM0Yjkh/L/gSXiSdV6CpMwg2ClUjM1zuP5sp4g8kNsP3OUJtEPOb1+z
1cTnFZ1bYeE126R5CXvOGAll6YlN2Poq3rKuQWRbi7KU6YpSnmo6G+vTmY2X
uJPM6pG5o7+8lzuj9jWh6VpwPYPx8T6LftQlK7WbdYOhEmZnj/iC1UrAhjuD
KukVqCOq9CVyDxIUDi2qzwcGJwrn0V9H1XT3zUxBsxnt78bENRNXHyfgS0Mg
ge1LKIKlDWDXPLUH+ZQuYRb+Porto1JM3ev8ZzciPojvyVmA49pYre58YjHN
cYKdbnJwwYJ5wgpjkSf8kmoBmkKw5hOGPbmVN3M3vV5+kzzFliKqNAbwBe3I
oRbjBXV5bxF+7vhR1A9+6t1Z1h2mUCEjkDBXIbLyCFtbYV6Z7X7oHZSROvnr
Ls/Tkv4uVSgesh7cQnnhlGzbJfAA/zInG4d3dc7rXE0HFPH5pKna7m74pJ1Q
UTwgNhtP56ckg3P+tEgz3X7/STIOuo2EVWAORZGoUyfONBAXC7dB02FKRb21
GA8khrds6GSIl/h50Q94R39HW98b+9MniUJpaQKyJ9IgK+knalC+AawVRKeH
Lf8gTH2GgIPHXl0b1BDXuWbeETYcw1JFdepSrqHL/a4ST2y0b1jGc7XE/qOM
5kla1iqVUMEOWw4eHS7khzW3kx2s7d5/f62s9St/ZiejDAWOZ4jwOkdHvqR5
M8SVt+K8+Eye9N+BjS3ouQ5V32r3ro60XWVN49l+hqdYv6my/kkbELjGZutF
Y6bAQ3MtwrRdWDceg9Pxs6QeGvJU6fJwI+1yrrbXrJSxBgyq+NcT4KqylNyZ
KxFKZsQ2qwo1Cf1H+m1zj79IU+Lc7Sz6jY90Bh1uW5A1YTi07pHYuxc1eY9b
/vxvPeHM7WP9U8Sn3Te2RfOtdWr0pgs1cwRRQBD1XnwPxXosA27JH67D8R8H
TtKB5lVRHdtTxZTAoEIwyiY6620n+vRweC8rFvcACjI6ZBGprEZkxx7B3FpE
WToaoTV7Tr+cbgCfPYEIk3EWl5rTj7/hXWIyywsFialP0pJBFOFYWnYJSl+8
eMk3yMo9wqJO4QK1FJKOmfZN/Bq1k2XYOr+DM6TfpwpaEe1U6Bb6RM1BCcCK
LYLDtsvtpLHmh6httuFHlztsO5IaamAS1Q9sHHytNAR5ED5YUtYVJQPd7ZIb
/K2aAsYGwF8KFYAH+g796jOiq/Cu+EvBIgATBe8+8MuTKSuF0TS/H9T7iKBT
7II3+1wPsMl2JvnLE53HEAKgdwsT6K8nQefNLeeJB8fhIm5qtmOjlp5PLCT7
8NHNvLUWJCP0N2QBH5u8nrBCBylDbhAtdEzxEOPUd95IeW4lv2UOiYdDBt0k
zQqQHTRdWew6jzSrmdyMrzrBynMhqBsz8ZTVQlmBqmL3QKcxXyPNTDMpHc1l
nYwvizzCkUOYmbu3vXXuLmhHhFEFC7YoZMaNKUToekOTAl4bIHAuDLDY5XSi
mKrw8U7DTo48qOtIT0eHnrt8CvcB+wi3wSA9lmiutKWzB0joE1woHqyDNsN6
hDrrLDQpmUHSQaSDcmXMaiC2M1wbxxpED8ej602BhUjXQYF9NS8sIA2T745Z
hb7LKsVtUDWS1VNSqXr46nRey0Kutq5HywZ9gifEC7DWzkRJvflm9b7Dkjsh
y97uJk+Zbjmwwf07+4NKbQHHG6l1My6Brt/CeNx82k4e1xPlXwDZ76VBBilu
nK8mNjw5udeIevoJ/2U0iYazb+s4sU4eb0lf/GLu5XKeMqVxOxN0kXEi2Viu
UKLWkOs0+0JbbEqjs33H0pKAO+bmufvl2cprJv7YlcMe/jUMB4RM1cnS9nK5
671vTXCaOLNGXgrjOUBEb6KoAf66f+KGwyxQM3Hw7EcUCHWEZ9pKV2EKi0iw
oUvgBu9meFa4eJhHf9dFI3VMLK4ow4K7Er/uLzrV6M+iKrfo+W9SXuCeeO3h
bqMEJVHgUnt8eHdGBrreG33ZtG3xp7BZt8n4Q+p/yvHPRadAHZIqODRYt4Yw
JDPHKdca+I1uyD5yaCx0VPMDH60lrs6W+F6ruWnk7kzkfPBXWnVUGk1Ok/1E
F7Ucj5S/HPRZ8wffBTs++NELQUIL3d93Jp+gjWslWaS8CoHRGtVD0vTrRzc0
+aeySpAXsuAC6xyoslD3O4XCXqPFzhaeg/Kw6rsp0UdTnazWiJK233i6L8Sa
UkQ1RjD2pRNCiXov7ckTwsVS+k3JNRmUoA9RkGXBmsXJ8Icg7JVeYvqsVsFV
7zNEggegXH6VWXOT0bSAb4aBWw99R34EABIDkeoRr3Gd3JCb2GO/Wk00VlSG
XqJmiRTgawrxQOqCdRGYGwI8zHddFQwk2gG0aKMGqulFA8aHodBL5oadNyPn
X/o3CwgtIF9o4MefC2eMNFzZEue4GN/t5fmB6tJJZR+wPG+Ys7yreCTlz7iL
SxabRpIuajyyI+sxvcLMfuBNKLfZjDzQJrL0t1DN5JXh4+Ks+pq9TjL9Ap1T
dFaA03B2RSvcTkcu/XVXV5ZtzXZLXfC6+vKQ8ODnLAzqwyY9R+kmcAp5VkHY
IULbn5zGkKhR5ckXQyV2VaisshVZW/Tyx+EWsTHoDFOx80x3ZKje1VeM4gso
WcGDAqWzsT4n9B1KtcIADZQs7o9Ok713hNJpwq7PVyivXsV56MZAC3f7mE8a
xdUQnOc45HP9RGvtkPojxvBgl7BI5b64MzJCmA8Pnoc3ddV86IhKlurE2mSD
jMTVLfSpvMnaaPu8rkJq7viZ4as/J7U3dWQ2AG0l2+RVI7bklgP1v3gqcmNk
zadpPbo5fJoMen0ZGa0OH7TJssLbXP3DwVp7gpXQjTmld4rTqMwpe4DQ3nVy
pspsQATE01TgPbfPiJBvO2v4AHlnYVOdgy4qz98l6Z7PBB/PpH5HWvfntMA3
6RTuIAzyX5Oshm04itJEpFhsi2dU1Hyf3vnnVqyNYr9j7Vl15cDycy0pEzJC
COK2O0oOf/M2eBXAGhEtBpFhZoTSeNIq+ygQvBIEkbVMaU42/0D5TwEhQmMH
dPHXiazBIdDzOZmMieUNHQfj+iWtxTrmJWpxCeemEoEwvJakr9kvgHppLe+o
nM65p4uwYps3ZPo8a30gWfXoLDW1lk9NFgxQzbc3p5nYuL2SZeIXAStYQkxR
99l/GUlN2XibdJxxm6Q4bkv6UOgDtwYtXcM9R5C/fu6HdqPG3QajVKe5zLI3
LJqx4cPQj8UGSvyVVArDzXD+btoh3QLD2N2fZkNn8C7MGu2ILF3lsZ91H8Gh
zvyU60k802KIzmFe8j/rQJewquu7C+hLNicMmb1K3PN9qrpo9ySiTV+Z8w/n
ak2VqRrW7s9wIhETMJHovDN6Cq/0R4qBm6IUHTmXyeJbO5UqSznKGfphLJPt
f7Nt9FqwP4bifB8EPZg64eQvXUrfxHhsrec0rcGUkxtCN0BbOy0vIf1vs8c2
cTqW8VD4HwcbDdx0nT6RRgnq7MBZIqUOlR02d/Bvt8QVgWkmK5YCeA2nmTkX
BQW0YmUqQxb/OGLvym+XXurVoLuQseM9Dn1Zwxzc7a2/b9m4GTBPFm7HL/No
J0ky6JwGtZWQ8qo3K7e0Rk7SbSjFT5Ql1+ncVWxQDNfqE6ZvJyXPHA7i89If
/W5cDOCNWnoPmmY9RbXeeHGsDdZHG1UHiTraYappGwShr+BYsfqiAJZzmnGS
vFr53XGR4jkVQf9SlBZg/KtvzBBT4NmdB5MZ3BqfUO4Qtas76V62FYqmrUqQ
dlWLf7KRxztrs6JWuAoCZmQ8167GGf+GcM5Q4DFN2ew9hIxJxcz7FbohibiI
01PAAnuWsEZ0G/zKXr+nLUKDe8eUO1TZvS3kGFX1pnOvrs9bno+y/OQuOS1y
SoxO7Ts/1X+qIujLqoqZcK/zhi4YgMNskB1ecI9xfwPXinHFD5OrztrOZnxC
D7etApzCM4Be9mHHt1WKfHETD92vIAhkmFTwXAgof2ZctkqkLnXAxHru4a6Z
TMxfS64fIyg01tbFBoGrwRuyAh+YPq+0y9/moy/aN/yXlsX6xObG8qEXfu5N
hHykF0UL7DUL88H6xyA1hkalsmW69V69OluuAPTIxbUi+nlnoLXcgwptAwVC
aZkJnMhNL0MJmb7mVHNPeGTvGqwfO3zPrxwY//gPT/w0rn668FrQqi82bWE4
dTnNmTIWno//q/xX4mVbewPaFgjEI7pX4MgBIGoNlDrPe6MHWoRKrWBh4e3v
MfCd4aQ4M7Vy4LbM5SywWXFhzMRUx7W67bAgkB3xUNn17KjnUHXJLRw2bUbv
oPnyfIxo5vMUTl7QmKYO+RA6PYpa/uhdq/M5iKD3L5Kbaeq8UkS0TlFNAp7O
S/XkuGlxcHG3mMZa6wT65DOpJOG+DVtUiGFF2qYAu/Kc5/R9jXYke7yFkd2k
OJvdz9MhChBOIb4tL+J9OXSbQTWXCiiEMhl3E2I6MbqY5QCX7fhapwbEKB3K
LDC5pERDfw+CAlAGzFLV/gGPPehblnyrs7BdkQoH3xdXBHqAzKr/FVtSRESa
ENZKizf6ijM1mqFUid+2YMxtU1GVu6MOFIzKQ+GnGOlH8JEnONP4UCQ1FQg9
SgkNmF8ORP9agYI01ZM3IhCVhGNlbqEG9UNdWqlaeiS7ewVPY4Hq3q7b+gS0
lCLt3QmTEi34/rTCYFazZ75v7lw4zSefSWrQgfxXJJ8oaKn1kbk2DpcBGMUG
BFQx1VCvKOCBFoFGj/zZPu9I63sT3s2QYtxRf1PyCdRAFQOuXtpAtIJyCAaw
iOC8UwJm+CWnBpmRImuZtNeVfiB8b0z75YPqg/LybZBsfsuG1jgsR8xAnR2d
J2xGp6t+tpGREPbsyJXeLPhrtL+AA2uDmp0LV/kncVnFOZrJbQL+1BgFEAJJ
4neE2V/UONwcqLeGVPGeEAIy+vDQ+T4I2ttyrRXghieuTwNYKdvCdJuL6p56
5APDWrhCMgigntRHhC3pAQvRKckFvoV4XO09eCK9Z5iMtTjxl6Ulsx647Sie
DsCf4e6FW2vveW0ikIqVoiNzuHMHNOeU6OufojxLLi+uapmBVwY8m8ReOqts
B9aU+fk7psig1XowAZoAdN5HOEcYJDlOkXPKEED1sF0fXHja4KsIEamUQf0C
xVqw8E61XeDxTp/eEJD8fKcj2Rd7qBWxZqys4JhHVkioZGM3Lm9R5qQ4wKSh
5CUhs/18baA77E7u8/MO0fss6BDstwlg5S7lOeMnbEdNas3z9XfeAOJANxEP
8ND4GKFcLUn1aRZ13rUa2VLaaBhIcA3lxb0fJ7v9MaV+jz3PuyJ7B87DMZc8
ldsgTPzS6KbOA5ZI1H0T1wfs5oIdFzRPRlMTS35iDoo2TtiJBWtkTJjB2lbq
j3zjEw8e29MvcAS98WUISO2PTD57g/KGM5cN+fTMfQDYyN8Gt2iEIQb98ibD
7Nx2Jg0LNT74Jgu5RKWkV9jgpB1AyNZI6vvJFxtALgQ2j7sqaWGjT1auy5IB
hDW4CuDnMLMCSMgZh9IF7cTkqJATjqsuHzwwOXxDr8p1FJu1IlyOUu6PBCLn
Nm8elZidCLwkgUm97EPdwBd7qSP+8DF6NP5WaMB52Be3Yr6ntitWIG9R0/Bz
ND5f/sCBnC+7g/f8qI7Sza3/Nh7yETB+JQP67URoi65syDg/NO0JNdt/nLHl
TtgeTJqhjIT1orU4xdtV37Rz9MZWjZrnxCNSXdva5aDOFNtlgoT3JJx/kSZm
rxq/5/kehaChE388I+Fz8fqFPa27LlyEylIv1gcx3GSqOGJh3tuix0ppAnTK
ufpEvXQQ1IrE8C9ucTmTcT82Ca5cdK7M/GuQYdzZVvyBw12khG+fVEFW08AI
AP/meiKMCYbrMCcYdf/Jzh5AtXePsbRkBnBNVCWEuO4Qi8fpPU82H0SVJfwe
KycLzEs4O22JOaQoaEjhl1x8Zq9tdHdMOv86bGhc9+prQ1TqhIwknOt+m1vl
aU9K19tIOZnfAhYDh6GqwMHrYEWsnj0B5DNFPZYcGsF5BayEAdQqrr0xsdnB
HSwCcUx9/kTlCj435SKqS2BzxccDxH7VLVdIdCPFzcz0dOvV+ZJlOvxs2btK
haIJNmuUTLFl6eHynOBi9yVkqKluHot6UAUBJTUnrN+mZKy8qv2N0KeBmyXw
GDT3wFkzkM3rLJrUB1+34bUnSePAFnH3+xg0iYgmb9IbsbucoA2RAdSRmi7F
1Nt0AAPgHfLWwn7y0EBdcEH+a6gf5Vkd9CobwpU1P+PcNuHJ3pD7akindbT8
VKvN0MRG5OVC2e+hE2ZrVpDISwt3KfaUTz9zBZzuV38S/jwyPG2wHutCQS7k
T3kjgvTtmwd+RXkGYNde4FYHTQKby9M+PrVe4czVbU5HLOD+gPwFepJCjplZ
TYOCfd3gtPyNSW4JdohPH36dJt6+C8dAQl6+LI75WKdThQgvbnCMmqXwGDw+
ATkwuxQyroTL1pimInGyU3S/d+d/YeVGdBNSbex7YQ1wYxcWzjjMIJ9b+xBv
DZSKccMpRj9izVkSiSy2mupgWPGZAOZ3oCGiedz63jgrLMI9xfocOtcvGukf
Od8doy4ohCwGyPMnrll/QYtbRbJxqI3HyRqsmNVqTbAHEvp94FGU0X6VBIND
840tGwqaTu2T2PG2vaf3r43VRtSRo1UsjsAKTJLGt5e/M4AZj2fWnH+xnEHx
FMJzkX+7DN6JZnGry1iVOt3gJmS6WmjSJfN1gAjM4M+TqNySRl45lStr2YPe
mG32FBx+u47+AWmWj5gS9d/qMofIhmZCBfbvSkJzsJ5fsMa7cYQSbJ22+srf
rp1mpYI6QVlXzBVNEslLTqpV8zy40U70WwTg6pljx81CVyvuz2yUF95ZWzPM
0rh8hc6VpPcKKlUht71sUAPkB9k3WU7MZ7/kvdxUhvaf0gtaa4sSG5qb4hXK
VUNW5mxhFsib062nSCKg2g4KszZgxBJ/Ig1yX4L0xl8mllc6DLvy5zveOSOZ
kwc/t++7HjLIf7k+thMfWeKO1UUJK+zVkS1ykYDk28XC8zUOM25fcId0Tcms
5pHPN+T+/qE2KU030FECfysCqGKH6iIbaalSldAISr1RtrLTskl9XjRlDGzj
X83tbm+xKn7XQYV1QaKPDgrQ/JGrK1iND18Z3yloxllfMzewI4C/lvvEm56M
YKTlMNlt/oic/MKisDo5vsFRme3S6SSoPxvGMiXGOoMtVEwR5pHYAYLMOLm9
niyf40PxyVRdDwa5ItBaQ/pOi4/OclcmvDByCiEa6uoVUgQM8N+WR249LY2G
pRHLzrJewlPjkq8M0AvCoM5dOx5m3Q09SO5w2QoXUdgEIOcjmRIRWLO+QsTm
dRhkd6V7yAsDOPu9xQTgsqqAKBECqXWx7kTsyiIdfCMeF+t11Awlvgmx/XdN
Rg4Dnz5HVY/fueVa4EXL1hsTPjgCBQ+78+z5sazRTjE1rNpb9+FI+GOHn2dF
XIYcgZNMlcMvbLmjfSV4WB9fts/iS42vF5pVEWiH9Hn2fu9clUqPikQzDJEo
3PEZkGBAoFW03Kw5wmA5tTtGRuZ+CKrhWdZ05uigSmpht5bWj5YTQuGLbmy6
N8QmkMeOZZVGmAwbUDmeNozbiB4B2k/n9xsXccsZYzOSHZFyUXT4gxiSFpr+
wuKSgMo4F3siLWMX1Pzwm4U1eRd7UY5gexH2vHmj95iCM6uOPBI0yOddT2ZF
1J/UqL7rSKTj5xh3NsvNpNsZi4UqrCHUOaWqU/TgxgItDZ2qyneMoVu7zUQH
+Zj8iJRvWoIBjsk08fJt5Dy2dY71b8yNGd9lESSXnpX3uXUPoxs5HACQXzBt
4du/UsehfXIcsZfIyml+kNCrLmbJd3rmTlv7opP3XoRRUeXlQ0lC+soS19Cx
Jhv4uyT+uacghg80PzRiuwFKDyDpunBkEaJOuHvp0Fshfa5GZ2/jdCY9qo7H
l4Y6e5rV/HW9eafjf0xb7KystRcOaFQ0QaTeB44nUOPOybfKiVh5Te6ssapy
s0CWHungk11BL8o4ZvvcsAK0cdfmuL5GX+/9vi9wVQei3KWDy1Ljw299ciie
xs8Ukar7NKkulCev6OX6YKYPMe3LMYE48n4dAjzEkDU2CtfE2oA1ptus8lA9
I4ShTpuz2YC5pxGz6hOUYCaRvjD9j8nF2+xrAOIlwi1C29p3qCxMBGdYXKhi
pnIg+pRSQGFVefvIQd5ZWDSGNXFNAMac64nTmJ3ivIc0/kSKuVpg5xbxAU8r
OpEfzq0w+u2Gj8oDPN6g3L96Xk8IOTrXEem45xDsS0OfHsgrOcXkKo/bhK6v
D/M7LZe7c25Azw3Fod+m1oL9e7nNWcbY579wyHXClWZ58bdLLSd8i42BOVae
DV3Hd5yVmQRRo1cKLTfxPl8Re2E1Ieoy++U57AkMrF6F94z1n9pnB4rp5qSI
LnpVsRMnaG49ky7QXEPRbE3sl7wbHDPjHbUsELQXIbIzAZlesH3YURt2Dea5
jSLZFObNIhtEkt0rWc/U4rwQIpwBOKy0mB0wfm19CdZsU2mGqLOI0buqESkV
wM/Nmxzd0RTYnI4CE63HJ0AuIydl9BULPwoKkPLDA1xQB0vKPIePjYxB3Ypk
eOSq7v7FsXE2RQ3a55m9QYtE44ee/8PTTX07+j8tfq1x009L0evnNLw40F1X
jF4BfInsc+LHEIv3ZT3WG7UENX/qyssots1W/cBpvFAkcWtEcxH0HElQnO9E
Kk5yfB7pAwb9Kfk7Gxr7Gi1UohEIT6SG5ZayNOBqrUMfNEsYBsGUx4Z4vS34
fnPxxAY1HEZ0LhdJb1H2a4u63DHYzk9oSKiakWLbvhcTtPUblty7Dg96c4Sd
OmrENye81TGXEsFVLVyOFA0e9Lxu9vvv3bSPrDIZwh4JkCdC7hDcc/BOlPa9
eJy8/HUqwOIwyam8wnJXbeAE6KEFwmdk0bhmZ4tyF5mOD+aYbXRyWsjs8tNC
P+PnlwcA0J+hL1f26NkDjBa8GtTWHv0bQUhN0DXRvgT8uW82RGCmIYPO6oWB
nN5girOmJzaRyfOEVIuGNOfGBAXXeLiROq/0hsRFCoyLItztFUkZmjuoUYPd
bUJkadCjm6hMj0gMdhzRGlPGLA2YYIqIQNbwrhdcO9RGKe3DYyYdVlhO8k7Y
JiRyrKtDp45GYINUm5HLfgP4nPPwBcdhXfMLc2QZVkT+09QsdXLp5C5ZljjP
2VYTA7LV6cnpvD/1TsmjsIrkut4mHFsAQDia5FiI87vQkMoM+7GGboCXF9hl
+CO1Ih8v4h5jQzznH4xpOUWs6xOnAqdacIGbTFCnHtE+2Y8RXQWVaIfnnLZP
RgrMAro7xwm6ajVCDzNofpiu6mZCm063xdjqTojcV8MB15/uALFOqfmMLrGF
YlYPYzA5M6B4joc5yW+A4zk6B6axJjws2qXRdsoCglNyw13Bb2yjX1DazO7X
2+LXiwFUgNd7ISXpaIu9AP2hDGS0zXdy2fP4nENm8xMOwG87oLmegBKi4Yqm
/vc54Lk5FB4C7Ub13/9ehCLUDxeMZuhb9OLgBn6iYx7Jb3zBvtywBq9UfK4B
nmA/YTBnLn0llN+Udzfgch9DlPbqvobFJe8skiwJOx3jVpY3cbIC56Z60jKw
Qkz7dAcIZRheqrRKc5CJjTPHqflfUt+ujSJ3yVZJIiG+3NdKrL0NdBBySQo4
KQGq9G4SjKLn7v4zdkjpUicvmfrRou0+HRENEEwbktkSdKGXpvV4c+5ge6H3
P8Im5QqQ8MyWn8jT/X2CjqOHp0jAG6iSMMyaqcQKtsuQgIjai3elstPbFfdF
1/gvPCNkP8t4iJxPJ+b7xAC5UdRDT3sMqp5Gy6cEDZbCfuPH9h4tnDdab4uK
iTaIioAbR5CFOwcqk33ZEOi0F18OnRLbcZ3PJP1Na6v9qA2f3/4ofvOiYtVX
6sb3dYzUrGAWowWQeZEANg2lNV9Kb+vO5au0RV2zwFOYvqcuK7lKnwBNXuwn
Nv39z8vCOt+z896ZFA6fyTU/btE+y3Or+I/kqQpu5OmXssKtnp3YVjHNVrlz
/2pns7mmkW9orfaayQCAVEFLdABgPL16mglMx8VQaaRCeL6eIxv72LdhzX1y
lyFrvrN8DMu7nJTwu3AMbvh/vanOs3jg4scERrlEadw4bOizzsKO3nbxTjYK
Q4RFjj83pXs+p7C7RcRtFpReIgjTmGbttLg1w20APNz6yZAxPth7yvJErasE
8/AoOT4nLCFEeEsWYJLERmbsOLubL9wNp/Q2EjXde34GojMHpnv53cJQhIoY
6yeLKLxI5+0SdIq/mLSU3vuQoBmrL+YkObVuJPy54uIgbOVfbQQWM48N2OmQ
DeCen54CrYcv6c2OaoXYeLXomP8B2WBi3ZE0w9wSjYgNOph3HFZQ14nK7tnH
MynfcORLehaCzdCzg+6WrIPBIue9Ve3uUbn+Huz1jJ/TFjSmrD8jUXJOypFB
AUM1MDtu/8UIrrEfY4XhckR1Alg7X+tyMVPnzv2KAuSg+N8zCIBKm8U+1R2e
M4eaKaVXU6yZ5VBfUA+WHxHKMUU8ioXOC9m5DiHlbFp1aiTiARa+hbpNAlbD
Xn22ltTuk4WdfSoH7pKwcRIMgAOyEX6lretF62ZN9J3nzwlggv/uAlSkzKRu
9KgxI7wAYAYhgmoVVVEgBz86unhjdxmj99HjACcTGhafloQ58+WdJ+UX0N/K
dOjEeYlFOQIiMv811Nekaur1RdnQK8+wo2wiZXOOcTDnHmTnjOApcc4Meh38
qQ4+U8o7niNYkHRSnpZ/wvG9HO+8lVcnUTdrN1UIwIZvFEjx1+ZhKcTPxrh+
WWYmDzVNAdj5tCN+wclD6Hx4C5vESFpdwyT0zuQHVMT8Ii3WJxk/7x+iSHes
gZfHAb9ce0qpAn+8Fl9QaUfwXbk7UiG0gNUePD0aTX5u3yIRYe5Xyp871tgQ
2CXthQ8YmdG789edTEBfEfkMpsWESs4RGUxQhZmknC8sZTqxFY+/VwjqeCCg
50Z4ydZW5g3evNFfShGfiyOGoFVybqyuutULEMf+Bsa/4I6j2AhNjuc8957j
MH3/UiVHAF4qNu1PyAU8PXjCcG/LWqOlPtsLy3GijSmPRKzc8trKjOzPAU/0
z2Ex5Ja4x006g6EvQsbkccC/tahOP3rmuTakX7V6IpsKGu4yFiCPUznxqfhe
kVBJzWJPnaYDnC7ap3j0r4/fjDR0YvvM1IDxTqdWCq3mtZPrC6RO6CdRQVzI
QLlRDCSKPrK6GkHqq4i3uB2f9NqKo3T1Efj5n3ebzRRsQ9lEPw8YKVfYTQ3S
pRPrzernTLA2pWi7a6lu1Mn2ceQcvdlFRfZVLT1eYeBl1xeW1pc25Xp82y3z
8bSdxbNRY/rViePxGD5lZJFlw47mYm61/GbmLJe9rWvCMRvzGWkVb385ar+5
2J0ehreHSuXlRYovwr/ZeZKSJBDsXqWdzPpFzE5IpNYWtyH7l6KzYBe5P7n8
duQ5GWfYRhCJFd/oj3OgXnqjZv4gTFyWfSmOfqZki8yF35tnle6SBE0OLzjV
ct95t7z3K7K4AFHM7ShqwtYlWGaqBXzLHRK+JTmKchTdp3QiRN8FJFzT+evJ
GirAyKEjOnmSUG9XRnTXSljuIbKd5Wq8uz7kkUDzHRqb5wGY5DYtV89q4Gaa
JopyDGxOkdDpH2JRaaSlqL814jFnfFGi2YJyRPiitASSrxfSZVJblYPWJf7X
zsv40pBayXXMD2SF7fndNqHWItOBKaVvuv/Y9zda+gkkqjgQ/yX1Fpl0YCao
h0w0R7SGgQ4BGNYwKURtD6GA4Jr3I+Ma2m+mEdO1LGtHp4HdKD3jYFjh93jy
GJfmPdwTyDT2pGMCP6FtE802xvNhBv8k/3Dsk4QcpOHF97NBM52WFEk2bWhQ
yhr5xLuOg2A6qwVT1dvPCuqCy2xQfqX+5dWfNgzDLwkBlIPXLhZ5Ywi5uA1s
v1IU/knvu9Hb0sC78PMSzl1os75z5aNhsJR9vGnmrpbZDldnyO2dJu1kjLQY
+KjPnY9fcB3Ji6ljCAz/9d+JHNidSQ4G93+fEm2eNP5wUMubn3KgxH4l19fd
g2WpSKmDnsflH/ZF1rwJLgDTV4xBiXt8qkLUdrXmxmsFtxI5Oqd1/h7XHvyc
p4hmVOI4SL8IXcG0IRYBO/jiXYDXmkKncRVbAzGQSBW1tzawm0snolN9zDco
x9WRf8vVhOxukb9BUBO6SDYn7u+BnAqD0gMgfEg6BASdPnaQfUMpqPswrVOF
niGGWPl60LPCEkkxuvPiv6lBWziLArxpr77UyktzGBTtDAA96yP8hAGQkpzg
A9BJMd+3pjl2Kn00iPYxGqp6TPcbdu6e4TQ+oROGhUBCYn9Rxh5izplWq1at
L7bLmYjUK/bKsZat4qCI3Ftj/JX9uKkzYQNxKsMH/I+CJ6PwGQuj9COb3ljm
a9KDhpLbgzuUv7TLD1ybmdUwmMh0eltiM35yrVW3teNNMAkwEPb2dvXamuHa
XdSh98haWSG5hNNSh+nkorRyyX3FQUYyU3Y9sAx6Com52tpAs3lzTtBj6Iao
oB30nWUo/IPNH0hPoPtjfw9wK+TfpbO9QSysyuu+kuhtz9ZXse4EsadxPiCA
919niwNtGrL3xaVCbkIdyR9WA63SXI78VsZUV6orCXoYClW9Qq65TOr4TaNU
mc1D6Kq/DP8+CFsk2rnYZ9oFI+JBG9u4JghyIZAJuVOuBOP4xSRH6gfSTVN3
TVz38PN4PwUJu8szPbxpVu/mWVmvZBqDqw9ODRBl5ucFCGdciWW0gkbjv1YP
G31w+SYxXJNOeKpxfcK3j6/d1Xg0glQnO1vdY6BsML5m817uARa9Ft9dnKzn
5y3KbtquIWow+97jpcFTxhDXgBiip+FNf6mVBazFeL+wbPulL/pHSjx8WyXx
bX916gGGLnMvdigCTqcgGi4DPcZskfi2+MTB69cMsRErmCpYq0BEcAeFOL9c
p+O2JyqZMuLSzEW++bDPd8fuxU+nf8rM0rEa54AS96DRBMmuyZ+PycVBDKG0
0Mu17U9/AfUD812kJVcJmclP9ZRne52S8FET0OsleMHUor5YzsnXLW1Qq5Zi
21NOuroW9vu8HGmJnmsXGgUkwrJnGdyGPdDcQDfwnNburu9guTAiNkcNrvIN
aKCEuVwBHIhp14sx6DeYWtKLSkJLmGPCVW1ZiIXrW7EhW34iU0UPoSkOzjZA
g5f3Oz6yxsMo34pb2wfRp282EcwpaOjhXoZtpd3TBm/3nFhb8HeUmArIhdoQ
RkM8zjGaBcwoKW9Y5a1k35nFt+A3iqnJeIcYaRxwIdG1n+y5WDERAjWo9Dxc
0aBSTrvOpu4wqeARULtzDOmjIFy8d/IEynfYie9dq/KjgT+YwYWP3nGk6IIC
UHUgqBBl23+B3MPGQX7EuEzyaLC3zj7jiLdorx9sBFXLOLmje1LEeo2QTF29
iI3XhvqsGOc7ukRXGzPFn8mz8Vsry9yHHjqLD7neDlWu1DVl4szKHTcEY5HA
WRl+wCSP1T+sHJ4ytWrOUubRDbTCHsAzsGAzad0LjOT5BTxdUqCSSwsf+gfq
g7v/LE2N0aopbYLgoKjMLVNjIQtzPbzQPSmWU/NiLSAVyGY9JixVi16BMcLd
18bvbhnjdkIALtqILnJt0xNgjX6Lt1HxEGIvXi7zhjf7LlKTnln9+ZtGClfz
enBffNVzrGa9XmLJm5Nb+VREY2S/w+qGprtTEXLbyeUUk3z7joa+N3WT7uCX
rn4u5/rX227aT0MP5fnUsNBlTOgEqwflywgwuyL3JACV5KMHX3EQSMqmcn/p
BNyccxEHslTOdQ9/a5pzWHejpWAt2RABtEhuQG5GGrJmBuhg7Momw60qWOpQ
Rpb+95fxqrMZsD0ZBj/0J8WOonBON0Ftjd70fjMHRlF9aNlz3Uq2gHQyNHXa
yK+7vQQwvURbHllkcDD1mmYfQH9KWOC1NbYxozB1++83m+mdx9LqW/mAFH4V
uCiE8petclOYKOqIMx6xsofA2nEgnCDYXDoyYw7ue7r53OO/wpprxwhjF3TF
7nhSZdJJX8l9gfwD8wqdmahdlhWfeKi/WCFVSvznMnD9NEYgyf7YnPVVkNwK
W7fD00wQQKrhUsowsOpkCqn/0yD17CKKBGHCzKMhaeypXvHNXjDTx4YtGgjC
76A5a4l8Q2ftF6mR3G/Ziy2DEtiS7I/1+26JG1L8HtmzSgPQVHrbxf3VfYgI
C4C12Lu06kHJZKl1cQ8MIj+soTLetvaRsu5eDW0Nmlzu8k5R1GJJJGZzlLa2
1Rx5gf80Kjmx0MgHJHGEMqj5n5vniKDo3SrKIakGQ797NbWsHenOc/jDNiyW
Vvr+S/fIF+HKv2swzagk5B4+uQn6cHZdNkKYKQKCXRKwQm8sL5GPebml+zFb
wUNyuA3VCEmGBWbVco9hk2+CKhvN46eUjECMqNJpiHI7rMOeX7lkzjQ+stGz
qoM823DgpnS/8ERuquLQqv6eCOYn4qmUTHeS5mqhjMFxetfa6C7pQ12YjJ1N
HR5ifmzapo9uTZADcx+FwuasS6Drg2LH/2Jq+pCbumYVufvBv0uJrzrvbxo2
pRezXf9+ei5uEdkqC8Cb/GZuoV2R0FnvHK/TE+JMgVU+9uHONJgaX3jWwQ3X
uOCcq9iBgWILdjAKzuHIw6JimTo9ZvP9Cx6CPCWpF2O1MHZY7b8BnCv2cSaa
T+YrWc0ezYxWRWOKq8jtB4icwfluSD4pZeMumDFs5rdjbbI3jgylI72PPlMF
AnSBGFQkxDmLWrG48HxmpNIUXJLqXyGcT9E4IeT/ODYc8RKMZgP0We2dccsa
d6tCWLoza/HyXpcRs+Rq05qLAUi5qsuw2Ek5ESnaCvLQvv5Nh+6UMqaqWq5G
x8/x7aMmlF6mSQT3c6UOrWy3bNXaYvN5Khl6/woAiZjOse0TU7ehps2uib4q
e6rv1ps/4dRsQG7m4nkZybAsxJnYSRH5ZMcOkNCzW6FHiAzpfbglRr30a1rR
jWtndpWzlD0o/+MQgq46sNlkA4UySaEWzDWGrN1lIuIRo6h+MqB5TCxaArVz
Xlu9DoSFwohOOWnaKGNpySE6tZEZJ0JUSLiOV4O822uVG9otAIR980pWr+xe
tIB97zD0OksR41WxstqyiBtrcoCIP1CT1icVfTWlYMVH03aR5Y+Y1P/tTvcx
CY1ARUra8hMApnQniI2LXlxUnBcU7fWFixSDyXHxbDFo9lZ1ogbzZPOeMFrl
3QQEwq4bMFfTjuJdaVBcnK/Qh00w8JxwB1rGnuH0Zv3yR3w1DKrQkzH/tRkJ
y/Lsmirx518aXVN4h9QvWkJ6Foc0maOVssMOAOlOkvFSvnRiPFH8ElUcOpAh
QE7KNenC/CENccWE6au+4y8hAE+TpJE4UlAIwdzIHYpIJK7hGBxX5wJp5tsj
PC48YfZb6J8D33CAufNMv8gJejZxt7Q5Tz0V80EvxGNxQIK5fy9v/6P6Uz88
XOjY38tsT7R3xVa5p/OvDHiC3IngpA4tcH2d5xUvuXlHH+BgZyYYB4E8tvcV
n64KtzinfaWhM7XoHdoyVVPCTFaC9k6a0R3dG51CiNZbHHwqH9Lj/zGdVn2Q
AdaGfIO/1eoIMUtOsCinD0OK3zQH0dSjkGjAwcdM6WWE/l/Lp6qgWvvwIaLN
pKJyC5r+rrWCYy/jdDdYDxMEV1/QBei+vNsWMYEpYZdQXnlfk2iWS9wumEHK
aalYIPaTCoMVxTarY8p/X+hMHlGS7ef+xui7kF6at9T9O04r9Wew9kM0rZ8i
GbAFtuGmguOtSbEYwEaqYChqLn59Tvn1gIdUV+KC1TZSiasJjV/YYuhR2+EV
U9CMq3r5X3QLHR2uoiJaO37wyi1Vx05T4H75Lqp9jQB8RN/KV05NSxxEtqr6
a500ICx03Zu9UhFbXFwh8ltMd1HICn02aEuDZud+W2kWhyJeXlsEf+WoQvWG
S0DVL9QunDBFacOleoCGdoKOrue13A73f7+chzNaXWvQXMAQXN3RczgtBYHG
HJSneU9k8ycFca0sVvrbpjYdALRNWX5wx/EkEPIentmmxLaD6rVJ6tq95AgI
LRp6uYMBeb869wTXR/d/HOsvIiFb0d7c+xZd2Irk8E9P/AwSrBDE8pieBDTe
cF7y6ix8LuaDfmfn+kUAzAo2K0SVey6+J4GzCk0kwz97dtuAYnZ+lugKgWsK
H5zTQJ1oIMCgpcwZxYGUVBeiHH+SSdDPQlU+AqV5ZOllhUq0jkt4RUNUN7dE
Xnw3oJ9GCDaNrTHXI3mcXtFQ2PjeETzNmcDu/Ah752P6Gv7IPTHkU6YzEmiR
D2e6/TgNF3NCmOT01HNLhhJ5++tCBTY01Y41NULl65S3rdUUfW2nzW8wGFwb
ik/KArr5LBC6BtQQZgynUvEy/tQe6Ez2FI4WtQ8O3xlSkXVD51zY74NmE8+L
ivrD/LrraJ8Q5OFOwyvZl/hq8JPTTZ+YvCDvwg0DCjpz7oeXRZbv7Oxnot/1
rBscL2SFSh18VBNZv+OFiMA09h66qohcvP8iU5tKZBkWTGTA8eMifAfj1c60
i12BcfSd3G3oRCu6ohwFXDuIfAS0bAhxLsszrCn8o/fngaVdSdc2/Ox/37ut
Xic0GHueShFcu2KPzxiNGEr+d2inCf60rfZgOPMUqxu7WmYgDnw8XwYiryDa
d7mXZj6ac9mUDP8qP6sgbhmtVZ2f9PupfFxhDRxeG4LxovZMPw4sVvF8LNer
8CRvS13xBZcveT7/SSZMUSCmz1G725xqjqSbgyRJGiv5BOkx+ZYirfQx2aoj
8LwI0os1K7gInhEtLLF8rXSegjdOhlu7rmgV+jneQWrdpCLKwT+/INEsDnZR
73fe/Oc+2wNUO5akplzLpfbCl3uSfIj6CUC0rYYD6SUcqhmdz8AbnlA3GKJ4
eBjXQ7/Jc3HOC7QWjs11l1jxmVrrGWCYNv0NDFlL3i8nRUOx+eHNM9pMbv24
rY4Vm2acPRDXwog2L/0QWBsb1lsfIGM9H0vum08LoaEEuNK/mzes/3t05Egv
7KbDHSwhpFXj51Py+CIDl8J0F9RPab8cCN2kJWBkg/2Vub9oEndBQ50QmsZU
kSQLPJYO0Ued3eJZkVHvgQBYHhDX7408qcADAfbPueyEhvmHDTQCA7J6o2XT
W/vvnUtku8ZslFQ4vgrdt8XoWPTQ6lKJfFvN4zP5cc+9PIVT6vUohVqSr718
C/XLZ3v19n8zBVOBy2SDVSQ65DTa30ArpVac6FHM7LNRse0KEIAs6sp9qE+i
OUBj8sjrgHXyU1LiQOn0l2t/F9/2q9gB/jeDS1t3Yn8Kjy/3kGhjuMT5dZJ4
7jo3GoKZVW3gHQ2LY53gXwFRidiua0f0cAa9AXFM5S4cTb84l2QzRGfgb6l0
0wnWPbSBP6pwjgjAA+y4vnw/KWaDm/lN1I8iEp9wd8FKBkGKRe1PNkgO0XqA
Iiqurhg9RDuX/Ny/31e8ih+e2PF4cCnuPfNk5hWC9GbuTeDGpY3VgAU//EuR
1gWi5HEqiJ2bS7WYbm70gFTU7Pdvqkf7KhiiyiUf52CkEr94eJPuZkr9XsAQ
JcH9dQILXEBHMPKU7rQIQazHY42JAxiaFXmYr3aYbAnJ0M5bJyv7hmwQdnhi
n4fSlvt0G6MO1stONKat5Itj8MrFtgMLL/AiZmTKN37m9aEChaTdbPW8PcmF
3xwf+PIjFikJvo0VgfU7KOVCW9M1aiGMqtv9b/gMgeWDFrwBtfsx+mIA//Ts
8cB8AekPKKQ58zRLGGqTPJe/qrdiSl6LXOcg3WVRYagDoxABHPnbYkWGGHER
V0C6BGSMhOj3XAVy/Zikjv9ld1CQFdg93X4sZg1a8eMbrXVnM1TpP4zHGdgh
yDznlItScLDs8XedinrzNpFOygUB6PFloPrfESYEPvn48M6Zg9osSPDBXoT8
t1B+bx21L2wT2Vg4pjzFuxrR6XjeTmAVMuZJ23zrPpnCilbycfJZaz3adnHI
w7jUTxtYA5c6Dbo1R9/nNHaGLwC7jKx2lh4eC8tRf1G/hvTU91Jc92KvjMFP
sM8YJKS1uFDmjgITk+JYoxEY3Sm7IoB4UN2PLBwChid4e2FgtRGelIJPu72q
yunU9bnzfnNH/F3hWQHJuFSXPytqhh1k++j85ydkRSfah6HgVZaG4JMZGAQx
EdMbzUwndchsCKEKe/gTYQbAiI59jEb5XK7iTNr3c2Vkn0Kg1QDWXYeaBPfC
qFyIucCklKRzJwreMkVswlSqdQI8z1DiyTAAIj6kFhq9dQ+o+n8FQX4fjFPr
YFh3oESYGxGUL/zHZruAMEjsRkCEMlQOeVdhWume3NJM3pJybOjxM8MoyBHq
vcKZjhTgEVnwJ/YDfn9XDCBQK5Qn7FxHGGb4lpa8xfHhlJBizV7DeFV5G4Of
sDw9OXC5u32kV1zcVYs8ohAZJxzK7tOILH6tV/pcCh9tsGOjDqihGULm9ZhV
K+8zNT28OZoQFBENcDjqoOqQzPcWxn7oG28moelbsLuGSEpN1ovtook/xLl1
pKd2tQ/RfBKkctQCZqOmeAHyY6y1ysK0PsSm5g1Xl4k2z9tqgc5VLQqVTn6c
7en6dY1TINA1CokFViz+z6xopjF+6/oRi89N7UvmoE49SS2If4hFCQ/yGyKt
H3dhaniMaDNeovsNmQSnsnLG7u2dBhMD6WQZLRmcqBChkaNMuY0/tLsFhQOp
fe5PJQK3gS4n/1XVm1XaAv6NnAxmRyVeMaPEHVcXjwYLhfQ+Biys8lgQT8FP
2ku6Es5/67zBsNUajfiyjeXkRw87lmJLG9wPvn2sr/SaDAvykCnxzDbUKwr9
6VS0SsjnbttbI4bd920r47fe8aMBXd10wCsqNUVSq/L0O1zPf7sp/MqiGpbH
Bh68KKIh8x7+/9kE9kRG5hVGQUpkQ1PVhexEWOUXNfsmjkjn8Xiq+L02ZSjc
RnSG4o3Jx5cS5egFE+J/vhI16z/H/OFFvqL796OvUULiZyb2/8QKsqDbLuWM
jm0gy5v6uhRhCpEKSRiJKj3oG8DJ5yF+VuuIyvILFnm1ef/rAoI3iy8onKwp
C23kqD7i99xkZIPc3TOadpR6LO/X8C0Mpc0zcXck/9zemcjURLKNxhnZKfnz
rgrwtecGkJzdCdrvp7JNfSh6ojnedhW0Hn5ZCmrEzxoda2U36ctcpshviNtx
gC4jCAaL/9o+hAtXBDBqUZMVrS4IC6oJPuriAO3TI6RHOsn578a7rOE4rJRe
6SG9wgiIicl2efd7Pc8/PwjzjXKjAZ87yuhi9R7VC8jeDN720QF30F70d5n9
CmtZZAbYoumD1trcSv+dOWWRnv9amwz9ao5j2mV75k1D9RZZR4vkjvgV7f7/
xD/EJJltzJixEUX7wGS/pVpMU5kYSgj/gXD7J6gfaslrOgBG1uKdzxfWg/uW
nGiW8JAnoDS9GVdR2JZ5lC0B3CT+5Kj3YuZf6kzANppoHmpWx9R4h4mXpvK+
X4X548RXP5qcZlj2+NfelpLmarQLGb1UNNalIZxakF7hXDmodBSz0iPaHGCJ
J8IpEmiiF0DFqotigUI2NM4J0R+u38YkOYeD2iUziVJIbLWKOkmE3FN5qS28
Fr0gLL+xNIxVd+1S1Jr/V3yO0gJeGy8U8wQNZgyt1QXKdIezzEpGx3oWiWvV
idZHMz7VG8YWaGWAB8qyROKdUSvIxuMsIjT8OhhJsG+u2sIq3E5bqqkPtrl/
8WRvc6WE9tWE+sY9aGgXLQ5jTMpEM+YJefVCGKF9L7rlkdtRqYV6KZ5pAHy5
n69qLMvgjeWdUNY5l+Ntatq5u2u1K0qwu8vuvUaAc2CewOtWpEjm/hgHMvjq
n82gChcCYgsNne84GwCtRCLowTF2d7SGe3Nv8THndUuFOsau0tYv2PRU5MT+
khtNnrGYznamel/kEmM31Ic/DvYpPjjKcOzgMw5nMm2391o75oxwmS0MvH/A
dU9ESmMmj2quUcGOW9E0NZNgqxeV4K0lqi/1aHflL4d+ik6ixn5yleb+wuQH
pttwA50KtxxgLLpVVHJPP7J9m5dTl8HfgTbDangu/R+qRXqASmB2xPnlta5W
+/jMj9edfSJMy0VcrBvWLvyaNamdo+JzuYevlpTgT/XG17H+YWcEkJ1a5H5N
pa0P1/LF14WafvEypIyGFUV8hK0HO3lBL8nGwKBOswnKB53QQWwIKrxJ1ozY
RQH2AQENKwsbD8UrWCqj1KeJX7MgBHvLTtvNbekV9ybEu2LzbwrU+ACcK8f7
aGA1B/QZ1XhneiV4aaxmoT0bt3Y46Vv/+KuS7WXXKT0GOrnNUw9cfNcj97Ub
dnnFGynySb7O9gENpSIJMMEYG5afo7NZOgS3iaWoUoKxpL1JAJrUCrYhwS+7
pOEY/vm+79ZtVASDmiP+lv8hayM4mpSQKaPzKsKsmzpF8f7Zweh79Z9izwTh
5HJHZ9N/h3gHLMM6fiDFepLixjVKPVDjWaV3R8eYOESILT0fNEDbVyOgmOMV
oroYaVbdj8RSA9VIISzevjBK+lAdOqx7pMTAQxxdNHNcjP043o6XVNpGKLZ/
+ryGAx7kLArThz+S04FcKJ6L9OJQP8gNd0iM4/Suf+QnxBqaETzwD513eeIY
3Sx8g6/p2O1lDQ74puJzZrhc6xukFJ3AUAbZbz6nkorEVl35nV7NH7zR24oa
5tCnweELRgODi8Uj7W26JiFtdsV9NI9HInRVHdIWsfxR4S9Meu0/MO4xXF7D
PKeuVT9KZWXDHYTiLip6sPpPu2hpVf1V29pQ/9n1Wm8AoQX2VAtjV5AkoBxI
rz/WeREOzpCi0toczxhc6pYiEJRIeHqnfR4TDKJjYge9ls8qEr3AKTbNKX+s
XKF3lzgvkNTTK7gj2UccpQEB8G48KgePGydd0aH8KFQpD5BxCOwh7nWRMJMU
iS32mWbOW2kxg2vkRt/QPjiTS72k35W81G3UYgrV4qWYRtMqG6eRSCQMeSgC
PzQMXzKM2lY+KmTJCwNfbGMENsOBo7MHXDQtp0HkmIayZdEQWEJF5y6dYgGt
AEyiRElSuo/n0jAdkC9tnMAP3W0hl3Xl64cB3FUvCS9a5mUd374CyXAXy95y
Q6bmpRttBahRJUV9XUaAHeeClG91VQcmxP8/BrmmtwMBw1f7iXBa1phWI1RB
mBb5HyQWBisDpJ4cOAJ3t6hVwhYORucJNu1iGN2EFN3TnAeqIzq8ljTejYkC
/CYZKrOxiA+p9UfS3Zbgemdrw8ybJ345rinRzWedvGb/ySur5BlJNfRuLDO1
kkPfdUkFI5VTWEu9D05FCVDc5LdO75AUwFenorYIJY+aa0qSjf5rDkw+VVc9
awFOXQqRILCEr9EvFgrLTq/9ZbcxAhNIxaREGcEib/rqzAKknDx6WpffId38
9Ei4Hfwb9JBOlG+jOtSvA7ggBKBlUzm7lRYB0X46/186TA9orDA9J7Poq6hd
DESk54v+J/hSnHxP8codXQdBsTHIqU931CZ52aAOsNz7th72MoKxB8vaFglV
1Kp/YDd8jKhNpEYF68jglZGxfTskF6RTFXsS88rvGCcuJ2xtWaCjAJ/ulUBG
lhmsvr1UtiE1FsifaMpqjbJCYdLxVubscJEMmXGvXc8OjjrXLPIa+hUKaOZb
+ZfIhY6gC8vK/lYsM9j9zEJytnsrZnAj4F4dLdMfiC1SSyvedetkDdZ2Vxby
8KbIpdcVw0QMYay+qQ6+WjOF/HwfjCO/cVAWBgv1b7MnH1uI4630z2rp6Ztb
Z20TflMxPMf8TweWqfZM06AKnl9y4np9FuSpDp7fk+6PDvKDof7GhR4lIEgh
/0EPpq8hhLJQptCfUcqQeE6WFsp25c+AV5BPzcgStuKHNf2zRQ25kKF6uG1g
hRUJHp0UrDAg3QhXCPRJtPq7qpFKdcJLTrqhM9tAnm+YrFWWLNr0pVmq4ra0
+muRvuDOf5INErOvNAy3cudnyIqKa9WhpUe4ojyRXYvsDOnp7dDFA85Um78N
vmy5UOq80W9uWRl5EPfNYqBMqK+u7FuxQlw4KpTs8DWBlah/6kFGzBIlw1Lg
2552zoS7PYsIE+cLsTEnmr/4iGCoYXXn+W0a75NGQM4bGPyvckYEXLRmdhc2
8nC6WU2jRuvvkQZ4plobcXfRJ8oOUfvmjYwYhGTcdEL+SnrCq8GTxvBZ9ZXL
qCII/C+9d1cmM1a6Yg6dGhYf5ZvjMaJ77V3NX3qGF4PmNiASiMAg1loXbjfZ
xPlabje9dIFOnWtdVV6jvys3f0Hc1g3yqgSGGsaB/Nbi8wAhmjQgNb2CeuND
SlxR2W0y8Guwfy6PdYv3Nl1lfF2BpEgKesNo66PuY7tLUP5q2prLs/OBQNJ4
2MfXSdA7fn2bitOIvlkgQcFWbjnf4mY/zb6X+0mGMUbXi8DBFD6GAGHWGFYv
CVbFQW+ZF0/AwWhwSCuohW1CFWf+bLXWLFRU/pswaoO+NhaDK+m5daezNK+G
bjaWK23BAAV51I89gNNYxEC7cyDpbSAZCjnFAoC+CeKX8sp9illt/Asvq/ab
Xd2irJnLaZQFEhU1v7mSCya7Tk2g6YCu7bFrz4XZFd0lSC9AC3LQZ7xqv0re
Z+nhhkvnULGRd7eNPLBnyAjcMZD9I6W3S1pjy4thiAmOdvQ7kV35rs1YEqK1
U6qyfONw3uPqbat5oLWJ2Stuq+48nYEZiVvsthMCkgMgJh7T1bE5whnsvvg4
3fGuvmJPyhl+cVX57UleGwq6mq6CSL3nySkkmIdu+HlP8LpLGCR42RKDi7HF
LRHJB+MganRiv7LJLopn3fsyhQHd6g2qieDyaf6LMFe77CQw84nDvnQX1eyk
iQ1L+nYhMkv88faKdz6aUPhPX6wV0ZjLcvrjWk4gHXUvtUGFOKcytuSheFEr
tIv/7mgPW6JI785RPDjsR1gZk5hrI7sU5hfE7/mxrS7Ip1G8FTOWPan7cL4X
yMO137OgKx0hKeBBpcwMuRDxUlZW7jPXl2j0wmavlOdirS6yupVtdicy7Ndp
7J38gJ2M4TtsUxn9p+sC+MYBe1yTTtCvMaLIZevwTi14YhLYSTvBxG6r5y50
jhVcnX1+7bA/mvdP0lWtXjFFkw3m1QulXYcf41S0oiTsRIpYDVi3eRCf+tHk
49XfakJtN017Y+T1V5NI/P2mPcJwBH09H72lRnXmij17nGA4E4CRHZTjLx/n
9Otq7cXTwciN0T7P/7Utq0TR0ALLDiFUVw23y+BQ60vMP0iVs1T9VXwuiGXY
7IqkWNTjjI6VtuAd+bwSk44i0GfNuccIg9QiyfmR0qDgFzRJQseRyHNThBy5
MaLba79BSjFouCKWbravPyjVDHpj33mpepDnA9CQU/PJ+amOv1hkocvAL68U
GK41fs5TtAaq+ZZGGCdMS6dZXNH1z9DdfmLBYlGfAPAxumPDX9AyFjYFKKNr
rW3Wpo5flIeQa2RflssPKfMWk+fE+W7iBcI8CGE4OZiWBEkUqVfjMFdg+Ygp
0U/mqA6QLST86TgKdKIc6pzohvFwzFAXBrrQIyIc2iv5pwYjwinPyZ8b+9Qb
bVH4ZsYQGPfVrDWr+CjRKABXiEv33kk0p04Jr5vcwKukV0//FONuUgdlUlxN
3PZJJtzk1Efr681cdPW1amFCav51np5SS+4/nahX3+X/gnrvCrvLgm/HqvnV
LnD+6IaEfkTjyDYuYu/TnSISWc+iXmxOhl57yieeLcyljBH5aseFtP6r/Def
ik6USEPnB4oBZ4XMaOOCDtjkIsP+xuE4SLqk/OGgPoYjcyQQ1ldVUs/U//40
v8fbg597689vg/q9XRbl8+uoVxEOMEDhlwYARHdHfutCrHyu9n/+9vpnldWs
SD5KQkNmylhywh3hlZvDHsva8jtIIfmDo2B+yQJVNsXieUSuF/aNPcAAQZTL
fy2UB/91iq9tYBI6UUt73t4gO1lLgX5s+nrnzThZyar6U25L7LezyQ3E7nsi
e7bjTVPa+i/8SYbHs+e1oJjV+fax63wN5oZqPwUTQZ0s8o1urfCdIsPTgTOW
j3rZntFOmBPBkVM8fHjpDUix10ijncVrLjetDng4GctRbxXR7r5Ro8b6Tyto
SNciwViYodlZP5pQx8Dzb+yGvModm5TLv35Rf0G3jShav1zQY/dHXJymWH3B
7ijFaIWTEpzM8ZfsXAXxLZ3blASjCCwjC6CoLwAf9d3wIlxgEMTFjcjxB0er
oxrPWiL2VHVoA9+NcR7lj6Vpfc7Ih8RrQ4VDRFALwFv+lZlCHIEP/kRN3njf
romSN/nOAOXPVyU/4nJ7AYH9a1RMzIbKXZqUhnRwIuyA/eCn1tfkDzKxcWrk
yFOEEGU5UTx2Je34fdw/NkVAlzKJrwCO+VHAJhhabAsbS0IlJ2l4kRyoPBkk
3G33ZdYUQF2fD6f9vew9CrxlXGPnD4hCIZaWbCVo1Bl9UD1SQM9KX9mkynZP
Xh/O1w3+wHvCrzkCNO/tBUhd9DkBSvGHpYhIQ5hL6RAgHikHZaZFmxifQo5E
4MS/ddQspbhokslcfF1tkPtZBbJMH7WbcGQ3zqNHG0kkCEGcptvCBA8XkqTs
RMk1OSA71jsHdOApTrPvXXjTLBlc1QwaTIN37ijNQL8pRPz59B2uhbdNYGI5
EqmtRIw5gAIwuIg+rb9eJ4n4iP7GAhpCGx0hgpgkjFyCNMMHyC+3HhnspnBo
eo/hahOpdGDBri/ZP42QVT+moQwUQ+73ps+7iaVGkh7MYRXDQwXmR8DuCMJM
Q3acbuL1ZFDZaVefBfJwD0Q8LthV1ZL4v3ahe1Scz6hB0lyAgq1oE8oZsvib
u7rB84FT1DmUFcI7Bpbw0XCURH5tHYoegDCAMDOKKni+lmIQHYM6B3pICAmh
MY3yh6ajQeF/P6ItHsDxpS9A+dKey0D20zhplr2YlRFPl6SJh4OM06gcTPPh
NhMEkR+lfUMOIggQGnpdDM27MyBs80STLySgAotHBs/dpHXman63VQFrdjWU
BWn6x6L+fHfsipKCvv/pP1S2YbVBEO5/uta4+YCqhFT5ee8QG6Lh/tiHbFV9
vdB28t533wW1Rx+2XSRs2g2bax6QvXwE8g2LpLx0lqlyuxYwb60QegUOg/o/
VlCnztbShTfD+nami/N4hVvsjZVz0DYkqbQolhUAXmvBQSjJb9Nc0gFZDk39
JRiXWo2hTZqdOYQrs3pyeHHocPGMilHu4dj+Ja9SziYa0q/hzv4jKQeJPnd0
IkyjskSeGQU8RjLilOp0r0cqeVo+ST0ZyPcVNKE9YbLt8jCmywds/6T4g/Q/
bTysXh9LDeICSBQ5wCnMsZbTeIammPV2y0qs0As/aXEQ0CBSkMjeHvwbncxy
kQyJoZcGJdCUdfVq+9DbpooebTDK6dY+twhv0ZK5WOK4YO5KrR3JbLx8t4WV
i9rL7oTi4PnEKDz9Yzqw+QHroAGkRcmNtXzGJfyrj1skidQTAuUTN2kQqjUR
n2Y4DwPgxFzZNz9RZRK5ns901fKUNNy/Ful9Q1j4W4CSrIFJSPbhrr8j1DMU
yIgTTFAadb5SZwmMDuTnu1oOrNVx7Gs63cVYw8K3VJg2hJgE07Pcj/MuywSl
c5tAq6Yu6nMJp6vuCAqj2obpue2lcR73AdwdqMciGZNZMQ1Wgrw8zKuE+UH9
AVfJ23nruSn08nRoA5o69m53a0/UP5cKknuA2LiB9MdNhZVdLDYLGaWHF5P4
FGIXkngOXfpU9hiGMDaCqavv/wFyd2oTVO0pwg52kp5EmW89djUWiLR2YPWN
7nxWpDIlb+5XfGivPrOZUsUBo76JaWoiCdjB8YBRFCFcc4BOZhqTNntEHpCP
ExNb415knUgmLz8MUBytA937gA9m5S9joVrNRWanQlRKAfbtLZAxXIntJYnY
3sOWnHKtQt07cjY3vIxLSEEyoeOShjghBcBrEfNVmqp2bHOvduJIJAJ3SAJz
gXOy1nS72GWL7X3aNhb/UoT5WtSUImIIGQlRMoAJlg32V2bb5y6nNQkGb1GE
CWQkTiAuQ42/WhSs+jIQb/wuSGCll/9VfRExGXeD8bthxselh/jz1ZvBA4SD
LIpsacECAx2qlzZGjJEfFFoScw5/kShFUuc6Fdc0eSyQD4Qp5tzEZhOPlnGJ
Bar+qBxkvxAhXLbsmiarhX4ak9skpdRmmCssDPXR0QQNZhTk2uGJzkAwO+K+
Jtx9xloB1xc7CKNY3+LUTAxlf11OLCT2t8zgDFodmB5qKkmvVpXPI2zHrYyW
wZp68OHzgSw8yBsTe1CNTQqg37+a6nIJDyLroI6PDhlOef8++gTAsAWJtlXz
IMbV31xw5ODOApWj0m64SRfTHPjZTbY+0LNGzgSbMa+OAUdHSNQw4ovcFJZb
/Z8/7PPIrgrQNbndehnsLXXBC2T90h5lSKFREoj6UDLY2igN/HZRAfJRD0o5
f/eXpZd+3bOUeaf7ADUI1yr26ednk7QeK38o7+61MEbtrkCxCnqjZNjy4FaN
dzNcbz8HJuqhpTovNURcxcxG6GKu+h7CWd5l3KdrUSM5o7O9DiKjarg0l8j8
Be5cp4+BN1RxsHhploARL+nNC7cWiiYJo9q9Ta0Jl6sWQU657CC7cempdcXy
ykfoRcasWcgnenWgkj+ooxJ6qhjwm/fRQR7yBPkwPBFCaOBCA7UWeIqkqbS9
pMRMYHbtXFWHwAcGZBnCJmdCPOP5jssqdnUX38rc418s6auRQmFthcKUF0+2
yJXuTCAIt4g+Y0LiWpD+hfHP3LG7Ffg3DesRA8SEOgAmVvQK3BmUUS7EMUv3
D40FOsJLAF7oSzs5h9IiAZ/4OHMmqn1+2Kn2O0WpzSupGADC2kDRYiJX42em
UT0zWyls8rwzifc9PIL581w4CaliGIyHk9DtUa9iTixH2Pd/esdTLUShj1ed
GbFfkV1EBgzblIvDQwoIsIQ3fANfJ1ySrDGffKo4d2/ns6JM60UEEW6SZcma
pnO6WRUREGIUKemD5G4H/c8iRvpnwSB5xK2Pz8A10zUM49J3fK8Oe0rGUH5N
i5UT0fvVCRDlMd2iV21gc8eP0kMwBX3i+Nq2v7NWLphEHBuFrVVkR1oF8hmt
qEPeDg9NUX41k/o+ZTnmp+tS1oRDLTJOhVhkUG/z7rvlxtBlPIATCoWL32B2
wXj6IoMFIEUpp3IU4XwbUKKW/wT/RhLXbR3e11HRWeF++mLXfEePxxAYdQpG
fWBm1xEkrFxyY+xETmhj8GArCCGmI6E/O165F2kiIVsCLDB3olLIDumaihYs
NBSJQQx3pC+wTMu2ODTQIkp5/n/HAymCd30T6m25Xh0LvFUhKEtDyw2hyQTQ
DsaCNr5Q5fwxuJVndoT6MfZxXHMi6OMEzfIHdx8qxg7gk9NZGADwCQQMG3Pf
X+yuCG1KQsHuMI+nEVAKx2VfibN+WggJGsvMu3MWY4qbbmygIWQxBGulw6d+
+VxLDJe+0osTd7HnPoihYAcCwx7cYSlYh6ZU57JGQLXhdN10TaOKvJN1+5+L
gWxVRAR7BwnzURkLwqUMpVZTMH87rVxYA6IaAi2qhvP3nlGDMsOZJSNRRSKs
ZaxbsMOXFPoUw0k4pRbEPM6/LgvAB84OSpPkVb6kTYPNLhl4c0wT2g8cFztI
WAqCoQWuVxUM+O+UprfJ8ZTfz7T5DmXwIg6YdPtgV9eCTmY3BToBL3WB2aNF
47M4j8CJdGKJYW1qu4cyW2nt9kZy8gsvrP01kSY7/N6MUr08OGCUjuEgNLcJ
i+2TNX9uEIrdC1N2/Hbpi76IOyaCiTS0wTZkSiEk4CXKx5FGAGgqgTpCDsPk
aRT50qXUy1ZyazG9DSDMdnAr1quCjxezBmiJqJVOeRrD6JrHr8Kv59iWwYuq
62X7Qzt3S/RWWMsLIyP1qrrmqtM/1D4d/bnyS7mvfilO1v+lTTTgxX/Qvi4t
RSH8E0xid1F6Ll4mtzMM+FNYAHz+0dNALlAbQSR1WeQSR8KNPuKX/B3VZk9o
KZBU2eJOjgnD8w9yc4Ja/jOUhmKUyrqXq2Auyk8hAruwYMVrcR/vGeCT8m9l
pvGj2CvouDge194A0aE7Ql4SwBDgpxrQaD5oy7E+2z38AAKMuix5C9v/Fz5r
T6RK5TQKlbpNkfIqBrjRuAdiERyRsHr9444sFG8/BMotcZ3GMsKtu8F9Q6NG
Q+vmWQrUOIEXWdrP2BhOIXGD20btkcCrr6L1/DLTTUtDfbLn+G7SCr4yUsWd
7eT2vkLwy9hhkV84mcZ3jima2GrM2JS+EJyiaXCCw6KQPGMFwbnW55kWmvrU
nn1ayid5Af1P0na1SWxSxcwPcd0+yYtw3JBIgCZIu4OULSJk3TbO0Fg6A+T1
ZAOaScJ6VbmhX3OiQt+2t6DP13jGcJt+7eusWDjoOcyDx+ZKxO4Y34NiIY7D
eqRs+2E1ePZWG27NoOQeRkT+bNYK8m5Mc0vvIZQiQlIYOyd5JD/xV+NWfD3k
vofKjTOO7+v2XQ5MbTYUYQgWjsA/P4Oftgdy+K58mbnUQaZ+vT5t431y1CPf
a8z3HuM5M11lsU3/uraWqtVHqGstncvIwZEMjUFMLhhRhC6YIkt7dsG+YXBJ
6kFl3xRgS+0utm/adqw2Cg3N3DK8bxtSuDM7plJWhG79s+L7vPfz9w9tuPPN
C2mJpyGOZm20A7XeJwuGhMfzqhMSDIAN5axZ0Z2cPEpieXF+E/3EpOFIMdC2
PF4o0X3uCMuAtzIpxrb2JSbMxmy7ZVhh3VpXkwB6Lp8KJc3zWRBeM/WmMonk
TX91A18Oezn7jR5tXc+Nv47B7fILHIeZQKT1I1t/q3rfrqg8jw9d4iyJIe0j
M+BrZlsnYylA+gIU7R4xRSeGgDvc2xffbM7HmoO40TtftDXu3D/Oha59fhOl
6v4mfQS4EQ+JocEfTjYZYuVrp1TY9Ajpr9wkGTFHrXjpHeMLZKk/1Ia7kCd3
hyPkfamWk4e6ilnr+mWLGy8+7wUF+DP0qHKjju7P4DOWH4aojuI2d6SmEQgO
hYkiD4C1O8LY3mBr5kXdz5pY+NDEuu+M/1b02J4plw/O0/93qXeIhlvAWW+j
6Fo4h3WKht0y1bBQf+wliSrEFVTwobwrTLbliOtUt2XtHZBr9GeK92fFylBR
OUajeTORo2/A38+uKHxu3rDtsT6L1gaOSKGyf8AfpUwBKS8M02BCcCWEU0/j
CLw3zDecaRMKvRZIrTBsQuPAQEc539GwVlAL24cq6ucQojH/lQI0tvu0I3lB
u8O68ycjfWhHwJulD8q8aGcrTt0bsMixWKuzJuRw1QlFbakTPkrMbQvZNOEE
JbrP+N9dlQfvRalP7DNbpAQCK0EYng+jbbLtiP8N+4NGxqXC5w1ynna7IEnC
s1dkXlKkAEb+Gr2K9HbfMZzuJGCt4PHgN5U80MwGbXTamu+G0bHDiV//q5NP
FeUxsFPFSwkPXRnagYVgebOFlyltnq8prhVTbhH9W43Z7XDQuGpa0YfE9Xmj
dGPnmiQgZbOBVWix7ATtIz7QjqyqcB8pCdPnkEQ67DcdB32QkMg0zysfClQR
gz6WTdlTMVtCVaEp3EjN89pLTSjfuNWx0BFnLCCOz3CPkaGwqPmrsK24C1HS
XkKSbKuOwimkyGCShTS7cXiPL0pklGW5VYm1iZjCUh4hw6tZd+u0x6iMw1oM
JDgTfi8UNEtF2kj9KhVCOMKE6hQ8qh8PDw8ZkusHOXgWxnkovQ/lSOeZYZUj
FKw1QjHwQe2K7YCf1nNN7dVPCXAfSkLHWtd5X4/HK8/pdtAkEFJYYLblkjJ/
1J+YJQMNXxa5tO81Er4QHnEeASP2yssfH1GtBySBiuMcuRlM7yM4lWmV/hyl
VyWytxRBbCt0MZdpjJdl3CztrM8/FYN1MlFvTKTswyt3XiRe2trJxkkW44ub
pkTFwmPT6rnF/O1Q9hHaH42TxilqKKArtBENl/xMJ5s8MmK2FPHWvAdHSJlk
AmwE0REFjkMIWemq4kxoIf462h3cysBA7UWe6YxpcKEkhym8Q0IljIfcp9s2
wsFonVdt0wRcGlwt1DmNZGp2C3XDnng98g9JsY68yB8IdI+V4UyRJBjV+RRx
R6wmCcqDN0ReFT7CHjzhamimJJQm6cUkj0dF8CZb9g5LMdGKKsHp3Bl55pnM
X2f8RozfJWa/ViWmrtJe8OXZZT6RQbqeIL7ID8n18EMgs2CKEBnGC8iJLQ2l
uMb0wxM5Dh+1YLHf6hAGTQXkgLb0LhyS9kLh4p91DeoZrppNTbha3xOXGmU/
AK7iO0O9gnt1ptg/6/pxHxJlznLYf8znpBa+FF1Hm1TZVey4QD8zx0ojvMwR
CPgbr9FV1AWWeoH+0Tzycq/RUvef584xV68kxyCVOWOb1zi0W2lL/z8ATHqJ
3/gPUSEqNtdmEYnKFbwYII79JAvbXW1VRpQH00O4TH4xdjLbSj3anBCLNknF
t8QYq/zTVB2Xp80WhKyENXTf9uXPzqwCDBL6s2XFECPp4cxzI9S5DJokl+m+
qNBSZcROrn0hCPcpIZd8dlOddT7UmEOdp6fksIA08AVtqkDOsrp6mye5ckXU
UOS5EGNGf/dtEfoWkpU9urF9lV309xGZjJIa9apaDwIxEKUsb4RyH7FCbU1e
++R9HTrOs75LLCE4quoDUGZi/PVN48Bh7MX7qV6KemSUHSUQyA90AgzDqgu+
i5XrSQv+0hOsZdKZAitlUS0kt18KAP/OVKp4OVmqmvm8SYmftH73+hbLGdsf
YBz9FCryflXFjPOh6nCZNrc8fP+B+oETyz+tfLSvyEuFbX1jRu5T+GyvSBzh
tmNNPiuzgVXC/mhLe2hDPTN4OiKGOUK3FJsCJsCnlsyeOuXQNrb3VnYkl3RF
ieaZAItrUnjfP/xAvChtol06aEaepChRw6bBY97sccnnYL4dgg5mmKLI2AY9
J2ao/BeZgtzkxxshymc2XdbYg768OI4ydFxtV5cGXXEa3J6ghwBLiCUBFWrh
g9O13OoPxdpQiG6c5iNSaj3pT2KpV/L94GGmuUWUQud/ZXsBO2nIJC0VUbbF
2muNE0kRSJoPApdXi9wZrCLKGWnHVVMCBBAO3OvtEzVYNoiC/rFl34jTjgp7
ihXM2g1QyLK2J358vvOqoE3cFdUOIC7QiQpr73QQFpuaH23XFWjh2bl26scT
N8Uhd4en7MURriBbyaIbqYF696EAhNOT1zyX2oXr08TqQiNQJ+FfGGWVnz+G
hiT8Wd2XaSAeFufG1JJ0VxgblLzn1GX/0O5mIVdoIkbc9GUKaqR6ET8RXia6
CjzDm1a4FUfGUiB4FEnWCRhqLdtY6RHde9t3EG1EaqzVxY/tyIUb98gVfb9a
dA4t7q77rqA5uFdhXB5CZauJAF4Y3lB10hIn7dYWQP8AuTAQKOBOcR/uMAbK
UkcgIUl0kDUY0lUcsuT96NIxDAPsXXDT5unjNiRfUHlD+jtzW1+YixCcYlUP
iZbAckuWc1YPFsszWUl1mXERAyi7tnOJHpl0oFRflKCcXWmRASbcrkB34OQE
pOUAr7CY04sWqYgLoiyXK/mOMRaw+t6/lnK43bMh/MuA3u8zefIPR1nSqEX0
NPYTTpZUfnSVQ8P6R7ZblQVbjfFOkvcU44B6YqUIMIMiZugqwF51pood2Zk6
Mve87jDeqc+VuBvxNgHKY7YCSOuuUf74BW9Vy7fAs6UOa3Y2i+esniEcRI2H
Tu8E6mZtxi46WddsCyC2MTl/SqR8YTzTZ4ZZ2PD7B4yaVA4Z3ZBZyssApB0O
yMO1j29sQFpzFLX5qKVxwYvXJD4Ip+OqMviCwhsbLlhiLz5pCZDl+TEUvKkV
fXnzXt9oBWzNSEwE06sJ/oFezrUpgE4YlXfSOiGCFQKt63D2+i2Ki744oV/y
tYODm5Ipy/ZBt1XGOtM9uf1/2B0/y2eQ9d30wSLp7ktWwG6Lij86gZ1M87lC
Po0cVGcmpEpJJB/cYS6/+mem53JhTsmaIucPHCu0sQZYOtV9a5rJkHO3Dt3g
62zaRhSvxyXZs5NOYC7l68prEZHhBiOhQVRSDIhvy3vsMaeDhGwxz9/Km0HC
kj1AFNxnSDErwYgt8BO4ijgt8N151aftLN/xJWwav8P2pEwLoDh1mSSXsTvU
GTnArlztaKAw7+pHg5lILjeHkNnjELh4IE6jpFEv51+PBxXqPY98VUoHSeLG
0djDkUBf8pMouvztUn5YmJaMedSVId1PKfP7e2lqCNJWzsogaXvIV3fiVXY6
XiGegLQveOiSrFbBdFwtVDcypRMuiSl+4k/oJd6/cTuPtP1XioV72XtckK22
4xVCT+hqqztFnO+uRM5HENwcLF80xYyXXUDP4l90zrVjHKGYBjUyxZE+buSP
GBFWwSp9nUXMwt3TUjkvqimjUy1+JF/oLPADkDUCp6EJncCEJLJbPLQDXOEz
mx46wRakzAN0SJm9wdZxiTFMnvQHkQq0bYGkuae0DtC40P8pSY+08tErJfuR
KREZDybp1JmIRqOsPKH703TIvx72xheBKEwU8frcxfhp4MK4f76ds+3oipwF
irPrFL3464ZU0aG3Nd1Tm519h1Gs5JwmeFvhyVKJGHvxEmjp6Kszmhzq+R7c
ulAoH6QaXs600CNGWqM6/jYBJ6d2StIBiHTa8vcZDeoeb9XEvMdEt4lAWcRk
1Ln14jX5Uo1bj5HZjPJh+iVFdDjtlm1ePp0wX/eTbi7rwrwcpPpMY7385D1b
it6f4Rkk6aznXLZMhJANB6EMrYXrghS2KV5424XaeLn243Kl+EvvqPcM0qSp
HIsapAny/D5fepKCDg+W5xO+XV2SYOBMP2w2XvkEpi6VC1LOpEn7K0vVPCLZ
fCtz2OhcN1T+h5v7MI6OtKaBWdU/lzOz5cdyWU28euL2xOGmVWm4ZLKKAWMy
Hv9IMu5SEaCJzj9YZdYyf2Np2nzBuFlF27tj8/G50HRU0Ig8zG8k6oP6+OCn
L0f0EXpAyjVj3RN/GClVkaN+Qvq4T6h9CeV6xJv7iftLafeisVp20NO/7P0k
gbtoMiABMuqx2e3k3X/myqhq8Frj8IaKd7SP55TJE0EtcY9st1nnOWc6XXDx
BLmFeP52BTSP3w17YqOBbUZh7483Ga8FfHR/vC5IGee4IqR2pON8CUk4u9Lt
Ye5dD2rNTor6HVagcunpjNa92uPaT1FkjsLFQ2mOmYyyKouwBIHx8sMgp7g5
S+1XfIaXqxcYLUCAm/mg4G1kmz8QySX1rmkmH0XUfHapALLJsHgCF5WJOjPs
RV4fYZ2C7Ps+/3VAeCpxn464anfSC55YqVKrPPEQSYCsOZZk75XVg6JVsRcN
HnUVZs8L8KjxM25QVzP4z9Ot83dOVURZbEBLylXBrXcegWli3fUM22sjujEZ
CFfOPrtii0NlKxmlMb8IMvPBriw6cZtkZmzumeWvtGb3Q6alUnhinfXMrGUP
OKq1fxV5sPnpFvG01Cjdr/t9eMwk8Hc+72uQZyhlwbkQifWSRWa3hzVZqPu1
5WYh88Pfmj5qdToIALJVCMC6ciZNujKTvQF8xvt3mefBPFtnUv5QTyXwUhPb
6UvTCv1h/peHZ8KCRNMry5I5kJmkxOGM1dTs+ks4UdxJlJpXMsaMqCWV9Ano
WlkhucWbFH3mSR/e/hNHNTeKmmwzupkuGYSbRbW5LmJn0eee2fBlDun+NV+r
A7ztmQh+FzCywg/68aR+1ZA9fcB040D5m8nBLCbvtSoVSAa0HIfUl59ToBf0
RemH0t2wdoBwWjggmh1W/gjdo/dszqjLrdX/ux3o1K3AAGUJF7qAFixS797L
aUFQl2Ijf8db4PlGeqevu2u2HZrUomy6cFdNYX9GUEPdrV7fzJHoY8eIu6ls
8bRsvii4eJkJ4h2gWErMwQgEgbbwrgaZYbY34k6JvDOfmGKWbgiDMpbrlnYD
mGw+GwHEHmc6DTiaNH8FwuCMcaveE+VBd3tTHHxVoSp6ko1sfvb4e49kT0ey
pfdaxm75qW5CWu4d2mKKcc+QP+QsMX9jOCPlQSP0xJh0FJ/skmI4WHvuB7uB
DU59Miaje7bDOEI2KlaUBFX+gkSMM+Y7wFqXPcYXrtroYmsHEFZ5Dxyf8EJU
8Ms/2Gac1AkyRMe9GNq4/rMhJhJ/sagEFnY4bI/eCXz/l8otPbK4dJPn+TMK
9oGJHjVDs6v0ZDHWU/kUHxPmf0X0YHovmMf2YUNMjMfdwu2ttKISvVKq6wKg
Pj3ZjwragZviuSzeCByi1AdgS89B55O7Ri8CB8LXSSV7ycZUB5kZRPzM3kmL
MrQZgYZUHKOaqxGa6O6/8bq1n1NHP25RqyE7+eZ6fbWzE0U+hFSJygdAI5nU
DTeUsz4h4O8HTp1/P28awYr49NdMdNPcP2ZvIOrbxNh0+Qd31OljnouN8Lr/
YTa1tbhYWHsx0zZVwhfoBWQE1cJ8Td69UL+qQD5ewTeN8GfqB89SJzsN9r+e
KKkcDKcwVi638Uf02FjuzpqqHVIKaOefDje0x/naCUhQoZVglgx32Sa6lixJ
Vn2djtAyGr286RenrkTVI3eaiDRCzivyMHNdQroJPyRSvEVe/yygoUmWNHGD
Mbx74N8pnxzJUuYx8sgbLWxfeLjnJCm5pIgKL+JyBmQEBYshNTNr2JoiJAGW
4LvPJ7v8qC3a1xNV07H/0OnKqsJivNtiKF/AtOWzdjGzewrQzP6BPXLT7IOW
uG1UbBeKRvQc34uf/xtoSCQHM32uT3917LLheND5KvUqBdmIOWX3JQCGeWW9
Q6Tt7DK6rbjUm+cKdS6c7Q639kPXJEqbgCkRrDWtEG09/x+kvJKaY7B3Dyaq
gqgAnpaXluy6icp46ZGSHZBjMPLz5wq1STOrkpR2P+yrblT/DsxpXRBdyRlC
iOVRuML8NeaAY9inxLVzzw3BL+clhRC+h0LtCzGJyWMhActheoMj66F12c2q
V9JOweAJ47WOA3QMcfo8S7XNBVlbbP9VYLJJ0iWLtUXFYIlqzmrTJnmRsGvb
jTjGWC6rXlaMdXKKLUs9hK3PedVml0oe18XG3y165POYptZTZW2ROsgq5bYO
TKkwoF8rSQG9/POcZfwDvEC6VBeCBYqoiV/v6wcB6DLVMS+zYsCK9oE9liTw
3x7EboJtfqPE0yeOZ2ialQ8OM/XZ2JRyK5OVnRAE6RiOTU2tnT7mWQV1ZC7F
4Eg4BZLkmsrDEb0kiI0jjiJU1VvVsDCkFBe+kniD9AY15GFZE0ekEIm4cz9O
sRJNuD7Cp9eAE3Fkr/D084sjkfZ+UibkYGQYSU08DSJpzNmHIQVJYdRcrRcz
RxxccbMD4aPuXgKT4j1vmt862IgLu4NYv/wPR8C6HEJHziwnEAfSCT3lnlxP
KvFiOI2QsdCNiW3qk8/F0w8Ox5oiG70m0H/5zllEvXnzGiv48ofrTHFMtHBO
ABzu+gfhAPXnzSpoEv8+rFQYuXdf7Vz1owElEedtKS9NRNNJmtjEDwY+imNq
nx6/X6pOj58STRoDDzPX4ZEj01WcX17JEZ28xim0R8Cx3XdJk8SXkNkChGNQ
Z/jiUkeulfFIAZfz+3qhUw6U++DRoDrPOXvF6BL3Q05Atu6/9Or/8CGxQIHd
S1y+L8OpCih+Y5CDWke3XL/Zf7BSQiWWiExSrSjDSb04Jjs2YfI7MyW2bPs9
9Hyf4VhNy5oviYjmWkHq2qUTpFsepmjm2Io7rrdve5vnzSb9bO26odaJYWoD
S4bt+9aahExBliYQy+MeBJo7dZEjgc8pgVr/AHBirnc6DDUULHN9XdRXQ6wU
ZDrNJe+yTOv7rQ/tkrUOENbNxUSII9oYNWZWodNzb7DKb2FFTh+3C1BxRAjY
ty0Tg5fr8vRYt4OIWoSgZPt8Y0QLa45sXqYPQsn2MN0Tk4EG9T664/TLtdnj
5uSCYPVSqN7bN+kjUQTFALN90PIyFpgQPinB2N/2G/4gO2op/M4f7l4/JSTM
dW/pphCvmM928RxLiB6eK3TZwSnCxzZimDw4ZAyPvHmFDRNlTBhma5//ogpj
rxayuNINMnRZkL5xeXgAPXr3mPuMY5vEiKB5iRjWE1xs5zbgDNf8zk9cWDxl
CQVLGYpchGdd/5SHQ2MLjvocxylFk3YSQ5ZwoR34F67XENmKFNe0/lEn290O
Lbv5EMHk+Svrj0VLY7oa+0p25wo8O+2v+gpm6EHpjjPiSInvEUESdekdn5ct
SqP/cIQAOenT6El51nzrL39HFLwIPyuL7G+jyulrFL/hs75TyxRi20vRd9Dw
3IMt9+iZtZpynNo/RYxJlfjL6pjk1pLHtmRU2xdrfTRPPR7COjKuqa38slPm
g+UCncXHGWqdYoJaJOYp47YWKt09W0m99q+L5yP+23Wk5MJ6F8/1VzEeJw7D
y2sa8aBv/fFspZNhPwy5d/v+N+O9nUzS5I1MOv1oSTiLgifVYcGhfP9f8Qgh
VNyR+IZKgbHT2jCO6zIkYEfKU/NmgvgBp+f8oK/od7We850iIFVfrJdpivn9
Oi4ZN2faN8vTSSKo6Sd5xuaNEpBcZWT088YTI5jOGke0/Yjm1h4fxO2D39uq
pR56Q4r5mpPgJJ3nK50OLrVRAbid+tWvZFgTs/cCB1R4im2AKkjpymMcNDnx
WJMCJeqRXfnI6b6cFWAFsqDWBJqU54RG36g2yq7QknrxNqJ3x7bC6Z29/Yw6
RGWhYq6ETLJyketlC6FLP/HnMnOtS3pVUNhHme670Q7wyfdkjD43KfQtHZbH
3IeOQTKjpa+lhGnpaC2Y6b+/oURHIAbsHO6z6dwxIiWx8YGjofZKAWUXvSQ0
hWDt63zRgNgJDwE+z6vHbS9qY9rkkY3IfD5OerwPShBMAACzuz5Wy8FUyUgu
GMtsWlmf8fzDnTNMcvffPJXKxKvLtpyi2z1DNvMn/ZsAZpOHbe61BkhIYZF9
bwLYGLDVEJtbdAr33yvMrXThYw9iZhsfEzcpfH7SNhcnRTcO2SPKe4I+y/ua
vLKLEOt6VkYSBC/Eyba77jazgoG6WCGw7jOBHPJVq9wyGG7W4oG0lUZerwdE
CGi7BYsjbdiPGbqFz9H/NTIiGH+UsvZrZjfq0TisXGNQpaINm//MgP6ixNAV
KBcuV3WIG+2DJRYHBlhNbxCb2Q62AKzEp7yOnF49jZmtcNbOcqq8Og+MqeU2
Wl2HwPnmoeLz6+6K3fr6EkmCoDqflSy+vnwGXGwnIcLK/5C58nvcQVscSOwK
9o75ukdXA+wwdjS+ihcZxA3kOIEBrynUeJx14/1bWmcrDHWbjpxX7KyUT+eM
DAYpkU80EI8FQ3kSf1bIAPW9jDxt/ZwppOnUpFt/deb7UUy/GeyiyO5t76X7
OoLqdqIiJYqiAZ2cfPAwq+Zisz5KsIoT9qTAJCNFBJTNrmQc8zvBw7dzUYhK
pItj/3J1217KKZn9IRxktJXK/zE6X7zGftP8S5qrEAmjXwelONMmi74SbRpS
sUchQBi5iFeu1996ZFkVRDuk8mGeGqsXMVhr5OmOfTKRyN3sSuR+IXqa4EaE
iOmndtayV/mnTJNXaYY+Je7n5kl4YF8WOvF0qwIXRoXxgPYjDptvfKpCrfhV
5kqKKDj9qTMAPbtoauLa/egMcBTZh3dm5JBbuTv070UZZXKEeeoLJ1podm8O
710Ae+D1+2Rt7DYZ/LbjpxluIed1NP4Snf2e9FxLJ0a/Kd6fcuLAwZyeVp2o
jEK+JCBehL6lvpHMz4InyFphLMk8nWSvXEbUQna6HOviELERRIR44Dk3Pxaw
4J2s1azgk/OrZNChGb70tD8SM0+MyfxiX9Nuy0RUWl9JgTEn91WbPT4A25oZ
UrPTsVopsB1SPLJg54mPplj6S7rgySuLn1EESJsnxttuICyN+87OLt95wQE+
gKsQh5YdQiMmAZwKIs9H5l7rNeF6B1HSraW6mcFFRDQgmpi4kQlCPeTSfMVh
wD8eIekzfp1aAAuVgugwEPjWWhNM3h4+QsBXbx5jv9+tpO4wvD/RkTyqu48E
FCng74TOJr/W7H3fVerIy7uYC6U5eoyzJ9fKPQOZZ1oExL/AnbZcQ4nGhEM0
2UyL4uED+i9Df1S+S6h5pywuYFoFnZKPIy0e9dyVQwn7kYvGBZRIJN5MIbGL
M1gfB+0qiU6PwI9NmvuSACPNJNrfMIvHte9BNuVRxrLiInylMR6GvoxeQwWq
WR/Q+tegfDk4px1fkQ+3K3cgMQmtLin61Ua6rDH8BYT8pYhCCqV6DU6BhGKV
Wg9uwitXEFDbNZ9UvnJRzwi1brEn/CLZTkioyDZbfkwF56Am1qlf8BpDOaIL
dA1kQ4PmhS6LzilU8BmZfj17WhlwTf3nYoadQFYvmMn6t/nYUVGR56gL/FcF
u8nd8fEPnUB1I9CepWXvxKUIUnoWYXm8pnBBCbYicIw/2TiI78XcRnEICP+9
wlu1iP7U35OZ08qPEVfmH+smmEFN9Uj360tSgpsmF8RmX4skGvNuo+jtVF9S
T1NW4pxXQWxG4blcq4r1c4zcQFpL7jysonW0T0EFjv1HwwmQimJ+pHg97Iki
me91Ckpgu+9I0cjBxe7jshtrofiIMQ6fzFGqgiW01waNGSGXWOoFCfJVWMEh
Z8NOSWKFnMxM1xDEGwkd8jkeMgZ64PSG9O2Wdd8x7NUgb2FjxCFLGFgm3SLj
5eatM9JJ5NkiAkw3Yu+huqnwUbZ4ca7KsnXBSSv+TuVEjADxRUQaQIuwMEmH
qly05Q317Pu4ToSAKp8tz6rPOBg71cniCRlp67bCZ9oVn0fALp5jX+clAXuo
8ghgKUpSpAJw3z9yPCiF2v3Mpbd+2MyRJFral+l0C2AlO6aULRoFSzb/5nId
YXv47myvSEDr6HuVxHBVT03Prdp4hHcKS0Q1w6ZFwzVSjhEH2p2OPTP32Uyz
QiRkw4mPVp/rDV2HtubKb82RM0Hz4m/YXR9IbNMtoyBYo8hEGilu3hay7cIa
oo1brnsk3SkKK7UzRsEWjApik/L3DM4O0OsWau6yJSa24UqtmlIno7+BffGX
BO4prAUT4zqBKJvBHbAywycMXKStnoykmhP5hHOQZ1XFAseQ5g1v0cGn0Ng3
3Fg95x+eWCvj3fJP2J4YY0OeLy3bPJ9b66uX4zwcQ1Hm4RUAZSuZWHtgQa/L
mCIdyeEgglebKhZpcH2U4oaGF8nNw8+EB9hTz/IPFe8KATB5E/DjsxT2TH+M
Uxuqbb9XwLzd41YDsDlLX08g81/pjZXYwEhBcCo6OplizcLt0QF9Vrj1sRE6
NoJeAEVGXqbfihM475e8BORYiySPeKJ7lB8aAJ3ezUHyWW7Du773V2vwQkuR
ZdoBPl4ocWFa+RY2t/cDrp9csO0gBigiLfcNg1hDoWBUEZ4KxU6X7exJ+4Tz
6Hu9UgUMJH+L7GFJbx0SJlJe69gG5EcNFibOwPrjQPxGKC8d3OEH3KQQIWqu
FCKjOKZMnovLQ9rIB5AOw4XyOrIL1uWx+2+zaUfVypA1RXCdbWgp8dRAfe/i
0EqREegOHYDL2TTe7nW79NpkQqnNTQvTwNkDho72SFOyJj4bIdv/ikVpyQGN
XLkQfNmglWf44XfGRFYPyRzOfg7cTJTrEo9KT5VBRvj4A/00Z1vLO9edLoY1
gCMnBw+gtua88nM+++HNEGejDLDxR6Y6SPSz2q9+YMoHZfY/+z1gE3C9kxeY
c3H++Tya1/Dbj8EWvt7VK8pl7Sultwt9qc+tP1tqHq2KB3bMcR9MXJdQgqDZ
2YACaG3Mm+RIs7dBrXVym6Cfxo9Bt32CAnynBsQAZzfK3OZFaLlZmzp72zUP
gzeJ8BTNMkUgm8RxZ0PGLAFzfcBUwiPFTTVnmTNQI/7rWH83S66wug+SmjjT
oLfp0ih9EJebePjoes6WvKTRnwjRQIgeBs7SHK5urKoPVswZZqSTgtipo6Qi
DzACGzxeOlQXZXhVjX/LQu17H/suMxq6HfF1LGLmYQaUZ7ZajtGygj99opwW
AF62xVP9SXay8D1+NiQTnbJKYn0BuxnlopOH+Bq6wW5QlJu6LDReD+HlawAO
7TfflnfcHiZCkXvq9cqq19+7BpujjamB7ZsJ3pOvpLpMv7eX+aTZ9xkTiM+M
wtdHkx6YJpNUpO51y+mgx1L1fjlwV/bfqneyRjpVKpkMhMeH29qxDaFMvouS
f3jQm1/CEE8PyqRggfkvspOwRLRM+CWDeBDPriv6u4euvq6DW9Oq97bjE9rK
i5ZmVymcu3uPPSaxqE7gs4yHiiQK/wHppRkccahNUgmLV/xYMnu8lrRgAfqd
nshMzEfCJRLg9WsHz0cR1v83IQU7q10INY98/Pe/ORH0Xthj91UlTwSop+5O
XHtwRwV36qlW3LUmc230mJnGfhxnlYEmgy1zWfFrNFQ83vYxGj/k4BxkzZbJ
jmXUYsvY8jqf4bXY5CptdsV320Q2Ng7OxVE4Es5jf1Hc3iB0HPxR8ryAt4cT
laZd4aJ1y7q4p0fZbJwnNSgbdXs3ryxbrQlIgXf7XSO+/VYxR3Xz/y0JyOmz
zBN62myznsToX9PUY/CG/R8iX35WVwpjsqdisCx+h0ydMs6eQtY4EGekGXJw
S9PYgHwL3gwY63CsOZFi1Nm+EUXrY8vyDaJnm4zatOtT/KpAsK83M+mAdUnq
9GvqZ/+mTHg2yU8RQWVJo4RARKRMBdarCTLL2JjuymcnqCuOo9dMrZOTrrx2
pv0fYdG3r1vlHUO0iRdJMNNlA7T4C96OyOn4+jXzuJ3i1/V79PhkpXSrg7qA
WXCRwmyPJl5dXz1skxnyTUSunIMlcPJ/WoinjhrZlMKTwejFD5YMJNX5Hy72
gM9fUpQ53J3WIDsiwasUfyMesWn1OVUVQVmyf8D82nz20zUelF2N+XqoDOva
6dbFy1337ssREIMQaDwTA9R7J+TtSXd5VhSIsTBirCAgdmTAZXrkANh0iTku
QD+Sp92jJXpyMixsoyN6pKZ2xTr2LVj7+ggs/2Y+OLfTPNnOldjHl8fKByRQ
LDopSQkHonmTpMtytV3eU2ou8qgNiLLGr+6hgVex9igfzxJLMSVcVpQ0W1mF
TLfzuLcInXd6pTgGVpM0lHqUpPrKMi2VBa87GQ87Rxp0Ek298qkN+dPDc1Ta
U2nGATL29QzOB5Z/YN6eKANvnpMsRHDwWXFvNlvRMOSXSYl/B52JIZoYUAja
9D/nflFc40FzZtK+ACfNKkSGdqlswF7kDoVehIptBTaUyzJlKT6A1pCyt0a4
oUtHb1Yc17I0KDzVl7jUCVJyK4j7JXmetdoYBz8214+gQuHwlJ7Et2xpnHV+
UpCTSzMUreSGzlUrAhw/cj9lCV/IkVnrv/62irpLFam7tQq23lcqr/XzhofO
zMMzPTY0DCqnPYcxThg80H2urm8RAbav8SBGJ7ivf4E1/wPiPYNjqTsC/P8P
eihwnFdtSirydMwIK9KgfzAJjYX35U56ba5R+6MHyDGXtqEmS5F63Mm7QO3x
D61GgHF7PpLIEnsAO+HY1wPIv94QldkqpUte2bJXYeFQbHTzuvGRoWxCSl1d
uqw7q1AmZh6a4LccMq1Wi4mePthdgChCzL/sh56CMaaCgGh0Af9nhZjChFqi
tgvCt2REwGXIzxBx6mWeO4gddmoDJfZXW4NhBSD60jlPHgN9NY8h8LQfYUJO
gwe0D+n03/ciSBo3qWaDXQKeYBvCoO0JCAZmzt9pNs3f4/GCgsn1FJ727WNh
rMFJXqqyuBoH4UnhHTxcPWkwbrFT11q2AmSGSTyqNqdQxUoAzq7yWJEu87pb
pa4lagO/EsJSF8G4njko/eToJhsujatry09+hkd013Gwv3nLx6MVHVqgZzK7
tqspvCeoRf3G+w4fVRz8weGbXQGr5lk81bnh4O2dkg9VLYmRBhC4sSfu1tzH
doMizpQrzO/IhtfueO8W1pOq+CtQvBLZS7EhD0KWc+nxHBLrZ85NVFzAhLX6
Hb7LPpVHNf8aAjS5p0L1VPtgDZZ4Pzgnp2dfmjQAJYbKmpivS4+aVN/k8Ihn
A35B9rzJNElsUpsHg3yShoe2ZpEl4QYn7WTYLFfEPqJflq+Zd2u9+MzbQjCc
AZr/sUHf/unM0CGti6MXxbg7ijG/sr0Gk1XQ8rvkzPqwDT5WyKt+x2XCBf6k
+sls2F9pbmx+PyaaTEZEbnWI5BbrT4j3phTkSucDBpHA+USDUWmtkJjiSYh8
o5FSdmpkYjpvpgbeIKH3t+L2xWBLk5gxwAluLpMnMPg8qph7H0BGtL84mbMg
NVXCLjeFi98NGnNtk2uA8ICtOjwWAoFSd3SgIyFoxTmMVNhzC2HsDTXOsFEK
hB9eHJ48vx0p7TaWsqRsoF19zLz2zCBAtBfhAXo1xtpVEFlPjAEkWXjT+Vyg
/lkndmTyP21jmyrwe0usAdZEFro+0Mk6Qbh8DvA6YcskNHjSgIhOmgksG9T0
swFByWkYynI5lw0kUXP87qSG5gNb4gjQfnzdCLAbAO6QroF8qPMJh6u7a2r1
uKQBdXFIq/40+exAo/Hcwtotz7wQVeLowlmsNalN1QhTiJa2XtI0UVtbL5QS
adR8qryaBKppZC4R/EKH0eRBfAhnhx+Pcm8IrhQcQvQHN8tiAROXiw8kwIbp
l7fMHdr4FZo+KI83QmCfNLuHWiVztIX+mmy8Kit6k/6173t9daZjYEmZ7rgT
0I/TNL7c7M7HFw03eJDcvE/f341YDx2ssj6DX2SEmZ1VjI5TaihNAVxecjPY
cOdIZMP3l/BqtS7ulF8J2aJ69kUNXhAqhGzAGu+a4cIJwUe25XJeD5cke2Vt
rc33Rr+oyChGbyF+7t8UTAzjl950MM4nQ57LO9iFeaGAd31N1+EafwlzJXO8
XI3rnjJBYtRbEBzRjR4d5b5HfKHtI8CED9xLxb0NoppygkJFBazVmqnRtUhn
bED1xX22J0zaIWRu0fuEGIFV9hEIuLJhgTIk5WiFWvT3T40GIJpkw4usvu1q
qsQCjCLqsJ8IaBai6JX26tj7OP2dLcbO4gW79ztiSKoW/lGs9qYbiZinKX4s
wAUu3F9e4Rk0DcKMHd6oHyf/KegRr7nsPFyElw96jR0+9p4hbgAjt+GXBovc
mVboiuRCBSlbbXodSXvwvw/nWaFs7I4lkrbrBHImPWTJtiSKkUg6gg4eNw/p
jgH71hwdJMdE7sVzK7DF0tVhp+lgUCJlG92+3jNXHamDJv2U/XQFyEOV1W98
wEDGSmQURnRqRHhNUNswmCMi/6V3PRlPtyFDY2N/YAp/pnhCclsmiV8+S8RB
6gbKNu5Mz56Yx0e/385hLuoWiyNdP59/NLXhcfsbvIM68GhQ4CU7Lk/Alce1
SBxwUsTFFslz7hbv99jznYvj5zsNA4uNwLcFBKGUqZjIlPKY7s1GfNL9q1O8
uUdtyToY9mLa84wtxyo5UGSs0c0nhwKiew/0LJnYvbh0Em7jEaSaqidndBrW
ddqbG1zGpCt4JhW7HlzOaj58BnGWitBrRDBLv8EYqcIfXq2FEOakG1xtHoG6
GTqk4Y7kMOzSYLSPd2SM9mWG0bgiF7q2/4pcOmtDv6Jx0rFV/KqOFi4emdgW
nlx5pWyvZdMYNyMyXB6xHW3bvpx4Fm/apTtyk/6Q1r+TjeAe4AEqbSFa5RyJ
3SRqfOPdVTpdWNMVf4FeU7LW/dMSyQlYpRq3Lbu5JiTPgM3LOylVRwylPkKQ
EGQg+8n5Fbb5PdlWSWmeo9b03ai7ej1NCenDFg1cpVwKNql7qp3ON7dijCjY
5feNZ+rqBRrlgjVaMkLZySYgDDUqCIuVh+DmJLo11h5RTRjBB91cANBV6EPl
H7L+3RxOVRIHOPDDQHqd74C0omrRRkqKgZeaaYjHmHD01AYrd5A3MmNvvOhv
zw6xxEMnkRddPCo7Qks/K5/xZ0sJdsg8XVDAlwKhBEY0U31a9D2Q/7BJgk+D
nITMcQc1ZxGdFvEcL7ToStpoe8wkLlnfvmfwBcDf9wy6k+/b5/qaTPbO3o9a
g5eRfAbej1tCNgUCrb9XtWE3svKAegLzir9TMrSMKPOM0VIJt5d764O/QjJz
cLiELxjGewts7HndWBH/8Jp8ZityQVFQnk+DWijGSrbmuwAPDsuBAaFcmI2a
gSU05hmpC57uzeC38a5AdVjs4WJQYzJRXukcJ+o93BhtbLSkALnOKZCnBIve
Cfk0Vu+BbiaHKYWisHIwtMNj9RjtPRgGtyAKTiI79FaTmGKlvfr0Mmkammwy
YGhG32utLRHfGFsiBLxtmGoxq8GraIuPUPZ/Dhb96O+HPbalLhCdy4yI9SK5
ckZWGJTW2yW1xxaLS4j6i9YSlru8j6PwjMMCJeYfwCuWjeUrnW954vSxACYa
UqtOmK57TbkCRjjlyyYG/44fBUZ8NPKgK9bsignvqBXa73GszJtc/vu+1j6m
wst89cNceQn8Me0poeo6H9dyqaazjMrqqf+5b5W0IYgR6IPRqTkRro09ncwW
j308pKT8hjpBHTc0C2QmCy1jfeJZu5E63H49HFTZcrx0xho3kIQR8FhL+Fx+
vZpnoC4V8xfmIVAh8LcfWeoG/2tS2RAspWmNzrV9VdcwQut/0F1lhgOabbIL
1vbQsvCeOott+1h4/mPIlGua4Wq8btqgqYKOReaYWZZCE6hFE/vUk9u45zAb
65g7bnqm9CIE0uh2J1oMOdJpjv9xbJeHNi/1FsBOq2VOC8kRI/e+4GSxuxse
a5uQQVA48QR8teaR3OPKK1WEMlUVRmxNbR7dcivb0pbYy5L2RTfe0IffZEVw
NInuXJptecg5p/WuyvKSy1/1rK+/dwQ+rmDrpnTx9/3cVJsdAciHib577Vpk
mK9N+hpFnakl2RLYy6t9ixBe0bvCVrmzH0iy1oEMhcTF2t4NRisam9c+pipz
aUOC5qGWRcStmcNUgH4dH+bcoxhAx7zXPHhqK2xSpI+1lm1R6SSprop1NjZV
4sAPgZTdcWXTlCcHDatWYUE6fk7QaGiY00T0EmIvvZfzQK87aNOcKCWISNhh
LjhvL7FAUA5FIEP9bj5v3KOJJpIj3wrAq5YysQPq4qH64ic45zUtEsO36Wzv
veyOtbtgGmRYZv7NvRsSr9avEfvxvi89ma/+j8QdbL9IgqUzrbB3WqCznMWW
PxVatHfHZ5gpe1vHapwkhGfOkXV+A49xr+bGfuyOlmDJ6RfRGm6GLZlbxUgf
dC+vdyXLEHz4OY1T+kBFZ/caPcFDSX0jN/nZLl/bJjiFDXIDnbT+0nVaxW+O
p7/6839zBlZvehdpuQ5qc4KreL8dWcNYIft+FfHUYJnQCDVt3D6F2DhKXS0g
YS4dH7QrezMAskzIbxC9c72K5ZCqCx3wL3E/HPR25lm6JpKhXqBtKCtECf+Y
RAk54bj87zvhzS/DfVE5yNG2JcS6u3mAqtkjZkQZqtiNXI6Qr+kq0UTgIaju
5NQlUzc8FoyY5t4GHanU7+3A1eGWD6JPXg6EsAkzpmM/vu4SxykhOXITtPMg
k9K2ZpAlj3r6h19vMRxP2FXmmknIguLDnZL2CImsaQE6MouYtAztuIDstSrQ
pcFS1K2SMF8qMUg1NBrt+47uTjIEf0mdyiBWY5oZ375zM3TSmnYDeXD2vkCV
0GrCMYI+F7xnGNC6IHh6ZRISPbN2q1vybnQIY7wmQsoeRFX19hB016CLdt7g
SXVhfNbAvjqqBNOi7oSCTsyeFUXvEwRGX2Bxg2BPQv0w1JZ0LTsCAbzW0lA/
A3c+Y3mmAlVPvSL6ozTDUYlbLD198C8BgggTV/y/CiGlCKYU9BmScvWQ30zV
A1vs/xzpFnZV/o+WOZcBoyvYvLCUdG7h6bCeCmHrWrbjFuKJB9NE/bIbUkkv
FbpY3u7YpLSl/RJvuhQ1fciH15+meDYShjOT5vBlFijIdxYck6wljO448CKv
653NFZEA3eL+9FzSwVZl1wgE72HAdkZK8wB9bG3aFAjF8TyCIfNlaZsR2bXr
OsC61eMBobk6A7+wBuxlx/qLbvW+++Q3Pij+n0EFQDynaXeJTO3GHO3hGwUD
LtHq5eBUlHmoKWN9c0mxhyrj9V8IW3+wRB1FYUQXDIVeOxIQSRp9ec6gamfc
aDdY/SmJi/FN+3piT0iBFJmEJhf/3B7QfNBikWlnXlSDHYmhz7F5sfco05a+
94oWSMVXccaRSBAsCyFc6/ggrZ+9DL+/FV+TEgJli9qG6QhVHQObdcNsl02C
75WTBbvjm9BLEMYSO37nCaUJTe/DfQLJKG7ao2UZlrWgrAOn+LzsxPGcP8cD
tQPKT4YIHcIaY2XodsTq810X6eJqfWkQ9fCEPYox3WbSCMpAZfX2GEGCjbTj
P+G5zSIUqRbUSenHvk0E86Q8mzgcq5dUTx/bSgv7MMOD/0+KVkACnVUPqver
tjgdzl++gqb1f5vHlPx1vW0dVN5b/lGkRGQm8rzweAohSbJYRxAohkgW7dQJ
TbQKq10Oyc+O7PRCAiC//3VTZXU+kv+2IqZWlaOVceyjhfbqB8ctgnfe86O+
v9O54lT6/cy0Gcr1NYiCKA1oXpwXQ+lgj3f2k8Yh2SByQMvUqwMnsGAU/i9k
DnWZQMrdxj3zRNaiULqf0R7eavqUCE/XOG1MTFUwnMIKGIlVvKM7BmbnXAUE
ca2NSrXf1KFcPd6ixMJb3b3RQbMDfYriWxVjMAj7iKzU4yxRDEon0xdd2dkU
oXxWMxbyDVrfr2cK/Z+2w74ot7v1hCyHfDHaBVa2FYnyZRcwB2c9iOC5qYnG
elF1w9wiRAhk9W7kExgpDdwXjurIkCYmU6zvMdZ/TbMpEjSX49e39RBPIRK4
cZ3sr0MQlM6iDG2SLSLH1t9ZCVGJ+IMSsCbiQ6bfr6iGS+jBhYTwy9cuKJKk
DYBjRohGhOcaxKxFA1SBYPWz6YN0CjGciSM3gtAcyvr2Gd/wS/JzPedvcSKl
UsmMy9mSPn2sVpZlabMReuq1WRNiwGO86KxXuEexT2r8NmzRIRndne9LOeVc
Ovyhy3qy+VrsHKRG94CHMxtctkkj5wRO5+oEFma7GgrRm/S7Tt9WO4qwzpsi
R/JXlK/tqXsVTEnw6Cew7arRGNVmaf+GUdsqjImVpnFipe1SkNAU/nYgPPqt
mSTKZtB4KpZSlCAvyIctQOIcrR2JnLe4etfhvprsRfGNnGU9gEWWAoVsmctk
DInOYjBlxzeb/qy48VugEBaxpMP3hYYh1dXbB2mNm+7MY9rgNVE4YMeOrQ28
i/16VSLk2gqX3uuzjJi+e93iVAroMLXy4qkgHnLztsgm0KbetrEqDcQUnlEV
5AgQCBIBNjgS9sVTOWlu0s7d3NYCII9GBvjo9iyY6sz+UlGkUzCFIwD7IyBa
64zYTbAEJFtqSqeXsH1/IhDx3V1tSLcD0VnTYsHLM4tNZysUQYI9z1PfSvxz
ieDcLV7KeUQAcNBIHd41C9enDMLezK5GgOMjr6vVUAdf0+gU/nFZUAyutrDa
uaF4z+KvA2DJf25h24z1DAI/XawTxsbNqIr5SNKkqOa7SUgBEH0z6vuZqcZ1
CAzub2kqGETsvT781rPzQUqn6GZaPnUDul77oPvuTNAI5ipeMsoTJTMWf4d/
ziHbkZs47YUxQad/LT22wOORaFASYlRSk4dc82R+hdJBYMwtVi7Q76eKB/60
kbOUuWgpBBn3tk2w8TfHZLVZQBnVLQ2e+WdxcQUdvKNsqRvBVG0xn7lzlbYq
vlYY0v0ctOIjsMTnqzSLKNthi0H4o51UOYk5WdhUnqWrd7AH7XiR90a39jyC
XGsvgc7tt8Mcf8E1AP0TP5cuak1UCZQg84txCqhYJyutSWGGXnlXEsKSszCU
qHLhNvNPHXnqm1eq9YcxbG1WQGZeiX3stLmEomjHZwlhjgQayXBmQSTZeMMG
LjO9/eeB3og/2jbJfH++a8LyPwexwCSM0PiCSPx9GpkAp0vOUExwPSBzdSdW
kK4REt2iprCcVVZBv2bMosvfXRy9o2ztrI2MIGS2HtlsLwDbZPdim40idaVp
azaQZzFNLIiEg9ZpOUvEfVc6apUSCv8SmTh3oU6B4cV//fhSThLZ0dymbiqD
4N821Hz9d97SlXcomm3uKn8BqD+LdZl0fIRBYSC8SfVfUXGJuh7kwOHiDPmm
CWxawHu8/apJrxmdsIhpZovYBgzZovpF5hfTBAQcifCE/tCJJdboqrbRzAQk
RHc823T9wBNpbdHrh3XmefCTGM/20wbxSw2F3qlX/9xpSjHi5AbpE4iIgpWf
he8HCrrkftW6T1UHcE6gPHqWvlaAFY0M+5AK5eU7dNnOEv73ivgQdak97cZY
yFQGqGovVMdub4lsjKaK0wR2VJWDDNjXu9L0BLuBbb0paCPP/V2TezVNo7lj
br3LNN0t3cCA7MLkCVDU1ncFy/ahnKLK6kMMtUOTubxI/ofJB2zVfEo4QW2k
eW+jV1MxE4MbmV0n2WN5hqyk+CLKLYIv45/2DO/+WdylWPwlVy+01m9Mtriw
+0O9Gxuxv/3qaBD040OwkgaVecJkuMTLi6n0FXSbe0geMtGKaMYM1puUaxmi
mkI8U7XbbRjdGZQzOfsenSEZt6UV4htz8m+DfCVe9zsaSSsOFctYhgySGtKu
889J3I1uDGHoH+isZgGzMhvHg931Hbeq/SV/YG3E4u9+qKKQk8w58YLR6rva
S8ncHjohf/9GVO4j64i7Ic1WFZXdZLTK1sniNEJlvYSjtvupwM4pbdjmfa+J
cdUiAkJtxOsGppxxCo+/BUdVfrsFbbKQUuztpc1pn/QZB78Ta0UUxJMqGbKv
9Uq9bmB1ccOh3TGcP8uTcpMAhrazuCN6dexushcj3tzI/cN2+gHj9gkI75qd
Ya3QjDk4owA+KCsWMB+xrCFnvPPJEj31iezSmkPB37y+puu1RwtKJVpu8o4q
O1nmlNIU2zFd06VkhklqmOKiXdTVcfUt7VC4bdwF/j1shaA6Yh26ufpYXe4z
INwEtmX7e/AwrgAGViNao0EWSfLZk+xEx2UEdomALf3f+V81IDHVLc5WkBsQ
rniBDFp6k1Hpb1Sl4CAO07psQOp0gCa6zJYdkkcLxEiMybpw0Xy9UsmQWemF
w7F1Yv3mT5m3T7WZ8vDjMkz3Rwb/TO7AGeXBiCsc3gJtcN/UOsAhcE9jk8MX
QyUBtN+SdC6NDpBeZ+AoErfLw0d5CFF6OTUq+HHQgONkHEEnkwRPEi45Wupk
qGAE3f/NrPAb+8jVCGyycmPjkDBu/IftspmD7hIGjhAAOknjXKPyg4Yj0Ag9
Oze6tsPKKcuMkSM6J6c2gwKA2ZrXllSFvkjs7/X3rk5iDPWxWEsOlSjrgtv4
EgWgUvDcldSepfm1f1xfKxXF9GwTxw+xfPjeYjlizj2zxmlyGKLSqRU9+65T
0jBjSTIzoECezCHDqmk1A89qEhNtKfg6i+BTAb4A3dmGuZA6A6L/m6OSGFP5
Zbf6iGqx/lo7zgg679cOj7kWhGMAYKseDEC6bR7E6uP0GTTGtR6NWDZZeGb6
ytxkQ73Tye7cnuYIBaB+/0mP5NohveeaB9OxDIVx7f3j43dblOiF0Z8WumXQ
GPj0wbpgEsfntQMKs1H+Bz81yY4xNlqiNOVa6fiEmZ5MIODgwYrra2fI+XKm
u6LmzPCpZ0MuRcy4Jvk4rYNyl8jRjI6amlbJmPyaNwu452I3GEqBrueZZ4nL
wlpmAlgUo0Rk0bGuR5V0zQ0VetL0YduoUi5X8lip95syyQ5vt4TscgSDKTLG
LMi06EryQOl6aCzNbbUcQXCuaaDSbi3mQU0dQiQH1qnngtOfd5UtAdqXh+pv
Z26HiIi7KY2Qez1zBYZjOx6r06y7896nuykdpHYiYOvF9oN0dvvLkMqotUQx
ia6IWzbWDtXOiotU0LZV9mSTa/CdJ8YWuxvY5zgebLwj3rmZ1uMBDoRtzqpo
v49CkpJ8ePOWgztbtylf0OqvEwuM+dmSlBnAuwzC0jMyKTkYZ3GXfFNlhkde
1g1rntJ8BdWZsqjU2CL/NSQ4UJg0jzBcyW9LFK2BrtiwWMnDlUVxP+EKCJ/K
trfF/WJobc8xHZvzyaYg0pO2FPhaE8klPDmeVnd6RA6bL73xw63jBT8zVVav
Ld2c624DBXdhy9Gc7AOYX8htPxEEOJo7FJRSYy84V4TJDMChVbeRSJSyPgJp
X0tGVJRTVVh6SzCMWERwKZVz9tItQkSS8aCb3NmUqO96LlQVixMNgDvzwNrS
cwd/R5l+JwWDL1Z2ymKY+NyqhJanexsqcPBvtTOQ2bMBio6GJyEuU6lIdesZ
/R8PLmqkmr7oW4i9CZ/tDVJqEpoo0tggVqx7SyalpCLfo8o5A9XsHEkG+DKR
ZgxfhfV3WmhEunI6ZIlWIwpVbEqUzgl9cGk6u1gY5sa370yldOMWo/dMat3W
ASeFn/9evMsDePAkUCgi0QIB/2XTZVF8xFZQYD45+cv71XMe1ZR9TKeYWIEr
kOdghSIt3M6tMPanoCrnFrI+kseNIMgEiCNKgbZvQfs/Ek096bcphKGoOepi
lp23VNwt5zn3upmsMlSZniTQk4kgCEwt1M3VewxsVWVgBsWyr+B88GToB2Rt
X2Tl/i/eutqanRN5mu6/QC/umLRLq1KqS5hwNyQp1aFixbbKhdtr/pL+xRko
pXYdm6+XJFEwSM9OTqWk00m2hD0RQ5b7jfI472LU8wXapgCWXl1DYwwEGUnm
xLoSSHNvBCz1crXHubyHCMhUyNNTpz5NaQtPqvZ0+qVx5staaKsHfItX525p
nGIAFzUt/eYauuKbZNe3FPU5qCn2JY3Ay78KOecY12jQPbXapnbz4NQp/Fp/
ruBWwYJEDG1pjdGqCz5bY2tNGQbvXhM3+Ol5tcLVx06XCi4SpKYFL36yEy22
4Hvr1kiS3DenRVGNGrcBGJPUXnFcXBUh3KWH6puouKwFcLvQSOCrcloHn8WV
IQuvb8ICwQuy47Xxq/zG4lpsqq1ozJ7nHdiREeA26TMmF6zwpLv6iIDKEfsN
pUmV0kulZKgUhdC2KPd2xVPxoZUAQ+3+hd37Cnt5T0RFE01jYDY4kLCQ/Qt9
C9zStPyvniyOSWXqHLOaiUa/59YDABVp/vv8BSq7uA6ikdSM2EmBfmVtIcMu
GjfAsF85WkWQHxhrnI8kYHE16G9W1YzrMCcnQxtzfY8MVICfeRNj3ToP6XiR
ESbwKPpIHZxXg3kGf57Xixbg95K2Gk+OxX6+mr/kserZR2yPjZkvvDzKLeT3
8/FD26GlS3c7+e8NS3yGsucM4CqVOeMb6kygI3aBBFPNm2Uq+xQFvJe5wHLZ
N2L1fIxgaybD0smHpsSvxt7VRR0s2c1M9novzIj0Qr9hUQM5qMJ40FX71KmF
LQmHe8oBNqjvJT/2TZYkVT+qjkqzpItr1saLYPp1cNaxK5FJlMjZD3kifqSa
uB1bQAQJIGyFl9+/l3i4CdsWtoUw26hdJa5W59GpVumXtULaAS9NkK2FYAsG
RMPcpoUYFQi1BDY2tNxt7kdErTIwbQ6FRL5Mvb7px64L6w/VJ94z1fPvjYJ3
fOiiDv0oJSIkeLDKaxxC0R+Tl1gzjW0bDPq84exTgc3zrA76iNIXndip8KU2
SM1cKXbC6GOTVRRaixV94Rh2MMOcszwkquisClwZcI1wrwIYNK773VeQfbIH
MqeVTz9brT556ldgbOerooMlSJ/B91FsV8n5oTgR3UqBrFcsAHbTODLY8G/+
0xtCSOYeFTgjH1IEQUsVCsvG/WVKIm85vjjYAPVVMWz8Uo1QuY9qgruR9hO8
5OvTcR64Nvv5il+bZITejz8fgYtoGvgw/jt5kJUwVcMQ/5Lrvw2c52P5c1Uq
IVEeFQEDCB9x+JrW+5qxGmrGBG4+9WnZKNh8bBR5h+GaUeX4sFbECo2OT5+p
zETKCSbJEMJ/Xq67jpZO/ue8qBpPVOPntp/TY3PpWxDwGc9ukctrskPXYha1
4K+rX9lVTvvau+i0nsHU+Wsa7wIpOB4QBZzws8pyh17mbNdIRphtukUaYsrc
6J3E9H8RfcxkyKF0aR+fTYh/fzon5m00Fq28KM47zgyOCVczKWCeLSHmtF88
q1wxLSHAI1dE04FBVHrUeaXKHpRQ2gw/ALmyCZhIyDD2XipmTh3m8SxRCr2K
eFBf+WTIRdODlTWQwx3Tkwi+h6+WGY5kqJZ4uh0sc1ockx/Fz7gXyJgItael
72srZzWuLcJCJh3gJCn/3I2KPATfr7K2dD0sQVFLcQ/ZYqCc4rz2pxVuiETJ
tlzLSBxzCSjVlsxzponUv8MNFv9N8GCbKZLP66Bea6xbRNOJMCqeIW9DC4jP
Xq9twuCVwTIcYO6SlqhgxRHQ/aQ9UVuMQYxJtowN0NKd4sBnHIHktO/xNBzO
y+yhu7BZX+bKsgS9hV3yiHyBh8DJKCfAU5QVXLnWZAsZX8n2OTob/8fiv1qw
abanNPjbLzN140klCT9G8f/yd2RNUBca2RAOYJRvowb8KZCoPWub7uVJFzOp
27SgZdwf2L7midEdync+qsykX/B0AWu90o0apguC41Ar4UhAzlz6NWdNfT+z
TdhkvKQIPunua163+C7aDb6PEhFJUfgRLzc3fsXZgm5iz5Mxkiqd7qhUB0vk
lA085+uMI5CoE2dUQajtGZ0jw0dOvhq7eJ/bOeQsLg2sm2z/I0tCIs4br9oV
GhUCSjZa9uiL5i/eHqSFOpCsn1KNyd403m3paAX7dHr9J4TY0IWfPVyyNuAb
aUPhzXQTq+B+XUCU8EpkZjMrxj2oUGzUumS1PpYNbrlt7hMgZYBybrTtUSQG
x21yWo+Z8LT6KbrMPaWUHslaBbeAkRRNPDE5oICYeF1zoi1nUjab1pevEWRL
EmQAL0zNbNfb89Aq/YnutpXWe7pY+rSXbs6MVkfv1wNa0e2iSGVxpHpI7JQL
L14s8Vw6TMrzjlX8ZG1GX7ZkoLGXkEdD5/RO0hQbePNrGlAMPSDOFSMsqzwt
vKsXyPklr2a/ojx208l4f0el2YclrevWR4wAKfh71IcKZ1wu2L9DX0TTqBuo
HyCwEUixBQU8HfXoBk4KWUXEKkH4W629QZjK+mKlCrXAlBsl/6JDiEELy/hr
4PnT5JYeLgbauZPe27ZMgQ1lqHj5zty3U+SHVoWJl+KlYpmCo548ibUC2MHH
7owAnV1/tHvNRctVOUrUvqZdGAThbOCPj/tEFWPJSapYlUEflfJyMVPnbA3N
FBa4XcfiXrHYmbOJVq6OCkhrbe6JIMqfCT+PCHb8/KtlHZxVwWowMTMWBl1v
OEVVqWMY+yy3vh+B+2j08/jMBgmzqsF4aEgvrdpZuwNCuEJkSRKOOGj1D0m8
375T1tSFb/MPrEcJA6eSLUbyvQyMVIwhSvwgtKC8STZ1elDveyY2Y7zINYl8
UyZQJBOUs/V2Jt/aSLAYsorgDBHxXQMfXcg0lKlV2olhlEcZxgDNI/bVUIyM
tOf8CfTDjEu+fFnU8I3P9jAHbmHpyUjQbkcn+/yY73tWdiQjHGHeWxsiNlJg
Hpos3lsjqmaFCE1GdzIIP9kxxkGh10dGKFDMRRoPwjgK23zBpU0lc2GAeQc/
+b5QWOL3O7pbGXXjz5QOEIBV+9XrSACtDEJ8xco7nrkFEHo5GEsXynD293yY
vHa50AbcO8l01YEr9WqykIu+WLrzTBDOOvSj5/VfBCbTPpnZf1I5C0jnwhIy
dtd5hXMCDUt5YjRtnmnyrYTnj9+MQn3NUL5k+ZGWvkP+9Uc3+aj84/9WR749
9PLaY29K+MLaVRraRT9KW0xjgGlkffediu46OHy95cb/s1ZUrsWmBzJEHOax
96J0FpT6fIOhQJlgQMrV1V9NB0fz/SIPM9QkagQsfAUnT42Smj1jwZWXGCOl
LIgN/GGpCO1C/GugZgAbn1Omx9rj852HEGG/NvICelFH8zh1DmFc0CI0QI8F
NjPrG5YHtrTGBgUUYY3PgAxiToNzZBuwB92R5e9HDYlM+O1W6glyOv9at8lG
FvCBMgm45VbrGal1GWKbnMzM53OZHMRWLwYH/V8YwRnXgOCMaXSDyQFIBKSu
oZsdHSQKJt5n5KbU1+BQM8jVnhPduYqjzueLHVVFA2RCkve05/VrGglxbQuZ
S5PWljcHZsVNqkNkdSGY6h7oJMbhlk9apRZy7kvCZpnAK6szgP0lSdN7XSli
kMIUd38hdWnxr7+aEHZhyREbM4YtRoqc0dLpjSLHnIFWC8XT5F4ZyUNyztR9
9vHBUYjFDkZxwd9MQEEkKICdcya/LRyYcE4H5FgntuPqKyKXEfmE8RXaDEnE
ax1tsmChaaPuFyIImNxJWOCdIPV7mv4o9eefGoZyEZ6OoVdHbZTiYRNsBTKG
e64jfaW3NcohUiDyGid43cDxn2EgBBoLGsEB+mWIGlFVwFSRdxx4PC6disR/
izMhmcarv5rCTj0XAjAIds7YyKxsa5DpE0TQPavwvI3es9ThTi74hNNzcmNL
NP305tJw6/chezJsBAVmzqAMHo8c/8Sy7FzrxdROGfpmNeymdkeHzWH9oQwv
xAaWC7jtkqoydNsFxaRbSJgXAqxebjCUAjuwwkk8vkgx2Fa0UXyJHknCDEbG
d9Wkt42w21RuR2DTil1Jz1rpUcem99YIGSGoNK04tu60DMg9K26867MYeihb
BnKfRX5/XsYR1xobu0uQRsDJzmlagLWOoc7kmX5k4moq6PSqTwj2D8WgWwuJ
mOdj8mAPX+124F23dZRZA5SY9X56vR8mnfpF8xvvyOJKDLagCeCtfXxIHnge
A7MATC3AecDBVvSwxsVaEdCJGdkjw0/5oHxP8abFeZGHbkxyz11CDmar+kPZ
lRXlry3BXau55Is+4idNzf0ACx6NzIxOvQdFYC+rmQkvHKEEaMjTiUT3dWKY
P0B/pO5UYVi3a0u7AUkZo4AMxF9xMXFZoOdVCSCFdwFsGuEuiA7zVxgIL2sr
EqctPK6ldtIUn/Z2TZtJgZF/LHPnEGmZ5SHTfFCYE30mBgpkhK07QtIkgHZd
crmkGUNvRuiqt0TZwU2W3eVlpnY7CGXwBz0e/YHtiTSUnSj/3T1OyuQyaCtr
R4AFAYLq56Dx7CQOkyGJ1mAdxMifKpaexh9mxqUKIlRECysDMat0iO6j4xzK
/lKPw41ZrOp196qY5aPqi4cvTh8tXo6QmTOobPk3ArydjFaTHclrLvbLRfXz
UAANf88DA2kCP35lRBsqmQVpHJpaJ0niP49Ps46NgxAdzj3yl8yj0Lkfu8DP
zZj2uOIlkQ+FvapTj37Q5TOMBObTnjDpDm+braQsvsFxqlq7dxHV/Z71P5qY
VHwp4ttmNO1DP6Z/VBOqnuda8H6Jwe7uLRqs54x/Nmbj0RP9pr2J2WZ1HgpD
6WyPj3N3sZwuU7/pG35IhZFbTVathGbUuD+3D3ysrf6FENRXVsteTq8hrqgO
CxbPShaO8gAINTF676dNQdkUHpDkPDbw7j66y6/ftDFEt7We1xUnpE1WRk0d
GGfuHTA5cFOLqOiDoWbkmaqAU0jHAEWqgf8dcidZ+lTEhxxaDWHDsUUKxu1r
FyMaj6bjfK3OnZJnBnlFdIVLCWj0ZGWTX6dFfxm87m5l5jYiI8inXQEWbXha
nTzXm9mJLc07yD5L/ce6p5wpEq1evAjkptulKr5oqwLCkNxbhtwnV0w2LabH
nLSrc5FGwqZLpuB9/VAu7HRn4RMsD7P2aKGV8ZkbQwNUZXqRl0BwnktWPLdP
rbTi5cUkmTrlYXZ56R6kQTrrQ9VWZrNNkg3QAV/Bv/7sfgQvftfvWgUHQnjG
J9a0De8d0vvYk/6TQ6vgIhsYPy62kNTz20L6uGNp7sE5gorO3ewCXKgFawJe
L9xMZCWmJ0SlHf0NBIQ8hYUBtv1mZU9FEOZ1wXb29JUCDqauVcl3ZA3PXG1H
Zsv9x4l8HLnh8GLr/rfOsOiM/iBCEKsH7XB3vO+0MhcTMPAQxzRO2eD3I7A4
rJbAVfHRkHAkBfki5aRztDfrpFBhFATMupj/8TZc6YoP2wEHpWhZXkz3bnDr
bKXiQjg7VzoyoucIfbxxXgY2z3feija26eokkU80kyiBhREMFk5u/o84OPi2
SIlk70R7SpsQvuZM1tuvvsABQe49MlNX1udF3n1R4VedasxfmW3NjoL4iG2f
6FRljJ79py9JnHdItw6poGVm+enal3LdYaOvybhcowC+Egat0XFHGq0kEFQI
9SZgtezzmbmILKTDezQI0U8JJGRrGPCdJcsJ8klVSC1/k2hun5HlU4ZC3ebk
R13D5jglm/z5l2o4CsqsoveY457lFd7IdK9AWJJbZiD9/oIYwxDGXhA7iNVk
bsRSVxeR2tcgTol31DGZXvpPwJeTDNNy6PZMDcuRz0qZgglcxNFtJhrsejus
kTkZfUh0AxdPYuAL89Ah6xhKA9x4CxoVC37Zd+qumbn0sEgad+mfhUV4oQB6
UqbwRz5RKqwvwfbdEyM21W/osOhQCtUwT/LOxOBvdOs6nl8BxfBAd/8zAjvB
rQVQ7e+2fTauPHBIPS1ythdTbmD8Ep2GOQZXrxuQlKD6747A7/egQY3VPQm+
Pmtl1SSTfmM/FKzAJptGp9JVxsj6Eg0geCcRXBfTrloQdGav0cSbaZc9R6d0
i60+jbyBGNmY6/70FYd86+qjtqY1d0rdSwKT6e2Ed54g7LlfqnY88Dof7RVt
IWY0XG55LLleLtEt5VQWTgJydO3c55FjBtRDw6DLJ+i4xK41TiZIsj4eGcg2
eIQAshZMp6/zPPaNwDX2VoKEokk9HR26LY3phX84aR3HwiSlNzpbPf2l4Iyy
lDFPlHpYLw054Vz+unbeJ+s57PYqw2sBU0CClOZym5PdAe9AH9lucbl1NsLk
putbLV/0S/otxWQ0/fTjLhRNKd+TiX1CGKuslbBTC5vCWzfZusiqiiaih83W
QxeQ1PraOl8+BFDVqkNtzQCY3WMcreGL86mm3dQrF8r/ae4igl+hYZmz3Pl1
urDIRK1BuB/Cn7Wx+5Tu+gVo70Ue7wRt2jHwjPagG4uVOKvHD7zV1CTJVdVY
UrhELEAntmAIGkOvHtOMr1FDyifGGyO7Y+aKXZ/CTz1pYwRlG5ZkbdWmeRXW
MCRzxuqwguK/7FtnjYWU5PZN8Z5PFIL8YD+/qp62n3SLuGU/RIaWndTNGPKb
LoFBHarWEjRJDYrdcLuB/Xi2XAlxJyesyeNBX3dD1xqtuOQEIi/0+n2Ycy2N
t1fSGm4TK23Nemy4MJVWvkWZS5DQwLxjEcquzBbZmIcKY91XFZQltaKbxGZQ
IlX0mUH04Gkc/6uFIs/Swh2FFe6hPb93Gyqat+D+oONCnDEDlNuAXxkdyA8c
0+7OQCakMvKPJM+PD5GP/lo0BYpa++EVmqPgP6HLqtrJyk9FaXjsjpFO0+tE
7fTkRAl+nsnUuvLewuF8HMfH1WvxKtaSEnEbaSdY+8vBaCUvHyKSDqcGji42
WDoXuewJ3eiJqm3otuloPps0fMJ2O9VpVKDYPJMXFaZw2lZxJ0lTUtlS5b+P
xhu7+IVAr972mnooZ8OWZe17fjtl2D5k9O36EJYGoEZ9NUOOQKphRHNDYFje
84RUPIzz4PA0pn10oon3VDMJ7LvIWGK291/bWu4FAQOFE/fBLf+vRJPjso4J
bfJYyp/tFQO32P5k3aUVQRvIBzD8U7hTwZHbxHrmi0xr7GxhSyQtr3dTy1jW
e5PdxDEC64ox/1YVcl04e0MRwqn56slrIj1ci/Xxd5zTSIT4iRIBG733A453
SfhGZNIeM726TImYJ5bknnWdBb3kqwFMjEQL1LCOQyShe9TiiTyE0T4P00c1
sa1Ske+ggxSZTJYky+IXVj8lYcDXy6jWCEPe3hurJMD/7zFmwStRDABWLXAe
lS10JJSJkv9A0mS39l28qm6YpF3l43GhcGJubm9bj+e4IaWE/fJI0yzbfbj/
7Sa8ECt0QfQ2UV2Dnee7k/FM0IDSZkx9kxmrxSCAOqzzSLzZ0R8w+6GFNoYV
0S8Bz5FdCpuNx7lH4SidFd86AGp7FXrZMSZTSoSRzc+7wQ32K78CQW7ZCzYH
x4F7YF0f0Z6gg/RRXhk0nJmcBUV2alSk5yJy18G8OgLJRq9YOur/XEA49WhF
5ns5fwD0NEASY1pIgnXZo38xjhfJH8rPcqfP/x+6ZpS/vKT6w9HiGrGwRGrB
pkVkZj5+rIUc9NJLyO/IBTtoxkMrwFjQFDvVy3VHJvYvICSI/a5QXk3xeAd9
9XDKw4dCu9JwyvaFC4oATyjhlGvhT9vXKzqvBM1NUkpCXJ83tJ3RLXLCJTUg
6pC3UIuG9u4GbeilwshgIP893+CYpb6xPdL4U+cFhD8RwiHR3925LJEHLWgE
+fgGEJ9N4UuPh9Om/FoDSlMu/nuhgpH++fs1uAq6+bh8IZFC4OgakGo8Xr3y
lUvXpZRCorpOS7uUFDoTcemxswNAfbSjNVz8TxdVXnQAeAtKzrDmrSi2MoeC
Zo7oMw7Xs8xbUJE1dcw/VW6kfh+//MD+M8gvRP65pmKmJER5Oj7do3CNHDXV
6RG1fqlTn5WXI0IjVtAlb2wSEUzuaLVDs0QC/tNaODB3YsjPQzFxhXob6vvt
xfG8lH/wyZ7meSFbBBSQn5q4f81iAyqCCCx0uVQ6RhIworihQ6rJPlPG3mK7
958fMTYS4goSvfbxfCHXkit+JJkb+Fi7KiYCG2BPoeAl3jzoFYbmue67N2fL
LeKTv73oee1Q+dI3Knn+mGKLa9A93TtYOtrErjkigOePIkTPGUR0BJZmj9Ag
kBbBne4oYktJGBJpk99iLlbXuEjEinZjKwC2tfP3hqF93Gb5kBqWwl/nPTEd
lJY7r1j71Xvgka3OqvRibh+erQtKNqidMpu3zb1y3vivlnmk2dQcEmEGUhOI
8ICpitQtui1Y31lytlEXunrXlwEeWt5+Y1DOG/Ga4IXlSwWooISJajolyfDs
XrHJK5q7PyGW34GAh0nhOlooN/ZbpJiVrYNpl7ANJ/DKt+Ze2S8tNIQAjRba
mchSNx4wKaWnpYhdBhhbEiUlQ54vfwQ8yLpTbDQuyyZMu58bHU4qbQPGMqnD
BfmW0JdhTYxP0dvL58KWppgkyzyvyixLByYZs0xmARvsGfZ46JJyLO/MYZ5b
3pmZFgd+2TBMsREZd8qJdR+Gg4Y/h7aAfpuR5ZgU7rGHorFriN2rojvs5GbF
CWlAAkoGwwCEDTDoCMVNY5si5tX/hZAiqjaDBY1guKuROmjBvK2QzkVyEVXW
2+MM33J2P7N8se5Q1la2PVUCUx2CR8W06fkO7wdNHDn6IULegDUyVTs7eoxT
ZquINlPJOoEbTZ2/zzalQX2Svyy9BnVy44uJ1dI7eL3ktOjcRlS6G8+wvtEA
+NC5PDeAWKfr3NZbYX9/JyAQPDXwpW7y/U1cnfxyIIqAV3JsxyrbksS/9h4m
chaJJIuC3zHHrE5YJqe0I2mccauNVSGUe8MENGy1koGi+UVkFZa011hmSENp
otpbW/B50mlcnhgd2tUfTqFKqosx/wUygzP5Yuij7Extnc+Ld2bI7JtSBO69
iceLsWIfDlhF1aHmcBY2l7+QYnuU2YwNuUP2wikXeq2Xjzd4/sze7Grz1X8o
lfRy5SzTzwTqXbGOimFcb+ZWSByRB9gfQrDY8WNrj0bptopRb7c6cgyevQzB
odTYHdP1tFkBAXOAHx5aC5243sJRBYY1AaP+ZExzCWnpmIe/pGNbp1qARd6v
lRgYWcdhGWgdMJrlWY0s2chfYPBX9qSC+3omQ8w0wzRYO1lmh3Cz3SH8AMJa
mejbjN0irhg9jlzYMpzBkDyVKfFK4662WSqGCHIKlwOmpdONx+JHBIDEjEgx
Cjr9TEb8E7HkT6MsKT8zlhGYTGeuk5Z2ldp2fRRwdmOzgK4SUv/afvc9MmvQ
2//dPY3OO/YSe+Te/iZRolAVlf4rQnpXV17oQtKt4+WBFGA9EjXKVTrxN77l
ZOT0BKsJ8oREE+l2RM8NeJZoodh7JE2YvWMvcFzSMRBKzvCq7ARV+SA0G3zf
qQDR4y3Dfie0iwkeXe2Vx8bi0PLBHLsDvwg7ZoOJyA4BiIyJCP0sWQa44BD7
cfv5cvBbhl3zsx260xKjcFbVHeMzCdlmO4f/Sj7EDPHBE4UgloObXAOZQnXG
InNifOiVMx+HN2wBmXzWbi0jIqYn5GxO57mR2T1LfAigP/vknIeGsT95UUAC
g3igojYEvEBppMUVIP39/IR7IcV+KrQWF3sQjxEWmxGao7QWf0ApGT3idLgI
IOc2omFCq90TO9xYaT0BEhEUWbEO5kVcE4HODDEB7kk8t78bsNcW+ppE37wO
LnZxo11vY2Y++GSnSHac0kRyIZ9KIr36OF4PcCPVsS4qRTGu4EarB0bRwNjl
OONKcnu5dZGjQN6peY6ItiYO4HLu8anPdU/tYT3Jdqbk92xGavp8OAT6hqyB
B6S1j8yFg/uC0fSsUbSh4QUbqSLj1yUnVBZ/6hUXlcKN6NgG0yyGjHEegqso
4QGd7bbxC2fA9YOyEHOMeDR1pp68oCADRQT3jDkJs+I/+Ry2oVnSSRnBbZsI
xp5Z8T6inTaP22pEHUUlgQO17O8pK/NqtUfrgIAWzKTlQwNiKDhu3QfB/eAV
x11MNcD8kOm0I1KRzeupxVtkHmuJyZbWVpLCaLDfvi6sGvrgyFTAESoloxT7
CZYIFJAChjKpQ/mF58gAe8y1r0814gpt9cGhn+hk0HeeFUtMF8BpJ9sjlReA
f6VXNHxNJW5fyIYQ1oB9799skitvYVgwFzC1UqQUXCYQYPwSYAtPQMcZBTuX
YYjQl6NeQYUxaz0V6JT9+ItZeY4f3vpkrjLssdi9b7sfOS1MofNEf0RUTG2a
URgWMp3FH82BBw7ypip526BfWfDPXdiIaA5/LGb6fKp8BA3GJcKt+yePSpAJ
XLrleU+3WOdQKvb6fAvrHulHB9ljcAqlKahcAKMPEbePQ+BXfW5jRakPiFCn
8GrFD7rAhHXbNw78+JLyylosSYBfITe0cEL8OEnaXz8OI/mtqxtcSXiz36a3
GIBeD7mYppZMtSbCEcwYuxAKGB6H0h4gl5ZFCOH7iwF2jhlqUYElQbU2hhoe
Hi9bJWHWaGpfAepgHleSyuC8hVGT1EKXXswWmaBrWxaWjwnZ7B4I+cNCK9bB
VL7MvcCK/+Q2VhonY/bdyUcXCn5dUxcWMA+CLeZmve4bLPI/RNxrn9ndaPBl
hXlX1x9D4/o/KdhXxX8qIt/bnrjIwCyPLQdfV/MiiA/xGuwtbbyiHO6xzokW
IJydcJf6HAabu4bovuHVi3I/nRTXDBz1g/01oRyeh0/wRvYAPcClfIfbhevp
ratTwg66iGn3eOP1zwkGGV0I5z3upVfIQaY4xNzifrTx0in20wIFmsU6h9Ib
EgyiooTLDyMwvizj1AiAFNpTICzJjCmkdblNlWyDYFjL6pSQaLBKaZrW56yK
iOj4b1GUAZuk3p4vhl8Xfk24p8fp2BekCiqT/LDGbtDmnBoOp6JLon+/SVEU
zGELREnxqlnCTEkRg9ditDxSEpHJBS3Zf85otd9mSBhDfzqXXIlY68etU/77
CC1EwklTCM9bihG6atIWdqBMpWQa9I/UzqCAB3d93kXdsSEmDfgcquAIKxUM
0+Y9fewBFsZiOzQGaOeHwCX6YlorojtwNTTI/MFNORun3NACDe8Ia/phemGC
L/5EfcwLEI3fL4vHED8NhmZHUaLmbMvkb7MMXrUctZza8ey5H3483HvUAh2o
4DbFoXKu4ng305A82+y0uGD1FtjpImv7D6dFMPc9ikqJdtxUF0YgNUkYBE1N
GcZ1H/8tvdqxjcFQQSLuJKUud5uSqFwbgAsz3EIEHBYPjjxW9byGl93eUKgf
EsekNdlG6YujgaUcWujpxONjiZFlCOTU5W6IX8xDFFj3sn58zwF9ul2bBIH3
4EsUxXfiJ6b5s4Y55vU9V74K1XrT3rGvN5UxXGPyXTL30XfTwi55hQQci6Co
bJS43l4udC5960L1mPuSMhJg+4VqWFxKRc8kWboizxaRIIeg3Vwxk74hFl7m
UkFODsZlxfiT9RGD+sevsqcX3V5KenPE0ESohuccq/jHYkgH/eVJD6JCIn3U
zjqY0HZGDXynIakOOO+88aAVSs8chsrDGRpJ+Kr+RLMep1I2NFNucDVX8jLw
/cHrWQlOav4JfM50bKmRVrzBQueK3V7FSoghW3q1jVERsD5PeufHsbY9eJAv
1FKt5C2dZNoyEprfVLXvhZ40dG7JyZRe3kVbT8uM1Mn0GWfVc9+1cNehaXSy
Ev4Lf35YM5xUidq2hSorJ3SwHWIyRRGGdV605j1moJHNItZAixbzSpvYsNrI
9vqgMDHXB3xzxbxgx49JKn+2lH1to9qCO0EP2V1T+zSgUfFINVMm5c18XGac
/XJgug7WXJY1ON1Ir/zTUd3QRtPB1RQlLDSFYBxQcOnQM2+HqHH8qkWtItIL
GJWxeQiGBBCeGYKzufyKVQHnhkhPXozlGBArbLzgFXyxzca8vRkRX1jwnQg3
fq2PzwOXVDVlHLD24KEiJbxGZqwRdpYCTlGenfd1g/QKREvYT5w1gQCgdsbU
+oVLf7y5Ij3KIbcq6D553TLRmF45KKMKbvSqcmi11YEQIZyNuU1svehaEIqU
sk7PGRRhzDLNEDOtKb6g/AbwZx+C6Ez1gRl+SAEBuXk0uH9RbLWHIgI5bvkM
DGaHm4d8QmH3XaMzTODTJg8yPSgA6SJZ8QmAnPgSSXR/W9LGwyZ76EtzNURE
fgsRD4ZhQDRmP41Tb2++NwhDFvqtb4S22ITNTLckhyzkbnEXkM+9XHVYEIqd
5uV5adea2ClaNYXW5UNvX+yaUCKeqieM4jGHOWKX8jFd6Iv3p+1wWfE6roqR
aLL3pS88oQjys3XJCdDQfTfQH1r/Eu8g0tKQ1MY0/nk20tTlEObsfQqKvaiE
RtQJqRrYmGqBadXAINXXQd1wd8WPp/bx2TpI5zWTr25xG5IctxzBLQjxKcak
dLkeFIU2ygbBFDDdH3IKgNUg87ONqobuYI0WbDj06zhwfEzAV237mA9fbZFA
Pkmcq9vH+t8oavopF2HVAJwHL1/PRBkbGIxYgdgvBrS2EVAOhecQyrP3iCYW
JmvKsLxgcpo2XUiJR3Oh8kop35TU6py8h12EBtGNTDB08NkwKu2tr4mFI0yc
BJ3tZMy3IFWyg50RmQMiIGHIHuHO/RzKCpsuyM2OPWN3PKWLQJ+heVaXGOah
ky4dTL6q4E8c/qw/ttV+pUgOVcNPJKuIMqKY9Kv+PZ0dNqMOVljaOmIBjP+6
Uk8hD+IYiOk+DTWFGe7xG+b3VdXZGI1AV+bmNy+tJiN6pgXqctbfc+9tyFny
3ITwpRgd3R8V23JMQiyseqtqrbXKmGD/LOeoCdxt8uerYF+glil9TFkGaXIL
snZ4Rctd5gpkJPgx4ZfQpHULGkDnfHwU58t5tPyyjGcIMch7VBprE3osw6G2
uyRvgeXldCfUZMAdnAf6lxITWwPuPg9rCnHpP62zksyr46eshR3Tn1luMNFr
6gRjtQ1796nx/raxJCMzu/zD9kkCjEuO2nkVvnM4Ux6pAA5Rm4pOUpT9b7x4
Nhtcpzm3cOkCxhgb6AcqiEtGgEQyG/glRftKotfwkGt0ZjGJjl/RNNxCYX0W
FQ8AbLgx+kZbAg1nN/axQ47QGWH/brQjHrZSibbMJ9oo4UhbIf9gMXHhLV7o
ZFyrQhVeeG7eiBJ0DzmXFtfq+vyQbCXP7XLghWTf4SZcSFZXO4t3IZshJ/nw
as1LELnCo1Tt072bsYC8Q+br2j8oKOPqnokFRRvud0r/ay/PsnyxFrhqVhfn
UKhlhxGjgqNg3Phkr0/WRN0oFViqrPhHQMoEahRlWBd/2deBYBQYZrhNUlL9
3xRTuse1HOAKyZ8OQH4FenXNN6gXzND1/53JVw277WxURpUWZOT8gFafPkxG
7TbjEo5jiT3QfFO5wN/dXWfIT3ZnED2aAdC1kQOkEkCikym0fsqcgxIUIXxA
CuCRKZ5c365J6emdJPqBuryEnG0FqAx3f5FN51BossDAa2m8Tv71A1SzGMIJ
yIB9VU+qIGswMXa1CvGgyLIczYJv/80eC0eJyNAwUR1qighJTkGLiVczqrdU
oLrk2VPyQkUEEpmDRF1VcP2PHWNnA9fNbnpyMj5JH7ELSKac0tJNewTEfss6
kCtvCgeP8npZZnVCDIShQNLtYGjWMmHWX4o4rt4xW6Yaccxvc3+WW7Ib1Zda
gMNoBBZz8tV2NWse2CCsY75Ewm+RAlNR6O0sWLeqLTy1lJR35D0H1ei6D4V8
sqjCX1sMa6+2tEhi/hZmMCiHF4AMZ+Ao/JruBwPyaGcFEiKj1G+rChkc8py1
tVjblEzpxcaU+pFNdGxQuHwuDRW7DZaxlw/uxxnD9wsyXMgtScLMzJLqrzUT
BPJ7Nh8/raQjfDaAyxtEOPhHlEXf11xCMVcbeMtmBAnoOoQo+ku5nWyHLD1r
tIYF97blYp8E7HLLNyY0Qd22y7YlpIrRHdsdRDCyZ8X+4Et7emcEhaaJ6lbY
Cgq238C2sgbH0eQgQus7SFy/xUJmAnQMXtvqxjntxZlFhdHKZ+j8mDcG/RvX
WiXS+akb1NRJ7Gpuiw/SS/AdCAHg8KoWhYVaROXEb9QO17/SBuFHwvfGoKFz
FNvd1iga5bIT7vbflLIMAd/RFVxGnk1Gdpc/PtpChErS7zYAlKBsf+JY8Ell
Dxu697xen3xa35R/8vUJ9fadIx0UdIZo8juYACZtiIsH3Qd5qXg7m4+UT7jR
WP75+sddD9J2jKJe1fK5ZB1Q+lCXVk0mmSE5s1qw1clzM0AWbke8rFPd3A48
aqRZ82KpSE2QgVzFHhIHRFxlkZ8f3etKr3g0fUXVDH1Pnrp07Mtad2IYAxBW
+9IVnfjPl66NwkcGqwIBkbVbkzFAcWL5D369/FVODFqTMW7uZTjQI4A5idqD
/DxawGHQnEpHp0v/Ad5djmuN7IwYzDxaA54kKX+++2V1AiVo7pjQDndGIBwy
DFwzUJKFxsN4HJiT2/aayLkpWrsyrni2+jVp0qoWykl60cSvLdirKhrFRPBS
eBZAkrACbk3dqAYtKFe/oc1xyydFrBCb0VN4zlY6a+rRY4lINTPo8cillCx6
JkRRJxZysKibHZYGLtKRHuIOo+8he9umuA454Ut8nsyoTwYIl5G+EVZ7j5sT
Gs+W9eufM5YmefWLfu8qo5kGSSePh+ozKbglkbZpYYGpCj+mY3j+zllJHzpa
VXXUT57JO1HAJyxoGRuhAV4+T8jYHS/Z243E7hbv5yu0jIY0wJgxwLodoyEy
AHKtzNOMGhIg6OpIewjfuqQJcrkwJ8dkalzdgA64pmXQaLFEo/UplNKARG2Y
UVSIg9oMCXMvUGQoOHdGMN3mcX62y+CpqAXVPDathj+jQ+E60CjuHDiLA8pZ
NXu4963vu73Sw5+DmGrohFWvGrbT0lB8OMWtlTrJ2AER9flbDXl0MDXN3Zke
aF7C6YKtDtChOl7d9qYabJBsLN6iU9qwDJy9kPWtrQ9ukOatdd6k61DkJBWZ
hHqucB12b44DqxUPu4qlKKho7NcFNHg2winzNQhP5pdax0tH2SYa93EGHZ2u
D4kmYUH9SAc6fU63Y1nkTw+JVVAqmcsOv91JcDG7JIzzjB+UH7yiYO9QrsPy
Cl5GCHSC+2JaFUFdpdFhgNtW6PUL2+vFxJrayVidwkhIhujV5mvqu52fq2LV
UQ/TxJPmFLqLMM47e8Hhuh7Qzw9vV27TST6XlPeW0Tc/EvU9PYbF+tMkCdga
vvnfzxEY4HBU98D6SHO2nbZ0pfdGKgalVerlDr+apR5BcoAFQketqzAapRyL
3vcQtGYvTdAXs8VQbJJcpiItBrQIarffsxtUWlx1FBLFwwZ0zzgCjPUxJnGH
n9sHQZG8AW0KsGtTwv6cIlxTK+raLerhIhoIoIXl+fJsLiGyhhSAB6PuLnBQ
fcW2vNUwdZirzo/kaj8K835eyMMvqoH0h8h/qpYXJW80kty9Q1OJn1IFqWGk
T3IHIS0zShlRYG0Hdmakgo7/rP300eJJbj1gu3VMrtMkP2PNggljz3keDlwR
wy9D09FniXh0kXkKV85hvVkYVN30ZmqRUOm3P76T9qwg5zlbjxSMNVzbLQea
DPnwSp/TS+Agt/1Gg2VGRDEMrQqJPE27SZZuMsSVfipdoyh7XsS5lmppOzVi
DoKFFH+dGDxIut8Qx2RvO/65k6wvP8SD1VkA9U+x1sLXC7Zfu6JFh+DRyLJ/
DOeolbimx1INU8gnlH3H20DZf0YNa2VELNrYX+BdfWRjlj6CXGJY5vv9em1A
VuB7mFXj25a5F1mca5nroNyXbYuqtLM0SMjfm3MTF2HA3cLZaWm28ZrUjvbc
ZEfN5KpGzlg9CA1m5x2DOZm4MIUN3XGHpomUHC+deeI4qr5ibUijsWq67Xq3
Gj/lARSC9AaukAQS+HisKlYPOfp4frgFWlZ4dUfV4yZ9Ee1kkgU/+PrwBykA
d72i6c7pllnThUFKTpqRZnA752D4WSdseY7GThTft65k9jkUKLuOlHjzRg7s
yolaCtMkTIXYrSmzzJ5GUlZ+a/NuLmvDHwjT8VcelScKk9LcrnJqlMw6rTAt
wteokn+o33wk225gNYZRPvX+eH7FpGBQImsbO+4arS0HLaIrg9UO1/BxjKo/
iO3vU9ZXH4CYMHBU2ifV50Yzf/OKWI6yNezi6C/McdcwmzP5kF2EuHbCV4p5
wuXPBUfZbzK7xOH4GPs5jBu0/43aNQ5kFcPF7bjEGcLbSD9+1dJaa/PMjwPA
+DGphkGp5vNDNwIqagZx1JeKL3LE7KcrLagYk9hSdYx7q8hgpxSxR/jzribI
upuPDOYSLnqnmyeKzBtzHuVtT7jA1Lr9YxnWu5sON6MvSiwI9oTIbjfi3XKI
ww2rWssWaQFSmMLkmhlhFPjmS3jc1aO+Hu+uCOESv990n5EtbIV3XexT81/p
3m//Ps/OnLUVGBPdC0mqcnpRSZbWpIfyHu9ta7YnPayW6R8pdwmOj0DZPRtR
s7EjGu5IJ61ALe6LwAI82U0lZ2VDWJkZq8iLfS3mY15Re97FyCNOBAChxdV5
/xYj4yy9k4jAlluGx4KYEFavi04hA8d7d/9wrk7N2ub4I5KKctuBYXYhObNr
5vIkHGLe5yuq01JBZS49g8UTIOHDeVnTYeL75FM3jl9x7GdmlSBH7h7O2M2k
4BpEI8E7onSgp4PbfAxEk4gKPQaA59cqeSrSqIwHPNCDrlJ3vaSe1WdIK0ge
LvHmdsoQtMaOKEXlf/lXRiTzXbo3+geOt8BInRxGV6c4oDILZs4Ka7XWEHRY
DLhRlMxCy4IKRdHrDPo7M4kgedVsxIh68bPIZ58RrBVr2+6vek3ICHac4Dre
xmVu6x4H7ictAks+jKeXTunl+TVUXJvDN47blq/FmmCclv7ZU2laFFVp9MVa
WEGDujCGLUUFOh/lFSOgEuU0KmgCqbs0s7oBp1vXKyrWlKMrsfp88D2dixmo
YUpnN70/4vLbH9fe5DF6i9jhndDLn9FrcYCtycSCGytVWuSCG5C0zZ0vF+I6
mFBpuiPHe8r1lXh2dBOcVRevQODjCnyK35IoN0lzmne7tt85uXyxforzdnD4
43P6reSxmer6ygVzlC31qnLNoiC21meQod3CSywC4FN8lfhRbChBmbA37Ilr
Dl/IMtP+Ur8kBrn/X4XtrF1WsBSOl7Pk6CwtnZMJdnNCSpY+cxD+hhHYk259
xmM6rZaqTbpxBZjQ7RSUUR0nUA+hOWxVMFPPm3VFKuGxbrO+NSqwNX0U3a8A
kKRvUkIgY744BIn9tNtnLSULpSMqkTA49JCprGbP22iIiR3yJgqN3S4O745m
AKEcaTe/f/TyfueCU6GiQ1fAhCDN99SV1TvTnbd9ahjjoV4mUELk0hKOZza8
QkYciqczsfMDL7+eqlWntbSv6z/07lZo6hg+JyljIfiRlFa5BO1RZOcq5hI9
qOuGeSrhArcl6WQgM+mZSeDYg7rf7W9GHlwW5sc0kPi+mHyqHetFL3uj/TBc
Kb0IH/oBB0kTrIHJ35z8Y5fHIVmtphONdmbLoL5chOGtCBW5zAqpqz5TsVzB
s1YXcDdtatdj7x9I2uFDKu/cRipy0fEBmDLjM8EY2472RHB7a1p01qxx1r1Q
m6kfWiyDg+9WHfgZvewAt7eE2vo8yMbFrfuHpwcUGF1xAyEdqdQFTsJaM/JP
vR2kyASFbdmHNFL9vPDqzRBqoLWJAk2Fw4gu6qTg+6zFkEWDoiWW8cZn4ONS
QB8ZTeOVR46wivexIltAEN/1c1+mCwH63C3Il1yWB45JeuY+/68znhoD+YH4
UeDPrk37D2HG6kAiCG/8mUUlmrRElUF/XCryIUhgqK8QsRPzMpEOh/bhZxIx
PaOhhj9Xl3yegpBH6G32SJBjtbLcSJlLgg2D/NbbSrkvBcydwfMVYakgQs5U
ROvujY5ims8LsrkMArSeGF0ODJtURLgitwdmTY01a3K+3JppXaqvW/NFED+V
RP9uzU3eFiaWbcjZ0ha4lGmoR4t3qc964T5WAhCcibh9I059MCvps90Z4rNu
4FZnhrrp5pBZXJvnFkbYL/6ed+I4d61r4UW5CaOQeg+czbo09llgxCNSg9Uq
VRxdWwHrPj7vbwpH+x6TP4P8u30Sag6QznG+j0EgQAlzCTNvNlUV3eQjXUsh
XPlma3mtFJtVOV74UFHHwsvUykN/7OywFsKcxiFutsiNuHfKtt8gghDcH0i+
+H/9KPxkGmHCGUL3lo0UUwjdJV5gMWlGUagTq5Lvdak449HbWWdVX0srSzo8
wHot3Y4PmATRKobNYRt+zTToBq8R29GrHU7G67fuHOYhZP7ff3w2uy8W4Ml+
gogx2tqnwpQAIDgDEjSPgyKURnIM0rDB++dAwxAaNUFdMHOkx72wngOKca2Y
UGz93tTqNjUYHbj1DVzWa5LLehyMJggJ76j9AvgXF8sq/oDEMiwWaH5isGXf
rvWubK0xXZRm1y0GG4utHPwSgTKACr/u3a1pMp/3JHgzdLRkAodO1ja1qswU
vRGmHJCc3DZrxuo+1LOpIrINhy/eL2qILeH09/Y+q3QnKOLyxYsjbsIwfmo3
gOgVss60MlGPOt6CTjs5NlviblKGSPqZ3TbqjMNgwuBNkDnAAMtlq2lGO05s
HkQ3xRNqLi/8IWqA0Af1/To0nLHWngjZwQVLFbz4F5VS7wxO4qlWliCbmfV/
Ao03BuuQm6J31VdYyNgy2L7gsXNeRqAF6kzpPpB9ms34y74U49rnAShtVoY7
lzA5Cr1jvNOLvLEEmUKSdrl6OL14Z3pCI1q2huGygJcIm0X9WDW3ymt7X+zB
EvVvui9I8tLiqzY+8XBEZICUY+wS5hXhkkxwx9uX0oZT2iGrbVAJXQw4bbaS
l4ShHoime5tOq5H+h3kcnsiX85IdLl0TCknJf6RstAHupTT8nNBmneG6jd5p
iermJD8tM6WIMhW8e7FERpO5SMaBMpqBmYUUocruGWezO0LOWS/XvSUv65ta
dD4C8QYUBvk17H8PP8DTs6UF7Ha8BBnzf2KS4GX1PYwAb+7ALAodZY1PukCL
4y6tdO3PzxsYyeyLFDk+AAlbrLiVJjHvbi8YA4pPaV/0WXjm3cyKbcsRGCym
LhWxho5znZ39In7B+YycRw9MPozvPxgIx59Cxh2CylnloPK9jlby12XQhBG3
/T6fRneRWu72ESctZETVcWO8kJObDsCxEGrnTUulKayCoF7uEmplGdqEtLIX
/O0IIUBMJfNeOlLpiBFRhyBWSStz40P8vouBkA2dY9H7Jj6u2TauJhtSIvbx
Y22bPrc6EClRwmlYL9vywoLifcDxrRw1zIMLdZMQwzBdCbwb3U9QsoCRlc1O
fx/b0vmUVes74qo2xRb0zrjM/NgZ1A+7iyUldjQziCaUvACepvGivbxSApEj
R1sOc6ZQUnDCYHaa6wRCm0RBAgWHNwZEevWNqQOOYjGOlJg27aUJcGmlC1LB
Ozh4RS95MNzWlJYEGOVQ/LzjCPaBTJIamWONCszSjm+rlCplrRcZb9iHgsmk
2UX4q0yA1CXlTxrB/z3XYj1TOJ3hlOl2qXUHFzSvy47+XuJ8Cybh3taAPTvs
8Eo4nYq6IAxXJK1j3dOdxWAB/8YgdHcAOiCWxUJWGm8bHUdXLc0SZUPcuNK5
pmqo8XUNBuYo2z02oeG0qxwqptoa9AY/71vDM8vetSJR66v8NCUivpkCBV+I
hnc+8lXxZ6g5hAE4P5vqXRIh5ohxsYPKUxaIIa3V/SXqdB+6z2nYxtH+1k09
HKYxmsVdtxytg7wavgwnRfOxWPphrmIrpl1vcCi60sD5XxZy06BY/qVTeFuw
1nagQNI4/bSTmIp2X9G0HzWB/Z2awyRQi/2vPFIxl/4vaJiXtaKaeELe6m/M
FJ7sjy6EXRmlRwboJdR2r9IGLkcKYwwF/EH0DqFUw6CqilyXlNxGHFFUQuh/
FvFCKrDoNEd3mK8W/wIq6qQJagwTGeGrBJMDJx7ykXWR7zGg50rpgAhhTpEP
HNi2nIcC3h5R7MOh8ZN7+XI+h1wWTSqN12r28UpH+tMsB4yl1rJcd1M63mbM
ijfKqjHxxtCoMXT9pgSY/xytDuhXp/4QVjApO3HEMZ+Jjfl9go8xBWSvRMJn
FkEjXlF2ObafpF5mhV2yH+iu+tEalKoxTH78dsVh/O6dPflH6OhyXtWdYuYR
m/JrG/9VwPWH7w5HHEH5UB1HX7G0ktH/TkHsON47AojRUnm9GOEDLSB1sWAV
2APmanltctowSR5fQYZYcILx8DFvV7GBO/4DAnPsokEzpKqnsdJnUURTg55V
IGhXfNbKcUECHggUdZnxrDzRKFyz8B/EkkXTq0tyvYFto4Ov2LxzPfL5B9pe
d4FJl7zoX16W39x/6fxMbDRpO6J5p8CN4jODpxvrMWMV65W7oK/RlDNDWuQm
kZ4CQ8np4flwQ+Wzhea4h2rUNDhz5LAUSJ6CC+e/yXRslNc9K4J0qO0bP1kb
vNY7CTEewtOmp+So0f/trbTGQqUjtFwRzPp/j508vXgvVdENE3+q+QY4GaRh
YoGyjwELAJTiL63GX7a4fsAdJscIj0Sgz3QmaEQeqvsjR/RCYqq8vacYVtK+
xqVs80VasZsuvdT7iWODfw3PYRp9PQGEUw1KI5yt1wfGMKtBPrMCkcTnNI5P
ssARigmWzuStEIRA0JTZJf18WX87b862M1myOVHF2trD5pgWL0Jsp+/KREPa
2ouj26bkrpP8O0YVccTOYQh/ETgyGQfdlsKHJFxBFJaQ6sg6MFVqvSLjrYfJ
4gEDrmwPQ9tdzWDeWEDOCrBSGOVH4+P89hiKrm21EnGwU+fu5czv/XBnztNL
0KK0k/+TFRBrt+cuIOeRzkNJ3h1eU8r2CEf4ajqjHcnSCwgvisyeQhuO+aDO
pen0VKrke4w5BOljGjQsdAundf2urXw0tq/0UGYToo9hzq1rG7C+o1aEPviK
RPAPjDTUtFYB7cK4ktiI5GXL+TY4kvvAk+cFRbXr6IWtXqFXro4FMDXsAGRg
pD/Rg7tmNlN8QYApfAYYo4RZN3uvU1L17IHIZ/DwVHPPJi5CdJpG0Xuh9M81
CFcVkwyZqnsZpOn2OdLY8zkOZpO1W8pbMdV2kdcwinz/0NpbMrTLKGcyiKz5
WBKDLpLYUGe+Vj8TYl9gZkdixLTRRgxHeHPLPCmyu+uXzJ9PsAkgZlJXbtET
b8ukDchBhd6MaBtQDCzO7nkfMb5bXW0fZ9y56NfBVrvh53AKNRIACNjLltap
vFJ4LA+MrFkfcFAlb+4dDErpsg+dP6WOn1JbVsnjQGBSv0T9LatF6vxsQwMh
U76br022huW9thz8otjl6iF9I4+M1SJ7H1s65MIOAbknS2dYwYQdzj0xtmf/
UNsyH9VsmLOD4T8yjiyhT/MW4yqVGTvxgzw0RalT0O6miRZtBKphoVyKBkUG
uSXmxJJ3O5IlGkfHc8B4uZRcCWgt9xtOSFg5JScIRZLWWEfubDooj6CtfcB+
fXZVLsYsDs4FsT0w2UXj4cvuJDXdZ08PJNprHRAWmNgSfGJIFhQNNMI0XFCU
YGUT46nKsm8cEX+PFy/KWBvxMUY8+h/05oQbn2TxZbURI0Pb3YeRjU50RwMy
b59qREUZ8lXefEMCVbQ1gQ61DzxVnZvMMr1Cna0WmPtJrRuNCUmwiT4vN9Kl
v9Tf6A6m5jW7afAxObqE2aiH7X94yP3bLcKV1LT5wM41OSfSq1hMF9lBNfnC
H0B0V08qn2QTaR9ERLDho1/va2dG/dGsGTCK4aRx1di53jZQ4yUHe43kaUZU
eAxu0VJ9LtWKh4bzeTqNjNjIU4/Y8OlXZgJa9xSzTACPf7CxKr62u84ADOwh
iUR06QZeU4k2ImE8R0CvSZlEZL7Pm4Sx8LAiIzYjmSbJQXh/qeGJIOAa1Zjb
iLfQs4eQg46Y/R8Zz5NuTqGz4aZ3pHmdBt3+sdF3TaLWJDjzgryYVoRsWqJk
HWTKfuGiKS5w/5C37v4aVIgpdHyish1uw2Npv0LtN3E9mf5R/m/b9CCWd1DR
yR+uBbbjatqZS59BmnIKGn+w8J1Y6znfVEbB/p9qi8fPh4tBfeBeq0FA/9JK
D1CL9Fg42nqKtqvh7/A+BpLhbBg7GyGdNuqVLn6tVTS/+HidN1OFfp2vmPoz
Kh5d/oDdwXBgHx6rai5f78C/IJotn2QRLzHwRSd4f2h/Q9vrGB4PZce34Rem
ZqO4SwdfxsP9atPgwZWWM4VFB7QB6CX59dty8sOfuqv/KO0FtRT+oioyw9+o
sqjBQySGn3BTgfwgiphHNkz9R7zepixRZlN8qoIxdUKVZ9LyCV3RM+/amfEu
6FftaUuNvP/P/ficlYPgUlpCljLo/w+II8OG9vI15IYNL06DvgGGL0snZg5H
MNTTmcjHG0gaBppusSR1F3fHzEdK31MyRC+5SgP+aC7j30n5kPMyeG+MQzeh
Iot0ULERMj0ZbA2NC/n3vwJAznLc5vzG32sLwRxJErAZwslks/a1lMQq3bPd
JRRqnVJgORJ/WyU7VagSFALNP5/iqyK0eZY/HiQgl9dRwTOrfZXU4L2YKjZV
UQEH67pUpKzMlsLKwLjsaZY4d+MjBMFQqBZRnxKVS0bD60WsOU9ca5xTcfRj
ocBoe6clCgpJKNLvWBamnKulKDz1NWKG/H3QLEFaISRgI6wlEusW71JN+JR/
5Ow6rvZssX9m0fAWA0Cbbz33Mm5PyohJj9bLSSiPQ9e14YfPgYZLELyaUqH8
dGLSnXEZ9iRjILhCiC0VhXpD/PaVDGlYQ1Xis3vlvg7jFVQ/pcKukbtvUq+B
1auWkeZjmLxUaQAFZSpn0EpCpEOmV5KxyJNKoXttFGGtPoj/IAeWhY2uAFcG
PXzUMW4zIXIgjv+c9wkyKdIPsoCoVBgMh2LjlvPN/icQZSPQUQt9z3auvkRn
QbjEyts+8Jkwo2kiwqhJqJghrZjvq93Rmg86/B5UE7sFO4Xr1i3nhsBnbFsk
dvmb6oYW/PMIadKZKgerri7LG6NDzmpz2ZTKG6L0wo6bePs+BlJNEy1s3jq4
6Qt60RS7lmpj61QIyqZ4I2n1IGq/Tfhg/icjMy8OO5jOevdgHhhvp+SgxMLi
tLFb67Gk/mBW6cM+ByaJAl/4WzMwDWqd7YrVAkrVsJaoYKWXFg9ixXGDXICa
L1stKhmWfZwKLiqpjKBb+2OdQK1m/kHIEJ4NbDDT9i5no6Hs/cPaoqYjOytp
jMuLVLX31PIHG2mAdMOQlKSKA4TeCJ0tOfJKxfuRIsl9km8KUxPImG9wvYUB
PdMxvJR7/LviQ/0m3QWf99tR3X//iW3DQaLQo0V9N3Ij+m5If0DkZ6kMljuH
9+cfC/3SVAJugk0s2ARLvNagvJUsjM7lrd+F5Vj1OnpWAhGr/avmGfGuQJmM
G7l1P2N9yb2R5ZSeXxCtgOGzClwQEMgquFb4fFPg1DP9kTcc+ps7Nm2JnJxr
scLGZM1wn0G8cnwtBg39cL5Ch0pZPa4z7OT/eFLCULRUsthM9cf/6Ta9i5HM
feglp8xEfzVOO+K0iEhbuVZHT7axH4dP8AieDeb91GC+UdWwpMCCsjx2Vv8e
ak3fBS2W5cwHMoEG3SzFjS/VQEfvhuozNyjpmqgb5PfwaSI56dOGi++iZrvr
9Z3083nInBPjVIyVtQxf4ipHtPPJH25ZRXtvGmKBMLI1KvPL9LdTH1Sp6nhi
lXk1iibGoTdpahgzhruiz75WcGVl8WzLu2OdsetdCtVnZ71EsrCqcl8b3krQ
RF/xuFo08zmc64I+lv+olvTNV1K689C62UQddHRy8xVwlaYgFRA6rAqaX232
LMmuKJepQW20jj+MSWvTphFh+kzWX6nr5GM/aX9rX9tpxi025/VnQ5p4QxLH
4TdxMmV+PEbWwXW5a2CEM5wuiynGqhNvJZNkLgkHsoe1pzyXmjr4rTolwNuK
H1B0kbv7NXHRacC2X6/DSVWs6XQT+UPS2k4lR62N3i18IKzWSMXgf70TV8Fz
XWf8GqWbQ6S1tCOOFQJDeN1yJyv7ca+BwMAa95b5/n7YkI+U0MsejuFfe206
UC5JLJ8/p8327pl2+hd0E3BQaaqYnneuSxYexUe5BcWoUiq/xt7JfHFJi0V2
48j+pGI8P4vZu2dx0B2IAOA25UhmMnsnsh17sVF4NYzd1tHZpovvSNRIC155
EfDOyTzt9C8OpSzASvhXcjssPTS2nGxZAIvJsY4IsuX1YUbKO13wuxi3UrzP
xmH+gdRMb4I6ELoKPzKY89OHg5V/DslIzCmyllw/0vcMol3/KaMx8FF0vn8z
qltE3JXpngm+4Xty3asEHA5BMaWFXFAYqMjBORYa5Iya3UgUtYDsnz0Xnoqp
iuwlrHwv+/fBQVTqQyig/v2d7ZOAjkGM80ZTai46l7AptHnMEdMWfPQ+zmbu
j2N+I7F1IulAL6LL11Nv0mhlwt1ZkRmxnG/GC7n42a+0pbtjqeOHISeiPoz6
WFb9UrqtUk9OjxzmQlGHET7Cf7ulhFu1Ou8O/QSxhsSSvc87D3VgXrwk31Yr
LhxHw38W0Yywh3tZZWQ5idGBpt9QrLHKmhJ9WcI4OlrvmOEKQdADjgQiS+z5
cG1IBKTFBCC1hWaVJ5B9D560/Udn2xMfOqGFHrm9OQxH0uihPn5VbKQaxzmu
EM/bUSuH59FOrz/jvWCaOplB1IXnzNxu9LcBUoKp4ETETU47YwuhiOFI7liK
4UJw9JA+DYtX4av0ayUTbka5qFUQEtzL5sPGX0itbbmU4MWPEKY0TWfuj/jT
T4g75xR5oAel94nzY66rzez+jC0IZPs6LHwHvqBDX1Hk4exm4slxRyURTWqi
XWzhoEHFirQ25strHs1wXjAXqVOBE/CA7QvI44j5CAhlPXJlyLbO7S7GzTMC
UIAHLIMJaNwbDVLpIgrvTgaVaDMLCV/gfEPCqND93h7kxvfCQZXxD84TbSbH
u24LJzDMBYv/D4gUheEu+VLH0FEByrIOv6uw5VY+tT4/FfH6m6IAZSUDYScK
wirSAKyIMQXV6qwO7z/AgAPAiZEmB/2yChz6AWRez5qASEzTqWFLqL6hDAuh
msgHygfVrOAYXrSvXAQgp6YYeS1X6VfOL3uaYZvIipTRIQLUPbs2PKfKSvcf
eSQdXHznk1zoRCmj2Ai5JJYhzh4cYcfMcp2r2YQIDbwb5PVdWlq0HEKXYVoy
DuRLtiFXHZT7DCZM5LDYWcevTl6enzGDR5AXSNEGPa5fB36ZP4+ZcfWjoEUp
ZeuBln9zoXw+dzT5noI86hdZiPcon91qXqxAlH1CmbKfxL5+IDEO1nrUf3tj
Btny7jk11KGEY8iq88+kjxKM8+2zlWhB5m9vWQxXevNJH6fP5RWBOqxVprr1
YZ0dsPzZn94LELeJU0w8IYTfuDjYogbnls73gXK/LCBA1n7p0o7sQQjle3iM
Uj2qyBuYiGorfv+gD3RbcwAkBbFaXxU0hl28BP5bj3IMkVlVoVtyn5Q2USL+
99maGye0ddCqonXfjMSgznnzELbZpXPe416XzhgJq+iZJ9Dc9RlCMegjSTt5
iQlja9oSl/dkkSIRJqjTdaqUWMfkWBWPfq9I/tdKnkI0yZu0MMU/Ig/pI46+
LlrveFiMc3ZwLk8szRnT0BaUaPiI6+2f+OpfqAoROhViialxSpapTOqQ24LZ
pAZAs8mqsfTthjZSsrUbR36WMUSADPgTZw110vwzNu07br3pbPVKFUlMnmbh
Cj2Bbb2COkfuuQej0kO+K1IjEdlszGMGj4PZCpNc4q26dCg1ByhFdrroX1R+
tD8nEJaGFZq6vkahGRKF3tT4FKV03fJmelzmTXK94XJTa37oX2P3x5quNrnE
+JglDphvdu9ISzpbUTu2+5XfeaZouzqFoaJA4mmQzk6zKZuy499HRflFNpDW
N/IVxKfeRLOehXQE++1pK19YMQxwMk13p7Ege9BWfSfAA1rGVfhlltmJWBIn
K+VQxb3bO24wOdFTLzbGXmWmGWb+wWIF4r3LRh3n+KAR88QPB2foU5QJBvbU
+S8fvewB87y6C1YTQ40js9mifIjGyy/6jHOjVYPGZ66n5b9nmKQqTdeLz16x
QXusgdgC0gEDDAduYXdp2ILmsKywq+rUiuA7G3f8GOJXN7Tke7+sUz+rvwo2
lzi3qzd1jqFPExYd95RFXeD/XPfpioIJsSXSRwiYFO89P+EpxtVsHHxAna5w
sze7kW0NIeH5u2D1ko/UQOpCOENwja9mjLyhBcOkLlM+YjLV2FvhaVSDysn2
OgG51E/vSiFY8XKeN9ksZPNR2YVTLQ1NLpFmO4VyPBTTfleKWxXIgNmOvIOg
+BRddgplxOl9IcrRNoms/ZrhCOBwY0BOTJ/uvDaC3r1zb+D4OVl/6lcEBfXy
dYcyeS2hpvpPqx6HBkccH1iFndfeW19mMDQTzHAANlGWiFHv2jzBNz4LtxKp
5+YB1+CSIyh7EGq0CvrZjoZOeCGOUSAmGIpZz8Q0GWviWKbrADDtavHBPDh+
+adljT5YCFR5blNgU4O4ta0G2/xG7/V5u0oWGDBOE8tnamw09Ggo3yo/B1ep
NgEEx/5g22Qq4l6zcfG+x8j5pzUpUbnf63w0wd22MxteZN5sJIBYpFesntwb
usYlx/cBmjMcl3eZyrQmga9x8P0VKsKzWL/CWpgrXrQKcj9PDi0SM/4CzOAK
dkA4bj/9084fpT8DNUzTOe290sX3jF/Voyw7vhoDpP//A0obtXA5NhWK+aQQ
3ZE4LxdS30zKBWmojlJAuNNhuvhAJ9kfLM0XwRqXWh5k7VyQMvxGr742AvHs
60v6haVfVkvLYl5tAhmZDJheSTsDVnGO8tQ5PSm36RwtTstW/W/P0dGniDYj
8PaHSyxsCCp7oId5wr6xV5fh0WtmCXCHpU3usrfuu1brO1vwELQLq/2fKJCP
BS/deqh2IPwBnAlj83clC1TAckR5Ui7xkOR/r+K2a8vPalYIePZnvmtzJAs0
DZZg82punNyRuMBm6oQHAL1aOFCbDlRzcag9t70XhcsDB+z/AEZjeAiZ9rfK
A0VYOanCk3z/H3s0RM/aP6oBZROiHzcUwDGCp0C82SfVEkSMBlk0Nr0bNp8s
UJ153rNu79Rh6/bozYjEtSLqFuMcddYE8sjdVbtu7WNYuUwUgedqswnPVVZR
RA9QL/A0ky5y+VHC6DvwT/CWv50MKAGr/jWd3QIgjmaS9SaL5thU+rprmYnb
eXWQjC7Ydan2gm/6zjeCZ2NIoRULV+pHZE0bhGa+rU9IC+CT+JY5/vZx3GcY
Us05x6qdhSU/bK91wtHx1xa/tKDsRqLCxX8hD7R8Vs+Wftsx2ceV18qb0epr
VsqUU3o3kAFvjy48x2WVyi06oj5Dtcl+SjNKgKsI3xNsu+H88CvMvCkWaMKU
AvoyQXB9WlEk5aUzmFqS7XYrKhifRtGEGMhLSwM05/8Z4/idHJQhlvMJoVhI
gZnAcLTY7sC/U2/op+yORRgKLyUO9Ufe7+G7hc+zsM9a6FhU3r3MYDzJ19cF
/0tzlIqd+vnUxfrSuzaze8IQ41Whv4g2PNzpOv9uzImMFXLCbXJfjzJ8Rivr
FdnIV+iDzWDCFzWopmKbBlZNRRpOQGBm62/yMdUSI5XjYMADZILEVv4E2gEu
ikw7CkKLh8y7jfrE8kSHrbpMA68VLZvvMkq11hneLP5u6z8HDiTw0fEzzX5x
b4g0dvzU8ovVW434/DEI3i9KT6b9A2kQ4S3H927AN+oyFud82c70KDGQM7qY
T+Stoq4RGxofJxs79uGUhf4HZdHkT3SL/1FNQePF+nYvUKNKVsy5Y6A/bt57
3JXHfNNPb35TeqkjPgA62Amdl588Xaq/J+9e6MgFreEXkbZ1AFxWC+4CCVpE
FVca6FUl2ZZV7h6B+wkagCQmJscWiPPulNqFL+YszrsL20WTa5XFM/Can5Zs
3dNEHNeNFgN9UTxZ+XOeGeGvvu+DFC4PBiiOXi74Z7jO4hzI6ndJXmpXcO7L
KigINTA0Bfl50CeXu54O+tXtcsRBPaQQTPBBPxjNivfMelopkbsAQNeo67pN
yD0GpZmL9aYnE1RF5ynp8Qu0LX5r/+wN7K5NpZ1uGsgJSLt/u2Ancc++/P2v
9JtZDUgrYhOgPRG55McewvPjaTJCN2tV9SGkvvGeS733CMlLqjs+wJoLF5+7
zmQ0woHBXczrGkVqY2Ew1EvJKL7BvaLOTIzJ0lX3I0wZRFAnK62rwOUAyUyb
pyXJadlnQ2kp19pi8vUeXTwWqwcE9HOWxetOiW2yqGK3XEZKYxyZTDg/D9qq
hkE8aDaucA+nRBQCrPTBx65XglKzmpH2RyT/Hx7ZNXlii70d9ZVvgeT+frs1
xxJuOJ9rRU/8brmxu959EtUxWQ9kAkYv2RPsSs5k+9krnHoYQInKRESnKSuy
SdpqtIcboEP+MYt1tjaoTG/fUP7o82iR+ajutHw8FhCEhZmyPrsoNje7V3ed
xd+y6Wc29RmALNESV0m4stDSAIxfaqAhiKG8bHSTk2kD6ia2XMEhBxc/KDRu
TnZ0GC21/EsO1QF4uGsmOqp8NKrnOAK6dWRToruzwfwdfjOJO0kyV3F21pOM
EyC5IILB5cnfadu1YLoAda79HWWRO5mPAlo1s1rtNJO5YJ0jL2QY3AIrmPb/
DgOoTVWYXb2+LyqrsKCa//5pmoc2cKJdy/obuMuhnuUnIdazWpCGw8nLQ1RJ
JcEqjDEEtTle2fMDtEDMakUK5UPkPhS4B+XbrN8tivhJhJ8Ylptsm2Fxe1ZH
F+2etl7fdQ9BIod/P5nUSeHgnpOd2Fx+qt/v317LSA8ZXukcHFWw1drfmY/Z
dEK43oOGZa3nZ2C9p4e9R2IuIVUqWh0gpnMyjPj9a1ZVZeuOTsX/YBpd6whm
PKM7gKU+s3i41hYV8FX73SeIT74hUAKJwQmz7CFvg4bzip7shByvBxYMGWQ5
OwX7K2JMY5btpvfBz6iHyzAQOIFNBRORg3+rgAJtUizqyXtAnXCa4FmE9l8J
8ljmsuFTWgMZDK0+JErjKjPYQsk1CbNr+K8DVpBj4mQ7uWCXeE9CgS5ypXS8
weN6mLNfljeRdk22j7oaJf6dXE0v1LOtc4vUkzMUtYfLOqa34g1yWMyge0bi
v6wRTNOnosRcvU12fPqeYYfOybH+KgU23rmH5aYaRh8H9/OWIDd3JM2j/Qhe
kNQ0ywC2klKZZ7A/cLJ5nNVTIC/8AQyNui7C+Mhimh9xaW/zcQ/D6zTSeVDi
n3BH9FRCRKrhpRNfHhtTOTtjmk3AguMZUy92mc6TjdyIMKDBVIeE6SPnhO2i
T4HG04x2Z+glgO0ts2SWup1xeT0oM+9AR+Es5vw8roo7uEjsnnSkrOPELnN8
ruanqCwbkdLrxvMHOdxmIfNPB8EoATyuQSzEoRR7K8p9XC7hG8eFpXljXReH
9WK3qxk7XWH1e/GiIQyBWZ1LZHmLYmb9rFel9U708zMH92CfOBRJ87LR1N03
e4KTaCu6aUvHJdbHCWesE6071I488qwDAZoEAM4PMPAH2eZa+BhrnMHEOqpA
7FJeZP2um+IBIaq8gPAekA28I3uyj1SoTkk0Iaexpj70r//oTYW1N22z2z7h
1QIs8ELW66spvmDlxXjZjpAkYgY0vQKeEqd51mILVcGSDIg4M0pvb4apCYWI
KeY6Pc2oTGq5DVxD47DMIkVNq/jV4NI0nR8im2/Exq/xAyruIblXumR6Z+d2
eeheaSPaRGRhfRCWScDoJIxqlYxr6Ss50e4zVjeK2h+RPgEuAuTao700JLMZ
KsVVQGkf7Vev/Xp6jA0C1zfqdDLstKfTwgFnD8qNywEpOFpfC6UxeyFkP2fy
1pDxWzyZd1dYpQytEkyqZtRWjNoX29tzh3iFehI5Shnp7M6JpByIUC3f26KH
SE7VsTkf/DITSro+We4FAp9yNXpBDdROhN5G8oCLKYvz2ffjJH9hRBqjO6+5
rG8Yi99+0d7pxHRYC9xajMnPKLi6aWQSfQBBDRAdveCM6vQ9kgPlbeGnTpRm
DaVohFeiQdpJvEu20WEUQR1W3MOOZr+spEMs/nVPGl5vcV8reggLbzHQ+VG5
wNMkQL1Tsc6qbGoaMScB9A4AwyX0wurvTIdmIEYHI7ovyXZBpceGgDCX5v18
FHLfs5WACCmkq8pZVqP4y8cwwJZmP2xNz8REfVq34dntjBk+VY6SrzRuy/t4
NOxQTl07qqzyfGCRSxLFW54VhugHzrnVotSKL+xXJ7SNYYAup02FuTcA9IgU
7H6woXi/NL3PqbNWY1Qtv+UH3QbVr9daGqwwpZRD2iD6PGx7U+JpNGyVVnQh
I3N7zrBP2SMcF396D+vvwxSrpwvTpgijvQg5SQuXlQaZvcWEw+eOB0wleAux
6ZUA8ukYJAM/QsA/S5iOn7A1B9AMhF7/7RFn40pGdDinYSFJ7dTIIlP0whpd
zPsTTy9jahbp/PHVMWmE6OHruXc+cxIyFF0wLngyx9U4MZOMgRdJ6tr1lUrB
+w7jvjEpW6JuASVreJmsaS+8zYanoN+LpGvO00CClf1VbYRMBU4gv1h7zOaa
3Zjjs3jCw1w+37LSG5DDDp3LZJBa7jFcfBvx0tFqGwThtcK6VWjnBsAy3bbU
o9+d832GgkL1X9Je45+YEicz2pSsSX2DSu1laA6LEKBiHe4dZbjvP2Z8MjQH
ouqlnB/7n5ypyTkH6U/XLpfz4ykWWwWm3N6hdxCIzI8gnakMnXOEvrEnci+U
picvDYi1hGqWgximIcW9w+hCazv+xfyJTv2ymZSHmhJI1JyPsKEFDY3ODPLo
LoAS16rYx+Qo8jVJ8v0ExFH5vPGmr6eFUoXtgbKZtU62WnuDhvQc5Gp/V3mm
9b5HZZvpws6g3+u0HiAAf3efix7i7ECaX8SDZj5Srf1TQo4ae2H9bkNIfPYu
ws7j5sD0maX+yknXFGXdmnKcCXyv2wlbYGfeMxGoqEEP/WKHkO1JFpJhlj+K
e9Uf9GTbKM78Hs27YQqIYWCib+C+HNkWQXr5o40eUw7H0PwqoRhfLTTplra7
11o+/N1kKFkrIpHNHmD8+XXCxrRvlLVHHqlWfKVzyDrHPUwe2ckXEsDstZVD
Ykg8kupqf2vZcE0GMyK5HZBa7rURChj7a4YfKQ+RS4cfyoo8zb38u+ieDVc9
LHSpxWuzB1yVQje4stOeuuil4Axn1WF8kQWPhJzihwuqKAieffnoKfZVG3GP
3HEyGM65UVMtSncbMLv4tAxIzmc2io++ulioslk7FlKn1UPv8YopexzgeeNn
ytK7zO+zPD9iHoLEEcB6A7fnEvZiWWBcyaAKEKZduTXRwoTIEugtNzzvp62z
SGO5E3Sf/d+/bO3vc3Cpkbd9WwiM+AdxxaapuFEBbmmamx8cy7GF/zkclWE5
LbNoyP2jW2W1qlcCYm+J73xdW96x6YurXL2Oug+Ou14FBKK6cvZ2s8hN5XBB
Ejc8Zt28sE94QsajBnkRbI2mL63M+kWRtotCQYkApTZTecxBLQ7EcuNOoJsf
iQyA8Qow6Dl3PyIs4l0+Ao3iMWEQPjPJ9x77qBlEkH7rx2jg4hioDzRUheQ+
BD8NduMQQWurnjjm7fDPK/yuQHzzDOEUkky9Lzp4LJxAgLhccJErZseiY0IK
ssFjGHAf3blZmmpJ9LLSFXPVwj4GGcwTBDfLybhdqX2JtZJYEVAH7ofy3kCM
wT2oz5TPNoXNw6WLJG9wgVnuIEQcg20YlHzrCeoos/Jho5ce5annuJYpYY9z
OK2CETwTdQLeFGq9/nVW1m96w8kr3fItvBScSpvsZRADMbhr1AfLZO41VYES
oFvFx5IFlZbeZN+vsFug71E523o6HKy1wR+jwcOA4KVRjRwW/dIQi0ZOp6Iu
rXQSscgSEIlUBuAzAioB0wAjHstgQ9LD2+txpoO3OUxSri+5H7B3aWbwBy9r
UUaKoM3qATuZKOLUhi1bd3OXe+m7PSFvJ6u6wY11wfXcn6KVKoCBq1hkyQMD
YG8LBAqNr7ycHaMMIhiufyZInqwAcm0v/3VDjpjd2eiygK2JZoOx5TkxfMi9
DuYRuYXRJZWhr54dSz33RZa46A65ySxSpuJjdWRlAYUfovKZllXdzteyb1lG
yq97A38VhjePNRkp55hXfdMv6K4LukOkQCnT5Jl1NpbUIAfkGu80FERCY+3G
9GBvZrpUZYiTV53VBVgaxy5HAPHzOzH0z0Wv3u3BPgiwChJe7p9eQU953VKr
0HQ2ZuMGS9JM1yfJpGFKh0c1BGune61rF7ghLaAyUPPuYtJqDNaCHVtqFCvW
QsNYnw4wg5PlUXmlahRocZWGo2lk3hfIwOtVVweOLGEopaICkrRhGNMWh8q5
clKxYg5L3yChu1R8kb+ggp4DHsjkLb5kokvJWNgaW0iN91LP3xHhRqzUpU51
7FSQZ8EpiXB3R3f/5aIw3MTXt2kvtktnWR+jhNGf+TOCGd3X4PZ5W79pmAM5
wvcC17l2Co3t/kotAnCZww+iY718BvCJjW53CMcHfXSyruW06mF4yckLM8MS
HovRsf5anB0aD63zaqMfinvtfA7UzYbz25wmNNobNrE0mumge5CWCCGdWbVQ
HByb1NCYIBlPSwvgSg3k+RlaJ5sQJsl8QDSYrifNyCcDJDzl7is/6COChnxT
ZPqyYOqiQYjKdPD8Gg+LGvL1xlE8imk/KfeMxp/azu3cCbWgeZCROoP9cXQi
tsSxKjwmm4pVieja3qvpyrd2+gttvmAKfVYGz347hcZjUxkzcGUT2HsiryPs
H0nKuB+EVkyM3Oqsc80tF2KxzwLGzIRZ8P8BWXXSo4puUKqf0YJJVew8Xag5
0zf/DyAekE8DxoE2XS/Xd5vdeWR7zAV4PruUa+4Z9sitUofMus5/G1m90mdc
lcUf/LzKg0LpWaeL4S+3RCNBEMK+qm3wZqauco19yUKSql1iLSyUqNfqldS7
8Y+TABbEl8NhQ2y7EjASneLO4wynt3fDPhj+pjy8HbkgTLm4l8ds9uUtc1Cf
cde4WgBdM47RWhKYsKGpGiRfXriuZDZUWmALWrKOAafrL0Xm9a643xJqx3yU
16BpPjjJhA9vIAPtjQG+lE6iRrjrdiJbikZOz3h8CD1Igl6JzKcAn2n1MEm8
pedtJes9+S06wtkq6n33V+iVOrZhwg4CDkKA1Pax9OLKx7mkZ93rNXeWHJwE
NyIt1ymoBKWuviVssbYyZ2zMHUr9fLtOaMt9FQwWp81W7nfvgzMb0MCrNieu
9ydNVPEBYYYZREe2qWJXWFoMUIjFg68iFiXylIV1Ilodw01ih8uhvDSINx5x
DpAhahqRRInes3hHsa28g9nY4O6BKc1k9sWgx9trWMLnbboErjBrFsKBtnxj
WlnvJTqVT8Oa/A0WMLWv/Ew1WS+4d4dK81lzLXNyDjPBdJ2OXe4iWvl/gBGv
HBrQNYOQfHU4zoiLlVSjooDJ1/L3pjuGBvtbQtwiQFM+Z+C2ZiYDqpbodLei
ugZnqBnCH8L9jo4osE8Qyj/jK20yZSg5ZKitUugcho2hbkx+tEGvY00tXrib
xrep8sIXjm8Nbtz9xlLU5cP8GWr15BZLdiyFb8p3qBEps2CeUw+ukK0hBee/
kle6JdDE1qKTRvOmm7UwqFFaLsH39ZfLNhNV6OJcXy1kVPqPJJIznQoLoy5o
DF/nmaWEy1WxFABuB7A8lu6am6yMxATWzZdjkza6WSLIHJupVpnwloJJ65SE
989D8gm7wWjBoA6k8oyxRh+E67znEmQ7EzSMPNgWq6k6/2Q0RCEyWOmG07BJ
fbdRtOLdE4IyOj1tXXupBHr9UcygSRzzuASzFh8PnIf0dGp6nGr0BI9yaSG5
1WqkaEtuYcGMYXLmONAFDk6zpKbX+OK4W42YmHUGd0I3uhWNFs60ZWXJc31g
+q/Nls3tjOVHuP01CShggfXV6l2oP0TjZeft+JjpssprlZwbuIPcBkhrEnk6
+G/g3vpHsamZga9EtApP+vZUYJiedhYZirwpEh5NJ8eR89/quc/Cfp0OKnLI
84lbXPlaYzTo8eBobCr25vpajf8y8Z0RevroKs/Idau1lYIB2L++YHh8EjUi
A/Z+/5qIRvfCEI8mFPLvFVSzM3y5je20MbM0zb/kOIgK0CVtECVr0T4K5NDz
R3TgObfmaDzI5E9mYK3IyxURetGb5w/j/xI0sYnoFuKB+nkyiYpAUAo6Q6KK
nfXJH+PRJOE8Q45/i60nX/eJR3LQbCxdgNkgo/QwSJ2r7VfLmDyMpaUSA6p4
5gQuRGAEDhmCqoJSGj9+5Rbgm9VE5gNYIZW/MhG+641tQxU9378WBP3Xbwho
vEaStpLiw3rVbG4cHmcU68PBfRkoYSZORG+rVXqmiENyMrtQ9IBSHwzim+ws
Bs3ZOBIiTGMnx53848xmmIpcQnJQYjUpGSI4muI37CZpcj11ZGvl/g/8bKo0
EgCFq0Zoaw0GauDAx7tSv66jjf7AoECQskIMr9cj1ej5O4wYFVmSbx34WOYx
n1oIIgFn0ebvIGt1ueF0hDtPwtweb9SGtAJUKgumXkfDPUP+FSIcnA3L44GN
pc/1yiYqUT5EqJfjFgcJjQKAWD+hRDrc4LHQG85FML4MwZegr63TrtR+KgD1
LoTgSEEBqUoqCTgqMZSixgieCih/c8dQcpZUGa5lSn7Hch3PPPJVpAauVIxi
vG1UK7GVFN4QXZtTFpz8DAtn4y31rIinkmD8rI4KvluOJ3HB8fBEdFhgN1Dz
8ohO8iRT1dqmwatOvuJF0GespPMeMhT4gZtBdbZ7JNbEZyCg7N7ofQPrRAsy
Z7r8yP18NDoQ98HXIAwRAetxQw8uB+kuSBMfjIrHAYVH5LJgsyDxkTjywxVt
DLHlWnyv3+CWFJAONLCzxs7oFoKDYnFNSH7peJ3N72XzGif2Og0lK+YOBzWm
wtr+MNq9F8TzgO1c9LU7HHMsoG8UUFxWk3oVduqJERrgKsBukSuTV+gEiXLq
n4J2QeDE7aXmhKfqhSbYZKmwlQUxvAWLErtLGPUurZxXrfnSvHNoNEI1Sk/8
WLijNbQZhqQDCPpk+6YAA5xIy8wO8ew3p6xna1kgAYplhkqQ+IiJHluVBDY2
M7gdi87Wvzf5z77lI4l1EWQ18qjE4lhsdsuHNHeVYEV/BGpSJnFoyEg+ZXVB
CIM0HHAajw+ArkjlsYqqSrh+6rgjuhOmswtN0FP+m1gad6TDzxSD7dUryiAU
GjBCWB1YEvav4cdWqz9eXuJhd3hnCMLmpPNz3jhqWAMjBGH47Cl01AX45ioX
NlqrH1+gQO9gFdwHE173emh6yM5+Slmip11al4xqLVBEPkJzbHAO1FLAFOeH
/JmBL2cezQMQQMSzIUsuuqNUU+hkiA0iO2Lv8a4N3CdDU6MFIV8ndn3JWZBp
VI5OSz+CycD9svlBbNAlO6tTSsjsGUyA3QQXZ5Y7TUmxve8KK8QTjLAxMJRL
vBT82OCFo0hcq13ioLi/FsFqp1K4xmmp+8IxCAYjaSpX9lTESFL6PgEJ0j87
lk6bdhLZV/btkNyu1pi7zfc9OKjpApTUlyHSDFkVwa/iUJWWuzRBMAGYz6+8
7U7vZzh1fyq07uq0RzAEjGkipweta1FR9c9MODjC0/3FqSBZ1jT8hqNZGTdL
Cuos2DxYuQlSBx75bp2Pd0+A0bwHdCQHsiB/7QFhmAwS8mZZ8bwym9mAilci
6kxQgESrmS0QmfklrZwEQ4LgGMFZOg47o+4JePzQXpeMaDNiiZL7q/P21iTa
tRx/+7y0c/JhJTP9hrLIgVgURRKUXzI63Eb6OwEImNsFWjgrh6W5HBYuQCy3
oO8V7PgReAx5ofHWi+YKw7mgekJjAk70OE9bSviaII2Pgg1kw4t/PP2/aUam
S65ZBKklg5TVMyg0zsa9mjNeqfpUU0w5LIcIAKY2Zij/x7G6E4P9eybflXPQ
vm73qmoSX2ZXDEAT5VGfkL0tQx/2iPjDxxZxzjbpCAd41T64XRhguzDth5At
223Il4fQmPEpKjNH8QI/Z3NJOcDWWaRMmosVVK4Zq84Kb2nB48J/0l5sucHK
hHboQVpcoScLDVnv99xvY+AjAxm9imTQXJE6YXvq/CEyGxZ+OoKZqCatilUV
Xha6L1S4xo3qLR1QXr4rurb9o0Zbtdnzon69sUAIdJjaFPs6hqaN+fJwBjJo
sNW6HPh2sVYHnMlyh6BlAdtniDRSuRA7a/DpwXjMkfoM3sWLZB2szNE2RZDa
LJn7M8ga98SayPhIpyw9/H/Wrw+sqxAIb5cFFcNO84wgTvYzd1VHuSsz2JHE
i7oTywZz03IYmI1G/1wCltTsGZRnspznFOncsBcKDgxTnSx8NZrbqjsAXZYs
/eJxNgAA1+CDV8DSYmq6Bve+FGPyEJC9H2Xj/GPMNJIiHiW02GwzmLf1zAjF
8qXKB2Wwqxra0vvXHxmREtHqtb1txYf2scX/F4siEiL/Vb5BscMWzVe2JZMM
u8vGQluAAFtmRSPl8+YG56dWtmN0K5d7VGViFKYUVhF6LXCqPU4hqkZmXPu1
8OdN13wrwXMAYAdpAsA5To1Seo8i1bYzfMlDnDPGSnUfXy0CDk4TIUU6zSJS
lsbwB6KhkMNmrXOgcsfeV8AOiARsYGSSYTLiLTV1sR/S3iArr4yrrrYtyvQH
0TkDEZnTK9WC+VDP9tpucklZf3ldixv7gfzkl7Ibi2IAjGnDydCp2sF/oo1T
qutlmam2Ah72brvisEwe3iujf8T7DuX5dOQSUoCGZWeOWZ6Nhia4IQdZ4KQT
A1f27JY9g/3cZRwm9mJQ3tn+8r5zVpqXYqmeo5GwIPd/60BqQ9jDLpAMLeYu
19iUxPjxUUAIxic8GZNFKk0frlRg5pnc/mia98zWEzP9H9lMlZ0HTw1zYZPZ
qHEnDpYiDnn84rfrVtv8n5oF7fkk6+5VbFgSbLLdWdUHWHuT93oPPXvcYZT3
+aStxMGu8/A0Fu6b775fLTzR9mq/DbF2WMZlLCqe2zas54+YPMiGBO4OeDh2
BVKBQRXXVXkjpiWk6m7ZnQfP26OGtcpiTSNOcDUN+JBCQQnhJ5JUVp2yqUXA
clb1RO4z4j+fYy0RmajMa9YWQPJSfyUWMSCoY8itd1rwFecSaUmMt+2WIDRS
4G+MoL9UiGfc9wjiFZc3LXxBckZcvEJUGFwJoGea39Z28XpbPOw9SLkTwGhl
KizLgwN1po+94Hg8X5qy2Xa4j0qgERwCEKxzXGT/E7f5z0sA6iH3CN0ZRi7n
gXTT0Q8hi1VHeVH5/6GBHanxVogcP1GMgPMik4Jig1X13759aaooNPfB8ccI
+JIUTEEew9I930WvWpsnkrhX4QZpaWnVFcvMADZOx1qY1WEe0mJBlLzeEc3m
BHTYU2RwRDzjB4utFIQeD5X76tQlQ386Pm/eTYLh1bVo0HP8NCVbMlSao+8v
Yu0LlgqueH8kdcB9UVyrVKMOc3y+ryDv8s88mXm0nLMe2n5voBTILXOqbIUt
KeWR4fJrKnRlqUHMpGEgVDb5aqAV04qR+W3hW/B4TPsZ7gxm1najCQtCE5E5
HTT7aQkf1s6GvLJDaYDCeaqI/IRsCjnAohzyXNU7CMAQVEsmERi9I7BKcAqR
04ytA0sptU2m9AM52L99bNPdJts6QzgY38c1/9nzbrS9B5dfRQvEpbHXKLSG
zWg7TkDWmjff9QA/RJf4CRmTnR/mm6hzckbFQLHTbw7xQZ/0zSL+HkCNbZA/
v/5Lz9zRjf9+gPKB0ugsRdXIuXuNu2SlsAU9Tz91qEBE7va2qVUATxYTRjUt
rdVwY73g9eRZpMv+fV3xOSGH6YowcHcjLch3bnyRY1wu7mPGXZDWCUVIXcMC
gBYTzLFM7OWcWoWXovVdcWAlPm5ED5I8Co8E9fbyhP3BPlDyyQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqe4ez9BQXb3W3KYy8CoQDLH7+mXLduh4bvzfPMgyAk8lY73UjmtzGwBhfulxr/gWLNAi/btsrNgt/nk8edH3P9QdZIYGreSt9HiQ+c4lqXgvQSzOfBLHd5hIkWTLvRK1w2845ZI9BzsVuw+0gDCRcMzabjSpUrvpvJ+cg3gYRA4rKDgqOl2lN7g7/V6rDbK8jeujS+QQyjEqBSuLzdPpTMEDdGeVwHak6jaLuK9PQBK9SdiXUa8rYF9shRGWU1w41SLFOwSKBbdXAcJ+NPoYCbb2NKxuoG40O9b+HiCKHALV/OxLythLZxU6b5ASjMd1sYgQ3BWNDRNwaPxYZQUQWTaRiu5AyK0z9o6hLMDm+bhjT1eTF/pmIjiBk/6gieHpUWu+lBq9bj+aLtsn4zgVAOLTGdbpFddxrhNXIOmvJ5driv5Ey1cK0pkOQdXjwYzo0FFXV+NipXELkqYNlOX5BFv6giZmNfpxdq2YJRwO7gkUdHqbQsD1cYK9imN62IDTgkx0Lm1LYALsu301C8ljjHWbIs1mI6e69hO3+pxDmrAnXpere37p+G0ynZTzls6hNMvT0IbFE1KCJVExN1SSszbl+1sIejqONE5QnghRjDIthtbv2hsZE5TjDgmnuEYq4gGSkI4Q56lUtQG820tBYCn7rSapS6hJ0Ce/WVVT3zTUzwuKlnG89Kifi7K4uGWA3V79BJa0532Tv2CpXkoE8F392ATCOCjRwdSn5dgevbDNeJl97oHkpc/Je1CIIR9TdYz7KbTrq0Za1CN062uolVZ"
`endif