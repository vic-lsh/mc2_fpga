// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
1WuZ2eX9sqypHUVVIakMe9c+i4bxbM6cg775rKvBMYqF+dzZkAHgY6mb2lXx
wPX5dxj/9nEVkI3JuKXnNDYtnogwFA4SyGqUXS7tV1fLyxbLDnt5K9/spfE7
vU0euZ4g0Z/nAgJM+udIcy4OGTNFVYAw1k3d2OifZDtdpRLDpJPgpuixN9pY
n32VVp0HEmIDNNEa8OmqCFicsvDPBgta+OUifOKUx+afaLaB0vaIbgxKeYvp
svnt9X5i1KPFz52L4xYSRz215oRHL38TWUcU2DHBhNaUYVKrN3ZoHYvF5wRT
+9A/2L6KeADYowe6HGUAuWwkroM3hn2tS37t8EWXDg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fa/CvQ+9+Pk1W19LsNdHYGhpR++763Kct1hOwqem9KyTUz0/PkqLRNaHUMde
xfx++Ne1eindX0qjxdtpe/Bc3e6rGx42+Qnn/IjOIIpZC00LaqR/IMFwmuA1
pzLO6hGhx96AU/k4eIkZZ4NmwhbWe7nbuq4E6qy5EKJ5TDGNGxrbazl6/Dnc
o5iJFbUGlWqq0to6pVtE4SkQTUtRcbmCuv2oxeqKm+4wPR/l8VqhLgIyIJXN
+lNDkXdB2nJO84l1wIwdsC1jenkyGts3KJ521nVNiGw34zpCtO12jPxyvujo
oqtaCl1FMkpf/7xZ/EpaQoS6CXVHj/GVzuZi/4N1rw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gwLVeVga+472KcUav98/SVPJqRydeiDSoS0LgnXrXW6dP2qyMKw238BukuSl
g1hjN+tbf2jMl3lLxZ1+b9mVFWZB9QsRKs3D9+WFCb6ByT9eIqSqldDL9V1x
FZ/zHE0OX/JWLFpqY0ZHAm8yLyP7Wd9MgwWZGKVJZnpLTT8avHHzSBjKW6ij
bEMj2FVOcOzE2nVIMSQOO3700TzL0xGR2o/zbGEOynRxZ8UME67QUv161aqX
5xHdz5C0SW4QL/1ZGH/nzzBTRrD5w6rqa6hKi9dZbYjGJ/UUS5EMFp1djAKt
0E52TkCsPHXab0kgcpE7WaTU1o5yZZbiNVn/Lrc2rg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JCiVKdPlxvQOu4UMfLBvQJqM2vjkOlTYcW9bJ4dxtOBmOoiLR9uPe9OOZ/nI
3C2tdcET0IKeKr60QlGOQS7oW6tzvmFNYurETMxgZxURWLRm5dAR6w/LQ+13
B07oVjoH1R/BCzCJSA516Y71N+sUaGECoR4SBk5vcUNNFF/z2N59Cv9NShwk
/yuiB9bQf1sC2BqATrv0G/fh7gxidgfP9fVq2fmnJvrCZPNfTlJRPd2CzkmL
aktH2ytLJO9qlQzMv3KIJCF0ZjkZ9GLKFlWCi6fjNrjSagVS3gXMPP8X0Svg
/jjFGLlj1n6bvHR+xWSpcXH3YKPeSIQSuFAUCBIgDA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Qd78kTHilNO4C9xVyvhId9UlNasBgi9CQiyeYB9fusvme0CG+I4UGEr0AVKr
ZW0QiMXq1godn02MGuIUMEHxjoY4DIztyxmVoTc+yKosqho/gtczpfDqL4b8
UtuJjmgZs8PYq6OR0xYhWBauykCKUqU3Xn/qAP0tGeXUFhWpClk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
spCCGR4uoOfquehcm4hwRX01v5PvMauCpbKrY2i5/o0cpM5PDH/86InFaSas
lO3kipL/SGhUTqkbIL+TmI4UchY+7Ptr+bglY7UTP0Ul/fMAqL+90xcsc2hM
CD/bHvXsD1afw/gLfVNdcL/5AbFOm0OvANSkOAWwxpxsILU/Pdzh53ed94+y
Wxg4KwCs6Dv7AoJHntwm00OJIJJ3lXuAbrQUA1QWKTN06xWf+TwM/oAkCf4d
iZqGuXCGj2Mbz/I0PbtADqQjuDH2pYORwA9jIrULvWtcVG5i9u5Xx8p50Vd2
l7Ru1YXPnasrhuJRsTcMKW7UXu/43fJScqWgQX5UexNkgcNYC2g0vDkpzVuc
RB/hQ58kJbuTHGb0+A8nssjk/+SKuGUBvss8AR0c970EUqZ4JDM3e5njny2j
roKambhX7h5Bl7skxfX6JstSXW5jfSvazyDDRFQSEUeDfgG+cSu4CAovbviq
L3MVK4tOl9+9GBme/rkqkPL2Vtlx3qLT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BlD2zqzgKFbq0Xj7rbpYFM+3zx/S7FY5/3APblwYMzXTFQkMG/oUH+LQenpe
HhVqTpf8PH0rhtrbcQA16TU1S8yx4AkO+8c+taH134BmdNA9BX6abpBpgGBy
pxac0A3WS7Cloqk9sCUUfn/ooPMh8ZXC8FM2/r+2RG60rjQd80M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BCaMhjnUyf3tU7GrZOL1OSVNkd/+LMDrddQClZXGZEsUg2KXDBpDTucB/0ys
0R2R3X6KHKl7gYxiKbjVlve9Bg4SJlhnlWWNEm1OBaaLN+xyqI2Xdg66Cj/D
N3EaRYHagEimgCw1wdPnTBUNaSApnXb9RMeEXekPDy7qAZECbAg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3264)
`pragma protect data_block
iVgMGwS9OAT8fSh+WV+ciQMNrK/hDkRFD8pxnNs8BFyFBuw1XEPQYfxE6X1U
vxP5Cwm9a5Jxca6ZPVbhLwRwQHlqFSO7OMxRmqFXYtzx/ihihdHZo5G60aW1
xNyD/vYlutVRoyVH9Yg6VhytOPHeOhAl563ddhAYLeRXF8wtfc8OFqw0Ewle
e/pqxLh4ldA0oBel1vuyiSlJb59kwVeg0lP4VWhc8g3HUdX7Pn0ab6rWM01l
pcxHYwxMc7ZZwEcLvUiJF5oiZeLlU94y663bcYVerk/zNI5AlocVvv0UsNk+
Bb8J+uIdK/WtFau8DrSl3q1p7GiVSgodicAXBKgVr+lTpI0NIvTDVLDiRNfv
SY2Dp/CZavvNMXdPrPMiyXKkFpPuRvNWvMNbLbxz01DaRIy0C5eeokhsEdoG
f2zjXmCV64BVfEwcHW5P8ZFVckawlstvvVAATie6hiA+KcIUv7nbVMSEI4OP
zCrASt3HQZqK0gUJedT9PbXMuaVWLQdcnFlYoFXxIlCky9BwjJKr3FgdoxWg
x0ZbaEbaG+8VpacMrcVd7bErXom1/QnGbeB8bOQrNCptboPMaLqk5dSYzGUt
RguGnuraAXhY2VRAzMCEaZvGO40xHvSIF+nEiL9YBuyK6tGK4/hPAshXAOR1
p4XoOzg+ku/mhEJyGwjOVl6Xdh+K7z8rYMFJ5CPnQ5Qg8QgwDS3hye1aQIA9
k6dAD0bPCjoDlxQ30ys4IO+8DPZ97W6WOPIE/sdYLwtlAjv4CKNgu0EZUMv7
izOduZme99zJxjEUw0jzj1Q02oFAxeOyUvkRNLzhRBXLNXCOGj1QxJA5hxGt
+/wqm42+GyLPhg3jqG9eqtZiikLWYrwRvwz/sm13qh/ldZAZ3+fYc7Xx0kFO
FJILc+4cDiyDLGQ4UQok9utlwhqN+sujxZ+ewO3xhFB9pjOMEoigIYlEosqV
Me95R8+hNTu/FrcnTHZWlS9JdkOakM0PGnsdnImPk9T5RSEzVyAGvkwYtNzj
kd/69YXOJ0XLMuahSl5z0S5TaTiq/1K6asJAsDKGXVS/oOiBt4OadY1mb1Tr
fIQi0wgCnmzGAdDDHD8XqjLdQEU+EECFsVMfQzu0ur8H1PhGbeKVHV7jR5E3
8/o4/m4mELRAh3nuCu3spAWr2U59qPI8dXX6ni611ndC1Bve0lvPtyc5QghS
RVlz0a16e//g49oKbBKYKLq+u9A/hfqHtR2HHKUl/qbfTTFNwI6/jfUz1upg
DCmK9QWWz0sQyg/IBO6Ch66CGIcJPkxysHlhRXLQ4I5WHMlKr04lCcVcBwAP
hjXxHYB4zFGzz0Zc1IjHuqwHazanm4z8C8aM/lpZoSLUgZgbTGx9zYoFtzjW
siUJR7RaZaSji90JT41CvBMw5B0FgC1HipM9kIVFgb34V4H6vnXJPv9G9eLV
GCrJ/oZRcY+lI1pmtJpdFNYlqBJCo+gUa8Cswp3NQbopduk8i+mVS/jeFzeR
68SYNIPKKweHVTD6QpGQVEJfvIIbO4cEE+SLxv7r5Xa/o4Mpx1cCw09MPsND
JpHAJzed5UjhIGGc1uO2GOxhy0gtyldoHHbKjC3rRHYK/0rONTbvmaSIOKMe
9Wcr4vfgCoUooWTjNhTmF544cvZdgm9Lt6pKKUWFNoqWJNEmh5e7UWPIcUPD
ReEdiW+vzc/9lIGyyCRHgGhDa9qjgSonK7KtpzXvtaVz9GLJLDsroP/yqxLS
xyqoVt136BrHGejjUxZYpTHl6Vd1DcWpVyxG4OWFqQsB/JeceUtNtxAj01bg
PzUQU9Ak1nTOgjupvxUtn6Re/0OkyPMfS42b18OPYhGw0txqD9C1D9zRwkA4
sfJPvLdiGgTq9evsJQ1yI+XoPFj4dTeQl6pgAKZagF3v5s3wOLGPWEm+qTKf
ASbHYMVwcHpXXrVsOdP5KBO56SVGKgSV3La9GungvKX9Ik6PdzxJ9xma6n/S
HWx6L968GUefZkR3VS6cHWCmhBAorfD2LZtVFvMZYRIgtOFHGucuXrTgPpNf
HqZiDgtPlihPRNrKJ0LU7xguaoY7rRWdtJWOpqLa3b68lBKx6qdBX9xwUjfl
Pus3ifS3k01GZYn/djzITO+mwsB8LXbjODP4EkwR6F2L3UpWMpfka8nVRZ3e
k/YxYl5jrexxAamK9ZNhPFFOwTy6Lpvb5vcPCRm2fnE9bmkwGZhgTlsxh+Xm
gerhn470GnIlyOupPArq0p4uihtvYFHVNqwlKGojCmLfkZOQqXh3xIsVJqFo
7uDVXsxkxgO0s88iC4bR5dRhc5XS14dxtVqBeckEcK+Sz1WgB+RklFQFD/Nk
UqR3BM8JMiv57blOogH7ehP+7L9wEnBOi3QTES+tRro+ptexO3YdMZIVkZXD
yOD10K0zZLHEjTDgmy+gAYwihSf2v8dQsuTqFhrexy1iI7dqXns05TrQ6OWF
oMx28lrjopsstvbvG3V75CLjUPauxiz+RNJZkrDXl9yFf6OyjrblDTLhMYJK
nXZdz/nIBBaTSlsDM2FNVNNq8VIs0GQUS7PFjw6fRuxUOkuqRVeJB73Og6ZO
YdRE2ULLYKucCMVDkqLeDVj8oZMdcI/gWZwllM0k8bHL1yRljfWnnymBKrZi
k4g/kB7jkJXN/q3WPtuTca8B7+hBJAy75MPLInBqYhR7yCXYTtKqdhJURDeo
/+liYa8WjLgs7LQftB+IF8nopgrVtqi3dr8c8xCbuOJDxL7YPr43bBySnbXP
Vbbki78Ytf58iKC0QhKsmrEfRYlOTs4utgBxFkG8/XwDwZtn34/iK5KVgo2X
anbCQHKd7PltGmaN2/HteXB0FGw7aIl6/ZuKVciGNHza+eu18V4uLpj+sfp9
uTkomoIffbFyKVFY+6/wajh9Yje6jozaHNj7g//EaDpNEUDeYwGMVgMGCB/p
sBYqrlqJy5wH0x33sdWO0slg9Nbfss0Pkz1bgj5fbRYLcSRYqC55KuHbzOeT
AL7LX7K3EtSwzAvKIYD/3DhMDrgJlJXr6Dl9eQU/uKch7Svwqlatyu1nd0Jv
UeVZfvlV70giZrm41exgtEfp5Qdww4q21VU/uXQ8fFDnIvkxaBs6j/30nD2s
i3HW0SieSCeth9yE9scw956rzZmKateVWQEzEtd7IT1Mp9YtOqt0CDBVrHnR
7zUWKm+ClnG4+f/wy56eNvxU1pkMHTs6i6AgNyCBNyj7dn49hjKtpWd0h/Rw
yfONHpRVBs/oKkuO8SRMwDEh27fx26SNxKa9wqvw6jDMtJ9WzCgZEeDC9nbp
/ntoG5Lja2lHu8WgImyfpwWSHaFI6g3jIXke1CHxnbXDA/iWhGjIFMbnmR6o
iIqZeJZB/s/Pra897c2s4ATz01E8vhmnJ2oSqw5OOtCXVsL+Rr6fu9p+pVC2
lMYjyeIX3KiyGKL1Iy2hbUnDkiftUcfJZrc0zcoeZrGQE9AuAigUR3ZEzpO+
lSlIJbbaNMlKxXsiRWZrF0XGSS1mALdjB4cmI+7yrMN+10aYex/RAOIHAz32
s40E2w62CJl3Ce+gOIFVCmWlEmO14lHA9w7S/iZAUEZMD9X5hQS9ki0RCOr4
IKe3Eg/SJdDTCS2g51dtm6kA5O9BlB8Xf3CJO0HLQHJdIS2NBY22eCm9TVQL
gko1bG7pep8ZleFu+C3Bz9V3WdUEsXQqjJN2TlUqGay7P/qokOwGImsxJr5x
wLVg1QVFfv+LLtUkokWpCmyLpIKf67siESwWnrTtp4wIwtuwrc98SpCzSQg4
MFp8iby/ArW8ZfgvG3hc69dcsEe/a/6AJ9Ycwq/MFUsCQXhNiCm+/ecXZar3
JNaa8PGuBNdtMQJZrOOeUNZxLYmEr+qvJpXhYQTg0G+aGeFHduenMbzjY40H
lwFI1Zci41jVKvZAWFh3oOM+0vMiqctMO7sO2i9NPA+IF4CLWk2730HvY4vR
/F755CYn77tW/C7gTlxw4I65Jhczp+DR6kSzacqBpAED+8PGCxJ0PRYwghGc
4nUw0rxiz4d7vuB2LGmLuG2AGFgpaAWbsxh3mtzh1h+CRpYyyN62XcR0mMx7
OZrqmBSZGgtU8sYUj1gfArciNBj/22XlH1v0C5IgtcJ8XdONwSTiUGbXjPnD
2xhl8HDoaXoPhLtmrZawwu1d45FA7Su7tQ2Egy98apf1vbgVFXEwxYd7RBVs
Z8LahEh+edCf97LDskSmw6rVc/NOhENRvyl0vHGbQAFRoQ3AydQg87SWaThB
aoBmX7MwX3/qzLmBvD8y6JWPa7yjoLCrNrJ/b0eiQm9YC9+DkQNOofxO+6uy
kHYWDehARMEXMk+VKBryyNMkXBpk+OZM

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Eq3Hk9kNq2l8D1QCUDafqvRSFzCgqTqcURrzEtzSC1GjT1xUevOeHNte9Aublt7LIJHnTmoJJHLmkC6z2ETPf08AiBDTOs2gFUnl5+W55Ei95jxGxf1haVqVlRMrExfmgczYKj+OY7A+7Z5GyXUzjRhxMGcgYK2YofNDlkMQOFYhG3wQPzmxRs1GR1CN4f/0Kke3M2cSbPOKHM6tbSj57UI0xEkh+8BsXRp0YftoumOr0DqP3ZMmqbMHlPXFJp09US8V7BK6dSSEjhqn2uLn8Rz7LC2p3wiC3/whZTOs7S2afWxEj87men5QwCH6JX3VnPBJa0OSKu8/ieyveU6/rHVbg3zplreKxOFeZrNaE5h+tE4SgTQ6gWWJD7BE3S5cqw0sVdxR6jgKOMgV+LLdzm2RcQyszKimdxzhWXo4fpvf6QISBvU8kSW0wXnQ1FdWs7vdygJddqG1Rf/X/QzHHKdkTbCAsF1DXfgjQxnPRqfQ+68jNdn6WxxIa+xo74nGr9V3csjt36rl8sSPNntWr2m5cvxCUW9s94wAV396hxilmksiAB7sP+nn8bIOUAg/QeJYs57s2b1TPsHfBl9T/8QJaVecHMAaDEEcdcSacq8JvA76X5PWUGEVQMGQoXDdGRGEgKyDnQTSaYWNB55YwMkYWNAWanV/nBtssWy6F6EwM5EhdRNQCFRsJQBoaQIy08rVW8apj/vkg52oPzy6cgTwl8+vGxVboDqc1hidL5jyeS0925kaq/SCZEhmwxhdcVuX27fFz4/lUBkks0KoaHu"
`endif