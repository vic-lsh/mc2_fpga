// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
1C6Bfhif27CifqtoB4t0Q03cO4PLOScq5hIntof7wNFTR3bEOtcoTkOvKcAf
T/h9+Taph6LIK8Tf892CCmVyoBdfADfTtOoxiXDfiks4ukhux/aFkvRhNkYe
WWaNmUiiN1RBQNHKXdzeC0b8gFh3jskj0RZCXGQADcbaS9Le7fmPiPZZCGea
iZMDmD8ZdC7kjD8jyc1WVOmzIEX6QL4L6ENRlKLGcOFxRrTtS8LlZBbRxQiK
wlLEvvuqKLMuqJ4o3GX7QBaClXBTDH5U2vfiu8sg/RlBqRhgnqsdjhb6aciC
y9mfFI6A6v2vKLhEyG1tLquTRuaLW+grPXz5+LstTw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b6CDBr6yUNamycZkK7dLeju36O4rO/XD+cb8h8vvx+YHYb7GFZ8MOm5TaTjh
1DVhdDw+5aw8FKgSN/wWCuqvRE/wHYSASm3IRPwhwP7ts9wjmNNenHGw5PG7
cu0NSX0sf9T+XWe7jJq4q5kSp6izXVrtlK++rzDSKjLaH19fwkiZKcVoHt7i
hDdRyPet6Yu7ZtzxfnhZmaPyEs64ozWs+XAUDGP+yWKExZ+u+Qkx2b+Io3Qi
atk+4n4zKJLGACjv1f3wTvkW2rsnYcInmKe5mWgCvcol7tizl5H6gbTnrfe7
rgMeQZDSEDDFAd9GLCLlwlApnRih94l3yqHo12q2Ug==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jlt0m0tQP0V5PLxxrLY+f9Nz2XRUgUh5h1MpEfFgE/49amwcn+zkP/T1boZp
hvTgS6qMdA48R9S3mzfIRQmdKz/+w7xN4hl6vV/wODuhwykEzP0qB+BtFbsC
O7RAB8of3SHNBRKVU82bg+Nf59Dxv7fccEiP41A4hpIticikD7zqRdTmDRHp
XSgdAGgSoyNDg+CMWgDmEFv3NN7D+tePexxeoN4b9NcMuhg8T4KQP3j1xldE
k/kQVYGoVfqpZRtchJr32R2Bw4jJPGD0rpdnSPJ6v0jQ/UaQ4AIA1QVFVQuE
stANRwlK7SzsGJSV+jL+c1PV62dFJkoeA6lXKazl8w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jfpy1GzYa8fH3tmmDpLrd9hpozri+TtKz63VZHTDDgM2KhI66nnsm26isvSe
hTv6urDkBjptVUF/eJiOf05UwxYHZ0VTEotSbo9c7iyamhVoV2i9YzCO7Awd
sQ4c/i14HAA9Oqpzh9UyzIEDVRzdl3fEXcPWluk73uJuoCPLZCVMAkrGkWM6
mzH3rZW2ClH4sf+F82yltbjzXIbpaNh/S1vL+1YjQlIT3ntx4+Fnry0YGdix
F0cYbq470WEId55lJ4AEBQdNHYLhejIiG5r4XIoWVtuBYKqHnF40m0Sdfe7M
KDJjMwnXcuLNiHRHIEAE8gRcdOVepyPJ2mcH5AvqPA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LCSxr3VstWPMy0n7vZZk3wyDEz42L7rWa0MUROeTdtcjrsXnNYLGQ2r4/MVr
B6r2uwiwZ5dQRA2f3jHZ28HEOyMtYmMMAYLnpEFGBzX6EGbLKEIvswMRE+bW
Dfgu+vpMIY9Wb60OYc7gRtZ4nh4D1AAIqKFfgHCdayopgfchj/w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mq/G4mJY7I8avB1SpmyGmysJTDVJ3qDvLDCuhpxMaBLrU2l4jlNZi8EIUbmw
rOWgRjk5wK2AFMQUaCJeKQQsIuXyIy69OT73B7/DvNpKOcvHkVvCO4w1KLic
G6XnwMlYmE3wWDzI8FIJWSeLKOw8YQiiikVqNb57Kckoa0R7D8mR+qT5J0pO
Umybh0DVM5fjGFaskkUj4ek3u451Dpuf3YZ1aJe7eqg0kRYSV4Wb+TX48Qdy
2YlMo8hQN2OrouM5U+3c1H05vP9fHL3oRjK0QpsC+OCoyVJIspIQjVcgL5iN
Uv29FSLhd6Do5/qlZTMdbKVA/MkufTfP1t+vUKgluCaodNAaBTGrYF0ab1za
aEJv2O5+l5hgQV+3oVd4JXusosJBQv0mDOhEj9i3WPRxD+tiVc4hQL29S0iV
tCOMgLDyd/JMfwKVXpceQmbHrXmyLoDLZcDiWeVv4PkohQLnDQhaywxY8CDG
IIRDt9X/QTg4aROI0T4NXfz61kcMo0LN


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OOraeGmI3iNt/xUFFSmpjQx8YeqL/ZCTbtYqcEs8GZ2buu+bdWDSKD70KN03
M1bEf1zVO4AdZ8LfQSz8QROh7e03lBgUs3rcM9SyxD72tNiyswBu9ayJU5fy
JuE/D4TiPZz2qNM5FtHSdX1hgTGbAsS112CIJm0pnxxGxBPHXos=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kU8wZ33cVATBdVijevCTWke9vJwmIoLmeCCLe9Th3AHucPTdaDQIo1+g0G0a
S1GS7KEuNxq3HDrxMwaDtY87AiqV7IT6NBvV/hHozPCz3cZ/6gzWU4cVbN9G
3FMgF7VWTqGrUjYBjCXYjvDeGjYTvrFBf6OtEiwrvcULxlAi9jg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2784)
`pragma protect data_block
ea43EoNdx+c7zlyaRUMCEMiSNSYCXr18HuLLQtZifnSU1n2IS9LJ5tGlElQ8
xuDFPkdRWw6HjJdtyDMicLy7wnrF30BW9kjs4Zvyjnq7cRRGKEVQtLfepCeU
t/Xw+iRkt5DVvKh3Nk0I1ZZw/9ScxYAXesBaYzoM5Wel/4u0108BgdVHXNEH
sNcvyb0MJ4vHSCDWq0Ox7MITxmomcS4f3D2y+tmV9x0kBZ1pP+YpZYISiyxs
yP5WbAshCL+60RS21x7sozRhQiWngfhQ/0CGpWTcoYhypkvfXIixnWz8fENM
HS1Jt66Pnb1xD7T+Hg6Jkd7jB5bJzXXvnr9BQBB3JGCnexVw/FCM8gHGpgsD
gz6GqTPrDkTtvbokh8/tJc4a/cz5ZEnKre+H55i1oXtf4ZtiRGGY30F5npsf
aR8Taczyh7T41YGlLz1e1aUj+5K4fpADyHsFZ59oYa6Qb2f3gxe9yda7qPtR
UmxnLcOqS+cnrn/8P4Kq/H815YKnTheDAQc+2RkO6LZoiMT/Nkp1cTSr8OmI
061ou5uTNHlRfkfyMRgKs7+yM4TzNWW0SebYKCzLVjbsgxKLJ+cIlMANo1YW
QIzGPTyMu1f3yB7D1gwdHackEonjgXIqd6TX6gRlcVJuIfhg6p8dkzIZVDFI
OZeMP9c0q7eVLahFdsAQE82luH+uvQuFk8G1Et7T+pSn5278WdDwsspmudkA
ClWU/MpMJGUPODFLZs6fSRz3lsptREq7qc4TqwX4wQSs43Cmm5y3mDxJcv2V
IPOVaKINNZSkB1Wck+MHaaKSjlpsoD9SKRttrWn3N+2FX8DykgJtJ05N2tgw
guRwj74CqYEb25R32w85Pb0a5XN+JzmZlIIjb0Jnwce4o8oJPOtdp3Dnwl7S
85tlDdzZqQ7uSVq8cFQg/DyBftYGqL1v3ZfQGt1T/sQ0MmEfk2hC0GZr72e4
oBIsT14emTAFcXXsztQWJLcjH8IUb9ctQx+mVVOaWjZSfwmROGhb+Uje1Heb
y+Jr4e033IL+258iXqvbh2Au4UvU+VpPM6MOUR/4kdjcbH5eDpqOQAXEtsge
NJ2LdKBYlAuto0ow7ipZb+TgQnMHKf137980EFrnFXZn1Xv2aHEmfHNqgdto
Walp5DRZJ5JjHlUGPabEWtOk+p5NaMWKBcTxIXr02/m+8lvwhf8ETqDKFM5e
lA0RVVyzafhwZqqMhoNnQbOblDx8+mTXGpFzfA0HTTQs5PqMgEmNAzvaqx0d
fHUxtEGHsCD8bOChFqEycq8d3LS4ssKNLt39C2WufjBMMCShCVDDb/pBCBg5
+c2YyQlGollNzsFDmjetGHQBJgOR41LMM8N1CXmI46wwPa+WKqyXubh3TKKU
OxgUl9AhPgtqRVHJGLMj8cpy69kBvvfK5oXC/mw7xl4Pbfm9g5EsWUG311jc
c+3hkxmVphqxPma/zeascpFZEYmBGsLVFUM7R8HoXce89g9e7W8UQJlgvIH+
O8Iw9czqUCRQy2QYQSyuhlBvwzDXPasGv+gJiYvJ7E0ombW4tdhVU29uEAA+
q3wzNBskm0gF9CamJcFTnQkvjVsvjtccMRtJGPaskQ6obPISyS3neA/JyfVK
EG6mLnytkjZu6G+8qNDrCvR0IcCQ0Q3suyYobMS8iqtokAl/6Su9SvKjioDd
q2Kmo715eZxnFEPh4Fcyl2OKahAhUSKXDTJitUZFpg726h1Y5kDfSxR8LUkM
M80sU/w2jsRChNUtVo08kQWYMRJEKGeosPXpWALQV4EKrlBnwV2QN4SQrzjH
XXoifOv4jPSMekTRQpcBT9uqyht76H8QjN6FRYlIzTe8IuGo0kFl4wN63mOZ
jIfesj9x3F5r8I4FgyiWLOQMoY7dHbYBt3WNiiuyL/q9SsH3kwDAOpqP4CEE
vWcdIqQw9b3SScrDZQjxmV/78dP+bQaOPbDCnnvBM70WOpFeHjWfA4YuEqDy
f9xFQ+2qs9Vf3yQ5LzK5BTR/pgO5/01ll5OFrs446ZIaLBPD6O+r6FAaHRmr
0OL4BMsD6OnGqhonognk/TOYA7jcsF7Htn8aX5fpQSfk9X+629etdxADSupE
m9nMgLhd0kN0HEXOJ5mXhLEJCYGcVz6jfZrxPWBASDAqzYSd1/adalyvYMRa
K+osv+0wu4IcKzKTeTSFKLlcyvwwjQHvvfKeQkncoTnRcwWerHmXJbhTrbdQ
69j1u7ufBUSMq7lYU4LsFmjYAgeXt6O8WUimhfQ61OrcgEifx5bV74/1a7n2
Z99vS6S5S8fHwLdDggFbF2dfOIQxHNeZ2NreD4TqWlHuoTS7ctB8F8KX/B/a
n35oyR+5Ya1rSOrcDyHsTQNaDCE0wCxlQ20Efd1ksp2V3IOE/m9KBdFyo0Dj
UdB915KWP3ecfS/FNPsKf1Jgbdf1DcjSscwqp9TEWB1gGjkqohyzk5Iv7mKa
cqKhEWf4VOVfrjtLx13EHrxfo/aBylZ22axUbOd3j5MbwyWAr/7Bamp6F+5+
MjmK3KscScGOywHmgISFsvUz+mECZXKNL85u3SZ8p1w+J2KJgQ6Hbcyb8v5C
x/fuU4BEquj2Dlu39GRbHGm2DaTRxHrZ5iTRMbPWdqCjoRhFyM8+O/bD4cBM
ESQkloBD48EcIzhMLZUuBhlEPktMprlVMlfQX7XpR2EdWrKL1K4pqcNIzJzF
Dhg3ke8rKmvLAqrenjc6YccEUulx3NgijSzB4N9nPwTSMwOQ7FTaiHNldDCu
oHGnBh6TLjwz6WYkNtHZDELfmUHDL1eJfnBvBccx4o3WiRi2q2Bhyw4f3K/4
Gt6SFrZqowo9Ut7o6IW2cWKCxY18oL8Y6aFxw8Z6MrNJS88g/4DlNTZ/tgyM
CBGuWHy+BwfZKCuggLVCn0oc9mF7AS693P3t8pVlvSb2NyAyVw+dW6xkkzCN
y2zQRtb5Oj9zJEuvusCEJEiHX+EgK68XbiSQZUdrgY+Gw0KyTcjTKfAuDwzH
7Rs78MNaMEmSoSM5FekSbM6ZkeTYKRjAMTogS/9/4CD4m3S4heX6A7L01d0G
6GXJg7UbYLhMVawJkgYr45GQD8itBguDWg8mICabUEniPLiudMtgSjAZKyEb
4zEJUyc0U7Yeywo+uTCpW7fH4+ynNsumntfautqzhAY6uFhhgcTeqgwX8jfy
zOpcua65LvyB/fQdx6MMJkAKwJfpt8tu3wvOX08wELZO75jylUqGTxylu93E
tLe/uI/1JpWrYJNZ0hEEqBksYrm5xL5z1l0zf0MGchewQuAS2Zs2yFMyxnj5
KWHvKNIZsxBJpNMl3LOrjDrtTMZ+lBDgCl3khPLT75ukn3yGFRtfwY+XAWf+
Ygcjfhl0tJ+aci3tuMncFuGinzvrfzQvl3C1ovU5iUlTpjDKh0egnG+2zgii
0o33Fz6a6O+qoUXsAbWW7LNF64do9Dt6hfd2D5d+46AbOKDrcF/BxNXYC7DB
r14JlnFWh8OiME7YDBbM6aTuu+CHYs1eWG7wcQE6U8KCTPvXvUkC3q3N8rUh
xaSeIDYihmxd8u+1QYYtk4jykd3AWCEONVAV3o7GarIvldkH+k3+egIA38vn
4NkY1nu1viseFakJcLSixx2Y/0cYmFvN68QQYEyz91tA8OrMegqXE5/LFbmR
ByHYUuJO8riJ9e2inIzVyHXhei+63J8UKQMy75Hq4HN+Xbw1yHeT

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1JLSPc93F4oNjWwCvbm43fFvZ2o16UONvcTZ3NDmduINTDynG5x6FcCkgCSwTVIzHv9EZzguQj/lQUphCMs3TlEnrApd26wy0PcvCuPwfrqo5NCJiP9PznXDIQ5TgK0YTrz4a7MGBdMbw44feZ7xZ9c/GEtxKtkyw6f369S9IOLwfeTjBKu4o6dS3LmGbtTSlZMEOkcfJqAJRrpmJCR3ayrQuQothDIHu/PJWKctdTT8TCUPEuLp0ZVogb/uukPi7PUZvKa6NqHwWLeTtb4qhCejn4ECN0d300icwsgKkXyFGSrkyfqX1xn0LPEpZB3A5tetDnm0hYoK3QGGR+eY8CZTYeZUO6/dOj2EONDkN83aNZ23aSFmSnMhj8vvgwUVgpaWqbXbUF5oa7p6MOdccVtmFJEnf7amT+XDHEc6Ty3C7CyY36p6I5GzAr+wT9PGWqmCqkc6bU2q3OIFudEVHWuwfwKlFjw4Q0cakRiJEBpKlfw9fOyY3HOA5zJvdcU33VhY8PtEi8ideEJ4YQE7vsJ6XjkNtvPUdi9nZ2RZhjmLu7AQEdRDyOlLNIyc3IDKjMEAr+WcCZCHj0f0OvpiKcwOSz05tR49EYyS046hYFw5MrhbxACMRz5r5K+75m3welksQwapMSQk/6rkMy/+BoWZk9P0sytseTR9c0miiqPx1qqyrdeWPTjlNSLf0HaX5m2VyXiDA6M1qroNzPzA57iW9MlYAWxSouW8NBBkoR8KLT0M0JVMsinQ5+pv5//yifwCjvYHdjkkUR0YSM7C8eT"
`endif