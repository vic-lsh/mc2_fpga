// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ggTnV2G6hRG02VxhTxFHoTy91px89rm49efbbJ//oozXZFri2pwyzICmxTir
50pEYTwDiXq+AzwzznrdFAuAH5yqAeLIv6AxoZ33TKXUOL9m3yT9OIViP5l7
geJzT7RDD4YbDQnWtyvYyYg51xzcx2fIwE1EHeqj6bNKv7kbanI+Uc+1zgBl
LvlA3rHdA9OGKuMtVztcM9JeqJma8AFxCt1PW8lO4s52hVIzldLJUMalN4+M
4dzo8SkKBeTFHmG4zX7PEYtM1uBdYv+iUcCcb1Hach5nFnKKps6/bnbRY+ls
29OYBgidPlc4vky9+88XH8FftnFCI66ld5qCia+pBg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kpVMlZlacQECK6BkUbdfbjl+nI3W0FFvJQ+Ijg39r2sbnHAitYoGBrso6ceS
SpW9wtE2sa4C0es58wzuO78cnJ99+UJx2UfRKhvcvSJjxxpvmz1OLy3/n1dU
EHJ7u5T+rjNl59WNIGDPu7kCOSo5XM2W8de6Ndhyi80uvrnB6b3DK9T9y5IS
T2jtFiqkPTatAYw8huT5Y34EBkakKafmP7PAn0DaKoufC2XdehApbGAFHTjS
MIADLLpT05yux3/MbDx+8o9BaHYsZ1U6d1OUuS3VBrc6T6ZHtAMZMUXdz7U5
TdjE3DbxLA49xSDLZ08RizRrTB4JfJ0ldhnMm3WMAQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OaespgdckrZniVcArekGrZn2Kwr7zmxlg7VY8yL0eud4fjyvV81vbvqT01vA
NY0Z9gqyqYJpVtl7I2Te847F+WKQms65OwNaDZcvw5VOP2rcwUqXGCuuG1ue
rz3jfIjq8v95Y6ynLF9xdJeGUgQxXjniCU9ked2xVadI/HT6AXzKegQuqyaV
xMZCyoBN0umOhvhvJyJ4+iVI6qJLdIcxlLCEUM2RY54wpFdptAAyOCwvovSS
XgaFz+bbU7FQSHy0/3pBH9CMyYGCljijm3L7htNDvxJHgVL/m6OgvS6I5t26
jz4xVIfIezq2EtQL6ygKopXs/jONguZ5OcgUTd3VQQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jwypG10GejgKMbjbgB1BBZfwOm9AfPiAKpb2KYAuZd1SuL39HqrkQLnT71mz
fTwxQUTwIgyuUM6cOb9QeAz9GQZlNwON/xBOT+ds4jd4Ok1QLByg0fZPakfa
X3oGrsSvQbCEzCFVbTwFTERMyb/TaTvSG8CvRZMVmsjETZc37QPQ7V/t45fr
jnEfgGdj/UxTNAlm/zsjosT/BOz/pe/kPuBhzCMkxyQR5sS1M1TXt72+jdvi
PygLoOoTUGC4uLJnP8MuQTtfldiTL5m61wq37H+GXEO0sKP/ZJjSJeDNUvus
56/On/4bThE6xmlF1h9vntrFtL94Iax53jmvp2RYNA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lxmMsEnnu86gTGUg0zR5XXZi9W5jw1kSKEYmra0Tl+lEfnx7dSBnY+iv6NiA
BiWfk7kbTAZx9dz9mN56UPnk6xUCUrxFGg0kMogP9QDueTxJnA9FndjTaKfK
QrvOEp2zIhP845i0DNzab/nfyIGMtZZEY+6Own9p/8C6luwQ9Lg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HbA8O0nprQBKEIE0JUkXy4uHPmwkWGzO7H0jBuSBaMi6rn7wLelsOKXCNUfu
esZl/A/btDaNZxkvLPDiyrDDsDZcLoYHxDu62G/QCBraMYVcK+c30obclKfk
LyL1ARunB6lrcepRodmxcG4fqfJhmoTygwcIpPZqZrK2F05E78O+Vzmd1NN2
OVJ2dgSRVn+zRtppwgN1RFUOXYP6TTJEJGMj8LlHnw3G6+gFgRdaDv+hByeB
H/ZUDcRkS/Vhk0owMWXp3WcvPbjRtieDzGGPq/XL1KiYGifp7mTw8Qyf6ypT
HBMAJEu/+8A8Dw2pWmOLYf1PqHjn92Zivp9yG+IYQD9MMbioviZcTf538PkR
s0Tv+z/XdJzigojlQ1TZxKqW0fum5/rDzESu84TvhDizRuxGjwthDgooU+lI
8j0S9Gb8xEttFLbFzmRarDdEEptxG1sRWja5NrVhAO/QeRDM/JNXcHTJJb+y
A+qB/Vcg0BBKykDdTQiEg8PWvcJHzG2u


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
j8ckHfvF5z6cVNgINFfyoQ2UCiYLNaH/L9C+pIl5DQ38CDRSxlIUrUtkD93a
t7eIdrBGWd3Hr4OiPTh7lPpIWaOLDF6jjGp7esnsIfFDbYjDqsfniq5Lm6iL
DMjcO8ufKRbribNvLREn/n4snwn3d660Su/cicBJYEPvT1drsHM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B7EDr1WoP+HU8bn1YrDeqlsoh5UMVh5hc9F9cXlMiqmJthkt3tkti3a9/EiU
805sXtToIBkunYrfPf45AlPSganpJsWEyxppkjnzRXAIemNlmwQ935B+KA/l
5eCxhVmXL/tDtWujXZvE7McGrRa3MjuU8CMaycyMQ4udvbAJFtQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 36048)
`pragma protect data_block
ARRx3EkHkkOzjp2K9LIIZgiKdOnTI4F8oQjBrbS6LP8Z1NdJ8dDNqIHc2/NS
c6PhXc/X7nOJhUFw+xm3dajYlurcwUHNDDr9gOPVEIYPH8jf0Nvq/q+GEPWO
RYDRktdTowHvwJC1+FzmHGfRln0W0c00ZJ2VF5VMFdlTDVnENMhFK9r2sMt6
C9RN3FbAon/9l02X3fUBPGyKUhXiWKhSx+U9mZ6RK8c+jZgSZ+tZDA/LVGds
wwJOIbu1r88W6rL1ePbXr7zBLJ/3AQR7zRxrs3hP+KUmyNqWqRHwWyU6YErN
Y2veLHcppH7bD8OYKfY3sb9MtiZXzrgK7dweajtp80MiMHHzqH8/jbGq1R9l
MIYz/mQR1N1p9Zuwd6NmqV5ih2dQ2x+fcX2iXtFcKOnLk6uwhU5Mi97XcPyY
8t5gSSpY7MxprIoXNNQB56uqUtK2RT86RAcKLt5H0nN4fzfzmxYfBpwAlE0+
+0GE2rFGoL0y54P99H59Yd24qZZxABHqk2Ge/Agr8u02N+eDs5dnNnoBx3TE
S1Tt0mdXSddqBpT0ws260Bel0j+qOICjlB4O2pGgU2kc8CfIphMy+NztnfZh
DsnmyqDHPHbrgwWCELXdRGU7p4KlMO+sNnZx/zGvFjPoytszYFtpB104fz6U
TwKen6gbZo3DRa9tt3oYF++y8kwaHQNbuzkhnsEgw8YE6cm/+5VNyAD0UJfS
fUUJnz8dfY5AfOOEzTn9bxLdCqODi85CQeaCLU0sC+rDockm6GYgQoobb8LF
N3932kif3WN4NEQrYk2OqktavPDShEwGqkSb4jZ3vgvF2E177VAyTmf02Ya7
q7tbVyByxOviR4SU9eZTOsXzOkePqddZpn44BjHHBOXA1LworPrQdUBwYDPo
eqDyfXDXlWGVFEoe6/enyMs0FYxpgSAoVOvclqyatNXyM41bjyrk9z1/cNSW
ZPJutbFKymjVIKLip3Y9iq35tAp3T3mtL4Dn2BVDPEU7RwYJC33433rI6sBO
GlkdOsigvagrrnSw3K0M72YsIKXbSYMq2hashTy5/Hfd3SMIeIQbslD2VQ7n
4LM4/+LqNsQOLnSuiGoTSDicDpAeDczeoqprmmnYqFUsGP/5uSg01KvkcG2y
SI3h4PcY9/q7eI8Pk4IxRsTiOtRXCrc0vBHh0Ym6Fd8fmuenzTklLdYvPBt9
/xc6eTl7dQqxkPWKVh4wEDnDfNm9uacrQNh9MjUsiiAeaLm2Emmfa3IY+eDj
Q4DySK5Uj4zI/BMhC+JixFTjyVC6IFKz09sQE/FiocIbp1chSfJ8iiyjpseS
N1nryB6qabf7YQJGhKNviSc3HfdkhSfrdRsfpfPR/HHhGzIZ/q+b7WHHHPHp
q5ThupGKCoxG/i3vmCrb5SmruMeTiJngRZAiq7y1+5QD9TOZ0Kw/vOn7B9ON
Opdr7+jOVL9f8+DxfOxv2BbvwUmtIE3DOO5L0G/0UoSsuvFKqfKIxKBRduIM
qTHmAhvfjmOzqMspHLP1lcSsEF15xMmlwKjMmazkkjpQx+TZPhq06Ty5B1jj
5UyaDTUF7EMlNcIwvWkWzmlAcNj/xVdWaeg/x8Tl6g86T37PtLDIIZDodIHI
VQN5biGG1zqJzCfCrviC4QcwUtzvbnZKN5bhjGeTV3pqLOa4/o/QlnYJBQtM
01xATKRx6R1gH/CbKm9HVo1+h7RWCET2qnD5x6zRw99tcvNwjn0suk93unyW
FewWkKDJbbbNKEo+tr3xqHUyYSkQh8Ae41LGtKeEv8o3w17fudvrY9qGti/c
q8ZClcpj7aDI/+JDWTtAQyqskZvLJSMaWcrVziKJuVqjAvuampflRRMNUhgb
5WtLQjQU5hCKtpJiS92A2DgWCvWQlylXg+gPpmYV+K9DdnYojiRFZkU/qEwd
cJr8FmTIE3Vh/hsIPfryM7yE7/J3lxeMRsNVgel+974Ha9ipQ5xG0DZEkswI
bAR3jB9nZmyOhaNqvzY1q2OrbD27DYs0uvip0jaP8Xp+z9sDlQ5Eq71skBE9
3wYc/jxyqX/54PDBpePblDCqPEOLES89uftAu99s9Ynod3QqmNi8w/entWA0
2sgxXp9QgpH/YbxsMDjej5r9ZMXA8r3LpiYwboYFb7FAVrRbgUqLTAWZd10/
9SN8TXmuMJ3/Y+hFO4wA0xCpP0BV35/PoZACGO118SQ4+4Q7ErdHZSwLzyqy
MGVu+4AeVBgGcYGifJFy7aYSsqvu3m0pR3qqQ7RkuDCc2v/5NyP+dTTSrcBI
vms40VAwuIiwp4/FzCXIqCrAodCDp1HRCeSP04NcfTJ5H0u5BSYKLm3oR8YK
M95CJjYqhQpmy9ne0iPe3g9kGOZwfLz/WyrDBRpqS/xvj/PbMZwSMQjl85Y1
SSHt59+Hb7nizXABWLCojQfKMBc01f/zuD/v+610V1NVw2mfhpTlKPaEOgjf
yiVe5hzINTAFQk5+1kMRPoY5O23urm8ba9I9gVb46V/7oKdnIZ2t6dem3sg/
g1z/0Vk2Y+APH9TqMy0vd94NZhwFxwNk5GOwMem5UncTSRPGK+dZInN+ilJH
ii8csTmNYh9wOzOEZ3LZ+t4F+Z6NVzI25YyJjnGC8/+CNTBkdVwJ0hM6lSst
YvTHoEbZ2MntJ3ZAuyhAuEqTx3S8U/tzCIy5Cqpo7PooJs9whpL/lBSqjEUi
uPeP2YXazeblBaZp+YfLYoC7o03Uo+wxGVwCvXNlbawAQW6IRcmGXKFv3tA6
D2FFS0G89lvgVpz6nJz46+1CcJuNnYSv2x/RcLWgEcEkt1TipfYHqP9NCKnH
v5i8LWBBFWXIVtu4imJxxPm1SbhNxicMwN4xPI5oEVWNjzkvVsKwZ+/qkIN3
zRavWLZX/RXzjmtzSD2WGp5OUx2jDoUXltAvrazpBnl3UclIczQGOU/5+/+d
3UWuvm1CSDEhSwrbliNXLK6iLT9f+qu51oWNllU6nlBoLcLienM7GoHVUc8i
RIuO21kVShk5571fwolZv9S/ECJd8479EECoZkt1BYJNtAW2JaU3DXmc0TwA
IokHeT7eKryb9QQI+rgd7cWLTBj6Bz48WjMKxKf+bcdS2s5AGzcsPkxuhpim
MyLewB5rborh4+7QTRTvddUrIM0pBmiApdxASLJjDb0Ix2+M5Lrw4Ydw1FzM
FZGoAWzLxs4Dk+k/sGbyqwXybBK74TYw06/Oi8AOP/EH53OVxwtwSmPSl4N2
ykIMV+Qai3+8XdE3WMDQsdUfwD6+t1B1uYUQN5ZY3fSG0dsrCoE/ZL7g9yMb
nZdNU9mk5dIrDv0dvbU8NpKlzVv+JFta0DoCpNqsW/Y0FtHtZNqRAVBpFMP3
YiAzm6bVrPJI3Ohcaq9a22PIzAXe4BRyodbeJFdYpjvLRVOKN1ZKPSkyW9ra
hiXHlOaDRLEkBhmKcRezVMx8OFgXSbNqXi4Ck52BAVO6AVe5gtJcCcfUFXZ1
5EUgn3H76WlSwonEDsGCyZVdDs7BKqfBE0esxaUTMKgCAkLJ+UVsffFIMHu6
zkGFRAhK+u77APiS1BBOE+3efj4Zr3cN9OPKE8ZHhgzwN3+7Bhrir1ZtBYYZ
qvhYU9VlLxHCxHBBNKCbnitMrz7eLF4tUe/KxeijV7vxNaxL3zrAy/aBiET8
UHRWb5T3W017nLQbbO+kL4AN64vFEiKcGE06rcH4umU1PuxUbRRLcOHo0Twt
O7JLicZeBs2+NpRJctcx8TjgAYJQT9feWcGWz4/KDdXKfOhwUAi3d2EHlbL9
HorZHFM7PkYWzoJ0eKm91xst6zMIMkr+i8l82MCZi3XQwUMpXjGcH4aMvi4B
J8nFAJfOlG/0Nr9I8JtoiPTGxGExSJfdEdTi0TCbAsRwWAnE/WwE//b8WK/m
x9QHaaT9IC2Vmm4CoziWYfzYPSmiuZWZyjplhCttsQnlPBkdxyBk/b1fXrTa
6sgyj4W54naIOOxUi2kUoOSLWFiNngjMl3ea7POv8iCMhi9dki2oQzaYktzJ
KLhra/cU0427NzHOjWSmRx1wyr/qtrkqK99byi2tIJcKCPv6x+qJXA1XpRSU
H9XRXQklsx5IcTkouGFGTBdoz3GZszqfbITgT99AKMTneKmlJqUZlD4JLQLO
lUqzQYVDLP9FpsDGhCFyUXs/BnzNbP0yq4SH3aHxT3xSAi74PPbaNcKxwTje
uEQAcPd1X0irmx6UG8ip93AxUV8hWnqKVuI+hxSwvZZfBtYRVgoe4lp7GH9R
c51wXM5KrbtBZ36tothy/btHv2LuF8HW5l4ebdw3Jy5C3OdMfwo5rncZ3/XU
P4ejdMs6gHWv1Z8JqbrdUxytCURHZPiLasNZjbuUFdMMs9hpU2Z51I5+IENG
kNg8Iry81oKd2b4p8bXKu+JEqHElyvUXZALXxXtfDYKRZwvPXexthZvz0UQ5
kiuv23HhpGpbkBiuuAh8bIB2EU6cLVLAV5ZhkaeKH/zqQb63NisolJwEiOaX
STLMDBJQ1fzXd4yotdQqJZRJpncRnpht8rGeiPdlK3a1GvjaeRKuMkPBnmZ/
3TMwpKiEkMdMzV/NIRmgiIOe5SwHDHonipjExzL4XEW8YJDoaSJ5gEK1TK0a
Yt6nQMtUMmyemm+MCei9e39QT9fFCNmgOfVC5eGm3LKijccS4SFIeGqle0mn
Xj1j+AdW9ZC/QFJsv3G/9ca7e8ht1sbJrF4UduLbrpEkvsiR2SnlavGKcCwM
DH56a7CzSpy45mZ0DAFjZwUgD7Y+OpmM+nm6pLnXxHG1K2QW6VoSpAZCe17O
x7ZgBDgnU79GjxKUc8ontM75vLu+yaMc+j5g9aU1XJc/GIlIvp7/X8PIhcKr
4gz5ZrPu4w7jAevQNt2nNNZUDi13+X05NSxHsYZWt0Dz64bW643dixmksIv9
dQUipK72DiE2u2Nd2GNufGBfQSvuVwc4XwfTlYtMR53+/nw2Ue7fZNUumRTi
DN/bx2o6jPPHJoJmMFBKIkHoQkqxQHBEs5KaSz+qD7X48yEW9im++ZVSEpDx
ttbC+465TtHWVhN8xYk/CWf9cUyubtXpJ54aMBQtu0G+W2i7Sl7+jHxLKGMB
deRi61DsV8cDUO/tS+BZbLdmoTOgf7WI0n8OjHrfb7/VtJqbd/Np/foGfOVE
mXdPM0uWkhF7r4qHw2YJCh6IIYAvfrepE7Zk6W9MTLS2hhSaw+F8uAAu/O3O
XGTwIHXeSjalUirxveMy6OGPqQTpSP+12wjgnwgRmCMx1O/FP695Q9bza6CK
OCyWkbKeskjRc7EMwmK9ppXRen/6A7e01zsOuy8BgUtee/uXSJfMDBvC8edM
11NBseaHwCoW04+kbZGivPnYY+o46lxWoFDqkROSKtidUDN2jdUAce6X+MOf
hxbu5ZkTNvahlo+1Or5NOeCUMf1v8o/ctqxZW8NhzNmEh8GZZNatB93Aitue
X+UyX2inz1NJp0mBk2UnKh0VgE4+Bbj3g9uekD5CrPHAJpBMqC8puRHfAsnQ
3xyh82WQaIYinpC80dSoVXlL/vpNhfGKZeU6syonlO1nPETRXEcNu48h8F0N
M3VXgarYG+Hleup82PsuE28lyWxlTbeZqakd2zWAM+i2rWZBI0fF8QEils8b
sdP2IJT8bOrbciYzYQK1kISxuPSJK4+0no3qW8YMdWW9qKC7tAhIIi++Hsn1
o3zrXIYMZO/i1qeMaDjBiA+r6OG89ozfYldx0FjyVcOUH2tSXrzdz6LepvZD
zk/NfOo6h3rjzC1ZisYxZ0QGhTu+OxxOiCM7tNulMivRJRuaDwGMRH+vE0Ur
/2s5fxJIfKAeunwXEyZFLRafZCMLEyUly724MExcb4TDr4uZiM/N3OzIYsqJ
R/1RotfpQDc5o8xbFy3WOPE1AsaweG+YDcLttQr0/ahzLTEXENB8UiQlzodC
LVfpopho3SnamFqc+uvSgWvqTyLtPAuZqTyKBrdQNC1VZu2Kmj7nHj1KpKOD
yz/rk9wwPXjaf2oBT5E35GUf5DSs2gmUJOLQIMZ7BHJl6NuOJ7YzWf1f4WOM
GnXk2EYqvdK5X7QzLWvahSz3tYZ9A1tkZidzkLAxerP4mwjGj3r+54wFqKmM
XgWkGcbnmUKwyWONRdL5cbnS2m0f0P6r1EwN0xkKpxUDFD6VkiZOxClvMsdE
5/a8b088NkOTxucl2TrGQlYsJnhhNRSJ2pgx9/WnpTp5D/I2UR2QGYUlBiTx
boT8Gsa9U+c0WgQO1DaS5/Lw3JGVlqj93TZKXj9XJQs4tVpzM+n4sG+tfbyn
fX3gcTm80c+Oh1qDQaQw13tcz5mQWIWz88iKQ+H93J+n5mH1VEFIDpFMLN1s
zPCnQir4j4HVjxkaoQkhMEzJ/MOul3Hzh25B1VMe0SOtOX2NllD9Th4hqNoH
5zeSxwv1FP78xsGOmw2OxM3w4ep+5++OjXcueWamMIIi8YopPaplG1ebpTg+
DD2V3yqSETR3Ra2ZxUWu+FcrZkcruuq0bLxqRIJmauUbGcRcjodxp37W4VWP
VLwez75qxb9gNhYUuSiPryALiwxM5sZrJEhBHdRezJ4X0rzHC614+z+fvnw6
SkrI5ze7obtEU4NFicOZOjXBSbJww78Nee3zAtt2j3rgJUThNJIkUVtx5yW7
SavavJBreIC0hLKE4UUVQk1DQzudj5IEfe6cLhYM0UKYsugm7vhBOsqxEYsz
+eFZgD6vd3Ff9rSliUCwbJ2mAmFM7N28Gxo+1BDqkPkSVGZp+vusL/uK3VC8
uouLVoSPh2NHcD6Yd7o9K8u5vcO/2MwZhDgckNI7/LSPCyeanFOYTGkTk5QF
u5ZETaDc6QWYgSIQ380Al6xzWTxUrnUfw+X2UQ21aQ0jVW9TP3KE1ZuIcGC8
zfciavoEFxSVVR/tpZcep9hpJvxpykt+8XFQCouVlfM5FUCQE+7iuOBAtuEu
4nWLRzLnKcOV2JM6lUWNR/9LTXm9pk/YmyxEC0kMkMAfcfOpsvKkRU8+Zn35
txQQFraLj4NINi8Seue1Sug2oX/j6IusPAI5tBrDX6yvcOznBmj8g6+t9KuB
u0YHNSYhEzvhETPtyuSRIwib1++htIssBKo0CiyuRqsunE/eR34euXKS39V0
q37zV/7wOeKCBHjOc3oYDZ5ndv0E1dQuVia+lKniRENcV+b5ESKZb6xwTbjo
akodnWNzDrqKLt+nnZ44rrI3q7QpNc6tWan9W/BbgRNLV2yeYVMsgkb5P32U
SC6q3hGyxF45l4sGMhz20RkIxaltd8zoaefMS2CxM68ekYGyM6wf2WUfA1lZ
LmK9uW+QSoOcD9ICLSlqDTmRFHdno38432sC1nm3SjgZBoO2FYgoRpzz0uH0
+BVLJ7SnT3l00eAI7z9RLyTwSCvTP3kGPQhdBQzmzP/yuXIplN0zCwj6xU74
du/QH4DRyq2CTp38kY4dd/cWvMOD9REZW56wHywkpqHxTNCF4BxoY+glVuKa
e4/2NK22uQHbpz/4hZXA6luYYayLNqaiKyI/cwGD8w65cixHuV3Yr1gox6jp
oKESB5FXqPxM+uqv+1Q1NnkD2V1yz456PBtilTuFs/q8JCchX998Vdj2qTQO
GOGSUNLeNFOtAAwdaPguWmnEsnVmQ54xMGHFBFk2n5lPo1oNMtMxxQZ2FUxc
TSUkW0hXcUlPkOXZP6t43w5aVC7dyc/wjyU3n8U9mpjvCyJhF0sq2pWFQyov
wU7YmX0/Qb/fFhQzSQIkSBVef9pcl4vugoGH9abRB0IexH9Hx6lXZEzHDEjV
EjphSgu0PChCsVdplMQraJ2jrEKoX6hcG9Py8N3t4jv1m+TPXCYy27ydthjk
FMWsTgKw9dLyBoNEa8Zo5ViJ5AiiqCm7nCGRZZsaji4At7tsAz2xWHL5tZif
w1EE9y+pYyymPouQuGRHRFOdokQfhOBYl3XrcNmArBhmmsoG+dTVT1dV7bz5
Qgd/ekEC51Z+ONSKe/Rp8KdCyuttW4lcF8KHYIYXBhgXr8lLWxJGnhMkyzhU
rG6fj4Mi5drus1eSJY+PbWsj1hllJqDCRQQzfIjz0R2ECyHobC79HCKmGUwR
vE/nwdSPoCuQWBEU7MWeG8JIvV+DdxrCXXn/CLNXpWmMlQbaf6hlDOo2kXA9
UErI7+ZcW9WnZAYXutCtUA5L6UBfqlMkJKonYNCyYwfKp29zmwoCNewplSO6
HzqZc3vKF/n8+urJUBYq/qv63Pc6/6XLnfQK1OWJMsVbgvonqbAeDBi0BfDP
ilk+2saJT7cefb6T9v4aAuhmwK3vql2qnbVHLIThZWYE0o8W17TwTZMiA1WH
qmSBJ18ru8S8hHUkCMBj4uqcWKGKe3KqCQWSgr/bhTMXmHUAH6KF4nDdAYeU
j09ABgIA9PNttoS4TxSCtLoTqdafjWDvyQF2XP3+Jo8DTtf0QVjcZg+rM8I0
p/qoQeKAhiYz5Qb2o9XFIPLPPFgMdwgfRfC64QQuU1LUUzXpijia6twkdP9b
L713jWz5GaVqKwDJW/jTYiv13VhCQADXZvM0pIvYWIPlNT0h5ShMMulBKLUn
1Jie21ngyFNVR2WDK78HPGmcs8Fp/zG908SVgS/ZOJx06aaHvvdJarLEqXkp
Ts8pmVoT+AxEYUayH2oL43Nin9Awneo8TkO/7hXpd+GiUYiza2WzBfTIX3lq
vfvyvDiiLX3R0FQTNZvJBX7+i8tylOnX4NxhG49NSfJQ5n9/kclWc5MEQaSc
GlrhY19Nt73ZqeGtfxza6DZR/CnyHEkabzRgp1u2v0hVgtgo8P2F/6dhmcN8
lKKZgle8DLqyGFeWsR2rarr55S+skJTuAb9G3nTmHXgb5yp2QdBMXQX5lS9b
nq+0Ozd+Dyd9sDcDv3CBTM7gt+KQsnJtnyHiXmFRBJIfov1wkHcQ7NT1y+qm
DgY1nXbEArGy8o4XoImrT4E06vgQOiElqjNLdS6Rw1hTUUcVEdpNwrWXwBYD
wDHH1jocLlzKZ+e/MpycGc7J5Cd5v1qzqpCV5h6+/+I5AtxQkmp++kG80JNQ
FttVbQskGl9AwaLHeiYT92Il95MuhyRzP6cZ2nJjxvBvhpDmkgykFJnqCryt
YZ+7iBiEmzhEgcmYZ0xz/dO10epvLPu8Sypk+JN6om3o8g5GV2C2TS81Xb3o
FYRELxob2ykuR1eOvO3uZEdyCOYo3qS1cNEZVh3fBKhiK7psTHjYIHJnfVZI
fVwMNRe3TbqhWjNe6isVmNL9NeAJc7tQJgHidK2zphLS2shGZKOEX+Ro+x8S
COWr7V3huoQ7vJNADUwSGCbbCaI7/41fVDze40KV63CcSHQc7ycZrJmv7Ach
t6g0gv09++8Ym6GMQNWQmMo3G+xinJjhh2RETMjlPhn9oKMkpf5qvg/3FxIm
UudOKrhoZthDtUf2/iFNA/tlDyMXhGOBOecpQ6b6X4eptYl2XjQ1uozBny1j
fSLc8th/ejSFMPwYIbvj8jgNybfUo1B/KcLnlcescLwM/T0OT2ZVlljA5MWC
z1pYDHe8LSi8qkMTc3A1jXWsnAGRC85Hu5GYGoRfZ6y2X9BqbT9t3Gptls2E
sXv5McHwkBz+6/+9UCAwQAN0ucn4tNHtNG4FO0UzSa5y1GCU9BAEtyRDQebn
OZVEf1+zfA3Bn0iC/KG5TLrP9ieQe2Y6wOxr9a7ubu7RLOYhTDvoVF03wlqy
bea+i1yFQSQxKftY6+ZvZjQuZxg+XPSQ0Ndbg0EXqcpNisRN6zQGKVk8ZFU0
bQ8QPWjTej91DXH2ULjjtFBDlfHvBIRt8UdaJMVUTLmqS/Ex2vANJpu0eglB
as8zIVWQp9wJ6sztT65sutHpgBkfXH81eRTQ2cT/wFMJJ0iJJuRkbxUIhBqj
OLQuAXtXn/2Y8aYLdTJg8Na/etfo4LGQucTrPCWMgsZnsmeq6rOqLxl3BypS
nRKabM6d8mPzL0SUDq6b1I/nJTqvhTb4k2K4CKsP89cKSnWuAhfmXY/ZtbNT
6GoUUIyl0s0/RFRAlVxhgSOs+Wk9ZErmySGogDgQ+uqIsY6MpfDL6WXYiKjx
RNmRI4SfqxvLQ7VCJh8MY5IVbkJ8t3xbNvzdV165SOuYohCeGjz5DiTFkbZD
y49H07gBSzcWfWQW6TnLYwWZezDcTtfbmyRgToP+ptArz68mQ9GJNfI0kThF
wuLcLGFzq+y2k5gRjkrKZ+pQZ3n1+CaVSJ2hSd6n2dfnAnlrI6RiK7xJTl0q
ZQE+mbnUVn3t1skC8v9zfq37s09cKeEecKQoQ+Y3mAi+BfnT9Rc73kUOe3Iv
6kK05jyTBgYYga0jyTZ7cqHZuqMNii5GuNa0MJXEIKgtrM2yJkJlzCiM2yag
fOopx4RDsninfUixH1tByyk33bF/cM7xNgRAS6Ai7htw7Pko55VazSB5YqDI
panV6bRl/qfj7gihbbj76sPZtZZP+Su7LAo72ZfQDJjfmGeC4raooKGsmPQD
5qO9Q8yaGnICdkER0nQTSMyKoB0jb7kW+LjNlr/NgFUW3BS9fGX9u/OTItz4
axQ6033YI088LSY9dXqxH5kff6q66RJUhptr2T4y92JI0AhBLxdk16jWXU+A
/wUldSYsgku9V70r8Ob9HMert8fkWp5DiubUZ5+Fs2MCYGTMzhhjMnFKRb81
sLI8mJ1ZTVaUKpQCfuw6+NVxrg4PsA2ibDsI+8qynZPL5C6cvjTyhcfBFVPt
sQbUeH8Lbb4vNteoEj9Wt9VdNoXQ8q4EgBrsgWgRUsiMKCeXOr9ASqtEeS+m
XPKaHWCQ7gDdMAD6OXlNC/dG+p6wsjUsQtWN+8rSVUQOI3joe+Z30yY51XEM
CMJnn+QJqd586HZfmeSJWPOeEDpMFXeNS2CysouMaSrozgBt/1FBn7VUJAMu
VzE/L+rTyorr8TuQlmVQc1F8jcUflcdKxhMULr8g9jfoE4YSdMf6oGbwz+Gq
rqXl7M73/oJDes7AXvZcUthWl5LX98NDjRctV9fFDEZJH5CBzDPy0sy+is/Q
7jSl96ucpQwItZqLRYj9A1mATjlms5Zk0iN/WVjvaAMNeoydHdu9roUlMM3q
DiWmd2iBKY2z3/woB4aPx+E7PnpE4zFBgl1eoWWPOe2AgyfNsfm9SIxAz75V
UgP/tRgOPtGiEGgZxmcTi4j5KyqDgqJ5xE4j36vFobJ1iO+VCpr4UXhxmtkZ
kUbf2cJ4UbhWsW1/aveC8WJG9yA3gIreRYQ24uY1pN1JFk0bDGxJKvG/Wff0
OjSAakH78iyo1mRTfoc7aq1I955NGJqPkkQl6Cs13sasRztubikkFzwY0DSk
g/tjqhlhwlotrJwxd4FUM1ofPotpphwSy/9YT2Ap4bGDcn642Xo+es+WqHMy
8oQEfGF+uI3IlD4hpkCZPd0lVmjU+UHHylDxMN8ZdFltwjWOMriYSxG+j/7Z
DdEdOk5GobrcXI9Q1LLsRhTj3j1dklsFygJpSAkBlmHFXCZang6DF2oQfZTC
zrOYZUeUxfzpO8n6VkCGqJM2xx9p8QIIewLb8rY23PmSi+5vMu7wOTyLuppX
Jj0RI/pqJCBEG2XZmept0osG9XAAWEErQi54guFZ8Nek6W8icGVJuB3QUu0B
og4HO3eKHzd2ZaQ3EFfKNeIoqqk7QmJfwR/UT+MLBzfMYz+P2ONioER1lIRq
zI8KVhog/VUXqQOUf26uzywVOFMM2+YZujHwP/cg4LAMu/tgjhZN3tv0Ns4c
vOHekufHARvHIo9TgCW6995Bc3hMyJAP/zrku8ud0NEDJ9OwLLdDIwx1OcRt
3deLjc300sFoHrBCdvjx9tjfn545trEC8//rn7HBFLAt/VpHlD8kXtX3qWlm
hTJP4waZIXHcXHcRWbAi/g3oLqLpZKAjak7KSBXAqlHUlOmbEUUEKTdhSJCa
4tdLGpcZLep0fzsmvgZdYbdZWlg8ZNUIrhRf1dVTDzHENnPz0XDuG1dUzGfV
wNPMui0HWUwevUPzhQyGNPcoxQ+aGYvP1wyGAjtQilFoOxwdF0lpIkkqKrO+
aKCXI40vmqA0eLJcrjTq3WSCy751yiOSDGAImOthyw5PmZORJBy0f+WNG/Vz
Yly1YN0nvdZzl1q9FqnD1QmyCKPoeTHCRD/H+vyu6ajIKdJamYYbB2MPHYah
HcNCXz235Afdg+Po8hmJrFYmis6N9YHN/T2CQI0MQziBjElsSBdS2NGGD/RN
oMyb61DNiTYJfPm4SSW/pqlIymlzYlF39DxxOv272DDwuvkDNvjEZNMPWpPC
wbF2m38ECz6AaY/jag3lgUn+JUCR1K1/6Yr5BnSZdNfccFjUR4SPWFgDi92Y
ilK83DtINJd3icJXq++KPUbXGypt5jJXbZ4dHQra/bSOiF0DfK2OS/Z8K+wD
aFzwVN2ZlIp8zOpKGYKwVAvt8yBJAJT/cPEOa3RIJe/Zczo2PIT5kp0o7RlE
VEOp5G6tO7MGlSJ7ChBSKW6zkTn+8grK/0ApWveAf59FDGmFg7Zq7kV6B+bt
T3eEM1Gm5jesfqDkBywqn7gXCSg/tzwVWfiUvt14TEY8PdxIg+PgpGP55Mmu
l883aB73KdedgbkE+YzKPj+Km8InSxV5ky6rnNuswtKDaUQPjJzKugs7t4eQ
dcu503GRMyXIdIxFWIImLqRlossFnM7Nfl6i9X8DVu5DRUsloTbzfZccIaxb
LXSrR5weT8niyUoNbU4XaoITK5Zp4sdo2uzh6Gh2OqWiJaS/GNU8Bbmy4fnt
iEpG+vQCy0oZXw1K5MzJCe/Cu+ojlQDtSIb3kOxc75g+eCYVPkmglo+0vFXB
qrEixxyDvfOK2XWPBeMGJvxbuRQetAHWFcWShl4Ox2dcp7/AlxN//ZNSFcli
38E67NQvUfSS6CBs7YHRxXxa+qqa518MgRAhnG86TZSPYTssnS+GglWH28vp
B876JSD78tvHoqMsmkpr+GaJ2bnXAMOFGLzzcc73GylrnotyJ0Jy9HcraZnC
ww1zsskXVHtxyMT7tTneMbSHHIetLDiTuLAt/B7MD/BRYvAWDaeMi/Hmvk0L
nGmBMRfIOnO9tPwDvL+qCZRI1a4JKq6SVwp68GzJQYozQgPUs99arLFwGZpS
Zlnq754dXIKNaPLukA+e1NUalIQUdSw0HmUhF8M4Err7cx7ncTdMSoA4D2Qb
x+3MoiwGHf67R3f7kmCSp2tEH/ykymWHJ8YCO58z0W0IpyagFRqEvjbOiAqp
GlHQ96AgElX01BMx+1cPE/YL7z+TUxGy/1qF95rRXA7BfwDv316tf/uLcEuO
qhAl8ScrXWm4sdC/HXKy9KQdXtMapvekz5uDkeN9elSDF/lYkDkMKrweUBwN
yParjQ6jYdDA08UjN2aYpmSGM05ay11+b7kwmHlJ8xMgod5kmlD0aZ/WZvFw
//34i8/1kyAzH1/kgxKfJ07ArpY5YzkTiAYCS2zyIaYCwH+HPtioXxJmZuPq
3N6rgkZHHzAu1I+sWncdv2KWL8weu7A+GJcXaRRF0xnnZeoEa1RafpYiuqZr
rwA4CyGAz0oaJd5RkxVDtTBAQnIkj7DclTwOd6ZF5fU52bqba7GE452VtpAJ
hS7TBCEpRbyvz6M7Ikg9EXVsm65Ldfev06yv+96gVCBXbiDabQJ9XRkPyPJj
sEW3BJOqvpyh02MW6aPml1AOs5gRfov5ev/Ypc2Y0Jw16HNfgLexFsHVjtut
j9g6SL7mpXxwvd/KhkVTQzZTUJtx0pDIgookEvO1hrYLhi8sk6zwB4882ZYX
FAJq93Csq+GH2AzwgeeLL12F0H6MFtnDvFJbbc044CbSSWbl4WtbLDrApyVl
NQ/yLgpomIGp9zPx8ZrCwFzK0TJvo4KcnHZNierkiMslkhCSnEJ33W6z/83M
177YVNk47xw22iDbcp/i02lAFDMb7qJhhfu0uUdY1Hkq7w4vXNkeNdHlKd/V
+044Vxnh5oUktQFEYkmHNYjkd9Nx6UAdaGLmrCzCPkMQ5zmLqZbU9Ddhv1Jl
tzS6Tfgk91LGhEr1fVneMhOsg+v+mwYikd2YAVmAa0Lydve7E1HY2k4f4mb3
xcEfTdk7g6VeFEKe/o9it3rwMDYA2mMu5XKehi5sqtBrRGO3Tnz+1+mMuo7C
Ph841zaSflxK55gX5cQCSH4s1YOpLmC93+3NUkKuBEaCD3FkR/lhK7dv/KOu
QhbLb+DwcadntqbTnoZzX9TZcnKaS0H/exHgX6gmTGPsmwowsADZ8zfgEl6N
TsmZG5T/3a+ESrQHyRDz1LD3hqCViU/qQJ8ZVIy2bFoYXOl5xaPaSI2WPRFE
XkEAMPL8wTI1/iYKyxyz8WEDiVXsHkgWCg8jxJmoaLYWT3QA8/bI1nibj1VJ
VIqlZEGGmT483OUhwMrOeTZGX/jscLwryfgRrrNVswyHFRxoiuELD1HtQnz3
i4G1bcH8XBOa1lJRGtTUR33kW1g7PxrAwE+KVZv22U9/hbbGNeqiG0SohAOo
itBufh/Zg2srv0ctH09CsnFYsKxYSFqb9L/tEEnPphQw227vT/GOo+AUlBy3
ZjnuOQJNsvBVFBiPBQ71FcjDbq7bZ5BYHfI0uZONprT0Zky1Aq3AdkOK21XD
ABe7a50Mx9J11FJyC8684119xVK+IXdOSzncl2UE1K46YYgHATVAuzLhsgWR
dfmlgI9UjrpO+8egr9bbzisjNadnFQR1NoeikBQSFnXVtWxCgelSpTqEMbSk
8Nakkpcmp650AMbpE4h7DOliG9Z20tLcpYAGlhsbnRK98wq1q4Kp/UeH9Hj3
KYRiKPoStZVQVvP77nSUZEtRcBUNtQqARFP8t39RNSnbpuZ6+tB5zD2WOSG+
1QzcfFLmGNsxerBfczuFcumBOBz8dX07Rv8ruYCev6yz944R1CsHwh4Yatda
uW4JqKDjUTR8ocUVgCbo7uFaiL7ZFyeE73zpr1S4WHdtPkiWRjBY6sxr6bdY
e1X7iP/4QtUFJYCTM8bzxgZO30VlaabB78P+iv69SbA6OlEk4DviFO6i2L0h
hgwPsV3qZ7ruV54OWqXrhoea5KPnkKeArbD+74aA9Rzkkfbd91r4+YFq9W5g
ZyVmgbFfKt9c/o2zliQZ5tYsAnLSUrYo33gQiAx3DqAnABoTeH5ghTdIzt1e
7TrFLCpPwkfOlvZyAsGvHTPAlgmeG7iBlW5yDmpmMJpifwfaiOOvI9gIVxlH
2fY0a5LBrMbSg6WeGZm88cmT34Khbr2+YjKOU5EtwTzMxqv9M1JFT4Zpep4w
kZrDh0fOlyZJ55e7JphbmwmE5567/BfEQecY0qaocyKqAmpVc9WIB3u+UjCm
z1g/PsoBNEpD/d7SX1KPCptJcNUIuqSwi440MR1pO6mJL7OAKmBovvRpfYQR
FS8XxzuDumTb/kOB65fdqnTO2PK7vnPb1fEN0p3Oe0zlkbQgPJX/QA00U09p
QODvSw6BXVMuvl2pzO6xF6A1qlah+QVMMPyAgg5cdojpNUKPP+8HEWr8zDoT
dS9PjpnZa1Rcj5cQArSwDSdz+yv4YAbA9j03cSKCcoWb/3jAckGxEmoTd2Lk
Gs4c9hagINbjtqmrP6vY73qKULtsZnbOQwH7w8rP48XzXeJLS8ALSqtbA7KD
Dm7vEMyebWJdX3/pBNEeIRqxrNMt8G1qIbmfFzJL2cKMaJIM1M6KSVvSSljg
GsTXUUY5WuKrAty5ZzC61yHV5qHCp654QEqNOt6/YDbovNjxQBDJRr8oKaXL
i17O2swdey6WPcNSBMF8Lmo2lNc9Wuicd+aZKzWP4ugTyTkKUwqQm4YrDB+m
JALbLzkJumvCVqiftuyBePAXV6+2vNp9i7DUpd2a2HnsG0fIIPsXJSyw8Trs
R2xPg3BII7f/ZtADRPd0AMtD5SzMAIwAT+AvuFjj93B3NLWdKTukz6EOJFHu
/kHSSZ3/MgZ+gxaT6hp3baFAqizttHfZluQTp7p8e9fIqbOj4C39f7mVvmsL
iLDaXoJnY0UT+gQnOsCjKvGsMHnwBa4BJ0u3RWGlH62k5RH2gLIVgHL9S+Bc
YU7fbM/UYkQBDFOrnF5xreUG89owxARjVjxL/CbtombXWXIAvnYA7YcZOxTJ
htV34xn/tFbLqAHJzbSTzn4+dHQMWqdKBr7BbVbXzMtK95hBgXnFmAOOwSNc
3SxyQ1d62WsdRyTt7NuqbuGnrd6nIg8FCEWx2LUVXCgYPZJNfs4koUas++w1
7+uXJ2Ya8JglOr1+OvoIofAYF5cQNptmAb1TAvj8dQLzgU8c0Hh6R7XP3tLc
lt7gp/g/NuIixv3NQZkYems9OnFbP/0Y22dVPhnebjg9tmxWxwcDmeGW07GY
//EsgrMUF4KO4cypiENgPKvro0ePqj1Sw0d1YLRlhQaYotc6VQLtACBsz5K5
7rlv1m462stJ0kjTDS6yHJNMNkG5M1nKdHj3DWAATWwuz1bQaM04z7xtNQEW
1+rJket/jQ6LrEOki75TierEsdnfWkigVzANBedrJ1uj1+8iW2UW+4PQ1RP6
FD4mQ4oKGbFVDL+ryCssnAUi+EN+evbHzzOz2cTpRMhY12FfuhHgxSnyuCwE
kKM2bSM0hvYQe5EIyim5IGq6NzDe+ETqy5TjMKpbLY3ryYwXAY0AsnYb0rYq
8lhU/WoHDGdS+3xEDxlby3y8WWqVcXhGTUVw5mbQ2Ay6STkqcLF8AHxT9kF8
0ZDE2PIT0iM9SagIWxI//ctRJPrSg1u+v7bQ6fIQNbDOpTrBDM6Q3dxXt4Qb
VFzD9TWxGadtm8omB5XsgpWwRBQXlNTXyw+tReS5uK5nfSqT6TKuAGaNzrrg
p6BfyRnqLyjtjV71nFrq2+TpJL60U0wEPp2aB11p/+bXE1JgObHNd+BcV6pm
6A/DFlH6u5V3F7lZs2jmWsWp4baet8ejel+opqG/TrPKiuDTBzuf/bH8MYFi
aJkh50UyO8VgK38WFGGcTtk3kTbwv6RDCeN6UfXvn938g3R0bPiUvA+HczKZ
HzQNGnPy9uAwBXTeIgSTyQ9A5YcM69E6jWrKVQWLuznV/g2gk+piIbbTOcVT
V1QibnrKX2vVWDJaWZyFvJYl711bsqrobPdGrGjxhWMDP792lot1gKydP53p
5Dy9Y2KARgUljDOV9O9Iiqu4NXAFQAnDFHwxTqy7mVlDt0QwbIHVyapTVZai
5fYyV1tcR26qRG9WYZ+qMhMi+BE5oA3ZXWwi/rQnbu8O4reZ+AQ03dw3DyUv
7q5y/9dB9V7gnLGeTvG6UrZHSc2qTBTRgUMO7do2liqBANV1fmC2V4m19U3x
CT2KfSzCBFQbBsySWUDc8y6HViZQ+4cVvh9IniiXWreHCNg5uQZRS2Mno0Ws
Iez/+QIqK2yJtgx/RPY82EHdL0aY+PofnqlGHDKD2hmWbwnYpifeq2tpG4B/
L953arF4/2DP6HtDnkTdATZqXM0ZfIEDa+AUckt6CoL5rEUhCSvHMdnTT4fb
rUhiiswrXnb3g/GI/1DUkzgOtx5nyxeKcbZgA74FyCkAyqrubAMt11/13BFY
wafusnyTNtmo/2Z1KhXpRbnHaffqRd8Yf0Bl418ff6PeUWnVc2JsUUTryQ7M
piI7GX7jHeXFmZ2h90oMTvh/uIgwNsd5Gmbl+Vp62RVOi7dls91SvMhoGW2P
eMyf26yOCoqSkf/zbG9t3D/349qhhXiPAwPIYQmWGj7nNW+FTjcJjpopqbg5
YI49+j4o5k792wwFu2GrHw59RHjfJaLgy30+nL/E5vDeX3YgdIfhXnJr/Rwr
k1BKSa6GST8YmceASt1/THwFJ/pGgghLMJhtwmtUk9Tf3iWTAu+cTgtUA8Qp
BBii/i8QNpt7DZLO7aRDKEVAc4y+4fmb6zELNplWj+UeegAuuUFPsVnqcfJ4
XXzOp7V+v5JEJ/fYK/rSEIX7XadyaAU9ncAe+6Yw7Ul/YWtrDymhAttt6GK7
9LrHpePOwVbPZcBjrXzGlkPD+dvCghhrFfavqLicE272eWBIoH6Elhdwkf92
+GUGNIBfoALMaDjIcIB8L6D/muP8ICTJQmL7nloeJeY5KRWZRk2vPABMACDD
Q4s8mHo1/BHqTkYKWFbH+mTp5dfCvSFlgl72bpZ/WyMTnzKCCql0nIcsndvb
S2I8FJPyJoYNGZvwmK3nD8BFern55K4Lla9LuWkm6W6BIdFfVnIncklpygqc
eEB0uOvdUFEgAwyxzfNis6ey6tWc/li4SHZc5/kdzNwCmHEYXVeZhNmMK6CC
aq70/CjOYi+kuPiRUguRrwyb3dOgDT1uiZ/GY6Sx2j1un9UQEPoU8s/wx8yw
UHNkmVlNka9rkwQzl7Dwciu3trjJP8SIRs0P1a5yW2I70/4nw69s8ki/yEvd
ERCn5+HYvH5MgFy11S0wQ9ZqLVLiqkCc6oby7SualC4T0ihEag6Y3N33eqyV
e9KksjH8/wH+RZ0R0fKUt1jptEqiUeLGeAAi+VsJcZxPjy47Ur3OpRWC4k0i
1eAKSIfyKoO+ckZBjZ9PQaXCxM7FiMT9ZveX1KY3K12MILBD6MH6fuK5h3pu
CWrB8dQ4SDJj3VLL7VorFCrIgoxfm434xUnSnlZC90vO8WNdiMmS4DUECyYN
xsMvmdTpoZzkSWFg1dGjRfYR+o07yhMqPkq3hY1pN6RHLL0UrPSgbtD9zJeu
Oh0Zm/NoTFMsIuVRoGbM7ztJ5zcbyy2Z47Xb88gk0116+da5IIYTvjuNWDgz
sSESE6Sg6ZDqpcHWfojI0l96N4jLEOJ5D3TSV6UVVlu0xpIk2qO+P4lJwAKQ
R1e2Dtme5O4Z6doQSmz7qd0yKEOaPksK4pGdHJbOT7ffOTb9NqrCa9PYNWRh
vN/jZ46T+RWkP8CGstHWmUkHXPK+oj/i00NHSaZgDC9f/lQ1pAvTzq1HsJsq
DXwwMD23/Zjzuy08pn9hZfFuyTylzSV+9YTV0LYrSD2B7psR+pY4WfSCZFbe
yyRjwSerWq+aB1OlJFwL1i09PR16J+4tqmAp6BhXIopc5XJa/FJCgoRi4PpU
LKbXsqiNcll8LPUWhzVepne6Hwd6c9q6NkafyvxfPTUij/FuLX6K20TQDCWd
WtvjrqUSmFg1XUQiIqebFmahOmAPuOVBQ8+wtjNAvRNXB59Pys2Wd32/Os8I
zjm5l3dXR/keJR6bWqu6qwZeW9sOjXi8DOryK7mQ/bdS4ffA6LuR4nPsXmUZ
27axfPMWC6w4vNJSP5nN8UsTXCKGrYPturgoyGE1AkWSksyul7pwVctGocie
ZHd0hCMSqLttP/Pa0tFIWXgHOXkl4svvwYvg8whpTzRqjV6QowoH7+7EIfLh
FF7sBZYlGg2AIm9+oGdSPb9ChOmxtCkMtM35HgFeGZscvNIWw5kOCFeyh9BS
Bu9eOjugZcKHdKsVb0/c8lvWf/E1Qfq5t68ykVqHvq9rnWMZDZ7ds7/y934y
kCzZhHP5dY0Yr7m5qZVSm04XtNRosNkyCE+bCTfvE4WpWHXJ/Q2VOeSMKXSQ
Zvu38tAxKbdl+4H06oewAGbvpqRBmkyST0JyyHz0wyrWNx9VpijtDgrOz1Da
VAX5/x2TPQTMvNKo/AdJpxM71HfN5xBnHPj5XZQ55DfYs8HjBFiBHe9sbWrU
CXydDuk9G9ZnDim57uFXZoZxzzvI7nPRq4Ca7/slCE1woIFWa5u3VNlN9xF0
CXt67CmrMCNf8cZkxqdKhH7d0cw9xZ3tpIdoSqg6EmDRKxUTaritKwvKXhzV
ACOg4KX7nfShsYxRa13FiClqInvrSplxRMzsqWjRYXbRGorntAMb9aQPHTrv
6048QAQPez8jSUMTpegNzswMDTDzdnwpsr6xzgITOTAwDcgP23y10frQaqbl
ICmmrkwZZMnTJ1IwKvzD//BVGhbk09w4sblI2Kyyjqdd3Ldlp7Sc8a8FuJRf
KgEniRSt2klZbJQB99dGHHkPBJtkKda1ttdJ0+EvwuldykjBPQmX8D/XXZri
RBLA50qXWXQiWkkq4gfobVnMKdyIeN5Cs+JdOoW5pbms97eJobBgupT7FDY0
n9M1WSmqjcam/f/mR2+D9vdsqSyGNIXGuz2I2MAQN3VKXWgJ4CwEjkyDjJDr
jWmwJ6cyuuym8eXTqNg5SQzQw5SzftGatbS4rSKsmuDjPQqPdMlPsvCD+LdV
KMzHvugJ9/d9Y1z+rr3GPxNjWjB9dHvRCjB+K1QsaZ2IO+8acUwRLQlzeVg5
us9guUad0L2wiOaehZm5auP0Jg4a08bN/j4t8oPXCirzny2xZS/5hBYuEpXJ
XdhJGIRk5XvFCqvx7hzTa7ML4gOOfSehFC9P55iJD+kpWJaQSV646r0i82x7
Xe4E29zm+6bl4neIiEoGyXkN1jrq48AEsJO7huxvBO4UmjQLVxSjbN4NMFpq
yxi3MCA6w0+rcq6a2jB0nUt/qk+L38dQcyLu8LOWsbC5F0+aO0vH4LTMY1SU
gW1nOYJdEFPRpzaQq6zy8OREzTrr15/+8fRIwjoYmyP8P3+TVestZxPoFsf7
T1woSDwJVWcMsyQx2SE8OME1vH2leCLkC7mHlNr8xJ0PdWi4OFDnvs+LTt2u
HlkrW2bVB2bY1rD+84KaAircegfm9rX3p7tvgYfHMMZSQT3WiM+d6R4Z1W+8
L8Ho0otR3+t5qj6gEpkVaT9OPTJdcBpy7P4kQNMenFcgMRPMjR22Vhjb65nN
FDR7HzEKD5983iyIICr7pjUCv4hdGmrgsDdKidHjZuX8+W4yk7HUlDpmdUyk
inVq7wWNT9aPEFr64I5/cnd7zT15JqHvXZFLnWoOZIfAXmCdngSZ4gtobUch
URtbxn1SO5YQGKMDCzcGOsfe6RuseO62JaWwL5X1aH8ImGicRod0AsnShOLJ
4AKN7YTgZkjmLNON3lXCEtZo5F9c/+xbJk3DfUkD4+sO1Rzbt0077DqTNHd1
++/jA0OcsWyuIsbyBzv24jRetehF4ZGoJmSwMHvM46ogmlFd60PjZhiF5Afb
wu13WNv/4H3oxZKLBDmfbI2efX9cuR/ePdWkWE5qohb+xzFoUlEoHH6bnjoT
0FzapT4LR980pQshkwDqM0dYSSJlZClpG91KnRcN/auTkpK2vS6kVdBHTOdt
2AWPyDIGKvvAFyintsxIyzu6aUzqweuDjvFQiEnjA7Xg+aYo9mpnWPiNwRkr
qbh2wraMtraB6sjSMAIkUWSqDBN5zo2QQXExJze8m2b4lyqjsBZOT5TITcOB
43pgf0J84UM88vI3BrmvjAUzLkKqvVqFCIesq/5ruQrmukq/c9Smd5iBsUPp
a7TZiLb7U89e1DVh+8fPoUEmoq+7cBsrpOM0O7WW0fU7/fzfSdXm4Bcsvqah
m/WoHmfMuSLO3Hcfe+8erkxQxrkoyMOglvdamGCe2OP+fEn7wHwoNWbzRzJH
brAWVs1Wzn51Q56NnkzDxOlW4lW93a2kXEJRvOXHsYrigRiZgxSzQhINmv9z
zheZQVee/LZ7w6SX2p6F+ufNtZxpxoQ2I5SyB9rVKsq5/xOnLLRTBLd11FK0
7+NFYWYUQYNWUkf/dH3mos74eJuVRvuQHctRqmuEK4vBKlZLMV+OS/+f1Q6+
y+A7D46hbo9YSd5WTvdgrSGOpG7mxWFtsdUFNwM3NdjFHZiSCXH3BwQeOvjI
hLlCQn/S31p0JhI36prdmKPv3ejLc/5o5QXHMhDH5Fz266RhQEIZlRyoMI0j
XixnTP3ly+DwWygSHkle+GOfo6HZksaeuErZBM7uZMGfyD55jRmsequXViEl
11PneJCDuonWZJ2M6Uk7NGMEF2v+Gnuj83R7s256Qqrr8y0jbr/fxRD6p2wc
42PMBKM0JgrcmYcdWez3xno/HPZ25KFwkq87jXz/zohfjfIRHW0F6FnZwQLO
KMYcsPaHXZL+1xP7nBSD74b6NfH3U/m9Lt79FuUe1ndxq8r8mkgZo8XtweCm
IV3uJbY3OAjlEshNSdVh+/ezIpIxUGi1v2LMX56LM1TT2Pib5DvjTc+GdNeH
7oXzmhFUuHJ0YHjxrZrJjUSURIMcuk2cDTVZg7NX9wJHgfEsTEzwGBaXCHh7
qZf9Jy8j8+52QgQ9FzGyt/uiUyi86PaNB6o1bwgOtIVZ9bgm6BAQZ2rooYTv
JLkOnfkSYCbj7+CvFyVfY/mTHInD1kaZ8uciHRp8ZPYXqtu4UiAVb2DebyYs
N9M7U+2fX/zEXcr/UeS4Z3r02SuziL9zVYn2Fuf1xu1tjKCkPO4UsB4sBLGw
4sexlduD0jshD6dF/LNApLv8tUyneHZYKQ1u72GmQ10tdK+MbCsw/kxD9G2v
wdiJULf11EYjmrr8DhNJ5NtYC3mIWyL+qzXh+hIYPvhJMy3defXsduiPAsr3
np329IVze5fPNi86AYrRNeqE9M52BLVba85gEo1rOjBLVOEzQBj5bafOPAkI
dWRe3/gBN80gqMDKBVgDo21neNuV+nP9a6DP5H8/w8v1CaNZOOkS+5R3CrhB
Scz9YlyBCVfSic317BCTxZKCVP3iahhIPlxcAMaNCyonE4B2O87QJyYZZ4SU
GPL44Cy2oFJlIaXNcdF2D3vl4jzxpeSmOy5t3smlaJFhsY3xUPDaBpodZwsP
NIOMNzqdT8G3RbIT6iNcgHBvG+R/y4odaBHRcLMuwI0xNYwnSb33LEk2OTuh
mzNzThzitqt02qRFjUXfW4ibvhX4tWKVj9klaJJQEYckLJamAHBlVanMNAJO
6QJ5xG99XZWNWqVuEDgr3ukY3ZaHO0zYep9xZ5ZBV4b8Rr7gvZIoWeMvS570
A/sLQq7V1/0kU1mvRmFFUz3/9rjKB2wu4IqZJgKvSDBG7CrkSANgsYvWo+2h
aL0JxrJPo0F0yn5DPR58bCSO3YJU7dPQnIrEfEULNotRSrtaC4XkijMKC2z8
Dp62258/OH0H1NFX2/5CjViyK8rHaLdc97KPWkdapBNA9FTdS++SDYiXpTAa
k/jlX6LNalvMrPMOhivTvYKwIZKgfuGP4bApc2O3zBaYuLPAaJZm2Gl0qEX/
Ub4SqoT3clcS+KU6QNWyiuEZ08FQ5mlfk9CK+a+1med+pwZWmqvSYYhz86dl
S12g4DFyM8OjiSeL6HwY49f3FY5pnukCRBWFvlLX3u0fA4+/8BxcdB6xkxfo
I+hpTLPhsYV2mf7FvZwJRjf1/5lt9uVKb2E0sKWNVM5eNajH/kgj6GRDLKoW
Pw02g715t184Q/+1cOj/3OXwxWdZ19Bv8YgQqBzU8gKPno6SYxAAR4JKFPZu
CwSEJnddNVLQw1vLF92fxxZhRJIVIAtLhz5PJCc6cGoB9GZ4oTmMXyebNCe0
UaXADFTknb5P5hyiwSjdjFdOVMZ8Nvz5RpsxjXLyWxNk1RPSoBGMe0KEqbOw
pbi/+OJfARdoWnhAvrC/NPBs48wQJpg77qaV/VnU+jVQhKX/MQYpcgyrn8fA
MNyihO78fFCYivQaHqXI4pC97X37Z9yzI1uCnCqjkKhNZYQgp48RYBFMVRtP
2+lNbIZvkdyY5euOetd5l+Q4nfe1fI5M+ZMclpLfLFvqQSHXndzeJVhx7Qq2
NaBittc+7TYi0nMt8KIznUBh6Zzxf9AR/Pw5f84/Lovc8qTtmUPIFaYatjWO
hbAuFpFqZugWwpFfOEuaukS2KZBAuKLIU5AqRQjX7Djos4RSMgOu3OVkanI7
N+N1nk9VyCJktf9Xpfu6gdLf89i9J43wfLfgZ1DhhCRt1Ue3KRM7V4z69EHI
0zaGHrJmkgy6pYSlhchUHthZW6fMmtlrH2YWtWt9HGEU2gF6iStl/GojUcJZ
pMsuEXCYGWkOky9MhtEN+sTN9394UXoVYf66cXa2G0TztwRCTy4uq0XH50V6
hyDnlfaW6HNk4cqRHTuXSPri6xYw7LGVBDKZ6nMz1dh7OE6wAnDSxyXKdnFi
tOCX7SKyvp59Ma7EJIe6Y9B0gu3Sk5jbGFzM3akAp2gvX6hnwhfieeLbO1hZ
RG5Hem9deVH6PYgxmiQK0asZRTYqvyY1GO2fYH0rMe9JsRU4pxiLSZw/kz2B
vlTfOQHkltEsqJNVVwugrdh/+XoxAqwhInO8x/vpSFlYVjKhP+3iCROG0QVp
eY1skOAKLsWs/jXZ37svkQotYbFSWzzWa9G0pIsEdLFgFBoiDZTlNmIiFJbv
SQvVFCEM4dvuuGyXqsguz2rtDut1mW9uXJG7HnxVazW1nFpftiJ/n3RZnShY
Q6PwxjXiZz5OWjXz57Rf1qIiXqy/+69UqWrJ2GVvxE6ThNVneLTyFi8aL5/x
CTspEOBISm86ovXjEdFxdTzYVoaiFq6Wwbzu03ouRcG1HfwNz9kCUlGGDiEt
ogQsJZ0tVAh5gVXc/t7j4DVtaTjdeT4t2UmA8/IbK4Ado00l9ka/EhvShRvM
qfCqtWKqqwXMONcIQE4CYTE7twRJ4IqHCcHzYk3Vt9Zu1QwsOTm4hzj9p49w
IZoPIjyX+y9hWO7ZK8WU8yCUl8mjwi8kAS/hf8RMUFZEJehLoNmZpXja258x
N6e4ja675671JLzdUowFDSz8yeTknsW+yHeNAtMhKri0xqeN7tMhxUvwnjkp
SjBmqs/sVUtGQ4vprLgIksWxKhfJg3ZGW42U7kQZg7PDBmp0fEfoH1SU/ZS5
+qalSyZBuKOyRqonGrXViYYLvkd9c9KGbL6cGmxkVQvXQYGJRc8iIBlngg5u
T0G06obAylIwAN4GTh7nC50hCATL+mdvAjVGMqDYgoX7ggKPKtduemHhpROr
Xjx2d2LMRCEovr9ION2d8IUba5WFb44rjfPCW8964HTGcmK27GM6m/waH8HU
J06qYORJFoJ+RLZ1VvYJT2n87XcAMm6GTDrfnQwuqfcEtROoPszqOg9Ksfhv
eDeYjLgdplvjT1lN2RnjMCN5UfPUEsuFURY30ZLd+LNn708xY6JtwIR5qpEZ
4i7OJtq3GxDZ/gjYZ8IfHAfNN0auGfzSEBiycngUaq9f6Y99E9w3ZnVmoTq8
11Wxj+OUMjE4AKsVckNljOOggM31p4Dd4oUDIbnRJvYu2ovWfPYmR8qPgTW6
gZywCVl+RckzGUMvk8rf+XMVgowdOpeLEbtJv753utXTjPswHCS7z07Xwy5E
kSr22ANTodWpW97nMvGD79M/36LoXKSqOV7Ku8wqxVffAsWX5kiixTBlPwkt
A6NPo/hQpDUwZ6a7f57AmtzFRvWmNODa638PjkrvlNFeNfslKtDkmVDyHcMw
m2rhYUY7ey4nOaefrOl96HHpYyjpOVKKQ8mJ+LnjVqw976NEr0dBLT28yJJU
UERWQbd6a35gQ/ywS4MwGQeJl5dfj1VzfyLDq7cYGYWck597PWJINHbsrbX5
wjncczXBiiGoInOCzASMjmQxyhT0k6Fh+FPv9LwL/SgDZ4Av1LI7eaAR08Al
aOtc/NbgYSKppucxZ44aWYmEoRTdepVSI7vQEFFFgNOwjz8MzQv7pbXvYtrY
m8TfEphO4tCzw6XDy8EVXexCbFAXz130iXWPLGDdpIyi4j3NglokDBNxzONf
Ei2k0HbpiqRZ03qS7fmIxqo2QNaDbZk0QbiYU5g684zXztLLGKuNoe02jACR
BQw63+XBLo6oPW3u6eaBqQJVEw6nnW3hiicZBoz8od4L6767dGSKfnATzlRG
J4OfcslOCkColR5yiiewv0SyjoD/SY+U5dgyKiQ3afIquAz3kND3AsZhrJ2A
OkUvyn3PsaM6LHTgXccfVwAv2EFnuh0xt5+r8zmWqidGb1CnFaUgbB60hewT
iBXPxnPIKQOpqMnyxqsUFKiXhNVVuq/WV1KKRVthvvrwmp9KtTTj48/UhshL
9GeK/K5phTx1Fz6vQFWrwhRZTPWe28VlU27YZWQIffQtF7qk8ru4V9dhI4xl
WdhItW/rIDr6JahvY37OxxwkGNm4l66PDeTE+1bNbKFdQTOCJsFc2l3NWvBw
i4xCmmXq6nRmd0jK1q7P3TtWTDCPZHCBEGdM9igNfh0h7BuaSp1NUgHCyiOx
HiwIqlAtKXf94K/iQ2dPgvQmi5H7ujzHA5Rda2EnYWK3P28J9iph7S1BV1T4
YzhrmZUGdlyehvBso6yZ+GKzJPPlBbElLtMp4L/5bPvCdibB3pYYkNMegXyk
KhuqYxCOcXAoKCoIMFC4nUk9aEf2y8uxgybEwVBpoG6eFkL4T5u84HYQ5TGE
4VwHlD323IOQujoiVDZFd+PL22oCoGUV9f10Xc8fpJM/4p3uLYqsfKeZgO3+
HtAAYrTjSaWh+IKcd5UrOSP1ohOmbEdSn+Wum3fSMIZWkB7A9it00rfZQzuO
oPUlbGxrgPOrvE6XXekPbQ5FtIuoxrvNWE1oTMSq57Y8v/GVYMlOaRauOtF3
OStXR5+miQKJ0wxas5yrjIKhLVHTcjWB/N3xb0MTxan681+bUOwwUQviUbcT
/toqkOAkwiaTzP32NObmmwq9RNy8RIcKjL6s42hG5T60AZA+v95rXkk2NKUZ
s6g1NxKLHbh0TxewIZfVddhFb5QMFYvvfjtyJRUGJqwaLGOw+thOX4eTuqPA
zH3p9a5rmSNFJB2be0uwG/cE/FrhRr/T0p1QvJCZqtQ5Ja/PRkLhaGk+8fm8
6StsSLxmXY1GRADMO3MGL1QhMLlc8vMZfiSb0rzQsy0X4T6UYuFFWlVEa9oe
um1EqQi53TX2iPtFtBpDpIt/R2Ep4EEjJpP8lQ1mOqScG3sgH+OuckK7NiND
7lKDVrPDo8GS3ktV7h15xRxESOG8hZ04z3iA9c8eALJlwckQitAGvQoFE71J
fPovxqktYBnSHo9jV8FRVTTivVj6HhMSP5C93v09qBTDMebmJe7hNx2BkgQ+
pt/NrKMQdAHhznPC4qvYMfl7zktipx4Wz15W56PNAvk5/RzpkhNLrVvjrws/
/TDDnfzvETGIt3VNajipx/7/31GW9I+limFDjqe4TOTS28TZ/mWtGvP+WGkF
xADSr4DhJFt+bjRIMUgT/qIO+20ceRIN0oCFdJTQKwJuTSCxOlv7HH40PK4v
vtSZv0XyXsWdJA7Eosvgvwl1Tc64vjK4huYQr6m8FWQh72YeEU/+Al3xJLWC
rrMpSDuvVatDY1fvUsvOKJMTuPP+qHMxM7MWYg2F3vx3ELpimZ3r7pU78rFx
xM2zARgBx7Tz63RwtzuHTKJYWrSHcVtAh0MRC+/An/IPbVFCN6x5VECvGW6q
qYvGBthTGNjjit7hiB3LBQtC6X/C0ivojOP7owQk0aXbsOdZzts2vPyI8KQM
WCdt6ieDbj21GJeHYxuU12DjFWy69xeml9oDr3vN9Z5CSls975p3XxIP8I+K
j+46mXV5R8hzC0cwUsdHWiin+VKYHuZRGZj4st1vOGQVbIa8vBedQ1QvvHuw
85uX019OL3jaDmsrkrHGtecoV7rk28u1vTDsmtAWWQ4iWj6VH/LwQsNiyMzE
cKZxqUoOItctruZHzjw0x8YTrwNkFOgIwIfsaQOI95AL26ik07dg5l4d5ENe
XHZLK/GxSjPmcNHcifkosQJPhkUJ7orzJXquU25L5g0Iuz4ex2xe7sgHutrr
J6SVF2qvk0lagBlAZyLHQxh8XRdjOuvHy8z61tDRvWigFAYgFOUAJ+zT3KUE
KfsrEXaNuGK/eUURRqFLeXElug5Ei11eY5mix3WmYzVUS0cIHlC7vKKj8qq6
k7Y9LgIw6LAjX6wzR3X6BuZyuwbhfiHoJ3eP/iVEkUAwM7WuqxtniDYGgsPQ
teX1sc4zSxGG0MhQ5xMV6o1C7SnV2YdwVBqyLub8AoF2exYbglJ8CWwe6o2f
qv05ghjbESUo1dR7kWGY7AYPh8V7aJBm2l51CHC9PBWg/urFS0GTEcTCKXWq
l4tv0OPQ/Cg7PmOwyba/ckAkMoZeniyorj9KnZoee07JJ1Pwtnl4ageVsPNL
0lzyt/f2i/D88GkuNCIoGiGa61peuUdtQWDeZmkfb/R2nvYrHCAH+kNE10qJ
lRKmuphI9ItF760V/mXOvpz+scRb66kWulJystrDefEZ03BAy0YwYrcQ+Ouz
LxLzBbmRW+FD5UDES6Y8YhDgp/2OersI2szH2CdDsa8DjJgNY/dFtlRKIrsm
FaSws+ECsmn3mQwc22LcLlJqbUHFVVDelmxOYELI4u+4jlKS1/n739ve5XWR
JG0rcqVURhEk6qIcqoN2e7rWHIwIoE0wz0vSMTQEsHwNKnuldoFrPo9aLRKT
F1VXqZ86l5JGCRjDq/iZw4p/YUivQdC3MP1hpqcV5OAietSBqRvyQywkyQMx
CS/wYnHZuRVvs02usnK2pVYPDGUBIqDcqJETORx3REkT5bLhJ+4FNKdDcOXw
EU1Vr7/66mQP6mqg+dw4oHOZPROqbWRLRerCQtfW3Ktf95Yr8ueKZyy5OL2t
f2cu7L/NlOD80kLm9ydGLtVtIJtRt96NTCuksCpcxgW1fXBTF930dg7ZswHr
9UMdZWNJ57bB6wY7XqPOra39yzSgd3NBjOJfPXR4WBHSKVlFhYSOgmiQ007j
IN+0gueNkD30YHkxfSpGvxRNzo91HJOLWD8/2hEG38ZPC/7COUa+kZ49/nHy
XGc34CQgUAmM0w7zu0CnTnD6WVyRugWZe+8dsWp3hCAsK4JXcOWKA4xwjBCn
OuDlKgusUwuY5rlIpEgyxdCYQEgGYhwKi0Ta3KQAYciZMRvbRpcfh2T7gmvt
MhQ8tUdWmgUYJvyxKRtA2i/ug8oxZNJK9672YN9teBmn+Y9bnVqq+zWJhLvV
vlZ8qdzO7TzUc6pxdYFfgVKt+7IK7O34cTbP74Xd9nyrImRUeUNsRaf+IRwO
iSyboM3NkzbbRg8JOwAoYL7LCR337ftLpBPLmAYAEjM2ouRYwrGhW8Dr/BNX
K40m0KvUWcjxoxkU7O7bsFgrXAHF0BkH45a0PN+iQKpcrAtHHRfiYhV+dJDi
eMt4z6RTZ6ki9VUhPsugwpFBl/FkxGRE8bXOa+4DNBryGq7K9msZV/fGQVFs
HuczIyFa3skXKul3qWOcVNkfpCHJkW++kMg5HcF3xfwTL8A10/21AKWxdWI+
rwqEQUoejoqSv3vKCiaORZzsfefC+xNXcusWEYAgyvMe1Rtw/s/Ot6T3zzQq
bCvGxnlfNowTncpaMe7qQBnrS9nh8ZV3WUWViLraxMRwdpc3DcouYsi5KNvg
C0/uLue2IAificxzIpZ5iA+TxWJ3jTZ4M2/VdjfV9gFnaKTjvw/RlkJXRXCJ
sq6Vm/nKd4A8ALddy2HAhDxck2hw9dY3+2kY7QFAzDIzbroJ2l/PXqfBDt1B
7nnuc999Wnslqz8c3jbvPr0+g5YiesryFK9aJvxKIqJH4qzoqJqMZPHt4iqm
e0oIUoqElA4vjC1vLPIOtejP9704CIet1YSjG4NpgMnIM/tR8OT44paYjESN
t4GJu9GkWSC3D8X/lhH3Y5eRkpHhiExsWNTB/r3OpZCws8n0jMqkC8XGfogT
SRw2jojymfVQybQwybyDYrELn6nUpKCwQ+7ih8shZTuXZ3DpNLPk+UkL1F3z
VHJ951cgcJAL8qqR7mGnWk0mW96bCk8FXC5oV8tiHLIXki0gao8LpCVUXtsK
IZZgagpOLc8Fkl/CThHV/09e/uqNXM1ogYTUiy9diCZ9gGpsq+knHLy9+3yn
Is4XD1aCCPc4cankk/7O1nzyoC/wDd3uxvXmu0Bib5z7DpfZ2aRf041g/S2a
9ZojJ2qCpsvp3+T9d/+jOhvuM45krvWQeIAzvJwriEsY9CLu0ulnhUsZGIwQ
qX1pRfAXcFllS8FbJePbRBKDy+FwVAkyQHfk5K6v5SzwdDqedKNMprd3n/y+
csIdRHyqHLyLWZqnp5dHOpTnrrac9yh0C4El2B0ed9sszc6khZqIPqP7Sl0D
Ptmraelcs55EM03zjdhY2MHLS4jHiZDmIbYKp0VduT5TSuVbFqp2GyCuZsVi
jIFruldvso7Lh/kB4eaJIZn29HN2TZ+NXtWEXkceUkShZL5UvkmgR51axeVj
ETC/4q3PDaTvYIL9zp3nmMaukqZow+ywp0ApbZf3cSawq8X9IbeP+wiDt/Ll
CXqhD7y5feCbRDnamc/WE6eSw95xL0sp65ZpQ3vmT2zP0g/aEQ/tOetM1Thi
+QExH4eCYSOdSBIDABt9clJnzhUwq5WnT61ESBiXCtRHZ5rWx5oE0zS1lV2j
ed7EBgLAL3OPuX+EUNc/R9nGUSJpFIV5ZN27284sGmWR+ZVZg3JG28a8Vcsx
IkDDKaRQn0+9nQVAh8Ngp/PdvVVO6tj1EAxYllmtfeEUasnd428kC84/2p5q
0OYbPcewfdWo3Gvz/jxSL4LXHIvd5Rj7m2vxdIDwrCNKorY1ePIprCi/V1g3
gkLGRLf4TiEMAU19ko6tG6lkg0VP/lzrrQQ18Vq2PlzbxmDI6km8R4k0p8ot
ip8lxcx1nfgNnzpZaUaRHy4mbQR0UcRZ26FFEvFP0hFfdJ/kQKCXwkRHrjk5
jK389Lwj3rSSyBt1cVxwx/MTgtFIBbRMEEkXSv8oU6Vfwe9C7Ex91boRh8Ra
JzWQP6eswiEWvQTO0ZIhmLgcXAqZpBcb2ls6uc/jh8vSLR5XBsy7bHUuohbb
GNTwwYQyasSiaerEX6ynDyNRs5X8QncRxgKBohZJsF5WTKh5WN2W0PCyKdBb
tm0jR1Qx6sr9W0C9LSaXKcra+Nw49KkK6A8om4Ao0Cup8rcDgYx6x9F0GYAD
kjm94Uux2JvnFYEFAhDCiMbzvNOXWKL0HtxCU2/kCmRwBwIDM5aVmhLaBAtr
tM6ui6JboIECgOByORLC/tJfiWJUau1/Etk+eAUWMfYLCyAeZFQzyuWsN1PV
K3MnPiJ4CkggfsCpJTRppNJWcIA1JPPOm/d7G1L1qp9bP1XQ0fZ0XxxfEPmm
c1tpc5kLZgzCiC1NjGffrutOekatpK3cfsCK8LLpg+MN9I/W24LofgFe+qEt
a/FuY0ZduCrQw1DM5mCSNT/TNbEkbWpCe7W8GGai/vhVWjDuBp+xuO3Y1F4U
NozxP3WocS9PmOGwt8USW9yegm1vCYxIuSejdOR1lT3b5U5UuTQJBAGTVs1y
0UmCFpsYL535cd3AbY2LC2NTnlB8COViEYiTANkW9gMbIDGe21t9AikgiWAi
35m9/4iwrJ+A7U+HtN2/TWyfJHNhbLoeX2TcWnN6bwI9Dh8kLB9iJikM9bo2
Vr9DyhkOPB2LUY1SJydB35RF/JbIpftqG4+8ncgYyxBe2w5+C7oF4Gb6ACVS
WOWQ83VhiRNiywLc13sqhseKcTQqrbJPbFDzM4xlrf32rqGWBCggqWMIRWUp
0HecHU6rZmn09E6jOajGQM0q1VaBfgIeUxDugN66RVG7xV08lCfXLLiBFSzk
QMQMMJIILUrVXkUHI6oxw7eEidiJURPFzSf6De5NeA8cVxsKKxH/b5Ztfpe4
Hk8cMUzUI1hEHBzeGIfayQobITs7/rKnX/ymI5qONgvDEOBdZnofb5EquLGT
TaBW1lVXVjMBUPMtpgVHcbLQ6YTMB0UW80gr3bOSoOIwyTojsmvMaC8TeVOp
0Tw6hkMH5IYf3BV49X5VAgIPc1XhOrc2Z+fcL+/g7ij0B4DhUn7CYBW5dIMN
EblOJ2oLkg0t/KS5KDxNEqT7IM1VWej+SzfSVlV/AMQhHXVW3Qk1dyrRQH9g
X71Prj7tWFiaJFEg0GN3/nVMyywpdqCUV79JPtX1Hd6vMc9Vf9lIcBNYS25h
uiPSVB6Qne3+ja5BM9jOciVwcB7NR/TdCYOKte8tGV3y30QK5Fe+K2mCQzOm
5CPWzwLqlWDM1jrdlrwskOI4zG9KL9n0OzOBRJJ5zz4WLN4A7tCSWOb/JbF0
sQImhcPINBWFKVghoN+Vin+KURk1K/mjgxCvSmFabY4LNWU1i6tEPt1dOfnb
gxMi9KK0LpWcAdHFmo8190T0CEoQUFbVocbLaCvtoEj0Fmr/AZMfslnE4aIb
fx9MXdDxwtQzSPZziI7CkByrluLVMo4PuvvlwsmJl3na8j6RLjWtZRDqmT8K
x5HYpkz2hIfn6Ecd2LVNn210C1OuHlDkvE+HvZu0sMzjZCpul66u4FFPoo25
A1gFqiYu+tIJ3dcrUEoQvTxLFyL7JyNWc8W/3Nkx9pDM7AfGk5+IgmPrqfja
jqy2gVp1/1alPf6yh+X769G47tm+Jf4eSVHUKNevLBrkGygq+YsBXDBdmkaV
yBENG8wlblJ7yoqtTiTSp77osyTm7+hbC25fmxR1MLOEglDlutjt6qZuDil1
6j0FjJqfk9DSg3ODefZ9Bx8GsTc81l2g9gViHhEEnF8xJZk6oPMRwB8RNYr0
ImYRcMGOabmqMc0jR5eAwdrdJq+DIP4i/JD/PzAuiEvZKhrsMOF7YSH37h8H
AsRN7ZzFiW0INkYAOfwhg9WUr52yc1b/lozlIXMnPTmY8z6AGf4xyWgEbNRR
nId2xy0eddPY/8mbeDEjPHfTtcJ9oOx5ucosgh+C6cVlG7KXzeMUxLfIk6DL
G+TpYmhX0oDha3RXgwg1bmY+M9uCIxJuMJyK/s2LRivLIRRucrLNDemcP/lU
BhK0U1ch5tw42+rSw1Z32gGC2ujeJMBZp3uRB+jmwrpS3oA2jobGDgK/qVCa
z6a/uTREFss9FtH0Y0sxhMSNKTFQ4F9zDKwVH0Sfs/P6EtZahVfmpbajRUOO
y1dQzpiZhukK7LcFoxhaJuQpWU2dZCN+8mJ9nnTqTWcs7Ir1LZ8cdSlYEEzu
KCx8K+x7bV49YCwCG4qCrBuNUnX8cIETC5D+xZ71mx1tzEnn32oqfRsQLiqG
2ay9D7fr/FLsajcY9Oj+rzQDWNOnCsxoDTznJsw7PtH0cJoxvzz4wJSrmgBa
g4+BH3c1EzLpSqnMxou4tCIU+E9LUHv18cH9IWykusA016e28uhvo0Nf23le
01dknhWIkPvPQmOAYAP7xwwoJ9sGSy5bCxlbnlzupkYiyv+d/tVPk+RPAlKE
/NCT+9gaUlADtvQYxNGJG7HgM36pXqG6QqGQupFp2ykcP6QBfseXte0r7nD8
n4UY48uXUb+uRjz2jgFY8gZv1snYDavHHb2zxmCLkh4p8HTvoi97gtATdgRd
M4VpydDQkV/n2VIRMVTmin7NmzcecGnhvYGV+hlhghG/s4fC8L1/YD98MNa2
RGsZ3v7TUGD8wUpfe/sHfs/I7SkZAha9zXrw2sNZIoFTsQdyZJEkbCbufIjf
mvFLwRR3ZU7LKPCr66jRw/zvfcvyysoRqMppNa6ntLjgR9w/YYXIy2CTLe1W
eOipPi/SIRFwAbxKuZcJ9J0Y/msk2fdCVJaJaeFd5Wu6ybg2n8TxeRbtqkAe
Fhq5P9nodzKKhA07JlxoYtH15V8uD0JLZzvVt3f7Dk/W6znF3SWK7ZRAMR/9
IAYzltIlKPY8PobIvYDwFB9nfcJ774fsIgCnMfzNRxnRU8hD6jWT1zW3loZj
k2clL0dZV1OKz2IYy9+AlMp4oj+fwBX1kSrkfuQCssAOSywVaFHPdJYjBNfY
ZqT9GeovFSEEJr6fp8FaRILx1wiLl/OZ4AYGXd0kSHcmNgIlxq7xVPLTOaXB
WCnMy0HHd/OAzfcPTrzrQqQ29rYMKE6uJ9aCD3SoWujs6HI3AfsghcbPOczY
OIMNuPtTXnsirEYmolNQc/5wQnrFUKiwAkCC28H+QDVMFDkJ71vokR2tq6PQ
NI0eh5zq0b5K8UpWRrZDJT1JRHhaNG12UmbEgwUYEMPy9fefG6i5serHJ7U6
aXq1CV1rJ/b8XMF3HCsL9ObZNtje5ys0zbaJKlRvaAkCcnjLJtTjoXvkHhwb
JxC8XNMXgyPz/6BD97qpYSbYpgFY5ye0V/MrcBPEZCqJKjcJvcwK0Z/oX/iH
0hCyeFS+rVmwqwGcOpyvpe3p3iW225u4Tka78mNMP+XzuWFMsj4LGA6WhUdS
ha6aBeiYwc6WA3r9EIsgTfUl1Li7SxVA1KXXmqfNkPMIY91ewQXYVXJRYRk2
r2Xwni32TKv4Qq5dkJr30oMLoNmpdQ5JF8MhhRnMFVXIBrV+qYJvqIIRjsCS
Gn3UpZnRp03U6iDlk+pa1gunHMrmPCB9h5AXLymrg5NoVsgNTVLoAc7uvWKK
Bk4F6+fC4WycyaDgRityGYNedCDQWy86s6bVtZsWXwGIRC9zXnXn5eYFxfcO
BxMdBl2+8FG1EWCmQzj8vOpxVGFi3/y0woFzTtt6vlhVAV8GUM6gNF+JVjjA
bE7m3gX8RQj54eUuyT51dW7YJMrCNCrmbu+IyEY8vh92w/nhBuoWz5SiwP+7
8aVIF4Ct8S8JLpP1GM7AJm5DxI6xR0d6JdNAkZaRXAaUnjc2wMixbeLKiXir
Psu3z27lt5tty+gEv3TnzkAbJQ/AOYQgFCiQw9gQoBWhJeca7cnamrs2/amE
eQlHWXgL6ZYsWXJHgHeSyirsVoybk+x0InGiezSTAxoq5YBhI2qpTkhfmiiD
EYGzrnx8VzyjvmevtlXHL0oHejbEzIEcyUssB3vnnEbB1xfLI/VOUATprtpP
54GDnTW0yw7AF2hGyDLEIkFyd3POmih4vTtWnCB6lI6Uuuh4r6kMc8RfNObz
z26DrrIiT6dtPd9Px0Qcj78OzHVPDp/QyfJhhwkxm/FJx9ENKYWmQMy7Jttj
0SI8eyDxQIiAp7/SBvYSdscbRXqXwBMMfGES3rwT+LXP0/8CJQ4RJ/fBmPxd
sp9VKJWFWsDO4jR2XBqs1hdDnIdiMmFCjkTL6FqNY371Y0RSwwdvj4A+/ndn
heqma64TUY0UhoJarv43CmGwXnanmS4/PlErEvB/9sjyLnvUB5rpYmoi5EeZ
Bs+UpCgtWPN5WAxTHuK5OEFx6MAU47BcgeeEX0fcWPt3bsipk6lNzl4ZJbBC
yeeREmz94roYdbUX6vkKqSgk7anMdUMg7df3uq8FGaSH7aDrHiKB/NEtJzMW
VtioGzw8iJyAJkHCHaVmk5JoDlM4wImSXKILvg7FUNG+w6Tu2fop479n8QU8
SGLtO0danZ2lGvnSvxJ/7xaUPpE5xTP9S4SAqnrzkPhs2HERNo+VJdfFGAY+
TKkx0mP0MlgmtJvreG2ibk6EQq00ZFWzwGtR6aEk2V1ebHWYtTueniO/pv3w
J/Zm9PbrgPqPfedtfsEW5Vf5vYFDVDUD9wyTLWAoqID1FSC1HkCdhSJ5LonY
njqPD8+XjGjW8qdKP+W/piDPb7gtoWMESpGjtM0h0e55OsiNmTnhxCQmTCL4
0QJ5ZTQ51eGlXB41IQHe+nvMQ7DmJdZOepGJGI6kcawMiG1gIx4GCPbUZAt9
E7yckb05BKpRVau/ha5YgHLSzCmv4tGPcVRaOgHDF6aDHMR2VMenL5P1Aecl
2iAKPUs2613sLbWor+T+zpeOw7dlt99/bF7z7Z2GuVvgRIdFcaF3LagEZZSn
1cNi3pFpqeXIKuSWzPWzCMHGpjdrG1vy7rHiEul5FbwT9+pYU359qtNXaTve
S5ABxh0+bZvDXFH1+wCgjsfdFrn1J6a6EiEQ8eCxZFPfFMMl7wOgQ0JhencA
E3LLVRTURLXNhmpXZqifgnnGgGyfNP1TsqtEBLwjwT2NRCtvAvWKgg1kiMsC
Zf397XLfZczv3YTQKA9sMANG93NpvYPmLHJqIjtZBeAGgBHKLDX8tlYziil6
ODH3WKTKgTSsGRZjQmiqsRON4UUC//P8u4rl/SuoA4eVQsfQ+1sU+JvUlIN6
IQiULTHUoqM3+U3wEWnri1JaffmQvXJl+a6hTccZNPgWLlRRgeuH5F+ZgBd+
h16NJNSwHHoUjItxkfMW1ffD5yWdpF59XEWcoed7gS+mkNHQdxJfw4qpD7Ry
sHwtum1JIeYO6/NnFkZzAyAZR5YiNtqLBFMmG7/a/qUWZdWX74E5Z8ePV6NX
vlfEhApz++UqHnKfflm9Gjguf5w3xl/CSOFPY/k7hnD5p+sfkfjT0NZDHcEM
DZVCzU6cFC7HatygBuc4qCQ/9nY0cyWrBW9Zwdo8F120sho+l1eKEoTJ8y3T
gmd2LfLkH1REZdVABUySDQOS96DLp9sngjgrvNe6wd3MJUR11Gg3UXFweocG
9ZsCYNPXwmV5ekQN5CY84TjbmZzR7eqV2adrIXwwOInJFLKj+91o2Et5+g5z
PGoRBkBhoiqYq0IH/cjGIJbB8B9BGz4mpfupi6zFk4spaBAcQyCtnWNeV3oH
Fip0Bju411RhdJUdcLTQjW/iNbOxQ3IL+o+ZWqCxXBnAQk2nQ5uvgpddO+pg
CCOTOOd4+AciDFCOuMxw5tiIEPwS4NQLl7lshk1WYAzL6ldu6kFqQcP0L0om
AbeP+ZCUCTlb3V+xzOBzMcqNs4EL8zQ8LS5JFCZm+y/flB9oWpgKVzGymbPY
NQtXOZgfv+ync0bU9jYiJKs0yy6lFWK8/OolFN/LT4rqsuMW4FC4/893+qli
/+Mvg+F3cemB/2oZMZNSix5S8lKrtx8Po1328dfc3JVWV+sYah5op7BHBX8R
hf8dH0cM7OUAJXiXd4OskZYlkfA9oHp839rPWl4COodoZ8w4qte1Hc79rmQp
Xl3evJryz7PEAErwf63/q8EDvYh2TolnZ1qe8at2Bzn7a4Q0iLGSt0FXaxCD
u/7AUWM59Ahhh0eT6OvbM75UoofW8cTQqJwYoyv58I4pNckwL+5im/lYeq+A
iEjQAzuFTouH9/Vjg//mB7hvrxdYENDwIw6TvjpFP/1BIE96f5t87nx3PV66
mgRIJQrDGK5E+hejnP8NM9EUthlpx/ytQQqvmXob4GpKPi4pDPQWb+SW+YP/
gSEZnbtE+fRKiCNrofIFLPx3n4MbF0zzKzmIYzLYTeiKfDcrCuKj1tGsnbIs
vLhi0OYCqS1EYBgUqSDtPXZ7r9dgkGQTZlAtp+R7eufdV0nXPARvtdIVXlv/
GIUWJyzq6v9zSOAcK5sBoAQViLII7xL/MNDMueVN2Uiv+ylyI3/FlGhD3eDb
lyegVefxCEAuYy9S0zqYYgbqB6bEdyh8s0bWSvVgKenJe6K2dhoxFGPx/3I1
Ot0pvLG4UQcB8UqyvAvy22YH0N+3Ybm2B8pwUx/8g6lvFfNeWvNV67T5IgX+
tfvXFu5MWBYsZBECF2QCKroEP7D49sCh5p4KiS5HYp65XkGZNVtyuXz8PjvY
SGsfAbUWs4HpSUh/BrON7iBsU4byBkmBomnJan16CHds6xUPMvJXgpWunRS8
kD1TZOkLS34WbIcqa0t9u4sYNUyQCYbOEj9p9qH0nxXvTsWwuwj6q31POtqq
aabAKbIj6VumMwkgbaq973UvdSvQ0yBKXYm2DNsL1sn2bdxLe+xU3OPqWahe
aRPqkqx/XmYzsgAmTohIa6Mo3+UX8eXfX6xRuGJ72iOID3MoIS89nOSAEhz/
afBuqEPOFLQ9jtbe4dD0AiD+E2rhagiJFWQhDMhQfaDfgZsvCAkgdtuTF7dD
UXJLYsfllBZNkDa2O93l7M8O1bl4LQbs61YZskx/mKycfXIZ0ABP3i7fHbB+
XtXPg8DPAYPfcOMNBWi1XPcSYHezWgJEGdb7ODmw4Onad+ScIyYS8GwmH9ha
6DHZk/4W3OodirKrI+NRsjTqVrmuSy4+ZEh/2+o/o6f2uiYWozn+xioVeX9J
0hO56CYrczWzaRa6gZDYNnDcNJ+NOiLsA5NSr19yF0HmRI6/HyfXatcnxwk/
u/Cmcodt45J0lRt5eh14wwPFiF6RxoswLAh6dUzXBnbRZ818FkVzGZ1YhdOP
XEtRdqX/p2f6I6g/onuQXbqFQCAtACVjP33P4ySbqsF96JdNoJRtc4u3F8gh
2g59HaL8fjN6SECGY0thEKIU9tLDuwdQDb3Wcol/g0ySr5JlUaVXurtO6oNW
E8vkJ9q57+NrphlMntW00L6ihjBvuH+FUKvkXNxursnw6+OzawQ2K9ArLADK
Oy/1Xf+6Gh+caK20yxHiVaSlU3u6k6MxN5piMQN8szOLdDGWmdRQfjM2vXXw
60pCVuryF5ZgSwQ6BlI48fUQdrxOSSOkIrIrElS2dfIOZ0J7rl8POKgKyacS
NP9X/UloRUVZqRiKCpYNB2BADHmsYSbj5piaxoyA4c/xbrEMuXUE+KUpJr8Z
Yy6I/xnWSOdKXfUZGtf70sEBAzI/KZOs9UYVShFUbnN3cl0X8EsS0oJaMsOt
0IJcKQdX5A30kYwL52rMp85ZynBjMxv4Azw++tN+htjF9G0gtx1FPVoki25D
jJs9hdWhFvFonLDpzvi1a2n8uR6aX/Mb8ttr7nPdKOtA0TeZm+Go9puoYXhh
xx3+nJMXDn+xj53rrRh82O+GDCZcJaosa/MGjs0q5YTSUBLsbi2XFJ9woEz3
nGfZZhZaLDNGaY9BjEi2qEhG/QyP/+cp7buq9awwOIGn889MvngEMiKuU6H3
sA8vjFl2nhhdg/Cg0z5bvLgMi1rxbaF01ZfyIzrDiNBacGLqsOMmy7oP2eA4
TyUmAXs62khK3w/8EhpsQ7noPRevFOH1MMKIT71VbDaT61JA4LjGWhTqxRIo
b2NKmfRwC5JVL3yYBKoSeFAPYDrFdSiz9yU2YwkUbEUMXiapO7rfH3D53T1F
Bc6AJ1oRMlV3kh6p4L+kHAAuytznA3zG8RnjcgZqBVHnCeUisFShXgWPdmsG
CfKMZTmm8IJohJ0yZshDK1P4a+ptfZu37HinLRz347VbIPbD4JXwqMg26Rfr
Jmp8Pmcikr7xNyI+2ZfxNdzeZrFsjSN93lExJlHBfHjL2f8gg59uFaHaPxvE
MPyUBSVoqesYM8E6QlewRZOIfYzRGIbLMpynzXzGvkK0+VaRaJFLmmUarsP9
mp/hpAvialCwidxmcoiwRn4r+T6VUSwAwNhvD6VOsi+zefYU649cMBFQ6uaM
owJiULUBQA1gNS1HnlRbkXCE2/nXwCRX6iDsv+ybTgzNUCzpwVX4KT7r4HZd
2Ml9wYKj4ashNPF4eXEJn/rmBisGyXpxMwcl9vTKW6H4CIZYxjbiyaWIlv3a
Az43xqJVIRPKZlcabfx0IGb82LE83NZIMrJkodSbJWY5sJU2rXaB2qfghDzI
IapsgnndXNv6SSUAsLSlkL10H3/uxA40BxZfYnO4cd3ZWv+e3VPPOiAKLXva
YO8jXpIdghQTQGF7e7t+sL1ByUAWaG34ObYktfmrJ6IhUIajhQhtFMDG6sWZ
S9HA40BznOQbW1/73zDxOZiI8m6eC+3yZoxdaKgED8b00Uae/tZveYI9nFyO
JD8PTPWYaHAO8QALIUJx66hWJzz2nK9/+ZkIsmQAnFGWJGpyk9vVoOdrINUV
EucZPXrnabJdbm+MKOyWeGh6myvR2uUhM1AMWgeonTiFXRqdS1XQdi/cfiGc
yIfI+V8ZR00iZAZMx8Ngt6vgIKP1Clv01+OlTCsKouUCDfONaoXS+57mDDCJ
X6KZlqLynwWwjb0AySggLXEv3Gm/2rJKN5h24T5O1nZEiA6eO5jDCca9koa+
vxWcVBQsSNv0pksc2SSkU+C0D76bIYbK5bceC2rT6k8LXzwV6UGMt2j+hnHz
KNBer8jJqM3rjquL+gCzv5JcjQ/FQcgnPsUcF+dvK70fWbNMsJ5o2SAUHB5o
n/fTRzu+bbZSldrk5lVaf9AIxjVipH66wr64jLOGsEtLPy6wCuFZ7sjj39vG
7vhKM9SEgm+MAq9jtjXoEALQTCyHSdTtpNF+lqRWNv8KSMtsjsX8m+QyNLiy
4eIY7N6X0W9faqm8uk4CfFQHWJq80kvmV5iDPcqfGG1LdH++uEhU8LP/+Buo
rtTM0E383YA8EsCkx/dXrG5zYhbwGsIj5nTDsUeB7oecBFnLSGnz557nrF8N
X1LsJSldxWO9pSeutIiBytMI/leiUlz4APV/HqfdMehemW4+e8dwrEY+SU+y
K/z2r2wNDeYOVpb2MEr879lR4jjrySDIx/ot7P7kCxGaWTNbzg3xMVpeh58B
1X/tuUua7JB0NrmrI+JyUYpObQL63lMsJy9yLTv3XvmGn8mIowVSJ8u7ikiS
LeGSFpo7tHMdBsp3lJ+YYWZiS9e1YDyRwqBHSpN8Nb6MjXl43PT9AYz4eTOQ
TmY8d9Kg3VZryiCJY48IDn1Jq+FxRXg5tuW5vI3Lm8XLLqRpMXa/UnzBGucw
O6wYTqc5LcsNCyIDLBxSOtJmxu+e9XzHc2TJOy/8uy94iRxcgSX1/0YW2Qli
tm0HpcEVzlOY0WLuywv/ccuHHvUfNNpSUPNbmP2WSWFWK7bBxg1CUyEeBLMu
HweikwX6XNWnjWVLoi0q5KYRHqeajdRIp/gce370jyixrHlPLqDEuohtJzFD
9aylS6U10/wicEgD69J8i1a1J95nNAaKehrEI4S/p6TVmTe9HPUwnsVnajQd
a4UTcg1bROXnctD99aG9VcBwJ+eg2rue365WiCIQISnteLBh/8iAImUp7694
DFsAp6vm45h0iLhq0fgVn6uz7PqvS159xAmSjTtnipjQS5CEO7ZcimWClBaX
q7e3cNWSAUkHFxcJIsUsoWB3Xfk5iUzltYRSmxyskVCJWzasKj94d+oHumbs
6KaxQa8yepko7cgr7jwBpYiZciXlNKHxGLoMuN4v1lfN6dVtA//EQZxofFPy
q8sx4vuFFSpA3Xmuyb9+RiZ+onGaCSgo2nbwpc15/J2bQDGW6OdbcB+emuES
wbyYSg2V0ZJ9jiwyri3GGcLR7Qxi+1Ah44Jd1Pr4Muzrq38J9k6WZmE9rlhg
etaPcpOBaVXP8yzT9HfWcHU2uL3+DtXi+vGvV+j1XO01KLa3dEEX2Cai8NvI
m3zL0zC/DsQGLyeab5qXhfsFxGevAmXil5HkvbFGf/L/Yc74SIBum45Bmtty
2G9kA9EsQqP+BaB3Ohnh5UHFU5+cb+uv30/46dx9J49id7/cfxE1pJnOHdh0
+o72eqhsRP6BGKY44Xmc1abAKIeERPefW5UhYzUU0zMPX2HlQ8OVl52Zh+Dq
S9iGNkI0ze+4UL584TGG1pK0Y9fbjDmRpxIBiVX0IVkpXaBoaIyAX0ygxUOb
DnEoYkis88B9C1eRt5fyE+7GEKn3i/VsMlHIxANaxXgTADJEo40pxaF6Zfi+
YmEnaWPJkhU0bTRQ4CMRMNs4qcMXv4DvwWZA4A4D9LVKHWlSM0odZ0RhSId/
E5hU/TzdPGCntZpExd77eRt/z6xwiBMBAduFtRH1dNhqDRfBTsP+hqM+D2r3
JY0HA+P+FSAHKQ87i8hRV+FkgFci+fMh9ONhrFbPLpHIwS22BDqoVMnlXAem
m9KfwZFoLkf7A3hW8ndTtiGZ1JuPmR5TqYuFopArGmqDtfrQ4reZPmdCqe0K
uXDCBclor/GfrlKcbGliLCClLLFiHhfAMVSjmb0+HbnwwbC+qCUtOohnBVIU
4v+pelfeozvOCg3TR1CwBaUTzTEEyDjRlKQzs52vfVMbylwqNUuEvtNGojhz
EwWjcVCzFNt8vHiLN587tK4fNQng6ZolyCXRCvc4R1uKXRH1zJVqJxIa3Xbw
nI++6wj2hAJmewgjlcbJ0eKe5vXVo+S8ixMNwhz1G1SufOHPa6S1DwqRt9f7
WzEHAcOUmauEzsfREgHD24Xj75LliiAE6bIurQGNfbYA2148bJXTLLR3BRZ7
+2e45vnNLUkz1Xsah8M+wGdaMn6ntpaXsa+p0/1Qd6jgKCgvXM/s28TjzujA
Ow8JUL2UwFvueciMZyoApVpAjv3hU8h7rqwe7PMukGozYGP874t+0Ud+AKN0
xF1x/EZ5qY4jW8WzeNKqUjUc90MuvH8nWWIpb/9O1a9x03u56V2EmJUwK94P
gqV1kTFluT2dGh+rMLnqumdhi6bq7bPKNteh1gOQyt3wPzqAnULap5NOs6ed
8CAEa8aEomWV35SpSF/+fH71gqzZAeWOaHQebZi2MRHN9H723LPeeJH/r4RS
9FpF0jQZj12u38iQ6vkXh0dyxtU7Ebc+emZNBPW6GJfLtz7C81PUIc8ddCoi
3xgtVnqHzg3BH6nKq6VCT05Y7g1jh0A85jJETcHqscX8VeTK8iJ3VkRlaO7R
xq2NYVLE3jVgJ7hWqDRYjVg83spw4jBzXKVF89/3PirEJ7aPkUgxeBTnYhym
z3RanbJ90WL+wtkPoFj/5h2rGSFmqZaSyikBtQunhDcBC+BnXLzdAQB2EyGf
ho5qye6TUfDwM38Pekt7WZqCkxMKMoyvamHETO/NU8BvP4fEaSPXEc00L9Ir
YPJ/ayMX332GUhS8ecuoIBRLpp0cLk/6aDzxP60o66kcHGK5q5tr2VT6waMH
AfeClAnfmH2LjDE214sMNFy7sQT8rnYes269vy1v1dEstMDODkyV2UXmOGu0
+PaYXJslOcb1yZlic7Z1jW4CWlU9MrvFqCB24hLbkhfsWqUPSSYTel/0h89E
9xWUkHnJwvr/spZ7a+m6HIcRZV2NbARzSPAOt+e8IPYr8lgmXQ94/GcpLyHP
Q+GevW+PlSokdtF7sgZsbE73BDwoBDSb3u9ivNGFG1LjImEEBfP9qc8W0scQ
StoQdXTRsgCmJievxEG36OM9bPRzTVrhBk/BWwLCu/9ynZX2bEF1utoAUXF3
ujndkbVMLdfc3+r6NoTE6EwgHPl0iHU2ANctTauP0ZJ+XDFfWQahZXhbfpYJ
9wC5Cfd4B25f3zGQUHRsqCjXAJkZtbZ6W7pOvWDEBZPedpahUaLS3lFuQv47
iGZw6MMHxFP/IyKuDkRhlCKhVSooidYXpmqQGgw1hv+Fy8oA0DRS5uiAQuBc
VkdVxrqwZ/+pmuVwqavN4MYJK6FYRPJ8S+/Ev/Tzf9NTDYSq+sAuqNm6IAws
9s0z+1fT6mKMxKOfoBKXNWlGOwrdh0llez7L8/jM0ZOLU2gwbuZMBBEoFBMD
ntccj5++mSlVFu2Sdp35ai61A65UX4N4G1oiaCX0sjyo9Ckc19LpLEOfTa7f
MpzrYBNFYED+hiRwu+CNN3vtqUecCC6SIQlIPBkcbhnDqxRj45ayKl4vVicq
1wlalbWp4FlTV4RcyOZfMipggghnX90G7wLUjZB3pp8wIQl9smBZDOf82ivQ
vrf2ZKiFDEHvAi1eEggMOcxJYBCxnKQ1Q9MuFruMSEs6vXyXuyOn3PxZ9sNe
ODHrf1pOt7s9CAJ2uv5ZKJtX9LEnXl6vxGAmGbmGznx1p4ReePOtE+OummXa
iMqdjrbjAG74VkPY1nUG40KAFDr22/Bz8P24fjY3YPY9ElXqaCjKLWc21j1B
xubJepuQJ1SG2OILZvtgk+dk2BFNFa7fax9ARGx+kg9VHVJjbmSRquIBd0Dv
XLFCWMXdSOWeJml4YCCAvjregvT/o3Z1ifOidzDJJawF6UvGpITVUrhdkSYP
8BxBoyfOA5FpusqL4TZgiTHGrWZbzJfx8gCI6dBi7Mnp9In3/Mv80SdOn0V9
NCy6Ug55XaoVJl/d8fNf5DF2XyJGozIsLiLNJYS0iQEag/M864+GSc4BHNGw
uURW/qpUbmbRJabNTYNeOtltwEF3q7jOa7uBabHSrX0xsatBbJwTu7X2YQAb
q3LOkgy6PhsbCjTcIW0tS4Vj30A9Rz+FJtKAIwm9zk+uvGkhE46GvCbpHxW+
j/1fQbDYvD6lWothYRnCnSeTeWHlsZRsF19bJC2cChoRoFZvmiak84fzlVZ6
bAPMddsfQpL++OlQb3hNsm/G7rPsy05TiIbbHOplwOFq7Ngfd3DqdeyIxxxD
NOBjEauLNhG86hZVIplq/m4RiYG0HC0+vVEnr50NrFVQUO5DmWJR/sANPOO4
ZZqZd5VszhxMR99LFcRuyhUbXdmk3tG/qRw+H1QtmGqhGXvuPQxbO0KxuHW9
QrjBoduICehWBUvzCnnWIIYYm+oCJEGyxD7tClUD5XaWReSPchlJhMdp8MZf
UYO8wMx9i2nL7NTTSTDHF4q0XSEMmOquJBOW1L1VdtT+L67P0z/cKV3Bfwpt
db69B0NGUKuf02+u2+TXoye0/okCmep060QrDIUJghPkut4R2cQygiQ4w6nc
mIp7o1CEnZadRmBXNlor8MZkric0DC7UlZoMX0wKE8UZTvS2NTXN3HhCTtrD
bvKOeCJYj9Er9HDdlrds0WkToctgKP7vPHjkXmg15rJr+gqSccWvrYtfX7Ew
+qPYcZ/F/Ks075oBTHbh6064cZ2J3qMWzE05x/lI7VF2JeiCkTWYkXzWRQaP
BAIS1TpvlwpoHZ3KSvYtJdpivP2cZDMj1nv5O30fxG1CEhuI7dKAnwx9r3NR
jJ3mMdzoPJ98wo2hR4yppXdSPp6M066aTVhP9KccFprRAR3w7oHtFkFZoMMd
/A7fkV8aEBOIY7E1+jBcOz/Lh7jZwdD4e70wy9IMLqWdEFC8GI8OugW91zzC
/0LBx1cDGRi8oaG5luH73sWjwEDWkys5TZoEOu4SpV6+QmQA1xanqyuDO6ms
ntObJIfOWDOlb3B5ZvbeETb4HqElZKtq8XnVWyyYRalfHMlgK2u4yQ7Eb8hQ
QQXkZtEx0kG2ruGk7DDwfRHwGicckAqh53tA9cQ91leq4BCMq3DHb46R7IuY
Zvvv12wKZeAZ5xFFjak8BGJV3SqLKqbFua9D8AioKJYUei34pPAwo7QY8Ua1
jh+DEW7yqkcTme4QDAN6H+rR2kv/FwBdtcjgrLBJseuXsyFfHjBrEN81T7uS
KS6+nihpfP9KBvnCoLDnuCgE/KJFQYtl60d2vWJt/IIZ4mAF1PWN7FQikSZO
AKnC2dEJDk8ikymRkWOU1CDu/+BYcWCOO44QN29+TlJfO9rH4S/xKZnu53pN
OGH/chX5fnzgsZDwnaTo4/Opply2ma74qpiALsOkqerB5RLIDQcRYZCFUwVx
xfGSS6JAcnnMBdZWWkZuwxtFVCxselvOOQ2NdzbN1IyYGJWRJibGb+pwnx8h
eJxa/4dammqlb+jGqL+Iwvrf3mxpt5s9mOsCdBuAKulZ/zzsqY5PZ4p6KpoF
Ez+ZkX7/2UMlCfiKCLRp71P5qqHQXfMjfcooeKrZ2rMzNDnNaeNWKqc3vTyn
3cfADEmkcWsLCu2yAlUGwkOiYPAR/+8RefnSeJFi9WAlzu18Cs6Q/4+P5/SH
dNsxHSA1W87aSQTE1tFdkpjlSlieA+lguwreIC0LrEsbPEesAArAXZ2CSe0x
+I0l46/66nEqXhWOrgv2NmKw6AkLPfu7Q0eWx+hZp5VeaUuNATHa1T3DTn1V
53oodrPvefZSOE0H6ZF5I2pOool7vFs5cpwJmeXUs05yFcm0qj+ppzZyESSZ
R7oqgPWKg72hpYOxfIcZ6kq3LRJ+yO0qMI/YmVL4LNWaURLDxIL6YlMrZ3yL
mREJAudvY8r88bnUS7PFAz2mJnf5TFZvGFWMMoP/c2wfXNCR9Vjl4mlPMSBJ
PHmpcgYyyk9l2jcOg5WsDPJe0QHifcFx2KSxEjj5Hmv8Gl7oCCOMZFmfd5x8
6+5s1gi/BSfKBD38g2OMTfL4x8R5XTkQr5IXcIv72jw3o9a5ADf4S6AIO7co
7V2SbUuOt6hTt2Qo0qUiD96oJPmrEcfLi8NdX8NTKZmJ0XxUQS+RRoEBGIVc
d2888npGiu8fpPp2RLi7inz9ymbkxW2AiFpIXpjixNpNRv0qSsPtz8z7zE2I
pqprht3Hj65t+llVzRLSqm2hLoj6GL5fwk8It6Vxl0EM0+Be0UgJtHGsrfdY
Vd2Dzzvu4jfa/lWHXjd9fAPT/qjOyyEk+fbvB5BmXSb04hnouZwY+jF7srA4
gkeeUSckjgM6+tIRqFUR+0OwqND++MA4a3gxg3TVkUP5RbaJo8o9g1zOgaf4
ScmkSN8pBQh2va+TL39jkYsYnys9wfdfb9RVYuHxHpLXDJHq2aoTRFSwe+Yi
Exo4TH3NeIReTnvj2fsbU4OE3vXHJm06/21LM1c8kpIsawupHDcVVmQkdPpw
hfA912hcX07YKAfhUSQmBPy95Yvv4NLpYUUqIHYBSCN03OUKkSNo5h9xRuXn
Sf1fE8dp32W2wjLics0I5jJzDPyZzjViNEZAZFVSBnEnHgOJX9lOKlawt4ko
irg1CEIBpmewkYuNgMd2eKareQkpw1kXbt1BQOkjEneK11Kvl6Zuj9TrvfFP
w/9JYJkt0EaqaqJKdSzTkVbB/g9Vp1ZRzPKvmBaSu7H7uTtjqbxY1G9x6NVj
vGIksjSD15h8AJDbIctXRSr/9depCUjc3E2/edQiRgnIFV+N8rTzwXUCH5Br
pbxpAjDiprAzHYxkoyPqlHsI2PV58fLywkNfPD1IYvkmVgUaebCEYt84k1ZR
dhcN55Z2e5HDkaLiGCSALhLfpBvkpvHkc44jW9WphrM3Eng8cI9IfAcLvOqD
ueXHtCv5I00MwG2W7aXpyGRNOkDdH1rDzUCExh5k/GM4NqZTOk133UVM1OIt
XqSyiKiR3VLxEyfBwPbr6fjatb3M2EU1p7UhdhKe/h4cgLUZp2UqGV5AnQRI
RU7tRFtvPC2BXOUjWEBCjwPEvX9Nzl86RZmNB4q+76P/XZRwqPS8lhVxMMvw
KqDbcQkXW+yPWOl+7mSW6FHr0TmWTHpc5TCY8CsvM6fe0aObQRpkK1Wo8Zd2
8k/ldewtV5RIhWfrFGf8xoa02Oo5aPYq4uKD7SNgjeBUH+6StoQvZVB5CAxI
EzDl0PoPuEQODykf0FuwNaEiwimF678ibV9LXaFICQihCjg/UYPrDoddBA7e
q1NJqxD4sDIRG68uY8mJtdZkK5IWYENbonPM52xH5AnXMo0WQ2czWa//TgyX
NEFmUubm8URw1WASH/XTNs0QuUtXFsDWmlwAP26phLiXicAyRjmIZqaNgMhf
H27Gny3osjQHXJsFY86OudV4POWqEqYVG1znbsStt9fVUZ+wdrV7FjD7Ols6
k8ec8o1Qbb7LE7xutjwR7GDX2hl1smBcT8UNRD5QK9wsgjEHcFSy55ysTdxN
c6BvOS6PhFOkJ2xdIrRFdmemeHNSc+9gbGFdowXX/En24I5/ga2nV28q2Qs6
IbTQzvcnUuJPi6UI+fWhG1WK+V2h4fiSQcBb1Uz3EYgw7Y32Dc32zcwdubim
hgWF/HK610OKNGQOuwhlT2opwAMvsO0lawl7oebIUnUk0akdHiarf0QO44nv
1bSNt/lgHMSkqXLDIcBuZyzwFA0Fm8jU4VW3njtl1xfZcxZvdT+emX52LtB3
I+qHGHDBgaHUmxOzbv32GYO5qJqbAvImVLyGzzfkS88uoCcjF73y2CU492Yz
pIDlO3LhijfjszS4Kd6nXG/TyMf47iSNMwWnrE0M6TOZFFPQZEWyWC4AV82i
we2oszRpT4OkPQNSs8nzF1SAfOvgTznTmBy6+DeRDLJF9OZg5jZnKAYTLVWz
aXjmfe4Hm5pHD+lEIhsS2zli4r/9hrFgs7VV5H8IaP1B/56r13ydKEd5a/xY
+UHjEr2gLNKYWLF0vVi+XPBEhwCu5tDGhLFpPoW/x0NCXA8BHQOgzc32tPsM
0FqctMmkYP/jgAMFz8wV4EbmAkUzhXR+0eGcUGoDXD4KgQ/60bIsYUquVjJi
fJ5xMAJJQKl+ORsvBb428Gq8u2KZzg2yTTfrgQphk4/g2sA+mhDQYTztQHiV
XLiesfRuwaGoUEhf/zYyyWX91LJIB8S0RNkj9bUsGR0MK2zYVeKXasUL5uGy
qES60yx/PoyXIw50PZzGcSGu/B9D4o7sdrz75PaoE3RzLW7uGFO1MqnW4YrW
Zw1cArKD3sv97bpWViaCTJ/7XxST136s3XGjslljXXzOItrsbO3k6cC24q4T
SPpIojUf8qmy6fAgXETTFdEEfGjx2/dxQrnmmNoTb9vX3B5C0Sf6/9yN1RPc
Ckw6

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1IVfKCQpZykOrjejVeYteci2Jn8PmnipTPDUWWsSL2oMR3vpCqf4Zbf+ALhmG0nsMbtF8znsEeETzNa5KTdsg6gQuJFGcxWLkH2oQaZLJaQjHNJ5sAk0lQYIyuG3HzQbDYJ+HBCtzBEJ0aAX9kJeVJ/26/4OzrlY/WyDLLrm5CiB93ZLIy6+vp23SD/vDH/uWLMAVoCX9tdJMyaJQDwv/L1zP4kcTF2rPzwS5q+dyylIgKanMRT2HjBOqRmJ6lTxLKW+PgFUZjzMb9HDzcgPjBx5KbZPvFYpRTKagwkG4HjK0vYF2R+tN04h+I2D6Bmbcytr1KzeRHP6wO5ig14wE6fM/JbhwLmQQ+camGCxIM4BnMZlQfte6RmIXrxEnbOIkFN/Z2AxzjJdBqDtBm6gcUGsKHj4quEMMmjpVKVV4ZRGX2bJQRXHGLtk319IXMcAohN8bI84hHwP2t9PPkuifxO8FrYoOLth3Ahedc1xSjiKlP1QY05zVvU3m2t7rD2TuoxhL15G4sPK0ydProAejkabWBXiezqobnl9eAXIde9lT6Ot2I+9JS4BIawCRg6xRJigXkebaCmY19UIwo5+0Lmq3FOeAN342OqkOOagZ79CnaASgmj4zytNg1f10w3IANIes8oMEshFfBtgFP+p9GmFc5smQDUFMG3okhT/fZyvRjcNYl3kqmx2rjIVw/KUZeCWDWRrhrWNGiMOOISmXUywCeQx1A+WL6RVohJX9vGdWW/VNBCGRiCKCIv2PoaBTSJKvRAe/DVNkhDvUnVip2y"
`endif