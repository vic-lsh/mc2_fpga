// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
s78QcteWTRJZmstz+ODay47ISYJLQwzaAEjN0gk12qAHeKYYmz9nT7OxCwmD
2ss0eZqPQk/t1YDS4gMloVXYSEAZajxo+MdEHuLWTfOmevIrgRzXqBNfdvws
+mM0A9o6AaLS8Za/pL7H4Z3bznDrngm+EI3jtgiiFK0a1m44bEBU72MxVvIp
Xi4YOmH0AkmNeY5iv+RjFqM11SDgiHXkLejhA2JJdYgoWz++2B5g8iuv5ZUU
y4MC4tctbTqrg4UepZ1Zr4Kzm8idbXWnjVSpIPPhfA8eBkIeGpxopY7xj8Hz
J5GObOI853e6Bzgq8yE+Xmvkbtn+KkvG7MyonQ7Yxg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ogXVPud+R7qvUChnyoeuKw5kSDJh5ttF3gaF4vQwB2lRvBp/3AhdoesR2QGG
D5oGmc5ER10afH6kQhCJQfwUwvkDL9ZjDF2Dd1/kOlotLiSMQoIxu8J2Tzy8
3GxLI8P709LI57f82Ap6KVJl+ERqq5PL1/7VNNGVx5xzYARLS9V7PwieSOTg
iONSNf+n15yY+lPz8v1d+Sie/e0siav91jLM4sF3+fd0Kckix5U5iyl8xwYe
WTGoByEI+6raPQzPvMgRnaBx1ImZTMhwjCD0LX8556AAZ2WJabu4KwjmIqiC
3sCIShAhOgBBVuxATG7xtSNcqnYS+pdJ7UhTnaa23w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vb6XfdSWP2nTies3EQ0vSXSye7nSxZhp8G3vdt08BHr5bFt5ELLP/iGO7Hvw
5RA9XI1PjWI+ZWbTNAFQ22+LKQwcVuoozCg9DD6tX6bUMhemljdx0I/yhHHt
DGLkbxaPwbC5MDrwlLIf+8EIzJ3hEz6PGMNwHFW6WDc8MFIf6LDta8QL9xHb
XB0qRIFCEPeI68PWLTwzXMczMPmWTBCrAJ5aNbaZ2fwkzXBBJ6/6EhDoFVPE
0dL1sAkDe6GxTm7YYl4/TIkQs20z5we10UR/0lBKGv6KNB+ZW//m26V795KG
8C+1U5ZzugE7yh94iToYgd0eRFFSI2GD41+ejI4Tfw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PMsusaPwpfC4qvDIYPF+5NDv566VAdDS5INC9PW9ZDrwNwJYAlnzxBOhoG0m
UqzDdgdVlw2QSpqre2LXtXEJNWIqlMzIJ/fb1aVc6ab6LRR5C6w1DziJV9n3
4abjy4i365ydurjYdg8htHv4IN3O3wXd6aNIrUv8Bfb/ju4gCiSzgMlLVcqH
U9KVX461t7E+q4/Ijy2YL3qYjiTLtByZ0bXHu1Sde+AhB46E/YO4XsbxeAQu
94HJXkND2devFks0SICzRRq6eMHBukjTbVDzCKejjvt6viJe5QbNRMuYenlL
3meBmIytQBUYJJOe8KDg1Mve8hhzlbu83xlQ2/WSoA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iP1Rras1kWjNrOo1LyfotcneDyxMTdQndx3XJSRURTPkqvbDbimXYojYA37G
Ou/twukv49Zs0R9oI6U7qiKuDAXMisS+Gl8gwVrqwopCW772ao9ph2/BPwfU
CycHXgD2BOcwuTj8xCjl3rK19QIuo1sypDji+6FoD0RiWHG3Lik=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NM480EToDg+SJeQysBY+0DSbTVC/xw23svoi6xHNOBbrM3R5lk1fbmB2uUQx
RIra8SwlEFSKekZ8s2ZzYSJhGHQzIMIugQUzIycTu49fOe7HzESOzBIaD+f8
SziVC+weFStyZpwXJRvqgSuDNI+8W7vCtWG1rqDoe7lSs/yFcaAgyy08zKxx
Sx/4IkxM9L2mIm3VuRNqekeDhdPcXc/o0I5aL7S9GszNnpnibEoUO0fy0PwB
h5IYRfNq+nzwDJke12UCudbdiTPX/A+6HYuwioOvzcvuRgD6bKAmjjPE/cSP
lZSaUa3GjCvEvDmmDieyK4RrIVYfoldHnMLODPHGZfGp+EKRi5D2PzFuVgUJ
QpVsuOBd519h4aJoSo0M9nmGwDknPeLHqtjG0Gn3NalH/p5PbbZvmFrGjxWE
PVR5+Xwl0U3k9qK7MYliUx+KsccUKlVpY93etZW9izovC2fvnZ/1lBhuc9eJ
cRORrSWsLeteM6ruEo5zk+mqgB/4XvIQ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nfgoOcBXdF8/eaMn4X3LOUFXdSsNGzxPpClWNA5yBnp6b4KO/j12uJMCmaaY
vTSpNEhh7YBHsmBkbgcIt+qHmmVnrGeElmVd7gghvHmeasgJPHx/Mzbjyf6e
X6MNk0V2qAT3z8OjDOcACNlQ8w7SaxTA4zsxcUz7a65+3l6Y5wI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FZN3Hukjed1gD0Y2twkJcQ3nMhH7lwSwMo/ca1vC8cf1IzQT1Q68nQc27kDK
P3EclPwlNxGKKMP2pyZro4DD/CkxAcCTFvMd2Dcuc/OzZreTvb2icBxZO+41
eBpXhAPN16zU5zjc/gtAALV2uRw3ALwLlBMGmlgKwTOItOjoW0M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 91024)
`pragma protect data_block
lEuB0VuVq1BJ1YBRI+BmO0D3zAnrXpPy0dPbj/10FNUvey10YAl61Wykclp9
3siRKPcbf+yNSiBvs0y8elgHAJqQRZXqokscV6DbZaR4+LaFZqCzokyAiviV
zDTG9ORYX9ENgqdXbv0ReLOEUPdWrpdav+N008HdYOOK/KR2iwvIXYuOFUI8
Bye1/9U/pdFIg5six/rDMEBpSQNXjZvcxYSRZVyPZwDuh0llpDW1/PA/ZfQE
FytNAgwxd+vHQWiTKpGZWPjV2HqR8ShIE1yGkOytmLWXrmj7D3x+HtHyYTCi
6L1JGj9J4kO1LLv+fNZSsDTLJCuqfqZYErCS8zuozZWRdf+J65IcjbBGp6vA
0IyknrOpLzv2BveVtyHgF4JJq2V3Qf3Mon4b05GjcjokuCxGA7QoxEB3HJiq
wKBdbnUzVJIpsfUZydA2RecwOvN1Jp55ivm23j81EAhN3xXQ9KGm25NLyc58
hvM73q4epTtzlU3zYbN8KL4oQ8k3ADWh0ho9fhrmWkLP7QYz7WL5570DTgPV
M5bO8tzECPWUMMk0L1OzyuERVzqA3UYlZ0IDHBGaPn/TSf9clzr272BlQnXl
NGacX8uYABOIusPo7yCtT+G3EczVO2ofJAFBZrfB0f2UYegzu7Ydk3ShoRQg
Yl+9qATc6d7Q4bk21FXgpcEyVWtdcUHoU94pIvQl9IUO6zsafs1xQvlZFL2+
np47PYxETc1Ok7QL6zbvyeZaC51kQKYfDWndp3m7hMEhY9SEnCc67f6VGLb4
SgogXKjFHprnH3OCSctioPgT9duiy0yE2NE1opssvFSuVQ8ggfulcrAYuopW
bfKB7yGV7ryFJ4s4KhdlEy07bJEQnQg6h33QCE8aIUxXapfygpw7G44jIi38
7YCqtsKcsqmaoUzcCU0gu7JLabOn9tmrlP7UmRicuSgP2KFm3cxtUc6BOm0j
6EJncSIq5Z4PhXUAK6vy1ynhJbOux25bbR2G/qIRlUic2crbtVs9Y/DH9GpF
6G3ZYz5BRWYjSEEkbypGKC+KgRtalh0eBpGR/Tg1AranyQE8uqaAUkHOuRCk
68qyaj9y4W8/2ftSGHAZRVqw5x5BtgjoH6jQSZDpPJCtGcap0xWRc5wapxHg
Fip3V8skCq8HThU+m8VF+1CG1F1nmlAQnvnhe03996LfTBK2nWlvHOKd2Vg9
eRaQ0IIjFxsvs1UDRYJzCLfntuulh5JFi+cVz19ZZQzWBt0yS/K8YZUkmBMh
Q1YAZvO387HA0Z3XLmbG8tVDXN64ly+ZMpa5jtnxkt3dFmv3LpQ2A/lbNypB
cwjWd2mlH8TgpftqIYjIbliIgwzRnl8rCns7gFbxUsEgWJTuT+nNgpNDT3Pd
Sj1JV+kfPC1JSP9XcTCa+YRXs7UvqCX6NicNs0dJ/1u8ChCNkklMTITFHjvK
TeaIQGb4ojU1Fvk7F+3IbJw1AJzv6z5TysYvMkHmvlNRQ+4DoXKzc7x3suH2
21krFrf+IHYI5UCdozDBT/mHcvrVD1mEhktR5gsmsSM253cgKAnId/MaYHqB
cXjf1MzElVkgdcoOtC/FkI7KduFnIobeCavZrzAN+n236TuS6NO3Q8/MWl7H
WLnOPQ8PcyRCc88QZ4lXH9Nf51QHFXjH9KckQPZtiDZa7DVmX1AabsUCKeI0
Tn31pUjLyhP0u8JQQfC5Ks69qe8OZHjYOaHLY7Xz1wP2cbm0GoS3Y2DHzLIj
7dbhchfbd24pkfwIyRijgxuK6neenNufM2NAMQlz1Aibb6NIvbrOFHFVWiik
3tRerW9dz5qR+F1WLFs4x1bif1A5S9gJTHF8pQ9SA/u5yu/cBeeRBFuay68Y
LoOIKdK7AJJCGiV8QscDGr5OBd+iONUPQUlqu/7aJzRyM3BOojDX9axQw3ld
7g0Xc+2qf2fgMJ3/2KaSEh+YpMR8I9Eplr6tNSxrkLjQ3YhhNyMui8/uKasn
rPDlgQY+34IYIonL7dyXPmgGV6DrrGi7lNMV37uKlL3gEYjZ6NuKo3v+z+Gj
XFVL//IBAfGbd2Ay6svY9V69yHjqMxd76e7EYOhxDwJcjhU0xzTftFrHSO9U
soTaHW0QRzyELdSTrxxR3tNKHXvpATYkoh5LH7xikm+CT0GOddMirfUNXDZp
cyASwDeSaR9UxSRApbMks4xrEc/Jn2L1Hg/2FsbiIDNgH1HoMZfDlwt/rNlm
syaTbGLj5WiGiEgTGIncAH1Gd9fKaVz7zCvynXf6NgJrQxKSa3Lhc+WqAL8O
WHzoKGJDxH8pV5/tJ0nfrJeoA02n+XD38H8AI89RfO40b7yBU04iEcdOTDiP
NuV0AxvZ3Pf1lXiRSaF7iAvpSN3MDgNh5P981eBamelpiKVN9Ri99bp1GeLR
Myua/R/dFPaL+7llrPq53Ct0PpQfGNQSNDUwVg4LrSrcN109cmO3GWmgi60h
fnajMYeePC17G0IBxxlm5FVZ2n/XZONQC/Qe/npv2EkL27DU1on/+8dJVTsJ
2fporsrur30SCGwfaorCfvOCtTnyGoy/QdNB7GllhbHlvqD3ekg3BDU/gz3m
ujPTQsKuCPvTVoLnf0WrRMTPZqs2apm8oyaIA6XSMvqQABJ+CUFvOeMfMFK7
1TaWJQ05WJKP4D/mccXhhNVs+D86Vos6wMNCPYvApAxipy0ahFQQ/UWUlete
UnmY9D+UM7t90Tc3Jdh5PWeBLOjxiO0f4COqhTEPz55p7FsJ8m9ndVWJ1IAE
cake80lRq7Qv76JPNyalAUEshxQ6At9v+MLLLjauC9kCjchvEacR6JdNthCN
ppapZeocgq3KAW3nng2yfh7xM4IINS/1/HRlzgSr/t9apR1rlIn9y+PU0L8C
w0iXN/O116sjennFPxv6aIeiC3rmeuclXZ/SxvQFx5+FGA5kkct78A1zELcl
+YRSSF3wLlM/l6ix76BLHQtLgxPo4tY9uNMUdUBaIkQRcfGTnKsLtxZYDCeq
u92ktZ3eMA4YWEP6XUBdROBSe5d+sjQjktl7wk+UX5DYcZ0SiL0+HBVpUMHc
J5tJzD7ZVX7dOxNMiWiS3QxwD3PDlxZJV8qHIac9yc1ytCKyFmaK9AmHdTUp
OXKHSLr90e0DRD8WBbNVJ3wiDTyh6druJbCNyydXHPHf2wWbMN2HwGovw6L7
YP83jpx9lVCib4/XZvp0TFORYZNI6hWN5bo0nEhQVcEdsp7rHoLwAnSP2WOB
iG961usB0N9WmhCE7tLyx3jRlUuGws/e5RxpPFjpS8e1a/Hpri9XNZpNPxIR
IZwo4GiFDji5FCpmIj2jwoOEfYAs0k5nbiFGl8QIIdKYJhUR5fQYL8fIc6MF
5AoDYoaeH+wOOlEgckaXzqeFKVnoLccUt26PVWZK7sjsx25nx6kV67ajLiqL
qCRSS/RhhRRoPuL22Ht8RmB+DrZWTH0thPlhonGa5lOq01AJ3Sq0srhhLV+r
2u4iaTdyqnszFioGHgs9NcFjX38IYF7dRmyAG1BfsusWn9WPzbBYx6Kjx3ro
ibcY1lxWeJYSM/dSNzwtabgmS1ZCKp8m9zFTgl5qh0DXCwcNvI0ifJ0qAp2F
cuohuWtvf5tFrVD/gY4InWQ4d9bwS2g1REwEKbUtBgpUeSXmOrEAyPemRG22
YiUGAsT0sBxNprUquAocJmRljukLakPOFh4N5GBrhdU8WxWz5OQ7JVuOq8Rv
JfiBY+5+be9F+bglCVAALlXjjIVJCmV4g80HsP9qHEWetae94hAGmwKFe6m0
AXTltSbHuZ5Kmp/B+ZZmVfR/aGqlNmRmBxFyd3pfPgPOHyvrPSFKGuKXDLPi
6ntcWA67ZVGVmHD3v1SmexJOSVfLqlVJzxT+vkwGAgAXzPaLhCksJ2JQMdDS
IeBCcwKHufZdC/sQwgh15sijTkuEN1bnxFSCSTxiqmAfpxsSis7dbT96nqG+
np30DhcXPG/mUzzUVK5xH5XTc8sIW+mZyj3dAmxd9U6e9PacFWiGk/dVnbKM
9OYJCfUGW7Savrq3y/JfZ7HDWgrpIZO0aQSdp5W0EmUb02+iE0T36kb8kUl1
974edtEapIAkq6vYUvK7txp5XdlUtJGGRjpAu9AEmy9se96IDveaQKO0AWaR
NCrRaZMkHE0qbD55xLWX80ym+oW+uop42hESrKJ8LXoZiU7lfxLsxfAzBWq+
wYxiW9zSRDjxnpMf8KkLtGl65FUEXA98+31EZ0p6mpBRo+aTzUJU5+6QwF6p
6nO1QMsd/3OeI/bpcO4xGUsYlwKhrrcSfIjRdGWteFdXlFtI/eruKt8wL2Xv
FYoaZ5iS9UaVHrjgNFq4JwjQheYI/HD2RLzE1+ZEieAEtA4RUfaOkpb1Ijom
d6AasHjOo3dnKNHZW/3Na+PclFzqeCF2eMH2x6FIDIkLg8mn3HYQBg7GGOZu
7Ek5zn9YytHqEOOxVMIe34QUvDliPO51kbvep7/P90x+RCVICh5PKaCwmWi2
cqAIa9+Vw6GMPKfLxg/25kOdujVQaN3KHfuxWKVoyNV2kWI4u6KMmXuVyBCU
gdtpR4Sq8zQqhErRtMl6UXaEgt59nRIQVBm+TBneWj/DDhDeCTCiAvCnJfFV
/G8MCdXhVNiPeMfdyWLu5lGsvv5SYQscI64hX9WlTxVNRggi2khY3uebgT+I
Lk6Ue+sigJ7l8JAykeDwnbvObZmTkiEmPvz9NaOZccvHhnZQJG9E/qG9FFD0
ppxY2Bek4F5LJ/d2c4Z5jrbMX6rz7fnLKRnvuizU8tTRmnxWgGn14UKbQ8hj
b4k9v8WNIfQxXIeItw6g+2mqYk4xrz9nJYVKNLLlrMkQx5LJsrob+5B7cp9J
gYnNrA7fp8LId4UkW4Plc3tPQP033w1WVI+/rkL18mCRvgVlKyYCCRlMp7Zp
UQyzg2ptYt9Pstro7G62bLK3p66L8GM5KaQMnpKr7wy9DmasNofCom5HVxLL
eP1sAkVIxKUzpcOg3y20594DCJRpzg5d9TPnLdevH8UeW0xrbWw+Im47RmRb
2ev00/4luj0JVBCYJ4iKJoZezsgHmKNUPCAw5kaGu77HuivkOK6YrJxl3r6b
6kkWhbY5Rapvn0CnCpef8dUJ/Y0y9Cnxx/VF41r5jVN3Tdq9Erwx7BwItk/X
naRPHIUXHLGbbwKkrzwIX3hAKIBGf+2n4k7YcD7dpWd5KD8G+z3lSvkvomPu
2ub3NaHyvMZdVAtmbWUpZdcCxkTeDZomVRGUhX6j5PGQGg8Eh8vB33BTjZUR
ZhPiFHSZ2jVo2EAifIr/exyQhW5PcV8ggKHak/ppelo00XHNY46T4rJx1xEn
1j/eY02yMg4XI1Pd3LaoFkFEwiUeTYC8Zb2kqeLrOemKa6kES3h/R3DsmjYM
+w7bb4EHJWwJ3vNjJOddu2RksPqctaB+Wvjy1u0/r1RpFdGrJvEo0sS0cc4e
xTlaps5Ot2+bKNYk53iSxiDePEdRDRs8xL7egqJjhkA2d8iuC9xJiApOZQQz
ZS3MXv/3a0XNSQR7HHCUl5hWV4Ju0r12Kr9sD/qSCbz+RSI6sQp2TLVeASit
JDoGQgo5aEV4nDyBKH8Fxn2xaHK7DC6gCyb6aD7DrbeN28mI/ZAc/7ZLmSHg
qVo/zv65+nLipYdzt0K/fZhwcanTBFVbyryeg2eWN+0XOzWqIiUQUCVm2RzJ
bBBKv5FqBYtaZN9whlEskGza94fH9nH3SLILhP8Rfpf2MtlhE0at+uoJjtX1
jRgnT/vhsJReP03sI3LGrgoomIaQ0KklDPStQxPJF2Z7FLN9K0/utlFGc1Sj
1glKl6QZvuYxEOxko359ciNh1kWx6uvkpdmo6p35MsQPsQRbIL61zDGcrfFv
3d1Dw3qhkuDx3Mt+uIrAcHj/WtOl1AI/TLKBUMat2Rw/a4UTTYmZjAoiIDSK
k1U8SCmXZ44L076QG/GqpGdhpOrTNqonYCTu+X+aNYxQJEyFnf4cmqjHHRm1
7gogcj61CsZkZNffcrtydF6qtmZA5Xee6OipGNk9j2D0VA/V/ZlklB+FsxIM
9Y7h/DGsPOddUklUhwbh9lNDK0oVj0i77w15aBmqMQyqhBNHW4wpIIa4Q68P
aSdZb31/QtaYtmzmcnwVi0BNx1SfMjdl+OIWmqY2jBJIbiBPSc2oVnEqhD2o
J/i2u1/Dqh6gx0kN8qTNcK+ya/lpxXjUBxgHeiOQna8E3iu/6YwaDw1pRW6E
HRX6pZzS4gyTq0fXb4TKBVNMBZphvRbrpEEoYN8syThtEtq2q3j1CHC/P49c
S2lJtwxRogExXyAuIxsO6crITNaS0vLhfyDdHXHstpxbqjlTBnCzOZRA6Lpn
HYaXtU2GLobVI5zFgXo0nHV94bQAhDwRvdODZJgiPi543xnA+xh9pq95g3jw
NjkOWFfHnOQ5DRhjcHhHhbeQTBbQ4v77Jy7j7SlakeXIA1JsXCjOMPXpXpyl
9/ahu96L6X+6S1Y9Io1MEJp6qqQiSC/5qd0h1zZjjuk52l9sGVrS9vr8ZpCF
y+fXMGqrj2Iah9DqWgk/W71zjdD8ObOx58rZvzo41ILkeX3HDw8MDEulOrY6
GHmjynBMh0PQs5YgAeVjY1BPSO/bFF4boUDWtQ1fNurLOoNW2LCRwbszzziH
9PDpJrWJZkpZchf/aHAXEhAK2Wk4q4BFez7e0AfjRjpzuTvTqHsRT2SQDZ1q
eWMnnVM5qpKl7GWV+iBLiDHbccVPfRcA4dt1tTIdr1/lyzVfY3u5v+jERB2i
ZRhV7vwaRdiId9iFDkGEDClKu0Z1ED1PqXji8hPnWGi+qI452vZHD7OInGjf
JFJ1QvVil6SNx+28UbizPzQynr/U/Jj6QcOwaR04uzWwe7k/cjlOjzrNDiGw
yJU7tvziDnj6Ka4xfLr2i/98n5GftrjSGRGqq20ppJNXzUq2D1sQcyATgdFK
814Eb+UpWkWFqaBYamYOB4rLIirdTrdUGbG7DqY1Ad29Gir7AXY/yz1RUb6N
4ltbMigPRrBzpE1OnJqw9pomuTzeKeObJkL+Y6ng/TZSNql31NuZHVfsPrhj
DkDJSzCvUqz3V3ZKN7HJ0/w2k0nMDmCLJM0lbqlm37uuxJuXpf5pu7LxsLlj
MHr3cUX251e/tMYoB+D5jx1IpCtnVkXF25NpJw4EE6x6R86+A1pwzazgaFLc
QR2KSeIszYM557PrTof8jPrv5r+Ux5EBz93Z6PLTXEcsZ/oXoCL6eHfrWRpJ
66tymTcew5VNMxSbrMyTg4FU7HTR2yh6kTvgy8g/wiwROrRfezUrUV/9H2Bn
Oklj5zlbeyFGDBnRQbE3/1TG5pSCvRk3nHwg6u5FHTyF3tAjFKTuBXt3ygUy
AfqVh0jR1B4vuE0m+YkHyS+R2o/8AcNM5jFW7UOgDoZ6zTouN+dvRybgjJ4G
QncZimQ6ooZZpJf03wQ6e6n+N0QNVl5UvqCXnguMWx/FT0z5dRy3aUX3X11t
HEn0jEfkJg07vLoLnlusdwJFPdHjBS4Y2J4pvIQQo8Rio+/KTlC3HF9aUrsh
g4wis5WEtOTquQViIM0FnKPika/IXLysqtkeb9WmjlQVMfeZZQsflE8EhsH7
Xe3iVdaJN2oLhVVyEd65GI0PMeE7U+SN9xdRBOcVNQXJ0pVixJCl36mlfvmg
VPYRx+ZGX0c74c1beryT/d4c9pwCw6j97m3tGuycfyOaFbInPLMfxlKY+1Ta
ZpIn+HSNActmqnhohNAoVyLthmPwlJFLrgNwItnBfv8r+VacQi3Vz/vVa6lU
fYapHR6GlvewcAih3zrJ/n8qZ3MtVci8T+WVio0VkzrER6NleE8Cf6+Gaf75
n7KKyTPlFEwGwxpmM17eFOcb60+7gbZRtFEi9SC5IUNkCbLUCHaJsKlGAGZg
u1z68sr4Eu7oMRQChdrdxiuJA/x7/o/DQXaA4dwmG9OdEunJw4Mvf6mVWaXQ
KTJ/rYY3R7iZnWPsKSPK5KDa2fxhIJMWabFWjU1MrOLO1RtKes+N9WLkgKa5
Q3ccrJAjApApejZziPUuxf36Ep/i18o2jF5EHuXskDe8NMJ0ILZy3JxQGi4/
fTgngzivjr8jm+ILQ5WeyGhvD7BU797EMopVqX5NlMyxepxFhA52oSoAgdXv
mMeo9yJKGeUexFqfXPqF2EYGhn04DiuhLh+1N9WKM6JfvmFijgbq1vEQWWk2
8b00PH6Yzo/XLIXh7/HJfQOpR3JIPqDnwfAUfvXc381F3d4ssMWJU9zpa6GC
tvzXKei3A+5oRMlRTJqBHezMJTPyKws4Q5LwME1ffTFihip0OVeqsTjTloMb
741OozcMVA322rMH4nQj+z7DtKAF7w7YIfFXR9Whcbe0R6LTktzhdSu08Q5K
pdETXyi17xY/n+Sgv37qWrvsaYi/+P6jff+AXrByzenYPMNWR6t6aolbKjwp
cxqEY1hRllTogkgW89Jmb3EuVjUPMUFa3KR1cOoQYjSV5/qsOOHDVaIdZUP0
xg6Xg7pmb3iYXD1E1TTBj7G1l1dAt4NF3Ronod+0UaFyJe1FydOf/ymDv6mK
U69r0PiLrsNdDHbXiRRep6pzb4ZEW6QHZs2u/ejMfIlXFy2HfSZzezorwZYs
yHjOzmduIshmv7eb743iW8Y9rIZUbglgxoFsGywoPd64piPa4Whsm0pBA7UV
3PZbVP6jfaV6qEnZoImYgTlsH1rd4bfV1xYn5e4XKGSe49oluxUcF09DwCl2
wTaI21KCcUxqlTz8sS6JEtdb6hvyeQFl6fmkIfTJhTExH3S4jGq1NDA7zprj
lLg9uVmu5yGiAXW5juDVu1VWeyQrQI9i13TndWfbhtB3WcpDyoYxc1UCGffP
/IL1ZMfmxtGKzJ8M5Qmh0Gyh19U75oKREYEnyqXVtGomFrMZ4iHwKa1WbFmX
RVOjCezi+4g+8JWW8kOYijVsGRI0iIVmmGF2sQ8wAxbwSiaaWJUMY6n7MABJ
EFq03/ElbLlmXO/IhbmqbJjNncT3OnYJvrPxvAXcOvd5ycgnOYgInR6f5en5
+iZBWIC0j1WpuAzloMWnXpQFlgkOm0tlicSvOXpOakLSg40xGvUW5PEHgucF
CKZ0SsM9CYxwtPNpjcdLATP/4pedM8zEGowY7/y9tp3ef3UalnGEdfPo89LA
2bJxywtFze2p9gQGWZB5C6mf1Wt7V8iQDc0ylrzVruQXZOaSRqob+CCEVvzZ
KM6td89RtXYyvZpudwyHJRe5p3/YpVd3PIHJZfFi0D4SavT60N8RbSdazf2K
d7JPpSNP2oPqIjo4z6oqtWG33kOGlearJrUJdieZ3KrbFLVH3LmkLc61TyXD
uN1fPEaeE3zCZ5jTT2A2grAR/ixuw0aUguj2YI1e2eYmo1vUxaF+P5++j84N
NXFQ0gtQpL682zR30It+5ITMhRa/fiCsCCjUFPV7Mp+HRZkSmEaVri+6gTQ6
WZSSNpWq+MZWTB5rN+K328Qw3D6p7wRnOhBK1zwa/1VueJJMHvdqHP9tSTwe
3QTVqLJoSIzpWNUUjjujaDGNhBEeKMQ9H333HUBMwU64uxFsBCRMl+xnSVTE
B+KeinkBEuVQtwgueHnIoZct5fLoAeYDNlXk53y3hvxKfjNSSCbnb31WaXjC
3nMgjyV6SWUlrVzxiI/5yOMmxQKJuTOYEO5ywYfbvUv8LuVyhJYixlUsoN2/
GMZGfJo8HqM7kuln7D0ouO5mfZz44l73lBJrz48ZgOsCOetFNVXXkwZr1Kcs
BnfJxV15u+BIXHjOyyApti4DgG3l189NnOfb/MaJjU+wwIp41I+M5v4+EN3L
HWiadOXG6XB/lENl/FeMcpx93vCi49DdPGBOix4nFXnj7elQxHUBvJQPKWjm
7VnMlwtL0MavKGpKisQIaW+SKFSHu3+82491QHALrdMjCSriSVdOe0qoBint
Jh14bTcacC/YX597clris2zYq0QOC0YSNMie/37gMi+Y1YdQMOcXKWog34uV
JUY2HSkpgrxWdPwHuHWP9yBC/pfFW/RRKvF0U2blxcmac2NSivu6qykAj/S7
qPNINeikoBAMX5VK51RWau3dUt4lY25HjlF3ji2GsYchESQkwwUposq5S19z
/Favj+ptJvwGAMj1/45XmF58XsbTOTg4PX4fGNrvXEi+fxaroVVkseiSLd/U
mT1+nn4HCocBc4ilXMqFVDCg8XQHZYNbK33rnLRKHN+LsBu7Vd8NNFjQGEMI
cRSpB+iIsSpN/FFBP1S2pZIjH/EocRWxx9g82P16h/o4G53hSdfwMAuvW4wu
UVGtiDhIW4+2hnmAUhninDk37p539/a+0wUDdLMxQ5FmZMByxKhJA4wy4pUL
SJD8Nq9U1cUIPjoCcUQHxG0nn3XvRiYj3fMiCBtOsuzcal5/MgJQCJg7vWkS
ajo8VWq41zsYggkDmg5743rIr3LsREQi0i+fH2orJ8Zt7UMNXTjK4cKMVYbM
dcpJGjQVrpffM2KJTq6b96t9GW/OFGaFaT/SlsK1QuyIApx20rF96YryBtfc
xTIHStLoOXKyQVA/aUzGU7uOjJe3al91lUmacmJ7d1cVpXfmp24JskfoYWt9
n3Llvk8RFeI+q0ywemU6cOYkj0f2IP+AqHUMS3Pkg/+RHlzi3S1Ls6idGomb
ifUuGu1aQ/8vv1Ft+CIFkCo5TfKeuFbGnJ5H4akuk8SdWvpLt4F/eoTAhyA+
n7g3oqiQ8fVoyTOMbOm+GbaMd7GcK52WZxF1h16W8RRFIFMHdbA+k5vyTezq
BbgQ0cP6MoGUVF4EVZ6Htj6H0mfOkuR5W4WXF2o81MOwYcm5B7o9vOnymYwt
UUhY+HQim3ukGRXRLWa5HFimsrkXfXtYPNrjGHDmCf+6WlcSGSQ2z+9hDz7Z
esycblyWhHHK7Xn6HVlCwo1kHiDbSM5isoF4KClRjBqmZTbRygtj1DFdxYFh
5NDz2LbiUax4NPL88yYd9kmJ3tJZVaJtTBt2D85hSJygU4KA7ruQ801DV+an
PEFe88Vs2Zrhu7VOL2MbBJTz2MvMeCMCYsObPf3IaSp9gk82MZJMtWXdC8ES
3n6sxsf1+wJObLYMrgH7aLgqLGsV7Z8JQSTNhuU/7+lPE3j13azgl+bNdqwn
G5Kavs+2VuK/obIcBuIhdIk0u1jcir6402V5EyM7WAxUV9ZVt2ZQGsHNHsUL
jHS9g3KX74yF2QtXQ9BchrvpYO/qkuTJLiS67a8GznUk3tSEQ6opB9587E+C
OmtTNew2r2JS5ndaz8GghInar8GQLU7GI5XJ2GPjyx7B9QuvIKbfQJxNv7G3
UhQnYxLTu9/djc8Q5cjp6xbI/wEjxnE3aRXyQYo0/bmzcuf2jKeKNazPjW7C
5i+FIB3Zu8mdSB6rs+wheQrauvI4qwl8jLuZM06HpdXVep7OPkRZhnpEcGvP
c37ZDCmrLMz/gyQ8lEpCfdNeKKEicCkZby4gkfWkbpVzVRi7zvqYTFdYp6cc
dBc8sUpY5YtAV/RV0EgPeia4whWzgHnDxPS+msKFLCXOC0f/MZgABFFNumwW
D/88tsLCYGMX7wBTnF/LZsY4/Fo37pU8+bHAF4SGxvD3exXZoq36dELnQwFJ
06Tk8zyVqflUPezgQ2eszptbcwfDeUJIK/xJKJA0+GAe7sfYIftmTuiPMlPL
KxxU4Lw+kRP6W4wh4HCdXxu+7z8uqdmG4y0ggqrSlmkXnAMkj3baWw8SaU2O
P0Q8+z2LDSAVR6jOxH+6re0gp8qltBmeCdbvYRKoLrtpJ9dwSJ5KoTdyLtBd
23YK/4+wKIgqKjaJutu6hqLAV1+j8EDKBSe22wHTOHz90r34VxHmiKt+o0hN
hztL/11at5rVPsitrPzNNyvzKx2Nu612uNkMXGGJbSJeZOo3dNsA+ILMW8Ve
XQp/h7MLWIqZ0bjXjDJSGpn32w6C96AoHP3T/tAAhFGSws7gf4PZ4jyZUGhy
MZSCZkcqMEKeW97KeTak7sk82mTxn4E4UfX9JNzMTqA0CQ/UdoR3tplh1pCL
/+edZtAxT/x0/KTAK506iMOarTeR+xJUl5S7jYx2D69tWsImm+aR/+oPrYye
Kl5Nx5IVhoMA7I0ZYCFCzhB/b/LZ0cwCsB+FwcHG9FI7bO0v7RMstbIvGysR
vmZYCThu+787EtBBfBWifLoi5VytGZ9QPSWMg9TqR56FOOFRLCNyYhTyuMZE
SDdq/f17XnMc0F9oij7AGNARBMd7Ja6vHvyMY1VyPPFT7Na2Pmy4W1p6pJs/
4fuI1Ymmf6+7J3okMFB4+b3p7EbJiNHFhfY/Zyw0pTQoyDz2kbVlN0GklCov
dsl9QMSRDYKC+q02JXK4JxDDiqlcu3cTtPELa9CaZWKq5pe0Hgz4EnQglS6H
OdymL51PPadTGGufPDYqL2NciLV+k19spAKu8X1j6DAWjj0W1KKoZVLhC6+L
6fDyvp5D3oURAD0L0xLQPOt9c5+i8w+FD42rvfSBd543ZSZ5U75kmfUhmc0t
we2Tpd9cOg4L8vJcuJjhtgHd2fcyP/A+TVkLnXa/fJMVbx/hwTIGIzXxqI9l
UEnYrl64eMuDLWdb6HeJhkgEGpv2Aq2ZTW/VSBNI1GTVUrtlTFvhcxDtcp3q
nTXz79eJsUUdzohsjGLzYogGqcvw97KTHEmxB2sHoh+ZiV0Q8B5rQ4D7cDa3
QzVENKjcBLnLEoi5QQwwMaDzltYwuZUeIw1VGGbl+NmDEDUuyvyPEmERxozY
C8b4SAl8xuAfA2vElwDIA3gsVOVK08x1VqYgZs1rsTQFWGavw9T3p5OaD/Gr
/TqobxB3/bLiZa1B8j7/qif0sYwpFycR57DZLQJ3m6YbuLMFlfuc2gTH/CRG
WcR1yEkXKivwN4pz9wGzmbX/jb/7KdegFpBQTwSAg8Sb0Q9o7Ni1JHmwH16X
PnFatpDuhMHtr8TNwdrKa/5+xQaYCW7kblyelup9bldGfEN08KLIZ+W2HGYj
boR8kxw4xwDxIt80gak14KpHx3rOVo+uK/MVc8atk5h158VTbwFFbfVsHbyg
HyPrFtYiAL9GvzMzCnUhtHFbnMDSLVpzFQOjxcWObS1EnfLcAI5BG7ax529v
WMfi27BhizfWjTPwggP5sDKZHWdO8J53fbY/cFEJg45Tz1A65fECqoXGbjmv
60JsqUBqOZB7NNLI4ixLxDc65TbrfuS0xPJ+yQjDoLSAFX4CUTGjFISB+VnH
c7OcMv8AAUDztpuTTJwP2EP5FBm4MdzYhxfmMvJoMTGnZWNmQC4nCC9EksUX
sKZX4FjNQfRTtb3+OPQBc7LdrEWwnUvWJREGGgebE9Oxci2iXFcuOea/Unqz
cGUE7uTezj8XzHwM4KXQRlj5Piv60Zgi0zTyqmV2scPSM5YE6nx61agqluNZ
fIKIHtW40VvEroVRiPYdNKP/KQXeGQQCfwicpDSybSPst1BdCo+C+5hyToui
wJCBJZsO+D0R3lV6RFvz/mheBemeQaTfDs/lTjg4Kdaggynm6/DRmXireqev
Ttik0Ynw1GjhvWrlYbWbxeXthgTDUQgPphTEQA1Em4lGjKNFPJ60ZJrq/NOz
Hgz1aOsCF/FDOrnSrIqbgaDvekKobj8zMUHE7xkB1B5fqWFxiQsitfa2iL+K
Hv6go17CrUYmixOdiyx/7EkEFr/GXTdli7qnrqrWOThyqNQVxNjLCUxVcETy
DUBzaYN+A3iArbFbQWk7PfDLhc8mpYwM5m1ewt1HUAEFN2TDOOKPW2wK2B/t
DNz0jO79X8sbFyAn+VgdhIfUIj1XcUZGiOokQVrdWyN10vFqKmI7pas1oDb2
gbFf+wgWKgefxTm9EwyCvW4cJDxB24Pt4hpdPzAyI1jn8VOLvvIhaX3e1Pbs
cf3cv4/r1K60me1UlMEb/mQnSHzUaMNko5Fpn0fi54JjSpMm0hqo1KSqn/mt
L2L/8yunRfOw2jko+0b37o+VWkQeCNchmbVgP2OegLACnfV72V4js541YO4Q
lJAsFgW5fYkhinMEDxrX/36YMRMkuS1H0Ad9i/lvJMAk78jM96iR957pgH4o
SEyND4SGvTF8d7DGwUzZ0AqlmYOPgLKrHEGbF/vqus5xbnESJB15mFrOpaS1
aJrSjQeJpGLZVfuUO3TrAUWyyYuCI/Lf4bQGw6tunFRulDD9/bh8Vr8aliMQ
N00JVtBeEzcfsfxQU76ZpMcVG5ntkcAgMt4/angLTcCNVHAqtWY0ynifjtDi
drdmDXOf0jbNVWX81AL8h88GvVyadj52R6RSPYNXdYL3h7hHiGxTkqh+omtS
CPgyVaJS58H8XP4JxMk2GcTFjmKhIjPWIvu430bMLQcPzIdMwejVx02HzmXx
yxepXeZM2UsHPFq04aWJPfE/kZEoc4J24IPKnRYeEQz+XYZ3pRrIDPlwHWkv
Kp34bW+CTzVUnbEyquNSHjRZ+RO9xp4EzWkJk+3lglAr2O93HM0NBvt0CTsh
jushAsp9g8he8FlGwxDJchKKrIh4PumQBtmXyt9RXr5zYHvh0jUi8BaaPFwv
C9exhxgtxkZckH9rUgDy0SO6qNVqyrua5agYMbqOZec5/Idqd6sTNKKnTp3V
iCK9kwxi5PdEG/CCvmEFRtGUUvzmxG2tX7YJA5C5+6KXFoDhkam5thdAX6LF
c/dlmm2poIu1JXDWk7JmseW5IdRC+JaI89HuBbIFJ7FE6T+1TQQJhYkNQQks
M4CscZ/glTLUYd2ONTaGmUMBvAgDwwjqxQkdKRNfmoy3vhww/q81isRdIKVO
lRkS/tNCecRSfuoBY66tcnuPVw5PSPZrFT1xGvxpJ214aoI7JiFXK4Sa5v9j
WkS8zp8AlUlUB8tGCr4KKXxfxGMNCsbSgHfh3JxKbw5R+C+nm+fWS3FI81E9
QngXn7cDZpXVO6+SwQ1T2EaY5f2911CW9J+sATrw9wwKYGshrgzgI+P+lN2/
0DLNKScaMvvFjnVFVwvKRi6ttdvw+45wV8pzJke7GzymcPkWCMDepPIl44/5
ZY3XDsX4pewWJVANh3lRoJ8cB43XczmCdo8GxJffdhXn3k5ORiyyBnGSRVm/
kZH2VfFwkSo9T9UeGww68uhSxNbrE7MbNXSrmq4SLUYOx3acLs0WBXemOtOx
1PYDHeLZdO4dyaiJMzIDgII2Rv2ldbFIwAluUmX0e9ncMm+oB+K/sKbJ0VkU
Qri8YSxpZOrdYVQZujWbhKJJ9Q5FmKMf6APFg2/Y+xwzLZURhQ0bcHSg9xGE
JZioxdHp432R8aXorEukFqBc2xTr+1m6GycwH26VowXPkZyNc0TyGpsymXit
/j151ahOAf5aCmjY0uHZEAU/rK7MGWgekg1mUDT1LnblDSF3Jt6fpot8sqRS
+nFybTYhUA3gW7004+2GSDfeSh1sdxrDA3jQbzmavN/lL+JE0+/woo7er38V
UxUujrATlpK2ck/xfryeGzFcsipiF5ntzFOhHUnWDekCo4ZHaR89IYpGCLsa
I8b6grFaBnv+KBC9iGZKJNoWDzCsKvOa/sfclYaPpXUXrFLwHBBNZWeGCcw8
j5fIhpA62YotZY0b/KiFdFumzCWHDAmIqsLuiLF4Vlyyc8poQzlmSBpgmv/R
RKNfOQLFlWxPOClQgtghvHKq8SpIQD+5xpwIhy0RtZ+N21OEPq+T7PydUhK2
0FO+numW0pb/RZc+3w+1CR1aQhsHo30l87NFHKGN4kEURmXJyGO3QDnde0Rw
PxemnOnb45lmueEXm8QuHJFcYfana/FpMt9FLPzRrellPuEthtTV/2bwiRRz
JKhZXJxFI50zzI1EAiuFTaDwd6DLo0WNIEBTrszD2eHdRvaBBcHtsYjv3qC+
DEegc5yJpRxMuA2flM/nLHVd53+9tvVQyaQRoOe5W5K8KFFrPNfUm1OLRFos
tIfTYnyy2hwdE5TLE7Fpw5Pu0TDDZ/sWYl+cqjCwnhVKMZR+mqQZw627m1Qo
TACYlk0jBuRXyFlW4pfi9ZnioVQXoAhU7PlBLtrA62zLAnLNghNCRsW74usJ
kQCZDxeI6eKzOlg47f2IxHwQwpjEyicfNJTMZXS+A1t4izbFHRPisXz644Gl
pokszNECk9yHlFLfacCiLGgyMURX/RnwM71UL6UBz5JghMHR4QzyWTIrn1D5
IFcy8ZuKZtuo0RM07OC+f0MQTev6/IW+UMq3nnoQD3E2UHeoKicvDJUlkDAd
a8eRd1RHimPTjqT4636kydw27ErFhW1IU5YSPRh0nXJDIx8FxEVHXkzhnZ8i
4ead50MSRzOfN+JCIsjOFyOgIlmmbEdesuzvHa1V8rn8MWA3CPFZF90Q8mMH
7e4hHr9bGDW+OuXVurr3m3uNwPr+oghXnZ/oMnuaVCFDXetm5uL7gQiDCzau
Bo6pLzHidL2JV6MNnPGqe+X28akDYuRw6RZq/dl0BU4kWoPHDzEz59kOC/gA
xT4l1vtQy19gG6jNT9090pRqvikTCTwKa10Hr6t6MSOLpPptD0NUvswrBV5F
zb06cV3SP2IQ26xo1p3aL9I3xyOGSuFgNkSwvWNUksIfHhI4NgkBrfy5Fxho
M06YwMiGKlrxqgUqoZA7EdcKovbB2uLw5jWhVZNSpjROdUyfXkWr4rZw4Pzd
JHYFi21vjC/O0xSboZNRfkV4cXASK42m+Trnik5Vzs/kaqSgLdmVKnfrKoYY
dPah7ikqQ2chlBLf075cwOCD6OY2mno1hA/MnAmCzsR1Qk1TTZwbOu9IqPlb
iVDrWOJxqFojOuloZWdwZpFT9jVTTWtRXXGkoBxEWWmmCKtIW3CCAFwOQTXm
4XCVU4gGqs6vlazerTNSMyTy765zavFGeXXZGkWMshdPEtRqvXZFYGQMal1E
4qmZZUM5msepvZ0msB8XKxvPYn3yamcWEavKh8Xh0Zv+KjyRrt0lAdS1K0Jg
4TZUM+VNJz3/UWhkH8N238wZewChjxIsux5TScmthmxfsXHYPKJj1VhOtx/Y
9tBex11fwFKs51Q/LrLTRGhxwI5+nrHvBoHK0ai6QLWWXP40cZBuO1PaE+Dv
wD8YlRXlXSHzb5gH7eE3p1lRK+unoQZa/1QteW/uJ+gFX06sKF9PhDtWKWzu
eYKhnLBQAE6TFDXRDo8TtVDBCKnvOtCXK0TE5IH7XGPVDUYc0BnmdefizDk1
7npke2EhwEkpqT1n+zvgYg2flwM4Y7okZjay94Vda5XPVRUxMD2nRgyZhTqf
xabn4I5MvFjIucoNmecC52Tqn0YL6x0NNz8Ms10zc4hEf4Six3W44UFb/87q
jgc3HppvH4y7xs+lSCQYSQuj9klLAkk1lMwXQV3fzGBx+85nSr7PtO8tbgQH
hAMp+Y5MKXoC3U38gpNp7LdFOg7MftTfL21GGV//1DKAemob0LbLWJG5l1qf
0FyzXAkrhWVMaj7M11TF2QlPe/Zcg4l/hkhkfkvEy+vTpdM5LW9bJYT5nP+F
uVgUIdW+ewPlXWpYEwnFjjNi1RorLI/tLK/5R2J5nkqUVPHxluw5oCOZ0zca
Uo+l5j66VHZ3OAyNyyerbJRsxwC1ueveX9naACpXFNXL3+7Z5IwyKWoEVqQF
DRyZqxI3+fBznDqV5NlQxxydWIr0AxvWugd6rVuY8PPqlRkGWr0LbhtlwkgY
uZhItfOM1+Q8baiv6g+wV5WB6pKC67fRDg4q84Z3b/cx5HIOVajDcBhm6pJz
ocd/sKs2wLHy6+dVCMAuFqUtWx9CJIsfLRH/bhtDuw9QmL74PGUbrUvkTvwG
Im94TJzkKF6Ylio5WraldgtfjS6fYdSDn30cCSwcIoZg3ewxY3moUo8/FxJw
+TA7u9em8Xb7qkrzNlc6Ol/ARcHzqIAiXqaZ5SCtPJXUFMqPjF3PXXkT/0Tv
WOHdZncMb8Jn2BjHNLGCSerTq0TYseNiEqp8sKUx03AOzNkDHcpSGGeA24Vo
KBlrOvgqN4w18DfAQsULkFTwx1EctbN7ThjTKW883SAnoCcnL5gQy9jQ2uJi
qMXA2BF7sER9pNKCtE2+QgOzIp6xo8xMrymP0vxkOK8LeS2NCpL2vroUCM0T
esXagvlaGcUVG0MnR4akPddpSnIernF7LBHi6l18VQrM/5m2PdtDunbeE+XZ
u1u0/UAcvjT5SReDuUziJhZLHXnMUftIgArbq8j7bfJ4TojVcxVvSVe/Nb0/
j7Bjsmi25bbOg0pJFdMJ1Nla+bonBXaBZKTwu6xcq0myFglWAWRo01L524+n
mf6OZm2KO4bWNu4K74Ow2FRHrJGIPrzeI+nTleKEJ5eLOlXDTBkfG8R+B9g8
2yk0Ew8voF7aAYFqUSnrN+5DVHJy6lKBRX4E/krUZ9Ih1hZil8ZvpwdHbHx5
1yoekgVTyWxBCqywhBf6i5czp+9txN34wUx93Piw5/MmxA+cZUrdolUNrh/e
hypYNP55XzNOIGwAhmrjKAscJdZL7wLvnJOY2kYFxquGPW3fWquGacTZD6qD
yld2ATu589zOUTxKwk0S0i8kKrcKRSDXVw2gfx2cXb5VFODjaEYcqHmoULoX
7LB5m2vrvGVb5gGz6yfA76YvbnwAU8jYL6EU5bI/t1avigWXAC/zxevuMKY3
mqaH4CCNV10YnZxhapnm2Az/pFNS47rPphR/TkcpYuFuIgYNRAouBYboYxGv
d8Ayra6E/bTdymDOVt9T7LHL34ePCd1cF7g48UMe5M9KcLsbowPMcp1t4tme
b9thJrqn2OnYLOil33y1MnHIwU953gnw6cui25GCc7efa0d6SSM46z4iTvG1
HDEOfde48QVFFNKNm/Hj4YTChlvbF9A7fDd5yipUR/Hp4bwoV1xg3xyWIiZh
Avp5QH5fgkVCP+fut2QiJg/bcGGH40G5ZV8VHY2ujJvVEnVB2lGYp7D15BbK
/NThoRTuFqqkqCfb1uxJGLNcgNWgd4RDFOYb7lp6A6I0qK9fRRKp0EigJwUH
MDFMCKN+jZqwjmXuzAOPDVHTrNmX51b9BkxOnulh6tI9QKyYVxB1Dm6xT6ye
bx4LslulKR9Q4JixMdPDZXDRuGWPvfc1GfD4dN6ET/PCPWzejSHy5jHESrO3
MdrSmBRPlyn3o6//XlVN0+h2Pijmsg1qMdn86qVkW8LAeigrMmrc9/R5lH3J
Z5AF7aMI1YkPWzQo/JJ+DKIwWt7wJJknVraO0oocRbd3zhkHFwq/GvZZCj+2
q8eNrt93LDm2ba8S3a/k5WumtPHKnZ6gnk3hJni7MsISNn/MC0g9yhBGCcOq
rqid01jlDAbNS9Nj6RfqBd/buQewZOfq3si5jLxDmWCR/aQeJXiiUn9i2bdM
Aaqa9n4C7brHm5tL0cPDJh/YZFzrrO9q73id55ibGk71+vXjBU8Sxnupl0Nh
qXVbL/+ysbB2hMHsY+Syu04Gvpsm39FRXD6RMdJwSJSy9DJ4+tpX6FT6cZSL
KtQ353ibMZnmiq2kvYe3pKxR0pS/DtIvXluPdzRDq/gMvs7A/FCtCOYtzdet
PoDqVT8W3ekrrQ41/+oPS1D/uHUwS60b62XeR9l3x9R6Xy9fIpOp1NfDGXWa
FpFtE3V6Ho+FuMdg2EA2NZRfpbfl218ttivLZYyKRAdhKHwEiUi6oSaX2iGx
r7ad4vi2LogDKMVH7v9oBfEWTDV61aq8xGasuUG+ONVure/CvCH4moTv6k9Y
pcRt4HsVhim5Qg4SaTu5VvvXv045DA3/fFp+7/BKQT5U1730p7T1r9/EXnog
YYLiyeZ5KapT2pIFUCj8wQc7PXhjvoJQy51AMsoaAX7p62gEGF4iGCQvlnO2
klw+YTnnwVkkggGibIF/jI/ru0ae/sSXDxmuqagziNbUdTcE4cVWjDRhRXGI
3DxEjnqqXIgj4FEwYMnUwVRHXP62be3FHsVs/sQBiIiHN4uPFNLFsWr+2mOn
jKqFT6ne+WlvXkJ1ChbYuC8nXuztW6EycyolGGg9wpVxMkKpPuGj8cdOV5kf
f4FIR2emJ+cLF+pcd+/s8AV7j4o5THyQZ9MWQpCbJ3EsTVwNnpgYGnYK9ize
iyc49JXDMVpQP2Luy+3buVUNm8dwj7DzYDd3/kBA+FHF31AIC57YMz/Gkyad
NgxkvbI6CoBAOxmFppbMZsM6D73ych5di6VSWKqaLQCKyqNuQVnwMiOcPAcg
Fwyw4e9oZXXiQ96grhTu04SsosQbcEf2pF6NF28yNLJYdE/Qyj7jocjHWKk1
E5ljD7kr1miyhucJddpUDItTmPaMDm+5/1czum6z20l58u8GrSRnU4KSgx7C
SeL5TZ3szZ9aCXJeNHhLhLHwYTgGOLxrbdpW4iOZZ3Iwwyyhfp3yYlu6ZQuD
jtAylWBlEnOzCWo5oj4sFknFsrJJLDphHH+sCo8atNT/Qo9XKY9lIVgwBTq9
i6Yc5e+c/JMp1/Dylfv8e03IcaCHpDgqVkUUXwYcnx5NvKiIKDqtqJ0+XklH
ED8J1oQzq43Rp30ei7hetqjFIWpvJsEh7QjTfwk2q2Zl4b4bLFRu3JR53CNl
kvSKtErWwrZIznzmkee5oPv27WzwJ+Ss5v9mYtKO1tGiXNwJrUSuhaZC6O97
06sU6nAecLEQA6peDzCnNFJwJ1FWYcFVMMxbYK1/f53xjtW7wph6qcsnO1c8
6gBR6UWQJ4mEJeSpRuJzXz8rgiksVbP+MKYE4ew4WdndEBsiD6fMffhpJdfm
qXUyJleKNtnQV6QAuRjNOQjR6iBSsajcpIzL2Fb2qO+JvZwW3yqv2aLiQhxc
YUpiY4qHZL9MG7r1zDFl7MnaPxXttQNkihxvwxLOvkGJxTu2wjCMKzI8PBIY
Kh+x/aJbKDfewKiA6/RtXonh4YPTUJliFEVqXKESPoHT7fD9G1Sg1Ub94/mx
RRVjrhxRfaTVXCS2Gz+63q/3RZgS5X0JiULWi2HkVBDAq4VAwZiUj4uGCCym
BdHU7dBRCz/rJwGO/9/LDeBePBTVREWrG/AUpiU/sj2AH7gfAJcPTXktNU5/
JmOqLTauRleEqbNd5YQ4vXxhFW3Hj5gV3mStP8IPKHu36izNNQe5ZZyyaiJp
VkaSuXmBMkCIH87m2G3oviHlUGcPJh+aKDGgJeV5KaUcG5PWvEoiFHv6F6dA
JCpXFAsueZ9kEp+F75Fpp79uzj/oBUafmk6e0uIJFn9IwRzgA3MvTtbr25W6
GUfRYWKf/gOUT8Qp+JTj/AhSf8ocvff15EU9vBY8/BWg6DaeG8HHi5e9h2H4
UV8gxI8kIT5ACU5gA2cl6JtwEG/zxtaYp4zgRe3TpJHafhl/+NImQp97+Gt1
+5/YnTJLQ3eO4joUIlvgoDlno+zwYqPkBYzWinl7xiLbeY1orSL3uvAKGeCk
fbSgTa4WJiMoq9Ox+aKfkciZaJDTbZYP0SEUvv+K2w3+wICHsX0HhlyIwQxS
Pwv2tynQUVtg5dVKs3shbKFSVbGpaVxvNWBeifdnKrFXkjb4HguwPD59S30B
dcfQGfD+aw4zRq8VeISUPDl3CY1w6HkpYFul9QUaVTueWYfU/8ngRCY9va6C
6mreX5ipon5+nSHLcYULI7ni5SmFsqFw4HmuD3CVQwIhjYucZpUqnLounE1n
9gcOzP11ngOEAadgZl/pmSIfYCE38SACf7igF72/wZuAvLvbJSDt5Q2BEpCY
jJ/EYdsmgsAUlZoagn9y58y7HZOnXvCZduprO6XId32P7XxteJNKH3mm2ydv
m/7lIxYo4z0Z6yUbiy6H+e6wC4fXWF7K7IUjwNid5UqAC4XOqUtT3gP58itR
EhBhYShxx6YFu+wkb6c6/o3ohOQbL2+pn8nm74gOqhZ0z/YGXFJQXVtoTpON
mkRdiwMHV1ddWdTiTvrY1xzlXf2cVVlDM6N8GPks1AzfAeYXkzEFqB94/aP0
qkJFTsofdLMVHR4efnGlnGTPVI8HlwzG4DNBStBpgEJmGqhNLMs4GcNc2ovv
a0f4UpmgPTrrA5YtnyI2dzbBxicLPW2p4+tdjivHwh54pZUETGzb0cb/dpk1
hkqcM0holjLpIG2OUi4Me1JkMlA6E3NCqe+f37iHocVhOkwWmB+W2FuKUp5G
9WLJIo1bw5GPrcC0cl1x2peXsvV+zqUFtaYTg0wMVIm02zw6gi8Y7PNxvYzV
fG/MoTAJhSCBNE0DWyaqYenI7laDgc0kwUrcCJDKDqvIm73mCsDgTjy11DuH
wwM3nPr0hza8O/5cstO4enqxvsO0h8ZT55vPElcYZtlvfVFGRXtGdWb+gTPC
LgDLRqzFM+/p4ttjdLbS+qmkXLjv6tt6//OU5BoF50oQLBqzoAQMczrTy4xe
mM3OO6DqBgO5+ZthmUZj8CM425wYgXXsM104XPUDMeaV3HLINxGKPHL0Gn5S
2rChK/tGi1JTjHZymgATUyYMBJG9h89U32xIQVFrtx2XKn2JjThJjktXGSvS
9TQ4XIZ1cJylrEaThMLhE+ekFX1uQKHccfLwiFpovJ+O+tfaY4U8d159ThV6
bnu+09TtIKrGxfqOVNKshG9MSDHUsI6e+xqL/FeCStK/UFzAfiHCcCAfbiWX
59NLDgy9/LcWbj6bTKOsOvt/IgktmqjgDTk3Glk6MEbUcIAFtM8iRvdQSHhi
qgcxv4EX+27Rbksxk6sYfnRQF9FVNkeSzyWOczwJM189dXttXBJtbBEKezNT
Haib5oHDGO79OTU2JJ/R5m2PamjRWXVWq1sly3NBV/VIB4WNZ7U5a6aaqUUC
RK8tY6+IqRAvqwFILT+IeMKHzwB+3h0ezZcffIP4CVhGAa7VDs+w0IsNpOvx
+19fqMpKoeFDjU7gxs/+5ZdSWufA63FB8Twz48z0in3JN3/veKp1yqh5SME3
bhHnEM2r2Fu06ag3nMp5x9f5Q/Y12pix9/dXMHj4NYNZrljl5HnDfYLIJ8rC
9DD6+fH3bVvfSrPS39FRhopeFW8vLYvGewPPTNPpUQG5bF7PmVgvzcyk4kcQ
AZtsKOFo2X9VPi0z8rMP+KhQqZBQ3yPIhWZUeZck/4PV6yO1rYZgaY9HmTPw
o6ybm5gm3nZ69Iwzcr9H42Xb+PoEpoUCzqnI8QJexZArPXevj1CWbMVfclSq
a8usrQHFtR15UYUBDb3hfKvqnp4s1dPYikJbhl96ZJQ2iawhVStw/jOsyPXg
9GrWOinuVPFRCvKvHW3/3IROYpc3WfV/6tvQJAI0LcoWCzka4797xzaXOdkl
lFcid2Qj7m/hHzIfyHQh7OzB8ppky7ty/sTLn7/sqCSyvuLk77vUltpIWNRq
Lnb6Y42W9/VTdxkv3qaChNkQhcMZPsJaoQIp/gCYL3wbNXAN0a+ALsxFjmzA
YC2LztO/3OS0GKhWQw8KvMNyWDeEXqTiDWbkvTV+axal+JxHNbG+C0w4QEhX
X6bD/cnN+s85qv7PBCsKTpdf/IQngyO/O9sufuyKZ+6ZqpMXbjgAtX8XcJpV
KNI9YUZhkk9Babks3NPshxfyBVs0F8HSoxd0fQqIoOaTeGF/v7nQ334hz86C
CYaKjkzdy1HawGTGdzDHwuyD3U5tVAWVs1AxehFGJJS5gaH2vvu7kpOkpiNA
qNrcvzN1e13mM1Q2o0L2WdSuOlsneZZyn790wdnC0iiLCleEE+huGiVFpJkq
N4T+xCFoNcRfJfQ0IYQY29S8mrqaEBBvQjQn3Efw+nH1HgcZIJNnCu+M8Lou
6pZXqhZek0/UYKaFaSaWV6laTI5OIs7E0NWiejQ+7s8iyFNCDwGXjY8+hsnx
zlZjIzRQCfqkAQCdR/+TWZ350Ow8C8EdxM0YC4QhJ5b0gLznaOZE6oZxpTOL
XViStzIfrn47qYVxBYpDUCq2pLk/lZNSG7rvhDlmlt1LCEKBA1mnrR7R0W1a
NsNTE59QC4dMCVnKUgehwpPzQHyL7OmFoekbEqh/IPNCYgrCAZxEFW33E59/
/qxEsJM8z/lRs4x/BOvPxLS9eT6OS7WmIA/dZOpMDvOscwlaYOOTXZ0KfxdL
3MZkbiErWs2HxT+woUYbWz6wa24U49I4SG5aXKkolau/fydTggh1AIKQqNcZ
55jOj51TpRN5tzKUbC/FrwHoGXt9tQ+czdWvrnGzmPFSl7bzN6Y+zxQNQuy3
5zKc3Vof7TfT4vxVPrr2iSbHdMxNWf4tKivn1rSYeil3FAaGuxdoxFpgJ1RP
OcZh+K3aYpiLC6N3WhpdrPK/FMj7wmC5+S2/jCOZ34MhRBWt+Kli/Su2UBaC
zPKt0AuNWHTzcmzqypAPLSfOS+3/WWu3nxFBT3DxSZ2Z5wDSJRAAfJiW3ql1
HrJm8ENfPl8RWrCSUwXVhIK+Rkb4AtNJhO2J3+4d+mBOlk//AwwLDnSGJbKI
7q1CG1bwIb7brMbnjYIzkaYVyVzw90tWjUik6ApAny1FOtAzX4lYylAhPPhS
oHRjDM9Fd2QfL25PXE9BA/J36SG2EjzyqOMfX1Yx+TAsfH8BBcSwepxmccjd
DOZpWFHwEZn9mhXGCFe1P7YlsJmlV8foJe4FIDpPgO356kwQ7NY+/k8nsrfd
03tSGb4iu/9xcG14MaBxJz+iMckPLCTyiUZfMoXm+nxBXmZCAUWQ4otu+odK
O1H5lR0EpCIr28XZHh3Yzo9+73h46qn8iQ73OlgBttCklnXPef2+7BROjbcO
vf9/uBxyu742ScSu+cSvbw1rQlly382gmJWkVpKuef7W+m1tU7K4Nx1l1Uh2
4wHwTHvDqDTAMpyNCP88bkc9uEuYhbo3521h5COHcsn03oxND0DnSnfAyrzY
UjzL2o7r6HccprQYRvdS3VHa9Mnthf9h+aHnhmVZlvQTN5s8brfG44qrJaDz
lpYv8tWimJRVrwoKsNXBK916JZrAE1FlztSAFbmpjAZOzYFFZZbCJjRXclGj
5Bgmuej+R236ECbBLiCo9M2qSxyoX0uodjh29c6LXrZbLH49yuJaMFBAAUMN
FFo8HgzsQo11oiTVVbQ4c64xk6If9wSibb1wf/3mS+mdPeFMHQS8Dvg+UGUl
Rkx5elG6iyckkmqnuuvgxAvbx4wJdeGL082XyuZKhLBPkEr/94fNAvlyjeHl
9zw55mUaj0PUyjFYp71aRb/PG1diwHyH0vYRrr8D7TTbuevolxgQ5wPKzDCz
1OxozG/5Jrg+kwKIUZxiUc1H+rsmLghE/Yj0Wx17IQrRs2jtMFK6ST7xIMee
Cgn1VtJW6l3y3DKUAO/QkLQOcUdL7qLYXlx7EhjbGOlbN0v3DpDQAvQFhCHP
zQ0OzHKPMEZS9gm77ht5LwhFeSdS+jF/yue0YMa9rGRLisE0XSKNefnEDt4W
ldDXTrmmUaXoOqHR+2wGgx9RZ/xPnSykpwYxVW7ok1mdw4ytl8AC5+CYDnpM
zhzxy4+SCQ4Z3mQbeCfTyfKQYd23MRYA4KMNN3dE3pb/CDMPW28Ywv1yjcj1
b9t9CaZFY0yR1qUhHWXVjdCzMPmuzB9Xdhj0RgNwYd/XNBhLm4lzcWKNlnTe
j6zmNl9Yri6GqAvo4oNJF/G1OFFWswtArmKXefYVrbxi0lXSWvS+mo4e5udZ
bEOspKcde545v9fWvtyY2KY9hFGb0heGvxrxTDCCp2J0Puq5DD6Q/3saeiwz
6xKbEd7Uh94XYFZ3rPqPZPV2KPTakWslJT5JzMfs9mhP8AHo25Yped65snEj
5OqsOXyjfASkWOGpTmEjnGeqldcMIXsBKIqNHK8jEVjCUvzg5uwk2IoynNE6
Eom6eLcWTXKClyvpdnhURLxHf/LDYsgRk8R/4LQI92A+YKTJ5zcLZJkzZvJZ
Is8cUYc3m9peyGnS0bMJk5SMRGGORw9Z5aVWu8SmqQb36ypCOLwLsv2MxBrc
o7MUQFtVuICWR5XsPsmDCfprYmRLfTtFzHOlOHqIa4nNLiw8mxKrNALSn3oK
5xMw/7NBLCJg5HTEREtU6rFAV67cAAr7yyKzDsDudz9ZK88Z5v90lCGfQwkS
Q1YTJxMnd369wMwQr7bF7LACEGqdvwRCwg8pEmjd4u/rLbR5A6HwqnivRVBf
GoPQ69FzYr6exmbe1FhIzIFkOLkGloxj/rXhF/M4c9yHTGg60N8ZWAGDurvQ
uglN0GcsSlVshsleKq7lh8gpB87l15iAW8E6mrqExJhqMoLXjOIpxeZGulQq
lQ5jj4fx1fNmRgGNQd5dV5uR4iDE1YNZh9/ahlhHYSi8UCK7iS82fuQzkpWP
R2u0BPccRUe313vLElLUZUNnQU14LYXLKsCXUZBZTnCQ92fNwUHRVXptoH+x
7RnmCIrlZfjr462WYbSu0TYFNtPHdl7kmg23iOyiJD2S5mgT9rSHwilelxm3
CsCtb/Thvj2BKyQzYg3uYTBMB8Kw0AYhKVviY4cJ6XmKsFmGySXteY4UgK9X
fyiCqat6jPX0IhDlIwoHtI2ZwvpfefjZedzEeE2mMQIhfNp5MCV0Fsahwofh
5CgSbWMFnOQ33+DGIRe2kHKRLc2cF5NJO/2+lWt8fIvHeNLo45ktW9ABaoPd
/hl8721wXOY2j96w3VSVYjGgUtZ/V+akGhZPcouMnb5jhJ2dyAYx8LYtjQBP
GKx7I5t9qDJOQjzccEP7/lwEEyyDxSn2RSrOeNaZFO0bYFRokrC/lCZvhI3m
3aOWDWb4i85LHTCK1gcGi1jTxAeQMFuoV5d2rLj8UFrjvc5k6E8Owu0FF98f
e9A57pMScs6yhPaMxEdTDVxEqE2q+nd4/N2TJX76oMLX1ZeF0HLpPjVcF/co
WAM5jtg9/YfW7md1nJyLO/T8L4yDwD+Q6v+zRWX2yuLoVmsBUEltO3rboaFp
i+1e5g0ZrTQ8rYUA386FgsR8xACnF77Wojbk87ZhkHLUr/IWD4kgwSAcUWdO
1qQ921fb7p7dLKfWAkoK8x49cDlWFyyo70Ebjv0s342ahxRnqn8NXs/LD6vr
75M4yJUQ01Yarj3VzNkxC4fReK96AIUmqh58zIfokCDakc4rNJjy0CTHurtK
L+0lnL5qbOKj41eYFTef+q5w9c8VNsOOO81GcFAL1hSODPAG0Tn5NsVxTWHF
xSqmCsspJ35kp/Lc6AWNCD1OO0ncz/XcfC+mtlddwF8UX8bgKLa6zke7YBhV
aMu0MYD9XofDKmg865JKraNckESLUvD4zvxDbAM4OSoZe71Vh/ijKJxI4A+R
jk3jivWwawQ3luD9cGBJJGkvPPDBdADy3KD7QT8QyFcI8TyRmS0xZGXTW8uh
+2UOCdjB81vXXdUJbnXzyYKyuVuw+Av7G3uHEQEbveYecENAIsPeGTOuvBYF
aR4m3tE9K7tSAA+WbLWHfS9XUzjWf5p9A1o9dD6uiWG0jgpnR0b/QEQyf4/P
o3+LTsxmTtm+fWb/IQBDdmuciSstzrtV5jJyw0n5WvsJUsff5MpFpuTdA4Gt
5knoO2/Qcbs+rfGzPTpaaNKdgTrkyX01mwVjSqHKbcdMDBvQuFbIvg25LXaQ
7uw6m0juelzAR/O9tJ3iKA/g8h5yLXFJob6aCabzXEiJhgaxHoy6RwA5Mmzu
cFasaCQu07EPxoh7VIcAUqJVxmxPcpPzOE8zg+oihtgrfdiEM7OqecwT8aZQ
8EalWVbX+y7eUdKKGNSrqKVRghYfRtsbQ+GFkV6JB4MqyNWJc6L1wXGZvjQZ
P5GfunPXjdCMjY/6iMu3v+jSJyhOQTFe2NFekRlnbGWM9rP6pLSN4yeMIdSm
Vxamq9bMeb5o9nDiW4rjHpyD7zPrmqFeDtNqHFkSfLpWYRpwdeyrABxOb16Q
isRpoFqQAOwzRZuXK/mWExoOmY44rTxhKRjFWYEifbxkD4bfSs2Cd2Riifmt
fik3AGTCNvo+GZqEFn43Vxr8u35oiQUfTMtgjDEaHKFSsy77riyi+mH765cJ
B+31M0Ql2GffVTkRiZs0lMdVrrS94FkgrQdGO6uTr7UMeH4wQ855FXT9Kabr
dQgjDfNwf+mxttgDCZA/bwuHSljDV5/vQrCBYSJqy3EYSHWLThS2bosHSCF8
S7wbupAsN9PZ7uYo7aYY+v9LBB4q2h6gsXTQuQsXwL72Bq8WIktqYAlvXJil
KIuaT01Y/EY2l/y1P4sFrMfAzhnrG6c9697EFf387QQssRzrZN2V+zGzO7Gk
rREz8ZX9uY2VAB1Djynp9bFy15aMQFQzn/F0V02jrWVZoQgsVKGHm5Og44A6
3FU5gJT6T7rblcgfPTSz40Pa+3SmSvKFen/GjQ5h/81XkY1gKFJskAd2qJL+
hKjMPCehZd6iQoSADq568vr5YU+MAcBQYjjWaCVnmlX0igBG+quPle+VlOiM
ev6/iBeRLMAYyfNAnV1dV6X//UIPRowtyJmRxfCeCFQ9VVYCPHImo7SpYVNn
75K0YmZ2ydHv+sNaHvkJZWXfjnCKCYu3P+kQqQz7j9Vuz+sWIcOAV9Yhgkah
HRtKNh6pAwE3u/K3C+cyqPp92XCkPrduCEZMZVkC+x8rzQMBdGdJm4SMQAXT
PeAOqhA7E4V6mi0B88AwrSTpEQdl1R4daU0JYmt4WN5XSKCKwrevYAa3q/Ue
3dkLHdJrtUfTcIA025Jsj9UyGKnbL/iVx47xduVAi8IdnL/8pjwLqwkgaGOZ
75tqmuHA3RBzPzbiDuQJaxUPYzlo9LgiTu+29L063PHkAl6WQITXgAwTD1eH
UCQEKBET3rtAxftCovXK86u2Dtjki8npoOaDRmekbuloVWiUnG9KIAhAcZdd
uUa+YUY58aEMOur1HXQQwATpuAfaSHluhgkC1a5UpG30h9eFObRNcA2smiIs
UwOVmTANV1xJalUtBdGLPGOYLY7oixA71hbzhpqgqfeld2y00LWj+SLMjDvD
bxE8MIJXfisIfG9JM562lZH4utkzmOPgu+iObakdOLDK9zAEQIPsTFC6DdU1
kKUYXaXPraaK4NL06tfoaStSW8XGFV1FH8cbQa/8XQVFqJ5QsqNVDjHhnuyr
X3GO6hQ6xXMoVbK+XceOLSYUEg69Btd2C2zmcMQZRY+usZ2JLrSQ0A4GpAAK
pgHuZONG7GyMq+/Kh1XQGNAY0oaVvCb0qPSopZzJeX3drA0UvYaFmPjtiW99
JPkluZA8lWkT38oYtCAVsKwHczloKhLxON3wCH4O8uIcmNAwGHEmYm9Nlij0
51f/fEt0pIE9DB20BEOxwMwZaouLphuG+8KShnoQ1/m+fmCm+V/2cacDbXrI
R39MOqatGN6dgtJ74xJbX3VW4nkCGy0O8lnOaOSuyO5rNlMuyqYJg1V/qOHe
YOm+WSjcfX1SfdoTVzwq5beCtTdNwFVS+b/zRS3Lx5+ooAupRaLGQU1TJB7p
xXgoPsyFz2n8YvG0A97AgeEAh+r7aH2eHvdagBwX/xdlqPJ7tRRwf4O075Eb
TkpHGxKBlBnhJ105l7FVujSTre8lG72ZFTRRswg4y7NdOrw65DqVhGeX6BB4
k8h4z6QfAZQhaTGcpQqcSVytqsQLqsaBOBUwlA3sm/HmAvXgKMJGm80r21w8
GvJP4zhf0jBC4aeBvFNEyJxFl4Zs2EHOydRHP+8CdVUp9x3zbxYdPysys64U
79uZMLD6kxAGpxHxpK3xfS3mH9930ceLs7Ji8VUYdEnSSYEEIaPoh9pDAIhl
96cPOEZNbEdpqicCJOF1EdTeSd+3z9Z9oTFIh+mQTh93Ci1x5RJucvsggXpW
8Gvb7z6LAiSOKbPBOnNWI75Q6x8HAviCep+dejcnOA31BdUZpKI88cJqBQQr
gQToE54cuPZ3E9XbFsCdTi62RIqK3OO8jKbThVvvhJn/1yRDsTdMf6v2GMsQ
ICQ6wFVXLXzzmzhDXCaHMdd4+lGLNkmgIc0Y/IbLdYD4XCAWjYufHTSqvL75
4ZfC9v4quynAv/aSOknaNzRyZNVwg1tl2XD2kgymJmWmd36TRn02o9EduerT
0Pi9usSdV2s+rhQNrb7yaVG3MfoLmHcV9f4w9AYDwrLeZ8uuJDM8ZFvbwuj5
lgLeqsxsBVugHV75Q8gjyuMwuM3EuUDPfE0fjDJqFyuWnby2KsptofAFX08d
sKY+Sv/ivbsQ/9npqB98JBN8leXE3kBaskeabk7ApVg4nv7vMk+2JO6FA7da
J8e6M1R5LEVL/qk16WaTxDWs+/7lbxlzAOJbPz/N+9obBhbDkbHCJEKwA9+p
iV+jdd+RGPx8BCExveFOHCGyddN0Qw7MO/3lFlRoNORp+HngPvgXCcX+Dc8F
X1vkbzcp0/i3PvlPyyGzFF2eBqieo+ZzEo/vyViNpOmMJX+3EPj/rmyiounG
XSH+GNzpr+YFolqG94iZEnFNLSwNVze4ED936nxK9FPEyyu5IfLL5lBmp/Xj
rDi71cNyXcdD+jX4GJr/xzndvNhojSmwPATWhLoJhuNFwVwVFVw9Ct2YDU0o
AiZ9E142bXYhe2q3Ofgid3AgY0MvIP2bsmM8LomMHA+cOq2mRrza5IvTmKTV
AFcMxggbXvmtqKy5drXh7t3pxx65sHB/IrxekSi+/VtwUY3mIt9tCE5zr6EF
uT68rp9rqJrpC/BH+dLhOBZ4SJcf3FCD6FEesl50cODYyJYbMveb6EfMwo7g
E4rwABZq81JFvkOnGDmvmJR3TJQFL8jyHrmKaeQXTPvzuMiULqFMe7TQngEO
knyqvpJSLEPwVV1xUJljgflf9f23SDpDvKj8KuCUGcYxSsCl+7kihf00ed4s
Nn+THKIam6+Kxo4mtBUfYlmVmGtOm1Wvw4Y/qyqlbb+VWZG0oGtOCLezSgz2
vDB1a6eakFFkQbX2Bu7HTaTEfTywm/WY4rAv0H/W+dY2tf5y6By1bUMiZstU
O1GPH+emmRkHRv9eVXFtbNQTpqqIXO3BsgaZpWqsHBQ0FIlsowO4B1qbNUSJ
FrmjSso69DHi93/5rvdtm+B2XSedEZ4MYkXNDzDL1z0jEP1lzaKAey8m7/JD
J/SUFO9TK2ovO3FjDDtNln8pdiE3W9InJMQhlnBi+1oH0Tyht6EVq0bvemSI
HGr650EcptfBpUj5rZFXBL81BnEzPQEfUsGNgJZQMzL3J9qpV8StUKyC9sNI
jpRR2r2xO78vUXUf0hbchquYMuY8S4AJOHYBKT+OQRSpIV34CJ9CZK7uxmxo
Q0I5auKwpsh+x3AIS38bgI4JR0p7CO3N7WQ2kMOFfxNBd//Mjw7Lr8R1tMqC
m4DD+K6dTJaXQbe8ZIu7XyGL15djGjObOynsAmq2aqVGygVbyG/m1tSjPblJ
0HIj+yMSbOP8Dqjt4tqBcGS7HCDGRH59AxaxU7O8ESUMHLwEAsDLK3TXBqKu
uBSSOqoJF1dHYi+exvgRigZpzYH/0PA6b4UjmeouT5lazrboo/rS8C/MK28k
WxbfktTXyZ7QPa4NeZwX4cNwCKRJd0Cuou4YAOUJBScK6oIA+hmuRQf7KsAf
mjF30nRUWZ3iCCm7zqgjOGLBpyFKz3U9FSVnNrnZjQaBnSTkC6lxr0cyUtA3
fwOZJwpO8QgRp8lR7kRylBext56n0yxJhTbuKjstQMtoyELZrEFwrm4sW4hd
Iih+DRJy5wmgDPzxFk18ZJaSYWhpZO3+idVPDpmpqjfNOe4aFRZSk/54p47Z
k1iT0rTbHP9Jn+bUKZIyZtU1EQ/a6fDR4lUNJl6QL1oBtO5pS/qygGmGkth8
m6Grnh13TFbsGF1Pd3nBZO+lCNmyHYQAgPkkXta5o7LVrOrE7mtAC2/taO0H
ekGyomBZtC0rsNMKK7s77yi2tjffmwn+rGPXKPIXOsmma9eAy24u3FqK5dqD
y8N+Zgg2Gu/0iyZWkY9tSGztUCFRiE5rSfvklHdD8rEFgQNbiR/zQZIZgT/E
XhcVnjPVywhNGVArpQ1yzICS1VmHPEfkNAYgTmzgfU32/p9BYUHhjssMeXo6
kXaUljWhaa4GDt4zwotnOdfTYl9Bb9xYafM38nc8GCckk0pQBbGsRG/JDy+t
ann2S4Xi6HzQqMHDWioOwAbhdbsa8biBcfhIZPuuMsPOFeZCuU1b8Tj2Ydy7
Wz1Vuwt0VJsvFmnrIvQeptsSX6Kg8VufxRuqrawLvqk0DcNgbP50ZFeo/ciT
wOYIcF/7cQBwY/ygvM55ML6k1BcIPgrCgPcQ+9q/+c3ekIkcU83iJPE/m24I
zX0+P69LfDe/8TanNu5e3apHTEjK4DuRorx+tdU+O3ScaxeahVxAkQz/O2aE
W1DgY4ek//B0hY8jP85QID/nNB8o17HCVA/cd3rS80L+WOwAgoO3cRb6OWQS
tVAAE862bqx/IhjSyNtge59l0aJNZM/K/Shsk98jXwKoSwYe8FuRhnzcJzDE
C9YHXD474EVGVmEWCYzxY2hxGn1ubuVnEPYLMjP0AVhqQXJUd4eAHmQsoPuu
K8v7fBDKu5UBcxFyTtchvAp8GzrRfZHDLZ1Qts9IG1z8QXFPYYyfTvAbR5YR
ggTZ99ChWnfMEdh1icyTG+AtBcKcEPHny50vlRfEjQWdPweqg3eOEa6uQCop
g4WWWoJSK3GqZoYTm24VqqRfQlPskDWUbTszC1TkEJUOV7Yimy1cs7f+aWRY
+9Cf+4iXFpbCLmzLDeWTjPi+M6AoeGCUvaJxMyb1D4W062YSBkfRZuYVAi8n
EpYiPr3XCs8bXu+wrwA7DHm1yRMgYJqjhmanVcVPzhohgjPrM2XfQ9EoGPx9
qCPWtQf6EbgRrFI/RxcA/tdyKa3RS2mnE6Z4mKBojyHbHdJSBuFAhwgLeEpt
FLrrnsZ+ByxSOZtJPDY6o6SVUxhhSm59qNPH2c/7klEOs0O4sMlYbT7uGS8/
oPvQx/RDfUg7ZVW4e1emT4GKotjfxc72bR3qCady8yAh7vyrmclObdWK2Qdl
YTdn8uarsz/8sIcunrhsQNx9Y189VJ06mWDlQNVNzJRVGpw4q2ThtzaQiiRl
j93E9iiwpm0E1HeGxFyYswcnZnc8XdzqzrEc7eiHjHKLjl0H8Z0mV7amH6nK
Kxtd8EJt/h7LYQMRCKknzq2XG+Z8rQTNdNmG2StTUxAJusx4TT74eioAnR/V
YFTYDZpJOK5Mn9aCjs1l7vKUn3LFDaSwVLCn5YsVoYkbmeq4GIR3N+YvLGxH
pFwdc1ksQAxW9+/HFD/deT4wI6WKaKOVngG3BPQ2LV8dR+fISASo9NsRHBYE
0pqHuLdDMFhJtLhbWQXLwX83GtWzuAOEiuBNnWiB7yuioQih5Tlol5Sn+I41
2mKmu5XHNIOc88Vm8UlM2U+JCHMGFx7FIW/YHCu2CMSJwBCg8EPSe7OyceX3
7hcJ83DMBwa7i2Wpl8LNa/GeJF7qUcuOVlLev76vnBXkM8bjKJ5TTRiMHeNo
E6teLPMnT3w5/nOTEd1TA9cAJtm0BOJlGhcfbKnXcR8idmBiB3vOs0HXO/xd
4VPDwUeSGYE3kbgKXE9O6+U1VlEo2uVKNTNCDRXftNNC/HUItulN+pE2psbe
IHRpuIXdu7Kk7uiAGAVf4cJfJbakrQhuC5coli3A/TYqrzaU2iXeR0kH1T7L
sjLsbzppZsq6mITwK3v7AvNKgVJ6aTciZhRpCviVYvo1wlvQYq3gPW1dD4Tn
cQ1we/UJDogeIV042V/CXIq3/VPbbhOFif2PQQwfr5d4kZSA3qcH8jlDZ6lg
9sRFga+yJsIDjlAMtre8tnE7gw8k3KHn07MkYai/Sl7kWO2uP3PL8ek6FJeS
tRkMD5qfpWZu6Mf0v9jMpwn1Sy3XWR6P6sOIVTffQ+9RSnX128dIbRzK1cd/
N6wrIwg0FODrwI+NpnNkPsSGzQwRdQ/qQC/2MuS1uL1mTh3JsEAXr+97pAtp
7pDruReMKr7yRKHA3YUef4bVzO7cf+AHcJF5AzRdz1hDTaIm14D7QUWuD++2
ytNOo3V4GcWw7OSsLi/DrV+/yX8xVlAmPe3HYIqrnmuRur65z6dpG8ru8vIi
Joh7GNI3FfPvE7mICmCL29mebcWyfAqJY0VpgkiM2DW0lqNRLneDTxCKl1RU
jj0dX6aGYXZ20l0dm8xA7k9TQXAJPS8z/EeJAbxZp4Ns27vo7ziz7QF8V+pE
r/Zv18Ygi4jAr6tv4Pl3oNk5JmKNNEePiApgsKZdjDN2MpTzLN+kjBn2RTj+
4CUn6l4XHx8X6P5gOA96LQSIk2C4AnmH+tuP8t/ym0o1GYPW7cXdrFC2fwlm
gvBlxsIBAefpyS4MVcgSy+Gb5li60op3MfrY8EpxPD9zwToX6sTIU/lFEC3L
yse3zbQ5z3iLe2UYItYvkABU8WN1WVZ7GNTfV2kBWBXnCRKzV8wt3VsItC4X
RVWQHKwAqYwN35yzIc3MdieU7+eUbqrK1lBdNXaiGUdb2iJQjEAd3kywLVRS
1tjE8gX9aRICMW03ijIw/GuBPwcS+wZ92CA1JovNqmdt5qPM7qTlxRx70rba
HP1ZrYlFQB1PzdzD2LMVN/vZPVLiyvS30VA9fNIhbc2E3Y5EBAXFJlTFT5aA
KIaucjyzGWY67LucEQMvy1qvR6xYmCULVr8GGcLK2ItMg8sCiyZC7k2wQF3F
rigXLHqf4O09BSTEVOZm+4DPdVb+hu7Jt1xxQ+rIU1DmE9oXO085pugph6i4
gpyK4h9i2H9Wgg1pMH1RqIpgCA7daKPq86rIf07B/GpM9+ldm3yyj52yrOYD
aA7k33dDOmOsyk4saBh6k0E4Xwj6/uQbESim4VqyjvhWJGg+SzQC1pxFUMJc
rUfpRp0S7FrEVuBQyUJ0SmbQerfVhSgfy9GTE8rT0x135b68hGwrc/R1fytR
RWW77lYORAoS1z0DiY+hJ84dxtToTEFLmK3HWBagxJ8nOruWc9QinvRVljti
ONQjDdPXcgV7T7peip6aFF2WCwxWuE2uCLkJggh3JLm5OlrZXD3VVA8+gi+d
yNy4iNg07pyTkGZF5nG/S41gl00DMYnmHuZaQ3NBmMeZU8uyVi2GA4SM+1uJ
OXPdoZK8567xOuLUZi8FoAG9Rk1sm+pQZxn3meLoBWWNrCdePjnfGZE81SRK
lvn7mDcLBdXFjFPPuB23bI6L45IETTQWXpWZsAQpBTZB4cGJTnJFTC5NkptD
UbTrBvboi/Kl+YeZmxK84Eynx29+mmUeW+54PHcfSS+vd3mC5dZYEr5NY3AF
44Bpy5NMGBay4w3DwecPDCVXV9aUzh5eexZLVpra/xgTZ35P/ps0jzmC2bZ3
mR+dZCDgUUAw6cAUbTW5iKPdIMbHGj3LqeZivmDN2CgfUFX7H+/MLX82sAOk
/nfZDoXfNNzith5D4hbhXaUMtStRPUelTAqf0kS75qTDoJtTZIGriotENcu0
vZIWibG+Q492x5O7cmyxyq2bPRMeBpVoXXSCuiqWQaIwXt0NSXR5mao3rVo0
5YG5D+6x7tx7IAw/nJOtqbPGXB03DT2Lac6uOgk4pF3W7bCWeTHJFt8Brj7i
cvyVfHv6fI1dCh/NQp8oQ+enbSkxwCzkKjposzyIz0Cvw+4obN1gRCr/MvJj
Cp4t1qGK3Q7eNfPg7kcYEBbUqdMzZoonC0WZfyc1QOV/UFAAUI5mJ5nDQLzw
zcW4CJ7W0mNqarACrZqcFC5WuZXH4fIero529W6jSl1IVVtDOJz9w9QlCYqZ
KVkjWOMILyhZ8eBDPYI19bQtvysl7uCJH2H4JzUk2C7Lq1tiigW2KwDREj8v
4Jom2JAbE0fcbB7KC77Op4VDr8qnqEmK4T0PjQZ+INyGSNFBSKM3rU3BTR24
0/vmG4J7SA6HjrR6C5X398AKMlQe7t2xPVFkGz0qwm3k9ynPZIntUXOrFMiu
men+Z6d81Ze4/gnRaUcBV/EjdTryTNz9LqkmRDB2uBJqPWmZXeKzGuk6C070
8+Kv5dpLX7Hs34aWAQJ1hElmeLeRvlZ9zM94StuJbbx75G65p6k5Ms+Znq4Z
a+gHrMe2IkoWyuDC03tCXgrBKzLc2mnb4m9P1WicVMU2i3icmWec2nuvVWDR
nCkh2gY9nhtfmSnJ24bjmmx9R3NL9rzjU8AeICKF/hsL4hTh+hJ5+K1UrVc6
q9ItPIVS/VzWd7Jw/+SmkZxY2bwRdCxWU0mFW3Ark4dzbl3EsyyHjnaGwGXA
RsaSTnA2HTp4N3X57LQdPogezqykDjwdyJTMVlmBCmvfksNi24tSHIdfdx0e
swxIaWeZe/evSvHU4znOXy/uCnpOkqG1UhLUKYJLkBObM03NcbpC6Pn5fxQU
NWdY/cR71S6i07nVFr8F+xVpf2tIVdKzLRrfGVGOwURLYcjLlW7NSuvG/dpl
pTNMzIXobH8JuTUBkjDTNzUicPUXHKb6dvzRAs7OF+ifJ0ln8IaP7OEppejy
7z+yeCcPCH9KgEKLsBrBb2+C78KzWmlJaBJhKgQ5JzK/K6XJ9sX2ucOGpDJn
re+f70x7bmEq7nyk9pLb4yEhLGEU9cpSeS8LJY25O6ALzK6f+erQ9ZCDUSkh
4A5X/Mh5Bc4Zj4muMz3SxUaDErX1sey/HHa7ujYUJIcGKDlCSFaA4Q0DxKgV
dJLqZWzSO+SZRbo4ecSaffjsCJAS8NEukzNpZQVjGcsA7XKNOvuqRnWDcNsK
PbVklfHsQXU58Up81UmGuvXFwNRiT/ZS/seoqc7kJexrY3zT7f8Z/X2Yy5xp
AR+zE7SQbzBBtO8C9ru1eKw7Rogj6TL6BihMSOqsSkvJG5tuTSz3mpdx1Xmf
gmEQWIaqPbdDIvt9KBv5+vPOS4wfW53AKSQWj1XAMZdRJA70RkIVb6LuJVZu
jC6dLqFeb8ZMp0twu1RsNNB2iMko3/MD5aOGlXq3uC/TNyulgoPLQCMXw+bB
Pyh0+qgsWYw5vP5EgK/p9miOuCqxVyaeNkQPMxT670TKyzo7Oe0wEKCeEVSF
1xcyNiPOUgAfUNGwXSQAY390rwqvul/FrGWOkytdZ1Yzq3oAt7wE1oz3xZcK
Cwn3dtVNiDZLXBl2ybqm5htaH+gUNv7sYqxuDSBteMbScqVPQiov468wf3dO
VayxVqMQ0W8D0ijC4JfRUKqeun9vNIANrPkgN0VOslNSnBZVjaFdF8D3q7Ep
Y0XAmxPp6Se3qkO4EvtEQ6OWIf3efd8PFqGkIZT+m9T0+V/ijcMoWkWg5Qdf
2U2SU2uxNtSvbKqc1q0J4W6XynSYULuixycnBb48e25qzWWx69VjdfNoW4oj
DPBXy28iEGjoaeZFAgcLeJ9WZ1P49gn32jbvPY3a3lhLCrtvhNDRkuBQHLp+
7c5l4LxgIFBtbHnIose+LosO8zx1siPUV0Rjh822jjASsjOd56Yv/TGOCJBo
4wDNkJrW72EE+5rX0VFQLJHvkwJa44786DzcIVbCwgumrcURju5MiPCZmPnl
/AeiUFxftkrguDUSxzCosJ2dG4d7Hkvhig/CdVqhKcSJBGltlBp8DsBPRuCx
thqCLSRgZZoSrjh65Cy7q6ZCTlYh6YjpTwmAcSwUSBNIgqV1CUONZCyGXtDV
NgGlYEt1JRNYME3Lb5+mjJ87lTkaCe/66EvYgnBSERcjgyHVjsEN7LMlaviQ
RG7teJfhcyObcOGiFy3Luv36KMEY6BBzzMwJSixwvDgehxwqarGyU/ebXTeL
hELj01u6gcpHPVKQCyANeGAd9rSHdKOJL08LeqZY0MzcoxtrHCx1SuBE0/J7
gMWJXkaaSKLWPHEYgDUK7Utrk8FOyKaBfhIb45qbCUdHC4Sv3SsyydWDXvFt
EiIrjKsVeCchzvkdMSf7g+kf4t2YC10NpK7+VhOYuzOdB+EujM2dvUE3HhoM
wj9i466MGA2YPEJs7Py5VbUxhCg9ho/zFk8y+pFzMubPVf4DHxCpkcrqQV9E
IMpJkWkXZHR6wStBTPwn5fMGSRYX13kBJTwav21CDRmMVT8HQk3UEojs3zD9
dMebmc4imxxdT3xp6rJeTCln3Z/JGJxJ3CC5FhyZyHAsJDlL5A+yp9bc65Jz
tgqx3eWV2l7XbBDgrybBJx0Jdx33Xuywa+rzyYKZQp7MEvxwtiGUpad7hoec
Ym6/qZsbA1yV6OVKBzkQxG8DgSL9YRQNdBp637nvrXcF2Mdgklr/FNf3U5aS
v2JPxcA1G3jzg/GXmahmzHRBnrDhCUGZ1LHJEieoEfqw9GPEiqd3NCc886CY
LVCyRkxHdD5YlZChKKYa18U+IKDqLWEO0iJJGJaNv2MzStYM45E7eHfkBuUw
ABjdnM71ekKKr35piuuXoT5hjermJVoxwVrsYik1XcA8GaOWFJMta7UICqpn
DvCNypTGUjkuvdn2PUwEBfz1A57Lcf5k05Q19iKbwMuBU6m4yzZDJ7USNN6Q
rsZnGgTKCSVXJYoLub0CpbVgOcTer2ZDU813neTbwfBMGYu7fNtJ/MuTRgyC
bz8ITZnE9lWTCnhKo4leofie19o4h57d5s1pAZTCBPFWaZjTGZzcLz02tQcI
VW+4lmCTiDLcwt7+co9H6fUzM5R8eugf2yr0TVj7IawGDxH6xZJBYc1HBL0u
5gVWeNDFUOddTdb0RgoLJ52mpmIONmMwIcHLR//5qwvoUUEuZrwt5UZBmqp9
Dw2mNbu6SF8/+4XNLAXMX068m61JZHfo/+N9nHSdWTtIpa9ba+aunwihVGmK
cwxrs/oL+e2oS6XRCsxzWLa1FkTUk8gClkSqDxgNlZB++WYA0njGQjloG+D1
IRqlHms0x+fs1JIEVweVS47iRmZ7XLegWH4uHBF6xZmwgecN7M3QPv2Y96BX
lPtW+Yn2VOFc1GJ6W8sFtjVAcnQAtqhV7aXpHhpFaX0W8iuE2CGjb6XIFek5
YwQIVDnrWNAAUiZsWSrCMiJyUdsojvC301qIe5gfmp2Bw9/PCiqq+UskNZJo
72+AzwpGkL6ie7cwT5uhZVcSe6yVeK+xf3XiAslQ/f6xaope9cf0zOGUB7JA
+VDjpaDArOhBjKkXUT+dcZGvC3HbbrycET5XkJsnhlsf5KOZmjlpq6vlgH8Y
T7QzS7d8iXheSDEBJDsw3xBdcqTQRDwHSejdU66mFMiJ9mNpfWkLXf72UTrC
1Y2QoppD0tVUUVbbbx6BFDJ/IEqSBEHEgrJ7Of2JTUK7biwL2dHihTe8paJC
U1iO/hPlwO9yPf+YvcpcDpjIPJ2ofmj1LPk+abPI0WOCWw90oBjp8co+Biu/
mjSB/m9B8MFz7cfhA7FBZl/8W3SZ4H1n1RUpfiilW1Sb3vOm6nOMSAUCDvSZ
EpDFwA+dTb0qfHF93cRJSeRBvIJLxKqPO1NHM2yP86svPVe47SpDeil6FS9r
tlphuBd9BGJ7CgSMwBIFkjE6BAnXsf6Wi9r4ikEirHhScrPF1Bj18bbqZfsn
Vdixx85kh7h4PLWeUk9+H7dy1Ien7RjMJsnsynbTs9O57QWrPBfwuGaOyAVm
pR250x6NiuSm0+hSXrSMgb0yF35xFBeOaiut7/GRYI205iRUSEzZF3Sr+yAS
nyitzqcnofwCT3HwnES6kV/f26sulqW9quGv94zpOK5VFwrti9umB4K/dN0d
lAqPgG/DRMGuCZFrcCHAi9lmrNtDd9/sDVdsVr2wHb9yMjMLPZY/6aos8xMp
i5idZEfFM/Gq/5exOpZIK9GEP7PSit1am9jP7QWQWi/MNXdlNv5cnwjRH/In
ofM133M5O0loZRaSFh1ORYG93J6FREneguFJ9wRX5Li/vukQKcH/HayNJ2xL
lHwcNRpFVdXIEIUq4Pqh9XcOxM9i5m/7jHG+H+GLnZO0kXdWUKs+LHaqmxq0
lmQPR9s33SZD2QSrd9aJgJTP2tv/es3egSELijbVoqYN4xCGfzKH/YHOirwM
ticppFr41ehEq88A8s+YrsQ00Vge6MJXBxNixJglsngjQ5CAVKNzwm+LzdUJ
uyy31yKzyrVpNMycq9rMrxQ0Hpd3xLCPmLXJ/892I3VJc5N3U+m6x7n8nEYv
YwmqOrVsXGpYywJTBmM0ocWEJA9m15F61oKdIIiImBoDcW2c1bXff7ptboiQ
E71jFu5UrRlA4iWSQbK03fffG08gqf90jfcAm2539MmO2GGkQFDNh5u0Y4qC
HadvKk88WLrMf0ClW/ZC9fJwwTyLObZYNvctB5cgBdLoBzLgq6d2dy2ch0+i
tk6oeRwPsEAVD6U0yDwk3DpP1TDj7UmWtXx/dEmaApXt8OevaRE+9Qm9JJDr
7i20UE0lLARnv37P6am3tPSv5lyvzIgZUTcNpGWYkm4lCwsWOQQbAjbcehdC
Wb92nD/n12OYP+LJbpBpQ0ZVWLvmirYqjh1oFFTR0PQiGurBbXlSYnYdNyqc
Z9NwI0JhNlL54Pk3NDO6t24gOiroqPaupCqOJkApDGkS/1ti6e+BjMvosYAQ
iiVkN1l1BDBQvrGwqK/wVF2yW3RCxFAFq4c7SuLXlIh7nvxtaWTwaCbRQAWX
YAfaDjHvdOp4bxz2KSo7JusJQW4RXXspgWZjYVvE5b1c3JB+6gDkvdt7A43Z
T9Ek0DXl9HS98InYoGhcTtyYjXXB8BpzhhMyvqCAV/5oO5jQo1VtPwOWwu9A
TyWY476msys0kUorS6sGcd3bw9EtEc7kglHJ663Reb2BknqwRhIt8OqIqgx/
0284IQ7lzjH7lHxVvSvP8GudPDprCqUxF8HSGXNUM1zfvcGGuwkKiSQAeCJ8
BVCQod4Dvd6EDMltBzSvCwPdWhzIGtTTestbiDAW13DNLvQO+DSs+Zb6DJco
qE30ql5+vZ+4/mK/NwoIJ4lDLuSHFu3aq1QHek2biufIUO/9Oz6nk7SfjPPv
epPrdi/cCi02zCsMo1IZuFQ11O+8YSkQAHVoYPX07+Qay6Eh1dONyXBbOy1T
jmPpglUSfMfB4LrfW1DUbh+VNXZFrRDxnIuD5yf3/sY7P74Fw/b+nyu2i+Y+
bgLr31RGcSizcQTkHwgRHSqhA/4uWYTk2Day7kzYcvHMnYheP5+UTjLfaqpZ
Zm9DnWn2Xgv1XG28WZV2Je6T6DJzegFpmbmoklNlK9lpwuVKh8sCT994Y/b0
L6SA9Oy6Y3qZClNZzo6AA/QMnfTa/00Q4Hqa6INEPvkpzGbIFHTloFx+BwzL
bjGiV0P4p+ak+nwcJyAJJD9fWmMcIlIUkYx1vgpRr0zINxY15fU+R98MBOrM
9tY0gqgJdCwSu601MD09I76WQ9gNAskHeRpDvdCV9V3AscqRKYTz2N9k1CbC
cIVaLpDXqN5bFQn0DVhSZ/FzY7Crjt6c9yKPrLKo8OmjpPrYQQrfMzAqVvD7
evREIlMc7v815/OOsdPZs5ChAf7l2RsZWxohO3lESauB3XuHAG3UP1pXj6jG
id4kfRh2stvDV60ZOEk0WmjWXRw0yrtYc6RKBqzML+x7AveOfxsNGZwxepMD
lOis9fpluxamX/2SNJejHjJeJqZ0ryVIRiACTvSCO+2SBj4Vlyxls8tzGJCm
pOqya3t/HdJmO+dHKjOuQAmwBVlCTvo5CVhxhyGW+aeUzM6o5Tm4ughFc+WI
EuHkW9PKiaXXHHGqN7hxfk+FE0s/+VrlCkkWnytRNdI5ZAQmtQT+ucmGIMIK
iJYtGQmvD4CelWKS2NVn/gNRSgSavs4GFI1JcVQptUuH/DCbA+ulSTlp3541
IkjOw/ig/0umqsFH4z3xiQvU6nC0c3RtScosMPcA4EEb7G/hvzs/7Rxqw+gR
cRrv8k7/Isgaj6Udk4GxbKyntqXQKMa8s7EKYJw0ygFEzggsF/M07rd7jrcz
8XiIVzG5RjLGNHFI+bnwMQVqrcDhTNOqXEvnEiSvvKtDCYaOujRDIEvuyosi
RyEoIfijwgBtFDVLdHeqD5jhQRu0jOpQH/epmZdPgXAg/5mFUTIkExNwfVyI
+pfQjKA9rJr9RMGEj8i3ErNEcH1al4rvfr5EDjpbpQC3BpV1VXTZSgkutNmw
XV4VxQm7t74vDSlTi+euhqBKqq5OqRqFDE2HrOBqnd0e9O/xQxKkvgUKYrQi
RKRwB6cypcKY3UHDIuLoaxgQC45LujL9QOwRRzWOYKmDdoovtZI8aiXQ8+aq
RhC4YdFcEih56SfO7XNLg8E1IxeJFLYy1575/PuwaATlMXOgvsFK5WOHjm36
v/D29ZZ2wdv4XmNN9CFvqvytPajQX3AtHA0l4eKUv4L1IP4QvZ9VT9decYEp
Dxsz+vtjoiCE7HDfHcBVvL6fumSxXw/Yoh1g6UBfX75305ltJ3B/wpcB4i7U
R0nKHGFPEG8MHOa2K9nQl203IMNLViT/gcUO5UC5rNw+BSJL6ymPgyHTwCkF
YgVPA9KkNw/IDhGwBsCcDyIYcTgMyUlxLTFRhHzx7tsgzqUIfMozucpLxrE3
W+jP24iXLbWKpOf8rd8KrupLLS2wNHFdKtTVr3DpnE9rl8DcAoUfuQMVWnkp
+ukIspowsP2wBM3QA6ntzmF2S9+5ja9X43hJImhioy+ZloyspmkLzOrf4gOR
7WzkeHqxP4p58OvxDgJNemT93dCXVNrnbQ5FsLadzkG1nPmTBgaBg8tJ9/5K
IkDmNsja6men1H1AkKSJPvMML7Q9EVpv1r/TfSOzB0VIVa6Owl1TcatNwcm7
GhiajNS8JCb8vUbkPGResQDkg4JcVED3zmKrB+EdAho5Uggo+peEpBhNKp1J
5i4RSHkOzLZ7vJ1TW3E6BM9R764RtjncZl6MLndnNGTsRTiacRHAJnYcPm4A
Kkmnuvv5w4F16R7cdWIq5tPeM/zL2mmcSPYguMP5QOomqTzdjN+vFypWFPce
v7/t+EreOfpsx4IbUd8dFFNN1UijtAko0xKyG3A7MmwYobYX0Yoj+TrSCP4Q
oYjw2zlxvhqbnskK9gmT9kbpslW2VPQn05kiFSydF4WFcVufP5YccnSavj5B
KTPSYrXmnMMuF7m5Sl5NauGTq1D4oY4sS1dXfUB5dMZS3fgYIZ2/CpDnbt1X
sECy0uveirGanzWmmZgx1gK7TvmpiT0fWJ/GYT3wJwm9EsdzZI7HMJl5y3z4
7eTQS7uTSkNTzoyS1TDOX22/9fq1b4iKXz9plEL0aaHqjh2CwJz0TrH3V81x
MrFIqsDpw0wUr+o9MG/+ARHF7asOyNzcNTgEoeTpbDWnl09+4MUM4j/AI7Gj
DovSbk0vCx/6zMvjjAwG5RVUgll98P6SQUsuvgKQLhQ7xNIJhTKUG1u/lCAh
RNMb5gaYqcQb3kjYhdh9nHXpctVBFwPK9wdULCOSQvyLOVGzESHbV1cCOmHr
H0v42Rj9uciPOMEzxPKUJXimNej6NHI+hWNDjL53XuvCkyFAOBVy8C+V61Uf
oacEmH8newgRzKdMvMlrE8QOj8pSYqRZTd5r1ziLg3aNRjTRY4qoRPU84KSR
f5I2M/qmReTiNiw/n4VOccbxW3b5lwKEu0IrZwQ3oEjv8RgUhuRZ57Rcd3S7
CTCR9svP/y8/yEPporK9MvtWu4nrPKQlFmpRFggZaf4ZcfkSsCsR/Kkz3ZL5
wPHsWPv+n6/ZS9EUBMhddysi48tnVEzl8F/kuJP+yUZavNdHRXYeXs4QcQOu
q9EnhdJToAl9JhDL8iPCsIdV4c2QEIK81IZMrtKCHHf4wKkPT0etSo0n/rsp
Y0qXpt4sJcv6oxPZHvmEIKExLzPOd6qCDz8YpiC4lduMDr3hddRaEWmheO00
G98VNM+geLig5xT7cAqacMGpUyvSfkYuqbcgxE6Ek2eBYchhzYwb8NJVH2JT
PTlOB0NiMNx65QoqoR+ta0yGU+tN1lHD8sysTqLKBdOgQLC54sYfbC9QGyQn
T3EUEZZWUy6yn7ovk8AdPj8f5zzjhOLbGRHHMv2lw0s4yrVWCpVB6mOTrpdC
PjqMlHmWAHOTCskXmo5ouy29kwiQ4ZgAVNuTKtrRNAtJ2+fwbQXqetLlPYM9
K6NYG5/sf7G+BDy2x2byspIXX2ptE2aYC3dbYs9Vyrr2lkXCcZmebQbNlgZ5
wERmUHTmZgi3sqkwakTxdlH5HwUmgagIiMThQ+yXCGtFTF8Lxkxm+ucFCNWR
I9ksceAQFAckvjaIy4Wc/GuqgwLuVhM6sQAtF+gpVY7czEZmNtLD+DCPKrLZ
4HPWPzFfolNLXY2T1vA6fx5a9cdos6p64DBqOTp5082/vqdVPuq9W/ZKM2h8
AfWIoky+OgkpjE0Z1NWsC4csxxV353Zhj2aQmMy6xzB/1urZFYh4nsK695zZ
g5xHzTYtHm0qCOYnQU33AuBnWgiVGql0r60jtaG+wx8/cieqchsptm+1hIU7
FjPzSNinjcxnhWPblfVe22MJ8QHxxIrtI/Lyy68tRB3F0jyCyKFLK+awK+AD
hEAeAPhEyIAjYQJY47piphk+C0XEIIJS/ddV8pNCNJWqDV6P1LlcT5ZIxX3F
kA37wu6oAsxKMqJH5oHUYhi0dR/PQuGT3WOtKoxR/OlNgCye64/ybGIdCPiS
s5X57/Rvr2V1Rq0aUHFsEvRTpxDHsdJSeONGqyd9vIhLVw5dZMTQ5dVvJszu
1BYBb+2cMDE7qWQypcPX4zZ8e79NbKd8iLK4rdz0e5NXK2pG14MhEJJblgRd
0G2JzvRyf3I3daVLTEXK1/se9f8AQYbn7Vcu5ViXwtuYRDsXe1TUzP/gbl5v
u9r4j0K3t0oEMW9TkwKQ2GPuPA2vWTRxrjNBvl/VPHJEreByaj/KXkz/QWN/
3ebv1PxdCjPT9boK58fIt3QKq1q6M4Wq7dWVdBTzr85QDQdRrm+EZSAhIcCf
N/ImQHUossNGVMZyCURAG4u4qX0AsN25A65K4/rtF5b9U0Y786B6yp9DNjAz
t/GfIo0bhUevTEWvHEG9blpMbzsxVVnx+tDNYhffVfD2habicqCVZToQbUNn
pwn9QcCWm024EL9ZxjhoTfTj+OTWezI8eFF6kX9mLWcAm2Y18tRECcq7YiQM
0SAby/1sShmhddwBtO2LQvihTRgDiAD6loIDXWmtdgqYU0tSUAOY0vI3thQb
OBR8sbWpK2TmXzW2jI7iwNvIBo8wB9Uz3iYA4hpjt0Tm5Rd5xZ3coO5V+u6W
A8FRWpqQbRbV/5TPdi1DBWN4S6G7itnhvo0+O1llykqcc7g/U4NCiXlJxUT9
W1oBmi7loeqo1+pksf2sy5koYlHCkmKva7IgVYruuyyuR+wGoMRuouIy54xC
I9OvDIGzMM8jJOFoP1JsvgzyEFFA59IgzocbQrX6meb17dCOqhM3JAHuplXJ
2Tb/CAkGkeMLW380IKMkwywd3IYZWnFRFh4GeHr0moz2AkkkgJAov6n9HC9x
eOFcQnVCiFC3MADqEVWJTIvsR8pMUMlLItqduK6hO8OFNCQBhkzIy7cpCrMd
P3U722OB/5Au6ZHulajak/1E2GomqepdjAfO5xNnilNBFE94qDTUDE1hS8Gt
gqE03v7ZCyDhCsXk1tofG9U6aPm2nLJJJwc0LFRMyzGP5+/ftiW5EqssRhK6
TDWJtvgln35qQLnxn83u4EH4Re10IZON5MnA9S7eMgpQ06Ze/ZFg60+eo2e5
Bz7MuuTmWpVwfk4BLyMyjKdX6/+CnzlmUqAk4p3DxtSwrmh1pOA1IwkOac31
LVbRPV9bvkX/2nSbFX9WGNouz5SJs4cwKnuXUybySz0bPRBOxWUIQ+LhRSzn
P6I+/ijtBvi6iGf+Z7Z5ppNI2GhsvbhOL0xZ3GT3mPiOZ8QmdJCA/lkBz0HH
MGrgheZU9iIgV+wKtfRsjbRSHBWEjBcjIWxoqDJtaPDFVmgJbWw3HLElzzhQ
0KpggHebtU5oLaNgYsqAw1FaxWPHeIy4IV0elkzjDjxQBvpe8o2lglPvYllJ
hbjobMH13ijRtwPceGVRkY8617f6x7z1ftFXn2mfr8D+J5QDmheKGfJVYtfq
C77XHtDH3HG+Ge6zBhxFAzZqv2WjHxSlGUURW6HxVH58klZA47P4C71JPQqc
c2N65YtBFBVp78jq8zhh9dGgA4oYjCNG/WPRMNZH4vR7o8T05Erz8n6S9pKL
rPmfq1a2je8yWbE3aWonltEtlbuvri+Ow5HGFiNSUuc1RFVP4ittIaYQu/WN
vLFChFm0nRBzpTMRqP70aFksDzQn6sQetM4U02GKYfnJ0siBzJ2PY4wbINT2
W5YTFeFNqs+wfkVQDMbMdnPnxi/F2/LzFSNhpGVZO6TootjrCPzy4wHwqAXy
VmmukfuFt1R0d6lVhqMad+4ysGcWJboQi2k+xURnwuSipwTeXtCe5qf3aYDM
J/GJ2YRE2M+T0W95qdw5BuVGp6ZQAaKAyyeU+tve4ztKaPpmB/AOMkrTzhcO
SM4KBCU/SSIdh1daJIQONOommAuJMk7EZd9Bv/5K3YrY+lZOU77uoDEJDsa5
wxsLLh6w1N+SC+6U8fTDrPZ/UJ3wQkb1D4vLoWjMcIhaO61JnqOnYhf1CXTh
fiZOaIWKTuIyTqqZ45aisya1l2ZQ7UFh+9vWGiemaMR6BddzQKeypFl4D7cd
xqRshjdbfSBKLkzM13TLhD9CSNUojNI5+s/lKFG7G1rKcE7FSbFWGWiXYnJZ
W27nHKmIMewD7wXSmVPUkZ0dbqhuywzpxdDb0LytPCDOXyGI5+dDdomySrCl
dE0gb3KMa8CiiwnazYoRSeW3uajvoFhm9qOs7VwVQW5R5FwN1KmHLDnM1tZl
BWndjqlpUdQ/OkNt3L7Ffg/FRQYNCwHm47VQc3k/7NqigSEj5JNq6djJJD01
jnjxDR1lRVpuJ+MNnM5BIIHUkE82LYfLsKTve/YmmQiFvF8qUb0RAS0HN3sK
6zgBXzbl1q5Bq9WFzAIXczeiV3jLGjZ5TK6c5er9A1c9ExfzAjZFx9Y9pQv1
8efrk4ppmN5DKjoXncb3hbpj/hfoDgigTNRc0rwDvXlZZUhtpmePuITyHahC
hi6L0GULkim2Y+8K6LxfP4iyMZNWhC16E+foxqkRtgK/hYNZtEb0s2VgOMlC
q995NBioXtvloPp1PYQpSwzu+YUH7KZiaj7QR8f/UpGBVryObaojkI0eSoRx
syOFxfk0L1Ux9VbvE42qG6zDWr9gDF6WKoM9sWxYPRjlVrhrL/Ge827nHDGA
wZb9yPyjXnCImLpLb67ugH/dd7anLt4WPBz7pb9Vrsu9GJIgRqFw3ljiO43v
vkMmdVvpy/+qWRieMNuXX5Mwll7trluqJk0xrUAV4UjBqG1SKo2E0GIO5Eh/
yKcfyHTCgvC0p8kZY3q9NGytIVICW774H6jVRad590S44nwim610DNHsZPKI
R349JBJpPJ8A+8xxZJ7/x4S3a48bftT3wOqREjfD3MDjpqHmRb9/1VLQLVzL
mYBIke/2j+L2TZRytln7mD1X2QYYoVS/xOmQgluDu1zXxFqhQhtYGHzzwelb
ZynHK6H8w8JWuDAUA2jtaKLQFyiKZJukeSf61D9CoynmeKskB6ST++7a3WCb
A//rG/Q5f5NA7FIAoTSjnmns+V0mZ7n0tsKosJDGnQPlgSaShG0WIiF+ZWow
EKtR+zLGEbY0oEYp9wtpdQiDvU04bXcUjsKw9/4sObFpgpB5wcwqNiUO8DXx
eq6/e9/+jrOYryJ1FhTyS4chSY0JmddfE7tE+UTdlTbY8Zceeqjnyeen4cJa
FsdJ0tM4o9CuAVAASFvUWoW7Tkdsqm4aJuakeuyJB41hU7rQHrFYplYm8aFa
6lrZF7c1DWDvtm6lhHhWTL5Q4kjPeal49WRs0b6KT58kEyFIcNBXytHNkmgM
5HTH4cgsTnIHEI/udO6KUWq3G7u3/pcUJWYNBk5jS+SQNnVVnIWR/VntbHK7
ESUxpf+/gm/CduijjBSg9hs1AuqipJBxpojT6dm9qAHUD5BPt6vtc5u5mcSC
hkhM7lRSdTR4pulFWlbxhLEbZpD2ts4LPr9cbpH106iHRBUcsYR2YUWZvR7I
kesnPMAlw5cV2pg1roA8513lIHKMxRzAVtRnO9G2J7qdF73OeDoCs61jq43N
QsP1cBPpk69a+lqLmpt2dcdeVwMKL0F2e+GYr68oflCW+rGvgmUFxwJqYq67
KUISHu4Mpxytor4b+BRpdGyFh4alYAm/fwasb0kGssIhoSkkjtRO7QyZctaJ
j4zeCMplAYnin7zLcX3tkxh+6hi87RpAoIuy0IszgsoW/m0xQdIT3i1HGbUl
VDla7w8euCxSe6uy5vTldDplgSLTq6LiTHZqWZaaTydSChKlIWhpaFcynJav
AfRORwSs47WZttseumFxNs1XNGMVrHbdA4ZssCBnhsoGxvoqF7pt0KftcAJJ
wDsyqHDZK08Pj/s5miQeoPUc2IP0JHWrwFubRWEZk/IGlYyfy0BjQOal1sMD
mOSiysZ4bficGFEiWyqZ9MnP1oYpMdsPXkuhPI2RE862p7C3lh6qitjnsMDn
k6RoUcRx+8QSRntJgQqeANMSfKAu1P6HlKotcEgzNsWBwTnmjd8wyzAKJNYb
fFOos3O23CxhqMbvjXJroAnDPQmQRt1Aq8WpQ3XJryqiC/lx3+WgIdYT4wMO
RzPrsKb/z45cVh4quxHiYNb4v7dX0YkZaR9AG3xlM8rMTniOFtxeYATgkOeg
RBXqYcPYxqywqZCFZ9w7tpv+gochQxkLL0z0h47jiLJXUkXtU8PxMLps0Uis
25usy20dpJdw4jUUuYqFvMBMxrQgjsR7nvdGqhHfTgrxFZqt5Ok0czuCI0Yn
bCWtYz5+IxyZWs3x5oYVf0VZq8rIv7RKN4S0i9VhbzP9Fk2Is+67/hNbDtWh
MDv1vjQlM9Mvj+n2LImaGcpa7CRCS2c33x+IYWMpbQBYpQ3qSh2smkHd3RtV
z1QXfXrnsC/oikN4EeKtgaC2fosL4rOQnSIsi2K3c3hB6JCQjYY93e8vdsbd
mhVLyyYN5QLg2qurgxEtaDCUi1k5YCIPiY27yUJUFIVYY9/8uFKU2NLV28g0
Drx2JI4PxDi3/gKA8jlZYsjfGQhiYQBNu4AINCuwSIKOg9JBP4D7Tzb/VZsN
llfeLToCpbPi1r3e5aAsLZgKmkAPz9g28ALIqVphFG79gdEgrVePsS92o655
YmDn81uQZW1Q2GCymAB9MsG+5HTZvYWCsUSKVW5+R2MTDUrqJh0eMUdZwQdZ
f4Q1E1bs20G8bg9VS5UyHa+sQDDaJD7DZ3MkurcHiglAhf2ETdac7YLopGzL
+ZJWvAc4GG4Veq53OGGyB/omJ2+gbmVMGa9fI4jPXwE5oj5zfsyHoQqH0Q6W
Vo0iUV4UAAVyrwlP+RjHUDqmSZxFPytbW7kMl3wKK8WsHBO9wHHrU1c/7NZl
zP6uQ9mgItTbKXyiOnhFIhTs+n1KbBclQf++lyLsl9eEw7238kc4Z5/6rfwR
ILY9KFrmUPBh6T4405x552R7tEl4tVIsyFjjSF4ZXhyuFijzaMmsCM6RHpIv
lzGVnAdqPteYvNlQZDE9wwyE15ctGt2gLyMH3ztjcav4+QFpVyMTm0QBYnon
5okPD5ZRe3cAuG8I5YpUR+HcIg9qq4LFsXCdC+57SXCTigDySqw6NZPgCYXT
Isx+/0wSiOn7hwWT/LxDJVBFgUrTVdcs97AjAZ0/Zjn1M9gycN5LYeHxce/Y
diE5qSbGxdTyo6FkexbZ2nFybLPi7BzmM+8ukHeGLwapvy10A1J5zL1hRSeE
Fwm8jkqPuMBkYTNMwDYm8ZiprH2VaTYAOCxmsik/8qc/KwugqMtV6PgKds+q
D2KxG20T7wrV3rHKXEWvfRimx9ENtfYCWDQ4+GDHXmCMpaizlskIALLJ97RZ
ZLfxKY7B5RjJVc8iDdUaobnzVySpRKY31cGc5xTXqTaKgOVhkgydMPLwnJaM
V9s8sUMKvs5bt3yN9y0mpo1fL/KPNB2sYA06tdprEWMDtK444YM1qjZ0IKTV
jbTDsnYDp6j+pC0kpQdapqbu+l5yBlk3nAa4Tjw+5KncYU9djasBTFvxQt8d
knXkz2355f7npVOvImlWxzoZkc2Zat8v8r1YBhHtX17YDGndcbBJwfnPneKX
XAhpuD0/FOJge3QBhJS3bPkM15XudhiajukMVlDKBxI558/0bUAfU4wgZK/3
c40LddyQExESX5xExWGHYc07BpAn1ss61xYlZzzcKmhPCWiJ9pgPAn+bLpGB
hYBgfv9iaBQXWLHzuxTwWO6B3LJkj9sn42su1xREVHJQEKp5zMoqP8wN+Dwj
23ySpyt2l8xIMhtHjs1Hq2vcO5c7wru+0rsbbDqLTUqju1Pc5vc8pYKENiR5
2v/VN68n/YAwnKV+9RpNKT0Fbbd8dPcytqnvfuzv54gW5CJVDOFlBguXOGu+
uUFAdhpvvHQ3nNithR7lBtvwtBvcxioV18t74kPdjhc6eYzNA7Vj1WdCkhcD
XAj8GOkY7YJ3mmc5FC+LHIdF6cgztu4gvazXOmua48PLKOI5Mw+zYIdBslEE
6fiJfAAl0s4jUYNUWm+q1KV1SKiHGdVfmvunQM2z+p7IFTuieg5LdxZS/LNu
TC12NLnwWhfdBxEv85HA0et7xZgkAYsdQF4063e72F2TvJiNRMh3uDiQWt5Q
hPDyopOzbHOck7tw9Kf1VAAijRJ3zniG8edLc20MPiBDRCaLJoNgpMdVdlA2
OKWjoyLLDrf7vC1GUDrAq2LEa3+QZ1mOn16q2/u6IrH7BMSB+yjRX8aqw6KJ
sn7EMvpRI2l2iwRjDddA45hbYu7l2BOHMG10O0L4+HhaFcwd1Crtbg7ogjPG
A/EaBzpFyC58X0zSKWVdPiqC56mnXNBWO01n4xpEx3ghzqsgwWx8XxO5OGq3
cQXg7RUGtVps1KZd5N9XwyfEWLowWyImwH9VvOcmK9zlVQtqP4rrf/rY0kZ7
c5WWaThEvTziAd3pXHIUZFx6LgAW/k3NEfkBrOaG0E6+IJ5jIQa5QtNR2Wor
VccuxtHHMBsq2sL+c0BAsyB/MuasGhFKzyFu2j4tVQ7561B6Zu7CqajLw1Qd
dTuJBihNwKSDuFK04iRtdsmb/kmD4csVt8nG5K670cXNYYa1ZqCBZHoBTlkg
/Mx3A+l5qoDoNvTFA1oWJRbRGD4kTbIfM4tj0q4lKB+XWD7fXb0CLmVvMdir
SBp8trYVGNa758ST42dddyeUr74oTA0DR5monJYn8JQHfCuj2WBcxftRg113
5xGLESdm53N6PtuXBA5GAvGNYVayg9EvGx/U8213KCukj5JkytpYCok65w8V
mjhQdBX1Z2CCBniCoSCiBYeb/d86TTmC801qGWQ6IU9B+huEez8mWn82PG8i
jaMgkU4v2XCMVjZsjnxVXhrN2mzJGVhmOVe0LsTHDogA00Q7DvcLkFd2fdRI
sKpYJ4rwFSQyQG8ZHiZqjrXoqMlNN7uC3WsgcqZqwmsV3eNuzk/l7kijv6YC
hiHhxRoRHErcVHOrUutM/NpJqFrwL/TJIqJULbgscTH+0fc69paxjD2xlytN
amVLJwPAGPi+M50K0NA7FOND6ARZ22LzKMV1Bqlv1lNRWTVFUpgV+iHmfBpB
0KavUEfzz3JeYwRpf18y6dCZGswe35B5Tjnj1M4gv9TGxKEReEy9CVi7BAI0
t+5TrZ/2pdpK9cRlGer31VKSCp1YGVlIYLYBqDDfOM+yjU9z5JJUmwbX34tD
2lEHfqGdxyPxOhd4eYFjq3daIGLlszuiXxvk+DS6SKel0DTc1A/OifEALlBD
S5IKE1NmXRPl4oATcZOU67qAixRu3oE7fZWiW3Lkxz1IZ5fyGopIgSDTf96s
TnISkMslm1w7Go40YHjCm7hqXwKJbTZaNAwqeclGjDr0CcRfdXXvazmX80j9
HKNBhK1hZtyp0ykGLegEBRa55tBlZdVzllHNILs/ijzpNJsbaCvb4F4mm9c5
L0vU2PV8BiFGwJFI9u9jpLSSrOC5Zc4yAuQ/FKrnKnrbFQ4iLCfX1m4jFtmI
c9gv8OTLezd3EnclTuFlq8eBnQru+7wqHqWCIB78pyRdTJW1uSyVnY16FKI+
cPhiMIwUMIBm4YTFgDLCfUcxMWp0jM3NlqKvZbWiuCF9U21kzgEKaNC4+D7Q
zZnNYfT0F9HpV+ROBXNAKqLtltjHA8IiEPXfSdmKO8QkywPbAGWolj6QwbHb
0OtztBYXma89xciSd/WtqYsEVuOKpCS8z3GNMsVjSeurzXJkvKPSiMxk7qQ1
Qq1KiOcMGLX0rroQj2moF81s22AWaB9kmXHGwhcpaTvDb1bfiDQcat2/yuL7
oxZJvUUji7VocEB9brJIc6TAE7hC8hCnQGo9kFlKJ/B9n9LcHweENXl8Migt
PkizPmyqFFWHjanTf7ose/mUcYuy6PDR9cDd8+I2adVaq5cvFm+RdsIqntRV
s9jWa2pk7Ua6qCgmHIe+k/E23AE+4rZsq9NwyVnDd/wcZ66xL9pXWDNbt/pp
McgRwC/VRN2OhyDKvtZj+GHtzXifn5CZHylMLrYsFA0NhA5XsBOb2tEvX6xx
nx7q6icc/DYwJx5b2wgWqiOKtxeDpk5ghYWA9oeIVMG96ukkwDTafVtAB8yU
YMCzoKTfR190A1w2hP9EhSfhVHV+Rn/kiWYDepPq5s9uxuIRVMVprQt3cq+J
gu0SlFY0ta/VBX1Z5hME4XrKavoTdv4eXuePIWpl4CuQkn1aF8kiF/iTzaOY
ZvraxP8qzOHKDVqZs1NlZHQo810OLhcLou95FA8xg+5VX+AZ9E7mpy6RRxD6
rVf2+gq2JPNGGTrt1g8LtMbprVGxcQm6r+XMFbBez/db0lTmenjvFPMGwfWL
6r7RJ68Hsmr6iV8h5bXSJs8ZjVAZZ/DS/iZ1Q9J8JBjOSP+H22zSz+H2OjzF
fucj4HGQ1L4Anfg6ARDjYwb5l+4uYpIHPjDSTvlEDi9ecPIF0buQOMHzsU7L
6nRdj4PTqw66nydxANuKa8XYEe1DystRWCzDvGlvlWIscPenLZkokbg8PXIU
bJNHnUyWK18fyljObDCyVR8v68q9lNPChh5zoWnO88Clqm1NCHCme1a3LnkX
hfga0V2BxQOlzwQ/NbVPrBkF4Y19QOynH/c2r2y8W8VQUcqUAFY3fQlV5ZOn
+gXXcJcr+doceDb+/Zkjcbxv7hHaIDj7oZO0+MJF2P/h1aDJEH74QHDOyMfr
sGoySXPSUMEQ97FujGEu2oCWDdvbYXMF7sE9dxJzoMQZ0QRUrrYq8Cxgj63t
JaSz4t7ALCaiK5SpfKrVupKAeySOakJT2pnXPUbsZ1WLZ4vvbW2BbNyI4raU
viZ4adg6MJOX29E8Rs2k/BLXvCkfbzNJFm8EC3aMRNpCh5edzlp9iV4hIJBq
pclGS6YpaGCpio0lESDa6ag2k+h6O+PQZo7pt9JoUsThlPFL+C4AT4Tx9q6T
1JXv+BtyvP/6KhHF0ZjKk7kzAQLfbhOdpSSFPOtZ4T1nR8nLYB3kQMUTU7Pa
1xMR2wDFbz/x/djr1WV3/Wv0nJh+0VuXSX4e+PwpXTKmerrNebVyIAoSgpm5
VKdIcIUI3oODbS7fBks4lZYfKSQTr2XbniQkHYE0rF9Rm/TReIl2vzULMhfH
qKFWguwG4OZoKSnUc3lz/JRxVZXgQhizt8DaqxzGx5MAiH0aRxq+xy3fdy1E
JGDkK4N7qM9RVR4KsZ2xzzCZn2LIdRB3QZwUIWe/DSqcXydXbbE1Ku9Q+cmf
OR8UEvkGF7u4+Olz7cC2ZUf73sHQP6eILSJtbQ+Oa957ZZTt98n9sxtJ6rQB
eTQmHCh39LQKbX9i0yeVDfKfZQBJa0+BBqjITHDGutQZH5LtP9MgGgK6+D9I
MPaLLOarjvekac1/puLrmsUgfXggk1MDB1LQPsuaE9tT5t8sumgodS09x3Rw
nTUIndbKcD7yF4UYW24Xzwxre/5E9BtD0cobEV6mcdGgSc2UkB2uq22ycjXy
cvEbU1paDhAiHiXKDMX8YmnB0+m8IhSiWWz5Pu5qcdTPg5TvYreXdGZCWqNx
4I8jA0XbpNtN9nA3ozYDTlGUHb7r/SwxJBGmAm9TCR2OdhMyKI68+WeemSHF
23A8ILctY9TCcbQa8qK8zfaHbHue2+oPECeSzYjd9cDgFh8S1r509Sn63lxc
pRSTmKwsA37wd2ipWIjHps4MvrAB3mXvTLpZTClz7kERVpf5EczQW2XPkhFz
O7Ab6pJmT/g37bEv+HrPAvIIZIkvNQI6m1yyHuWYYvgzxzZ41cBIhElztVu2
m0GgpBkBkVupQJme8cIMjg+BCuuqTccPr5psSMZ2BOsmaf3yjS1/pWfQTd3v
Vjoc1qqSOymt1usdGb1rSXtBRg/BfpbGkvvol758RvmZ6VO1J9t8g239IIXa
G/6/Jpp37ISmrnv1p00C8Yyd/WvOC23rT8EFGo1+UuZD1mcf++d/NZBpgVE9
+5RgWf5SuP6ADFpZmlGMAcTPst0KQvqTQuOZMgZ2rGAW/jrLyb33CI7pfRlW
VAGr5hEJtDsUeJ5ZFORBCH5VYLV+6lvUEwfbRlIBk+vWVZ6ZZX3YHc+0O7JM
NqDnYk1KkylMfnSK5NI2MtqvRq6M7FJF5NRuZXWXChNKEknYAjlt6oz9MkxY
uj/sixtirYSIH8SIcvdc/lDg4qGQERZAe8c6ONROUQewQsjsLg3K1qMdOgmI
2ktig558cLvIccDDx1FtL4AAHVfc2GHUxvqusLGA0uTq6teikA/G5SEGgC3C
5pXSQ5Vcq11wmw4dIDKj00cpsnkmCnhv42QrZ+RUiTk577ODExzSdkNnfoK+
XB+vi/TGLZO3uTBVMpZxfaVunPT0JIhhe9U/3upAu9TIEiznXjdKhIaQyAmO
hT+WtxLB5pOovwEt0LuYb+F0qquJ+5tS6B5Em5VRTSUunkQd3VSSoZkmm2wk
JQpUktRdaFWe6OVV5kghvzQVCz3UTS+MC2GVNJErh5e7RebKxt88GimpCLHZ
lkIC/fpqhrnXYb983m/9B/n+EEC1cQhksAKInf/fIIrHlGs7zVF64YlRoupO
GD4KWl0coignPYLvlcgtVS21MMm3yqgZakocivn9WihMTCM6srvK8w2xxSy3
etROif/yDacLwQxVik8UkBw9PS8TglTepLkPPtlwlbbs5wkHLTK8B3DB2WCk
RzyUG2/kY0FxpX33cCsfhLtvuyzvnb7JPNT22S4ISTnCRGz13FhYZBeLXGpB
x0qwOv2v2xYKzygem6v1rJOR6OENfKDxNtZdhB5dIeUsI1faT6NNnxLhKtwx
0KOGwZWV8RaITqvOgGMPVOzwXEOT+bclhxpq8v3q18WHs6IQ5ipd8ZBu4nOY
Tf64D683+1TnDF6ulEcp7nGXIsk5XYrwWf/KvQQuGlcUIDZ9PswoWzxIem1m
SPTxJ/xcjsIOPG9vRk61XmO5LP/egTsOWsFB+pMsv3JXG7u6WHMNohVosd5k
2iow6BD3Q1roVv07fLWemegk/ur/NFJI3kRHOsoTEVCmv2/4gp90McGcQPQn
A6CmzqOHINjoq+BLlAAavPlJPq4iQ07zfwftI6/OCP94ynt072OujBBGai7r
0Xkd6Zb0wpE+B4WYAxYtkakL5mj9Ai5NGfLnTvlyRrERziwHMDneb2FgG+/7
T8VGSxUYAzv1Y+NSYvGFr0QEP0+INVMf1AFpUGHp5C8vHe1syELnOQqHK78U
qsubMwi35riecOwRDnqABL/3QmoSRvCBPMqOKFzqHIdQZWG0+kXixj7Eqczo
0nh4R5HUarjN+UWL41cdonSyAmSHu153PmiMcl1hFARy4skhXzrzNda2bgWY
sszS8gA1JjpA8xO6ftrz1EYLi+cLv/S9oE+DSwyP9h4lktDqn4QKE5c7sECX
bmKqmGzPm4e0FhDq3vdAwEwLSQ/dAmStxGdEW+KaboaWtdteGsFG3A4UPHoQ
QLjdgWFgdTcS5jwn/O67/lLOdy6QT52JWWGUpbahOBxJCfGjN5echsJ3Tmz8
PAhvuvvBNMkJrSXdNPGYEeq1+1eMmXEoq/m7fCVUVApRrAmtu4KTyu2JlAtq
o1/C6rruEsIe1cfG+aare/2JQq71uNJ80jZpN5cySlV/6c03llG+HKYcQuF2
Gp3oE2Cb1pjsmdQMB6wjMZ8856yi15LO+RfCVrb5gqU5ry3E7nb78ddZDrDX
zlNt55ilQXoIqdpc2EaRnaJBjK68TXF8acNuASJr8odgYvpICUzpq7Cgwudw
4Ci1LFAVPY2l8yEtwfUg6G0mMbokl/xtCpeWRdKqMPVgNnqKBrfTiGE3vQuN
Jya6qOqYoWv0GSKQ8FE+TtkkUoGNOWc+oMYYDIgM13c4PuRfgvL6LXdJtO9S
rgdidYUZDHDHxk32aMGcGk4idVmPnOFQ7+axWYFfhey+M54f/ryd22H+3QA4
P8GTh7yI5B7mVv3gl70vzNMDOc4ImKoYpGURW+ZoS6nW/6ArE5w8ClYIsrYK
L0xTDiyB8+CWjTdRGv8OeDCtlqHd0QvSP5gk2q0ySdHCKkDveezZXuHAV1s/
HnZoqFRoqLpZYrZivqRm8TaFc2Y77mVpdWIOoVm/DLvQdrdCZRMTEnIjOFJM
vFNQ4goGiIBh/Vbsl8JFrxJ7PVjC1rhxuGQR7M3nhbi9jW8RiJLFV4yKCL6r
LdDPr5pK8iPi9w7vxpxDZUweLU7HuV+x1IIKi5c/D9A2qKM3kK2kIPH14gKb
cYi+eMTN2QNQxIlRAlBIwka6mTEWpQJiKegzZeSBrq88TTynE2Hh842XDs2T
dFIQi9TH6oStLB/JFiW5bpzJ0qEUX5vSSCdzwXT5lmhK1Y/X8RHbg0YkB/Ok
sKSE2gW0ClAArflTOFI4LOG16fq+lFvCF6ooCbmPS8aZAsjov73oF/Fh0lEJ
ADK5uWayclNlBrZfAKS3q/ijURlvPCtVPA4lzXujtdFaX+4rYEYrY+18MEx7
Dca0gCptX/9Q3FE5c/3ugSsNQLB5pqAa2ymAskIOP/gyQGQ/8O0+Swrq5PIc
gcRd4f9sT46Go3wo/+9p7ojA/LP9QZ9l+wHPRO3xIxyzoiovIE+fJ/e0Nb7g
eF/D7VywAw5ruV0V5xrs8DeCItyGZPZ4cZ+dYhoT7gaINl15WG4tSPPw37WE
WMYS3wTTiLkw75sIp4bLpdMifhT9fEPcFD7mD5HS3YELN5KCQgDHm1k6RUpz
/8s+zDAAb/GIJeaYPqwKm6C6QsKE0CT9g+B0Gz1i4HDkX4AMIPOdKpsi452+
sxIGPhVHlZmzXaL0a1ZGqeWAW5D/+qhAd7CPJwJBMoxg0XN8YiytdZ4mMv8w
Z4drsWi7gfSAF6DbK2s9jZPkMgNh5fnKmJXed8yTuk2NOlh4IBM0g5JZFbiA
QSTCsNRljY57Z4FabfuDJDGUwhZLPxPTXlHxbWoKS4KiBX6gm0NF5GM9jv5W
e9HRVWDr9rYX46pYZHjSIut9Man+JShF/yDOVYQ9m3q0QvHPW9PcqvpGiEpw
0ia0qgAbXag9MM7BCcqNZXCRgBwZzr08etBBuXkde34jL9Qugid/MSTVdieA
WFxNjCb1GuqDtgx6qJ4f7FxPjdhzcKq7k6AyartPiBd243fyo6GFjRlipK7G
3Ev/0n18gEgTkSCemksshUQ1WqHKusK9D5vb3MM/O0YjEDrCi/Y+uo8chw1p
Y4+muLTNO88zXFyotH+6OqTFa++xPTJF1bYplgZrHG3Q0YXbuabRw+w9DtCp
SS9bLJQn9Nk/FURC8vMsunlohNmhnw6YiicDOa8catOaLSLrkndSWj3u+714
XAFb1S+rC/Xlp42LuBbqaUNIJlrL2EJlEiHGTTjZDREPZHY+rshYDhvLNpOG
64OcYn/ksKLSGR0mfE8qsxdPFMda+V+Xq9pC09JLP1KO3WQAS8UOs92ahanA
yvX4d/4QWTQeurscTMN+I5YZXt/WYDq9QHjPvgAk2fBV81Zv27NzwRwJBjRi
+r9vJg4YUkmnT8ZSsaeyz0O4iBjlqqQ+9/JbOi5w7RtU2ioMUA8sFhAAyLW5
swe+Pj+N1ZVQsAduGOEuvN229wAOs6vGXtsgiRlMwxryZTJ9RM+UA3Ojd067
nivILPJQNGKaZsQlxtepNEQI8SMl88ArAMoIDlLPb5/Ick0kZQfNth/PK1fB
esIWOzlBThzJWjbKJ1Q1COib+8DWKEeU6aX20KPP+LrIuY27NNyuaL9HJJUO
zxP0+a13oQF/ubD3AZk/qcbR5LHjK2ZNG4VJR+s5Lgjk4SYpIo15ZHrjITgo
gJj8e3NwzBk5PD/9BnJbcopACNu0UedNzoPXd8aCOPtgU9wbi/oiDFnh1BL7
wZNPVvqMqLrcm1zBn5fd3V4QKmamIe+hgvZwuUFBj7YdIKPEQg1OERXKMeJi
X0l2/kel1MgNaDH05Z1XF3D5drYaE31ALlcO6f17fzkLcPu9CzVQgaarNZKc
kS8C2JchrWp3aPFkiMtRoGVW7B5v1FbV/og32xv43CZ9NENHp4hZm7XAuUOZ
7ft1oxXlZZS2q732DFXxjEsK04ub6s0sjxR3JOzlUrUBQmhAUKuFzxeSw92m
AnTq/nDRpB3eNcECOI7kL+CZMOrNyi0ielBkXWrLTkvNsAuK+1CAwYH5u5YI
CSlUB5DFlpF97GFnut0fMMFclYX9Ph7IJ5m8HvZnzmRLxeV+C9JconMNOTBm
lZLZ1eAfJAyKQRrmjikiLFkXk3ISaqJHd4UZeA+hEmRXbJ8P4QMj/tALrKwR
oayolqX7YCoizdcarWY9NYcad0MNwksoWBNJJxHaLAPLFLdJO+h513S31kll
VWzSswMTjtL/jIlVeD6WofU+CFWVs59N+kZX9r6MCvtkDAK7AlLa+c/iKwNE
CM5x9XQ6r3lWPFvgyAnFhbJHb8GogZQgFT9muLL0X+hqwXdUhOmMR6xWQqGF
iWvwF/fw6AErDjUcMBHC7R7KEcKnz0gOQv7JUSETrCFDFK1KFxo25FPTWpUM
K40Ymu51OamVycdGRPFnKXrc8HpAnjeDU54ZSnO1HbiU4cPJTtjdZJEBHPsl
JSqouO3TAhJVFaCAITa6hPVkdJ3PJvn4g8xSdYET3OlJQm+dzvCPztT6QU0z
2A8YoGfQ3CEIrtqi5Ap3M7o/DGRSWcGRtZhvlG2PuOZ2l9jdAj8gX8rglv3w
0gOpr/LPQO6PvgrP0d88NkWuMfJ9Gy3kYFs2LTitwcd+Eb/PUjQKD2EU2Lwo
nx27vPn9ht34XY1EVGrl6IwmhRtmRTqAWSLNEcNyBFekkLRclq9QZzVsQ/+i
h3pY8aGnixcGQn40vhQRoqONXmwAqswI/dhxrqcis3KnWfeqjI/FFhLFgHuL
CL/oydaDQ6JMgZUSIgTnRNNrPZ34yKhMoTFqtttI3SSH+XpO0NTXK4CmN+H3
48h8bRb8BYMDaIBzTjPY2VRSED8vxURRED6737a9KNnXSNrr/Mq4wRzgR2pk
PQ3sYdH3TwANNKy0ykdDz6Y3RzMoSHBEGb7x1uPXJCp3ExYzp11qaUDCSNEq
qR5mU/0hRxF+oYdm7bcTRKyCGbEZ7Kwf1gsdtH1Bx2md6PxH0upRVGM9wwIh
T8ZxHQggXYHK3kPoU1P0d5F41oQ+qvDN/wTIjEeKWISkxmd8l1kmiN5vqSvs
aRbrf2iBdHlmOQptJgypdvKXMmLqYpMVKGZAWsI8HDJ0wW2ZThKHTMu08Fc3
GuoAH3OL3+9bnjD8MsQDKMbRB+QQvqqMjIGFINplnsfyiJz5kfq5hhrxmoQS
mZdzg2iefeWWo5isUw2PRdAxbzSADhZHHcsA0WX5N7NBoUrj6QFOqYVRdb0K
F4ZSjaCiL+keZfxp9ZFkyZBNndgA4Vw/LfT6TCsQiWDwi+0v5ukhlmsq64HM
siVHQhEqfgTzofSC20O7xESNhhIIVCQZie8xJX4P0Mv+Saf8rcio0KZCNQEN
qOP+xwdVqxgQWb8ZE6/QErj8L1C4zmhTjfcuFMXhamwX629uS0nZO8ZfKkBV
O0ItSjpV/orLjYmptS3nPMNuc72B2M3T8W8Tu7ctJU7vinHB0WOVVA7cb44M
Nk74HsaPMXM2Gg/X0skWQriBL+RLihRBydg7s9fFOVcwcL08J8gI94pPhMgz
kszyO5YBLL5uILajshv61vAbA/BTzeKNkgCKzaMjXUVbuzbDwVBFgnsBu0mH
1RoeUp2n5Su43Musql/GVrOzfa4uk/YpFkR0M7x7v0X/GWI325yT6fNTrO8I
NLRgnWOU36YWsGHc9lyJwSJSU1dVT/+277Ps3G+vaOqhrBb7qOj1kMvGYBdh
W6KgjdLaVSo89D8vSUUQfNiee3u0liORoJl3HP80cNwIVoT/3othMpsbDSlA
LkLW6KW7qJdv7HWQH5dWGHtz4m2eqjnYZPe//ztZPop+kpZLftvdSF1TN3YF
/l4mx/AVtB/ErgyYmV/aW4iMvDvagaKmO9AyVw1HbNqKkQWC1z9prb4Fy3XV
jVIw0goJbYi4+zTdXCe3yCQBc+097qEJzKKD11LClUCkm6bi42v6RYdkmlyd
HCocSVvjaa35jgP5s2ZVyPgk3qMDUewGjX0aVs2GKQRway1d9hIYuUhl/Jvm
jwRIijX8vrfmSWolDQHkDo1W4BpATK2sjlEkLYLIwLpSmid4jzULRk4Iu+n1
DSrW0bqAtIxQ7boB3hQFIOVCgGLe5UrUlI1mtjU3jD2IsedfBscHDdmPXdnl
zTIKEprr8iyfw4DppgmfrXXL7aKimayZrTfzKgxbiYlNeWYzLwKVCWomrBms
CGdiwP6Aqe23VUGYxRkoMBx1UDTbluSl57wqNwuDghRNISsTQuoDAV51UJIe
DZDrrbhCWn+2JDmLz1VMiMzIdoHrR9s56nag6l+xwMaq7q+feqIn353GZKyn
XxWeVABg6HdL6OP8lj52LGJjoPJrbJh2jU5D2gWe6UUe9fmVLOXPA/Zn8LOU
MeG4NiQmsZGLqMlaX4j6qt6xUar/lQXcSH7QlfZCwAtheQ1OdjdCIyBqKlqn
X/c3cCgpqArkbJZWRtZ4XPsjNu5JTpzeFUhSp/mjsE+jnCUJfzuBGygXLFNr
WWHcnBmWjltEAOYqXZr8FfcpjvrTm7YIy8aC1ftkgTeLHO6z7L3EC0LPQ3fL
AMKHNemOOqNJG1QUxYaB8jRvqMUnEDhl6m/aobLrVy3wrd1Cik5XJB/QoatJ
oSWNDirKkgNU8RM5frAFCsH8Ef9kbjcVggnTL53ik8xiZw4AB3AciiteUQgs
8rac1ZX7cBeJGMAwsqaQed4CeTDcQ/k2I1MOx+gTq6fhHpQoicW36BEDpPAO
UOibtpNbc8IaG6XjYFNteXt+dQGjBMbcKLqKYX0SOtLAntPzZoOo7LF30J/x
+M2DEIIHKpfKIgo6/9e0ufnjhKl6Wa4cnF9uEUyqAui5jYcL0UpPDUtlwbYj
ZAPSznqZd08u28oqu0j7b23f0DP0+p/v6q9GWNAFlQWn2UUgVl4sH3xENJ4V
lsBIFaf1Piv9jLgBaYJ48QhkG6dxBb1wrTlkWWq8mslW895SeObCHdZppSc4
dyiL8rUP/K1NSwiIHY436U3t2s0rwzB2gTb7UWYrmTypyYuk8Idz9LpUAXCv
f8EzW368F2P6vZn9dzYHUTQ8wVOrZdL8PA/pU3nnfRCZCCw0gA9QZIPSgmBt
1xQy2pBd8ygMAOofMgvOvhlomhO5XBYJGP4evXeX+8tz+fVjRCuPNmx6MVDs
RUHnUw2Fyfw1eqammCMscdVrAbp8xQBbiznVgkXVTkJIMPnfUM7ppa4HyXZi
hsPaXl9UMKaVKQ5S/e5ZB69/1uqG4q1mN5WlyRMFC8p0w+c4yonSd32hQi0w
c+0yjXhKGW0Zp7kn5/MUOtmBNHEhnNU1WUlBgcr+SmxNZkrB1ck4JvnM3acQ
sKXtEc5HjHReZLjEG1iNRl0+cwGhvGitiZBnQbkGFrMFYeONMywj8xbSCGRf
TQ8QPAoULQPYM8hRQXLObC6naXxfZfKZJ3/cTtfNaQpH9X0GakQat9aK7tVm
hZ+MU8iBq/p8OA4JSFytvOMAr2m8521VGgg1D71i4JIsg7HYoNMwMiiLiHYE
Ug2Yc2yHufquIuMSk8Jhlr9ma2f24yE4cA0cukK9ZZdmyPy7Y+Myvq0SrkcR
RWog3wh4YfFXdoC66xAm/IVguB7SQNubgJaYNaTuvIRsCbo9d/a9HOgrKfJh
DxUTQ116VnknZmtnhW+68CgJDaa5dvJb8Jvzf2cGIdUfJx4hJIR+rL2ON6AL
2T3ZHI87mmqRyT7HWKkON80hDBS1sm96RFzpKVWaVKUM+8ONSoy9uFF7kuCn
399YKfATxFA9bpDm2R3E4OPdMaSI3hM3EqSXqT31uw8ZARG0T6T5biFKekBp
AHi8XGwRzdd+SIMaE6y3Hre0xa+8u0bl6m4yaLqdMahqiY8R/EjggI6Y+qGj
nRW02chV/4/+I6OSzFt33R/l/itendlkUyFHHS1SglBI3OEI+2hMUHdd26Zd
X9LbQpgKtr6WLfBgIGdyUa5AWGIz7T0ljuwSrCJP9l17Anz6TGNSXSiX5ugR
wPDfQQnohPo7r9YS9PI3MKpKB7d/MDBBkzUT9Jp9/ITKAAuiUo0emqQZp+4S
/G+V9kpBIaxLmsJwZuvQ6AlfkVXF7dVzGVzL1hmAGxYh0AWqmxku4DitM0qn
2R35VHpV2tTK0+B5mQtaI9ua9Th+rhMQoVwyldaAQkSeWUI9yxl1fy55YqX6
oVrCxssoBQ8i56YhSks/MqX4Zaf5Oq8J2HI6zjM3EdzackstUSEdeqzR/yVZ
RoIzKQbbfBbx5X3DAXWhKanRslDYpIKJWbLlQUxbjyIk2rJGRNrgwhyKaQc+
tKabApAY9vzDFdYEKKjdN5xPWz1SSzWefzcCGR8B0IUGv1kzlMn+Nj/9HIDF
zsNs2aHADbTuA5/XN3OL5OiHskULRHt9qRmAuU1dm7t3nC05MqwPH11dH/Lb
V7KnPU11y+NMez/urct7FJVksvaTfmpU75SpOMR1s6Pg7st4/kuQD8EXC+J1
QYSNC+StSMYWu/jqYFks/uQyNKBFHdP/F+MwXW0ZlytS6yfsAM90OlDxoInW
+9tt67ATNHvYBOkYp8oHrSVyG8U+awFIcvhcSU35C8kBDLJl3ENZmhkSYYpd
iGQRnl/FU2zSkYrWXR2nE3X3ve7D9e8jK5nKrUaWMZHzLH3au+AkpGpGd1BD
gyRCn2QVFOTGF1SDpOmQBxt0WLN0X7BD0YIdKUxL5FgVmtCcY/iwBCL5X2jm
YEwt0fU43wgiIKXqZYjB3Wfz2crJjJGAXAV5e9cv2/B2TMxgk6gS0tMDximU
CPkPzuMWcfwFUQ5fULoU05aMZUZ5UluPy9uEDVfJ9r50DtNvfoi/m2WNOxTh
fBDQg6zVIvhw2+cicKxy8HqpHTHZsJuNASFqbHigBX9r7ZvSYec9XkdTPfSF
lvr93TgSWy+yatHwSAvEa70Jctj3z0Sz19JmUUN/31wXPLERwLokHP0JQQwZ
Q9j2xgu9he3HfaF4qSXmIfBtrUYfNpvpWqmw1L9MKyMTpH5LKzzFiKgWraYp
dkpOkZOWECcWujDFkRpUvVKDFv8fw5a4BijyCvP7Jktrn9Q0cgsTVe4NiuDg
78L8xD6f/p1R+cu9yYdez3hofgC0sZiudjA4+Nw58Vy/EeCPfSvWjFEKCKIz
DRDWovI5GWbWrqaCDwuatVqgL6AcBuTtCl1/nrgI5WZDj5yHhqRJzWLjbnbj
m8z8nyk4JQU7iTCKBim6butMXQQJEbmW2TI1SSwgOJI3LiPl3upsjNGaEBXc
J6y0eNcsoTo/D58oz4g+yiMf5czf4lukD42TKrbmqRFBHNPu/qOCHgiy4JLl
V2TmDjS31n2flm5CPGP4XLhfQ90NRFMeWL7Hvj40L11P8Jfn47A/scC63JtF
ND8Xpa0FGs+Uk7Lxx+Xl6K+P2c8Q+pCqoHq4+Q2l/beIcz6ipJ0GldeCl3hC
0ApvF0DhAavDvJKdGcfAAYAgWvP1vJd6eRY/AhusSD820IHtvyNzJ8OEspRV
DSmhXZLg4g1HFs5/bl8hELf/LETcp6htoC4qB0ZLcMjHW5mvMsULwOf6nelJ
asrOQl3jj9xd7yPeOBK56DyyAatLjyD86i1LlThsO06Y1oor35FDXOj1mGD1
CuJrfcqWGK9FR3jdC9N08fwz3ssgKoEORJGb3UJGNKcdLirX1aiPKAS6SDAO
OpyAvbLVVACZQDOV9qJ0D55WID07pi/9BeMJi6yA6h78z4P6+/3jP+Bys+Kp
xZFwpuIbql4rJ8zO1EScJYhrZujLXu7vvObp1F3R+wBVCkGJlw2Fyfrjfn75
1TGvG5BcJ+4G8/RcuJStGZrU84zWpKyVpvD/KHkPjH1NGWI7Le0fBPiYAijV
ezC9JmjYp8Kf1SUOjoZnrQTsts6IwPi7l5JpJCljgSX/y7n89MCV6QdHsc6H
Z7myQy6N6fXMXc40iGBwYwDsC2evp7KJv/pyQWcR4RWAj1YpCAmDYsP5JoVO
Gd9h9vAKGEzztSfsLqKjU2b7/R5+oFdBciO5KtJPl8E/cV8aNShZUMJ3njSM
J5Qh50lbBwgW3RYJ9/36TJ5x6BSY/udhURnS0FjToFgxs+gdA1pEA+LM7NDS
ipn1XrYQiWqFCY1eQozsIDfMnD7y7yuyrmdOLg3qn9WLLi2/P9P8luQhw8ZJ
lPPEqCF9IapfrqcmwDcY4RoLiYMq6yh6ZnU0fhZORqD/Ct7DIuwCGvVSunr0
ANiwFRtKD0+jOi99zMeiQOJXaltdRcRiQE5yjwfOu3Y5LiGevVMx3UUI7HI8
TRa2oPS1Mq3su9zVRmqSDkLJo+2ds9tLtD4PJlNwXaqFegYhsMPN+IfwVVcB
JO55Ikdxe7ji5LULo3i55yYHSNjM+QCx+QJR9RZXtbl8gNUy6HhOWj+wTdf6
fbbJAhSZj2iJSulYoqn9GWRa0kZPWSFx3Hjz2pKBwIxCAeh7nlY8y264auM5
GFUZYBWIXV/NytVzS3M6X0f8D2AANK+zwTWAfIOvUCxQ0zY8KV2SzVh7Ji4a
axkAK7UY+K09Y33XiaT6Xp0WXQ9zyR4Gpw7UYZyw2tqbuvKEbWwgiWh7eamd
jOWRj0zrKKlJMIrgh5ElssX032S2wclflbdGD8A1oJXRqvRJrqyr0VSEzT/l
UAmVQXc3mfYe/0HjvS62ynW4gPydRhe/W5jClz5Q66EnmkVp/UhcQX4uEpml
TiN6H7IAbxx4+eNrf+n0z/Qkg2QL4hGazn2j8P9zKWpuUH8mCjVTJ/lriXPm
9b48qj4xn07WahRqEhDFSoAsKLndI2tKOmClcnjVyIHvc9DkHbLbe7Td5oSx
J8G+vwaTmBH6sH4Ktr2cdSTSanhpUzlmA4XpXmpum7HtpR3n6hVKjs/c7u5T
u4/kvUsVaW2rYiL4WvQeSnrf2eJOheoMj+8jOHOvbI2306kON3Fng446isCb
kItLcJi23VJF8ACIlUHsh8Bd66YRGqKIOtZz7sIfNO/25jdXIKRpub6XviuD
HFasjRj/n2yoDD51/QzLB7g0EfQUviErZENnG4KlvV4H0J7q6fgk43EQkSjM
YFvEKYA4gCrmny6vxmJdD/HgrskiabycXImDA1Rr/9NORgyC7FqQrk6Ee8EM
XCWuf5yz1Dyzu69ClnfrxSA63gIy5iNWijkodfJTjAwQJGf9Vl7n27zAHz1X
RYENNJJNjFa1tG1d5ZuRHxJFQIv26yqacNcD8k1xnUjbSpuutkBjTpAD6Pb1
eLLNhp9zg6dBewueqRTYVeVOGdYrf+bZX5gvGomWsBIte1zdzwaUs+jL+F5E
3WU5kW5GbnfA3yxjKXTUqCxQqOjIX6OSBRFPWX0qVA80avSyNHzI6n9aW5Qf
f7oSDpqgQXa67ma89TPyrYHyAbkyIX7HwngAc9tHqbXp+zNKhdyF+PsUfQMQ
fxGCcYQzRiS/c4hRI4ieaA7tTbMA2JmWwUic924ZdSWmmIPXUhe5cl4XaJLa
BbrOzL8zXhgzA2gMO20G9PMWmTFYdXdNEBV6LF995BF7EmkoNL+brM7AoDPv
EXnKLuKlNO2HhGA2XuV0RkNNSmL81sS+JiLE4fvwilSIPxJj06V8gB/y8S6f
eDyvBMnrEETNDD/acS4oSudM0liPN/7uFRsdQRBRdGMDPEh3Uw3tjCHHkjtN
Ks1xJ1FccQgpXWKpUlFsZj0B6mRw8GNqHbkhMlIYBsl1d+3wpnVZoY+jP+wc
SS7qXRms/F5lR0uaeCvir9nouXyOpkPLcIgQs6xyYS3qxhQJf7ocTmxNaBLt
nlJxNen1xFvzzhAkKcfwX4HDa5SU+uvBioTjz60HAV/nSj/m6WCK3RUzJT2+
5ePt+NkvBxUZ6zQMykZLaTa+oVCW4hmT5VNBa5gRGZiUXUIkC0aLCXq3ZWIw
SrquARNYdEiAKfUZu9rv7C1GstjE9Q/HmnUA12bIXLms5Aj5iDry2wQ/7apU
5XkSkt8gbXTZcyDOiR3QWyhXP5o8HL3egC/ASzEE319UsQlgpoyDW5ZDfEZh
mp7VMHVd/hgqvj75u7Fn214cmPcF413kW5t3LlJFH1dT5DyWWB+v9t85+BL/
A/jmsU1jxFhjROtaogqTqUYHuFaQF4IholBuZ43eaJmOIC6ws+CldqDuie0Z
NDK0GsVfyG7Nz60mvBPcsYceaRKdGOQx/lAzz88Zv2/IMWpAdlD/iRumjVzQ
OnFTyqZZzkRhsJm6ifj3eOmy+TUs/rGz2ZlsfaHiPwKdh03xLmrafmgWOM2t
+BcfBrpszhNDh7OxgeHjE4FG9MR8qt0IoU3oca5AFcMVRJLbfQZq9PUOvGKe
5NEylAMck//livhrNdaxgOFgycMibq56kniTseF6uRd/rjx4f648xohEUUz9
25ppFnRL5r2+BMAdTUDZlo0euqCLTi6yJztyg649SDTQcGgJECBmqk6ifz/3
KybhM/rE6rPSyqDIIKOofXMNae+VHSWy3k5nWlkzyj1/47WgYV86dAK5731f
IznF9dXzVRwiAg+OFJ0FiI7j/RBNkQbKSi+NIKq7ycqax1Zo6v/usdZbWajT
mMtJEXzEc0cqAAYKXibcLcnpG0TASiSg1nbxPlvIAtRK304i6mGwNOS5OtbW
o+k340XO45/587YZhKfcKxU6pTQWGKlE5hYB1Hw2hfHTmn9bhMYDBMTsBUGz
+A+bl4ip68cEiCLcJxK9wgGBbFPv7cIKXlB/OMd5UBzzNXGe6x3i5otKKgF/
WhcWXuWiFbMTe6Fux2VURLqcBoesQ9lWHJBrRtRsmCEaMn7n7ukNJbjJpPOa
+t0MQytdJgA5bCA+dw6oKdufmcQp3XyUm6fLUo7XpfJvWjxP4eOhiFPzxDDt
ieGPXhk4BHYgZEbkDOHSEF1fBRZ2yV03mFn4t+kwFYkpQXm7MrKJgqSHkwfu
AXOpvmxUzsUAt3VWmHIGyLx9U8PNDOKDzYvyqzuhG+bjNTH/xq12R82sX33t
LWNgRDV2qRzXu4fwN6TzTZGZd7wdh7toNufepEcbP8Eqomtn8eiT8QWUpLc0
KB7MN62kniZNndKTpoWTDrmkWKuglVS65PisGWm/y24osySH4soLtxX4ejeo
jX6DgIW9f8OKTSdq5G1hOq1kCmhb28VKzDtjp7owDOpYsfcZljip5d1uwW0/
M+GXSyGWKejGSkYaSzIvzQPs9gwkKInMJe9KaOUlnd4sRf2bSts3OWr9iVTl
EB3xe3gmhus5SoKoSZSER0TdTWiQJUgbno3yGaCnetC+FeWkZK6b1HpV8cQL
f+No/0Bo4nwntpTTHWLSs5wqzotN2y1K/R7PJ1aIoVzTyOyXvQ0SZzUKUkCa
fY1q4I9RSG5z3M6qBUlXawifPG5SYuZLSHbWpcWLDE9tTEBjUgGUdstrh11R
4D2ab/eqX22Ar95+xPK7QEFAjiowL8gLKfm7Qq6KhDJEWVMcg3YfzYVbKuiA
mhUObqWFv+2p0C257X5IW5UhMWWhs+tQ67B12XI0+XoSMXEJjLr6pTy5udvJ
ndmH0jP6AZSprbpUTHCdNfVfp6tElJKuIGpe2yc27dN5i/mcJYpLddzu7nGl
ACnz2/RvgeY/NGbFhqbiZR4d2JMIunL6cUe+p/F4JcEfpMXH/hFDX4JwzlaF
XuE04SX0XAZnEhdQWwBuP3rHSTs+rOhxBH1K57ApN/fLJcSX2aoM2J5f3jE2
YhspA3vfu1Msi0ZmFaBCG3U/Iw4kFawZKXixbFeVEMhVMpvCKUPevj1zIv+U
LW4oYEb8mW/QPiiRYSQQaL/QV1u4q9rez33Nx5AeZZVHMdGGOgmC2BBRtxRK
IKO4eejwPMGqH/E9kpU4NHNVSlqeteG1QkKFzau45dHOcJndPoFV2h9l7Htu
OpXqLIjC31YG1nQmJzXNuV16PrcZazD13TDd7c1P+e+YvBSnzkTbUWixt2Zx
uQMeXKgGk2QyVetqiET/vuneaX4OYLlqA+a6Eadwza07Hb5vyi+LU4BibG8f
5NvOGYg5HviKUxLKif5IwbShX3zQrETXeizUaR35dYDsvi39ZrcKOs0A7DSF
nV0IemMDyIXTj+ZvKkMF7TU4WYCHKOxXsOyah8Cw1iziWgH+YsV9WJPODn/J
2N6JL8dE3CCmzpnSI+fJwo5UiPcgy0tro8Rpjyd7KPcLoCBHHDlk1ITxMq4C
2NjEX1PCNq2l67I5BuhpOUwwnuk77fOEsFx1IGlA1hkdFLy/qHmi7/JJM4hO
I0dT8C+IQTZcIBoVAILsIK1zeGdLha3+Zzn3nHVsWdKbqdchrP/CyBdYyXPy
BRSZfugDiPqNDxaOQUlXjo7q8cPkwctCmc+JWXhST/TlvMhPBNDocJ0YUkvO
tFg4SCjpiOy+aZwPlE0BkC8rcRA99iZqalaanhB6WT25cBEnMkOZz3ewuTGW
nWcHWj9Hp8wcYIFJHnvih7p7eejH0BHXAB6C23O+1aOA5QMGxnjrD0vpNYiU
U1vJ+WdPY707s0S3Om831xnQOLoIGYkvfEzBTf41lFcDw4gBpixljE0X1BjM
WoDfxZMUEKqh40sAFP+JMEbwQMgT8do7tqj15UAzm6jhKTUiXPXTA/TzkIXL
v9Y5hlfUaBCBM5ntfsz1HwRROQa5MQ4SOqDRtUHxBxck4WbGS+QW1qaVJavO
in4nesxOTQpRgSgcgUg8mvIIbPkQACF+8qPNj+WpWcEyVpeVlgfFd/kdv4lO
pQZRShTmSB0t1WuF52+NrCx4HRynRp3sC96LtZAvMMZo+hAMsj+ENCbP39Zf
IpfY6Dk49fBmCGYQ3HgIHxW9Zs4/kWz6ZabimOt3D7qwf5FV5mGrobDaJcEv
ts3mo7bgHhmlMadPPY93YdKrtto/+Nt/cWPEA5Oup/wE03tJojiF7EOCA6ml
9UZ52CTSXt8udz1IDAJDeaiRrSLBBS0+yoGJThPWODkVH3Z/VJskCK9VhUbD
KL/W/GxCGaSD+CfjYAcehqbweQJ9g8QvO+YSY8WZaKaZz+jDLLHLjwGwF0hC
ZVI30d2NmJlkWM1Y9OHuwfL9wqIcXMomCwvuioSoHTheJyz4CdRrOBzwD+az
ZD7wKHfwZGhbs880CJkQMDUkegAJtK2H0S77p86m53M6e5FTadZembERTKQ8
oYgixWIGsNlOHlkQZFG2hzzb2QuG2Yrh3DSKfMI9ongRJoAySgWMNiRCK6TR
FXNr7Q4rJG49bfBmziX4VH3ciAeikxVVJvj2NBaxYWbD8NV18Ylhnh0DhaHy
BepQLyp9hqxXlrGRvcbdkSyJYgSlOTgQPHzjoLeKDMcjmeaBOXg5bJHeQm2/
HIFdm04s0oUVIYuTpbGEPYC6/75BbHUnbzwUNEPJmBmnYeSR+PuY099SXnml
bwkLSD3tTkfxhW4mzB05Wii9Df/0er0TQoYxHZ1BM9OchN1vsEK4xDoQKKrX
LOr2NgJsgQzXTG96TIA5Q+SsT8GHmy+bxPcyX+jCSUBBgAk8ad5hjj1VFXvp
YFvaGYUy4M3Lli2UWR3cV9l+RbF/hDEXQ49GHfP8qY4j0RrzJ4xTy/l3sHR/
tclHnLfo19mbRyCu/bLC6i/voMBjeqtiU0dZHVIKNOgYjckBziuJpIvwvWnJ
1do0oYiKFcHcxNaHfg2/J2JkgiV5pLSJhClyuX69qmXm4V71GEVseb33DLY+
f0OmGdIMq8Qc8RjWzmBJwW9rNdOL/iBlT9/0u4zQ9wqKRbqUYXJEZuFegXeg
hACLeQ8/FyVwYDQisSrBfhK9sR7lyhNAnbvtGZbR7nb4bP2GwhByZT2tMewl
EbL78vISnFbshMlFzRtRtCRmb01/DMtr7Vo/NTgwUO9optiWTyH/kO0rIxCu
HsXkb/E6vcTmlZWMlFHIMafCNBJoVEa8a1cF3URt8+3AlP0xWuyUwwj/Ryuy
2NZflIM2LKQPxpKkHzE+nTTN6IG4HwJvYhGv5rrQraYM62XN94r9ay4wT+Bi
TuJP14wwOxwRHVfOHRGt1ijnHsx3Uqwz6qxt2HRn25tnM37zDWmCdeKT/4Cd
hBzAbp2pvCwwVW+JpNVqpYWCQ6ZYVNF0t6VqAqxwlOtPblGWEZBX1u+kj0KI
VlJ5Z53qIhh8Ch++sfUfasqVAgjaz0rOpKt0cgjloS4q14Qv15wzYhuLGJMD
D8ZCt4mh0kx9fh3QpP7b2AMsZ5sw65UZgkh7Gw9NKJdgBdyZ1ayAbrgXNplZ
aovPI54Bmv8n6WXjAoLWRCKQQS+Xz4kMFOq10XbKiEqRc9GPU4nz3KdzLLVK
PBqBB3LV5Px1DK5g9RunpMAR8zR7nVLGSQEZIm8cJVtyiMf3K3kYEKxEMTKh
LC9kUUsqH+IBxc940A9OIQ1rHrw2b10VNhinDAil1ToadPUKi/HzIjtI9YTk
djFjOlSPLOLhfgUze3PQKKvsqlek59H8fdVAcwuffSzkWx0Ljw6OjMDLRWxV
OOz6l8KUfZ1PWFH/a2i14odc0OLVt9vTQhzyaNBkY03dZB323jwFTXqw3UZ3
meuJ6cb5VSy6z3Ut9DOGqzQnbjpeaJ2hBL8DV5877NYR45tjr1EKXPehK5JX
sQ0nFEpxOKBYMh+jvdhbKV8hAbMr5B2XDetWpgghTNGdCVobQpEwlcNMhoTH
HfiMboUHEo9mQqjL7P0BlGdF7FRD02fc+R6OEVb/k9BxRM4bIIdJNOkTbJUL
ZIAhjfwDopjGauQRSiu8dDNF6vjsWxf/gieL6ua8lpamo14f397zqodte7+Z
TTaTxHsW0WSRLDQv7XJVs1WlPxq1uLVnr6M2nUwKsqT3/KHFiQn51ReYNZte
xNkruoBd4fZ3Lk+y8vMRKv0+L2nyPBZlGwTpavB0L6YXplEqFpwA8yh4rVar
Ttqr3xrbW76N318Hoc6MIPj+3Jpi3oLCgkbpHq07bbM26GBOZbjAJMHYtaeX
Au7VqdZZPXzaL/AB+QkR+ajrFg3hlf7IytvCEs2hJP/sKeCgliA/X442+Xkd
Ss4DsTzo+O5U8e0XesVfW9RCwC/xNXlcu5188QBgPgTEKsxHmbcihIGvjTFT
6oWeSpGD63dFNszA65FHd9hpVqEJZ6vrEzlmm21QeI6TRxRIcXv119w+zGKC
Np8D8Oqmw6+LFxvC2QRRyxMHdmBLqdPR6JBLPgvW3PV1u+UgV/3BuWe1BHdO
TAZJ43s8oko1e1tAZROei7uckU+UvUG33sVrg3X6fDL7Pe1KUBWHKtc2OOCB
7a4VjtX1zHWhnsqiRdeJgrVK4a18j0Ds/xaRDgwy+mweKAmVG1hpLb7mu0Uv
xHtTC124uK8EqD/l9SZg9fBx8nzYV3sfpgpzEp2yMh6gYZyEFBtldakB+9o3
YB2yO1iplJ3K6rJA2UMo+ecMGYzB3qTQ/HS/drgpowMBjW0WKbPBM10oljXe
KT9akDVjFzhYppMdUBDCr26J0mEym4iivo0xKtnMdGZSeCyhSMw2LD6CcUW5
XUQ0JqTeRN0iX6IU4z1Xf4nF01gwX11bklIhHoyG2jbnV+o5adgcl0xgrBmi
5cYTcywvGzPmT3MKQJnA5EVKZ+FdhS1L1wqBE6k8pKKqK4Ce28rbx5ug8d24
BX+og/xuzJiukDgTg3RPRapmypUUUuJZi9qRiOTWbTRJj4/NZjPNVYXy8Mi3
dHJ/fNVe74zblWu1KR4y9N4gg+I2EIKETQsd67SYs6r9csJjCNEu35kcld7v
fbb1AUJStoMK/ofb8KfBxx4TuMUKnvBq1f0BzRwkqRAtBjb0U49d6WxdYRmn
MYNDQriK+sDqoMt4bsBokfDnskHKVczoouHTdChp4qYOLeZne9QsHWtukQiM
nGzRy/f4QGNDdiBt3QtjQSUfjyclKZMUZBodxXKUeJqQx3AD5UMQYe27OIDY
GFEB5nhSjsTLcXzAxC371YJIfGM+Kb8/fPWNVn66XVLFNMq9+7OBSCWCOXX+
TG0AGRDIs5+oDhnTaEmDx4TGuaoEv5pdgUO0orrr8MA9wIYRLswHiuIUqQA0
m5wS2b7/cxS0PjPkDrhZT+KdgvhpEYi3SMal9G4ptuVPRnf871kXrUO121l8
KWa9gT33KFfgk5CYbHhY9FrFbPoCH9AP/KfEHMywDOZHX5ql6m+CNP83WDTT
xxiaTdoWBD8AvPbYbAjKrPg6YDY9iVFn1DOHcKfm0+raUEteuxcHVupuJkAk
nR+EteZWVLfdgGNxqIa3CKspHVglg4AQM72iUo7yrNNUotAsb7M0H2VKL0Be
RBGWhGXQRlywmKmCH53FF2R/Dbhv4fBlyd/zNmjmS868zqHMl5tUtyxe0vsD
ytu2XQMNOY0zGblAWE6U0S58PZOX2AmkXowEfNAJO5MEoF/mRZDQWDgCPEVm
C3xfs1WssO9ayp3p9m6hi2/2y+TLXYIMws+iqIPAa40KTyqVxsCAv1urpX70
S1if+LMjQt1KMu5AFLhytNSmUqkg4C/LrcIKjl8pxafrZwp9A8rzvsfkbRz/
U20JODiP1iTaLBWHl1ugj/1ZoiQ8LBxpDOEagLADLHLRKA9KyBkvwVdZ3daB
5nTO1VwGRUKf5UTTldpqqihTPrFZz2I3kic9/QYHtubdBqsZddy16BNiXINO
L+UHkgg0FI7wKXRM+9W1nEJYRge8EznejI4onxXWntYL0E7pMWXpLOAxUO32
P1yXD6/mqrXbwqhR67hqj+riOrK/c9rNaZie5QxF+sBXkeaAOKXPtgh7nqpr
V0TBU63e18BjxGxDlOEnJVqDgfhW5RF1ZNaPTaHKJVY9566Yy3MvvXhTXDyM
s/D1d9/VhB9WJLC20KmoQsND4slQjR++HsInBVvt/0P9o9G5O/LwGRWaUBXg
8PHo+I2kKWVeULi2Ve4S+v97RrCMx4fQLYIpCH6yLcPzL+RGjTvNhF9tr3oa
mdqzyGIVyc5VLRZT34xeDZVvWHkt1dHQlnY9N2VzEoWGX/od65SujHj8fPC6
eieu3xLdNQ5/NZlEaZBdXnA/nVA5BaM+Ap6QTC9R6k+QaeN8x1mMI/Em+RPT
veDcxVQuWpGFwUOwtXlIh7pTshKmozJYGGe3dMFcEgh0cs8q7wgAdi/boBmY
wKpt4DLQeiQ9tnex5SOmaDbd4REl8L52U6+D5LbnYcYTh4t5oclGw2ZKOmX5
qqt5EDrB15YaURq7c7vRBhUbPhj5AY06aB5fqpD6d+GS+KkLP4OzbI++PC1J
hmbPo2sRl71nVARyaP1V5j3JfrDfIpyZ7mEn0io2fkC+MX/l02aTeqdHaFpa
u7JIblyHgvsj/9eJmegaJ1Du6c2KfYE2nDfAJ5UUpnKCrgl6wF4zhJQGbBr5
6ztr0TiZQFVqjoBLcCwf3tGCJ3CFhiG8Ka4ZTceE3RAQ+BmAJKsQ9+lN+I+8
JfHhSzWbsB3VPRfgobP+1twA6krhk3Pal7nN8fsqmvaUNTi3FWmIZ3BJKWi+
mIxymoKnpl05h6HOJ+vR9I+SLi/xGXXSTS3hjgYOTH3XHXbK9yFi2GMylB0W
ZxBP7QgG3wkcBk0CSBqDFoFo6lbuzuL7b/fxM4T6gg77FdlA9BFuCNJW/3Z/
XUS0whZPhe3YiyDjl7aof//54Exixq9dY/sOJezGr3coRqx/82MX2dp5Tkgx
mDdsfYJTapIdAQn4KlsHy8wM10SQv9KhAK/ZMtKFS+yDB+asbZ6n1Yn1+gkN
jhYonySZV6z3bfKFSSDFM/PhTh9rzsI5GBjhHZbF66wYde0Eqf+cvD+SEIdH
xqGXqCJXGCgKgjUKDA5NcEwoIdi3I8Pn/qQ8rkU5H2CQ0r9TLap+n5FIfmG4
9+SDFMowc60+0qdIzoYlxkEbt/7gQmyd2fUyydmFOq93Wcn6RdDppYZy2wda
UEvPZsrnGDj7qhSgDR2gP4cROwkQ0kJbvMs9fOl/fpyzUDVT4JtKpqVAqN47
407wpyo+i6CdH+OrQlYZLml8rcZXe2ZjVDd7Y1TWgL67kwkuKNU9q2vYl8Wx
URt8dvAg3VDfA/SUKUX3hbIg+MoyxL/2wSYVuSW5k8KUozR2anenNIsMlYxy
X3sFvSB0uqOzjCcBEA2JVWXxKMbDOTH06I+/SRVoo3wVG1GB5RpWstk0Td4A
LSbVlNvJJ2Xls0YVkraH8N/BR+/Se+iTtnwdcXi6r2HsEZQxSQrec0AMonb7
MiKSyNkQhA8VxIA+mM2Lr1Un81vLQVYCvTRKvO0PD2q8EgNwKCar+vEf9lq9
M7sDtalDrEgQ1Vh+1HT9ycp6QS2bc8q6UI1iHrrfimcMdt56EQC9OY3ROfM4
dXriY3wdaWCKUzPblPGAicW1dcmxhOTiz/k2k9NRvI2pI5rjXYs+0pZTbyYp
4O0QlYjdyuBJ2ZYf+sLJMHDwWyzsyk1q6uzr5jxGinePBLYp11XoeeOzcoiZ
TAthFAhgiLFSZsnVSN4aIjQ/hCJp9Asn7zWkYzpDni9JmS/eIwXzCzqGPbh1
/784GHRtKLJfqzc2EdYb0QXSTRKZ16Lfnf8qUbI6bPPgPFBiN067KGE5WKkB
Q07UrHBLWTNL2fF4cyyO6OM98Yw4tCobx5O+wKNRlNqDHdlGCniCiVBm3tJF
Jbei7aRYehSvNEftlevq/2NO6TeRf3dRfoXP3JNiK9bWprsn4I4FEC+gJ6Bg
WLDQlx+ApSxXm+Xf4Y6MvxLLaB0dKxToO3PUtGMvTz4Iz0g9wPu+vWjBoAfe
jJdOSb9ZnH7JJABlDKRe8I7V2Yb0HXze6w+aP9h3ODoEFgaYo5xlrzVKoW1+
s+ySW+Zza2TeORadV4O8ATmu2e6kFOq6fGOFvQ9YUasDJY6E2Lh2OpfJ3Wwo
0otNPmPhTpQbSoQreX+ZIxL7wq8OWtcWmdPnfl00n8djgRyLh4I0N305otvb
S4v9s2kWnqankVFP7wvYT7js7K2z6DkNhg2l0HfHgi/9x10fWatYxi3qj12T
Yh3Pgy1PXedfHJjs9drPYSNMr8fYCEm3niiJsheyl5/Ixet9R1OMcYneYidE
y+JSjY6zTx/AiqxcWZNEa7Q4VFR1qF+FM/8Fy71g6HiuBMfnRPYmEdD1KLQI
FbVH6TdQ2hcYRakSB7pAU4IKJqaW9t4Z4j5tKhMZfVcwABdnvMWB5sb+6eou
Ec0UQ+zu0vBGSwjaefedUReUHKnKAXBpZyS2cm1LakPFo+YmPDslEARei1Pv
4dMF/B7sDeDjFhwtf7MTjjEMKfolhCooq0RhH8F7GY6FepUn1uKD/TBTFyWY
Q6+WF0I7spJnJ12MQEJWsZ33Kt9ezgIPVdZIznv0phdCKK4cixjZLs54RNjF
5O6svrcW9w50pOzysnScgHDMzwkLgqj3Uw3dp4U8mZCsUuXnrV68qO5xkjuZ
nHrS+6/Fee/q1pmOvebMk1gTfw3KLdH24afGAQxioosoYeetf2ZjdelV5fed
YTIQKQTnkCO3i0cX02UXAibdTWFBPFD7gUG2YHJstcEVgAmX8PD1Hyhd5KgI
W3x+9XfLtb5scCpfMCx6yYNDGAI+1i0XYO2/O7Oe/4mi1KAXrsbZARnYSo9G
a8TqH52wRhAUlqn3OO/1Hzjio9+qMbuSi8LCO8U0ffizB0poG3aEdLoPuKj5
dGLLYXnx+0UGpo8D58x57KJTyWpXxcCJedgBUbN+X2LqODDGD9m3EMaxV6Xo
FxkLH2h7c/8f4qKhoR7txsisc2yeUF6PHpEnUsi0LNrbndodJ3FyxP7Clc4Z
/14FzDXj9a962UnBoC8/4aA56lejMCa1coPuD18STyxjXkr7NXDUlnOq5cfs
g9G6fp2IG2ixvgaWNdU4BguzinY3bf9mVYS+pcTJLmCHRYFUYR2VpZ2CMQbI
yS8SW2FjEpixpGmBx4Gi6thhHnoU+ObncGPhO4j6PY14acHKj3r86CRNUNrl
QmVdNOzavcdHGmlDXjpbYFQk06babZmhsNzgXkxt65XB0QT65tFkkpwYZSoe
uDgErALpz35yWFxORJhXOrC328u6GIcSuih0+bkpp7ndRLPprYMW9G8srHa0
lMQZW1GdSNxfSjFmX6enjRhkoRVLRgLbO6j9DwQSExJjjimM471+y0KcPFZv
m8leMxGSTNp+EpRxB23lAk5+FyWTTxHobOyHkSXhHq6ZcCZXvKXXPrtLO9+n
3nabigwDgjeHkTNfEYZ2kjgBtw9TidCA02WmtYkeE11qPSn8lNmmu8isE6Oq
75r7VCdk6zHuDLmmlOGtRjB44+Fxnn0jo/4kpbJWnjUTj+IFseiIXDWwlJPz
IAnjBM4sBJUCWBGXmEm1mtN/RFOGov/0hvu4sQQTs5RG1rK5NRKrFKl+eAim
SgFOgJuErrMb2p+tBnWpdexKwivaAIQ2D2xqerr5HcvvqIEdq94ZNTiSYd+d
++WLTKvaYqqf/qAEyfP/TMM7Fu39+yV5g0LEqZl0yEzC4PpzHMDOUudxFB71
XxK8ou3NU5RYN9DhsUWjL1Yrlk/6rtBVw8cSmcbUzemcFGgOaD8/gdl6+pwc
OweYxE9HeFHUVCQJGy4/7IBs/keC84srsqDg4FGhr2sO4q6JLEcBaenuCG61
u3C/GADpG1YROpuXTEcL6cs0mvUwX7t6IcXjHIkWaCacSvYeD3EJ7gv8zH5E
EEq/JAP6EVaeODHiIYhzJBLHGw7ULxDLgBTTHMmbVLw6l7Vgu1vVvbklYXDO
xlrWz1VlEE5pPjsedDFd0Jf8ny8RfradnHcUbaJVpKdBRAsey3AaBidWypp9
yEeUfdhMc3YxBLXr8b+cE1leqk/z2ptp6iwN/e9F94SOsDNruqDkA4QZ6iLi
YiBsnmxbXjq3XkGIuXwXujXpl9TERjLSBk+doRd5SgSo8Gyu+r7z6BsKv4+b
I6DUVdx/bzWcc6fFigF+d5vEWdYQTQ1oku9Y6cz7fJvGcpW8DHGFSAPHYMMQ
FoUY6nvIYl2cxZWDiURj+4VMo/W7TDyMJbfzWtQIgQqMmbK+4vPo1tO5DUzT
gXHhvMcTP5MEptDArbS+sZd3uctBqU24ag9a/DdsBHafq/qspf5bNeHwtUKh
OLk6Do0387HGQf6tyC7UbM16WnH6JgHfjOFYm2wVaT8S1agSGivTgGXal0Yj
aC9OTzSckEj+/5/Y57SCmTBiYSV/SCY8mstEmCEnC1wuPzDpRFuEFp56o837
bZF0vGD4Oinf9vEPJMD5nnUFiItQMu6ryQAElEzdjVsM6Sly0KkaV0RUYSzR
n/VdejPJRxAoLwXy/e/NCpEf50oRJa5YwriegmJPKRUY0jNgCqKCzCl+XhFY
itqJbggt4Z8j9u4Z/3kgNZEMsWaQG4RtlpWcwdUWfsev6wvdV6DxiZ0/kYBs
kTiKzexY6wU4UrDTZRmGNfUW3s0w1dkUT988OOnRgxr/ADBL87NmVZpb5udR
SDOUhz0AZWtGrguyfnHZ9CgrXyJjulrUAnEH6EvjCvlDmbbLmpfAD+1CeauV
eeEzRMHrrTn70g3GAf2Y31Lio5CwhhRewYOebYNi2HGkveEMvvwOXSCwlpIM
SwNhdSzrKD7Hq3ztzTIr6UeoB8EB3BKZTIluqDcsQ3mN1r/D7JDO7MkkV/NG
YO4HrqfIIVB7HzceHxrWT34BGacqMM7/3urUgqVhQs7+sGjNrEEr6hYELfiU
Q3szGtRR1jC+aG4I6S663yN2+mbkyH0PDVKmKXFTCV+ZE8JiR3+Y9Ycl/TvU
pYs7jXSBhT5w7G1tp+DTS87hX6qIpJGhfMD/+mj2qiduinSRB+0x5RvP1Kc9
hhFZNSLDOehdlCYTjGLz2jMRo5x1vSv2g1cLHmysXC0MusIggt4triOcUNsA
TD22wAszUhvS3NKFRhYGP01SGRGgrU6QZCNpLo9J5ZiYF6+COqe8eeeIEDxG
dxk2zQ5tgB+cQFUuRzqRZ8I+fx2t/XGhP1c/fIDVpdibG2J6Q25jTTNC+td0
x8ylVgs4H8K0k5CFZSBOpWSATHs1hB5fnWeZYAeDbCA4gfWfv9ELTVZEoPCI
05d+wb2wqnWdDDwDMbYMQc7Tv1QTOuf3cpY14s/9nHtVnUKoJCPrcYKvGWtW
lTUHCEiPD6HEDqNc46jCWsRODDcgo1q7cbbuT6PHtN4yMnGE1kaZJTGweSiv
ePDBgZXbCVpackCDkazq1CTXfylUZy3rgm+CFJAtc+eK48Zb82aUOcLyLpwA
7EJLUiaCWBP89xSDdQRqPVw5Dxe+SO7J0uzGoU4sEVcE+zen9hCx82p7h+Uk
guGHBs4RznRczDQqIPsLMKGg2ACc8LNSdx9IJ9vXq1abkt1OBcA5iwuyYyWe
4gz9NBrSyVmZUtykrFs6VjFeaeIIRNAfwrAiYmx9D+ZjVoXy24X3g8jMXohU
H0HTQPM545hDj1wvvYpkzB9Mqh4DXeHsUohTdxOsifOPE/sjSkE4HvOPeCAf
0PIUd5HEdJZvR6vtk9wIoIHCGIfnEtr+A/i7IXqHHSkODsG5CfzbX2nGZR4+
+Mwxd62oNMo+hkMm8tWc8q44K/v/gpoTihpN4WFZeznF6k4jonE+mLeMm97e
aoL/bbtsBKYKY5lwJ1z6PeWHbosUCD4LomGVSIXT7lN6jMmPztRjexRCraf/
i9CeMohWfTRKE18gcgszkxBW8fKP/wTdkm1wvkq4IPnHbXbzVD4RD5K5RmBF
u0DgsM6bQe30KOR4dl6D5/1lLiwdJEhb9wpcLT4hFozlHMdrboG5nc8LU+rj
txZTAJ0NVk7LNOBR96eWPgyi9KzGpqrCtXCqhQAsYfYkmLV6Cxt3+qFJw9XC
3OL9NDdMhq2GW1G51Rt0g+L1if+Xi+m7PvqDeflNvdn1dUJQtktoYq2tlbRV
0sxLMPub25cUgwD0NMfYDO/1Cbkj+4MLSn4POWWFBddYFw/yy6l6koL9VDYT
G8H7QWqvGnc6UDdi9i6sD1uOegSQrQQ+RgWpmdopCVaFtwzXlpW4l/8b2xJg
T3dGUjM6/XBV6O3UwFV59dE3v7wyDr4umb8BvAQ5I36ucrc4olJ8C5aLtcLW
yFNgOua7W+M+wNiDljg5zDX9Py2zKf7hwV4DQhZD18usYkQyMUwHNqHZHkbp
MoAPS9F3AOxUelzeOhc5X91yd7XquyPgQapriWpvEtnNFI1VSRNknsgbUK9a
Fu4w/HN+BJz/lbREvQm0bjedWE3N6kzdkRGpxHMeVEwAFfAdtWVLPzJ9z0BX
01rRvcdGh3+Pjy9raByYe9O7sKEWv5884liU6gjhT+NYHCSdsAzkO8fi/uRT
1862c2dpPDdLZIb36dJmvnknEWxOP6QM2mBXFHnfqXNvOZwI6WBbALP1bzKm
U3z/5ltnwTt+rdEakF2FUktlnRfoY60yonwYDnVw8NSbdxiI+4ZNaFdZIRZU
R6xH0oOdKAu1o4o9hLga3WCi5Dfr79RyreFHyVVt/CitFbhtLtNU4/cavY8f
8RxJ4mLzGCaC6wMWjwKtXl8dx/H8yv7H63kNfC4OLgoRXSyrljfNlQNFJheS
YCXWvtxUu8dr6zgChI9T0eArQcvAprEWO6QcLD8SdLebSmgt1naOT1GPMguC
NdfVMxIpRMadT/BhkLquwgYqaar1cMLFhHn/fxtY1TutRDwAtHNqURYZ55ek
uLEaonOZreCAt5JGneZxDA0YMzJtAHgoiwbl9MHaQ02xWwjIoc5C0YM9Cgzd
37LXtvg0AMifl+pxT4CpGIFJzN+op76Pl6mfUXlu1Hcx+23VQIjrRV5ufNHf
K7BS8qa+qPsTxKoUSwuHU2DXI8tyytmgqdSf271jFimu35YxPvdypYelvlDd
MRZN9J4nisb4ZUJUqatGHu5wPZotFYpcdGiVbNn3HLkVJVvmlQKE/i6ZG/Ok
+km0W+Sk4T1wpC1k4nTv31KF92WErjAoRgag0+A5ukPgdCzPPUauMUPMFEcV
7xRga70BEvofYXJVkcXeXC31zOzpkJmYHq83ZsvLHGK2LKaiuwcbjiL4ojx2
5lem7pRwefvVozltCRNXXI3fHqezSZPPy1Up4N+d9V/3mUGH8U52bbMg8ywf
zQ36w4yKtn3f5kMjqDVPRlInAwMIMCXGf2jXfNEKGhDjfm6sfY8wyzYpTDIh
9upGNN8c8uhesoNz+oakouRVH9Q/P+G+kxtIm3v8aTclVc+pyhLXkfrQOJsO
7KVgy3vx+wkN+OiRneUKaO5GOFFJPjKh6SSZzKMjM1066TI9TmM5APwf9ke5
jXFuUufqbRgYU02fj+Ak0+8vSF3tovUlq5waZvtNWwrV5Z7aHawd/qOGkyjh
dxnIMoK0soJ7eMfxaE0XavDqoMqnvYYbqC2+wqsJqoiceuHIdv1pJ82V4ViG
3ks0Ei3VxRzkEUc4B9SJkYAxsEZmLyNiaPKpLWCmxdqCK22A0UYRZ6mbUxDM
fCvhjmexAmAprXdJ+9YRZ6MGKtQtVqQ/QeJlNfv/QrGZQEIGBjWyVh6h7IOT
ngsFRbe1217Opf7jyjde89pfIVcFlrTngKBmDwKmzc17WQKRhf+28qi0XlRT
VZL7Idfv4+gxRomKU01vsFcuAyb8JYGRr7q2ueRg84Zxr0vFgtZZWCizNhiM
d7B/gOtZsS18KFjKa/DapT8FOsHHsN+PBlkJR2Qr3psH5p+s5Brpb3rEFdCv
lS4b/2XLIDa0gmiuWehyVxeOhSmJbvWGgdO0L5Qf+Hgj3O+CJBU6BeV+WIcm
MLDNN6JHzfXNgHVvidv9kufbSzHrHCIZCSHAL0bdWKC4sj2Vh9j+jTD7Zs1j
KLAa1E8iYRXXrh+QXELs4QNKxM0VorCN7dOGl5VVBHBsnNo5lfXdNh9PGv+L
gQvuCKzs2vc83mwrnqJrLHnySH3Nj8BKM/y20xzep7Zno3nuinYs0oGofgYO
dCnt8s5aJW2RS75IekG+1FFYaXcTzDkFrZZZmo+wDD9FinNpvHQpEwpp4dU2
s8L9Aq6MeQ5h10GZ9Ir2tF7XaUs9i4VsiwFL/kx5MdURZrS0OJNhbMc3zzpd
lZvGeiSj8ktr7qrxFgOXMeYtqpdgWfTu1tk+AeidEe6h9//4JKKldgzoLa/6
R+kI+hkfv8hicNHf/ZKsHWd5qNw77OqRlAToIVXCOCCfkRiueR34O8SRrmK/
eNQ+0RV4ejISRVuJ4/oDGEDheNpJpx+Qtj031SYWaQDXGPea6HvPGHlTG5cr
ZvcpvBus0uj40e7+c66hAa8SEaXGmRzdrIzDYbg/9/t6tEtA87ad2nOZWG9t
PJ4XQ3VHdG98Y29tYpRNVT0ffCYCUxGWk6ekn5m8KtR0jD+/xbIDGTO0tUPM
MQxSvT3yRLIrenzTJVhrhmZteA6aUSjnYrTv5Rio3SAuoZ2vFokivmpWh4kW
+jWQ90M2zDUunnQE3TI9U0BbstzC7p+I7Wr+KU7R2uFkw6hAgHut2nF6lAat
cAoWflFWzdDXIYP2tRlwu7t9RVNzMt/zOW34w8hytSh5WTRMVDKYDw9XXcPo
JvQ9ju+KJskDQH8axVVFch7VMGcZ11qvhcciwo+mrUh7eoh1PhhD/2gaaPcZ
hHHXWRWw6T5CjjtutjHtxR0qKKGUAIX4YEZ8XsTkeXrQ5O50YK9W1VI//8KU
zJmGGtJRNi08bWLm2P7S7+nWb3wV+CR+3BI0NJUaGO3rxFDpnr6/I6xPSGfO
WSH/m8O7vfYK+fBb1bXJzC9iR5PwiWNQ91vkbEHLM5yj2/xB0fdGUFj984va
rF6FmqtmQ91ZtP1q2eDviuYxCnsXmjoRM4iXQuRdiavQcAMuB0GY8Lpv9uiT
M6GgLXWE1zwrMT5IFGYcf9ALOf16dhk0JsLdcAiI9XVSeaUeMZiMb5d8wiyF
shwVgRvxc5VZOPn5ezqE0n469pm2icYgRQZqyTRn19PQ+6bkzFSx5mHRsI7X
9V4wd5gd6lmn9uICSxPxdN1eu5t4BnMd4o1ZnpvGxgaEM7kQp/bKhvlR1N0i
UvlZSlY5vTirSwkohJShpuifYcjP/wDJK8iSRoRhs3sYGmwySJrFowU11Ts5
yg7EATlJ55EFxpvxE05pO3fnDqtY5yzTCqr8STUZ6skKaO+v0sADOjyQWlOH
oRIOedc3cqBdHCi3TuWgVs86g+xQg+jsbg8yBD/5s4rvdmNAWWGNSh4+1//R
LUZU4nBh8K+JTpv86xN8LfUcM/oOGzbFG7Ck8GA2nXO2EeyzqjC5+53XY8h/
uf4u5DAy9DyLIxLvksJL0OkdvBGM7JyDfOnJ5r9rhx3MHESAcLRvaK0Cl5dE
/GvLDvm+cfbBnsfYluvWXbv0mt0+bjrv7odMQf5OfC/jnb3QIkhDEIH18Qx7
sxFL4YqJiYhQb1zcFzQJaqdDS2+pP7DyU/0EM/ddF2k+PcDZihS1mhFrgYlj
vof3sFZWJNyusROmXnAFZdivPxrz2DgpGZpv+UTdMlons3hY+bsuQC13KiSo
kVMGHYvY/afE/oqoKf96jASthFpYlx/UqR5ggmAv5+Xp/qjJrM6xkHfIHstd
n2EB4foIgKVsHi2a/7AOdpd8YhdJxX6GsbxO0nRuvMTM7sR19wR5F9HC6LlO
WkLRfB6Ohhev1hGP8nr15FbjXpTQQniWtxvP6Fe1qgvoGwvrL07gv///OR4y
3h6r6TwkF35lDYBXFlFnE5H8RGavsl1CJj5RVt/cqWtPcptBFWM1x3wf2cP/
8r2Snw5F284RfZIaRAWh7Ge/Lro0CXfEYXa2DdnQ64N6G17ILXiKNnf71g2i
faqUGBUBT2jmMT/CTXou8WTf87xf6BJ7vhJtgg7BC/XV4p3oDqrpX+kH2a5f
UYOIzpTaHUmHfRu6XLmR/ykdtklqb6Lqu9AN5WBa5zbFiT1nk0ljzeNGW0nK
x7E4CgMfKxOJKkjylOf99pk6YaZpQS3mCVeaUI2ga+0+6zX8++wBCtJEgV3o
9IaXipd5H7oFywSgxf8bxur799DDUN5GXU0SnoaMJiY+ZKvzJA07b1kge06I
CM/3dI3ZOr9qmZo89k0P4NZco0GH3P8ozS8cBZ1vEkHq4lr6pLThWKeDtKpD
6T8O0CYTtbKYAbV5qBW2u3pwm3tPD4Lxu3fCBTWL8W/Z1/hGszvRZY5/alWp
N4dd9C/bbG+UVc6zMM1cPmWoOspa+XbYnouCLCRAG0jmJgm+3lCJdgRNiakN
KWrzRe4zfjp9WQLQFpvDcj0RBtIdjfRXTAXbSmJhEOInfOxeChqGDRbp7xHW
SR3i4nPzFoqNrBg+4qLFYcb2BFB226+ZfYResdOqPJ8i5XFbcCJXz+QQReGc
27Hii0OhpWJ/L9T61ADzeJp77PgptzCnWhoJdO4ghFriteb9EX/iAsjfFnsD
6iET/6o94e4pDiQLjqJxVXoLFpwW2656jbyRaiM0o0Jn65s3DLIIT6jxMiDR
fGXi1CVbnI9iz5Dq8AHPfCHd3QEBCIw+UgiQSYl2HsGwHNhFhnWW4FGAAD02
jwL3tvduCgBL7d+3NKqToGiP9lx9nWh1sfviLHyuabr08ccv4+JCJ+yFtbc2
lmE+0NX83yyhdgIaDvXXgN/r5VvhnYdXCLcSloqL1Ke3ciFKMt4whqXt8ao0
pmQsaFBjt6yseXSuMrLWUopE5elwOEp1PP7ij3J97CVif6QLnVNyVA5+Tf7+
ZDM7xChllLmx4Hyah49KjYhATl6hdb+Usou3v0wvEcV5ySu7e6O9QE7wK3YN
Nv0iyqtirarxrsa1/Rr7eOxx/KUc27cKSNpuuuXDcYrAsDZV4qUPKZNRH+O0
V65CVK/ClxSefkHTk7kEPFwAQtRWUDOlDfUw5zOsv1BJxXb00nYeM8yzeS1l
W/G9jtU+czcXOC6ts+Si1/Qjfs+H5GNiDSnhQ4YVxiipRV3lSSDOzzOPvajL
zzxXtW7QOf66OiCfwoK38Cp8TgtSCO6xJyyjCX5ikcBbz/FkOuIoantSOCRm
j+106m0TpyA4RcSvr++U4kukAeUwc9QsBPlxxfrKnP832+l4+0y6KkuOvP1I
5fpzC3xEK5+eUw4qlU3XKnGaxkEh89pzWQ3PTevHz01IWvJ0zRUwxTG3U68T
7xIrAoWvxyO5Tjo/0ZOQNISytZcIeb5gvtIsjUIH+5OwSC3kCkCa6Vrl6O1W
tLep0SOEVKgOmmfUT6rgdMT4UHGyT2FaTwy0wegaTzIie7n7jzEPy+GSF1ES
QveGLElgGM1NPzP+4Y5cQ9EDk8Hdh+gfLnkF80jxkDYWYC+ndpoXcXAHr7/R
x2taNvPcEXgExGQCl+4NKuSvBdO8cKwbLqtF7RZjg7Ql7AfmoiX39/N2Y9IJ
7pKBm6KZdcr7wYF7iYObi9XdtSTylrDItdRK0DvUm2cscnG1BrXD2ASLgiK6
a7AjprfaEzmWwTleS7mn2pWLOr6GR3aY/3cWCG3yzK1wJuWoCcmrCaV/Alh3
CH5ieNDznKY7PSVa8zkjxJJAeMI+mATTByr2Z0+cvVFc2uccNhiCR+QClGz0
0jSEu2L32PXuybBJUisdNnfhicWzEo7s//FP7vczN9tTVCF/+blYLKq1eBdz
5npqs5Y44U6rbRtGVZgzJVgNTHgFvRNVArpgcOgDvjhMSC4o6hSaqJt6rbxK
nlWQb5EzALz8NCRdNwR1UzDqUNVz82Luy9q2BwUJsj74zbFSriMQgRcrBx58
rvQXdRUCiTgusRQdFb/shVEtP7M9gM+9WA1lp2nWqNJROp3tzhtYEBIpW8ed
1bYBZuQPCY33bDVcLPUMTHRo/36ACX0LaElmwuR26gmmYAqbO9raDYiIADkf
nC5eAj1pIXaTHwrl3BssxekU31Lu7h4lrcBrc7CAHeBZVFv0ijYEpj4rzA1K
kfwBn+tS6DtFynfEb/cYRFbpSjJC3dPM58J/Veg9+AKESwaUWZLzeTMVdoVz
q3uoxl273tJRFoRHTJjFJvP5LSGGwBf/AAjX+GS86HyomDlJpnzYNmNL2eZe
U/lG5XRk6PwG8GiGnQa/N9axytPotnwtIUhIzmHUAiVb2JR1YlEwes3Arv3o
adqRpj5bfNxUDZ7rr16DFMayd8cr/fztP+LRCPZ9qnEC8rMq1F7YWdrMZ+9X
W1ijUr9lpOPJlYE8nhW6mVKqD7rCeeRt3gd9/whCqCj3s2wvtBEQQkg9sk6z
IGJpl28HgT4So4UQwCUnSo0c/CIi9lw2TR3Wvopv3cAjUlWG+gf8SoByVis9
H1klM5sT6/0bjoPbWuvI+w4CrEYrDPpjt4/oxv8JWJtjvgIxlo2zgCec3ov9
oNMw/8+ZsZ7rF7/MjOR8Bfc+sF6Q1yphHpBR1to+qFGnVt6qcWMKy8nuI0u7
IbOKVTiGoxwNELr4nbYshq8u2EJKOm9DzGCdZ48v5uy6yhFJAc1VyOiZPGPI
wrQqMuK4BVN1cx5F6pJX97nJ3UU99/rmd4PNXr4XjmnPHIiaB56rkJaB5Efr
okkm3AC/yXEGf4RthCs+mOX7cP26NgjKaijGPsSVv/kMLOA+aH26F9yePF7U
WvY/l5sN/66rsaUNV/Jwfql8UxOTe2SH34p1i95B/cITuAMDjCIq9bnG3mol
XBLcnth9stkEWtZgptqHXAlRjRLEsQW3O9cyC5HuzE761jwbxpNasgjjAe2G
2bB5C7/6Jkx4flzC3xAHLUGPGFOtw3Umn9jc2yvYcLQiDar2zsxogGIctyhz
2gYTsDwmZBa+myJm99obVNUm71HzUfCBkrWsHkiewarj/sZI1UPYdIftOtmf
wOG7jijdxgv4JBusFKRamVNkogURQSbTXs4mpBr5WyQ6LSGBCDevOaYk6x4M
CnJTNxNdGHNYjXTsmh5QKZ9pb1RaDi6nxK9iWewIjx5vWS5uuIrMRdyMoBkz
Ni6fqlbU6wFLauF1Q3Bzi0EQledw88GZQaXGh8oO73iWtq64/nwcjKfFER5I
OxnAjRve0qcAa/UvOX7LYqEUP7ph/bN2JUu63nkNbBCbuzY1Ch0Apbe2fnyY
gCE3zBD+T2yzo8f9EJQlR4d8xIi8liSTCcwC3QsKfcaP7z9yqut5GxXLy6Ao
+1k2giMGDUyAEa4CIo78ZjDqRbxdpIiSpariD05+01XOyo5Vhj51UpGiYbVi
OrPwzFYuXjVRky4eXfRT8/opFCcts/b/tEA416Nwc5xrrLvWkY9OZdVsIITa
3EPn/5HaSW50syIEY/YGMWkokpmgSBQne1QLuqDjfaDkAT0/Zjg1CgPkHYu7
9uaE9esu9txjmSD/PRQ2ATwOjq52uB5HpCssGZ7tlso5FaMCI9dYjszijQJh
eUsQ6HYchaXqwcgZSE96bMF0Ggc9v0udwsZHbSxeqkgekRYcUlixdhytCaJT
8eJsf04cnP/t/emIHRztYt3E7xdNY1cjkhRRt5CPi2vS/6Se8OlQzgjqFXwA
mjyx8v2ggheLqleYJQdIrIAWCb3MtZkGlpn/gX9tgAiMjON9jt/rpmVe/k9R
A6Ytb0DwQKYTufPW33ddyhVzEgGDu4P93vRFGDBFshVI+L1wVbBo6681Kp4/
wDkXV00s3xCQKPUJrF0YffwLwvZTp594abHewKFCMBtcmECYxIJ846v0tvz5
WQ7GTnZC362lViZO2HbQelOATp1PxT1WNgaou6a/GJLPJWDfTQ5wYBOGA1hT
qkpRu/PDF1xvfXUw4V89uOeYfa90GtGBqwf2vpMjNPMpqTgKuqOwuyWhPPHU
+8nf/qv/d1n8wch3vzVshON2Ao20ycy2oc9pqcnlAXkDiJZyMX1NZfUNlSgt
EkY0YT8wViyNHDa0yWygujAtx95Ev10qTU4+PvLR4dUqmE5mtCC5OVBagjrr
Z4bWCm019WsRs2RJDaDDrSWvplHzXzvWaKDSWS1KUSRGxPGddiZ/AZGIbyY5
7plV1zLwkiWpKG6Usjf8PNykBsv4JRWkj7++dQpC6iQ8rxx7ydhNV5i3IwzX
jcz1M0APBy9liNoK97lpzWU9ly0ZK/nXQdmbi7SnWlJ6wQ7v9xzKLcj8JZGn
uO9xUmIoxFX2Ea+XdSjcUMopAg9hB9ZGbbzeX8eCTHVgNI8ziO3tKHFrM2Ua
EmX0dv38sELBIV0EMFt4wkPmBNz4bOryrH7cz+1C2OojCryN0AuZMPsw/r3J
+1dKGaRH2PtCe04V3rv+GwpXNgPnhB6lqT0SYI8ADHo5Zk1ldy7xshXEXEhg
Ua5Jb5n7MHQlp0UedcmsOu07NXu+oHfRmavLDQnntA/BVbGTOyG5FDxiWg8z
9uFmx3a54aI+VoA3UQVbZpt1Iab0tmoqddzMIi+4t+VG1xUfJqaBUZ93eCrp
nLzelEvN0l7eiqqL/Lr8K845uLXxE4Hcoa1IzC66BrTL68W6aGOqpHzldwlE
Sqp7RGyj91KaSC6QWNx0KkmkELfNkEIwFPfSsHkYIr0uT3eqTE6JVbzeKfEy
hSYbk0bVn00z90vl2WSTPvrFr1++JzaF59D3OVgeL5uKEDcNSFw463KL2BUD
bq1A3qw6veg7hl6vwDOhqRMWSzEuf2GfUAqg2anUkXeTx9u3incJ77ceERBJ
/zoNkbDtsL3nrPqi3jw3tOPenxaBI09hAT1DbgcMH+gR8noJ7Ksfpgk8e27t
HBYuvaBn77GsATRTPOoXNcKxqqDoTUPO0IipzINLgUudzF4Z5UZ5FTa1U0Kj
YctAkfxD0Fq0C4/0EmGX4IS31NtauZKd89qfV/cVcPVqova27nrfRdExhFqZ
+uYUZ+UvG4/S8oIxYBg/d15D3oNT+SBzTPTYnqorlGs3bgLVVUA2DKNkGdn8
MsXRwlu4tWBIF7PXJFAnaYkjy2IN+E9TcuJ9VNhBh3C8nT0DzCLbtEC/Edg2
M/+yB1PSfocJdEooSIy5fMfQt02x6GK1904oPVeA17S59jT6wtUHs/Dyuee2
ZcDvc4he4SobefeEoyjoD+lPvOd4HbqXiLgVZjoUcRq0sZigXqBUnTPt2vMl
Z7UXOgZICdx3zoxd210OG2TUOVcf80lZOCqCt9xMIojyAkSUe1QW3EfblZW9
SWOH2x4glIBrQInr4H4SCZPlr2NAM4MPAzoKkhs+9b+2z8/wwPnX6ZuCCTCG
XFPTZGTHOpXw8C3L3RbjhBMxbq0G/TTp5I+8mBUbJwXy9Iyj3re0YdL/Ndwd
LZcneFS35kTuVMqR7yax4Bh6PgCkJOah3LpOP0gdvcm6pIzw4zdNBMD2ZHGj
388kNUuJO9P6Z/NpmOV43vgjmbgvpCd0buQwSziqkfskjW/O8O6tJiw/uuox
yoCvxMs9lujewtnnxc5UpHfmagq+FLe6j6gVULRWneoG9OBxE+0is+n3kdH1
6+ygSlTidlOCvOSVil1z6NOP1zDfMiTCx4auP7FcewhqtwY2Vngp7dEKjqvc
EisKJ54jbNqei2olxkAIfJWmPIYJTNMLothA8OnIbqgSOHjeVHGlVQHzESOH
GfEKFBUH1+9SYKvxQ5x0CoY05MllVMyapbLps5HFCtxjxRmHQQ8KC5SjINYB
SeVBlWfLcgyXs9kQF0bkFDV/3AGGdjsJYav14VHHD/RzWKczsmnxl3i+7Okz
wC8/na7OPLI/9p7v2+T5WO+4+Lr20I7QTmhxkrKTxAHXFnh21qXhJ/ZrQ6Gu
SMJLrC2pJ3JJK6qdEbwZ3ddAGMdN+QdIAIiJnOsc2mqHwuEq0jtRqgoEr88q
IhRgsIjrMRFDYtD+lZgXJ8unstPx8oKoXJbNGQqMJivrVb1bOzSNNy0X07pS
vY3ZRq98lFDClu7BDsTG9z9BrW0FoHSlOehnU0fUbVGRAv4dTNyPIniUPYDI
c2I1GqdmcttZFhmar0O6kIOIPIOSffIOgeJk95MtmaPlDvcAwx9GGxuCb/pO
QH2Agox/cO9qeJWV++28zZ+lZq1e/s5bIqvKVOsYl4oOPA1hIiC5p3f5W3Ku
wAY1qBE7dXMy1H9LQ/gouJLCuPblRvDFAVAPYscy87DAZqpUHp37wO6pSmLf
1MBUjpdxdJyWt//EYlfia4SrBcQNrxw1+OO+yGd6GP0epUFE5V7fpNMDH2QW
GaPre2qERkuYMOxT6DR25/MRp075NmLuj2NUUKxNPJe3+E7IsPR+nf3HlGFP
9Fquv0eEDj1Dvq6y+iUUaqIHz40JzLEp5RdJ83JkgEDXU3vg+3Q0tDKFqFN6
eZz/A6FDSzdmnhWwo/p2fR9vyESzDoXV5Xxl5Z0/4zqz4+/X8QZdiUzorT1w
0ZcAORcHds2/2ODkAZQZZbm6OUEzxKpsag1nGzWS3dOBSEVq104XEDeyXolj
iZZmhIjnqS+gqL+44Bx63e1eXawgwVF1dHL3n9x3ytXsdBEHDX5EPPEFXUh1
QzqEHbamlBnaNJPtfq6iEqhaTmBe1IN67wQaOM2NovZL7lw3WTgkepTr0AWc
ppwPUoanvx+Ln3vfs7RwBYgYOS+JROumEnDgwlfzwNaMi5r5EKm4rb0KthBz
XwSaegy3JOMHE1ISdFZfibYBB20AnN43uWZJASoi1PEvFXlIuifg0tJF/+gr
utuTxl71MfJduverqqWfvCzLRin/dfFbWiXGgZ3v2p3BLzXSvWYnvcseNYtr
C01AZAGOBRXWhfk1j+A7N/gJHnt9Sj9HKIEiKtFjE8wgJ4VjPqWTL2mxMdXf
Olr4jzqKTOndOM5QvTtgofS0K7sAVt9YrnYbbIh2bIh1bxsWTkf1qVxv/EX6
gZtaI84DCULNCKlQSPtRgMKduR6bcKR2yDrD84V7RMd4aOKAXL+Aof9q5kVh
VqYjv8tGklRGYrar4Q4EVOEnMuKhz0HruQXsNf03+LtpZAq++vUwPJW9ZFgU
qwhKaXsomGW/j1wnEnCSllAfKa7WJ97uOY767dWC1oUbh+njCYAJUaBGbHpD
+u2wTyuGYIJDHuvoJuWCkFe+mnmpMIPoJOMl8L93VHDIsYg+nS3IKRRcUF7J
et7+bRxdz1N7UrKAfdCsAbXKM1FODd+5QHHeHkpQiKapEedJQkdZM6h+bHYJ
bPp0ZA3xrQqqEDCW5S2F+U4hjrElpeMj9F5yCxJHVKDhtijW2kSsJ/m0hN5x
qhW2x1IgkOVXAtnb0OCDnzEsogbiMmt+IiQogVysYNLbSxcEpOgPQvJKawdH
ZR4MPN0kMk/VEpjdyi911Xd6LHnfIws2c2NoOqHhcgfCzLUVQRumftDwe5Mq
EMqfUmYPh2xzFy84cHe8CI3Rk2Xkkcu+dlHgXJ6UXyVdQjKCvMA7AHS9V59n
sZ1Zi4IK4j3Y3Iu7OLh4o3M6xdKRD9vHRb56ZaPOHUk0f7pSwAp0DQ3IA1Jt
Vn/CtM9d3+KqbeLyPlYoT/vNVoY2Flruny58+PllyfauvbOZlNG8r+/hr/GX
GA5keeZCZj4WvZ7PKiCDB2l7Pe9jBGX0QRcDarTTSODDO0l0bthQ9EL+cmV7
tz3cpxvdaFwA1CGwatwHHKyAje3yUrX7Yha1meL9o6+VaSRz1cGWoViKRNUz
cLFkn6G+ZoHjlpOhV2nNI/3O5ayndaQ9fGER7YgndIm8bb9AR8A1GGp83Szy
PurkVrwgiWASktcZglDxsOev+gVPg2P2k7sea/jxlsmEq/Wy+xhngRyMrGrN
ioHCGFpkyzdfQficmC6KH9GhjEhoWdxTB26a0ORGboEbQlE8aqvjbVvQSo/s
Pm93CYgE4JoswZwm5ajIfe6KOrKrXsytHd896xqev9F2qpZ0R3nsEKpg51pT
PQEx22/qiMo84zZbWExhTZN/EXEDEnUlqvm6nEBB4jKlnBBBZTo0YjYvC7UB
YJG63A3DwaWQQpzvnzkBtYNZhpE4xtiQdqKFlfd3d2j6oFQ+ie+zsNu4FCiD
JnvC/aiOxZTaHn2ZoRug+SNrGtbBzQOtayZcFNIRwFnXMprBL/1i5i8MQrn4
o6tXFZYQbU0pnMqvCnciRhhSDj9s+G+sG4nDUnZSXxWgJXSRko5kz14tRaxH
HT+QMGSO9fW6FRC5mYH6JQlUm/rQlVs19y+S/U1hiaLMNIJFt4XNP5F4WThx
Jtkr/oI/4+rUjPnDIeQ/XE3hTdGzDsTw3YJgBumKdrONV951bxI/6AkEmQ9i
mjexuPBNKHYV+vDeLQpQ6VEWgSaeQwIi/dZwEIoqAAw7MPOK5dSvtHKr1FQW
LTGc1fTp7Z97DQ/UyZHXDLfW2T3C1SF5Ru/mSHmGEkO6vdMJAtWpOJfCtGlr
JAozeUJRGboB2ljAACtPhLzFW2h9UHmGFtYunBWaa9xJ/i3whdbrjV6pd3If
Z2e4PpQUalxTuLrmpidtP9OMsE4aOEEmwS5WU32kCXITdCME8RAAUQq9R5Db
CoYbe/8zeXzNERo8P3SrJn2i8l0v8Yli9Z7PQveZ422GIVKsi+GYR7vkPKYT
jraOp5W/2dk4aHU7OzU17JMOvnIxjDpMntu3lVWmxGXWg71v9AWhpCla5KUN
RuIrV+EwoVZJEIMABh3eIm3UHtYZzbguR1fnUR4+clsy3HHAZ3wbYeQ0ZDAy
TlMhVxfeiFBxiB35XM0yFZ3ty18thLYj5kwetViT6x9dUhfQwpygNMmfXEsn
qr6oBBw7EzFG/lX/3f1rvkbHDxy69U0pamAYcvhLi5MHd8PJ4XZEx6FBt3ta
VdWsUKgtN3B8IAr22PoEefLrPWgHpMuh4PT+my4Cj3KQHosFlpGb51JZhPiI
y9f4izdTLkjIil/AW4x5TP2HO1WF3IiNcVnYUkGr1Z8vJNTDl+XlGoVnu5Do
pcQHiWLn4U3GUO7viXLbTOp7gIY0NwRqAL/V5YascYvnge0uTxodOT7UWldN
QGpPFSUvqa+HuKgQdKgIRGeJTe570bg3154Fx36bfAUviQICXSA38C3vwCgP
UbHLzHcgUSFH7FIafpK4D0W4mFPCgb8SNb30jCO+drmT9f6p3ha4RcQMD4v+
679uE54Jy7WQtciT6VLMmOGaASvyDq/8CYOyA+c9SwpOjuPccscXYizQYhO/
NM6gWXhxKvYzOH3GmyCCuXKrz6OGovc2EfJKujGGhu6b/l4zgAXj2OgNzMyT
MjezlNEAcmJ4rMRSTkBJMxR3FvOHY0ARaitABxTjuOtgeWCG54ZwiRcgzu1q
p/KcSIW3XeyhNjS5bMuoKFd8kSSk3+rRa43lSZRZWT0RhFGe86Wlqjhfq3Ff
/CcadMVduaQdNYgFGdaq79vIGFowFd2cwKRk7BdcJLAg5s5KDKMIC+2CSgUE
/FvyVVGjc8WK2mVIpws5xLdQUP0TyWfoJaSoma5mcTguq94bN9Jl73Z6WH02
cJyvVx3bL/Zh6xmhZTbfgE3LzU+ir1cjgR+numpmMNv7q6aBdZcikhzpNe14
TS3ivch9n7nEUci+74AYjmnDT/N4D3O08RO8mJbHjfaOvEhonz2fb9cJpA6e
kjWnN2zj8RxZHRxCEXQ8BGGCUWdR7dRbwRW3zHF14PMoAyfTWcVDY2yHV4q9
zZ6C0JqPAcUtIDsbEzanouus1d1IpR89xU5WikRWvDjwIn1oVnSTSDbOAuQN
xBmRbbh6G8JZVfpnrLbbRBrJRseAnNnVSqOTJTafCbdR94kBRHa2qFhdB1D8
XLX9qy9A9jnROaHrIkEWE/FtydRaMC4f4PV8Pnpp4Ecg8U4LOlzRnQxWccbR
OjN7GtMLGOUhv6oH/pl/THNIXeJytebqAtcnZAbnH5t6bvSDftW/z764R+PS
PglNsii3X7K3UCqSwEYWGGqmKKpzY1PKB0F4QIL1++oICL/uG6Qfo9MhMXVB
FgxpKSr4gzmmu1S4o4Lq2Mfb0XYNm3ARbz8JmXkApZpD59WK6RPEonzj1EFF
jW6WWEjHJkzPfXKITfIlvM9m/cwa9synSMdyx+5HglZRKe5O6EdFUfYrkvUd
yZr1a7aRq+HaUV59cm8Wan3glvDYGpPDvWlzCwnbFatPFt554xLRIrsI3erK
fquHg6ffZl0wpAsFLyk9+JosQPpT6SIuBpVj1Ua+/cBB06e0R7GENKJ10uNP
4g5KQk9EZLiSA9IqciJS7NhYvkxK0XttOIzzMIYEL8jKiIDK3QpeoNLDSA7m
6DDkjRgaZNOJM6ZZmjG9epAOSKMViNiRZTKoxY+Y79iMMifMt5dG7s1fcdOd
N23bi7cMCU5K+aYW1Vh9Doq/Rre0g3JjUXPVy4QTnhuqQnk7z8OgQvM/g6xJ
8tYpRc4XuQxspU6yU7zVCQ3RM1TSlGMvAx1syGYUCJtCWKycjVdhYggHIg3e
BgRiy850HfI1k2dprxY4bhmUT2S3kIik1Dg5ni16dh94FGCk04iybax5P+3j
3p7zKIhRkUc0k9BRx+vGkiEXC1tykgo2DCkrMd3fVy+GLMRMQgTfncWruxa7
YM8fNLpOyBSFBJeB1q7jwFn+ogNMHi27HVd8P/tt/bXUq2p0zqap97r7y9j4
WK/u5JzqA5uxdo9sx4h82K8rMzXIXgFvMZsLo3oLd0C4boEpCuyOz3/7vs+d
EO13IL/E0giu47KBGimGmEx/+61Lo6D2fRvgppWzBId//ONxRdWN8NS2qfen
6Mv+7uw7KJRhZVLGjVlw7eM9lM6r1jm1hT9TVQuVnOcgqi0eguzj1urGX23M
Wn5Rk4Zrq4TBRPxKhYlQY5vANWdCI7hN5B0Cg9IQS4aq2QMdXtlj0OIehvaA
R1zFLjBPt86XmQGXv154OmWuy4bfodz8MvuCUgPhAxcZAGuLYemDPb5G8xXx
xhkvKtjqkuE/zsk8lYbiZOLO49sPAxrKV0vhTw16YV9XmZJjUNKIqGfM0QI4
piV8J5cPCam++MHXhEXTy3Y20DOoMpPyc0FS91CTlXL4FDVVA/Wu3YbYdfxG
WCOuDRZTOwCnG5KS6s4Mimq3QJtyd1x2I/Z4sAeKqSW/UsiiToFU8yCFwHQY
mIg0N/FWkDxVmYyjiR51dHPFR76zoqSptdRgYRF2z0MVPaNQfSUM3GG2RYCF
Zye/R074oj3THNM7F00ZYN1JUiXcahp5heFaKj9n1B0FF4I1hn3CBmyvHOKR
QVu8Qdp7lYJOPXyBqo1dEH1R81lYbstNs4qE2SBP+MpWVbHLkkzZ687fViwb
skVElqHxRsdrQO5kEBgUbRMhLn1o+OUzy0BACBHXHK8c7m5Wo911hMPe/zZP
dw2NRtpSB6wSp2rMaYlYcw6W4YJp+8S1CmOC6o35BMLXh48A3kMVHiOuWh8W
gzFlKwe2UApxkAMSN3aph6YEJxIGdbZIw1gc4tOB0eSsq4zx2nHrLI6fE7X/
RKh9EzOu8b8OHjsNvvOublNesjIHQM5WJF4kPuVfKETEbHrFvIiLQhVW/ukF
CpqQxQBGhMzcsUzEh1XPyJei9wOrn6uTMnCUDr/WTRiQT+nqUeThTpEF9N+F
DP910HEvhMcChBgYMF3YRbCBjg9aV/RVEa6o36e0mFBFbMj7WbzMq17APqA8
ofF536noxE3Sdrk24k2DqR52/RP3ZuZlqFYOGAGLBIi4lDfENo1lvw1R/h2c
MeRnMqDs5uEQcudwicO1LNd9J2AFHRL3mPMv4JmBcatf39UbCdMy/H9JK7a2
ur09eJ3+3FKDkVfhGLnDYxaJFWzRhz7z0Kq6Mo0OGplqwsa6sk4OeFEzPy5F
Pj7mlUpzs9KU59M3k07yg3F2w+u1hte1XJXJQ6PnZlNcetJ+m4AniHKyAlfH
K5s7UxdvOmpZLnEnlDfwQ6dj6HKZXVACF1k9ptnvbYO1+3hjJcuGhYujr8YM
w0EeRivfdaxS9FfU7YmH6yCbZ9R6A1ydMR59jxpUbflMejof1EVD5SF51wmd
5ZUEWuiso7ffZfVPBLbnqxTLycop3945Pcn4cxK3HTjF5whih1qGTqWmnATO
dIixDRZ41g8b8EqGhGqBSclUFrQjOafjUehopPpCjVz0ZeqeIZSCf8ljDxll
EkoDOk5vq4cEYZX/MCJQ/xGVfdXB5+32tgpXd9d1kydBAAR5/76+GvToaK8e
YJ3GX5/cS6JcfaNkVtRGtgrjEB5s6ETu/B/7cFwAeMYRpob0/uqv91kDzsTb
USseS8WIknnO7ZDsOvIWHR2koorrbLzfvp4LacnzoTp70lBG6vMLUCkTZBFd
F23+2FeWbeJezkp/qdEJXIZcaoWFo/+Rjvf2dkH/tKeOAsl5p+FhC7ySINFN
soQNHXfAETAtxv8WxTvwSIC9xl8HLbkJ4+/RVyXpI6dYwcyRZp1z7oNso9iV
fsKKKyCZeWjpsTGNOPBU0lGOxYcqK2XIkmmAZUfykENZTMUSAQ/OwqytoUku
DUsJ4w16Mn4jY01bPIvu/jOPaT75HCR4uLInKGYRw1qrU8BcMWsjELR+XEoK
EqmbD7D+qklqrScwdMB6GRDRfZOM1DquUqqUz7JJhoJBOC1qZpyMIa9XZOyd
SzdKHRWB+BAUHxdFP8B2uBj0BeT06Qr/QK+jKs7iaBb6PUSwAFBZbvX5a4Jw
P2iMX8KXK7OnC4tSrXMuRCLBrrjtGbr6Qm6VidIQKqpVUltngjdGqnBdqJ9P
TQppT6ryM8KD7f8EiYAFBI6rIciv2fV6DdhrvTWrLoAOiMEp5E6ilJm5B3BT
4qGcPuI6lIjCnjFOiKzkTdd4v2IEf254T64gZA4jfAGxKr7s9vIGMx52BJ3i
BnjktD25lkYt5AHg3SBAFprqTpzh+qYoXxVRdyD9kh7Yqta+N/aiMOkIyk4A
1JH2drwAEjOtAHX29UuOP0j3/gCO0CJOhwQBv+SFgEdOVSNLEK9/rMrt9F7g
gNuf1InQMmj1forxoyO+MNvkiqgFx9Hzg8gLt8J3S5RidyBD9tVV3fZgDuDa
x481VuwGGrfl3i+NF3S1Ix23UfrpSHfIwqvftgt+4mXvo6yMwuwXGzR2/hrC
p80+j9E/cLOT/XX1R4GXiNNEWconBUGDL2w6eLUuhuFOD9dJGYGMGRY8SACp
2Or+W8oBhSyj9aw/r40nm7dNfQOxlHwa9MqlGnyfE/wae534zWZ0VKlnVykL
viQBiY5JlkLNzuGvPN8hXPlZcEhve/9Y9iGLTYHq+lckCMWKb7onUrCrU+XY
b+7bX+brM6da0WAeAUkCzKYuEgm7sGxDOUsolBCn+SsVFs+NVafG6VQgeqB5
XfnO4hhB5L8/mKJuY3a9SGQihPLeU4mL4twhTyHn+U+BvxKdxgftyhUJ5xNY
uSctjJaB+RkpAPVh4+/byrEOND0rqOdd3nLsTrALrR+/lcfrq/ULM+GWWWVQ
A89JFkljz+na1JtOm+9bM4WfCRq+KLWjAsmWp+S8D0d93RQIAmU96/IvZZWc
SURY5UMZr1oz1CXa78pAe1gd2irSiIJ8zdCkv9D8iH641MVV4cqpi1xsDQJF
Zf0cJ1ke5gxbBFpKQmSO4ZBeR+29f/UPPiQnPsIba/dcZA9N7i9AhFAetRWe
g34f2iboP9MLr9gaMFytQjpq1Jfvfc2LTVDmE5TJ5v4je/1K9nScYyR6pkGq
i6euu50jtlba4nV/UlLjB+6SpyJbrfAgc3GAEgymQ3p/ijNc2yYKNHwWt16X
Olb0+7I5BY/xkc8Xa21UPU4A0x1RAnOTPgZg9JFGEqh4jaeaNzVMGdxjixqX
783LRtJYe/p8HOBGu4oeWezYzp3bk5mq2/VmQXV9bF7XTzvNDPodvDYtEgbu
kNL1IoLbVbO/TcvxwsQ9d2ld0c3el22tjDwbicsV9sWLyQ/1HTgSVb5vo58b
zKVyTWetY+pS+z/S9YF2o1Lwsdwx/i1+UIV4E16bEc0xip3T3rbq2cyBHkPT
/lG6hl9tBgVN7BRm3/lckXHuV6tAipkRxuBSI3taEfT/m4MWzh/pBrATQsjV
rHoMsjG6WlmiY73IHyStR/7Z9SvkXo0Mco5YBYLdDVcjCAhHGVDHafuO8N4p
xgYFRQ2aThyiaBsoUv0kKiikn7lNzaNrwijIo/1YJmQH9m/NSWrlnqPfMHBg
Fe+fZ6q9T9VzX923O16b79ofmf6jLqibK6pSlwKYq7YkFj9k5Ajicognl0fF
lyN3A/nPY+LYPRL5woxboe2jDvA1tU2AEr5kw3rX3AzGCDUTTkh7fEATLLcU
Z+kKO+qAgi4bI306XQu+aOHFKXqgSEtBi3EerL7jozW5tEsL4j3xSPV/snBB
nMyw95XgpDn49G9duw1bgQmLUUzxnyJOGCF+HIYtLUYiykLi+sDHoAm40NeN
bmpPs8/puZ4njPlQtOK6GBSX/eZYsSyZ69+liAjluhtfR+I8sRzA9l2lS+fP
Exn8wGg26AjmugANQW+2TW0g1kVdrCk7Ws0kfsAE8wDvEheVHcwEQuerqn1F
eTYfpC6CbMG5myqubRZSBwgC9MQb3hcKpIh6tj5awCMWcI5Z1kmto4yCnpLh
pk8dME6YBiUDy/yZPdkFf+OptxrZuSUGXXYbhr/JyoyMfYatxNKm4F2M6sr3
z3xn8bvaMxPZtu6SlhRYZndIw9XPv+m1QcPcqgRDF1WFCvX2iTqivq9FJsqr
Xa39+arfw3Eg48h28Fv200jepovOhfW5TzdaGTZcO1D5x5dPaylqF/QzK+dJ
pPuVkrcIrYARt9kJgFVAXLGSfiMhH2KlpwsXQJj3GmRw7mj69OPmSXuu0POM
bbVdxW7nAvAxb58EdNCsiD0H1uVg53w4nYlgZYx3eQTj9iXIkNfGQg/MYSks
FKzfLs8z595pPYcgidpG00TXfcUZvO4q05RtKmnMbKDGiPXYKznyFOinmvJT
+zUdV25yUD5cN3SYtKzGNpd75w+xfG9Op1u8ETaVk61zLis1Cy6fWKSwnobk
VGx9hHT8/rDFhg+I+HikjmTWxlEjvS9jGCkG87bvtkOWJrJsxhZAQ0uKSDTD
0HTdV31q/ThaiRhMW3ByGr2iZEQYaSES0M3S3jDsEKqJTraWluKhnVBl+xoq
k85saSGtZDdI8xG84LqjbYIvhISAty6vGW2V1aVkfADiqDTEMGmhardd/DFQ
7gmDjLbedbsqxrr/lfWOesftuJ1zVOY5g9h9sdBheD4y/Y6OTQwFLS3Tuto9
YiVwysVhWqzlRXxLXWT+h2cSaxKY6Bec9Xg8A46ILnMX2hsFmhN/owoOGDlc
2/vjpjLfTeGivxwBlqu2Ov8vbLRv8+4lifqQ2ya+v2t/jwefB6hBJqp7xW4s
56NSdj5rTNDN6XgYdL8oSj4MCYgJIOFT9vxNQz8N2+5f+iIpMKqUBzUtUykB
v2z665+NkZsHb+xm/ZMotWI0SG19CB5OKJiS9H0EfosqESw9R+0xZw2XPoxl
TW7iWi2GvuQq/3AItNlaiEK6jGk/k7cq50Nv9SMFDqwxyYKrTabZX3YHHmkV
wPBWyerir0usZBpmaKqbRG3N7x/BIPD/gusiPtcDb1hezoJm3xJk5s3VRbgF
tAhpwjgfQYjHgQf5441huUEX92Sp/fb4PhO5A70Mk1fdLs6M4FiwI31e7gkT
9ExLXdJbioTi4AVd5KnbwN5GYM29NQ/texhs2xRaZc/F49UIlYABVFtkTa2R
Pe28P6dMgbooT9MeUIGima3jk1J28m7cswezUk2y1HO59e5QjQI3j0qeOquG
iVcqls3Nvb3wPyCFN+bYMHPUftcHPl8DJjnYqR5eRUCG5myZ6fwGWL/pd/XE
Ar64u+3zgm6+uy3D96tLbYtA8wpOfus1FJ5TdO8O+XLNG+FopfhYpxKfoId2
Gl46I1T+CAyC1IKvPz57CZxY9q5ve0G9BzFBTSmMYAEekb88YQvYm6CnucY6
DdYbNh+Y658Y1fLH+HAw6olX/YNpEgdNvGzUkCoeIUqHlenV4aiB69KDXZOz
Pa8R0IOlqbGEzZTVW2/dKNewrFaXQlo6luli3LoFLVxaJTWNfzTq7WCd/eo6
ZOEorXFpV5yRW7PK/6JuGmxsCgujVHGUH/o3lg4hfw3fWmtHIrFj+xSf6d2x
2wdjG7amKyHUr9ad1WNygzyG//pRT04TEAIa3S0xywjqvEXvabIPoDhwHfpZ
bLEtZrwGznkZ2z2rFHaQ0Xq5Ol3wmh3cgRw9de4NGmJb8WGTeIxdXf9LbLZ/
1laCmDpYdkdjzWvoqHehTjDEioY2puvsqMFFBwwAunZx+ErzXqNVANkh1TUg
9Cff8QENXctjFnn/90TyqEiDgdUGZWmDvDZOeyiH0a46caDBbu91irqaP6X5
LUy7oSqiJvF2bfWxByW9jzmZcJ3zzrmFAwRr61WBDXQydUsVhvNNEwz0YNgQ
JIyKlRyNbb39b0v/CjwTD3/iGdpUzlZxWi0Wtwg+B24M4O35HRhWNjEqDEWR
bbWxhanuqNM0cOvXFkm6YTpa9m3RUPUofS9k1EtR36k+ACTPExlvu5fXkCbh
ABFsF81Jf1vQdRnpRcmIklalcaHY9G6QAMBN6MXBBbkKRFpAjHtdyFLFDXqU
R4Z29cas1ITw9woS0B5EdBu87t+y9cpA8sy3cFFGs/t7SNlnU7HbcdXU2p37
Dwtw8tg9bO/hnF3PRzMyaIGttudiVmHqwUkAHL7krEL7NTvArL/GXMN3LCRM
uiqjUblTXinYXquY8weQNSCAg9qNePBotGKpfucnXC193H3Wxc3HZFidFPKK
eXmWutSnl01Ped8o/sCyX1caT2++EPGk2ONWAjLZMJw2aVqLt7bkPiAdu8OH
KiaivAaWBlLSHG2MaBGMiT228QxWtfGLSiLe2IrX4Yauhd5Iel6JCc1kSLjc
E4eTN00MPBZydMtRZSi0PP3vHa7TlyssFTFHMBrLCwqWEHDB2VOKUkYbtAlX
FxIF9BaYgf0BQN9c6WgKPhGu0FwQP/QE0cD/IyQfcw9CDYMM6dpOA5/ba3/J
4V6C8pCQH7blJsPdTKHiCb/l2izKvEtbdQ4FQf1IV6MQtp0T0W0UJTM98EC3
9aq9Cy0MhltuQ0OUK+xVEEyvp0Auw3IQvfcxNrTIc+aEUobumkgX1+jK0zXh
b8uKlmv9I/42AQFCU3fUayGQzOC71KWosgvpFSK31oMgh9XJktyD7Yk2p3z8
NGV9jnftQvmFxeQNXyhXfEwXIhRbZRvCW0RnfyrKgf2MkZL0PfeJDhZgqTDu
+kbPnG+8PoHXtjKGuZX3Z/EZ1vz+LVqMm0fuKqQziPWytIuZ5mTUjiA9ITCF
qzxfYOWEQvh95pdZlWfq57A2QmRwdkMScOhyDDQ4FedovjfmudMTTRJroyVv
oeNMqbF3Gp8xRmwOwvOircWekWtyr6dplEH+tce6vJkCy1Ercww/8B1V2DVZ
+XKIiEJmfLSAkEKZWmgD11BXvZIVUoQ8EVDuH1TIPDk8WE+8fvOlAIVpOil1
Aol92uL5GXlWlxmtZn/oHahAM8SX6XMVW4tZI6oypqVycDj8BDo+SPtDk3Rk
bomTbb/8tiAgBYE3giRtNvwdE5BY7hdk2ng1ZgP8zwo3o4JPXrmkawNooz/M
1hr/oEdDUJKg0dLtczDpsjK9LLtq8sd0F4feSdZPHOHiia2Fim1C8zneNbZB
vYGdMnc1SFPmxPXmzYgmyrNs0AdgDtM2BxufhleqjIba6f8NykWSEquPrfB0
a8qQYf2HfpVH//5h7321/eCEnnV1v6qXFDYwNlo44bsCgEeMGw2yyJGkvOPd
d2xKjARK6qy2LtpaveewUtrz8ZfwwVbn5RAbNSfGwgZ+OVQ6gw76rrZUOnEj
LDYEUPofqf9Rbgy5oiRUP4UINhLLSaaIzXLw+e4k5rwlbWb+efuJe0IzNE/c
2UgzFjc76DB4S3bleF79lrO+KICZ8e8PrkMhmuzmiGTAuF/WSqyfx3ukEDca
NKSpC6OqcCwAVPIEtMaWN2lMdQzcEP1oe7IM1NaoygskoX6TVH5NV2duWghm
B3IBfNJTnNPOFzbJBcsqtc8gfgoDRfZc++BEWvjqCeAw9ONB6JWAA/EWFbQt
KW+udd39vL6GykdpEoGsXGHi6Oi43pFI51iZI//J47sforFuMylWEQtzKQjg
bvfDy8U5syZby+8qzVRNZNzOCq3TimToMwks3z0UY9P6sLmgtzAeGCSe4bjO
XszS0xuGal76bqZCN6UrxmTb+rwVlnZ/xFufjE7epE3KPzR93Wqhzt+fGmm0
ICgArTwIJGzS24sFFdQO8LUmaUihN0IoWIxP97jQPpmP9ka8ZC9QcluGyv6Z
U9pDq3LAcDplNK/LhXw9eI7U9MvHkR79EBeKRJYbHMHgeLBtHxfEwSDav2hP
PH8waeCbuZlXy3kM94pqgjm8DYTz91JHx0kZh4xjX/dYhtPA54h4BieLezCY
j/S9S4ecUshhdMb55y8FHzD7ABNU0BrqQnZXtut1/MAmI5bLKG0wE1FrqJo+
vwG/MBv/sNPnQcofFLadLAUODFJScJ3lZukT7Qw7OhlxHpYbc36MO800dw4m
FXHfW/L92MxWqSphOb1xCnLMqBtTy+u2k8h3AKGM4eHUZqEl7L192cmIvi5g
Wf4ARd5YG8jccMi2vf0ZbibN3DwlG53hzi6OpJgpW6hDqGr0/EKm9fWB4q+N
PZGqiSD/9J9tzkCfpLVnOHyLa52ZnTRCPBw8QJIzFK8gbcEmruv/BE5T6+4l
n16xojvAYY4hq2Fyxe761bmomPZxD3abKKvz/NssSTb8vv0uWuld5hMNfaVi
zgqIx5oBASEGPizbk3D+6MMP3n5MXb45nNXO9tlUwELuxgUlzyS3YQjnTYWV
/fpPvEgrIPFf4ZBWcOgMk5O0Y1CKoNNu+dAxx3/Q4yiZ6R0QIhUiDUYBWtQN
QM1EqKcAPplVAlJ7yxraxAOw5XlhoxjMrvWYJjOK+NI+TWFrleSYcKApp34j
WIBFxVnC7tJNo0WwxyotnQ4tYrW5KrDOMgaLhJsRAuf/l2EBVuhunc4H76VF
O6TJ2V8CbOKmIoqCrug3lS8eC0qUT8+O2HsZdo+k6+7rMM6lIMSvcSFGc0zx
OwqWDH892Z6V+bPt1cYObKOel/b37UMwOQO/kdDoaA5Ic3Qahc60iW+qhstk
qlOvVGvSNYvWt6G31AelsCI18rjbPqOrkKir1PVJ1sn4MMB98nDrleu4wF9E
2fJaZzNncz57R6IBO/44EqSaUUmEhQkITgUqRtoNV+eGe1EspgN7IC3TXcYP
x7BmZlg5n/sFuo9ZDKknZqwGY1VdZ0IlamJGI5NWu5n7wDKN7pvtJ4dEQKOh
hNLkVN8klVEEC2dS4i0kbtUMpoNPmjLIEvXvsqEFvww5iCbM2xEWMKpzeGla
bNB9dLBDq9/r8sGCFFzl9yjQgVaE0s88TVH0nB/7By8OEDLJbOq+bxWzEkLk
6TLn5i+TmIMcDC+R8Jbx+4xMwbZXi6tZEOLynz4/zNBhO516T9y7Xq/f7o5V
jPrsH6xRiLW3iJs1gdwZoQKZ9Oni0elYCLnU1CubKedchzd9zRPXzLTw8ZAi
GJEPGcYv196LOTxYP+ljANe+IxUWkthI8K1V3rNj9Esb3R1NcJcEoCIgoxbW
XOFvDDV/jAf/+/y+FQA0rK5YCnJyOFU0wJYBrpWuK269MaykiEnAnQDWNJfG
pFzmF/8ZVZ3ff2agYc1kmvbPM8udzgGHlBpE+zkZH7ChR4GoEOOyc6llWxpp
9zTMo7lzN8xG9iAkSNn63sFwibqSf/wwlyyMOF05m7RPF/VtYo8eqkzJao7S
NHDBjw516stNU85QDB1WTn+GG31sQgHwi5PcluEkSEfZBitn1TFFxEsBlhAX
tVaUK3LNISRzat8KCoMXW9K5sf+Ps/suqfcFVrRiSGkv7tXKzxgU0K0i6nUo
Mtufvlpd8Kx+Yi2rUAVSU3PzOiwSY85atml0K7nnT9aqlwhlH6x7vlQvnVWZ
Fm+jzIMLFTvJfBxVxN4VvWq9qhcXm03SIwPrA/GkCFa93TF5+FJ5yY7hmLvM
qZ4MRvx/0lVS16rXQMhn0SULmkOdT6fSxHFtak0ypVtAAzRWwzIeaGC2UUFv
LoGDSKPThCWITBSOYKGzEHIdda5zW7AWJlKF7dCPI3jve6KzSuxWfvAmZ7ja
sUBURTniF9lLxNGrRglQDFPSCWMknbggRNbvAPER4/AFEbXNd5uRHfMXHFrC
MgK9JynIPWoaJAtGxG7hSVFLv2O97mLMVQBH0S1eTOaywmmwbz4OLUlk+ZKJ
oZSi8Dfu2ry+QaIvVbWG6WyyJnkIsIhIAr2gaI0QlbY8oe87cvBk0tETT0QS
7VPdqnJAHTcA08U5r0UXx512ikgoMDkO4ubyzKyf1bKgKneGm3xigGccO7PY
8cJBiWVNmhsEPf4eTThxNk31Nd9i71cuQ57RDKuj0MxeI0EO2m8zQwZ+6DJH
4PxbGWzGUnhyWlopv74JMtSoaASHvWYriba/+o2hWsVPe//Gd0CCfSbv6lJE
ih+hIk5V4WIILYgNdPQhXW5b4prHNTK1OssLTeI/8gs4dmzkj/Wn/C+pT06M
tGOq5CKUWv+J8JwnBXXCCxFsIUHk/u9bPhjCZI7wCwJkyejB421l0tGnmYL5
W1HmgSXh8AR+v5AGHTwvw0C7P4PIurFdHl0WvxRG3GN3cAX07sJ2cIgaAiEZ
42nth1GvTiMNTqsDLn4mRVpryp2c0VJ9BEe23dfmTSAv7yGwYhI353fzVy+7
6R8CHYR2DB0F4JsdNSYOi81TCNP5Z9RErxkUMK2GRbvLR1FMr3TWSwI5QX5E
YmNOgKHk9+fvRG3Q6yJC/jGjwcGvwBtTgc1KF+veiGe2M9a52UYNV5wUBakw
mGHO0t+ZATEFdgcyCYzxjidGsqv5OXEtSO3rDZMKh6HiczJGYp1IRHgQBFQK
JqVT0iqExoMJdWorZXnCZMCvin59mU8nXmpZjCjc73cS16wKb+GrpGk5cYFR
LQflmyK6YPdtn0V2pCN8BhsUbL9v73WgZzpOvtpDhGOvRkE3E0rz49mJP1h1
UhMc4AMxgw2YZ/6TQue3UnK0F75zRimn6IWrbzjiFWq+zR7jDOegV1VihNLN
0sIMcH5sskNfBY7qbc83dyCQgneaDRS4Svd1wCmjQnPyfoFXKhlbnzXf6sZF
LSWpIEOJc6KYxddoaiyQscPEx6Y4nvIoxIorv61VGvJHRSOG26xPUzyitxWC
G74LaJHZXiHB8LiGwjaGSMgf1czSMKKTPK4jDWK3ToXbmEscAJLoSr/7NW5G
XYflNWaavkLGdslJi46PmEDaIgG53cX3qxUSiZeWIQQZpbbrMuSkqMCBCpWN
3PTfM2ddd03fgQLJau3UuyW/xxE8ZlauN+3KZ7P4ePfb4RnOt29EkcPGJUmp
sAfoPA//ofi2pWRpbe6IFPqcgKeYqVFcSXuhn3eL2C+/VgK2CNRC4GifieZP
oJBvoY+wYWOzt1Ef6BKWkzW5e06CZtmnyiW7lY3GoNFvalKeUmzvymuG/U3F
BXFA5DVyNDiCE6LFdJG8NdH76ET/ajuwoeX7wGGuD8+G2VP03GZ2G4x9lgw6
MZpGqn+0f3LlxxsuhthDhkDGfX0sjXRgsLUi7NNZvZ3T5QM0XsKEzODhEg/g
A0AO5SxHngacKbZBJaCWQsKla5OHT2IDq2LlUV6TVvo1xukou4hnx0r8q9wA
VudAtBxBBV4tXDTqEo4UDwOLESxYf69+uEuH69c+4Ez8HCp6Hzb4QDUZrcU2
8Z9STvFVcvk4yZltsI8NGsYDY7rx4O4VORFWscxMnEwUJUHxUg2R7v0qrIHR
Kz3O0/QQ5Zns7iqnZYvABQFbe1hkp2S2dwDAqektjixYd4m5frL5MMF8EUzA
jhNRjRdaYI3u0y0fxOxRjQoha8fofy3aCJncmjfZezedHyYK8kWJ4rr54QbW
mbxRkFFBNb5DcUc+WnMdG1er0SvLnLPbLvNgRIhh1IZM/f9qWqAiz9J/ptYZ
ZSfRA9ke1trR7lXyZP4TfZYJYjWyOIC767jDhTkogS6KsitBJSvUeXeJTR7K
TMR/FlXtfZHwRn6YfC/O0HbXiRYqyQXcBhksjeM9b7X8Y8Skq1RvQTNQ9iRj
VZtnEwJSmuRgpY/aJXQt6Hvtb1lhTyJxrq2fJtZflqpVcgu8T7OvREUrzRex
rs2XnR2R+2kKk1Pg3u+lfwdk9YEU8vgZYscLEMkHQdalPpC8i3GzwGmbwXnd
D8ms79MTr/O+V/ge7pF7WnLxDIoIUkOv/jAZh++6og/d+ZE7d8UKw1nNMmCQ
v8gwnHcfWIycYWOQFoGEWgz1G1UPAUxzAULDWSxO58w59LqfS7sllJCs1tpg
bBUkWG5vdCiBLC3Fw5wTSiKeyAaCPCvL3Z0HmjzLoOLIN4K3xY2hcGruohYZ
DxMw/AdfLl+4cyszBr93phoBzziWroIg+u6cP9lnrovonHF4+Qvfg2pDRPV2
wqolixk4d5z4fTkdKDzavtN4YDvB1uu7xbIsPf6pNQcDxA4YIXGJGBV/qGEZ
D+eGLJon7lFjd+tuK9z//B88j1JaztGGnhZj99fUn9/Q+xDOngYD/wsCy/Sh
r6DJDdmhLd67xqAhwUtxb9Jiq0GTLhbeJKeNIKVU9GxMDxvx76uWJUXciDP5
L0x5LnffJhXaxuD+u+RDMqpCxFcA3zAquYdk49ZojJGnzxnYCSIXPAnFrP7v
+6IOqUpi8i0Zed/n7zK/XngcjLIWOg5Gik2eb7T7N8lWVKUhgtqsbWL95WgQ
EMKBqZavoNs2fGqOJBJ25PiJO5cNfMyG6JI+bPZdcnwHAtKams+K1+qwyMFE
1y0GG/EVn4B/Kzjz25sVEShAXkeWZKNhSefn4FN3ogsftDWbmYUq+dAoY3vY
4fh5DITYlIJpd25/EJQvW+wQoWQz4yanGTKrXMJF/iR91sEv4ArnxFwLJ+be
smy+I6zNC+C00FVfXDk2Pp9pJoyFLk0k1Xce7Rm1Jye6uUwLOerLmvSdFCjQ
4iwZI/HCEZqTCE7L+ztcfGnIzglEXwfKFc3ILRbAIsy2p828j7bPamTQvjQ4
Ymsuvyry6fuYGe/8Xh6J/b+ypcQDrvcGzMeVdzu5My75GWc9m3OKiHuoOnDv
7zimkkCEh1+N/0Ktjo/sgr8gLOxRRort4n3sHkyRT6r9M96P88DV3NHV1dIh
2HUiGWWLOe2T3fZ8rKH6V5YDDyGuiyFauEiI9ZB8rpJfhbnzVSFaYRGrLkzE
C2YVIw5OTy+DZLFUIFqJ50KwzjNaXDWou5HMiT7yc+Gg7rXx3MHzzA7j8Mm7
Ez5iPjjLcc9WxywgtyoSC7NHKXyYL8wviZBq3X9PZz+cB2KrXwtC3e/rdvmI
sTC6/X6YsO/Jl4iRrP5+5/CdAKeWWXYmJkTBhmn8znPz3CM8YWLr6gd4YVcj
JnRHqRcgKb3N5B2WEkGzA0OvCOjBETOkE/OLhTKEwaiL8QltesM8YS+rwm5X
w2LPN+ov5idC5foCtBi5wOiNf67EXBzAP46FIt5O+qow+Vt2UvmB2JaOHWmy
haR6+dSabnTdVW5r+uDKYE9Z8cfsh/+TN9ocKCzPNmaPIoF9Pse+0is2KAy+
uvElkn1fzESBbJkeUThKjl3OoZzbfS9hVDSrCbj9j8gzBjpbvWT0pn+uoGFV
o+o7VjgwfKYyLBTyDyJhDZaUvSqhOhR7RTGAIOzT7B2ygInj1zJ1WhBl1FjF
EhdxCYPL+vVGTmI8RgFIejiKC72vGB4E/0dfnPlbM6n45ZVWwD+FVeD1hgE3
11WE/0d7uAU1MexQt0X42sMQ6P9Unej7opV2yERe1sQR6pMSl/UcpvZo6mKn
m4tT/391BiYBaOStL4xoTjXT8YmfWi7EPOupe7e5Ydl8mIBe2aUOs7qMx1zE
rwrjrM710cnNn8jqCPI35xjcmBNSVy7/HryP3M2oGBaGgwuqoe2vwKVi2ywb
f1V4ZAbR+IwedemD1NWXYswIVZCIwS80ad76PR1k9iAkX9OXacqx/MngJMTK
z1gXk+Z2HRbLaZgBkfxI/xyLvus4OTeQ1V9qxTnXkMAekk5HaZXesVr2TZkr
6RtYUin3FCfgmENOSmOyotsfnugJL7wMe0xwSzIMl0uvNx2r9hY0G6mwjt0j
hJ97vfIHr9bn6G8XLv1BPUp5XWjl/UP0J1h2VOLF4Dj3QxfWgT1OUhgkKJdo
vJg4rBbDSneV/CxP9WAzvwY6Hm0pHCxVCj3AHXYaXGmuMrrr3rHQNjUtI5d2
9mKsRYYun/hriKMIg/DvlQO9ncF2GsexYBDo4CtFzQTM6LASoLUBRcJa4W6I
cMGtMzcVR0xJkUGLdGakjg6ylWDceH25O2eCWv7c702E3X0oEYHeVkOx77iQ
loh0zuSB3mPC0R5mD4nIvBACCSkfw+FEAvfOXkGk3JRmuFAeB5NHNw3Zy+vA
ezlhx8Ui6xbTsE3KWZI2lIITnbb/QEjVm5t7DxZ2Jf1K7h/fQA4/IvmiJZ7G
hXrx7NAldCiko8Oi/mRR64zBfSd+n9r90piT644n3KXlLueUVfNKb6PyYO5C
eT+/57ZPrRKb+2iU6J7E0hXajuP2hVu9AbuPZjGWX6XNBc0NlA9t/hnYsBYN
Q38Z5CgGbqW5IJAbEMEN1GhYwTcc2vxy+klU6sbeR6c78dgjRuy6gIP8ymla
KLT/EKLSyFBL05QsdBqjG7YVa+DoMyiLHe4qiDSRzz85mld8JXjf7rt68sxC
W1r5o6XlK6MVz2Ra1aWE4M44VdsBw4/hDDoNFYcnVfEauWkEjN3cOKtHa5Qf
X8pqJhn2Oz+GoT2kZDS5HcX+jFh40eT+8mrAtbzp5wzBhv5ufWRWsGCxaVWA
n24LoP7ze4E6BIXNYo6DP1baxxGGLm0+Vo56qwarXLma3LXscphHQfcVY7hl
8nm5uXtYWaDf6F/0rFaxZV7toR63Oix4Zuqa4peTSHFValxt6by2z7iGOu8i
7J6XtKRBNe9iIb9AHtBtZdTElgiKSl5w60COPEe4NsbQSDuu+7fERDrwIvKc
X8W2NPw8mwONT90U0jn98HCvUgMOcQCtkHGPALxx0cwR1INXBYfPZFAZ9BVY
ijukm+a/2uohP4RoTYEB8ph4DwDtmQ7Ng4Iysnnl2XgpuweSqC+r7bSyY6si
fPwF5i4trPFlctVkao6BbkocsWLPqzqSUCuOhCT+TUC6NaMMNdgzKNPfrfE6
xIKPom5hEo9qRWGXkT7whG58T6rO0rIFTwx/segqh6UFaSbAUoFYALP9KF2D
PQPnBF11/W6hlA01BMUYCGghdRszk6e2gHYRrnzXxPUiEYY7qfwjLLllzN5F
vCDcItJpLG9PcztgQU3BINWkDgo3sXFOrcg/7J1RchvEJPkKqdoyZr3VkWGt
2JGpJqgvJektERLo7zXnG/N7tt+fcfKsDPS+C0hpDouR/ffHW+eNNkllKiFl
NOtznNOBo0fADCRuink1pKL2bRDliyKIrchLU6bW/x1rgUA5RO482X3FKPPx
IiOIscR31OGIBnxFr2oKVVJo6Y2elOnC7sUiq1eZoVBG7t3pfuJX6A1F+0YR
pQutVSrrstG6c1IMKs7eh2+cwlpioxJntjIesAnf8hPt6fUPhJHoVowbXsqy
l+WRCJdTZXV0yPfrcbCc9ZgEy12oi+Go6hQlFZSlZKypDDeBk3B5UYNW+rtg
yd9wpk0oG+u9xRkTdZ8FNJ/+ekms3xPbCuCQPbw9SCHLOSsuAhLk0a3b0kYM
H343pR92i6esKQ1qxBRpWDO0v8Z5An7fZOwu51Pe81J4W1ON3LAtphEO/6Vs
l/800UgK34LYqgXdLoAkoHJItb8rTCZfHIzRPh/eeUc69YPEbUwwP/Xas9PI
0YA0hZQf57A7XMiUPPNUJL2vZB6zfvBEvp2IMQJR2OmbSefLEnPwJC0Nj7Z8
iJT/GIIeVgW8BHggg2IwtAfTi+geVxVXNMv2RAgMoQHs4A/kTALUUcgtdP8K
4rzEEANv5GtMCZ8pDDFQtIahv1wZLxGqdKS3Uh6DUo6XCCdzkmKr3TtghS0/
RI8BtVtF8M7KGey78xu8J8vkYxLgCZEVwpwr+Nr9ry3C2IeQJ3o4cvDGxQb/
ovGalgf/d+FWqXS7WTRumo4dE3e0SlFos5+MXrWa3HdmmNxFBLK7ZZQLfD/Q
UMZe79UUNPxHRZS7/czKEcHp/roXS2zW/BMi49bPkCZbmnVjrbLIxKg8mGiu
mBLIJ9QEtoH+huh2SDKhmHLlE6hJ9zaGSpMFz22BbYjIM/eYpBTDGYDhrqUu
x2ehzHGlKkF/8y/UkEtRJrTyX/ylyx9bXYdRHJWdn9ONvp2ZydO2r/M4EL9P
V2iFG1yzwCwFod65GqC+Fi1h8c924Fu22NgVtzTiyQQuS9yvu3UnxQhrbzFY
pL0/bXcl6yL75A7eKgaz0ytfN7JvGgRkdM3uyaRsVrAVx0f/Nj/eNrbgsHsW
bt+O2GnKxeLxMw17W0ZRZ3z0Q4tN8Gyc8IIhcDCO/ovk7XXRKhj6PmNymUTk
TZtLnaFHOsP3+je4GBQ4ANH89+9YlP5dBX4oG614DcE8uhsSgDHqnWNsWtK+
8ELGcxXwB7HFl1McN7ZTK2L2VjMQAPeeoYV1jSmyQ36gc03G1g4cPg5UGr4S
E5ulIcp4K4HMjVK31H2vcTu5b7q0gI7TrmRaYfgnFrrnZBIkYZ738IpxBCb2
fLbBQCHIMnfhwnPSzwn1myMI+3a7r0aXDPmK8L/8n1UtzZcsOlQMl27JZepe
XxWTouxZ+xOnMZrw6+tvchigit5C4B/1tKVR01s+bcpCxVanKBYs+iSdx0qX
EO+CM3kxLst+Z9XXHb5uyCuBgXnPfON3I/AoE3P3sED8QDmgygWm2wh6f34T
nexwpSTvb6MpZJ3AE5f7A7btJSbmUoRE67BA7H2zDLsz93VbERoercYPIj8f
zj3hbHJGTElJOKaagDFZB2L0meFw9mQjjqLa6ikG/aJgohUaVFUHk+MGU4Ov
4Ly9R0AdWVPXPeRhyF6ciOu9aktaxe+51AyuHGSCEIt/WCWYgNh6VHRPf8hq
0UeNg1+nB0wE1WFkLdiPEcHxTev4t4mseEXpzugJicpryiMp/CxmKy8HdgYZ
kVHw0+SBzrRZ7HyCrrbMZZGs9zsTaYCjogBeQbR9CVVCkksl3xRHa9dvVfX9
KrAi0xEfmcmnSRQ/dNWhFxcAyMBF4klOjsD2ljbTft38Tx09/Ax9gi1FufEI
Bh3Wyf8+w6CDS5VrNEjeXN2/vaBn/JQmDydjph5cps10UgWRdXEFNi1eWhPO
GcjdfhHBwNQ3q+YIcRDIiUds4a70pEQN3DbIkohcn9/fU3Xo6OGFdan3nTky
ssNOn9rYMirj9AEQ+Hb4vwHIOEyUOsWHRy4AHyQmHbiLatIzNHAnjqOKyII7
IzpwlAKvBPbzx8miCEtSZZgPzKXik5dt/YFXRRS/9j9aDlczYIOmHPRzPrFZ
1UUjuKDA3+JHuM6l9Zcjly1bwATPuLfLrn4zXKGXSZF+Md8dIvZUei0D8wS3
mk6y71RLr7Z5f2r8e9nOWmV5ixnMGs5YtiFMP33JWAqLDP8HznwqaSncOZ0O
9hnbVOpR472BtS1eP/tps+eXOcksMqKfSJcsq0+ngR8bpi5iJc2dhdduP6nk
z5/AxB77J2RV9+gIBnQfKPXnZyo72EQTqr8pJG7BnxxyDQduBS1WWxAGamch
LijG3Qg//zZe/ROlBaWk5juQhCtK4X1SUywyq7VitiM/xi7evC/1MItgV31v
mLyk6YJi7b6NY5RHPF152i9wclEqY7gIvdxqiRCAphdyamJty3mvWSm+EYnM
Am8RU313vqxlX9pb7wMkA9hnZRkEp/0aEPIX0iQ4BgrD83NMRAbglxQ4hr3Q
oV1xPiW1/Z89qSSqzdoTOOhx5FY0aqbMSn9iGsBQ5U1NdejudkeosLEXxPXp
y4dBtjRmV1p+6KMu7reymKdb7nOtYpaHOgqsE+cfkQmItzrGKBUDomYva//d
liKMfUNSyi4i+sKKPlleTRZJ/YT9LX+eiFdVHtq4hjKO3ETvQo4DO2ecmE7S
Y5rCAlTwCy1ReAPH3aM3MntotKgbO794gIbiiHtSkMqczIzj+xYKC77skjjy
tkiiOKKTYYU5bHCdXLnhu/SylHupD4j+tWB96T8mFWI0cxlFnc2XupAeaChm
gKJFeVq4i89wEzznvB4PXB0e3k9DhqDSE3QtwOAK8unoMASvlWbZkkg11xjn
Pcuegg1LTBsCrJRrwnTS1xsTp8mRhsDnj4RxX5YmIZ1hsw9FUg4+gBtUbAmU
t7/B9LKBrhBXE7aP7cfPPBPotHJvxzaVzPmmbw8Vxm1TtWW0dmmcZ8H6NztK
Jt+0zFUXKRMR/U/q0DT5Y5GdcNLJSeff77U4mV7j8WmRnuYP0H6cg0J6hhNi
eze7amOKaf9BJZjwz0W457irWZbXfQSBWMTvfdyL4FBMRnMzLeEzSrY5cYpR
XMBlM/fvmePq5OqM1eBQtsdmHz0geKb+w3GrVhqgFTByH0oLchVWvd2miDaI
CHdQTiQv0sgj6nVHYkNkENyEgEIA9CiTh9M3OkLR2RhVVhy2fH31eMsi+LQR
63+3tKbs1iy0bAXv91hZ+arI7BSkkwXjhrrEIza6VHIpHyo6uYAMwagRA74O
/hrHRSC7VQqd8HJypnGh4tlKX3QNd0C0VKbFR98wPsYl+isPIEd8cXMR2viW
+n3Ef2jb2dA1dcW/EefU+RXC9NsM8Fy0d7WNGordm0bcgDtZl0yuNYNiNNI5
yzLH3sQqE0JiU2z+7i/wPaH6iwV+us1afq1Hk5vdVzjFgWDVzXe0FBgrWPje
t3XGy7cf/NOQPnmUCar9/NERVIZMeIGJ0Z/UPNyA6aVaolQb9Itq+gaBT1rr
NhskxBOzXgjEBWIsi1QeUPHabB56N2R96z+xEMDuekV/f9g99FQoFk4rZCYP
K6ZeBr3KoVpVWFvsymrTJ7zO23oegYQ55C5JhHuWI3purvrvdFLSmUtaBQW2
1cI2tClqGuyzAHc/xVRVCtkloekldx+KHveEa1TES3tahnhOKunI5vuEtI/L
43FMtqipaHz3AVc8FsKOl2W9ohMU3zh5jGBM3GFoWyUS2Ii830eHi++RFbWn
1pHVqs2w3uhloCSuvo86dJTGSpvRho4WCSIwBOH2CBC3PF23KfjfrxKUrjWI
JMMA9piCEbONNmta4tbqqzTJcy1ynPE36cWcCl0PM919ZfOmmXVurGfTD0cD
FSY0ZzZ0QfOdb70SGAhfDDJOBDnvdGxi0Do4Sioh3STT7oVmIqllU7WnDWXz
Gj5ZVOf1KUl1FZu3WNiXzfFJQXv4qCJHYm39/ViIII81JSBqs+mdU4mERa+X
qPjVhg8KQRw4X+RecBlhqwA6CljyGtds/w1IhARD7lupS5l8U+O5Fm8WxvdY
WFLpOOsiqR+MWME75ypVm7HqFow9m9utCxglDsNzU17pMKyf0SjsM4rZUUu+
HuJjqB0WcjtN76KZ/gDhe5qM8NYBPj6Rs7qwOR10El8PZdM5dPwuoIASNggZ
nt4uZHDGgODSY5bxt8qdOm9PGw7tOcipaj2KnPgPINfuV62nifkqyMS2euZA
1QWSTIgbQUra70A/iVkaIIkSGqDWIUQ9L4Omiw0F5NOqzwLpf5R9Idvi+g+u
uwdY8E566lFyrIKO0Qh3JKvKq3VP2Rlz8RfrKZ2Re/NAz/fCxqnIBKr9m/fQ
gQx8L1r1kyLh9NXtoXEiw0ezZ/nrsmmn9iDhJkns4Jrh407SnSBfoqu3bWq5
C3XCqZG6cMPkpw/gI9sIHs9/adplz3NbJ2vOTjSNbQ4skMfxS+CJXsKZDHbC
g8vsiyGoWt2zRpTy6pM39GeVSZw9sCbX4O5WuVjDHXM3M+hivwsCOOQ2IX1a
tf9AK4JnRIn52dt7HuaprU5kuTP26q6PcTwlZ+2I8OyQQSjE7JEa5PEwHm24
zoTyFtySsTNR+XyKtTU3C15ySvfTXPRfpxETrvsBhiIssBRuTUX7UYMmrm4L
hObM8WOOkfp6WdafBBqCmBIkZ3q+Q6OU7rqs25e/JZBJTvVEr8zX9KbcwN74
vOQpEKqQRUKMMyK68FMD+afosP02CYbVqwDEac99SYrudorYXj8KxyjRg+D3
GOLEGAaNuVobMiM6spJNs20jq0lUMkiQIOxLBxqeirs4MWPFg9JQw4tK/8Kr
kh6qr2Rt5BiW/BLPb8Lv0ULtpxxOOZmLJythjwSVWU93dJiPoZI/sz/nWSFT
6IPSQskS6FIP/NrJd9+iPvw3cY77Shbns+AZR+AkhK5xSxsw5HvwZFsut0dW
mA0Kp9HF3XU7DGcSyECkxHYdNZvJbbfctzx0Clwh9CvM/cdxIYoGa0l77xZS
hrzw9dDBFfJsgmHLI1bhSnZ7tkGBpDXrSmrOKGET3xOqLvlpJjOOQqeItEjt
pBGLy8EQP4mwek0kpLmbccV99s1ONy9uKQ/qWrPrnhgeRbxPfAopORCXB4RT
lVx2ZbtIlfGNMdki4EAWzLASi9aB+mdSpSHwYn2p8YaAazafg+SuRpwyRo2r
agXqFTSF4FilnYnuPzL3OJxIqsBmNEw+YtPJt/gzhy3Apr7yYcDjwRRo/jTJ
px5fzEIDxl67FvQUcCPT34qTurmO9LntwOGkTAaAy32vxYsImtZUzxgeZF/K
TY/+jXbmj5cPJUKuNKjshgxRhuVKDK3xZPqzMhJPvHPGJur2DqxAsD2gw7Ln
U+1odMDX8JwmTfTjMEdSDM2V4QEN1np3ZSg7CuzbNH/7fpvaUhp+UrAjEO4h
X2KmmWzOppZD7m2bUTx+eXLP28CAtuNl4txPWJ0Pj4teDD7Y8q4bZ9y/JGU1
S0EDRFIQbuDxlD5BuSuA6oE1sjZxqxyjzbhKaZxYpwAFAa1oHascYKBGwSQE
qNU7cq1xgCRXsjB2UwUTXw9RmYWzQQT8JSIMluerFcRihxKm+PTe8udeIUa5
DlPDvcCEiMC2sqcPZUIerg5w8xv4VK7RGj/VY04of0/HaBZpR5gVl1o8wXnd
/pfOy4o3EbDt0+ItOXpp7Z3J2UeGsR73xiCC8CGAd4zKwP1x9lQoLtchTXUB
7MXLHn1R8o+QR6T7J9gB5ZRQBgWCqsooENE22jjGqxo/pIDGJgLt3k4kZuux
ia7HOXnN3hSfObMm5qAclMokyx/WImLve4hy9mScnGQACiyvkoQhVgb793sk
H8CocA13Z1zQ/1M2RtfLU96NfIbnJtquzx0BkH22PXUo1z4q52560DB4TTN4
qVk/EIk8EpllMv1VxvZfR+i0mP2BWQSA7rHO+mSVuDliiFVa+6X46p5yMBZc
jAZ6By9oK0r9QWajXXOQs888PVCTLz5cptS+Q+2jQsbFHr7NLj4VJgkhroF8
xNjVPmIHONLE9vuRaOKOJlj+55/WK9mkDF9lKkBKk2BSvWL+a0HVrtwASetx
nvotVcZBPhpAkdJ5fZeiR/V01fUzhsyYsFlFuPArXiPtIxrJmMxSlgGCHX7u
DpWtD82QIwIYvuSrVadXMIDlW6UShRjHD946+E4CYjtJNEmgtjnYPItPhGbZ
OVqJA4rH7oFPREd7u83lwfnkccggDlkTZcIDAdA1nTqpJnGcNyYSLs7GUvWT
lA2ItNG16eQrnGXgGJ1gTjV8FjLgRuWY2LK8r+pizOLNCzmpYYQAoXknNYOW
TXoNo82OQBdZYZI6/QI2/+J8Lz8gIovD5cSIVkMqSRtXBUZRuMnejvyIoh64
eTzWQevyWLx3h5uCxMxBmBmwuuAx1nvWnEjUoytAS4dlOKy1SAshsetnqKZF
YauLwdzU9CF/F5qWpuOuS18YIFtEe0YabGiSacr1DUNgIE6uyRlj2vHAAiTa
pNalaV5rDGeHB1SyeD+LFQDJQnAWXUFP2AJkdlrqR/6CDJkHOfrz9cUYNm/8
kkf/dcbLIlMA2XXdxTFPYFR4EsOboTdeHgJukSZG5qJB8zEdPKY7Y0Gmm4Ye
1s00U8eP2a1+KNuo7tL/8yP22OyjA/JoIgvWSworD687F7a+kbWBCmUxYebL
ewl8vjHZdqYrgJISaSO/PZ3TBx1pv5PNI9Sq8unRJMRi4YSCpqW8oQPjZpje
Cx+4SYg3cxqU4YpJZA1yCOFOoJRoMkfgEx1oa9KS+gogKJsShdPyf6h+lqeS
EbFd66gNOuyRuPoqW6E0OKeET0Pbg6j53TQtNAbSvAvBRARE77DPiBRPnbwN
YTGuQFf/tV+nAvyxxeqjDtxCwdSgvDOsO256McJ+YFpi04PvroCWLc3MMU/1
45ZNgAbZTmF2WgNLBmh0sgF8V0si6LKZ+ofG29LYB7jREJewaGswhR2b8eyx
D9zKlhprnlvv3Ld5Cch3l+gnH9N6vY9flO+NINH4EUuK62hnwywO6sAvQhu8
EqljHTCXnWbe30bkHGCGpT917h3tg8PA/ESjwsiAo/RuUhdBWe4+imuI8rZB
pBVxI1xqWdYvcYRP1TqMtnnFATgEz+E44ImbPN/eH5aJ+F31GuY+xMpLBY+X
5ecI2D4uscl9TEw1gyded2r1FOFJMvDDmj7Fm/CL+/O57IzL7FIZjmKeJRc2
Ig84VlnIoGequuTy6/D6NVcB3tp6KcBnwohsNkrfnljpd1Ohs0EksdBCmKE1
ipj4+TH6u108yDnkB+lMPKefXT9SRS0kqbEeJZpmFF6ij/BcfN7h6oXapFY5
wvgV7DpzmguG7HevKGcvPADSSwhLa7bBVie8asr7NVdU8vPb347CW4ULoJo+
AejKVWJ4MgIcBj2P9/b/uN1KXEEOsxns/ClOAkPkrkJ22hJRVDE+uv5lSKR7
4T54oT1Zzre32ZQGsnyyAU1lJemY8zyEQHaas9ql1jWl5rnjIGuivxeb9CNt
qRE/eIF9JAmvPpw7MNwBkTNh9/XNvRXmFtHbITVVFwxEyDwE0550zGZu/ANY
KFs1leJDT9r6kLMgFjkDbC/dYkMHf0tF0go8F3J6k01SN7/xwzZd1R8FpViC
BsXySHoPYbou5FLpBrg9dUpZNID20AhdtlYxfKkumZ3B/C8pc58yoPJOPmQO
N7K0xtomvDjivzHNnRDAyjis/wQbO07SLgFu8Y8OiRB13i64mkyfPDQTroIl
dJu2fleYNRTkiy4lgRhw8Y5WNOykltcM9LsoKkJm+ste9+0IAX7uXvlLPpqC
5NTfIe8r6kdi0d1T5bh9nHOpXozsRkSEdgX563X7tD9xZsHx5GIB66xnE2qT
9biOdgxjNfGy9MhJ0kDoEi6Gi77xkUxXnohLNu4aB2BsPz/5O+iDoUfHovJ8
CQFLuppZtwyKE+0R5puOB8EMYYFhfpec2md0h9ioPlMVyzj/0Kgc9BfBsZMV
CSZ42t39p/AZub2DR/0Sz5tN1TsgLVRbaGDxmybWqhHbVPAjm2E+A9bWsAes
cMWpoKWE0NflnwGfu6uHu+P8y4p9sCcIzcs6wUuIUXwLSsr1MlulMbolvveh
VjKJ4NJlbfVxB/sEa3CxQY64/R/1JG4ztX/6w/hmCYDvRJHO8+dfSQ00MGjI
dlTgYyJ4wP55eCEW+NyhPEEM8k+zcWap6XlItKtNii47oJoJjlKgJBsACBz7
gvPu9e86q2jLb0CbhSHVPqvERrWltlC4/ehPwTBEpfcK1qsmTWphoJ6x8C1J
JAOYBzUP2hulSANaVXihcwIg44qYHWMN0i4S5SztIeaok8+q3o2R8+p2oX3Z
PEAUMN36FY/mq8NYCC/AyBV+Baiya6F33Z/KmtuPlPZ8etx3o9L0wlTzOp7g
bLZwrW8JdNq/CONr0+3fmvg0xrkOCpKzzq/EnUxIs5bbfahLuQ/0SAef+f0p
lN0NZYwLJ8jmXeG8BpHefXTKF04U4STpkJebfzH9ge1dhnxhHOb+S1XpjLTO
3s9xEFNZi5wzHWLzPaeGnLzJBKx8uQOUEkNF2szThcLKsXmT9H4FWKaIwg+b
gr1owcaZ3h98IYygm/MDZobD6OVZ6PoygUP22P8mruB7BNjPVvMPvBMTNVJi
/9raxWAGSPLp36ry6k0+NtCmLMbCqmjI6J0ZceZHQiNT/cOPX65lQOj4Qk03
LLo4eSFrMCBOhlYdkQy0nPlUckuMpKMBt32SCPaUf82uWcKKJng6a+BtQiKw
nCsCaBG+Qb6ZxE5K6MTUc4qFEgajLfXsKN7M8y4wMj6NPkh8H4HkeOmgBns+
aTdcxp4Tuw5HLEQt3zhJJx+NDAFUchrJIadZt+VT/wo5ZU8HtphuJCxOzKbn
5lSkguoR3kofUbYA0liLladZtAaBpRk2+Mo+runhfClcb+dOSTgA7U5pnfMd
NW+aOAG8DwHnfbHoRPC5Rw7acDgfxB9CqFvmqcRkU6hs439ww+NAF8ZsvZlH
zhoABUz9pV1/9ubGkdJErSu6OBqpfezDm/KkHYy1HNtKBMYvEJYWWwBnI7RH
9iJKOJ6WIwePTHgigNi4xkdOD8YDTdipooraJ/fTYptkjro0Fv56sp/th0t2
MXx//GtD7gimyUnyvjgvY+AWMQsTbJmsNJq608YKozTM8fkOuc9LAVWeQaY6
e13MVUhXb4F67pG82yRGbBPYj3AV0pBEK/2IjbAlq446LdmEJZAZ6pU1LsDP
pCEITHReo6T7JJpLqKaNeXKcWLuxMfuCD75LKbuWAIFKrYFBpd75mQ2gYrUH
i1xpA6N3ecsZNag8tageGV+cH1DQjx3YWgtWOs22tQWdJEUJm8oTSUdDRrVu
bMwRQx3If0n/UfzC/rjlr0tBt+cccLJMpWg0slvv9BebSkcqG3LbIrMxeulU
m0iupqiwYM3dkxNqV4LVyYoeyQv/elxBKM63rN3z0Up6C8OBdzeAFV5wkOJe
6RGzIv80DsAPQ+qROpV/1PWXB5S97j9vuDgT9otBSmuuux3EJ0mmbP7+yPEH
D6azZgAcQb+cI5vgyYG64LjBMoaOSPPboaVZgJdl9cQEvI7M7OIoisk/1l4P
A06f26H7yPdcZsVwtK6znShT7XVG9Auwkmeib8w+usKmhh1T7XpSojsTYnY/
MuVtY8n6WsgqYHmNv4OiOMmTJgOYjq0wP1yc2cqALqVymEO8XA6Dv/WYkuMu
vvdGbsw3lkaa6I1jGaLU5L+xzL3YMtE8/ts4UF+5ocJW9Tt+X20G1MPHI5e5
a+HYzxJ3LDRUS6ynSkuece8Dep5sOf+sWLdrunTjg6zvEQ+EHqnvK6bdvNWi
3+2mUuKvnLGjitTbnpXt99bsY/lfzrE5goZSbWDbcpouqRv8oZwlUPscwzG3
N56S7ncaLxoSJlxNlu6jUeDsUNA2IEdgSnM9G5vGzX1pHPZehEJNSl79lrwg
K9YmgAMxZRn663e5EmgtP7IMHMywmWXW2XFMKHeMQuFAztFZy9kl8cVU3BbG
WBARUx9/CkKMQoxJebf0c+cWHXMpLzP2Dz3fujCMeBSR4KNC8Luo1MGPRhHY
ckSylNWjyKEMgdLEe2CxCyU0soLt48CveDz7ksm6LzQCKO2EosvKboXLlD7n
oiJ5Ugn0ROWF+idrXGhYdudGAta+KXo4ZXl7BeZmDXdA2SzB/jAfTQj+wUhT
bB9W1WZwZifOhGVlYLJNUToqqs4FSJYel8BE9mCWjEjbfBAYnoQ3qCyR6XC+
vL0TpzFBLMSoj6mdOkRIkzuBw9GCbER8X5vtdo0uo9qotPDg7/0wli0WI031
otyFrEnNB84X4zyR5oqkBjH+1MwxaEv90+1JtZg5hn/fvozyUBjV5BeJaJ/z
c2URyclhr4hrnmci35d6dYsSzPeOdms6owcO66alci+bJOL+vsZojCKbJvRC
rWj+68fUCzQKhhXZyqELem5lRf0CGkbPQf3KjJoz9HF4MKLWEGF5OnlW5oDW
eR+jYTmIXkSt9DfwIA2qpua5xx08gez22n6VGo7DQhFsQwM6rfK4z4A/qzio
ffVn1QbInnkmpGI2sH67bGC/gSaCqKnJQ74vpvH9VcG/KLDSOGstxLtiLcWt
W2YF0pmyAVZWZBJrQWLqUUjxlUSDV2Rrudbb7Ev+wDiel6BwslueiG4z8sde
abBR15dSlMh/TwMAdRU0dZ28W36+MZAOQgLPwmnfezOqgWd1Hy9myRlm1066
z6PGXNmiePzR+vV3ZMMELaX5hyFFDOXSWFTU4143qsapwMuNdYpQmkeYXnVa
MF83igVuv8B9f5tAER0KZAebiTJf7an7nfnW0ZhosgTteydgEOjyYopKII8W
1/+j1HpP2xoDrQym+vpwwK274EVshoc11cWJAS17WRgVYYbEAokL0GaLzOik
6osaEGLb6PvCyPWtj0Z7XB3N5veGeIk0E+IsGr45gP+pAp1H4eTQPL10LbHc
KVwc1AMd2i2eOOmVRCQdREsadsBgLrF+kmes1OrJNUF1svkbHrt1w8wL8GPg
T9MBIl5LQ62LtCeCjRRVOgpdORUKdCt65mhndeMQZ3rAvwd4Dp8kzRPUrLiT
adysl1qKrO3AScvxsuwHUH0OOafflFrlS+xU2pRfSIRim04EF2vjvhY2wNr/
wnP6AIFuycCVtIh1VhKMXUQF3Xrhb1urWXFh7+/lwtr/q8pMbUXXAxVSOSCT
xuzKVnFfTUGGADqLhkl9Frf4Coe3UqXWYLl3hKUBj73DB1r9mgv8yCrMhGPN
+U416b79L5lAn92yPWhu8nuuzInN82hn91GMwbCX4qm3JgTXO+qKqvQDjlpV
YxRBGdn+T6iBbAXi3P8WbXTicRJ8D+GMrTUmu3mz6/gEjQMTlvlwFS8NdcgU
zkvJfQauCZLbPFdWl4LB+pFJ2S7L8+ZwwoXxxdmWEsOSHeUB/a90qSbVuIrM
2F1HM9SJh8oDNx1IeECIkYldpnVGRseZq7r+H7FeysP/ROzgvu2HGQQkpcu8
jSezF5WRz12vc2f/+YB2OB7zMtAgWJ9cMUQjQifGJ1Ytzz7rP2BIQFdbP5TY
cGczREGaOd5FB8D5CPrQ9LLEYdFjmKuKp+Di8xT3ggFmR4tyR3KmYtj7ynyv
wm978wNfwnzdLmRWTHm4idmdk/+hCtAoYfr1ATJD4osozBrzt80ojDfXRYVh
rIHncmj4szdGGUGURVFY7WwJm+UTNuVIO6Mt7wpQBeGU7F5UB+LZAPOdlRJ8
8AaMO2ry5VudbyK1cg4ZGQ0gF5McOrF+jD3jfMNEuPNCUcOUSKPEveMZH6Kr
2WuytkJ27tH/9Pr5CRwLlOqWkgDMT6K+FKMC6sQrepBkW+Hx6GRatRBIiuAt
b//kq8hN0i7FyWWDgse/ay6dFRfXK3RSoUVjCqe6KaVRyQg05rkArzrTT1kC
0FHJ0tJVmvPvwQvy0PVCuxvoe1pLW6Pz/pTYTuBTmQbivlvOh5aVYSks2BJN
RTUECsYzvcOeIui3X3uw9z4O3BF+vjVyP5qLqa2RaiS4vwnT1tG4zYTNiizK
oX8df25svK6bTQf6fKsKf3g/qNI1aLzFzhUYJSfxyJfmKcq6ZrSKJXK513Uc
EmkY8C33ZvJGxt5nVZtfi1mQnXvbg/4kZnDCtrMhNnf/8HWiUYnmLftYFD6g
9BaP4bzpbe9bXZCGg6+HHGGtQ06FDCkskOXBiFHosZVovhU0WlQ8uqziC1mU
kQIhmRYs57JMNhNc6cRPMggNqVF5jQYrTfFYt+qMwux5vlIAodmG3TCATd8Z
VEZ7UyXQUJWqZkpa69Gx9XTn2BuwdBYZErQQAI5vDu2fPw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpej4BFFZ33T1XgzV/u6BkHAlmk5IuDpeppIku48O7xGe+YdNvv9jFEmvpjJdgQ6VT0INyzfXh2JvV047HlwqnYSrhQS9VO0bVSR/QfkaqnrwPHIwUFkStR3NggRZFCKbUF2TeAQ1XATesPA7QbJU6hL7tH6W1DoAYVCN4Zo6RspJfSh7qjtnBiTjVmfIAunlr2iVS7QBxOulj9QjrpFrEK/tYiUoAIqhJvFcZv+08iRXAD9xA5ZAVu4l+muNHJn0u3JcREva9XJ96ccEYXBC64HMl2Hn+Qw4oIFsH14fn1nZhUigQhBFNMiAFSwVoLK6pYMs1DTrmoRja15BQg28XwkSz11eO0PXu0sSMkzk8iuYHRFSCwcwYLWkvrBTn+DVqCywMe/Cj7zO0euyoUhnZ+jVcYb28yt82aeMZ8/xcKEuW9NaWkzYbketch+XTplKRk/L9pvvE+B4zWw7f7PqjqQsJX2jjPqmSXBuQrQ86tDlaLUJ1S3S+Y47F3+Gt/gWU5ubQ0R0o3KmK4HtoSuSu8bMSgwukMIuoSYI8CZfhzbWQSxmLBKpavYrSz90T0aRFpi40BORzQsj+BIgcDgf/Sl7jCCFRyF8bviC/67OpIR9idZHVUEWT+6FWCjBSN0JmlhyJxhyWWisFfBBvduJyzq2I3+3hIZeRPr2TMK/HwONgPIHR0WDMdjx7ToECbbx+hD1APlrLi8xgL9HpMB/DWxl4qiyXjQhrjbrQMlrK+FJK5mUXdJQRSo2oaAQ8tb7JqIifVMLU41lWaX27/xS50oU"
`endif