// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jz95SPX5Swaej6MuoA6El+k7o7dXFAW2q7IbmDs7ZQB9dQ190eRCEstOA5o5
PZhXBeI8ZY/qasxFYsFVZq1GOe8ccNgBbG/M5AduY7P4OOltlRHnrEfeZm+X
1CJuhXnhenUQaNb+bSVazufRnv5iznkuhzzsH9QrTSfB6LdEgYKcAJmPxbgQ
i6kSNH6IrwrcV1wXeU7h3zDWQ0dDdF2a83dqn1EJSLyuwtzqfBeJFUJdQ6G4
cO2psJY3eK5AhODweq064DtaapQDxUfAV91mBQCAKQ+R+YcvoGxuA0uRGWF9
fEYTkkxsslkj9acuaNYNy/uTlD1ro54gkdOeJMKC5A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ROV14VaeUvKmYQV/krEfBCmvphG9CP1ZX7VTw9/PXMk2AXPejsd1osdpz+P2
xpsaPKJIfQyvLn2IDwXOw0PV7RhTordcB/hQtqawXgUP4igESkO/LDqFt0Z7
POlh18u6b/msbyUciJtnkCOzi/oBanxU5zHCzR9lMzB6QDEQ74qv/pbjuYnf
a+077C8uM30HWmOwLA1Ma04ZA6jdeqcTxpZfn1QOL46vDy52mICBDJCobaes
tk9l1HGwz0GeYfc6H/OOEt5eYHitbsRDlvgguBfOOdA2fP5CCNsft8DdnsEz
BRXvlJEL55+jbHTCmz1OJ9+TPNQKoT/cDmjLIJ2qOw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aJqYGuBspufnSbNXKRZ/bWTerRUjSokfInJBku8znm3MzvtcWIo7fH8uUlMK
tfUt3BbZXp2FlDvPo4y7pYnMMeUS0ReZQw8GP2envF8NuGXhwX19egXAGE4q
HKp1aSmMJ7cAN1mBP0wwSIugAolAJgTCj+XeLpcXGWt8BvvnpE5dfNjCesKf
ncuOWSFGfqiRCa+EOa5jBq/xZO2yK8at5ktl4R+dlNvPbqGIThDfufpAyjDt
uGGmDLr35PyByIH6BU8yiqq5RHy8/qRWuCZi2A34W2RRGRaRPbXTokE6qkPr
oN+EUblxb2eWN7PHX4T3OEKGvP3jWNRSFVLFEvuVoQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
byPrrogYUXKVCLy8p68byjDU97yrP6/7DiJBipKlb58YdO6H1w8b9/jhXpEp
RX2F21uDvzWMPnebhj/9f/4hpNW6SSf1FI5xRY2mPCUhIdgB1ypIrktzOT3W
nan8xYyM9bA6UA5+1RNKwNbTb9U/MM+jQaf9uxzvzdQHAR9avMdsNy7dz+aY
NWvFyHhAbyg8prQFVsHN7Y2oRnl7TEFcButf4sAXb+vlp3Gjyx11M/3vvT21
FxuvL+OaqnSbJV1f5oxYYthTMNvsqjC36a8wQX248f1uYCeAn2BexrsnpXpj
B5LtzMSnfpZ8laTRQ88sy2Pkr7aJpy9ECI1pP6eycA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Px0j1G02YuWdI439YW+rsoD/D9DfgXAilrJAbZi+6AKal+hwIR3WUuEsc99a
I0ycw8Y59qpJfAAdwxdpAwoItek/UMBOCTa8eByrU/LxT/99uLav3DoWkWXw
5giRlKusRO1Bt6kvewcU6bnaasfgSilxI2RqgIvSmNQ61xkH6d0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oxeHnpSCu6dUGEM16hBg9DFnkWrIemDk1dE5RId7NuuzFRJnfoQOiMzB08cV
wwvHU8BsXj0ZjAY0jS0ZeQzUVfyTZxy5qvSG0NcIjN4xmDmwbpujhmq0tX++
ayIApotFT6KroQySoQyECSe2McNa53+2zyR+kvgmjKewPkrtn04cdKQubZzk
S2xiE3sqzJzfAhSHlDjRRVsUqrN6feDwI6Mx8LIQ7MlYkTiHlu17RHnWwJLs
Hrc9QvqO9+3QjzfnMVaOuBuJvMMRSJzWflaXMFpdYcOQqspC4K+HeRm+CI4+
SSdtv2x8ordtb6jHkZvJf/6yTMeqUkvW9o6FL2uhl9nxMTqSNzqWaFg01m3G
eNHXLGHWDTvU49eu/d1pQUHnVAOMRNvqDfSwN5O3LUrhEPGurHYNmprzd4Z9
wd+jQ76TM7adgGyzDxfpH5Eq5LQgIS4ad5T+yXsNAWeS8X6Hs7MMK4C9yBD8
vywngbXmIxZZ9KqE+9UdeOQD45YwuyYZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lLfQlhCjMGX2otR3p9CsXqBImPtbPGUUQOvKqSRHSIghC7+m5v6j9nlzQBy7
fcnLNbxEsnE3Le+bo7JZXYEBBfV8sI0SrwbbA8ik4GY0f4KRlEp719s2FSEj
oWVHGp+kEO+mNxW1AEqGgzwwOVTAB0Rb41aHPuz+qo6OXZ9YtIY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RyjxXjeiUte17YgiuULGScAz2El4KPhPaxAHFxO86GqpryF0qgqie9zkwmAQ
vHpbKG3F3RFxfgJgeDxendVuOiJFJ4JrBl6CIUHp6182CoxXXYfXtOTDK/LY
y5D6JAYkoyqj7l5mdyN+8hvC+D6SXkWUb43KhqtsmfBMViutGIs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14560)
`pragma protect data_block
qOq+Im2T89Covd+JAoQ6wv5IXfHYqwhyDSnd27VgYlyD2Wug9AmOIdJd/Kd/
72BIl1Cr+nGr5cILBUCykKq/bMVsFdUrjl0KzUppmHwAc7hfOT7Rmo2GH6JB
jEMhLh4hvI/iWRfekQuYJyXIcjGjQ/AmYnyd6EdwA2IqUJWrHSpxdt/H3SgI
3QfrjypQ5uppn2M3hvv1tlTNf4sjohsvOAP4Op6js1bKpKyCt2xCfZ+jKR5f
X4mmjZvq/L44JVflcFyCWKHbi8BFZiOZCBQyDb6cpBOUg2/ehWO5lcJg5IFe
aK6ck/RVvLY3fXryabI9ZjPLGyUnG86bBQbRLeCNAkD7SyJNy6cKHWaOPUfI
r/Lh1oTEor5s70C6KrRPeaJ2enEzYTQWLjb47Qck3OZqZltXmNCjd6H+uYH9
1uAsFoaEmCWCh31+qDSNpYysVmFN//KaFCbFrHPgoU9gYDelVZUeFo0o/gRB
hAbyVUjTXWoD/ZqDvqg/T8oo0xxgHANe/6XhPIIzc3lyS8/LI9SF/Ov+3Xxl
yzPtxNpZJgb6maCmaASZT6ZOUXfm3fs4IWmz9vZMjOMMiyXaMOrjlZyIfYPB
7BUiz8GHDsBbt0bQCvCN+fCTDK+tLKFFINw7IYCFz3YwUghdSr6SzFQn2LHi
fbeDgDxv7Vgl38JqyrkNf+uFVPv4bAvvpsecbF+7KGfrFrQtUlNuJSLPs7Tt
zlIIWfkiSV0ghOEtZ8F7fwKUGPR+NgobTZ1NHsf1qmzasR6Mz7w7hQY5zAN4
pCRYrZRelLdX7C2tGSEh2kChnx4WUpa3Uut2xpkR8outh25cA9PRMjU5mlqT
Ensb0eArERrFqlx4v4IjWyAUC1WjSTlif+ky50wORpYV5UsMiYB+vklUJ0EU
g1ydjxxc8uicFWix62A/Dm/aeB43WaqpisDRsQ09Q1gzF4RLxyPmr8ZTHmYA
NBRFu4A4NX1yc5BAwI8B26mvQV4PQ3J7ryGumPiCyOcHcmiL77bi+tdRNpLG
jg8gBJ3HIbGkNhUBXMaGxUUAZWp3/a5npHOpvjmoMqJtOhqBG6CSZRYnYFzT
/uzJsqtV4G8Ze+jeTIM7TC2msOZf9RWa8DXSON1sP7vGP7j80Q0SmrSeHN9M
IIK5pUb9P1NulvRJ91fADo3RRPvxhB0oMRZUKfTFk/jlqPOJRip8DxgJGU4Y
sRZM7Vvl/8xbGQsQC1MeCcm64Rz/MfeBLfbUsbayvbj9R2BicqippfDILeLP
9J4VUMY88i1VrKMtqAlQRahFlipUE3avWRXQ+QgOjsLEaRIhPjqBfVv2CQ/w
J3EKyR9GikpeyIqvQs9kONRq8HEtj5igFtzTMJwJUAMfrjb227GJ9c9PfVAL
8D0zwgvchGlYDxaNxHFUghf8BkSEsWl094pETsusXOs0LkBpcoKW5eH6cVzs
3bGQGn9ppXOeAiaFj0ssG+xPGu+5ObqXa6BPrvICtQataaMO2fwfKCRxQV9+
XEfTQkezdyj2MaA4CIl6Usn+I1YmpEb66Cu4qQnEQyKrdVsd/w9tshkdW47o
ziviKJxbPfwQtoLaAaoJ7t5L2xBntWARjUDQwLRYlNjP9H3lctktSrBSno3e
qHIibnxZeu+N9LD1hxysJcgDCTvCs/qnchUuj1f6Qgyi7H01zOwVVUozPwfA
fGxr1jjThDdoQA5tPuB904tbgOsNO1IJYkp2rJ+s7r2B5AM/l6I50sUpDeUL
PEwsBh4I4MMiFeeViHCxDtHkloV61+Y8orB89+fkFwbinVjC7pmvsHg3MqiD
ulhUTvBDinX/1iAGaIIp9vKBLOdGJB9Mev4WW7BXpiY0wa2cnmMabIbwUjQf
scN8LQOvfKS/bg5CZ77C2sfTCBnQzf8msgtCJS0XYdWCS6CePnzH52D58AvB
YZ83LF1sbBtrcPgtJmX2gZmsw3TGbr0aMS7MqOkCAXw2bdmn13WqhI+RBqt5
XAqH0GF7R/zIV9bA9la/d8J9V/GLCwjrhBEGoYCw7UYZ9eKuEZIVR4mm44Y1
cnmN5RYoA39JhmTvAYXG7AMZ53w16jmhUM38RflVvHknq/CyWGlOoJKoAYRT
fhCyvkIUg6R3oUmx6r42/zI61GqYzuaURf+gmidj5T52TeYPYXsgPAEWj3be
Lh6jPSwE5wkUXbIT0vSNQsf/nvMZztzfNxlrNNTG//vX0JrnLwCwPb+Us6aZ
yRiuSuDksCIQyYBmNcJrfz/wcUO8rTNVTe6plZ3I2S9AHq1DUKB7EoC8a8oG
GFyewR+izNaf6+vAD9nKl7jVIxAxEQOW6fC6jBMZpNuD5abtpJyhGWDiQKEG
j5ULFu9qy7Sc7B+oIZbm7ZZQUhU9oezo0PdWXm6PnYA4tMSHDJULTIGVUYDk
O6xAtReLjLZW6bNnZ9P8Eow/A1aZReILFaIbJebIXFNtUIHUIQELKq+MB5Hc
VwA1Arof3sySD5SXjkitEeEp1njxGBg3Z0hig5IfAluZom0SXHVhDqMxOKlk
lfQDycOohNfmSIhxmvBOGTQPwB8L9QSgq1LUxFURckUP9ZGrLFARk4WDEAdk
AtVAZxoxMemQQLszHpdiaaFkDjXmTaCbTh81O5fY5SAWWSEMEGekRFAe9jmg
IzjKNAomn9rOQHXe8eIccUray9Wae0usWU3VVqElTxhxcBEO8z5wjLR3vD99
FDPVw92LygvTsvXVGIIWj98GWX/xCBpAqLzEVJEJOpohgTjvv8H9eNTnzfpV
7ZhqKfr+ujAKN0W97MvKfLTXKjlA5hcstQR5JHLHmAtUue4TVDeLpL8+wWQj
gKlejQOjt4XBbm/kvED7bEN6yR6siSiyhjOwox6WBgjmdUHFG6/V1w5CmjLn
0x9QA4bJOPGKix8EILhwkqN09sHi15rfJzDYRB9rTf1VGRBBvlLdY1dWsdLC
bzQFDbDf0+wKZrr/FPO9KxwUkhT+tq77/jxntlwjPe7SgEdk5Zjhkjuiln3y
n4qqDk8ufozOoF3dDqG0NGSgR4unhTNilLGT33C88DjnFaYXEUkIaLYI4d3a
FrFvovNbKf2hBGB7DIuXIaq+UFBqnOesMZN9Xxwr6sb/zxMmkKyl+m0B8KAQ
EYPqmXItUdCYj9fTA0YYZhaK0kL+2lsPRHRgKL9zuZl9eW3t2I5z7MLVkVrj
YQL/WX9nmuhuZN0fYHVr/KrDjdwZdHZwxZ+ZT97IoZLx4lYPLYIQouUSOkrx
CD/pfqM3ls44YIiY8relp6VN5DgeMfmexKopHwnUuevKEqKzPmnZ59H7Ih7c
okf5LriJOqxW5H3wRQ/0lJbiqwthW4QUMV0NSS9HN4kacuY9rR5CJPX8W4/E
CCpMrS7umhKnzA10KdvqlVjC2tMkriu99hyGj0ySBOZ2i90HNVVNJZV9XfMk
/of0Fvt1Bfyol5BrVWSUcuCmdYX9Q6amYq+4cwAI1q0FIej8c0/0Jsurfiq7
XFHJzvcPqGvco+q9CF/NHnAlgOTUJq+5+4pF2HKrlCfdhQaYefjyaehdOCLA
NFXq3TAijnjuXVbNmmJSfdqO71gn4c+Z7r9r9QWppUybTXf7/d3FAeKMSfYG
YH9GYQ1W+RzqhZKyUAgk23VAPCGF1edIrHnNkGQqlmYAPjFjKo47ujA0AISi
SUo/qQwwMaRCUN9CBHH85Y3lPW7xNzUtA6BqF0g3O9b69hgZUfyv/EJaQ/jP
sPqS3jsOQyqNB7pkxrWtHyrAOgAAz+oZjcNeeAjJ6BhQqFxA+cIbDZu786Ik
KymKW1ZjSYgxW1Ycah2eWxst4j6N+HGADtZgwGYWBLHqiNG/cIMvOQRNwCUO
kEHKC+ld8RQN1OJoz7cnAaUEEYjurdX1J8CxmZzIoB3TiI0H9GuR5OS67SR0
TlwuoN45LhKjmY+28KfmlDQVEgjjU0AN50Ec2TmhWYiHLTb5lt1h22rFapHV
rUCAg+DxCu5eHXV4nxJVLEgHnUeoWfOAgEjmyd39dAiT1i7cKLk70/d+oZVO
FL3FyFI9b8BRHPwzIPRgGJm+d6ugcZcKQTirQALZ/wqdJvlKoHhMnbCaQthl
+TxncDVewmMAP4Y9RcNzzQje8u0kgo9CGGQbC6b2ufPrQcjp6wH6gckOEht/
hZafdyiA6k32tebOttHjRHxTzanD6C6ju364LE+IX84KUiZUiXhLo9i+uL4M
aukgTJA4+ufOla6cbMv1R03C+aVs7PWf0urkVnC6wIyRVNmrAb3j2vghrkdd
JkxA2GfmbbghkuBLKyX1hZnV9LlK2cHeJTmvDiBZCTV+86v9hA91xjQLVRYa
UaFtAWnG5UJnmr5Pdb/t8zUhmG5B/f66MuHZ0eKgHR8+eB+x4QRhNzGLsNrZ
/qE5JN3yZxmlmqZpVzUMo0uFgL8HRxlmjuyt3x2KDor9CvQ8KhWgRH/I1j11
FFwl4E3EZ3xDTZTS15nfMxQjFSBbfJ52+aaM+Daw9GfXxIQ6JyROpCloLl0v
0W459cjRaq7ZUpCpuhzX8qvVezwrlTddtUZ+ISPhxb4TfbP4IrM69M+fyyap
3JrJkKs3hDkRYtKP9PyxebyiSRPUhNYFw1S8C76ggHsI/ttSgf6pgvYlfIMr
pjeoKQverU3ZgQqN6xjTJg6MVyCjpAKwbzKK2ak6E1W/QaqqJo7nrUPPdjG/
nYqUvOT2NBJFXg3jOKWwu6XEedmtX6+e+dBU4S3Qg6NJgXQeiXHlS3xdXvyA
UuLJgwR32pjqKBq8wuidfnk8fz+PUNNEOEniOBe9AKMrMwtRkNtIWPwTpDFl
cmfJgtAgU3F/wobZGJTslfm5oDO4avx/V+I6Wlnys/0Pe8ovu8t1FCrmmCiC
twPG6ADOu5KIhh67xDpc2AIseinEW8jKlL1LMQaCRnket7kS3y9D9CvdKC2j
VM9RxLA4f0mlWmXITYnl0OQVDOh++wExdkuIs0Yl77nduUDXLpL76IDdnC2k
FNS6ggkqSg1avIyASQsiV1F+iWHUYr/CrnDRh5HwsUzLABoIW40/pk0o2IaI
mTnJrBB7fdRz2ptCsSk1D+nkzaIHTguSrrOYSKVmZcOjfpxQSbRxRIkPBXG0
BfS5HpBMvAGFeN15oK7hWOSAO4+SmTkKHdqP5ll+tA1zIXHNguN8gv6ij5I/
0z5JbZyJaRCcThIt0YVTd6OGINGaUlroKFzmOEbzO1nNQtIwM62gnFYo6XzA
+nr/GT79nqdJeZO6Npy3o5WPNluC7sPKlFdJ7+QjjybvR/0+3gZeXWxJhP9t
LMN2Qbq4zWj0fSOvSu5apPdEt4dNIHOKspnNhqx6C5pHeBR9kwdeJySML7jX
iuuWQq4Jp7B3knGoXaciy1TfKU4HO4frdfhAsSDupmS49YTs2y0/2BNLGLuw
jGb3cBYpoXdBlPeQnbGIAg/GtKYjrY5x6rirq82RtaYMUA63XtEm980Gb/Y1
I1n5AM7r7j7XSNsvaalsiYdnpQ6ba1mf/zGlkK46S7xTB9MMNcPQS/5rC+zn
cePiL8Mf8ACZq1oOYqRqcmXtDXSjroQIKYEDDJb6YJBhbKWEAoyDe8TvRIO0
R6cacpaTJhy/aZS5iezIJesGcb+I3BohO4V4RcEUPUMUjLgXfUX6v3hsH1Wb
ds56B95/zlylx1RvYDnzIxox5X9ZI49Gra/bpFLLDrcoiXnjp5yuCS5tnDZN
I+TrXrDWTSVBbezsAmP0EU/rLLq+uHBEXbY9PMO0nUJKXpVfVx3i4w9ujoTI
32KxRY+5t/BNOe8vPC8TvvqNbP/i7ykE6Oiw3BC+uzZOQ2q4IEZVxwCdlHvD
ggk2Ph/WjxuMH5rd1MVo/Fy5Qc2ZlIDR7Mbc9CV+LvzodZumhbhsy8vtJynl
MZpFTp1ubFxfwnPhojVxTMUEW8X516zYeS10BTAXsocex6W+9fomyYrxg06w
MqycRoN3S5mH9aS8zXKd7bnMSW14b3akN73/ZbehJkfkmfV/grnxfPeoQfFg
lpFG3iSRnPglo7Ui2B3A1hjFaCACj++GXB5cJExDn9O5cGUT5XY4FOHkR4Rr
KQ754QGODAxOfo3Mz8wS8SOgKnRsfeZMoclmb9kcMDhie4a0FKwiiNyjyIXO
MTlX475USHIESzqjY+unLtWaihI1F3WOARNKkC5SFzsn7OBbRFKKt4e7IDzN
kPBMFyikiidyP/0iqBWBvCRh3f17HW5iJQErf5kxy1Injr0Jc8/Iu9//gzTw
IlH3XkzsF9NUx66ekhNLyLF+ca3ibk2TCYdgHwymX/KqzzCbk2ycUlWDhDOn
atK7qlkA8m0QmA2iyXQhOa73VCRPUeEVL9k2gdeWQNd4kPQVgeZ3bd03yK/U
vqre5VDQMlkQslN2ZZOFZ0Frbe440DPY7PxV5oQWlCvzTI/gOVDn5EHkUpr/
uijOrKJwF9M7Z7xgh8u2RdfqhWWhSx8rxpZJZoknHeqSu0f/7XjByMtlLHSN
IkdEvKt77jYGz5TTf8966cltKcxFYg29oqQC4yD23x/Bw8qg3hNbzuXbU7eS
aklBNVn4x0Ya7VFOZDo5uPd4QyrBfgZElTlHGuUpml7ddFFpxyuv3LSbOlFh
JR65CUpNZz2ffccYQoDoVQr60+E9KIcH/Qiem7xw3ohshlSjkBH56L496tvA
L4y2cfIbn8JOoB7JxxV0noQlQRjwX1IAmSGS4y/6C5LTmWto/6rsf9P9aeDH
vIv5GUbJWJl2AFKRaNgG+SFV81LiWD96R9Co2/lz5okR4sWoJyxp9DOTjGAp
RJtaT5dCLLWN8BVdjfNyc7PoRsC9bT+W9NphaAu5jzNOCYH1TUAKpeFt8C+S
hh8n4pjDgrMT3AAFr966jK0+DqIqSFTYNVr6xz6BfzMP5Xi7walwq7wOI1a5
BVqJFSwteNsRa2erkmZVD7RAUMxptxE6lVSDMXi5YYT+mC3d6HjFYknkuHzx
E5+B+E+nQXCUQ7zG6DaFk50xLfmZUFyY1XPgSsjKqb6BI1REbP5LYyjn7K2B
bARYs2nuYFm1kvs5QnGONMGVcS98UuJE9y7OP75mqpwhSLWSHwX+2fJrcsRb
wfE71gbNYony00rRUceSByLwRcXSiNzX9h8W7MovC/CtK7VxESXQPfEGmHCL
4qJpHo4pmUVYs6tDw/dm8AvN4ZngcZtetf4T23Sq6ODdvT7vj3gk34nGUqSZ
401j3GeHFZawkyn5ZnDIzbpPdjK6gFbS9aemCcXXSorRjjYt9AR+H7xUuTDD
t/UV8/WtWyodpkyf1HQjO9Klf4/ZV/wNeDrLHrT5mbh60wY92MbtyFzl3VBD
0/MLa2wgpb65f/3ugyG8Hh0WaxCVYKMP2/IGP+iCtP1nDvKPLGV1aIns+YKW
81eghLkQuVljpUZqqMilZ1r9ZTKqkMbxoWk+0ccGR8dZbmGVUIW9MjEeHfxj
PRYiP/u0SmirH0L+mSSzpwy7+TY8KQdY4xQ1xxoo+8OeXxDkV8QExtKe5iuP
ZnaRV20ikebs8ZUMs3WIpexTkhVIvIY2qmbZ5R2fSO0rnn4AQdMczU2rZ99R
8hIR25jaaCjnX9zHIPfEueStzQATKbUk3Knu9P++YPuHbamPPWPaRLAPfCLr
lPARxacud3/kl+9UfPlsrUiNkwS5rxG2gxpOM1H3qWLlT1+r22FwsT3rUvkJ
LhX9AIFJsp2xYxCv4AJsaGhYaCo2+BviTH52S8lLi6VE0UTBRl1b5NKgW7Ao
Lqde7AcUv5+tRs/xIJyXT6jEWhM2wZznJKdfkW+Yt8Hal2OOIN4i9loQOqVf
oBQ2MqMyZ+ppbfsZSwBFJaE10Qv71KnJJ3CqWmKJzeDVUBanlzFM8qH2K1rb
SIE+lOkSuGAWJoGKdRlpQz1iOBECdOLPxZzsy+eVubf0ZBFzbehcOvyLB4RX
fF4iMdiQNRCqv21rhpflNK/KwomjN61DZRvEuGfwICL2YHkX0TE0G3mYVKj9
18JdqiSUJM5j0tSb5W++dekk0zJux6zHiOH5h+VMYSt1Xe4UVqSQ8KzPvGrd
SYITpxKVWNc+KPtve6NyXBjf+2nl0NMyJz/rTIAQds9DK9U+2W3jCQnmOaTY
NKe38NE5jrdHyLwN/navtwycSQL6+LihAq/kol3PScIE+01lpGm1tOzQOa0a
3551JitWmAZ0ZbxIGV9rUzQqjKghlKdWg0AC7BX0p86XMII58r8L/HPGlVT3
5a7GGqdmUeVy4JUiaBVffsDuBBiLsOuSp+XZ1IrSkuXVW29Abz0h4jqNa9fo
EJyAK7sFk8ayGdu1wsTcYPXzJYW82WvqdXr7mzXFhAuzhkUzcqrIbS+HgbBP
d+UC66AQbYYrIHi/wxML4HwoLVOaBBGuGbDbmKoaT1cbDg7N1db6YSPOp8MG
PEzEMveS8EArPGcUBftgr1OEZtrE0uNj+oMxqTVsUBMehQ19k8g1+nSDDjIN
TcaEdN9Clb4aZ0gc14TevLKvTX41jm/QT6YwaUR5VeAMQHRDJsNceVo0PEb/
Iog3hvuDkPojNsMtF6sHUGB7NFqf6vs+nsDl1gd2LcRW6Vq+fMwfdToXYlCj
suI9vvc042xD9yz40SiVWPBqQC3J/pUZ99KUJM6Z2s16C3jweDCFxdYfZ/B5
ZE7EYl5eaGBBDQyJXzTjCiG0Fn3JKw0K8f/YG64ZH8ZgdHQah9NU8MqhXfi0
bwe6l+aldeqD0NlSCEZxS1ao4x9o2hGjmLz2ht7DyPDo5Jo0qE6/ZGunR00O
HZSmTgofPBUXxyI7S44Stce/WZjfVOfSrN+UFKoo+ou+deAuJuVbs1nPjbej
MPz4LjgCSY02xizvEGXZDs3XUxabEWCCjKCoZ2+7qpUpQaIGOZdue460NjaC
VvdqP6IWdGAfNMa/9GugkTP3oPdOcsG5+YiLbCiaqe/44+fK6W032NRjng+C
Q+6f0pvfpskKUMBOaxL6Z8p9oW59Lz7I4LaTBNRy5VtBaBweNoF1qmXdimE8
gFBNT6h27t6K5gPcXTPRWVSWRWnfAWJkj8VYD+0gEdYy6sTGMPFzxeeyo0Cf
hOyRzyDyrfcNdV4Am+ss+AYTzYWw1WcZrjmZU85iGr6s1t2nJURQXFligEo6
bMzAkR+cbyqEsmYU1Uc3rle+/VgCKh2sZapFsLhfETb76bIpzJcxEShFEwTc
NJC4yi1n++keytsyNFkOQwSXe3WBW73hMgk4zzQ5wPgs+QRrkaGYcT6YK2Cw
jCZRrOYe4omNTCfJNY9sdMq93m9AloRjTIJJ1p/guSswuZYaN7LhK+28N5+4
OYSqmo7MNi8MJbjonJyOciSdgydREw5a/FVSdUrscup7R6NQz2YFbHtdzm0J
Dvlju/Ybk6knEMirumXNihIQVUHJ5qFySSN97p/a0D5hBxK+B+dWhQWv1Ria
Ns0Aw98NmBsta9AKrYfp9lwSse2Or8h+k0cDMKco4lYM9ibsV1YKoX7NCaJ4
0xLpgxOgHJtSSpaqN9QcP8apEEOegcJGQGfdco2mrBgeUoZyV/GxaZtGz7Il
u6y8/DJj6tgt12ucnpPpWcH22MIxE7MuKCGcMAe5oCMz5aWG8BW0Co5nmMS6
x4cnPQA3FjBlp81tPnf9C8QRoK6f49Xc2PlwQAcxeKM/6BQU5kYCCld8dkZC
Fo28gmY8YFeK/8GDyaNWpq/okbrSyKNj6thDLNl5EKXs+jGH5vtcUakbZcwo
Q7C3rHIzt3aYOXGAbwe4qVN0/BOBxe2fJU9eyNum2M+jjm+IsmxweckZk6on
K0brOgqTvRM9qmJ2h9Tj7JsVM9MkWUPgmmHXly3Zk1avqMRVWkiVEwCoo88i
9iFpVfVETXGoaHn5O6cnO89alFycb4V1jNXKQaX++c+cMD6S8oQJQY9OzMzT
BSc+CzJMlZgVizS7K1nZNoO4BH1Yq/gSHojn6VHP68WmfkW51mpYxkU7SR3a
rZ1szMYOhrLIhGfmRVVl+ei/kU2U//jlQyNyKSSF+ZClXVNRbwsGw9fNnL1w
D+rhGCjLu9JwbO1DbaI8hK/NumT9RZb3+7lxeOaVtyzVBjIe6nl5F/SJtbrM
WvkDRq7ZciYzOea5Xu4kv88CR4CfrB33LtbthS1J+uI40zx2prxwMbol3KXJ
gscN9Zbg+sTQCqNFtWmrz14R6iaJZAkRYmoi3uGe9itTuF5BJtBWa/otcoUu
fgXWRpyX2YTRciKraTY+ao0SkRQkSIFQyW056/ew/0PYLfAlyUj92r0B4F3K
V4r4Jk/PHUmsypNx9czL3u1QoPS5a8YTEqwV+T4s2s+jMc1YCK6TP9BKYVbm
S3lcUy3/pQ/o7mLKDKozmaHoF0X3EyXpYVCLY/F+bgeId1OjLpxdUBy3hSKK
aNloqojWN3UQhQXW52WkDx2qxC8Thozm+c1SulnzIkqrh0SRAFhsRRFptdNS
/RmNHBfZwSpG4y+i6UkupzzmhO2EUnmNEKQKjcw23quZRBZH/5WU/qFVVLjU
HgnRJeW46shXHTwCk2frAA6UjZ9EoFMWFD2XkQnXg9nFOT187Jn2GyQvquTK
8byczQQpSl+/2MbJCWScP4yRM5P+9Pvk/iBFy1tsF312MZKGlF/FyLiTPiEQ
XFHPdBGd9Ysxtho/nC+UEQR2oE5xEE7S0j2HMj58W8kH8qKf1tTMLsqUV3J+
lWZzeGPlXFfUT/59Ma6HVtg9xQm2Syo8lCpGFVldIFYBRjSNeqsY6S+D6tsv
54w0h+caOAQD9AUoE6pSZvsQ0J+6EcVvkdHDDHkn0Z7zdfPYTR7wuJDvlUe/
R5MdN7TXwNZQiSiX8ARACHef5aS87NlI24g+W1DUt30WcYxW8VZMUELGE7Bm
6Yl5f9WbHwyCtUCobop6haob0gY+b7Z7q/ab3fKZ4ZUXSrBaC5MLhS6diPnd
JNe9SCgTbcHJbBRwnVhn3FmiGhU3aDfXDhA1PHjIEl4bozoziFxe28Tb3oRG
+VXbTwbhcpvKOeG954WvSKUwuDeVptuK0XeN9ZUr+N+tYsOatoGvoL4PyYjT
u+e3CsDZqYPPVTF48vpcBZO8lRT8WFheIIRQFVKOAJ1MjhbmEGt3KMmSAGGb
TNbX6tpWwzl16okHu5uPBvR+sSETxLupLw/uu4tcug0w9SX5GXWlh9lA4gdy
E7GChoSd4mjHPAA8sR47oHwc52R5gmHrHHrgkr02ox3vQipHaxlKz9OTr5Qb
kPx+ZyM7x5bo9Hpkp4imH+f+roViAR5VqAWe0YEp3xkap0z8B7/UGThhRsHP
ub7ZiqlraZhBWffQ9h+2+Teyw3FSPdfjS/bgwjD5bwWSZ/U4JEcihfh9A2Ed
ANLbuc0x2aWWtbo4eXayqv74hwbZnXjpcE2XZ+lLLN8ZPyj335iX7R2CQ11a
F+VwK9H1DzU0eB05mnH8GQ+I6wJ9obVVn8gbZU65FburqQv7KpT6kxoZz97A
ucUgVrXU4frE64Ow6tfc9JHOa40RbYqbcmzY9n2y1qWJL9yKZb8RvkcGuU6u
ycbnALAAXUhZISKhyxNU2Bgnqoc3MOHoVxrqeXknLE4n85IQkAqS5Gwg7mKm
hx5hOjKBQaQrbu+Hin8WS7ZIyMVpn06/R9IPQOIg6CK2ZOdoTk6AcgcTEHG+
E6xPE8TpAHhA5phT1WGVlfGDM5S0vWKTR2Fbv4BiYOrmSHQGDbhrbX5JB0JR
SMNILqQoHU/i9Rq67o96EStxb5orURkLVKEbC7VRFH/AGuw5ypL42O7Xijny
43Qo49/zqxAMgm/RGnyzStcOaYh2NoBEQA8GqBbQwVGnaXW5jXenjQHMwATZ
XN7Kxstot462JMzTrYiD+dq4xacE/0ClDJ+vFxdwY6dC67bqJ1cycy9/AjB8
Bs4RgBAdS4peJVS+EC1lmN6eaLC2h/zNIdR0RUAbyMSBwp+rdNBs5Pwtio8Z
2ik43WeljjGTxd2VjwI7y5GiWLP5+9Kb6EWClOun6i7UAQdmOv4ckZoy1sfo
aHWP7q6RguylXz+iasA62GUS60+OxnBv/mF0CrYWsLAmvf5gRkWJWjLvOHo4
pRYKemrmCZsoyUDIg1rBcSLINeEn9nM4eRyvvdTvpLraVGrz2uVhA7nbQUdU
5cSDLpBcqZHJ+yV47wrqs+aeCQHwm6Mx+FRS570x39OcPQZt9P1tVWjMXdkU
gZZKOSmqKcnxiIJ4QLK5OQhTacLjS+DQ018xAM7oqWSVVCujwoqlp3qJ5dF5
FIBG1K0tEcjLsoJjECvSgC9FG+BnZuxaHvtNS1qxjtghZ96uxi3QEGsf1wcP
Y6cnjO8J7WShoH5BuF4wqmx9sgUIgRNXOg76ainxE1WkokvnQM5+qG4Sf240
sD8SaoGp8r/Zi0NUhMU2jrdKGvq4FCX16mxHHYI7GRC0dk7DQCrCW0dKqqIZ
F8v90Aybq6G28e5iIVXVjWeCE9iCEBVJl8xMDbN5OypylJSz2MaxmpAthk8P
EOocv9/srqLJIYxa1zZYgscoOvsoG21LquUEBRupouDHuefnMde26CMLn+Xn
fbKnaBeELzp8SL8VW4f47/s8q0q2pVLdeJOaJ1jCLPh0F9naRjB2+VHWn4dQ
kM7Q2VwZC+7yT3mltdGI4YvCn+K7AL3P8OW13NJ0/50i3T3OSv9I5xemIIet
nLI7RwjJm67N3y5bGFo7lhmTWOxR9+QLv6YZlcCKBsRRN9RIo1q3BsGUV0zB
rjxU+KZmF/5nW+OPkEFJJiAVPEgt7E4GcxtBzzACefuAYEpCW/5jaF+LxW4W
tccs2FLC9jfoWysyz4vv7IuYCmj6OR4HF/IU0F0LW+nucIUXTLoQwfALxMPP
zCCnGGNG8YTFu4Hbzff5aOLFqif2MuEuVsxEs787Gi83jfZWTY+Wd/sPff/x
oYQozZGSy6SAL8WY93JllGbNytU5JXhT5XAYQP5lo5NiQXkoknfE8mFhbgoF
8tIvefyttJY2u+VB4cgBvzink+uaN5vI+p4LRhA2/Q6w1nmUuZBJ41UBQFWp
MNty9Wi+7xSfwMqkRDC+hS/cqEDJWZT4YEPseYyJQVFfn17TZONEnMQKiiqq
q50KysvYaqX89D60zzNoo0qnZe/e1drwcIUMqjdJb+6Juuar6xdlG6DwbQok
Y2dGXx2ye6NU5/RMeu8yRwe2jCyX29NRqI4cvJ52PDfMUMwfQ7BL9GiUpgBa
fUsxkBauhpIXCaQRXjytigN+cG88OcdeOqHJ8lml7A3AuiLhzm52DY69dO5V
PrVG9gOa8JlZQddoy3r91zIQeJPE7yIJe+7tTN4/a+TyTgTObIQoamou7JBd
8EPsmo/R7efqanD/S3cW4x+PnMhCcxtksIyY2mvH/TwWUlGI9I5TZjoBlbcW
RrBDKHhipYuglQJh9BJuMbdL6jDTkigxz4ArpnLaPZF3EUk2Gd4EcgjZ9fwp
T7SmEq5+MI+QbMPQBDw99JYKFRb8yJJHVKEh02sM5Dhb60UQDlQ1hu1T1PYG
bMHqNyh92vGa5pKaSdW+pQY0Zun1IiyGm1k5fzVO8QyuahkaH/uT+nUXg/q4
AQQmrsecrWFZMJ6OH9YV9YJ2Xuq/jQ2acBivKrEHO3UpNYdC+rz1M27G1Qgv
wcSokxkT+92veJlgsEtWL9D0M1jAldeuuHxwuJiVZ/vtlFFYU8RYZ4/POyj/
9POJYy5ZshHe7ti/8t/TXmWfCbu8EjJht0HlDX8cx1IZBuVYZolHd8MwBZ1J
NpaFNqwAbGOrCphOvwpDYfNJ+3MZ6Br3hu3S5lzTgwLZn9Zu+PfHGiLqtWaf
vk36wm7+BHLIPvJ0msOz3C/ROPlLRXBl0uM3lWzZxh+COw220iEMsMZB6Tiq
QMh6gIVYH/NqxyapeahkX5Ic/wSPlRpdcHtzo7W+be7MK1+Slt0AvQ6HqjE6
WF4rgW7kyrezrzUbKEGa4ZXmlyysrVRYfn7y5Q1/+A20m17gCnmlgYZdpy45
Z1UEfFTI+ViezgDArrjSehen6RquMA7/YXr/tL9Oghi6HZMdVjMJps2cO2Xg
3SyihxejrZGq3sd/5KlUrnHIWph4H50Vl5ZGhWUhyPgUwmgweY//dJZWRFix
OrDFcQWJrtdJvWNfo5jvQCBtcow9YvKspG8utUUSjZo7dbTeDQ1V9+kyk2DU
K+mIXtf411C5++Uz714FgGYNeeKJrtI/TBvq1bBFUhWPSvmYhIDZNE5ppzd/
DwRFdY2W4DkA2T4ph4GTVyqMZAJualnpMA5zZepMV/JAPQ2fgYThYzGGA5DM
ygF2gX/eoRWQ4aax3nErWrNWiREXTVxEhJM66vXsVYwtZpzbnKYnN6w/vkes
MIB9iGJGhc//DY5PUqAgva/EyZwO7vGFvpwRAcsSh06Rm3H3/BfI8vhe8pWk
FNRo+2W6OWG81oj3VYQbSwZUAfKesQd2hMx6ZctFxQ0v9z4efM/95ISmdapj
mu8eM3bX3dGVZdOw5AdGey+GWde1yV/kHuPm2iUjETjXssiTTdUIkMZFRINO
oAXNNRSzh217lKTPM84F/JSmkmFQt4ZAjSzKNoA65x3aYNnaYAq6L01LhjsI
AjhkQaonAEVwYK0FOisv5yjZlVTtQ1uXvcSrKI908T58wfnfZUxUnRCoYHfz
oVdeVHOhFCnZt06Y8wyfTwl1nc85qU7kkfGzLsXEEgC5HCXUxoRXrSxEmw19
VIjkrBxg7D8n4iCgaYmnNj2MwtfXMScxvB5ZX598jIa3v7Lj+XsKh2nXZqGR
HkKReP9v/xIgn2exa7wiHhGv2P8GY5qp6ag9arSVbodPXy7LMPVKIhdUx39b
ZUAG89OyUbnMlwmkKsP+srjiX8c2C4eVE3SCzgyRSqbiQPMjDcbW6hXAm0MK
e2COJfFdIbXWW1p3F79wfLfiO7Og8cN6y14znF5azQhZHSgx8u/4e6CDUfni
jC/qRgrfw0Ddc73d/CK0MjhWG6y7xuR6uxp6itdi47lJ6e1a6ASyFjElHzT7
A0O2nQNxBOZrolUygfTZMo+KdccyZDK9UF6doP5WEEEibsTxx4yCY49J9kBs
rcvhVm6BCRwjYUAQ8d9N2j5qeNcT/fhuqd4VV8r6emPUJU2+5Yr/vZBAl1GA
0+7ss3uSBatMphlADjyoS9NzpgpgS9iDPK0tNR4n091jr0sYa+Y0lONdpX7d
eJD0nNqlba3RFqYdS0Y4qdCczLvbEB2GDH79nxQmNpfrYkLCEkSq5qdekYHK
ZeDi5OvFIuBgICRxOdK/C8qOCcUerTvBxbD2yJt6QKiSVXCTGR+PsKBkS0t3
UtTX6xkR0S6baW61S7fk6XlDz3N4ayRYlpTDIBi0lfoogSUasI/FOrC3JxYL
nucMivSMFLD0B1KCEiFGtdmglBfnOP6wA8T6jLyHYAO+pvjxaY1AuB3C6Tcd
KY77cX9jMY7qS9E8vET1YHyrFHy+6yLeLJqeUUzrv2CvMt9RY2aJGe9AYtxu
/SNo9DsLmdi3hdDfsq64z6A8BBO+FK3/S2ltEjp3ptGfjelgmI6l+h4f8dsJ
XAygOs+L7ARTe5sK0caWxqoEcjSh7AcsfAzciH3+lEwPWgDJcZOZjLr9QQ2m
pBEo649s6IYc/+meE/m7V3pvMI5jeWwtyxO6n4YTszbKf0t09uGuaWNoFEFB
doQ/0xbOJousvVsLGZriWVFON02qFkYiMvO5w3hPVEErA/5DE9aOL4qq+lvk
ytdBvR7PRot0TkcP/fGeg2poa1wL0fgPPDafTVB2G+hoPy1wj2r4EKOpyxUf
W/86QYvny4I1UaDxNZfKg1lKXyq56iARwo0QnHYR6oZJWjh2DQRy5q/qy5Ju
dDJXyH1aS7XxhzJ2JNTBp/+u98xyPfZlA4Rft9G+l3JMuQQj7Y84r0VWW2C9
Oa6uUW7SJb768PRvv3KZKzx2P1nIqTEahL/yO+1NIs5TF+FQ3cil4RAB9e2M
IYXV82VTNqDX0uhRiZlvzzuTAsdnemQhJ/3TYd62qNHOoQH/EhqgVygBZG4x
gIMjJJU55g0haljjiuHphvAfzz5q6vfcVR3CbJGD9AnnvFhr1tylz3zJK01r
lybda/uDFbt0WR66lGqRbdPHIUNIhSWy6Xzc15F3uHiKDOpgWRqbo2H+YWZg
AkxfbaOwQoCUaoXfiBRrugtStHU3qQZi/eiUmOxMlG3hq43EnmJmnqTosKY0
LpsmkQOEJ9/KIdNq9OjVG75W2FGJAcu4QFhtPbGFRTXLjZ4z4ZH9FnJrbp1x
RIs7V9VDZcxPpHEUiPO18LG9yFMYM19cu2x9fq8AWw3E4Chd0zaEfBtQJ8Db
n2a9p4n/TZ5aWO06zjEZUpQuSC/cKXNsQ0CIpriyYSWy4NcueS67G3UICLns
NTZ71r5cwFAcvmMflPQ5Ru8daePAE7lmW0Ys/pCRuq6D1XBNZiAtyIssCP1p
7uQR+yROlaoMvccN00XvVbd7e0YeSJfO8SGm/TOdlIpFNt7Vy/wfYvtN5q99
4tQNnaXTDKX3N3HiwIoiu5yRhTXAItgym+SxAdbkHksaYCVhAm5WCy4scLgd
EG+gJRZOt5Ndq3BS1y7UwtA09HPYrRATSPtG3UE/Wh+ovScSv6BcSBmQJpzG
tuRoZXWWiaybbWSWEowhZ/A4W9rWndQvHrruNJDSbc+J47RnZM7Je3L9Ae8O
TkCX1fF2m9eOA/Thfvu72TGWbsNKuoTODn/eIX2hVRqJyMd5na1a3Abhlje8
IbaLgui+YUj2UDHl8/7rjykP/Ijrm02z61+ruFMGd7ufmz58HAvnMxgLIAi6
n9kcJwftNApQrFzMBsHWzQsLRxdjITO1z6BoSmXmiAIsXn/82tZxi3ExtxZ0
PEfnUWQ54mbDixCwt3nzyqSZdRrWGuxZ95Yb9NQiRTcQFac0o8RogC7J4Xhd
Uy67pVjDQxl6wNeg0W+moKG8OXD9CIFkY3UXeMVWHMX0xrhy7xxLNSN6sK+A
scn6tYvBWkluZaNBfHI2aTukgwC3MGAknh7pcDi3z5jOMUii9ivVtNNmXYdq
DrU8191WYiFU6iWCj4eTi7nvBocvRN8q8LPemEhbfoT9pN3SW9HHH3pRT2Pi
grmrRcrEBbrjIMMNAVedTXqfhzfrzozUJKpnxlBp7yi4huTy33t/cDl0u78r
vRwTQo9C+kIpVqn7rUKVlh3+uShKV7v8WYz1sj5ZcHMeqjD1vstXMYWGmAd9
Ax7Hm3BqDkE5/b8U0NHtl3tSTSuNvBCRMl5YPcEWzNtP1EgGMJm0Qgtaw8jm
MC6ZseNlLAJ9jqboamz5CL6BBjhz2viynx7bKRN2zjdnmqV6Jexfv3mvztsL
2Dg+WF/Cixig0buS+Y8hiJrokBdL41nXAFalveaNi8Na3etJUJpyMDcntcoi
GOk9TkrxavzxRrbe8c+Y4olpwvD3/OKumkK7G6l0TBujsk2yxwrPJMMnHP2e
O8dItMmGY0vdCQSO5NerD1j0rHMpq6h3LMtWHhMF9aeSqDqZ+hyvn3/3EmW+
KZt0ZPlraLVik26zqLLQIE3tZeNR2DmwDSY5rhAH1achOwiH9pSHzFv93bS2
2KkrXhfM8OETWmpkwJ/NuXrGzXGzylwH3YYGtjcv48oYfuveZK853DVB3pfh
oUYmegtWE1lLHjE2zmVs+jbms7gNfM8Nh4IS9BFvwbAfDNjf8xavLVR1JEjk
MdCEq357L3jJDBzdRl2HbNnMVnNOBtpUuJ7WaR14Oj0UxYTcx3IegEkgkn+L
DSIkf3feZYbbN/smyrsez7Ul6zLCqSeTgEs8IxwHAp19d20VFEqlCaGtFtiu
85eAIb9KoInH9pHNDZ3KApzVefEIp7F8D87NthKIW/HP4VfQGsS2aGssxBg9
i8dEvXpbHY5BguNsxmntf5zoSCw43R2L2lpxFvlR2a+eKDbvBkKDHbqfo38h
/0cYGR1wm46lbElMcmFguD0krjuC1IEL7mSeJ7fFl1D4VE++hUdRH04P+tYe
0l+GTMCBhc/Zur3PEjXc4AWWpx71txUa1a1GPXWt+XOx2v0abE007oHR/6Mt
u9KufqBnUEW0iA5hIqUsC/UcRk04dz4OBuiLXxNUwWuEnCXfnrn6SsVtzaob
Qps152HbRYAmNCfFLo/ZpWOLtlGxjyV3JmfZIN9BK4ZBaRRtLApVFHLrDQNd
GPhQmdS8UxvOc64TKYt5FXE0uonR4/JD/HS7lxbzT9Y3AtMt/JgSyi2OHa2D
WQ7d33C9+sFgjPQYdyp0rCXnyVfE5NSDlT5vyP6N0lhFx3cwc/qOqzF1EbL+
iFTkULsQFXheWz/SxDsumJkd6DcNtZxsjxb+sHWNc0PYKZqEToloAfPW+Xug
wS5Z2CF670x0XX+AUBa99Hh8TAoyl8FM0xV1HU2aSOGwPjj/nC/PDCKsxEVb
rv8SF9H4rhlNDVZdUvHf//R+ed4+qVF5YNWhAbtGH1d3cWLe7oggG6pTORV/
FzSi9dvH+w60aVG0P4NT3TmRSu/tI/EgrlxDlqNWxEjwIRseguZYHeUqmesq
Fxut1TYVgx1xkrwDRekJf37gsHeo2M0K5Iw9sM2X+ItoZLCfRxy9EhENeiq3
/GfrXrecmzoWcdl2RCf2wsXp8dNxR+/Lj02lxKFYrLMsEUv4KQEdHn8kF/l1
5OpjJxtLVHHCfmOKXM/nYrkhy1r81G3CdKJHaBlgsCcCp7W0+pZQuBXTQ91t
O0j/sTDidnSoMg0yxQKykox7eDuvQIVxTBdb8X89d9QRYRB0C0Fyg90yoPK/
SGYziEECrLM1p6M06zkPxD6mm34HhkkyLmdxOvhkpZ/nVfAcwNPi1C31ozam
CD7JBmuM9Vbw/+XPoF3hGcVwrKkL0b2FzCxQmA27jnKjjkpbMFoWu9Qg0liA
APS38A94ZXzmTaE4T6UnSGMcQHK936nzTz7oZQk8JmOiG/5szUitx0mPt+JX
LJom/EqKS0hnQuk4Z5UEYBKvQotVJSJjt02bKbuGc2xrFoH3QUkVU5hR/nW+
zhLeRgR3/MIEuctsI/tXAFr3JM5Fhx4X1Sj79Dt17zmzG8Fi9JrrRlqWbOhf
HgvPYJkrGtwTRoq02xX3t1tuazUrU8eKmpDfyuBJM4UNXItBskC+FbkSHQg9
ePzw5sChVWd4poRWVpoG+V5vPUG7jJGsar6yp72Lf0iT5qBTSyQTA1VmI0wx
9XA9LcrcuRNAy6tSO4PBn/r1f2WSXhFUHX56LkAkFvEIuKlY2CyTgwh5DODv
9DABNl8QzO+VFv1RvaCDHdGnFB+HoIv/obSOQK/l+Ov334v7QSjFobKlRWCD
+jG4dpoNPK7PkUsCIcsIaDEBJbei6fca9XcKsIq707IRZsjNalCf4XpTTmdV
eec1qiUicW8V0fvFwXJvY8NL9znTdzo3+Q==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KCm5s+SfdFrNc/xArBCfyIxaP+fTrsnglbzc1CNd/Uq2SpLHZJcVTah5S/3WO2NUeguT/PqyLSPS0MbE8TbEDWsAgeULxiHFHYJ591oYy1umMSAWUDOBFPSYt6NllSM0WW6GrzTWOHz/g/4+xRA7a+nIRaT77l5TTojORFMUvjNz8nlt+Z6TARez14YyQft8AN5LpKbZpMbSEpnvk/o1JOh36HsqRbniSIXoHPARJ3/hld1E3JyTHA73YyApv4nT+8Al1NtQBJ4ohqmdg/95VaIbZjLSekKwu50zroFWvmWB88STVZQURQ96f6QOkYi++97RqpbJDlUqzgfo+mH68rpO70OljCC5YbJOlBD/vKQVkX9eIbaiXzhJijhc8+Fmhy8Gute5tiWCvNfZW4JPFuRmmhMld1/iwzXZBUG8Ab/MMBcdzVWvR2xAbLzZuWc4PdS9wgFapv138MWm9FGvYZLl+KvRttREqrvvx7RrXqsghUbAF8mpV/sSRQ5q5AZJnAp+FzQtIZ1b+xYoc0a+gzvIS1TzYBWvZnsh+BSMMl0a2zYCullxjLC5262ruISL168XKU4j7HigBWA3knDaZUA5JeI+UokRZ80tWNPJDQLP6uASagNsH3kT1hsaDEgqQw4fc6ZApVblvwB1cjpzR0BGqRceXtak65qBogE1oJwrfXPUHOn397UOb8vmzfG1/TGvkmwlEe3FwzF3YKj8TOCHdkQ/ePRMvCUNxqqjv4J7Mvq4uvfS+vVP6qYO3giejehNGstt631N8nG9wWWBKQ"
`endif