// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FZh/fqIjqgveaRa0IjVnGkg1aBxASHvlpjESXj9cFVsJ9kAsHlcDtOp4D/cG
Ga/W0n6O3cUf/0knCtfp3V2r0LrRqkj7vNILRK+MF0ap1V571+AyxiRh3NV+
LCT8BtdsykU/3A7i4PWHoFlwPmDTmIVEU9p1Rx6POuO9ZY1IPwH2N8uFvssI
DBY4wYzblliwDfkw7708g71Lczm+aTzfk3xzYe6yPrHiKzlGpZvF+qbobrgY
UGSHdZUcj5QpZ0HS7icnXgKNog43YwcOpRgSTC0XrJxFi8/H0NQuLdkKhmHb
a0iE1cJSNZ3eBoPngWTQGMHkVIa0gWyZzMeeRpSZcg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lhyF85Anl8JEFmpGTiMwBnrsMhZ2KxFUYt3kuPRISVCxXC7cHZKNJrqLzEll
merZqczr83zfqWP4zIEmPVodGqjWbZXQfnwYOYvygIy4pLEZkHpOm4IWKp3Z
P+XbjlRKSvAMRL4mtb0iposxLc6sHm8qtVYMAHD13+iilNG44Zkq1W0F7HpK
kb0DM0IlVz3XHh8yS7cMC+LmI5Zr3DAksmSQ6FeN9HRcYwC8GzE5eVhwP7JJ
3QO6894x5SadjziIttMYOogleB9zdE4c9gqrRNUND9CG2yUa6JGlUoEP9H06
CAuAaxZLVZWieGJL/3EARUHHkvipFGGPlXiNtUrh5w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dOY6Pdzs44gHOSy0PrwOBva0dWZcCe+vlL0o0MYWsa3GyJxFocH8mloVDNGt
K/dfcoc6sWSrVicgYdn7buy9Pm6L+FQrw4uxiF6BRq8gLjuDqo0kmMEO0a0n
PbjKVQA5esBfCQIgdfufUYWg1ZLpSTz3nomRLl191wpPqJ4s03dieIR3NI8r
655BfzSgjgtY8J8J6YMYAg4NLa86gN93VaE4yQmZvKulAg9zhYE/fw9Qp3GU
BBPZZyK31skSFdHExsIsYifx/7vXpsotvM1FdbMrOnCWHa6EJtEphwB4dCNf
rcapS9cYggHnD9lztXFmtWiVXS9XrQreGU21YTXQDw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
htW2HOjSGKxl05QBBfWv4IXwlY/+nBQ3jEWQ7vYk0dDMuLe+2iWGBH7etr/h
W/D1fRMiFHQcOjwN7L5mZxnnt7hxNq6aG0byh+V5jU0BtJ85DbKo8kgDchO9
NkTWXIA5ITL5/f2ZbbvIjnAgAIyXxcXsfP0SBrjZhQSr5ouHxtbvu0JPQY5L
qTGDJvvyWyV0LZAQterhmUtXRTL2FrR6NwD+/nsbRxaol1/U5WRXyWtPgXRK
6KiuWQC2k6S4N1vep37o8+50IMUrZZOuQ4FfYy/GF1FDmp8udP/8vjLefp+d
1LdtvxvkqGLQHWGFFI/0gQsmizggL3lKhWTbp6p1Ew==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZhalCNCP1FMIykz2QellIgzTTKum+b8TRwwhqfuzq9/mnkQs9ybiNWdZewBK
KQNC7bBH9EZwz/TQZzKJBdtdbPbkG/3IPaB4iKFwD3NbkPJVuXFiiuo6sfYP
Xna1dUf0TxDPsPQOtEWP6uEeUbw5cHhkGSa/OW52cWFTKctztB0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
k6KY1NxkBsgR4HXnlCLidY4/cMWaonsM9IEpuq7B51ywW2e7F1q4Ea61ytdM
Q1cnmiuyCGPxWY0PHQzZCgeTs4VGQEW1hNnxgrZZgJgGdSjqBO95ABEqNUD+
LbBJwumqcrO3DIuWKfaSgeSVv6v4/+6VNKD+lZ5TfhLdBk7JqJh0RAAHwsFT
Kt8WudGqbyR7n5l7Z429Y1+M/HbsdnHyHpOtIh8r9w9gz9dHLK2QH8kQAhv5
A065+vozZGys1/0MzLl/0P4FMTKFEqe5f+UJPjoyprA0tEKRsNkMBNW3/UZn
gnvCRHlTwgnhdHIFGF6z6shl2aRVKNVyDFj9Glb1o3PRdyCGWj1Byu+/SBkz
92gp0nTtnQGxqXioN2JmLGkm9QZ9yJ+484+Tjob9zDFCclrbQVFyKXA9+nae
w7w2zPmyNCquMCotDocG535LOOp7OYkc3hyhSpwxklyo8deyvpISU1SGRFuX
8aGjXATQJWNC/I380n/my/a5kizfyVek


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LJMUsbCU8WoPjltxk2Y/OIvKSvUMn80qCgxPJHlu7cTjIS2WqwOZ4vas90oi
yvG2vkkhUThSaSzArekh17ShzA44T5IeAe23pPPmkJwPFnAMhlFij8UyYACI
Cwbiu6kMRrV31he8V2OhOIIGR3q1cqaGrMrsH4wtRTat2tx1AZo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
coEGJoezPF+PuYQ8R2KHHp/yTsL+NGC1ICyCggBvzTPCDAOq3KWiEK71fIc9
JA7vpkbOUdPw9f/52JsEf08Ukp7vjJbdmIV9wOPtA1beqlaaBJhZqoS91y8D
DCEVT0JqknxwaICTQxsBf+yc++yBXN+y2d0d7UjHBM89UOCqOj0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15904)
`pragma protect data_block
axQaAjZqZf75NVDd5Yzlunk50DcIM7aq5H6GqXr5I3TvgHhbzoIqXIM17W3r
q1G+knO6l2EwVUMWg/Gmz/NAQT57Y+n5Ypk47J98vylAfZYKMAjHg4aBvlxo
aZ4kNqt0nrG6RKAEIM/dseXi7KlETrboW0XEf+YBaFYs4yoSZemThkpRX7cT
KGKbp+VqbgqNiwb8gj5Kst60mY+l6ko8M1ZdEzEv4JbxYRwxqyB/+R4vz1Kt
hwxk+v0wIsBd9czpKeyd3Hvm7p0SaAqL86Xh8FWf1As5tN69uGigbXnoC4JI
+g2MTnQQqj9VQjvIneEhl2AksdWaUgC1EuDCETwrPD59t1NvNg+DJw0gO50d
0wTIdIIB0Jc3TcLEwr+9PS1Ooe050Lah91EnI53TGxizT/VY3B36btErLvEM
Z0SWqWB7rG+76Ho27Scq1DFb7kh/NHOj/LilKjRD5lgPs7XSRZlH+HrbazNw
pvHpJfWCgldwS75eTC7rggcJ7vD5QTZcGejsRerFg17OZyZzxhH7sQa/+Ilg
/EVMhxq6npP0AXPxxQ8uHRUXtrQwo0WAEMjR1Lcn+ZskozZuLKGQ9plzR1An
+Lz91KMKN+/l4MLb5ap7by1zrfR5acVygBRMCpGOK314v7DYsmjpJpeDIjmh
dQMyPSxTGlKvwyK1EBd4Q3Z6F8AnA57e2PuuRGbeWi1RbA0l4bzutunQHI0i
4u+TEKA3aVgteil9YlHYfKFePFvnJ+XI9q7f6g6FpU+QUL2lmooVahpve6ro
EemgMgnKy9/sd4yk8BrhccPGrURLIxyzyherGwY0HZ6DIqFvO4ui0UP5q7yq
D+HP9Ehj6BtwKkzhg7JEIXFwacIzn+R94V8hz4WMehmw7n2i+o48AcPWDBo3
6pGoQKUdDBclEwBWAevC6klGaph0Dkw46CL3CE9Ji9UF9kzivqeg9wnh7OeN
632EoQxsInfBD4t0Wblik/d78hr7uLXq82XJtosz0Ctyuk6i1WzkonpjlxjU
En9/Ri8UxbEnqH0bIDxR9w4RbQGmJ9tK+3ZFLuRinO88iMOmsnOQ1aGUL6oY
4yU+ixSF2W3LNSfXQZR06bW7h1fCHjCAnEHpAWmbBd2SkWvwlPeusHNwvA/h
Qur0WLVkSRAwMcKKOT+lT2ByMJvEpsOQ7f5dGMUQ8RGKIJV35NjDkSCt90yb
Qv7p8CcvtMYbrLTtw+YBp1AFe2qg3n+HGQ4GxnP35ef8IK6o3nQxbHdnRx16
8KTQAvBULez+2tO5CXzozqCK+01hnMzqWujtynXgARr+n9rC5AXLgasmml5R
niydP/xgHsLktDok13KHxRV/bToEMnZWF1fKSVRWwabYwrrNEvO/u8wXWusr
hnnzGIHafaABySNAld2/TYNqdl77Uy+2qOeDypd8k2YyyOR7EvV4exIFqXQy
Uyp7igbOrrtBmhceWok64TzMUYqrpYOr8W21DMHX/V+TWEMIOdqfkWUONZLf
oGkHmffqlea3wCHWGR0SFuelz3vRcLkkC7/G4nHcKjsYjgr70UCwDN+vb9AX
rXq6NhpvuaYoL/IbOSMKt9cljCGFDkvMM+O+uLUMxnlrmL2DmxucKtS+uQRE
sTqmg6WfNXMouDe0rxP6oKOk+ZxUW6/zUcyBqimzCuYLEVvpSeQuIIOvVc1v
866JjoB7JWJulz77iF5VLV41c2nOp+ODKpdjWh8ONDzn++ijFL+AUucsLuaN
9m3z+Lvp6QGoO0APYNHKTIZoQXhJ1dvyIzwXl7UU3Pcd8f5KB7dy3EmYSOPY
cE4K1z6VQdOkRpnnGCijMXIe5eAxt66Y8YVQWAWNr1wnh3khSYTMmWIqIJaI
vXZgoListkVUnDy86OZygfVNmSMAaC5jnraPp6pZLDrycaCvosbFEG/80/GY
PVGr2FRh0eB2BV42o0ijmqFppYDtxf8Pvof0NAGmsYSuvDwxoyHXk40c49/S
NuynGX8tWkqhyXQ4iODIFZllMaGqvvrKWNSIldChw79DFHQZcHGGs3aAeuTy
USbvg2dOEJnaBMXGAefHX0X2+cBC7leogdSkOY3XkSSTkiL/aR/Pk9cTE750
1d3Ak/NMv+iSMFig0lBK/fuXndj1lD8wnRTXSgBAw2EUAW1alXMg/Nul+RMX
4u4f9AxksFfKrJLd3Ou7eXMh0IZDRsE71imL4JdMzQnI3I6PUshthmpiB0Fr
AEojg0miAsYqzobtCp9XKcARGV5kAOUCCThqQX4+raob4em2Kz7Cc5zBbPMk
G9t8v9BtNIJ8ZFm0d+m1lJLyTMbATXp2FbMVfveJK8HYgxMBozIqz0GMYgg+
MqcgU2qfLAwkCA2Ya6YpErxUAnpirjwh/4K3A9aGwBIkX/Z4BRQf5xwWynB0
QLk/b6d1PtsNFUs5x5gYOPJnjchAeq2+bee+43eJ2hU0RRzbkiY9nhtGij51
xXeyxX2xOCeod+5U3M7BvgZVvnO9lRBPIj2rnPCl9z5gJErQBSfe5XMqMrWH
9tQntr3zDU5su/omgI5X/OXAmlIEm90b6xzfWtVycurDhPDB5Syh3he5OrCi
MWTy473kK0KISRqCrXMLxxvkS87P7MtBDzb6vOzjZJrETCwPPmdL964vcOt2
/ERi9PFtl38+xdQRkORsAWV+jRgJti7wol/6QefDnD1vm0u5bWOEU2WSPtsU
Eu6itcB68Fu+pqcO7GSrsxLdtl8VRQVGVANBr+GdBQLCFOnOx4P0P/POci6I
Or7IWViRIlasZkwYTF7hi+iRflCDTS5JzgfrZeoKW33U6Qo4OOld5kvMW+Me
Ek5KDcagyuVi7jGjLQb/3tQTbE6dB/73nJkWIzwNHJY6KchxM7OZ50ExFI58
9cq9LSqHSmaiksY8/7QwaeGw4F18xrDpsJXKAD/0xWelP6Y+F9446m0e9Gou
x9WNC9wIucrEWxzwNnfqN9qZYd7KbAkceeWu3RT73QtYgpfwDBaE96fF0tTw
7V4KtcsQKwsh9Zq2OwDPilL7qYE1DMWZOsfrc8kUdjlimf78672JzxKD5ruA
NjnsUqHHDyRDJ1jHCbTsC6V74jb8X0J91FTIb8rBlWbvPANQzPUrCWh/wi43
xStAH17rCqtl2a5JOayilU5v0erfFIl8g2sdv2SuvZ50FC8vXPQLTK96UTMy
yxXfkf3d3IGrRhouVDte4GYnuXtew1WPhvEZiiyDk3P/qDYf2mlJGBvTk6mg
icNEbW+oKkw2wXgR2+I8Yqy/t5d76T2QvkkdIBYY92fzcheoyWiT7rUxdbQY
cSKzCTSr6yXiMCRqyOo1KtL4C9ryuNDy4Bwghc1zDo/p5ilQo/UaFv0/QFHj
DWlIolpIxQtElI7cPptAItpV/QWKMcEC85mZV9C1ngu63adCCmN6/ZWR7zHZ
+FYTJQza0QYDseyCSxQJstIUkYqCsjyd7NuyLDwScDoNjQlOXE9m+v2TlEdd
H5+egqehIHyT9MfOR3vqQjSgWTbpKlqnGebcpcZRR3EFM+TtGzlZVSWHgFhc
6Ttfo+Nd6Gj3w3F4kMRy0YkqvkpLsPq7ZVO/E9QSxv5hy8gYtUHwjhwJkqwO
lqOFSe5pjgw/q3hzWhavgkIVsQOImEIGasZQ1WYExH1Hde8yF5yUHfb7LP8y
+JotcoD2HuTzAg/ZfG6aZXTeWIfStYLrwMrq+ZdojL52PUXMdievoFRnsh9u
0JBN+NyzhgDZ4Jbukm2rcolHeBlqB3/3gBVDE+k/8e6Nl7p0IhSJj2kMNO4a
vfjbog5Dmmd00SbViZUS9JspeIXKxXUUVoZVKQC2kmPOM0Rq+jqrxRwfiTDj
FRhtiMALfTAaXLgh0cOgtAfPqslXTdpijWAAMbP8vZn69eColiobz7GK3NaY
ziOVh0B7+2SDyEFqU1T8AoFxAifQkTBEXSXI57SI5LZKKhXseYKra+poGC4R
SFkHIK0cMSMfmw8FTdIY1sz+gstnjU1gysdqnUPqLhM/rIGt5Yfq7UXWkwMf
Gb98Hq6h0/5cbB5XVKIYT3p+fjYuetHjZ2Ff4qsX64lwKjFUMzvbiPpYFcnh
P7CLKeTw6eOHlY3L21uVA1jiBTNJmhYgJ9Acx0ywq+9/6ok93vnXaGSZF5qR
XPKDLgqHMRla1BwhkV4x9j/VoCSFkZbOX1y1yTtKhOx9StCcXIsimjvsdsj5
R9WlMobX1xj7S51Pd1vCwwrrxa6ZCJhUYe6KZSCyQ3fej4maLBMVlpJ3wMN/
PyJz/QGATu926py85xkTItc3lY59qmfH0rQvi4V0hQ9J99+xT2vVvYHg3dZD
NCWnuhNPDSak/bL/NcseRutGCrozYOYjBJVMme51TSeUH3JsELuvBu2gB69i
nz4c5J4HHSyHlgmCg0F2nsjiR72v/1/7VfAleizvZaFYa+DNUGguEoCez6La
AMo9+67hJuhnplVBhfSIKYz6sKgQvBwgOlCm+ZCJS5mfi/1gybyKGDyrOrUn
3nlZVDpZDAN5iIfsA8a96qcR/voxGb59Yoq2ClENs0fu4qewMa8CUsNJCjS2
hophq8WkmLHIFlFsPPltpcAZLaZ7T+v1HQNiA8YkPjEBrgQadigSn2JzkYEw
nlFGQEBk7DG7wPWznua2q8e/G7o4M17NilYw/bVTcIKZkOJMydl7fHVEBJxw
UUEh71KriapcvFQgxJD+1vQ7LldJ1WVKp1JY2Pl1AtsWpI4o37y3r2hvzidu
iZDRhsVvHA4sQvLRRM9EywKMjczV02Fei8Q+yfOeC2/+FSVws9W33OA9nPUr
K1xMqFliate21SzieS31Pn44J6dKIaRxTS1TeX2/t6Gr6e7hwO37cYVn+Q87
vKMNoYBauXeFD3CxUqyuiRZtpDUl3En6tZwXBUb+xPx2dO5o49W1NeDoFCcS
aPuAnNTiaPjMi3TFReSCVN2qcqbUWuQ4mMeelW5xDvTjqU2h8qn+mYZeStIG
tC0k5QftAMbhxcolgG96Z5SBu/qXMwnS7Wky9RQEBYuPXYDWy4Bm81ZPIY/p
z9xzEtKGgVwlL3cTPNNStItJDCM6XTgJAYYj6HjGK4Nv2qAbT16teg0nTuVh
ipZA+tahAk1KR84z2/ZfBFf30PMYxUYIk56kw1hKK3bt2JSuoFZ7dKdEdbA4
ipE/wJ9CxsdbOyruG7sfY4QK4BGMQFYIMmuNGEMJIXSa0JyM6SMRAO+kmZDx
IZdJrNo8Dvb3DHhIvilo8q7n5YmICo/PoH+KYaa5vqWPv8VqPMsoLarHB1SF
cPd5LAsFewEcerSWqb/rDzEvKVOD3n03FzUvgoaaugd6vFGVzR5buqEHpuO0
4Wb/6p4llIFEfYqW6BdMA1yiNImpp7RtRXreROTxYoMvTRPscMyeIPbqN5c7
mWLJEmqtWvJj5PBo3obG68gMtFQ1a5v5mw7pif72kHY9qjh6JQAFyT04BKXt
JbVfYybJHo/Rjj0sYGj7nsXoRWeQhbK7Cz+eDut6F4fjGQKKoNY5WKxrYlM6
dwNRmVi8fJ3jvi+j/evKSjCOBBTOCZe4o5lVmIXO95+cNPYVN7avf+R9dTbk
osj6U5dBPIlNWHEjChhIW02VtwsfTRujadFnLv+mv3M7/lOdAOahyozXQI+W
dr2FYloH8E8Td/N6tmDtSbtPwPtT5ZN9PpGNEFH3APPymnp1jXEpQDP5IUyp
JKT9sra0M6qweU9phE3Bam5rqaQAeHYyR/7fZ7uNwBcoKqIHCZH9vHEILi5d
WNINp1YNaujegoicF642s88EL3dW7TBZlo0FMu8AKvmVjcJy1W88i3Z+/eOO
IzFPZ11Iwf0sTfpsnDEE+jDvvMemFjQ2w4euYj/k2k83tYKB+N4nY7O8GOSs
otmUM6ub70OQhyqY5I3TYsB2NqU+YSGJ26I8zgV04/76fsxY5U28utPT5Fd/
Xv7IUeGEZlPoDmAoF7olmHgBzk6woqlrmj2rTjsVfz2CKZJJ3jDjhI9BWs8w
Y5flubpHSShZq8dO7dVkA5AhgGJJPMZVYNKDXCc4oOaD4cpZppOgX3A5DxFx
AvFhIFdstFWZJt77Mx0SJbL9QTDHDvefbnSi8/hQlLu0LFusO1Y9rrepgxAD
Byb+FmUTLy9CYbsrMT8rIIzbb4IiVzy6ARYtfKRtac7zQTuEPZTLFqm2mku/
Gmy+fikaoIyq879R2nhQBPqj7hSSy9ys5b8CZ6CBw5oDyRDPRGdbu/ukTLNE
SILNJ1OhD3ukJOO4EOzIMZb5CRiMQ85bnBfQdEIj338AVq4JOfdI1tvWKBI3
Gem1k31qA/dU3oCYhj36Xp75jtCRBaSmVOhr5TWEvPQh6xtfBwgf0+rh7EHO
kd5iHVcOG0uXeHRKD5cUGZCyPflZ4v71kVQ8C176C3KvEqYT4N5kMTkzH96q
+gf80GXFcOAUhFa0yQYGXrGzNgEk9qmQ02fZR6ClVmok3kWeBIapQWOMtWvR
bQI8QJwRJ48xFChkc4e9ZAWUltSQsJm4LFlNnYRV8KEmPu5VJKacztIcboFE
j9osowE2iA12hD7fegp6rj1Im+Z1ze/dwLhIE4uyLfLTso0EQIDFx1fFvmwW
IT+j+Z1qnHR16VpB/zhb1gjbKN5a1UEqH2UEHJturM9mm4AMeczsfGJQzmCZ
EIjLp/ehemTSi3cmk0c+R2rph6rL40CCGJglrCy0PlSIHfqWfdkQN1TwY4MM
uf6kmUKmIhHGrw+Q7PktTiYy5KhjRVNKklaHkPdihcCpIaOXNx5Lddkw4+TT
3S/zMcWGMvEtqT+xC66HgHPD6eSMvv7Fft6JGtmHwltM84YMW02PrT6QYTLY
eVGBTR9uwK7+6CUECFVubADf2FK2eRwbY2EocjFqYxnqLMtgfPrBaxbR+M23
BGL24obNhEV/ZuzxkYA7VqyeXzP6HwGbQMJ6IVzmBr1BvsNNEibcepKs4zUk
tRr/KZ0xNtQmmRRWPXKiWjfySPF+BxFBV8vMYRqLRmDS3lgt/jzpIHwWDV1A
vaSekpIYj+/xD8jU3Hy/c7eKy+BnkC7DizTf8ewUKObaj6YhfH3F+B+NQ4wE
iv0DJKDQLSCYhQaDrczkX/OTCA6v1P80k/pCddbQFad1cFnzN26R5Ae3qR5B
PnrC4LiL7+Ux1QQMvsNDVQHP1hZFfMXfk5nfbRR/crSFj3Cc9I3Bwkt65AiF
fZ196eqMioIwjDHMJdUhNBGGDV1SQ2J2QBgvrY8DAjzju2O+FMS6SSb9o3qY
vyHv0cix5IWGl41AnyuXp1RT5DYoaOhpIbyuP8J5MrgHtTWo2LtZqe0ouTDg
U1yrN0Lw7XTAlWB3qzTvSBv4p05Te35CVHTr6HH2YeEUszKtNLqjZ15ATArO
5HzCI1b9sqItPUeEg81OosgiTqqZfpF/WAY/3Y++jxpo05bshQWqJvHt0Nnf
VoD1ildiQAGDSwzzz/Br4J/ycCLRlhMEIVkDeWfYRwBzwx2kp6cZSi8Ou6aq
nr1ePeg4zvKoHY+xzRCuAEGoUY/gQFqmFt+eRB30Xm4dXMjyUiowPatPDaGn
Pc34WvMQK99dn8/fKGZSbSztsz7mIlq2qeSX5g5jdFYU7dvIFEZ32Qq37ENR
aGghj9rSYWHlfcxwmVaPP85aBLcQiMUQilz+A3pMZRtNwiXWEMcNKnSQmHQg
3jbgHSHaa778+jPHaSVeQ+8sgD5eSltTFKTAj/X+M1doiVOzWGRpIfZaXLTK
+IIFubLEZKhmBU3ruDkw1o3/1cPl0OsNuF9c705wHmXMPoVFoJSug1Ar6fje
YwMSR0fivUKWIPuiFETupW4onkLDW3kPfiAJItQPeYguvaGISaL7wQtgN6bg
vTz4nqCJ6mILtKO+sDCAClxQEXTDBAFLJuLhTMCEyCygpNM97X1bDZOs6UOd
0o2vRVoAG7g8QeDpjfAoeH6kUDWLfU+ZJqExHWfupUXpHzj8Zd2L0Il/N2Wj
egR5QwFzGKjNLU2M5LxSjgsFnUIUoWgxzND8Dr59iLvirPzxi0P4SRZn+ozh
vX8csOhpgjc371GhGWkCcgxOyo1jdRmbr9GEC3ZMoRClKTAwA6AqJOhTtU31
J2Yv4LPjgBs7q4P0ETkTX94+zfHLrWdsFamox9hYbZUAYMV+6qQvc4cT8MPg
OHR5T4Lo7KiCa9qBj4PizhVEpSvBLrih8TS/Of7OcpcJfHahbKXlxLMEKqXf
8UvqVEG0dZXTvnlVoeL15aWpHBoJK23Z2KaLOIzZhXz07J/UvwV3AOP6q4ix
5ps3oz+Qz7jPs0kHwkvGL3ECVzQGblD7ia83Uevy+NtzZaf3Ddhr5hC1+zB+
sR6ibg58EDeIBw5H1CGpUqpTyq2/zLeU6rUnRxlJPAAgDB6lW/R0/UJnlBnf
rGFPcxrolUZ/dN54jmNhLzDD6iZp0S0loi2ubJAtIvv0PHSakIK2i7tZpdnc
tqazdrbId9VsGS8XLzzhH65C2DsQOgViXOhjPZ9pqGMCf8ADDeEqDx5SqL+u
zprmp7/2DEnDMS1n/b7Y+OZP67lE/zQH3q2dRumJLCqAKlfJ2qKEU4MhQdEy
f1YvyI4V0Igp9pYJXXpsDqpik3cRvPPnS4AW2+q+S8q0/BzSQTfh+W4UO00w
cEq6ohiMYQkVpK6EbI/z+3A+UzecUFOd6G2SQVGhShF6p1RVOiCBv+rvWOFI
Ofy6ZcRG2pJ8ULWPftZQVPG66lcYv7CFdXzSEI8Le+cjQTCpLtF2NoOQA4hJ
O9RGTzVcyDWKV+sy2T8syWeJJo/yyf4CSd0wxPNzqGj2qpvtJazZj5KZV751
vOp7QtJ0V5tZ97oM1hz+BE1wnJy42K775GGiUe0iHDoC7pu9raCcA+pmaOIi
EVZTEzZmODjN+PUw2YZRq7lm4+uo9LEVB4VXQFkLlnbugB+gnq6jE8NvexYv
uvz3fBdt/sPwOsuYt+N8YdtYypyeN071YStGyW9Q0NE0J4eoIXFCVRv2YlCB
RkQk77xYwXnI2nimtyPcQlYS+hkEQvqnLJKvcCgs6JTcBKqLZLwtCU2CHrxU
DvUTYAdge4xxlnLsftOQ0+RegV66TByVZ1LxV+7xDF9tkdlBmfilF/N8MBug
T2RlMY5OCFhz4UgyNSiI5U68u+rRSAhiiq0n/gr7LeRdGBv82JOLYSK2pH4O
ZPoF0stkiXv7St3PQZW89brde8+1iJqVBdPCnhdpD02nkNAic5rHFnwcDoYv
p7RItb/UZIQJgWjEKCM0bFuJ/PTf0sKft3qXkfvdlj1BCTFhdfyh/7l8HBC1
qfVK2ppgIhYFzLpnAQSFNWxdgSHdjVzinDMixNKP+AGZWpCxDGX7I3KRA049
kst84UDLC7u1ypCPgycp028ZnW/p2FiXfwczUIbRkW6gsN7kF2zV3ZZ2COvw
Wo4URqxtx0zTsGEtKeVovtglXEB5lyGjGhp2ZsaTaifZ3JayROJYtX4ZCmab
YMs7ThI2dmp2cY5Ac0uaPDvxhZ1d9mTDt47zJRTrHoqdDzLEQOXMWrT85r3l
JDq0r2whBxdPPzBih87vT/UHczQLVf87vX4LcifuuwhOgiMlYSt3o2OOl7RQ
hJ+EN9YgMoKhpL6JeWu33KDzJ0rUHxt1lk6aI5BrcpYTsGjRW2xUZNDwe1JC
e5srNgure81h3oRnWx+yVxC3pA/7jRYKLtQd+lIzAEMQHvAwhzY/7pkIlRID
WNMvD3WT07u0cpRu1oUAm3eXx5zflDNKeizy4cBTX6rxUgrZyPfSd8UwS5nG
GLcQ9mcrSl1fAaIzqcc/ZIEXHpgWDhqsdryp+vfJaLvo4PaUaNZq4wz7UNkU
NP8zW+QUcvvZGmm9osMRzzHhk9H8VugKu0qtJpEaJC4rW8EkXOPPXgtIrC7L
IAef4pNbiFmGZjRIsGIBQso7bueUOz9scBw2lc1VKG6zwBgDDVzv+5RSB8Xh
TNLTJL92ObP4zVyXAR9VqC9DAu3cCzbjo8HwP22m1mx8b6QO5smRbUmSXX8d
ybzejXZehrriLDDHotn8zeXyHYa7iDvScbN48JAxw3Yss8/h9ZFuaEznpYLg
zU4KHFvWovBIKDalgPvOIGcsmYgSUlh2n+ISRfflGd71cWaIozcLGKtmJdpR
w9vcY6Lb3JxM1F7xBCWoVCDxDNlWhUnQ8qqOzPyg9TH/vL0PqId2CdtFn1n+
wtIvLt6fM9cveNAHDL826GRIXTBtBZbAGF4WWzy0UDb9jNNsTdhnpO4Yn9ec
sq0r3JfeoSzm2dhEC28VsTUxk+TUBDJrDEKAXdtyE2jWr9NXqGxJnINV91wq
v7fscOccrnns7meH4dY7dG+I/1JNXolexeBEALWdq/fOW2z8Gnpvw35/gN7l
9P4oFRldtoPMSVFhsqt9xgKTfgImSOkrzWP057voBXrXJV3npxf59cv2zqfl
2L+e19q3+tlqosrgwjdgp+U8ZUsLBou51rm24XaAD31z1SBJgunsq7wAWk73
f9Ic4/30n0Vn3dwWIK3D1j9PfbBxlno7ho/MW+5FgQyadUUqOZVEx9VxLtF8
YjV3CERqaQ9gsEgGsdlDwQN5SPMG0XC4DnSbH4togV2AlMMK7GT5DSHRG6Cv
RtE6xmJ1UFLL+ouSlFXsVr/U7QG4NHJQubYD7HYfzRzrgJMhjszEEwLj11OX
AtUxj7LFx57V4Z7YQGxMQN7xCplEyxqF07Ot6iPkivJT2Q5r5AN1wkOgRPWW
PYbc3FynDyd5I27lJNJjog+nJ+5RwZDLEMpkwQrJMPREEDktoPVcrvod7bru
179QNujQ+lgDY9eddNXFxA4i32wNYYzbwhHhagUV1BbxC4AQ1Z9QPoo9s+7X
T4Loysp9PwdaOdhwwTfJPh1C/CSamR3D2uejoWTQKlUdjoHMwibfGH3z91kb
ACLqCX+i9V6VSYHc9WASR85TZmCKLaUSfyL6UF7N631gVg41yhtLxWJYMOef
b9JCtRv2aTjwXZDuznbFlchTYYilyQd0GB0Jf/iwngyZkGDFETWfhZQkHvep
aX+/xw+UZbTmElVrcPckKlTrU0HFF1vBKNJ/9aOF/aLx3D2n84OuvHjaZ2u+
UdYJ/KBf1+G1F3SvO77/xCtN3v2hYXApdtmeRk73/bzz8yQqFJO0rdwlsSkx
wxbUjjiYBrQzhHbCaAKokYUbz3h803GtjakAimowuh+0TPo5lr5Dvq5xJMhJ
CKJytrV+IwUkXLqt+bEhpk/fje30eN0uc+LR6oDSN0oXHz864/4pDanwjbrC
kjYpvWU56bw5JoZDTQvnLHzsYqiesmSSgId23KxnVbidT35OxUSIva7DHrQh
bs2jeE8rFBKNhkQIxsl9+qsWFkitWUdmOfyqYOXUH0Y3nTB4BrJ8T1fsWFRI
c5x9f/YQz6Yg0UwS8u9IaRJwpQVqHeqbwTWdM8X/X3n6QPV3RJ92/X3tisbo
x6S7IubeN4A4MoQrmbhyyzcMPr3LNpsGhAPxVD0kpDIv7TWez3RNPjpD7ydg
0SUXuD1p9Y5zKl6FM2oN1EcGHX/BlO4psKFwfIgGbnbwvgnuSkajgbcozC/y
Q6OFFoB7/KfTWA3FLbSUHyBHQUUxgDDlRpyjwJGeWtS8Z0Y9JTkk62yMDb4a
31QvMBb8kI2rWijbHuSM5eAT9bUUpvUddhYzEYOEX9Znc4b+2PmK9PDYNPWe
TDmTLhl9bjqigckfuUsvLWUuMKb8te65FsACmjSt+C6XM78RMQznFEFqImkd
OkYJ/aYg4Jy8O6pLx+RUkLeB5onZGoR0xxnorL7mvmto1v3z3YdwXUqSPeTm
HeeQLFX+C18vuTrJs4b98i2JhE4R/8nzFaq9tZl1eqcQ/EmXifrI2onDZNDY
KIo1JfSVBy27CptSLuUHCqCE2v/V6ABmW48PL/BcZxnD5HH+6gB8+n7XGAsj
kwNe81hfHxb5Yy1WeAlzugkEmZ+xKDHGKxSorQV/2X6Jb+Beq98AIcuRBChq
1pPyTMj/GpNWybyWe7MLAEaFV5H8vc/+Ys5Aar7TM4uJk5fkqbtNaHZm7iKk
jLvkl2FQjEHB1p0AmoNcTVOORjpvJ2OizRt/WFVaPXgqVoF5PB1JMRvntwKm
JZWOIT5JVn4+pN2gmgj9BCBuXtNe9sauWVkEu0zcbJ+FTtlRbmc135UpYZM2
ROw2qDqZPRFleP/DytoCujR/HBUggyU1tZs3mymcXzb/KEzxHIt+YMAAcGyU
8xRmpHioce7WAuxJqSkWZpnsA1EKfxqDjAy7mKKBX7L/mVVN9yWRcTFoBovJ
EcetvGKvILMh5/NOSlmdCjQi8+Af0TGv4hCqj+PaXEFiUJjlGXXAnGwL+5uo
FeVcwY8zGS0uJTWky2l3GqJssy5iSxKI2Y4rp/m1YctndBWvPgplWj0mTZEP
xKg57LF4vD8b36ZcVd1CBWhAjijF6bgrw9Z5GwQ5CLB1xIxQmi0gkgOiHyxg
LZHrBrGD7BeAb21GUZToZTNnwVopPYpqgQldDn4g3Odnt6uwZ79wKzVSa3np
oCk72gLQAcPJG+oO9VDHm4/c4k/XPV+NPc3HZG/dyeRw86hrpnZBkjAnn5AL
30b4lc1Z4sS4I6jR39b3THAxOtHVxKaGgEzvmE+9lyqAbCkI7Gg1f+6AVNM7
JtIPWMV+6k85eDe6nZrRTwRddC1Qs78EZ15cd2FWsAcB8W8N/pNgYiVKunA5
PqovHDbJAV7Uxx93bSClURMoTRCsqJxcvYLVRt/+M8tCaI+6P6O/kGi0yqho
6S18IBuFiVcsDv+hjKgnMnczG+GHPwqjktB2HVf6T1UkxXZ+beVq+qxqHi0a
FTi8KMbLiDq1w6Jcpz5u3kzZ5sYXTWJsAWaLVWBEInIhfRb/YwPCv004enro
nBJW9+OO5Y8Xo5GjKMrPkGILwkLp66IBG8Cm/Ng7W+544JPIpUcU9SzAWHSi
xICIBRyjNs9hNo5RxYmbqDZQ5wCowuIHl32UVgnLeI5JZv94rlC3x9qaI67x
UD6sXT6dEVhngJUjGhBPuw3iKcHnxaEOeTpusTq/P+rwEf1IzMPuVTNyPyUO
awFbpW94yvUepU2pYuJfGJfHS7f+5/TE0j1LqMt+RYsrGVp2Mm478x/6AZq/
jduFEztNkf4lv1HxQqjs+wgQxFVuPmyLLBjg3wSkNfjAIrM9ZfO1EC/P+rBp
6tVxtWvuLN5KZK63LYSS2dz3rkmGmYEqCWqqgsm8diffhNO2CbuzL7PNfVAi
AvPNOQAcv95NnHgODb3oySr14S3knjGxaoJyQOMlKIy7CaSe9L6dJABOHJXc
N+kqmMNBtciDHPZfXD+8/53EETq7MgoduNczV1MCexrEnL/e5zl/q+nVNqma
KB+e3a+1gCkoRYu6mIbadjquiQJfhYb8GQJ1CGGD3yNY4RCWvzlwMSmtxZ2j
SbESVArx/ujZ7hukZB7qvyqpk33+HcghYld0Gd01yoxZ2QAm6VrsfhXNoU5V
aiXPTqo6MEnc4yekoEjTZ973kOPWMCf/bi081xU2t8ONQYkLbWCXYricaHAy
oSwtl6RzgThNre/TninJo5KYhtvqM8elqyXw5XWFw51SuhY1Qm6jt2CIIX9x
JFi/oAy0T0BNh9+p7TEAluLsX0hLqmqFi4HXwtIrUmepOWJs7VdRE3uqzyWU
ePV4zFWVelZ0QxwBK+bLbGOSu1ZoFL2FnDWDDJpZCzgbUtaA1cQtwQCZO5pn
U7Ce85mLEkoX8+gcGEznjgGPnmWbvEY1Ng5lxd8dAwXwTjc5Tu9Gy9JXWAzs
E2Vpz/ZRCqtQu5fo0MJfqJEj3+RchSJTr5fX6K7s4hPDoZw/yof85J/4I0r9
xKscQIJ1bvWFapZtr9FuS5HQ9zY1UeoXAwEh8WQScL71OLth5ViOqLyiGk3f
Re4195GnoJj0qMRGCumAi+TBa//zhdf6l2NIUWs6EaXYVYtKZoNZlBh2ovTk
V10LNrF34dPvYv/Sm7zBAW7ghYaZk9/YQGMb+T1Ld4nXibGqF+BtzC3HLwvI
V103P2ZWD/fMr1ZmmvZsd1zCCKbMw8ho5o45rwbGFa0qpWti6au4j6ACPXKV
2AGC+VYkwVqczJS5/bq1iqWW0vrYS4PfWkt/ZLFXA0gQB/JAzzYChDmKzsVF
vH18RL6poAx0b+87zedqrIlUqYgYwZsHnrfytE1DbRDSlgHGPtELhiuaiOV+
N/z9YaE+K/F3Wnh0zaBP6J54ERF03K8sxd4jUNJaiXi8umwgxpubdywr70PK
v0VC+8CbguCvqUzpCSn4JBrki+Pjr/XmK6SDW8i/te6PVxnCcUMmtMs6uxfA
lhCR1rMbm7f/KuCtsPy+ZERRRUOTZ4TCZ9fLEJIRyAWyMcRc+hyB0H2FMP7k
0s2EpKg06qWqwsulGdS7EiTW5IGg3Oo2dqzj9op7pMFbYP9O8a9lEjmv3CnK
eiEg/dz+GqjKmuLEvRGFCJgKbXMLDm77VHJzpJs0sJ/gtEmGm4bQI5JVL7Qg
xkj9OUc/+1mlw1U6BkEQ0YheqSF6pUQtEi7RQ+lKfWn0x3bAiu48lnFaJdkX
2P4uM0AIF4oz95hlbT6yonXsVxKseJFz4YE51MRnwi8C6Ywnhiril44neIv2
7tobtymaMG3ZiFqYQWdn4mtNhjzCaum8GRzDNyqXMkJ8/a29ra9IZD+uBqB6
QZIgTo0jJFxTuCArQeZhf7ybJeheLGqzDvTOZTAadqLSzOZWmdm2ha/ZF0ym
v8mOmDiZeUHN7UxyTHx7qaFNuT95ljn1wbTrmdrWoEykzgNxtvDobsgn0GfX
bgQzFFzDkNnXkxpoysHNnCdwLgvJTCEM/sjfLswXxDbV8IBmM3iLB8Iw0nmp
ZiGNgyY9tJgw6XEFX/5VSKcobb2un0zdpc7sjwEPhisKmAnkZy4sGx2hl76A
T3E0yTle/Sdnxq/yV7NLtPbMqNKiS6NN6mHw0ohsQ+PhuN6ew9HiVr6GzsAj
DJhT3uCqBGIOBtTYcO1Ql81bDDNmYOTyVtOe2EMarTnDjhgVFU48ES0eHNxc
5QjFtuZE53HokyAAzl1NYvrfgUqXVQHrmbREIamc1vA/09Xy93h2TUxmUqYF
0FOTHjAScjP0ohuqhBpcwsLr2pDfmEVcbfySv/oiBA+42CIIzqWoJqeg9Ork
dhXpBfTA9Y5JTU/e4gkCiIw5zQAXa4uLbiN42zm6uchR5rMniB8XARZQ+DqG
GBMgky/M2tGcfipwkx6qW9OtMWHPQQFkWhD6tb8sGTgWFtRtjwgUq5SrKS/H
lzEYjbY8/bk2RlAb/Etc8lHLA+U+wNPUIPr4ly8arL17p8n/G+AbFnnvyOv/
Xkb6LAmLWL5oK4KzpvILlgFKUEJ5z7BxhatCDCzwBRHn/9WvTie/4qN5OH2R
skaXTapT0UBVMjSd/pgZgk/D70ICbPTAaDK5II/4rFnaR0xsJbVjHRDWmEZy
sjiQCKx/kj/H2fZkj73uFnlSU/KLr2590VuhWAolgQy/ahTs1lvnXGZyShXx
1Vani36PQIZyxbrJan8Pu2pT/GZlN+7tElQNaeBugBVuFdHjXbeSwJTgWI2D
TbbB8ZApbZaUZrSHXoL99l7vKm+QvHwdLHaf6knxGnj3s4+Adifz+tW7RjzA
EzDdaL6Q8tMfZ95t9TCuunG3/y70ogKx4ICnzvpNKqLsdv83/MbWKDkrjvo0
DbEl3FIFedEPfOWtTNPbRqeEfrq0EuzY7gvdE/3cLa+fjuVehzgsmkA/Met1
Rv9jjeSzLqAO1dyc5BynC1eSYvhNfV0GPjE1wzSE8jztJlXacIsHeMVTGD5H
1hXm3fGJFoqx2i7FT5AeOIUMGUKbIGOVYj8PFehaWD2q5aQpC7vVfbpxOQlO
WWOLmoki6CBPYLsdJGjuHyEab68Kfd7f2aKKfhjpsLMJ95y+HdBmpMWgetjC
tlpEXzwhtHrlu2VsJJRFgXMcHiwW9mf7bIOMHscyE4MrYDSGaw4UKDJBuLza
yCSDmlKXki6eynEXe7m2z9N5/lFXJx2dICVH8vU17DrdUeGKE1Gv1dIfOW8L
gTpAjSk5ZMukxrl5xVqmbkX9IPoDLi/4uYIwP09Wr/7izVebih2VOWqEn2Zc
KQ9buYeKT63Zza18ytkg/WAgjUrhIfXfb63xPdpDeoqvC9W/jAbTpILiUV0W
1MuKI5GgMlNNx1tY/otSgSZUtTgShzwxFC1UIsHt71WF9+0qpJfCNe6/PYik
619Vewt4r7MuaXF6+5xEa7d3DPWJJWyvvmkeOSNyogvMgwxfHfK1pDjfJCgy
3WaUTpGgzF9lNEJlJFDcDYj2d91heQLovkRalkFlOcZYmCpjLFiwpZshFfCH
osWy3AByxV49xEdEIustR2nAHbAV5W5ErwX3Qok+VUcwxfGJd2i+CaNZAZUR
AE510PsRgT/Vb9oJn6emcgwDEuZ0y3BOPHx6O0oqX/9z4/M0XM38737bhz/9
ZqCLCTqCTGKZuFYbS/WNR/C+C7fOUpwVRdlkL0Cl91KGW6QybVyHzuz10mWx
zvE8FYRuMOujz4upq22T+IS47yrohCRlxjz2fFCtXQ/aclZZwcIhU7JFN+q4
AjxGz/SLrYuxXbrSqvd4MLY36Z5cm1dOhPVLwRej2T2iMKjznNrdUDFcIUf3
GHMIiXwGYkRbD2GxxYOCnk2yOOivNtqN97lmkBFYnv5O4qAC/xkaoXtDi7sl
/WaUvdxR6nl9Oj9wvgQgwRYqq1/D1l2oyfjZi0Rhlm/LqEHT2kxYqfWvNtj9
+csrdzEwm/I8UqK54gdkv+FtTywJH5Rp8JWthK2dVKwQSoAi2wxPyT1A7fbw
qbd6kgmz55OyA48c2B760d/5VBGwFLPntdbj0LRYTO4cLpBlrbDvHoZyTjiw
eZPp9s0vsz7d0yM+xvVwdTrZTyxYIyumJM8aNvEbqrhUYyFISQf6rPZtLMfz
XpZlSJcLpT9iC96dY5YZDutZhkdySuHgn94ZF5YtjcWOJySHugg2rwy7dFez
ecO3FyC0ovDV7NPZ1dUYQJHlG8YV8Xfyl42MMG2YAv9r1AOmtCUkeBIOWBd6
m1vipCNQqexeAXq4Vf3cUFwZMHg8pv1SGXXqvhqNI0FC55Ha76Yrrh3Mbc/R
wSJooogmyH1IKjrB6xsvQMqAbPHup+K4aDEw5MzZXjWfxAPvbfDQnpcufjjI
8euzPAwjjKcvcbC+j6ATyTLMAY00pMCpiv/v3nfHYQuXjVVy9OxFkZ8TiMqL
4r5rMowFGhV4B98DfKeH20I8+mZaNP0RuuEOjJut+zbbTuYIRvrpY6ksbrQq
rRxHtWg+i+GaQH58Bb7mdlFueRWUpuAixLUFafIW6l+Y3VbKCOD/+iL6gOF/
qYJ1bHU3wOIX5eHXCv5ac69HbKJ+RD6Bl3sRTFdWiQ2HkZwnnDQfkDGoZKyF
qX9Ir0RvAwfBSYjLQgnxzftfpqkV67lekA7e2RLTRGRYeKLwqqldwaTh3GRz
FJslA/LLa9CbTnevJnbht5S7J2oTvPIrlq7hCBpJA92mUwVLzf6sTfjSIpkp
IKqGDPjY+r1OQOW0xsCK1ik41iUWNZFK/YKy5fgpqA4kXY2qaAbk9sctDrvF
aTkwMX3zbGxESZI4yA3RN9R5a14pZd2urgMhDlYN+/iVslFdPmwcSDoCASOH
vH3MBclf2JDQqtrLlcIGBRccQ8/9UNtmE9vg5BluRzJUEriMgwcH4DfO0JKh
m+8shqnRn96iIkK4Gh4Mj46GJhNiWKF6S2l8kPy9x5IwU2F6/n/GmGfpUIRC
Q7GV42AsKPdwD136vhyRW+5uGoEeW09wA0wYYSCIHg3xuKbSb5ccTJMXHfu/
YrvamIReWi0ArA9C6NZOGJeJYy0xY4YJx1WKiJj3i8yHlUCnjF6biSpuCwas
bmsCV40twth9C+d0/ELd6rTjQ5uTxIR5a+qUi/vWVlVkVVK6YnNQaN4x526a
JTIL3iDoFCqV4qwnIl7+mZqSVne7CMMrEjNx9JGN0O6pje5pxahCrD/t9N65
67oGW+CrGUSu2bDMU9wyMqMI2reL8SWzCOjI0NEj4uVkEQ994xdZMVU3nomL
ELhdvvtgvAWSbz9zdMo6NH8/v9X41Dx7aZJ8s/9UGppS/qpNCkf3QFteY43m
5b9UQID4yw+tDrU7fOS5KWKPxBVchSLACm+uCm0xuxv4WRtbsNbEAKoU2NQo
7oHxKEnHzj6sIujgGtiXjXiDgLg9VZ6DwXSc8MUqa+1QoL2rPIgfB+xekVVX
cxYsNL72aLT1hJITfL+drXu2rvmcz1YIHYMMrnW8exawEaePhFGga/QtbwW6
kJXrG/B726989XFizMkUSBnHJrBLgDq1eIsmbwlLzx/lHfVuAJ16w2PHZIbd
Z9ixHfG9jiOLPjTpO4kleL8Xz12FwQ4PsPHyZG3xWeEVcGCYsvUBblc/aa4M
TkWPvZp6yctg/2J/I0kCO0IMk/0Etrl/KDFLlR0Sq6DGKeU/outCFXzgHeeJ
+TkQxbofP7xjID+Jf+9tJcHT8RPfLfv3qb4xg9MKi12kpNdyzzBWGHVuBCZI
L83L2bYQf7MGJMZcavaUEyfTDm5e+V5v/e9S+lAsQ7awxC7kBGBxSVls91YV
M2cWrC2w3+Rn08TKcsg4YEaHNRbSRJfFkor6kcXGjDfBeZaJq/V82JWTZeCr
I41KP+5R3ZTOMuc3nKYl6w3UUEdxE/vmn+KiD/7HZvtnZJilIFd3z3F3gG2P
mcOfM+Rc1EOSF5PIVWGoY+U8sjBuq9Xitv/wCk02ps0IRjQwCTBRwohLW6Ty
YyqjZc40upqBXOqp+zKok+0s+ChA+/THXCgL90IBOSof95kimMZS4+xo6+Zt
K1oclMazPsG+3CS6g6vZsgyny7av5V+DjtAGyoTl6yHcFwd/G56vQo31+pmX
VMaKZIsQwQPfzaGRhC0nXEqTziaeyT34qznmsUB1tuYHVutwsanfaMhkZlDd
SQnm0mE9D9aV1dCNjhfyfMig3LBTy7g4vkCa8CEVhEnhKBJ15JOOs0XUvTwK
3a3l0gXhbjGxIQtYe91bswORhN1mAavMIvcCFgarP8XFgt5BNU30dyL9qJEC
QT9JH0i9owEBcXFYeHYwCTYCXoaw+9ReVdM6tRVp/hzRohV80pJ1XhyuiS0w
meS91ocuI8S68yNCISAdOs5lr6Ml9RX3mSkQ7R7TO/eml3l9OkLTxnQQDM/P
eZbTnAecg90lCuHUrE0MazYm49CxATXJsnxqqR5wcDVig1T3VyRoNDddDOsV
yUvtn2NqwAMI6puTdEZgSw+q+kSTzsnHIY1ZFBuajQrnFvRqZVcev59vG2aN
iedg6qIm8ufaTUJIDhEL4MpUVeJsMlNhUy1pSDLMeACa+O4pfpKmL7dNn/lc
PbXlMSwbXkwHGbGaEpVRc7689vVo83N+Zzm5MjsA3k/Zpq61x9U/Q49xDQgG
wjj6/MCNOZ+TwZ6aC/1iyQOiUNUzZCdtKNdIIPYwzhkVH74n6lL9qlR53GyX
YeVo8bijQrftJkowirBlM4EqGUBtsjBK7wxcvFedfl2jOJoKVWxJO7xnyKqH
d3NRtHxwxnDZSnN5ruVBuTaRZdG5fBQpJSMvNAayPQbM5gKY6hQlgktkhMEV
cb+GdQX6TrC/akdEB3I1so7GPtag9Q2tJXGpR1IgvV5PVIFFQ/NbHAjW5lGZ
TULQqeqMDUC6IjUODAor9LFTSmoVmhCt+vyzvjZEz8gYJfrHvxucrk1cx0kd
3lfuNvtVm95TbIB4ozbhvmWZGjkO7+GT/54pSu0zTN9uzjmDXGT7GA87EWXj
4f5yXcVAC7/6gKCl8o4thvptSS0YQCPiXjk0m2eDLVRq6b5mLTgAAvr5E1eT
IgC0IVauseXDCuYD68VY+mUP4w1NZHKtVQN5nZyeHAb0f6T0fZqzDdWsgPk1
dVHhe/SNP8ZO1Vlix6jpTPIJ159P92ZTgU5KE4YqqIp0VBvcIxBFragukvGa
LPO2E4i+20pd4zczEX6ybcuBHfOKGIoWuDlbR33+t4Brs4P0/RCsMhsTJkl9
KHf8Xp0VBj5+mrYqQPFJ6F6Jow1SbdCo7Raa4viv6EcNeuh/33OP3VP9aCRI
FSdOIiv12dNF1su1CopCFQ25S7jgzokKnQkkm9y25smqCebf0XYhQdiZWoqT
QMIYPBbuJ73qEiZmlE3bC5ozeBbWX1cTs72ND2DqdLz4z2zSraDwHwaxBDZf
eE/yodQNgB6eUQx1daE5xgrrH36md0QvCI2I66/MORlh7gavsaollHIdGixX
SsvyQ5NybPiCeaS4uhauVkKJXIWtDPWQ9TKq+IFxw3R2XwsddNiz0Yjy1PF2
/q0y8H1yw6qtgwI6pB5sMJ/e0NWvWpAIqKg8jAlbVslZvk1ENw/4S4RLgRIg
dYWDbvTYHD4zLgqkPCrgIdKb+loYowPP8vXeTYrVEfkgNEw5mnAYZhquqDr5
HUOleLlIOD4z1KjeoYIhxxrQgMWx9bbGYYul2q3B/k3E5tMkBVq0LatYoJ0A
PsBEFV8JPF5gdU2pldgEcyX7gbrp4SvA+jLCo57Lz6Z40Su3wnhHbX8k6k47
pXATU3b1imiRcDKNyUYvxti0MBSIG8DH+N2lgZ37qrVBe64+QgcgjzQtUxrt
2mKsJ+wr/Ampp8Q2VdnOMkLF1qByxnuIVJzzXJ0USXVujplgDYM7SmtstzSB
n4nCx8XCBjSDTVPwhbvPOPTjnz38Lm/rmeZbyERBh1mPT+lToVpsayxhbz7b
Dz1ALny3/pUflsSfubWrzyfWCW5O2czxSznP61D+mdtKMtAZ7vlJpY9So2QU
zMJB2Lu1aZr7TXNpsCC4tDPGdiyWM6JlxrhK58fl7yT7Vn0t1lEfX4uiX7Uo
Ug4e0M8xK9K99a7eleVapX+r+vwhxdVNsGKHpczE3L5hg9Af9zi/PBKE8LIM
PrzfeNFqNKp0myht5Y7yGNfHQTUbCSHKHHnOMeFcsa1Fz8tspe0XTQK/TkUv
siZNqdBHLhdYpvrakGUcZMk6XyMmRrItygVzLdmylMDcPhYwZwW7eLb6cMuG
jFHFJqxCewGJ9cGLlwzeJ4KtP9sGjWVT/qGwD7Bj/mvuCzBtB2I4eUJApYvb
uOMEUg2KxgT4qTx8ZPg7Im/LRg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1K+/EX5OXcq+V2I+RV+3ozppllcoapt91pFPybslRxuDhC7zOc7E0kwQ/4ph4nwIOKhcNcqaScnXulZZTL8at/15dU0WawD2zJLTJfKMxYtG1D3h1saBPW5Y5j6gVfvPATX7kBSgR/4nc0amCKxGXxKGCJcTmBbCFYa0R7gFDA+qnJRTpLNJaLPT8fEeVsiVuoXtWJ1dFRd2HjpXTWtw4Esfp16YT2pMY+C1Rbbf797J+s6trObi6/mgNaOtum5QxlyL9l/KX0N9Bvf4JOdCRZudoPg0w13tcLa0EGLxevto+W2oZvhfQYjr1rwRkvzgWoPdYf8uVk7TwcFdmwm0GonQlr9JXPseaeJx2tPXEdOVliPWvwS+dollwJ6ZKT8WTVrkn+xIEG6/qBoJauq/gNJ2iYEGTOVRVxlL5IxeMB0IZF/UZiEEwOqq9HAy927FLOf6CHeAV0clFQQNVhLSZT9C8iscm7fQDcNyZ3BPf/1sFod2R3XmQdkVacWD59Jxcad2CF0NsEkELzMTpeE3vlUmatjpSJyXX1CX83NsNp07dvUq21y2AwjeOmvPSukC8EnFOH92IXjEYj1xP9qcB2sZuW3ToYz2cmsR+D+LiJk2vQBVUQjuM81val3Qt81AMKhI751ArUqPxdCC5jeM3ssfgSlX+IUUWOoEsi+kGkIXOhYsmZoQ7TBIttKxKSZsHU3Z1YDQeTEwfRLX2yA7+H6wK4Cmm9MXWa9oKhziEVgosi7QkSmF6dVEMlubY6e/CjGsMtMxjTosr0ZxLKZTjKA"
`endif