// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0sl5MAYi3V9Wsx1ajevVA4Qvtnk5mOh12thJL7D5xTYogTzydbm2GZXX/tlQ
mj+lqkn8+BIgllM7f+374cFmnjBP9KJiK1kxOkP10m9k5LlbFj8ROGVANgmQ
+ayIS4AY2YdDG8yI++qJtRmkLmvhj8wfFlYe6wxsROlujxP14raaqKr7xF1N
fDudpbPPYo6CCDvNf2kIki/pA3eyYEaeTBBS7ytTViDXMrbaF0g+oLeL9PuU
3He5YiY0uFQdFSMoRVZO2YjEcmO/+dzEcuJOUDHiJ0nVI7EstyqswzfJM14l
nnwXLxfNgxBT1DCSiagkjn4UdNFDepf/2NQfq+1Y0Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m8AcjcDDgpM3KGqj49hAnnjaUWsrsS0hQDk9maF5mamYSEfI028UG7goFMz/
6qMH/PcUay7HQQgXEqO6tgOVmDv51phdH+NvkCTFO+essQiUaxEK26vaqNF5
1yBrbji90tzIV4VOl8mnXq/cbW5uxdYkLurRrv91pPliozq9bHi028yLUj0p
1RcSYt6FJLJePUdGlD6ROCGFY+XgKCj7hZx0HvpPVhFHOFfuODO1eJa84YQI
i06kaSGaVeaDRhPadU6CN14Krzir4Ki9Xb4G1mq3Mz/n5BqFRWLEPPXHWLCh
DF1x2hddi9a+tb4pGwFlZXyNbotgLTeJ4IDN9uvjQg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nxkjyhPbKkPIcJ69hdXjKZhj60SJD0mGYpsDeLdwKNt/X4Q4TnEOOMo383LJ
07EG6SBD6DOUJNtnULmupSyz7HNaa9M12ohDzmiLIeIGBBYZo5dy1I7KMast
idIsrF++EuLSrSyJAAI9NY1sVeHLuxFqQX/PMMMe+ylpI08Y6/zgYDmWEkjk
4kFKkXMSHblUUESq40D5RtSUYxmuyzsxTkRqLRl3p9iZPplFraJDlDAysYd1
3YYHOiZLsmSVXGC/TJOcz9hsfNwF0Xh1FOdbZmDXTYnzlzGB7BHycdxv4g7P
ZpQ/CTV5vCSOFr/LneAwl4/qfyYDn6KDVcBJhwykaw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hDw7NSpGITTgm8qSMCDze5NtqZXVvB9Kpxk648YMsHrd2eoI62iPdbGpkUjG
kyx8s1hXZDWGJE3vuqCb7UlxsaHNkbAQFhk3hFtNcFg5MNX7sIEQl9hlxyGr
sByOAo33c1qvBSO3Bqs0yrcIME5Bvta89hw43xKf6/mCJxbrVcNmy7Q0/mBL
3ZtrqnRUqvIF0mCMTGrsWoBLHwMCPw8sGhddm5OeIlXo04/yP7yzxeRkjd7W
0thBUaUn7A39805xDd6OOamiJsjbYkKVwJLoLU5rHrYi8g84C7W+tiWInwgY
GfQy1DL3q/rtHlpVLLLer8MEx0dxt+ehYnoLFmp06g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hhgVrlqZNcXs7Xf1uZl1tmWkeCpTR1XiikVcFFsUmX0YXGKZaP2RtaRsyObz
cbZaJT1SS01y8mB24s61hDyi2LKjSAfUY1YDLXXN4+ZHqcjpcNRSfwV3qcci
ljiZdoN9Z5sB1XsW98F/Xy9aTqrlbKcCQYKbFbxXA7vF0LnuO3c=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
tOlSN/UqsgLjLQkz2l+uB1DeJGApTRDe/2ndPK/D9nX9eVUlQ31NgSMBKfRa
3REOqRWgTTJfc3LFkBECFcXOJOFF0pl7KujGYwtwmvN+0ewPrOGt1ONRnpct
QIV3A/OJoZ5rG58z8nC4Ml+DxBi891gTIZL+sseK4MOwmsPxnwHeYPyZVxIn
fAdFaJwYcLH4yxbVxbLj0vk4e7Jra2HZRB7GrRcjDyh7Z3aKwQLcM42TzJAP
9N4xqvZqmf6kqJyLi8mcakRW0AZmi954PAb9oLbaNQ+TPCaUOZPnCsiXPvVv
u8IWDutrYlaAseIfXBKxpdGczaJj2BtkUO2cc0nODp8HVRA3sDeULGhlY+fk
8kmYjonNggPbk20ZPgYWCYHa1TfF36Yfyl3AXaS6PL1/puE+lsUXepFZaCG2
exPZmJhh07XVEh3ZtAUcBbLT5fDVk4/HHgCnv3ITH2jlTfYgauLHXiJ6LOY9
tbQM/aW3Byubpm59+KecETYk+J8RfPc1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZiTTiMA7ZUasnWhmcRVvNOpj/RjIMfd0JcDJA7oHX8nA2F64QrfiYt3XYCak
r91PoapyMeJB9FlELQIQak/kbSuYYoEneATsL/AAgfaR2NqSaAtO8xE6e4bf
WR81fTRgV7a3Xkwh3cTkSSC5joskWQkgMo/uG8Ox8gbWVcbPUwI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H0cclL7knaXUAbh5KWJOPd6cmly16VrNddMEs9Fmr83/TDxCw68GCbP/KBGq
z1peVvorc0EtpweYHit1MlnhyPc/tiDhV8S7/nL/iCQju4+7MqYZKbCYKPy5
fw5ZfqNDlxCRMCWrTtbzP3PQ4ApQaXstgejHfRn+YpCrXFv6iFY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21072)
`pragma protect data_block
ITuFQXsQ9MFgDxadMIpXMwxBwOTCdXe28bkzRDThkjHmWAnSpGpBjySwOLg5
uABLu75ggotQlu1K3uEHq+AQ0WKa0Z+DO/9blIyfhrS3ck0vGYWa1PhZU7ZO
VPmN7YQRSX/YAZtBA+2iYpKdgNyS2e5Vm0TK6co19sM9tj2zSweHBJ5SYZq8
ZaNK5MjT2z9tKHQTj8jZZrF5VaPj+v7m1ktVdziDSI19bTdGLqwSPiYZUc+I
7YPrS3iM4ipGba04trQBMd1EjJD3V/3l28mG5vA8TB/2s6wWVsTm9bC+XZ6Q
HyGw0+VHyH+rh9KL/1LcELqlYonN7IQBmCah2Y+qU6Rn8yw9yNcK4ir2+kKO
ZC6cozHZznHvY76RuLOb23QHRRPNfaJpGPsKo3Z0n31RtepSZshM4W0bswwL
cKdfhtcs4b8dr+fyZR+ZWGr+99QkEj/ytEVOnIIwyJhZ1Ukf5ZUhJRZTblO0
GFOOppjRI/Zeljl1JzAUQ5udYusYN9QAh3hgoDRD1S1q+vwsmLxcRvOhwalA
DeeFuhXDrZTQN3ORwRPDzu//d1LH7RbSSvBvNQaAIS4ugNbQ4zeHrKsOmDa1
IwxbzeBBMu5Vp+ke2cTQhTQxFOd6+fbekfMJRp5YJviZfuXhAlhmRkyDPiKB
5lQTTz29DWlhM1mnJ+BfbVEpytk2CXkKdi1ICYvqTFdj3XPXYf2xyBRg/RaZ
OgddK36qbNrBGFfOKw1cgfyF1Zk3SjctI4CeFPPTKDQSHBlmfgdjTftXwa7p
Npoc5U6/1IDqfyuXyeciTY8B9j9ifQ4l40RvYkzTYq5XVLMj4oAQLlSfrypZ
MBChYRL0mwpoN5scffgfX/3AxtE0+CSvmKPWgRooH9E78XZUYwRVU10DRhOH
WQ+Qkv8t5WcLIb5sa3C98yQodutCpO6HVplgwvlZt2NHHD6oEShvaLigaLDL
kC0CZbchVupi97cxIPxILNfV5JOgAZByeAAAEelI1LR+XoYkPObD5bBvECfL
aXCG0K/JRJtf/ZvRvB7irZKOZ5IhhtrWpncCv6qwlsHyEHn2AbcgB8dZ2fou
TjtTyFUYPopmzrOYT1RoS17UUxSE2yY5mdy4sBUC8WP9NgvAT6TfC1QKvE5R
Lzpt81KgYHSYx+CJYXwCMvaQpfGxTrbAwPxc1FY1kc0As7CiDAIb4Ad/n+sx
/f3gbHsblF8UrmoELYBsue9F7UT3wgScUWCdVk0XKJ54Lv2s20J8HRtxzQT8
RImd389dnhO5JJyB7VcqquJ8g3a/I6MphCy5C8x78cn5TVHfuCvVOCXOYMk+
vHR69h97ZF5kFXFEYoGzCiWoyCiK1GS6G3VOlfN+Gfc3N63jz+2NF6qCd3Nh
SR7zM4jmGh1nslpoKuWtv97Khxm6a6+ieXYMRpENHmi6cnvIJEbKGLS6VtXm
PkvwvxX7OtC88gYrs4oCn3C/x+3CpFogKU+ggFoK+RhiBThgajKDDCajcsUk
6jZZ02o7WNP759qiciQ+5MsI/jLaCAAL7ak6yjYllnOLLFBIRTGKdrp64g2E
ypYF9g6Kagcz38SLbz+FK5lN2L7Uv+OwKE9fAdfiwqlumEFdiox1shLx9N9M
Hor/M5xZADQIo6x92yiyZ/Xw4huCKw9TcPRy9kfKvDeKeEqBHNTSE6ZeClWJ
KA8SdkLuXvyE0YTUk6cy45dtmhn3WVM3jjIjwIRA7vWCnFDZSSxPZaSE1gRh
OOSsmSKZLwT9wDaWEtT1Y5gG3ne9zrY05DbIvI426VBdQB89eXNwNVUrqEzp
cJqRRsW11fR4q32cJ3FvERoObhdJn3ETotk4Q1ftcQWJiYMybceVAcv6Ui8E
gHyHnlIJlU1tbmqnm4WKp7Og/pkl9CYRn3worG3toTc02K/2OFhpo5Pb9Xlh
GYpcYLGuM7emPnC9ZQB+qdOFq2rkxcV+xrTW4bSaX/mRacMx3aEcHfWOHlCc
gtXOqovsiyoxBMItPQh64Gw+73XBmvSBMEyTOpKdv6W4y/wJepeoEmpLjae3
DZ/XFM3Q/UfAX71lxbZngkw06ttLaaw4KmhzCLu8jFMVfmLwT5hwl+88uYfz
EUaBrlcq12DREJ6Cd8LY8CW2s3y0sw0I26qpKJh6U1XUqa+7RFlXuaJ/5Wdi
GZ4bKIVZhzwfrxczsDYui836WrTEEhTYzu6R7v6+TUVt2fuQRaGHt5WFi2/P
JAkLpUmx64mjoKQHOWKmQCR7dAXP/4HIDRFVvZYiC00JTKM6bGMeMa55lKdf
mL1yhI6gFh8ITS9r/1klH3YJsoVXvV6C7fSm6F+vGFIrKVGPVXO6smUQFNal
ETXS8+qSS4enWXOejbef52C+aUgaBwe5zlFTRcTiOLuNyU0PIy1iUCtvjet/
waNVo9WQyascrlDhYepXmL0E3rlbP62g1pyG9TwOXetTZy8gIwSij3FlJC6I
5cIj1+JCpmwzqw+xWxnyeaIxuceS/d/Suq2tBownCdtRXGckmju8MrKxDGqH
RNmmoBr9r6Vrsk13X3cK1XR0/y5nxt+ud1J6TAZ1pCs8Z7HuTMSLuHWtGQC8
nKFNgZTI8J5eLieuTJn4LQC1SVahQHJq2Ju3zg5tXgTzGxNuuP+7Q2UFJPGb
wyR1iX66o0S37Ob4mN5qAuNv7yBKmDGWgsXxd5ridA791ABrmYEA0/vdbZjV
J2IWJcGYOwXC60ql2Ym84nWIztNUPuHr74+c48Cu2onUx6+JETSsc6cVyV46
yhEE2K0ailXEDb84PMu4CgQ80e5IssG7+lbys1JbHOhE2RLlfHqoLmbw82k7
PL2TNSCqTU32StW3u4/AzrRK6ly1LxQ1ZzTR7S6Lo8Yt50+omUPxl0W2W4Z3
ZSWwCxItYtcruewrXRLZ41CK6kVzTolOuRdtNyilT5TEp1Lwf0wOlrvlPAnO
FmX85wbXb2Qr6g3A619TsEo+ej8754P7HX/dDGosLO46oPgu/L13djI/bEb+
j2SPaKqJzNJ0ik8mR+ccv3hJUZVPUb/gvOMzHsaZJom2AnjCu3ePrx30liKQ
FAC125ZM7E4XT3JGpAbfFRLhjhjAqQzLGz3HLBMNRjWI4mT0Nws27cFaWiUp
yDvclQnZuEFI+8YL3eKxhT67gmk/XQKMpBRvhhqHK/hCY2F9OkjaieZzVQ3z
afRJbuncWl6esAetuNzKvfxtGyRgoDYIEAD3WR7PKsf4wWlhjoQSALPaAPtJ
Ba3NJ59zikN6oneOiO8Ms+qC3MTIEiSIqC2xI7MLNFIUvjMTK7IfKJl8rpni
1zcYOqHjQBenlfIlbPJnUjGYEvR5dGK/6M7WOmxMP+Yca/ttmlc2pab7BJoI
g8UwVBkXW3WCG3Al4EKzT+JeBiG7z6kmK/CIxOPz+BsOaX7xkfJJ6p2b1r7R
HHhnJU+4IOIMkkLlRs+waAENkGoO/3ZfJ1ZQopymQ12Hb0TlRK7rnBfAng/U
AREg5mnldzrAV4hwgBmE+YX+dbtzONmmndndzDypVv8OQQv5yaUA9uGGSuo+
FJPSjjO1qgv1YB8HUW7zj2k+StlK52w85ISgMOOWZt+YEzC7snq+3OsyJgrD
682i6sVN42qAMZdjJcc1sckKqa3na57uWZRmFpmuEMNTZABZAj4VjZeQnoOL
V+tiloEP7QFnJUAqct8jPXew1sW9LLhiQuUCKoDBkNZfmO33tTaR5xCpNFsn
/ql/HQmUpI/WhlfoUUlV/rUsiS+Lfhb62dbWfi7nPGJs5NvwAt9PUDbaHJp7
zL5KxyN3KLGLDqQplwwvPWBnlhpGRi5V3y8UaWhFUbakG3otCwyXJOPOxZa/
KHE5RBbtBhXAbV6D91Y+WoK3qgsHs2+UhZPe3N3FuVHetjExcH52KJKqPlbr
5dB9oOgM0qPCX5UF7ZBdyOlXSN4C3FRXKWC3vgyBhWB1c9gvILqIOZ/TdDtg
MWr/N8haVJwEn2cG1AEmuxbpahkc9TbwdZKzANHRTZtQSw8DgBEemi2Z6kwG
wXIw3HHudVrCTthbWmqzWNkILpNcBF/N9JyHcsj4I/TWCAi/xgT2D0vvIkkn
BIGFllG2LURK/5TqsMtpAEeJI4BfXwnda/RXFq3HyhWl7fRsm4mWWwv5mTK3
OCze15j1rWptpGG0LIDeLscSvSGGbFckvwQwYE53KTHYPFbS3cnhR36swiD9
zGce1jgdmjq/HWBdgOD2hiNVi7PUqAzJtazXiiKoE/F1ZQ5NHKpaq7EtdGru
LU5P21IWdRnY4i9Z4Su0I1W7mxUmzaWA9kyWrnrWWVjrZHmd3OEtHZEoNGk8
UJ/yvYQtotBNv5kYYsvRCC0yu/8FJ2EqbCU+itxatjNIeCczkIgWkkLNk9Q2
0C72MbxwrRfE4o6TVK6otYjY0IYwl9W2/uatmbjKUqtIKmCdaEcLm84hOhuM
xCKBKguaMDy4ZkBG+J9nHoDrqEPcgRlY0MguMo/bDFYq3D3kf0NA0/64UVOO
tOjEtvjTZ96asur6LjmmrmNANzfwb7N+Dp1HVSW5T/4oh5bFgrhOFkJD/vPy
CWrERtX+VBY9lFl4tBlsZe/G0UNxpig+5NLzt7RvWQvr2bDP3JHUBguZ1kDL
QIQu9TMj8Sk/G1dn2uKROOVK2E51pGZdTXoTiXceXxAulZ+EPUoBAlbOKa/S
c7TxtCJnV5WY9NOMnsObKTHlf2RwS74giD6w8ne4JxqNKmBTgDxbxfOBDvL5
4MBeM4P5qCOYWGq+Uns8BthJ6oZmj91KRTvNeLuFGwceAoidVT2hTctF4Zig
YWozCqgwfzZYG8plxqFenPMchg9E0c2uI5+UwgIgl4Ih05qTCwVgpEJe9nFX
8AuHG3HuMtUpudhFzxW1vaesKUzaqihN5SROkke5tpsjuIiSZFVEAGzC+4Zv
MGKi/ScU6f+nb5Z/8Ml9MigJHZBotYSiHa86LKPfN0Ps7/P9Yx30SY5j+4AM
JrTmwAwkobVhWdqhx854ohQoXsd+kC6a2rebeddw6Vkf1K0kR4yI8w8SMnho
S4C5KP7UhjsBmooo7igMSw6OzUfP4pOS/CfDJl+p+WBZeLQNBg30vJ5OB4WL
C7whRdJj6pRsUcI7zQ/a6NRsDq/eVye1VRiGjSoDdrwqHebuDo/TV7By14Us
FNs0MRC0o+kMIdtWxYCyXHO72EgRWvppAFenQvYMjHmhus5tBDsFfWo6Mvhq
5FFFs+PLxk5GdvSFNiE7sS1OMHwKy8oggF9LXhMOPsnFWqfZSS2+J7MFP7xd
x6VoiNAI4SR8wXXApshgYb/xCeccrWwEgb8qHMNW69YUVHMZMp0MesQnRLte
4bjdh58fuKvMWaHq45b5KXv/fMUD9gKRg7sv2whsBl6tA1PEyZrjcdBhONTo
n4VJ+JYvGqHIFNmJwqN/slST7LuNDU0JCDlOh8aW9lMNRPNp9oPsbd5BR4jS
uIGPhPxzaXvBCfmha23TCfnNC5mjGy6dFN3ZlqdA8li9KVPACvu+aRnbGd0P
zfNH6frQNkBOiTu2yoXHryCiaG4jiby7CWIymviS+m/qsGnqtg7Opwid33Pi
jx66f2IxkN3d8Dw0aDAjv3k+wc9+YSZcGqwVRsH2wiEd7YvKa34LUqQ+0mwM
Yoh8VLHmSQzU10QI2c2+/3gaqxSPbBM3dSzzItFGAglC0EJap6agm4BwXKCh
1Xa/UKRM2hyzfuD2cZSVZ4X8UG6gV8m379OLCQgW1pZplSNxEJPbG5OlxdkU
GUtgoyfIpQEVndbxTePMuc+2buwYrZWIhzkpbPMkfuFP6ftGwWjc4Mxa+UcG
An6lja4q9eE2tUseLrH1xa9WgfGskVTzzxGF7U9jg0sntNR16U8Y1eyK9bAI
ZcEH5sl9mADkhu9yTDeagFBsyaZvzrVotToup0KL8D/CZYHA0XV4rrGG+eEi
+lJp0nmryJoLfnd7wyab+dW9JX3VX6NWXyjHsjoEqt8Of2ChoF297SESspdJ
C/1A4CjMu1XOt92xSXQzkBPP7uSBzinPCyQl1uWpttBwYUmKmR+L9vlRh8xT
gTx3AZBOPpqi91Tt9PhQ2tdMgiY1wMTVH52YR6Oy6xNjVWjC96RVBKIQ45WY
7bQqKLKpSuh8ji8VA0DBO3zINZ8Aj2wP6GDQqyKRRZbWmlilu4eeavnTSkMC
UYGrD9qwDtlbNq2FlX0HrSYLsWmYTsa4iAU+HAGLBfuzCmFoq7U9pg7I/wmZ
XnYp4QAq2d5nxyo0h1YIGU5+snHUWj9iweB9yBX8zeFZt1uyPvKqLdVT8eKH
1GcbdmDiQlyYwRQMGuk3V5IL6vqZUvzp1x1Tn0FaDtpGmRFCH0nk3n4P6uMw
yRJKMz5vhDXUaaAU3KqvJvEI1EsxJMloKEhg6DqwmHvj1xT39NV3uNCeinCZ
ute7RAcg4/yMF2BWR98MZHmOneHzVq63dzLCdC+odSr2kX9P6sDRVImZMBi3
ImIJlCno1XTfXTKF7Clqr3DxWdmukamZhea4hdTHQ+R8jwqt34qysw7ZsFyv
BvEwzYzNXKBHMivdngfQIaRxq52iS4FhuL8JnaRODGC/iFf+voeBml8Gs0st
UX4h4EhcTYoOCdN7hI3+6t7nWseooBEIkzBAEMuM0jJXO0FFTup3fH5Ezw6N
eBQceOZL7XUqoWGzl8dX+xr2rj6ji2O3I1IkPqIY7aKp6/ESGlJh3Fn8MeWX
TyFCKgYhu0mIeqHiJJfNuSr5w30n9FSSpX3PCM8j1Lgp3NVp83SQmWINrJ6Z
jgkjCmNGqgwRZs777B7dWeC4auKkvBUHBrp/P1/RPqa/vARxc3HPPa894Kl3
AMkvOZ4cPW2gsTkuD2X4h+WCNspfFqgd57GN3THEU5s3l0biVXkEjFJlgTS+
mAvzpXNUoBJ3Qu2h7OudFUrPsZmxLl3FUvAC8ytPGIMF4gGGS+45SFwUij4B
xprzG224bFCoMZvsvcdtEhWbcEo63ViLR2NBgOmL8yBqiHXGrO/5186ybK4Q
Y0I8R8fVtFKCCm1PFXRTeJR5ItElwZryT5b9IQwdA9sHEMDsAxZ+E5xo9Vgr
/3qaAImpKjXatnpJ32Zg5Iln07dX5MDTgXXDWu6hIOtQ+f69wIsTOMTl7sTc
1ER/qk9/BdYPtJur4JcnBJGbwPmBzReTRxdbikHluiKVp6euJqENPoa4ODFF
sw/gqFP2clLM1wBso9EqFvnkGHb6s5hyIxsnSx9i+qNla/7YxMOaPilEUa5/
xHoWquKc6QGAkggonUX+CdafH9tVPvldCZnuo7dvHdGyVykAY3hZRQQc1s83
JCGjwuYPemQ25QW4jL8DJ3Cei0oEhrwiA2/BjTT2U5+wU98jk9cjv0YQpcpE
a5TRVNkczVJiMMYXZyT9XBqUV5szU2d/s0C87GOXkpLBNh7tvGCyeHQFSHcn
0Jf22pqtR0dTGOftrkcGbd4dfijM1p2HOxWIth63PrR6SRJZnATEn4wYGsPr
LyipECFdU6505pmrFzddM2lSyY8JatsOqqnRAEoBOuC+pFSfaEo7WG29oIbG
UU4dLWAl9eLEk5g3MLpSDbqfIglBl4UiSQNeZ5Y5IyB8IrffywJq6z7/Gw9k
mQcWrb1ugRaW6VWhFtyNsYWPzFR1k62pkbFhddrDisUFZlHa/smlC2R6SOs+
9T2v9fJzLTptqZ42zS44Oee+RzlnGeX1Gu5tGahE218pHkkN316KV/oW7h5s
ax86VCDbNyeu+JDx0ebasyKVOE3qHeF4rcxZNkSFflPvpexIW4YUUrN2gQ+D
kr7eS2DWVclQ5iV3mzL8M6L8+MIUDXDFIfm/E4gOFkbkHaNrlURF4h6wfOWl
O25Vet7z19/OoWGw67ujFBfhmG0Qqgfg2LBwoUT7EpFdIv9z0llbJET6lv+X
W75dYPgSOnumxp0XeaLWVqXDhciMUnpUX6gkJ7itk3Q7Xc1uOLtUdZTJG0lM
NI6+zKpdppKoWIF2amvC0DnxMXqOy8XLtZDCx8yOdMNtExPOFyaUxyiGVbSK
RlnxYK8+hjbwnwYvK2E8mYpY+8MvDnch386APdaX/81UGgxBw3rZyPvMBBGL
D6XRnjt/qh0TVACSeSoGfr6odiyLKZxC4r9AZZcrOo4e+OfROY7XUxBZDQ5y
oD8wfW/VjmsRvHUrb/wSbpVhfxSHN38bCuTFwoWq+fc8EFAJQKhCVdT4KDyX
1xUzdXZUHpztZ0X02uRrkHpqiv52wJea+6VQ89OaMeYJRnfE4wIjAcJqk+lV
7q/EedBq9DNL7qQhoLXysOvji7otoqrfz9xQvX7Y5DMGnjkwp9KbxolG+x0R
HDnDzhCua/SBmCZ6dnKe3Kkql/CyhT3OnDt6m88OYqlf0Lmfpj5MD3Jaw7B5
paw7A/xTmP+EDehM3kC3OPMzZ/9RXtTrvh7nw0Dm0f+DEJQETcJQqovAbqLC
JfEb3AyR17+K2c6SmqynzHc9mRQCJO3A4EY3EuLg2RxAPkE1bJsck6ilmJpM
MElQK3BgTuehefhqYUxWtCndDLsin7HIfGZf/CpuW0mDFlfnmo/Je2HmKKCV
7V4pVgtzztag6CPWAwlwh9Okn+3t1+geT+r10ZtVFQPvDgkicCzXhcaxGNPR
arVbs8kk25ROV7p48kBT0XtlE0YhRe/SG8aovP/5unDIgFq9+5208p58q+i4
C5/TYVZBJwdMUkyPpTmvL4siuVHohRYdweBcWxa6xagFP/MgxT/0Khrn7xKl
eIoQ/hKM+H8vXAdOfVtKeXbixd+h9PyJ1AFNSE5KMkdh89gvv7jkk59sRV1/
aijbgm0A/XQXU6Pk4plb0PIO98lcDYGdqNJP/S0U8sJ3Lj4FnEGt7ghvfKed
S704ggkvl0Xkpqs5FSRpkJP25/zUE/KFh5GS6bY6hXq+8FJ0XAUbsWWN3/74
vXUwSWaDrawmz31RJeNqvPvQxNp12Ub80LxwNyHSOQPPzkPDWmLo7Jol9daK
1jDNG9PZXR6O8rp562VrfbIvjnZsEbAweva2Ftv33Xi0exQprmDAVUEmpp0F
VO7oM1CNf/Ylk1oSmkWqRiBqsXdBfKBuF/6TW3pTNJU2HCWqsSoKcNi/78AN
pu+apX7Yr/r7SCU/36ByWkVTZbBIOAopChLeyZOGw696z/020QFV6q4ukQeB
LcG72DHScyrUAAXbAbqf8ptmz5N/aoHjJ0dxfS4to0Ytu75mkUTvvDbhVzPj
9/4wIptZrESoX1EoUIt/PGfCq2+ct3PY44uOHwd3fla622ri8LKd/ffgyTtD
gb+yqIigEvr8skvp7u1L80EA3MjYBSSvjTT4it+AMpar/KTzQojuqaObqa3y
98Y53bUYMkfjNntR5Y98h71mxvdkvgsvPosHV5SFVDOto326sNoWiiXPNclX
ZVwfiZiyG+UqCK4HmK/p5lUdUAihhzUDEmgppDXK4/2u6PPqGhd7BtO3ZVNt
U+CkitfLZbBsUlXLgcWhAgfOoQnhacE/loh3K3UbWZlFzrS8H7mHzxX2RkPw
x/bmmvcX7CFpI1NXI5skbPnDkbniKrOlJcsQ+d74WgTgAhrG+smCGUXoBIos
5tvZ0cZclA0da9U3abl8UNIVR1zezfcp/36ZFWBj8QBA0vwQDFoBqPqi7ShN
IiRe2lpdG4Ra70OkD/CGXasKiOWClaRBgMsLq0zHPxXbf6ezXSmocT5k4ye6
c8c6Js1p7ktNDLz80UWTXQnfBUN4srjzJd9lzDP5Etnj+CEFasJCti+rcTam
qtHiVsH06Mju5I8vYG/WaiG2xvzHdCfyzgqf9lNoKwTGhK4rLoYo4CguoCm2
AO8sqABd8PMR5hx8rsO/pdEbZgPuXuD7aSWif5yjkRvK8kl5V346c74HsNQL
81rhgxvrdJpS2JzqC4tEbERiikbwd7xjxIioaC2YxpXmbpr+L36pqbqXgTvI
r+hRxjrQ5IvWloG3OBuRA+BGMyXmGHD3DaIZSZMn99knaNze6xl3YRFYKX/4
ujJCNDY62C/RHCf5zD7DeFu4eBpaRMvfDhrVQJFscVq9jUpfp36UDJM8jN5G
cklHIRSNtMSt4G/V7uzhlVAzT/hh1e6w/idbD9QzF1vCKkg2Mm2k+e113XHr
01BplQ2rZBNxQEN61+58MHOjP3rm8XiYy1Byqbj4mBFugYuWe7hiRE1oFH5Y
bS56T88Z4kVjKaQJTbT5DGr47xg5YLUbjYNiDYy++XwH/wfq1DK3s0u3Bq4u
BZHlU8J38PC+5eT9I2cIshOJ2/jLaSlyE1z2w3gzWfaMc25k0dE8+t/+DDAv
aZChbLpLO6KSZbz2GcMTORmNkpv70Sd3hRcMz5+J80yHIpQifAfEosDq78ov
yJKd6CqdH7z9d2boq4MrspKsTlhmvyaXubn2qo/cQxpD+C5Z+EY/Akesp0q+
NRp+EJCs7ho9eU3Buu4kj4D7MGLK76q/R6WHKnxJAxpSTO8Qd3ddbX5uAE+C
A8R3OVhrvjij8SYEHv2Au9eW/LdwGOuzs6po9+wg6cVrGtVZUii8fU/6AN48
EjIQwLZRUmulXPIdpRNF+9WOJh+pwsZme478PiHrwMHtVSnSUKHv9OTUea7B
OS5luC0F0TXKYlG8zVJMHXOIRuI/Qoo0V0PiRjSRYUyNglbcAxj4O4bQUTzD
yFPsE56KLInwGMoo5qGlrBSc4W57iw1gSTpc1h4/rjBVJs3cYRQ0ebV/ajNj
Wlwfej/KwrbcTsu0GF0foLJ2r26ZPBeqfIPzSmpoHsNPWQzanem9+AEV0uRM
k3F36gOeBvf64cpRlAtzjkdoLpPv+IbjvCJ4JVLmHax+Xf5SlcrE+RkGJinF
4mMGr6qzs+QqppZqb0BQa6LKIk683H22VeSnCpPxGvfESRsiR0E94TP7De/J
C9vV/TtncxdF77YTeOp7M8ZgNygZwRCuPiIh5cPCtDze2ojsVAchsZGGfnbk
wPrZRlfPyBvoN5RoOChRDFaLgq109ZKyYsyeKto/DSTx8yc27VzW/t7rOzi/
xl+jFHeVAuWZ11XhkeFc1r2arLPrs+7bwbLB34WwgfGnUwky2KMn7txBu5e+
oEXQHz2CO6LgMld2rkS/mkwST2/PhAJqR0cmeZJU6ZElBrnq60Zak4xjVheq
zY/+0EX4U8JAB39sEMwtupJyiraxczEzsJ0dXq8GXZ7rzzo/UiERZwTIslzD
bKKovCJkuc9DVUJ6h8mz/d442xTNT2QklbJV+0ZfwgviRJv8ZM75UylvSsde
5+rUpo/76qvxHzRkSf/AJ3wD1Q2K5t/1a8HOJIRWMa2HkojHMY7CcoNSYceV
ORsUmoyIKdj+qHGsYv0CEcSOgn47cYLS9RU2BN9V0tjzTqDk4yQV6kggWtCM
laxtwAwesrU4U5i5OLIYSetK1guPi0u5QCvZTVy6AKZXCZJkztHG16DiqIXL
30tNvqBRDe76K2hkcmuaKgODeTNWCvMfbkOqvbDRRzzUD634GWz5V/NKoFs4
Cu7bluhDFnqOwceOv/8zJQRgjmc8+A2dyrRHWZfcf+CTmu1Rvk37KNxElNCj
+nNOFPMRUUgoT5iJ71kSH9LDFPgOEH1lKT3e1Wz+KhiLHxHsQwHKxqg8S9dk
fkz5JtLl6rEaPux32B0F4iw9VojjJJ8+X5LvrThZ45AFElvCmK55hrkx7eCx
6Qq+1SQqyniJtc8nzjWqrGwB4jy+8jeRzWuegk+GWVz9H3vWBdrvykrVUWyS
iEa/iLNw2SOE0OWxOkJWbuKlxtF35Ko/LikNz07r3J7gtiBRcgUqq4Ejt/54
NqX5ady0eiikxliUTFmDHR26DxpQbQjBsc2e0ispYchOqc1YZbc245h3s2/s
rPh6+jMnH29QQZ2gLstZl5kEnIpFn2SV/UTCxInpmVvKtsEV4xZ0zL5WKj4X
X4dR7OiQb0nms2Uw5JmJbcSGTzMNZ5w976sFvGz8UuSYzQPURg0J5wjj3tqK
Q+XiDd2z/pPqBysv0JmvCnVvtnrW/PRkp9Y1Q+JW8RQTWCTeV0gzNwENJ1Yf
sIpBVTDv6RwggjyQA4stifadCi1N66FjgaKGCrict+NI9ycvOesPpdYuZty5
H9cdXdE4Q74+/hYJP+Uekpkk4ZNeNOjzhp5hoNTphw1y80VZjUkmmmYL/iVB
Q2aOv13zQbrmSwFVosP9kypAhfB+LZtTggbai7PC9Z0YkiokkrUlo+fYWGyy
xcBi88YZfKL/o0xHkBzJTFjDKqg69YUsGx9JCDTWvuSYTUAClpXaovxgKR6M
3YRdYaxQLlo+JP7A6uotOyE0+9YORXrmw1HGEFMEUjm8w1ie8/fI2pNq4GAV
/faUXhWi3dB/VQ5nDLlBAABF4NQXq27YCyryYK+Qm1GFi0ec5w7PoyAQYvnW
T1iW/tbvJMtJd4Xjstx7yxSV//FjINCoYkKMNXcWarfqc5C9WaKXWG8K1s3B
vTKMK+Ko2qvvrIOaJLKR7+lD4iMqSTtrEsZZdmcGbTaBvymEWXY1DLRyohZe
DrDxd1rGMUmMLW0GRyV+R/x2X8QGWh230UOxc9gQ/PKz82YPrpRRKp8SKLk2
NrOjiZRSTiiLUIowL8dn7WFr4fQ61IukPaso9Fzxg1r93xUqXp1UQR8+Uf6x
WOW+yiivQ8df46Jt3FJ78LIwSaOX1/0tjDqG8BzpFfhWyArJqXHAP7KPXOTH
h72NxQCK4DKQmNgIcJvl1o0Ayk6fH9LpyuIuSIuOtHcCoL+Xxh4FLzC4p0x+
ui6+G1RLDT6a8oKV7MnCuEe8fqKEG8n+pvrrmF4lV/E6Xg3+gQ9pb6nsiYbf
OFfHx1rJJfqDZ1JjxxvSi6ebD/7AYyW1FmK9c2NaE3IkcRCS1qt/CpEt9LOB
/UKBzRg/XYReax3p+EAh0hYMdKbfGBVJZJ19e9devpgmpKpg4eGhPY4NHd8w
qstZYpjflLL4Y4fye0oZ1Uyes8kmWYHRNbzfTp76JMMyAZZMsAfUmDR6BbGD
e4F2UDpjSioesmK1aRlSZNtnC20RDsTDRlM+NSv10JIhwJKIjsONLPuDiRNM
P3/mZmRVKXdyRjsABgpr0ojbAOUn8EKa5KmVTIy1AUrKO7d35WbcPUfnQcwa
/uJ1aFZPeY/GQLuhCuVnnpQY/9GOP+p0dlvefMMWzcBJkTAvFnwyMeK4vLqD
yrUjVYmxEtN0yKMDBnbrpd/Ef2PQ7DnTjU0FEDY1k33UySmA06JB/SH1eQ1o
C+pvqIS0iY5VgoicpuUZXOyL0ypOboVaiojrxhxwAt8m3/cCMkijuBm9nGbh
KF8/eDhFwzHzTcV1qZyet4vsLT5roCQapMQD28l3o/+T5NWmuK6ppSzbj1yJ
yIWNkcW2yAFjQEIsWusgQl2dUT8i9pXlPIsWCVRZC/kTkTPqEyjeWXeV7jMh
bRj8TmDiMDFpE9X4N0tTOCyi7tkWk694uLvBPdT+9sOQgHAtpYSccxc4a8OK
IcRoP3PyywMfZIh3EcHcgeoK1OlZiKqH++ySL2ggcS5SfKKNI41e3WxuzAG4
P1s8Clt3/pQZFxm3rvh5+LiksA+OEJ0PQD0W0PqMLyrCnDbKxp+NFQn9ilAV
rgj6eL+H1/8AyTd1WDFLiSTGRBjJuo4Uih3nyW/jTXNFgxgSV1oiqBeOMKKi
JGu5a5fcJHgfk56KvVvfCz+b0UtkQZlsceuM+CoDPI3pzVlE4lks3jf5vSIv
B6doLJKvvBy99BeLaG1iD2cDG42XQaNpAhsQ12feaM8CQigBjUY1SYu5AC15
3De+4H3+lajSBsJAlPzPKCBocayt12sCpUyec8Aiv5otkXPlSZFWDEiOoJKW
x9GQGWi3y3ssVd9imIgNiCgxcs5hFhyjtVgHYp5wMlyksvX3PQNpZfbLqWxz
3FcVqRWT/A+umyhaI6HHPijIEG7dsKtHCc/7xby4sfNKVZB4wtZ/u7XrIiYk
l56G/o5cJc3zv2XMVPb2qGvFrbUH4DJIDuJqBuSTSY1EF2iWy2UJMYTa6ZJf
LzNr0Ubm1fw+y9a2mc1o/KXZY4pl5ybQO07TwMwWR1i+6Od2zlA95/Z3B9Q8
4OneqKpVxa4+bXxh/YnO/4aqI+GX8oagGFV/YotWl0dDM2kBVKdNY0viV8FT
qVSTr+DF6elDSK1OIIjGCGGNpivwpEePoDP0CcIwZpROivENlrqgE6boSk12
zhBiQ4N9gPtsVoVcsVUMFI+2ve8qptZ9jPBR0QWgTHiG03zViX1nTASRSvCV
b/Lk6L03DUbS2qAA6NAl1LlXXWKX6INHS6D9M2Ny6bb5slhperCnPHBUSxNU
zDUbIda22pbUyyeq9/l2kNE8BLyexwJW3Q0NUyL3HmKFInaWcmeRB7VGaER7
IBvMgpGKcobLbSTbUflK0YuzktNJXS5cNa5wToBhXX+QsRCORA7xFXU0s/hI
O6cmgsGESG0HWgthDEp94HDVaGeKQ749umfJnlmD0+E3bribuUC9nztzXXLe
37u6At5223v549YcP06zdr8D5KhOfRNIStEPFGoH/hX9w5LmEq0K+zdwHmkt
1/p/ivnW5Msn6yzgGAZ1KrGwATYCfGxaRUMQrsTbr5BEXWtcB5JaGaFW/RoT
/CBjrBKx+sn1V/sLnCJfeBsFfEFJg/fyEDB6LnXduNIKJCac1GvEuxq+hMt2
wOjjpbWqdNP9+wUo6xet28uWC2mXNN4/m7/eXVBvCMHgv6aXoeTvT62HRJkk
vQ4RZi3Grhl6ECEJaVyHFI2IfLqTZTJ4eTMUZHsSIvZHjlvycDctWuj6xsLY
GrzWOiqp8L2ooJuyX83BkbfumE/yM4g6IlVzMuFV0DGZNDeO1wNsy8xwmIPe
467H7PodysxXFCMywQoddy6kRRgZHxn/9ri9hoqRsG8IevP5Fhd0LeNMY2XN
DNySaGvjusVLLp1Og65ZHvVznhE2uvuBLFK1p0r+xOj5os59jRcMmveBM7fo
OUMTFd9dAI8pWG2Kt3m9P5/nMFyjUyve8PnNUdxIE2pA4s2bXP+zSz4ez6Wp
ss3iOyZ2q75Le8qw+osKvFV7EW1BBcoTjgy/xEYE+QF8z1/UyIS4DogygnM+
JKU9S4OxRi2ObfYhfFPMjonn+KCfYJCw1iJLlnlytk4Dg8EgUdG3d1ObvlX1
3FF/qYSxB4G7wRkjLBAjBIPwFzk0jgt2Q9P9eVl0yIEgp5gKQgqeHj0R/g/E
IcTqX7IQcH1qWYQAwRLstwU35UH5xVCoR5G21lzzQwXapmPrIMrc7vT15YYI
GEzMajP/5cVk6Qpw7PKAtceyNhUIXxFO0tsMSf3uqSMt85vBJju2lKLWi5ej
XmWuCsjb+H0Y0Ai2eOfQWVrAD0CFwOI3g9o5vOMqvy4s1DDh9ZMpoRfdGlOw
p75d+QKTr7esjqihQ8R76+O1esJMWxIIbCWap1PSsu6gjgr44BdX0zn0lvG/
MS9k1oz4cAjKRT1JiOtUENPlmVD7rt5VDm8OzzxmkcjSh1SHZFh/we+lpH/5
Bfjqk0P7Dp6MfqO8dAKnzwAzIaI4AsCf1LcsHquIPZQQm3IY4Ik1JXJ0GCI+
RWMo8a8jpra4fS446vKw2jfJ5cd58YNgrUkQsJx69YD/70Nxfw3tHzPkZF95
qIhlC9aYVCD0UE0upaH0f8YXY3C//wcBE6RESndAVEUWFBBRV6BVdEzNPUKL
Cu83M/2blpxmRgkIQ0h6rJq8aaKHuBoMDoMEqGxaasosnzaGsbL+cbphJRq3
qaN5oWwxxfXPlFRzT3OECvfSn2sWjsnV19pzjlIuM1HsWW6hJYxIA1G9+Faz
bjIY/8QydEhQCsYlA838FHTrklmnv7U8HLYtKq7M/R2c76ldkNWUumAVheSB
s0nten9tNUBSXZE8N4nRYiRsJGf79KvN1//1ttkWOM39oSmloE25cMxPKvsH
KnaT2b562K8cTYT64RZa3Cnp2HYf07rxib8nH7O5yUmXqjvHCDar9JMv1al1
rGc0fv1ROKyctEdXlUdJjkmQ47WRjaiWO3NUn1S8kz42oBg55dR6EWSwaiw/
dzi1k/A/VRcX+n3742+5+vt/0m7ktviGy//J3EnrzjAbMbfC+9OuDe0o0hNf
43segsZZ6VtdWfpneJlTWPDZ09VcgZ1P79GWgCHSoUgb8Dcjy5UwcbJTnMBz
i/UcuQ4PRD2F/6sJ2S2G/LDokO0ewLbtvxQ0eHq556raUvFPqmIjPc67yHQU
J5p9mDn7icB+H5v4ryGBPYrIKIMROAHcW4j8of76nRFNQatgNkVu8ITiGidM
GrO3pnWLWztKuP85qMDPnl7XXiLoBIasyGCqVj+x5lJHzA/9Qpt81EeOHwTW
XiQtGFsDjKgeur3sXO76gEYoW8HrwlEQf6/UMsrFuS/RwOTltW9fcfg8kenh
PqEjLKwFERDv42FZfk4t5EWO6TTa8eGA/LeDGxAAy67sC1CI7BD5mGsXDfVD
Dr8tJIq8eHw9M5+jZw6y4vQnuk9hWZmeKP1aDqWryuuWiaHfxF1aJWHmpFL+
5w2NhG2iJ7rw50B0Dy9YbtMZxq0ROpa27I9lwcKD+EgU2E3xf1N/mFAjla0p
Wn+OvACxBdLklismy7sx0d+ltpaZ1BerPBgwuAX4FFH09mnisRY8XF4jqCjj
3Asj/QWiJPHh/BN5jQjPnI3Em0nJeMJ8niTmxZfm4MOwz7olVC1mB9F37ykT
P0GyEOscSd9OtA0ZOOcHt3MVdLMSP60lQ6HUKxvK/ykk4taVz722GBg5vat/
sNdN8OZBjUjy5Y4p5l6ewPNegJzpe/zlcn2vDJUB/Q8r8e82HhOa/jTpvd/K
dSlQnrOza7V05mDF5txq+uWvSmNLzFiFNtISIsC7B4FNbJHJ9gOxp/gnl3X3
57YteIPLS1vksC7ctWb73OXK4AhUuybDMw1Zbr5UbIoohb5geBEuqjQ51MAv
nszyFbhNYXCRygAEzFI1sA65NKjiWJfgFCgBEGw1TgUytwQzj9ssxjIAzxsn
FhWpK/ULAqbyQAFhn88RorwFTLQQiI3mIMTaGDCN1/0gRYINnJcNGsLeJ1PR
L4mxWWUTonrfDDc3rjD58iV+poVZ0HnqNshYALF4YMh2I51VX9xdxCZPExGr
4otfg4yAQFrnid3tH0GedUQlyGhFcQHy+zvf4UU1F4gJ4kAzA3GLyjtbiMUp
9vm9/qHO0Nz2y5qBlsnpId6bE4osaiTatH5yleXfWUOWuCDeetz6NUnr4ssV
IY041wTNdQ5lmnFa+kb3ovoBRU2uuFBBauhEZHiPAISgJa9JEr/wNs4uKysW
/6BNQ0i0zYm301pUs9Eh8YJ3+Ynn1v8q+uXEMAKamL0bwnh2HNUnBB19u8Nf
lanSFbXx9EuedVgMU/PZdVXDMkI3d2PJcaWAqnaqcdfmJfI3dQREZetaXvHW
1XdNkxrFCWqQhs6KtYSbPnI4uEyBBVxRJOn5Y5/T4wiJDFkD3V5ai774mnCj
9WjTMI7HhIJ5IK//LqmMiSdI1biti86kwWMRrz7asA9/cmSUwE6WC/cilTCw
nDL6mq1J/Xg5R7bf03qcoOQolAxg6E5CKPDPK6vY1/KiqA9PHCXXGqsCeG04
Mk9TEwnpTpzjW8uFegsZDETLIQczNke0uCaVwxvieb+bh5cYcS8JiQt2abGA
ApdzsemXJmSKIX8ABpSZ/SM9dwb1/0FVOOdtXYgZDL8ZgesdZzz4M9u7TqRo
gpkCbxj17CcZkpPkSbGGAppp/NJF9xk7vA7STOSrXWT7I/H2DOSD/1Sy+0yD
2QquvS+chmjb7Y5EltOdBXg4FcSc3f68ai7HyrDE+0z6niuRDMtCOn1+dlbc
awueyy08EkC4CJPAr9vuLyHn6prLxOYl+dV/JJCzKnfIEL1PbQ6mgMs2b5q+
QT4xPPmYyKCtJTk6MxiRM9lwLLwGs4dG0Yh5dLespOo9hi3tpUfosUkidL0i
Zqo+31Z5Mi5A17HN1ejG5RKVc2ymTA3L9vfwDYpF7Ml5XGqF1EIN8gVygDUv
B+SeKYGFPN61Du3KxguYNXsM5rV/MtBkjLHzEO4utSgW+1g9SfeYi0AEOWaz
gp3nivVcBcgseJSMiik91NjYxSwRLk8dfIl/KElW8cORmbl5nskY3pMYf4qh
OSYUIduvS0N/0INOYWbt8VAODmKVXVSYEUfY/nQoKqUQhmgeryN/AKuZ7zNS
tIgD9RbJYaIUHDMhSLG2snkPYp78FE0mLzL02w7nvqIFzTu2gdm+v0gDMbAp
Rj3Xlev7HYj+nPL+tzauudSV1SgfcQR+TOgID0p35CXgQ8e19v/SYTxcgR2L
T7QC3vDxFmAosYu1wHU2m0IVGY8dOQSHujXLs7s9viObBvayJsGejUUlXM3w
BTdsv1hQd8dgF0UpKHy2KHguAphpqDwoX4ETZZF1Y9qKb0NuRBSdRAgt7U/c
znPwbWs1oKB8chb380PSidtLxvw258J5zldi55YgRDlhx272cZPP9TJkYdQG
ip9DkHzJ3A1OKEVo6z26O1wj6rEHhF7+BwTcXSorW38yPhA+Y1smEjbul3K3
V76UYNy/Ab5kTj218p5KcFXzycNHJwESktl0PM6lLAAYRMffb8HYFc+MZVK0
uJM9zZ5zDgdF+tRZ8Vxm8XqxGPqfu7cKko/u6M+ec2395gTlO19b05rWh/6n
EGEM9n85QfsNGJ3FlAOAftkMJyMtfiyTaOcgUslOfzLjSZd+Eg/pvbhtkxzY
SoF/YGOoQUOLz+77uRtLflpTpw8TIY/oOXr9qzPm+V9bl+pTIecdlu07mQpi
OQBC8T6Tnf0opEkEjo/4L2/l3bDxHhKfYx7LCzW7Ci2Opc5Rzp6RTMF1vt4J
wchu0XOF3vQgfjZCUOgq2PlF6Pe8J/MpOguWrhEDirz5ZIHdDBDdVUmDv6Gd
iVqhCvIVTW0cNxNX63VP/lCeNZIeyMJeNIOV6k9nd6rPFROTGuMMtJZBFKAQ
eHXAXahgm/y94MM+Z9/BaGM5CFoka9vLA0VnVxTZQKJRmpF0dEEnBBl17X/b
l0BXIKq4RlCgEmmSd8eIJpA0ALeNGi+UDl/JwbBiL3ssx2CUjMQQHwXIzsPK
Q3gVr7YZMxrQ9NzzDsmzBfFsOpfjylKPmQu18Mc5OuVQsfBZdokYNOl5d7dP
gQzfcPHWbGethljz3mrnkzvBgmtlqErcDWThxne7zFXt4BcdeykaPHpLXokX
U7ptfbQWzAM7N452uK+bmDHxCmtXJDvNNDS6okkCrLY+E5YKlSzsB/0TMFWi
FgkyT0mJzA1LI9v4HMVlhE1DWrlX83e/z0bAtiLEMZAvSdnR59GwHe4ZnWzQ
fn94VE+brwpgz8uh3UNzZsKXUMF3skX9JCuykZ1Ruo85RTOvSyL5r8e+xK81
JQ+Y/2J0qYih01vXtd2jIPI9LEZnFsdnSP88qdeWgxuticQA2arwEcIAhT5l
szx6NIkm3eET66tI5Df424YtD4gFYi+qyc5KPS7Ji5diXKM8or3HtrTAA5HY
hg2/pD4+RNQL9hckRMY0aDDM5kDZfBKUTLrUxb/KGqHJOw1ZrO7cpxeCpsGy
bfb3IVjVb+2EiyV1oCZuZFNrWHi1YpGTHeHBBU2ZlLsexWYyqQHFlRFd2has
yiQS6l/v4wjKZx7hdmXtAxLLlqv3ZRNFp/hXPpRMnkOfndyD6hyFUGcHgRBY
9DouCVOK8rOGmpI9KX1mnI9eA32JC+F967sQEmjuhvccyvDZn03iZegy+vEj
N0b8RNnbe+Ab//z4DL4RI8Oq27alUfXu2x+DM069r/lSzlT3WGnkxuk8ALBA
L3UDTIRC/10mxJLnQa/sAMB2Gf6EnNrM9VkPxWiWQgU+XV9xIB0zzgNseE80
yntHuKV4+1/fwrV/8GPfEn8wJlxXHgAh8rGCdQVNkz8b99BWO94rgFjk8wlf
oZGty/2XuDBpLk6ZGiHS39Rd+zYv//SyBaW1/fBbsmpm0Yb7sOo829sBPIAn
l9XKh+BvU3lTXwXS3wGxslvXwj57eNu9lQo1IoLb54rRhrgFkMIvzbg11FWq
OGBMBD4WBcbEE/2ZnlAGZum9/g2knHc187E9T+X+cbU9va8S2K0XMapX8ilL
XIsJKOE6F6of3cWoYuwt6mg1BOTfoxO1gh7IQDGEF7R6Wu6oFcH3GRwPYSAv
4u6P4KxH0w5vYdq1IT6ZDjeklIcR3FLzGkH2g0NmNPEKBkMPoVe7IHxd1zWG
qVyJLMEjg4tHYVXC4AHEON9tg+Ctehn0zBvMxQBSzUqkvakA38RZCIYgrdcu
2fqEIRTmsaIsFyl4iX1T77g1OTIAEIvmajswLaDpxIkL9xLipcZ0CtZJg+6n
Lav4fyu2O6y9AoEg+hTnY1knxc8Axsu69FunzU+o4J1dPb7yZihdhlpZpi8c
VFnzVX7iOz8OUzEMtuaKUsjyiHy4SVZ/bij9zmNiyRNs1TE/7rpj/zd2q8GW
uuoY2JGGu6ZHI5kf4/f+rtS1f9blFN6LIP8njYEUXWHNgGFiICwZHs7P4HFh
W+ewpNF5qJfBICuB1403TEQbnn6nGdrgx05/QL0kwyCGfZx2sYx9ZkW3KfRY
eJEsXKGzOu8SAnVaQKnfpFusaWcCtkdccVxJy2GWXu9Cbz4kovqoTUmHhh1g
Xi8zLZfiTC908iuzAavqZlbqcG/CSuAPjvIFSiOKgaJmzw2go1MdZJUchblE
7P3Gm/844C2VN/lBK6ju3omDU3JOsk193S8x2PxtHfU8af3kwvety6cBFfOV
+8x/HOrVhJ+YV/JsfGnQP8ltK28kLOAowQlxBdDUcy3wrHnmZrx5qe4jr65B
U+URqTw5hayx7RcpxFE6foGGzGfwZvXN9GOoSXhnzryR0DoOuvtdttbIbx80
AKMpTLga/tjtJt8QMl0DKSEKIH5OYtrNfvrT+znqRkE3uzir1McZGrEigt09
5zVkGVIcn3/XbUmgP69npcNzceuGwUo0l/nmWRN7t226B0o+SldCtIGjqlBG
xHZ9+ukYo4GvQzBUX3klUeUWTBqSxXCiYYGkodpnRFhxgWausSJ16388ER9o
L2Qrx//bIs/zBXZuCtcmkKKIEGxmwimELWfqGkmLlj+1TaVk64Rn0A9lEMSc
JtboneyvVc/hWKJMtLBxs06PmZEQMdoep6X3Zvi0KikVGW4rwm2U3Uv6kD1O
H+uib9CSUpHkGUuJF7drPcHydm7POtfSLKyCx57LJU/rGce5MEnjo6DGb0Qz
RKidS+068TXK/+gf8I4UQpkk9Hy/I6PlXXctJyPS/0MehcUTcqoQ6GksI45B
Qq5Lkyc+spRyE2xIMZlhcCv7OHJ2LC/ppPUqb42Hmx5/EOkVPZuIWFaUoK07
G9xhO/lxZ2vHdbipcX/aZK+IHPyqLKt2/3mCvE6HDkbfTO363DsZNbtzsSoR
Wr4KqpXj3T0FdaZk5lfH/BR+kE7BRfgr9dv24GKeeuI0xs7YggVtjmX67JE+
bbWoB33wWK23adWZqv8Y0DsMBAGC1VsIRcIk+zZNIWDE8nn7pUawEqs4n3Cu
pWFvnaVSFAp/yPdaY37r38eJsj6aKvkkkh6TnehA2WQghTURFUBxggi+IECR
Pp8xkXswHgRf1EfuYbGAgMevJwoanm3TK3Auop26SPXOiXohfDwdzD99vowH
M0kYOB9b3CWJNXxXAN6AYM5xR5Sg4Q7xyDK0g6fGhI9F6VfH7tJVQz1vYBkr
o9hCcdlm7ir1tTCUYI9831Thdoigvdvu8RSJrisVe1haAf/GUy0VBuT5+/z8
gxstpiqP2IKruIuexEFqmqRKsNRXTAhLkTs4f4vFkrX9lbJurP5MQ3PmpiSr
PHpGYLncTHdTIlWAVEYSZoLIoGsT3nEdlvNsmqewerkNzvTgiUwDCCAoS+hs
VVrJxGy6B2EUrVQYvP240eadugua5aM/7Z4lFAgzYMUXrbITl+zOd9khVpNn
DOyYtOSuV8d2Rnfpdlc2vz3YUihKOwV5ZExI5p2Lx1VMhtKkP5Fj6Vv4wNxG
zr94AkXYRrdH85WPZt4eboQbiVk5kPlmRIr4SVi3U3pJrOHsZaSmQQQa6JlF
Cl+SZRSj5kZIaVcNjZQhbFVFCUADkHXNIWnm7mYnA0ghNoOI1Z+StbqjNNEP
VS/2/PKwCRDFU39LgEQT1mDNkunABJJ938FgRmlI+rSgwPX31iI8f8bCq76E
yDy9A4dtjV2EN9i9lw9ymPGL4i7LD9vQkpKMRcbD8F5vZThuzz0xczFVfr73
7sq6m30KQaf5XDKR+YP9XL9K3ohpW+mXd4IebkJytwNf8kU8i5bGhjFjDmX7
C40UypXjN0h5HfkWZtSQ79IGV1gVBx5usXWZ/KpjI2oDE4uU3/3t1uRBsfeD
G9aN4fzLY74lsOR3AEBDnDUCoTdqTn9TgVzqEQw6Bss1LQaOFBJRkCPRwbg0
ETkKoj7lAN7CvQVnabZxOqKmOTX7/gzQuvzs1GiWhuqoj1q9sZVY0YF5MijP
ok0i9LlZ2y0+RQAkNDJ0t00yBhayXeS5qF4mq4UTEf3LF9QNY+mjqDE+H9sC
V9B1Q0m5mNy2zFgLU5eWWEvE898iZbamxGFHNxfYLsAL6pkfDM8P0OZRj9YA
/SFJjCuuF+JaK940Ft/e0C3CVExj+5xltyTop0g0KoZWcyA1vKVkiryllhke
VW40UiBQTB5Gb/wD1jAq9Y1I3Ohw6LGpKw5SdOE560NnHsWweHM7ANYLIXO8
9Em0OZSs7XlXU6CIMmll0OpxW3FNAfBpQ4hz2tJJJrLNV/mgLbGHhfRo+GlS
LEeLSFzDYACqgKu7Uq0VeQuw0NWKIz2Pkg/F1e0fdOU489uCno0pvDWVlzrf
TcPdm9rzY0IyI+jZeBqEv4RQx8eYB23MuSvwdWADXuRmsPu3beP4gBarSafu
Md5TwwykQVwMY4DetHONyBm5H5qyXTWW2g8u1ohD0duonwwChaZHg/il1Fsb
9xxiIQzjvRmOOE+c1R734JbJD4Kf7c0gOS/2T0MH9cnrLv7cpLvFuN21KZl4
MW+He8FmFxx3APedI5hq6KkyVUZk02CjLDiQjN0BMEvj8qsxRDj9zHQSPDwb
MvUw2o6MywX+68w0mV/aKFMmc/2VKdIAwDGCCgqjUIXZHnI3jgQBVzFd4VMs
svAHFrYWnjsKB1HxSJZn3Koc+STbBbEQU4UZg8HLKd3SGXH43aUjpkjqQB2N
b/p4Mk25q80SkHa+vQnfYAEQlVgm6DlI4t3U3iRn+I4AOonkq6ht41X9/eXU
5AnDjaqD/QdWZV0ulWXbWLhj14zNoXbBrohL7FVEgmagSmrG+Dg6CgOYEXC3
mwzbjzqryU9jR3AowMdQC1AFXdBQ8THsJwb5Yy/jmq0lSS5m58MiyrCLoFmx
rFs8+fQk1JRVBnWcZ7H1Mgai8pQDixc7rtctxHQD28yXWQLjqm419ZFhpjgy
a8c8jvPu+zkJtJi79a/c5e10BtOVQ4UpqfzouyIgbTlJDdTEclJwivks7lbS
nMvSUgehOtiPKubO7Tyq6VAIblgtysL9j2VWZL6FSPw4yI+rojw0Mo69wW/f
vztLmw08GILhMP9h/IgZH6UYLACQLbehiTUUXEW5rz1ArbuOrAUBdbwf5kO2
3LV/9eiIM/9ZQMxXP7FbEEkP/EUqldKf8orOdd6xLjyC8/KRVIS0W72FoiET
zlgPL5ywstODOpwNw590BVFU5dRe9WP27ebEhKmfDP1XhCw2v/Ar2BWtIfvJ
lg0Pbqjqik/EiuVemNMllcq2o2qkB3vCVf5KDj9hpGamw+WxnruDIzpre8Z9
0Bvqag5xvHLP8L5gbUtIrBzytO4IfCjXiwqfn0Q+z8cm/ahD6/fn3PySP5qf
jSlcGGt30Ic3Wmg1ijgYPMGUnK7F+yS9zpdqhdognoQctpB+edklHdL4dwOm
9QvXn96jesrmuqVO9Z2YYhhkk6X2ZcqzChcLbfYbf5nXqxiupQbTyL4235wY
pDf8N3pV4rc1YlTtBEqBoWAs++/DEFKf0iuzFq+tgv9/xNYqqiIfI3JB68W6
l3cEOqkTYk3GbPIp1n8+7gtPTkzK/pnQ/K7TyP8sLps9d2S+S4IxvZIyEKO+
2sHvFrSjHSSKWFIMKDMj+s3z8e7PmbtmEK57/4TkkhNZ8EgoP/vOXity7RmN
Ju5hBY0gajPWqVRBcsGrXAstI9IvTUErOyaI/nhCfMYaEtL+HYwRZgjFJbqe
21VK33H3BxQjggwczrnJmNVJ+/+MJ2bQXITEGdvKTZtl0InNIdgrE00O6tyR
FB+7xEwDu3pZh/+EOoMEQttgB1yJeoPppSJS6C4dqnTC7I/I6Gn0RvkdvjHs
N25UztqZ8W0zxrtEL32EnRJPv44hjXLv3XD+X1lkl8m5OUkHwdwagZ9m1J6w
ufjjJRNHZ/wdUEgLUuHkD9XcLGLoNobnQ9ATo4hWGa3asZbVvx0hUQl+UsdV
X4/5mWrx9y8psCiQYTYAEw36IEoHcCopJneFDKfx89oKiR4MyjBzmkoAUjJI
UZctAh6VnZURSHFtyk4LZtDhy4E5YXztAbF8WMH0sSFLktsHgyAxM48Wzo+8
yctB+eD35yCZOE/fy9mebdDz8QBTgN+PMhtiBUWuaC42tJJTsBi5d0ZcRed4
V0b9vT8msLEYESCMPcajYKSUM4cSeSKdeXPYKuborSbwntacJpAyofHaisbH
RYgL9aApL0tjKcRTozRKigUiT90IaxgkIRxMllx3wT084afBiSetBxu7I0M2
WyI63KBBN4xHEQ0vdVauXUu3fT36M24Rou5m/RUSdI+1oYDJNF9tOfzPC612
D34E7HMJXG5KPprozjopKjKex+Rf/NkdIEXF/VRfBQw3GgYXQS2ITdmIjWxl
2gTylJJjxKRBoR4E5tggdHJKFuVMvqPtbN8W3gSntsZSC++patfurA02w4rr
PFVkZ+ksUtG1Z6wz0mLU6ehvfBxLW4VOBGBd8yLciU6oSA8FwxcswHVKr75H
0+ZYlOuFaDOw1mbvsMGBcLTViH9fJcoR1faJ/TKBmnxdnXHIPwpXnG1IrdfX
H/G/gTpz3IMmCqbb1BZvtos1bsmTMVwqPcj1gyCByqwrSDB0NOmpgSUrtR66
5mpylKiAva6ud76+QRtPlZnOWMybO52+V3jodSKVKNpsmMJoAme6+DB8ivMg
Y6ZmwDvSUjcw7V2EowSU+fmox8VEj6ILVM77xgSSNxn4pLwzNBnrSGM0CYgj
Z5bpkcfT8alXXpd58789K3/wB4DbDy6uXNjrGJgWvtMA7xyx6eqchpHIpz8y
uI36Tw0oc3h1QqQOADB4PYk9KkN6f4qNscMWmUtshTaTU7oxl7rbXZ/c7by9
t2+PDJix4xldUwYqS5UIHWBOwglEk0ihTY8+owtWUWpOiKGV4LSanEZeChyM
o1zIyny+Af6nZzycDwUt2BItcimrCJJm9rk+/x1CeoouwEjTWP9/PT4NZT//
ft8YRh6M9CwnZv28R22uujy1BIsPz/qL5rSfwJvTzV5Cer7iFXX6sCXQ2FBR
zy3s4+vv/M9o6/fW2QKnRVBj/nhXJHRXpTV0da2IxUCouhy8+P7KK3WP3PR2
FT8iA2MwcoBMGeNtNkuOvFxXCzLtdJIJ7EVs61iDSfwsR0fnfRKL/JBwENdQ
VdU5ZZd0I0RGapg2TGc2uZgLvq1GH52vMtk27kbQjDo5x721YX5wk4JZR1ms
U4c7ziZB3bb+naVOMWw34HUT00Q9gkC7OH8gd2grf/Feje7cpB5sY1EOOYH3
m5P0xiNG5YQYKVaxRKhWDYT3gTVLSH243eG7X7l/Ub+7TXUcX1d86QXbB0yP
o87Q9H7a3NsUmliiEkBIGW0Dp4nPpiWjpnJjYGTSvJERDcPeus2t5DcU9sSI
e22EMG6CTIG6Xel10MkeAB3z7cKjuwuKXEApuvGs8N0CZJz64edKoklXv2Sc
pvavFtO7dDEllXnUJ7qmswrCRsGCaDVwudc4Y87QBosWZobwUqX+pm9aZQCU
JmZnBpQUd+I5hzGgZ6hMbn0yMBUKYXiCD+9snezZ5AR6vsboK1lN0l1/RqMD
sbfqomwfsfdVNaBTz31JHsxkkSvCv1v4gYIpgKUSxt2dv8AsgeLCPAjEeFyG
XdhnzCvGvh36ofkTG0FzOOcuWRLzbw/DTbenqUSCfP5pBAvU1ehiXxJfQ/Nd
nZl/jVIzwhPNKhBUhxg9sxmRG4sdJzuvrPEXD8ZrJdSA9r4yO83jycZi4V7B
z4YKQJIN2bdxKUX2tYIxce2szaNmW/Xy4zIOIFg65P1D7QsI1EzSKP4VaPr9
O21x10jhG/huFT3A2Lz23DKn3SFyySg3MeAp5u27QgoQddJehYuSzQ9nfTc6
wdkbpKo7lDcj/R3yX36woFB8dmZTsJ2eB4cc3KchtpqOH7R38CymuFUSbcZV
8YVoDZBoHdGNKve0L0QFnIng0S7EeUs7SY2a3oovz9MwpUIjChvt8m7iruFs
sRFjtF2+cfvw6YpXwsaVk3/2FHBNh1scU4Zd8xy2NYtd1IcCYlnHoMCqXsHc
y+zREGsSRUJoeKFEJRfrB0xXmEj6Sm0VMeqgGoM5fo9AXOV749VsSlJ5tIzJ
fNJTf7rJx07JOpnd0u6kc3mf4JAxLw+QHKi8BRBMGrNX2A/BpJjsR63FKnLl
vtaIxKjMBrvN8t7hTNES3MFSjPEYH5+QArdpTkJZ1hSB5ec9txkfJrD/yRkf
6NorIsBXbka5//uiIilxjkkhei28KRaUYPtmqAd/dICcQt2hg6M765+nT9gi
rEeNfdNLpoKv0GjTV2u+1BXKNaSrdr7MGTir7dwLYKt6Ewsq8m6gNEZUUQkD
ClmAvBMpDcE0q+KvUwq9q4B0MuPlkmwfCc3xDhEPrsdy7csqA65vbQfAjTp9
iCbhbsJLvqO2YZ6/5cIaJEG0HRcwUE4C0V+jkrOMKd8Oe2bQyDLhvKce2OQ0
vGVn+gV7hh7Z5g9bjIU3w8io4DG9ms9eL5AHODa8Q1XZanAy6LCyt4HUNEK8
881sJyMC80azqcFjE2Wr7pp5yZndgcoIfzcEW7tB293bBaZqyzAQbbN/lMmn
wfhz91d3hGGgOtNTUhzbWTSHYm6+ZiM0rtiaD9FGC71KRUTQe7FDWCJKbUik
t3qZpTZDsNGitavUeeNA8RzLKTuhCWMPoRHkQrYdrLhzq11ph/uFO/k/hBzM
G1kviF+JESyzHirGwK3J206/TMNjldOXJ+ytsl2cTdeMOoEmlwUFZgTnqkB/
TgksCfRYf4UjClApdA8n0w4J22H+l5wmSM1XKDtcAhysXgme2Qr84rl5W63M
2vzCQdKHx6SZsmP5GFxX3Yn90+Rqhsb3BcNVNaLATSnvtRXp1MaoU2y9MDVX
dGArDd9uarofdjnlWsT9PmBrs8NL3+sQ+PyKW/WvivvbFD6rqO/N0dkvqe6R
ysa+7+6prLag06IJxFYCG1E1zmegHo6Oo4gWg5hcwIFOq8/7YvHSxObf3Spm
DrBcrjKEsusDrs8vhhC7NSoQn53Rqg3me1Z1DTupz7LdJL4ckEeKNQFqq2AJ
7JCQjiBrg6/tN7MpcVbfxAjKfQ1LKkUqMLJpbLB8AaSrM3CueATIaHnq2Uiw
KhCVhj1sS85rWSyfMsTGVTt0LrOWHBbJMMyybwVizN/Pw5QOxg/u38CTQxSo
XKUHhcvph7jDQzovHWtEcXuc2Ka2n6za8DrOIJNM+c7TEnCLDWBD9Omfsxf/
lHkpACE5lISTo7nZ0TwBPefx5DFcBiukNpCfVf+S0YMnbQD0+Rgc+NZFc6uu
JSEtmJCwlCXiP7Dj1vQWiZvWIlTG4Ph1QLgYF+1FIoa84w6Q6sPPhR+Znm44
byNAWfsByNIOsiMQle9RJawqs7FRIiFNOt8AMv5ClN1/AUEZVjEAXWPAp5oq
H7gWZcW6/ZLgAlQ9y+ks4cN2RTYwc5uHcmpMqLHbO7g+5tbRndsMBTvWNFiS
i/Ya913xol/TwQN7

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1LmPDHQJwrR4AI87KHlGgtPllL3/irn8p4+5dzxQU8hp4tI8p6NQ6LmjtvcEm5wb4E5tWX+pt06wvSpPDwVTSV/RpxrZSGHlw+DN5vh65yaoxkfDHUqULwLToIs90j2ci7zCDQOMpiPNUlq0FvDNnWFTmW+osEDNCZQqQu7Z5W1E3cXjZ8vB1SJMeZvNRncZnDCr9NzrqY2eycwYbw0dkOe2uo67dH6BC2M6JR95wln1g10E52ldl+2ongjwewjyVtNwNt3SqKe1kPvGXDNuUs2Kx7Z5NBdg+7Kz3f3xLw8Y04Ueyr2SCmNubo0+9fOF18dUyUOqt1s/hoCI+ug3GA5fUFA0PgbE2NmSH68zMs8EUDnozn+YB65gjEets6ol3XEr+KVbeOZlWi/BCtimGD/xuO+rXXRjphT1T/WDbJCw0K3YlfB6S8GQtvJ0tD6G+ybWlQddjA14f3AAu/RlZYGTNgZsNNOOUPt+1XgzpQCqr3SRHxIqW5gEs3dSICBvHagIRne4I20qCGjPBjRRpANlxhjcFHwdv6Oe4siGlveHv5On92h3D6maE0CwcdW44XS7beDa4NhVFTAAWdR+d7vsQ0G05xnWRIs4kvo8p0wMGGs0hIrqOSrXF6FrmB5YIewxz1uAlUaxlxdZ4nRrXsBCITz3nxAZf7hu26uDFA2FnUvJA/nYAlbxzzvOI0EmpGXGRQzAm7hYoA2ZS94Z66bIXAxxvvNgGeaBUP+rNGIgTJaxZA0dhfGaJKgNUMnOP9qPBKCinXiAW2WnT00mQP2"
`endif