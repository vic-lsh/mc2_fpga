// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MRv1BA/i/HGhIp6OmFKU0XXC+vjTQ1WEk20JDECzhQsrv0SKwdf36WJlJPsb
G312cDfnMDuaLuUhgqbNVPXTtlyYPyspVjuLMRnpN9954q3AHgADDCeJcuZF
HYPAB8IZS3jtTCJORc+NenAWCdbBBulzK7LUMbBwCKv5fjukQTdipTT1FhHU
SpC8PvPPR3VkR6sDaXtSMUbNP4OISsuDh2AijtEdnvWcwU+jVm1GMK5pz8eq
hD8dw9qHtsysmfXeztu/E8xAtqGBtkKbmYAwuvxWYxf8gIZdZ6AB0Dzi3bW5
3IcHA9Ns0a0qR9G3hkiccweh8UB/3ov8xotCPO0cZA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mijCpT1wbRxg7936HLUC0PfBBdqvz8CbIgWDXNE+6tY2SHG/3YKHwDvPssUg
zz8x0gwqAcqJAGYZNOzAmoMtZoiABxekTUrVgSRcv41431yes07ch686AVSG
xdF+ZHZ9e9t68jJfzUVVN8Tl0xQIWlUOrIz3XuL2RqbOp+Ig3nyYU3CjEGys
I7t1v/Pt3zHLrbzuOLxldTVcnDaMq5JkSd90uJ5FeyI9QUSv5VbqHIOKOeBi
mSZ1VjWGwnRNoVVgtzcXfN8Fz5Z3+7EQebbyu9IDYDsUGXNR6EGoEfktMyV+
FSjnqV74lhx8kUo8ULPFfEacjYwoc1Yxd7NArah3Ow==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aOtJGbISW36ko1H+oXJC4BVEEUjICBeNeF1avjVtuOUnXKesRpfvMU95TSVx
1jsYGJK+D+FUGZIwGdzkNewFNGwzad14ZLIupRrJVTfvmN7Pgx6Ad40UAJD+
3x/Bl5AyZiybwT097nCaO3FIyz0E9w+qxbk1gWxETnjCflZrjASoxhSpGgf0
h8lp+YIz+9R0vkKDarVaO0fITm6DZMGNT79J7tEUMrYNYbcyfNKtS6xFoiMW
ISx9gDl6W11R7VVSr5L5pMDxIAJLLt2GDH4Ngt+0OYXfYtvcz4Y8gVo1OPsN
Nr+82coU2A677S0lINoLljTXF6wABYyrjI1GWRg17g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nyYdh4s70aIZIkMDDMm0WU6tz4hJe0Ec3FxfmfIBClLP1A7eOyHL3IUV5mbQ
ItUDTg/WZDXpBQL5lZpQkUCQNPuJUqZ2gKuWrES7p9AhgWCNr/FG5Ml5ZSvV
lr9au8U9kn8x7pY8Vd1euAVtg47vfQ2KpiXZ32jpyMzMce86aOYn8txxf9LK
yEBea58U9iPclc+wadU3dpfMnUK0rQNul0Nh4BNF7AtZMpM4KkZY+iMA3bjh
vaDIS/WOOwlPhIcZWHA1kJqySAGTGhJHjvlM43tOWAYOt0SduatLjidg282t
uFuFO5y7I88o78LCbe5m7nYYMOaXCIGkpyTLQIYxMg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jMozA6KouA2jay5nJ7s8oV8tLwnUZpBt5ct3bTMDJ6j5AdpeGxzXgRO7EhK/
8YLw0Kw9MigO0b9nxEG3kXXD74NeaQb/sr5a+Td8U/1ctXPalpy0yLax48Dz
E9flGjnWY/TmGOYmmmYTwZOUl3ZrVxvwo5LM4nONlhGxIGnqAdw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
An9bxd2oEgTNvkamya/ktdovrbUTmS9hHs3MEoVZKE8bP/4cmJLi5C8iWAf6
Fdsel/pqJGIlZiu5LHibgXHfLIVwdI9WP0vFG7ZF6Cb4V527O4DHkc2ymIP3
bNanYPwHZnjSIskaAjGuRB0WjMKWSyi99R2LFFPw79uxwa7THPu4Q/dr3xxX
78e6kI/7Ijx4s9awJlmnTS7L/6sm8H9sHJZe5zI75qTxWinvKZl/m+1/5mUY
Ss7XSQauW4EBkXIX0BF8/ekV+PcW3I2+b2CtToZDPbhGOmXmFKDkrC2+k03f
U287hbN2gfTU1nvmCqESFx1gASHGb66TmuoqpxRJtsPJ4M34vT7lOVGLAQ98
1I8ZmAXOrGrsb1/Nyjg1o5ogRPeTUvld6LKU5rcaSW6Be3Qyq33TVmSLQJl6
YETeKcyfIfqyiIr+X1GLRS99l9CN6co/vfnUqTjPFH+DPLOMrxNA6AkWnqXG
sUXjUedlDBJA9+xicV7oaKnfmAq4P8SY


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cyJ12zI656QqbEMbNBiRdyUV2xoi906dawakvQzqDSsWfp4JdiVAJdI7SBDu
X0NNtAM31DQEvH9CSdCcz5sbnVw/wVgWPAOesaBSd7+XhH15lF7Rq+9NXlO3
D7I4h6scvu7PEfrtWPdq8IY6mkSUc8RoKWm3lgU4XAv6sPNOMVA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fco2GrJLc3MQIkZu6/HDm1Qd4sRb91ZrhmB6CcSkc04TJo4WUXqZ7b1YF1Mv
I7y/L9KNetg/6DJ7v0z1vFxCKwfij7Iw6oH1k2S8/onq8AtNAWWq0vdCXv0v
ZlhUdgJ1X1N+O2UmvNp1E80VNLT5ljOuxZd1IJE3R3ylDrzLWxI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 56352)
`pragma protect data_block
sis15S9FcSjPyEQv15xLeh3fysiJTqY2iTaafFIwrSa9Da7uJgB5/Zl3gopD
Ajld8aNCebtxcmH4ClOq2H+YrDpSGDNnRowzExfgkMCQRw/GH6RdxjGinIj0
PdFg6MCMagCf/XPbeSIZxu6MwTzdR1+2Ci5Go1VqYbfxJ0dGlny/Ht+5hvk/
K91BIAjekkPWIxdtIq+UlxQRneaL4tLMSMq+r/JFhOhhvqqOlqz/ZGPqIluX
ai8AMDtLZ3TP1Z1yR4vF1p7h3GOE5WSXdgFceq5Ur4JRd+nBL3vaNsRvvDi6
tYRIS9TnT7vtlyhwNKeUKns+73Lbj9uB+sqCgzfC5IPVwdRxeBl1c6UwuwgV
Ewioooqjhu98aWlhRTSTFIAM3fz1THr+GKIud7Zs7VYCPq+U4f+21MsXk/5Z
0DBjW8yeV/olZfJijZvs+hc2IJOcMYcduQiN74rSWCvZ/LWvkDCoPvCJ6Bey
6sctFKbZESFx9tkJr97TC7ZipIARrz2dJNjdZ8pwZ8PIr05uVvi6BLC8SASi
+l1b3r1+6sl63prpFHGaVGVqehrvKzLaf9fETy6P6TWd/XCSlcxXQ2bj1j7M
gQkYt7DCx6uh15ypUdJ/mAhN9d0hppShC0gqS+5SJoGv/i2lrEtFzyHM18SO
HSrA8lwQy7pVcR8casgnhS4XknJ6anm3Ua1KFlyippmmljbFcJpOE47yn09Y
13t3tehmSZOa6gfxYWvLouj4p3BqGg8RIPn8cBzR6mJW5RbHLegNeZ6FZZGz
vukP9vuw4XHaO4zoZqlp7t0HKf1L9qTp3RuxxinVftxS843SYa3amlqGf1cb
+NcWIsHOz0Rjw3/qcOmptBHj5AugYO+0Gv7K8hSjDZ+5y5CRLz/lAoCFYqU+
1C/4PPN/2jex976QpKzxEh5ClnfmtwH5taWEC4eaYHzWZxE6iRxLdYtLJYsf
a0XI3cIPV2Y0EZsPLFihsUQhqTHu2V1chffiCcdKjwvqH6f9ki2WvS/h/zed
QV/MXdXh0hGoPCHza2RiRSGeSj7BXSJg9j2044SGGJ+k3p7UjyRQ3yVZ2zWy
mgWUF019G2rvSI1esORR9IabBNciC39ouGFMQLD6Hrawz1MFSyPcRNalTu6f
ESLSxT0IFRe8yqv+0Sf5/+8q+UiDYkrtjaOz9lMOsvT3kO8IjK5BnG+S91ZB
/kYuC8Q8JwiLmOekZWv9YKonDe+TcWfKZRxv+4QlOSR4FgLDD//7MMx1PvGE
pWjC0AsRuaBY04BdS0kcWy7qhN6lIN5QUBQcFLKKsjGCh3nJiMLeXXOBXAQn
k/J2oSaHP9jJQMkXd+bjs2Z/3s069CvUl6e2R0FQIdmaHsv71GRic7IMUU1H
PwY65gw8jEgI7/Md2npHm78+JqvWrzQxq+HwK/9y9BlH7Zj+EPG+t/5LGxRe
+Mh9vHNLD+XX+eSkanZajvWYppu5+9hZLxnNjudBQp5HgT72qUnaAMxCDfWR
hbZYQgJGV5XeFF9myUAzW9t8SqO1hu7LTlYxbr4JKmKi9S/QpQHma4DTNYAB
qWJcrL7KaZ7ygVek1H8ZHERRXi4RM2N9Y7kcvVCeoLvP5tc2KscTQjbwmHp3
PXW4XXDFE/qCEcFuoozW0dOSih6cRgtyIfh3Soinaf+iT/JalFCDroSN0H9f
waAv2LZS1kMRPTo0vhixlTDp5KU++4f1gnwpegwOH5l2mwMAH2TXPqaGkpdR
kiilbEeBv22Lj81vVaXZzgU/JVwYER8qMkG8CY3YxQm8/rX0wtWBLXliWxxI
eI2VRfRyPq7JSAwl1NWPVjongtxN+fY03OIstc8W+DmCXmGhCbJ10oaLQjxM
JVXrv8Z8A/GATDO3mvOWlHVpgoW5tBq/vd4S8x2jdK27zaDBuEgVTF09B7VJ
7I3SlRUaAdIRqiIQ1W1VAAxNQ3L5+SpvoQvVkdc8vw3ffOCJqMBdZxGHs17C
abtXOSao1RfoNslmjOCwGI1R5E6k5X00OVO4k6DCYHSGOcX5WuB0nq3oEqwZ
/Uj+8S5H0WvSGI898cBWGl9kkfk+TDnrrtbIkyQMRr0olXXwsmM6FPbCN5MX
aUNH0iM1WCvFOftXYo3VsRpfdCgrXr2uFc3KBebDffhYZOXRSCqDQQ5CVD11
CrSNUHhwGBxZfh6/sL28+1r9DwIlmj9hA6wdRyDrUMrKJtEWx7Y9mOEPLziP
hoiNBPkvjbTXho6jwLQAsV3Uathy3FOm794QfKpr+t2lirid5KPpyQ43EIGK
KQMehX0r8h3NC4ECgiRMqXDAwn7RwL5BL4W2Yb8ROY51Dcn3BCS0cmh1KEQY
ObpkmYKlskQNssaLxoNXB41PifxKg7KrH6PfdUbfBYyU1+B9w/xx/ZPATmb9
Sp4b611mhcnII/im2RJpF8B6Ig+J3jcOAjQtehog+dkW0hLH6dLirIqx3DAJ
ajoyXenvRXDw/WQIvC2cxwPz6hYD2pCgVMuxm2HxKIdO9XaAN1kMq6Hb2CZW
2Vuiw/5uoQOoTBIjkOevgwK84dXNJsfUs0DvBjpGS9cASRHBbihjNnngWgor
/IY4J6UxN9DkUHnambOtwqWdr3b8hb+4Wz8Mxej2SLc3p2nNq8zFLdBVMUed
g6Kv23bJmLl3DgEOxJcT4Ucmg0ulTsTpIGJ3axdd0DF7ZPpJb+kE0H3yIg8p
dY8ZpPvcZa72j42t8y9AGi0p/ESUWaGU/WpVqzeFwmZ8Fnj0X2B8qv0rkS97
s3ns89HtsFypxCeo4+7HrCjSY2SsVmPDh+eB0EXK5nHcBPlO2U78+4shfpc1
PJuejL+FSlH9Nw87YdRqoaZz0LXMht90ddXjodXR6VoK5JdnWaXrqDc3q5Ry
ugYtw6SPvLgZfBvIcsBKyPGAN2489nQOOWAnNRv4rLF2z6CDvVDQUQX1r4C3
radhJwqfDLv1++gyRhmDO/KdnHNDCp5bO4vIRmMtizb/7lIJPVLgcfWX32uJ
OwzoDRndEEFKZ1T4ZgJslvsOjD87weTIkcwC8d8rcgzN+RS+v23Ns6ZYMXqi
obIaKYvQykThwYFPf/VwBkU6C71k7e92bX4wdPvfGZxmfVT9uk3KLbluVCoC
7nBRTlV7tE/bF9n1ES3ImPVTHEJB+foiqZmsKLZsWv3p/eb2EJgLmDjHoTy/
iqdjNiE4A/viGn5MvcB6ipITHUkH2SkHrvbYCSi3fvMlp4CevJ+2g/zMpvCC
lrYx3ijP0U5Cr1c6l5P2w8UOKGTDQwOQ+xWymr91vR84D5ISEra8Dcpe0Gw6
67WPz98TAJWDTl8M+Rluolx6MCHJFlqRcebJHQILoqMvFeQk1awJdLm6jZgd
6P0FdJQPxYduaRWcPLguUtHkoht6Ltm8HtJ6zhAeohwaWhzvWCMSwIBlNgmd
C2JTkUVqixWMSp11mZvSzhbeSekD+nAWekueGJOyjYgq4L2s0HCO3604qu06
UeaMXRjhTrEiTxnYUMmJbd3gcBp3KxlbmWaS+9xmRaQgaNk7FtIobwZKG4Oq
6rSarOW0IlZIRn/yMeLiFotcXYBFiXWnGKgKG9U+wRuQGCAATtFxy5tx1ZIc
dF2FAdNBHJVeGyn1l6dNUPK31Es/DVM1k/50m9AQ2N+shPPhv4uVXLJjGQAz
ia0FvSOeOVtSUcVxBZwcBEz2DuT0B8IxhyheN573aWT+Wc+QGsoazuJrw5YN
TH/W/ck995vv6aE2lywNpvk8LSqNUFp+70xFviOdYek6b2udHiny0R0NPKK6
SUtMF4CEFdCgC/5tD4Pwm6QwFqCke+s+kyvPRA0Ho+ZhiJ5Wd7eInGwTNSwV
6EfhuWrzigCu6Sx5SeQASuXVb6MIio8n13Hk/OGLYcRcyW/7Z86K6X3h4RyG
NTRWbRfrdhwjwv3Qt99ihT3H3KNXsDS0UGnOZ4j7OgzkkHsbuWkJCqQiBrZk
q7rxYmKENDkMGby29cFqIoNgGzlsuQGlkDDaO37yWhfiPgZoAUWk3VHv8Tmz
HJLxumolq28kfgFNHPl0Uxm+sJd4UWFvEAgg6UMFKC0Gj0DCZUnTXU4dCtOG
Hod0p4dVYa4lNezCb8nHQpEWGj9B417hMzVPdvH2zAJydEbr5Z0rs1D6xnR5
KMtRHLrire2rhKnhNFmY5f3McAs4y8/C49r3jLhz/HFysjDzu4scZc4B7Sd4
xrA6yftVlkF6H0nRB+QwL03Ufe1FvgFMLKjcTSBC2B/sOnUZAtJ477HE5QMk
4m5sEbqak1vpDHLt84UPVKanQtIk0q5WbOmacFXLYEfPL3Q2qmBPaL1iCaFs
a+1ZQ25ORJ/0bY1EHcQcSrzQLAro++VFVt5/vZ6WTu5AqRcNbdlwI9mvgWpo
wozlD0Tk+oASEGYowwGBTUpX/Wfz5GXDG2cW2GIN+vb2l2uAwIYx6eihXC++
7HSzwwgWVymtt/SNhsvmyk6/Rh7oC1HAvPlIYm7JJv1ne0tPYZbXW5kBe8da
zQ/7CMlVsghwTP5yBlbqzWtXpeC+Li/oTIF/MfXp9iGdTzuMeuA4wDLH94Wc
43NcDlB+JwCqudhPy830rKKRzz2L+F28QKXDwyStGKNDc3YD/cWeDSyVlOJU
SmsiKWNKA5iXPVPenURxupvWuH8uL57kSVwLPMv5iLiJ3p6PAiO7xfq0yLmB
Ti3QvtmAbrGby3wXSEernSC00S4XWGcPJDUJO/2N4dBthDnmYa2kf3EiwHab
KYnijVBR1gIrv+JzhMlXmYZskT8gS1Kr6UWm58/Cd75ckzfZ5mc/blvfPJoG
5SOxxfLGNtbyb8+w4EVz26pa5Lid56hoLdOH3SLKcIRD62Q8KQg1YiFcq4J8
tZeoWV82mK797MCYwqNYnAuoRNmrBtN3WCmnqCpuRbPQ7tw/TDVLYa4Xr/WF
trx6EZEQpHmZMDBBNtec+SG2UPDNdDUSYjYGuT72BCdfST5fyYQPEiYshu19
hVFDugVpPJaRxfd+kNFbYo+JzAtnClnc0Pnc+fzwCNRm9uBKQ6iCpVCsX5IS
oTL7t2L5M1yJyc+t3DtiuROhKWN9MlEd431+vDUSs/zE7JsnDy8bfQBLSuWn
0trtwPJDm5Z2aFVDp+n4vMtjcHB6Qca/3DxtVs++gEqdfnIZNsSVxK+h/i3t
Z4UcAaIdetFqG26s+DSs3936rnYS+CkCLp8heXPGalg2rCvZW1C0ALtfHebM
xGiWvZPuc7Z4ZTgHdBmgbSdEWxxlF+Resw3r9D1/182zdqMgjAs0mszP+Hsb
xaFnomoIawEhue+K3HHv8SEHeC49dZlaKa1KnpU6Y4j7MeC6eyiECLEX55cr
Iw1RWcqqbGtlZM8LYD7XgfeiwJOEfUGhWNuDZr+Q8Vik5ZjybNHaeQ35amhA
8nzB44kTra9s3vKjkVpzm3rrP1Mpg2ulqUrNwU6WM/8Zyz0AhgNSJ5ql5eOf
e01/r9iIAtGcKKrF/4I3Pq68V+Xoqy6L8PgqH7ZWi9l/+707ONOZyQhD2lTI
ZUZc8wHpDroR+HOatNHeRXJDNkL2ZGSofFbKj89geJqJbSZ23htE2Dgsc2uc
0ByvWmScjQVL13DvsotXINcSP32Srr6AGGZPfX9txzfraTlePvPBeWlfmyCO
CaOAOhM7QuJIL1TU98LR0KSc7wsiG4a4ivrTLXIWzxth5BmHsXBce9Oy2LOx
lNuFiQCQBDsXBh+rHyRjxvN4xH12ZmnOG4WJTDqDQ7OIWAYCL/cOR2obD8rB
6Wd8b4DghUcDFtzPhpiwaBRu8svSJ/MWuikqHGkXHTYQg/n+W26QjWu7zNQO
fll9G1cRkzh906p4mFiXKIf2xKqQ4Z1noHhSiHLCfkmxr6S+uppDH2R4fqWj
1TF5ba/BwTXTLWlY51dwaS4Nth8Mlhc7lb/fkEtllJt2JjqWwnwUMOk9itO5
wNk9tuaivlZ7zek2nClzfSx/LJd2j4J+9v+d7XInnym+4OoA1IqiD8sZeht3
OzlU0X5QlrnhVhM14DQLNYaX8rdUEAqs85t9xhjNuP86rBJzBepZAOfhGhRj
/T9iPDg8zAnvhWHqDqFSvNk23qYwBtzp9b6zd3yigVpyv5vVaxvTAa3eh3QJ
MRPm3G2mwIS2EW4y4jSAy0Pf0R0PoMKurf1QOudTCYEixaRzqyQjMEm75IY7
vM6RQrNaLcdnx27CCvC34qPycpuuggUcnDZuOYhM7p6Wqu5JYkqa3SFE6oyc
5WdYpwxoEapiOObz1gVZCkLtZSF0HXiaeZ/ZI0gL4Qz2J7ZDmV/ABHxhJbDi
YknJmZlKPnjHrAI47R6PtXRCC9w21hMs0hUF729r5mvcm9HXG2mQ/hSdrAj0
6v/scHOvJ/ELra+AM/lKxVz1q+sMh8R5+OUVqdVPiPYdJ62tGDR6VWcPDbU1
sP8Wl+NP9V2C/ZvHDSOxC47X64cTOyk4YJYAuceQoaMi0zctCVsuLxU4DT1j
M1ZzZ4WT+fdkR37chopr7nbUTzUKLYW7eWVVzooi9v14vkvfsRNPHKYNuTDO
OEAwTM7NbixTTCcybGuAsy/i+F02QVi6wnzJ7lqHd41LqWu2HcwY5TAQhCqV
1OkmGNYhrZsHo9syQefSoEcBc7tx3XhF/y66c/xJPxycSZ2XgmjFKPvk/ybj
iYLKta24qIEz49rZzm7iYBRZZOaqSURSsWxUvtUhH7mTRrKj71OHq2erxFIY
xLzMHMVK5IUL9ukPk2n4oj+j+Oro/pi/GzteCHR+F7oRa7bUsQ85V6MrMVkv
sm5CeUCHLY5dDKzG704FYNE/z7QrinEj8m1nZcYvIsRBdLzhUVSktvQS1EdX
gLwFOzXz8arQe3b4PCcs/R2SwT1N3hYvq8va2TmQWXBu/ASjHO5wclEwXlrC
tjrYs9bl6sYBmOU+lDkliOgGeJCv3a67MrJpW7KAgak43W47HpRu53wSR+iF
Xx0NW24fBDTsywigPsOSgbWqD6QjAIRUqcZ5oiFksQar0UIzUEQzqNy3cvU+
W574SYzodpIMlKggGOBvgrBerNlm2HqjYxyfWABTG7pymV2sCEsr4Li7JRrv
aJVzG+V+LKbdvHjf5+HmIFkuxKByOFH2qnWNcIWg0A9FgHeHZea4csnJrKfF
BD/3ykb4bYIgBZcPwB3bL8EvxgZXfmaCy8l9hmCm5ylPXcrZn88Li7dnBnz5
tFEaxCYCekBh1y144em+5M1z22zxNc7Ls81qe1HIO5hN7Ok7Np5FPoSolVX9
YMD2jS9Tdt6bZI3xZjNkHaVlYaXzDCTsiRVNVWp6ZSGYp34bkLK09989soET
/az/S0hly79Hrv3sfrC7BqzJmJ6NOUldKlP3vGxo7S4uVliqkG7FRTEvlzbs
XZ5xKPem65b57kC9rdHwfgq4XqFQJ6VLTGTqX7zHEGXdcMdAtZRE2foj2qW5
SRiD5Yj5oX2IOBNvXKDvJInPzeBN0Iw+9gtTp/aOwUosLR51wa12kA5Ot7ff
gUUaxP2LKoQu49797m7kf92dmWmzaX6fB9Oh6J6I4Jy8ohPlblSo1xRBQcX0
JqPSxPRJ+H6iupq4Wwgri/Gtuy1C1JFYvBoxJN66mRBlemvy5VQ9ckAI7GeL
YneGnkcIaN68kOmrbODaReiidEf3i76rGnQmBFkl/QoTBhFnyXgw18yRTahK
muNdGIF7t4+GU5Y3oo2YXDbFAv8fzbSJ50QUr11+Z0OEGqj6Ppp9Hhgd3q8r
9eau6CCHhFCHkM+Zug5Vm14NuQX66cNdDKtxlQ94i6bsgVLG1rkBEQH8QQJD
rlBhvtPLZzUHpvNizX7XoBGmS6Ms/SiuV7XaOxgfR0LaQ5fULo9IoPZPKMUE
Z3otiDOqIibKuDwc/+kzdUWy4OxNotkN018Fl6yaR2cLc9XVFg3c1YWr7CiO
pcoXbSvGVDjTRL4daR4HQjdo91qnJ397GLOJkpKvISOvbiRi67jeNLBi01u3
RBEBtmOdkw+4q/KID0f2Q0+mw1hENWrwPa10ckyYYvn+qE+d1/4u+AzTMESX
EY1/5gu7Jou2GKBbpa7yYeZiEmtLiwdxLC/3KhfiPA2cVUDEsztkvYmHdIll
Y0RWNhq0ElBO9WgTtAwG+RRWA8ZXLOafhzyUiG0ryKZX6LL+LBQwq5q7pArJ
xu/aWQ3ZXiv9/MqAzU/aa2wuueKlc010iU0tia3vhNfjsyBflr1N/Oks6DL+
lqkuYnv4y+ZvTmkyGQbT5fpXfoFg5obPQu6qgV7FBK7HyOrNW7oZDay2LfD+
1b9W7EmyDovvj8jcebhKfvPTDHsfQ5mtCO7/lFe7RyWeRxTTlNilcBo2LTpV
HROYFNYzE7t4fg+FN9m5tiqSYSKVZbEeWaXSaTTaWHm8Fcu+bT/n359/+WSX
Rv7P52Ka3YrUG5eU2YNZWvMwDKDVHaYu3uZXDGoS3sTtI99LHknqnWwI46oz
2VeI+p2e9eJopqTqAnoRUJzgRvKGC7H+JrQfsYIx+AhhCBnElJPQ1aWDixy3
5YOhLILzxIeUT369FUXliJfu0LWPiuOS3R6q44kAtJHhmS1m6o5sIB5DvjSE
903mXb0Rjp4DHgVL4Q09pmkch8G4vKIx/lVFOdLNaNKCLXnIYSPwc6H5TJRg
y0nteQ7ssQ8Q71OvzuERcpFSxqwv7JI702XzRFmv896uy6RJ02aYkqV405D0
qvnH1JRWuKjb/yjW0J6aQvVTnSfR0qJweGrEp+1SAZ+gkT2YYHXbrchjAjbJ
3xYuj0EghmO6rXwkrgaAbG9ubAD0HkfjY0fTF7m+fBVDU/+rr/rv3/bTIQAP
v80tO2yUtmQ+Y0vcE1/T0UOlaU9sXEhI/qiQOY3R4a7yMwNACi9z5WHKtuid
8MsBK+Dp2IvhuBRcX1iFdMKn1MFRmjybHSrQp86NCbr8If02/isYEA5cnBT8
Jg8srvhtcHwnisb6QTnS0kBexMV7zyVWRHz2jfOhRDveMzT80orvoe+6Ri1s
KKz/AtXYXeRzL06pnFjy4aQSMe9nQs4wRvJp6BF2OALFqp28Gdd0mDi3DbE3
dXo7YV9lLQU6o61m4yT+aamgpoe5pvgpDLJmWKVounfzhvESRe/Uey6C9iz/
xHwG3EKeoFcQ/uskUTX3Kc5slt8M/02c6FTHfy+enyIrYUkcRwduBbrsXDW6
1Scjx2kzH8LPmV+uxV7qCP4Wfx7KzcnqwI5lMwXKYnqulqRafWfz+7E/fn6H
b5GdyPxhVmKnvDVHBoGhn7T5uWovW5U2yjKWmprqyOc+l39/VpVHGJ8NrUxK
Ych3YZ2ZxJAP1hiU4kBJ0S/pXkBkkfQyiWGhDfO2VkK4n2LcgkT+zYKYdpoF
DMz9G/jHwFQOJalnnvOB50Lpven9IoHZZu0zMhqgZedGwqe7faBq8SqNNo5v
JqEyP931Yjplj4s4rJ0+8xYkJGLAPPVvz1uHfhcMteh2OgKP7KSonD7iHDNL
/bBPk8f/S3SL5L1hHdpTNAmBE+Y0vennSV2ebmQwRtep+Q+tRmyXtCpjYflS
8XFo3uKlbmDa9OlJhXNXPck/oyJqljyDNupUXxW1wNfJvuNL41DCMVCbGT2R
Glpf/5gPa+B/HvRoX+JXExhdNaHj2sh1+vRqLX7CfZC9G40lbyJr8SuI+JsW
X78uGwayPZDFy/r7eWLBcCHtGpFpwnhh1FIZpl1QXpEEf76Qt9daz6tinIYP
0PzMMuAaEMW6xFHA/IS/8aZFhgAVU8zXvMbRDN8MmCdyIiOvVg2c9SfVgr1m
FnYBwRNj9AR0q7rOMy8txPD0WXXYfEWfqZlQ8xZvI2FmPaudexjWXPV14aqT
twoLIlfLtQdwFHiL/3Kxp54tFyYhrDMx52B9dDcwiLA0KkfS4pSTOeNgOzeZ
nGxVqSpabYlQWLHjlVjH33mt60mXqqkBRNQlKUZsjbpbVFKF/yaNKQ13jctL
3haaFkMhXVD+ZzoXTgMYsS13DiPQKJ8qzA+Xvt1jo9LBuVmGkrSyZVVQZwYp
Pb2jCeTlDJxLBr++DR9ksDEAcmeKFnQnd2gfwrV4ZLWocesWgJXtTbth4nUt
EKXiFwIqaCp+yGW2wq2fYl87R6jk5eBVEqqSFCXffOL2BcUJzMEMlGjwXXEd
7O768ktUe6qT/q4fg7KtLCxPijb6WO8qkOw9+gKxSGzI8FFOtL3BT5/Nfwar
YWmdr3De7TED6GnLpNBIwxZqKeih+pZSYM5G1aq4+WNbmlaoYx3NmG1KdX9U
T6xP1iDxkwJt0oituwAaNPQvDNJq+X0AL+gNiCmPHUJrQrpA0T0UJsoIT2uw
LoftgJv1T/U5kgadic/Zy4we/wEKnDZQocOvqKV2MsLiQqAhTyfdnBDXYCe5
ZRvzFduU7/PaOth8TzJfW2eTO7gXwa2Lenb69vcS1HJJ5ULQ3jMwzoCgBD+N
RKH3bw3VopBaq7RJx4abBbV+Jz7nkV8f6mE0B7WlkQd9zIJCAfZ5Fp6hiyKx
khAM/fdw2obe5faKpnXHB50fg4TecF68AQ6C4mBASrwRlj6/Tb/AD0qt2eNP
dq6OxHd+6bV+RLomdBlKLYO5uPtbtqpFyaVa6oIF7rBP3p5RS1xoYlv+QTS+
CoSCqfWgYPbKyhra6dIY/gHFbTLDCqNEf+5A4mdCQxydGk0+cK+Q8WIA0RVy
yn4Zq5MuHxu2/8f1Q8cLAuzCDqdCNi4d5iyxXTyBRXv1QcqN/7ecu1r5hnzs
N3ssQa6ZbL4rAdWCO0zd0lTnpU+G9chOoP5SzblYW2lAoo8m6emQg8pGusVi
06w1/iBmZm7aZfI5QEG1pFenezB7jdlr8mXOmLu/nlakZl0AILydu5+nBXVp
8WTBRjdie2k1VVphqWIW7I7ZCXTp8JZtDTxJ1jbF8s3wYk1ZqV6ElDz8vy2t
PlASDMcyy8unOjRgkkDN6aDacg/4Ry7xHFiLSTT7s5EjWVqTMXkh39T6rIgG
Pst3FecWPqLvxx4UnZNDHQa4yTepGXG/pEsBRG7rV8zNr8gboJ7AAzb5wQMe
Q2UJAeqZbriia30j1/sBD4LYdM8/2MoXPVh+ghLNwacfhbstfT7Ourfel9ux
AUvVA9I5n+6jtt0CnWnMYCU5vMF1I+pyPOxbBR3+ELInERs45AuwclooLePO
IMVZlyWh2eyqtvG0lX/CKdMrY2P26sAuXM2DZoUY7b44jSwjnzdQYPF7abJA
2M/iM61mm+TgoJJk+2ZhIyYW7BrlAOVOGS4umUk2YzfKoAGkhxWu41ErU1/X
eF72z1z39eA7GWmm4keP/sWpdMNX5Jr8Ek1xtQT0oWB64ouxnZBozlZygYbj
kjuqsbh31ZF2xfA8iZT2R76Sp/CQ/1qTzug7in0uE/1Hib+ezfa157mCf3Qz
w7MjUS46EJ0BmFswrUIRdSfH/bjBtaasJ/b5v3ZOz5M5Hbswt/M60JqARKmw
89chVng1z1viacbZ6O3kyBz51c9lYkCWxbvmHW92/MX+DfCXfrX6YiyEAqPh
9oH1khGZFQQTLy5xZgEvJrHo+eqTsUPbE/WmTF2HXeTPK9E+T1fzpivAsKTk
CWWYs+WrrzU43feDQFsSUJlmcbxHz+pEpE6LgHAUD3EB08Rw2p7Yv8HUMCIu
eRMWB2noBbODol6Md8IVps3dgXij2dPDaz7Ye2HL+xzQ8CDWP+pQdW8rUjQk
ymduKLzri86KqM/9EtgXtq8pS6QEKyUYDOFb+a6EoMDcIcPXoaT5Q3otH550
dNTw6YoAFHw1A1EUdBRvitGd+x4+4sihGfoznb/IgmZ6EulC6oIAaNQnUCw/
ehtKTruoQM+OCEkeRw41ww51jPRobhiKDpKnsy8Hz+Jo56doy0eoJcrYotsa
ewXCjp1LO0gotCfXWnVXUDPk1E22fEcbQXz2AZmMBWvoH0EUeA6NCaCfJoG5
RwMdxOMIJgCHgH2nxrVq2XrmkJ4aXrHjopvlP44DniNaqCLF+LZ0Edvolook
GRuxVKxP6Dc0hflOZBRfjxSZXhJ69BIqzcH+aaMcqzV8ciKVUOpdEzQ9VDov
B/lfwHLKT4rzyexaiWyQgi9KCtEJidBb2eCpiMSuVAWPrDjEGLt0X+CZfJ1J
L2at17gE4Bd8UCByUnMMsUy2RA81l29j86uQRvtyBpQZPn8Cq1XqRHTCY10M
RDtlFiXU09HcgKES0QqmOD8fp50T2sAEGElG1ghodmG0ni4c1M105Bb/rIaR
LV4PPBJZRox8W9huZ96TsjQUhSdhs+hVBj7RuE1i21smdjvucIUIiT42j8FT
aNSWJgfGyosIZGzHMWuVkAMhUxSgARDqWQpgX2+HBPsytMJoqMCTJp3m/0me
M+uX9EeeG40zJu23EkpyJNOypvYAeuXu8EyEvyjamFf/zIBhwr4R3tYy0BDG
zNEKjWFAvfSG6ytB+8xzA99dv8PzeWF2fpkHuinceHREcHy5be32qkjJIrLV
TIt2z4YHDrVmF0e30NZvY2ZiTNZyDf25VjeuKIRhoPUgFQUm/J/CViN6plqA
3f54/ZTGTzy5KZEws89TQ72iBvDct9VNKNHL1jyOn+NYRyaLX3fXEnOWeIPL
+zRhWcuVQdsxjMwF4T7WW6Tm2JoQFiDFgkQbfq8ivo7fdKPKpjb9Oss9UN9H
OVoY11KhhJo97mxaERHG+Xks8VxXtHSpa546MOcOthtMVjq/LXXyA3a8lERG
bXxQSM6g+IuGwj1t4Y3v1DfXKhx20+SN0JhOONftWIPITKcz+k1ztrFFi8NM
37iz0eDntR2Tqzr6374c286Dkih9ULW57pMCZe0Ojmk9Xwy43AbxJnphzxLM
x2cQ9iSM1x94t44TyFquf0RTRgowIpGhDXh+LPZlAOnlzBDSXmPPy60b7stR
u3wIpzci++YNO+qLRBABQ1/36L/GnQNBT9zrsUQiDfFbZXRRxD1Z0vdzSv74
8w+Qhj1FHcqXM8d/behsEfuz3DRIbC14fY9R71mY3Mrk+zP6aWo+8QYW0QJD
ltMZmSXblOZQ3siOVsc54XfT4un+Xld/gEMwBQANXsipIhWaw4P72P5R34OV
kx/DMxyg3LWbaHGbdQuzCZDOomDAd8CFpGWgndP943R31NTOYFK7Pt5ntAuX
4snuvVPWAUeUPLCrwFN9eRQlFvjVHNPYs1ZmZKLZo5z7ZkW4IMeNmH9y5drq
eucBETWlgGZ12xgF/oNlhD17RlODweD9HaXllDwYoVr+yP5H43QgN8pQmutY
iGTi2wBYBv6xe8K8rqUvEsEPjnWEvEjOnguRIypiA/z3uITabGiEOxMmtQAG
HCoHDW7khumwi6ALBqQKstEDOJysUXFtJ//lw0gO2imcn12RU6+sII79m+ni
0hF66qCvgiZe20gREq2uqCJ5tN3cwe2rFSkGr2RNVddstAAyiJOfENpNwy1p
fPBA0lu0Ig/vz6UN1gW2ErVxfOpQ8mIHfCJ0lcJs4Rb3kZEDw9vexCKKlYUZ
hrEG+ZN4mu8XxiRNGrgFj+Er5xpoqDabim8yK0XBQ37SqUPJQzpuyeseb5zm
1KqHRaq0K5QAlT1a1X1N6cChYbVbaQQ2kMZSciGNOXnU3pa8czT4ShJ5T1xE
N/5jGoFCKWvIb3av1pPTfzWe8h9mG0wkFvcFnepI0s243TL4q55B1fyZlI/e
sa3ZnkkDRMw9/vanAzZj2TxivgWB2UXfV2fC3pAOTcE+C1IPAU8tU8ztrSQJ
CmuLtrnaGYLcREK12+jU5NQByHpGtms82jDgkIE7mhU0TBPFIR4aMlC88839
OeCyYJO0XjllIkGTu/6f/NW5k+4VjQyxQpaJCrL8Ad5oQaVMewh5GRzmyItB
tz2O7TOp0jBstFuIa0Bc3aej6F+e8t6YY+l8P6IqfjcPIanZywg1AxI4TaKS
iPxHBpX17DZ6JKHx2MQ5VAklFswgiUpuPQPUYZUn9KGnrazsH5Cga2iUWAL7
/O8W7Zq9OgkaaVJmJg8X0TG4XIGdr9udB1w4ltJs2kOhVJnneLO4Id4HQgsx
TujkV9VpbCOeYx0B22x9S/qnJk26yoh+OeJZ0I9M8k4bjLMZLp/LB0kdoTYi
Tv3xNVL97DYS3FRA2jargIRExrz4DDWuX/82Z/HhJib9nls/qRXpGUnsll7e
NYQfsX+/6KJOC4lcYpUNYXMLY7x6pGBqvuyNwglNNruOJJRNHF+cnhDtKEG7
ZV7h2ij7VMYyMUzw3cVzgdwj9yiQMtTvpsRYwR9iNKE1U4/alWWgAk24T2HP
GhK0M0Y/Q3UOuXsmQj9e2dmi4ispR4uriioeMqOm9H/uv6eO8nHqmqT28ZT9
WZiDKdkBBME4vmG55thvgds+hxH9WDDyCucXhoM9+4qgnvxmXfz9BN2n7K5K
1jiF3+cqf7PL2iU2ZmBQPXqxAUQacF6MG/5lNbMoBY/qr3+ZGf55MLXqlO6X
KmEc71+g8noLjp2R2rE4/fBqiAO9pATK56yuZlCvj17sijV6/8fLn0Ijge+I
1TvSBFWhY7atYZiHC59WQuMAT9pmZF+qcidSas0Mn0A7dnUr3odxA9K/ENHr
gUbJSsSnZqaXQCQf+oOXdGT1JTzQJpA7zzLYYzVKcyimf/S38fFv9nUM+E5L
q/KzKMPc7ri7me5C9gPiTrgs+Gn+uaMy/p2O7iLjqylUm8wunEOWmHDQt5Tu
5pRJEdvwn2DyeuEcKb95Zwy9t0ulk9FIdoYK8mzFQE8I7bxz90pOPaxAdzzX
YgzVTv8onoHv+GMsF0rYrQQxypuw4DO7++wADSXN7Vhz8ZKXmDgzYvYN9YMv
jZpDOC7aqu8YGLIi2LYYlE2T0dRhqxhfiQeUzkK4fzFP/60xe8SHkLtGAsUW
7NY6JfUU9UeBv2XHJwDLW7GJDeqKzf+ZIt9EVHKBwCpMFhmEgi6Mz/0Jcq89
3PGOG+Pt1+CFI1naRpePmqhvy6QjYWj59o1bgmAn3WMv+a88DfmeKIsbT04n
JPWIFVRoUwrATH/X4ojX7YIP8JmB9nTx9o8FXUGE8q54laecGxWtJoIq3T7D
RaW4vfUK7G347KoeTUj/e/MyIM382FyA2PHLfXvemWCb8+t0p0AWVF//+DS9
xJREbku9mQnJvCrEsBChqGJwxqsaNTIc9yGnARFT1EoU73yC1SMptFZz2exU
bqJwGLSfJkXzw/eLbOr1hkZoA9S1EfgZ22p3e+tA1xRb09M0Wa1tlRKLaQPq
bGL7sQlf+CL1JJh/3Kx9qfOV1RKV3mb1nwBZPSwYyoM6rAEdUn/Gjx3lNrV8
h4M1yLkWnmwg7JXIPMxliKx6YUunU9gVVVJONGujEjoezLzMzgVRfU1cFfr/
NQ+jb3AECvg52BIwl8QyD1YMTLtyjMe/7mPvQbCoJrv/t+xLjBiCpCyrUhvH
2cbfqRksQg0NgBoFmJcV3VvT80AIPIsgN7ARkHUc3hhchiBaIIW9YinzmfEh
r6gS62BkdwvS64wpptm/Fes7N3SbjvlHQtJSweCSZ1akoXa/ngycgGcRAvmr
DkqNd3PhmsgjSdZ1NXC+4maIUnFPtllPIwwISTdf+WBTp0dBVbFhzFYl5fZw
PaA+hvg+vkvKDrlDc/xCvqdohkCD7naxQhyQDKw0iUjlemx4RKVrUaZHI5Ui
TIf0THRQ3A6KuZxO7kMMqOgAzGe5upx+27S2QyZkD8dwLvt+Rz8gTnn+H7Vy
f1tTK2qNl8G0axJXZI/fnGrt1eZQnzNtRIMOAQW0lNdXbckGFzx4mLqSRl+Z
XVhQT72n4OeUVpukt2n7TpkquqNNgm7aAUAqpAFsbtI8CPjlJR660JzaEH1S
u5LttJf/EBtF8AD+L7ySsoEN5VTykrjed8khEDIiLAFJoE8ro2/E67UGkrCu
r+JSE/D8KF4nmWUblTdVxULIqWKbcUXpGrB8Vxkgcokgz6qaVNnfBSDomTW5
6B+OPmCUxstc0RLDh2NowJxQUem/zNor3Txrdd/Cc6RHVTywXK3tTsWulWJE
43ELAc6uKvvUVRXXJYumzZIvjW7KsD2DUrfXOgjUAY9JunbqzZJE5BN+Fm1U
OQAAtl5Hv+uUsFYTg3p6tCGasqpNi9FS+3Zw/E7d9TSXpYGzrAT3dVCfUz7L
8wg+EnTSrWYXRiPk6oxoq7W01F5HEvzAa/Rt5BK3obg6Iik3NNYzQSKEW2Ie
hBUPxWBHdUcpxe7TUrmYy+gy9DYkyPyoh2RFLTib2RICl3h0wZrpMa86RxIN
pMJ9VkPJidMOqefdgqqaQ4Pq44mPWmkyl/i6dBt7bxK3iqYzvHmfwNIj9jGu
N7ELempwVb71NwUqK2SemE7e9gADItYZRtUrUlRGo8Tm+w8WJrPJuoo9VQ2m
EWHHet6efeDtwKZzNNEJXcDwge8QHQW/i4xL+vdvsU9rD8c57oh84OP4srzX
XWY3t+4ndQ5U6yl/Cz5n1GaWtnvcAvZAJclV3Vllm11VMsq2BgUAIwEhjdbu
UDxOaDgIvQzE/c1NxpAYiD0XpIDVPsw93vi5J8EjB3I9DrNhIbrRZZuZO2J0
w865DwzPPYxhS+i5sq7hjxKD2FzBFiVX7XavoEMwrZnT23bDmCLhoWlCyUP3
WQaNs3LmJMQuN1GyiuyCdFe7uaybKJWUdQNFzG78N1GkIWud6BXk3ATUX5Sr
LQI29iOgKvLbS6162+cmHokwZldGJF0irAerJAoi0zKuX+lOskL3rVitQtv/
533a5gLXAmGd8sss/tOWTtXZlXt7IMUuL/ELiXctDTOk25wOYGT82QELvKQb
Uhv1KdDBJAWQehExsaDNWz88wegqY7Ex58hM9WlpGGQ9DybBpK5BtA4QvKmL
HfXVwtlAzSjm3o6W9BBFTMcrCbkhf5g4LltMrJhEWj1ikhViaimFWBWcSfxF
jbx4nZQe0um4bhUpknMr9GsHbIMuNArrw8iSY5gm91d5OGm5McDqp7V56xO1
GNvXYwUUSN4s1l1zu8MKO9jTvFSiFrz/sYDnddBxOwYS9l2RYNd8JG+iblnL
7doDZfitJ4PcMW/a4ZiO+RFHpmcDy1E8fuWPswx/GSdgIsABeO/284qPqEUJ
joeWPaLNs73MEBuJnqyOLZfn2Sm/R9NioTJYF0PLBdnUkqaPhOw6eZFLW+vD
HlhZ8WVXu5bnd0e7XNeHF4mBEtt1EbbpHsRN1EdVAFjiYKluBSpPNf1OCabV
56zsup/3NUxzMdxjXp5H9xq0d356aVM/K3rqYikVW3L0IgVJAiCrwW8qFG1X
KkicK172Rb/8ww6Jr5Z/4Lq4xpsPSFB51AWc5GuHVhOVqMElpMPcfnzl9Px7
l9SoNzqagTUsEYcX154KxT+PMQRVSJ4y/ZUcK19UbKXwjK54QdkgFaQUrEBp
EL5FQupzXOCIQB1xtbzyalrN0H07yUcuf0ssq70d/m4i1Upucl+qJSW/rP26
Voj3O49DxX6Nw76y2EpFNdnN3dbeol2P6FP1yg8/zneF7oKONrKvs2VGpPCg
h9G8NbE1wfLvhA23mql8Bm/zGsg7mkCK1YK2/JBZO09r+NLjbCrjRGPVToyB
0IqZmyz/3G5L8FoGZnqsowvAGzjsZq7bsrMRD7swuqi42Dg5uIGMWMC6No0z
t0pqd8NNq3ld3szxEshSpJXsZg5DzSNCV0Bjch/L0XMJJ7qprGC8Lya7XmVM
vTPcvWu0qa01TjXGherb5hadmzPTZoEBwl+NlOHcQCk92kNwqYa0M1J/oCqf
bNbrxiui5PIBucw+49GfC85k1ZrYSOdEGCDBWrlUDqK2jcpjxGCEnqwy0G5l
HKAO2YCAz47N8iPEtCWUyJ46qVU3G42Ebn1DnzyAuKTdXo2faOxH9CLDTAd2
rAAN0B8/MKbcNzP4fSnZzylPA+PV4G0at4ukLTvNqELjy/S6Qs03SZsMSOTo
otBu2K6pD22RE8QaTPso8JPZrCLUqYmLZ+uV0U5ppTmXj/dY1erIUdG2BACF
sLZSOu0ESMAyELaMf5ZQm8zQ7GyTeeo4D2tqSXDtAbBPFHLIEj0JFMN8XdD9
As8J/JxyuhNLQK4fKH7XpW+VUGFtJGaYmA+trM5I2lOyjB3IiO2u3OEQlL2k
+0NqeJlEp/nauPMQAIyB+T50K5krbKsxcjzQLXWeaSIiVZtkZgfw1YTgDHjF
mSIlN8wFjFQZq2axAgApw1GVB73JU10w9qWs9HRvT2meokKCwjVEuQ6p1hkA
RSL+wAKzU8lgKq/WOO/w+Zj23vRJ7LnlhHKEUZ3yJ78VsVHIw8PMyDlr1XM6
OWiIBvtKbkDWA79QzjjX3E53jAUMtdbl+kLLR9JvOriTPL/BU3ZfNVngn1wZ
kTNlOtQ7NcdWfKQ3EuMMwpIMELkafuJ4eVhWJPQb+majQWvzW2DFDlTINU0a
2C+KZrvuRZARDbt7K8Et9dUFFGBKt6BnvNJlt3RfsHA51v0ORuFv5w9YJNjO
vxeS27PebfZLbh5Lg1H0T/Veh+Zdqx23VMZV3Y3/rNPWBT/TVdyIaGBK8rH2
ibTTciT08UGcd3HRdm4Iu9jU1b7jN/yhjNtAwz9gGxzLtrQojSuAvrPF12Qz
ZZjrS0S2PMLbF8eMyI4Rxpx5XjxZWTiiOatQuQdtiaywRIFpPMQZ8Q3mlVIq
f1Oj+UOS9U8+jg1dXMQswTy1HlVnSjCesgG9I+7zZaV6op/RLGJyu9/2mOJZ
Z9pxNsXHfeMahbrEdgKkx8tvg6lNqkf1AulysVUdOJvGmSnhv2BEvkD3HatH
WN6fWs+Cgpo1U6E2HeFd9wpzfsaykjHmfkd+/T0Re1SAFHNAhNS0PlUKd3Tt
tYvOB8s5jVFzXJkU3TopyO6jG2MVclEdDGXlpXPiItrhksD15ZM/vbQMSW4j
n3OJsLM9/+QVY3cSeGYeHYNHMFiiBi5EgCrG/oVi7uS3hkt4phCSaAbbLa5i
hVrLWEASURz1dvq/GMIp6BTH/afyOmtFqlPHTx7miBE/jZf6eF3b5SaUr/tS
Hc2zdxB2JWCrMh9aTM4ryKgWq6tWl+QmrtFCcH0F2Klom2ivI+3InJzl2qzW
GtFZeH3Wbjp5EyFkRWwdF7B7VtZCla2FcVex0Ye/JE7US/SQ1JwUlOanjt6L
4x2IaZSnniXwWrf9EYiqbMlr27e7yMo5n7QvwYnhDU8uc+WkbMHTSPutbCGK
kCJHblHBdyQmGY5MUoWx330QJpQ8ZDezkLUkCaL9M5sCmiarXWarZyWmcxh2
ZqmnJg2+fN21uivENdNHcNG0JSgyiINDvU8N7PSdexk37wZ9kdntzSuMLSY5
ZK+JCZ2lvwnU2gHSCTLrmqV+lD+B6F96x17tx9et/EeWUgl/zfE1rAosmafO
FFGT0vmYGJWZW9zuSYOvq4Q7uVkuDbgJg7Zv5XrKfrK9FlIp8aiUnmcdnke8
meIxmfAntNzMGDDxSIVthbNI5SJ2qB58D5t2MAy7+t9SilPTiqKhEPzlBy6I
bRqS9teVP6ZpA6jtipx99ZPnwZdjHj8e05DJ13Pjz/hhkGlpX4bqyX7JruJ6
BSOCwYNs8r46r6DxRqAqlUGYkUuwBUIFaDqDmZ6uwHEn1RJi15YDzEsrfvt5
yjBQUnynQDrBiUU6BitJfXS9uOmR0p8Ne29q9qA5Hg5WVTGNMUeJ7ZoCPDgO
AOlKSdUYt/PjIbDU7VFCsFW576z2On9uKFvf40ecr0YTfaTo7nQS5+2PLV4h
kP9Nnzir3HBpAUvu3u1JUAnDXMsuhDBeADodSp5ub0siTzZtpPKcjuxb9L/Q
N1UftXmbedpACiSvWWhPp9xovlRONJQCcM793QQD7B2egvyUh+YYCgjhSGWm
qzalb8saf8cB/eO1dBKLj+yK28wizZKCWywHWNI/V5Whl+MvI4YuI+776XEs
HU8BQVjdLPhTed7W1//GdBlzO1mtVF+6kIDlkLkGifDuusa+qCWNqEGw53T/
30ORjpo2RqR4w1L1iHmjPDLT3CBiUZdPAorU2OV3fau6Mt6YBFZU6vmCjCcC
nwK0v3QHuWJ63LTbREEZAnph7qK/tXkpGSOmT1++n37uyHZ3N/amB+MYL355
YLNSrwSIpnl/SlF7++AJzwvFzYDusiC+AhnL5NxlseP7fTBafs8z1q9vxidL
mxL1/o8Zu3P2Ks/Llq/fbFZPgV2v1Czw6fUh9fxVxZ3cO+Fg6HxKoSRnkhsw
X/yO9t/K/Aa9+P+gqOna9mQkTxp0rKXh4jvyWkHKuANxCx/2QFB3kiYIM6bz
+xTGIrq/iYMbzvjHPdpAIzOULHjg0KxfALRo3xyHlEH4XOHMpGsGR3AbQBMh
BS+PQKiidJbkC5Aww3gwx9CwGOTk1g4mSieHTmhNCSQQYVhNOFlLwqwFZQnX
qsv4jrtus6XEZJDoQrhqkX9WcSmYfEQQmuQJaqwdcQGQEJMJ79Sf8J49DFKX
V2N8suc3h5YCaD333B2jfFBlP7DYWkBSuVaxGZpjdsPSBhA+bugiLpyLVatH
+/MAn4FqFo7phIp4YR9O/pF3O+bNjeE/po7K2U8Zy9pmmbrY8n9uhcm9rz2s
puY+ku2BBm+LJKOw9F9b9t3OZ9tQa4b509nAG50XVE9ijHfSgYT/2hOP1Vv5
w5/EXrSeN3wkiZ8914XmAgdOCyMn9Uydec0Suq68BFVg5cJaj6LkY+10pCUc
kGilVlKaa2QcaHDlsxrHIFec+tP/IFUsxZ8Jx/wyJ7CJeRj2mIfnXEq0K8VL
q3sIVLnJC1zx9EV7UPElqgXP82gTaIaeK4FqNPAicFwUDyKqAMI1JoJql3An
OgnCxfBs4ySIdJiFO5XFZSV0fk30P/FJMm4g0+Q0lzmVBzSIS1JN+6ILQhq5
o6dqk4GFBzoUH2yHKJZmYBdyJ0TUu6BeA2uTRFHyuHqZhzmd5sT7E0NsNA4V
8RC2IXSrwLV0FgVAp0IFTg7oZBL170HPllAay/nxGWwEffwn12z4eWsvRwLk
X7RUeF84cB9yZczsid31IHgaVDs/MZgvAoQtjW1jGpH9UWpR5SCW793G6Ok6
j9Xv+aLgPoyp5hOEPIzIF/fTvtxlg+fY9VyjY2dzlEt06v9N1EMe6xxQGqRr
QDFIjmAAfWnE4qsdYupmVj5PR872WcpVF+51ytaEGeFhB9mNIYjIpg/GcRIO
GudBjF94siWtawxcGH+06BFEaXa5ZSPFPpXdRjEt/NmuW64V1SAPL7VKt2IS
Gtqgutz6NOC7LrKCtwfplS/EYm6Ul9A16SzuukFryZdUVNHXpeyQIsXpv0cl
YD1zpsJJmIg/0DTxrZZopmc9/kYV6aJqCJIKihnLRtJhSUygNHTVcRmzdsDH
waSK4+InOpOEy+WKfoDZRtXGgS7TcmDZRNSpRgJSzpLEA9luanDpbGJ0VXxb
If5Wd6koymKotCue2yXcUDXWjd5QYuCuMzeZVshsCbWIOREMdiT3bdbJZtu5
jAwloQZKUpqBU6b/vU/b9NTIk6Lsj7oer43KoVP7fRNpkYfiwQFSGo33Ah/C
nMglLPQaQM1UCvCF/NWp85/cXWnFAzeu04f4PG6njI/RSsJsfVbF8e5mSIGR
lYjvm/Itb/bg4SE5RowF4YayIkvkxZlBH6BxYz1MH2aSn1opw1jMQ63MDFYo
oKLvybWSflNoJYgnTkn1KGc02nMwYVu7k0AJ9lIAiCahIf9HmxQjXID8Lrbl
TgazahI5c3lENeyXa7xiYaupMUCfu1IoHSBXRGC08dcjv90dgam3ijXSdtc6
sGl+DK9w1Xuutx/cAwn/sTsaYXX0VJbEOqGUwA+P+3+EZC+BGXQSjkE4siHh
l0UKWPAWHKa8MjtbHUaxtCbz8Z8Kiw13pqbPaCh7t7dpRrunlrfN+xeCa5Ad
hv0MrNbhdnzjbKr3dIu5gGnhMjy3YUO5Uj74YEZNSkjueYfrvd1Z2yl8Ygg7
fKXYrv1kzJS/wZqrnXmX9dVFiNPCx8ujaOXYSYSc00i0D9AVJ85P0u/aoeDi
JzI/hzyCE+wAWiGFedZ6JPNj2F9MF1O64LaN/wc4nM68Spt4QrDwr1uIfsk+
TCjG9d4XnQd2jxGRVxD2wlubdrSk6x2cTUsBlc7f+5BGsG5SIn954bksa/rs
rGojs8h5wdU6zZqnhxg9dEiSMRpW7K1pK5WBduomQI875PPken3YOlI7bew7
kYU+/XzdpH/j4zLG487kHXzIWaLZe82hMjgVdBfpY+vs7XAXI4UUaXAYoP1v
rTkqBYJJEj02RMioDNo2E9mcnPQhRjaI/2JQcvLM3AGBcs6FIbL6rhFivN6M
tgYTBoOfCHiN9x8oyDNMf9PLfHC8UqN+ttYsIBBYyjV0dyUOrSPndaJ1IztE
JWk/0epU+/4QCkseN30qwhiyghRC8z1IrMI4aNauZ3xClF/3+xngo8bvHhmo
TkqJoxlHKl9CgxkGuxdU1RjLjO+xg65Fdcd2IfQRyMUyGOQZQLBoUtF/b+EW
N2Y60D2Nk+hWJdPqeBfnlO2brAakIZqpw2VZuoEF2nWbuwbcitdXrNHBv4p6
h9b6yb8qzYoP0KbrZydAf/rIpEuUG+Lg2ZPvoj4Z189LkPqYI4p0pJKxzvNi
LnZiQIWqcTHd3TqoGEO2frszm0C3UZQZjJ3yH5dTvun/kFGIW2i6Ot6kh/Tk
cehgDv1GmuVtEmRuLdedorKio2h8KT/CMWLTS7aXvFyzFRD5Q1ubwfCfT9qy
joCxmfyLPAFV9PCJBtkgnf8V7Fs9KTlzluP2dePanXGqQIATMFqce1sF8eg/
OymSX5RERn7xtYMsZkd/bizcANIc2YP1wjTpZsWRD5SvzGrARqHKHW9Ah3qR
jKpM6RIeLO2Ae0XGNFdLSf2LusjDvb/syeiA1Tj+2yMc5Gruhx77eV+Kl56G
bB0scotw+V+nL1UiCbEcTBWwZJ4mWlbYjZC3h8HyGLRneSGzQdvODYnwB5vo
C5hUDggdmK7zEkHAGQGR+SKHLjPRnFdFGrYbwt+MogoX4kvayieY9cUBksW3
IAV4LDbL+SsH2gNDNiYpeZudsjj9Y+GzsAWENa6ZBjM9vfQ1dRo8yPBYyyKu
wxR1UJjGRMuB6wKLXFQAKyvjaw2dLfguhbvuKl17DUNIQyc1aQ879v7W0+LX
zawCxm7fCFQdQkB1nWqPzkyyn8VxHdBmbkWoS9qxk11ZHDsQ9efyxPzI5wpc
7kid8e5mkZHcjfhHXEIGE4oAN9P4v49mgd70CDGUKsAnC5LAR1w/Pbf7wtbC
IUVlVmrAs0Jsc3quoLqFyuCsut+beaZSjfzsHFEaEx/yb3nC4xGKtIP0MN8B
UYSpjGek+4ifXe9ehGtBB+phf3QdFw0ftSrDLBAWuFjfHSi3NPZoTwJhY/SO
ygzCkmnQJN8Xz3mjqwI1nQ4ihjiaxn7+9pVxsYHtEe3G7gLzUqG4Ogmwmxv0
fhJw8zma91XDVeNsfySgTZ4ZvWJbmd6cpyOwRc6NNjn8JqLYA6tuL4JjU1t7
5oSClHdKhU0+40Q7i0GRhLtgPMeOBCrgWeIu2W0v++RVR6bHaXXESp0BKk0O
CyVLq1ymDHg1aBDth8T6T9tq6EWuXmtcI6pAdDYPSoACnP0hk3XqK02VhfHC
f/EQApdZlyxHD64+WbKhwn7oR9253s/4fqbnthKc9Gmji/IlizvNYDzlor3t
8/7Udww6slm6gmqbmEJ/jO58cTyaHZxzUrkFn8kobrPiJZqw3K3z9xqwsF7W
L7SJi6TMcOhHohh5IAeJLOY6HPliXYfX2SLOQycWA7I7dSJ926eQ52wT7QVl
aP75lwHgd6uDLP/pkeURaKJiuTwku32lXiV3CYDTaJbStzgSCKf49P4Hlz+h
pTirV4EaPOQYhsy93QQ+u7ZmJc7++1Ur0D5AIpMh8Gm6VAd2bR/NpkCuRUO5
P4qJto8almRUAzf21GoEi4mnjJUYJuV7vUQ0zYQGsnIBEefFCXQocYkEXWXe
QgfYSb8fwlA/bDMOZ+i/+ZVvmkjCegw3Uo9eqVD8HXN2RLyL+ScXl+LkSjNS
hivGdoQBg48K8b94j9d0c4fSLCuOeC/iXaFQYw7HRLY/VBnj7zKlOj5z3KDP
RrgE9AEbsbuwk6UvkJlNtSyH+qTcOYlYYop89VqCPOEzhcVCKPiyeUWdcHQr
R92kaWglsDiIXRH812XleYim8dt5D0Yr5YGeomDbTdoqvBTQB6kGf5vBkTUu
Cl34qWhgCFoWNulpdVVBQICAMr+MgPQuXvYxwC/Zq4+B63h98CxNgCZSUs2W
XhpWuE0v2Ju+LjY74x4mAokNr7JoE4k7Zztry04EEEoPQQdQRrc3MpxBR78p
7DNEsJv82gSUyEmSqmF56pG4vnlPQc/o+Mkj9sWe13a252YG/Dxf6CbY5NyM
8ZclhpjfH2MKGXb4W2NyB5+4MaervShpNUA0yyq8awsjHf7madA4f1U4brN2
/lvZuezIWZHvUPSRfBzphxju11tHh6aLHapYLW3CwjbbJzOcb6MMXw6G7uDE
ThQ3OLYD3OhCOZxh4JzLaNoMH+mjY5p7/bYvZ8e+TemQ8cXVHHTzAFymkkVY
vVPrBhD4FnmYgKzpn6FzyAxhCEEQgOkXrfvJEsyECgWgpkN/Q41T/KI91O1U
XwiNOG4TuAlOVUERc6zXv7ls7OOqv6P6pqysRJhTukSqNm02ko4Xex5+Md0A
OFdgmXNRFXtUrGHxlQCzaj79JU3ij7LHWBzAmVRcQcXJCqYZsyFP7XI2bQeu
AvCiGaJnYpmW2y9xIolewjL2z0V/W1JclpQzxi4eLQFTUUgWrDmXvjElGjnQ
FlK6gmUUwJlx3d9SsKlUKrCMSJNh14pm7Dqz74QEvSdTvixaDPNmBN428OOd
cR3xt928WFVuVKehgChrZvjUqxP7DVD6adIT80+FCBsvwxxc66MsuGnOgbAw
AV5pOo07O40eipw1PoIL4d1kFtV52sCpJyxMAbgclE5IHvM2kj6dQH222zE4
kLqIlGMILUd3kP8j1P8GvlOWjvK6Vj+TNOutt5vXOQzsTaTdHe05gDZwggqw
PohkgKq3Czihv7TX64zofxZX72MkfCSf1knZTnRNcj7JZ3VnSLWkl4Deg59S
gBelm7MfD7ozapzQ/7Pcp5dVKu4hq/YmS/dUebzyjnaM8AEIRakzJ0QfG/Ju
CwmHirWvI3psF0bvKQrXbBDcagWFOCoKL4hXrryt/6qfc40VGc9E3HPRQ/pT
WJvqLVUDmfy/X/ozZAojsCWCJ7twa3otRKHQGCESS5NWOgS54cLr8p46sY94
fZtFF7820q7Hc98f0e9xexlq5+2e5TfkMUndFRbS8OyYURksoasm7NWBPPHb
5OQzxSzWu2+wMp3kN/WZ+sAsz1XdnbIPvStV9NPfF319qOWYCAmoWgBDzjgQ
KAeF8KOrX/VYK3QCY4m8rLnH3PcboQnUyxOOJiztQ5rGiRqp3u1jZXRLB9PD
2ZvRQjFopWTXaBfWgGpD8sPpgGKo6a4EQzN+BRKP85pO78PbI+X53iJzYVT8
JL+23q2+zK5jaq3Bow0a3zQ8eFh+McQ455tRjMG+u8OPK3FIrct32BWWUoZF
Ut9xfYRMZxRx54gz8Dw8qF361eDkNeGEvz0vNfIKykK57oefODQvglvJxbjZ
iguQ2zZdffO7HtPe1VSJ5p4FpeuxdYoXSbZHqh8kPGQb9kWVtpD1Y3W9Vjk0
QB6QaQZ1gnJeQrGUxvy2lewJNf8fSCvZovFROoiB3ImVpyPo7jv1OYKz9HJh
aUX2iw2ChpVHNGPPmX3MRaUtnlc9IaoaEnFzt7XwrwGGUOTFrvLWE1JxcGHR
CqTELbeelq2lrepxMvF9g0ZmtBqTtBNuye94/an/xG91GtEQRt/f9hWEJFVj
IpwiQrv7X2yphSuzVTMYQodLUPHAnyGeMw+Ecxs0Qpfrdb3C6Hnk+sc5GBir
L/a7x0VHtppK+9moXrYYKbRaBlAfVFP06mHgSBrEx7dBW9dIBshjnpN6cSSN
K9ADYrCpZtkYOMxc0ETPRLewDyvkwrk1DAeVsSUo3dibHctaXCBFir/MgZ33
LUuorTgeElULud5EYK/SOt7la3vk9eEVB3BtfNNQIi+dHB0ApNm+YEui8ihS
KRDHG8gClRyx/sZwHP2NZtgQ9ngKlA6ydky1nmuYYOjfQVw68a4uXrFhtXEN
EvpnMNiQ/z5JDhU6XMsSmZ7qRbPELUKXYEtOtonugLO3ECJiOmRRZpJBGQ4N
oeecKNfRtctn+AGo8hfUFHVrFI94LUHJr8ozmCjsljhggAq3kinMVNL6LdD3
LEwCdNyyroTFYbgHDPjh4Kajn6kqH77wfz0nt4u5SMHTr+J0WOs0JfKayA7g
oERyVyH3a+KLUk3kWqZUrZCHEufdo+HEHAtWzV4mN+mGP2os+ypzOoratBWK
ylbTWAozHzcPFMQHg445TO2YvVy+bwW9IvvughsHih9I7G76esp66BPzDZxZ
eUH0ytjUNI9VVH0Z4v7pfgXeqZFiP3kJbEVE+9/HcdnuHTbz1kokVyZK5dCd
a9kdOofVHZlzDkDe94+aRsNLCEzmBvrCVBhQB0AdFTrS/Wwfi2BNvN3oXrPu
dCv6nswZfgBaewQCuc91VCg/Gl1AWVwNKvqOFLxIouc+pfsmX92Z8mKcPreI
XCdf5emF5FI+jfPCUXagNhE9XlH1nAW3XWZUQAlGv5Ut5yQhTsIj6mb/CZ7l
WFcjHyhXcn8XrRxC0472OgQKamQ5HJhL5v7qJAwXP2adpvhA67l0D5t0a7ih
lAoJlr26hGl9wjITUtT6vOGuQJvEnNjTpujCgESqWsyCNaGXjGvMYRpOOlyw
2Rtoz4iparpDWcLsY0XfOK7JD1Jnwg3scOWKuyec74BUJJLq79RonSMY8/jn
mcDTiTw0zeOC7gggbsbW5Wb4CLht/icMQUzd1fNaHehZYLebr9KCGAQsnf4M
FBfvjPqSifNKNM4+Zrm0uYU/+wo42jMgelb6eufIbX8Xn7V27WfCo4aEmPu1
9N3VD9U6fMq7dtkA86IoJ5lYQk2p+kTIJs4O5k2Ykp+nZLHw1cO7zAwOLrs9
rYyLqVQuhy1B8FCwWzWzFabdW19oaJgQPRamwLE+Tf4TYnA8gTiSlOnTLGX2
DYGlSlT/FEr9JeViWL5odX+N20uLxAMHsLX1vtCGSkQ7a8m07R2BgovdM3In
Jn0ttAebWixX/NRrjnpL72z2L0egx9vnoNCkQo93gG8DhpIy3uo6FNnOPSKb
qmrpguBYfNcQuKis1BYd2eazpWpwoAQttnqHU3DNey81WVDw0v/QNd1KnNO+
ZRrJjv9xNJO4hxw5t9JbNMGAO6JP8Fd0awGZX8b59zSJZWd8kWz5Wi0D3tEm
+2nj5Zr2pXzIGOGoOQL2hruhueuNetNl6pZLNGpEQ8MtC7h2/+zMmHx4lUI3
zQOD4L6JfOpUhm2YFpaZLxzlGfsW7yNpd+1vnydLsDkhQPhZPu52EeLJOeCk
Nc1LH5UaRI6P5CdCrlQ0MwCJ/k5IgF8vsW227g7Wruq/cIGd/XQvuu/2neDl
NQX5YLFR7uPvE0pq+GWdDZaIsS7urwBHzdotZUOmVOIKDZB9RpUWT/Gpj0IH
/ywhor4eCLqF7C6ZI+2awvaLVP2pc2VBw0vMTYCBEvHbcCe52pEsMgQzcqaj
myvJB6e4dLR6/S4P4zXfi0FPssZrXIZZ7s9Zj5zvbXpHNuTNcDqzeuSG9daN
q7mdB8XFHVBhFGFxb6Waaq28mY3qP3ELClNK4u7+gUZXEt34SuxNmBGeBROw
xrbr4yv6zZxfFtd1MuP1BzBsy0eOPnJCSM/zm4kvJaAxW+N0wPdViaN3fLf2
uBaEJL7TYN0Acq7hbf/NEUlQWcavcCtYn5uxgb4g5aGoOc0TjGeRNTz+/ZsX
3GXABKwVYyhqdd4Yb/Qs9pKiXSAap6kgHm5hcwQjn1izohe0AI+F8JlWrfqX
5vQ1Nz9q65DmVY6vzI4Uu/n8nt8Ij/vgcytm7yRZxLCCkrGdDoKSlgIluqfY
7szNFpA5mOzjzlumcURxpI4TLolE5hgdiyTESyrINFM1NA4OlhzmFU956PmI
qw9cnuAsZkNc8eRslfOidi78WgcNbcN0k/CrybL5goLo4gz7K+Acb9BmeGu9
qEV7NTPascMnLDCh7gjJ7aN7n3tfdr6DlGDl+jwEhPTsQEJYzV5I3g00j+HS
p4MrzJZUtzrU2Hyz8MceeQcQdlMXtVgfGQfUJ3RN54l2+A6fnXfHwsDXfSoY
gwyV6b2S95cg4gKteTgNCYw6hl0JnoY8RA4XjMSwEvrRau8ppN6krKX1kLR2
VFar/d4TeyFikoBOLYicvae3BRCKmlTA7n214ASiMKFHtmKdd/zyVgr82WBH
QFxGL14LRIPa+WxLVOfrhNhQfKYyrn1de54W9QDIrlVwTV4QPOWmuUP229/B
EnOdo5s7R8jI688ibuwES8TL9qHRL47Pt+xkQUdQRU7hrGvf3T1VF+ZJI8UZ
UHbOlwMyn54TlSPISKuviPhMr7nIV43GSs1V3P3e/028gcEvQs14QpAddTnt
Dzx41cjLU159CfEo36m5hM8YwBi7EWW0LieA/EQeOlmyoWYFwsvYmjXGtShi
9k2kr4aWzX4e6R55UoN92nT/cWcyhzRbX163t8fO7WymxCDBBE5YHj+wtGtz
niGneMlJvFK2LWui/wxsnHmlbocB3zoA0NTbhtw+gXSvMQpEiLey1Q+sDtME
1rM0rKaUJyZmZ3+Yr04Cp7A+T1fw3GIs+oUycC0lRlbcnJWD6QbKjS1vZ2pn
bXdJKnmiJSKtSn7tjskZPsm7rL0Al1GqlHgQaB+Imlnu4O5Ue/lJDdaizbX/
lPrZd5wz76VHLaMde0XYF10oeUrwP2Xax5Y4uR/AQjiFOYxDpmnBGMFjbbGP
f1DZjuagV4r2X3SHIx4RRt2M+K8/LIJTaSGhw2FJrSG04+Od+LWe3PlclTb4
imu+bXmSek8tkV68odZOVcoUwC5NrwtggMc0PAABW3NDE8on59V6Au6a6oeC
0yq/3WdB/h89P6Lu448iAcxbtfNyiL14SnpAK3bASzsj7KpbT2bHoHGQQhzD
ENT2nD8zSCyuxB50uI9hK0WLSxyHqPgQ3h+vqxif30N17X62HUFMv+BuQsuE
26fjwkfac9titBkE/O8h13AMkgu7sIQpd0+DsZD2jdlo+/jKyPY6MZOF64e2
jYZKX/eiw+s0G3VcATArRuWXtuzoO894SDG1ZotcX1GuaQKRlzdB9meZ7+PC
PNkfWbgEy+Uvpp92uzANUNO2hQi1ZsQaIR3YxcYozl2PoLRq12YKWIwkC65S
en9BiL/8UAzcVVQp2IZyhCEFzFEh+ALv5oeW0jfdtZydRTFh4x3e0lMnBTRe
36RvJDN7vHKA1zc8+UTYDeKxQ1g6ZYuPGgFXeJlymfhVKb+NyVRYOIbo4lyE
2fpr9+NLonFdErnLdOSe3tnciEhINFwBNYaUf5Ta+wOz8PrTPDgIWuk8igky
Z65wGpcW4Kg5GjXxetSxiSbjrLAZCTgqoncqc8A40J4QqQzVyeILnvpDq9KD
ZOUInwvISQgtMPKPuQUwGtdTenF3HR8FjXlQLGFA7H9xthPBGA0dH73QNcZG
2TogJZada8po1yvqvxS4wpKJDyZqJv7ozbzfHNqUafCT5xBWSC1367kSUqqu
gX+HsDP2yoGdHpeBEXNTxnUpn2JcbFBryvJyCm2gIwLu3sVuoQwpjVd2MREH
Im/awXfFXuKpNrkOxeClUfsmKwJ+iD3zcvVnJeEW2RfzIHrhweLZV4WUGvT8
2KX380hzCyuzOT4YB720/N+oOMvobr7hB7BoCzgzC7aXNSSLit8aTuiY+UHt
YmwW/YrK4Di8Rey863YynM7vrbCWy2eE8h/O5NtZBBOW5gwCAWMuIdu3OZrJ
r3q3hcohmpTjXUVgPxADkOk3O+0WqzwFLJmBqSl95NNEelpIjWp5TZkGA0+K
t66K97CjFFKM25n5zzRpBqUUglEA4ZTtDJCRFyGBTZ776PQYG6JnEDQARQqE
JrZ+k4P+VnHlZtEM794myM2BHL4N8N0Y3Zff7GPruRa/iR8uXF931sofcOmU
ls2qb0968eQ2lHOUZO6EJCmIM7lkFnBd2zgS9FIEU/9jT0tFLs3/k08E3vOO
hM49V2HvanvmTQuvaYBkenUkks4p8OhKAHeH97H16J2PDEMloRIVQ7RnprWP
s6+Ppt/KnUI53GZ6/pR2cp1Y4nlKadmEtdszVQAMIVH7zvL21Wpb37r8iWo5
K6s7UeT3iQ5eFYQWD9quF2Imr/l2x6vpdCVNCSfH70w14EAZ+F6DMJY2xdGC
taclGHOl3Fio81c7sk87gvWGvm5mj21lP7ZDkqGJe/SC9mec6BElB7yxWKLV
xDAlQGHwWE2yP4Qp5CJVFoD2wpamOJjEyc3O4eox6m2oCjn0w0X3R3f8L+SC
I/4+aZU6/hoYt8f8Yxr2ikDDIBeYDTxtIkQjDFV+4WjDcSqm2EfZHPTpbwGy
svaaAALYJ6Mrjd7dIYqkCjvyjgQmZpXwG+t0LZvvc2Dj1jpXe8q1ZSJlV14c
5AgRz1B6nD9WMWJ7RsOn/0cZvTMcKaqz7IC61tDIJjPCYNFSlYyg9SL5n6xt
qRvV9shv2mqPt6ZHv6KfZlXVKfluHZdaJUWgrsRgnZVc0JKgtCYbXTM5ZdoV
VXf4KMfGbcfXMsTDu6qvzfyLG/Y7LgWInrM72u44zODwAEYw8Du4qQ/6tN6X
FBR4x/xb7Xf6+OPr6siNk2MW7OdGXaw3Sqi4aoc5eERdE9wfjxxklWY7RIbi
kDfc1y39FJe7KEiNLwUxGpHbf6nbp/TVRRsp05UJDfE7E0YCt6rZMqblUxUf
ZmZue1NTPEJ1u0My/3fW2hrLfy/Ed4iH0WJ96BCg015YkeanYySNluuU0Nyl
BrXAXBwujehC5CzjgwQaeDVg8lSUIyMd9sa7yLojXaM12iPOh9BuGKg3kdea
h5iQ2eQhnYeeMmFO/52biPnh2R2HOecJHogqY6GKepA/ZoXqYxR3+L3YR6Yk
e1z+Scyvu1V0mUHpTS38cOaAkmmvrf+bv7fWRdKQ+s1oSKejsIgT1xWZ+uaX
2saFW7VxC98K4DbNrmC/ZHrQzJ+404h4SaCRW5ka9r/C0HuQJGrJrfPitQE2
ICq7yzTLnaU7Ee2oLChpkyM8xGmDQqxkY47QDsqu07t+WrmLaN+EHgBZ2dpT
KwXV1DM8/ztktTxEEXqCRMDTWhTW3dFq7MWd1fLA///In2I69Miohl9LSq5u
q/Mqh5te3j5mxrmQYtJ9+RLCDumshBr+mPJqx7AUe8xsge1uL5Nkr8bPD25r
cb0oDO3SBTy3IavxUS2OPvIibShzzB++dHVPL/vEY+bIiB0JKabMTj+uoBiW
WOcoTE39sHNVxOOgDz1yIrrMHqlLP/QQM4N1qZvcL6eoMcOXFehtVx/R35Wv
QZHAcPU5+nIQwuLk36ia3Lef6Df8F85F3dIYUGRZTkIhd5EGIm5idVEHtSe/
ZdT+bUob2VGYDwS7D422FnWTanthFnDhS5Vjyapk39UvBpwPGH+XjRJjt2VZ
ibLpLE5fQFJFhqTrMZK27EzZokPevRLctCA9ld366vOAXH9GCEWddfjjORPI
9YvHzEBouh+UGw05VdPIbM+MYLuShaTETQ/32wBLMdRkWpDTJuyS5dfhvT0K
1tYAj89gSzCHn79pQvjnyq+eOk14S6oWkLv2QEJ7isiYJV1S0XrXsnkU9Qjr
qOq3h/d8FDdZ61illIuPsz1gi5njO1d0wLYUtAxYgxsm0ajiR2A5YCR16vAB
e057XGbZsH5ahClrX/sS3oeia/bf65LpFe7/BUmdgdVoa9TUfO2y0HJj2a5j
T1N/OA5StOR9oXaycGhOuG1IQAXOHEaAQsoJIzlf7pI4i8/lrv/BdJvZa7dv
h05U11pNtYdB0F5GMndEv+0jzTlKu1eImiwW/fEX+gW4nkbjUcv32oKQ1+dS
EVCfeGipiVEUtIKQHRLKCmIV4eCIIhgMe4Fc+D6bZitpGgn2foy1GCoffOfc
KM25RLZO3Puo+P6FMyOEBzCDzELCbP7yQBmJg5Kdc2C10SkY3I7DfKOL2ePT
OtwziRVQbzOtglTJVBpkjr1moUleWgFwEkccZj2d+9HVHKW87l/zcpTmN8xy
jbNzWFVgSy5WaBtGoFJjal5iT7vP4bwWyg2z3LAmN5zqI0ivCVr83Lf5hDLF
YmPAHbEAldc8u7DA7bRrE/NSyoIVLloqzd88z6EHUVtwWFDaFtpZREDp3w/v
e+YGyBkJ/P8brJuMqD8NbrdLOp6YtiBVoOyJs3QTiW++IZ0xgGL8hiHPCTIQ
NiGNH53ZubdtCF1CkqdJw7MRgmvB/X5a/I3LoG0RMpEMJDjRLRpGYvlSCZPO
F1StHmXsT1eZ/8ChfNF7Ii1J/9VeZ16MSV4JsLeH2WebN4iRdSnUSiLIE2la
QyiWPzpiMtvbI7dzN1io6fzTVzbXYin81En3JbsbFQPWU4iGsLMaBHaiJCiS
CtNHEBizJsUD8HY8s3MMyiqbqUX1IDRpmtWBi+Ze2Pd8JtwZOmwD6RNJxTta
E5OkAyOhmPZDFamcLC5Ydj8vEst7Ql/6vcyKYg4IURaPjI4jQ88378dAHJsC
9QodGVsRbEyz10/T+8SGKyXueoAvKpQS9eRqvZBXCpnlJaKg8R8aX2iyh559
v0MU5l9Ol7L/d20VS+aJPlnsWi7kIioQOe9aFyRIIETeCAzOBcUPAQJDnSeH
EyRMLd/beY2yU424Io5kqS/rQeYfT8eRh43uLb/K55idsVJAAT3v1c6VUdp+
NVU/IFK0d9qVrFTsLHBbv6pCpAtbfb121ft++SHqYnyMiFW6kDQTiwT15Dsm
X9hbUwX3PO/GDth2t8ASA73QiywGgShsAYRcpA1GGfS+IUyQfuJ5JLJcrLUy
2uc0oAUGFxuWZSGDhR7EvBlegcZnZK7iup974mMmc4LJD3IOWIhVkvuldggW
yoyfNbYv2lJ6wdhL/ngUAuc1szUz4Q3Efa8fAmgb6SaTSW8C1sq4c1JobcNE
nCcIcbKwahVkNYqB+PkDUaNhUcE6jFmYeqtPtS6omlbf+I67gABLpRoPrRF6
aOA5gTx9Qj94Kl5WrFsejFGZHkDWklKVlCaweus21p46SPgZGxw4RpES0C5b
IxpnOYWtnLIHahqTvAalYyHRgzPuPH/HiFZwTBIHqfsP8omCzesAgIdprAFg
fHeD82/XDLvXhzBdZLXhcjLQtk8wVQIuVY3pc4JeNryI/9oO1gMAjsLzt5/z
55q4bjLFj21tISSKOncR1TpAdehm70KTJFcRiTFZQvLeBOaIzI+gCEXc3YS6
cw7pVrIItc0TYiSQ8+3VLgkkCZu4VWAeiZz/ZU/9LffaIgIvWS4WDp5cuJKE
TiaHWGuxSc9QxNNUOtiVTt3O2Nvo2pmLgtpU6y1t/lnEPaj+tCFHcvnve0Ud
YIxbMc/dzKFJ5TWPWenMF5ZlIzC5q+n1gNqFUY1Q/HDQC9lrrNW1pfaJT1F1
p9Q6zX4CVs3xMVYxcqRm4AtFP1zv1TA7YuGo7hao3p3GJMx26k+SPrREVCMz
oDkj2vOnDr2g2rCbDGySRB/YBTpPR0vxlvZLKg+nEa1p0Ep16Ob5/qOIKbX2
mSE3Jse/to3Ou7V2G7O5XZ0r5XjcndPRIbwLnhVhnnoyq/DtKeAFiNDmOExJ
6rD6sj/na+5s/Gw0oEWccePgKsxaTUYGigWpIIRbMde2hJdyrOBdNw0ZTy4U
LJLOtDBcQ0V5CY2LuyezGBzOAVLAhbcuJTYTtYx2Y7GGly3TA/robMBtB/UI
fqgdGs/gFFA3Ez+XgVquhcaIEJ09OdhxofBtzbqnirKNCCyk2bVvL3+7eLbj
FcK4MQarcu3FEkmGsO6FxMdcyK/Qz9uuhVAbIXgTFmhjPdlR2f+VGird//RW
lx39Pp4A+iMKiJhkMpvX+jSZynXx169gz7kXMKKvwsmTW42YYWcRgReRtR3q
XkE0+jlcNYwFwDJJJOIsnbGlNSRjyHU9eU+o/0mhR1E2HCS0y/o2HkHyt1/W
Cwl/YM1vmm8OLhhl/lAC4avo61zjdobe5HmgtCaNyTZOAJoWjaHEGF8Itoch
1plBC/CUyz9ogfSPmoXe9ln3gydO/6E8WPQIe52qSja0ad8sULwa55h9kIQe
4wM5BYqnJfnGjxA5jWQVWb9QFwrP7Dw88RRiMqq6mbvVVWJSsBZ3wgzua0X0
sE17BuEYgmFq2XtvOZkudVuHmHc0q5bS+0a4OOpC7aVpsPxhHZYHbmgaLqec
rnRHTTta0AqjP537F2CUCOC056lzAhVtiMeq8WUnO7sXj8UtXAY/2sHdC90J
3D2Awejb4jlXvVyTdQF2fkRulD46JpAa2DS1kAolUIeTAiSLFhmsQ/jWTPUX
dUQ1Md+IVLeq2GZY61RLW89diqhplHG6ddpJ3odmkEbqgEDlql472pIUMFaU
qqo5b5tV+hV0VDwbqtE/5kRbeHthBuMYDcchjeOTeGWxKsPfaE97rI7UbFHQ
k/R6rEJlDbCNyS5R0zY0YluZtnYvhArcF8RDTECKycxibY1Zs8deXLPTIHdh
n2HqLhdwzqf83jLK0O2TyaGmMfphFpB7+1bAuH8GxtkckKEONwnmQBVWU8Ju
QwyDqdJ0ukBvtV/TJCNO7NByhauTck2yNNuM0Alm7dum69cRrUlkbGpl58Z+
Z+hOQpziaMv+D8y7YRi89ucVrBTBvGZxyBXk8UaxupmFS+zVS11QBjt7JufH
DklT8n2JAsbBpme3BsLiRxbqkDYrTKV1cjfp2ccvNwYL1Tb9yJh5b6iytKas
Jc87bgQqC5FPbwTFgdyqkrSTirzJQQ5v98T9f4QLenHlmS5U2UnQoHVU2N1i
OofrSmExbA22tg2aeStPeCSSUb0U984o0Kgmv0HlRAVfw1Lk5gknmB+9Pj+K
a60G5ywKYTlZkCW2sJ4uN66sc7OyN/sfOGs9LJFABPcSFUrQu2fD7WMv+8Sx
6U40L9WEpfqCMmQv3z4lIxelrQ4tF1MotjjAGmGQHNWCT1/pDiNqca/GPnCD
I0QC03aE2THb+tJYbNa5Va7/ZKH6rXgmEfXQMBLAbrplMwQ0r44TfFBejekd
2bhO3aDr9qN2xCh5xb0Mln19XTqF/rp3ZCB+oxtzuY2G5gcb6ueuvqo1lhsn
LMe/TXQ6AAt27DzIKm0V42epW0b2e1vf3/2pVePAvlX9BgU8chagiz8ShYFv
1RqAc+gQmt8XvlG4mdr5HguqdGxvUTKBUlRMDxhsSdKtiDiTcPAk8YtJXW90
tt1y+PHOk9yPjq8wutYOWLqG4vmjx1FZCkU1HmQ5LRCq08rWOUG/ct14N8Bb
lUzB6YbxB+5dcC6fZ9KY4k0vzgroZCuBhFT5xdB0JN9DwIhB/lPMsauLvWn1
zxJ+kERp1wARhsAvT2tPn3NMPoO0aZUvfmXhCKY8qDFvmNbapoNVZbYA8WkY
E1AuM430fwNcUG83eVPUs94wGKTL4+HOkZX1F+gxRLGMj6WFKCipBOJZ1YCn
x3+s2DLJFAQSXyBA9z/Vyce+i4ysjvvF8eFosZ38bHzOsDuwWj8uFMERugSF
LcwZkPtJoSNkDLHBIOjrwKC/XNwq4k1RDcqDJ9kNbcveeuGNd96DSNjDl1Oj
BzgEgu0jOoJSF0ty6Gyu47XX1QbN3FcXBgTraM8nYIq/iq7XblEe+tnwKcQh
9+7m7gCt7PmKTAwl3FQmkJoLeiDdC+Duh1ElCbghZcv1NBfjOOcaoCaqejiq
M5vCerI10rGNYPmTJkpk1M7/nR8hDv5nz4ucHLxWjCjMW1n2jbiwcLfu/XA8
uVvNh9oRV/923pBAH9a90RaJ9GoVapadANvzjvVIa+cLFgEZzH+PbMN6GNSq
Ciz6qcBQlf0ui6x6sDMwmqrWgVut9ABEQteBkfkszXOqLdxcNYotZgQRYWk/
04GTtF1PbwjQYC3EholQajWAQZ7oGiZv+JVZgfZeoII8WOIg4VYme4xmiys3
VKUmpKqLOwtppV34eRmk3g0wruvLxp446015ypKoJ3nnlAQVdVpTIWKHjHmi
Y1H7cswlcto2KETxqwT6sYYRSHHXeluSmXmzkuJyLtc9DiN7Xr1FV3omQ9GX
Dzsvqqh9xPsR5stwjaLndgCKp5orhRTihWMoLWX0wPyL/23o95ZoCoJ2cIrn
oIn3/CqfSBkjOVcpozWlYJfdEL9Hr0imN8dY88mnSXBccs7mJnhyMlOsXJWb
RFi546weP2o5wDBFAwybuMbGqAKAVqDhz1jAkBoMsPwLBkZinstIEhqixBEd
DHnsY0EZUkZPbDzdEJ79gfhHKJyJuquCR/tm4shDLc3XyUWtAP4/r2pA4/HT
M+UmbnGhmGL9do/tYqRnuE+D5jFkmkNsayiDtmiSbAil2VjnV6sCFkD9VwJ9
2AB7IOwrXHw882hvc5QEFDEbiAOvAK3ngjzYKmqPpRvpN1ETH5xn76CB7zIT
AfO/q1ZWjepB3QI9NLZ/I9+I9UicxDBTBj03CwruNBd39VMd0nr3HH/7t8B1
m/9QBVVGHZFSA5d6wvuq9C6BMQpMEio2cuHXZtFJZbnom3AqGHHdGYUXoDT0
m5bma6ggB2tfaoguMSCnk3CyxvA44gcqWChDhc5tc3WmYtpiTAAQmWoYselk
n5esx5Kn7HvnJahvMCJm2OW2v94YSBzIsGwDFKoJM46WuvqcWPT/pReiN6tg
LlXO49aCGvew6TSh4j+ExN5D3ituIN09Nd1uRdxPnz8Avh+Ewcracpe78JIn
PKcxmEG/OCoYyaOI11w9+eKiohykd4rJUaMc2HnyFnd3mGeC26AvQiwltAam
P28ILDYVQMt4tjqRSfngRrx6bAR05/m98+aMMZeGKRW3OgdfVUDjVJAkrGmv
o/7r7+iI0EVfzv6+74oTHBoK2TJ+HHj468UroxY2VRJIyZgNDadL+2iQwAG/
5sI9uZBk5UmwTPD9WCOUFAU0ilatuyTu/MWgyXk51PErIu/3sKCVS7AgKPL7
JVagD4YeKisB4SwLGnIJxGac+iMoBW3REZEN+dwAl0j1ifhENKGaNk6uDOvJ
qH5CNumLt8gacYGh5HcsguFbCG5Si25Hm9Vkjn7eb8ZMlC6c6ckjbPX4hj/i
Ee7yIRxroSaLgww1gEDiACIxhHafm2t4csRlVA1E6VNFPuSWs2+o4f7CfmFU
9z+/za/lNcR02zQ5Bgz6woEe8TESl0ssQmwpkI/wp79zC308tk2DzHV9rc46
mvhejRmz5JiSJh/PfJoCDZH5/zX/FPo7U0/JH9cgqSTQ1B8WiHUjSP+HS1/f
x4tacUe3HhaIGpFa8FvxnAXCBXvrnNX+1jgpqMzIwuppbDZ/cFEPHV+aoXCJ
RURnY4MC4Tfej3JYjnEJaKLLTqkdLvwNH0cjYhfgGVv9Nz8VWbvHJCVI8aPJ
c5p8qOJAOrrp57m2grQvqPW3FxftAbkjco/6lgLXkOtDgp1eMCTMnVMWKsJh
zU5lizKuf9UjpasmTFhvNJojS6PBWkchV4103n0RBUM1gtV0iFjAkdEXL0hI
mh09rRodB1gfCEJhGgT4Zh6ONVhm4HrgumCwrrfTWEXAfbLnoya71h13JReC
bK9r2a9DeqGC0LGf4c1iHE63JRKghTVpXLSR4YOEndbvaUXLMgqfIFFRWrzD
x2NSdDmQ7jGzexETKm9LrPc+jZDz6gaWGuT9YcaaxJoiby6iOLw28ePJ7Bjg
s1WB/+SvoYJGReCEaWD+zGKQO/Q2k5OKG9ELzlOia2qRacfCPMMmbUWCa+lb
2ZGe2q1k51nE/txVAH1pqfzX7BvVUOztLjyqYA81Dplv4PrrKdHBKPglaCVx
2f8mPKr5q31xZnfz17CVIYeEOjb8iiUtm3rYauJCEzkE3+NrLRIk2/WtsGTy
UVywybrKeYmgyZkuLEZaAjZvGFKU6jKJj51LlZxm9/1CPzpjhpXrJYGEbE9p
zu0RTltrv14AKo6d5zVpmTm/BRYZOInbnPnkKSIkCL7hJoQeuDnCFZPbEOGF
5gPn/tP0L+GggBkob5Y6CZQ+uTpo1SbWigXtI8fp8rWlGIlRlmg5Q0QYUvII
Kk5d0DJsl5yWh07zTtTg6NeQvUGTWgluvJi47IFLVCF2VIj6rOLOZooFvWmY
w7gdgbW2hz4ORtijPY5Jn9RokMD4/1z0tnqpWZQjKJl2NlB0Pq2CyopvTQel
tZdp9EGLbH0CoBreB8ce5+3lDCNKcb8nOiWDf9DICSsf05aZKxp+6JL4YzDL
lhd5sf9O32Q4SZPZvsgG9MmSKD5WvvrMKvUgSgQF02g+LD9Hvwm4rx14sSAK
dAe55PHOvcoxBaA0WAwvWHeVB2J9VNZoaj5uo6RsdhbcVuFjmcH5fzxqzjiR
h9KM6i0P7x+XYlDaRn8/Kadw6NFGAhs7nabfE0Pi8+az2dWXs6lOPQEqMmwj
HkCjbloALVmctvB4jOYvR7qAL+Net18zRgewsfhVFRzLZMwni9pR0l0KzrjO
HFDTzXtwcVfyCsRJqtb73X6k6VMf6xF+jgSxAK1AAsMKoCDJQDqsUT9ZW3bA
O8jumbrBw1Iak4xmCh4prJd2/C0t+DbioP9LxHx7y52EZOxOLHc1JgbBnrN8
3XVhxaBbH0onX1NeX1nl+v+OG2bJVNnz7VKMftsvt50izqAxXJDnyhCJn3ho
yizNwpQRhMlGO0UZ8vKaSY08EqsxEzKDrINzP6rJQoQsyy9YZMqWQyyCUrEq
I5dY/AbzttTW54gD/qKy80o6VdKOY7gbaCI2pqVZyPmx+3Gpie0ZOEDPVrdJ
ILlpnLjgMFdidiFUeDCVhk7CGrzQ5BLMsxeAAeTeDzCJkbsFy5kWtwZjJ++v
Zgs3jLne7i9+OQzN1L3bos/aJ39gMZPgeWFj1gtKAAz+GhLYQl5AIKvoyh29
6UXlJnDaZjixTeFRC9IKO0G8beV21Rfgp/OEBgj9lKSbvAnIhILKrxzx8qjB
juTqqFfcJYrDV3VqmzdkLvshCLzPBWgzsaRgt16u4NBJvAqfk6mMFkRENvvy
0a7G5em5oNkeN8/ggXekXr6+l/XhsIaZF+gUEymyOXa3+CXpZwXQ+K+vGw2Q
7PNOBSVagC41GdT6OZFci2fCc7tct9+HADvZuwAeiBx8j3mpLWFUdjU4l2Af
fd9smu32C6UhX3JCNMBSLl3txriA+zxwOm93QaYpCN43SHPU8wGcD3UY4qXc
QNHAe5Rlrph2rQMRe+Z2bX1VCRa6aSaHNWxxNkelCCBrZ8GzzKhah2YrPoLq
rbCEVLuHWy4FVK2PlVtpbu++QVnqR+/vtWyw0TwfDI4CQQRhvmUAZRmURltJ
yaekos2qlbdYe/WOuBjKROIGng5OBCDXPaP9f65/OU0xICk7OIVPbR614wsn
9PFX2CHpROflptXlzyjBe1595e+OaK8X1iWdfAdJfZSJdaolEe38caro5y5/
TBnN9Ci2RB/wCMYUsjMF7YYsOcajMOMiakWwt3kO2k/UIfzHj9XpTHbyzN8e
ol4AexUK6DdF2LAbGHpRo9Jp6SZ/tUfSl0mqNmaik+ZLtyLXmMTh3netBW04
hyG2AQt2VHLiJZOS/Mrvq+h7kKIzG80sZdS2+BQ6LQfq0R83DCyLBtJgQv2G
tk3/BMyBHZFf7BfYZfoey24S7ES8u2crh9GhUWzylV5/YndwAczLqX+RapEt
3uUYlvvEpyqTOvziDAdJzXo5B9J9UDkCsZuNjROn+ELu6IqZFtFykr5tEBT+
DkXfbB+M5LDnR0FYGTB5UthSTetqgg9EZCeB/q/5v3APHJuB0gw4utuiiOep
nKMPGwlZyVzZdNqUW1l+3wnhmjqx4VZ+qLVRlo/IHsTsL6SVgneEhPk+6y8O
RqY76yUim0ZEP+EqUB8LpIb4F8PT6djrSrbRPUWRG4kCKvK8PyhstHh0Wos8
mMwt7prE6sVVVM3OU+oEbxZpzhWINKVgDl2VVnSlcXABraILj+t7k8aK/M9H
pmZE6KsGl+8VBRuPdCphlaQc8a7j4QShg1w/wVAneOIIEqj7LI28UjpEd5ZT
XoVbBrYnBUOswveBFEmm4/JdtBiAudXhHExkQrT42CD0EFY0l7jKyoA7TufV
+ctQU4u9JFJHjzMn9gOdhVpKY/ZgybLJncWwfqpaawbEjJ3R7YaGVBbJ9XX4
pv7qeCXMQDlbTC2Rm8uSu4iw7OEqkh+CZPaTVKJMjP+0jHMKvkdhKYnjJv1i
yM6uOweMLq6D2AxfQT6AwtAA7PWY0Hp3QOxGMJarng6TnWyu31oZs8wRYdaw
WFjD2JLVsaCO92GojSvOs5/Asl9HaA1v8cHrxoRzvVZ8+wU8W9dFnos8ag/X
p/GmqWXuBGLPuiSkVCxQ9Q7vfgdBWX+Lhuo5mrcVrohEIqvO8/OyZ5+Rajtr
6q5acxPj/1pIlxDap4wGvq2ZlrH886JXBdaIBgaVQ+nQ5WKa5wzkTlVk9xAa
3KOdO6fPlEGfrlb4+C/kh5q3iFzd9AefbzdOntMGog7ZvqK0X1QUoUhSLS9G
F2l7i+ltepK2MMH9gFJFeTX3PhxmLP9zhk9yPNzJtT5itXGZIUZrFaKnOEiT
f68oWWN16lPRadTukqTaYJIVaMu4aJ1VeXfDMXQVunyKD+wg3k9oDy24OPeZ
Su4rPEvB1vtkRm12OYiMNQR6mTfxomNfroFNxVxJqokAwbxQQ02+4wqXcV4O
HyHWT8BtV6RTmMjEBOVYdI+jeJU8D4GynU+6D7HnGqnMMZAY2Sy2W9go3ZRM
HZHuNqhEGFXU6TTaEwlv9/WiBCrnQ/yGb1utin5AKXMaU25cHxsDMxfVXQDI
fs9vvtPwnXXiN88qqQO8uNVJkG7xxHmew0+XM/mx0vqAAQYMf+0vcdwkqMSw
LaqOEBQb9Hd2zCHOa7Z/xrS5f0mFxiUCUreTk+uIjj46u2UXvm3f5QBTYKqA
LAnOHQgegRNTFn8urx2gvlyRBCB3aatJMeD570JYyjmywlMex+LWq6encKhX
XltofV0E5UiLOE021q1+v6zzdPsOw6oF2OaccI6XiXTc6ely8/6b7xzqH5Dd
EqTj5qKK6DOv12TaAdRNVAQ5bfVh/bBsLKU7DdLDEaVOhP1fOmg+HKYXVBig
13cHw78a4EbX+eP6WRv/jfj6vvJCg5zvxQFLPyNxVNiPXAfnf6RQSkUsW5Pk
etaj0lDRBSy09f8jc7mr3WaNkTiv097w9NGpbh0XAJl9D/0a3/CoQYv5ZB93
1vURsfJGDhr7AsevLc7GAtJkbuA+JzqvRU1I3999AocvSdjpk6ZdA+m2oDwk
dNE+pMrKHi9DNVZcg3mZLdvOOAX9cN1nRDbaqTDUoD+tg944aGRjejZtQ3HC
uZln6O1VioEj1JR8ri/Bv3Dn0kRX0rMgWYTxag1TUIdEA0cbO+9MikvV04Vs
VVXlw1BEUwcdgkbWLO0nbr+clqgGgQF0aPw11oP8oFn9SuXJITDUhPWNi2S5
uEruRyQgqZKowYZYY6RbNwK9AcBLaYnZmp8F0Ey4Mh9CTOnGHK7ELsAtShiK
osa45eG8qJ+SdyHhffMbymmWMiGZVSIQbNqVgiKfUoU2yW+xswZMgI2O1Vl8
TmbimTaoLuQDfyHF9wizYuG5hPsCLM0F7Bn+h23T5ZWv7+5Dg6E84zB02rda
Q3YbQEZVTytimllUbKbfuUIaZINXGCKa5Xe8JlgElX3/UaYQ/vf2l3kjZ8yJ
EueLip3V+iZ28thhN4swFPXX8H0pxXUeWXjZy2BodgRJ4aYcZWcSQXvbEBCA
A2Cf4R6jcVhFc2rVl4yviXeuWvSo1HQIMUcgSn2oRDkZt3HQdJJMyjiP/8SD
yAFvZ0Cmv93KKO/vhAfBpzzLrzZOc0ByPJ5r14qqxn8GI6Ul0wv4XiH8ZIFi
sbWB4WqKnMVJKcYidkdd+m+6jhwfWZmsuOS0TaWUL1v+aPt2eLghvdcUe119
XQr/ZX0f6CJuZ2QLCcxK51Od7MOQRQ7aVsyQIXe7KHvIyHf0P27LmcvYunqN
gHL89gFvtLuofGj1LfRIWAVSZaiMRtQbIA9ug+FAy+ZblKqaI5XkhcCN8sAr
mpumJzWx9WTG41ctc1gAXPPD2hw6GNVfDBWE19JrbyAjSLKHo3WbRp2fZtLq
dcXyD9n+Ht5mbvBT5aNgTd2y3/t4yeFgQ103x5sdTKI2NuczNje1jVJEkGeI
uWczyCKU7ZBW0GKfsHOo6vfb8nMwAmhUaTFX9BbjOULe1Q5+2oDVShLZzZyV
R4IyYXRhNTVx0cDOovJFwKgWx1tFL0Vg/CAGPRQHtCgde4MwkPOBWAmd9Zew
3DpfZ9LE9czW1DEEiRijRzc5sgBZBZg8pGHESaE4azcpW/mpvmtLzyK6nbli
TPNulFAC27BPapQ+PYgr6BaPlobQ13bB9EK+hw3WxfB9nccXkhkb0+dnXZGj
+BfV49Vo8CUXvJdSvWdoOaEz+bPursfkBfU4huCsSeReBmjFXuj3mwTaqbYl
wbWKg6pjyXqcP1B9Z7pAW+od011z6vcgTnkVnJtE5c5cAarWGhsfgFMJryaS
Hqf3vQEuGqU1L9GwnvovUz00o3fiap37AIi0hHQUw5KX6W9iW5K8tyqAj3Oo
Mats5MOZEOPT/6jmWuDb1A3Ng4+wfASjv1Rk6dSp61r2mZ1VNLz6vwCGsPRG
hVDOy+b2qoK9SkGQ0e4VV/Iu5imJPbk9KJkaSt5dZ9WVyxI3O0g1gglwpLQn
x3LnQVRetVnPpnmjwf/JC4a1cwxtBDvIP2KU++ZeW9a3k5Qm0CnZjdhYOuw6
lswo0gSbCsBoZobtnc/a7kc3piNsgXi/Z+g1yWLCksaRsKmYJqOlAohmq0jq
I/R68Bm0SpEmekkExzisijbCJXsn5RgYG5rufNGr0viDGU9W1dTfVCSoK63o
bSCr/QJN34Wbei42X1it36fx+tXcXTqjIzs2jvokC+R03bQWd+jn3IXueZGY
CpWAxLaCuQ6AtwwBxMgcsYDBVepFUu0JTq6snB8PRQMKp0xewULKUaVPCr8f
ET+Jjvkx99g6qnXkyC0Z0+W8+1f5DrmJp0k+ykolcEwE7tpylL9xve/ahiwj
b7Y/t+4QfIWN/gMVP39bXY9lySFqFGkVIhexZuhSYQc99gZvRYmEBj+lVZ/x
BwEXAxjDXr22VOJK04e38J6Rce5dTx+OAtiktptErN0MY+iHC/S7X1AQituX
l4xDc7iNunx+X1PjTyGPBgjF9nvu9Q0/QzQLXaiFuP32ljT4Ktk8J1ubJTUh
9kUyqO/Hw1wnvbcYU+wMaC35jO81qWDvr5jAuHYPfBeTP7UnuNMnxTzO38Hh
c/m3qwwrwPd5fDGFgunAbfS43DUHTIE0vpvHvLM7o1ekzzWVoeB3XwCxSix8
AgL9XNJ++hASUwYR+2LlQ25NyiAL8xMadhxI55kvJqoeCtJNO+kwNkurq/QI
e/+N49KblsNZJh+EADfYg2lLyph0Z5RJgTrOVgbZrUF6U+RFhXAUMgNGw64J
IAi18xgXh2EQpaxu+56sZBWAMPwOpUC9VtPvLjTlQ4ftwwptZiJMpEeV8OBN
aEl5dub0R2K1K37dJqHILATf61Ym97ZIaQJQcHzcf1b48EN2+NM8lexHkqO/
41KAmZ7ZSdL5prjZcQec2u0DbQBh+xkWkGHZ4xqN9+KzNkwcVe5ZvWWKnjRx
IvX+yS8JGX8QrddX80AUFCjMHLdPSwdcpTw1pYlu3JU0j97u2ULeSBdlbK3m
quDu8y/J56frVn1xMd2qZuo76ye5iLjZUzRoSlG0b6NKwWEn5Gi8rBOr+7xj
hjRpsEjvJVbTG3m1wnfv3LWCkdgGU5mgtGRJ3Tzyn1LsXMAO7aMlCt/O9Paa
7ME12Efc4I0BypTNwGxL9KNV6FvAS64ctEEZ/ocI/dIWDreVvjRbORJuIMGY
4S6+t6jTvvolgl405w0Zi4vaZtdxt9lSPjPTJYABb4K57LY2LAUyKm1VxTEL
eKB+sTHYNDfcK7c4rc7bhLihT2pf9oznPihGd302uXtIJTKhT2gmxVqJgnAf
nHGlqadruiCeDKtee14MCwGHhYsi/WkSp4ZNj48KCgN5iTD13NCY20DLvseX
DCWBWaayP6Nl7dJS6UKDmtAEHkcVFWm1DXtgq+j1QD9D1wymHIZS7k35U9Xy
uZmrBHQ7WsfFc9Ye1L5E1o6qCF8J0gA2csKILVHqrZ9/9UVAE6ctX43xXF4a
CHncaqfA/hV9MWZc7uRnyy/aD8G0ju7cWSI3AObBtR3BJasH3TVM1/LxPYgb
5iymPACnJ+KO50qKX3IHOcCVVQkAP88KMGQDio1odeM6P6zn8kdApkniIBlk
eDsYnqZx65rYjtodooO1riGfhyk76DfvMavbKJL4OiLqm8N3n+NrqPgBZtAp
NaMGi8HmV3cMADrkbAutZrLA2swMl5AhApYmLEYNw9g/6MWB/5hqphyGo6+5
WNW0HEpN9F/26PEwhqo/OUvAo2RUR9GXSEc+71yvy3gAg/nEijqTF1H3rA8o
a7EbyZKU9N3GKQLw3JEaTv4T5h3r2WarsFK8V+mRfD2iagiyhKxaNEkPvYg9
wQTRzjGiZbxzj1LENJlqts0KexobPzHxoEnby5UjoQN4cG4sbcYihSo/J4Zx
jSC+GDKnDWeKeqGejxiP2yu95rCBd29D/r+RUcKm0K2ha3VfCVn4TFOP0msI
BM2NEPTcbyRTUaHQia+kFVkTbGZgw0Oi2F5rtvlXpTUhpjiJ8yDFOsbbvxbb
2NmxwYadF3oDzMmlHacpmWza9hwhWTmCiv3pHlgg27gb8tbONbb29mJStO/4
Ga3bxaUQkiy88VDR/gFSo/uGzC4BKjd/VPRgwsDjWwVnznzu3IFc84I+C6yk
nVP64K3cIwnIMwISNP0+THK6VrCD8OpUD9zHxV30kUiHzZlGQL+YOZM8GyYV
qrarZHvHZcZ3I7HK7fNgHVfpJRcpKqVf38eLMQ5XDe6a3vJCngf18EUZbV+S
b3ASMUBeX6OKz20RF2miID2sNJ0wLxfFsfIRBKm85vQfo45LlB0tzPlxrePg
EJ8APVKem5lTGXR0w6yOOpdCaBC69kb4KHWQ1UslzmDu3Y6tqOp9xtn5EBny
6oeRod1U5E/E1TGoz3mkdb32Q6pT0G1JX0GHoTTQPC9K/d08MOMzIicixn8B
xr9NKM8vxNOUpQLHaDE8rviEwk0jUukSTcZJTfbiXe13sVOTrr9QKWxVEwzH
HdpnhsszFMZ/fwZ5IBZ3XBaOvFpWjRBeGtF0NUMKs9jTCI8XdxY5frsomrpP
BAMEOLvtk0+Y+qgTT/XZEhOMmJq8yuW6UWmV8cDZ2bkXGjnEI18XSuC1q7Yl
sqiUd45ndiy+iG18JaH7YQL1TeNUkZHyloCmEWDJQCtaO3g0eSa0r6kleUky
znothJ7ms8SLD5a7dwiWucdOySX0DGWMFeySRbPiRysfNYX8mIMibCzBIOw8
NbjNPdYBTNEoDC9ODeNndbEceFsERmsYd9qgdQho2VHWfadOIDWyB0mjzXqN
uVIQmrDd7PfNVtgQcFp72Pf5AN6WaQmE3sov47mJK4c/2n8uXFl8cv09Q8SC
ZNz8eI3F2g8Ei7QlPE5nsOVZaMzkNkLY8+zY6A/ehaSZUZUCbgscpp/iNNca
yVWauoeeaFVElFVgd2R0tEVoOTUpUmP3gmt3Bj5RW/COt47N9GSN0pxB9kaT
z2TXKmWdsq6ikvwKJdMHa9aNevF/nVStkr77qvI9NmhU8GbczQfZSq9LXcUV
UUfSGlMUFCSerpU/spNpJ9XyfZzxez5r8sYkOCbiA1q3j1XK6NQmNRVcoGza
2GVXEP+DYLe4f8WUB2IXiV90sco9uvDJFcD4X1Zomze72m0mslm0WsHo/fFT
JKRd6x1t/rylUEha2brUXwgShJgK+MFn6+lgyShDSRZadsGpL102DExrPdSN
YRQM/Mp6AsVENsKJWN0jHhrOdQIylxie0244eEbhxhoBrZJqiFMfuf70pD63
cV4HN2eIbRBaWgUuKDy3NgVfzaf61GEeBhCQKuQSt5MKUdgjbamXOQJsOddO
t6TSc33COJCkalMBXCRVMfjjjFL9cjhi1R5heKZWgCf6JdvvL9h0DHQX7NJc
6EVBXTvXgR/+Ez4CqTSfoRvGuJpq6iPItABnYLwUtDQInJIFazKrqhwLijgL
KTShyOqp7nqY58i1+fpLmQpS8Ml0qRW1F6gt/HZyzQhLhCV5RI7/cmSkxHlE
f6wibKa9nGWobYqj78hNdP2lombxNX7YbY+ksEVNn8XnBzrc8fgRhX5m6HrW
t1IQq9UHwK5iIyI/zZcDRb7V1E0Exv2TyJqJlrZ5aNsGhHCRC9B+zabgmQB7
/TtHg4aFi0i+qvKTiNOLwLPo/VmeEZlsnXRMd04WlzLIgl7Y+75vcslah37c
pCumIaSAQTV/0G+U8mUgD4to2yNM0ijhjT1CZKTSuEJpSn7v0cO0yzUf4cXW
qOMvbwaqXNVVPceaJ7v038sOEQLPv2CWB02iBECBpvX5SyH9fRqNPkGjs5ch
nSXgV8ToKfDdCrp2oc2JZvi/JcdjaD6M/6JSQU707pxa7Rs2186omQUaqCvM
fnlaxSwCMkb+dTZHrSm5bIqXmbSe4c80SKZgpplExeV4V3aPi2VjRhOnC34A
SJ/yzZNlv7zvLi5Zz156nJ3M3tZ5FBvewhvg9g5+bQ/ufjgqgjAKN2rCYjZm
Mvq+YVV6i857kMeUloXvDiAGgnEzlyYpRnt11FBuLGK+TVMOZ2JqN2+0hlkv
k0jmCPF6APye7Y9pWRzuUegz36eL/LDZLqttgVhJCswKYtq45c7R78T/O0Lq
ll1MoGXdCXcJtAdOUDY9DAo+o4Qu85aNSQzREuPPlfhccM25rykb502TY/I6
1jVWH4pI+7CSooUQhMFBHxB0hBdpqS48FFvAxbpkDLn+rfoQZDwNFOJxiAY9
CVwN5V55vrvbXLA2rzrjCJ+f+W+9+mqqV1j5cE5KCkJzwSpXkMkK9d/KK4bB
NOTtRIQmFC74LpfWrQkVxy0b4aBELSjsuM3UA+CljjH7ia1l8HiHfdnFJVZy
lcWP9le+KsVaRLtavrFW4LVj4IL19a7duvpAhp/2GQ8wM0QUwJE1IRffFZE3
oJv+lTl1V3frskTUSlHYIgSSTQJ2LOns3wSDcZsGSIms/4vtVF3P5VdVMtrR
sZOdJwg+3gzKKHcM/0g5Ibih7SX+H7hlxAngPs8Frh83sCwrrO5aKot353eV
MAJXEWgAfWI0BlhWbUvdQLrJFBT8zWlp80WdTtynGknTu876jpbPdx3Bs9Xp
V00jZwwfp4d4wWNyzJUgNR691vFR3DIycEFq0FZteG7j0COlHpZ4AtRqHhXx
FYb6CoL+MqheYA6BPGB/AhfPjokkaa3tHajmse8INAqx4mPQ/rygzmwQ+XJa
P4KfmJCeq8S0Zk0uABdmAwtng+SLXY4afdaxGHPOOp7xiC14IY4b77W1rlvE
OvssclvZtxXgY4/munfHSa3UhbpuFhVaTmmiajesZPrg82JbqJxsRT0MHWpJ
22jNwqqtG06k1NsKBRoxYmH6SfigbboUbeI2luA+9vOjJrDTLR/dJ8I2hfnw
jtRXLphLgmzEdbsjaXDo3FjHlJ8r+2uIYa85GdVnMdNJ/9MmrhQNBe8MvXI7
21X7v/kajaqwEE4c5QQ9JQOIxVVHPchvRG8DRfDOcNGEZEOsOi02oqy9yzkK
FUhT/sDzQDIrb2Da/yrQhSsQJhFb6WD0MDeLW5dojKjFhfrGNMOGdFMANf1W
wh7PokCAIeijvfEPgOMwO5bBf4YJ+sP8uBnj2hg/G+OyEfX5B1KGkVdR3eff
tBoM/q4UOGAYVyEK+0FEdEdpCa99JlMI/uwrE36oxfxQcvI0EoKK2E+z8nlm
6UxqvwxcjewTPVOxJDJfgDUNbm7pEvruBuMLhoB20AflZmwF9WrLRY/so/wN
wQKenW0k94084AR8crIWzWz8fpvZzt0HQdZDRxeJg/dLjIXRo6taygmMnbf0
GwWdlAbiLV4rQYpfhByzbRFp1LZUsqC7DeSNDf8AUCEL4569m1Pg9hlcPmEt
/jLHWYootaWKSoM0rzOG+UlSF38X8yjIKL2GYkS0HP82oiF29y0ewiK4aMjg
MiPtZZHNPS18DWpBRRJFVuiXzGdWeN7QMMdjOp4hgUESeG37rKAf84AVmCl+
HKtjCEJc+X4ugJq+3p1CczMIxUdhoPeoe5ppcierzkXgtTc6vOjEPt/H1GBl
nqpcNF1IAgWA5tWf4V0eMjBMdjfnnO8U6QTk8s38fE4pNRSSvIQ1PC8o8xUp
Kx1loI11TK2SCHwdt4w/nd+Pk5aTYq4nedZMxQUT5fMqz6Vpzl93bKvwpKg6
tavtBjenlDvKm3g23FvEceJCoiSZYf+pmPShIrVL7qKp54FNM8JR+5LT5LXU
etnbZRVOV2R+y3fqDdopuVJy1039hPQASvb4jQBSpbUnVVJBffEHAreasLhb
ZIxwcB/lebK30P72IRcsC7ytnIm01zG+fBchDk73x6HWLdfVHS9d0oDiMqeW
UxB+YsBHHpOQhnC5yueQLbpQ+oN5YQWTnaPbF1h85d8PqIOUYOJkhidieh+p
gd4N4+/NKx30zxHd9gdZK1m6zlXzVHw01ugJYMeyzrLm1OeoIuhiD8vgW1ED
yY405oN1lCQMmy1ZMdSPaWtD/H7UM4TaEPP+T543f0ZD3v7LIin8Eeh9bBeo
yVnCqXrMhoIBzfzC2RPl4oguB8gHqq7y+al56Sg+4GJFsAsbJBhu4k/qbAgF
phNF8e5QFjKcj3rG+NyCGOJoO073SoHegSlnmejPzkd6ENSpWUL8P8PznenV
xOK/6mT/leFSElk8r4fvpnkk0tyApkgumi3tBfGRw6TR1JMrzX6XP3Uphnq9
wyxHeAyyBhQqOOUbG+UkZ4G/GS0+ZYNO4FaKxLR4FTCYmVqdbW4jhSQIVvuK
x8KcIEqw4g0bD6oeQNQgbirZlCDXJn0Q36sX+x3Gzh4Uy8JktBdNWs69PPcI
ag4acae2+ld16Gn+l2fdDPI3yB23gd7hlVM5Ah0whFwSltOmqIvueZgpZCiv
innM2HBXVCuX6YMI6y0OKCW4EvscnExr7Ktb2MuWGZQTZ1UaENW6K3yjU2uw
fjsXhTq5CIdDvx7ivNhG7DKt0kXtrTh84saE1tOSuvKiY70OGJdtUJIrSd33
8Gj03nIF2V82/vZgRbtS5570wRYOgOWnnsV8T8lqjdXsuI/7fctuqNdp90YS
dymB2cMrWW3D3Rishu6stz2KRWhpJ9r+UqMDR3WwUVQHkuNITJFJNNrdemDW
R2mDQX0sjzBopqq6BJjU7Mt1oqw1wmQuH///Y9nNJ2ZHJ9vIOb3RSzUz/638
nHPZ2lNswcRCUx5urjnKX6f1g7LsaAtaz+5G52WJ5VfIRc9zZQaRDzP5smJ2
leyKd+zek/jHIwz0KLr3S/zfPyyDeItOmQnv61t4ZB3dlyeEEYvKZEl346xZ
0UR5DEC2ckaTGtGoWz5ZNvvJXFmL2Ioj2rNVJNSHsBc9VXnnllOSx1A78gCu
oX0UkEQftC/iQog2Cp15ZluTfPsrwc3+Ule+OYvl121K+nd/Wrw9eYQBRiIg
JkjJT0w3lI35IT7GOtbG01cm9HF36oL4HoFj3kUrOvrO+ZxGMburmsnBKNwG
XIGl6kcOGcl02DVDy7HH3euWCths06NMpNwP6H409Oxj407M1My1NIHxLNKm
Ld1jarzaJSu4496G6VzxBFiYf92A4nRRtjsroZjy/02e94mQ30flgdWZ8lSu
eXL1Eh9CQy+4I1uOP8UggEjS81AaHMZ6x6Yp6p2s3F0qT3Q35tDGwaes62sl
NYJUZjtXxaTGwDrdyE6+c/zQ/cD1ViJtFseAI+xwEZZDjG5j+F+ha12gitCE
4SXnpCRMzB9CSYuHfXn4K0eOd4bnRVuS/68yu6Hh0RO84nUamAAXT76Qp7wb
eS7w58FcT6RBT92XWarEwi42V0sDwxKA+A/1949H5jkwV1mj2tZAuN6QLIQw
wDh1NMxPQ+Vu8ldn1DbeIyhulhPXKmefyAcKBly7iZUEUdBJoxhlevvOLEyA
922hU61of4mXGVRATO5Ru3394ZWslW31W7GTOGdUhmHTr6h7VLIJRqvpMfuk
ShRqct3n+dq2PvbrRt6HYKrc7xuKP+qAefznbpiDEx4AKllZ7SkB+jM92Sqj
vz5f95oIW5hhQtaYGKW7WXzQ5aK/yFi2F4opuGhwYjYeInSgDl+vPZj8GpMy
X+mdbiljBr8R0p3qQ/tEdTDFWgPBw9cHMQVnTkGMrzd4BusDc23ej22VTLWu
vFJXoTIY3q9AYUJLm4xYMyAoW8HoNI0eE1NeG71QGpa8XxJ2XGkGh3DPP9xS
uPftExTJzeOjmrIgbFsZtjUqnigYOdtCLT4WP2bCUYrZHbBTTU2FMZOWkvUg
PgXOo2bw0G0fX/cTQ464sEuBLSMGWq4cY4HWOyWFGYincER4JbE7nFkzLIqb
78CY3ZNVMwR7+iEB8oqzBAsCn6Ey3EwrBjUCEHR1OoL+j5jUmYhX/kh7+204
+pgbfWqzvBxfX6+40sX+AMznZxRcan3beBqJomGR6OvkOvOKIM1ycgHLdKZJ
Gc16DY2w17q+rmWnZuUBBuLwp7hjkhQvjr5SCPYbXkarity9q73bLJUbN3E+
qtxMUGADo/7lfvFxeCmp8KIsh2CKmsl0oqP5rFr4Nrx1f/iUBN31mbhKpdq+
4SrklYDbhnKo71VUTuuwYyLiBqPR6x58KfhnTIIA7Uk6o24pu59spN/J8lQ+
rJWnPBcovY0bpY3D6Os1QJbMmITwG/XGys6Fw/IoRrNs+/6Em+qDNTIRJfDO
21VjpsGHMd4aA7FYsBojk8TAC+F4IHiB5/+qXe6UyX8Kgq7W3Ue5BKorGljd
B7qWFqE1ZnkySJoRtPxtYueqdF1PjONBTuRyRqJFJSiDz8o0ksf3HiDlpXIj
9ThDHy+uv/z/JbRFkXMZgjwoApana7w/y2tu3IryNSNP8NXQMZB8/16ye5T7
+HfTeyNw/a5LvuAuLZikSaGz17Uzz5GpGvt+o1ZdpFNUiEJWj/W01JAnfuUF
yx/tsUtzf1dwVGumFkZH3f/kYpWWH4AvdNAef33Aw7raqwhahMVJET2D2/Je
Vp6+H3NsyWwSjFZkfbiaDqUeiIDNxsOeaP+0tAoU9Ax3Xg85+ZRJ/K290BCQ
lJu0EZh8RSOCp6ekk7kmx6nse2W7fLXzu+f5pc/jBoW/i/BdnWlB+2Mh+iqw
vfEXq/32LjihQqnUOsE0oRlHvAmL2n7xYY6KGyoVemrEKUam8en0iMMeDJq5
EQ1SSfunsS6iJFmbjhgZtOrBE0PgJUkl1GiB+Z0inA/Sy1UiZtQpDin4XZS1
A8EoZUFjAau5Fo7j5x+tfWv4rKFqK3WKl1uu16QpIX08yewMD1F4ecYC/+aG
+LmjowGCfXW3CwpWyK7jXbM1egMkozOyufSMM2eV+HhTHBW/GPEyd+8ChHz+
D1GpCAGxWwmI7sbMm1vRZd8BYdUqNSPKahgbaqkSQEueYG3VVcIK5+a0b1h/
LNQV3dNQPQ48luKr8nEQpadbQqbHdHPI+c72h6JVYiUTLWpML7j+R9cnrBws
Ht6J2vz7RyYDMuVZ/tgGvd7+VDUY9kodfXWVnz+iH+12cMEMg4Fp4fmRseLW
i2eG2PsmLj6TMLkd7uiwOOur7yDEu9hYsfDRAhDrAPxV6F8STGjZvArWnNav
FdqhGgKG/Wtup1m1U0vr6ruVHuPE0a6NYan2OU5YqFzmSt94iyLcEh2zNeno
gHdwcJyH1NXXo+5SmFN16oKpqj6idfNdGbobEneQPKVdmOVF2SpPK/M2PdVN
CZTMQtMfn/5fdvHx5xt8uk9ZD8R/H3Iwck0tDtrrt952cqCPRXfxx9vKhbPU
rQocVN4bvaDa6rWJDPFcZBL0a+ID861oIyT0sPDArfNuEEjUC70co+qnAec8
0p8wNkenl/ZG4lawYmy3waL+MaQWbAI9a61VkjmPGwmlT5R4L3J/jDThe2vp
NoxeC1KG+Zvyjwhc58FcaX0Vv4zp3r9+m+lcqUm/nge5XQqpJBxOOQVKwhfg
B2xx/aF43EjJFiE1iRqrXyd4ifzaNDz3HDZkHyDwpe1bhVZGocvE3ice40f4
GvugPs+ELw15tN8NA4Y+M8Kf/K3D4uG/8E4QSYhZoX7gVGB9Px57ZTMm9a8w
FzoTybQJQts3vMAUDW0+NrHHTkXQ1uuZjd0b8giwVAUUKFPQDHv13sMzRuL1
k0xXCY/8gVRYaW5ZNqQTh4EdBaWvUqd1HUBTsoeNVC3SI9Q8F33VK1jRuYfu
xubqp+v9mY7uM+ULsBzGZbKcUhUkZlxr/zK06/BwxZEHBjnaSBQq4IyolODJ
wyTgZAvYq3ZbCXt3QrOtTcq0KJ31OjLw6ZqYZXaQsZxHDSHwuEdpYUO6zPZb
h3btLFn5xXm+tKzgRmvqpJ7ONFUAdVzreVXAqccexiJpH/6ZiRSvS7L/v850
YlGXtGrasbH00n2/wfIE0xqIr1x2UqZcCGbB9E6LOollG5zKgGsegFzff+2A
S3ME4oIlF7+qSsYg46qqz0hXA8HlmDvFpNkseZPovYVUljz6TOVYS54NcEhu
o931qn+QjK5p++tHbXqb5g2wZ4okP+OIM5HJeQpvuacK2Hh/XzT4k/frLyoa
e3jgU31E3plznnqs9FxKZRpCbfmGelYLENPZrFeKiNshCI+sadkfyvGPpACN
eJM6imlrUmY899YQqHrV2PDmgbKjMlo/3ll1ZFgk2sOND1kTADj7oFhGSrFj
0pO20ENBrUOXJJJTW3h1T09mAWVxae/WtRv8A5NIfgNP+S0FKb4GWGYM/ZDP
JXy1BuSDOTVLWQEjerFQoe4aCh8WnyW8uGChOShsYH/Z2OQCR4T+F4elilua
wRdUz/Wu6CHafOY4+4gf3lUghjqAFSkfd8229xc1B7mMrNkUzxE+9x94FH8+
yqhauv1Ho5XWPSOeeT9AR1TAhBIo37G+Xh3M7VjAGtWXgkcoNTiKK68OvhJc
/FTgcvWKaKqYjM7HnTUtbRhz4Kj7kwVn8jcg79VctfXrAhf9KgcNEpdyn/p2
pekHNQzscOFNzs9iIsbYlHAz5Z9mAOgwvn7c49w15XbNkIjImqa7ZYHIXtNF
/K4cH7Zt9hmQthHwP6xp2yKVKJ5MltyP/L6+hq6Nyw6ohuR6P6Sgh+M8AX+u
/rYZJ8MXNRHuzfwWyVjUuJ4CAx0gqp5bMBXOJBCU7NliMl1E2PtyenkQShqO
OnLMsxnvgq2gFTZlwctH7fWr067jSsLo6CqBENVtOL+b0tZKPlAay4qmFgH+
3JUy7xaAfefa2eyk7P7NX93FqT4GLfpj4sDsK7USxXJAn9jGLt/AcYiOhwl2
tibpNMwa9zNCnn7zYjI1jOtzLZaNDPIwXSRHFOCLiAvHzpyILWfQ1vC5jab/
5Jcom+WHJ3dR1nsNhHt/htFz0y5cmeciFMgxDfwrOZrZvUzr17L2wZm5h1aG
h7OcLzNarw2jLbR4jXpJXKOJV0t0ZcLuM/O/n9A0vcPnRXScu5Tmj8rYwRyi
8HqgUJ+C0a4jK7grgi/DRc4otqKsyz1apmPOoOwLPd70yn0nO9OqytAcajU7
iqw19cEwfHTd0Qk0XcD4SXPQAHRE40N/7nnmU/FcFK03ma1DckJc27YrF3Ha
owoK+jw4uZ3b/bfjR44mv6kukDdEpeb3agP8xV1P3w33mU2Ra90DU/BYjDQY
hyTjAB4rAc8h1oTdlkkoiYG9sKRdnMzcJc5LQmVzAbSyqkuQJ4PWGWRvRhCQ
/GMvMKZCqMyv7t0vg56n/YYLqJewdiy7P1zTUdk/jfokR+xWuvrr4C28DQt/
b+pfNmcHjZJKIVCVCrGnongtSFeBNCmNRGq0bIIC3vtAJbvoPRYtFuS7le77
QVWdXrPbncKgEQluIM2PWw+nHvDZ//MnmH1kubeBneGTJM4P+VqPossFgAXp
AJfrZ34da539PDEA/PBitBLD921LSjB9FLqFFDVOSYwhQETiEkmibd+PjLra
20TlJpm54XDWbCXapM13tjehQogqmyLrFFfTXyqzHirX7FdvtYbjaO5ZvynP
havSwhpfDTKoxkhTh3TD1wBeO2lPxhVmmcsoEVkQQ1m2IMIHOS66dkMqt8+T
wtRzRPXXxSK0lzD5PWcYozaGXOZhhwCj+JfGzfXKcj74am6WFqfmiwGMfks6
cx3Z7MNgss4DAOUTF3VTLliheK6zT3YCzKVBsl2gxOP7epCbZNb4FGFk1m4y
EYUwJxhk5pGWAygWfEMwlsU2cPk/62tLgHN/4VVryXRz3Hn8msSvrOHuHC5r
DxyyDJ0UjA41tikOCGgqXe3YGPukKare8sh2z3o//RcqmEKHUyegB0K9dBgN
wpNRZ4zQRgWqowXlRdJ1f3HUzlP1jbCY27mz+6pQ/+feKHGK9ByXwyCuq9HG
eVMGT64lQ7l1AupEE7KrbhNRX602whPPWKb6gD5PhzfCb2yjwUFKOsVpdjiz
9lLX5zNPXlLzmg2gJILjHq3AwofQ/Z3FWN4GokUqvCo1STQ1j74QLALaneBf
7eN6UZhzgTsJQUbcFneHREbMQ4GzfnvbILTULRdBDw4Kzn2XLjCuqaVnAmfP
Cqu7wRHAYNeGlb84xGcV1648GqgR1aePP04Hh0nK3XoH9SRn+0rjZHl+B/Y3
+H3wIsAd4m4SFcTyKQ3AX41vIIdemL9kxU/Balzk74LycGpaBvdfPHyzD9Dz
Fmtbxw9YmeC5QcTdH2uyVx9pNCOM2vC43hAcM6U6lMPDt93EfLuT9AqEQYvY
NVrxgXpbe8B2knUte2D7nmp1iy6+fxQ8M/ZvXn45vCX/60//42t5OB2aPT8l
tBfXW/LPYg0xN3isY2dJSt6KgkqCaULQz4ErpZba8RyHjHlOtj/jAuNcnMxL
RsN0RJ/RrGBkvcbBJQJVvaBJnddY7qZ9n+HBGYcVBCswaZaRYlxdXmq4MTUA
OMNSWnISmIZuZIls1FbWASujD8T7oTbraWI9VQzNIw3ggTAqRxleMOzWYv5m
F+TBjaXIXuCFawIetwGM0ve8FsyoWjnf9XP4fInqQKElbgwzaM+M9DlQlt8b
pady3ezHd2q5P+SO9+ZBsbAIkwyRNH7iIwGLV78w+0UR2dQUjnGEBbFHzAle
ZE4d0P0uqW0Yl0Ey8SuV+uBScmfks6Acfse6bn2XSRZ3mG+4nYGgxv2E+wwT
miXutopGScUKZ7CuP9zib0cBB6aGTe0AZYKD/7FrpSE/3UXf2t5PSFtSSowc
NMoI8dB9IcP0NVDQPcu4SLOWPXvszie25L5vulMh9/5Fh/K6kP5kFHYnUSF8
/ZFlAALrzhoDZFI1DGhya5Z9fu82iyaOnq6cBW25lY2lqvSK3vfx0JZnVHzb
MKWKqjZIduA/F2szHv9FnvLSK4FyGiFLBlMEkOmlBd7L7XIUSnccXVob/L+T
XeNGZPloBEFeBKC5vwiOOb51mCpm/6bSO6W7t5bLJJ2IX7g05fSLayQnmwBU
VKlXnwsZSjWpY4KLtNLLTAdRHgA3s+V6af3KDmOzLfw5gHUGg4hd23TVbHWr
Rl6Lhj6yDyHPXKQecWJ2TNtnqnh3XbZiV6DefcWG4/WkHm06vgjNcvF6cRwG
z3JaDLYsggA6DoSyNtcGcF8SaTJVaMPfEOCSO3CSfi6nQ/opPl9Oky7hDYei
vcyXPM9lK6O3caINLfCRC+mIuhl7Y3g+i2uMr2VsfPQHfsCMjP1/ibLgamsT
0FWjOF1Qm0mNxBSTmzkZccGHpqQzegPzjL6CH6auRNLNWYTWjzDf2CQn00GL
WK/gWHFRrOOosu02OUPifU74Fd6x1yejZR7ZxpdodU4JZrdcAE/W00J0rjKL
+2PPnEKaD52qy+37HX1cf/Em8ULfDqZ9PZqaDeyEPczyWryepCuzI0ukDfCw
QcO43aUNY1z0635FJU8Tdn6Wa8MD76VES3BZDMYhYWkU25QXid5S1tgFQ9Ii
QcMkoa6UbUVC5W68lqB4/MZm6ntJcGYJ0At9es3A4fDMNKU3FpQjw+UelhHj
xsmdyduqtSu3RaJzSsxQatrMTc+wU9TiplA7ivCa3JSkaQtOkw9QTzstJ6EU
Ve2EX4V2OslgQQBv2L8qVt2HtW3BkdZhzG3qECyKNwQ6HSB93CNbpJSykeus
9rhGbeUOjLOBpXravUmZPdF4aFb7RKI1JoDvzgnDwfLYmgYPGoXDEq9lk2Fz
EdLYElHHah6s4OwQUbz4RcW3/flngduaHdR4YYArhux1J95zu+ANnWT1qDMN
QPN//DyiQmZk+kRux4JWjznKLwoluWRUCopYpMffIgm7EnVBLBqMFF6a56lR
xmPMDJQtD4gFpv2r4t8zhU0bKeY2MB46/nFHhH3jIF6kvOi/c6d8NMySm4QV
+j0oKgc6+g6V9zw6JXVFL/k+AZD/4Pw7l6OhGt98xmSgZu1AGGz4XUEpe1fN
XSFLKO5adTeTYyEwAURXKqI144de63dqb0oTLDQRdX94vaLx80dOY4Aq5fhW
moeoJxuP/sZkFMcPHkf2hGlatGrS5hJ+MQcMTNtj0g034f3zvgR8Bubjy3Sx
L4hjPMoDajMz5vm47yN8b+qgCnUUUxJRXrRclYRTfxtgbsZdB0AxSxzCc5oQ
L1lgAIYm30+Ig22KGX4o391KIuKue0f5EcEAph1q6gBGf2139JgdvTcjvrDS
1nKd0Nj10bPtZXXBZiCJ6JUzE+sOayTBMHnblvhrLoYFcv55oi+oAuON2jx3
VfqcS2SoN2pvVafRDNwsZ3GUbgj37UjCujI4qsdt8DIsFl1+v5Du74bCPkOS
Zdpvk4i4fFWSlhcCAoiuSc8t2pXb73bS2hSOaaYg5ld7QS2oJE/EEZ+7B1+w
IOqNjHjVuyCr9Z4H/fLCfxg/PCVnSLQQ1RfEYJJAP/gU8H7X33Quuaivv0yn
cnz1EG4L+cGcej+bkLX13E/2S5VF/UZ63btn1Hfb4DVAPqb8Y3/vF4cAS1k0
Z2bM9NuPuFFRUhb8aalbdkLM9a/TmPOZIsUbK6ws6FKE0mrgKGzVISQhJa1m
1ydz0NsJJ3QNZBRV7oNRFiQQW1U+sXRO5Of3qlidtoNTS0HfGLEkst+PKDz2
Kqctwe/vQsLGDktkQuCiFQrwnqSQYMHfLda8xt7ll24iMrf2TaPHHSjmGbk5
Rb4uoOseZl1gNTlICDdKMP1mFLZvsh6cO9gGgFs49/gpHCAtISECApKXdc8K
TCLdVR4ycbZp8drE3nV8E1GeSWmJ45GkT6ehL7HXQYbFCJxUheOcy4LOnn49
8TOSXngtkQWo9Bs4/915+8bi4tzxKkXrRIvGyIRsGS4UUeBsXhWxQ2ENDk9T
lmXTyRs+x9HAuXot2cWgIn/wKjwDdyW5iLXOE0FtMKI08bhLPLaMBusCN+PQ
avXDUcAvMhlrvGehcaSnzpWJrC8MBeK8g5MQPee6K3armPa079LTSQyko2fZ
mprVsR785A5Xmj+WsfGxsim5xRH/uSbcgyphbdjw6iihHGYs2vKWaSBcHXJg
xRbFAzkPLOQat7/j22VC3PLymp5JC7uJFt0Vm+TyXRq4WIOlFQIM2ktxW7W7
QlCPxpkJM6lsuzOwfKR3BhFhDsZZrlOIc2zBc2PM9d8G0pIV13wafi72auqx
TsRjb7tRAR7JUGhrDCVIGE3VLeR4OLtIjtQBGiW5w5XC//dBk3qWKO0huP/s
qi+Mj1mpz8LDgZgJTCwEjcnlXB4+lRt04VnWAAKMhzJjCf52MjsGoZ219u4J
vB3plQTc/5cIV8+HR7Yx3T0h/QP/4ZGklPVOos5ls9zIWYqRu5951ffXvI/2
qy9hZXid7XEO5yThkZNqDtVr9ghMEvXKH2HNlcy/fEblx6al/WQTrNR7J+nA
NTgvqCa6ZzO1Nv+vhUUNPmNm1/zfqUufvu4/jPe/x5gGr/eDTW3gYyM6otef
nskG4kU+55rE7hN3lJxLNQweF97FC0hyadw+VIxJgY65qZ23ouDaJRtZf6Pm
C2mQkd/5OL/LGw4KwHbo/8jDr28299b22Xvkr7YzpRyIWBy2leVVi4LTFf8V
v1SHhBYtHUW+jlanXJ8QZfDXyxUeVCb0Ur9J3K1n5+c66D1B2k5P2qqnv70Q
3rdt5XhqzzJD86oCXV8WIBKxuUQir38UT/pLnvdNb/jk5l3ACt4M5EwQNklP
0Rtbfec6OgSRXQpozgDvt+JB2P6g1C5VwRWkE5W8fHgK56aPmJfU+8snpkEo
GyJ/wb7iLmdj8fhQNecLkNuvHY1XCjoLTP85Kt48H5feytD58+lGT1yYuuX4
hLDrYtujYrYbVuzoTOuEOR/gNsJo0d2tXoSo35spelDakenEVFsd69fSSSLn
nz9LmdZlbX8rWFT/RwI+9aGo85fyhxsslw4pdLlv04dpS9HuCtPbUdFz4O/0
K+dAVDeESa3MVqvxJw8tGaI7cAaVdXPdOU4M2Bkelbzx6Sajd6p+rLiZOkVm
V4P5IMZ7hTnKEUyN3R4g3WWhPbL/HTA340mUwJjxIQ3olLsa9ZwYzF96kB9b
2ijToqHxjmMAEImKHMJoVJqHkUipZ9IgJMjxQBvkzfVflqM1bIcEVE9uPX18
P9+E56yndP2MtpuhM/YmgYGfaL16si6BDS0Q+YCgN31H/YTzO3Zm0uAZcEw9
VhAQfqTvb7Juky5U1XvKzkGHfozJcRcSFDZ+bILpbA60nq1faicGINPMR7we
WDrqF+FFYc5WYF/asTJg1Lx1HOoPEao8Ke7TzeL0bzyJBl/+HKbzvS0tjqrm
pSq3ppH7bdaPn8e2A4BXSp/cqCzkGMMh9033Y4cxgOe4kYjMnEHLJJ5RfaM3
6hivPPRVm5Fdfz5jCJ0PitTzHTWEY+B6QSGgoGF5OTGS8kzKZEX87h33PD0X
URSR6y7zq5xmbW5juPPJrZj1fhChaoOc5oGMfAJggDPh6n4MjA+cq0V+Q9Uz
WwWuM4FUNAB9wPuxI0+XDn2QfqeiANdW5dXZi5/Ha25JPRvFjs/axP5VsM8k
7Uvq5JtPLbUm4k6RYZOVIgTUkEQaKjBVbuI01Z6KkxI2WcvvsaUe/57w65Ib
/FiJ9cD9K6oJbOFVnwJCh26Wfxp94lVMzC1ohX0xAD4TFuW6TlSbj+A6dPU7
Izqz69KhOFSbmGKk31pHf0aMcA8wcI3fxlsA5PqlyxeaNl5TwTGpc8A68A+3
3ZQfW+Qe0Khtgg6ly2ypORbwmbH1S1sTLKVMXbDDRsJGlR9XgbOX3CE5q7X2
1yNpFTl5MJeVnmxLAahcjbz1eBR+pMOzpXUdodPMbdUnjJFUlNB+0QixaxS7
X8mnoA8LwMlz2BjG16sYercFwAp2vhXP+2S4KLdtEJnO/BDI1c469p6zcjO9
2Oxvb4HBWeKztNTiw8If24f5sTtoCqGaWentdY1wfOnUAwMgBfVxmjoBxJyX
+6OgntStNEqygMeV9eyIYglgYcoKaupG9sZsUcsAotUsPSNYGX818HBsunzJ
d5x+5/WtPaFvqeKpJrXcEEamYgpHAPQWxyFE/Lgcs5e/1vxtgQtf1AseEKDK
pczFTm7FJT3fcb/hSQqepWszbe011nVTehp/9TqFH8dS242X8Qo9SGzD3BGi
sFZW7t2oynxGVkVrFuXuGlDtrlBEYVu3+CyArvrBxHQLsCIJ+jTnA0E5qK10
nJHMesxC8LJPhJOSHMsNM29iKXPc9Ivd9mIZzngjR4fDQ6CrVhwVxiCfQVcm
XULG7PnUz7Nwy5VHMn5jXAJ9m20UVtDO9ebB3nEeDE/McBOwn/QzoIAiSfYL
oV3c8alr5xLk3wuOoP3sWoUeQLP8K5kHle0cBN2SsTKOaLWsEplQOQ5YJqbW
+A9RBD+DH0aVBWj5tkLTub8wuWhdkwo5xlXZU6VK43xXY0+ajMnbVDcfO/oB
Xb6MeNmmMayXjGg23gI1108reZRNWtAEWTQEbGgix4Ep85b2WvciYn+DBpHS
ZJ/mOIGaRc0bApIOf2baXGyDe9K+s/1xMP27WO/ozKlbTjNhsmEEsW5siVHn
AR58NLuwpNsQbOBlQgxo21cMk89N1AfFVaG8iKLj7ax32My2fWvE3N1znfVE
gY1zd7fnu25R+BgT97wKj1J/3LJrqHqVb/NYMvJdld/jgLEtg0cM+8Ox0gnV
pwaN4uwK58lS+fF7EMit6ZAzg2BIXHrZbjzHwotMscr1j8c1UbMjFIRR+EWo
z5UVY/i13e8Ap3aShz+4eRu1EfgwPbQECQRMoOlSL2vEZafsP4Rw41GRL0Gl
oQEqEKubdylDF/xm0K1K9zU5PRaAlTeLrObUH8n/wYn6KmPlqOJEGSWF24DX
63IyOVIkscs0scKJ0Ell7DJ3hj0xU8P736pJ+xPljylM7ntZ7g7CX9m3P6yU
087yHGWRY4XkkkkBEgCsBxnvtWolvYDO99xRrjXzCOCqF5+ZrlnolTAIoQ8N
Bq+bLThtuxjRH+FO3FKPuIkDu5PMQPMyClkhmU9jCFBhjKDSUxTD2guf2Sis
5DxiAjXuh6viwDzLgWbiM2bEY7ashoV8PXAS1dly5BfyCg3DLWHBQItMdcLV
HoPQe+WPFFhPpu587HSfapb28OP1ysiPGtFAfuYbS40Ygb4lPaoyclaBpF43
e/66HwLZagnq12W207dZtRKNf8/NNPSX77edj3iX9zWNVT3YfYF9cZg2EU4L
Dk+kjl6wsQNgEPiP3hUTJhOz/o43OCIpM7c+zDaCYKsnLr+FkwtwCsXiQqgs
RHasADGRH6QOdaOdas3tPeBvIT6CiRlIxd07kxegb4M9gzh2BbpV04ay+Agt
K6gEAjRgARL7xEYs0d/U3nMucjztRtn2b6PpqDr5stEMvyJlh1ye4i6JtfKg
mYO17539EM5BwWfTQBQTn/A1nRw86nEoWP+UzQEDrXqZbmYgdd/4n1hMmK6G
iR2P2iykjdyl9201J45Y9cELaHd1J7JjuNslYdQtVB0ChoT2VKtMbB23TYpB
M4Y9KFM9LaUNGkeQtHgPf22TChsO5LYDobhU6Zn4Xp/YYXQo/nOXLn7TCTlL
Kc5/lBBoExKSA1tF+4smj6TXS4jelG0BT9g7VGS9EQYOGzeLRIoEwOYPAv6f
zPt1KiXeHjUUHyfRJg6f5k6wBC0Q42nOY/fWqy5DC0OBsXP9ScnI4NJcMhO/
UBkwoPAHyj17h/G6igycPgj5x/Ep1mfknW2EKhBcY9JPsvSIkMBm5GQHoyZm
B3fMsimRhYG113xqkGqtXJU/JuhhodNBrnlaDgvuKG8c52IkOxCfJCVEEK0L
s9fU7w9zH7dprmCZ5OP4YldKr7tYNRN+lPj8f5vYdxy32t1TOXNs2H73l8dt
azitZTVEcRhh2vKtE6+kDRK6kGrLDLpznCZTxg6xxU/m+dcD4d/BSzOqpfxR
dFkzfNhRtCeXoRNhPkleZs7Htn+pC4+SV3C2EreRjxcwV/elAxtYhKax4ERq
fhUmmaQC6m1xn0Mbi/HxznqW/lnxYhY6VfPuL8PYgcGtyEkHHTCqwDTBCo5x
QVEULS5Hda/S7Gd3g1X4L/JP1WE6vIezdWkJxVKkn/robeC1WPL3VY80NZXY
Z37kNFw5PUB6LDP/vUqpTOY1ThCPbtcIIXccN/x+G6SlmIAXWRFa8cM6EQsq
pXTtdtqDws5BkORMAGYQ7unxQp6M1sxC4bo2+6VgaQcbxdTLW4b1/7MkEUb1
SeTFqXWR3XyyatZk20TMr77gr+ooEGtEGIGNLlgnT+hLSKKIMGmf0ZtLhVMU
2yLyPbkk40Wi5lpzJJC1ImtEbibL5QFSs6VxNSraD46fIjSlGkdC3mFpvQFX
WGCiOFe3anQt7ZGDiCiegqC6x+gx1irzUF0yVKBeN+rlnslYSn8e/v5fUQht
nAYvIFVOtWJaShnxWKSmwItWhZdgUMRp+6iwrnb7846t+zGFdfsRkh6VuNdu
+NDiG1SXjL+KjVlZlO0LMnRihTud/8IOOv3FWuDkVzXOiaXxNRWWVvCZ2jmg
R1CZMwp3RdypM+36WCeal8YLz83NP2ABSQZcWClnphdFEw/hxEHAm/tMak2F
Z/Z4em1Cza4kZKG5ikQ4SLiAdqSzHHnndQ+p/M/FsRF3tAvZ77JeQQBq3AFr
PAbSqtNt3h/hcsOAZASRz9+ScEh/0EO9bEAvrUEc5z0zgaIITbY8oHDY9YKE
6aHpA1FWlTtbNfmNGX4fCPQo7kOguoYbvwDpj1xt1Bb1gXtobG73UxmLcMDE
KOL6IheNzeM8Uun9Ujdfg96Y2iQDrNkraY6m+/eX1W0eU+dNsa/Jlx/m/yOn
FffkULVitH4LYCbvOaHz4+dm8I0O+gXPP8mwMZhJJQi1YFRbUWLv9W213jkv
2mJH20IaHL92TJ4TwicWvAVd6CMHeQyypKFhbIRi4oFNfhXkTy2PCuLBA6Ne
nnlvUtpUugyfEw9R1nkcvjADx1BwyOhLGypf7PriyZ34TnidTaPospCsQI4J
NAsiej7n0K1SQTbgOOSMngX7UN2mxXBVxpPR+f2MhDtrzjzYVNlcTUVpYo7L
jBhFoo/wvXQktMixjq2Ib8S3ZbLazSntxWXfq/sQdvyDHd35Kwjcq6bhFvFy
3NNWvnh4LXSFo4+XwkhVj/Yw7s0cb9aCDXzKZBuOmnGZRBJUt2Llfbl5v73T
AfsGQe5QEoKX0TC33/i3dZylgpCFVdfhhSfSaD2nAY6zEkZGgHAJIz68FUFC
x7HoTYWlPucGpzN3bmdQQRkPdHdRPV6uA2DoJQyl1VsJqgV5wuis228kwHBp
UIO8g1vGkgFxBj9TUuCznr8ialbvN4ZGUxZF15ppHsRR8HdLHYf1uipQZ2Nb
Ed2+qcvJTPzW20tfoEoP3DjH8uYz2VuYxGw0+FRHiVaGAaaJflYyX2Ew81nD
Ike8M7dUwxodqIjc+PEwqj0bbUeYcZjRBpE6WY+33grCIdiQPIwPO6yPPVhc
svKRK2jkUVUt440RYdPJVOismk8ziWnZL6ZVlwco8hc4uIUUnMNrKFOBTebm
k48qQ7iH569u8h3FHLQKie0Mk6+LlHeEcCuAJUAfOL4u68V6rMh9Anl1ZofJ
8FVVg02fj5NI32gUzSKYM8IMguMmKFxEBHIud0fZ1hr/+cMwD6FpGKezNb8g
2FKlGnIQjh1o6Wa3JLpZhzT6jP42OBA9srVZLCkVo/2tZ5TQizXEeL1C/2X7
gypD48wBKprBBvnQKiba0HbkchfabS9w0DAppvL+F1pq77P6L54+8Sxpqgw+
4lx53IIsm0vyZ7H2hbegSfj7wIg2hBwWx9tDTyiQbuHZfvfOELDaTBstt0ee
DRmlBEvyuFtSA6/MjCnoEp8Wcff63IpGJ28F8t0XzRHaKx/pwr4eAXuM/MKP
OW6vMugN/Z/S1MIdBc8hPR5ztNjrWl1KwNKQxJ4WRhMztxkBFmbChgyzHCX7
Us/2zTtAValYsrzVftmSAZKeiCjC3CSuwuTwKSaRXmjawcwC1K8rgyS2b9Y8
fqNbYmIjzeEcwssQVCPuywlGeLil4u0be+l776zyjGud5ttQ6PfQbyAHuJTm
/dtlptv7EKoULvSNtN618GQHWsJhNetlRcCzSHj5IGRrUsnYRnXlr6XnY5TS
fVuMag7+9JEGIxiz/lOsgR6GlP0SZHISGYeUkl2XukZbavTgsXbRMcJGhTeh
iJjtAyC5SJgSvaWhy5Xhdrtd6ocOLGF0ek+ro9B4JGMJDFQO/vE910xLxK/C
957hhQpiEOnCAmsAGV1e0coscRqaIX9nHxrCYoDwGwYNkpDIRGQndgAO22xp
xGND83v5fWjDZdqwRmvCOqMBF2gVjk7Sve8xizVIQtXVPMXxqVKOYVmp+yy6
XCA9aF/q2J9I7BAvh0jqL8F8jN03ivGDpavGFVioF4tTxGQKflY4L9cabFoY
oNueGU0DY+ymmE7lUms32C5AbykSaAKXUg/KuK8keRuNPYVoA0254hJb6YrE
Qb28Z0fpHTXrJ19dMpY8Kb5HadVY4c82onhQAr+jPfm/vHAzFfuaAErqOhAC
e01MmjP5lvUI7lAMs2NPgEQgSk6NFXLZOcPfr0v55ty/YJGE12KiVk3I8lpP
Uz2hNMAq+OOZItmx24jFk+VxWmP3GX+X10UHv6jEItoUWtfsha+FN18ScpXy
yKDYO0kxJJwfzoRSq97uYlvydZSvn8RDRdn1g00Vznb/V7GECFW+Z0z1XzBp
1zQhq4MSxyyC5xokYwF0I3EDFmUSppXVkzJ0HAMThz3jAgqYnk6aINe3M3BZ
qrw0ipY+h3AYmd07hWeCTaiMasRXG8gNsqNivF9tg90J3ULUzyO94gCpYUIL
ugw/6hHogRt2oKCcrsWhQXJEB5y3DIZbTupyqxQbSm+5JoJjMe+jG199EgBf
oGvvIN11jVag34pgXfEclp2dvctX+39kwmFzGtgHUkipzWJt6Nx3O+b9gX3U
K5ivEfLpLQi+om/YYNQ4RmACx2rBkuiFV6ifdq8g/JyOSWDlHxxfkq7aUleO
hSzhJXXQHciINBqKFjYjE1i2uit5xYqIHojvDz7clrxqnuHnX7U6qUATM4QL
U8OY07W2sauUlCoex8DEGVx7nX9qIDRQmknOFjscuyvS5MfxOC9UpzDocuES
izFAyL3CrLsjbs5NmQc6kkJrQ6SNet0OScuTg9XAQyT1l8UGBn0hqSiSpdU7
7ziQfO+sHqMWMD0d0aaGj8+2/rnkSMXGxGbORznLbLVeGgHa3h7AtM53FhVm
rJmART1PWIEgH6FARE2RpJQYe4MqZXQFMI2LKEjcEvsMwzEWLNjea79kAkmg
YI1NQzb3y5kglMyhLhlXbJQO8M8aKauKCiv+qD9F8wxKVxwvV0FR4J6Nn9xQ
tSQz0TJXse7ue3D77BBjfkMHIFH4fegl7zFvCZYHg3QD4RyRxdxYXvDxMPw1
p7xth4axpQI1H+SKmif1kTC8jmC5GpVYci/+hCUUP5Qm7wlsULc24TJQ+8jd
6s/6GjkXfmuxYNrzy9BuoNbuIRNPK0bX3+dMML6OjUKe7Ys/TpDpgePLW292
TiW8CjbHCNJApj9XcOoe1IFFxkEdv3h9KGl9I/f8iy5fFc+J5cv8BgY/jolm
+iHDVLfEGRTdbLK1wRtnORLh17hjdc+8EwCSwsanJky4IZqfrCwySIQvBlq6
m7y2WiYR6Hr1C+dUYIRYYJyW7weXEDbdAJ3t0+c6KrK7XL4DVZCo+sNa/7Ra
kbn+SF26oDzj6cAbtZl8m3am4/Ya4bXkPbYctf6wgVRZtDKIGd9JNGq9H0tz
SBcfmWzeD7YoSpZ310YRhij+KtSTGtu41HCDWWailWaB7CpCrIvb4PRZwA/j
G4M5iFPzYejXFQoJ2Gb0YwgGNekaxlU2fC2vlMgJgCmkm21bi/9DWytsr3GY
AKl4cR86RJpuf95zkAyfHG8ifW674ce0DExfgebATiLIPjtqxzkGZAMu5F/x
4VNZoOyru1N9nVtrS/oaL9wKdESxSr03eCZC4evanN7/eohxquZnClZMU4nf
sAaWbiH9RYg4ADJ/wyFGF82py3V6wKlUOETBEfOcj4+SEg915emNmZfViYyn
ZHpIdWyLDAQ42NDNW6HiRFYz0Ats9JiGA1ujt9pvyTxtyLAe3BawSJbyeNZe
QTIXftjRTVM9Hf484OqgJg4ZZ7gzvIpKFPk0vi5/nkfXu6aQsQPP81GzqTKU
y/P/b+1R2wycpZPqiZrMxcYv1cXGYNYw/JZezJYIjgK7lCV7B/4Qm7fLzx29
aHIMA7VlhCCajuWonHTB3Drgi4xLllayN4AVyeuUEtBADPtRSYdSr6+GYovN
CPCxQCbgAsFZypezPstpCFdM6E1mWyO9RSM3NIKw2f5grNOvPHrxpNYqiPJt
6fj/MTd5ELSeZowYPNUtms3Opq9GT81yODrV7IzbGt1m6/pvUzZRwpNCIOmH
tjEjTfWECY/UlWWreTT2ppeJSW0Y+3xaXaBSGINFWpl3JNinlLIQCsu2inEX
7PCHxDwRqv81N5yAZSZJTsndCF4UHOciWvWWuFtiAu5+It6ZsGwfDcDKTyLT
ZkkEybyLzbYjmmHtUUtrXg6Jq1e3tGt1ffRhHLnZHTbJrEeDsiMIbdBQ87bE
T6K4+ONugEeQBfG0+zsVAIDPa4ymaUvprWkKvooeKMAb9OhzzudBQ68JSzex
TRnAQzGjnUHL/5iRLVxx+HypC3SrpbU1lAq+uNxhCRln1FU6+GQLT8+Qh9S4
4B914pxKcSSkHeBV+QkVyLG7OZBfTXEt3T16Xd/aeRlc7ondPuoClfBlRzrb
3ZvTdadlov4ExHzHFuGPAYom0+hXYvodSJU/vDe6lTZDeRBRXpTvZ4FUWNOi
CA9l9WijJfISRq9dbNIiGU848PwWvVxOBifi/GO0DQ20MKoFHPkG9Jr8Bwkc
WyaDSs36fIRKgiZWVOql8JZ6n4bbQoLnSb2nL4NHJ5pBvuLygNlyOaRjriWE
WrsTx+RtYfVXktADbRxP7oOPQ261L9VzEv7uT6UbxJOfMM1aTISX3U4bFlsu
XlOnA0LfQSNke22rr1nQYME/Bscr9zLVizA1pzg1q8qsq5k1lWel+M2SY/65
9dQNbmahVQi39yh1uvp0bU3OZMiGgt+j0NNOcy56Q8YJut5D2yS8v7qSCRyH
4tpx50ga16La1uPeTO2pmk5pyk+hBl9Ral71QFAjdPz1XYRMt4hTzTEpm2jB
azQSupWoCpv2z5YGfamoP5rVZewWf06HO6lRHpiF2VcvZGVS5Gmk4LFYdfUa
VmMKBaiRS7m1MZsQxoS9W0BpmvECOeHK3Ak7JBi7KM7NOcWX7PcWnehBeT4j
5iBoApk26ict+7N0cpg5zdrVNt1tYo+IdJzbpn/mqUUZefZvpDhUDqDShLmG
K2BSKVL2DxO0h1scZRqb+VMCT3SmilT9a3c0FlNkaM7BOCO8xQUII9qHD38s
2ZCnz8uqh07jNz8GAUCsqPBFHXpTFKjz/fbLiFADEILZn4FXANxOG1idRioq
XPCvWN2euUlztV9Qi8dOVNpABgg0zyPBecKc2MvfwlHjaJRX/6Xf1yrtogXN
IujtD3AMxsDI2Lioly1mGQy1xm4APqdh7q91jRqbFhS5y5tr5YP726tUkhTa
9j6kY4qzcRyuzbNwtUkxlVkF3BkcVbsRPlsHUICefV3z5slD4yczNdzdEkJs
6LHBOvgiBGdodj54a+alf4c2Z9CpEAVNNXkCnwfvDjqoVQgdWK5y35yfSwm5
XnTjuckwONvxyboGq+3ydRZQVwmysKeom1/JeO33SMTx3DbkAmt3XL+QiNgF
ePDpOxU+/f42jQUqD9Ud3iXdJUPx6iqZAYDbgsbVRQHD2u0fFADjMX24YwxX
wNFwqwPTeUhRnedgSHt/8IvnsdR5XYKsU5286oRjNCzRQKh93q0TvF4BscZ7
mqRU0AMcjUoToj0wq4zuQvKfmCC862BsmWvZYxHLcdY2So3ngiCGBiFF2lTM
mRzl5Clivjz7KX77h62AbMlx6cziu3ygW8ruA9rk5P2tUj6PXnz9UcEnvkhB
DCeFF5dqCdjQOxSsqlc+VgJleq4AbWBrnTIaZEy4IkcRLe5RdBrz+/2HG+lx
IzeGmOwUwGpPmBtPcwXzpJZiC2LzcMKhYqPt143dXNtzGmGBQfAqkBtXr8h2
dz52Q8vL27gdv2H7PlDOjhyjeCiXFVqlm+jxtxS29iWAjGDJoBvWNiY0y0Vi
4I4iPNdXtEfljJ+5ySl5JOvZPnPU7FWLi1Nmx7JeAyhhALyxEcvV2gfsWeP/
r6AbqngWrcTRuBONvt/9yiqKKqYeXm4vT+2MD5X3uaVLqPDXr2kf2kgQPQQI
5M40DP/sQ4SmhD98I10evktBs+KLJ5mprC6gMSXqGgrx0CnpTbogslYRAWWj
ZGWJsWGXang7tfKgpqypyPsd8CWxMV7aJYBbxz4fA2QckARDQ/QPtVlixgJ4
mNi+KCYZYYnZfOSwPfLe0Bd1LsbLwdza+CfAfmyMYkLdhuKdMQIEm7uszBwc
6bWRwsPFnOW8Iao9K9QZ8rtBYMWVnszCoRHY4PQ4jlIso+OPrH9bzwJtpDbf
kkMQcA/ddM9eQ58kGaIsPd9ACR2sWd8hIUMcv2THWag6fG9YFC8iqkA20MUf
BG2IDHjnQ+qts/H7gWj+1odZkyJspTRBR3O7HPeC9lushqG4Yj88VvlWIUVD
OeZvIhsaZsO80JxFdWPo+qLjbm92g7gs7XGFqXa4FYpqlQG4y5RIoCwKiCSo
ryr1hHtRFqfr03vkHeEbneGDOVqRwqRPjkuEMIdg6Ucvw64HyPfZTRRgKa2t
0ubqjiiS1wl39BCLHR1UYy47hzXpqt6E3MFn2BF8fy4BTMVUaNkSa06TV6Wx
49B6t+HcWVykKg2UytEOjg8ZVqBO3alt83VQoctUugEdCRhj2F6qUCSrLTFu
v58RKir7y452Ys8piGEx+VHMldSDFFHP7PUXRa3FFCVIXYKFswOJ8AoGlExe
p/AbrsqfQSt5v0bcJJUsUo06Oql6hYWasD9fZmOGH8jIJXowy0m8TEv3aSa+
roimYp0R3kQcucRGoBY00H9/goYfDFurL9XqeFY+hcNzbJbHnfGzpQd6IXbu
qR7d4gTeuF/2pStXhaE4XUqQ/z8W76rw+U9oNpF2kd3YsLfwZi5DAHh3OguQ
7fUuAm1FKzygwhkE1HN6832m5fYN6JuMJZa/JN27v/eB14kZtjQUNFb77fux
wh823+AJmulmr0E49axwiQ6fCRPAh6dUrkaGHMVj7UZmIT5Sx5XRVfMoLNXe
ky9O6mp5ilhEdpmIcd/zFaKaYyXHa16H/+fY3U4QVUlTb7jBof+MQXaMOf6K
OTfD0kDMXJwmxKoo0siS2txheBQKyEkIOlWNrZYszAk264xb/Bw3zX+SW1hs
5W9yA96SNJvdiSmkMjnYIR7sUDjeRjDxeUF6THNj6h97jAsabxFp1gakuEUB
e9GcRBvJp7/jcIeyHZGvnzAY3kjQbWaXEvFABbvSw/KNW0ZvYKpMPwxuoIpY
Xq3D1/PmI9UNOO27HxtX1yGmtCQm+qfNyp2gbBfjXTIbrs5vGIh/eSYNjD7A
FN26ZP4QC82wus0cj1zgqAQVqIe2jIbmlitFj9T64LMD08//OaqvCk1S+Uau
3tsvXUw/v8Db58Q6VFCYsOGWnuNTfSx0fSl9VawQQKzrzXNGCCNmy4Icf8qM
mZYNm0A2Vg1sjRHRUtbLyh8xyCmB0fpChE1hxasrsll/7TtoqDXUi8JJwpub
TltOsvQTjtI77kJhzDiBXl6Y9szoUqBP78jylWSZ2oAoWhXuQ7+fjPecqLyJ
cfEk9sDkDS4LoCdA470t1cn2+EdinYjugA0A91bXhx2UjlcxdUDkHADnCiiw
RRG9F8VajaIjvVN2oZY4/Qxsn8PA2OkIsJjH7r3muAXmNvo0u2RLDPGw9W8e
U33KAFB4bshv4JztA7Hy6jA4odbryscaDsA+I9V4ZPq9j52y1bWHhhWl2kte
mefZRL8ktcyr5zb7sVhXZR3BL77/2xUNkbARnMC1EGGrRdRdfO9FLdWIIwvj
gNi3GtX+8OXao8PBdJjt2nBIy9rOktVa21ZSZU+LiulRAlpfIZgwgntuOhHR
mVq2lxw6p4qIHClZPr90OK+/+hNbiadq3hYO5etq4qF9mlhpws+ZzIfyefI5
ouvrQxemoT6N+DizZAahOEoLtgJ5ghziYrIaEGpwGcv8R3VepJuP64CdHSE9
/UTBETG4ChwlWMIW1/taxZWotzKgeAdL8LgmsDlLRH2rGySBOyWS/iaYOZxh
ALHXEN8vlKfwErFG3/XbdKplhnKTaGfUjHhYLX/QQCiNonvUxxpE1w1VaFo+
5DgXZVxb/61CVdG+VUNq5sNq89GbVw9mov7a77DLN+mGNkcMh1rAUAbBg8dT
soqY4QQtTXdK074CZJAKgTlQKEZohxtvgF6H9RBCwVXb4MplE4lsb+OMASed
/JsQQ0oAFonfCEX5LvZren109FcKhzLgsoTqwF82OLEsNDJ/4SuxaAk7dI8v
YYUSm5bXJwMn1pCD3hPXOSvz9dE0Nz4fpEdQRb4kFzKEJXkXp8IerwFgk691
A5XbqOKVoZzXX2AzCPBxs+CKbUpeh4uy9uoxGFSmcasrDwo7ZJqd++qgQbhf
9gZnDT//PFJ45VfxghKlwOezmKcHt/AuPT2BSNjL7L1ps2i7gjxX3b5RUiOG
mYZEQJKtgpKGnrObNzNiF7lr+Jw3qG+rwD3b+/pbunA8mL2HxhRC8EfgUx49
NLj5jcoprw6EthckFtzlm/81WsrgustQenoIiY8MdpNfSuqyJ8CslqudCT+m
iRiixJtuylOLyrY9LR/T6s0UXDjvVmJDMoaczTN3H0rl1IS5tqh0G9o1qYMB
n8SU/0y2KnIDcy5Q2ZO48WmfsaMCJgIDjg1vQ1fXpFcqZDNfYWh+RO/mEPRC
vbw3K32LRlRwgxYBlHO6v2zj/araFP48DjvhgBWWieRm55YO3xGF4VIGp+Is
Y1RpaXVvjutOKXAzB1OfBEQvCY9ozztDetoamRfEH9QLoK4g3V7JvZ0I4h9T
zol3xgcG5KeaWUiExI6XEjBBpcCjK84bd5n4DYRNtaWADpTk1I/LaJFFKfGT
61ILpX72GgZXgKsDalWHxfCU6x3IhyXHROSb5GA5kXIIjm65Tki5cEQCEnmb
G25ZtXCxWLwNxJ3f8ZsMmytFjP6v1y4zZcTQa9MxzpwEgfbFb1DgKjJK2eAz
Fg9Mm5JcAE1WYmLnQG+L3MWhXDr8dDp4AeQsTLAIJjEh36bpUGLgHuyVB4gW
ocxzkaYzL539Zn68TNmKZ1KnC3kMm3g3aJVwbJWhjaPU/sHG/erW2b9Qy3Fs
czX1ge3xDhdGwF9O0pKQiqTLnbRzhziuB1DPNj4w0pxcR4oxNR8vV5hLi7wK
P/h6NYp0ja7NrEqaO7EDyQRZQEjmlKqvHgVEk3m9dcy1xeP/8roNKTmDBoFX
A0h4qmE5KLK2OEP4IBYtZG3TWUZQ4xrFtJvMyrKt5ragJw8JqkiJDxKoiRj3
F4849RYyyoAg+JdSXxQztwDwZ0Hbr6p1BXg5q8e79VnEqS8FrhChra/lgGnR
9iMTYDT0AWgHLu1BfDm9e4GnUGUW+BWax52GPLO+zZYr+gePdQjduFYa2U1l
+xg0aJlJAwMdMXwJRDuHeXZw9lniRaJzQS2RjHHpMaBNkboBGXHxRUpgansV
XPGwiSq+BHeRPaR4XzeFKNDpbzQl7dtBgVS6mTdh7rK1AIty+/EEDEsChtTo
1ORmt3lTdM1wJpDaeMJ6N3SBF+g4fqH0roJ1+wGYpPHKMlGnKd1NR4dWC3Lq
HNlcIwFxLPVAagOjuxVqX9bD8FyPrKIHMiJ+hjYfdps/KYml3jkoe6E57dMt
KKrcQRXEidlqG51lzKCVnLIzjRIid0j8pMSmyWOL89ipIa7yRgaGPeAIwzr3
k2pda4qhRRQ9xsZza1rayp4PC0yLFL/3TV87f/socY5a/+JihMJUDH1kh3Su
2hAKMfJP4cSA342+Cio89yFaGAdhkK56hFjafGfF+RJEL86hRy2Fk47fWaMQ
J3wjMI9n9hDR1MsQJNAj9MIMDThcKYfoYADYw5ghvepYxQX5ebYJWx/EzyxP
mKGqr6JZzqh+FD/dGtoSv2yFkNSYFmr1kFjb0KnnvJiNX5mys9O4YxdsWAuP
WN2lqGa+h1+UY39gfMRjgtJFw5vaowej9MnDEAB0pPoOgCWbbgyiVPhLlesh
NiKD38IhE4QCgGu3lAdyAJnyIjFk/zMOc5nmUmRlc/3ya9ZiD19p61a+BGPX
AhRCS5rJ1nqA/JUhv43K2j8ihD4oPVI13OfLgrgZZCP+4sZ5lJhDDwzLaA2G
xb5KJ1WrqdwwZVCGYOiylsbjkCKoVQM9DVj3B1A1p5COnHDDOabfuf6haCmS
1uvWZbXYsshp5ZEFNf4HsWJt6pt/JQLvGEJXthdG6/Bczig4bq7JzoksWArs
qeFy7pP+2bDh+R3iYzyN4HT+s3x9eTs8RCBY6I43ef8IkYMXdWwtNaS9wHzp
zN1jIG6J/NKqskXoaC2555VfPg79GmbAtEJr0WjLWM5RJO4fh29eCn81brCb
e5SA9Mz/VbimrK7Mh2mXawe6XFdBmooca3Yg4xDK01pw+BzE5/LPPc1Fww56
EwrYDr8yLTI6mPobb15tbmd4waL6cEyJ5sZhym4ckt8eOnssn/rmHgLdMh8B
g6Hk/kubGayyd/xgZrqpnHKKP2wkkP9A7Vae9XJfSyj9WVo2BKEQE/FRovSn
R022WlfEWezAcQVLWaDHH6kN4+ZiZZVq7COr4bxJ8jHdI5zPHYPIEdhPPw1a
6VIEKFjRWBuoamzrBmub22JaCZT9ShMwLChVLJ6PrYUqLNhw+qZmU0TxFCWM
11lNBQrka7ob9Cxk/sBALI6lKfRGCJ8nqJASMZ1aW0pCJ96NxG5YlqeQKuff
FDdKh5LsPb+tsFLPp2vckuzwJQVMprAr1sG5l9qiAcmLLSel5Xg+3Jxv1w6A
UomH3vKzUQVeOAKYN5/icvvLtiUwM8WOZfdjW1VqWOwtns5yk3aJwSjL/uor
YW5rs3ZT4I4vT3UNt6uWtJxnYqmKTRfwAj11Y0QtoNkyoqk6e+sDGBpK00e1
ik0+faKU6Q7OHSshB2dNZDcMHn+SWetTvEjSPnDlnjRQPoNzgGKCwSn1IzJn
juaoXsJz9PVjHhNfvUQdzxAsrVXd4Iy5LK7WRAQIx+0aO+cUDmSWNl3BewPU
/ICM9ynhzrH5iqP1VDxpD9c+Nq21DD9CKHOS6JTRF4i8CvAnfzThFGjcW3Gr
u9OSa07r0kmDmoAVhMBCWB3b6siPfVo2SeHDGw0lf9q5NsVMXSBvRaKndP0p
1BuxvZvOHOTQayAlBTWtfSDB4WeDR/jHNmpdjeumapswed/Cr8r9BcLAbcUX
eWw16rD6ffJFXQUoabJCJ+Xs6I3NAIsFeZpxu/w4ZTcEMiMLi+qAlhuJ8WqG
efE9+7KRz0nWAJGIai4F3KtXxpcr6svOnSSAyLLbfx53FcYc0zZQBPRFOu7/
A5pjksruktEFkJ922rLp3x2Ucc7gqRongQ0jrGUTZb6ApGAnTalZHfnrpYcY
M/tsOdQ20JFXZS762cSlittEUG8eijs0nXmKXRz/jtdNdlwbl18CAJ1BWXPB
+nKXRNBiejvrkaZz3YmoW9zlzZqw6ZvEIFlARv7udtxMQuTn7mMbvZ8qxkY7
gvQvRX4k9BNkPiT3PHBQm+k2tzFtBzzoboU2rWkxOMqGi0OG73qQVEoCIaXs
ODU+rwDhwp/srDKlDVWDpJ0LBJ/bJD/kt94KAYrEhUKliwaSoteJUrtogKz4
v+3uMpTM1zpWwwxkevZMN4sRz5vXnEJhKjtQYwj+85ywWWM4Z1rmaoh2pgz+
QZ9GGhDqHmdIQxqJTksqmSciW5A2SLSlYeTSNfZCkwxmKjZS8Bbvj/mkakHV
bdXvkVckIv0nx4QpjIiyocal03QQb3x4DMIW1+5eeifaPpTT+gHa/uDxPfXa
8rgTMu0VeU85HgtNLiSngbyXRP3eU7FnTWWLMN4usQ466nJIcijzAtY4U41f
E1fztBbbTl6eQO0ioDsGNU5Ku1LC212O0a0/xFJCZwXV5BzYu9WNYW5W9qXI
KUaDP9U5tiOQq1/CAcsORpycdHDp1xrMOZ7m7Bd6ds44j1u2ErakZXirm1h7
Qmrj+IxD6EdILZceSen+kEMa3Jnci43QEQWmeDratHHD/U0ZdfyQn8eqkxPi
WMbrqL9naaKBxLvBvTfsx+2uXFwz4r5RnX5BNMnCUaPSLudVPjHbgirbxbZv
HCXfXBNVnRBtmpECPMwxp+h4gUMDo7qVD7MVYC9blycf6nIf8M/VIzfHI5jG
eTtg3GXwSt4hlEVDLJzLL45ZnF8aqCWCmhYK3UMhQDA+31JwbCbohPzzgke+
ZvMGHIXV/oHzh7CbJF8elyhfT7lXI8dA31ipzB74lZMvmnwGMh9AbwnBJkA6
0JCWzYcNGcsEYsf2mqQ7x9lHIrf7vbLQFDsNo1zRBoaF3VWKu+LETuPg8DfF
ogcY3ef5L+u0uzzK7XGnFhlgdXA7LQ722bJv4oqJoaUTNoMUDjKlA4axGFEE
R65oabhWo0WRwM7iETWt60AJyZuV/sZB5RLV9mQA6tccoS8FQjtktN9Up2K+
a+pOKqrgGzHDb/XTNwRNQDT+3ClPIz/nX52Z+PQujdbLGojA3BM1WfNU7G5i
+2p9P5BJIV22g37un2qtQY3apJNKPpBeUI7AoxdE9BHCQJVKRX085TprpxTm
upk43ehfPcFEY1Nh6KLClVYL+K/Dw2S/DhdODG3M/yHSMANvdJg/TsSx11qH
DWAlPxeWmvJ6p1xUKFFjQ+p/+R/r5x2DinRbBZiYQBZjHgNM3bc+x6kYq2Px
6hIgqtS9/QLwZbQ/q9wTY5uStHmRpwF59wqiTXJ7oVKvf8KZJoxVACkh9pbH
7xgfDyuD9q6a79n0gwBhU4WQS68N9mjsmFhEPnnJ5dIOPyVS73/M43bFkQdz
1pxrSMN3ovBZsiFI

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "hmRb1hCms2kg5lxwgzvVC1ojkYPyZtVhUZroYIGDp3nv41l/XQfn8gMXcNw31HDDWBFvru7tQ/av+VlNCOY8CAEc3dS4tSN1iCLWoSLzjcf1An3u0nZDKunxPUWY57wMTkfTn6dFEXYBYGQG/cgNqAwhgy/sA9kmZ+yrzAG/xfCgRlDUR3RpN+hQPPycj5HNM2pIgRPAeD/5T2qj/frBFu5c2+SfDL19Hg79cXZFl7VCf9MHdzOHzpjPM9YtpdYj/zLxeVbvXwcnqpeZNphKQMWKrwtsK5WkN+7V2ynYT6njeNCrCLkK10J9+apkLojBJHNDur4/8ddItVZU+oFa9kXgkMGHi++6I5HG50LDVa+PfOZb7gbyUUnmkkjTqIk0OQUvk7bNJ6pOfvrQu8GcyMEoksuJqyra/iyaMj/VogllBn/RE5+yEj53lX6Zr+AKm/WAxQNFb0EtRe9QZIZZ6MUeq92D5BHHzUlOVcw7t57KWQyumU9caiz6p4/lwc2ImTsUpgxX0Uqds4UAL+MFyf5x2DFFdG+td0wpSqxDSUorNntT0d6VMgkDALkbc1FMBn2Cdzy1beRMsQ8E4cWXJc723g4P/sV0lYr3t7JorHN4ATP9E8vf5imdbXYrXmWK87+Je3l2xiAmpPsFoB8+HiohGsRlKmkjY2EugYTBDZ4fIuI6ACYExdPIHF8rOpwW2u25gHYkmPpmV53zsv42bQazvzm4yiWzDe2i+eqbaahzgXuvX/aJPs5j/ubTWvOoaDwYdG1vAokCltyuYn7T6/GPkNGYus6arYQJZI44sMnerP4z+Qz8ZyVQ9CknFbfVQcge+NXes2ZAS9rul0XTN/7G2auIfqBBOch/NPNcnywmx2f9q92Tpvhsu3f9/4O4GZ7DP83vYVSEazAOF391MtA8x/RgrRWJ77t5J06sMco9yY6QDpZ5pJhOgrCMX2q+purUEa7KmMPzLW/8zD2VBvtZS7fYeIweZ94fDwCb18ysvgv+tkZi1CZKfFUgrA+1"
`endif