// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OSTbNkjoOFNCJGP+xMFnGVf0wpkldVnDBdfID3BNLCUmeTJXe8EK3AwGavCq
1jNm2BTkAnGUAsIct4DvneRvSNmlubkArZXCt83bPvfiirNg2ij1grsuuFf+
pqHBvWFKbYdWzEz2yry/vJ4bfQahb4eBdz6sEwfs8IwNzXDMSFyhU50UzfoF
PI0VK3jX9F6ZofT8Tbw++TOWNIXKbWUalFSlPytiXS0kZNszFp/+Pfe/0JH8
LJo8t5pIrC0N6R3ukWYmj31f/bV3OoG/7aHNgekDqVrfquCmVkurWJSP8F7l
dTyF9AVs8ELpxm9tMne2D5YmSAGzWCLSZlf1sC92KA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iXjJTwObYMhVXVj0udA415xbOclJ/RyEz9/9PqswrryY1bqGRHwtNv93G3yQ
UaONhr1JfmZRVR2LGZrmaWXqO2jXEzEcqYd9CQY8tDR9KloeVkKqwWeV4y/B
7BIBGcirh4sI+X/689EU4s58VEwlyDSovd8IM+cHLeCazopab6CjNawKwz/G
TAKpptr8Vh/Ig6SWHjJatoovgilYTbJF7sBE3e1c2qgO34i5uK+74fB0YTEB
sFym11m7mnguXBOesXrGh0Dz7yvDsDE57laxSsuogoyaVueh7p4YrbpWwa5s
xt+EtE0g91MAj44rUy7KNQNOjhgvdo+YHzQm36C1HA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LODzkRVIvwsv1/Vpste/EvMBVFfz1aokAi3ivKhPS0ufZ6EGbefFPDHWRal6
w1AlJxKl54/eoFY02kHKDBUEaGth0aOH9sfTPoYuoRX6bymL4anPkiTpwdA0
4xelHHHAOYy/EiRWGeUipjsoLi0QOe7EteGcc4iGC8nWhPkZRJFOcs7MvLob
WumV8kKhe64HI3xK8ZqGzM9rmJcL1/D+vQiGWUvekCMrgBcdcwuDr0BiwusE
TdkIGHtv2BPWR+efc5bjeAZUrX0r8nYzsXRc6ATON6Q46aPYFb7nizf8Ayf9
A3KfGX9jK+Qy9+54yAIGa2EAowS394N9FGLwKBskLQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ejtFuxmzCWtGqgwZ2E8RVrCbguC2sICz29CRhK7Vmuib1UXP7Oogr3XLs/KZ
/sBy1Zp3JmAH3FF4Ta+OWX4InTDJjjDOBW8/CqcUnpiSTP8k1ODPs9x/hTpw
1EmnHl9k8gHGilg67SoX307Gjc8iMv2SeiCNZm0aEO/AYWkm6OJRsEuGXUPV
U5343Ew6PMGv5IUX5AxBF6c8vXxaTfQgk0JqCsuqv6VpW7WPNmi0QkZ+IT1s
HEPbBU25PBSL2FibSwf5xOJDLR6fh3D6r0A2GE7ypA4BEgSXBkSDGZrxOVvQ
iQc5uz33r8iL/0vQZvbPONxr5aJJBf2TX9mfUCV9Aw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Xk1vZA5/WZf9sBk4RcAI52u3Dk9zDHnYukgifJ781LM+0+bT2aNqNMwYo4Id
UFd2i6721N4Zcb3v9JlNoRi+xW3sx3DdxGGJ0YXayMeoP4ofBXGf0cs7sFJH
xua4kSFUc2jvfMLsQLUmp/F9WMw9PPQ2qM3sX9r5Vfz1jahLSTs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
dC1fV7KyJSmEbN4AOfR58dTLg+N+jyQWIvDkyXnpnZNas9wKHLeTLf+Oekgu
NNvCiHskCQDFr7JbMhMfinAx/oLr2WscQXnVpSQujcM5yzDL7IOc/HsaSHWw
uOtEOkZB+9LnruIpMyuAJuGHv9fMPVZkKhiEyD+0B+C+5Lw0qy0sQcd79hPk
Kn65tRun+T+A3uZ74OzgsRhso8WTMV7I3zkNTXmxpLHckpLpEuntkx7QPHO+
DCdq277YZI7Ynvxjdur5iykzqWSkhHa9s6dfRy9POWemzgRftLdesfI3Sh12
0uixAx5o2gh7wvp+SBKi8RS8/k4nbIx1kkERLaI2zGnRCour+gDRsWPdAvOK
Or6fRdTDBa3sKBxixnnYQJSkORIcZbrXMQCXIyjybUiVSshQj+zfZ0mi+3ht
SdFUwN8rqyD62C0neYWry97BtYeafel4ZswNVcgNoFo/H7FWblNJjsntVTCC
oidy8VM/MYIUtHkGO410Twalwd2Krb1f


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qb77cN2W0jMb2X6pnsx71cFcslt0R9EuLN40vVhiWl1P4MRQ7L4SOtvHb8CS
SHyzp/DyCwZDMJ3MnbGXBzSR+E+SE7Q8j1Qx2d4vOUU3lcNtEbrLzDHsVCLw
sZrUZlHSB3uyR9S+DCHGDFmyE2vDDoGTTguX5lF9PuaJIO/3f+0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bXeaOYKAA/tjRykGl1ewMz5arZa24Kpk1NdNQZQpOlDY8L4NuMI5RWKfqJ0f
C4KKCmFaVHQMVh5lUtd72/kFtcXf72+thHScQZU72rdNkvwRoZYuPH/hKJvc
jrTsifxRmvmMqZKObuMH1y7cJEQ8swGJwAqeunSClI49S32XpMs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 57344)
`pragma protect data_block
yOj4O6KlQ3TpklQB3do30JT8/Tj/yXZ134ast0IefsjAhchpBYmczbIeFnQ7
Ey/+HKJY37xM8vzuNX2cNkHWULTWy1CH96JqFRGUxjMCy3dloFK21uCobpi8
JokqZ47hONnU4vnkmdS9sdS0xHSxbXv3M4yhC+JYIrJ3iigXKzyu1tPgCNUI
jSHK2rFwQr2lzq6IH+IIMU22KXIGcGzZICEwac4pIwhlyF/CshS6qB2wjjva
MicdrmVtKOLANhkRYzLdB0WMaJDGff2xvPuR33s74fXpZM3GPmBho10i18NI
s9Mics/LuhdebAMASGsfgnJVB77KhDguBssYAIMlzp5yPEdUVo18f3IHhMcW
Hmvq0CcuCX7q1zbcDAbcdsiUWj9LukKAGdnO6sIoDxnrusBJBfds0SBKssZj
yzABUpuLXCz2Stx90TogrqexgOOd4w1f/gyL5H5PtJAmKSrcDsHI1RcgkKXN
y5ONWgGlo1bkK3KIQ7S586Ra1hruG5i15XeWFy5XqDdRC6TW5ZHMdpamtL01
oV39sUipn5XJ5e5ba0f5jowrfP9p9kChbZKpfv2jI48AgRZgVnBjwXmaYRAQ
fFRier664fJss2bIf06MwuTiSDPrg8qME4P5H0QaOSwoTawkkwl+7TU/fPb+
MLbCsEyrnhEXmEBQCGXTJZqX9iOhGfBJ8SPBkNMoo78oZXXulJqGzGRDkBun
I0JWjL4kfu/L0ffr5Ht59pN6+J2hk+kvxtfwRnJ3GkswhwZ1cX4vgT430Eeb
VRi6vMlwejK8OTWHXEbnXaY9KFh6GHFapovqbEJUGBT76OUgUKyLrmWRKWrf
xfy7GmY4pizUHaTRHnDgUTPSwQ+tiVSps+WOrFJE+rnXeur+RR4cxOMawJoq
QtWCWB42ytoXe+E+fdi8kjPbPS6gDB/WZceR/S/02227rwV1THsuNlNxqmi9
yUknzc0LUa8NwGYMTa5/W4mCiCFKfxhS+beJwZnIodObXk1bcOqB92qkb3Rq
Hq7OHFbhGiPOt0PbdrSvGYXLORl2AVzmrIGmfGdR4UEQkXuH5jmZkplsVxY5
llDdg8A0n0wX9ie9DdnHeiebuJ0/0dHURKfrxc3CuwMJe8WSEUEemU/R3K7D
BEiXA/C83DkkmihWeL+lD6C6jV1C9ntm02p35FUCqgHXSCnSkERPoO0UeQoJ
rmtHykOVtqidjAUyU0bF48tVe3SXVfa9cJolF7sXLSnF33jUUYRCwt7UeX8R
mDTz721MAYsyqF7QqdbKYT1jJ9SC3Y9dDT9EBI3qCQNpwHIINpgTManTL9t9
PjzsI+B9Q+hWZC5LONXA+6/auFOmxnSABeeBy/+I41H94lwcBpBB+Bj98e8N
mTRoNjvLlnUMIUwbufcytcHM4aMTBgTVTWxWtsr5VNqNQzFJuzUQweI+TgUK
KzSrDJ+gEDAvcx2F00MwRTj2LMEjClH6XTRnnMjzRbxWOR7zVtJrraoafR+q
mfjYOewvbSGVHRZZ0+3+II6poBmsscdXse1fWz2EN5PtDciNGzUcapmJ6azo
lyhd5e0e+ziUw6Ltjmc88OQ/TVZiJdr5GMV8NB8ozKb2PVW+OJUDAqH9ENtW
qOy9Tr0Fk5sDx2t3Pw8jCkHl7MqNXapOGGcU9FG08LSFl6zX6rviss7aCb01
vVznSruPGIrwGbFoDpna9mVpeVGn0DIYZUDOKbbdSWAsFN4rVDWVfLjlG64R
ZF+IhhIJyHYRC2QX2eny+DxcTRjZpocKaGimGDct/PKVsHCWP15rgxIx0xkL
ZEv7rxz2lz32Dxp+VPVWPAZ62DNXKe2PeuAkl7K1JfiZFtSowftww4KGnX8T
qdedHx1xMEEH7dF2OZnwMq64TFWYru102TbL6TsL5y0LmdilUQrEQ993mOlx
rRiDGB9M+R5jLTOIR4mUNZuOnjALpSMcnwtfa0tFp+7C4MN5eJfsEbYCnzKh
GqmFcqyFA8qFXGXbvHSyH6Kam0Ka/oloZmWbqUENPgZIFAKSDfckXZi83QQd
kUHFJZftTiedx7jm55lRhkddrArfLKVqKeiURmn9gv0ae/94FVWTfs8ph/N3
Dma0HjYJxDedccZFX6qs+BlsCt2HZG3vB8bhfe22CYLMTbAeJ/REjA2wVr7V
vGIr5M5tp+d7ZDg9NrzrhpTQh47XloTAk9vyZLstbPIlGAFLGIH5AZrX2YF2
m4a89y3JA/fumN8ISJ0Mu3DXatIajZyduLNYpBgLA0wZK/F2h16nkadzRnPE
NKwfLJ6h9lphfHPyTC68dBZC1FXsmK8TCetcppvziCf1AUhNAlA0F0Xo6wW1
U0+/Ll7YP6tHHc2SkIcDbkEf1jRPXEzhA5WM8aabVf69ss34cZ/+FtGmwLtA
RaQPCwSUu/bOBjYOc0KSFADiDGyDG0u+9/BGk/FAlQF83laqvvHYY3s7RN2D
A7tHQ0Mmo1TU3WUGuIGQVmStw9mfsEekwnRJIhRsPvb6ET+2GTdlvcyBPSAD
1Ds6RLVkb4ItB2UdWfFRhNg3ZJOwBoEKuV22ZG44LYMGR4Py2I874dbvmS9k
aIlJg5XDVormaZaB15NhrlhouYMNST9F6mlqwd4LH5gXkzk2qN12e4GN04JS
Ped87m6ZcD0upw258e7ZXmHBYZjNgJLxnpaEJ+ZHPjvyjmvT5/dEw6NWLbKt
QnEb7dMqOE+zzwANapk23NTBjzkd1q5oOfU2o9yv2oTvoQ1fcp3/gwzNO7CJ
LcCIUuiWFsePY2GCBflIHqbYfbae6tU5owEa5kv3F2es5xKvO6wn66aUTJqr
vBo3HWlkhTSyooSrcq/TXhJCLvWSq6RfQmUCTjQpLJVTaaB6daZ4r+MqDUeI
My2vFIUtYnqsXoaTpkQKDdqmwXbgHW9Xma4dzMK7ZDYsdUPy2G3liwplDIz8
kcCgBvga/AtmK7OW9J/DMLki2fs8GLKn+a0rHUivQYQnV8WAavyUZRV+PGuK
DuYD9wyp6TRckwFMp4fPdJQK33ZYtcByu9ybaPBXw7amAwHK84+Y31LXD0nF
22DVN3f0TE6hH4XsSqVy+1Ke2V/V2qoOZACYS/0qp3b60PxxGYNNSuHKZvle
2cccMWIVBSpZ38btD+Z02NMl4l+k17Jj7h14PRUFi0H4Wb/vExcVEbZ797+L
WNTqEMmS8vshIHbBZ3eFUXYsFQYK4b0O88gpu3XoilEU8sk1HQV83dMOBkEp
sKfRIwyZV/SL495NuWNtSPnq392a0ejbhUsKeUyyIVfq4pFF00TFFgEhnHMy
/1PWk22eSjktF4KQ8XIulIIY0oaQGbB1O1pn4dg3g4ycHdj2HAur1S84KgDR
TcbK6OX2Wkk9JwTJ7XZmcoszQ1qgyeMKl++nZsGblFFB2yagANBzjFCSNuGd
xoQesVmj7j88PCEpzvO/HDgZbM7EayaoZCAEIuwm/68n8C/eePBAw9/lB7pN
sVf+zP7/tEKYj+uyOK/mgyDLCcvrMZRRGvt41d24mG4Z7pWUyEbN2IwtjjIs
FfEgUHZuk6d12t5wMRC6K4FBSBuNr7Ey56fHV32SfF3MHrCOKsYCm1tnAuk+
SzTzgzf7MTOON7cd4o0g8Sjy0MkLHqWyXiZjHimyzYsOpHr7p3NVIJjYKbMk
mcK+gof0CQF8bzDm/pfeykZv+p9Rvp/4GfalZXWWFwHJ/Fun7fhLIIyR4Iba
1ZLlcBpizmeqON7oE4JKOojMRolCNnmJY2bifciQ3I0zm7YWCaeDH/yqJoQL
DkS0TO6K0q/3qAisvZEwhPbTlV0sWa40P4n1V/NaPj8wBMBdzoR+YjAidiay
YsKjUFWdHyoSs6RR+cosIu+o+ikAdf6RptpMftzvrMIS097hFNPVM2TPZcnr
gCoNsW0Ey51Ed3bxYCupoR2RjkaNj4QewfMbsa++Yz03oyffnoiRkNdJ+zqI
U+7TWm3M+S9ubq5w+xIQlGXC68dY3sj2fZ7vJeChEKCgsJ5Mj8wImLdcgt2D
P1PoN1YzC9jKPZt35VDZR9iNY2G8SK/MyHqgk6k209tlPg8gK9oLJ11Brz7f
HH/3inacdXPm3gza83fUzhTLKIYeS67gqXWY9INOeT3xWvkcjn0JCudFtZ0Q
iibNwaSmq4eo1tSbLqdp39blh0P+LTHtHKXf+9Ly9FMtFHZKTNL+bXsCi9wQ
R4+NOI+mUMe5sH/E7tOaerIyYtz/ltIwxkcRmEtzUdFxCtgBaqWuJr8kG1IR
6PG27YgfvBO+VnadNSOOLHsjsasdfKHrTIOOrQsZ5F03tknA08vxEN0AnAol
AqLJiV6rQeo9Fh4SFWJfy3wO7LJ/IIvodDjnw9rpJF7ONfVnobDhsXeMeOoE
Ou/1WSwIZdGuRpfkORMtBLTqXXnt3i9hqyJgDyYRZjbZoO8f3iZ+BHcJR2zc
CCxUiQyIKk3REpQD6vVN/dP3ofEVdwtIh4yjpol2iutfCDvx6FEv7HPIgFRi
z1uzPcT12rSHgJrDXxHDCj0I6/c1o6WohjxziVtKowPmFoPgHdm4Eo1xxzwl
SpvhmRUMsHIxeNuxSt7M02NainYHi+tgLDCCrbvh2JkIE4t0hDfeNE/5mGXU
wem4+akldcCtTc698qbuYQIvUjOV19SJ5YMFdM+JdlmOKkOOzKSumMxMjsyW
ZeQj5cHjTnaV5BNymI1kflhl8koWZQV3yfp8mJPhZG8+Rh5PcBVyCw97EDL6
/iJzmoTvYQNFn49YRErWzZqKFwI/jNGvErEY8TNZOGnlBSJ/++uFrscHBQeY
FdMKkq0r/gGD2V1wL+wrqLllCxzGC6pGw7ai95hXg1Is26h35/ypKCpG68Xi
WudvP4FfzT4NNHcdELZamAFDR84sVzX5Wj3sJOFq5Xg0ly/Oe3gJObgLb5Vn
1YVUopXnRP/TesySZV8Ru2LOkWUdA8oekxMXO2kWlhfYJ0AQRkH/hqB3ByEH
iSydJHgxB536+nyR90IUDEjeZY1vuOA3QjcFrzq1NmNfN6Y5kkzrqJcV66+W
6nLnU7loFzSMwThvpVaIsCQ1HrMzqAFWff2mKPheOiXrU+JRFKNyHg4zax/9
ihYC++LeRvMcnbaSwml+SCD9yEvnKZ2tVmjlyzur22BpjJCYpQqdij3iz7Ge
wS/M/VI+s5vUgai5bSQsEFrCiX3cBxDBN4qIX5Nf8jxa6FFMpSZLH8yiBMgM
dEZNnLfPU8RD7gx8yD2MS9E5mT0JZ8HbXO0roNQPqnddJEUed2U8QcoWMK8b
fa9zw6HPI/nHdNY2xAN2bdrkW9oX4duWM7VB0K71E2ZX0jXMVE71IK9CQR/K
dS3fdukNiI5awxyeG1cvSXsFF1NKw8tfIB6CtILOxsKuehhWct3ElI+kw7pM
KDLXfa3nOVOWagXn3v7UkcGjb4tCxAECf/rAFVqBvug04+F0jEWGlFA0Iix1
S2VPM+lynEcLvlFpWXW8E+2GTqiMpS4+l9AFywEt3oJu5YlVc17wjb1NE+Dz
bD+vXwBC1LjinntjzmBd+XH2reqAZrErjWN/JMQqU7OderckP1IkGD5QMKw7
jy+7AvNWFWZBmQWbw09qRqlB6eI9uOwyTK8sDGXrs8gdEJzFCi3hbCSksApm
4q77ZYVWkRL+2vifoboBH/BfUNzTXohVYoQNsR5/O9VOoSDoDyM3lhryEJGo
fg4vTYgUpyuJW+QH6tAD8fKT8Egp46yPZZ7bcEvP1QlP47Y2XyqH8Yu0km6T
Y9DMI32q++BL8ZyX5ih9gebNkybtuEMaPjsT62tPY9hGM6JRyMhrcjLmnKTx
2eTci0tG+3axYOBbEzqckn3nVk1/gRw2FRWKprCRNbPitPWWpkJqnbctlZ29
Kn2JAehKDDV51DqGjzs2i75ecLW85HmbMjlWREi/NU1cRZTSOokrDEzbVNkf
7FP9/8LXHGCtmqCn/Y8AEtCaddyq4hreaAKky+1I2EoGsgbHPNRj3234h5Ic
WpP8LKO9lqNFnTCKUoJnKD9CVXzPQAPxQNk6I46B0A5ef0CiVybmEYNw7GHF
UmgIR5GV3zzcGstF1/g9Xpe0WOqWCoJKuHkB6UYu+ANfG3/vJYlSPd41+Ash
Z4VRo3HK8tzO5obcZNOffed8DilwPK/PWn75+XW631Kln2MPuNnumglnzn8E
bMgpXh6s8B8Hhut0/V1ZfkgLubNY9uUlEZZYhTMY6oFknrn6k1OGaPl6OGnR
jYFQ2lhwYa22YnWSG6M6RM7UjQdxeEV0pyf7lx7Y7LTum2GcVNfX25FWKPsY
60jJE0qaxtqI3SABlN0vlH3C99o1f5JycW3TNNZNQ4TSo8bN47EwVRH/KOPv
yLZi/xKtMBZakve8Rb9h+fufYXlSP+59paqKUjw3KqlPH0eLxDC4QGQN3Z8R
omD4i8hAgsWhWms8v46WyyPgKxvouLkNoI8MB3Ped60pQ+KQCLhP6nAWKy1S
E59YK1tDWr98Ns+jNvzxV2h08XJS4//PiLoHyGl+LCMwEq23uoP7YD4xIo0s
LuxUsYO1+HTW4kMYstV0DWWe1UE7IV2BMD3AClzxSLZxvP17Wbk78/Yhx6El
dzRfNgj6oQgzSilc0YMtkYiDy+0A+2KcQZy1qmPVnfQKzNVPzLaTSnsDSmNn
8z6wh1dcUm3ql7Ei3iklLJch1NqJwHQWPlhhSFTNf2mwEC20E4ZZA9VB6hbw
t9y5QF/EaZGpJkTEPwj0H+BxK58bgOLV+37rdfreUj8zuj+5e7quALVBuH95
ke4q0bzKxkypl6HNuu+RT6JtwxB2C57CBbavGjH4MNfTat0Cc0CwvIXuc/54
ouqlKIu10OZW4FaeWdTuR8MCtJjlwloOvAHJrrqq+/B4A3Mcjvzntv3l3Mas
2vC77HQS4KBpvSoeaNh2NNP5p1Z7zszjnB9kZ2e1LBC6lPUN2n5YjzK10woi
r2+16RSsiABSZv7ihvIXU8i2IKFsEiUbbUf/mJfFVnYb2tFKgPdv6Nn5GKtK
zZ9S4DiRRiJ6066o1OTeIwKttq9/EWQypgW6hSKz2jqTL9fgn3YnW3BVvNyg
GAxUzHxHn7qInQxl63qM0AIA+7TRCAEPRbpdc5jY9UrV3fM7mirkuAN/o7dP
J3EEc/pY+mg/sbgTA84Aj++oaTqtmJlYzM0U2ylGdphXO1KLL0a5d/l/NF3t
40kdKp3/jre6Tf2fBSwzCwUDD09ii2cXshxfcrSP54ZGIjKPH6SF9dHDDW4c
f74BUA1jmc+FHSYf3M5Rzrm99xwkbZfp4IwNqakhkmui9fWq+vAGwAGzJVoe
/MBa79GEE32UyXqTjw3eFhjGPi10PAGFhcfMD9xfCOalW0NSExllwGwRfmG6
dKnLeizsAfpxezz5Ae/D+90x5OK/O2/n9rRAdCzIKBLFrhGazN9J82+ZJWY8
3gEkXmP44hUgNnVj8Gne5nwZmP9jwAZ8WxEPLUWn3yJ870ksWuX4R68Pl0jy
fJOAA9yTpKry2W+njIHbHrRiGBgHtwXOpzSrtuFOnC1Ok+jwLJ8tQf3/YBoz
HZvnqMrR+MpojybjBC2uSVAevj43Mt7FDbTecbsvHAU/lMNOl3bCbeTBhwP3
OnY6tFKSV0uc0Wz5oR+q/G8OOd0fIzwDr3pbtJ2JUQOC/mEQjVlxEtk3IXm/
o1jZJuw1lEIVqB3HnlGQkGe7A8EYir2Jr2VBVYkQrGkeI8/XlyTycj9l8H/x
miEJjZ2OYYAxY1Yhyd8neNxvSGynXd0u4LghzW3jH+tPUobK7RppMKXqHFvf
dGySYq7SQU6qYaSW3IDoPAQogXHfK6NfxiG0LYfekKqNUxPQ5xFjqtNHQAsp
LVVWh7z+hRcVMDu+DpWMs+rfJK0yUk+H9PeXbLzWoaSr4AIFImbgRtPZbZm4
FZVNiSDokjBUMIcL2K1Ymlz4yIhQ9K5oFrpYinTMpYMEJFkrESziL6AQu+gI
qObTTkr3CN+zru5DQbsfYaHVtv11qyxUxuwOxhcpd0fQzcQWgMo3tVUBbatU
qon5mgBwd6Ql2tUNebyjUkiholpkkX1LnMjflxf/hRshh/xG3vi8LEe/VHDV
oN7vxX3BRRA4NjCIfAG88e84ghv5PUcPgq22k1X1WUsE4Iy1bpSzC5SxDKgc
42V1IZAhXNxLV4DUuqbPEC706r6YDI0YeeSXbW116cniT1vt81VeZNFlefjG
GkFYNfWaNs+GyWODpxcCGmNuZU36OSapHicBNqg4OM5l9Hfb2eeNc80ov53S
UOODcBjZx8BobeiWC/8BIVrG/giDHeoHMguSXhAHsWv2vLcMS6JiGz7piKEy
+KlY8A7OXmv1prepLeek6oyVRMfd8V7H8zIeurXXgVOXCvcUWBc/RaYCvP+E
y7S5sgVlHb6FxVRlxewfGm6u1QZqySFSPD26eRNdIoyZXYPL2Dwnq65xYVdu
26uAvxM0BWc+MYK7l2dqgk29vSWcqnbO6QXd0Y1iaUI3UOxa7cRvG2C/ZTPr
lL7+T9sSTL74hfUObP2F8srH4p3Qa1Q/SZgsUqH5JF5gmCtVBtw+nUO3IAa+
BTu91J789Vfcp9e5s/tqk58HIWtPTFU23yb8G0b43RcOA2801RImnK2MbD4i
HDMc/3dfEiwu4CA8pI3RaXwBoewWklI0x1ObJqPnPo8EPG77pE0uBdjC3Fz2
8PwhfIXrIVhPGMs0xmCnlWvGP/KlnHasBgfUMW7ebrZJk7LSY5fn2W5U4bns
MJsijxvdQnnbs7zAHRvPrPwg/XFpWgLvzEUzovr2nghN0a8vgrrFn9t5SEzu
vqwxihYiad2hjXDOAYL92y6EjsR1L2+Q7tWsMkKJD7REoT6/1PdY7duP4E/H
xH8qTANNW1U9chc6ktmAYPbxkmDRfBTrBXuxfH2ctDKchOyjJLcYRYlbS2kL
NUEuP3OIvAHXPrfSMtNGmLI1A/eEa+mDJS+J78UkWTRxgICxcW3ZxU7InoPn
9o6FoYJOZIaWfpWaUPc8Q+HOVZtdK+gS7XI+1YO9vGUzv014rs4ME9XPhuYu
Pcs1u1JWr7LltTk9HKX8UwErz3D1ZeRCm+klBzDwAsYmbWLKBxRzxtIp7U3t
RzVqzSgDE1wGUA8LJNAS7HxXn22xh9KcmIIe968Ku8+jb81kwV9nRJbtMz2x
sJZNkjgKN2ftjAoV+a7amjYUF76za8A5dLt63+vn6lZJsdddKU28U9L9igZP
aHj4mnEcrea+jNsXmLwxZDhuQhXTtEQuVmCHcqKvF/ZBDD0sm2vOM7B0lufG
jZtI0d1HOtnQRMJk0GdL8VnIRmKeZBHZvgh+c/hrVJBhMipB5r41v33DJdvY
2qTsRkAzujMzQ1WxfB3WNxuzqekaUQDTLVSIdY96U2xoOfhBzKqWsX9apxYS
gD+hl8MA3mDb+K2BsxcVWmng6dxraILoViC4aItG8RfsHtmikjrzUS8dp7SJ
7tW0Nc2Aq/l1KuJmShIKIL+BMbCGUoTC4Y5f1HUWT1W0Cy+3Xqw1V3jLB67L
/LdVIaEyfSc3ALskAJk6vGWqGMlRvsfzvMencFpYHMLo9ZPoPqSS5V0HtTrx
oxr8o+THi1oIIt3As6TMEE/AbeS1OH/LRJPgmzLWLkp8zFCSm2Tut2aNcLa6
wU8ejdtrUzsLAklYvM0NYwqJGJ/67zHFzAQToWQsVEOFErIVnY5Vb9AxptVb
wpVqZE+4BDO6fJXfCPUtsRafcaYj2J5hEY8e8B6hmMw5oS7+R7F3/BOuWywi
OdDOEeeUT9F7B8c26+dpPUMFoon+cwqNSkDOkdWeD60WETzcTjogGiZUlt6i
xz2X+q47arE6udcGjLV1O2S2q05PyEuWEBr3rt9umOiyE/Ef3aVSRcuxfyk3
ZqiBR/vxq4EvHOLQIadVfn2B1h+pJy4wQeFZRnf3crCkVignhxj781gqO0gu
Ke8OFYrfKa7H3a2lhZOY0hiTPznnYgGlBvk/q8sgDm0YQNvkpMBBeXf45glL
HNpQKuTNoEXEvG/cBxGe29qN1eD1bLPKzX8CKDIFwQfAJJNRTcgckFysDBS8
0tcrmVTZlpLnfgN3eOMmyxrHOVlouLHEEjBkVoGzIxhm1WKnig9MnPkLju55
+KTjBUmj8m4QtrKaHs597PtXXvkmlsnwuDj5Ob7hFaFKe/fqxaNi6RySe7Of
bdgNi4i91VQfPbeU6fPulVXcUDOJvJi0gMfb9cumVPFDs/+otjf/y+cwpJwD
NTJnPhM8DKiZYJ6zlEm47fNv6iDzUX+TFSs3UcuhLpJqf4xQHDUohVLFlYoL
k1kmXNM19xyEXhqlEFCNI7erLp0AQOIS2MEj41gzkr9GKYtC02aYKABcr1pb
z7QQz7urZBK9pDxrb1WzA47D3JomJsPBufJjhniO5ZxXRc+MJILrJpSCfiZb
Z7qcPjY+xZw0ry7cdklbhmfiYepwTVI5MMkejPhbZypOAEgli/iqcM1qod2f
wxlq0SkSEpjkTsHRthrOP14OOtHkTWC4qvTviMQUEIAGf8ImqZOQR+dWIUd9
Mwt9zuw1Lqjv00gRLNn8vLbyAqkwn3oFOHTaXumDZrgxlYwb/I9nIVvUMUlo
yvKMz848d/IUTrbqUrgQ6X9ns4wHhlK/cMJRp3STn+P0Kd3RELgrI19Fpk4n
n/apnPMex7gukuUgPrXVgRnGyb2CkfX8v//01sYepFgmt4Y2aAbUwXa4Vs94
97RoFTR9r6cnqZWEawnEE0iDTRqaBVjoV3fltXxri0dnsWgBswBvd8ma3kSi
OFRJg+iFnaPbZVxa6J6n54INslaKCLSWIImUGPRzpN496xiiX19Enz9tQfRE
lrBsN5yq4qEIVs7/7kkFhMgbbcO9/CDNWpXihMrb88HtMEDlbWRsXPbXIrX7
KeRHq8HHOy958eLauF54xQhJuPB0C6kyGEU0k4lhwBK80EbaIOKqqDwjRcqZ
b0De1tI296L3FKE8m88epuuk7oA8NZor0Hqf3X/lsQav+iC3wwgIxM+p5pfs
OkZ3ea139xRD70G87WtKM3vRCRLe+hjIp/MeNUGfPGwd/GEJGUze40vNGiAC
LGiqzdHZQk6um88aMI+g2IWJ/F3XtTyF5i9H+aPwZeEnPYkGCrqH/Xj5uvul
G0Ej/cQ+fcmLpc4l7Qch9TuqmXA9ptNkSOGOvzegKfQKaHgK3lPP2ZYtKuOq
nkwoI0LWrtoHwIpOlRJ7qMfaqw16czRI93oQM1t82Bu0tUR976YddvjiZINh
cgCJjig6htirf1Ej8rtycPnQPWYxty7n2EIYkWHi6mNzUJwTrICmzFAh7AO+
YzlqrEPbMfS9mqPW1Un35x4GKm3obhLE6409sVKqRgrLiB+XgSYavznTuZVI
XDfADNY+qM+U27iYHig5iiaCwOL9rN/mXH3fmtDHlQ6I/c1fM9VnnTv9VokV
RkxZ3Wxmz7zk2V1UsTb8kVEj3Wtkih0UOWtnynxiqLAj9HjRMV7tViZiEl+X
O4zOOLJgP63dugXCBAnaNtS9Iilble+v64G3LDRxEwRHigpvGhxVTkiEvjeZ
GXC6+B5batBmqauP6BHPO6nFbfxAP/OJQzzIy+cyzaeQng2QlMAj0GdJP5Lc
sReZEumbqh8mdRtNwx8z0WvVtpMNTSmVT47iCQIc5b449kOj8shNrgPxlPCr
WNHXn9R3TYvPLkxtWn5vpGLsobeH0KNbdo4cpxv07lR5CC3oGU2piAHsW3sd
U/QqFEN8zc8xHxayl6uBYCvti1D5mIcC1F3keKDC1WZM9Mc5XdRkiVo+l33G
ZIfJEaKwLDJnv5bznt2LFWF6KUzOJwp8BTbjd9Nw+G5yWKGXLuQtZ8Ro+l/a
RZUnfX55E2Tp6xVV0xfYSG9WCwV9u3BqNYhHqXjyBJu9q90ryRq40MvAwZV4
rxbSCtOHzithqBk5BlYr7mT0Poprk/NrfSzQSbmiPmNvrTVy0QGVM6adqjvO
wSbHeuzZT5/ElJV6LjbG3rNRg4GdDmvQh8FqDwRIDFDR42gSY42+m75oRP1c
IPxlzMOWbb+tOHS5AM+OuT7QEq6ReGNwI4B5nOkYiRXXMcH5IFGfyfTPqAvl
++3p6vvNmvxPKzSzVzpVjykgUZaHmVFFH06KWum/LqVJewmokXOdMpcApzNo
ROipQF2q/5i1toZBHtyi5AaE71MzbyQ1LlqkkcQl5DLYHZ3+n5r+3IDdmzuA
3vCOjT/lLsen7YDU/4TSPlPkqQgjNAGz/DvpN94jY25ExxMLcGDy0hrX5sWq
bhv3fDgkPSQlq/P6EtcF1aOmmSNx03oarF8r+Gqq8tOj6lqeEIGevIdljMgi
rUp4gZH+lXAv+OsDiiV+HyFVgGGWDP/sHrFr3/xiUlQZ/vJaJDVWm6g5mYI8
oj7szdATvkNpwSz8mWackJplDPBYpd26j+NbGrtvhK0h/oa6JvpmEbln14L8
LsomiY5lJq5LZ2iJmJwrxAdEtkZ9Su+tk28sVu9yQHlCvoNiGsgvKZLvqTGn
zGlWu6k+mO3gT/AWyjbJORY5tZY49y42wFzCO2cWIKRIlWU5JUmdorS/i4kM
ZtkQgDs3nTY1nKoMkCxeqtUDqXQugQD2I1qtwe1lyXaJbZpXlQOSG+F/FM3r
KFuxnn7KBbgs+2xsI7+K0flPhffoQ0MLWAwx20bjzZjptTiH30wAqeZBYSXm
oCZGGiRRKt+bGSKGI5VhMSTvELkgBAqs9a5Ug6kFtRt1DClnbRiQdoKSv45Q
pImwktwGcEc8e/XpyssqQjZXBz6gdfqzvsILMgOh/F1zIl8rtaD17Jcs5b/h
L5LpKbNZSJOejT0Q0ki7AQbbelC8cXP2KTA+xolNL4EjisfD0U6dr3fseJGC
7sFdutITE1PvZps3qM/x0juAyU6qk70wUC5aLuhuvBU9xNaw3u4VaTxB4hdX
WfY+5ok5lGyPQbFuxfE1SwgokWGoIzFrUgWBUb07idmRViz0I6pAwes6v1VJ
6/osuajcnOHt5FQWbzDEp5iqrSkDjU4VqqAmqBulgf1e0UfTKB0zOFGXOHww
8MQ06D2Dl+KZvcedix3fEnVJFukgNyD6Oszrm+w9g18xEHShdkLl2l0zcRaY
UP+jRqfwzyEXMNdHKuSPnhKFPm4pAoM8fCAx4FyGvITP7C672uYuKWFtzmT3
fdgbwKnYiJIWc657Qzgo4FgB06G1ps88CQIhQwn2Rb0OlU29AK+x4+6eZKjU
jZDDDkgkSONm+0ouBHSYB0wUHK7LXv3j2FvdzMa/DSHYDGM+BQ1NaviE2bCc
LojjpK2WnPZKcSzRJ297tmbQiL6EvLrbI7UpLjO+sANhhs3xslfCIBURP0S0
cStur1PCmt7PcedWAUFxtO1hKVmAci26s7HgT6Uwk8W1RSKEbWP8xpP/vaIQ
ZltAIW0BhMt5+ZTeYoz5e2kRBeoioTLyFQjN6mwdKjBfc61EfVkMl/AQxt0b
coBG1UjqdyqldC2EbXpVUnOjxoD/8shcs5NLkTVIirBeHllIuv7dfRH/K9bD
SJkVxZb7y5wXxC0Vh4SRDA5r5xMFhMt7NU1CR7LvuRnLnztMMSF5x3WwrdUM
TbCElV0SO+MJnpFFr/QOhOaHiPywe+ObxqcXaf1GFUoBBp/5IZsyLVKUKN7U
rHjYA6n0aXDhizbJe0I65PR8cZgZgVNgcyTRPaLlAK8mhzpZrX4/P0u9eMRD
oR8LzgB7UgUyQ9ly0Evr90P66VXpXB2kqVxISfs1Na5dHo8/7SX6S6s4Ovyh
1bm6DjPB87rRX8SfUF2q8UV/D1ZXoGZBE/JfQ5kPwQzDNTbMH/MzvHuOVOtR
AZJ9PXYNShwAM+1/9SVxzleCljHRSbXefSftX26RbF6QJw7eFlmLab+UFsNR
gexcNN7KGbqbxFJJaPWQFiAv8JF/IZZ4Pr+WXhzwNWw/BW9jjBYsZEEQsXbV
Aj8Sk7hkg4vd/IqihkdYQaLrxE1/uQen09k2zNl2E6PQQlhZx8H57P6Sf4Sq
3DJfZN80zCMxZ+WP4IlyJPOfYdrz4rC8phIChTMV2V2mZPdZ1QdG3Z2uxVlV
lR73p9RrtGXZvr2q3pDUyQof76xIxtNJf8qDkHO+gB7oUHlci6tGRFOlCErV
1nCl8+3AUWh9qN0iIDb2aUQnEXlPd2z7PRBogpn+YReFoy7wrszdyN8urnue
feuacV2y9kL9KotZgQ2tiuna+K4zupnmxaqvrRvfRdW14+L0II3x2JIvB7oL
opLju3Wj39hQGzjHpgrkZr7IhtNcTKiyYRfZH6qIFfqznF+pEp15zupDrrbH
g0iUXUroU0bfituddrdTgW3a7MlRWQsMje5LD1SySADtFqhgob4MQF4tTX9v
CZwgLACksMwkbMd6e2khk7kpBa5sZ5AHA/lgqojDX5Fbn55quoND+ezAgE84
B90o/fVXtCd5qUeP1vV8Uwgx4fljU8Y9PbmeKOeCGrbJaSMbLUHoZY8pBoS3
yEFYKPexLVVg2NoweXf9zKoZrmkf7pTJg+TcHJMO4MYzCbpKLvVuLXl6ZiRJ
5mlSgipEovbg49ARpRQs8VDn/dlDK+wF36VBwGGVau6KTumF6ItaKE3cslT3
c9/kPU32Wi68rxu3Al3Ycf51g4VEM/4IiYuuLElNg3ML8h856PGG46s4J4A0
AEZTooSzgI0cMbc/d5A8RmwsFbU0qR+YSJfSYoD0kdDTlMjsRmBEooKt6134
Sl1U6S7KNKcMbpdYsDuF/Pu6VhrK6D7ggOtkLvNa/fDWBFGRlPqbkrh33Ei1
REM7sHq0Tz7A7osiqxYCUZW69aHMiVeQtSQL1+5BbqeN/BWyeaNH2RrLPHf2
n3a40y6JxiTHQX9CM+WNQdJyQGL1OOjba7EkKO/0UQxDD1gx08lYVmNLQwON
/l8ofRDb/o+3JVdcmE5JLcRagrFnRkgRaN76Jvswz9Z84I5kR0RXQ37JuY/t
53C9FYIh1NvffHjqDnuFggoK1taLBgmGSwNfD/VosMkt9cFIekxvL2PBJsXG
ktLuAsvTRjlJz/SZk9nPH+OZ1H4KY/Fvzz+EH7GPjApo5EWSc5uHt3MpjO/o
xMrATPEsAMmeawB9DQNBOHNFk0dUCbxExDqk8ONxi2u5xWRHtMHxjZNrROwY
XxAxaDFRQKZEVIk4V+0rMH9ubCfTIaUqAqpKcsyuk8PskrujvzDINFRqvLca
MnxhllEkjaceZ4yxdpB+DzqRKsTFUE5hJ8HEcElmF7bHew0qXgEPliYn/Sl7
RFSVmfzmkzHTN2vOX5LlxZYki2k1/x41tI3DSvSlOZC4Qk2UfsBwfKakpVWF
278NYV9JvtSEu2RpLCNjcDmV9BsD2an8phx9HCZ7SKlQd+623EydjF3ZE3E0
pkrMmNjl0gbCHnA6nGGLTmz6OE5COEO9eeAfuXtTHKqWhUM298E6+tVBF+BX
eewQqKwS+5XFj0LuEHxEmqu4yTk8mFyvmqKDiWj2ZVlTJlcC2oPCpmXeAn23
wmCT+5QQ1ZvY3HxavCurXpVgrk/aesHGJPo4HEB5RS9yxQYbtZj2lH6DSvA3
zF7jNL1IlajeNRKtJNjWUTe5s1RYFMH7AGtUO/xbPBUC4HUDG9urILrJMye1
bCsZ/JOwrR+VrNZe3Kozhohu/CLSIFbYsw9xsAgO7lp0uTu4vpihlcnoOKsS
3/IFXXl9ytZr+Abp2U1B1rBtoUChWX2puWqvOffGQhpce4uBjbdsjUzyURpc
BXViwziE0x/2U90MaQcrBzvvTg5OOowph2vMbR9kZM2b2fkBT6dcknZuJqAC
DydE54jyN0Z1hdW+HiebYIB0r4BXJktPU5VlM5i28yrpl5IxxrLPJcFHP/Dd
Q5Ich6ZUdAuvslx05pmzAJI1nP+wY8BX9X96ITb1MHNsbc0Z2SCqXZPjvXox
8UsmXw4d3gt4oQlSr+9rop+VvyZcBHKQewps6+GySZssbFgFtqGbcJzmsouO
IUZrNC4NKnSvg6M8xXKX6THtArYGKeiLbyC3a8VedYT1i194toXupNFmjRwY
SYfVXAWEhDsWFVCqbI3IE+OjOJNV9njNsEGQItrK/uC6JraefwgP0QyOpIsP
f7znK6nMTpjUfSIFGUS8NddFvRxevTKUDbejrnthOTLGghUyKLXRQe/en+iG
+FZbIAy8brQNRUwTfBZ2wg59306lK4ky4Vhf+pdV3vWjySW1/Z2XKOT4ztyw
ou3GbdUgcHAtWMHHXY2FkaLY39nMgKhBDcT4nXP463w9+VfkuafC2pd50Gru
ABvM7Q+uic6BB50Vhaf0MJPfS10vQ+CvpKtFw0hy/cj4eX0kcTpZGpzQaT5X
FiYccod1X8Y7r4ycT8Qy4ifnb+jBjuHmssx6Q/iJ0kYJvrKwQCZXTo7yqZYr
xYfYS1r4eSuvWZvLsvtPPZLAMeXJmxIvGbnNCLqlkqCabvdphKhgBIucafzz
yUKonCZmgX+xAyPCGFGZRKZkflwm257uz5psApiBCK1xIo17hulK3+iccgzc
QuVhyebUPuG1GQhxUI+QWAUwSNZLCiNjRBPIkUWINM4OzySkP/XyBkSZ3VNp
6SYY2HdW85MDj88v2I0wd0QEnvcAIiVR8rakFPPWuSvXAY4Ks3wFJP3S0iSK
JYPlYs8PwQ0fx1TNM68truGopPoErNEuVwz2E7w78mx0/nVh7e1kc1jpZ4uR
zwbi567bg0iRHuXxo/Ptvw/05UY9SDB657xppzcGlN3ChUrmLy8mSQOehN2m
S/CK4srmHTEsOZerKu3qvbLvSAvQJttoiyLMaduORD9q/wX2MQQpR7iJznPP
NU4nsSzt5D3T4WNda3r3iTcjnNqHN61ds/Lcca2DaeZHpY0SpYlfyA6n/KMT
gN05RvEyWGGnzzppe55gIEYszWiWG+VB46TmKlcxCIpz89Zzdfx61imb4AHV
zDWgwZOGu1X1vWDC43CgLBBx9uRnnUDdb2mTUzda7i9myt4dqAc3WaKRXlPl
xMtXiCbZhAynK7XXHKOINrldb8zCLbfq16KThA/URby6MCEevSf0afX7mmdi
hVIKCqfdZbGY0FzWp2DuC/8AsCSAtYqMU2183eBpH1hRI3Xq/0YSRB5Xp01g
aTg7GgmzipykDnLxVp7+J7ccebzriL4GuxZKQmRMl4mlHghVv2gS6Nfs4bxI
Kxu1ym6EMLIooE+pc57SjdjgWslKClUO9TnYqJjpAQ7TULzllpXH7ybgFHjN
RiNy4EeOmMHc1457jSAYI9LGLZSh5Ge/0N3jiRzKuyejziLoj9gVYVDwzd58
OhdvlVCtDsNZp8Ixq53Y2N4GZt4TUjd1e17BEvK0EAhHBuc9C1MyGVCwv2Wn
psYzxCeGEsn69zN6oPsmSuAkr7JBEhPtXMWJMsIVQYuJEgEiNMyoBj5DQA+Z
ANLkN13Ap2sRlasayAzKG3EMXGwpwRamgyfc9SuOubHJSgz5CrWpxuiWgQv4
/iJ4YCXgDf6h49NQHu7vtX5qaIgl7wVoAiAenUET1c8nVJB1flp+52TIedB5
6jKOyoFwxG7Go28ucyKnV1hwr091DaD3lYdj68IK4DTd482uXA1wn127c16Y
8X4txU5Csfv+xMu5k1VvufY2S7nBA3US9OQ82A8beuaRNia4XUOyBafvjErI
3FqJyKY7IliFTNZ8DKh8WSAtb5/yHNEyOQXWAOFhlyrwXcX5KNeOGAphl2d5
IucJ6r1FhP8efuWdN7XSPgioOxWvr67BDXeZLv+CP1cfsMV1OnPZDFBO3gyY
BvMZW6r5oH1v4HHNpCNxkPg/XDbLjA8Seh7q6+9yxVvRm9jv6qL6B5INu5wn
HKJYEgM2SU62orsExoxikaaW71ovVBk+9txAQdZA1uXEqy3I4m/glk6A49pk
ufsL3nV9CfHn6IQTc9VU/Y6F7q+RVkSpHc0nfNb0AAlgNgp00FU0qAkOlDVt
XpkFSGVjoj+7Rjt0Ye67MYj9NCSEsf1lCWzvBeEtARsjmj07paqq3msuvvGQ
bsLfY/TVCRl5xgd5JkRmE67msF1cfDJIQMoAgvaX5lOF4kj914NDgI3PzpLX
TQjXUcFUbY62XPFfKozG6yEEO1yqwTHIiCfZgHGwF9Uod4Cdl3T87jTS3Enb
a8a/PtyBMUnjHj9IaoqnhifRPzo1x6i9JAm5NdxmEKZUMAWwZkY5h54F4r/z
pKXR/kyTTpw1wodBqSNgkoSmqqHAnDhM3L4dh9kF5sPae23utPJfD8I7JI8x
sNkXfL/pgF87VhNJLP+j3lNVpPkBNN5fp0gb1/PbyE3ZiBJHJy1P3kywV+BS
X2SqyZ3fgKxdvMjmOxbvyl15PlSRkNCoVZg67Um+BwUAdVHfPUgtjO3KUJho
08PH5xElo0208KCMBkzuJ8f279JQ2E8mj5XF110okcInl+t6pj7QDY5SEh21
wPPl8zCgYzEmyw4+CFNLIB4HMz5GGcIiK+kvURpZ4f7XCnpPns/NNXW/rftD
T8RhbQfsP6H+4mlg8/upq6wJPmtl07TKJn33rUrCY8tX40Gu0RlAPzeZQM4V
GTGagQzTHcQ+HxoWD6sf//4zM+0Zo9OS9EBTV5hmr44J1LMSf6Ho3N0dihjK
0hhmFgaORTgDF7Cau6cpwQJiGVszY95EUHkjml3N+JwBce8XwbzTxq2J/hEg
/lxO8q8tgdxqVcg1AgX18Am0HtY+te+DOR0PiCBdkxNJHUo3krdsD2G6vp2X
myo/p9flUY/21XLeNUFgOrdxAudYktDYD6hHQmh0Pf5Eknf73sh2nBmJc7Yu
hNPIs3X4/pW81NbmKHV6mZQaWiNbRYXRJFaVULp0RWj8yA0vzOUsL/yknp+u
e/yWUQczOkLYarPUYPqKu+A0ApzHsqLP2pR3joBFHVHJE14/qL0oALBJcbHg
xIyfsgpcnajLWu2ZxEe59Wp6MsXyMxaqevzkz4IggJ/W/LAg7Jpry0Vflcxf
1rPQbUe83GIB+y6OIY/AYIujtm95ifDc2jtJypEgzZ8en2HzPf/cIwGrKtWv
fS30qrosK8B3Yqcolhkf84GeOJTNTZbL/qZpy35XDc7pJzAz+Bv/jnx06bD9
RU/XDR+8XqteavGPZ+Yr56dHRkK2Co+XPsq87AvDmw9QCBeMtaNmlPD9eskX
ZdIalNSRd6en6nDbnTtPLwqpaqK93pLEelbKoZ5wCb4D1ATyO1g91hqvkyEC
dQwoYp4sWnIhOh6mOpjzCC8cgKg6MdRqflmUxqMdVuVrU8vXHR+lltHPpGhM
4uclyG+BMfu7uGCc66sTuelyZPkRjEB6GuaeCXsUgVNdjHLSCiWF+70J2HTY
gh7l+yUtEPhzpUdSJSAiP49q8SdPb1L3ZV2is8yJcbTENq24N/6wqPfoHtus
EYrH+Ga0L47IhPEJvbc05mTGxdgMcE+nygrmkHwX5V7JZxd4yOxL5lvFFB9I
M18OpOLNfihYXoUfBRRWyd4iYUhGF2s0kIWLm9WvHEdTW9/fXW2pbxX5JTYJ
HovTk+IFVc3WGMQ055FOELV0DZQjRfMWCGtWnsI0Gm7KjR2t/4dBz8CRXa6A
WLcZ8d9CE66fdHIY+cfJetd+tLHLoQGh6X1RPrJSDO2zLROgwCPoRdaGHyDu
b+xsTEW4LyKw6gD+holqCqMK2bC5XZRkKooLPkrNSwP9tvwq0i8AMJkPVo/0
NYSvq4BiMCiP7tVNgfeNRDliBaMrz8UwjMg9M6ppxHGRzJDGbZgWBaoxBlvP
HtnN9D00s5V45XQvv8ZC1Lqoe/CsC5Be59Gvch1ukwXUH7zkGyac9xvvmme4
/b2+Qaxp6K/2IYLyV99fDbgGRFV7QsfcxG47o78VjRUzAEE1QLhe4LERctcI
f8TzZbM7ilZjpUpt6Vhf+GlYhVFGANK9Ye8bIaBfQKbli6hDrT3Vtn+7M2eJ
Mhf0eAXXTCYkaARqwmWt0Y1cSJeKI2qmopniQAeDw9ttP12laVHFJYyulPyH
NEM8Pwc5+TtGamN/2ohMEmHtKkHeUNuswZYkh5r8T71ieqK5EKmNloPQl2wZ
a4iCmxkrQcQndvKel5uvY8l7qmG6jhvIhpoIkMAwZOIibRJtLBtCPVzATaff
MlKHgAhiB4RrnrPJpQN2wYSZuBAGy7bS8fnOym7M5y8+npgoUk2zS0taMm8B
u6bvKLZQ0zK2OKOZDxfeigagZWvqy+sALcX9AyqsUiBUY1ejul8UDQCjaGft
p2b6H2e96Y6L4KSxRN8oAIyQMuKBynnkJLVg9NpZD6lXtOHLxKMRbteKGl21
WadkW7bpKEkB6Ht92g9VUmCwYDXu44Nnhhavou6ttsBEdEkHRjGeCT5qjxPu
BxAAbs/584+e6JgG2Bpb9yu9J7OMkQ0b6SozgvjtsHRSBOMsFJi4jUbHvp+k
71xkIjVJisPUk2kbMDkXs27ORprCfcX7gtSuLlpHgGLaBsYKc4JycB3E56D8
zhwIRKZ1XikO7ZyRgmP6MH4uXI7S6ge8co4SfTsjV+Cr3GwPmIGhhkY/p1Vs
cL2bYs2pmswC0ZOIrTL4EDidf2Mcbr/QoY0LMBOPLVGG25AjVfFhrMfTJKaR
peCezJCUxR3RRvTccpAuik9dHTArLVDTR6HpMHjNUn57W4+C8r28mtl1gLap
OvFNG+9ejdFkHmcJJGlOa7GBYIebuBNizkY/SWviCf7XOjnpT4nfdEDRNHfV
JjTV0vMhxsGuSYbfisEOUMYFKUJwUdH3QgKtvYM7QO8BTm/VrvebyiM1sUUe
T9vkqpwFdYs/1Z+pskVzFKDn5aKklalhhUaXKOf2GdLNQzx7Eti/P4+ooc2J
M+T9rltJFpuX9gJAsyeH9n2qlF6rwgrSIPkcnieATQO/KnZjFa8CFHIPY1Li
Oo0VXIgGa52mcY76T+KsUokVNqp+ueL34vtF+A/7AaN4oth6BUQZ46CTYxyw
xM6tGJmu2qQetuUYlmJD+/wwiiTD4No3NaueRERs7jvvDX0utOZ0a9q2n2Dm
gEW+7c1Bu2XR7NmZx7IjfWqmlawww2DZC1ZN80YKwH1lzhXDIohz6zuVO1xX
O0/fCs0KS4UnW9+PEUiseh0tRe7iEXO56fI3SeGE1oh7XxIyo6+lpRDGEIyC
xLIXDK1jtrrsDEnX5mrFgSGIeFWc0rlEJT8z/xaO8IOOpOl8AYU/UA3HJWWE
5u+J68F/Gp8dEliRniGjmgRWOh3DBeA9QblbhZZ4I1FLDfvDYZOwZigtj2+J
5TY6CUvPVddyv1ddaxTstQGFFnVSrB0n+r4jS7/sbLgyyYBk0xCgO8yCs9ld
d6edDbgItd03x4dB2svS86FiCAX7uCKRD/4ToVKbK57F+WEfy6P5l18pe1yA
Kt8oyL/V4iz4roOalUfitvj0DxKEoX3ymPi1USVYsyftfYHE9iiDpua33n7w
iJXiGj/FYgMiSDjtLXIHcDpbFxtXkVN0ARYAvkQDmjgTiFRkl1ZFScnC9wJW
+f1LLWOI1/nTmTsqDY/XAuRVzZGL/+5DQkama4kSyW+VFORAUzAZfGnUhVA/
OvS0HavXExqHm7iNxyebvoa0PQKBG5dwRkFJahI8KIcU/G5dPdQDpS2dxIAc
7xSog5HQ9uSh/vRQg5/qD7Z3RgnjZaMH40d4g9NzeMGibDD324hgGSb2qW1k
KcYNmacU/fDTEpG/uBKpb7fTbzq4MnwjIqh+9f4M4NAXGidatNuk0FNfKYFN
//beHvm6pBqevlK1laSyj52Vq31CQPAZ0fwXucXfjAHx0kTLPPqycCf/t2XF
MpI5KBfrJnj/KALTO9JG4QQDNbeuWWaxLgkkf3Noo6chd7x1VW7ktJ4fcBIq
6TtjFNv3BltnpTxRlVIjzUPPGyE81TURmidJl9YNGPjvFpyBvtgr/qD0qFDO
iZG8MJbyL0qzJh6INzWe29/iMGMknV7jjFfhs01gwx8uSEfKmpWj9wxHhd9V
zHr5KLK8ESphIa7bqCkZDrX/GgLEnkHVsOqGvQ/jnJwFZCTnCj7ab3rI8UCj
sv8DbuZHWxNQbaM4YvvCwnA2u23S1mh1QRCBmrFpPsCG9Xby9s23G5nv48PW
XcjOxAgL4ZZKCK/aktNjmqDb41aRD1tY+69FUwXc+4gDmCfeefiOYKYBAT2J
R3mxg8d8TnvSE+JLFo6sJ7gHH3A1CAnaowwhuDcBVFNoWNXoKMeNmNgd7qH+
jZcv1uQgEkhlyQnym4piV6KtlnurNONo4WetflEO/8pRJxGgzyITm/wf6fxD
Fnl1jAWW2NPOCox+GnyjI5S1GzGSqzQw28qDwfZ1W+KS7c/VGcryzkYB8aOT
bmLr3gZkQxxFRO0Vpa6T6qcbv/iDLywkARBBJVPbEVPuM8HrBjdsXJAFlsyy
DwDxBlyQcIXqKkQJW2409GJcg/gxRWvmqXPtydj8iiB6D757zMq3BUOKtUDV
tALkq9YR8/NSQhn0wCxfPnmjjji+FF6Bllz/Iljmq5x7WmnkORZ1rwchD/ni
BK/pvaDmjNNOJm8IBlwKeGO4DjxMzaFx94KLVubsVj8nQYSQb+ZBEWDuwrlx
6mfRAtV5ZVz3mVVUf8ASaaCkQflSPmyZfvZUdGZRoS6Cb/TmDA1JPbR1jNZX
RqgXLXEh3Z9ym+oE4D/94GSaDmxDuMICuySmtDD40NxoUBuTz3Y4CFBY8ESZ
gp9PbgDnppWZXJVkMgb8I/QiJr9MogejLbaveYhI5jshZWpWB2jkxBs94j7D
OQN+SE0USpcD1Nt+SPgEkeOwS0dFtO9X+Mj51+EpFTNwVq60HbnPc9Pt7Gj2
mJPtY/86SVeu4COyfhBvZ5XMCVE/1178jpxuWNJ580mz5dkVBo1xO3FQNo4F
OzC+hrbGwa8p6anDwLWpUr5fK+kg08aIuZ8lzyXMN53r0ElkeEY2DlxAg0Y9
X6+Kc4ANj2uGezeNt9nZGEit5WYr51MzVFb9AFm/g4jceZkwK1OkHDa6Kyp3
Yr7DHZ/lmFLB+2vmGk/2DH81CPL1xgz9PqaGqZSow546Rbxp+hB30AyHrDvP
Oh8LBawI3SbJNwD4+5IZtsRm4X0gJ8Kr3x8zvk4f3IP/VGmd7Jx7qWQr0/i1
cKm0QPnuHuY/1lHu7V3xSu1pUhkgNonfF8DzBuOtvF6EKypKbFRCK8WNCuNi
qb+d8k7IJdw8jnruZ9fNc7vohaBvmEu3EItd/EwfkkAFWyEBUN0YcM6YiK/5
UzOExJQywgkzAffqYey2dLM868JbR7WlYz+fEWgA7+v9X+nWVMwW/hqOjqTU
L5v/9hp508FefGC3B3PfOEwpKM0B7fixKDUiu5nb1KrrANbsuiF2Wyrys/iR
RPrnfwtCG/FVlTcIV/qYsCa64aicp1IYDR3igHbiu2L9haj8QTj/TKXBCDoQ
2Hn8FlyAKiRoGr+CsqgeQ32c5BN7tFTbdMwsjXHWahFbEPnwKBCQt8fWZ3HD
hhUlMG0fIiomxqZMIaqYvkSST+B0e2y6yYz/6lRZmOOE7GQ75pruJqd1JB3s
4fdwOYJmOwYwVbPZrrtc+3OL9TJ8ZxKj6tAAgppWjbt6d8pxmldH8z4k7DAK
Uik2Z4qwOv2Tfo5bX3NNsVg7G3K4PZLPTnWba3phpXxKWumIoY84fol1VXga
JDK2uIM7c8Qh4xAIj03t/jMc09eo9yYNsvAOX0jhwbjpP+vL5YB//CNGV5+B
vaZCrzMogsPAfCjM8O9Y1p59apLvYOhjpcL4UxLqT2Gt9ogLvso02dRGEbs2
3i/klN7gyAY7BtopIn9JY2XkJITZageCROIF+oRRSil+9YX2GbpLGawP+/Ub
1E9ALLx9w4r2AvdFDBMgNqyENB+eNIERR0Z6JayH5m66aE1s36Z81uaMJLdS
s5htMgvl5Q5gILZrFiQt5uz7y/Ch82Pk67ijGpucuZAReLZYlf7RpWb5czhv
7lqTv3eeR2TaR3H+tx3qWvOyYkvFkVeAbfLggl5btqxgffRJwQ8Gcrewp5Eg
U7QXIT4PnLDKDUEFKoD8LTvnJJl6kE9/BAy/YbRf7YXd/r6av6gYtNt321h+
feDFhqYyC0DlbHfscvB1GHvZkFmF0IIwPtdqjuq/iLo7gjV52iEtuSNRuMKM
c9S0qZ4Ib3zhRO74Bc9vJtUFhYncOPNsz+9A3x0SlwO3T+kqc+TCiRrzb+wD
caRChb+ZO5GbgFd1k3h0tl9OhT619hrx/DRWcZFU4OZcZDNlfdK1KNEHgroV
+yZgmBB9TFFFin3rCUkihcA6LRmcZMENqXLJeGeq6shCr4n1ewDjPaqhllkX
Ax/uAoDthzDFsm0w2wf6WHoOcjOd6Km1+LH6Tbc+/b2NkYDgbzDy/xQQ2BI6
x87xDLv/c4e8F05q0UiYnhiJdtfIt3NNv8n4nOoDIkrIAnxWkFtMwENmX/iM
dmmrq8hU0/m0s/SR2c8pp22M7uRzFdDCWVtejcVhgRHQ/ljJVh9jTzkKc8db
0k7FF+Bkh44Taz/+/fuL75/q2aG8hZRVc2oqsxI6tQIzp0DWiOaU9P8rd3QO
pwVGsyfpLCYWq1fVT7B2BFbOqqA7SdtqSuyNjkR9K4fmOho5cB9Ubj4joC9c
peNDR7/iubujM3F+FPAxsovbkpbXgYYsl/ME2WN4Bo6bDTCVlDZDQ6O5Y4I5
U7+taEYyGvzJAr/kNA4BvFn6AFRNA0pwBFm9XmgEoUD2KAWmA0U0JV9l05Bl
Hjl1haVF8RmxLAw5s2JrZWdzkD1hQQTOenf3sZURLSpu73pVNY3v0us3BDMh
otjA12DSGj0/m5SWbn8jWA9fmszQ/vNq/ecbY+htsXWX8bWbJJZYAAHxa6pJ
vQM3bPvdEjf7JXsGSVWg6ejPCl/VuiAuKA4Gyt7xsg6d6/vY532Rhcc6e6qq
7Id4+uF0whaz+Imu6kaUM8u901XAbf5eJzQSe9n1Lo3inhaPuyqYkZLWdo0u
bNjysdPq/TF4wI1rCRYQg9D1hLq3/OCWntLbFexKNTvaXtwKtOaCN00tUTjI
2KAGwjnkA+tDT9q3foNH1bQV5qph5LNQwDTbD5d9KV9boL5raEsFemJAQjA0
XFTtaHlTRYvNOBSey+C1kf0A19dtxIbZaR2xgT+xi2uvgYJhpT/laCq4dMy1
x4KHUkrPcW8gTUsK5peSeejoVwhbKPi/bTfT8AmlionLc3JaU9Wu/mQJSk2n
qdESXbwPbMw6Ao2AOVn2P/fv7TxHtluFaA2BUTTa0goEcBTYHIDsYLNsg6dd
tYYGcRbsW0QPHy6qeS2B+W/XnP//V32oaylJzv+ZP6Mjf41VfslUxIpGgIvj
1Jp8M6plHRVEiFQMj7oknAm+/dLY6ySDJfMVx+znl3oLLDVCQ8hUK9HdmEsp
KMm7cUCE064pZbNi5ZUc8a3AlT+uundVptkTSPZFgAOQFGMpqRsTlhHCbI9I
XvR3fjIqeIbfkmXum80/Tq9PV5rsWkEALJEhCKuJQ9r1/xMhyapSyvRd4KkB
ZQxEz99tFHN6j4Pgtk6TJ8EyUqiZTJ1MBg491uvpo4Ig+fWlCN7owv3SyMhZ
8wfTxKoP2P25fJzN8EtMidZMQqXIk9jcHktnbC0GzUZEuiVbKbf2lt+G8mwL
I+Tk2yxSHA+vIpGG8MIOfXbJrMTSIOBq1aogOZyBD9YXGE6hnod5/Hn0toj8
oS8/874USgrkVa5Bq2DJ4IgBrRmIYqZtu/yWjZ5H36is7iuEdHLb+1as3Mto
+TJcMo/Ts9t/jG0GnJcZmBv8ZrP4mWdPdsNRpenE2WMhWZkAAFD56huXfH7O
2Lr3t9D4laBWMqb8El+IJBVFiC+NX3RZBEtlA6i/GUqufc9BWguql/zfD8FY
fKBHJFahaOi9wizm1BpPJ8cRk/71oqHF422sjI4fhqvPq388PsygUnW3A2Tv
ljRtihBYFe2XdqG5kWiSve9HBm5TqUJ1pyFPa130/rh8kPYhYIpXi9aGYPXB
zQtwF5ztxm/BJiN5b+hRXE+BTLvQIA74d+AtQ1uOyjWOo0rsYEo+HqG6Mj1/
6t37chOl72XEWMUyDh5gbn8wVBV+7rrvvI8J+rKPc9IsBhVE3gKLQ7dZlBa4
ZkuCnGcSeoxbviqpLuWUUURAcDO1XDkfiDAFHgWkrdRtlSiBz+WmynBseMW3
NeC1ixrxtXyU/jmRNe0e84crdBeYezxh+6gzQQ2CXbfxroTJOMLvVSxNhRDS
Ih/WI+OoqE0AoDjbNjkLXA2ba/wABJsyqqM3Dv856ihSl/bRCRsCOlTf1xHd
r7bP/opbl9u87jKSQGfr5xNd5GHE5h1sEdg2xTkqxJIBu1JjYpz4BOy5A5aA
SlNzMHgbXh5uIDV3/CN9eni602Z0E56W1uuYEW8CmdNBTn3K4/M6eIrpQJua
ciQ4IYdzOP0TDoM6mZsf00NITQDbHlp4iP2tGsZpx75jVe/JIakQ+BsUKZss
lggTgHBqlte+NKgs0yR5kwLtCscWY3U9Dq/iR0y2jzPU0jz+eZYsxDgsAKgb
Xzp4FAnVOW469k7KSJfrRSFynMNMc9KmExwv2/4tosEO4YXquJVKWgEP/77B
4AoI6cUm3ckDukqyxuT2RUbAyQwVaD4Kh1TIHKvQmTHY3K8V2lkbPF8XxqvR
TpAmZsuZC1778QUMF7HjCH44BrWqlQuX3gL3HVeHRrng1VbbdGfL/It0b60a
tn+Us3zGqFwumwG6x1h8EvKdcHx2NNl5xxHMyiyXqXZZzmoukD2+l1DDaa6Q
m60mafONn1/XRtnzknecoZSDSwCLRbgFIevVn/rWKkD/h6bBPj5iyJCXwbld
sr8nIBbdKiqPpVRCvAZI7dncxUa5q8DJ6e7mijyzHf/r2PfUqOTLeUXxn5WP
UITzPtdDyp+Okm6lC4zsjHuNa7VfhZr1c3xW5eqzJdolgP9woPz0pP5z+wa5
2XB7TStkLPYUvnxxsbJ2megYKgfVxca60mnnwTXkuslrJd6h0JHNzSZTDRws
e7xv7NctF+RoQE8zpxDnI++rClR6CaURaRoJntNXVl29yO5qXz7VPlikFiqM
+HYryMbktk9Au8CdHhaSN4VhXwaa64ZjmxxX+ltJoJU+e/e1sWAp8xqKdACU
PJqAIRCriQod6Y/wX/f1rUzzPu7QzBKmx684ANKYPfG46dXDytVtFm9YsJfG
DYbed5rHbNwM9DNYhujhKEtMjzBONGd2NNK1xtJtE9j78Yp12FKU6bNQzDaE
OTuL3t+QEjm1ImTP76MB/jlwXb0MDCBJyVJG6M5VWYWtERhpuxSmw6m/WNJJ
FjmbCRiQ2dx+V/4+iuvQwmLZggxpMPNhPg8fQXv030+YiwkX/d9jqgZaGNaz
HF+Xv2VPyLzvm15C839/afKCH/Y1XHMxg2Apd+yWJKVyqaxjRfwkOinFm9Ju
18IWLkraDTVVZ4VrULf5kuXA/Z1DIzyoebxaPiYVLuFhgO3gOSPsFvho5IUn
Z2SzcHBGo/ON5AaLQTU2KT3ZifNRi3UXJAC8s/2Dj0QiiqBXRKgJGaEgjz9k
hQr72ZLsFWrHSCMwrUUShbptsCLdG+5NWCHJQ8VfBhfZUSjY2KRlccJ0Xwx8
H6BaS6DuCJcQu7Yof6x5/kj4zfDEYH66W8CbI0yFNuEySVoIe1WJPlgIy8Pb
moW+V9TDcfPsEFLVExV4V598vvg0uo3yCKzux1bGO6xKpDsuMAKPZx1Dc7Up
0ZzDd56DnVgudbmpVyTrAe1wq29iI9u1DN9X6P0QR03R8gftC86tsDNreZzD
ZuiOst0bm70Fco5/hu7nHfdrAmpJ9iNWxV1Bt+vYUWzKXv5MOyg9aVqGgqAr
UNSzkLHyHxcF/bcjdjzlx1Wn7ZMFojiPRU7shB/h+fFcUpsabFacsGXe8mKA
/dq9oEz72TX9TESjkWCrdVC7+9REcYTBxg1ehfTtwx8uG0LpKfmgkHbCwnE+
rpxqr6Dv70EKPzh0FgYcyYXSnAWKjFhJ3iBNk4Ok+d6u0mnqTtZfcsH99jSP
XGzwosVi3zsNBDjz74pAi2OyCs0ayUeyJC7l+pCNIeo0v6Auzpp8GY5E6g87
R3HhkG0JMwth2JoDJhhel9rrHcNDcfRLnIoNKO1lWE8/GYheVRzvbpDatA3N
PpWiWvHzOOmYZm6ZcXtb/GjWyc3QemJoAvz2sgcau1ZlygypgDtUFmzCiTrM
RL6afqI4sGdo2ongVV2pXftmm9hI8uuoqjAn7bunj0R4Ti1mYt6tO3f7Peks
OhQ/+UOJ/iZzWm+pFbSpli/hIKw1aN3nTiPjaxgtg7AeWUJiMOYQrnChFrrd
sXrhVmsgBP41PX5GaeDKojHpd9kB92Dbw42keNSB22fZpKpPw8esP/2j6kUp
Y7Qa5ZdyqgxIY6NWR8sBTgqfrCUGuxvm0iEW6G68HHC7Vc9+PeUVggAK6jfh
80sddoc2iYvsHhpuUalr6y6cVd6dT4BUtyBOGIvL2QGKomf08a84p0sgKDTW
61jzVQRTHPq+Y4SdBqMHSvsKb3l4cUwBH3XnrvoSb4ShRHhmTBG9YwekzMjD
vK6CqmoRksv0m7FaCd4fsYs8UjtHqUvOIMqFUZrDajc0G5NOL51p9VSSV4PE
DJAadxs2dV4C8wh/T2Pvye1wBXCoj8XGGbNSrMEznU46mvXvu3VA9LOW5SlP
REB2gVpLBOpyxSfIl820NmD+pY8F2SEsfubSZG/O7+ZNQnU267tz3a0BbSlP
sXneJONRhwCyNuiBfNnTu527685CWxfaVCLdKiv4yrSzrXd7K17vEOecP2X5
ncu6M2alD32VLmwcTb1p4+KIP06v6gGZi/g2doeFQHF4ztWyxVqjh4TxqHzK
SnYQ4AJSvFy3rtkNGyLZfxfoXBG8kskdq9xZ1k5c4iD2TJ3AAaNAeAfzDdg9
mHnpR+R3l/tejJjl3jgqor14mBKrWDCFS7GuWZicwPJb7Rsa+jBHj8AGhx63
lCcxsUdu90fLACX2Ea9mRjL6+cz2R9xUB/67MJzdamP2vK7VCkVdrZ4eVkLQ
ese6FMgyI0XLvjLKxKvbU7b8E3eR9BmQAeNK0Pk28embBajhyw1bI8zsziaH
y/9sW9q3GfyiVIO1/JfBsV75EkWdS3mjH46NndJ7dkY2cwCUCmrYqnYYYuOe
50oxcRzl2Hiia3Rb7imPHQST293u2++FTbQnZ1KIEu+MiIgnJM39bc+zUOB/
c1Bfd7pV41HrZ8c9x6eI/kkT6wMRFET+NxrT4cCbhqcT9UBfMFYp5KLyf+OR
koGOwOVaVrruzTaFQimDZgTgAXwrXHGMUzTQFnL9yMd685jOe+CA8gtEYrC3
w3sjitdN06+/j2xzqSvLolHq3bSSvP8VP9PefyQli1zKyLfpIgHfIn8N+hfa
7XU2sINeLqCgzw9BhNmcpl4Ug4DwfS9cyUG5ytMgK9z44uKtfFL7FUhEyB0q
9nD32IZ+uBIxl4XQ6xb0zbzQi5jEaZODi+Qj/kwsInPvxRKo3xLti26VEFfT
rrXSiaRDsoGF3NtiVnkjqpR4Vqcd4/V9pPDKwZRFIG3O5qsh6VVlswYpaU2N
jK9Ttl9x9m27+3EvoJOCASj3CIhakilMaTvyT8YsxQ1Tg/1GlDZxW2DKo0Bh
VXBo21ooTX1e3ceBdtAFvmzD2gPno/5KvH/WFc31xUSsTEM7YaPL2VgcPgaO
8p/hW4dga5lAb0GsfZ3ELEeH5tPkSHf44cqHDwgFe/Y+LoRpMvAd6BZr+Fms
uZcPiZzaQv3P5lZJkdqP/P/81MvO4SoAfjNE8ti5FwbXPzUIYy4u0ivP1Vt0
D48pwhgIoZT2f9ItFrlZRkweVIXUIvXZJCO4kgXy6mt18ijTLD55YYp+5OiH
Z1Th4Mm10PqflKttjQXt8VFml4DpuLbxcFeDJXKSp7qkmrsW/I36FlryO6b9
WDeyfsJLZV+vAHqxzMqyYpPbBAH8QBtApRQfO9zMhVMkVJba6e6WBQzyXDmw
L2oXxVbK7MTmcvFPPXufn3yxlr9Anj8HvX3GeUVKx+E+4lIvKIXVfCcSMy/G
wOiNaJZQmJiig5nkXQxMMO31NyAhPBHocDugTnDclhHZczVEVYgbYRHEyr6W
jNOl+hFK0snglsG7Imy7AV8jb5uv7X3OffZ29Kc5/QnVpW+oYzcS4NMYsCrF
E6Cvuf8o9hvPKttWtDSPIexPQYeIZ6KnvMd0iuNVlea9+Z9wj90z9/rlOLt5
nWpx5uRqtdPB20FWBZnixP6J7UlxfAGlAGizhuq37bRh/ihEaCf7QFb9mQG8
kLkpoElQxLK5+1u7QGUSVx11pXovGkh2JSziGyg9qbbR4t5BKRWJ7pjO+A4Z
p5HoQeTllZPIqFjU1+s3O4atN5nJIeiZ/715EXPx9wkiBbhDxDuuHXzsL9TH
ZXIgcAs5Uof1rbW9lyM4xEJcm2sE4yE3EVeLE1OdYFGj1PoOBrVVo82aKWlv
BMdLJODWW33lY8Lqm4W8KiZntQNHWlvheu+8Oi0wNtMpki7XUNf31bIV2rbI
5WD2gg8bca/biU8pudnIB5kWFp/QZ03MPia7kFmkBCvqUIu4vYeoSVo3/0J0
p5+V1kycrsxNd522qJyVzbqQTW5SlL3mpr4rNornuZHg0WmZuCPGODvIfyxj
q7zLvx4DaOolX1hfy7JjJkwxFDh1p9jZZoCWuUD2oVy0NecOgQRhTVgIB/Hy
jdvtq3DFyUjLbhqjX2l5gepL6YQJlHKuji1xrBXR3reh3dK+2YVC+tCSyFHQ
91Ciqhib3FMwD788EnkgSIhMYGXv7uyi3+7I553lyYgjMz0u18bYfucazaK4
hs4HB/kLT6nL2puT/l8sxFEHySDfsQFvge0z2O+pjNhY7Rg+me5J8bx1IstY
4daTB7LmPDLoT2MfWOOHptg6BcBvSucGMW7HTU0PvzKOLr7BoQOAbItABgfk
1schRSnKw3HEuzfJw5bz7XzdSNEvQTKYhLg0JatcBxJOWR7IYB5HWZoJqWAs
X/T+aDvV1PEC3YPbP2jNR45CzMxMP3+HjKknx2qKc7JL97+Q+4upJMXjXPGm
hU5uBe8uTomGYmZT7KBMbkFyXqDZ2qBGjfBbyWXvbl3ESV6AW+RdviFZI1FJ
eo72B2uUktvQZqjxeN0u0W4myRGirgYj1OXn9pNBlVwVLBSbGkm2DemEsoXd
byURYlHxJSxMNIRFn5y5b74x3jsTliLw6jzJlUgs5P8qyvmOa8bSCxRaHDBP
XbCKDr2lTrvgTBsDo7/3ttXFTJniZGijI8HLZlXxVizsHtBuB/LzKikmRKVi
xXVkYnwE8Uzrnz1Qrm0LdgGWoT0E5Mhfy4IKNTbQ/gnJHCpEKtVKmIhRvDqr
Nooi/MSaAUyfVBN3tocRyq5cOHAPvSMobS4y/ChZSoXm9PvjO/yvKZquDLrY
xnhA8kihyNKbxmfSU0m3jnOfLEaeJHy51ORcP3TvRv7wbu4V99nqI6RWoRXd
mhN7v2D40cAhhEss2GKiAJoMX9Rk0vy1kotNcL5BeeKajw4au0ejpE7vOlt0
xyfWIxK8UW/+2u655mehoHYgSMUO95bVH958RQrHdLI0gtwPF5CAG3V98ang
iAVtYSgtiOf/XkrCP0G4B8zUF32RfZpGIhK59BT5jIMcsZLyY5FvwCOjA+ex
3OaDKO9jVzV5a+ka+ATIFm+aXIu+iZhrEf7BGpcfWWHUfT/rXHcvaTK1nKeO
+8EMei3scNBRgZlQQ0WYgA3R4dD8ATdC+K/5hFmUZpmgZOgE15fSbbC5pHLV
BOp2SFaAnseA+O7t923v5raKTJQ5VXT74EsboizptWNCzWogq6Xycy6UXQYb
X/vHOJvzUJagI4tqTMqrnGPByMT/aMpqjjlEcxpg5Ds0/uiF1jJGpSONe0sT
XqiqsBcHJsmtijTtlE1Dim3yyyz7BvA8bXpvgu2hNogHWMCxmKP2ITI8kKE/
iZ36KRVyYWN5XnNkMlVTqk7V6uC+xRHL0E5wUaWTEbeTjht3jJKhG0/TMxGN
TnUS2gukB1WwG2Ngen7Mz9dZpG2kReeID374he/LOZXHMKBUMkgCHhWfL4qW
lcogzs6mpLUm/rhAkVY4rO3DZVUbBiq7wHF7Pwe46aues/0J3f+Jth4gBnjh
HJEWEvuw2OMTq7bt2iFAE5e5icc9hdgL0qsojWLCiePnhZdJP6cANAqggLIq
Jj91uQs+cyVVKUI3CJVqFronl6mQTEGryqlMKdCSYRHiwVjpyhvfMhBrfLOW
rhYYi+IksEgKdUYN4dnazSb1GOsxmPfEGuMJ9JdfmorIJ7X6058rBJUPgVNT
kTb8k+bt/D4NdRdBj1YQAjxvCQykg50uf++yu9s4zjFgtDa28oF+X2vyNjxx
Wx/UdKvkSta3HTTSOEgWugOeppTJ+9WLdZ8HP0qVQa61I5klpF+dCPUKvfVK
eggQ3E1I3Gw0SFE0VwzMBjggv15ttUJ1BN26S+4XCa2JVzn7yYJL3gaeDm0Y
ZZ/b3PtricUNBGKbASts4t8XkD7xSL9HeKVRBTrI2FnvmEsOTSGQH7b++D9T
oZnfHFdzCENBFUF17y8w3trehlZ6q2T+n2CFTmS0OjCpIkS6Nr76/3JfjSi7
O6vayhNZjacXf+dLJ74Mp46LrB/z+dAkHR9A+wMjaa4xp7f9SakS5SdcHt0g
8eWiiAe1ymKvysVA2LTotv0/gI+XjseUIfcVK7XyBq+LoWGds13wBp7sh/xY
XduTHfLR1mqYQmv1ymhQdwuP6pnr4nngTE19T6LGw1e/0F1HFAFqQvMKYz4S
0xh+2VOGDhIgluHYunMmPs4MCIRHsJdn6b7Z48Nen7ak46cODCv0J8ekxeDc
F/P4Cufru/XaHp9s5Ses5nZRr28wTa+j91vQkhnRi3MFlNgFHXTlIZtStsIv
9Rieg1w1NONEDRCbv8MRKGQHj5yCcUxC9fDUseNpOnwES7rwEzwF7XrrAb0b
qfX9CyzxOCJpVcmqS1tTUGUyGZZ4mvCYMFm32X0Y2obhP5D4wymPmRk5C9Hq
LZwvUI4rt7nMhbHtpp8GqDY+e5k2jO3xxJBnFjtciDa+eJrTZk2it0Ags6Fx
VL4VDVD28vqgeN1BtKB5zOlds1mzmtqMqLIcwhd4Fp2SgnKwpE4qCc/3J2SU
VIxgv8CQ4VNXhU5OqGXhaqdVMpapxJ8YI9XHhqAzrV8g7Av9e8dqYEHJK+Ve
DdhzXKL2lbyr2ukqcdJ5iqw60DaJuIxgwdamDc5Z/EZ71dokMfFEn4Y1YO4B
QXy2Mqk9xF79BD6eoK9UrqbBA9cMYkMchh/Yr5bVGf4SIqTZZOV1c6cyjhrQ
WxjWSAavSnE67SDJg/PE4YeavBHw+nPmjwjyYtfgKwlbbT0xsf8ZK8SGyXAT
XmDQJGTZexFZlavMZ175v6zlVNWG08OEm8gJnhiOB237RZYZ2YS7oQMRFHHr
WIhEctwYQ0qdhEmaHIy+LwX9HuU0Ci4KJSTotqk8j9z2fA7joIHydC2keesS
38CP2EWxjdGfKQARqZjAmzrkxz2Fk/SSIGA1fpAYJwSVJPPHhP/iA0xgHt7u
rYi4WbwczC8jWjxfhIqV5pXTWLrBUyrOJhULEgYjHY5CkVDcTX2/sZIEM9Gv
tc0IPcXI6RWAmn+Vss6IMjZfPeH+8kFfyrnjqcGZxhWryhmGUSy0BfD2GYGu
7QSoVMmOJJGygbyF1hoehcQTROwuCz15jZy/Jz/4w8n+SMjbNmBvNealQmrd
A5RK5H2biQYzggWnyFNcPzBfckga8EIlqDMD55IMIxflFbA8nF1Wh2qamciU
mCGpxbkKMqWezAIqU9hpoYziz5yA3Y6/xx7IgUKnv6mhFQBsCp6JWRIxFMyc
7t9Xs8RPSN/vMpu2+Ho7w83kufH+oT93f5tDp3glsN9Yllftx5tAtqNYrI25
/bl8MTENisf3F1vK26ikTBUoE1qDPKaBjryUUhuRQroege9l0AmIxBdcsuGw
FK6X/dO2b+L3HiC1fxON/uug8cdsLeyqR2O71hS3ltAm5MHBrXJE+eR5Tq3M
vxF8vrEkgEOq8Qfo4+O6nlhApdNrx1PS3MSCNwyLNxNQA7wGx5nfkwiEYfHw
5nnowIuFTRoEtU54qmbX2GgiZ8j9NrCdLlVJ0bB6Z+0tsE0pft8SNjA/77vV
6GbtYyLVODLl8m0kGnUTcl8OB9smErFgLMjrIF2OKem7f1dlnBotisIMj/V+
NtKVxsy6++Ru1NEuACh/13R+Ev2JMi/ddACOIVgK3LRHZqVGgUv6GVL749KC
o+nHEO9aCBwAMPVxXa1QkKqNc47MxbJJlWbDsSJKsKJZfj1cqOWlytynFmoC
XKwMguOkUeHebV/uFv3PqEeB7xyv3HL0hmlPW+p4cwaaBuU9QD+sVv74zTgP
dnbwPvMqtM2wt6TKcyYcX4I4zrY2HfQNQTZbTsF8Z05IxEd/HWJlPOQ72/XJ
wOsUGiNg3NcVwCbsnrka1e5RpLYgcLXilalo2NNIljUjjsAlUI/6R53Fkl7A
FS69FT645QwUnp99EAez05NaxPLmgPTawXSv1S2UIUfRxg8UjElSftrJ+U3h
anQZ/hQv9BoHbw+KIOQb1A73T/QhCnw9emAvm8aQ5Yb3MTNY9yN0/jY3QuYH
Sfd7cx1POjMd8xD+zNGhw7TUSGPG/7TqrG/5/UCynVhvnr/v8eA9P8vtbVCk
A7ifxRm1YPxPKNLOa+PjCIPHOd5ImCmXmI6I4tArGAexaEjXQ4Fh9HSW9NdX
TlhacbN7TJxjJfaCnbpwkgBHjQtKKceCSZijtW3V4azWCtgDGpwG6LbJxHUN
W15E4isL4TKaDQlVjHjwC/DYn4qRqJ2FZ2cR8M7zKR3E19mWlphVNiuL+hV7
Q9If5lF3QAFwcr2/Bc7xWYsuW+dzxJUbnU+CgqAxUbrU5Y02hOqGxNn27KNI
M3SUzPag2mP/HRPV252kjbjPKvWQ3jGRjT5nDQ1hJqnySMzx8o3DRTByDK1e
tOCWHlW0q4rV2HlJPeaPEeP0E8MYiqmp2jFVHaLIFCBbKGZ62vPW87FY90vs
+4nPry/DGHDeJ5RHZXa1L1oM27vyjIhwnBPfX8p6Hdj6adqBKu8nvQzy61eU
t6d6Kr0m0vfl8F3rAZQuvjYd8RFAdxYhcl0nqbu83H4sNBVifGy/eyNdiGVl
ICSlR+kb1bY7cW58Suac5TXJjLdoGlsBg11At2OCd9MKQvKB/ZqEF4vheKjf
M2zRLyWn7HTbWxy8fWxMRXVbTisS1E09CrCx/FMhxvoiCtemuyWKGX9U3FO8
TvibSHi14Tg/03po5TXOfIFPkaPJOL2bENaW8yQgA0JpTXEYLRAOZ00hRmtL
H9j/PG0rM9Es7T/pTBNwSNUbeeHAzENoqunVBPjs9nepgvn4OfWg9Q8EW9VX
+/YesbUda4m5f0+LJkiWLUbXDOP5iPNTf7zdvjD10cctNDifT5N6Mh2zMWeQ
dfvf0cafVIrhphIX1ggnZWXt9EU7QTOB1DmXT3gISJ72AK0ScJX1ZU2IZE9w
hMc8y6VNNBTmHDia9lobpJJ5zXk9MWLB6JqMOUel82h0fQFgVos3dT0ArhXq
XpYaggTa5XQ0qZpfko3fPSr//IocJ+GQJzXvoG3u905mTuBtUBM22u3DFU8W
URsFPJ4KzkJrLXZjn5wnakBoc+t+OXi7dZh3VVyk3JxZ2urSx3rBbaqrGZ3V
D5PpXFwken0q3w702OyRR4bTOqDaNd6jDx9VXRBQa/lx+lqY/afVyXLrGnyW
Euh/nounVDLj6xiut32UCiOH+kH5ASDGZ+AD2RRAJim9/1QULF5YhYgxSyqK
hivvABaR2fIDQEq3srqE8zPOMA3a6sdepA5u7/S5NPsL2HnWrXANzMBM32FU
w0zJH8YXGAH6uJ0idyWlwGjP8b9lqr8qMGk7ovHIEV1mI7lKmskXd8KPrPnc
/Dy7kO8lL968QRODLA/8fAWWQ3AnVMqei3NfG4F0PnTUqq+LaevUtbfimKsB
WUCb0LKi442pLBWQWGZf05NMwMG9qorf+JzoJJe/WAGdWnYQILiXQqjfYiSb
J//dAgGSXqgW54rciJ9jF4p52rLjv9cTpvaqWn4dyNlHX445mWOIpaqUE8v1
gSsiBzE/x72AiZiFUCMuUKjrzTSzIzDXYnT7GNtszc6DGm0qIzay3b7yg4l9
ZbwjYBGZwKCG6rueD6qx2MRqv02PvkT0IIs40afK+RMJa24KZaZ9AJ+7OYzl
h8UqB7pUK15yhFka9ZvMHbl7newXdipq3FpLSOLGSoMMSFtz6gFZNe9jsH76
mUSPJ6/lfhj2MztOd3BDbdJIK94ElgpuaQp/48oDzHrcNuAOf95m/B1tAfID
pd3i6R7Q/jpXkcnf9dA+LO9/YVmsn1TEC/ug7800g9hv0thVF6/HyUd3q9cM
D9lGsP4+gHud6lP9nSlHCQAgqVOZB1Gn/tqhCpOoPZpz9Oz9iWfUlVy/TzfO
02nzZgLZgR43lgXRYZyvQ1TgbVRqdy9ZWaBHDPIIMPhMrDlB9Z3dySuQ/zMI
m+5KsWRX7Pje2FwgdhICOPXTDVKmzk0mnLMDJUFAqNVaPfFf5iY7o/DXBiEi
P4itxYMy8+djn+rnzIWuFE67lRP0aMU70QXtyywarkkPVZ8r9XRKFYZuZz8s
NOARCADd9IJGNYzQ/epinx7CzanmfSLda3nMURbbc92ixZXWM8A84RqXuCDs
35HCxmH7+D3/yyqXgCKmKD1VIneavQvy3tZHBs14o+Kue6eKD7NUS39nUBP/
H1N8aNOzJcAaRDGRudV34NXptSh9EaONHObd+gZZ3HesODalVLV1tdHHmDJ8
Z4sbudocG2U4vSGn7dvWb8dmp7KpRwYHQPv+gU+blJ4PWO2bb3Ez2dj3aAin
cYhohw9gdB2gSc4zKBp+gWNbPwdw5/9jeg6ZmlqSOk7vyzD4djmV8VSgKNMD
d1zH+fzueGWqdhk0aPul9IpJ8TWwZRcAfbqqDsFljZlhY3BtGroBTKRS7liD
wBlkpv0g1HhuUAErp7QTRjs3whMcX5nNdw5x+Y4+eNDJUVj+2q5mZAunAbmy
wB4e4dklcoVWuCutJp3j/PcJDGpgGfAYsaj6NdjIWb2ffCaAtlSmyvxYWUxa
tJ0PJkoJZmB4cv0WNPQIFEUkyokXW+xR+2UrEf2fwkc8sHTrYajNXrwX98yg
OxWcxiC6dY9a3ktSuALeXZmwNDTiNSbyiTrpjJfaqvSeWt3Qah3WTBFC5pvo
yDCrtRh47gqaRMliB83zcJwsgZ1UFQl6NoU4nScCsONETTADV657MjoYMeAi
mXK8HFh62pKGQlQmHUIfRRIpCEeTzPQp4/7zr0ZodXtK4EBPrLFb5IHBYlsk
Medd3HaZ/xEvs2qwPvc1GM2pS2ET2TemMJLyJ+Jypg0Ki3wvher8h6YDqLoi
8d7Z1JxramzGDUv+xTXUsNnhOMoIdDPadUMQXOLYlK6zWyB9dX99/ai7qmUA
g8u0OWALiL7twXb7MNYC2jStbq7vewjZDgZoXwqnBDDpvIOWOfsDJePlZIly
pYa3knG5OkbeJI56vlv7yRVgzHWEJLdB0Dv/YIL9cNsxOgAc3x3zFcrY4Ar0
cEje8rpECodDSNKbvTvVWflFJCilFW+Zg2LUnEBMGFnDjodLASd/8gv+oNrp
E5NHMPxGyGuNAa8G18aHsk7RqF+Ic2O9KT2LQY6gBn3sNbdhwf4uOJcJZZkk
wfXW7383MGTByND6lqGWT12vKr/HCJmwOuBloxcRPQrZF+EgV4vCHgGg9W8l
sCwKQ/bEbqwYW/qcqJSqevIbVtSKmFWv8yeC+xkAAUfUg1fYIn2sG6211TN6
EFLiApWK68DFzKCicvogKSkc+BouEYKmDpMqi8370fwxnwmphWMoyr2NpqV0
JJIe8KizStwmUpMOwqDr2eSwLNYV3FIruKbtVhKT5LriUB5FxWD24BG6Lud4
OeCLQPHaUiADSYvs1PYrcHLgz+6WnmdxCJWBpoFf5LU85INELIvWOKriLaMz
zObbvibxfXwTGoEdUXOgoAUOZRKVvoAWwERFeNWnkvbHvJryAsyewAEISvxL
9wSQdFk9gDedCTXg71n+KuHoKJNWei2pqoxeNUZ5cA5ULI60sBBP9yypZ0ZH
qEr3UxHvjvZB5bWI3q336/onc2udfmuN+bBNCoBQibluGku9N58P1sbD6scY
mYh1tcdMdnSzRVzZO74q7aMfmexBO6pkhTJK40sAOfUjpGuDXauxHAjwwpyl
jDVS05ddsm2OF1lakBBcUv0PVOdOw6MdakazRCtgTT7LyeJ3+k3pJebCWXSL
hL38581tqtvql9Vu8MJzZINFWft/tMK6NQnp4nczPYrdcA7LCJlwoosGCxzT
c4AYwOsW3Kg+yTNLqG8lHf2+1na6HOdZA6Jmy0UG6XTjCY/zTPCtKNWQSDPP
/8RqFPvriuTM42lR6Awmig5h48leVJ88G9FdF9YVjEU1/GR5bakwkrEsdxYa
qxDqEHxPNIeAGzGOuRhG5oOLpkMt3ImEf0kT6PkjIN/QWtlXdXdQwhzaluLW
3ghq4oefcP+nuD1/hoi6r/XPzX86aKE1ChMnmi837ED2/JXoLqEKQAYWHX4e
xOu1ByNCPYFmr1aqUxzpJ2816IZX7I11B4Ojdum3Pv5aa7gZH0thmhQRgmGM
RdfLTuRx16j5m19YX7DDIOzS/74bWzPf6v5Jkix7tawCWfaLVHhkeaDmeCD7
Jfod4E48tNw0qEn9qAgWZodTV1k/YlwfpOy/Oiyl1T6O9m/RpPIATjXbfkMo
X1ZWT3L+v+owmP3GRuVnGGSPqEfuQy02qlzowzGP1bAi4fJeJSfmHhAyG5u5
kU5RFQrCuwCvHjo4vGgaizsrzWtHWUr/yLTZPOI2Xd/400/DZRt89K3rH6zk
eGWhVcsDEfU40ddqinQkLEgXli4KQS1MaujUytfd5LF4mM97p3DJXGL7J4At
FAsk+A9XdhRItBMhpQY4K9NzP1WaGXcLVFXPPud5yclCLeSPWDplld3KaDE/
aF3K6fXu0Ws55cfAluQZyTLqeuq9qfJdRqQT95gzK6CH6/H2Qv1fGkKHUOuK
QQS9s+saySFSNiI5eQ1HTrdYl6hN1cMHiP0TLT21ZDC4XKNii94KiEnXiTVo
5wTTi4T9LBXfbe1kt7/4DG1maYOW03CQb8hQl0Kt95UWXm7Ay6G9Ptcg7AFb
k7Cuu3CdGyDOLKK7RrM3YolMK+H0fmH8zkIMG5x5gvsIrgeauvtOYFH9jzeu
zA7dmMkNMkqpEWsGIKdXoPvpTh/blWbuqio/VGRt0VF+9efrJfK8G53LXyZd
C5MIWfr/8hVLuinuYoqElfbML4c5z2j5luYm4g2XiQ70MvOdIurBBNdgiWiJ
KORjh2JllA7FkdUZ6781PWaGE7nk2C35dVLEJ3u7QBDSBWHN8OB3iEAa0b9l
B0ie6PQTcFxyAJaPwiAVAYdpVtkObdhuwUDyT5XZMmEacAIL42WWoUphVneJ
ArM81g80Selcg1HoocgI5E7TCLZ11W9cpi9hO/KD5s9AFVZyjREfWGvyBCF4
oXbQq9GDyohTXP6E04iIAuZwDF8inAu8ReA7VuDTmszIoo0IszAkc7VGc40R
4u6kDHzVBldQO0FdnWDV0Fvx2SEEaIlxr3So6xbxzHy7OoyO91DO1SXiEyTQ
pg2MZoce5WKaudFQEHwtjXUequq7PGrrh261ToOpyWUyuwiykGcyF1VGD9kF
0ar83NXtLN5sv+1fF6yVdp0rSj9cpSnxMzlnFrdxXrA+HCciC36yaqt66y6I
oUqtIf0246gSNH+HEypgo1Y+AJO41HYzKV9m8mdJWSc/b1FkZfdptf8yypsC
+Ukkat0HsbfFh+A4Xc3ksTy9gGqTvuL+e9QPfuDAubifZKE+0k2pmEnhGrTf
r9bfS2OIA6jx0rqcrWlvBwVwHnr/ActpFUyZGacsdUaXCBjc/cLxhi6mUvLr
5twZ5ArgpK7nCeT3uvzielYbLmYjZc2mhr7IuVkRREpnF2dWgx2elZZBza0v
O8dtBfLJWIFZN2gv7ZEeKU27BlPlWABt+F3n3GRM+aD4n872nuIdlvn4y4H1
8WE5VEycVqeHBZ9bq23p5AgURkjjEIXrRzrxZ9LBFVFnjJaa7OA0VCz3bqU/
7At/uxVYKQ3AgyqMEF9FVCpgnHTwNpWtLJAkqfSPkMKkpGinrhw0bzNlHdmx
5X132GeexFgT6/t4Lv3NgtpVatBxyyAxX31HXCgLeeBroGx7s3pZ6+fF2scu
ABdEzZCaX6hV99m3FFLrw4DzJ8ykfGWkirOaxKwcDeNA5x1iKdXxN64Hv5jZ
lckLjimGXu3SvRraGja7zCloW2z49oXvQor0rtUhZjBsBupqlsbdKLffcEHs
AgsRxXP1jS022/rWVQnxs1fkwDDCertdvcXQEVkX/cNqelYszVpGx+4J3heK
Ptz6OEtXR3/ufAjthYGTIYzESx7Kqso8xKtMGsIxsbeAEIfmWdJAJp1QDZm5
269ROCpGOcIf5hqKOMnf8Z6/DrItXLGIyJm1w9XhDfa+S/aGB4gJUB/PaJMd
3+cySuFtwEqJiqtcYiLg0AklCM9ti4t3WLjBPILUNrknadKwOlezUvo+Xfcu
hW/uKO0+Z4fttDmKwNQqyxlwTkcTO1YT0+e/Yute8dLFGwvXt+O1fAcFfm7B
mgm2VFQLP8dICe0sgegLS97DbPP1sbEuV8Iz/G3ZDDB6+V1/CfW5cXeSCt9k
RZO+YKEjoWYKwkYwObi+2JBuN9OCUMQJ+MGSkfM78SE0H+YhfTLs6Iv+CWUO
dj6SmnT0yfZ91hKEaPSjKDbzKnSD8T63d8WorqzhB3ULlFZNa9dJBZLCRST0
Nu4aqP3cSO6wbG3epPIXq2dSKlhsRPPIIT5fWmY8mKo7234tvhuxAbPWx/x/
+iFIBglO6ficvnefGUmdU92AFN+cxGl68KKjuaMxNS2qg2Neq8ODfQrBUUlB
JWhs1GDbqsiymRN+D5g40YCKppkn77Ixfr+dY64juff3lhMpA5n016uol8WH
pcKEyfhljcanIW9DcjWPM4HQ3r3f5mo3HVUG9qgbVwVU7yZ2hTEZfzLsUBdk
QDDNKBuUkokZq8BHRaOpYHXAgXoGJjmzlJGcvrTlxr03y6F55JpCMCV25+aS
NaKQGt69JdXYQxGmoqoknPolc7GJzBvmnU2zQ7rc1qICKCHk7q4exL5PU2fu
BH+G0S7edN/ieKmGO6OGxK7mz/Ywc9MAeL31hGsh6QVMYJg5mstnO3xGFi+/
4LgnngTaBj+LW8Ldq0G6e9ts/EGoTgOlfuNcjIoUSFMBBMhCW0aj+HaThI8M
r7GMkcAGYxef3jLiWymzNgeOoJMeTL+cOVTcttdBbPPq7rAfoYZ5LVVxprd1
QZxpYXA2uqtFFCQkgj3LhavfzCwMztZ8VwQ4vfXjaqCzQA2eJSX04EVTe3T0
sQy4xygcyW7OSpGNrKjFFqlJyhIg+xdo4Ve0TL0M5Zb9tNM5fgwXWeNwns5e
2iGYoDl9BFmWQu/9XkUNbePfo9M3q3IxGqlPvrVsmaedoLggV1rFQWpXOiYX
tlNqKKxtfBDy/qTHETixG/EbT2dXU/LXGEtZS39U2hhPVTox/Pa9Agm7BTWR
rF4Ff3BPVL0L+hbOO6QlzsXnpzzNBHY1ctjmUyd5mKTC7oNya1ACx1k5pPjd
SqT0yVGwforGozZWplIUvqRonWWhoHQ42zgXHf95zCX9j26IAnZ0VXrmxGwH
DpYRGdwrgVxhhrOQQYA7rvrguWK9/jMiaf1I/n0KKvAmRXVBzGmt8lFX/1zF
n8DxDxBx281xVwpRFm0c4a/XNDIWkb8YzxCoaQPquFdSzZJWbB4G9yBoKRg5
7UpRVO3z6LOKBBnaEkUUXoy2K/mkL0xhlXVExKZ8JTjKhJYe5gEjzAj3+xff
C180W0hdt1NF44PLcz6M3liqhHMJQnt01OyM79I6HBKF1KKoSWPatP4D/U/d
c3qc5rekrNjzFyL03bUKf6jOHoORX6pPq5Lt5tuLEnqmcQ7egUHClBbkQxg/
zLi3HvkVC6F2WCOc/wqsSsm1xmPUD9S1FRzhy6nM3Wc0BXWBlq/XeUDseioB
ubppiR82NxUC7eRaSy1PkWyx6riyoIZMt6zYDjVBL4FgIgXEoSulrelTSxjM
fiWruObtTpz/sT5peqFh+iQuMu7q5L3lyYitmBHevJuvDjNQ+nvbjXs9/eXQ
Sq+c/Ycy3w0HrgfzsC9c9SeRDzN+sbh1G6hnT6twPBDujd4iYyzIGISCxKQN
Pai0bzNXxCm0UxYS2KhuhngTheFaNaWw7ktPR0uIWLc31FMvqpwAj4Xc2cxv
9RiR2CbDXax4MsXVx/bNLOtpm0e+3jUYeSWonGtd/j448UhC2W9kMu8QCpjw
0wr3ldSw1YWCgKe+28dTqJ9g+6DSRmIfMZ5aX4NInKyFXvnPHQ0xAnmrpttz
yulxjymDYZMT+mCeSlGj0dVHMZiv9PzRApTiYHEJAFwQtbmlvB+sfjcGBFpC
4UhBoxyvr35weW1D6+hE1HMP0ThXkmgiLaEBGlhh0hAgcBXU83iLCoYtrOvk
aEtb4a72w8hVHT+C6xkQhb/PUNqo8IVSmXvd8lnO0U4kjYetu8RcuRiYNdXW
M3Km/dJBy2jDH0TMeeMdtdhFTiYBCR1k6bDcHGYgsqgaCJkSwE6EuRp/fis2
Y6q9VYTdZ8sBEhnw/rzATYm35V1JiCgBj0sZilxeoG/vGllLFePaWzYmUwOI
EpFi4CR6belc1hf1Im1RaPUIESaLVbNpyaDvKb5M6AY9iCQ2gWzDzo8aOpHd
u9VJecr0gJT4+xU9YEi0FiJHPNFoj+9i8ePQE972RQTRz3pgN9Kijwunx+Qd
31JIM4AdqQ+Vr72f4dQVUSc48hz5peSa7QeO3RdJrJIw5RveusENtyNzAshV
VBFEFbepf1vV/tfc+AlEykIVlISTbC9oigiEffZ7wJgujjIv/vTFmfOVXZXV
HyMe9d33oFfqetp1Pd/rjnI17xlGfknwgXEC24vaCh5ao1/dsSS/sC5DAzZv
hQIU3fNw2nr3kVJDkEk3+GSb2v0s/kCzwz3bYtNZutNTPy+UQ8/uIGzlBFwg
HiG1I4h0lFmUGKRrZZ5tC9wi0UGRypMgtyOKiLnk1YIUQxRnMmgUS2Q7Jzu+
n/2xweIlQ3EVURifYFFQvhsKhAgVEzuyzSNhzZA+lSNd4xc1jJjIRVeNIC4V
Rl13lMnUJIOjjxRtmo8n8PzV66EI/ox3Vk/sBRTLR/lO3IxB+qukb4csTlcU
6gN1zcJ0iICxkOcOYFZRuBwj2YRf7b7w4COlbBb/YOlqpEXCS6QVBMxpqFUO
jzPY5Mmy0reiqGwxKEQOEca9meEP/vQETZdzPAR8VSW/MyN8kJNFf1CGh6TE
zavVV8lucsjGVso/hhpuGhJBIzn7caTRnfI0s9vscCIBbfrvikyEuZbb4q59
f0mlpwERQWAkE3bqgLyoWGdrk9gcIqpTACkoimb4Pbvrq9m4lqLZ7S8Vu2bi
gFeWMZhUycv6JmpK8Hsru1e7VSuGwgmus3VcZ3MwfG1oG3F5lBxGSrigVaaE
7a1hHJ2zWbNc3sF7ArW0X0Pz6AtO492DCVjER9O7DaxhvvX/XYoy8rQ1NCYQ
XxsEjRcIhjNwYdW7CArZIW9a1rRvfVLCof54z3GhFh/i7a0cm1YiE0veFGqm
InHEY2V525CUFRUYgWwKx+XbYdCQsvXha2rk62cU9vuzXgkqxUOscC2vDnDv
9Z/jRTREnjpyC25rPBUyw9DVvltpN9BO6CrGt9lLSUR/HCT28dnqvLsXfdBE
608m9K74gh2XTzjc2WoZHlHbG6NwfHH36qVZnUChOhJ1LGe+f+mk2D3cTCRM
1QeCiyTK+tgYa3IJuO7b2OQ2tOGk98vdvUYk2hRlK7ktHYrnwsSAvF5kwvNJ
HT5mNrB1ptQ6RoFf5NwHFJ39AVr6yXvgLDCVoITEb0SuHSd/q/nXmzi8RonK
gTInFaDA9wWEwuH6KsTo7uk9f4+AzZZM+otGQQM/R+94TDxsxLnDI5IByKYL
4xMXlvlWYIMO8/aGUHXwVjLpEZWOcDZFrDHnOoO0jjyuQs+k45c1BnLYIAni
66ZiUy/3K7fi7RsLZoj9jFTy8CT/TyPA10zZOCUY/dgbX+wzOX9z6lT8pMi1
BwQtYxLM6iMn1y4gRMhYpn6WIhDZC6kY0eYglZG5QueZaxM89EljTuTrtSE7
7CN6B3e+EbvwmInSdnBQkcYZDM6sBrE6VoFts2i4t/ZEPseCsvwI+UaXmWaG
qFiv9DVrufQ2RoW/97K1tr79iFDv7JCOdw+oaHDTmE9pmG2lzXBtUpQ4yQLn
wfoj7Nmd5PKbVxY01wyxoxm0BJ0A2Nb1rTP/wOq/eSJ+qCHhP8nSkwrRfew1
UHwSsNtZjw2IcnrHKvwpZ79WmCSGQzQWKFCIRwMe5X5irhYvNkRdsUuufPvC
leGstsPWB8Od7Pfi1hwUHssQlZcAXcvlail4O5YV2/7XevTPAEFsCTW3MgN2
3izrFxwq16OeuO2FSrSbvVxvTtV1B8QUEi7gjZRbM2PZ8BwCnUp0fUSGk0uq
mnqKFQSpXPAMYBNQLg09Tu4gBMFxgc9DyE5RuDUhxATQj2jWzHTHS3HyinpC
JER8O97N11R6W0QAMRU86fuF0X4rc6yu/qNm/NdCPghYH9z/mPk4jgYITn+C
oRCQxZX3rdrbTMDabzx4M0dv5vDXdRrKNW5bvA76kEEpBY6ds4eRtbx4DAlH
Et+jibtSTnOz1RV2EmGczLbXAT8FssdEvrjp2xV+S1AfHtcO7TaaBa2f4WLM
EEpTuIAwMo3FWeSBuqIFW66dey+eZ907YXXoQvtj7sXmNRxr7yCCTiMu3Xvh
VieJ7FKcTvrvGbNJsibIp5RkDk/oSv69D4leO7NB0eK/Dlrpf1NgeJIBTnz1
kaCG0qIuT6ghAfWRh/OfBRDdhv2XJ1vEqiW12rXts8YDdvFc15Xt2/G6+9/e
jmFVmuEtj6y59QrlfBY1EFJ4K7LSSSdoqSv6Dv2D6G93MwNlUL9cCGiNqjGE
SWTzIe9vHYz42wil3SjrhxIkiTYrJBv5w7m12qmS5YNkkDgfLufgyFobeHQH
Bb1LHJFd4dpouXrsssyGfjMkb1FVGm8LAadyiIaftTMrY5UrWFsLmBpT15Nf
3z2LZYoVzckXQPwQ3WmJxR/CLVl9MC2RqY2c1hBZCK//P478q4P0drxb2wNh
hJOqr+1ZAGFOydNlt2N23xauuibHYHNDDlSze7dE9QV+r7/d3GBLA1qJJD3X
shXaJv9/wS1hhYqtE08cIqyKhY7vPLxOLeUyfNBY1CmaBibaygivD3sF6wdK
YgIXgTAxq/a+16ixF9ZqTDXrikDxX4ztfeemdaIJyFZGRFvrMxA/smmuPllJ
VIpFRfNFveRR0EjuINycwqJn16i2G8PU00q1IHTpfTMbOkvJ9F4Y9hIaz2/c
hc3XZc/Rl00XBL1DWQt82Upia5u4hvoeuo3k5TppM7QyqkHfMcXMRZGnqIYp
lWXTpVpU0srFrfKKIksFCIIcecQx8291OPt7Ucv6Qt+IPClCX9MsOWNWP6w/
EqGTns1dxeLIAhbSftcKmAKuG3y+FGI/lwbCq7+l0xnQY684GRwVIBLxndJu
fvefJD1RIvL0K2gNxU5se+MkTQgW69PL5vBeujglMKX3E3hfHP0XNhX97WBq
7LajKaDncGnkhXrO76/v1NtkAP8CBtayd/RuldAHWKZyEPqskBCHM0GZoYG8
RGOqtB2PX/3Zx52EdPpjiS/ynPPxlY01+ux3ThuBelJusHS1/HL7oqKwX7h3
2VF97bxDoliON8I66UpCD1Sxf7NjJWG4QrS+1CNJX1KlTPOjv54hzC0Qn9TZ
qMsiCdT4fTUnv3Zf4/avT1JbEyCU+zeuYIO3G1P0XwERI20GzVoXARXGq8hU
sYOnCAxiyIWNOBFA1iXzqNTVo4zJrpOZrS4ieyJoI3d7YkCbOv8ur4CbrXt6
o2pcme2fJ3OlWclfRJv0uw6M4GZiebzuXxk4MrBVSIxqk0Ze5Tqc+ONKGtls
CJDjGFGeR8MhvgJxNAL+X1pXvTvltBjE/qrorOls9ZAtdvakWkBiL2IdGu00
OpA5EdeVgA1VIm+xJlgkHLLnbuqroB2rq7cFk4O4u7pR8imqBna9rvMYJvw8
FjSHiRoBcc81e+w7RnNNK4lWIFtPK4md+Q9kGEWh43xnjgxfC//lWxQnDy/j
q1w+AZ7//bmlN1oV4K0PvtzDjYP19P6OReMG5HocW+uFiQ5Ihbeov9IZDJqP
UTtzFiX04KMvfZYOgk3ZhvMZmpGIpMfK5dhmCNbCwWiSmaU8Gp6Y1oMneEa7
8sb7VQ/xojU+qsMzKz6NLCR+6mGSoBTkKhUm3k/XiYcEMjuerBt/Sol+H3u/
N65YZpTXzrh/iM5lpAVEBiUkfHmOx3PhEe4fBZIAOeevM1hrTRe4vpPNkvjM
6nPmarAMgwUTgwQsq5UZOm7H0S0WdUMgg715eFwpWY2PRxE407OJY0xrFh1S
gySzotv1L5r4FZLJKXr3QBQcTwoOtmVEMXD3r9nyfaM4/TpcUqRpYNhtZbKr
Wgu1OfKyESc+PKPvf+NRL6hq/3A9eE024TwZpZIc3nn2Jc0pZTD7w49z57tA
siPgOjhK7y2ZAVYua4evLGPoa+0j08JbHKu8pERhJZ4bdY1McMx7LJB8PFCH
oNBn1E806BeDRW14vqWn+IUncPsGPfFVfGsVdDnpmiJkC9DJkWclba5bS/2Q
6JT2o3BcwjxDj/cyO2GdR/HuG+iBxwhlV+QMszyMJInuubyQVEJFOqlXQO+L
bZxFPfGAVjXE2YZRBL8Oem8GxBW0AbUQVs73LX0Z8I1RbAULT8w5l2sg1aAk
7IKGSCxEwGTJW7GOU7/4eYLaOHzXolemuZN1dg5VUnRn2m47bXpr4kcD2xub
kbGJx3jBfzalsMv14WI07rOFGDY2LirKgU8wajN4DND1HQU74tI2JhZqrOoF
99BSIzDZC6bN5jNEOfXaFu7q0vomfoZeQe7CgSTJ2Ri2o7RSTW5/Lhbl11Oj
3jbWxElTRoaWdsqh+xESj6YEi8K9G17O+4ZeCUi+zzBPOwTiSrSV9sATRA1a
JEWsjfw7kI1/VtIBMyClzi7M14c9kwAdF4DumXjsgzz4JIfmdQh3a7lp3MR1
CcJ1H/BGQZXJwQJ/a0mX21A+hQ5SdTANl4XvzTfsvqjbSkyODl42ctNeGg9J
/jq6grCSJNDkl01VYpW9zBDYf1k/GWcB203eAnuSHpByVITT45Qp5wqVwveU
IKmfjXhkMZ8CW8Dfw1s5sorMenHjoAhY4muyFMmkYytbzTw9YAYqcrfo09xS
fcSwsQtYjsV1Oxj99ALOcRkFYPCsP2pkfVWWKDX4pC5hP4iaCHlUyoOEmveZ
uit2/BgaxJPT6WSQdtrcDgZoZMBwuU3hfisTZyQn2HLDdMghCN64rznxreWS
3sQyCU289MKWtLbx7BuTz+jNxqORwRHwC2NSckUSLGVp7QaYp8+0u4zitO+F
dgwtPIq7KqkwAzYlfrPKQihgeUijkfOMA7rZXjpRULfPhPBQe1BmavtFOfKD
enwkcJM5NT23X8JZwRIACz//58sL+EWuw6zamgSklo1gn9yWYHEypXFrmRL7
d7AhoAQotlqaoH3AocX2d4pw18K1AaVUXxs82TU2fWANtg474TPuoVcB6SuD
pv0jq2o0qfT8hCodYN9nwwSQmIOLVSXFeyb4tN8BS/LqhIzvkMtijJJQLpT1
Z04DGAFiXeT5dtwzgr1aCagUYXcPRpvXtBY6WtW7t1yL1YjDI+OB/Gs+EhPf
4n5r/jR5XYJ0NJmRFPdvsLigCvgjVCUnA2EWoSq/gnMl9GrQbYfnH7/kO2PC
p2+blCT9vDbVO/j5bUJcwB64cTsT0KfKpC2XeT4Z29GUK5H9fNVVsHNGjpcR
Be9RH19NzsgV4P38bE+HBXrBzdIPPdHHnzMQn5TjogqiP8DeSM+quVWOgYU+
tcA985GnP/AfUt4ouObrPCr/9go2jpC0gXBYyN5/Yiq0lLQb6fMOgXkXndvg
cbwT3B3H6a0PBO96TLvm/rtXa47p1jVhZTa+tVq7hAcCsfdynj0g2f2/Tfb2
YfpUdrlPUdiEhJyGtUKa3qPfaL4g1fxvytbXb/dCM9Tdtu4QcRvcHTfwsS36
YRLZqYLRcEi2XIsmGLhq7GVFjvwBXd2wa/fnefjrrouFljkzlQ7rND3Dgov0
E46KmzsF2CEBHzryyG+OSjfVqV+XKSVsL7t3yplVqA09jDsAThqb2f0DW5Tn
LeCh2ICHeVFvFQxKIC5vfO/7021c0Tjiu/26QaB0T1FqO4Rmw4Z1RlTi6zZ/
FclXbDHgl+GwRbmZBaZeTXzx/AgEdCpFNhULYqO07fOCfBqAvhNwz8KxpfgZ
AgnP9PJirIC8PqJDFfp+mYRw3L0Qn2OIl+sVWCNwVcmdUxitVpOkyqCppB8/
isfDNZumvcnIZEERAumNhi08srNwsHzGmD+ksGPq8FYCDkogYHzSNDdZ/Hqd
V0VJAIQR1ghdJUJsdLYopVgOveyrOcAlLZDd1zYwr2YXqxvD9RHBTVjf5B8W
PoujQvKIWxhDRsAe3tC4AVa3XsLHD+9VuLKzhk4HZofOOmoL9rmVpfv1mvyt
o5m/XaOb6WN0aLNi2NniRWwD+Y35NlVJrBIGhvDL+GaazNI9qLfsFzizYKIL
qVr62U9eXLXFB3+T++ilBH6Hr44rStH0dK5o9qg4yH6DB7sWyPwfYD/fDLZO
M20ICcyyRoR6KH5TyjwRF/T9AwMCsBBdmp/MKA4Cxt20VLaqR9ZHTTNn7uZn
gQNIy22t8EOH3y42o/rFpxhN+w9bqegmfjQsbZQ8bEjBO3kvDqdH9up0ksEU
55Hgj/MAFVAZf8P43R98BJupisHhHDyb2F5ta9N2YJuGW3P2bQ8BB0ztjnBf
rafvkTM+a4r1aOhXNYd7Xs+mEKceZLFVbrv9Kt1Po0KBt85YKbxmJ4cg8BP2
UMxmL/tl7wex0Eb+/KkekRwbyY57pwu1QTQcPfntAfV46RoN7qFsh4kluTjX
HdoAHpsKvmeZcBWrBp8ubJFsH7bULqvhXj5HcAHbcLoFRzX3LOZpAtgwuZj5
RzIjkx2KI9aKyYQ9RC1nRXATQVoYermjtbZ1ZP2uGp4Uk4A6aVO9wfEzXPwt
bQivSRY6er/sNAj6fpqhDHWm/mB0zgy6FotAKv9CFpI9pW/9l/xNEWpD27Dr
4TeKHwAm7ZgujRNfZRfjGXlz72P4FJEd9jqdap7kStNhoiWQdyE9Bi/BUbNl
KboO9qZQKZGUaxa/u8Xb0Ek1I+VzdU5CE09hb873X82qsRDtkOdMKpXwsm0M
8IwzHtG1yUlR4NyIsmzpdOOhAfB6kdZHvztIRiBnpVEmLRalotDM0IukKqkQ
SrFKZxyLs8MUOBjjl8sEFccVXpG5H8EVmCCh2EsXwpz9JX2xhAIwqZxiC/TK
RT3NCgub8oEF+RO7482vum/dV7eB4juQBa4Nb2JisocDg56fvW4CE5p6kaHO
69zUf0jY+eH9Bslcs+ZPveJDryZ1bj6nlnIK0uB1Y0m5mTskk7r8yyteTRJ9
03DfE4ajupsW5giE9wSV0OPtEZPbKHz7AkGpf9ZC7OrEJft0NZb1F64TTFhZ
OXk7g5JBz7QopIbsOXCcRhZs+OH3mrdjHU4bK7DS30H1xj3ey0bA5gi2HdjR
TR2lluH7QxUoGeMQD+1gn2kA99tum/AUNUZ6hQessqPChoXx6xa0SFf25W/e
zhP8vrUxS18rG7YyYgqpq1uP/2d/AZZebZrgLQVjjXh1XzSkuAbudrcMKIvI
c8g6m9B7vvn9PS8BrwosBbs4E7Z6ufyZ65bgFmWT3k0plEu17TUWrx+UJEoA
8sJyq+xu7TpFTAodeodQsbO6z6wakBxZLCpj4glO2cO5t4FKZZO2aAYOVmEP
EKc91TB0kSUuV7A8Q7Pw6ba/mzuBNqLZh/RGW9hWRF4yAftITaY91xP2id69
+Ip/15wCde5w16UoXHVQfmXmJsd8xYZVFFPINXoJQjr0MZlo8affIewkbN1W
wIIUVqF6EC4xnHkYk+Tv9oJraqNIGvh3XTZVUUGuqZoxZcBzxnIc9ghpLfkN
s2HRBkP16gAA741gzVfIdz4rstpczvPSKeXevvOamwLVJt6biixEdsLeKB0v
rdDt1GGLP7VARC34KkVbxIG6b7UHPOAwLuhntbUplr9RKY+qm8Ukqk6i7GCW
TiquUw6vINgfVJ1rV3slkI4rv/gfl2CNo6rGZKK/zRqMFedQLSmUTtVkdQ9Y
OOAaj207I+aSjA7gmHaDYNEw82/i4j1vLFW2f6A1ZjJ4Vw3dKz13rFt6lQHz
wdX4udxCAmmT0ebmyXcP65nj9A40+bT315EGZP1MfoQV+VLSnNzOxv2rDFwl
F8ib2IkYZgaPgN/GKF7eONihRg4NbwZFwFlQwn+04p1zMpmBf7rcGoDUYohl
u5OxwE/DqSN6pbMqQzdyJ0APsdtQsyXdKWTmlKobIeZmz01GlrDqgJijtUtV
7I2FBGI2qEzl7skQn8ZCY0MqmCSQX2dMN+MR9cXW/xCFa3UE7t483129zPNT
ju4mlesOOcLEhFYCCnNVCgA9fDibwO3JKcmGOHGaUtxYNHN0YlEjPfXAhwpa
tk9YNHHnVO8xrgZC7oQ4E/wyiYKDWxCahOK2tp/oSFfTHTGiy+9BK0SYdJH/
2wnTNDkZY8vTvPZReFKM8ke9ppBW/r/Y3jbW0XRBHKbk1Oq4kxceV5DWoG+Y
1PSEBobPZng2AdkscHQcDzUbqkzUDMjjO5KSObgK9XzbmtLD6yc71JtbnLhm
1kFFOl7U1QWnBi0jiwGFUuKCqiq0bLW0ORRwRGcGUjhvvmXbudtB6s5EmaeB
XBIwK0gnMAmSiWzEi1tYkxPb2dDsTvc6CtzcaXe3Iw/1e2WCDCsRYvaDse39
sd529bdiifVssR+o1rM1uEUXY0z+ibMNJKAJdg2h8cVBaS9HCgFmC9GJAHuf
gjyFFdMQfYmtrBPfNXKpWw3liDPSrxRh3zAmY8MRoSZyxxL0WQ7cLmUqDdXb
vJm6Vhd2UYnVvVd53BYAtNXLhqJ5QmJN7BIg2EuUD3bpZZN6kECl46ZQoNUX
z3ZLxOEPWPaAGTZBM+D2DBszN1Lhg5hG+thqYAwwfwfF+ZkFSOoGgY6BcEMZ
vqP/UgJYtP9sCsu7ahCVZo1hyRibk8t1tKpNM9A7EQJ34W0B/g2TOLre9LIh
j46cLX2wCfdGLSFbxi4upVfDRyozqjS/fWCzseqQvC0DUJraPtmWEiP/MZ3Q
zXpmYt+pp6ndxesOlZczGUDNtICLvhJAYbOJiQilv7L65hajZjA8IjXARffE
zUaDL2fMMYscwAFgP6K8zemSannZuYTq92//IQDFqse4mgubiALnNTSsAxpg
b6810T9um9W29drLT37BLA4hxgyus/uVz6DuJ4NmSU+YuJTdEuKeEOlhtG64
5K4cHiRhtNj/Pymgm/9e8R9nv61jpo0d/y2Ah5Bo3xKdRJZiekX0yZjGaSSw
Z6M+ZMZtaeydKnqMHVBlj/U7kKYjgNUOp00taIjvPYqsSitVPRVhxzCIktsM
EBRzL6Wy3whKJNADefK+yUXRBLwKONi0tkw+TWM2olinpQxix4mt3DDGLBwV
V9wyOGb7CFYBDMMxdg6vJInSMkb8hCZYRneaZSkRjlXxsRFdsdZinex9XivB
UuIPlYR2uOfAn0/POXNHKtkC/61VVWOT2wn5U7Bz3kF63lKPCowpDYc7P3bZ
CywfCAimD+1jDxtb98uZANIE6OT8rpQXV2gQ+oo51BV3N60j06crfNxVz2Cy
Rn2qTiwbISm8v4QEWrQeXdnVjPlfvpGJVvCEJ7Aic4dR28YX0xoThAavgDsu
+Vzvp0aobE9qRgZFngDFU6e/gbJg87CVCuOXyESi1pd5CY2Jlrni4IIbMhCU
C+2zCCbwqGZbtLioqZ7Sah9EuS4PnsJMPS5+1ZbhUmvBULSZQP9JIjg9ursX
Wiw+YnsWPiIIPX/jJdClE5Fcxk/vKRfinOKghvHISX0b9lHTKPedtljo9Hqd
E2ezZ98BeOFtYXC3i5Bsn4CmO5Jue8EaNbsaCt9sFk4hEsJFu4qmnTG4rZf2
B1TVg/T37zn7DTwkE7KbbSSOZ8P/psZYUobzDXJBujUOcLcU5yAfFKZh/2nL
5+vu/QWcRzezIWqrjoYoTFkSkXb3G3rVWgnXou/gLti+O6V86+e/nfENYEpx
oE/4FPZY+UZZSxAW8JRPHKzXdqIfQMl0H9ZFYfW/L6huVFlnn0xoeNdyH/PY
Dqc1EV5OqZ7TtpvxIfmVZczGUyYGY04it+IUvUxXj0hkvCDtWXY3mnFIK5U6
41yUqnBss7khNQK7g/aNc5DZhEbMZalWGsuxtLYy0Uxk7oZyAfmKx+cdMBav
SYXblE2LSDOo9vwX/lJE81HTh5Rbw0qN5mDEPlZYDK7s0cqiUYnRkiodBpjc
2YE3RioamTbMoTiVeOHyFux6kvY705jgb+9LfPysRHQF5dlwW1y064q43cgC
Mr0Kq8OuHh5tcLnjaTxwR/bVvxcquah/2edvqKrD3/gkNzlWM0Plo+xgi8p+
z884AauUlnqPFg3wHAta+QZW2HbX73k2lAkX2tQ4Khun1fUEAhV5RHHkUwEe
EOEu6n/x9W5CdGuiEvnkpsjXoqk0eX/3sZ4vV1+gf8tl50WpPxWXz3/9wc7k
lGa6DzsVo+sGOFPbtPjUTZl6DUkuFplOtHRooAGNbEeT6s8qvVZrTPrTJJyt
KEe7v6DpYpn1UQTGK+fMRvjvpj1XOBw6vLzwYs5bQaPH/d4qNRAq8xYKuDs4
yWPAfvzAwfcYi2/tAe6Ao6plBIeZQ55upLE7iVE8olUW0S5ZpY0KePYSZiXR
OWWOX8QHQ4DPnQBlG9kd4Fn+sdqwFYFrB6qvOnN3yHxL4QkBTJ0Bpd8bW8z2
1mL2ANL4hSMF+3rqJz9Ot1ieK8Jw7hIAcy3InsTHafExbnbcCyXScSAAH05d
/Ywxkydjr74psSS/9Fwb7XOy5FY0lGU39R/a7dbkpUFquXPGGWp4WPiFKdP1
46ggzOvVEG8inq1h7w0xHP4doW8n6Rp38wsE/R1YJ3LJp7QfluiLTHkmVIaY
Vtzi61/LtKxdXYy+GhrtXEBkA+++SoZ+WVioypxWhLyIsigezh0IFASSjPeB
yja0hlemhl6LDR8LkjAK/CtmwxaijDMZPDTmSzM98+YVcjtQ3F2qB8vPicPN
YMmU0WLC56Wh06eTN7YBaeqQ0ILGjrcfSxC2vU/Q15dL3WPQjcMq6rmwUeKP
Tf0plMAPCz26e7hi1r2zovMZppqCWND6s6kp5DM/rQuJcmHjXRga3Nnm/wXg
2f4hrcHCuCHinc46qVufEf63Oou+XA59FW4SrCMYfuKXN0vfN87rTWXPaQdh
AkwFBUQS1OFBOsWJ6T5b9HKwHVF7XRSo/LmBOodY8U2dqZpeJsOvsw7PMOuO
pYiXrQEWW5cdSHuulKoXnw3Od2kFjb+vmVsDCMt5qGRmSUL0qRK6k36js8RL
yGr9HV4dpAaYjA2tNarZT+hcXT6xFAGTavMux78j3hVmh2PekTICozxM1HLF
wuTGtSnqBAug8TCYWKROys0MV6Zpu43mkOeSehp+PDbmz0eRMfryBVuxLyBw
YVITI5x4eUhHuTGCF6eBidsFqGX8YijFuSHflrNSrfzkui1UqI8OQymCUSKx
NHzPNgarwc3JOOc3IbBtZRTU4gAln9UFPRqeSqcheehJ1qZQFoCi5YeBUphT
9WtyL3h3fY87kF1gJCnVJLKMCpO8WglHFq6RMdyfogTjj1Rtp71sJ07Zb8TC
PCvWYyzz+gedDTSAFOPwMlFi9vfB/v/BpjwfRjni7PiyAOQG3CW/rkx1wQ/j
FRx9QfSEFpguG2xl0hESYObxMx0XFb8Y7u1RZF91iuDZVTW7LJplF+nPjz/7
LCY35pudFpbl1ft6BqRf7hCPEmP64WwerekiQiOpa8ePfGFOyfrkfVw5TCsa
WW2xR3gO0k0XCINxd27a3Vlu0KEbonKdIK2GwYe61jQg6Ha0IT5330bcGsol
fifptqC3U37P2KbVvmCwMLnJa278ijjiGbtGNxJrwn9+e6w+4zoROx7L9NOp
gXNJbjtn5q/FtWzyNURb6MYCdkNP85cf4FL4UPgvl6nNi4mxT5gnW2wgcVNu
69Yea1SRKWZZFGkdVb23qmsf9QzxMRoll2NEXJnL4bAntvzPAr52yDsVeeJK
WyrAwToPfKqQhnQRYwtHvva4NvF2RRmxBahGV5bNUoTL9+xMAbbbqtTvCb2A
SSaO/LhvNzgyuKz5lKmfrJ2x6c0DWabiPk1dT6mcbHPLxu6HYvpITo758HAI
dS2/AAcKWja5bt0D5AxYG00eZsAFFu7B6X6dyguKVSLfiuwuszA7+G2eA5bE
4XaU7meyv/4/CgN5b6duo6QXCsgsj/n58vMAzBW0fddZFG+ydluIzYSZUH7J
4IuUrIfb0g/fchjAnXoXptIdzz/kWtaGLRQDFwqFiKuHAKEJv49eDn+/qpW3
ImjnDPLal+0HZ6R1Ru327Bjf4nE68h1MEVfS2TviqIiKwXCFf9XfXQCmcWT/
/Qyg75oQXmJVk/RGzJaghSLx2FsNgA/2vHQMtb10YZAf3ueInIUVDTnydGHc
0WKyQ5DnKvQBEucC/pGw6B7GzDN8dlflIoO8CQqj+dN2ZjUpYdoX1EQvlTHA
GDo2SfZohWi6IO5qsCasl+V/7SdXVdi+KQTr5lfuBKcinzE/gTi8q5dJyd0A
K9LHPk5KQsWEechj3f473VBkIahF2p85eiHkEV7VbMIxdiwgGN1hBWTZ1WzF
iXiv/oigkgrfAuupvXh0J46tg+P9Gj0x6qMMZ4Vwd8feX5j+y3bl2J/TsX51
3j8FflSfEoD4tBfMKN8nEKvalD0GP+e1XXjpsR1oxOA74ppuIq0em4eLP+aL
Vz4lcGO4UcdPxHtEDinZEvNx6z4SAGsMzbBj9YE3YXT31aG2KUfQKTpPXaHX
YSwcy6Y/9ilHw8Yt3c/kCEQTlBgLCGEL7T5kJgHMc6jk20enCBpLVOJ4BkzI
sxGbifx4ca3cO++nedfkY5B6Zt+ZmrF3HBHGr0Hlipz9H/wiKmBk2kB9VcO9
TOkn/wIM7vxEEVtJGD8JPT9zsdrte1tyXMJPg0LBWVWAPzBI54AlE3lklu2p
L4Pld1Cm8mUYp8dDzfqoSyNZhM4+QYrgfNzQ8nxo2g1lX1h9CseNQM9i8LdW
R2MBBwTMkNGKli25FEX53693pfNb1iCFiEM4k17LlC6cpXW0deWj7G47Om/P
ABVpc/Kyd2AUf7Px6L2gQnaEpQ80JTfqw0JpEAxvs+QE0fxeb1DTKTpQ6lT7
ByBDF+mBDCHC1/VKTtfVLG4bCsgxYNVlzyq916Im5SiZ+CcHAwSmghpAOikP
QchVcOqlz961uFxhJ6/KR/8/vpTzbWFnjAcjIMQYYK3eXe/8tvUE5WS/lwwW
BdJg0KUHv827gqkNcHg4tyEzyRmFoWL49OUMEhGWY6b1P62kBZnK0VSE18lF
lsXwsX8NLzohJRcbNv7vsUHj7mwoIn/6UeoFUosMuPuZDn97XIBHBKIdTiju
xJuBTGVIyswWvAvI6QXMSawzjeKYaoidCLc3orO4c3o37SnPRIzU9v/Mu2aU
SYnkJphfNCXbXiyFQsfSiwVpRtzz7nkavoqw0X6LM9IBD6Fd1fl/lPi8cqum
KZDVYmzZLAfkF+SXyuS4iNBW6yEik1RfSBIFQ1+iy3aeYkJrWa5/AMh2bj3E
VNUE1fdyFu1fBuIdq0ZhqDm+ckd9QqKE/700+MJj0suVMzaqulErx27NS6RI
nvIhCYei077i+254B1h/bcct+urZR87iwqCLUsUH94QEaHpA8ye6boGgwSsY
RgrktAMZfb96qTN5ui/DfUZAvc0K+fNdvliKxGvRVmqO07u7wbWYNgqROT35
gO/A2DqRoLsDF7UUughcOHssME/C4EBxhph/kd7brX6U1odfAXSsmqQWs+Yf
r5SQUaFKC/64LluZf934SME8kBKZ+U7oiYK+Y/2Zq8JdXvnbkgx1zm/vDhrP
Oph847ab1EPchMiP8onEH9KwVbdMiLr+zOrNzWBGM4rmRSInFAS7UDotegCR
FVuH6r2w3C551eq7kMty3gGARcbEl47J1Lu57KuectxkRLauSiT8RWvdxgHX
GjRE7HT7dSkJZRBcuInHyKR5NDY7u4NZFmgJD/T10lLzpPvPZSA9V7r+iwEr
Rh8uoBOOIEaNW4ae/m8g3VIu0ioMl1tqRzO565dxim+koDrdUGCF4jyClB7T
Kh0PHL3rgwq9+h+ibzadJYTf2ua7O7shuZrAAH9MjyDwRDZR/YHktdpYG5nL
Q68kv7ksCuVwrA183YUl5aOtjl4pi3CGL8EN7bJ5kND9W3FzUpbjXpJtOzby
g5J5rghDlhgLsC91+jCIYl7ZVuDDky3d/bVKRlW4pAkDVCbEiIGQKGKZ5WTW
TN3Gp5yc5f6C+rIfZb70RvzhRGFxRSAkaNJ2aKTLUcilbEqeuEEf1+nGhrpw
Iz31Ow0kPcWQWq0YD9gK/2LTUg/CL5h8jnvlQra2n0vpDBzVMi0KVdUborYO
UEgop8v2zjNypbQ4iA5Rz1S2G/Rtw1g8tzd+PomplrVsCTMFS0ObSHHJ86zj
QRkFf1YaCzWw+jE/K76hovSd5invR+GGYcjbUHuv9UTjJKMAtBefpKJ4WPRc
IXqmGzxGuSUvrafJcJm3ccQZCfilYOzt+1T2Bl6f9NJ1kNzWO3lGsogp02sQ
LkWPg7xqORghxP2GkgtV3n882TmGZ45+tBSUSrYCaaOuIjtvGKMwn8iXaGqx
iqB/duMUQ1Lk4CSTVAMaEiRmewl5FYrIet55CVNP/0fXCscQznsEvCtTTnm7
8Zqf/XCiEzmJhQ3ZhKlZAujVTGmbQa968Ke17j2brES8tf4tTEsne3lQ0hXB
SaLtdWU3Vbbwuaet6FGIwdYqB+ciXyx8lZtyZ7gT2/n7GjpqM7fDp4wA+8Tl
nuaJsmRxYKxuoCp88iv6vt1gSAORoEPeQqhTC3wEgfejydeTapPnZd+ZcAKA
WyMunt4xp2/yq6ZFfo3rlEsfWBCeBmFP8JUUNukhcwn8n35n7b31GtUgQfqR
KWojdzfz6sewj0UBJdLqG9LsgSPb2gp8Zw3a2SHSHR5FcJt3XrfPjtCgY284
E8bjxaUJ6ywMoXNFcXcwtj3tbATQLZjcKf+3f9Y9PPwpyqkHh4Vo421xFfyz
ua2vHBgmU1w1DuFKGkDbw5esIZ/Rw/JqOHSuedn8JwLPbw15mdc05r3Gtds9
GEy9KJF7HSvI/qgcnRdwWr9lVOw1Dw7cuUASBxQKiWy0ANBk2inTHWbHzi1b
GUc29L0YrDOINrwW74kh00BXEFjvtKsydPyd4OyIQy7D2E3lCKg0zec6LRFv
M2BVM3tENurgB5AJpFmziWZALx9X61n93kcfUVC1gdja0GEOL2aL6krIFVqL
dTAz8dIhTtFqfzhwmU5S6ZK1s0lDxymIExOuAiXV4yT4PY9zcXiUokylv1m6
eUthLhugJKzv6z5vXH3hZgXrsHl0L1g8X+JphPbht4qheLDELt7b1BQu5Kla
uIwhtC220JvnjMFc3TWB9WwaakXU5Ne+slSwgSMvrW3SL5+Czrf7UjUFQvJX
BPyEIwz7j7v1Ap2F+wpR8GGpDI/H0ZnIKtdRMN5kAfUiMURgyCCIxrJTyJCB
FIwXdB5FkRk2SB/fPJxrHuPeqa5LwalzjMkuVtGZG5Ho/s4ZSGbzAXfIcmD6
9g4J4PPKdL2pt4HNyDH2dpRdPZDKNEDPg2j9tv+MiimxSr9ZQm94sKbAHvOt
mokFxh+aSkUAJPnpZFSVhZYRsWHVDh+sDNPDfP34xqLSO/+2LHLxyFhHZ6ml
603PawYxZjIrOVNd6J1hPW87m3BpRqXS5JhCJF+NlE/bkAdgodpVFg0ela3E
En6JLVQaX+iitAMqCJWe9S+dNbI2ftf8mWo9FVC3/iGziQt2YNjs6qkLE18/
6GmMcdJX7iLnoQ8C3F8zT/1SrERj0Bh+909TKTI2ZZUNNVOjBi2j2JqD8BDh
z+L2bTBWwmwxz2Hg1Qa4o8sYVWLvufAdJy6hJ6vxbsuZKKYXzIRRU28LC9wW
AVVOCJNawty4YJVfl3o+L5fDu2cyfnu4/q5TVTY2rElm4fDW8oMqx34aHcY/
EF/FsVe0hZ/o8U+m7jqxznVsDfPIyQEga5Ca3oi20QCPijEbuj1fHdkir2Bf
wALUX7CWXldoqv9/aalTHA99fxIqCcjhHWeUcK2pulMhAdXCeUZGOHtfSEoC
qJCFBsm6XTrZtrTtv5tAbnEMTjxLCKTTFLErcUnU5tUB9u240jy5msgCwwaj
NiUbZg7RP9xKe2qmjB+6U9GJuEf6rY/5L9XOiYmKAfD3v7UoaWRmZs/oTrm3
A1M3AOVLPv+xh24eqHQaNyFKhOGt06Mdms8AgZS8wmooRyJ/bXKsOALqlEiN
qJeDu0BDUYEhKQcRbhw2Mdq+rUeAv5E6lJtkiUUxg76AW12SBAGbxwBj+LBo
T8G493EgZkucyOvLokWRg9fQlviRGxoI28du/QfeMDCPhL7mufVlQqEGUgxI
I+XGnChdbnlcCAQHI1R0KP6/ihDGaKZaNTk4jEEoMIndI+Hv5ssGPbNJlXeV
pfkvIpzcyWHDhKnsGxAzpCLXu7OuGTv9SRQZLdRi5lW3irIhmtwCgmNyAT3a
a972nsuP57Y6f1XIurq3LGMPW6ipEDQtfYw1ioxhJ+iwsV3oQy6D43AyqkVT
lgCelnW85bK0JwEiQIdr5It80qm21hie+pCYwV3CXGqrE/6ubi7/k1P6pmZA
uAlksvnUK4AJVu4VTlzi7sD6+/tOleRA4AriHi1ku/0RmNvzKAuJts6zaVjB
wO3n3QQojHsVE6Kg9xF2GICtBl+WDug30M9u7DnDg8tEVJLsDH5n+zPLY3va
8HPWejRxnrHiKcnPjI6lukq5dYU9iQDumsyQzmkFOV3Akz0aO7b0eyehukpo
VhhuoVlObGqe6RUOEcXLGHquCn2zprH5zCX1Zor1Rp49x3lmoyeKG1bov+l6
JlJVCR8AdNFcXuylqRULBBjWM3t7hMzECBRpOwEDfY8TBS38bOaiYttr9YCy
G96CRgxR5II3C+1dsoioJsdHp12oDvl7hQbwKfJk8ja/cNGkZDG56RLrp3xg
IYnFDPhd3eGu0PSx6P3tBQ9YDYuxIsNJclUrC+ccluVN/YRlilaID7ypPOq6
63A3+gMy9u/I0kCPifuBh/OjNTQmNm/7GyF4jonuDpo3pda+cMF/X0QA81v7
/oz5QTBIwYGcQ/u2Qui8r6A9SICuTKZ+O8vUZeNsI9Z69EzV1YGRJRHmEv+7
9p3ifbEhH5Z/LCl2QyjUfyZCK8zbbBBtW7os16JlMbZ6BRG2M4u7MJP6ZtuY
+wQrZq42howgpF9Xb9KvgNPzRf/EZ7WOvUb3OQ/fwLBJ2PuGvwcFg2XpQmsb
9HC3yVje4RByJFgEYk2no8qEZk6pkQxd+Q40/evfX05zA2YYusRAmZgEz7eY
UGFNFFXY/TE9yQkXp5p4HJ0qcgOK1+2MCuaE3q9XlKCZO6dLhklZCWF/OFGY
6s++SCygcyMuvBVOrRIwYlQrYDYuZ+zigjCCMHblGZNmc5b4z9kO0Q839J2K
kb9RdrbvX/EUeSLHF4Fr3phemjeDIpFuW9QWV9tmakReb5yFKNiTV9Z2T1I5
gvgWD84pDeyfm1uwjuJEd5oeHgovO2OeRoTmF4KYLmV8Swav5MSCpdsh9qq9
NGuwFtxwEo4k4Fx7cHI6YqZBJ08WGAMKb2UKRFAihK06fG4i6E0rnGB+4Bt1
TY1/GdCPCKHr9JnSfieJ03ou/DKcdZKO9OAfu2jCEQ4nCBP/Q5leGL+12LAp
dHTNuyynChU3e4JaWLrOiGvEdaA6p/19s2FS4KuOBfPeIxXTFAD+FM6WJGD1
kVrCtscxkN7tJLF13MRjuRjT7vumVPR8ECfqvHecLrORcllI2uBVWHZsiNbg
cIU5jlPJRbDzDY7A6zr9AxiJp+oRIeDiTEECLGaDzR1jVWyrAWM3jpaqeq69
IpsCxMkxAETtDagvlIMTLB4bvcxnn2HoneVv+snuovw1Rspg5iRNiwRRA/nF
cZZhUZE59olDbuf71PRp0PhjFT4hD6ZD9dMK7GxCTMZMAjp97NI+03rO8Kwn
QDLTZGEFKU/enq6EMezwEw2fQ0c/Ovf5FVwzGpzvzsnDwzbOjy0M4GDyXnZN
t2fLgrHalS+stTzv2RH3S4sfLdjRTEAHSCgGyNnGbyucLEiVGPlvY8zYncfT
tl9CvcSrRYT95tGYftG3A8AWySIfLFpWhuNSacVpljuaQHGAEHOOb9sUjCIi
kxOtDBWrNKKDYOXYL2A2e+kZi8XruVieS5+JpEIlzWBfqoFO35Li2fEQbCV9
Kc7MJd43GKkLvq9N/JEgsmopodwm7NfLzfQFZD+x86fBZRW61VU3SdHE82cA
n5PhNYPLT/Nj9TWJb1o6cSnTChyC80BU15ONBA5up5o94A34BFwPcbIF8OqU
7cPXzu8wf/1w+8oSgA5Ppwisy0U02aMX36VVPaVdlJXUe9cq9g6FTAJqjPGg
1gpMQdE90b3OxOdLZGFkz7BKpUTegeZPFb7IDh3y0IJvtyqf8oInDP2MDoe3
SF4XgQoKWvkaLk/mn4udzcI+6slKJzXx35grp9UIIb/QUFCxCqtUPgfnp9FE
Tv6rIYC5ckAbwebuuodBcUFM2BT5XgwrcQ3m1vNCKH5jvQvv+KkkGyEgDFPt
RntEWpTErI8NJFb4PmgzkqOrdEa+pLglKnRYORJNy7t4WVh/ClEB5oDPOLdl
ceWU/Y3sZbBF2x8wGaqnzfjmPJPAVqWsKPuKm5rV4RZ1VhGLtFIffakalSLU
iVSQa2IFtqkM+penuVdZlDtF8gefdiwuEipZ6mMcK8P6xDvsppfMbAfgHyH0
vnCyk2bWv7PShksOAIw5EPB6dRi4ckFNoZudEmkkvOFVFZGE3ocnfl/rpDFt
at8l9spvPXSlsmfB9mgU8wwvMhFyWUlqWh6m4c/G9c1G3Y3jJa/j5kmzVEma
BV/7zemRTjIORKg0vjixBLB7iXZQhSxIS7quvtLLGm5J+fs6qoN4o7gmG/1v
e+cMuECyJGt33XOPdUDlgpQOyUb9LHFdlNABaYVEyRyuMf2adzU0zze+LZUl
6PvtFQpzUa/PStg/sEPppSPXmWOSYmOCB9MM2XSlZFYH+d6ogyclnrekXXUy
RxMaSasq5lPKxWXDWZ0ii+xf6hcBDYQANvfxBsTh9mtM1PZ+O7SSXFXRCBsq
IK96uS/AT6En9GPEyjZzNZStL5cHVvobB2IiMBqFsFocFLl/6xfTaqRtasEQ
xoojFwC4+hcufmEfoyeCc8cGVdIsRDaONe00emaKsk0ASR+txqmN47x91Ka9
XcYIOaNq12DE4g/ESkDbN1lQEJP/DhKgg6s5JTGeoT7RGz2JjWD3oKHiV+/Z
u0GSzjSaVMtuHg0fnTnYDXT6zJt7HJby0fedHk7vJLH2Ecjc4EicTYp5LuCl
y9annZDSJ0POBUThKrjNug/fI5TixT0J7/wKHhGu62eK2Pw1NkofN97i9YuL
MBwcB0w+RmK/x22aHI6lMUmBSnIkVwPQfgccgwbAlq9iJWX4d/JXo65xfeFe
jE/nf5kksCE5EOTeAUhAWTPUe5vsjz5harg6CirDF/dK74rf6bT/ubaLjiVj
59RU1P3pT6G7RSGmuuKvoZlF49wwqsHBqDVP+3Je07WShjD07ozhvWepLu/L
XB/L4JHy2ghkZJxaKSsJdRmOwCx6/G1RnlE9HVgXQ8dPIcJuxAjSzyywERg+
1bTUUJ/v205VV9ZEnHfJp9Uj/2MfxjBPtLxasZpHqVXKrYv2blXufEa/suf2
fUEu0IJ/A4f9jH6KQGEPWwQXsGccMfK+XPgo19dzMX2Le1+dHlH6HGY5Kp+U
B1+ZENelUbJlXoIReHvm4TpYzJELW9NJvYH21nSd/obrdijGf73pb2aq7XXZ
a1EZn15Jvh9CGaTUvfasmKWBe/fkHGTXyTEn0edzUkIynfQN/Eft0A6wwDmk
dMLXfYY8Z2wTjR0ykSxUCwAQeHse32nPL3aYWiBcoeaIr5isrBoZKArVy/2N
Puw7+tzXWUCggiuV0T8AhgX9Pzt81ZWz/mSi1PsxZUX5vrxTjCiuDMYmbQ2i
69y0aqkXsJ8OenndQzrpOfn3Kg7dbTQfCEaqMIJ9y5mIPNiNxLJJ4k7kdbo6
RKzx+k4OvUHTVfwtknJ/oDV40Kz/X0pOgobeq7gvsC2kxH60DlHtTpIroUKI
3qHPdIeHbYdaqfafZmEauH3oeIt1SszQclBCPUKwLbnPuOcC8fl2T/DRSGjG
t50oqpHcE6j1+jdMJfsHsSgeHPHLn/Q6OmgJo/6gccQiZJXFWRqCWJSEVl6S
bCc9FrfOQIA6jYLqsbBzcKufxt8ixzPF381w33Ddco7gcxm3TuMmtAiGBSHZ
MBtt9eC30Inhf8gvlF1tegsFjugK51zsbC/wOeYE3HabYYW3hYaUxmF/gF/j
Ol/wN+RSXFEWvPWOvQ8wR5LCtSMCLTzRz40Yop3UDuG65Ecw/ViIMmNn4VBu
9bkqyueZFsaAy69kXy883y0qdK0UHodkqwjwF7f9GDERJHp1RcDo7X9lcLNP
89zmOIzYiJ/NehAcM0xVnXFpbixgg081Fxjvnqau7rqTgwoMwe7P1xmwyIT7
9IuJt47QErQGfLv+dfez6m2MAThyz08mN8MkFOkL8s76z7DoqVE+WKnErNFb
EaG/3mC+GCP4t//T+hgqiHorhnMWfTc4FzJKpHYVyYLh4mDJGbrmSh5Z2zfd
JxdYwesuBdSE2geKfrw1lzHA0snjq1+rAkxPmVa/gjS8AVrzSIMFB0JWqod7
OWoTJ+J04E8DGnPL7ebK1ZXyVyc8bpRVz+waaM4eJ3WKX44v4Zzs+/Ncu9/8
QB0nD2aT2GUnuAulMJLAZYMi+lLCRP2eWsHVNJKp6wc++ZpTeaf+rtEsNAXb
IwhHNo5bpSOUWMz4dITx5PoEkinIil92utocfzMOWTQERfrpT9E+PbC9qoEf
sbaYlTRSswTphe4MCR3xgQi4RVpAkJfuJcosNZL9fXNIxp3OEZ7OgjQpbTP/
JZ+17I12yHnybspPBFZ3Xan4UqUV416yolM4WBJFicySC+zvkWXXB2o3slAZ
JZq7kF2FNcbn4Q3usavlbacftnEoeoZEaVZYa2EA6RBzSiixYJyY85QSyLCY
VkYZ4Oz+paTrviuIfJgjCaWjA2yu1KHyaF1k1KYrgdrZ0EY1W/cZCZVEkUBQ
HCeEBH+IQ3Mg8OUidclPy8bnGzO55V06BtugI5nApHD8IFkqZtJtEbmHjniF
AIEQfLM2Y0ZVS4zuceE0tsNaaAj25xkzMy8ecUArLyqyCJkskbu1Ah3Exiga
jW00BcGWJH4cn6J2qm0aKFR4G43kfNxH6lhq7oSoxjdQpDQkKIVhbgCWKudZ
pUM31xp6ofxxxBAA3HFH5t0STlmSWukGUuZvd5UtFyAQ4h8laidSndWPcWnq
AuhGHdTMIFd7HWEhB9AhT/qQET9iwgU7bAgThWq/rvbxJgoKJnHgVIn0fUvA
9C5KKijlAqh5P32TaRNFRR4gVWlh94UxK/YfY38AwbBF2fO7dhUXxnA2wXyo
Kobzmqg8mWjpv+0kphrmoApU6F2xK5Bf7mQUv51RTOxMol0KjvuL2jGou07D
kKVGA5S1d/A1SF5Aab3QBK08/uVgPwB+bTUofl4T6lf8XZ2fdtV4feMI+Y0x
o9GqwW1qIvUYVOhinHFK8q/TvpQwGkjf2+KIf6AMTwV6Q+sB1u8Rcerq0YQG
IVkdqazvO0Lhk/R92OjKseU2YY7pyUXygekGzVUBwrydHGjmaGhAUBt0X3cJ
O9Aad9rXo4QTSV2TyxV8e/9j8gIBINBkK7+fm5ZykFHw6tsy+s1uswcCaLsm
rH8vgfyqr5sk2UDh/U/Fi5BwcuUWK0BXYBjar6It56q5mzcrl5AARVgydLXP
fYDe6nQhQfwdacafjaoyvIS3138rn3YWy8G1lpecjFi84+zLr9OmW5/jvkUR
sXv9ORgDw9IY6ZmmVDQgWrOx3gmWJKpc6KJXpUqq7psr80REOiZ5zPG9zdMp
3bhubwFPEUran23V4W6xe+TYc+SRwUTVd1xxeuR7dox+vh5qfr33hE0ic80V
ALHCCgu9DqONQZ+JsDYa5CUmA3eUC88M3MxcEswpunlnq2c7v3QcMYQZxQai
DB+IwFjSz6uN47vTjK88TzUtqRmbEKOOY7J2HRqU9YIk3eqt+S2MvNnRLQm/
R6KPqkCemMzjO2kuJdW09cqWcGdCO2C9LgiFSBC5hkGARJowvfqAcSR5oX7W
shYpWIkUoa/QsuVOyv/BhAZ35aP7NhYfCUjHFgzl366zzRar62pTlLos+MmB
moGQKkVC8GU25VEWWrDpVww6yRo90dDKsszXU68TxNUINB9K0N2Z8mtXbFwi
J4rb53i5yqTqcHm3NUslm0iRwsCbUImYkIGztnOAsj/Gh0IC2w9YgJcielxE
uvYMADtazLddOX7yYr2qNv1v3EJe1w6jCGDVE6edgu/7ITPXBQy9kw7U+kZf
LH3BKhFyO9wCFh2s8q5KSx+wvjqhgptfUJ0kRadvJks3OUPetORmWWVOqZU0
V1W9BN64mQtGCUCIiKZHoHRtezPA2iQkuHC06i5eI43xQ3WTJMb+rDosdWzs
j+Dyp2e7xS80i1Qo02gATq7W3av5em5jOu/gtaBDcy6jedtoe9geBLSNfbBg
iT6SDCnRiyBh80Z6ITr4h2g15V9ocbIMl1APyjGALTg0hkJpj5hb6flJH+V1
XFLyp9vg622OQM0kYcoK7HHwiVDRCAOauLGoxX4ZZz37mBcGIlhJRc3/C3Ve
yNuVp9HEOeDY4FbcUzIRLdWZCE1DnYO49XTBJubFd8XdA1zNGCmKLAgBK4uE
v1kkdKJa68lw26u5cwKi587/Su9LeOu3srWcqEG8xVOeq+MgTSCxvZaPEy2V
uBlGWIrnQislmoLJi+z4aJWOa4bUs6i2k59xVxGR4M9ek66uL8RSXpZjGjgY
SYxoct9hgMVPXNg35XUeQBcVSAvAsL3HneX014mUOCkcTt+lvaNmV1V0KYFP
YikDz2eAjcDNphcsNe0H+4JjP4SKpOEdyxe5ctHvfczAhU/9LRdK6EEN8mZY
gLgk9tz0bi9kICgK3ONuBy5ZC/GjcbgAqEhq2FMIk2EH+RadLLa9bDxhadgl
pEcudzlJ+HBTBFJeSkuzlKrnC80Sc3QgyKkDLRaEvlPU1ry4rwvroY4LvkxU
Hw4vHUXdPano88crtMR/EMwCD0LzMxuK3E7tBZhI0FsRsomlL6hDjPCRdoP0
p7WRB6NdGD/UqBsviKAtM/ylQbuhyihE1ro5v3ZmbSFybCAb+4SR9Lk+bd7A
Ja9o53+n/dkkNnkv2FYCct/YcojqNamGKehQAcwGS8NZDdvkHO5R+/Dkk4ZA
NEj0hA5RuB/mjVS9dxs41jv81qpXKcN25ZDET2/PwHVqGRIkHVup87pNTetd
F1Wxt/1WyoyV55dchZ57c1BNhCVlc7msMW4deRB85q26CZ7mE8q0iip8/k+Q
fTzO6obZSgrj5ef88vk/6vp3QQq5mw1vMJZADUucivmBtDof/zOYbeAFpqYT
Gu6RRhi/sI0Mz69I0DujFEUbWnzM4JyuZoLYk7QeL9IvtnTQSC7GoW9TGt0c
hcTtRI9ldV+GvyrnKIUo9Pb0lrURc3ZK419B8UyZxIhzrkYxnYe9FPl9xeGt
o4EVjEvNHdp4furdKznqqQXyuz0DlLDeTmzzzRWgL0e0+cHIvsBqsGShpJje
cN12WbvLltLzPh/8T7nkTxaDL0tIiWTWgVPN3i59dScZw6u//93tNMQ5CLia
izbkW+tq+hylyL82plhLrDgK57ggmf3I/Je3y+tK8GHR02+oBV6edByIr+Vz
Xxgx68Lwzfh6ERDu39cC1W8tq885xA/Z9IgBWqLLvLv2mwORIV3RER0TvEpl
t3ex+L9hIQXBKkdh6MS7QD5Fps7Vcjr+g+D9zTrBJsxxJvnGH/sOJVsQkjZv
I4fftiapOpFPnjHyqMw13156AURGU+WDYrS3rrYAilMLWQtvvtG78609bSm8
rRpBf1uX15vhHGDwdXAqS9kkfB7M/fZorC+V8wMe1GlIAMtmfy1YQDEWwT4y
WqXyxwnRUUaRWDKt9mc+lWRKwwb8Z//lVFNNduzl1dhNIhd4RJ+Ty0Z5tHtF
+PbLGhLTQQGp+qNbbOuA8vxXQA7+3j0dtn2npifjPOXuexe+2otGZQWd6WPr
UsQuZ0YQlGpGpPRTIQJVxBohMgmeMHw00INHTy8mrQ9w5ORPDT2sLCnvzUkV
Pc5ryCYhWl3xMNAUuzm3WAWH6JvQlUyI1UYpf9xC4OSfBYawFFuNPPZF4hT2
UmA12YvRlUMMqTGcdSagTBEyH2qvKtQrhOZPVMRVBM8uZksQY5zvRP1Z+af0
Q69i1b8DNcCeaE9PjwzPdhy/GZg7WELGk6rzplRfBkmICzPEQH46SC9T1m9e
DJ7DqN/lhVJM3T2tkRhMPOjAm27x/of5FXJflGjdJVImxpY0WBd/MeP6G2ca
HjxPcF8SorBwA7Vi8uXO7dTRRxree0QozC2rEB+tOLbGTd6Q41oBIgcOemcJ
H0QtibTVjyZcAhcUAho7YQatLOjod6QoPKnx1SSxiEmcfe2f5KtW5TvyWCY+
fvSgeT9NeC5zLk2EEQWBp8QnrJHH4whDzWp6iuHcaL1wsumos4stpiWamm5k
WhUC5aUhIZux5t+5YAjdpjkBy7eVNuc6DGRXZ6o5wCuCVP5brmQOLnPiu5ex
Aueuw6nKIhnrD++k1YoFSWcyldhCVNkShvN6ZsyB4vdmwvpPnatBmoKF9zX8
B1c02t4EhEfygyV2D2X3WByww61H154zc7oek4Ald2stNyMoD0Ae6OXumxvR
huXV0P+kWE+TFU7EpESEe+CStE7eCwPIuD0Gv7l7uvkSLqycTc90557+Glyh
LqKFiENxGXELkfD1eV1rScW2gFCpQNOB4XSlVvJlPHHDLvGNq1Ax71q3Aqjs
NzA1NK7FPH6ZC8jFz1ZiVhGBBEYbH98eHxLoNXLPMXNs9dVjTgBLyIDpfGcx
kf8wuzO28IAirzGCyprYZ+DpDL3Tc3Uhbq9rFZNIfKIG7FnTI2QnTJF5P+sJ
yZ0jguAz5V+/Ldm1pawY/mU+BAI5bKq5cADGc3d9wT74Lbw8XyDDG6n0saMY
KkKI2TfWn+UA38G/elbLlTxwllVw0VdTR876T0/I/AR73bD1IZgYO3GD25vu
pJPCvqnOT+tEN8h7vqZcwnbFEP4TZJh/72QILBxD9neFqe7qX+MxsspiterL
Bcg4XCVLW7YaKSBtlXvadfmGxHDJo3ahfO3i73r6sH+p2jDRzEA1I48v5kCO
Y2c5RVDK157Ql4/Vrel8y+WW3gV67Z6nEuKmEMkameqj5KzvQDm3J+BITL2S
8NpXHyAKM8nhLfPyJvmAHljlSpJ/Fr83E4XhK6Sh0tlRRQHEeu+QFlhWpLW/
vIRYCNIrqYoRvl4tK5kR8xPXuO3vSyaYTNyX1eaZv+fRAh7YAmCm+7g4GFde
/oECADcQgKk32QqHEPJD4tjHJiO3kIZ0j8R9EinGOywEYk6ROiyl/XY3tMyE
YKkTbUUL7rNduSLqzt2T1Q/w4bLpQgMhDBgPFEO3XMR3C0CFXpzMklaHor75
IbaKZwlvYkvkPNbWVH8OQA9X4il6K0/EeV3xkqmreBNYAKv3blYjq0LAgoo5
RTAhTDmedaeYphLZ0AH7rjv1NH/VPPWtipg73swzzyYGDBqMV/Td30RhodJ9
zhyuHxYQXVpBG2aYPvoZI3oMGWmF8wOj6CcSuhxeKiot2TBRu8j44VmN9Vpf
tUg/C5YtM51Agu1j3qQInx04tQkLllapq8SYQlWgbU1b1bofmd8cLyZUlbvJ
Gdn4z9qr06FxP8wBJOBeP3mZvM1LcL76k6HXytG04V2NUQ7s6jQAm2NMzKfG
+XjsHk1+9pL3QJpGnvM4a/QqHwaCApBKeBRWfgDEe+kwplst1aq3UrMgWOK0
NqqbpBZfkbuUHxtUlSWK9GQ8V9dETFg/Vy1mdiKzSTt9gFeefnu2b0WR6B6Y
YJKC61kwuxbJ4Ml9b3PZ4ck9dYIjbzt7fJ7LVM0BHbYnf/k2c43qJA/k2jOL
kKvktQk9u5Z7Q5ej+ak+uPh6uVj/lflfnAQSxtUySO25PUItOSHOV5ikJNZH
6Gr2C37XW2qdgR2NwZutTkL/NnGu+vA39zdaaFK5RCKQ7IoCYnorg43Oz/+h
cuAmVjRnkebsvo06SFH/4u0DIvFUqPqqGVI3w+R46bDxtcbzdUpzvB8II+pI
y82tn6o+H2b4Gm9sB7mnwqlA8tUC8GJsag6Pc5GUhizRNsdAqAa9iLpNjgOY
BlPsCkufCuJhPrIRvxhgpOOunud5AJdqPWg0SywWzKs0Dvm9029KW+ifv51U
QKEh1Xko+SdTpRmFDUTi9PDGrf72Rf+ozGK6r2iqRQrbgLeG9dDcwvDLsD9y
586rrG/8Qcot0i2YDLR1l9/b0wsn2UEBDIJiHxwnFTJJNdzeLUwKH1eDttQo
UPszIPnITeW2Ye5VGL2efrglwKBk7r0/Afbd8iyB+H4I7AHDyykrB4oCuTSt
viif17MBbx9R3E271o+kmFVtFgRKCDfV5Qt+M+wJkO9bw3hSxzd/KdQz8uh1
M2a9/s6fKRJBCMB3WOTIP2M9ovu0yPt9LevjR7NCBRBD1dtfsHNGnj4Ecaqw
rf5q+BRGl+6qKQNIKDzgcQo1YL3oCDTPz3azMvg8Lm5UBfbqkwpd1fJ5iqBM
wKApZr+8dBipTTcTOq8ZMnX/qxKBfZ2sbUlYGR6P0Bf5Dnf2v3Qn1aP8WPrx
DwD9wcOMmP85kEdwTkgUwMNsqJh3idxTCnm9xZTmdloY14p4jE8yElyAtkw2
L1auUbBaWy5jYHfyh/0Uy4+MFvpjBN/biliSfo0HJPWlmA5ljn6k76vcqm7k
zFNuoMBUMbFKsN5SdjgfD5bG8n8K/Obw36MMKXm1XYHckAJ8wn7fzqqjpp1n
TGqwuOQF8czPM86dQ3fRokkVMfPKvUC6Sfsg4tCgD+SLVboCjTWsb43QQBXU
eF2Y+bQB9p1wNfemeG+906FjXopyAGN08dqRKTs8UmSzqangxkJWSPbQA9oR
mbzO6M7rxgDOuvpIHpNfOPs1UHp4eBC6KqIJsM+SShLcP15YIu5B6ErcvkiU
iC9R5C229pPvWocNFU0mLs5Bu4S92O2sKrSSk7UKWdOpOWuthcKt/ECgmNVG
ztSTqRZp/UDzM/UhWFGS4ueqsIv1tzXsPDZzHc+7tggo4oCfXaDKpufKW0yN
qwclMrj31lWBPes2u9s3u2wP/ay7gPTK/MdYXnJQMCi6DWf3Ww0viiywQ4Zt
u7pAegUiCgZ3Qv1dK4D14SMu11PMEPd3XY8F92rXvzvHcu/A3UGkALtx2iUK
ot4I2EHn5n5yqmU3JaDsdS8IZvtWQj6318JCu9pW0nnfwupy8p5rX7ekwTPT
esXBWuypVipKXa6QMDI/v/eqvZFNvUnUz+Uh835vJRO7I2fhunL/cIdhtQtK
52RJIjdhiweA6AF5TcFec0C7TKul0Pg9q4N3s4aWLC/IQZQxVamNmnqToKjw
aW1zX4QLZ3CvG0+gYx6i+3nFxqB0pxpMcfiL7LawEwLLGPMZKOnU6W1q+M5q
DvVrSTW2S+kcOCi7zsKSoLFFXejBYY++Ll2blWyomoxNFct80b3RIIANDXAl
0uPdf6Oo2v6jZfN3oAi8aUktVDuCmwpQ3WruYb3w5CTrRCXTwVo/JHey5IX3
GGRgIgZIfmtELWbmt/pcPxWtuimZbsvvHK9HwL02w9gxEJhHiCLVuFv+UUg5
tFMbuWkINGMz15pFRCoRtI0zG7BI+4zG6Wih8a/98bL6HkiuDyAymeWXdkhS
YHHHRW2SfLktju0nflclg0dCP7QUIaSpIshkqypvsBCPwG2RGEPXD1KO9FFH
YLOpGirrrkjIcQyjTT7Wxle5ezTievTPN4D734YvPttU64UUnGXAJqvxwBxY
fw03teAxfoj1oc/oKvTe302A/7HDOzWGJZ3boDMW5GJkIUr5yltSpLsDkeNx
jvIoq2hMkJQnwytB8ml2u6r1KnwVzD2S+iTYPjyENeZhH+G9pJBSJcmKF77B
cUli8R0/oz3m1Pg9qx22aO++qtT/pAk/17wvGNeIACNYTQx/HqOo3szhAK3h
EwwEkqHD5GacjM0ZPdald1bv+iGrXmR4pEbrAV+TEl+y6Q17cK4WyeN4Nx9S
lzP5mUaWM7Z0Em5fEgUpU3SQaCFa01CItHK6HJ21yfwsmMMaHuMidPvFa1mW
sH3uSIcKgf1MkS+kCbAeJMFjATJof4IPAqQDTF352b5zDJo+VGWRCgXDwQGr
pZCDHBycmbSvHc54NYLHXK/DC6RRP3ZGczDLGm2ze+Nya+5X+epM7lsxHHPg
kmPW+91aaNmTP9psSb2vjfN5j4nh04rhe0cHfxtftytYzvd3lrYmCXbnbS8Z
7OkmLgccDYudUjfE0ApGE9EFEiOsTdvkjl4bClhdB9mgblMnBDsHG1sAtYwR
+zo41oQqHaG1ycpftlkoCzcYhOzgfbRtHmpIgNx0T3/iO76nnf/M8RnChGvi
3tCS0pOxC6iwK7DH30VA0OsK8lQeVC04Fcfz1LqRGgmuIucsOreI8RlUxSkD
dkFJICsq4RoKwsHIWz6ygMjmOl57fl1ihD872CszUkwfssVJRWfgSH/7x7ON
w2NZSq+E/IL3zqeCM6EXjFZ90XaqUtCo/hN4FYsvn0vInkWJzOSjHkx/Ypre
iseifCoJivj/gpB4J8DagJRISdH/czEiziaqcazFozihEp3VMjz5WD16+EXq
knPUaYvNfLtFJbfOMamRPfw8IDkCMor0Wuk1dt3xK0HofEVR9EKYvbVLB0wP
aDOqKgTb9GELyLfLHILfIPqlylIe7bYukUKujZZVbqWGs1QqNonEZVjtHuyd
7IVXjVJgQV3Mu4xcARgwkXmKHN81YHO0eNN8xD3eFVsHjpBMT4UFOorFdG66
xIsg/FagQhqtfmo+REpUH1exSP3gP1f9OL0sYYbjVs2D0f1ma8RzAqLQAXJL
bRVhq8Ym0ZIs+2wYZNG9MdxNqqq48KKbLaHGcjjOEMAdN/FFEmauU4ncBLsy
fvqmZ/rw9Rz6ALEccoVKqMZCu+wf63AsHKuaZ3x5WE7ATUSrBW/ksCWHSWvL
u/ahQigAU/joPksI5r6TyY39JWBfQe8kHS1c3Puycua4C9DJAc86pXWltXEZ
yi9yOct7AMu0kc3epbbF8Gc1ox5URMXTfgZKCsAGXcYVHfz2VCDdt/x/ITtb
9UGwuiGpYgfp9clZARZtL1rrSVFCZv1iLqnoqcSCosTP+AsayYl/VZJB1NIj
ITS+mN4+bcmpgw27yPS+k10v8Ly3vICaZQCZi+tk7lYTBz1edDe0NrrBvBSb
/sCqkU7XThEgflZMKTmbYabDuEP2WS9OTtVoVuXjqLRkWxkyt7gwx5L2ML6p
jQk2qPmG2yase6XI0ageuFZYZAD5m7swhtWyh9+9J42vRUt+BcBbgTtcOh3p
wGjpeZqtpRAfJLNx1Spvz2wP7SiRnPjQy3fSVAbgK21IDhi2z0jYvv0B7/hn
XOdQtHjjlB+QscV2N4GqARieukO7+yCiWlVub3YCF3mlC2DYf4w/RvAtS4ps
Js6pPththZ/Mlj+ut4aZh1VlT6LSAgzH299oMfFBiRRpZnBHCMkeeSmRaTo0
W7gzuvv9iYpM+GYXM0EVcYDVGSw92ZWc6v38EOkd5h+0zWupy4kiAHmKh3pw
Oql7siOLoT7eZoT5OZG1NV1aUMVrHMqjsbVh/cxbB5IrA3e6Irw/MDxnzrbv
2XNQDIoC9rDDORC29fW1IZAYGxr0MsNcSfvV+1myZF+emoxsiTBzEawxdRx2
5RbnvvPExkNaGRpNBdUw2YG26L31DADhclIiGdD9bzP6QY+t2m9JnbHfddxp
InCPEHZnWRvdwghS9Jg8exIuF7DVUOpz4bSnwEDOkn1XYbApgFEUIxvE9Hky
TP1j9r5xY+gqRDw10i3KNvCPP+HK+onCSC8F3QJlQ7WYbfk48s3mH9HKsNRv
CW9Vt27xzRx5Y8bg4dZBiQ1LkKE9aY6HtqfyrXLaFXLcCmXYy+SMx93X2/Dr
jEEYfH7pLVOi+eoo8WcJsT5KPwvHwMVZuHVt64X7mCXQlX+pdHTpl9lVfJeo
kL2J3aQUdQjMdtPNozx9lhh/0oMKV20S9RDtVJkjPjLANCe/yVBZ/AtsZ6jx
j8laI/c+lxNd6ltnTqrpl2wv+4uvjnuT22BK7rl1Ffp4m/1Qec1c/jWi7oR+
AAG4aEO27feKv82JyKOGssrp5BhikbWirHuoRzyowb6Q8jh1ukWR5L0zb+k3
M/ongedqX3JrNBAcpIDzleSP7BoIaxT2vUEvsNKNNH+p80Obrb7O/JYCTcRi
7S86KZ6rbmeJ8OclnpaC/FqqYJAmc5G4W8QoyZDYiMRT5XDZum2Fq/TChGUz
KbDtKf5UxygrSdjcqW8D2QQDtEyy5sY8dT/bzfXEEPiwhVyupMo5jZ/7y5IK
vzbMICzQ/x9gjZsuLJsvcq/9165NmrUqATvAGqZgXHwr1X1am2Hd9UlHoB8u
FOc3i7Wqn9BT+v+sQ2LXB7l5DWiHqZmO2iUNo6ddN9xk5bnar+1wUdYZXTDl
AQ742PcwVyLWkOQgTGPgKS+aCt5Yf1dZkWEmSg/h36U5ropGJ4MDSp8HLJAX
2DBHnoe+tHGjxbVrGt+BHFNu16ril7DJvlHXWpC97A6L50eb/7bpvapdK8HZ
r0VSrI2jR3Y26FpmXGvLtig1YEpw0X5ftzYpwjEG6HGv0o8Z2T2sX30jcE5I
UEKk73WqotQP1+Lchdgz4XvYhX3MQ5CJLIUrfUze+X83RAIvmeenHsDLolr0
YtQuOMkWbWOhnkrpN627rWkxdZZaUzLb2elvfCaI0twO4Y0pEv2YyWz1NdYd
ExBbops4L1CGQWCQJ6KXJiMLZFDTTjt+TRWvg5AvyLVE11oCKJpf7Tb5PVK/
6yVVW8pzpaYhlYFaVeZ55Sgce1RN1bJ0fYbjiTPF4zBcrLPuWVYU3aKJRizO
yoz30DzXxplgkm++NEu8C2dVB3hPqAB4KYX1iH/8BSWzZ/05xCgWfsOPIPX6
viOU5rOozT5ZXBeyVvp2HexgVJdOkVQ+In79eN2Qp0KuIwuOAvh0nwkL4QPS
1ob0/a2YURaaZLiGjTcdP+MDIAXUC4jJjgEp1/uvM9nmG4b+ymPwhuZFts3o
K8FlIc9cbqw596+UQ6KZqlyv1cdBKTGkGYwezngNyNYdWZL/+UHkXL578cBQ
AbFebg4fDEDl1tXTm/Q11RwwNnWH3gOULfOpq90Cj85fGdEV0BB66Nezo38j
yh/AsWmI9/SH9ommoWF4EAq9jjxET7RRc4uC6ENgqHjlX2FnxIqPZr5EwTV7
mhSRFae5neW6WVH3N9nQh8/hymJLROPTnlOLUwPYJWC5KRu+i9Cjt8okEs51
wiX3blRqa/6vtG9mzJN4bIAAMFV+z5kb3Ob0S/eAyvIp8ceh8KZsblACz6P4
sfdnOwIgGIYMNpHMdwLxLyzMeF/8Sd2HAwF7SIPOeax2aPqJNW3PMVGO15TT
Nwqusmrijz96XJ9fX0T1OBaQ5ejnLyWDl18nr2gWVpJHlbVk8WjDLPUnkg+w
BuFCrG7lrmujdVMK+SJd1MfvDFL7YI32xrk+KUWl7FDC/7FSW3OOKXCPbrU3
SJ1xrPH9xY8fnpcfQf/tCg6rb9Gfjsem2/xNA8vmeVK3++uOunFXSWTUXeYx
kLldppcdvFBsyuAiXZV1sC0dVhnG0SApGgPNkqeseMwYZRysrUxzykQPixvO
5TWbw4XeeRHmbHGQjDD9av412B+t0EKL46MEZYDHOt9n0b0f4XFg22J69p5i
k/NtlUPiSLEf/668gT4ihsM9i2487zpnMkIfhZ1ra9arG3Qq7JhN8VqJU6nF
F9Ty3Hr+o2RdR/aYSy3lDMh+nB0g2JmeFvbQ8L9erwzNyAoJXkJpMiMf2ho2
G2l+tIP1/8SIvzOLg+UrIR6FM/ThRGAA6Jjp7AurqR2JN0itTWQF93HQlLPu
JcDRJoWg5W1CNkZ7ABBCEMAxz7WzDjEulZHJoGc0VoJ969Cqowb2hL/64TdQ
HobzoJlhFYslsMgBd9CgENLNBdw6eIw8HYsyxP9QS11Y0LLtdSGy+aEbi/l7
ss4EqtgkIi1a9GhHVS3a9eEI6QeIiTO1EROELWhjgvFEIKKb1KSFMENmAQaG
1wXvfLZteD32j57IfQCxknKOv1ORSmb3J3txG1InpHFH1eC/kbINhdw18dAy
DQSqDkQ6J8bbYbq/sVYL9NS3a5hdMhtjOix+6D3fGMlZPJWP7uh7TPoGKVRr
PVa58BisP43C67Dp5/84qsSOUdI2XzXI3aEatRe/GkfUQSPa3481AlhrhRQf
9YQsroohIZEQCYMZZxHllxFgPWPHTXBpPNJbwXbXykMf//Ew1GA4RQeJ8AWB
cqNNIukQ52Fjc6X8YgORuKsJugbEObuwisj4S8WU3e5Gm0dbqrrbkeQ1C5GO
RvtpltEQ+OOnGIUdtiI04eqnN9JDPfmOOrp7EB+CtkZZdTQ5zKtVuiloAuM9
qWPplkum2FcbhZkKgQVKVQh0w/gP97LSjTyekqeqBQmwiJ2vhnc1OTKf2ioL
w31Bu9ZLr7XCNTIWyvRV8wDH4OgwJlWTwrE0yBGNRbQRyWNhEom1rE8egaL/
KQLcZikkL0OT+MNzLWQnXqhWc1VS7EXNZXX19uIKmyYjx7+K/Hulg5F+O7/O
XWlDxM4IfnBfP1/3SmiyiNHTsKKcXSIcEKNaCUf7t6hFCAKbDOAH9TD7prqv
AFwysAwbFx3YxwKV9Qs55thL2tHPfNgvJienN6yYmwwkm6ffWgHws0VTZF0+
vn2HJgK8lXP8RKLnO7IHlSr7/PIKaH/PLy0b818phTbAdrKSy0cMY3HPgChW
OgOULpL/wOmsPfqgN3I+5rYAYa/X8vUbWmWyRU77XwXB9lWaDLEdHgYCNEmZ
lAImZ8JxePOnezyjPCzIxPBsEyppqghLe5sqD0UvLGATqUmPnjBjUvv+JjF2
Ux6k5ORvo/DukjD0wCpl7eta3JWDAlUEUM1w4b9SNukxck6IbLt/qX6Ke8Be
aVzaq3a/GQSX1Fqw3OR3wOUSkemgqrZsY0DT14eLovVtS5YUV2fa6ggVIiAs
gZNhqDEVJ+QY4iigHmeJi1aPTLdChys3vgVIrc9VgvlnxZLxS9D0x7HQKYck
0r8QfqXGN4bQkrTtNBH2e5joRTI06qQOBy5HSumT07rbh4yz/WcMBNIkjkta
80cHP/Yt/veS2VbOlUfi0p0vm+pBnpo+WFS7gONfAkOBtwnvQHaWENEmtKiW
g6PAAAmnlVcbEG+/O4Iehg3RCi9N+zcd4yxykL0Brzof0d+Si7zcx2EiLmHp
SD/Esz3kMzyTJK92KGjkNVBYRZY/nU94xsnBlV7ZdXdS2IGILi0WVgiYhIZf
hjor7wefY1mzD8MK2vOQEfI8OLu8smpRBExwCad0n4CUYILZ3jOGNZaqlWvb
AT1hXt4EGyc6p0A9Yq8=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+ErI6wiY2cNJZpfyJsxadriRu38oxH5cbeEksZ6Xc4lpaAn5sPGb5ndV1mOMsFI5dKOon6NTYsqD4rhxgsgOGZE5rKZ3qMzHvvkkWP8pKLWa/vfjKso8EGUx0Bh9rhTHZuKaxi3/XpZGquye8dBRaCetg4vNmrX7YcgAfJ+sDZ8NlSDVwKV865G04KAaevJMz8h4Q60cT4qXI6z0pPvy8PtyNknW7ks6gQZKn6GoLqo0SFMi48SRTBhwSmuCWKxEKi88Qy+g3yKn3bCvZgisGoGbAhTXWTNrW5GW81Y0T7mqO3d3kXa/nl9Sr+SOGHreSevugB/cMRgh6SHor9oRWekJT6vOhoRX1q8SAjKhBA3iOQtyyFjEQtCGzTlzbyzYWft/t6liGBO5pL15RAeLhSeZkXTX9EfDcCdfphi1lXCT2BMPhjg0Rys97/43fqgu5OBtYKs8kBhrUe8MomfDAv4SG/5lXhuPV8pmSmZtFbPxCdnAwmzp0WPiFaqy9+4CAgWAUlIBZ3a/vRqrwwElVvACuVL57G+FCp2ZDwDIr+FgKELY8in0Fo4CX6UuighdeFp39hp5PYTJw04Je27fHhnc9y9MlUccqSGjvy99WEX8+PDdsAHHU4Nrhvaz/KHMQ4sm55rJbOFTTz5fEZxelxS+4vqDYi0g3DrA/PaEqRN/kdNmyUKObLUL8gC0IF78OZ4lEgQ8HVgf+N7UeiCdJG+PWAXeoE3ag2l2yjM9GUxr29RDUNRTDE3+GIz3Xwh9QhJPmMbomWuET7cF4qffOW1S"
`endif